// Benchmark "wb_conmax" written by ABC on Thu Oct  8 22:04:30 2020

module wb_conmax ( clock, 
    clk_i, rst_i, m0_we_i, m0_cyc_i, m0_stb_i, m1_we_i, m1_cyc_i, m1_stb_i,
    m2_we_i, m2_cyc_i, m2_stb_i, m3_we_i, m3_cyc_i, m3_stb_i, m4_we_i,
    m4_cyc_i, m4_stb_i, m5_we_i, m5_cyc_i, m5_stb_i, m6_we_i, m6_cyc_i,
    m6_stb_i, m7_we_i, m7_cyc_i, m7_stb_i, s0_ack_i, s0_err_i, s0_rty_i,
    s1_ack_i, s1_err_i, s1_rty_i, s2_ack_i, s2_err_i, s2_rty_i, s3_ack_i,
    s3_err_i, s3_rty_i, s4_ack_i, s4_err_i, s4_rty_i, s5_ack_i, s5_err_i,
    s5_rty_i, s6_ack_i, s6_err_i, s6_rty_i, s7_ack_i, s7_err_i, s7_rty_i,
    s8_ack_i, s8_err_i, s8_rty_i, s9_ack_i, s9_err_i, s9_rty_i, s10_ack_i,
    s10_err_i, s10_rty_i, s11_ack_i, s11_err_i, s11_rty_i, s12_ack_i,
    s12_err_i, s12_rty_i, s13_ack_i, s13_err_i, s13_rty_i, s14_ack_i,
    s14_err_i, s14_rty_i, s15_ack_i, s15_err_i, s15_rty_i, \m0_data_i[0] ,
    \m0_data_i[1] , \m0_data_i[2] , \m0_data_i[3] , \m0_data_i[4] ,
    \m0_data_i[5] , \m0_data_i[6] , \m0_data_i[7] , \m0_data_i[8] ,
    \m0_data_i[9] , \m0_data_i[10] , \m0_data_i[11] , \m0_data_i[12] ,
    \m0_data_i[13] , \m0_data_i[14] , \m0_data_i[15] , \m0_data_i[16] ,
    \m0_data_i[17] , \m0_data_i[18] , \m0_data_i[19] , \m0_data_i[20] ,
    \m0_data_i[21] , \m0_data_i[22] , \m0_data_i[23] , \m0_data_i[24] ,
    \m0_data_i[25] , \m0_data_i[26] , \m0_data_i[27] , \m0_data_i[28] ,
    \m0_data_i[29] , \m0_data_i[30] , \m0_data_i[31] , \m0_addr_i[0] ,
    \m0_addr_i[1] , \m0_addr_i[2] , \m0_addr_i[3] , \m0_addr_i[4] ,
    \m0_addr_i[5] , \m0_addr_i[6] , \m0_addr_i[7] , \m0_addr_i[8] ,
    \m0_addr_i[9] , \m0_addr_i[10] , \m0_addr_i[11] , \m0_addr_i[12] ,
    \m0_addr_i[13] , \m0_addr_i[14] , \m0_addr_i[15] , \m0_addr_i[16] ,
    \m0_addr_i[17] , \m0_addr_i[18] , \m0_addr_i[19] , \m0_addr_i[20] ,
    \m0_addr_i[21] , \m0_addr_i[22] , \m0_addr_i[23] , \m0_addr_i[24] ,
    \m0_addr_i[25] , \m0_addr_i[26] , \m0_addr_i[27] , \m0_addr_i[28] ,
    \m0_addr_i[29] , \m0_addr_i[30] , \m0_addr_i[31] , \m1_data_i[0] ,
    \m1_data_i[1] , \m1_data_i[2] , \m1_data_i[3] , \m1_data_i[4] ,
    \m1_data_i[5] , \m1_data_i[6] , \m1_data_i[7] , \m1_data_i[8] ,
    \m1_data_i[9] , \m1_data_i[10] , \m1_data_i[11] , \m1_data_i[12] ,
    \m1_data_i[13] , \m1_data_i[14] , \m1_data_i[15] , \m1_data_i[16] ,
    \m1_data_i[17] , \m1_data_i[18] , \m1_data_i[19] , \m1_data_i[20] ,
    \m1_data_i[21] , \m1_data_i[22] , \m1_data_i[23] , \m1_data_i[24] ,
    \m1_data_i[25] , \m1_data_i[26] , \m1_data_i[27] , \m1_data_i[28] ,
    \m1_data_i[29] , \m1_data_i[30] , \m1_data_i[31] , \m1_addr_i[0] ,
    \m1_addr_i[1] , \m1_addr_i[2] , \m1_addr_i[3] , \m1_addr_i[4] ,
    \m1_addr_i[5] , \m1_addr_i[6] , \m1_addr_i[7] , \m1_addr_i[8] ,
    \m1_addr_i[9] , \m1_addr_i[10] , \m1_addr_i[11] , \m1_addr_i[12] ,
    \m1_addr_i[13] , \m1_addr_i[14] , \m1_addr_i[15] , \m1_addr_i[16] ,
    \m1_addr_i[17] , \m1_addr_i[18] , \m1_addr_i[19] , \m1_addr_i[20] ,
    \m1_addr_i[21] , \m1_addr_i[22] , \m1_addr_i[23] , \m1_addr_i[24] ,
    \m1_addr_i[25] , \m1_addr_i[26] , \m1_addr_i[27] , \m1_addr_i[28] ,
    \m1_addr_i[29] , \m1_addr_i[30] , \m1_addr_i[31] , \m2_data_i[0] ,
    \m2_data_i[1] , \m2_data_i[2] , \m2_data_i[3] , \m2_data_i[4] ,
    \m2_data_i[5] , \m2_data_i[6] , \m2_data_i[7] , \m2_data_i[8] ,
    \m2_data_i[9] , \m2_data_i[10] , \m2_data_i[11] , \m2_data_i[12] ,
    \m2_data_i[13] , \m2_data_i[14] , \m2_data_i[15] , \m2_data_i[16] ,
    \m2_data_i[17] , \m2_data_i[18] , \m2_data_i[19] , \m2_data_i[20] ,
    \m2_data_i[21] , \m2_data_i[22] , \m2_data_i[23] , \m2_data_i[24] ,
    \m2_data_i[25] , \m2_data_i[26] , \m2_data_i[27] , \m2_data_i[28] ,
    \m2_data_i[29] , \m2_data_i[30] , \m2_data_i[31] , \m2_addr_i[0] ,
    \m2_addr_i[1] , \m2_addr_i[2] , \m2_addr_i[3] , \m2_addr_i[4] ,
    \m2_addr_i[5] , \m2_addr_i[6] , \m2_addr_i[7] , \m2_addr_i[8] ,
    \m2_addr_i[9] , \m2_addr_i[10] , \m2_addr_i[11] , \m2_addr_i[12] ,
    \m2_addr_i[13] , \m2_addr_i[14] , \m2_addr_i[15] , \m2_addr_i[16] ,
    \m2_addr_i[17] , \m2_addr_i[18] , \m2_addr_i[19] , \m2_addr_i[20] ,
    \m2_addr_i[21] , \m2_addr_i[22] , \m2_addr_i[23] , \m2_addr_i[24] ,
    \m2_addr_i[25] , \m2_addr_i[26] , \m2_addr_i[27] , \m2_addr_i[28] ,
    \m2_addr_i[29] , \m2_addr_i[30] , \m2_addr_i[31] , \m3_data_i[0] ,
    \m3_data_i[1] , \m3_data_i[2] , \m3_data_i[3] , \m3_data_i[4] ,
    \m3_data_i[5] , \m3_data_i[6] , \m3_data_i[7] , \m3_data_i[8] ,
    \m3_data_i[9] , \m3_data_i[10] , \m3_data_i[11] , \m3_data_i[12] ,
    \m3_data_i[13] , \m3_data_i[14] , \m3_data_i[15] , \m3_data_i[16] ,
    \m3_data_i[17] , \m3_data_i[18] , \m3_data_i[19] , \m3_data_i[20] ,
    \m3_data_i[21] , \m3_data_i[22] , \m3_data_i[23] , \m3_data_i[24] ,
    \m3_data_i[25] , \m3_data_i[26] , \m3_data_i[27] , \m3_data_i[28] ,
    \m3_data_i[29] , \m3_data_i[30] , \m3_data_i[31] , \m3_addr_i[0] ,
    \m3_addr_i[1] , \m3_addr_i[2] , \m3_addr_i[3] , \m3_addr_i[4] ,
    \m3_addr_i[5] , \m3_addr_i[6] , \m3_addr_i[7] , \m3_addr_i[8] ,
    \m3_addr_i[9] , \m3_addr_i[10] , \m3_addr_i[11] , \m3_addr_i[12] ,
    \m3_addr_i[13] , \m3_addr_i[14] , \m3_addr_i[15] , \m3_addr_i[16] ,
    \m3_addr_i[17] , \m3_addr_i[18] , \m3_addr_i[19] , \m3_addr_i[20] ,
    \m3_addr_i[21] , \m3_addr_i[22] , \m3_addr_i[23] , \m3_addr_i[24] ,
    \m3_addr_i[25] , \m3_addr_i[26] , \m3_addr_i[27] , \m3_addr_i[28] ,
    \m3_addr_i[29] , \m3_addr_i[30] , \m3_addr_i[31] , \m4_data_i[0] ,
    \m4_data_i[1] , \m4_data_i[2] , \m4_data_i[3] , \m4_data_i[4] ,
    \m4_data_i[5] , \m4_data_i[6] , \m4_data_i[7] , \m4_data_i[8] ,
    \m4_data_i[9] , \m4_data_i[10] , \m4_data_i[11] , \m4_data_i[12] ,
    \m4_data_i[13] , \m4_data_i[14] , \m4_data_i[15] , \m4_data_i[16] ,
    \m4_data_i[17] , \m4_data_i[18] , \m4_data_i[19] , \m4_data_i[20] ,
    \m4_data_i[21] , \m4_data_i[22] , \m4_data_i[23] , \m4_data_i[24] ,
    \m4_data_i[25] , \m4_data_i[26] , \m4_data_i[27] , \m4_data_i[28] ,
    \m4_data_i[29] , \m4_data_i[30] , \m4_data_i[31] , \m4_addr_i[0] ,
    \m4_addr_i[1] , \m4_addr_i[2] , \m4_addr_i[3] , \m4_addr_i[4] ,
    \m4_addr_i[5] , \m4_addr_i[6] , \m4_addr_i[7] , \m4_addr_i[8] ,
    \m4_addr_i[9] , \m4_addr_i[10] , \m4_addr_i[11] , \m4_addr_i[12] ,
    \m4_addr_i[13] , \m4_addr_i[14] , \m4_addr_i[15] , \m4_addr_i[16] ,
    \m4_addr_i[17] , \m4_addr_i[18] , \m4_addr_i[19] , \m4_addr_i[20] ,
    \m4_addr_i[21] , \m4_addr_i[22] , \m4_addr_i[23] , \m4_addr_i[24] ,
    \m4_addr_i[25] , \m4_addr_i[26] , \m4_addr_i[27] , \m4_addr_i[28] ,
    \m4_addr_i[29] , \m4_addr_i[30] , \m4_addr_i[31] , \m5_data_i[0] ,
    \m5_data_i[1] , \m5_data_i[2] , \m5_data_i[3] , \m5_data_i[4] ,
    \m5_data_i[5] , \m5_data_i[6] , \m5_data_i[7] , \m5_data_i[8] ,
    \m5_data_i[9] , \m5_data_i[10] , \m5_data_i[11] , \m5_data_i[12] ,
    \m5_data_i[13] , \m5_data_i[14] , \m5_data_i[15] , \m5_data_i[16] ,
    \m5_data_i[17] , \m5_data_i[18] , \m5_data_i[19] , \m5_data_i[20] ,
    \m5_data_i[21] , \m5_data_i[22] , \m5_data_i[23] , \m5_data_i[24] ,
    \m5_data_i[25] , \m5_data_i[26] , \m5_data_i[27] , \m5_data_i[28] ,
    \m5_data_i[29] , \m5_data_i[30] , \m5_data_i[31] , \m5_addr_i[0] ,
    \m5_addr_i[1] , \m5_addr_i[2] , \m5_addr_i[3] , \m5_addr_i[4] ,
    \m5_addr_i[5] , \m5_addr_i[6] , \m5_addr_i[7] , \m5_addr_i[8] ,
    \m5_addr_i[9] , \m5_addr_i[10] , \m5_addr_i[11] , \m5_addr_i[12] ,
    \m5_addr_i[13] , \m5_addr_i[14] , \m5_addr_i[15] , \m5_addr_i[16] ,
    \m5_addr_i[17] , \m5_addr_i[18] , \m5_addr_i[19] , \m5_addr_i[20] ,
    \m5_addr_i[21] , \m5_addr_i[22] , \m5_addr_i[23] , \m5_addr_i[24] ,
    \m5_addr_i[25] , \m5_addr_i[26] , \m5_addr_i[27] , \m5_addr_i[28] ,
    \m5_addr_i[29] , \m5_addr_i[30] , \m5_addr_i[31] , \m6_data_i[0] ,
    \m6_data_i[1] , \m6_data_i[2] , \m6_data_i[3] , \m6_data_i[4] ,
    \m6_data_i[5] , \m6_data_i[6] , \m6_data_i[7] , \m6_data_i[8] ,
    \m6_data_i[9] , \m6_data_i[10] , \m6_data_i[11] , \m6_data_i[12] ,
    \m6_data_i[13] , \m6_data_i[14] , \m6_data_i[15] , \m6_data_i[16] ,
    \m6_data_i[17] , \m6_data_i[18] , \m6_data_i[19] , \m6_data_i[20] ,
    \m6_data_i[21] , \m6_data_i[22] , \m6_data_i[23] , \m6_data_i[24] ,
    \m6_data_i[25] , \m6_data_i[26] , \m6_data_i[27] , \m6_data_i[28] ,
    \m6_data_i[29] , \m6_data_i[30] , \m6_data_i[31] , \m6_addr_i[0] ,
    \m6_addr_i[1] , \m6_addr_i[2] , \m6_addr_i[3] , \m6_addr_i[4] ,
    \m6_addr_i[5] , \m6_addr_i[6] , \m6_addr_i[7] , \m6_addr_i[8] ,
    \m6_addr_i[9] , \m6_addr_i[10] , \m6_addr_i[11] , \m6_addr_i[12] ,
    \m6_addr_i[13] , \m6_addr_i[14] , \m6_addr_i[15] , \m6_addr_i[16] ,
    \m6_addr_i[17] , \m6_addr_i[18] , \m6_addr_i[19] , \m6_addr_i[20] ,
    \m6_addr_i[21] , \m6_addr_i[22] , \m6_addr_i[23] , \m6_addr_i[24] ,
    \m6_addr_i[25] , \m6_addr_i[26] , \m6_addr_i[27] , \m6_addr_i[28] ,
    \m6_addr_i[29] , \m6_addr_i[30] , \m6_addr_i[31] , \m7_data_i[0] ,
    \m7_data_i[1] , \m7_data_i[2] , \m7_data_i[3] , \m7_data_i[4] ,
    \m7_data_i[5] , \m7_data_i[6] , \m7_data_i[7] , \m7_data_i[8] ,
    \m7_data_i[9] , \m7_data_i[10] , \m7_data_i[11] , \m7_data_i[12] ,
    \m7_data_i[13] , \m7_data_i[14] , \m7_data_i[15] , \m7_data_i[16] ,
    \m7_data_i[17] , \m7_data_i[18] , \m7_data_i[19] , \m7_data_i[20] ,
    \m7_data_i[21] , \m7_data_i[22] , \m7_data_i[23] , \m7_data_i[24] ,
    \m7_data_i[25] , \m7_data_i[26] , \m7_data_i[27] , \m7_data_i[28] ,
    \m7_data_i[29] , \m7_data_i[30] , \m7_data_i[31] , \m7_addr_i[0] ,
    \m7_addr_i[1] , \m7_addr_i[2] , \m7_addr_i[3] , \m7_addr_i[4] ,
    \m7_addr_i[5] , \m7_addr_i[6] , \m7_addr_i[7] , \m7_addr_i[8] ,
    \m7_addr_i[9] , \m7_addr_i[10] , \m7_addr_i[11] , \m7_addr_i[12] ,
    \m7_addr_i[13] , \m7_addr_i[14] , \m7_addr_i[15] , \m7_addr_i[16] ,
    \m7_addr_i[17] , \m7_addr_i[18] , \m7_addr_i[19] , \m7_addr_i[20] ,
    \m7_addr_i[21] , \m7_addr_i[22] , \m7_addr_i[23] , \m7_addr_i[24] ,
    \m7_addr_i[25] , \m7_addr_i[26] , \m7_addr_i[27] , \m7_addr_i[28] ,
    \m7_addr_i[29] , \m7_addr_i[30] , \m7_addr_i[31] , \s0_data_i[0] ,
    \s0_data_i[1] , \s0_data_i[2] , \s0_data_i[3] , \s0_data_i[4] ,
    \s0_data_i[5] , \s0_data_i[6] , \s0_data_i[7] , \s0_data_i[8] ,
    \s0_data_i[9] , \s0_data_i[10] , \s0_data_i[11] , \s0_data_i[12] ,
    \s0_data_i[13] , \s0_data_i[14] , \s0_data_i[15] , \s0_data_i[16] ,
    \s0_data_i[17] , \s0_data_i[18] , \s0_data_i[19] , \s0_data_i[20] ,
    \s0_data_i[21] , \s0_data_i[22] , \s0_data_i[23] , \s0_data_i[24] ,
    \s0_data_i[25] , \s0_data_i[26] , \s0_data_i[27] , \s0_data_i[28] ,
    \s0_data_i[29] , \s0_data_i[30] , \s0_data_i[31] , \s1_data_i[0] ,
    \s1_data_i[1] , \s1_data_i[2] , \s1_data_i[3] , \s1_data_i[4] ,
    \s1_data_i[5] , \s1_data_i[6] , \s1_data_i[7] , \s1_data_i[8] ,
    \s1_data_i[9] , \s1_data_i[10] , \s1_data_i[11] , \s1_data_i[12] ,
    \s1_data_i[13] , \s1_data_i[14] , \s1_data_i[15] , \s1_data_i[16] ,
    \s1_data_i[17] , \s1_data_i[18] , \s1_data_i[19] , \s1_data_i[20] ,
    \s1_data_i[21] , \s1_data_i[22] , \s1_data_i[23] , \s1_data_i[24] ,
    \s1_data_i[25] , \s1_data_i[26] , \s1_data_i[27] , \s1_data_i[28] ,
    \s1_data_i[29] , \s1_data_i[30] , \s1_data_i[31] , \s2_data_i[0] ,
    \s2_data_i[1] , \s2_data_i[2] , \s2_data_i[3] , \s2_data_i[4] ,
    \s2_data_i[5] , \s2_data_i[6] , \s2_data_i[7] , \s2_data_i[8] ,
    \s2_data_i[9] , \s2_data_i[10] , \s2_data_i[11] , \s2_data_i[12] ,
    \s2_data_i[13] , \s2_data_i[14] , \s2_data_i[15] , \s2_data_i[16] ,
    \s2_data_i[17] , \s2_data_i[18] , \s2_data_i[19] , \s2_data_i[20] ,
    \s2_data_i[21] , \s2_data_i[22] , \s2_data_i[23] , \s2_data_i[24] ,
    \s2_data_i[25] , \s2_data_i[26] , \s2_data_i[27] , \s2_data_i[28] ,
    \s2_data_i[29] , \s2_data_i[30] , \s2_data_i[31] , \s3_data_i[0] ,
    \s3_data_i[1] , \s3_data_i[2] , \s3_data_i[3] , \s3_data_i[4] ,
    \s3_data_i[5] , \s3_data_i[6] , \s3_data_i[7] , \s3_data_i[8] ,
    \s3_data_i[9] , \s3_data_i[10] , \s3_data_i[11] , \s3_data_i[12] ,
    \s3_data_i[13] , \s3_data_i[14] , \s3_data_i[15] , \s3_data_i[16] ,
    \s3_data_i[17] , \s3_data_i[18] , \s3_data_i[19] , \s3_data_i[20] ,
    \s3_data_i[21] , \s3_data_i[22] , \s3_data_i[23] , \s3_data_i[24] ,
    \s3_data_i[25] , \s3_data_i[26] , \s3_data_i[27] , \s3_data_i[28] ,
    \s3_data_i[29] , \s3_data_i[30] , \s3_data_i[31] , \s4_data_i[0] ,
    \s4_data_i[1] , \s4_data_i[2] , \s4_data_i[3] , \s4_data_i[4] ,
    \s4_data_i[5] , \s4_data_i[6] , \s4_data_i[7] , \s4_data_i[8] ,
    \s4_data_i[9] , \s4_data_i[10] , \s4_data_i[11] , \s4_data_i[12] ,
    \s4_data_i[13] , \s4_data_i[14] , \s4_data_i[15] , \s4_data_i[16] ,
    \s4_data_i[17] , \s4_data_i[18] , \s4_data_i[19] , \s4_data_i[20] ,
    \s4_data_i[21] , \s4_data_i[22] , \s4_data_i[23] , \s4_data_i[24] ,
    \s4_data_i[25] , \s4_data_i[26] , \s4_data_i[27] , \s4_data_i[28] ,
    \s4_data_i[29] , \s4_data_i[30] , \s4_data_i[31] , \s5_data_i[0] ,
    \s5_data_i[1] , \s5_data_i[2] , \s5_data_i[3] , \s5_data_i[4] ,
    \s5_data_i[5] , \s5_data_i[6] , \s5_data_i[7] , \s5_data_i[8] ,
    \s5_data_i[9] , \s5_data_i[10] , \s5_data_i[11] , \s5_data_i[12] ,
    \s5_data_i[13] , \s5_data_i[14] , \s5_data_i[15] , \s5_data_i[16] ,
    \s5_data_i[17] , \s5_data_i[18] , \s5_data_i[19] , \s5_data_i[20] ,
    \s5_data_i[21] , \s5_data_i[22] , \s5_data_i[23] , \s5_data_i[24] ,
    \s5_data_i[25] , \s5_data_i[26] , \s5_data_i[27] , \s5_data_i[28] ,
    \s5_data_i[29] , \s5_data_i[30] , \s5_data_i[31] , \s6_data_i[0] ,
    \s6_data_i[1] , \s6_data_i[2] , \s6_data_i[3] , \s6_data_i[4] ,
    \s6_data_i[5] , \s6_data_i[6] , \s6_data_i[7] , \s6_data_i[8] ,
    \s6_data_i[9] , \s6_data_i[10] , \s6_data_i[11] , \s6_data_i[12] ,
    \s6_data_i[13] , \s6_data_i[14] , \s6_data_i[15] , \s6_data_i[16] ,
    \s6_data_i[17] , \s6_data_i[18] , \s6_data_i[19] , \s6_data_i[20] ,
    \s6_data_i[21] , \s6_data_i[22] , \s6_data_i[23] , \s6_data_i[24] ,
    \s6_data_i[25] , \s6_data_i[26] , \s6_data_i[27] , \s6_data_i[28] ,
    \s6_data_i[29] , \s6_data_i[30] , \s6_data_i[31] , \s7_data_i[0] ,
    \s7_data_i[1] , \s7_data_i[2] , \s7_data_i[3] , \s7_data_i[4] ,
    \s7_data_i[5] , \s7_data_i[6] , \s7_data_i[7] , \s7_data_i[8] ,
    \s7_data_i[9] , \s7_data_i[10] , \s7_data_i[11] , \s7_data_i[12] ,
    \s7_data_i[13] , \s7_data_i[14] , \s7_data_i[15] , \s7_data_i[16] ,
    \s7_data_i[17] , \s7_data_i[18] , \s7_data_i[19] , \s7_data_i[20] ,
    \s7_data_i[21] , \s7_data_i[22] , \s7_data_i[23] , \s7_data_i[24] ,
    \s7_data_i[25] , \s7_data_i[26] , \s7_data_i[27] , \s7_data_i[28] ,
    \s7_data_i[29] , \s7_data_i[30] , \s7_data_i[31] , \s8_data_i[0] ,
    \s8_data_i[1] , \s8_data_i[2] , \s8_data_i[3] , \s8_data_i[4] ,
    \s8_data_i[5] , \s8_data_i[6] , \s8_data_i[7] , \s8_data_i[8] ,
    \s8_data_i[9] , \s8_data_i[10] , \s8_data_i[11] , \s8_data_i[12] ,
    \s8_data_i[13] , \s8_data_i[14] , \s8_data_i[15] , \s8_data_i[16] ,
    \s8_data_i[17] , \s8_data_i[18] , \s8_data_i[19] , \s8_data_i[20] ,
    \s8_data_i[21] , \s8_data_i[22] , \s8_data_i[23] , \s8_data_i[24] ,
    \s8_data_i[25] , \s8_data_i[26] , \s8_data_i[27] , \s8_data_i[28] ,
    \s8_data_i[29] , \s8_data_i[30] , \s8_data_i[31] , \s9_data_i[0] ,
    \s9_data_i[1] , \s9_data_i[2] , \s9_data_i[3] , \s9_data_i[4] ,
    \s9_data_i[5] , \s9_data_i[6] , \s9_data_i[7] , \s9_data_i[8] ,
    \s9_data_i[9] , \s9_data_i[10] , \s9_data_i[11] , \s9_data_i[12] ,
    \s9_data_i[13] , \s9_data_i[14] , \s9_data_i[15] , \s9_data_i[16] ,
    \s9_data_i[17] , \s9_data_i[18] , \s9_data_i[19] , \s9_data_i[20] ,
    \s9_data_i[21] , \s9_data_i[22] , \s9_data_i[23] , \s9_data_i[24] ,
    \s9_data_i[25] , \s9_data_i[26] , \s9_data_i[27] , \s9_data_i[28] ,
    \s9_data_i[29] , \s9_data_i[30] , \s9_data_i[31] , \s10_data_i[0] ,
    \s10_data_i[1] , \s10_data_i[2] , \s10_data_i[3] , \s10_data_i[4] ,
    \s10_data_i[5] , \s10_data_i[6] , \s10_data_i[7] , \s10_data_i[8] ,
    \s10_data_i[9] , \s10_data_i[10] , \s10_data_i[11] , \s10_data_i[12] ,
    \s10_data_i[13] , \s10_data_i[14] , \s10_data_i[15] , \s10_data_i[16] ,
    \s10_data_i[17] , \s10_data_i[18] , \s10_data_i[19] , \s10_data_i[20] ,
    \s10_data_i[21] , \s10_data_i[22] , \s10_data_i[23] , \s10_data_i[24] ,
    \s10_data_i[25] , \s10_data_i[26] , \s10_data_i[27] , \s10_data_i[28] ,
    \s10_data_i[29] , \s10_data_i[30] , \s10_data_i[31] , \s11_data_i[0] ,
    \s11_data_i[1] , \s11_data_i[2] , \s11_data_i[3] , \s11_data_i[4] ,
    \s11_data_i[5] , \s11_data_i[6] , \s11_data_i[7] , \s11_data_i[8] ,
    \s11_data_i[9] , \s11_data_i[10] , \s11_data_i[11] , \s11_data_i[12] ,
    \s11_data_i[13] , \s11_data_i[14] , \s11_data_i[15] , \s11_data_i[16] ,
    \s11_data_i[17] , \s11_data_i[18] , \s11_data_i[19] , \s11_data_i[20] ,
    \s11_data_i[21] , \s11_data_i[22] , \s11_data_i[23] , \s11_data_i[24] ,
    \s11_data_i[25] , \s11_data_i[26] , \s11_data_i[27] , \s11_data_i[28] ,
    \s11_data_i[29] , \s11_data_i[30] , \s11_data_i[31] , \s12_data_i[0] ,
    \s12_data_i[1] , \s12_data_i[2] , \s12_data_i[3] , \s12_data_i[4] ,
    \s12_data_i[5] , \s12_data_i[6] , \s12_data_i[7] , \s12_data_i[8] ,
    \s12_data_i[9] , \s12_data_i[10] , \s12_data_i[11] , \s12_data_i[12] ,
    \s12_data_i[13] , \s12_data_i[14] , \s12_data_i[15] , \s12_data_i[16] ,
    \s12_data_i[17] , \s12_data_i[18] , \s12_data_i[19] , \s12_data_i[20] ,
    \s12_data_i[21] , \s12_data_i[22] , \s12_data_i[23] , \s12_data_i[24] ,
    \s12_data_i[25] , \s12_data_i[26] , \s12_data_i[27] , \s12_data_i[28] ,
    \s12_data_i[29] , \s12_data_i[30] , \s12_data_i[31] , \s13_data_i[0] ,
    \s13_data_i[1] , \s13_data_i[2] , \s13_data_i[3] , \s13_data_i[4] ,
    \s13_data_i[5] , \s13_data_i[6] , \s13_data_i[7] , \s13_data_i[8] ,
    \s13_data_i[9] , \s13_data_i[10] , \s13_data_i[11] , \s13_data_i[12] ,
    \s13_data_i[13] , \s13_data_i[14] , \s13_data_i[15] , \s13_data_i[16] ,
    \s13_data_i[17] , \s13_data_i[18] , \s13_data_i[19] , \s13_data_i[20] ,
    \s13_data_i[21] , \s13_data_i[22] , \s13_data_i[23] , \s13_data_i[24] ,
    \s13_data_i[25] , \s13_data_i[26] , \s13_data_i[27] , \s13_data_i[28] ,
    \s13_data_i[29] , \s13_data_i[30] , \s13_data_i[31] , \s14_data_i[0] ,
    \s14_data_i[1] , \s14_data_i[2] , \s14_data_i[3] , \s14_data_i[4] ,
    \s14_data_i[5] , \s14_data_i[6] , \s14_data_i[7] , \s14_data_i[8] ,
    \s14_data_i[9] , \s14_data_i[10] , \s14_data_i[11] , \s14_data_i[12] ,
    \s14_data_i[13] , \s14_data_i[14] , \s14_data_i[15] , \s14_data_i[16] ,
    \s14_data_i[17] , \s14_data_i[18] , \s14_data_i[19] , \s14_data_i[20] ,
    \s14_data_i[21] , \s14_data_i[22] , \s14_data_i[23] , \s14_data_i[24] ,
    \s14_data_i[25] , \s14_data_i[26] , \s14_data_i[27] , \s14_data_i[28] ,
    \s14_data_i[29] , \s14_data_i[30] , \s14_data_i[31] , \s15_data_i[0] ,
    \s15_data_i[1] , \s15_data_i[2] , \s15_data_i[3] , \s15_data_i[4] ,
    \s15_data_i[5] , \s15_data_i[6] , \s15_data_i[7] , \s15_data_i[8] ,
    \s15_data_i[9] , \s15_data_i[10] , \s15_data_i[11] , \s15_data_i[12] ,
    \s15_data_i[13] , \s15_data_i[14] , \s15_data_i[15] , \s15_data_i[16] ,
    \s15_data_i[17] , \s15_data_i[18] , \s15_data_i[19] , \s15_data_i[20] ,
    \s15_data_i[21] , \s15_data_i[22] , \s15_data_i[23] , \s15_data_i[24] ,
    \s15_data_i[25] , \s15_data_i[26] , \s15_data_i[27] , \s15_data_i[28] ,
    \s15_data_i[29] , \s15_data_i[30] , \s15_data_i[31] , \m0_sel_i[0] ,
    \m0_sel_i[1] , \m0_sel_i[2] , \m0_sel_i[3] , \m1_sel_i[0] ,
    \m1_sel_i[1] , \m1_sel_i[2] , \m1_sel_i[3] , \m2_sel_i[0] ,
    \m2_sel_i[1] , \m2_sel_i[2] , \m2_sel_i[3] , \m3_sel_i[0] ,
    \m3_sel_i[1] , \m3_sel_i[2] , \m3_sel_i[3] , \m4_sel_i[0] ,
    \m4_sel_i[1] , \m4_sel_i[2] , \m4_sel_i[3] , \m5_sel_i[0] ,
    \m5_sel_i[1] , \m5_sel_i[2] , \m5_sel_i[3] , \m6_sel_i[0] ,
    \m6_sel_i[1] , \m6_sel_i[2] , \m6_sel_i[3] , \m7_sel_i[0] ,
    \m7_sel_i[1] , \m7_sel_i[2] , \m7_sel_i[3] ,
    \m0_data_o[0] , \m0_data_o[1] , \m0_data_o[2] , \m0_data_o[3] ,
    \m0_data_o[4] , \m0_data_o[5] , \m0_data_o[6] , \m0_data_o[7] ,
    \m0_data_o[8] , \m0_data_o[9] , \m0_data_o[10] , \m0_data_o[11] ,
    \m0_data_o[12] , \m0_data_o[13] , \m0_data_o[14] , \m0_data_o[15] ,
    \m0_data_o[16] , \m0_data_o[17] , \m0_data_o[18] , \m0_data_o[19] ,
    \m0_data_o[20] , \m0_data_o[21] , \m0_data_o[22] , \m0_data_o[23] ,
    \m0_data_o[24] , \m0_data_o[25] , \m0_data_o[26] , \m0_data_o[27] ,
    \m0_data_o[28] , \m0_data_o[29] , \m0_data_o[30] , \m0_data_o[31] ,
    \m1_data_o[0] , \m1_data_o[1] , \m1_data_o[2] , \m1_data_o[3] ,
    \m1_data_o[4] , \m1_data_o[5] , \m1_data_o[6] , \m1_data_o[7] ,
    \m1_data_o[8] , \m1_data_o[9] , \m1_data_o[10] , \m1_data_o[11] ,
    \m1_data_o[12] , \m1_data_o[13] , \m1_data_o[14] , \m1_data_o[15] ,
    \m1_data_o[16] , \m1_data_o[17] , \m1_data_o[18] , \m1_data_o[19] ,
    \m1_data_o[20] , \m1_data_o[21] , \m1_data_o[22] , \m1_data_o[23] ,
    \m1_data_o[24] , \m1_data_o[25] , \m1_data_o[26] , \m1_data_o[27] ,
    \m1_data_o[28] , \m1_data_o[29] , \m1_data_o[30] , \m1_data_o[31] ,
    \m2_data_o[0] , \m2_data_o[1] , \m2_data_o[2] , \m2_data_o[3] ,
    \m2_data_o[4] , \m2_data_o[5] , \m2_data_o[6] , \m2_data_o[7] ,
    \m2_data_o[8] , \m2_data_o[9] , \m2_data_o[10] , \m2_data_o[11] ,
    \m2_data_o[12] , \m2_data_o[13] , \m2_data_o[14] , \m2_data_o[15] ,
    \m2_data_o[16] , \m2_data_o[17] , \m2_data_o[18] , \m2_data_o[19] ,
    \m2_data_o[20] , \m2_data_o[21] , \m2_data_o[22] , \m2_data_o[23] ,
    \m2_data_o[24] , \m2_data_o[25] , \m2_data_o[26] , \m2_data_o[27] ,
    \m2_data_o[28] , \m2_data_o[29] , \m2_data_o[30] , \m2_data_o[31] ,
    \m3_data_o[0] , \m3_data_o[1] , \m3_data_o[2] , \m3_data_o[3] ,
    \m3_data_o[4] , \m3_data_o[5] , \m3_data_o[6] , \m3_data_o[7] ,
    \m3_data_o[8] , \m3_data_o[9] , \m3_data_o[10] , \m3_data_o[11] ,
    \m3_data_o[12] , \m3_data_o[13] , \m3_data_o[14] , \m3_data_o[15] ,
    \m3_data_o[16] , \m3_data_o[17] , \m3_data_o[18] , \m3_data_o[19] ,
    \m3_data_o[20] , \m3_data_o[21] , \m3_data_o[22] , \m3_data_o[23] ,
    \m3_data_o[24] , \m3_data_o[25] , \m3_data_o[26] , \m3_data_o[27] ,
    \m3_data_o[28] , \m3_data_o[29] , \m3_data_o[30] , \m3_data_o[31] ,
    \m4_data_o[0] , \m4_data_o[1] , \m4_data_o[2] , \m4_data_o[3] ,
    \m4_data_o[4] , \m4_data_o[5] , \m4_data_o[6] , \m4_data_o[7] ,
    \m4_data_o[8] , \m4_data_o[9] , \m4_data_o[10] , \m4_data_o[11] ,
    \m4_data_o[12] , \m4_data_o[13] , \m4_data_o[14] , \m4_data_o[15] ,
    \m4_data_o[16] , \m4_data_o[17] , \m4_data_o[18] , \m4_data_o[19] ,
    \m4_data_o[20] , \m4_data_o[21] , \m4_data_o[22] , \m4_data_o[23] ,
    \m4_data_o[24] , \m4_data_o[25] , \m4_data_o[26] , \m4_data_o[27] ,
    \m4_data_o[28] , \m4_data_o[29] , \m4_data_o[30] , \m4_data_o[31] ,
    \m5_data_o[0] , \m5_data_o[1] , \m5_data_o[2] , \m5_data_o[3] ,
    \m5_data_o[4] , \m5_data_o[5] , \m5_data_o[6] , \m5_data_o[7] ,
    \m5_data_o[8] , \m5_data_o[9] , \m5_data_o[10] , \m5_data_o[11] ,
    \m5_data_o[12] , \m5_data_o[13] , \m5_data_o[14] , \m5_data_o[15] ,
    \m5_data_o[16] , \m5_data_o[17] , \m5_data_o[18] , \m5_data_o[19] ,
    \m5_data_o[20] , \m5_data_o[21] , \m5_data_o[22] , \m5_data_o[23] ,
    \m5_data_o[24] , \m5_data_o[25] , \m5_data_o[26] , \m5_data_o[27] ,
    \m5_data_o[28] , \m5_data_o[29] , \m5_data_o[30] , \m5_data_o[31] ,
    \m6_data_o[0] , \m6_data_o[1] , \m6_data_o[2] , \m6_data_o[3] ,
    \m6_data_o[4] , \m6_data_o[5] , \m6_data_o[6] , \m6_data_o[7] ,
    \m6_data_o[8] , \m6_data_o[9] , \m6_data_o[10] , \m6_data_o[11] ,
    \m6_data_o[12] , \m6_data_o[13] , \m6_data_o[14] , \m6_data_o[15] ,
    \m6_data_o[16] , \m6_data_o[17] , \m6_data_o[18] , \m6_data_o[19] ,
    \m6_data_o[20] , \m6_data_o[21] , \m6_data_o[22] , \m6_data_o[23] ,
    \m6_data_o[24] , \m6_data_o[25] , \m6_data_o[26] , \m6_data_o[27] ,
    \m6_data_o[28] , \m6_data_o[29] , \m6_data_o[30] , \m6_data_o[31] ,
    \m7_data_o[0] , \m7_data_o[1] , \m7_data_o[2] , \m7_data_o[3] ,
    \m7_data_o[4] , \m7_data_o[5] , \m7_data_o[6] , \m7_data_o[7] ,
    \m7_data_o[8] , \m7_data_o[9] , \m7_data_o[10] , \m7_data_o[11] ,
    \m7_data_o[12] , \m7_data_o[13] , \m7_data_o[14] , \m7_data_o[15] ,
    \m7_data_o[16] , \m7_data_o[17] , \m7_data_o[18] , \m7_data_o[19] ,
    \m7_data_o[20] , \m7_data_o[21] , \m7_data_o[22] , \m7_data_o[23] ,
    \m7_data_o[24] , \m7_data_o[25] , \m7_data_o[26] , \m7_data_o[27] ,
    \m7_data_o[28] , \m7_data_o[29] , \m7_data_o[30] , \m7_data_o[31] ,
    \s0_data_o[0] , \s0_data_o[1] , \s0_data_o[2] , \s0_data_o[3] ,
    \s0_data_o[4] , \s0_data_o[5] , \s0_data_o[6] , \s0_data_o[7] ,
    \s0_data_o[8] , \s0_data_o[9] , \s0_data_o[10] , \s0_data_o[11] ,
    \s0_data_o[12] , \s0_data_o[13] , \s0_data_o[14] , \s0_data_o[15] ,
    \s0_data_o[16] , \s0_data_o[17] , \s0_data_o[18] , \s0_data_o[19] ,
    \s0_data_o[20] , \s0_data_o[21] , \s0_data_o[22] , \s0_data_o[23] ,
    \s0_data_o[24] , \s0_data_o[25] , \s0_data_o[26] , \s0_data_o[27] ,
    \s0_data_o[28] , \s0_data_o[29] , \s0_data_o[30] , \s0_data_o[31] ,
    \s0_addr_o[0] , \s0_addr_o[1] , \s0_addr_o[2] , \s0_addr_o[3] ,
    \s0_addr_o[4] , \s0_addr_o[5] , \s0_addr_o[6] , \s0_addr_o[7] ,
    \s0_addr_o[8] , \s0_addr_o[9] , \s0_addr_o[10] , \s0_addr_o[11] ,
    \s0_addr_o[12] , \s0_addr_o[13] , \s0_addr_o[14] , \s0_addr_o[15] ,
    \s0_addr_o[16] , \s0_addr_o[17] , \s0_addr_o[18] , \s0_addr_o[19] ,
    \s0_addr_o[20] , \s0_addr_o[21] , \s0_addr_o[22] , \s0_addr_o[23] ,
    \s0_addr_o[24] , \s0_addr_o[25] , \s0_addr_o[26] , \s0_addr_o[27] ,
    \s0_addr_o[28] , \s0_addr_o[29] , \s0_addr_o[30] , \s0_addr_o[31] ,
    \s1_data_o[0] , \s1_data_o[1] , \s1_data_o[2] , \s1_data_o[3] ,
    \s1_data_o[4] , \s1_data_o[5] , \s1_data_o[6] , \s1_data_o[7] ,
    \s1_data_o[8] , \s1_data_o[9] , \s1_data_o[10] , \s1_data_o[11] ,
    \s1_data_o[12] , \s1_data_o[13] , \s1_data_o[14] , \s1_data_o[15] ,
    \s1_data_o[16] , \s1_data_o[17] , \s1_data_o[18] , \s1_data_o[19] ,
    \s1_data_o[20] , \s1_data_o[21] , \s1_data_o[22] , \s1_data_o[23] ,
    \s1_data_o[24] , \s1_data_o[25] , \s1_data_o[26] , \s1_data_o[27] ,
    \s1_data_o[28] , \s1_data_o[29] , \s1_data_o[30] , \s1_data_o[31] ,
    \s1_addr_o[0] , \s1_addr_o[1] , \s1_addr_o[2] , \s1_addr_o[3] ,
    \s1_addr_o[4] , \s1_addr_o[5] , \s1_addr_o[6] , \s1_addr_o[7] ,
    \s1_addr_o[8] , \s1_addr_o[9] , \s1_addr_o[10] , \s1_addr_o[11] ,
    \s1_addr_o[12] , \s1_addr_o[13] , \s1_addr_o[14] , \s1_addr_o[15] ,
    \s1_addr_o[16] , \s1_addr_o[17] , \s1_addr_o[18] , \s1_addr_o[19] ,
    \s1_addr_o[20] , \s1_addr_o[21] , \s1_addr_o[22] , \s1_addr_o[23] ,
    \s1_addr_o[24] , \s1_addr_o[25] , \s1_addr_o[26] , \s1_addr_o[27] ,
    \s1_addr_o[28] , \s1_addr_o[29] , \s1_addr_o[30] , \s1_addr_o[31] ,
    \s2_data_o[0] , \s2_data_o[1] , \s2_data_o[2] , \s2_data_o[3] ,
    \s2_data_o[4] , \s2_data_o[5] , \s2_data_o[6] , \s2_data_o[7] ,
    \s2_data_o[8] , \s2_data_o[9] , \s2_data_o[10] , \s2_data_o[11] ,
    \s2_data_o[12] , \s2_data_o[13] , \s2_data_o[14] , \s2_data_o[15] ,
    \s2_data_o[16] , \s2_data_o[17] , \s2_data_o[18] , \s2_data_o[19] ,
    \s2_data_o[20] , \s2_data_o[21] , \s2_data_o[22] , \s2_data_o[23] ,
    \s2_data_o[24] , \s2_data_o[25] , \s2_data_o[26] , \s2_data_o[27] ,
    \s2_data_o[28] , \s2_data_o[29] , \s2_data_o[30] , \s2_data_o[31] ,
    \s2_addr_o[0] , \s2_addr_o[1] , \s2_addr_o[2] , \s2_addr_o[3] ,
    \s2_addr_o[4] , \s2_addr_o[5] , \s2_addr_o[6] , \s2_addr_o[7] ,
    \s2_addr_o[8] , \s2_addr_o[9] , \s2_addr_o[10] , \s2_addr_o[11] ,
    \s2_addr_o[12] , \s2_addr_o[13] , \s2_addr_o[14] , \s2_addr_o[15] ,
    \s2_addr_o[16] , \s2_addr_o[17] , \s2_addr_o[18] , \s2_addr_o[19] ,
    \s2_addr_o[20] , \s2_addr_o[21] , \s2_addr_o[22] , \s2_addr_o[23] ,
    \s2_addr_o[24] , \s2_addr_o[25] , \s2_addr_o[26] , \s2_addr_o[27] ,
    \s2_addr_o[28] , \s2_addr_o[29] , \s2_addr_o[30] , \s2_addr_o[31] ,
    \s3_data_o[0] , \s3_data_o[1] , \s3_data_o[2] , \s3_data_o[3] ,
    \s3_data_o[4] , \s3_data_o[5] , \s3_data_o[6] , \s3_data_o[7] ,
    \s3_data_o[8] , \s3_data_o[9] , \s3_data_o[10] , \s3_data_o[11] ,
    \s3_data_o[12] , \s3_data_o[13] , \s3_data_o[14] , \s3_data_o[15] ,
    \s3_data_o[16] , \s3_data_o[17] , \s3_data_o[18] , \s3_data_o[19] ,
    \s3_data_o[20] , \s3_data_o[21] , \s3_data_o[22] , \s3_data_o[23] ,
    \s3_data_o[24] , \s3_data_o[25] , \s3_data_o[26] , \s3_data_o[27] ,
    \s3_data_o[28] , \s3_data_o[29] , \s3_data_o[30] , \s3_data_o[31] ,
    \s3_addr_o[0] , \s3_addr_o[1] , \s3_addr_o[2] , \s3_addr_o[3] ,
    \s3_addr_o[4] , \s3_addr_o[5] , \s3_addr_o[6] , \s3_addr_o[7] ,
    \s3_addr_o[8] , \s3_addr_o[9] , \s3_addr_o[10] , \s3_addr_o[11] ,
    \s3_addr_o[12] , \s3_addr_o[13] , \s3_addr_o[14] , \s3_addr_o[15] ,
    \s3_addr_o[16] , \s3_addr_o[17] , \s3_addr_o[18] , \s3_addr_o[19] ,
    \s3_addr_o[20] , \s3_addr_o[21] , \s3_addr_o[22] , \s3_addr_o[23] ,
    \s3_addr_o[24] , \s3_addr_o[25] , \s3_addr_o[26] , \s3_addr_o[27] ,
    \s3_addr_o[28] , \s3_addr_o[29] , \s3_addr_o[30] , \s3_addr_o[31] ,
    \s4_data_o[0] , \s4_data_o[1] , \s4_data_o[2] , \s4_data_o[3] ,
    \s4_data_o[4] , \s4_data_o[5] , \s4_data_o[6] , \s4_data_o[7] ,
    \s4_data_o[8] , \s4_data_o[9] , \s4_data_o[10] , \s4_data_o[11] ,
    \s4_data_o[12] , \s4_data_o[13] , \s4_data_o[14] , \s4_data_o[15] ,
    \s4_data_o[16] , \s4_data_o[17] , \s4_data_o[18] , \s4_data_o[19] ,
    \s4_data_o[20] , \s4_data_o[21] , \s4_data_o[22] , \s4_data_o[23] ,
    \s4_data_o[24] , \s4_data_o[25] , \s4_data_o[26] , \s4_data_o[27] ,
    \s4_data_o[28] , \s4_data_o[29] , \s4_data_o[30] , \s4_data_o[31] ,
    \s4_addr_o[0] , \s4_addr_o[1] , \s4_addr_o[2] , \s4_addr_o[3] ,
    \s4_addr_o[4] , \s4_addr_o[5] , \s4_addr_o[6] , \s4_addr_o[7] ,
    \s4_addr_o[8] , \s4_addr_o[9] , \s4_addr_o[10] , \s4_addr_o[11] ,
    \s4_addr_o[12] , \s4_addr_o[13] , \s4_addr_o[14] , \s4_addr_o[15] ,
    \s4_addr_o[16] , \s4_addr_o[17] , \s4_addr_o[18] , \s4_addr_o[19] ,
    \s4_addr_o[20] , \s4_addr_o[21] , \s4_addr_o[22] , \s4_addr_o[23] ,
    \s4_addr_o[24] , \s4_addr_o[25] , \s4_addr_o[26] , \s4_addr_o[27] ,
    \s4_addr_o[28] , \s4_addr_o[29] , \s4_addr_o[30] , \s4_addr_o[31] ,
    \s5_data_o[0] , \s5_data_o[1] , \s5_data_o[2] , \s5_data_o[3] ,
    \s5_data_o[4] , \s5_data_o[5] , \s5_data_o[6] , \s5_data_o[7] ,
    \s5_data_o[8] , \s5_data_o[9] , \s5_data_o[10] , \s5_data_o[11] ,
    \s5_data_o[12] , \s5_data_o[13] , \s5_data_o[14] , \s5_data_o[15] ,
    \s5_data_o[16] , \s5_data_o[17] , \s5_data_o[18] , \s5_data_o[19] ,
    \s5_data_o[20] , \s5_data_o[21] , \s5_data_o[22] , \s5_data_o[23] ,
    \s5_data_o[24] , \s5_data_o[25] , \s5_data_o[26] , \s5_data_o[27] ,
    \s5_data_o[28] , \s5_data_o[29] , \s5_data_o[30] , \s5_data_o[31] ,
    \s5_addr_o[0] , \s5_addr_o[1] , \s5_addr_o[2] , \s5_addr_o[3] ,
    \s5_addr_o[4] , \s5_addr_o[5] , \s5_addr_o[6] , \s5_addr_o[7] ,
    \s5_addr_o[8] , \s5_addr_o[9] , \s5_addr_o[10] , \s5_addr_o[11] ,
    \s5_addr_o[12] , \s5_addr_o[13] , \s5_addr_o[14] , \s5_addr_o[15] ,
    \s5_addr_o[16] , \s5_addr_o[17] , \s5_addr_o[18] , \s5_addr_o[19] ,
    \s5_addr_o[20] , \s5_addr_o[21] , \s5_addr_o[22] , \s5_addr_o[23] ,
    \s5_addr_o[24] , \s5_addr_o[25] , \s5_addr_o[26] , \s5_addr_o[27] ,
    \s5_addr_o[28] , \s5_addr_o[29] , \s5_addr_o[30] , \s5_addr_o[31] ,
    \s6_data_o[0] , \s6_data_o[1] , \s6_data_o[2] , \s6_data_o[3] ,
    \s6_data_o[4] , \s6_data_o[5] , \s6_data_o[6] , \s6_data_o[7] ,
    \s6_data_o[8] , \s6_data_o[9] , \s6_data_o[10] , \s6_data_o[11] ,
    \s6_data_o[12] , \s6_data_o[13] , \s6_data_o[14] , \s6_data_o[15] ,
    \s6_data_o[16] , \s6_data_o[17] , \s6_data_o[18] , \s6_data_o[19] ,
    \s6_data_o[20] , \s6_data_o[21] , \s6_data_o[22] , \s6_data_o[23] ,
    \s6_data_o[24] , \s6_data_o[25] , \s6_data_o[26] , \s6_data_o[27] ,
    \s6_data_o[28] , \s6_data_o[29] , \s6_data_o[30] , \s6_data_o[31] ,
    \s6_addr_o[0] , \s6_addr_o[1] , \s6_addr_o[2] , \s6_addr_o[3] ,
    \s6_addr_o[4] , \s6_addr_o[5] , \s6_addr_o[6] , \s6_addr_o[7] ,
    \s6_addr_o[8] , \s6_addr_o[9] , \s6_addr_o[10] , \s6_addr_o[11] ,
    \s6_addr_o[12] , \s6_addr_o[13] , \s6_addr_o[14] , \s6_addr_o[15] ,
    \s6_addr_o[16] , \s6_addr_o[17] , \s6_addr_o[18] , \s6_addr_o[19] ,
    \s6_addr_o[20] , \s6_addr_o[21] , \s6_addr_o[22] , \s6_addr_o[23] ,
    \s6_addr_o[24] , \s6_addr_o[25] , \s6_addr_o[26] , \s6_addr_o[27] ,
    \s6_addr_o[28] , \s6_addr_o[29] , \s6_addr_o[30] , \s6_addr_o[31] ,
    \s7_data_o[0] , \s7_data_o[1] , \s7_data_o[2] , \s7_data_o[3] ,
    \s7_data_o[4] , \s7_data_o[5] , \s7_data_o[6] , \s7_data_o[7] ,
    \s7_data_o[8] , \s7_data_o[9] , \s7_data_o[10] , \s7_data_o[11] ,
    \s7_data_o[12] , \s7_data_o[13] , \s7_data_o[14] , \s7_data_o[15] ,
    \s7_data_o[16] , \s7_data_o[17] , \s7_data_o[18] , \s7_data_o[19] ,
    \s7_data_o[20] , \s7_data_o[21] , \s7_data_o[22] , \s7_data_o[23] ,
    \s7_data_o[24] , \s7_data_o[25] , \s7_data_o[26] , \s7_data_o[27] ,
    \s7_data_o[28] , \s7_data_o[29] , \s7_data_o[30] , \s7_data_o[31] ,
    \s7_addr_o[0] , \s7_addr_o[1] , \s7_addr_o[2] , \s7_addr_o[3] ,
    \s7_addr_o[4] , \s7_addr_o[5] , \s7_addr_o[6] , \s7_addr_o[7] ,
    \s7_addr_o[8] , \s7_addr_o[9] , \s7_addr_o[10] , \s7_addr_o[11] ,
    \s7_addr_o[12] , \s7_addr_o[13] , \s7_addr_o[14] , \s7_addr_o[15] ,
    \s7_addr_o[16] , \s7_addr_o[17] , \s7_addr_o[18] , \s7_addr_o[19] ,
    \s7_addr_o[20] , \s7_addr_o[21] , \s7_addr_o[22] , \s7_addr_o[23] ,
    \s7_addr_o[24] , \s7_addr_o[25] , \s7_addr_o[26] , \s7_addr_o[27] ,
    \s7_addr_o[28] , \s7_addr_o[29] , \s7_addr_o[30] , \s7_addr_o[31] ,
    \s8_data_o[0] , \s8_data_o[1] , \s8_data_o[2] , \s8_data_o[3] ,
    \s8_data_o[4] , \s8_data_o[5] , \s8_data_o[6] , \s8_data_o[7] ,
    \s8_data_o[8] , \s8_data_o[9] , \s8_data_o[10] , \s8_data_o[11] ,
    \s8_data_o[12] , \s8_data_o[13] , \s8_data_o[14] , \s8_data_o[15] ,
    \s8_data_o[16] , \s8_data_o[17] , \s8_data_o[18] , \s8_data_o[19] ,
    \s8_data_o[20] , \s8_data_o[21] , \s8_data_o[22] , \s8_data_o[23] ,
    \s8_data_o[24] , \s8_data_o[25] , \s8_data_o[26] , \s8_data_o[27] ,
    \s8_data_o[28] , \s8_data_o[29] , \s8_data_o[30] , \s8_data_o[31] ,
    \s8_addr_o[0] , \s8_addr_o[1] , \s8_addr_o[2] , \s8_addr_o[3] ,
    \s8_addr_o[4] , \s8_addr_o[5] , \s8_addr_o[6] , \s8_addr_o[7] ,
    \s8_addr_o[8] , \s8_addr_o[9] , \s8_addr_o[10] , \s8_addr_o[11] ,
    \s8_addr_o[12] , \s8_addr_o[13] , \s8_addr_o[14] , \s8_addr_o[15] ,
    \s8_addr_o[16] , \s8_addr_o[17] , \s8_addr_o[18] , \s8_addr_o[19] ,
    \s8_addr_o[20] , \s8_addr_o[21] , \s8_addr_o[22] , \s8_addr_o[23] ,
    \s8_addr_o[24] , \s8_addr_o[25] , \s8_addr_o[26] , \s8_addr_o[27] ,
    \s8_addr_o[28] , \s8_addr_o[29] , \s8_addr_o[30] , \s8_addr_o[31] ,
    \s9_data_o[0] , \s9_data_o[1] , \s9_data_o[2] , \s9_data_o[3] ,
    \s9_data_o[4] , \s9_data_o[5] , \s9_data_o[6] , \s9_data_o[7] ,
    \s9_data_o[8] , \s9_data_o[9] , \s9_data_o[10] , \s9_data_o[11] ,
    \s9_data_o[12] , \s9_data_o[13] , \s9_data_o[14] , \s9_data_o[15] ,
    \s9_data_o[16] , \s9_data_o[17] , \s9_data_o[18] , \s9_data_o[19] ,
    \s9_data_o[20] , \s9_data_o[21] , \s9_data_o[22] , \s9_data_o[23] ,
    \s9_data_o[24] , \s9_data_o[25] , \s9_data_o[26] , \s9_data_o[27] ,
    \s9_data_o[28] , \s9_data_o[29] , \s9_data_o[30] , \s9_data_o[31] ,
    \s9_addr_o[0] , \s9_addr_o[1] , \s9_addr_o[2] , \s9_addr_o[3] ,
    \s9_addr_o[4] , \s9_addr_o[5] , \s9_addr_o[6] , \s9_addr_o[7] ,
    \s9_addr_o[8] , \s9_addr_o[9] , \s9_addr_o[10] , \s9_addr_o[11] ,
    \s9_addr_o[12] , \s9_addr_o[13] , \s9_addr_o[14] , \s9_addr_o[15] ,
    \s9_addr_o[16] , \s9_addr_o[17] , \s9_addr_o[18] , \s9_addr_o[19] ,
    \s9_addr_o[20] , \s9_addr_o[21] , \s9_addr_o[22] , \s9_addr_o[23] ,
    \s9_addr_o[24] , \s9_addr_o[25] , \s9_addr_o[26] , \s9_addr_o[27] ,
    \s9_addr_o[28] , \s9_addr_o[29] , \s9_addr_o[30] , \s9_addr_o[31] ,
    \s10_data_o[0] , \s10_data_o[1] , \s10_data_o[2] , \s10_data_o[3] ,
    \s10_data_o[4] , \s10_data_o[5] , \s10_data_o[6] , \s10_data_o[7] ,
    \s10_data_o[8] , \s10_data_o[9] , \s10_data_o[10] , \s10_data_o[11] ,
    \s10_data_o[12] , \s10_data_o[13] , \s10_data_o[14] , \s10_data_o[15] ,
    \s10_data_o[16] , \s10_data_o[17] , \s10_data_o[18] , \s10_data_o[19] ,
    \s10_data_o[20] , \s10_data_o[21] , \s10_data_o[22] , \s10_data_o[23] ,
    \s10_data_o[24] , \s10_data_o[25] , \s10_data_o[26] , \s10_data_o[27] ,
    \s10_data_o[28] , \s10_data_o[29] , \s10_data_o[30] , \s10_data_o[31] ,
    \s10_addr_o[0] , \s10_addr_o[1] , \s10_addr_o[2] , \s10_addr_o[3] ,
    \s10_addr_o[4] , \s10_addr_o[5] , \s10_addr_o[6] , \s10_addr_o[7] ,
    \s10_addr_o[8] , \s10_addr_o[9] , \s10_addr_o[10] , \s10_addr_o[11] ,
    \s10_addr_o[12] , \s10_addr_o[13] , \s10_addr_o[14] , \s10_addr_o[15] ,
    \s10_addr_o[16] , \s10_addr_o[17] , \s10_addr_o[18] , \s10_addr_o[19] ,
    \s10_addr_o[20] , \s10_addr_o[21] , \s10_addr_o[22] , \s10_addr_o[23] ,
    \s10_addr_o[24] , \s10_addr_o[25] , \s10_addr_o[26] , \s10_addr_o[27] ,
    \s10_addr_o[28] , \s10_addr_o[29] , \s10_addr_o[30] , \s10_addr_o[31] ,
    \s11_data_o[0] , \s11_data_o[1] , \s11_data_o[2] , \s11_data_o[3] ,
    \s11_data_o[4] , \s11_data_o[5] , \s11_data_o[6] , \s11_data_o[7] ,
    \s11_data_o[8] , \s11_data_o[9] , \s11_data_o[10] , \s11_data_o[11] ,
    \s11_data_o[12] , \s11_data_o[13] , \s11_data_o[14] , \s11_data_o[15] ,
    \s11_data_o[16] , \s11_data_o[17] , \s11_data_o[18] , \s11_data_o[19] ,
    \s11_data_o[20] , \s11_data_o[21] , \s11_data_o[22] , \s11_data_o[23] ,
    \s11_data_o[24] , \s11_data_o[25] , \s11_data_o[26] , \s11_data_o[27] ,
    \s11_data_o[28] , \s11_data_o[29] , \s11_data_o[30] , \s11_data_o[31] ,
    \s11_addr_o[0] , \s11_addr_o[1] , \s11_addr_o[2] , \s11_addr_o[3] ,
    \s11_addr_o[4] , \s11_addr_o[5] , \s11_addr_o[6] , \s11_addr_o[7] ,
    \s11_addr_o[8] , \s11_addr_o[9] , \s11_addr_o[10] , \s11_addr_o[11] ,
    \s11_addr_o[12] , \s11_addr_o[13] , \s11_addr_o[14] , \s11_addr_o[15] ,
    \s11_addr_o[16] , \s11_addr_o[17] , \s11_addr_o[18] , \s11_addr_o[19] ,
    \s11_addr_o[20] , \s11_addr_o[21] , \s11_addr_o[22] , \s11_addr_o[23] ,
    \s11_addr_o[24] , \s11_addr_o[25] , \s11_addr_o[26] , \s11_addr_o[27] ,
    \s11_addr_o[28] , \s11_addr_o[29] , \s11_addr_o[30] , \s11_addr_o[31] ,
    \s12_data_o[0] , \s12_data_o[1] , \s12_data_o[2] , \s12_data_o[3] ,
    \s12_data_o[4] , \s12_data_o[5] , \s12_data_o[6] , \s12_data_o[7] ,
    \s12_data_o[8] , \s12_data_o[9] , \s12_data_o[10] , \s12_data_o[11] ,
    \s12_data_o[12] , \s12_data_o[13] , \s12_data_o[14] , \s12_data_o[15] ,
    \s12_data_o[16] , \s12_data_o[17] , \s12_data_o[18] , \s12_data_o[19] ,
    \s12_data_o[20] , \s12_data_o[21] , \s12_data_o[22] , \s12_data_o[23] ,
    \s12_data_o[24] , \s12_data_o[25] , \s12_data_o[26] , \s12_data_o[27] ,
    \s12_data_o[28] , \s12_data_o[29] , \s12_data_o[30] , \s12_data_o[31] ,
    \s12_addr_o[0] , \s12_addr_o[1] , \s12_addr_o[2] , \s12_addr_o[3] ,
    \s12_addr_o[4] , \s12_addr_o[5] , \s12_addr_o[6] , \s12_addr_o[7] ,
    \s12_addr_o[8] , \s12_addr_o[9] , \s12_addr_o[10] , \s12_addr_o[11] ,
    \s12_addr_o[12] , \s12_addr_o[13] , \s12_addr_o[14] , \s12_addr_o[15] ,
    \s12_addr_o[16] , \s12_addr_o[17] , \s12_addr_o[18] , \s12_addr_o[19] ,
    \s12_addr_o[20] , \s12_addr_o[21] , \s12_addr_o[22] , \s12_addr_o[23] ,
    \s12_addr_o[24] , \s12_addr_o[25] , \s12_addr_o[26] , \s12_addr_o[27] ,
    \s12_addr_o[28] , \s12_addr_o[29] , \s12_addr_o[30] , \s12_addr_o[31] ,
    \s13_data_o[0] , \s13_data_o[1] , \s13_data_o[2] , \s13_data_o[3] ,
    \s13_data_o[4] , \s13_data_o[5] , \s13_data_o[6] , \s13_data_o[7] ,
    \s13_data_o[8] , \s13_data_o[9] , \s13_data_o[10] , \s13_data_o[11] ,
    \s13_data_o[12] , \s13_data_o[13] , \s13_data_o[14] , \s13_data_o[15] ,
    \s13_data_o[16] , \s13_data_o[17] , \s13_data_o[18] , \s13_data_o[19] ,
    \s13_data_o[20] , \s13_data_o[21] , \s13_data_o[22] , \s13_data_o[23] ,
    \s13_data_o[24] , \s13_data_o[25] , \s13_data_o[26] , \s13_data_o[27] ,
    \s13_data_o[28] , \s13_data_o[29] , \s13_data_o[30] , \s13_data_o[31] ,
    \s13_addr_o[0] , \s13_addr_o[1] , \s13_addr_o[2] , \s13_addr_o[3] ,
    \s13_addr_o[4] , \s13_addr_o[5] , \s13_addr_o[6] , \s13_addr_o[7] ,
    \s13_addr_o[8] , \s13_addr_o[9] , \s13_addr_o[10] , \s13_addr_o[11] ,
    \s13_addr_o[12] , \s13_addr_o[13] , \s13_addr_o[14] , \s13_addr_o[15] ,
    \s13_addr_o[16] , \s13_addr_o[17] , \s13_addr_o[18] , \s13_addr_o[19] ,
    \s13_addr_o[20] , \s13_addr_o[21] , \s13_addr_o[22] , \s13_addr_o[23] ,
    \s13_addr_o[24] , \s13_addr_o[25] , \s13_addr_o[26] , \s13_addr_o[27] ,
    \s13_addr_o[28] , \s13_addr_o[29] , \s13_addr_o[30] , \s13_addr_o[31] ,
    \s14_data_o[0] , \s14_data_o[1] , \s14_data_o[2] , \s14_data_o[3] ,
    \s14_data_o[4] , \s14_data_o[5] , \s14_data_o[6] , \s14_data_o[7] ,
    \s14_data_o[8] , \s14_data_o[9] , \s14_data_o[10] , \s14_data_o[11] ,
    \s14_data_o[12] , \s14_data_o[13] , \s14_data_o[14] , \s14_data_o[15] ,
    \s14_data_o[16] , \s14_data_o[17] , \s14_data_o[18] , \s14_data_o[19] ,
    \s14_data_o[20] , \s14_data_o[21] , \s14_data_o[22] , \s14_data_o[23] ,
    \s14_data_o[24] , \s14_data_o[25] , \s14_data_o[26] , \s14_data_o[27] ,
    \s14_data_o[28] , \s14_data_o[29] , \s14_data_o[30] , \s14_data_o[31] ,
    \s14_addr_o[0] , \s14_addr_o[1] , \s14_addr_o[2] , \s14_addr_o[3] ,
    \s14_addr_o[4] , \s14_addr_o[5] , \s14_addr_o[6] , \s14_addr_o[7] ,
    \s14_addr_o[8] , \s14_addr_o[9] , \s14_addr_o[10] , \s14_addr_o[11] ,
    \s14_addr_o[12] , \s14_addr_o[13] , \s14_addr_o[14] , \s14_addr_o[15] ,
    \s14_addr_o[16] , \s14_addr_o[17] , \s14_addr_o[18] , \s14_addr_o[19] ,
    \s14_addr_o[20] , \s14_addr_o[21] , \s14_addr_o[22] , \s14_addr_o[23] ,
    \s14_addr_o[24] , \s14_addr_o[25] , \s14_addr_o[26] , \s14_addr_o[27] ,
    \s14_addr_o[28] , \s14_addr_o[29] , \s14_addr_o[30] , \s14_addr_o[31] ,
    \s15_data_o[0] , \s15_data_o[1] , \s15_data_o[2] , \s15_data_o[3] ,
    \s15_data_o[4] , \s15_data_o[5] , \s15_data_o[6] , \s15_data_o[7] ,
    \s15_data_o[8] , \s15_data_o[9] , \s15_data_o[10] , \s15_data_o[11] ,
    \s15_data_o[12] , \s15_data_o[13] , \s15_data_o[14] , \s15_data_o[15] ,
    \s15_data_o[16] , \s15_data_o[17] , \s15_data_o[18] , \s15_data_o[19] ,
    \s15_data_o[20] , \s15_data_o[21] , \s15_data_o[22] , \s15_data_o[23] ,
    \s15_data_o[24] , \s15_data_o[25] , \s15_data_o[26] , \s15_data_o[27] ,
    \s15_data_o[28] , \s15_data_o[29] , \s15_data_o[30] , \s15_data_o[31] ,
    \s15_addr_o[0] , \s15_addr_o[1] , \s15_addr_o[2] , \s15_addr_o[3] ,
    \s15_addr_o[4] , \s15_addr_o[5] , \s15_addr_o[6] , \s15_addr_o[7] ,
    \s15_addr_o[8] , \s15_addr_o[9] , \s15_addr_o[10] , \s15_addr_o[11] ,
    \s15_addr_o[12] , \s15_addr_o[13] , \s15_addr_o[14] , \s15_addr_o[15] ,
    \s15_addr_o[16] , \s15_addr_o[17] , \s15_addr_o[18] , \s15_addr_o[19] ,
    \s15_addr_o[20] , \s15_addr_o[21] , \s15_addr_o[22] , \s15_addr_o[23] ,
    \s15_addr_o[24] , \s15_addr_o[25] , \s15_addr_o[26] , \s15_addr_o[27] ,
    \s15_addr_o[28] , \s15_addr_o[29] , \s15_addr_o[30] , \s15_addr_o[31] ,
    m0_ack_o, m0_err_o, m0_rty_o, m1_ack_o, m1_err_o, m1_rty_o, m2_ack_o,
    m2_err_o, m2_rty_o, m3_ack_o, m3_err_o, m3_rty_o, m4_ack_o, m4_err_o,
    m4_rty_o, m5_ack_o, m5_err_o, m5_rty_o, m6_ack_o, m6_err_o, m6_rty_o,
    m7_ack_o, m7_err_o, m7_rty_o, s0_we_o, s0_cyc_o, s0_stb_o, s1_we_o,
    s1_cyc_o, s1_stb_o, s2_we_o, s2_cyc_o, s2_stb_o, s3_we_o, s3_cyc_o,
    s3_stb_o, s4_we_o, s4_cyc_o, s4_stb_o, s5_we_o, s5_cyc_o, s5_stb_o,
    s6_we_o, s6_cyc_o, s6_stb_o, s7_we_o, s7_cyc_o, s7_stb_o, s8_we_o,
    s8_cyc_o, s8_stb_o, s9_we_o, s9_cyc_o, s9_stb_o, s10_we_o, s10_cyc_o,
    s10_stb_o, s11_we_o, s11_cyc_o, s11_stb_o, s12_we_o, s12_cyc_o,
    s12_stb_o, s13_we_o, s13_cyc_o, s13_stb_o, s14_we_o, s14_cyc_o,
    s14_stb_o, s15_we_o, s15_cyc_o, s15_stb_o, \s0_sel_o[0] ,
    \s0_sel_o[1] , \s0_sel_o[2] , \s0_sel_o[3] , \s1_sel_o[0] ,
    \s1_sel_o[1] , \s1_sel_o[2] , \s1_sel_o[3] , \s2_sel_o[0] ,
    \s2_sel_o[1] , \s2_sel_o[2] , \s2_sel_o[3] , \s3_sel_o[0] ,
    \s3_sel_o[1] , \s3_sel_o[2] , \s3_sel_o[3] , \s4_sel_o[0] ,
    \s4_sel_o[1] , \s4_sel_o[2] , \s4_sel_o[3] , \s5_sel_o[0] ,
    \s5_sel_o[1] , \s5_sel_o[2] , \s5_sel_o[3] , \s6_sel_o[0] ,
    \s6_sel_o[1] , \s6_sel_o[2] , \s6_sel_o[3] , \s7_sel_o[0] ,
    \s7_sel_o[1] , \s7_sel_o[2] , \s7_sel_o[3] , \s8_sel_o[0] ,
    \s8_sel_o[1] , \s8_sel_o[2] , \s8_sel_o[3] , \s9_sel_o[0] ,
    \s9_sel_o[1] , \s9_sel_o[2] , \s9_sel_o[3] , \s10_sel_o[0] ,
    \s10_sel_o[1] , \s10_sel_o[2] , \s10_sel_o[3] , \s11_sel_o[0] ,
    \s11_sel_o[1] , \s11_sel_o[2] , \s11_sel_o[3] , \s12_sel_o[0] ,
    \s12_sel_o[1] , \s12_sel_o[2] , \s12_sel_o[3] , \s13_sel_o[0] ,
    \s13_sel_o[1] , \s13_sel_o[2] , \s13_sel_o[3] , \s14_sel_o[0] ,
    \s14_sel_o[1] , \s14_sel_o[2] , \s14_sel_o[3] , \s15_sel_o[0] ,
    \s15_sel_o[1] , \s15_sel_o[2] , \s15_sel_o[3]   );
  input  clock;
  input  clk_i, rst_i, m0_we_i, m0_cyc_i, m0_stb_i, m1_we_i, m1_cyc_i,
    m1_stb_i, m2_we_i, m2_cyc_i, m2_stb_i, m3_we_i, m3_cyc_i, m3_stb_i,
    m4_we_i, m4_cyc_i, m4_stb_i, m5_we_i, m5_cyc_i, m5_stb_i, m6_we_i,
    m6_cyc_i, m6_stb_i, m7_we_i, m7_cyc_i, m7_stb_i, s0_ack_i, s0_err_i,
    s0_rty_i, s1_ack_i, s1_err_i, s1_rty_i, s2_ack_i, s2_err_i, s2_rty_i,
    s3_ack_i, s3_err_i, s3_rty_i, s4_ack_i, s4_err_i, s4_rty_i, s5_ack_i,
    s5_err_i, s5_rty_i, s6_ack_i, s6_err_i, s6_rty_i, s7_ack_i, s7_err_i,
    s7_rty_i, s8_ack_i, s8_err_i, s8_rty_i, s9_ack_i, s9_err_i, s9_rty_i,
    s10_ack_i, s10_err_i, s10_rty_i, s11_ack_i, s11_err_i, s11_rty_i,
    s12_ack_i, s12_err_i, s12_rty_i, s13_ack_i, s13_err_i, s13_rty_i,
    s14_ack_i, s14_err_i, s14_rty_i, s15_ack_i, s15_err_i, s15_rty_i,
    \m0_data_i[0] , \m0_data_i[1] , \m0_data_i[2] , \m0_data_i[3] ,
    \m0_data_i[4] , \m0_data_i[5] , \m0_data_i[6] , \m0_data_i[7] ,
    \m0_data_i[8] , \m0_data_i[9] , \m0_data_i[10] , \m0_data_i[11] ,
    \m0_data_i[12] , \m0_data_i[13] , \m0_data_i[14] , \m0_data_i[15] ,
    \m0_data_i[16] , \m0_data_i[17] , \m0_data_i[18] , \m0_data_i[19] ,
    \m0_data_i[20] , \m0_data_i[21] , \m0_data_i[22] , \m0_data_i[23] ,
    \m0_data_i[24] , \m0_data_i[25] , \m0_data_i[26] , \m0_data_i[27] ,
    \m0_data_i[28] , \m0_data_i[29] , \m0_data_i[30] , \m0_data_i[31] ,
    \m0_addr_i[0] , \m0_addr_i[1] , \m0_addr_i[2] , \m0_addr_i[3] ,
    \m0_addr_i[4] , \m0_addr_i[5] , \m0_addr_i[6] , \m0_addr_i[7] ,
    \m0_addr_i[8] , \m0_addr_i[9] , \m0_addr_i[10] , \m0_addr_i[11] ,
    \m0_addr_i[12] , \m0_addr_i[13] , \m0_addr_i[14] , \m0_addr_i[15] ,
    \m0_addr_i[16] , \m0_addr_i[17] , \m0_addr_i[18] , \m0_addr_i[19] ,
    \m0_addr_i[20] , \m0_addr_i[21] , \m0_addr_i[22] , \m0_addr_i[23] ,
    \m0_addr_i[24] , \m0_addr_i[25] , \m0_addr_i[26] , \m0_addr_i[27] ,
    \m0_addr_i[28] , \m0_addr_i[29] , \m0_addr_i[30] , \m0_addr_i[31] ,
    \m1_data_i[0] , \m1_data_i[1] , \m1_data_i[2] , \m1_data_i[3] ,
    \m1_data_i[4] , \m1_data_i[5] , \m1_data_i[6] , \m1_data_i[7] ,
    \m1_data_i[8] , \m1_data_i[9] , \m1_data_i[10] , \m1_data_i[11] ,
    \m1_data_i[12] , \m1_data_i[13] , \m1_data_i[14] , \m1_data_i[15] ,
    \m1_data_i[16] , \m1_data_i[17] , \m1_data_i[18] , \m1_data_i[19] ,
    \m1_data_i[20] , \m1_data_i[21] , \m1_data_i[22] , \m1_data_i[23] ,
    \m1_data_i[24] , \m1_data_i[25] , \m1_data_i[26] , \m1_data_i[27] ,
    \m1_data_i[28] , \m1_data_i[29] , \m1_data_i[30] , \m1_data_i[31] ,
    \m1_addr_i[0] , \m1_addr_i[1] , \m1_addr_i[2] , \m1_addr_i[3] ,
    \m1_addr_i[4] , \m1_addr_i[5] , \m1_addr_i[6] , \m1_addr_i[7] ,
    \m1_addr_i[8] , \m1_addr_i[9] , \m1_addr_i[10] , \m1_addr_i[11] ,
    \m1_addr_i[12] , \m1_addr_i[13] , \m1_addr_i[14] , \m1_addr_i[15] ,
    \m1_addr_i[16] , \m1_addr_i[17] , \m1_addr_i[18] , \m1_addr_i[19] ,
    \m1_addr_i[20] , \m1_addr_i[21] , \m1_addr_i[22] , \m1_addr_i[23] ,
    \m1_addr_i[24] , \m1_addr_i[25] , \m1_addr_i[26] , \m1_addr_i[27] ,
    \m1_addr_i[28] , \m1_addr_i[29] , \m1_addr_i[30] , \m1_addr_i[31] ,
    \m2_data_i[0] , \m2_data_i[1] , \m2_data_i[2] , \m2_data_i[3] ,
    \m2_data_i[4] , \m2_data_i[5] , \m2_data_i[6] , \m2_data_i[7] ,
    \m2_data_i[8] , \m2_data_i[9] , \m2_data_i[10] , \m2_data_i[11] ,
    \m2_data_i[12] , \m2_data_i[13] , \m2_data_i[14] , \m2_data_i[15] ,
    \m2_data_i[16] , \m2_data_i[17] , \m2_data_i[18] , \m2_data_i[19] ,
    \m2_data_i[20] , \m2_data_i[21] , \m2_data_i[22] , \m2_data_i[23] ,
    \m2_data_i[24] , \m2_data_i[25] , \m2_data_i[26] , \m2_data_i[27] ,
    \m2_data_i[28] , \m2_data_i[29] , \m2_data_i[30] , \m2_data_i[31] ,
    \m2_addr_i[0] , \m2_addr_i[1] , \m2_addr_i[2] , \m2_addr_i[3] ,
    \m2_addr_i[4] , \m2_addr_i[5] , \m2_addr_i[6] , \m2_addr_i[7] ,
    \m2_addr_i[8] , \m2_addr_i[9] , \m2_addr_i[10] , \m2_addr_i[11] ,
    \m2_addr_i[12] , \m2_addr_i[13] , \m2_addr_i[14] , \m2_addr_i[15] ,
    \m2_addr_i[16] , \m2_addr_i[17] , \m2_addr_i[18] , \m2_addr_i[19] ,
    \m2_addr_i[20] , \m2_addr_i[21] , \m2_addr_i[22] , \m2_addr_i[23] ,
    \m2_addr_i[24] , \m2_addr_i[25] , \m2_addr_i[26] , \m2_addr_i[27] ,
    \m2_addr_i[28] , \m2_addr_i[29] , \m2_addr_i[30] , \m2_addr_i[31] ,
    \m3_data_i[0] , \m3_data_i[1] , \m3_data_i[2] , \m3_data_i[3] ,
    \m3_data_i[4] , \m3_data_i[5] , \m3_data_i[6] , \m3_data_i[7] ,
    \m3_data_i[8] , \m3_data_i[9] , \m3_data_i[10] , \m3_data_i[11] ,
    \m3_data_i[12] , \m3_data_i[13] , \m3_data_i[14] , \m3_data_i[15] ,
    \m3_data_i[16] , \m3_data_i[17] , \m3_data_i[18] , \m3_data_i[19] ,
    \m3_data_i[20] , \m3_data_i[21] , \m3_data_i[22] , \m3_data_i[23] ,
    \m3_data_i[24] , \m3_data_i[25] , \m3_data_i[26] , \m3_data_i[27] ,
    \m3_data_i[28] , \m3_data_i[29] , \m3_data_i[30] , \m3_data_i[31] ,
    \m3_addr_i[0] , \m3_addr_i[1] , \m3_addr_i[2] , \m3_addr_i[3] ,
    \m3_addr_i[4] , \m3_addr_i[5] , \m3_addr_i[6] , \m3_addr_i[7] ,
    \m3_addr_i[8] , \m3_addr_i[9] , \m3_addr_i[10] , \m3_addr_i[11] ,
    \m3_addr_i[12] , \m3_addr_i[13] , \m3_addr_i[14] , \m3_addr_i[15] ,
    \m3_addr_i[16] , \m3_addr_i[17] , \m3_addr_i[18] , \m3_addr_i[19] ,
    \m3_addr_i[20] , \m3_addr_i[21] , \m3_addr_i[22] , \m3_addr_i[23] ,
    \m3_addr_i[24] , \m3_addr_i[25] , \m3_addr_i[26] , \m3_addr_i[27] ,
    \m3_addr_i[28] , \m3_addr_i[29] , \m3_addr_i[30] , \m3_addr_i[31] ,
    \m4_data_i[0] , \m4_data_i[1] , \m4_data_i[2] , \m4_data_i[3] ,
    \m4_data_i[4] , \m4_data_i[5] , \m4_data_i[6] , \m4_data_i[7] ,
    \m4_data_i[8] , \m4_data_i[9] , \m4_data_i[10] , \m4_data_i[11] ,
    \m4_data_i[12] , \m4_data_i[13] , \m4_data_i[14] , \m4_data_i[15] ,
    \m4_data_i[16] , \m4_data_i[17] , \m4_data_i[18] , \m4_data_i[19] ,
    \m4_data_i[20] , \m4_data_i[21] , \m4_data_i[22] , \m4_data_i[23] ,
    \m4_data_i[24] , \m4_data_i[25] , \m4_data_i[26] , \m4_data_i[27] ,
    \m4_data_i[28] , \m4_data_i[29] , \m4_data_i[30] , \m4_data_i[31] ,
    \m4_addr_i[0] , \m4_addr_i[1] , \m4_addr_i[2] , \m4_addr_i[3] ,
    \m4_addr_i[4] , \m4_addr_i[5] , \m4_addr_i[6] , \m4_addr_i[7] ,
    \m4_addr_i[8] , \m4_addr_i[9] , \m4_addr_i[10] , \m4_addr_i[11] ,
    \m4_addr_i[12] , \m4_addr_i[13] , \m4_addr_i[14] , \m4_addr_i[15] ,
    \m4_addr_i[16] , \m4_addr_i[17] , \m4_addr_i[18] , \m4_addr_i[19] ,
    \m4_addr_i[20] , \m4_addr_i[21] , \m4_addr_i[22] , \m4_addr_i[23] ,
    \m4_addr_i[24] , \m4_addr_i[25] , \m4_addr_i[26] , \m4_addr_i[27] ,
    \m4_addr_i[28] , \m4_addr_i[29] , \m4_addr_i[30] , \m4_addr_i[31] ,
    \m5_data_i[0] , \m5_data_i[1] , \m5_data_i[2] , \m5_data_i[3] ,
    \m5_data_i[4] , \m5_data_i[5] , \m5_data_i[6] , \m5_data_i[7] ,
    \m5_data_i[8] , \m5_data_i[9] , \m5_data_i[10] , \m5_data_i[11] ,
    \m5_data_i[12] , \m5_data_i[13] , \m5_data_i[14] , \m5_data_i[15] ,
    \m5_data_i[16] , \m5_data_i[17] , \m5_data_i[18] , \m5_data_i[19] ,
    \m5_data_i[20] , \m5_data_i[21] , \m5_data_i[22] , \m5_data_i[23] ,
    \m5_data_i[24] , \m5_data_i[25] , \m5_data_i[26] , \m5_data_i[27] ,
    \m5_data_i[28] , \m5_data_i[29] , \m5_data_i[30] , \m5_data_i[31] ,
    \m5_addr_i[0] , \m5_addr_i[1] , \m5_addr_i[2] , \m5_addr_i[3] ,
    \m5_addr_i[4] , \m5_addr_i[5] , \m5_addr_i[6] , \m5_addr_i[7] ,
    \m5_addr_i[8] , \m5_addr_i[9] , \m5_addr_i[10] , \m5_addr_i[11] ,
    \m5_addr_i[12] , \m5_addr_i[13] , \m5_addr_i[14] , \m5_addr_i[15] ,
    \m5_addr_i[16] , \m5_addr_i[17] , \m5_addr_i[18] , \m5_addr_i[19] ,
    \m5_addr_i[20] , \m5_addr_i[21] , \m5_addr_i[22] , \m5_addr_i[23] ,
    \m5_addr_i[24] , \m5_addr_i[25] , \m5_addr_i[26] , \m5_addr_i[27] ,
    \m5_addr_i[28] , \m5_addr_i[29] , \m5_addr_i[30] , \m5_addr_i[31] ,
    \m6_data_i[0] , \m6_data_i[1] , \m6_data_i[2] , \m6_data_i[3] ,
    \m6_data_i[4] , \m6_data_i[5] , \m6_data_i[6] , \m6_data_i[7] ,
    \m6_data_i[8] , \m6_data_i[9] , \m6_data_i[10] , \m6_data_i[11] ,
    \m6_data_i[12] , \m6_data_i[13] , \m6_data_i[14] , \m6_data_i[15] ,
    \m6_data_i[16] , \m6_data_i[17] , \m6_data_i[18] , \m6_data_i[19] ,
    \m6_data_i[20] , \m6_data_i[21] , \m6_data_i[22] , \m6_data_i[23] ,
    \m6_data_i[24] , \m6_data_i[25] , \m6_data_i[26] , \m6_data_i[27] ,
    \m6_data_i[28] , \m6_data_i[29] , \m6_data_i[30] , \m6_data_i[31] ,
    \m6_addr_i[0] , \m6_addr_i[1] , \m6_addr_i[2] , \m6_addr_i[3] ,
    \m6_addr_i[4] , \m6_addr_i[5] , \m6_addr_i[6] , \m6_addr_i[7] ,
    \m6_addr_i[8] , \m6_addr_i[9] , \m6_addr_i[10] , \m6_addr_i[11] ,
    \m6_addr_i[12] , \m6_addr_i[13] , \m6_addr_i[14] , \m6_addr_i[15] ,
    \m6_addr_i[16] , \m6_addr_i[17] , \m6_addr_i[18] , \m6_addr_i[19] ,
    \m6_addr_i[20] , \m6_addr_i[21] , \m6_addr_i[22] , \m6_addr_i[23] ,
    \m6_addr_i[24] , \m6_addr_i[25] , \m6_addr_i[26] , \m6_addr_i[27] ,
    \m6_addr_i[28] , \m6_addr_i[29] , \m6_addr_i[30] , \m6_addr_i[31] ,
    \m7_data_i[0] , \m7_data_i[1] , \m7_data_i[2] , \m7_data_i[3] ,
    \m7_data_i[4] , \m7_data_i[5] , \m7_data_i[6] , \m7_data_i[7] ,
    \m7_data_i[8] , \m7_data_i[9] , \m7_data_i[10] , \m7_data_i[11] ,
    \m7_data_i[12] , \m7_data_i[13] , \m7_data_i[14] , \m7_data_i[15] ,
    \m7_data_i[16] , \m7_data_i[17] , \m7_data_i[18] , \m7_data_i[19] ,
    \m7_data_i[20] , \m7_data_i[21] , \m7_data_i[22] , \m7_data_i[23] ,
    \m7_data_i[24] , \m7_data_i[25] , \m7_data_i[26] , \m7_data_i[27] ,
    \m7_data_i[28] , \m7_data_i[29] , \m7_data_i[30] , \m7_data_i[31] ,
    \m7_addr_i[0] , \m7_addr_i[1] , \m7_addr_i[2] , \m7_addr_i[3] ,
    \m7_addr_i[4] , \m7_addr_i[5] , \m7_addr_i[6] , \m7_addr_i[7] ,
    \m7_addr_i[8] , \m7_addr_i[9] , \m7_addr_i[10] , \m7_addr_i[11] ,
    \m7_addr_i[12] , \m7_addr_i[13] , \m7_addr_i[14] , \m7_addr_i[15] ,
    \m7_addr_i[16] , \m7_addr_i[17] , \m7_addr_i[18] , \m7_addr_i[19] ,
    \m7_addr_i[20] , \m7_addr_i[21] , \m7_addr_i[22] , \m7_addr_i[23] ,
    \m7_addr_i[24] , \m7_addr_i[25] , \m7_addr_i[26] , \m7_addr_i[27] ,
    \m7_addr_i[28] , \m7_addr_i[29] , \m7_addr_i[30] , \m7_addr_i[31] ,
    \s0_data_i[0] , \s0_data_i[1] , \s0_data_i[2] , \s0_data_i[3] ,
    \s0_data_i[4] , \s0_data_i[5] , \s0_data_i[6] , \s0_data_i[7] ,
    \s0_data_i[8] , \s0_data_i[9] , \s0_data_i[10] , \s0_data_i[11] ,
    \s0_data_i[12] , \s0_data_i[13] , \s0_data_i[14] , \s0_data_i[15] ,
    \s0_data_i[16] , \s0_data_i[17] , \s0_data_i[18] , \s0_data_i[19] ,
    \s0_data_i[20] , \s0_data_i[21] , \s0_data_i[22] , \s0_data_i[23] ,
    \s0_data_i[24] , \s0_data_i[25] , \s0_data_i[26] , \s0_data_i[27] ,
    \s0_data_i[28] , \s0_data_i[29] , \s0_data_i[30] , \s0_data_i[31] ,
    \s1_data_i[0] , \s1_data_i[1] , \s1_data_i[2] , \s1_data_i[3] ,
    \s1_data_i[4] , \s1_data_i[5] , \s1_data_i[6] , \s1_data_i[7] ,
    \s1_data_i[8] , \s1_data_i[9] , \s1_data_i[10] , \s1_data_i[11] ,
    \s1_data_i[12] , \s1_data_i[13] , \s1_data_i[14] , \s1_data_i[15] ,
    \s1_data_i[16] , \s1_data_i[17] , \s1_data_i[18] , \s1_data_i[19] ,
    \s1_data_i[20] , \s1_data_i[21] , \s1_data_i[22] , \s1_data_i[23] ,
    \s1_data_i[24] , \s1_data_i[25] , \s1_data_i[26] , \s1_data_i[27] ,
    \s1_data_i[28] , \s1_data_i[29] , \s1_data_i[30] , \s1_data_i[31] ,
    \s2_data_i[0] , \s2_data_i[1] , \s2_data_i[2] , \s2_data_i[3] ,
    \s2_data_i[4] , \s2_data_i[5] , \s2_data_i[6] , \s2_data_i[7] ,
    \s2_data_i[8] , \s2_data_i[9] , \s2_data_i[10] , \s2_data_i[11] ,
    \s2_data_i[12] , \s2_data_i[13] , \s2_data_i[14] , \s2_data_i[15] ,
    \s2_data_i[16] , \s2_data_i[17] , \s2_data_i[18] , \s2_data_i[19] ,
    \s2_data_i[20] , \s2_data_i[21] , \s2_data_i[22] , \s2_data_i[23] ,
    \s2_data_i[24] , \s2_data_i[25] , \s2_data_i[26] , \s2_data_i[27] ,
    \s2_data_i[28] , \s2_data_i[29] , \s2_data_i[30] , \s2_data_i[31] ,
    \s3_data_i[0] , \s3_data_i[1] , \s3_data_i[2] , \s3_data_i[3] ,
    \s3_data_i[4] , \s3_data_i[5] , \s3_data_i[6] , \s3_data_i[7] ,
    \s3_data_i[8] , \s3_data_i[9] , \s3_data_i[10] , \s3_data_i[11] ,
    \s3_data_i[12] , \s3_data_i[13] , \s3_data_i[14] , \s3_data_i[15] ,
    \s3_data_i[16] , \s3_data_i[17] , \s3_data_i[18] , \s3_data_i[19] ,
    \s3_data_i[20] , \s3_data_i[21] , \s3_data_i[22] , \s3_data_i[23] ,
    \s3_data_i[24] , \s3_data_i[25] , \s3_data_i[26] , \s3_data_i[27] ,
    \s3_data_i[28] , \s3_data_i[29] , \s3_data_i[30] , \s3_data_i[31] ,
    \s4_data_i[0] , \s4_data_i[1] , \s4_data_i[2] , \s4_data_i[3] ,
    \s4_data_i[4] , \s4_data_i[5] , \s4_data_i[6] , \s4_data_i[7] ,
    \s4_data_i[8] , \s4_data_i[9] , \s4_data_i[10] , \s4_data_i[11] ,
    \s4_data_i[12] , \s4_data_i[13] , \s4_data_i[14] , \s4_data_i[15] ,
    \s4_data_i[16] , \s4_data_i[17] , \s4_data_i[18] , \s4_data_i[19] ,
    \s4_data_i[20] , \s4_data_i[21] , \s4_data_i[22] , \s4_data_i[23] ,
    \s4_data_i[24] , \s4_data_i[25] , \s4_data_i[26] , \s4_data_i[27] ,
    \s4_data_i[28] , \s4_data_i[29] , \s4_data_i[30] , \s4_data_i[31] ,
    \s5_data_i[0] , \s5_data_i[1] , \s5_data_i[2] , \s5_data_i[3] ,
    \s5_data_i[4] , \s5_data_i[5] , \s5_data_i[6] , \s5_data_i[7] ,
    \s5_data_i[8] , \s5_data_i[9] , \s5_data_i[10] , \s5_data_i[11] ,
    \s5_data_i[12] , \s5_data_i[13] , \s5_data_i[14] , \s5_data_i[15] ,
    \s5_data_i[16] , \s5_data_i[17] , \s5_data_i[18] , \s5_data_i[19] ,
    \s5_data_i[20] , \s5_data_i[21] , \s5_data_i[22] , \s5_data_i[23] ,
    \s5_data_i[24] , \s5_data_i[25] , \s5_data_i[26] , \s5_data_i[27] ,
    \s5_data_i[28] , \s5_data_i[29] , \s5_data_i[30] , \s5_data_i[31] ,
    \s6_data_i[0] , \s6_data_i[1] , \s6_data_i[2] , \s6_data_i[3] ,
    \s6_data_i[4] , \s6_data_i[5] , \s6_data_i[6] , \s6_data_i[7] ,
    \s6_data_i[8] , \s6_data_i[9] , \s6_data_i[10] , \s6_data_i[11] ,
    \s6_data_i[12] , \s6_data_i[13] , \s6_data_i[14] , \s6_data_i[15] ,
    \s6_data_i[16] , \s6_data_i[17] , \s6_data_i[18] , \s6_data_i[19] ,
    \s6_data_i[20] , \s6_data_i[21] , \s6_data_i[22] , \s6_data_i[23] ,
    \s6_data_i[24] , \s6_data_i[25] , \s6_data_i[26] , \s6_data_i[27] ,
    \s6_data_i[28] , \s6_data_i[29] , \s6_data_i[30] , \s6_data_i[31] ,
    \s7_data_i[0] , \s7_data_i[1] , \s7_data_i[2] , \s7_data_i[3] ,
    \s7_data_i[4] , \s7_data_i[5] , \s7_data_i[6] , \s7_data_i[7] ,
    \s7_data_i[8] , \s7_data_i[9] , \s7_data_i[10] , \s7_data_i[11] ,
    \s7_data_i[12] , \s7_data_i[13] , \s7_data_i[14] , \s7_data_i[15] ,
    \s7_data_i[16] , \s7_data_i[17] , \s7_data_i[18] , \s7_data_i[19] ,
    \s7_data_i[20] , \s7_data_i[21] , \s7_data_i[22] , \s7_data_i[23] ,
    \s7_data_i[24] , \s7_data_i[25] , \s7_data_i[26] , \s7_data_i[27] ,
    \s7_data_i[28] , \s7_data_i[29] , \s7_data_i[30] , \s7_data_i[31] ,
    \s8_data_i[0] , \s8_data_i[1] , \s8_data_i[2] , \s8_data_i[3] ,
    \s8_data_i[4] , \s8_data_i[5] , \s8_data_i[6] , \s8_data_i[7] ,
    \s8_data_i[8] , \s8_data_i[9] , \s8_data_i[10] , \s8_data_i[11] ,
    \s8_data_i[12] , \s8_data_i[13] , \s8_data_i[14] , \s8_data_i[15] ,
    \s8_data_i[16] , \s8_data_i[17] , \s8_data_i[18] , \s8_data_i[19] ,
    \s8_data_i[20] , \s8_data_i[21] , \s8_data_i[22] , \s8_data_i[23] ,
    \s8_data_i[24] , \s8_data_i[25] , \s8_data_i[26] , \s8_data_i[27] ,
    \s8_data_i[28] , \s8_data_i[29] , \s8_data_i[30] , \s8_data_i[31] ,
    \s9_data_i[0] , \s9_data_i[1] , \s9_data_i[2] , \s9_data_i[3] ,
    \s9_data_i[4] , \s9_data_i[5] , \s9_data_i[6] , \s9_data_i[7] ,
    \s9_data_i[8] , \s9_data_i[9] , \s9_data_i[10] , \s9_data_i[11] ,
    \s9_data_i[12] , \s9_data_i[13] , \s9_data_i[14] , \s9_data_i[15] ,
    \s9_data_i[16] , \s9_data_i[17] , \s9_data_i[18] , \s9_data_i[19] ,
    \s9_data_i[20] , \s9_data_i[21] , \s9_data_i[22] , \s9_data_i[23] ,
    \s9_data_i[24] , \s9_data_i[25] , \s9_data_i[26] , \s9_data_i[27] ,
    \s9_data_i[28] , \s9_data_i[29] , \s9_data_i[30] , \s9_data_i[31] ,
    \s10_data_i[0] , \s10_data_i[1] , \s10_data_i[2] , \s10_data_i[3] ,
    \s10_data_i[4] , \s10_data_i[5] , \s10_data_i[6] , \s10_data_i[7] ,
    \s10_data_i[8] , \s10_data_i[9] , \s10_data_i[10] , \s10_data_i[11] ,
    \s10_data_i[12] , \s10_data_i[13] , \s10_data_i[14] , \s10_data_i[15] ,
    \s10_data_i[16] , \s10_data_i[17] , \s10_data_i[18] , \s10_data_i[19] ,
    \s10_data_i[20] , \s10_data_i[21] , \s10_data_i[22] , \s10_data_i[23] ,
    \s10_data_i[24] , \s10_data_i[25] , \s10_data_i[26] , \s10_data_i[27] ,
    \s10_data_i[28] , \s10_data_i[29] , \s10_data_i[30] , \s10_data_i[31] ,
    \s11_data_i[0] , \s11_data_i[1] , \s11_data_i[2] , \s11_data_i[3] ,
    \s11_data_i[4] , \s11_data_i[5] , \s11_data_i[6] , \s11_data_i[7] ,
    \s11_data_i[8] , \s11_data_i[9] , \s11_data_i[10] , \s11_data_i[11] ,
    \s11_data_i[12] , \s11_data_i[13] , \s11_data_i[14] , \s11_data_i[15] ,
    \s11_data_i[16] , \s11_data_i[17] , \s11_data_i[18] , \s11_data_i[19] ,
    \s11_data_i[20] , \s11_data_i[21] , \s11_data_i[22] , \s11_data_i[23] ,
    \s11_data_i[24] , \s11_data_i[25] , \s11_data_i[26] , \s11_data_i[27] ,
    \s11_data_i[28] , \s11_data_i[29] , \s11_data_i[30] , \s11_data_i[31] ,
    \s12_data_i[0] , \s12_data_i[1] , \s12_data_i[2] , \s12_data_i[3] ,
    \s12_data_i[4] , \s12_data_i[5] , \s12_data_i[6] , \s12_data_i[7] ,
    \s12_data_i[8] , \s12_data_i[9] , \s12_data_i[10] , \s12_data_i[11] ,
    \s12_data_i[12] , \s12_data_i[13] , \s12_data_i[14] , \s12_data_i[15] ,
    \s12_data_i[16] , \s12_data_i[17] , \s12_data_i[18] , \s12_data_i[19] ,
    \s12_data_i[20] , \s12_data_i[21] , \s12_data_i[22] , \s12_data_i[23] ,
    \s12_data_i[24] , \s12_data_i[25] , \s12_data_i[26] , \s12_data_i[27] ,
    \s12_data_i[28] , \s12_data_i[29] , \s12_data_i[30] , \s12_data_i[31] ,
    \s13_data_i[0] , \s13_data_i[1] , \s13_data_i[2] , \s13_data_i[3] ,
    \s13_data_i[4] , \s13_data_i[5] , \s13_data_i[6] , \s13_data_i[7] ,
    \s13_data_i[8] , \s13_data_i[9] , \s13_data_i[10] , \s13_data_i[11] ,
    \s13_data_i[12] , \s13_data_i[13] , \s13_data_i[14] , \s13_data_i[15] ,
    \s13_data_i[16] , \s13_data_i[17] , \s13_data_i[18] , \s13_data_i[19] ,
    \s13_data_i[20] , \s13_data_i[21] , \s13_data_i[22] , \s13_data_i[23] ,
    \s13_data_i[24] , \s13_data_i[25] , \s13_data_i[26] , \s13_data_i[27] ,
    \s13_data_i[28] , \s13_data_i[29] , \s13_data_i[30] , \s13_data_i[31] ,
    \s14_data_i[0] , \s14_data_i[1] , \s14_data_i[2] , \s14_data_i[3] ,
    \s14_data_i[4] , \s14_data_i[5] , \s14_data_i[6] , \s14_data_i[7] ,
    \s14_data_i[8] , \s14_data_i[9] , \s14_data_i[10] , \s14_data_i[11] ,
    \s14_data_i[12] , \s14_data_i[13] , \s14_data_i[14] , \s14_data_i[15] ,
    \s14_data_i[16] , \s14_data_i[17] , \s14_data_i[18] , \s14_data_i[19] ,
    \s14_data_i[20] , \s14_data_i[21] , \s14_data_i[22] , \s14_data_i[23] ,
    \s14_data_i[24] , \s14_data_i[25] , \s14_data_i[26] , \s14_data_i[27] ,
    \s14_data_i[28] , \s14_data_i[29] , \s14_data_i[30] , \s14_data_i[31] ,
    \s15_data_i[0] , \s15_data_i[1] , \s15_data_i[2] , \s15_data_i[3] ,
    \s15_data_i[4] , \s15_data_i[5] , \s15_data_i[6] , \s15_data_i[7] ,
    \s15_data_i[8] , \s15_data_i[9] , \s15_data_i[10] , \s15_data_i[11] ,
    \s15_data_i[12] , \s15_data_i[13] , \s15_data_i[14] , \s15_data_i[15] ,
    \s15_data_i[16] , \s15_data_i[17] , \s15_data_i[18] , \s15_data_i[19] ,
    \s15_data_i[20] , \s15_data_i[21] , \s15_data_i[22] , \s15_data_i[23] ,
    \s15_data_i[24] , \s15_data_i[25] , \s15_data_i[26] , \s15_data_i[27] ,
    \s15_data_i[28] , \s15_data_i[29] , \s15_data_i[30] , \s15_data_i[31] ,
    \m0_sel_i[0] , \m0_sel_i[1] , \m0_sel_i[2] , \m0_sel_i[3] ,
    \m1_sel_i[0] , \m1_sel_i[1] , \m1_sel_i[2] , \m1_sel_i[3] ,
    \m2_sel_i[0] , \m2_sel_i[1] , \m2_sel_i[2] , \m2_sel_i[3] ,
    \m3_sel_i[0] , \m3_sel_i[1] , \m3_sel_i[2] , \m3_sel_i[3] ,
    \m4_sel_i[0] , \m4_sel_i[1] , \m4_sel_i[2] , \m4_sel_i[3] ,
    \m5_sel_i[0] , \m5_sel_i[1] , \m5_sel_i[2] , \m5_sel_i[3] ,
    \m6_sel_i[0] , \m6_sel_i[1] , \m6_sel_i[2] , \m6_sel_i[3] ,
    \m7_sel_i[0] , \m7_sel_i[1] , \m7_sel_i[2] , \m7_sel_i[3] ;
  output \m0_data_o[0] , \m0_data_o[1] , \m0_data_o[2] , \m0_data_o[3] ,
    \m0_data_o[4] , \m0_data_o[5] , \m0_data_o[6] , \m0_data_o[7] ,
    \m0_data_o[8] , \m0_data_o[9] , \m0_data_o[10] , \m0_data_o[11] ,
    \m0_data_o[12] , \m0_data_o[13] , \m0_data_o[14] , \m0_data_o[15] ,
    \m0_data_o[16] , \m0_data_o[17] , \m0_data_o[18] , \m0_data_o[19] ,
    \m0_data_o[20] , \m0_data_o[21] , \m0_data_o[22] , \m0_data_o[23] ,
    \m0_data_o[24] , \m0_data_o[25] , \m0_data_o[26] , \m0_data_o[27] ,
    \m0_data_o[28] , \m0_data_o[29] , \m0_data_o[30] , \m0_data_o[31] ,
    \m1_data_o[0] , \m1_data_o[1] , \m1_data_o[2] , \m1_data_o[3] ,
    \m1_data_o[4] , \m1_data_o[5] , \m1_data_o[6] , \m1_data_o[7] ,
    \m1_data_o[8] , \m1_data_o[9] , \m1_data_o[10] , \m1_data_o[11] ,
    \m1_data_o[12] , \m1_data_o[13] , \m1_data_o[14] , \m1_data_o[15] ,
    \m1_data_o[16] , \m1_data_o[17] , \m1_data_o[18] , \m1_data_o[19] ,
    \m1_data_o[20] , \m1_data_o[21] , \m1_data_o[22] , \m1_data_o[23] ,
    \m1_data_o[24] , \m1_data_o[25] , \m1_data_o[26] , \m1_data_o[27] ,
    \m1_data_o[28] , \m1_data_o[29] , \m1_data_o[30] , \m1_data_o[31] ,
    \m2_data_o[0] , \m2_data_o[1] , \m2_data_o[2] , \m2_data_o[3] ,
    \m2_data_o[4] , \m2_data_o[5] , \m2_data_o[6] , \m2_data_o[7] ,
    \m2_data_o[8] , \m2_data_o[9] , \m2_data_o[10] , \m2_data_o[11] ,
    \m2_data_o[12] , \m2_data_o[13] , \m2_data_o[14] , \m2_data_o[15] ,
    \m2_data_o[16] , \m2_data_o[17] , \m2_data_o[18] , \m2_data_o[19] ,
    \m2_data_o[20] , \m2_data_o[21] , \m2_data_o[22] , \m2_data_o[23] ,
    \m2_data_o[24] , \m2_data_o[25] , \m2_data_o[26] , \m2_data_o[27] ,
    \m2_data_o[28] , \m2_data_o[29] , \m2_data_o[30] , \m2_data_o[31] ,
    \m3_data_o[0] , \m3_data_o[1] , \m3_data_o[2] , \m3_data_o[3] ,
    \m3_data_o[4] , \m3_data_o[5] , \m3_data_o[6] , \m3_data_o[7] ,
    \m3_data_o[8] , \m3_data_o[9] , \m3_data_o[10] , \m3_data_o[11] ,
    \m3_data_o[12] , \m3_data_o[13] , \m3_data_o[14] , \m3_data_o[15] ,
    \m3_data_o[16] , \m3_data_o[17] , \m3_data_o[18] , \m3_data_o[19] ,
    \m3_data_o[20] , \m3_data_o[21] , \m3_data_o[22] , \m3_data_o[23] ,
    \m3_data_o[24] , \m3_data_o[25] , \m3_data_o[26] , \m3_data_o[27] ,
    \m3_data_o[28] , \m3_data_o[29] , \m3_data_o[30] , \m3_data_o[31] ,
    \m4_data_o[0] , \m4_data_o[1] , \m4_data_o[2] , \m4_data_o[3] ,
    \m4_data_o[4] , \m4_data_o[5] , \m4_data_o[6] , \m4_data_o[7] ,
    \m4_data_o[8] , \m4_data_o[9] , \m4_data_o[10] , \m4_data_o[11] ,
    \m4_data_o[12] , \m4_data_o[13] , \m4_data_o[14] , \m4_data_o[15] ,
    \m4_data_o[16] , \m4_data_o[17] , \m4_data_o[18] , \m4_data_o[19] ,
    \m4_data_o[20] , \m4_data_o[21] , \m4_data_o[22] , \m4_data_o[23] ,
    \m4_data_o[24] , \m4_data_o[25] , \m4_data_o[26] , \m4_data_o[27] ,
    \m4_data_o[28] , \m4_data_o[29] , \m4_data_o[30] , \m4_data_o[31] ,
    \m5_data_o[0] , \m5_data_o[1] , \m5_data_o[2] , \m5_data_o[3] ,
    \m5_data_o[4] , \m5_data_o[5] , \m5_data_o[6] , \m5_data_o[7] ,
    \m5_data_o[8] , \m5_data_o[9] , \m5_data_o[10] , \m5_data_o[11] ,
    \m5_data_o[12] , \m5_data_o[13] , \m5_data_o[14] , \m5_data_o[15] ,
    \m5_data_o[16] , \m5_data_o[17] , \m5_data_o[18] , \m5_data_o[19] ,
    \m5_data_o[20] , \m5_data_o[21] , \m5_data_o[22] , \m5_data_o[23] ,
    \m5_data_o[24] , \m5_data_o[25] , \m5_data_o[26] , \m5_data_o[27] ,
    \m5_data_o[28] , \m5_data_o[29] , \m5_data_o[30] , \m5_data_o[31] ,
    \m6_data_o[0] , \m6_data_o[1] , \m6_data_o[2] , \m6_data_o[3] ,
    \m6_data_o[4] , \m6_data_o[5] , \m6_data_o[6] , \m6_data_o[7] ,
    \m6_data_o[8] , \m6_data_o[9] , \m6_data_o[10] , \m6_data_o[11] ,
    \m6_data_o[12] , \m6_data_o[13] , \m6_data_o[14] , \m6_data_o[15] ,
    \m6_data_o[16] , \m6_data_o[17] , \m6_data_o[18] , \m6_data_o[19] ,
    \m6_data_o[20] , \m6_data_o[21] , \m6_data_o[22] , \m6_data_o[23] ,
    \m6_data_o[24] , \m6_data_o[25] , \m6_data_o[26] , \m6_data_o[27] ,
    \m6_data_o[28] , \m6_data_o[29] , \m6_data_o[30] , \m6_data_o[31] ,
    \m7_data_o[0] , \m7_data_o[1] , \m7_data_o[2] , \m7_data_o[3] ,
    \m7_data_o[4] , \m7_data_o[5] , \m7_data_o[6] , \m7_data_o[7] ,
    \m7_data_o[8] , \m7_data_o[9] , \m7_data_o[10] , \m7_data_o[11] ,
    \m7_data_o[12] , \m7_data_o[13] , \m7_data_o[14] , \m7_data_o[15] ,
    \m7_data_o[16] , \m7_data_o[17] , \m7_data_o[18] , \m7_data_o[19] ,
    \m7_data_o[20] , \m7_data_o[21] , \m7_data_o[22] , \m7_data_o[23] ,
    \m7_data_o[24] , \m7_data_o[25] , \m7_data_o[26] , \m7_data_o[27] ,
    \m7_data_o[28] , \m7_data_o[29] , \m7_data_o[30] , \m7_data_o[31] ,
    \s0_data_o[0] , \s0_data_o[1] , \s0_data_o[2] , \s0_data_o[3] ,
    \s0_data_o[4] , \s0_data_o[5] , \s0_data_o[6] , \s0_data_o[7] ,
    \s0_data_o[8] , \s0_data_o[9] , \s0_data_o[10] , \s0_data_o[11] ,
    \s0_data_o[12] , \s0_data_o[13] , \s0_data_o[14] , \s0_data_o[15] ,
    \s0_data_o[16] , \s0_data_o[17] , \s0_data_o[18] , \s0_data_o[19] ,
    \s0_data_o[20] , \s0_data_o[21] , \s0_data_o[22] , \s0_data_o[23] ,
    \s0_data_o[24] , \s0_data_o[25] , \s0_data_o[26] , \s0_data_o[27] ,
    \s0_data_o[28] , \s0_data_o[29] , \s0_data_o[30] , \s0_data_o[31] ,
    \s0_addr_o[0] , \s0_addr_o[1] , \s0_addr_o[2] , \s0_addr_o[3] ,
    \s0_addr_o[4] , \s0_addr_o[5] , \s0_addr_o[6] , \s0_addr_o[7] ,
    \s0_addr_o[8] , \s0_addr_o[9] , \s0_addr_o[10] , \s0_addr_o[11] ,
    \s0_addr_o[12] , \s0_addr_o[13] , \s0_addr_o[14] , \s0_addr_o[15] ,
    \s0_addr_o[16] , \s0_addr_o[17] , \s0_addr_o[18] , \s0_addr_o[19] ,
    \s0_addr_o[20] , \s0_addr_o[21] , \s0_addr_o[22] , \s0_addr_o[23] ,
    \s0_addr_o[24] , \s0_addr_o[25] , \s0_addr_o[26] , \s0_addr_o[27] ,
    \s0_addr_o[28] , \s0_addr_o[29] , \s0_addr_o[30] , \s0_addr_o[31] ,
    \s1_data_o[0] , \s1_data_o[1] , \s1_data_o[2] , \s1_data_o[3] ,
    \s1_data_o[4] , \s1_data_o[5] , \s1_data_o[6] , \s1_data_o[7] ,
    \s1_data_o[8] , \s1_data_o[9] , \s1_data_o[10] , \s1_data_o[11] ,
    \s1_data_o[12] , \s1_data_o[13] , \s1_data_o[14] , \s1_data_o[15] ,
    \s1_data_o[16] , \s1_data_o[17] , \s1_data_o[18] , \s1_data_o[19] ,
    \s1_data_o[20] , \s1_data_o[21] , \s1_data_o[22] , \s1_data_o[23] ,
    \s1_data_o[24] , \s1_data_o[25] , \s1_data_o[26] , \s1_data_o[27] ,
    \s1_data_o[28] , \s1_data_o[29] , \s1_data_o[30] , \s1_data_o[31] ,
    \s1_addr_o[0] , \s1_addr_o[1] , \s1_addr_o[2] , \s1_addr_o[3] ,
    \s1_addr_o[4] , \s1_addr_o[5] , \s1_addr_o[6] , \s1_addr_o[7] ,
    \s1_addr_o[8] , \s1_addr_o[9] , \s1_addr_o[10] , \s1_addr_o[11] ,
    \s1_addr_o[12] , \s1_addr_o[13] , \s1_addr_o[14] , \s1_addr_o[15] ,
    \s1_addr_o[16] , \s1_addr_o[17] , \s1_addr_o[18] , \s1_addr_o[19] ,
    \s1_addr_o[20] , \s1_addr_o[21] , \s1_addr_o[22] , \s1_addr_o[23] ,
    \s1_addr_o[24] , \s1_addr_o[25] , \s1_addr_o[26] , \s1_addr_o[27] ,
    \s1_addr_o[28] , \s1_addr_o[29] , \s1_addr_o[30] , \s1_addr_o[31] ,
    \s2_data_o[0] , \s2_data_o[1] , \s2_data_o[2] , \s2_data_o[3] ,
    \s2_data_o[4] , \s2_data_o[5] , \s2_data_o[6] , \s2_data_o[7] ,
    \s2_data_o[8] , \s2_data_o[9] , \s2_data_o[10] , \s2_data_o[11] ,
    \s2_data_o[12] , \s2_data_o[13] , \s2_data_o[14] , \s2_data_o[15] ,
    \s2_data_o[16] , \s2_data_o[17] , \s2_data_o[18] , \s2_data_o[19] ,
    \s2_data_o[20] , \s2_data_o[21] , \s2_data_o[22] , \s2_data_o[23] ,
    \s2_data_o[24] , \s2_data_o[25] , \s2_data_o[26] , \s2_data_o[27] ,
    \s2_data_o[28] , \s2_data_o[29] , \s2_data_o[30] , \s2_data_o[31] ,
    \s2_addr_o[0] , \s2_addr_o[1] , \s2_addr_o[2] , \s2_addr_o[3] ,
    \s2_addr_o[4] , \s2_addr_o[5] , \s2_addr_o[6] , \s2_addr_o[7] ,
    \s2_addr_o[8] , \s2_addr_o[9] , \s2_addr_o[10] , \s2_addr_o[11] ,
    \s2_addr_o[12] , \s2_addr_o[13] , \s2_addr_o[14] , \s2_addr_o[15] ,
    \s2_addr_o[16] , \s2_addr_o[17] , \s2_addr_o[18] , \s2_addr_o[19] ,
    \s2_addr_o[20] , \s2_addr_o[21] , \s2_addr_o[22] , \s2_addr_o[23] ,
    \s2_addr_o[24] , \s2_addr_o[25] , \s2_addr_o[26] , \s2_addr_o[27] ,
    \s2_addr_o[28] , \s2_addr_o[29] , \s2_addr_o[30] , \s2_addr_o[31] ,
    \s3_data_o[0] , \s3_data_o[1] , \s3_data_o[2] , \s3_data_o[3] ,
    \s3_data_o[4] , \s3_data_o[5] , \s3_data_o[6] , \s3_data_o[7] ,
    \s3_data_o[8] , \s3_data_o[9] , \s3_data_o[10] , \s3_data_o[11] ,
    \s3_data_o[12] , \s3_data_o[13] , \s3_data_o[14] , \s3_data_o[15] ,
    \s3_data_o[16] , \s3_data_o[17] , \s3_data_o[18] , \s3_data_o[19] ,
    \s3_data_o[20] , \s3_data_o[21] , \s3_data_o[22] , \s3_data_o[23] ,
    \s3_data_o[24] , \s3_data_o[25] , \s3_data_o[26] , \s3_data_o[27] ,
    \s3_data_o[28] , \s3_data_o[29] , \s3_data_o[30] , \s3_data_o[31] ,
    \s3_addr_o[0] , \s3_addr_o[1] , \s3_addr_o[2] , \s3_addr_o[3] ,
    \s3_addr_o[4] , \s3_addr_o[5] , \s3_addr_o[6] , \s3_addr_o[7] ,
    \s3_addr_o[8] , \s3_addr_o[9] , \s3_addr_o[10] , \s3_addr_o[11] ,
    \s3_addr_o[12] , \s3_addr_o[13] , \s3_addr_o[14] , \s3_addr_o[15] ,
    \s3_addr_o[16] , \s3_addr_o[17] , \s3_addr_o[18] , \s3_addr_o[19] ,
    \s3_addr_o[20] , \s3_addr_o[21] , \s3_addr_o[22] , \s3_addr_o[23] ,
    \s3_addr_o[24] , \s3_addr_o[25] , \s3_addr_o[26] , \s3_addr_o[27] ,
    \s3_addr_o[28] , \s3_addr_o[29] , \s3_addr_o[30] , \s3_addr_o[31] ,
    \s4_data_o[0] , \s4_data_o[1] , \s4_data_o[2] , \s4_data_o[3] ,
    \s4_data_o[4] , \s4_data_o[5] , \s4_data_o[6] , \s4_data_o[7] ,
    \s4_data_o[8] , \s4_data_o[9] , \s4_data_o[10] , \s4_data_o[11] ,
    \s4_data_o[12] , \s4_data_o[13] , \s4_data_o[14] , \s4_data_o[15] ,
    \s4_data_o[16] , \s4_data_o[17] , \s4_data_o[18] , \s4_data_o[19] ,
    \s4_data_o[20] , \s4_data_o[21] , \s4_data_o[22] , \s4_data_o[23] ,
    \s4_data_o[24] , \s4_data_o[25] , \s4_data_o[26] , \s4_data_o[27] ,
    \s4_data_o[28] , \s4_data_o[29] , \s4_data_o[30] , \s4_data_o[31] ,
    \s4_addr_o[0] , \s4_addr_o[1] , \s4_addr_o[2] , \s4_addr_o[3] ,
    \s4_addr_o[4] , \s4_addr_o[5] , \s4_addr_o[6] , \s4_addr_o[7] ,
    \s4_addr_o[8] , \s4_addr_o[9] , \s4_addr_o[10] , \s4_addr_o[11] ,
    \s4_addr_o[12] , \s4_addr_o[13] , \s4_addr_o[14] , \s4_addr_o[15] ,
    \s4_addr_o[16] , \s4_addr_o[17] , \s4_addr_o[18] , \s4_addr_o[19] ,
    \s4_addr_o[20] , \s4_addr_o[21] , \s4_addr_o[22] , \s4_addr_o[23] ,
    \s4_addr_o[24] , \s4_addr_o[25] , \s4_addr_o[26] , \s4_addr_o[27] ,
    \s4_addr_o[28] , \s4_addr_o[29] , \s4_addr_o[30] , \s4_addr_o[31] ,
    \s5_data_o[0] , \s5_data_o[1] , \s5_data_o[2] , \s5_data_o[3] ,
    \s5_data_o[4] , \s5_data_o[5] , \s5_data_o[6] , \s5_data_o[7] ,
    \s5_data_o[8] , \s5_data_o[9] , \s5_data_o[10] , \s5_data_o[11] ,
    \s5_data_o[12] , \s5_data_o[13] , \s5_data_o[14] , \s5_data_o[15] ,
    \s5_data_o[16] , \s5_data_o[17] , \s5_data_o[18] , \s5_data_o[19] ,
    \s5_data_o[20] , \s5_data_o[21] , \s5_data_o[22] , \s5_data_o[23] ,
    \s5_data_o[24] , \s5_data_o[25] , \s5_data_o[26] , \s5_data_o[27] ,
    \s5_data_o[28] , \s5_data_o[29] , \s5_data_o[30] , \s5_data_o[31] ,
    \s5_addr_o[0] , \s5_addr_o[1] , \s5_addr_o[2] , \s5_addr_o[3] ,
    \s5_addr_o[4] , \s5_addr_o[5] , \s5_addr_o[6] , \s5_addr_o[7] ,
    \s5_addr_o[8] , \s5_addr_o[9] , \s5_addr_o[10] , \s5_addr_o[11] ,
    \s5_addr_o[12] , \s5_addr_o[13] , \s5_addr_o[14] , \s5_addr_o[15] ,
    \s5_addr_o[16] , \s5_addr_o[17] , \s5_addr_o[18] , \s5_addr_o[19] ,
    \s5_addr_o[20] , \s5_addr_o[21] , \s5_addr_o[22] , \s5_addr_o[23] ,
    \s5_addr_o[24] , \s5_addr_o[25] , \s5_addr_o[26] , \s5_addr_o[27] ,
    \s5_addr_o[28] , \s5_addr_o[29] , \s5_addr_o[30] , \s5_addr_o[31] ,
    \s6_data_o[0] , \s6_data_o[1] , \s6_data_o[2] , \s6_data_o[3] ,
    \s6_data_o[4] , \s6_data_o[5] , \s6_data_o[6] , \s6_data_o[7] ,
    \s6_data_o[8] , \s6_data_o[9] , \s6_data_o[10] , \s6_data_o[11] ,
    \s6_data_o[12] , \s6_data_o[13] , \s6_data_o[14] , \s6_data_o[15] ,
    \s6_data_o[16] , \s6_data_o[17] , \s6_data_o[18] , \s6_data_o[19] ,
    \s6_data_o[20] , \s6_data_o[21] , \s6_data_o[22] , \s6_data_o[23] ,
    \s6_data_o[24] , \s6_data_o[25] , \s6_data_o[26] , \s6_data_o[27] ,
    \s6_data_o[28] , \s6_data_o[29] , \s6_data_o[30] , \s6_data_o[31] ,
    \s6_addr_o[0] , \s6_addr_o[1] , \s6_addr_o[2] , \s6_addr_o[3] ,
    \s6_addr_o[4] , \s6_addr_o[5] , \s6_addr_o[6] , \s6_addr_o[7] ,
    \s6_addr_o[8] , \s6_addr_o[9] , \s6_addr_o[10] , \s6_addr_o[11] ,
    \s6_addr_o[12] , \s6_addr_o[13] , \s6_addr_o[14] , \s6_addr_o[15] ,
    \s6_addr_o[16] , \s6_addr_o[17] , \s6_addr_o[18] , \s6_addr_o[19] ,
    \s6_addr_o[20] , \s6_addr_o[21] , \s6_addr_o[22] , \s6_addr_o[23] ,
    \s6_addr_o[24] , \s6_addr_o[25] , \s6_addr_o[26] , \s6_addr_o[27] ,
    \s6_addr_o[28] , \s6_addr_o[29] , \s6_addr_o[30] , \s6_addr_o[31] ,
    \s7_data_o[0] , \s7_data_o[1] , \s7_data_o[2] , \s7_data_o[3] ,
    \s7_data_o[4] , \s7_data_o[5] , \s7_data_o[6] , \s7_data_o[7] ,
    \s7_data_o[8] , \s7_data_o[9] , \s7_data_o[10] , \s7_data_o[11] ,
    \s7_data_o[12] , \s7_data_o[13] , \s7_data_o[14] , \s7_data_o[15] ,
    \s7_data_o[16] , \s7_data_o[17] , \s7_data_o[18] , \s7_data_o[19] ,
    \s7_data_o[20] , \s7_data_o[21] , \s7_data_o[22] , \s7_data_o[23] ,
    \s7_data_o[24] , \s7_data_o[25] , \s7_data_o[26] , \s7_data_o[27] ,
    \s7_data_o[28] , \s7_data_o[29] , \s7_data_o[30] , \s7_data_o[31] ,
    \s7_addr_o[0] , \s7_addr_o[1] , \s7_addr_o[2] , \s7_addr_o[3] ,
    \s7_addr_o[4] , \s7_addr_o[5] , \s7_addr_o[6] , \s7_addr_o[7] ,
    \s7_addr_o[8] , \s7_addr_o[9] , \s7_addr_o[10] , \s7_addr_o[11] ,
    \s7_addr_o[12] , \s7_addr_o[13] , \s7_addr_o[14] , \s7_addr_o[15] ,
    \s7_addr_o[16] , \s7_addr_o[17] , \s7_addr_o[18] , \s7_addr_o[19] ,
    \s7_addr_o[20] , \s7_addr_o[21] , \s7_addr_o[22] , \s7_addr_o[23] ,
    \s7_addr_o[24] , \s7_addr_o[25] , \s7_addr_o[26] , \s7_addr_o[27] ,
    \s7_addr_o[28] , \s7_addr_o[29] , \s7_addr_o[30] , \s7_addr_o[31] ,
    \s8_data_o[0] , \s8_data_o[1] , \s8_data_o[2] , \s8_data_o[3] ,
    \s8_data_o[4] , \s8_data_o[5] , \s8_data_o[6] , \s8_data_o[7] ,
    \s8_data_o[8] , \s8_data_o[9] , \s8_data_o[10] , \s8_data_o[11] ,
    \s8_data_o[12] , \s8_data_o[13] , \s8_data_o[14] , \s8_data_o[15] ,
    \s8_data_o[16] , \s8_data_o[17] , \s8_data_o[18] , \s8_data_o[19] ,
    \s8_data_o[20] , \s8_data_o[21] , \s8_data_o[22] , \s8_data_o[23] ,
    \s8_data_o[24] , \s8_data_o[25] , \s8_data_o[26] , \s8_data_o[27] ,
    \s8_data_o[28] , \s8_data_o[29] , \s8_data_o[30] , \s8_data_o[31] ,
    \s8_addr_o[0] , \s8_addr_o[1] , \s8_addr_o[2] , \s8_addr_o[3] ,
    \s8_addr_o[4] , \s8_addr_o[5] , \s8_addr_o[6] , \s8_addr_o[7] ,
    \s8_addr_o[8] , \s8_addr_o[9] , \s8_addr_o[10] , \s8_addr_o[11] ,
    \s8_addr_o[12] , \s8_addr_o[13] , \s8_addr_o[14] , \s8_addr_o[15] ,
    \s8_addr_o[16] , \s8_addr_o[17] , \s8_addr_o[18] , \s8_addr_o[19] ,
    \s8_addr_o[20] , \s8_addr_o[21] , \s8_addr_o[22] , \s8_addr_o[23] ,
    \s8_addr_o[24] , \s8_addr_o[25] , \s8_addr_o[26] , \s8_addr_o[27] ,
    \s8_addr_o[28] , \s8_addr_o[29] , \s8_addr_o[30] , \s8_addr_o[31] ,
    \s9_data_o[0] , \s9_data_o[1] , \s9_data_o[2] , \s9_data_o[3] ,
    \s9_data_o[4] , \s9_data_o[5] , \s9_data_o[6] , \s9_data_o[7] ,
    \s9_data_o[8] , \s9_data_o[9] , \s9_data_o[10] , \s9_data_o[11] ,
    \s9_data_o[12] , \s9_data_o[13] , \s9_data_o[14] , \s9_data_o[15] ,
    \s9_data_o[16] , \s9_data_o[17] , \s9_data_o[18] , \s9_data_o[19] ,
    \s9_data_o[20] , \s9_data_o[21] , \s9_data_o[22] , \s9_data_o[23] ,
    \s9_data_o[24] , \s9_data_o[25] , \s9_data_o[26] , \s9_data_o[27] ,
    \s9_data_o[28] , \s9_data_o[29] , \s9_data_o[30] , \s9_data_o[31] ,
    \s9_addr_o[0] , \s9_addr_o[1] , \s9_addr_o[2] , \s9_addr_o[3] ,
    \s9_addr_o[4] , \s9_addr_o[5] , \s9_addr_o[6] , \s9_addr_o[7] ,
    \s9_addr_o[8] , \s9_addr_o[9] , \s9_addr_o[10] , \s9_addr_o[11] ,
    \s9_addr_o[12] , \s9_addr_o[13] , \s9_addr_o[14] , \s9_addr_o[15] ,
    \s9_addr_o[16] , \s9_addr_o[17] , \s9_addr_o[18] , \s9_addr_o[19] ,
    \s9_addr_o[20] , \s9_addr_o[21] , \s9_addr_o[22] , \s9_addr_o[23] ,
    \s9_addr_o[24] , \s9_addr_o[25] , \s9_addr_o[26] , \s9_addr_o[27] ,
    \s9_addr_o[28] , \s9_addr_o[29] , \s9_addr_o[30] , \s9_addr_o[31] ,
    \s10_data_o[0] , \s10_data_o[1] , \s10_data_o[2] , \s10_data_o[3] ,
    \s10_data_o[4] , \s10_data_o[5] , \s10_data_o[6] , \s10_data_o[7] ,
    \s10_data_o[8] , \s10_data_o[9] , \s10_data_o[10] , \s10_data_o[11] ,
    \s10_data_o[12] , \s10_data_o[13] , \s10_data_o[14] , \s10_data_o[15] ,
    \s10_data_o[16] , \s10_data_o[17] , \s10_data_o[18] , \s10_data_o[19] ,
    \s10_data_o[20] , \s10_data_o[21] , \s10_data_o[22] , \s10_data_o[23] ,
    \s10_data_o[24] , \s10_data_o[25] , \s10_data_o[26] , \s10_data_o[27] ,
    \s10_data_o[28] , \s10_data_o[29] , \s10_data_o[30] , \s10_data_o[31] ,
    \s10_addr_o[0] , \s10_addr_o[1] , \s10_addr_o[2] , \s10_addr_o[3] ,
    \s10_addr_o[4] , \s10_addr_o[5] , \s10_addr_o[6] , \s10_addr_o[7] ,
    \s10_addr_o[8] , \s10_addr_o[9] , \s10_addr_o[10] , \s10_addr_o[11] ,
    \s10_addr_o[12] , \s10_addr_o[13] , \s10_addr_o[14] , \s10_addr_o[15] ,
    \s10_addr_o[16] , \s10_addr_o[17] , \s10_addr_o[18] , \s10_addr_o[19] ,
    \s10_addr_o[20] , \s10_addr_o[21] , \s10_addr_o[22] , \s10_addr_o[23] ,
    \s10_addr_o[24] , \s10_addr_o[25] , \s10_addr_o[26] , \s10_addr_o[27] ,
    \s10_addr_o[28] , \s10_addr_o[29] , \s10_addr_o[30] , \s10_addr_o[31] ,
    \s11_data_o[0] , \s11_data_o[1] , \s11_data_o[2] , \s11_data_o[3] ,
    \s11_data_o[4] , \s11_data_o[5] , \s11_data_o[6] , \s11_data_o[7] ,
    \s11_data_o[8] , \s11_data_o[9] , \s11_data_o[10] , \s11_data_o[11] ,
    \s11_data_o[12] , \s11_data_o[13] , \s11_data_o[14] , \s11_data_o[15] ,
    \s11_data_o[16] , \s11_data_o[17] , \s11_data_o[18] , \s11_data_o[19] ,
    \s11_data_o[20] , \s11_data_o[21] , \s11_data_o[22] , \s11_data_o[23] ,
    \s11_data_o[24] , \s11_data_o[25] , \s11_data_o[26] , \s11_data_o[27] ,
    \s11_data_o[28] , \s11_data_o[29] , \s11_data_o[30] , \s11_data_o[31] ,
    \s11_addr_o[0] , \s11_addr_o[1] , \s11_addr_o[2] , \s11_addr_o[3] ,
    \s11_addr_o[4] , \s11_addr_o[5] , \s11_addr_o[6] , \s11_addr_o[7] ,
    \s11_addr_o[8] , \s11_addr_o[9] , \s11_addr_o[10] , \s11_addr_o[11] ,
    \s11_addr_o[12] , \s11_addr_o[13] , \s11_addr_o[14] , \s11_addr_o[15] ,
    \s11_addr_o[16] , \s11_addr_o[17] , \s11_addr_o[18] , \s11_addr_o[19] ,
    \s11_addr_o[20] , \s11_addr_o[21] , \s11_addr_o[22] , \s11_addr_o[23] ,
    \s11_addr_o[24] , \s11_addr_o[25] , \s11_addr_o[26] , \s11_addr_o[27] ,
    \s11_addr_o[28] , \s11_addr_o[29] , \s11_addr_o[30] , \s11_addr_o[31] ,
    \s12_data_o[0] , \s12_data_o[1] , \s12_data_o[2] , \s12_data_o[3] ,
    \s12_data_o[4] , \s12_data_o[5] , \s12_data_o[6] , \s12_data_o[7] ,
    \s12_data_o[8] , \s12_data_o[9] , \s12_data_o[10] , \s12_data_o[11] ,
    \s12_data_o[12] , \s12_data_o[13] , \s12_data_o[14] , \s12_data_o[15] ,
    \s12_data_o[16] , \s12_data_o[17] , \s12_data_o[18] , \s12_data_o[19] ,
    \s12_data_o[20] , \s12_data_o[21] , \s12_data_o[22] , \s12_data_o[23] ,
    \s12_data_o[24] , \s12_data_o[25] , \s12_data_o[26] , \s12_data_o[27] ,
    \s12_data_o[28] , \s12_data_o[29] , \s12_data_o[30] , \s12_data_o[31] ,
    \s12_addr_o[0] , \s12_addr_o[1] , \s12_addr_o[2] , \s12_addr_o[3] ,
    \s12_addr_o[4] , \s12_addr_o[5] , \s12_addr_o[6] , \s12_addr_o[7] ,
    \s12_addr_o[8] , \s12_addr_o[9] , \s12_addr_o[10] , \s12_addr_o[11] ,
    \s12_addr_o[12] , \s12_addr_o[13] , \s12_addr_o[14] , \s12_addr_o[15] ,
    \s12_addr_o[16] , \s12_addr_o[17] , \s12_addr_o[18] , \s12_addr_o[19] ,
    \s12_addr_o[20] , \s12_addr_o[21] , \s12_addr_o[22] , \s12_addr_o[23] ,
    \s12_addr_o[24] , \s12_addr_o[25] , \s12_addr_o[26] , \s12_addr_o[27] ,
    \s12_addr_o[28] , \s12_addr_o[29] , \s12_addr_o[30] , \s12_addr_o[31] ,
    \s13_data_o[0] , \s13_data_o[1] , \s13_data_o[2] , \s13_data_o[3] ,
    \s13_data_o[4] , \s13_data_o[5] , \s13_data_o[6] , \s13_data_o[7] ,
    \s13_data_o[8] , \s13_data_o[9] , \s13_data_o[10] , \s13_data_o[11] ,
    \s13_data_o[12] , \s13_data_o[13] , \s13_data_o[14] , \s13_data_o[15] ,
    \s13_data_o[16] , \s13_data_o[17] , \s13_data_o[18] , \s13_data_o[19] ,
    \s13_data_o[20] , \s13_data_o[21] , \s13_data_o[22] , \s13_data_o[23] ,
    \s13_data_o[24] , \s13_data_o[25] , \s13_data_o[26] , \s13_data_o[27] ,
    \s13_data_o[28] , \s13_data_o[29] , \s13_data_o[30] , \s13_data_o[31] ,
    \s13_addr_o[0] , \s13_addr_o[1] , \s13_addr_o[2] , \s13_addr_o[3] ,
    \s13_addr_o[4] , \s13_addr_o[5] , \s13_addr_o[6] , \s13_addr_o[7] ,
    \s13_addr_o[8] , \s13_addr_o[9] , \s13_addr_o[10] , \s13_addr_o[11] ,
    \s13_addr_o[12] , \s13_addr_o[13] , \s13_addr_o[14] , \s13_addr_o[15] ,
    \s13_addr_o[16] , \s13_addr_o[17] , \s13_addr_o[18] , \s13_addr_o[19] ,
    \s13_addr_o[20] , \s13_addr_o[21] , \s13_addr_o[22] , \s13_addr_o[23] ,
    \s13_addr_o[24] , \s13_addr_o[25] , \s13_addr_o[26] , \s13_addr_o[27] ,
    \s13_addr_o[28] , \s13_addr_o[29] , \s13_addr_o[30] , \s13_addr_o[31] ,
    \s14_data_o[0] , \s14_data_o[1] , \s14_data_o[2] , \s14_data_o[3] ,
    \s14_data_o[4] , \s14_data_o[5] , \s14_data_o[6] , \s14_data_o[7] ,
    \s14_data_o[8] , \s14_data_o[9] , \s14_data_o[10] , \s14_data_o[11] ,
    \s14_data_o[12] , \s14_data_o[13] , \s14_data_o[14] , \s14_data_o[15] ,
    \s14_data_o[16] , \s14_data_o[17] , \s14_data_o[18] , \s14_data_o[19] ,
    \s14_data_o[20] , \s14_data_o[21] , \s14_data_o[22] , \s14_data_o[23] ,
    \s14_data_o[24] , \s14_data_o[25] , \s14_data_o[26] , \s14_data_o[27] ,
    \s14_data_o[28] , \s14_data_o[29] , \s14_data_o[30] , \s14_data_o[31] ,
    \s14_addr_o[0] , \s14_addr_o[1] , \s14_addr_o[2] , \s14_addr_o[3] ,
    \s14_addr_o[4] , \s14_addr_o[5] , \s14_addr_o[6] , \s14_addr_o[7] ,
    \s14_addr_o[8] , \s14_addr_o[9] , \s14_addr_o[10] , \s14_addr_o[11] ,
    \s14_addr_o[12] , \s14_addr_o[13] , \s14_addr_o[14] , \s14_addr_o[15] ,
    \s14_addr_o[16] , \s14_addr_o[17] , \s14_addr_o[18] , \s14_addr_o[19] ,
    \s14_addr_o[20] , \s14_addr_o[21] , \s14_addr_o[22] , \s14_addr_o[23] ,
    \s14_addr_o[24] , \s14_addr_o[25] , \s14_addr_o[26] , \s14_addr_o[27] ,
    \s14_addr_o[28] , \s14_addr_o[29] , \s14_addr_o[30] , \s14_addr_o[31] ,
    \s15_data_o[0] , \s15_data_o[1] , \s15_data_o[2] , \s15_data_o[3] ,
    \s15_data_o[4] , \s15_data_o[5] , \s15_data_o[6] , \s15_data_o[7] ,
    \s15_data_o[8] , \s15_data_o[9] , \s15_data_o[10] , \s15_data_o[11] ,
    \s15_data_o[12] , \s15_data_o[13] , \s15_data_o[14] , \s15_data_o[15] ,
    \s15_data_o[16] , \s15_data_o[17] , \s15_data_o[18] , \s15_data_o[19] ,
    \s15_data_o[20] , \s15_data_o[21] , \s15_data_o[22] , \s15_data_o[23] ,
    \s15_data_o[24] , \s15_data_o[25] , \s15_data_o[26] , \s15_data_o[27] ,
    \s15_data_o[28] , \s15_data_o[29] , \s15_data_o[30] , \s15_data_o[31] ,
    \s15_addr_o[0] , \s15_addr_o[1] , \s15_addr_o[2] , \s15_addr_o[3] ,
    \s15_addr_o[4] , \s15_addr_o[5] , \s15_addr_o[6] , \s15_addr_o[7] ,
    \s15_addr_o[8] , \s15_addr_o[9] , \s15_addr_o[10] , \s15_addr_o[11] ,
    \s15_addr_o[12] , \s15_addr_o[13] , \s15_addr_o[14] , \s15_addr_o[15] ,
    \s15_addr_o[16] , \s15_addr_o[17] , \s15_addr_o[18] , \s15_addr_o[19] ,
    \s15_addr_o[20] , \s15_addr_o[21] , \s15_addr_o[22] , \s15_addr_o[23] ,
    \s15_addr_o[24] , \s15_addr_o[25] , \s15_addr_o[26] , \s15_addr_o[27] ,
    \s15_addr_o[28] , \s15_addr_o[29] , \s15_addr_o[30] , \s15_addr_o[31] ,
    m0_ack_o, m0_err_o, m0_rty_o, m1_ack_o, m1_err_o, m1_rty_o, m2_ack_o,
    m2_err_o, m2_rty_o, m3_ack_o, m3_err_o, m3_rty_o, m4_ack_o, m4_err_o,
    m4_rty_o, m5_ack_o, m5_err_o, m5_rty_o, m6_ack_o, m6_err_o, m6_rty_o,
    m7_ack_o, m7_err_o, m7_rty_o, s0_we_o, s0_cyc_o, s0_stb_o, s1_we_o,
    s1_cyc_o, s1_stb_o, s2_we_o, s2_cyc_o, s2_stb_o, s3_we_o, s3_cyc_o,
    s3_stb_o, s4_we_o, s4_cyc_o, s4_stb_o, s5_we_o, s5_cyc_o, s5_stb_o,
    s6_we_o, s6_cyc_o, s6_stb_o, s7_we_o, s7_cyc_o, s7_stb_o, s8_we_o,
    s8_cyc_o, s8_stb_o, s9_we_o, s9_cyc_o, s9_stb_o, s10_we_o, s10_cyc_o,
    s10_stb_o, s11_we_o, s11_cyc_o, s11_stb_o, s12_we_o, s12_cyc_o,
    s12_stb_o, s13_we_o, s13_cyc_o, s13_stb_o, s14_we_o, s14_cyc_o,
    s14_stb_o, s15_we_o, s15_cyc_o, s15_stb_o, \s0_sel_o[0] ,
    \s0_sel_o[1] , \s0_sel_o[2] , \s0_sel_o[3] , \s1_sel_o[0] ,
    \s1_sel_o[1] , \s1_sel_o[2] , \s1_sel_o[3] , \s2_sel_o[0] ,
    \s2_sel_o[1] , \s2_sel_o[2] , \s2_sel_o[3] , \s3_sel_o[0] ,
    \s3_sel_o[1] , \s3_sel_o[2] , \s3_sel_o[3] , \s4_sel_o[0] ,
    \s4_sel_o[1] , \s4_sel_o[2] , \s4_sel_o[3] , \s5_sel_o[0] ,
    \s5_sel_o[1] , \s5_sel_o[2] , \s5_sel_o[3] , \s6_sel_o[0] ,
    \s6_sel_o[1] , \s6_sel_o[2] , \s6_sel_o[3] , \s7_sel_o[0] ,
    \s7_sel_o[1] , \s7_sel_o[2] , \s7_sel_o[3] , \s8_sel_o[0] ,
    \s8_sel_o[1] , \s8_sel_o[2] , \s8_sel_o[3] , \s9_sel_o[0] ,
    \s9_sel_o[1] , \s9_sel_o[2] , \s9_sel_o[3] , \s10_sel_o[0] ,
    \s10_sel_o[1] , \s10_sel_o[2] , \s10_sel_o[3] , \s11_sel_o[0] ,
    \s11_sel_o[1] , \s11_sel_o[2] , \s11_sel_o[3] , \s12_sel_o[0] ,
    \s12_sel_o[1] , \s12_sel_o[2] , \s12_sel_o[3] , \s13_sel_o[0] ,
    \s13_sel_o[1] , \s13_sel_o[2] , \s13_sel_o[3] , \s14_sel_o[0] ,
    \s14_sel_o[1] , \s14_sel_o[2] , \s14_sel_o[3] , \s15_sel_o[0] ,
    \s15_sel_o[1] , \s15_sel_o[2] , \s15_sel_o[3] ;
  reg \\rf_rf_dout_reg[14] , \\rf_rf_dout_reg[12] , \\rf_rf_dout_reg[11] ,
    \\rf_rf_dout_reg[9] , \\rf_rf_dout_reg[6] , \\rf_rf_dout_reg[5] ,
    \\rf_rf_dout_reg[4] , \\rf_rf_dout_reg[2] , \\rf_rf_dout_reg[1] ,
    \\rf_rf_dout_reg[15] , \\rf_rf_dout_reg[13] , \\rf_rf_dout_reg[10] ,
    \\rf_rf_dout_reg[8] , \\rf_rf_dout_reg[7] , \\rf_rf_dout_reg[3] ,
    \\rf_rf_dout_reg[0] , \\rf_conf15_reg[0] , \\rf_conf15_reg[10] ,
    \\rf_conf15_reg[11] , \\rf_conf15_reg[12] , \\rf_conf15_reg[13] ,
    \\rf_conf15_reg[14] , \\rf_conf15_reg[15] , \\rf_conf15_reg[1] ,
    \\rf_conf15_reg[2] , \\rf_conf15_reg[3] , \\rf_conf15_reg[4] ,
    \\rf_conf15_reg[5] , \\rf_conf15_reg[6] , \\rf_conf15_reg[7] ,
    \\rf_conf15_reg[8] , \\rf_conf15_reg[9] , \\rf_conf0_reg[0] ,
    \\rf_conf0_reg[10] , \\rf_conf0_reg[11] , \\rf_conf0_reg[12] ,
    \\rf_conf0_reg[13] , \\rf_conf0_reg[14] , \\rf_conf0_reg[15] ,
    \\rf_conf0_reg[1] , \\rf_conf0_reg[2] , \\rf_conf0_reg[3] ,
    \\rf_conf0_reg[4] , \\rf_conf0_reg[5] , \\rf_conf0_reg[6] ,
    \\rf_conf0_reg[7] , \\rf_conf0_reg[8] , \\rf_conf0_reg[9] ,
    \\rf_conf12_reg[0] , \\rf_conf12_reg[10] , \\rf_conf12_reg[11] ,
    \\rf_conf12_reg[12] , \\rf_conf12_reg[13] , \\rf_conf12_reg[14] ,
    \\rf_conf12_reg[15] , \\rf_conf12_reg[1] , \\rf_conf12_reg[2] ,
    \\rf_conf12_reg[3] , \\rf_conf12_reg[4] , \\rf_conf12_reg[5] ,
    \\rf_conf12_reg[6] , \\rf_conf12_reg[7] , \\rf_conf12_reg[8] ,
    \\rf_conf12_reg[9] , \\rf_conf13_reg[0] , \\rf_conf13_reg[10] ,
    \\rf_conf13_reg[11] , \\rf_conf13_reg[12] , \\rf_conf13_reg[13] ,
    \\rf_conf13_reg[14] , \\rf_conf13_reg[15] , \\rf_conf13_reg[1] ,
    \\rf_conf13_reg[4] , \\rf_conf13_reg[5] , \\rf_conf13_reg[6] ,
    \\rf_conf13_reg[7] , \\rf_conf13_reg[8] , \\rf_conf13_reg[9] ,
    \\rf_conf14_reg[0] , \\rf_conf14_reg[10] , \\rf_conf14_reg[11] ,
    \\rf_conf14_reg[12] , \\rf_conf14_reg[13] , \\rf_conf14_reg[14] ,
    \\rf_conf14_reg[15] , \\rf_conf14_reg[1] , \\rf_conf14_reg[3] ,
    \\rf_conf14_reg[4] , \\rf_conf14_reg[5] , \\rf_conf14_reg[6] ,
    \\rf_conf14_reg[7] , \\rf_conf14_reg[8] , \\rf_conf14_reg[9] ,
    \\rf_conf13_reg[2] , \\rf_conf13_reg[3] , \\rf_conf14_reg[2] ,
    \\rf_conf1_reg[0] , \\rf_conf1_reg[10] , \\rf_conf1_reg[11] ,
    \\rf_conf1_reg[12] , \\rf_conf1_reg[13] , \\rf_conf1_reg[14] ,
    \\rf_conf1_reg[15] , \\rf_conf1_reg[1] , \\rf_conf1_reg[2] ,
    \\rf_conf1_reg[3] , \\rf_conf1_reg[4] , \\rf_conf1_reg[5] ,
    \\rf_conf1_reg[6] , \\rf_conf1_reg[7] , \\rf_conf1_reg[8] ,
    \\rf_conf1_reg[9] , \\rf_conf2_reg[0] , \\rf_conf2_reg[10] ,
    \\rf_conf2_reg[11] , \\rf_conf2_reg[12] , \\rf_conf2_reg[13] ,
    \\rf_conf2_reg[14] , \\rf_conf2_reg[15] , \\rf_conf2_reg[1] ,
    \\rf_conf2_reg[2] , \\rf_conf2_reg[3] , \\rf_conf2_reg[4] ,
    \\rf_conf2_reg[5] , \\rf_conf2_reg[6] , \\rf_conf2_reg[7] ,
    \\rf_conf2_reg[8] , \\rf_conf2_reg[9] , \\rf_conf3_reg[0] ,
    \\rf_conf3_reg[10] , \\rf_conf3_reg[11] , \\rf_conf3_reg[12] ,
    \\rf_conf3_reg[13] , \\rf_conf3_reg[14] , \\rf_conf3_reg[15] ,
    \\rf_conf3_reg[1] , \\rf_conf3_reg[2] , \\rf_conf3_reg[3] ,
    \\rf_conf3_reg[4] , \\rf_conf3_reg[5] , \\rf_conf3_reg[6] ,
    \\rf_conf3_reg[7] , \\rf_conf3_reg[8] , \\rf_conf3_reg[9] ,
    \\rf_conf5_reg[0] , \\rf_conf5_reg[10] , \\rf_conf5_reg[11] ,
    \\rf_conf5_reg[12] , \\rf_conf5_reg[13] , \\rf_conf5_reg[14] ,
    \\rf_conf5_reg[15] , \\rf_conf5_reg[1] , \\rf_conf5_reg[2] ,
    \\rf_conf5_reg[3] , \\rf_conf5_reg[4] , \\rf_conf5_reg[5] ,
    \\rf_conf5_reg[6] , \\rf_conf5_reg[7] , \\rf_conf5_reg[8] ,
    \\rf_conf5_reg[9] , \\rf_conf7_reg[0] , \\rf_conf7_reg[10] ,
    \\rf_conf7_reg[11] , \\rf_conf7_reg[12] , \\rf_conf7_reg[13] ,
    \\rf_conf7_reg[14] , \\rf_conf7_reg[15] , \\rf_conf7_reg[1] ,
    \\rf_conf7_reg[2] , \\rf_conf7_reg[3] , \\rf_conf7_reg[4] ,
    \\rf_conf7_reg[5] , \\rf_conf7_reg[6] , \\rf_conf7_reg[7] ,
    \\rf_conf7_reg[8] , \\rf_conf7_reg[9] , \\rf_conf10_reg[0] ,
    \\rf_conf10_reg[10] , \\rf_conf10_reg[11] , \\rf_conf10_reg[12] ,
    \\rf_conf10_reg[13] , \\rf_conf10_reg[14] , \\rf_conf10_reg[15] ,
    \\rf_conf10_reg[1] , \\rf_conf10_reg[2] , \\rf_conf10_reg[3] ,
    \\rf_conf10_reg[4] , \\rf_conf10_reg[5] , \\rf_conf10_reg[6] ,
    \\rf_conf10_reg[7] , \\rf_conf10_reg[8] , \\rf_conf10_reg[9] ,
    \\rf_conf11_reg[0] , \\rf_conf11_reg[10] , \\rf_conf11_reg[11] ,
    \\rf_conf11_reg[12] , \\rf_conf11_reg[13] , \\rf_conf11_reg[14] ,
    \\rf_conf11_reg[15] , \\rf_conf11_reg[1] , \\rf_conf11_reg[4] ,
    \\rf_conf11_reg[5] , \\rf_conf11_reg[6] , \\rf_conf11_reg[7] ,
    \\rf_conf11_reg[8] , \\rf_conf11_reg[9] , \\rf_conf11_reg[2] ,
    \\rf_conf11_reg[3] , \\rf_conf4_reg[0] , \\rf_conf4_reg[10] ,
    \\rf_conf4_reg[11] , \\rf_conf4_reg[12] , \\rf_conf4_reg[13] ,
    \\rf_conf4_reg[14] , \\rf_conf4_reg[15] , \\rf_conf4_reg[1] ,
    \\rf_conf4_reg[4] , \\rf_conf4_reg[5] , \\rf_conf4_reg[6] ,
    \\rf_conf4_reg[7] , \\rf_conf4_reg[8] , \\rf_conf4_reg[9] ,
    \\rf_conf4_reg[2] , \\rf_conf4_reg[3] , \\rf_conf6_reg[0] ,
    \\rf_conf6_reg[10] , \\rf_conf6_reg[11] , \\rf_conf6_reg[12] ,
    \\rf_conf6_reg[13] , \\rf_conf6_reg[14] , \\rf_conf6_reg[15] ,
    \\rf_conf6_reg[1] , \\rf_conf6_reg[4] , \\rf_conf6_reg[5] ,
    \\rf_conf6_reg[6] , \\rf_conf6_reg[7] , \\rf_conf6_reg[8] ,
    \\rf_conf6_reg[9] , \\rf_conf6_reg[2] , \\rf_conf6_reg[3] ,
    \\rf_conf9_reg[0] , \\rf_conf9_reg[10] , \\rf_conf9_reg[11] ,
    \\rf_conf9_reg[12] , \\rf_conf9_reg[13] , \\rf_conf9_reg[14] ,
    \\rf_conf9_reg[15] , \\rf_conf9_reg[1] , \\rf_conf9_reg[2] ,
    \\rf_conf9_reg[3] , \\rf_conf9_reg[4] , \\rf_conf9_reg[5] ,
    \\rf_conf9_reg[6] , \\rf_conf9_reg[7] , \\rf_conf9_reg[8] ,
    \\rf_conf9_reg[9] , \\rf_conf8_reg[0] , \\rf_conf8_reg[10] ,
    \\rf_conf8_reg[11] , \\rf_conf8_reg[12] , \\rf_conf8_reg[13] ,
    \\rf_conf8_reg[14] , \\rf_conf8_reg[15] , \\rf_conf8_reg[1] ,
    \\rf_conf8_reg[4] , \\rf_conf8_reg[5] , \\rf_conf8_reg[6] ,
    \\rf_conf8_reg[7] , \\rf_conf8_reg[8] , \\rf_conf8_reg[9] ,
    \\rf_conf8_reg[2] , \\rf_conf8_reg[3] , rf_rf_we_reg, rf_rf_ack_reg,
    \\s14_msel_arb2_state_reg[0] , \\s10_msel_arb0_state_reg[1] ,
    \\s11_msel_arb0_state_reg[1] , \\s12_msel_arb0_state_reg[1] ,
    \\s13_msel_arb0_state_reg[1] , \\s14_msel_arb0_state_reg[1] ,
    \\s15_msel_arb0_state_reg[1] , \\s1_msel_arb0_state_reg[1] ,
    \\s2_msel_arb0_state_reg[1] , \\s3_msel_arb0_state_reg[1] ,
    \\s4_msel_arb0_state_reg[1] , \\s5_msel_arb0_state_reg[1] ,
    \\s6_msel_arb0_state_reg[1] , \\s8_msel_arb0_state_reg[1] ,
    \\s9_msel_arb0_state_reg[1] , \\s0_msel_arb0_state_reg[1] ,
    \\s11_msel_arb0_state_reg[0] , \\s11_msel_arb1_state_reg[1] ,
    \\s12_msel_arb0_state_reg[0] , \\s13_msel_arb0_state_reg[0] ,
    \\s13_msel_arb2_state_reg[0] , \\s14_msel_arb0_state_reg[0] ,
    \\s15_msel_arb2_state_reg[0] , \\s15_msel_arb3_state_reg[1] ,
    \\s3_msel_arb0_state_reg[0] , \\s4_msel_arb0_state_reg[0] ,
    \\s4_msel_arb2_state_reg[0] , \\s4_msel_arb2_state_reg[1] ,
    \\s5_msel_arb0_state_reg[0] , \\s5_msel_arb3_state_reg[1] ,
    \\s6_msel_arb0_state_reg[0] , \\s6_msel_arb1_state_reg[0] ,
    \\s6_msel_arb1_state_reg[1] , \\s7_msel_arb0_state_reg[0] ,
    \\s8_msel_arb0_state_reg[0] , \\s8_msel_arb1_state_reg[1] ,
    \\s8_msel_arb3_state_reg[1] , \\s9_msel_arb3_state_reg[0] ,
    \\s9_msel_arb2_state_reg[0] , \\s0_msel_arb2_state_reg[0] ,
    \\s7_msel_arb0_state_reg[1] , \\s10_msel_arb2_state_reg[1] ,
    \\s10_msel_arb2_state_reg[0] , \\s11_msel_arb2_state_reg[1] ,
    \\s11_msel_arb3_state_reg[1] , \\s12_msel_arb1_state_reg[1] ,
    \\s12_msel_arb2_state_reg[0] , \\s12_msel_arb2_state_reg[1] ,
    \\s13_msel_arb1_state_reg[1] , \\s13_msel_arb2_state_reg[1] ,
    \\s14_msel_arb2_state_reg[1] , \\s14_msel_arb2_state_reg[2] ,
    \\s15_msel_arb0_state_reg[0] , \\s15_msel_arb1_state_reg[1] ,
    \\s15_msel_arb2_state_reg[1] , \\s15_msel_arb2_state_reg[2] ,
    \\s1_msel_arb0_state_reg[0] , \\s1_msel_arb2_state_reg[0] ,
    \\s1_msel_arb2_state_reg[1] , \\s2_msel_arb2_state_reg[0] ,
    \\s2_msel_arb2_state_reg[1] , \\s2_msel_arb0_state_reg[0] ,
    \\s3_msel_arb1_state_reg[1] , \\s3_msel_arb2_state_reg[0] ,
    \\s3_msel_arb2_state_reg[1] , \\s3_msel_arb3_state_reg[1] ,
    \\s4_msel_arb2_state_reg[2] , \\s5_msel_arb1_state_reg[1] ,
    \\s5_msel_arb2_state_reg[1] , \\s5_msel_arb3_state_reg[0] ,
    \\s5_msel_arb3_state_reg[2] , \\s6_msel_arb2_state_reg[1] ,
    \\s6_msel_arb2_state_reg[0] , \\s6_msel_arb3_state_reg[1] ,
    \\s6_msel_arb3_state_reg[0] , \\s7_msel_arb2_state_reg[0] ,
    \\s7_msel_arb2_state_reg[1] , \\s8_msel_arb2_state_reg[0] ,
    \\s8_msel_arb2_state_reg[1] , \\s8_msel_arb3_state_reg[0] ,
    \\s9_msel_arb0_state_reg[0] , \\s9_msel_arb2_state_reg[2] ,
    \\s0_msel_arb0_state_reg[0] , \\s0_msel_arb2_state_reg[1] ,
    \\s0_msel_arb2_state_reg[2] , \\s0_msel_arb3_state_reg[0] ,
    \\s14_msel_arb3_state_reg[0] , \\s12_msel_arb1_state_reg[0] ,
    \\s10_msel_arb1_state_reg[0] , \\s10_msel_arb1_state_reg[1] ,
    \\s10_msel_arb2_state_reg[2] , \\s11_msel_arb0_state_reg[2] ,
    \\s11_msel_arb1_state_reg[2] , \\s11_msel_arb2_state_reg[0] ,
    \\s11_msel_arb2_state_reg[2] , \\s11_msel_arb1_state_reg[0] ,
    \\s11_msel_arb3_state_reg[2] , \\s12_msel_arb0_state_reg[2] ,
    \\s12_msel_arb1_state_reg[2] , \\s12_msel_arb2_state_reg[2] ,
    \\s13_msel_arb0_state_reg[2] , \\s12_msel_arb3_state_reg[1] ,
    \\s13_msel_arb2_state_reg[2] , \\s13_msel_arb3_state_reg[1] ,
    \\s14_msel_arb1_state_reg[2] , \\s14_msel_arb1_state_reg[1] ,
    \\s14_msel_arb0_state_reg[2] , \\s14_msel_arb3_state_reg[1] ,
    \\s14_msel_arb3_state_reg[2] , \\s15_msel_arb1_state_reg[0] ,
    \\s15_msel_arb3_state_reg[0] , \\s1_msel_arb0_state_reg[2] ,
    \\s1_msel_arb1_state_reg[1] , \\s1_msel_arb2_state_reg[2] ,
    \\s1_msel_arb3_state_reg[0] , \\s1_msel_arb3_state_reg[1] ,
    \\s2_msel_arb1_state_reg[1] , \\s2_msel_arb0_state_reg[2] ,
    \\s2_msel_arb2_state_reg[2] , \\s2_msel_arb3_state_reg[0] ,
    \\s2_msel_arb3_state_reg[1] , \\s3_msel_arb1_state_reg[0] ,
    \\s3_msel_arb0_state_reg[2] , \\s3_msel_arb2_state_reg[2] ,
    \\s4_msel_arb1_state_reg[0] , \\s4_msel_arb1_state_reg[1] ,
    \\s4_msel_arb3_state_reg[0] , \\s5_msel_arb1_state_reg[0] ,
    \\s5_msel_arb1_state_reg[2] , \\s5_msel_arb0_state_reg[2] ,
    \\s6_msel_arb0_state_reg[2] , \\s6_msel_arb1_state_reg[2] ,
    \\s6_msel_arb2_state_reg[2] , \\s7_msel_arb1_state_reg[0] ,
    \\s7_msel_arb1_state_reg[2] , \\s7_msel_arb0_state_reg[2] ,
    \\s7_msel_arb2_state_reg[2] , \\s7_msel_arb3_state_reg[2] ,
    \\s8_msel_arb0_state_reg[2] , \\s8_msel_arb1_state_reg[0] ,
    \\s7_msel_arb3_state_reg[1] , \\s8_msel_arb3_state_reg[2] ,
    \\s9_msel_arb0_state_reg[2] , \\s9_msel_arb2_state_reg[1] ,
    \\s9_msel_arb1_state_reg[2] , \\s9_msel_arb3_state_reg[1] ,
    \\s0_msel_arb0_state_reg[2] , \\s0_msel_arb1_state_reg[1] ,
    \\s0_msel_arb1_state_reg[2] , \\s10_msel_arb0_state_reg[0] ,
    \\s0_msel_arb3_state_reg[2] , \\s13_msel_arb1_state_reg[0] ,
    \\s10_msel_arb1_state_reg[2] , \\s11_msel_arb3_state_reg[0] ,
    \\s9_msel_arb3_state_reg[2] , \\s9_msel_arb1_state_reg[0] ,
    \\s8_msel_arb2_state_reg[2] , \\s8_msel_arb1_state_reg[2] ,
    \\s5_msel_arb2_state_reg[2] , \\s5_msel_arb2_state_reg[0] ,
    \\s4_msel_arb1_state_reg[2] , \\s4_msel_arb3_state_reg[1] ,
    \\s4_msel_arb0_state_reg[2] , \\s3_msel_arb1_state_reg[2] ,
    \\s1_msel_arb3_state_reg[2] , \\s1_msel_arb1_state_reg[0] ,
    \\s1_msel_arb1_state_reg[2] , \\s13_msel_arb1_state_reg[2] ,
    \\s13_msel_arb3_state_reg[2] , \\s10_msel_arb0_state_reg[2] ,
    \\s10_msel_arb3_state_reg[2] , \\s12_msel_arb3_state_reg[0] ,
    \\s12_msel_arb3_state_reg[2] , \\s13_msel_arb3_state_reg[0] ,
    \\s14_msel_arb1_state_reg[0] , \\s15_msel_arb1_state_reg[2] ,
    \\s15_msel_arb3_state_reg[2] , \\s2_msel_arb1_state_reg[0] ,
    \\s2_msel_arb1_state_reg[2] , \\s3_msel_arb3_state_reg[0] ,
    \\s3_msel_arb3_state_reg[2] , \\s4_msel_arb3_state_reg[2] ,
    \\s9_msel_arb1_state_reg[1] , \\s0_msel_arb1_state_reg[0] ,
    \\s0_msel_arb3_state_reg[1] , \\s10_msel_arb3_state_reg[1] ,
    \\s10_msel_arb3_state_reg[0] , \\s6_msel_arb3_state_reg[2] ,
    \\s7_msel_arb3_state_reg[0] , \\s7_msel_arb1_state_reg[1] ,
    \\s15_msel_arb0_state_reg[2] , \\s2_msel_arb3_state_reg[2] ,
    s15_next_reg, \\s13_msel_pri_out_reg[0] , \\s3_msel_pri_out_reg[0] ,
    \\s11_msel_pri_out_reg[0] , \\s12_msel_pri_out_reg[0] ,
    \\s5_msel_pri_out_reg[0] , \\s6_msel_pri_out_reg[0] ,
    \\s8_msel_pri_out_reg[0] , s12_next_reg, s13_next_reg, s14_next_reg,
    s3_next_reg, s6_next_reg, s9_next_reg, s8_next_reg, s0_next_reg,
    \\s8_msel_pri_out_reg[1] , \\s15_msel_pri_out_reg[0] ,
    \\s2_msel_pri_out_reg[0] , \\s1_msel_pri_out_reg[0] ,
    \\s7_msel_pri_out_reg[0] , \\s9_msel_pri_out_reg[0] ,
    \\s0_msel_pri_out_reg[0] , s11_next_reg, s2_next_reg, s4_next_reg,
    s7_next_reg, \\s11_msel_pri_out_reg[1] , \\s12_msel_pri_out_reg[1] ,
    \\s13_msel_pri_out_reg[1] , \\s3_msel_pri_out_reg[1] ,
    \\s5_msel_pri_out_reg[1] , \\s6_msel_pri_out_reg[1] , s5_next_reg,
    \\s14_msel_pri_out_reg[0] , \\s4_msel_pri_out_reg[0] ,
    \\s15_msel_pri_out_reg[1] , \\s10_msel_pri_out_reg[0] ,
    \\s2_msel_pri_out_reg[1] , \\s1_msel_pri_out_reg[1] ,
    \\s7_msel_pri_out_reg[1] , \\s0_msel_pri_out_reg[1] ,
    \\s9_msel_pri_out_reg[1] , \\s4_msel_pri_out_reg[1] ,
    \\s14_msel_pri_out_reg[1] , \\s10_msel_pri_out_reg[1] , s1_next_reg,
    s10_next_reg, m5_s0_cyc_o_reg, m2_s0_cyc_o_reg, m4_s0_cyc_o_reg,
    m5_s1_cyc_o_reg, m7_s0_cyc_o_reg, m6_s0_cyc_o_reg, m0_s0_cyc_o_reg,
    m1_s0_cyc_o_reg, m2_s1_cyc_o_reg, m7_s1_cyc_o_reg, m2_s15_cyc_o_reg,
    m4_s15_cyc_o_reg, m7_s12_cyc_o_reg, m7_s8_cyc_o_reg, m7_s4_cyc_o_reg,
    m7_s15_cyc_o_reg, m6_s15_cyc_o_reg, m6_s1_cyc_o_reg, m4_s1_cyc_o_reg,
    m1_s1_cyc_o_reg, m3_s0_cyc_o_reg, m0_s1_cyc_o_reg, m0_s13_cyc_o_reg,
    m0_s15_cyc_o_reg, m0_s7_cyc_o_reg, m4_s6_cyc_o_reg, m5_s5_cyc_o_reg,
    m4_s4_cyc_o_reg, m4_s5_cyc_o_reg, m7_s7_cyc_o_reg, m4_s7_cyc_o_reg,
    m2_s5_cyc_o_reg, m3_s15_cyc_o_reg, m3_s1_cyc_o_reg, m0_s2_cyc_o_reg,
    m0_s6_cyc_o_reg, m1_s15_cyc_o_reg, m1_s4_cyc_o_reg, m1_s8_cyc_o_reg,
    m2_s10_cyc_o_reg, m4_s10_cyc_o_reg, m4_s12_cyc_o_reg, m4_s8_cyc_o_reg,
    m5_s10_cyc_o_reg, m5_s12_cyc_o_reg, m5_s15_cyc_o_reg, m5_s8_cyc_o_reg,
    m6_s12_cyc_o_reg, m6_s4_cyc_o_reg, m7_s11_cyc_o_reg, m7_s5_cyc_o_reg,
    m6_s14_cyc_o_reg, m7_s6_cyc_o_reg, m6_s8_cyc_o_reg, m6_s9_cyc_o_reg,
    m6_s5_cyc_o_reg, m5_s4_cyc_o_reg, m6_s13_cyc_o_reg, m5_s6_cyc_o_reg,
    m4_s9_cyc_o_reg, m4_s13_cyc_o_reg, m4_s14_cyc_o_reg, m3_s9_cyc_o_reg,
    m3_s8_cyc_o_reg, m3_s10_cyc_o_reg, m2_s6_cyc_o_reg, m2_s9_cyc_o_reg,
    m1_s6_cyc_o_reg, m0_s8_cyc_o_reg, m1_s5_cyc_o_reg, m0_s9_cyc_o_reg,
    m1_s12_cyc_o_reg, m1_s10_cyc_o_reg, m0_s3_cyc_o_reg, m0_s5_cyc_o_reg,
    m0_s12_cyc_o_reg, m0_s11_cyc_o_reg, m0_s10_cyc_o_reg, m7_s3_cyc_o_reg,
    m1_s13_cyc_o_reg, m2_s11_cyc_o_reg, m3_s11_cyc_o_reg, m3_s13_cyc_o_reg,
    m3_s4_cyc_o_reg, m5_s2_cyc_o_reg, m6_s2_cyc_o_reg, m7_s9_cyc_o_reg,
    m7_s13_cyc_o_reg, m7_s2_cyc_o_reg, m7_s14_cyc_o_reg, m7_s10_cyc_o_reg,
    m6_s7_cyc_o_reg, m6_s6_cyc_o_reg, m6_s11_cyc_o_reg, m5_s9_cyc_o_reg,
    m6_s10_cyc_o_reg, m5_s7_cyc_o_reg, m5_s14_cyc_o_reg, m5_s3_cyc_o_reg,
    m5_s13_cyc_o_reg, m5_s11_cyc_o_reg, m4_s11_cyc_o_reg, m4_s2_cyc_o_reg,
    m2_s4_cyc_o_reg, m3_s5_cyc_o_reg, m3_s6_cyc_o_reg, m3_s7_cyc_o_reg,
    m3_s3_cyc_o_reg, m3_s14_cyc_o_reg, m3_s12_cyc_o_reg, m2_s8_cyc_o_reg,
    m2_s7_cyc_o_reg, m2_s13_cyc_o_reg, m2_s14_cyc_o_reg, m2_s2_cyc_o_reg,
    m1_s7_cyc_o_reg, m1_s9_cyc_o_reg, m1_s2_cyc_o_reg, m1_s14_cyc_o_reg,
    m1_s11_cyc_o_reg, m3_s2_cyc_o_reg, m0_s14_cyc_o_reg, m0_s4_cyc_o_reg,
    m4_s3_cyc_o_reg, m6_s3_cyc_o_reg, m2_s3_cyc_o_reg, m2_s12_cyc_o_reg,
    m1_s3_cyc_o_reg, s6_m4_cyc_r_reg, s15_m6_cyc_r_reg, s8_m2_cyc_r_reg,
    s5_m5_cyc_r_reg, s13_m5_cyc_r_reg, s3_m5_cyc_r_reg, s1_m1_cyc_r_reg,
    s11_m5_cyc_r_reg, s12_m5_cyc_r_reg, s15_m1_cyc_r_reg, s15_m3_cyc_r_reg,
    s10_m4_cyc_r_reg, s6_m5_cyc_r_reg, s8_m5_cyc_r_reg, s10_m5_cyc_r_reg,
    s5_m2_cyc_r_reg, s8_m1_cyc_r_reg, s4_m0_cyc_r_reg, s7_m1_cyc_r_reg,
    s5_m4_cyc_r_reg, s15_m2_cyc_r_reg, s10_m3_cyc_r_reg, s0_m0_cyc_r_reg,
    s5_m7_cyc_r_reg, s7_m7_cyc_r_reg, s11_m4_cyc_r_reg, s14_m5_cyc_r_reg,
    s15_m0_cyc_r_reg, s9_m7_cyc_r_reg, s0_m4_cyc_r_reg, s13_m4_cyc_r_reg,
    s2_m3_cyc_r_reg, s11_m1_cyc_r_reg, s13_m2_cyc_r_reg, s0_m2_cyc_r_reg,
    s9_m4_cyc_r_reg, s4_m7_cyc_r_reg, s13_m7_cyc_r_reg, s8_m0_cyc_r_reg,
    s7_m2_cyc_r_reg, s7_m3_cyc_r_reg, s3_m1_cyc_r_reg, s9_m0_cyc_r_reg,
    s10_m1_cyc_r_reg, s6_m7_cyc_r_reg, s11_m2_cyc_r_reg, s13_m3_cyc_r_reg,
    s10_m2_cyc_r_reg, s12_m3_cyc_r_reg, s14_m6_cyc_r_reg, s15_m7_cyc_r_reg,
    s10_m0_cyc_r_reg, s11_m3_cyc_r_reg, s4_m2_cyc_r_reg, s7_m6_cyc_r_reg,
    s9_m3_cyc_r_reg, s4_m6_cyc_r_reg, s0_m1_cyc_r_reg, s1_m2_cyc_r_reg,
    s10_m7_cyc_r_reg, s11_m6_cyc_r_reg, s4_m4_cyc_r_reg, s9_m2_cyc_r_reg,
    s1_m5_cyc_r_reg, s14_m3_cyc_r_reg, s12_m2_cyc_r_reg, s9_m1_cyc_r_reg,
    s3_m6_cyc_r_reg, s2_m6_cyc_r_reg, s6_m3_cyc_r_reg, s6_m6_cyc_r_reg,
    s8_m6_cyc_r_reg, s1_m4_cyc_r_reg, s6_m0_cyc_r_reg, s2_m7_cyc_r_reg,
    s3_m3_cyc_r_reg, s12_m0_cyc_r_reg, s1_m7_cyc_r_reg, s8_m7_cyc_r_reg,
    s2_m0_cyc_r_reg, s1_m3_cyc_r_reg, s1_m0_cyc_r_reg, s3_m2_cyc_r_reg,
    s13_m6_cyc_r_reg, s2_m1_cyc_r_reg, s3_m0_cyc_r_reg, s2_m5_cyc_r_reg,
    s2_m4_cyc_r_reg, s5_m6_cyc_r_reg, s14_m4_cyc_r_reg, s14_m0_cyc_r_reg,
    s15_m4_cyc_r_reg, s3_m4_cyc_r_reg, s2_m2_cyc_r_reg, s5_m3_cyc_r_reg,
    s12_m1_cyc_r_reg, s5_m0_cyc_r_reg, s0_m7_cyc_r_reg, s13_m0_cyc_r_reg,
    s1_m6_cyc_r_reg, s0_m5_cyc_r_reg, s15_m5_cyc_r_reg, s3_m7_cyc_r_reg,
    s9_m6_cyc_r_reg, s14_m2_cyc_r_reg, s4_m3_cyc_r_reg, s6_m2_cyc_r_reg,
    s7_m5_cyc_r_reg, s13_m1_cyc_r_reg, s0_m6_cyc_r_reg, s10_m6_cyc_r_reg,
    s8_m4_cyc_r_reg, s0_m3_cyc_r_reg, s4_m5_cyc_r_reg, s5_m1_cyc_r_reg,
    s6_m1_cyc_r_reg, s4_m1_cyc_r_reg, s14_m1_cyc_r_reg, s14_m7_cyc_r_reg,
    s12_m4_cyc_r_reg, s7_m0_cyc_r_reg, s12_m7_cyc_r_reg, s7_m4_cyc_r_reg,
    s8_m3_cyc_r_reg, s9_m5_cyc_r_reg, s11_m0_cyc_r_reg, s11_m7_cyc_r_reg,
    s12_m6_cyc_r_reg;
  wire \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3435]_ ,
    \new_[3436]_ , \new_[3437]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3441]_ , \new_[3442]_ , \new_[3443]_ ,
    \new_[3444]_ , \new_[3445]_ , \new_[3446]_ , \new_[3447]_ ,
    \new_[3448]_ , \new_[3449]_ , \new_[3450]_ , \new_[3451]_ ,
    \new_[3452]_ , \new_[3453]_ , \new_[3454]_ , \new_[3455]_ ,
    \new_[3456]_ , \new_[3457]_ , \new_[3458]_ , \new_[3459]_ ,
    \new_[3460]_ , \new_[3461]_ , \new_[3462]_ , \new_[3463]_ ,
    \new_[3464]_ , \new_[3465]_ , \new_[3466]_ , \new_[3467]_ ,
    \new_[3468]_ , \new_[3469]_ , \new_[3470]_ , \new_[3471]_ ,
    \new_[3472]_ , \new_[3473]_ , \new_[3474]_ , \new_[3475]_ ,
    \new_[3476]_ , \new_[3477]_ , \new_[3478]_ , \new_[3479]_ ,
    \new_[3480]_ , \new_[3481]_ , \new_[3482]_ , \new_[3483]_ ,
    \new_[3484]_ , \new_[3485]_ , \new_[3486]_ , \new_[3487]_ ,
    \new_[3488]_ , \new_[3489]_ , \new_[3490]_ , \new_[3491]_ ,
    \new_[3492]_ , \new_[3493]_ , \new_[3494]_ , \new_[3495]_ ,
    \new_[3496]_ , \new_[3497]_ , \new_[3498]_ , \new_[3499]_ ,
    \new_[3500]_ , \new_[3501]_ , \new_[3502]_ , \new_[3503]_ ,
    \new_[3504]_ , \new_[3505]_ , \new_[3506]_ , \new_[3507]_ ,
    \new_[3508]_ , \new_[3509]_ , \new_[3510]_ , \new_[3511]_ ,
    \new_[3512]_ , \new_[3513]_ , \new_[3514]_ , \new_[3515]_ ,
    \new_[3516]_ , \new_[3517]_ , \new_[3518]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3521]_ , \new_[3522]_ , \new_[3523]_ ,
    \new_[3524]_ , \new_[3525]_ , \new_[3526]_ , \new_[3527]_ ,
    \new_[3528]_ , \new_[3529]_ , \new_[3530]_ , \new_[3531]_ ,
    \new_[3532]_ , \new_[3533]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3536]_ , \new_[3537]_ , \new_[3538]_ , \new_[3539]_ ,
    \new_[3540]_ , \new_[3541]_ , \new_[3542]_ , \new_[3543]_ ,
    \new_[3544]_ , \new_[3545]_ , \new_[3546]_ , \new_[3547]_ ,
    \new_[3548]_ , \new_[3549]_ , \new_[3550]_ , \new_[3551]_ ,
    \new_[3552]_ , \new_[3553]_ , \new_[3554]_ , \new_[3555]_ ,
    \new_[3556]_ , \new_[3557]_ , \new_[3558]_ , \new_[3559]_ ,
    \new_[3560]_ , \new_[3561]_ , \new_[3562]_ , \new_[3563]_ ,
    \new_[3564]_ , \new_[3565]_ , \new_[3566]_ , \new_[3567]_ ,
    \new_[3568]_ , \new_[3569]_ , \new_[3570]_ , \new_[3571]_ ,
    \new_[3572]_ , \new_[3573]_ , \new_[3574]_ , \new_[3575]_ ,
    \new_[3576]_ , \new_[3577]_ , \new_[3578]_ , \new_[3579]_ ,
    \new_[3580]_ , \new_[3581]_ , \new_[3582]_ , \new_[3583]_ ,
    \new_[3584]_ , \new_[3585]_ , \new_[3586]_ , \new_[3587]_ ,
    \new_[3588]_ , \new_[3589]_ , \new_[3590]_ , \new_[3591]_ ,
    \new_[3592]_ , \new_[3593]_ , \new_[3594]_ , \new_[3595]_ ,
    \new_[3596]_ , \new_[3597]_ , \new_[3598]_ , \new_[3599]_ ,
    \new_[3600]_ , \new_[3601]_ , \new_[3602]_ , \new_[3603]_ ,
    \new_[3604]_ , \new_[3605]_ , \new_[3606]_ , \new_[3607]_ ,
    \new_[3608]_ , \new_[3609]_ , \new_[3610]_ , \new_[3611]_ ,
    \new_[3612]_ , \new_[3613]_ , \new_[3614]_ , \new_[3615]_ ,
    \new_[3616]_ , \new_[3617]_ , \new_[3618]_ , \new_[3619]_ ,
    \new_[3620]_ , \new_[3621]_ , \new_[3622]_ , \new_[3623]_ ,
    \new_[3624]_ , \new_[3625]_ , \new_[3626]_ , \new_[3627]_ ,
    \new_[3628]_ , \new_[3629]_ , \new_[3630]_ , \new_[3631]_ ,
    \new_[3632]_ , \new_[3633]_ , \new_[3634]_ , \new_[3635]_ ,
    \new_[3636]_ , \new_[3637]_ , \new_[3638]_ , \new_[3639]_ ,
    \new_[3640]_ , \new_[3641]_ , \new_[3642]_ , \new_[3643]_ ,
    \new_[3644]_ , \new_[3645]_ , \new_[3646]_ , \new_[3647]_ ,
    \new_[3648]_ , \new_[3649]_ , \new_[3650]_ , \new_[3651]_ ,
    \new_[3652]_ , \new_[3653]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3656]_ , \new_[3657]_ , \new_[3658]_ , \new_[3659]_ ,
    \new_[3660]_ , \new_[3661]_ , \new_[3662]_ , \new_[3663]_ ,
    \new_[3664]_ , \new_[3665]_ , \new_[3666]_ , \new_[3667]_ ,
    \new_[3668]_ , \new_[3669]_ , \new_[3670]_ , \new_[3671]_ ,
    \new_[3672]_ , \new_[3673]_ , \new_[3674]_ , \new_[3675]_ ,
    \new_[3676]_ , \new_[3677]_ , \new_[3678]_ , \new_[3679]_ ,
    \new_[3680]_ , \new_[3681]_ , \new_[3682]_ , \new_[3683]_ ,
    \new_[3684]_ , \new_[3685]_ , \new_[3686]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3690]_ , \new_[3691]_ ,
    \new_[3692]_ , \new_[3693]_ , \new_[3694]_ , \new_[3695]_ ,
    \new_[3696]_ , \new_[3697]_ , \new_[3698]_ , \new_[3699]_ ,
    \new_[3700]_ , \new_[3701]_ , \new_[3702]_ , \new_[3703]_ ,
    \new_[3704]_ , \new_[3705]_ , \new_[3706]_ , \new_[3707]_ ,
    \new_[3708]_ , \new_[3709]_ , \new_[3710]_ , \new_[3711]_ ,
    \new_[3712]_ , \new_[3713]_ , \new_[3714]_ , \new_[3715]_ ,
    \new_[3716]_ , \new_[3717]_ , \new_[3718]_ , \new_[3719]_ ,
    \new_[3720]_ , \new_[3721]_ , \new_[3722]_ , \new_[3723]_ ,
    \new_[3724]_ , \new_[3725]_ , \new_[3726]_ , \new_[3727]_ ,
    \new_[3728]_ , \new_[3729]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3732]_ , \new_[3733]_ , \new_[3734]_ , \new_[3735]_ ,
    \new_[3736]_ , \new_[3737]_ , \new_[3738]_ , \new_[3739]_ ,
    \new_[3740]_ , \new_[3741]_ , \new_[3742]_ , \new_[3743]_ ,
    \new_[3744]_ , \new_[3745]_ , \new_[3746]_ , \new_[3747]_ ,
    \new_[3748]_ , \new_[3749]_ , \new_[3750]_ , \new_[3751]_ ,
    \new_[3752]_ , \new_[3753]_ , \new_[3754]_ , \new_[3755]_ ,
    \new_[3756]_ , \new_[3757]_ , \new_[3758]_ , \new_[3759]_ ,
    \new_[3760]_ , \new_[3761]_ , \new_[3762]_ , \new_[3763]_ ,
    \new_[3764]_ , \new_[3765]_ , \new_[3766]_ , \new_[3767]_ ,
    \new_[3768]_ , \new_[3769]_ , \new_[3770]_ , \new_[3771]_ ,
    \new_[3772]_ , \new_[3773]_ , \new_[3774]_ , \new_[3775]_ ,
    \new_[3776]_ , \new_[3779]_ , \new_[3780]_ , \new_[3781]_ ,
    \new_[3802]_ , \new_[3803]_ , \new_[3804]_ , \new_[3805]_ ,
    \new_[3806]_ , \new_[3807]_ , \new_[3808]_ , \new_[3809]_ ,
    \new_[3810]_ , \new_[3811]_ , \new_[3812]_ , \new_[3813]_ ,
    \new_[3814]_ , \new_[3815]_ , \new_[3816]_ , \new_[3817]_ ,
    \new_[3818]_ , \new_[3819]_ , \new_[3820]_ , \new_[3821]_ ,
    \new_[3822]_ , \new_[3823]_ , \new_[3824]_ , \new_[3825]_ ,
    \new_[3828]_ , \new_[3829]_ , \new_[3830]_ , \new_[3831]_ ,
    \new_[3832]_ , \new_[3833]_ , \new_[3834]_ , \new_[3835]_ ,
    \new_[3836]_ , \new_[3837]_ , \new_[3838]_ , \new_[3848]_ ,
    \new_[3849]_ , \new_[3852]_ , \new_[3854]_ , \new_[3856]_ ,
    \new_[3858]_ , \new_[3859]_ , \new_[3860]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3865]_ , \new_[3866]_ , \new_[3867]_ ,
    \new_[3868]_ , \new_[3869]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3872]_ , \new_[3873]_ , \new_[3874]_ , \new_[3875]_ ,
    \new_[3876]_ , \new_[3877]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3880]_ , \new_[3881]_ , \new_[3882]_ , \new_[3883]_ ,
    \new_[3884]_ , \new_[3885]_ , \new_[3886]_ , \new_[3887]_ ,
    \new_[3888]_ , \new_[3903]_ , \new_[4018]_ , \new_[4019]_ ,
    \new_[4020]_ , \new_[4021]_ , \new_[4022]_ , \new_[4023]_ ,
    \new_[4024]_ , \new_[4025]_ , \new_[4026]_ , \new_[4027]_ ,
    \new_[4028]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4033]_ , \new_[4034]_ , \new_[4035]_ ,
    \new_[4036]_ , \new_[4037]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4041]_ , \new_[4042]_ , \new_[4043]_ ,
    \new_[4044]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4048]_ , \new_[4049]_ , \new_[4050]_ , \new_[4051]_ ,
    \new_[4052]_ , \new_[4053]_ , \new_[4054]_ , \new_[4055]_ ,
    \new_[4056]_ , \new_[4057]_ , \new_[4058]_ , \new_[4059]_ ,
    \new_[4060]_ , \new_[4061]_ , \new_[4062]_ , \new_[4063]_ ,
    \new_[4064]_ , \new_[4065]_ , \new_[4066]_ , \new_[4067]_ ,
    \new_[4068]_ , \new_[4069]_ , \new_[4070]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4074]_ , \new_[4075]_ ,
    \new_[4076]_ , \new_[4077]_ , \new_[4078]_ , \new_[4079]_ ,
    \new_[4080]_ , \new_[4081]_ , \new_[4082]_ , \new_[4083]_ ,
    \new_[4084]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4088]_ , \new_[4089]_ , \new_[4090]_ , \new_[4091]_ ,
    \new_[4092]_ , \new_[4093]_ , \new_[4094]_ , \new_[4095]_ ,
    \new_[4096]_ , \new_[4097]_ , \new_[4098]_ , \new_[4099]_ ,
    \new_[4100]_ , \new_[4101]_ , \new_[4102]_ , \new_[4103]_ ,
    \new_[4104]_ , \new_[4105]_ , \new_[4106]_ , \new_[4107]_ ,
    \new_[4108]_ , \new_[4109]_ , \new_[4110]_ , \new_[4111]_ ,
    \new_[4112]_ , \new_[4113]_ , \new_[4114]_ , \new_[4115]_ ,
    \new_[4116]_ , \new_[4117]_ , \new_[4118]_ , \new_[4119]_ ,
    \new_[4120]_ , \new_[4121]_ , \new_[4122]_ , \new_[4123]_ ,
    \new_[4124]_ , \new_[4125]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4128]_ , \new_[4129]_ , \new_[4130]_ , \new_[4131]_ ,
    \new_[4132]_ , \new_[4133]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4136]_ , \new_[4137]_ , \new_[4138]_ , \new_[4139]_ ,
    \new_[4140]_ , \new_[4141]_ , \new_[4142]_ , \new_[4143]_ ,
    \new_[4144]_ , \new_[4145]_ , \new_[4146]_ , \new_[4147]_ ,
    \new_[4148]_ , \new_[4149]_ , \new_[4150]_ , \new_[4151]_ ,
    \new_[4152]_ , \new_[4153]_ , \new_[4154]_ , \new_[4155]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4160]_ , \new_[4161]_ , \new_[4162]_ , \new_[4163]_ ,
    \new_[4164]_ , \new_[4165]_ , \new_[4166]_ , \new_[4167]_ ,
    \new_[4168]_ , \new_[4169]_ , \new_[4170]_ , \new_[4171]_ ,
    \new_[4172]_ , \new_[4173]_ , \new_[4174]_ , \new_[4175]_ ,
    \new_[4176]_ , \new_[4177]_ , \new_[4178]_ , \new_[4179]_ ,
    \new_[4180]_ , \new_[4181]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4184]_ , \new_[4185]_ , \new_[4186]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4192]_ , \new_[4193]_ , \new_[4194]_ , \new_[4195]_ ,
    \new_[4196]_ , \new_[4197]_ , \new_[4198]_ , \new_[4199]_ ,
    \new_[4200]_ , \new_[4201]_ , \new_[4202]_ , \new_[4203]_ ,
    \new_[4204]_ , \new_[4205]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4208]_ , \new_[4209]_ , \new_[4210]_ , \new_[4211]_ ,
    \new_[4212]_ , \new_[4213]_ , \new_[4214]_ , \new_[4215]_ ,
    \new_[4216]_ , \new_[4217]_ , \new_[4218]_ , \new_[4219]_ ,
    \new_[4220]_ , \new_[4221]_ , \new_[4222]_ , \new_[4223]_ ,
    \new_[4224]_ , \new_[4225]_ , \new_[4226]_ , \new_[4227]_ ,
    \new_[4228]_ , \new_[4229]_ , \new_[4230]_ , \new_[4231]_ ,
    \new_[4232]_ , \new_[4233]_ , \new_[4234]_ , \new_[4235]_ ,
    \new_[4236]_ , \new_[4237]_ , \new_[4238]_ , \new_[4239]_ ,
    \new_[4240]_ , \new_[4241]_ , \new_[4242]_ , \new_[4243]_ ,
    \new_[4244]_ , \new_[4245]_ , \new_[4246]_ , \new_[4247]_ ,
    \new_[4248]_ , \new_[4249]_ , \new_[4250]_ , \new_[4251]_ ,
    \new_[4252]_ , \new_[4253]_ , \new_[4254]_ , \new_[4255]_ ,
    \new_[4256]_ , \new_[4257]_ , \new_[4258]_ , \new_[4259]_ ,
    \new_[4260]_ , \new_[4261]_ , \new_[4262]_ , \new_[4263]_ ,
    \new_[4264]_ , \new_[4265]_ , \new_[4266]_ , \new_[4267]_ ,
    \new_[4268]_ , \new_[4269]_ , \new_[4270]_ , \new_[4271]_ ,
    \new_[4272]_ , \new_[4273]_ , \new_[4274]_ , \new_[4275]_ ,
    \new_[4276]_ , \new_[4277]_ , \new_[4278]_ , \new_[4279]_ ,
    \new_[4280]_ , \new_[4281]_ , \new_[4282]_ , \new_[4283]_ ,
    \new_[4300]_ , \new_[4301]_ , \new_[4302]_ , \new_[4303]_ ,
    \new_[4304]_ , \new_[4305]_ , \new_[4306]_ , \new_[4307]_ ,
    \new_[4308]_ , \new_[4309]_ , \new_[4310]_ , \new_[4311]_ ,
    \new_[4312]_ , \new_[4313]_ , \new_[4314]_ , \new_[4315]_ ,
    \new_[4316]_ , \new_[4317]_ , \new_[4318]_ , \new_[4319]_ ,
    \new_[4320]_ , \new_[4321]_ , \new_[4322]_ , \new_[4323]_ ,
    \new_[4324]_ , \new_[4325]_ , \new_[4326]_ , \new_[4327]_ ,
    \new_[4328]_ , \new_[4329]_ , \new_[4330]_ , \new_[4331]_ ,
    \new_[4332]_ , \new_[4333]_ , \new_[4334]_ , \new_[4335]_ ,
    \new_[4336]_ , \new_[4337]_ , \new_[4338]_ , \new_[4339]_ ,
    \new_[4340]_ , \new_[4341]_ , \new_[4342]_ , \new_[4343]_ ,
    \new_[4344]_ , \new_[4345]_ , \new_[4346]_ , \new_[4347]_ ,
    \new_[4348]_ , \new_[4349]_ , \new_[4350]_ , \new_[4351]_ ,
    \new_[4352]_ , \new_[4353]_ , \new_[4354]_ , \new_[4355]_ ,
    \new_[4356]_ , \new_[4357]_ , \new_[4358]_ , \new_[4359]_ ,
    \new_[4360]_ , \new_[4361]_ , \new_[4362]_ , \new_[4363]_ ,
    \new_[4364]_ , \new_[4365]_ , \new_[4366]_ , \new_[4367]_ ,
    \new_[4368]_ , \new_[4369]_ , \new_[4370]_ , \new_[4371]_ ,
    \new_[4372]_ , \new_[4373]_ , \new_[4374]_ , \new_[4375]_ ,
    \new_[4376]_ , \new_[4377]_ , \new_[4378]_ , \new_[4379]_ ,
    \new_[4380]_ , \new_[4381]_ , \new_[4382]_ , \new_[4383]_ ,
    \new_[4384]_ , \new_[4385]_ , \new_[4386]_ , \new_[4387]_ ,
    \new_[4388]_ , \new_[4389]_ , \new_[4390]_ , \new_[4391]_ ,
    \new_[4392]_ , \new_[4393]_ , \new_[4394]_ , \new_[4395]_ ,
    \new_[4396]_ , \new_[4397]_ , \new_[4398]_ , \new_[4399]_ ,
    \new_[4400]_ , \new_[4401]_ , \new_[4402]_ , \new_[4403]_ ,
    \new_[4404]_ , \new_[4405]_ , \new_[4406]_ , \new_[4407]_ ,
    \new_[4408]_ , \new_[4409]_ , \new_[4410]_ , \new_[4411]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4416]_ , \new_[4417]_ , \new_[4418]_ , \new_[4419]_ ,
    \new_[4420]_ , \new_[4421]_ , \new_[4422]_ , \new_[4423]_ ,
    \new_[4424]_ , \new_[4425]_ , \new_[4426]_ , \new_[4427]_ ,
    \new_[4428]_ , \new_[4429]_ , \new_[4430]_ , \new_[4431]_ ,
    \new_[4432]_ , \new_[4433]_ , \new_[4434]_ , \new_[4435]_ ,
    \new_[4436]_ , \new_[4437]_ , \new_[4438]_ , \new_[4439]_ ,
    \new_[4440]_ , \new_[4441]_ , \new_[4442]_ , \new_[4443]_ ,
    \new_[4444]_ , \new_[4445]_ , \new_[4446]_ , \new_[4447]_ ,
    \new_[4448]_ , \new_[4449]_ , \new_[4450]_ , \new_[4451]_ ,
    \new_[4452]_ , \new_[4453]_ , \new_[4454]_ , \new_[4455]_ ,
    \new_[4600]_ , \new_[4601]_ , \new_[4602]_ , \new_[4603]_ ,
    \new_[4604]_ , \new_[4605]_ , \new_[4606]_ , \new_[4607]_ ,
    \new_[4608]_ , \new_[4609]_ , \new_[4610]_ , \new_[4611]_ ,
    \new_[4612]_ , \new_[4613]_ , \new_[4614]_ , \new_[4615]_ ,
    \new_[4616]_ , \new_[4617]_ , \new_[4618]_ , \new_[4619]_ ,
    \new_[4620]_ , \new_[4621]_ , \new_[4622]_ , \new_[4623]_ ,
    \new_[4624]_ , \new_[4625]_ , \new_[4626]_ , \new_[4627]_ ,
    \new_[4628]_ , \new_[4629]_ , \new_[4630]_ , \new_[4631]_ ,
    \new_[4632]_ , \new_[4633]_ , \new_[4634]_ , \new_[4635]_ ,
    \new_[4636]_ , \new_[4637]_ , \new_[4638]_ , \new_[4639]_ ,
    \new_[4640]_ , \new_[4641]_ , \new_[4642]_ , \new_[4643]_ ,
    \new_[4644]_ , \new_[4645]_ , \new_[4646]_ , \new_[4647]_ ,
    \new_[4648]_ , \new_[4649]_ , \new_[4650]_ , \new_[4651]_ ,
    \new_[4652]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4657]_ , \new_[4658]_ , \new_[4659]_ ,
    \new_[4660]_ , \new_[4661]_ , \new_[4662]_ , \new_[4663]_ ,
    \new_[4664]_ , \new_[4665]_ , \new_[4666]_ , \new_[4667]_ ,
    \new_[4668]_ , \new_[4669]_ , \new_[4670]_ , \new_[4671]_ ,
    \new_[4672]_ , \new_[4673]_ , \new_[4674]_ , \new_[4675]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4678]_ , \new_[4679]_ ,
    \new_[4680]_ , \new_[4681]_ , \new_[4682]_ , \new_[4683]_ ,
    \new_[4684]_ , \new_[4685]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4689]_ , \new_[4690]_ , \new_[4691]_ ,
    \new_[4692]_ , \new_[4693]_ , \new_[4694]_ , \new_[4695]_ ,
    \new_[4696]_ , \new_[4697]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4700]_ , \new_[4701]_ , \new_[4702]_ , \new_[4703]_ ,
    \new_[4704]_ , \new_[4705]_ , \new_[4706]_ , \new_[4707]_ ,
    \new_[4708]_ , \new_[4709]_ , \new_[4710]_ , \new_[4711]_ ,
    \new_[4712]_ , \new_[4713]_ , \new_[4714]_ , \new_[4715]_ ,
    \new_[4716]_ , \new_[4717]_ , \new_[4718]_ , \new_[4719]_ ,
    \new_[4720]_ , \new_[4721]_ , \new_[4722]_ , \new_[4723]_ ,
    \new_[4724]_ , \new_[4725]_ , \new_[4726]_ , \new_[4727]_ ,
    \new_[4728]_ , \new_[4729]_ , \new_[4730]_ , \new_[4731]_ ,
    \new_[4732]_ , \new_[4733]_ , \new_[4734]_ , \new_[4735]_ ,
    \new_[4736]_ , \new_[4737]_ , \new_[4739]_ , \new_[4740]_ ,
    \new_[4741]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4746]_ , \new_[4747]_ , \new_[4828]_ ,
    \new_[4829]_ , \new_[4830]_ , \new_[4831]_ , \new_[4832]_ ,
    \new_[4833]_ , \new_[4834]_ , \new_[4835]_ , \new_[4836]_ ,
    \new_[4837]_ , \new_[4838]_ , \new_[4839]_ , \new_[4840]_ ,
    \new_[4841]_ , \new_[4842]_ , \new_[4843]_ , \new_[4844]_ ,
    \new_[4845]_ , \new_[4846]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4850]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4853]_ , \new_[4854]_ , \new_[4855]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4858]_ , \new_[4859]_ , \new_[4860]_ ,
    \new_[4861]_ , \new_[4862]_ , \new_[4863]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4869]_ , \new_[4870]_ , \new_[4871]_ , \new_[4872]_ ,
    \new_[4873]_ , \new_[4874]_ , \new_[4875]_ , \new_[4876]_ ,
    \new_[4877]_ , \new_[4878]_ , \new_[4879]_ , \new_[4880]_ ,
    \new_[4881]_ , \new_[4882]_ , \new_[4883]_ , \new_[4884]_ ,
    \new_[4885]_ , \new_[4886]_ , \new_[4887]_ , \new_[4888]_ ,
    \new_[4889]_ , \new_[4890]_ , \new_[4891]_ , \new_[4892]_ ,
    \new_[4893]_ , \new_[4894]_ , \new_[4895]_ , \new_[4896]_ ,
    \new_[4897]_ , \new_[4898]_ , \new_[4899]_ , \new_[4900]_ ,
    \new_[4901]_ , \new_[4918]_ , \new_[4919]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4923]_ , \new_[4924]_ ,
    \new_[4925]_ , \new_[4926]_ , \new_[4927]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4933]_ , \new_[4934]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4940]_ ,
    \new_[4941]_ , \new_[4942]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4947]_ , \new_[4948]_ ,
    \new_[4949]_ , \new_[4950]_ , \new_[4951]_ , \new_[4952]_ ,
    \new_[4953]_ , \new_[4954]_ , \new_[4955]_ , \new_[4956]_ ,
    \new_[4957]_ , \new_[4958]_ , \new_[4959]_ , \new_[4960]_ ,
    \new_[4961]_ , \new_[4962]_ , \new_[4963]_ , \new_[4964]_ ,
    \new_[4965]_ , \new_[4966]_ , \new_[4967]_ , \new_[4968]_ ,
    \new_[4969]_ , \new_[4970]_ , \new_[4971]_ , \new_[4972]_ ,
    \new_[4973]_ , \new_[4974]_ , \new_[4975]_ , \new_[4976]_ ,
    \new_[4977]_ , \new_[4978]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4981]_ , \new_[4982]_ , \new_[4983]_ , \new_[4984]_ ,
    \new_[4985]_ , \new_[4986]_ , \new_[4987]_ , \new_[4988]_ ,
    \new_[4989]_ , \new_[4990]_ , \new_[4991]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4994]_ , \new_[4995]_ , \new_[4996]_ ,
    \new_[4997]_ , \new_[4998]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5003]_ , \new_[5004]_ ,
    \new_[5005]_ , \new_[5006]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5010]_ , \new_[5011]_ , \new_[5012]_ ,
    \new_[5013]_ , \new_[5014]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5017]_ , \new_[5018]_ , \new_[5019]_ , \new_[5020]_ ,
    \new_[5021]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5027]_ , \new_[5028]_ ,
    \new_[5029]_ , \new_[5030]_ , \new_[5031]_ , \new_[5032]_ ,
    \new_[5033]_ , \new_[5034]_ , \new_[5035]_ , \new_[5036]_ ,
    \new_[5037]_ , \new_[5038]_ , \new_[5039]_ , \new_[5040]_ ,
    \new_[5041]_ , \new_[5042]_ , \new_[5043]_ , \new_[5044]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5048]_ ,
    \new_[5049]_ , \new_[5050]_ , \new_[5051]_ , \new_[5052]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5055]_ , \new_[5056]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5067]_ , \new_[5068]_ ,
    \new_[5069]_ , \new_[5070]_ , \new_[5071]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5075]_ , \new_[5076]_ ,
    \new_[5077]_ , \new_[5080]_ , \new_[5081]_ , \new_[5082]_ ,
    \new_[5083]_ , \new_[5084]_ , \new_[5085]_ , \new_[5086]_ ,
    \new_[5087]_ , \new_[5088]_ , \new_[5089]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5093]_ , \new_[5094]_ ,
    \new_[5095]_ , \new_[5096]_ , \new_[5097]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5101]_ , \new_[5102]_ ,
    \new_[5103]_ , \new_[5104]_ , \new_[5105]_ , \new_[5106]_ ,
    \new_[5107]_ , \new_[5108]_ , \new_[5109]_ , \new_[5110]_ ,
    \new_[5111]_ , \new_[5112]_ , \new_[5113]_ , \new_[5114]_ ,
    \new_[5115]_ , \new_[5116]_ , \new_[5117]_ , \new_[5118]_ ,
    \new_[5119]_ , \new_[5120]_ , \new_[5121]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5126]_ ,
    \new_[5127]_ , \new_[5128]_ , \new_[5129]_ , \new_[5130]_ ,
    \new_[5131]_ , \new_[5132]_ , \new_[5133]_ , \new_[5134]_ ,
    \new_[5135]_ , \new_[5136]_ , \new_[5137]_ , \new_[5138]_ ,
    \new_[5139]_ , \new_[5140]_ , \new_[5141]_ , \new_[5142]_ ,
    \new_[5143]_ , \new_[5144]_ , \new_[5145]_ , \new_[5146]_ ,
    \new_[5147]_ , \new_[5148]_ , \new_[5149]_ , \new_[5150]_ ,
    \new_[5151]_ , \new_[5152]_ , \new_[5153]_ , \new_[5154]_ ,
    \new_[5155]_ , \new_[5156]_ , \new_[5157]_ , \new_[5158]_ ,
    \new_[5159]_ , \new_[5160]_ , \new_[5161]_ , \new_[5162]_ ,
    \new_[5163]_ , \new_[5164]_ , \new_[5165]_ , \new_[5166]_ ,
    \new_[5167]_ , \new_[5168]_ , \new_[5169]_ , \new_[5170]_ ,
    \new_[5171]_ , \new_[5172]_ , \new_[5173]_ , \new_[5174]_ ,
    \new_[5175]_ , \new_[5176]_ , \new_[5177]_ , \new_[5178]_ ,
    \new_[5179]_ , \new_[5180]_ , \new_[5181]_ , \new_[5182]_ ,
    \new_[5183]_ , \new_[5184]_ , \new_[5185]_ , \new_[5186]_ ,
    \new_[5187]_ , \new_[5188]_ , \new_[5189]_ , \new_[5190]_ ,
    \new_[5191]_ , \new_[5192]_ , \new_[5193]_ , \new_[5194]_ ,
    \new_[5195]_ , \new_[5196]_ , \new_[5197]_ , \new_[5198]_ ,
    \new_[5199]_ , \new_[5200]_ , \new_[5201]_ , \new_[5202]_ ,
    \new_[5203]_ , \new_[5204]_ , \new_[5205]_ , \new_[5206]_ ,
    \new_[5207]_ , \new_[5208]_ , \new_[5209]_ , \new_[5210]_ ,
    \new_[5211]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5215]_ , \new_[5216]_ , \new_[5217]_ , \new_[5218]_ ,
    \new_[5219]_ , \new_[5220]_ , \new_[5221]_ , \new_[5222]_ ,
    \new_[5223]_ , \new_[5224]_ , \new_[5225]_ , \new_[5226]_ ,
    \new_[5227]_ , \new_[5228]_ , \new_[5229]_ , \new_[5230]_ ,
    \new_[5231]_ , \new_[5232]_ , \new_[5233]_ , \new_[5234]_ ,
    \new_[5235]_ , \new_[5236]_ , \new_[5237]_ , \new_[5238]_ ,
    \new_[5239]_ , \new_[5240]_ , \new_[5241]_ , \new_[5242]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5245]_ , \new_[5246]_ ,
    \new_[5247]_ , \new_[5248]_ , \new_[5249]_ , \new_[5250]_ ,
    \new_[5251]_ , \new_[5252]_ , \new_[5253]_ , \new_[5254]_ ,
    \new_[5255]_ , \new_[5256]_ , \new_[5257]_ , \new_[5258]_ ,
    \new_[5259]_ , \new_[5260]_ , \new_[5261]_ , \new_[5262]_ ,
    \new_[5263]_ , \new_[5264]_ , \new_[5265]_ , \new_[5266]_ ,
    \new_[5267]_ , \new_[5268]_ , \new_[5269]_ , \new_[5270]_ ,
    \new_[5271]_ , \new_[5272]_ , \new_[5273]_ , \new_[5274]_ ,
    \new_[5275]_ , \new_[5276]_ , \new_[5277]_ , \new_[5278]_ ,
    \new_[5279]_ , \new_[5280]_ , \new_[5281]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5285]_ , \new_[5286]_ ,
    \new_[5287]_ , \new_[5288]_ , \new_[5289]_ , \new_[5290]_ ,
    \new_[5291]_ , \new_[5292]_ , \new_[5293]_ , \new_[5294]_ ,
    \new_[5295]_ , \new_[5296]_ , \new_[5297]_ , \new_[5298]_ ,
    \new_[5299]_ , \new_[5300]_ , \new_[5301]_ , \new_[5302]_ ,
    \new_[5303]_ , \new_[5304]_ , \new_[5305]_ , \new_[5306]_ ,
    \new_[5307]_ , \new_[5308]_ , \new_[5309]_ , \new_[5310]_ ,
    \new_[5311]_ , \new_[5312]_ , \new_[5313]_ , \new_[5314]_ ,
    \new_[5315]_ , \new_[5316]_ , \new_[5317]_ , \new_[5318]_ ,
    \new_[5319]_ , \new_[5320]_ , \new_[5321]_ , \new_[5322]_ ,
    \new_[5323]_ , \new_[5324]_ , \new_[5325]_ , \new_[5326]_ ,
    \new_[5327]_ , \new_[5328]_ , \new_[5329]_ , \new_[5330]_ ,
    \new_[5331]_ , \new_[5332]_ , \new_[5333]_ , \new_[5334]_ ,
    \new_[5335]_ , \new_[5336]_ , \new_[5337]_ , \new_[5338]_ ,
    \new_[5339]_ , \new_[5340]_ , \new_[5341]_ , \new_[5342]_ ,
    \new_[5343]_ , \new_[5344]_ , \new_[5345]_ , \new_[5346]_ ,
    \new_[5347]_ , \new_[5348]_ , \new_[5349]_ , \new_[5350]_ ,
    \new_[5351]_ , \new_[5352]_ , \new_[5353]_ , \new_[5354]_ ,
    \new_[5355]_ , \new_[5356]_ , \new_[5357]_ , \new_[5358]_ ,
    \new_[5359]_ , \new_[5360]_ , \new_[5361]_ , \new_[5362]_ ,
    \new_[5363]_ , \new_[5364]_ , \new_[5365]_ , \new_[5366]_ ,
    \new_[5367]_ , \new_[5368]_ , \new_[5369]_ , \new_[5370]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5373]_ , \new_[5374]_ ,
    \new_[5375]_ , \new_[5376]_ , \new_[5377]_ , \new_[5378]_ ,
    \new_[5379]_ , \new_[5380]_ , \new_[5381]_ , \new_[5382]_ ,
    \new_[5383]_ , \new_[5384]_ , \new_[5385]_ , \new_[5386]_ ,
    \new_[5387]_ , \new_[5388]_ , \new_[5389]_ , \new_[5390]_ ,
    \new_[5391]_ , \new_[5392]_ , \new_[5393]_ , \new_[5394]_ ,
    \new_[5395]_ , \new_[5396]_ , \new_[5397]_ , \new_[5398]_ ,
    \new_[5399]_ , \new_[5400]_ , \new_[5401]_ , \new_[5402]_ ,
    \new_[5403]_ , \new_[5404]_ , \new_[5405]_ , \new_[5406]_ ,
    \new_[5407]_ , \new_[5408]_ , \new_[5409]_ , \new_[5410]_ ,
    \new_[5411]_ , \new_[5412]_ , \new_[5413]_ , \new_[5414]_ ,
    \new_[5415]_ , \new_[5416]_ , \new_[5417]_ , \new_[5418]_ ,
    \new_[5419]_ , \new_[5420]_ , \new_[5421]_ , \new_[5422]_ ,
    \new_[5423]_ , \new_[5424]_ , \new_[5425]_ , \new_[5426]_ ,
    \new_[5427]_ , \new_[5428]_ , \new_[5429]_ , \new_[5430]_ ,
    \new_[5431]_ , \new_[5432]_ , \new_[5433]_ , \new_[5434]_ ,
    \new_[5435]_ , \new_[5436]_ , \new_[5437]_ , \new_[5438]_ ,
    \new_[5439]_ , \new_[5440]_ , \new_[5441]_ , \new_[5442]_ ,
    \new_[5443]_ , \new_[5444]_ , \new_[5445]_ , \new_[5446]_ ,
    \new_[5447]_ , \new_[5448]_ , \new_[5449]_ , \new_[5450]_ ,
    \new_[5451]_ , \new_[5452]_ , \new_[5453]_ , \new_[5454]_ ,
    \new_[5455]_ , \new_[5456]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5459]_ , \new_[5460]_ , \new_[5461]_ , \new_[5462]_ ,
    \new_[5463]_ , \new_[5464]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5468]_ , \new_[5469]_ , \new_[5470]_ ,
    \new_[5471]_ , \new_[5472]_ , \new_[5473]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5476]_ , \new_[5477]_ , \new_[5478]_ ,
    \new_[5479]_ , \new_[5480]_ , \new_[5481]_ , \new_[5482]_ ,
    \new_[5483]_ , \new_[5484]_ , \new_[5485]_ , \new_[5486]_ ,
    \new_[5487]_ , \new_[5488]_ , \new_[5489]_ , \new_[5490]_ ,
    \new_[5491]_ , \new_[5492]_ , \new_[5493]_ , \new_[5494]_ ,
    \new_[5495]_ , \new_[5496]_ , \new_[5497]_ , \new_[5498]_ ,
    \new_[5499]_ , \new_[5500]_ , \new_[5501]_ , \new_[5502]_ ,
    \new_[5503]_ , \new_[5504]_ , \new_[5505]_ , \new_[5506]_ ,
    \new_[5507]_ , \new_[5508]_ , \new_[5509]_ , \new_[5510]_ ,
    \new_[5511]_ , \new_[5512]_ , \new_[5513]_ , \new_[5514]_ ,
    \new_[5515]_ , \new_[5516]_ , \new_[5517]_ , \new_[5518]_ ,
    \new_[5519]_ , \new_[5520]_ , \new_[5521]_ , \new_[5522]_ ,
    \new_[5523]_ , \new_[5524]_ , \new_[5525]_ , \new_[5526]_ ,
    \new_[5527]_ , \new_[5528]_ , \new_[5529]_ , \new_[5530]_ ,
    \new_[5531]_ , \new_[5532]_ , \new_[5533]_ , \new_[5534]_ ,
    \new_[5535]_ , \new_[5536]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5541]_ , \new_[5542]_ ,
    \new_[5543]_ , \new_[5544]_ , \new_[5545]_ , \new_[5546]_ ,
    \new_[5547]_ , \new_[5548]_ , \new_[5549]_ , \new_[5550]_ ,
    \new_[5551]_ , \new_[5552]_ , \new_[5553]_ , \new_[5554]_ ,
    \new_[5555]_ , \new_[5556]_ , \new_[5557]_ , \new_[5558]_ ,
    \new_[5559]_ , \new_[5560]_ , \new_[5561]_ , \new_[5562]_ ,
    \new_[5563]_ , \new_[5564]_ , \new_[5565]_ , \new_[5566]_ ,
    \new_[5567]_ , \new_[5568]_ , \new_[5569]_ , \new_[5570]_ ,
    \new_[5571]_ , \new_[5572]_ , \new_[5573]_ , \new_[5574]_ ,
    \new_[5575]_ , \new_[5576]_ , \new_[5577]_ , \new_[5578]_ ,
    \new_[5579]_ , \new_[5580]_ , \new_[5581]_ , \new_[5582]_ ,
    \new_[5583]_ , \new_[5584]_ , \new_[5585]_ , \new_[5586]_ ,
    \new_[5587]_ , \new_[5588]_ , \new_[5589]_ , \new_[5590]_ ,
    \new_[5591]_ , \new_[5592]_ , \new_[5593]_ , \new_[5594]_ ,
    \new_[5595]_ , \new_[5596]_ , \new_[5597]_ , \new_[5598]_ ,
    \new_[5599]_ , \new_[5600]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5605]_ , \new_[5606]_ ,
    \new_[5607]_ , \new_[5608]_ , \new_[5609]_ , \new_[5610]_ ,
    \new_[5611]_ , \new_[5612]_ , \new_[5613]_ , \new_[5614]_ ,
    \new_[5615]_ , \new_[5616]_ , \new_[5617]_ , \new_[5618]_ ,
    \new_[5619]_ , \new_[5620]_ , \new_[5621]_ , \new_[5622]_ ,
    \new_[5623]_ , \new_[5624]_ , \new_[5625]_ , \new_[5626]_ ,
    \new_[5627]_ , \new_[5628]_ , \new_[5629]_ , \new_[5630]_ ,
    \new_[5631]_ , \new_[5632]_ , \new_[5633]_ , \new_[5634]_ ,
    \new_[5635]_ , \new_[5636]_ , \new_[5637]_ , \new_[5638]_ ,
    \new_[5639]_ , \new_[5640]_ , \new_[5641]_ , \new_[5642]_ ,
    \new_[5643]_ , \new_[5644]_ , \new_[5645]_ , \new_[5646]_ ,
    \new_[5647]_ , \new_[5648]_ , \new_[5649]_ , \new_[5650]_ ,
    \new_[5651]_ , \new_[5652]_ , \new_[5653]_ , \new_[5654]_ ,
    \new_[5655]_ , \new_[5656]_ , \new_[5657]_ , \new_[5658]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5661]_ , \new_[5662]_ ,
    \new_[5663]_ , \new_[5664]_ , \new_[5665]_ , \new_[5666]_ ,
    \new_[5667]_ , \new_[5668]_ , \new_[5669]_ , \new_[5670]_ ,
    \new_[5671]_ , \new_[5672]_ , \new_[5673]_ , \new_[5674]_ ,
    \new_[5675]_ , \new_[5676]_ , \new_[5677]_ , \new_[5678]_ ,
    \new_[5679]_ , \new_[5680]_ , \new_[5681]_ , \new_[5682]_ ,
    \new_[5683]_ , \new_[5684]_ , \new_[5685]_ , \new_[5686]_ ,
    \new_[5687]_ , \new_[5688]_ , \new_[5689]_ , \new_[5690]_ ,
    \new_[5691]_ , \new_[5692]_ , \new_[5693]_ , \new_[5694]_ ,
    \new_[5695]_ , \new_[5696]_ , \new_[5697]_ , \new_[5698]_ ,
    \new_[5699]_ , \new_[5700]_ , \new_[5701]_ , \new_[5702]_ ,
    \new_[5703]_ , \new_[5704]_ , \new_[5705]_ , \new_[5706]_ ,
    \new_[5707]_ , \new_[5708]_ , \new_[5709]_ , \new_[5710]_ ,
    \new_[5711]_ , \new_[5712]_ , \new_[5713]_ , \new_[5714]_ ,
    \new_[5715]_ , \new_[5716]_ , \new_[5717]_ , \new_[5718]_ ,
    \new_[5719]_ , \new_[5720]_ , \new_[5721]_ , \new_[5722]_ ,
    \new_[5723]_ , \new_[5724]_ , \new_[5725]_ , \new_[5726]_ ,
    \new_[5727]_ , \new_[5728]_ , \new_[5729]_ , \new_[5730]_ ,
    \new_[5731]_ , \new_[5732]_ , \new_[5733]_ , \new_[5734]_ ,
    \new_[5735]_ , \new_[5736]_ , \new_[5737]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5740]_ , \new_[5741]_ , \new_[5742]_ ,
    \new_[5743]_ , \new_[5744]_ , \new_[5745]_ , \new_[5746]_ ,
    \new_[5747]_ , \new_[5748]_ , \new_[5749]_ , \new_[5750]_ ,
    \new_[5751]_ , \new_[5752]_ , \new_[5753]_ , \new_[5754]_ ,
    \new_[5755]_ , \new_[5756]_ , \new_[5757]_ , \new_[5758]_ ,
    \new_[5759]_ , \new_[5760]_ , \new_[5761]_ , \new_[5762]_ ,
    \new_[5763]_ , \new_[5764]_ , \new_[5765]_ , \new_[5766]_ ,
    \new_[5767]_ , \new_[5768]_ , \new_[5769]_ , \new_[5770]_ ,
    \new_[5771]_ , \new_[5772]_ , \new_[5773]_ , \new_[5774]_ ,
    \new_[5775]_ , \new_[5776]_ , \new_[5777]_ , \new_[5778]_ ,
    \new_[5779]_ , \new_[5780]_ , \new_[5781]_ , \new_[5782]_ ,
    \new_[5783]_ , \new_[5784]_ , \new_[5785]_ , \new_[5786]_ ,
    \new_[5787]_ , \new_[5788]_ , \new_[5789]_ , \new_[5790]_ ,
    \new_[5791]_ , \new_[5792]_ , \new_[5793]_ , \new_[5794]_ ,
    \new_[5795]_ , \new_[5796]_ , \new_[5797]_ , \new_[5798]_ ,
    \new_[5799]_ , \new_[5800]_ , \new_[5801]_ , \new_[5802]_ ,
    \new_[5803]_ , \new_[5804]_ , \new_[5805]_ , \new_[5806]_ ,
    \new_[5807]_ , \new_[5808]_ , \new_[5809]_ , \new_[5810]_ ,
    \new_[5811]_ , \new_[5812]_ , \new_[5813]_ , \new_[5814]_ ,
    \new_[5815]_ , \new_[5816]_ , \new_[5817]_ , \new_[5818]_ ,
    \new_[5819]_ , \new_[5820]_ , \new_[5821]_ , \new_[5822]_ ,
    \new_[5823]_ , \new_[5824]_ , \new_[5825]_ , \new_[5826]_ ,
    \new_[5827]_ , \new_[5828]_ , \new_[5829]_ , \new_[5830]_ ,
    \new_[5831]_ , \new_[5832]_ , \new_[5833]_ , \new_[5834]_ ,
    \new_[5835]_ , \new_[5836]_ , \new_[5837]_ , \new_[5838]_ ,
    \new_[5839]_ , \new_[5840]_ , \new_[5841]_ , \new_[5842]_ ,
    \new_[5843]_ , \new_[5844]_ , \new_[5845]_ , \new_[5846]_ ,
    \new_[5847]_ , \new_[5848]_ , \new_[5849]_ , \new_[5850]_ ,
    \new_[5851]_ , \new_[5852]_ , \new_[5853]_ , \new_[5854]_ ,
    \new_[5855]_ , \new_[5856]_ , \new_[5857]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5861]_ , \new_[5862]_ ,
    \new_[5863]_ , \new_[5864]_ , \new_[5865]_ , \new_[5866]_ ,
    \new_[5867]_ , \new_[5868]_ , \new_[5869]_ , \new_[5870]_ ,
    \new_[5871]_ , \new_[5872]_ , \new_[5873]_ , \new_[5874]_ ,
    \new_[5875]_ , \new_[5876]_ , \new_[5877]_ , \new_[5878]_ ,
    \new_[5879]_ , \new_[5880]_ , \new_[5881]_ , \new_[5882]_ ,
    \new_[5883]_ , \new_[5884]_ , \new_[5885]_ , \new_[5886]_ ,
    \new_[5887]_ , \new_[5888]_ , \new_[5889]_ , \new_[5890]_ ,
    \new_[5891]_ , \new_[5892]_ , \new_[5893]_ , \new_[5894]_ ,
    \new_[5895]_ , \new_[5896]_ , \new_[5897]_ , \new_[5898]_ ,
    \new_[5899]_ , \new_[5900]_ , \new_[5901]_ , \new_[5902]_ ,
    \new_[5903]_ , \new_[5904]_ , \new_[5905]_ , \new_[5906]_ ,
    \new_[5907]_ , \new_[5908]_ , \new_[5909]_ , \new_[5910]_ ,
    \new_[5911]_ , \new_[5912]_ , \new_[5913]_ , \new_[5914]_ ,
    \new_[5915]_ , \new_[5916]_ , \new_[5917]_ , \new_[5918]_ ,
    \new_[5919]_ , \new_[5920]_ , \new_[5921]_ , \new_[5922]_ ,
    \new_[5923]_ , \new_[5924]_ , \new_[5925]_ , \new_[5926]_ ,
    \new_[5927]_ , \new_[5928]_ , \new_[5929]_ , \new_[5930]_ ,
    \new_[5931]_ , \new_[5932]_ , \new_[5933]_ , \new_[5934]_ ,
    \new_[5935]_ , \new_[5936]_ , \new_[5937]_ , \new_[5938]_ ,
    \new_[5939]_ , \new_[5940]_ , \new_[5941]_ , \new_[5942]_ ,
    \new_[5943]_ , \new_[5944]_ , \new_[5945]_ , \new_[5946]_ ,
    \new_[5947]_ , \new_[5948]_ , \new_[5949]_ , \new_[5950]_ ,
    \new_[5951]_ , \new_[5952]_ , \new_[5953]_ , \new_[5954]_ ,
    \new_[5955]_ , \new_[5956]_ , \new_[5957]_ , \new_[5958]_ ,
    \new_[5959]_ , \new_[5960]_ , \new_[5961]_ , \new_[5962]_ ,
    \new_[5963]_ , \new_[5964]_ , \new_[5965]_ , \new_[5966]_ ,
    \new_[5967]_ , \new_[5968]_ , \new_[5969]_ , \new_[5970]_ ,
    \new_[5971]_ , \new_[5972]_ , \new_[5973]_ , \new_[5974]_ ,
    \new_[5975]_ , \new_[5976]_ , \new_[5977]_ , \new_[5978]_ ,
    \new_[5979]_ , \new_[5980]_ , \new_[5981]_ , \new_[5982]_ ,
    \new_[5983]_ , \new_[5984]_ , \new_[5985]_ , \new_[5986]_ ,
    \new_[5987]_ , \new_[5988]_ , \new_[5989]_ , \new_[5990]_ ,
    \new_[5991]_ , \new_[5992]_ , \new_[5993]_ , \new_[5994]_ ,
    \new_[5995]_ , \new_[5996]_ , \new_[5997]_ , \new_[5998]_ ,
    \new_[5999]_ , \new_[6000]_ , \new_[6001]_ , \new_[6002]_ ,
    \new_[6003]_ , \new_[6004]_ , \new_[6005]_ , \new_[6006]_ ,
    \new_[6007]_ , \new_[6009]_ , \new_[6010]_ , \new_[6011]_ ,
    \new_[6012]_ , \new_[6013]_ , \new_[6014]_ , \new_[6015]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6022]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6028]_ , \new_[6029]_ , \new_[6030]_ , \new_[6031]_ ,
    \new_[6032]_ , \new_[6033]_ , \new_[6034]_ , \new_[6035]_ ,
    \new_[6036]_ , \new_[6037]_ , \new_[6038]_ , \new_[6039]_ ,
    \new_[6040]_ , \new_[6041]_ , \new_[6042]_ , \new_[6043]_ ,
    \new_[6044]_ , \new_[6045]_ , \new_[6046]_ , \new_[6047]_ ,
    \new_[6048]_ , \new_[6049]_ , \new_[6050]_ , \new_[6051]_ ,
    \new_[6052]_ , \new_[6053]_ , \new_[6054]_ , \new_[6055]_ ,
    \new_[6056]_ , \new_[6057]_ , \new_[6058]_ , \new_[6059]_ ,
    \new_[6060]_ , \new_[6061]_ , \new_[6062]_ , \new_[6063]_ ,
    \new_[6064]_ , \new_[6065]_ , \new_[6066]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6069]_ , \new_[6070]_ , \new_[6071]_ ,
    \new_[6072]_ , \new_[6073]_ , \new_[6074]_ , \new_[6075]_ ,
    \new_[6076]_ , \new_[6077]_ , \new_[6078]_ , \new_[6079]_ ,
    \new_[6080]_ , \new_[6081]_ , \new_[6082]_ , \new_[6083]_ ,
    \new_[6084]_ , \new_[6085]_ , \new_[6086]_ , \new_[6087]_ ,
    \new_[6088]_ , \new_[6089]_ , \new_[6090]_ , \new_[6091]_ ,
    \new_[6092]_ , \new_[6093]_ , \new_[6094]_ , \new_[6095]_ ,
    \new_[6096]_ , \new_[6174]_ , \new_[6176]_ , \new_[6183]_ ,
    \new_[6184]_ , \new_[6185]_ , \new_[6186]_ , \new_[6187]_ ,
    \new_[6188]_ , \new_[6189]_ , \new_[6190]_ , \new_[6191]_ ,
    \new_[6192]_ , \new_[6193]_ , \new_[6194]_ , \new_[6195]_ ,
    \new_[6196]_ , \new_[6197]_ , \new_[6198]_ , \new_[6199]_ ,
    \new_[6200]_ , \new_[6201]_ , \new_[6202]_ , \new_[6203]_ ,
    \new_[6204]_ , \new_[6205]_ , \new_[6206]_ , \new_[6207]_ ,
    \new_[6208]_ , \new_[6209]_ , \new_[6210]_ , \new_[6211]_ ,
    \new_[6212]_ , \new_[6213]_ , \new_[6214]_ , \new_[6215]_ ,
    \new_[6216]_ , \new_[6217]_ , \new_[6221]_ , \new_[6222]_ ,
    \new_[6223]_ , \new_[6245]_ , \new_[6246]_ , \new_[6268]_ ,
    \new_[6269]_ , \new_[6270]_ , \new_[6271]_ , \new_[6272]_ ,
    \new_[6273]_ , \new_[6274]_ , \new_[6287]_ , \new_[6357]_ ,
    \new_[6358]_ , \new_[6359]_ , \new_[6360]_ , \new_[6361]_ ,
    \new_[6362]_ , \new_[6363]_ , \new_[6364]_ , \new_[6365]_ ,
    \new_[6366]_ , \new_[6367]_ , \new_[6368]_ , \new_[6369]_ ,
    \new_[6370]_ , \new_[6371]_ , \new_[6372]_ , \new_[6373]_ ,
    \new_[6374]_ , \new_[6375]_ , \new_[6376]_ , \new_[6389]_ ,
    \new_[6390]_ , \new_[6391]_ , \new_[6425]_ , \new_[6426]_ ,
    \new_[6427]_ , \new_[6428]_ , \new_[6429]_ , \new_[6430]_ ,
    \new_[6431]_ , \new_[6432]_ , \new_[6433]_ , \new_[6434]_ ,
    \new_[6435]_ , \new_[6436]_ , \new_[6437]_ , \new_[6438]_ ,
    \new_[6439]_ , \new_[6440]_ , \new_[6441]_ , \new_[6442]_ ,
    \new_[6443]_ , \new_[6444]_ , \new_[6445]_ , \new_[6446]_ ,
    \new_[6447]_ , \new_[6448]_ , \new_[6449]_ , \new_[6578]_ ,
    \new_[6584]_ , \new_[6585]_ , \new_[6586]_ , \new_[6587]_ ,
    \new_[6588]_ , \new_[6589]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6592]_ , \new_[6593]_ , \new_[6594]_ , \new_[6595]_ ,
    \new_[6596]_ , \new_[6597]_ , \new_[6598]_ , \new_[6599]_ ,
    \new_[6600]_ , \new_[6601]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6608]_ , \new_[6609]_ , \new_[6610]_ , \new_[6611]_ ,
    \new_[6612]_ , \new_[6613]_ , \new_[6614]_ , \new_[6615]_ ,
    \new_[6616]_ , \new_[6617]_ , \new_[6618]_ , \new_[6619]_ ,
    \new_[6620]_ , \new_[6621]_ , \new_[6622]_ , \new_[6623]_ ,
    \new_[6624]_ , \new_[6625]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6628]_ , \new_[6629]_ , \new_[6630]_ , \new_[6631]_ ,
    \new_[6632]_ , \new_[6633]_ , \new_[6634]_ , \new_[6635]_ ,
    \new_[6636]_ , \new_[6637]_ , \new_[6638]_ , \new_[6639]_ ,
    \new_[6640]_ , \new_[6641]_ , \new_[6642]_ , \new_[6643]_ ,
    \new_[6644]_ , \new_[6645]_ , \new_[6646]_ , \new_[6647]_ ,
    \new_[6648]_ , \new_[6649]_ , \new_[6650]_ , \new_[6651]_ ,
    \new_[6652]_ , \new_[6653]_ , \new_[6654]_ , \new_[6655]_ ,
    \new_[6656]_ , \new_[6657]_ , \new_[6658]_ , \new_[6659]_ ,
    \new_[6660]_ , \new_[6661]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6664]_ , \new_[6665]_ , \new_[6666]_ , \new_[6667]_ ,
    \new_[6668]_ , \new_[6669]_ , \new_[6670]_ , \new_[6671]_ ,
    \new_[6672]_ , \new_[6673]_ , \new_[6674]_ , \new_[6675]_ ,
    \new_[6676]_ , \new_[6677]_ , \new_[6678]_ , \new_[6679]_ ,
    \new_[6680]_ , \new_[6681]_ , \new_[6682]_ , \new_[6683]_ ,
    \new_[6684]_ , \new_[6685]_ , \new_[6686]_ , \new_[6687]_ ,
    \new_[6688]_ , \new_[6689]_ , \new_[6690]_ , \new_[6691]_ ,
    \new_[6692]_ , \new_[6693]_ , \new_[6694]_ , \new_[6695]_ ,
    \new_[6696]_ , \new_[6697]_ , \new_[6698]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6701]_ , \new_[6702]_ , \new_[6703]_ ,
    \new_[6704]_ , \new_[6705]_ , \new_[6706]_ , \new_[6707]_ ,
    \new_[6708]_ , \new_[6709]_ , \new_[6710]_ , \new_[6711]_ ,
    \new_[6712]_ , \new_[6713]_ , \new_[6714]_ , \new_[6715]_ ,
    \new_[6716]_ , \new_[6717]_ , \new_[6718]_ , \new_[6719]_ ,
    \new_[6720]_ , \new_[6721]_ , \new_[6722]_ , \new_[6723]_ ,
    \new_[6724]_ , \new_[6725]_ , \new_[6726]_ , \new_[6727]_ ,
    \new_[6728]_ , \new_[6729]_ , \new_[6730]_ , \new_[6731]_ ,
    \new_[6732]_ , \new_[6733]_ , \new_[6734]_ , \new_[6735]_ ,
    \new_[6736]_ , \new_[6737]_ , \new_[6738]_ , \new_[6739]_ ,
    \new_[6740]_ , \new_[6741]_ , \new_[6742]_ , \new_[6743]_ ,
    \new_[6744]_ , \new_[6745]_ , \new_[6746]_ , \new_[6747]_ ,
    \new_[6748]_ , \new_[6749]_ , \new_[6750]_ , \new_[6751]_ ,
    \new_[6752]_ , \new_[6753]_ , \new_[6754]_ , \new_[6755]_ ,
    \new_[6756]_ , \new_[6757]_ , \new_[6758]_ , \new_[6759]_ ,
    \new_[6760]_ , \new_[6761]_ , \new_[6762]_ , \new_[6763]_ ,
    \new_[6764]_ , \new_[6765]_ , \new_[6766]_ , \new_[6767]_ ,
    \new_[6768]_ , \new_[6769]_ , \new_[6770]_ , \new_[6771]_ ,
    \new_[6772]_ , \new_[6773]_ , \new_[6774]_ , \new_[6775]_ ,
    \new_[6776]_ , \new_[6777]_ , \new_[6778]_ , \new_[6779]_ ,
    \new_[6780]_ , \new_[6781]_ , \new_[6782]_ , \new_[6783]_ ,
    \new_[6784]_ , \new_[6785]_ , \new_[6786]_ , \new_[6787]_ ,
    \new_[6788]_ , \new_[6789]_ , \new_[6790]_ , \new_[6791]_ ,
    \new_[6792]_ , \new_[6793]_ , \new_[6794]_ , \new_[7205]_ ,
    \new_[7215]_ , \new_[7216]_ , \new_[7218]_ , \new_[7220]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7224]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7230]_ , \new_[7231]_ ,
    \new_[7232]_ , \new_[7233]_ , \new_[7234]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7244]_ , \new_[7245]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7248]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7255]_ ,
    \new_[7256]_ , \new_[7257]_ , \new_[7258]_ , \new_[7259]_ ,
    \new_[7260]_ , \new_[7261]_ , \new_[7262]_ , \new_[7263]_ ,
    \new_[7264]_ , \new_[7265]_ , \new_[7266]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7270]_ , \new_[7271]_ ,
    \new_[7272]_ , \new_[7273]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7276]_ , \new_[7277]_ , \new_[7278]_ , \new_[7279]_ ,
    \new_[7280]_ , \new_[7281]_ , \new_[7282]_ , \new_[7283]_ ,
    \new_[7284]_ , \new_[7285]_ , \new_[7286]_ , \new_[7287]_ ,
    \new_[7288]_ , \new_[7289]_ , \new_[7290]_ , \new_[7291]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7294]_ , \new_[7295]_ ,
    \new_[7296]_ , \new_[7297]_ , \new_[7298]_ , \new_[7299]_ ,
    \new_[7300]_ , \new_[7301]_ , \new_[7302]_ , \new_[7303]_ ,
    \new_[7304]_ , \new_[7305]_ , \new_[7306]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7312]_ , \new_[7313]_ , \new_[7314]_ , \new_[7315]_ ,
    \new_[7316]_ , \new_[7317]_ , \new_[7318]_ , \new_[7319]_ ,
    \new_[7320]_ , \new_[7321]_ , \new_[7322]_ , \new_[7323]_ ,
    \new_[7324]_ , \new_[7325]_ , \new_[7326]_ , \new_[7327]_ ,
    \new_[7328]_ , \new_[7329]_ , \new_[7330]_ , \new_[7331]_ ,
    \new_[7332]_ , \new_[7333]_ , \new_[7334]_ , \new_[7335]_ ,
    \new_[7336]_ , \new_[7337]_ , \new_[7338]_ , \new_[7339]_ ,
    \new_[7340]_ , \new_[7341]_ , \new_[7342]_ , \new_[7343]_ ,
    \new_[7344]_ , \new_[7345]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7348]_ , \new_[7349]_ , \new_[7350]_ , \new_[7351]_ ,
    \new_[7352]_ , \new_[7353]_ , \new_[7354]_ , \new_[7355]_ ,
    \new_[7356]_ , \new_[7357]_ , \new_[7358]_ , \new_[7359]_ ,
    \new_[7360]_ , \new_[7361]_ , \new_[7362]_ , \new_[7363]_ ,
    \new_[7364]_ , \new_[7365]_ , \new_[7366]_ , \new_[7367]_ ,
    \new_[7368]_ , \new_[7369]_ , \new_[7370]_ , \new_[7371]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7374]_ , \new_[7375]_ ,
    \new_[7376]_ , \new_[7377]_ , \new_[7378]_ , \new_[7379]_ ,
    \new_[7380]_ , \new_[7381]_ , \new_[7382]_ , \new_[7383]_ ,
    \new_[7384]_ , \new_[7385]_ , \new_[7386]_ , \new_[7387]_ ,
    \new_[7388]_ , \new_[7389]_ , \new_[7390]_ , \new_[7391]_ ,
    \new_[7392]_ , \new_[7393]_ , \new_[7394]_ , \new_[7395]_ ,
    \new_[7396]_ , \new_[7397]_ , \new_[7398]_ , \new_[7399]_ ,
    \new_[7400]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7404]_ , \new_[7405]_ , \new_[7406]_ , \new_[7407]_ ,
    \new_[7408]_ , \new_[7409]_ , \new_[7410]_ , \new_[7411]_ ,
    \new_[7412]_ , \new_[7413]_ , \new_[7414]_ , \new_[7415]_ ,
    \new_[7416]_ , \new_[7417]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7422]_ , \new_[7423]_ ,
    \new_[7424]_ , \new_[7425]_ , \new_[7426]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7429]_ , \new_[7430]_ , \new_[7431]_ ,
    \new_[7432]_ , \new_[7434]_ , \new_[7435]_ , \new_[7436]_ ,
    \new_[7437]_ , \new_[7438]_ , \new_[7439]_ , \new_[7440]_ ,
    \new_[7441]_ , \new_[7445]_ , \new_[7446]_ , \new_[7447]_ ,
    \new_[7448]_ , \new_[7449]_ , \new_[7450]_ , \new_[7451]_ ,
    \new_[7453]_ , \new_[7595]_ , \new_[7599]_ , \new_[7603]_ ,
    \new_[7646]_ , \new_[7653]_ , \new_[7656]_ , \new_[7699]_ ,
    \new_[7715]_ , \new_[7734]_ , \new_[7769]_ , \new_[7777]_ ,
    \new_[7780]_ , \new_[7798]_ , \new_[7800]_ , \new_[7802]_ ,
    \new_[7807]_ , \new_[7822]_ , \new_[7870]_ , \new_[7871]_ ,
    \new_[7872]_ , \new_[7873]_ , \new_[7874]_ , \new_[7875]_ ,
    \new_[7876]_ , \new_[7877]_ , \new_[7878]_ , \new_[7879]_ ,
    \new_[7880]_ , \new_[7881]_ , \new_[7882]_ , \new_[7883]_ ,
    \new_[7884]_ , \new_[7885]_ , \new_[7887]_ , \new_[7888]_ ,
    \new_[7889]_ , \new_[7890]_ , \new_[7891]_ , \new_[7892]_ ,
    \new_[7893]_ , \new_[7894]_ , \new_[7895]_ , \new_[7896]_ ,
    \new_[7897]_ , \new_[7898]_ , \new_[7899]_ , \new_[7900]_ ,
    \new_[7901]_ , \new_[7902]_ , \new_[7903]_ , \new_[7904]_ ,
    \new_[7905]_ , \new_[7906]_ , \new_[7907]_ , \new_[7909]_ ,
    \new_[7910]_ , \new_[7911]_ , \new_[7912]_ , \new_[7913]_ ,
    \new_[7915]_ , \new_[7916]_ , \new_[7917]_ , \new_[7918]_ ,
    \new_[7919]_ , \new_[7920]_ , \new_[7921]_ , \new_[7922]_ ,
    \new_[7923]_ , \new_[7924]_ , \new_[7925]_ , \new_[7926]_ ,
    \new_[7927]_ , \new_[7928]_ , \new_[7929]_ , \new_[7930]_ ,
    \new_[7931]_ , \new_[7932]_ , \new_[7933]_ , \new_[7934]_ ,
    \new_[7935]_ , \new_[7936]_ , \new_[7937]_ , \new_[7938]_ ,
    \new_[7939]_ , \new_[7940]_ , \new_[7941]_ , \new_[7942]_ ,
    \new_[7943]_ , \new_[7944]_ , \new_[7945]_ , \new_[7946]_ ,
    \new_[7947]_ , \new_[7948]_ , \new_[7949]_ , \new_[7950]_ ,
    \new_[7951]_ , \new_[7952]_ , \new_[7953]_ , \new_[7954]_ ,
    \new_[7955]_ , \new_[7956]_ , \new_[7957]_ , \new_[7958]_ ,
    \new_[7959]_ , \new_[7960]_ , \new_[7961]_ , \new_[7962]_ ,
    \new_[7963]_ , \new_[7964]_ , \new_[7965]_ , \new_[7966]_ ,
    \new_[7967]_ , \new_[7968]_ , \new_[7969]_ , \new_[7970]_ ,
    \new_[7971]_ , \new_[7972]_ , \new_[7973]_ , \new_[7974]_ ,
    \new_[7975]_ , \new_[7976]_ , \new_[7977]_ , \new_[7978]_ ,
    \new_[7979]_ , \new_[7980]_ , \new_[7981]_ , \new_[7982]_ ,
    \new_[7983]_ , \new_[7984]_ , \new_[7985]_ , \new_[7986]_ ,
    \new_[7987]_ , \new_[7988]_ , \new_[7989]_ , \new_[7990]_ ,
    \new_[7991]_ , \new_[7993]_ , \new_[7994]_ , \new_[7995]_ ,
    \new_[7996]_ , \new_[7997]_ , \new_[7998]_ , \new_[7999]_ ,
    \new_[8000]_ , \new_[8001]_ , \new_[8002]_ , \new_[8003]_ ,
    \new_[8004]_ , \new_[8005]_ , \new_[8006]_ , \new_[8007]_ ,
    \new_[8008]_ , \new_[8009]_ , \new_[8010]_ , \new_[8011]_ ,
    \new_[8012]_ , \new_[8013]_ , \new_[8014]_ , \new_[8015]_ ,
    \new_[8016]_ , \new_[8017]_ , \new_[8018]_ , \new_[8019]_ ,
    \new_[8020]_ , \new_[8021]_ , \new_[8022]_ , \new_[8023]_ ,
    \new_[8024]_ , \new_[8025]_ , \new_[8026]_ , \new_[8027]_ ,
    \new_[8028]_ , \new_[8029]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8032]_ , \new_[8033]_ , \new_[8034]_ , \new_[8035]_ ,
    \new_[8036]_ , \new_[8037]_ , \new_[8038]_ , \new_[8039]_ ,
    \new_[8040]_ , \new_[8041]_ , \new_[8042]_ , \new_[8043]_ ,
    \new_[8044]_ , \new_[8045]_ , \new_[8046]_ , \new_[8047]_ ,
    \new_[8048]_ , \new_[8049]_ , \new_[8050]_ , \new_[8051]_ ,
    \new_[8052]_ , \new_[8053]_ , \new_[8054]_ , \new_[8055]_ ,
    \new_[8056]_ , \new_[8057]_ , \new_[8058]_ , \new_[8059]_ ,
    \new_[8060]_ , \new_[8061]_ , \new_[8062]_ , \new_[8063]_ ,
    \new_[8064]_ , \new_[8065]_ , \new_[8066]_ , \new_[8067]_ ,
    \new_[8068]_ , \new_[8069]_ , \new_[8070]_ , \new_[8071]_ ,
    \new_[8072]_ , \new_[8073]_ , \new_[8074]_ , \new_[8075]_ ,
    \new_[8076]_ , \new_[8077]_ , \new_[8078]_ , \new_[8079]_ ,
    \new_[8080]_ , \new_[8081]_ , \new_[8082]_ , \new_[8083]_ ,
    \new_[8085]_ , \new_[8086]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8089]_ , \new_[8090]_ , \new_[8091]_ , \new_[8092]_ ,
    \new_[8093]_ , \new_[8094]_ , \new_[8095]_ , \new_[8096]_ ,
    \new_[8097]_ , \new_[8098]_ , \new_[8099]_ , \new_[8100]_ ,
    \new_[8101]_ , \new_[8102]_ , \new_[8103]_ , \new_[8104]_ ,
    \new_[8105]_ , \new_[8106]_ , \new_[8107]_ , \new_[8108]_ ,
    \new_[8109]_ , \new_[8110]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8113]_ , \new_[8114]_ , \new_[8115]_ , \new_[8116]_ ,
    \new_[8117]_ , \new_[8118]_ , \new_[8119]_ , \new_[8120]_ ,
    \new_[8121]_ , \new_[8122]_ , \new_[8123]_ , \new_[8124]_ ,
    \new_[8125]_ , \new_[8126]_ , \new_[8127]_ , \new_[8128]_ ,
    \new_[8129]_ , \new_[8131]_ , \new_[8132]_ , \new_[8133]_ ,
    \new_[8134]_ , \new_[8136]_ , \new_[8137]_ , \new_[8138]_ ,
    \new_[8139]_ , \new_[8140]_ , \new_[8142]_ , \new_[8143]_ ,
    \new_[8144]_ , \new_[8145]_ , \new_[8146]_ , \new_[8156]_ ,
    \new_[8161]_ , \new_[8172]_ , \new_[8173]_ , \new_[8175]_ ,
    \new_[8176]_ , \new_[8177]_ , \new_[8178]_ , \new_[8188]_ ,
    \new_[8197]_ , \new_[8219]_ , \new_[8220]_ , \new_[8221]_ ,
    \new_[8223]_ , \new_[8224]_ , \new_[8225]_ , \new_[8235]_ ,
    \new_[8259]_ , \new_[8268]_ , \new_[8279]_ , \new_[8281]_ ,
    \new_[8282]_ , \new_[8283]_ , \new_[8284]_ , \new_[8285]_ ,
    \new_[8286]_ , \new_[8287]_ , \new_[8288]_ , \new_[8289]_ ,
    \new_[8290]_ , \new_[8291]_ , \new_[8292]_ , \new_[8293]_ ,
    \new_[8294]_ , \new_[8295]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8302]_ , \new_[8303]_ , \new_[8304]_ , \new_[8305]_ ,
    \new_[8306]_ , \new_[8307]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8310]_ , \new_[8311]_ , \new_[8312]_ , \new_[8313]_ ,
    \new_[8314]_ , \new_[8315]_ , \new_[8316]_ , \new_[8317]_ ,
    \new_[8318]_ , \new_[8319]_ , \new_[8320]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8324]_ , \new_[8325]_ ,
    \new_[8326]_ , \new_[8327]_ , \new_[8328]_ , \new_[8329]_ ,
    \new_[8330]_ , \new_[8331]_ , \new_[8332]_ , \new_[8333]_ ,
    \new_[8334]_ , \new_[8335]_ , \new_[8336]_ , \new_[8337]_ ,
    \new_[8338]_ , \new_[8339]_ , \new_[8340]_ , \new_[8341]_ ,
    \new_[8342]_ , \new_[8343]_ , \new_[8344]_ , \new_[8345]_ ,
    \new_[8346]_ , \new_[8347]_ , \new_[8348]_ , \new_[8349]_ ,
    \new_[8350]_ , \new_[8351]_ , \new_[8352]_ , \new_[8353]_ ,
    \new_[8354]_ , \new_[8355]_ , \new_[8356]_ , \new_[8357]_ ,
    \new_[8358]_ , \new_[8359]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8362]_ , \new_[8363]_ , \new_[8364]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8376]_ , \new_[8377]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8380]_ , \new_[8381]_ ,
    \new_[8382]_ , \new_[8383]_ , \new_[8384]_ , \new_[8385]_ ,
    \new_[8386]_ , \new_[8387]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8390]_ , \new_[8391]_ , \new_[8392]_ , \new_[8393]_ ,
    \new_[8394]_ , \new_[8395]_ , \new_[8396]_ , \new_[8397]_ ,
    \new_[8398]_ , \new_[8399]_ , \new_[8400]_ , \new_[8401]_ ,
    \new_[8402]_ , \new_[8403]_ , \new_[8404]_ , \new_[8405]_ ,
    \new_[8406]_ , \new_[8407]_ , \new_[8408]_ , \new_[8409]_ ,
    \new_[8410]_ , \new_[8411]_ , \new_[8412]_ , \new_[8413]_ ,
    \new_[8414]_ , \new_[8415]_ , \new_[8416]_ , \new_[8417]_ ,
    \new_[8418]_ , \new_[8419]_ , \new_[8420]_ , \new_[8421]_ ,
    \new_[8422]_ , \new_[8423]_ , \new_[8424]_ , \new_[8425]_ ,
    \new_[8426]_ , \new_[8427]_ , \new_[8428]_ , \new_[8429]_ ,
    \new_[8430]_ , \new_[8431]_ , \new_[8432]_ , \new_[8433]_ ,
    \new_[8434]_ , \new_[8435]_ , \new_[8436]_ , \new_[8437]_ ,
    \new_[8438]_ , \new_[8439]_ , \new_[8440]_ , \new_[8441]_ ,
    \new_[8442]_ , \new_[8443]_ , \new_[8444]_ , \new_[8445]_ ,
    \new_[8446]_ , \new_[8447]_ , \new_[8449]_ , \new_[8450]_ ,
    \new_[8451]_ , \new_[8452]_ , \new_[8453]_ , \new_[8454]_ ,
    \new_[8455]_ , \new_[8456]_ , \new_[8457]_ , \new_[8458]_ ,
    \new_[8459]_ , \new_[8464]_ , \new_[8465]_ , \new_[8468]_ ,
    \new_[8469]_ , \new_[8470]_ , \new_[8471]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8474]_ , \new_[8475]_ , \new_[8476]_ ,
    \new_[8477]_ , \new_[8478]_ , \new_[8479]_ , \new_[8480]_ ,
    \new_[8481]_ , \new_[8482]_ , \new_[8483]_ , \new_[8484]_ ,
    \new_[8485]_ , \new_[8486]_ , \new_[8487]_ , \new_[8488]_ ,
    \new_[8489]_ , \new_[8490]_ , \new_[8491]_ , \new_[8492]_ ,
    \new_[8493]_ , \new_[8494]_ , \new_[8495]_ , \new_[8496]_ ,
    \new_[8497]_ , \new_[8498]_ , \new_[8499]_ , \new_[8501]_ ,
    \new_[8502]_ , \new_[8504]_ , \new_[8505]_ , \new_[8506]_ ,
    \new_[8507]_ , \new_[8508]_ , \new_[8509]_ , \new_[8510]_ ,
    \new_[8511]_ , \new_[8512]_ , \new_[8513]_ , \new_[8514]_ ,
    \new_[8515]_ , \new_[8516]_ , \new_[8517]_ , \new_[8518]_ ,
    \new_[8519]_ , \new_[8520]_ , \new_[8521]_ , \new_[8522]_ ,
    \new_[8523]_ , \new_[8524]_ , \new_[8525]_ , \new_[8526]_ ,
    \new_[8527]_ , \new_[8528]_ , \new_[8529]_ , \new_[8530]_ ,
    \new_[8531]_ , \new_[8532]_ , \new_[8533]_ , \new_[8534]_ ,
    \new_[8535]_ , \new_[8536]_ , \new_[8537]_ , \new_[8538]_ ,
    \new_[8539]_ , \new_[8540]_ , \new_[8541]_ , \new_[8542]_ ,
    \new_[8543]_ , \new_[8544]_ , \new_[8545]_ , \new_[8546]_ ,
    \new_[8547]_ , \new_[8548]_ , \new_[8549]_ , \new_[8550]_ ,
    \new_[8551]_ , \new_[8552]_ , \new_[8553]_ , \new_[8554]_ ,
    \new_[8555]_ , \new_[8556]_ , \new_[8557]_ , \new_[8558]_ ,
    \new_[8559]_ , \new_[8560]_ , \new_[8561]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8564]_ , \new_[8565]_ , \new_[8566]_ ,
    \new_[8567]_ , \new_[8568]_ , \new_[8569]_ , \new_[8570]_ ,
    \new_[8571]_ , \new_[8572]_ , \new_[8573]_ , \new_[8574]_ ,
    \new_[8575]_ , \new_[8576]_ , \new_[8577]_ , \new_[8578]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8581]_ , \new_[8582]_ ,
    \new_[8583]_ , \new_[8584]_ , \new_[8585]_ , \new_[8586]_ ,
    \new_[8587]_ , \new_[8588]_ , \new_[8589]_ , \new_[8590]_ ,
    \new_[8591]_ , \new_[8592]_ , \new_[8593]_ , \new_[8594]_ ,
    \new_[8595]_ , \new_[8596]_ , \new_[8597]_ , \new_[8598]_ ,
    \new_[8599]_ , \new_[8600]_ , \new_[8601]_ , \new_[8602]_ ,
    \new_[8603]_ , \new_[8604]_ , \new_[8605]_ , \new_[8606]_ ,
    \new_[8607]_ , \new_[8608]_ , \new_[8609]_ , \new_[8610]_ ,
    \new_[8611]_ , \new_[8612]_ , \new_[8613]_ , \new_[8614]_ ,
    \new_[8615]_ , \new_[8616]_ , \new_[8617]_ , \new_[8618]_ ,
    \new_[8619]_ , \new_[8620]_ , \new_[8621]_ , \new_[8622]_ ,
    \new_[8623]_ , \new_[8624]_ , \new_[8625]_ , \new_[8626]_ ,
    \new_[8627]_ , \new_[8628]_ , \new_[8629]_ , \new_[8630]_ ,
    \new_[8631]_ , \new_[8632]_ , \new_[8633]_ , \new_[8634]_ ,
    \new_[8635]_ , \new_[8636]_ , \new_[8637]_ , \new_[8638]_ ,
    \new_[8639]_ , \new_[8640]_ , \new_[8641]_ , \new_[8642]_ ,
    \new_[8643]_ , \new_[8644]_ , \new_[8645]_ , \new_[8646]_ ,
    \new_[8647]_ , \new_[8648]_ , \new_[8649]_ , \new_[8650]_ ,
    \new_[8651]_ , \new_[8652]_ , \new_[8653]_ , \new_[8654]_ ,
    \new_[8655]_ , \new_[8656]_ , \new_[8657]_ , \new_[8658]_ ,
    \new_[8659]_ , \new_[8660]_ , \new_[8661]_ , \new_[8662]_ ,
    \new_[8663]_ , \new_[8664]_ , \new_[8666]_ , \new_[8668]_ ,
    \new_[8669]_ , \new_[8670]_ , \new_[8671]_ , \new_[8672]_ ,
    \new_[8673]_ , \new_[8674]_ , \new_[8675]_ , \new_[8676]_ ,
    \new_[8677]_ , \new_[8678]_ , \new_[8679]_ , \new_[8680]_ ,
    \new_[8681]_ , \new_[8682]_ , \new_[8683]_ , \new_[8684]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8692]_ , \new_[8698]_ ,
    \new_[8699]_ , \new_[8700]_ , \new_[8701]_ , \new_[8702]_ ,
    \new_[8703]_ , \new_[8704]_ , \new_[8705]_ , \new_[8706]_ ,
    \new_[8707]_ , \new_[8708]_ , \new_[8709]_ , \new_[8710]_ ,
    \new_[8711]_ , \new_[8712]_ , \new_[8713]_ , \new_[8714]_ ,
    \new_[8715]_ , \new_[8716]_ , \new_[8717]_ , \new_[8718]_ ,
    \new_[8719]_ , \new_[8720]_ , \new_[8721]_ , \new_[8722]_ ,
    \new_[8723]_ , \new_[8724]_ , \new_[8725]_ , \new_[8726]_ ,
    \new_[8727]_ , \new_[8728]_ , \new_[8729]_ , \new_[8730]_ ,
    \new_[8731]_ , \new_[8732]_ , \new_[8733]_ , \new_[8734]_ ,
    \new_[8735]_ , \new_[8736]_ , \new_[8737]_ , \new_[8738]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8741]_ , \new_[8742]_ ,
    \new_[8743]_ , \new_[8744]_ , \new_[8745]_ , \new_[8746]_ ,
    \new_[8747]_ , \new_[8748]_ , \new_[8749]_ , \new_[8750]_ ,
    \new_[8751]_ , \new_[8752]_ , \new_[8753]_ , \new_[8754]_ ,
    \new_[8755]_ , \new_[8756]_ , \new_[8757]_ , \new_[8758]_ ,
    \new_[8759]_ , \new_[8760]_ , \new_[8761]_ , \new_[8762]_ ,
    \new_[8763]_ , \new_[8764]_ , \new_[8765]_ , \new_[8766]_ ,
    \new_[8767]_ , \new_[8768]_ , \new_[8769]_ , \new_[8770]_ ,
    \new_[8771]_ , \new_[8772]_ , \new_[8773]_ , \new_[8774]_ ,
    \new_[8775]_ , \new_[8776]_ , \new_[8777]_ , \new_[8778]_ ,
    \new_[8779]_ , \new_[8780]_ , \new_[8781]_ , \new_[8782]_ ,
    \new_[8783]_ , \new_[8784]_ , \new_[8785]_ , \new_[8786]_ ,
    \new_[8787]_ , \new_[8788]_ , \new_[8789]_ , \new_[8790]_ ,
    \new_[8791]_ , \new_[8792]_ , \new_[8793]_ , \new_[8794]_ ,
    \new_[8795]_ , \new_[8796]_ , \new_[8797]_ , \new_[8798]_ ,
    \new_[8799]_ , \new_[8800]_ , \new_[8801]_ , \new_[8802]_ ,
    \new_[8803]_ , \new_[8804]_ , \new_[8805]_ , \new_[8806]_ ,
    \new_[8807]_ , \new_[8808]_ , \new_[8809]_ , \new_[8810]_ ,
    \new_[8811]_ , \new_[8812]_ , \new_[8813]_ , \new_[8814]_ ,
    \new_[8815]_ , \new_[8816]_ , \new_[8817]_ , \new_[8818]_ ,
    \new_[8819]_ , \new_[8820]_ , \new_[8821]_ , \new_[8822]_ ,
    \new_[8823]_ , \new_[8824]_ , \new_[8825]_ , \new_[8826]_ ,
    \new_[8827]_ , \new_[8828]_ , \new_[8829]_ , \new_[8830]_ ,
    \new_[8831]_ , \new_[8832]_ , \new_[8833]_ , \new_[8834]_ ,
    \new_[8835]_ , \new_[8836]_ , \new_[8837]_ , \new_[8838]_ ,
    \new_[8839]_ , \new_[8840]_ , \new_[8841]_ , \new_[8842]_ ,
    \new_[8843]_ , \new_[8844]_ , \new_[8845]_ , \new_[8846]_ ,
    \new_[8847]_ , \new_[8848]_ , \new_[8849]_ , \new_[8850]_ ,
    \new_[8851]_ , \new_[8852]_ , \new_[8853]_ , \new_[8854]_ ,
    \new_[8855]_ , \new_[8856]_ , \new_[8857]_ , \new_[8858]_ ,
    \new_[8859]_ , \new_[8860]_ , \new_[8861]_ , \new_[8862]_ ,
    \new_[8863]_ , \new_[8864]_ , \new_[8865]_ , \new_[8866]_ ,
    \new_[8867]_ , \new_[8868]_ , \new_[8869]_ , \new_[8870]_ ,
    \new_[8871]_ , \new_[8872]_ , \new_[8873]_ , \new_[8874]_ ,
    \new_[8875]_ , \new_[8876]_ , \new_[8878]_ , \new_[8879]_ ,
    \new_[8880]_ , \new_[8881]_ , \new_[8882]_ , \new_[8883]_ ,
    \new_[8884]_ , \new_[8885]_ , \new_[8886]_ , \new_[8887]_ ,
    \new_[8888]_ , \new_[8889]_ , \new_[8890]_ , \new_[8891]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8894]_ , \new_[8895]_ ,
    \new_[8896]_ , \new_[8897]_ , \new_[8898]_ , \new_[8899]_ ,
    \new_[8900]_ , \new_[8901]_ , \new_[8902]_ , \new_[8903]_ ,
    \new_[8904]_ , \new_[8905]_ , \new_[8906]_ , \new_[8907]_ ,
    \new_[8908]_ , \new_[8909]_ , \new_[8910]_ , \new_[8911]_ ,
    \new_[8912]_ , \new_[8913]_ , \new_[8914]_ , \new_[8915]_ ,
    \new_[8916]_ , \new_[8917]_ , \new_[8918]_ , \new_[8919]_ ,
    \new_[8920]_ , \new_[8921]_ , \new_[8922]_ , \new_[8923]_ ,
    \new_[8924]_ , \new_[8925]_ , \new_[8926]_ , \new_[8927]_ ,
    \new_[8928]_ , \new_[8929]_ , \new_[8930]_ , \new_[8931]_ ,
    \new_[8932]_ , \new_[8933]_ , \new_[8934]_ , \new_[8935]_ ,
    \new_[8936]_ , \new_[8937]_ , \new_[8938]_ , \new_[8939]_ ,
    \new_[8940]_ , \new_[8941]_ , \new_[8942]_ , \new_[8943]_ ,
    \new_[8944]_ , \new_[8945]_ , \new_[8946]_ , \new_[8947]_ ,
    \new_[8948]_ , \new_[8949]_ , \new_[8950]_ , \new_[8952]_ ,
    \new_[8953]_ , \new_[8954]_ , \new_[8955]_ , \new_[8956]_ ,
    \new_[8957]_ , \new_[8958]_ , \new_[8959]_ , \new_[8960]_ ,
    \new_[8961]_ , \new_[8962]_ , \new_[8963]_ , \new_[8964]_ ,
    \new_[8965]_ , \new_[8966]_ , \new_[8967]_ , \new_[8968]_ ,
    \new_[8969]_ , \new_[8970]_ , \new_[8971]_ , \new_[8972]_ ,
    \new_[8973]_ , \new_[8974]_ , \new_[8975]_ , \new_[8976]_ ,
    \new_[8977]_ , \new_[8978]_ , \new_[8979]_ , \new_[8980]_ ,
    \new_[8981]_ , \new_[8982]_ , \new_[8983]_ , \new_[8984]_ ,
    \new_[8985]_ , \new_[8986]_ , \new_[8987]_ , \new_[8988]_ ,
    \new_[8989]_ , \new_[8990]_ , \new_[8991]_ , \new_[8992]_ ,
    \new_[8993]_ , \new_[8994]_ , \new_[8995]_ , \new_[8996]_ ,
    \new_[8997]_ , \new_[8998]_ , \new_[8999]_ , \new_[9000]_ ,
    \new_[9001]_ , \new_[9002]_ , \new_[9003]_ , \new_[9004]_ ,
    \new_[9005]_ , \new_[9006]_ , \new_[9007]_ , \new_[9008]_ ,
    \new_[9009]_ , \new_[9010]_ , \new_[9011]_ , \new_[9012]_ ,
    \new_[9013]_ , \new_[9014]_ , \new_[9015]_ , \new_[9016]_ ,
    \new_[9017]_ , \new_[9018]_ , \new_[9019]_ , \new_[9020]_ ,
    \new_[9021]_ , \new_[9022]_ , \new_[9023]_ , \new_[9024]_ ,
    \new_[9025]_ , \new_[9026]_ , \new_[9027]_ , \new_[9028]_ ,
    \new_[9029]_ , \new_[9030]_ , \new_[9031]_ , \new_[9032]_ ,
    \new_[9033]_ , \new_[9034]_ , \new_[9035]_ , \new_[9036]_ ,
    \new_[9037]_ , \new_[9038]_ , \new_[9039]_ , \new_[9040]_ ,
    \new_[9041]_ , \new_[9042]_ , \new_[9043]_ , \new_[9044]_ ,
    \new_[9045]_ , \new_[9046]_ , \new_[9047]_ , \new_[9048]_ ,
    \new_[9049]_ , \new_[9050]_ , \new_[9051]_ , \new_[9052]_ ,
    \new_[9053]_ , \new_[9054]_ , \new_[9055]_ , \new_[9056]_ ,
    \new_[9057]_ , \new_[9058]_ , \new_[9059]_ , \new_[9060]_ ,
    \new_[9061]_ , \new_[9062]_ , \new_[9063]_ , \new_[9064]_ ,
    \new_[9065]_ , \new_[9066]_ , \new_[9067]_ , \new_[9068]_ ,
    \new_[9069]_ , \new_[9070]_ , \new_[9071]_ , \new_[9072]_ ,
    \new_[9073]_ , \new_[9074]_ , \new_[9075]_ , \new_[9076]_ ,
    \new_[9077]_ , \new_[9078]_ , \new_[9079]_ , \new_[9080]_ ,
    \new_[9081]_ , \new_[9082]_ , \new_[9083]_ , \new_[9084]_ ,
    \new_[9085]_ , \new_[9086]_ , \new_[9087]_ , \new_[9088]_ ,
    \new_[9090]_ , \new_[9091]_ , \new_[9092]_ , \new_[9093]_ ,
    \new_[9094]_ , \new_[9095]_ , \new_[9096]_ , \new_[9097]_ ,
    \new_[9098]_ , \new_[9099]_ , \new_[9100]_ , \new_[9101]_ ,
    \new_[9102]_ , \new_[9103]_ , \new_[9104]_ , \new_[9105]_ ,
    \new_[9106]_ , \new_[9107]_ , \new_[9108]_ , \new_[9109]_ ,
    \new_[9110]_ , \new_[9111]_ , \new_[9112]_ , \new_[9113]_ ,
    \new_[9114]_ , \new_[9115]_ , \new_[9116]_ , \new_[9117]_ ,
    \new_[9118]_ , \new_[9119]_ , \new_[9121]_ , \new_[9122]_ ,
    \new_[9123]_ , \new_[9124]_ , \new_[9125]_ , \new_[9126]_ ,
    \new_[9127]_ , \new_[9128]_ , \new_[9130]_ , \new_[9131]_ ,
    \new_[9132]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9151]_ , \new_[9152]_ , \new_[9153]_ ,
    \new_[9154]_ , \new_[9155]_ , \new_[9156]_ , \new_[9157]_ ,
    \new_[9158]_ , \new_[9159]_ , \new_[9160]_ , \new_[9161]_ ,
    \new_[9162]_ , \new_[9163]_ , \new_[9164]_ , \new_[9165]_ ,
    \new_[9166]_ , \new_[9167]_ , \new_[9168]_ , \new_[9169]_ ,
    \new_[9171]_ , \new_[9172]_ , \new_[9173]_ , \new_[9174]_ ,
    \new_[9175]_ , \new_[9176]_ , \new_[9177]_ , \new_[9178]_ ,
    \new_[9179]_ , \new_[9180]_ , \new_[9181]_ , \new_[9182]_ ,
    \new_[9183]_ , \new_[9184]_ , \new_[9185]_ , \new_[9186]_ ,
    \new_[9187]_ , \new_[9188]_ , \new_[9190]_ , \new_[9191]_ ,
    \new_[9192]_ , \new_[9193]_ , \new_[9194]_ , \new_[9195]_ ,
    \new_[9196]_ , \new_[9198]_ , \new_[9199]_ , \new_[9200]_ ,
    \new_[9201]_ , \new_[9202]_ , \new_[9203]_ , \new_[9204]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9207]_ , \new_[9208]_ ,
    \new_[9209]_ , \new_[9210]_ , \new_[9211]_ , \new_[9212]_ ,
    \new_[9213]_ , \new_[9214]_ , \new_[9215]_ , \new_[9216]_ ,
    \new_[9217]_ , \new_[9218]_ , \new_[9219]_ , \new_[9220]_ ,
    \new_[9221]_ , \new_[9222]_ , \new_[9223]_ , \new_[9224]_ ,
    \new_[9225]_ , \new_[9226]_ , \new_[9227]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9231]_ , \new_[9232]_ ,
    \new_[9233]_ , \new_[9234]_ , \new_[9235]_ , \new_[9236]_ ,
    \new_[9237]_ , \new_[9238]_ , \new_[9239]_ , \new_[9240]_ ,
    \new_[9241]_ , \new_[9242]_ , \new_[9243]_ , \new_[9244]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9247]_ , \new_[9248]_ ,
    \new_[9249]_ , \new_[9250]_ , \new_[9251]_ , \new_[9252]_ ,
    \new_[9253]_ , \new_[9254]_ , \new_[9255]_ , \new_[9256]_ ,
    \new_[9257]_ , \new_[9258]_ , \new_[9259]_ , \new_[9260]_ ,
    \new_[9261]_ , \new_[9262]_ , \new_[9263]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9266]_ , \new_[9267]_ , \new_[9268]_ ,
    \new_[9269]_ , \new_[9270]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9273]_ , \new_[9274]_ , \new_[9275]_ , \new_[9276]_ ,
    \new_[9277]_ , \new_[9278]_ , \new_[9279]_ , \new_[9280]_ ,
    \new_[9281]_ , \new_[9282]_ , \new_[9283]_ , \new_[9284]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9291]_ , \new_[9292]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9295]_ , \new_[9296]_ ,
    \new_[9297]_ , \new_[9298]_ , \new_[9299]_ , \new_[9300]_ ,
    \new_[9301]_ , \new_[9302]_ , \new_[9303]_ , \new_[9304]_ ,
    \new_[9305]_ , \new_[9306]_ , \new_[9307]_ , \new_[9308]_ ,
    \new_[9309]_ , \new_[9310]_ , \new_[9311]_ , \new_[9312]_ ,
    \new_[9313]_ , \new_[9314]_ , \new_[9315]_ , \new_[9316]_ ,
    \new_[9317]_ , \new_[9318]_ , \new_[9319]_ , \new_[9320]_ ,
    \new_[9321]_ , \new_[9322]_ , \new_[9323]_ , \new_[9324]_ ,
    \new_[9325]_ , \new_[9326]_ , \new_[9327]_ , \new_[9328]_ ,
    \new_[9329]_ , \new_[9330]_ , \new_[9331]_ , \new_[9332]_ ,
    \new_[9333]_ , \new_[9334]_ , \new_[9335]_ , \new_[9336]_ ,
    \new_[9337]_ , \new_[9338]_ , \new_[9339]_ , \new_[9340]_ ,
    \new_[9341]_ , \new_[9342]_ , \new_[9343]_ , \new_[9344]_ ,
    \new_[9345]_ , \new_[9346]_ , \new_[9347]_ , \new_[9348]_ ,
    \new_[9349]_ , \new_[9350]_ , \new_[9351]_ , \new_[9352]_ ,
    \new_[9353]_ , \new_[9354]_ , \new_[9355]_ , \new_[9356]_ ,
    \new_[9357]_ , \new_[9358]_ , \new_[9359]_ , \new_[9360]_ ,
    \new_[9361]_ , \new_[9362]_ , \new_[9363]_ , \new_[9364]_ ,
    \new_[9365]_ , \new_[9366]_ , \new_[9367]_ , \new_[9368]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9371]_ , \new_[9372]_ ,
    \new_[9373]_ , \new_[9374]_ , \new_[9375]_ , \new_[9376]_ ,
    \new_[9377]_ , \new_[9378]_ , \new_[9379]_ , \new_[9380]_ ,
    \new_[9381]_ , \new_[9382]_ , \new_[9383]_ , \new_[9384]_ ,
    \new_[9385]_ , \new_[9386]_ , \new_[9387]_ , \new_[9388]_ ,
    \new_[9389]_ , \new_[9390]_ , \new_[9391]_ , \new_[9392]_ ,
    \new_[9393]_ , \new_[9394]_ , \new_[9395]_ , \new_[9396]_ ,
    \new_[9397]_ , \new_[9398]_ , \new_[9399]_ , \new_[9400]_ ,
    \new_[9401]_ , \new_[9402]_ , \new_[9403]_ , \new_[9404]_ ,
    \new_[9405]_ , \new_[9406]_ , \new_[9407]_ , \new_[9408]_ ,
    \new_[9409]_ , \new_[9410]_ , \new_[9411]_ , \new_[9412]_ ,
    \new_[9413]_ , \new_[9414]_ , \new_[9415]_ , \new_[9416]_ ,
    \new_[9417]_ , \new_[9418]_ , \new_[9419]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9422]_ , \new_[9423]_ , \new_[9424]_ ,
    \new_[9425]_ , \new_[9426]_ , \new_[9427]_ , \new_[9428]_ ,
    \new_[9429]_ , \new_[9430]_ , \new_[9431]_ , \new_[9432]_ ,
    \new_[9433]_ , \new_[9434]_ , \new_[9435]_ , \new_[9436]_ ,
    \new_[9437]_ , \new_[9438]_ , \new_[9439]_ , \new_[9440]_ ,
    \new_[9441]_ , \new_[9442]_ , \new_[9443]_ , \new_[9444]_ ,
    \new_[9445]_ , \new_[9446]_ , \new_[9447]_ , \new_[9448]_ ,
    \new_[9449]_ , \new_[9450]_ , \new_[9451]_ , \new_[9452]_ ,
    \new_[9453]_ , \new_[9454]_ , \new_[9455]_ , \new_[9456]_ ,
    \new_[9457]_ , \new_[9458]_ , \new_[9459]_ , \new_[9460]_ ,
    \new_[9461]_ , \new_[9462]_ , \new_[9463]_ , \new_[9464]_ ,
    \new_[9465]_ , \new_[9466]_ , \new_[9467]_ , \new_[9468]_ ,
    \new_[9469]_ , \new_[9470]_ , \new_[9471]_ , \new_[9472]_ ,
    \new_[9473]_ , \new_[9474]_ , \new_[9475]_ , \new_[9476]_ ,
    \new_[9477]_ , \new_[9478]_ , \new_[9479]_ , \new_[9480]_ ,
    \new_[9481]_ , \new_[9482]_ , \new_[9483]_ , \new_[9484]_ ,
    \new_[9485]_ , \new_[9486]_ , \new_[9487]_ , \new_[9488]_ ,
    \new_[9489]_ , \new_[9490]_ , \new_[9491]_ , \new_[9492]_ ,
    \new_[9493]_ , \new_[9494]_ , \new_[9495]_ , \new_[9496]_ ,
    \new_[9497]_ , \new_[9498]_ , \new_[9499]_ , \new_[9500]_ ,
    \new_[9501]_ , \new_[9502]_ , \new_[9503]_ , \new_[9504]_ ,
    \new_[9505]_ , \new_[9506]_ , \new_[9507]_ , \new_[9508]_ ,
    \new_[9509]_ , \new_[9510]_ , \new_[9511]_ , \new_[9512]_ ,
    \new_[9513]_ , \new_[9514]_ , \new_[9515]_ , \new_[9516]_ ,
    \new_[9517]_ , \new_[9518]_ , \new_[9519]_ , \new_[9520]_ ,
    \new_[9521]_ , \new_[9522]_ , \new_[9523]_ , \new_[9524]_ ,
    \new_[9525]_ , \new_[9526]_ , \new_[9527]_ , \new_[9528]_ ,
    \new_[9529]_ , \new_[9530]_ , \new_[9531]_ , \new_[9532]_ ,
    \new_[9533]_ , \new_[9534]_ , \new_[9535]_ , \new_[9536]_ ,
    \new_[9537]_ , \new_[9538]_ , \new_[9539]_ , \new_[9540]_ ,
    \new_[9541]_ , \new_[9542]_ , \new_[9543]_ , \new_[9544]_ ,
    \new_[9545]_ , \new_[9546]_ , \new_[9547]_ , \new_[9548]_ ,
    \new_[9549]_ , \new_[9550]_ , \new_[9551]_ , \new_[9552]_ ,
    \new_[9553]_ , \new_[9554]_ , \new_[9555]_ , \new_[9556]_ ,
    \new_[9557]_ , \new_[9558]_ , \new_[9559]_ , \new_[9560]_ ,
    \new_[9561]_ , \new_[9562]_ , \new_[9563]_ , \new_[9564]_ ,
    \new_[9565]_ , \new_[9566]_ , \new_[9567]_ , \new_[9568]_ ,
    \new_[9569]_ , \new_[9570]_ , \new_[9571]_ , \new_[9572]_ ,
    \new_[9573]_ , \new_[9574]_ , \new_[9575]_ , \new_[9576]_ ,
    \new_[9577]_ , \new_[9578]_ , \new_[9579]_ , \new_[9580]_ ,
    \new_[9581]_ , \new_[9582]_ , \new_[9583]_ , \new_[9584]_ ,
    \new_[9585]_ , \new_[9586]_ , \new_[9587]_ , \new_[9588]_ ,
    \new_[9589]_ , \new_[9590]_ , \new_[9591]_ , \new_[9592]_ ,
    \new_[9593]_ , \new_[9594]_ , \new_[9595]_ , \new_[9596]_ ,
    \new_[9597]_ , \new_[9598]_ , \new_[9599]_ , \new_[9600]_ ,
    \new_[9601]_ , \new_[9602]_ , \new_[9603]_ , \new_[9604]_ ,
    \new_[9605]_ , \new_[9606]_ , \new_[9607]_ , \new_[9608]_ ,
    \new_[9609]_ , \new_[9610]_ , \new_[9611]_ , \new_[9612]_ ,
    \new_[9613]_ , \new_[9614]_ , \new_[9615]_ , \new_[9616]_ ,
    \new_[9617]_ , \new_[9618]_ , \new_[9619]_ , \new_[9620]_ ,
    \new_[9621]_ , \new_[9622]_ , \new_[9623]_ , \new_[9624]_ ,
    \new_[9625]_ , \new_[9626]_ , \new_[9627]_ , \new_[9628]_ ,
    \new_[9629]_ , \new_[9630]_ , \new_[9631]_ , \new_[9632]_ ,
    \new_[9633]_ , \new_[9634]_ , \new_[9635]_ , \new_[9636]_ ,
    \new_[9637]_ , \new_[9638]_ , \new_[9639]_ , \new_[9640]_ ,
    \new_[9641]_ , \new_[9642]_ , \new_[9643]_ , \new_[9644]_ ,
    \new_[9645]_ , \new_[9646]_ , \new_[9647]_ , \new_[9648]_ ,
    \new_[9649]_ , \new_[9650]_ , \new_[9651]_ , \new_[9652]_ ,
    \new_[9653]_ , \new_[9654]_ , \new_[9655]_ , \new_[9656]_ ,
    \new_[9657]_ , \new_[9658]_ , \new_[9659]_ , \new_[9660]_ ,
    \new_[9661]_ , \new_[9662]_ , \new_[9663]_ , \new_[9664]_ ,
    \new_[9665]_ , \new_[9666]_ , \new_[9667]_ , \new_[9668]_ ,
    \new_[9669]_ , \new_[9670]_ , \new_[9671]_ , \new_[9672]_ ,
    \new_[9673]_ , \new_[9674]_ , \new_[9675]_ , \new_[9676]_ ,
    \new_[9677]_ , \new_[9678]_ , \new_[9679]_ , \new_[9680]_ ,
    \new_[9681]_ , \new_[9682]_ , \new_[9683]_ , \new_[9684]_ ,
    \new_[9685]_ , \new_[9686]_ , \new_[9687]_ , \new_[9688]_ ,
    \new_[9689]_ , \new_[9690]_ , \new_[9691]_ , \new_[9692]_ ,
    \new_[9693]_ , \new_[9694]_ , \new_[9695]_ , \new_[9696]_ ,
    \new_[9697]_ , \new_[9698]_ , \new_[9699]_ , \new_[9700]_ ,
    \new_[9701]_ , \new_[9702]_ , \new_[9703]_ , \new_[9704]_ ,
    \new_[9705]_ , \new_[9706]_ , \new_[9707]_ , \new_[9708]_ ,
    \new_[9709]_ , \new_[9710]_ , \new_[9711]_ , \new_[9712]_ ,
    \new_[9713]_ , \new_[9714]_ , \new_[9715]_ , \new_[9716]_ ,
    \new_[9717]_ , \new_[9718]_ , \new_[9719]_ , \new_[9720]_ ,
    \new_[9721]_ , \new_[9722]_ , \new_[9723]_ , \new_[9724]_ ,
    \new_[9725]_ , \new_[9726]_ , \new_[9727]_ , \new_[9728]_ ,
    \new_[9729]_ , \new_[9730]_ , \new_[9731]_ , \new_[9732]_ ,
    \new_[9733]_ , \new_[9734]_ , \new_[9735]_ , \new_[9736]_ ,
    \new_[9737]_ , \new_[9738]_ , \new_[9739]_ , \new_[9740]_ ,
    \new_[9741]_ , \new_[9742]_ , \new_[9743]_ , \new_[9744]_ ,
    \new_[9745]_ , \new_[9746]_ , \new_[9747]_ , \new_[9748]_ ,
    \new_[9749]_ , \new_[9750]_ , \new_[9751]_ , \new_[9752]_ ,
    \new_[9753]_ , \new_[9754]_ , \new_[9755]_ , \new_[9756]_ ,
    \new_[9757]_ , \new_[9758]_ , \new_[9759]_ , \new_[9760]_ ,
    \new_[9761]_ , \new_[9762]_ , \new_[9763]_ , \new_[9764]_ ,
    \new_[9765]_ , \new_[9766]_ , \new_[9767]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9770]_ , \new_[9771]_ , \new_[9772]_ ,
    \new_[9773]_ , \new_[9774]_ , \new_[9775]_ , \new_[9776]_ ,
    \new_[9777]_ , \new_[9778]_ , \new_[9779]_ , \new_[9780]_ ,
    \new_[9781]_ , \new_[9782]_ , \new_[9783]_ , \new_[9784]_ ,
    \new_[9785]_ , \new_[9786]_ , \new_[9787]_ , \new_[9788]_ ,
    \new_[9789]_ , \new_[9790]_ , \new_[9791]_ , \new_[9792]_ ,
    \new_[9793]_ , \new_[9794]_ , \new_[9795]_ , \new_[9796]_ ,
    \new_[9797]_ , \new_[9798]_ , \new_[9799]_ , \new_[9800]_ ,
    \new_[9801]_ , \new_[9802]_ , \new_[9803]_ , \new_[9804]_ ,
    \new_[9805]_ , \new_[9806]_ , \new_[9807]_ , \new_[9808]_ ,
    \new_[9809]_ , \new_[9810]_ , \new_[9811]_ , \new_[9812]_ ,
    \new_[9813]_ , \new_[9814]_ , \new_[9815]_ , \new_[9816]_ ,
    \new_[9817]_ , \new_[9818]_ , \new_[9819]_ , \new_[9820]_ ,
    \new_[9821]_ , \new_[9822]_ , \new_[9823]_ , \new_[9824]_ ,
    \new_[9825]_ , \new_[9826]_ , \new_[9827]_ , \new_[9828]_ ,
    \new_[9829]_ , \new_[9830]_ , \new_[9831]_ , \new_[9832]_ ,
    \new_[9833]_ , \new_[9834]_ , \new_[9835]_ , \new_[9836]_ ,
    \new_[9837]_ , \new_[9838]_ , \new_[9839]_ , \new_[9840]_ ,
    \new_[9841]_ , \new_[9842]_ , \new_[9843]_ , \new_[9844]_ ,
    \new_[9845]_ , \new_[9846]_ , \new_[9847]_ , \new_[9848]_ ,
    \new_[9849]_ , \new_[9850]_ , \new_[9851]_ , \new_[9852]_ ,
    \new_[9853]_ , \new_[9854]_ , \new_[9855]_ , \new_[9856]_ ,
    \new_[9857]_ , \new_[9858]_ , \new_[9859]_ , \new_[9860]_ ,
    \new_[9861]_ , \new_[9862]_ , \new_[9863]_ , \new_[9864]_ ,
    \new_[9865]_ , \new_[9866]_ , \new_[9867]_ , \new_[9868]_ ,
    \new_[9869]_ , \new_[9870]_ , \new_[9871]_ , \new_[9872]_ ,
    \new_[9873]_ , \new_[9874]_ , \new_[9875]_ , \new_[9876]_ ,
    \new_[9877]_ , \new_[9878]_ , \new_[9879]_ , \new_[9880]_ ,
    \new_[9881]_ , \new_[9882]_ , \new_[9883]_ , \new_[9884]_ ,
    \new_[9885]_ , \new_[9886]_ , \new_[9887]_ , \new_[9888]_ ,
    \new_[9889]_ , \new_[9890]_ , \new_[9891]_ , \new_[9892]_ ,
    \new_[9893]_ , \new_[9894]_ , \new_[9895]_ , \new_[9896]_ ,
    \new_[9897]_ , \new_[9898]_ , \new_[9899]_ , \new_[9900]_ ,
    \new_[9901]_ , \new_[9902]_ , \new_[9903]_ , \new_[9904]_ ,
    \new_[9905]_ , \new_[9906]_ , \new_[9907]_ , \new_[9908]_ ,
    \new_[9909]_ , \new_[9910]_ , \new_[9911]_ , \new_[9912]_ ,
    \new_[9913]_ , \new_[9914]_ , \new_[9915]_ , \new_[9916]_ ,
    \new_[9917]_ , \new_[9918]_ , \new_[9919]_ , \new_[9920]_ ,
    \new_[9921]_ , \new_[9922]_ , \new_[9923]_ , \new_[9924]_ ,
    \new_[9925]_ , \new_[9926]_ , \new_[9927]_ , \new_[9928]_ ,
    \new_[9929]_ , \new_[9930]_ , \new_[9931]_ , \new_[9932]_ ,
    \new_[9933]_ , \new_[9934]_ , \new_[9935]_ , \new_[9936]_ ,
    \new_[9937]_ , \new_[9938]_ , \new_[9939]_ , \new_[9940]_ ,
    \new_[9941]_ , \new_[9942]_ , \new_[9943]_ , \new_[9944]_ ,
    \new_[9945]_ , \new_[9946]_ , \new_[9947]_ , \new_[9948]_ ,
    \new_[9949]_ , \new_[9950]_ , \new_[9951]_ , \new_[9952]_ ,
    \new_[9953]_ , \new_[9954]_ , \new_[9955]_ , \new_[9956]_ ,
    \new_[9957]_ , \new_[9958]_ , \new_[9959]_ , \new_[9960]_ ,
    \new_[9961]_ , \new_[9962]_ , \new_[9963]_ , \new_[9964]_ ,
    \new_[9965]_ , \new_[9966]_ , \new_[9967]_ , \new_[9968]_ ,
    \new_[9969]_ , \new_[9970]_ , \new_[9971]_ , \new_[9972]_ ,
    \new_[9973]_ , \new_[9974]_ , \new_[9975]_ , \new_[9976]_ ,
    \new_[9977]_ , \new_[9978]_ , \new_[9979]_ , \new_[9980]_ ,
    \new_[9981]_ , \new_[9982]_ , \new_[9983]_ , \new_[9984]_ ,
    \new_[9985]_ , \new_[9986]_ , \new_[9987]_ , \new_[9988]_ ,
    \new_[9989]_ , \new_[9990]_ , \new_[9991]_ , \new_[9992]_ ,
    \new_[9993]_ , \new_[9994]_ , \new_[9995]_ , \new_[9996]_ ,
    \new_[9997]_ , \new_[9998]_ , \new_[9999]_ , \new_[10000]_ ,
    \new_[10001]_ , \new_[10002]_ , \new_[10003]_ , \new_[10004]_ ,
    \new_[10005]_ , \new_[10006]_ , \new_[10007]_ , \new_[10008]_ ,
    \new_[10009]_ , \new_[10010]_ , \new_[10011]_ , \new_[10012]_ ,
    \new_[10013]_ , \new_[10014]_ , \new_[10015]_ , \new_[10016]_ ,
    \new_[10017]_ , \new_[10018]_ , \new_[10019]_ , \new_[10020]_ ,
    \new_[10021]_ , \new_[10022]_ , \new_[10023]_ , \new_[10024]_ ,
    \new_[10025]_ , \new_[10026]_ , \new_[10027]_ , \new_[10028]_ ,
    \new_[10029]_ , \new_[10030]_ , \new_[10031]_ , \new_[10032]_ ,
    \new_[10033]_ , \new_[10034]_ , \new_[10035]_ , \new_[10036]_ ,
    \new_[10037]_ , \new_[10038]_ , \new_[10039]_ , \new_[10040]_ ,
    \new_[10041]_ , \new_[10042]_ , \new_[10043]_ , \new_[10044]_ ,
    \new_[10045]_ , \new_[10046]_ , \new_[10047]_ , \new_[10048]_ ,
    \new_[10049]_ , \new_[10050]_ , \new_[10051]_ , \new_[10052]_ ,
    \new_[10053]_ , \new_[10054]_ , \new_[10055]_ , \new_[10056]_ ,
    \new_[10057]_ , \new_[10058]_ , \new_[10059]_ , \new_[10060]_ ,
    \new_[10061]_ , \new_[10062]_ , \new_[10063]_ , \new_[10064]_ ,
    \new_[10065]_ , \new_[10066]_ , \new_[10067]_ , \new_[10068]_ ,
    \new_[10069]_ , \new_[10070]_ , \new_[10071]_ , \new_[10072]_ ,
    \new_[10073]_ , \new_[10074]_ , \new_[10075]_ , \new_[10076]_ ,
    \new_[10077]_ , \new_[10078]_ , \new_[10079]_ , \new_[10080]_ ,
    \new_[10081]_ , \new_[10082]_ , \new_[10083]_ , \new_[10084]_ ,
    \new_[10085]_ , \new_[10086]_ , \new_[10087]_ , \new_[10088]_ ,
    \new_[10089]_ , \new_[10090]_ , \new_[10091]_ , \new_[10092]_ ,
    \new_[10093]_ , \new_[10094]_ , \new_[10095]_ , \new_[10096]_ ,
    \new_[10097]_ , \new_[10098]_ , \new_[10099]_ , \new_[10100]_ ,
    \new_[10101]_ , \new_[10102]_ , \new_[10103]_ , \new_[10104]_ ,
    \new_[10105]_ , \new_[10106]_ , \new_[10107]_ , \new_[10108]_ ,
    \new_[10109]_ , \new_[10110]_ , \new_[10111]_ , \new_[10112]_ ,
    \new_[10113]_ , \new_[10114]_ , \new_[10115]_ , \new_[10116]_ ,
    \new_[10117]_ , \new_[10118]_ , \new_[10119]_ , \new_[10120]_ ,
    \new_[10121]_ , \new_[10122]_ , \new_[10123]_ , \new_[10124]_ ,
    \new_[10125]_ , \new_[10126]_ , \new_[10127]_ , \new_[10128]_ ,
    \new_[10129]_ , \new_[10130]_ , \new_[10131]_ , \new_[10132]_ ,
    \new_[10133]_ , \new_[10134]_ , \new_[10135]_ , \new_[10136]_ ,
    \new_[10137]_ , \new_[10138]_ , \new_[10139]_ , \new_[10140]_ ,
    \new_[10141]_ , \new_[10142]_ , \new_[10143]_ , \new_[10144]_ ,
    \new_[10145]_ , \new_[10146]_ , \new_[10147]_ , \new_[10148]_ ,
    \new_[10149]_ , \new_[10150]_ , \new_[10151]_ , \new_[10152]_ ,
    \new_[10153]_ , \new_[10154]_ , \new_[10155]_ , \new_[10156]_ ,
    \new_[10157]_ , \new_[10158]_ , \new_[10159]_ , \new_[10160]_ ,
    \new_[10161]_ , \new_[10162]_ , \new_[10163]_ , \new_[10164]_ ,
    \new_[10165]_ , \new_[10166]_ , \new_[10167]_ , \new_[10168]_ ,
    \new_[10169]_ , \new_[10170]_ , \new_[10171]_ , \new_[10172]_ ,
    \new_[10173]_ , \new_[10174]_ , \new_[10175]_ , \new_[10176]_ ,
    \new_[10177]_ , \new_[10178]_ , \new_[10179]_ , \new_[10180]_ ,
    \new_[10181]_ , \new_[10182]_ , \new_[10183]_ , \new_[10184]_ ,
    \new_[10185]_ , \new_[10186]_ , \new_[10187]_ , \new_[10188]_ ,
    \new_[10189]_ , \new_[10190]_ , \new_[10191]_ , \new_[10192]_ ,
    \new_[10193]_ , \new_[10194]_ , \new_[10195]_ , \new_[10196]_ ,
    \new_[10197]_ , \new_[10198]_ , \new_[10199]_ , \new_[10200]_ ,
    \new_[10201]_ , \new_[10202]_ , \new_[10203]_ , \new_[10204]_ ,
    \new_[10205]_ , \new_[10206]_ , \new_[10207]_ , \new_[10208]_ ,
    \new_[10209]_ , \new_[10210]_ , \new_[10211]_ , \new_[10212]_ ,
    \new_[10213]_ , \new_[10214]_ , \new_[10215]_ , \new_[10216]_ ,
    \new_[10217]_ , \new_[10218]_ , \new_[10219]_ , \new_[10220]_ ,
    \new_[10221]_ , \new_[10222]_ , \new_[10223]_ , \new_[10224]_ ,
    \new_[10225]_ , \new_[10226]_ , \new_[10227]_ , \new_[10228]_ ,
    \new_[10229]_ , \new_[10230]_ , \new_[10231]_ , \new_[10232]_ ,
    \new_[10233]_ , \new_[10234]_ , \new_[10235]_ , \new_[10236]_ ,
    \new_[10237]_ , \new_[10238]_ , \new_[10239]_ , \new_[10240]_ ,
    \new_[10241]_ , \new_[10242]_ , \new_[10243]_ , \new_[10244]_ ,
    \new_[10245]_ , \new_[10246]_ , \new_[10247]_ , \new_[10248]_ ,
    \new_[10249]_ , \new_[10250]_ , \new_[10251]_ , \new_[10252]_ ,
    \new_[10253]_ , \new_[10254]_ , \new_[10255]_ , \new_[10256]_ ,
    \new_[10257]_ , \new_[10258]_ , \new_[10259]_ , \new_[10260]_ ,
    \new_[10261]_ , \new_[10262]_ , \new_[10263]_ , \new_[10264]_ ,
    \new_[10265]_ , \new_[10266]_ , \new_[10267]_ , \new_[10268]_ ,
    \new_[10269]_ , \new_[10270]_ , \new_[10271]_ , \new_[10272]_ ,
    \new_[10273]_ , \new_[10274]_ , \new_[10275]_ , \new_[10276]_ ,
    \new_[10277]_ , \new_[10278]_ , \new_[10279]_ , \new_[10280]_ ,
    \new_[10281]_ , \new_[10282]_ , \new_[10283]_ , \new_[10284]_ ,
    \new_[10285]_ , \new_[10286]_ , \new_[10287]_ , \new_[10288]_ ,
    \new_[10289]_ , \new_[10290]_ , \new_[10291]_ , \new_[10292]_ ,
    \new_[10293]_ , \new_[10294]_ , \new_[10295]_ , \new_[10296]_ ,
    \new_[10297]_ , \new_[10298]_ , \new_[10299]_ , \new_[10300]_ ,
    \new_[10301]_ , \new_[10302]_ , \new_[10303]_ , \new_[10304]_ ,
    \new_[10305]_ , \new_[10306]_ , \new_[10307]_ , \new_[10308]_ ,
    \new_[10309]_ , \new_[10310]_ , \new_[10311]_ , \new_[10312]_ ,
    \new_[10313]_ , \new_[10314]_ , \new_[10315]_ , \new_[10316]_ ,
    \new_[10317]_ , \new_[10318]_ , \new_[10319]_ , \new_[10320]_ ,
    \new_[10321]_ , \new_[10322]_ , \new_[10323]_ , \new_[10324]_ ,
    \new_[10325]_ , \new_[10326]_ , \new_[10327]_ , \new_[10328]_ ,
    \new_[10329]_ , \new_[10330]_ , \new_[10331]_ , \new_[10332]_ ,
    \new_[10333]_ , \new_[10334]_ , \new_[10335]_ , \new_[10336]_ ,
    \new_[10337]_ , \new_[10338]_ , \new_[10339]_ , \new_[10340]_ ,
    \new_[10341]_ , \new_[10342]_ , \new_[10343]_ , \new_[10344]_ ,
    \new_[10345]_ , \new_[10346]_ , \new_[10347]_ , \new_[10348]_ ,
    \new_[10349]_ , \new_[10350]_ , \new_[10351]_ , \new_[10352]_ ,
    \new_[10353]_ , \new_[10354]_ , \new_[10355]_ , \new_[10356]_ ,
    \new_[10357]_ , \new_[10358]_ , \new_[10359]_ , \new_[10360]_ ,
    \new_[10361]_ , \new_[10362]_ , \new_[10363]_ , \new_[10364]_ ,
    \new_[10365]_ , \new_[10366]_ , \new_[10367]_ , \new_[10368]_ ,
    \new_[10369]_ , \new_[10370]_ , \new_[10371]_ , \new_[10372]_ ,
    \new_[10373]_ , \new_[10374]_ , \new_[10375]_ , \new_[10376]_ ,
    \new_[10377]_ , \new_[10378]_ , \new_[10379]_ , \new_[10380]_ ,
    \new_[10381]_ , \new_[10382]_ , \new_[10383]_ , \new_[10384]_ ,
    \new_[10385]_ , \new_[10386]_ , \new_[10387]_ , \new_[10388]_ ,
    \new_[10389]_ , \new_[10390]_ , \new_[10391]_ , \new_[10392]_ ,
    \new_[10393]_ , \new_[10394]_ , \new_[10395]_ , \new_[10396]_ ,
    \new_[10397]_ , \new_[10398]_ , \new_[10399]_ , \new_[10400]_ ,
    \new_[10401]_ , \new_[10402]_ , \new_[10403]_ , \new_[10404]_ ,
    \new_[10405]_ , \new_[10406]_ , \new_[10407]_ , \new_[10408]_ ,
    \new_[10409]_ , \new_[10410]_ , \new_[10411]_ , \new_[10412]_ ,
    \new_[10413]_ , \new_[10414]_ , \new_[10415]_ , \new_[10416]_ ,
    \new_[10417]_ , \new_[10418]_ , \new_[10419]_ , \new_[10420]_ ,
    \new_[10421]_ , \new_[10422]_ , \new_[10423]_ , \new_[10424]_ ,
    \new_[10425]_ , \new_[10426]_ , \new_[10427]_ , \new_[10428]_ ,
    \new_[10429]_ , \new_[10430]_ , \new_[10431]_ , \new_[10432]_ ,
    \new_[10433]_ , \new_[10434]_ , \new_[10435]_ , \new_[10436]_ ,
    \new_[10437]_ , \new_[10438]_ , \new_[10439]_ , \new_[10440]_ ,
    \new_[10441]_ , \new_[10442]_ , \new_[10443]_ , \new_[10444]_ ,
    \new_[10445]_ , \new_[10446]_ , \new_[10447]_ , \new_[10448]_ ,
    \new_[10449]_ , \new_[10450]_ , \new_[10451]_ , \new_[10452]_ ,
    \new_[10453]_ , \new_[10454]_ , \new_[10455]_ , \new_[10456]_ ,
    \new_[10457]_ , \new_[10458]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10462]_ , \new_[10463]_ , \new_[10464]_ ,
    \new_[10465]_ , \new_[10466]_ , \new_[10467]_ , \new_[10468]_ ,
    \new_[10469]_ , \new_[10470]_ , \new_[10471]_ , \new_[10472]_ ,
    \new_[10473]_ , \new_[10474]_ , \new_[10475]_ , \new_[10476]_ ,
    \new_[10477]_ , \new_[10478]_ , \new_[10479]_ , \new_[10480]_ ,
    \new_[10481]_ , \new_[10482]_ , \new_[10483]_ , \new_[10484]_ ,
    \new_[10485]_ , \new_[10486]_ , \new_[10487]_ , \new_[10488]_ ,
    \new_[10489]_ , \new_[10490]_ , \new_[10491]_ , \new_[10492]_ ,
    \new_[10493]_ , \new_[10494]_ , \new_[10495]_ , \new_[10496]_ ,
    \new_[10497]_ , \new_[10498]_ , \new_[10499]_ , \new_[10500]_ ,
    \new_[10501]_ , \new_[10502]_ , \new_[10503]_ , \new_[10504]_ ,
    \new_[10505]_ , \new_[10506]_ , \new_[10507]_ , \new_[10508]_ ,
    \new_[10509]_ , \new_[10510]_ , \new_[10511]_ , \new_[10512]_ ,
    \new_[10513]_ , \new_[10514]_ , \new_[10515]_ , \new_[10516]_ ,
    \new_[10517]_ , \new_[10518]_ , \new_[10519]_ , \new_[10520]_ ,
    \new_[10521]_ , \new_[10522]_ , \new_[10523]_ , \new_[10524]_ ,
    \new_[10525]_ , \new_[10526]_ , \new_[10527]_ , \new_[10528]_ ,
    \new_[10529]_ , \new_[10530]_ , \new_[10531]_ , \new_[10532]_ ,
    \new_[10533]_ , \new_[10534]_ , \new_[10535]_ , \new_[10536]_ ,
    \new_[10537]_ , \new_[10538]_ , \new_[10539]_ , \new_[10540]_ ,
    \new_[10541]_ , \new_[10542]_ , \new_[10543]_ , \new_[10544]_ ,
    \new_[10545]_ , \new_[10546]_ , \new_[10547]_ , \new_[10548]_ ,
    \new_[10549]_ , \new_[10550]_ , \new_[10551]_ , \new_[10552]_ ,
    \new_[10553]_ , \new_[10554]_ , \new_[10555]_ , \new_[10556]_ ,
    \new_[10557]_ , \new_[10558]_ , \new_[10559]_ , \new_[10560]_ ,
    \new_[10561]_ , \new_[10562]_ , \new_[10563]_ , \new_[10564]_ ,
    \new_[10565]_ , \new_[10566]_ , \new_[10567]_ , \new_[10568]_ ,
    \new_[10569]_ , \new_[10570]_ , \new_[10571]_ , \new_[10572]_ ,
    \new_[10573]_ , \new_[10574]_ , \new_[10575]_ , \new_[10576]_ ,
    \new_[10577]_ , \new_[10578]_ , \new_[10579]_ , \new_[10580]_ ,
    \new_[10581]_ , \new_[10582]_ , \new_[10583]_ , \new_[10584]_ ,
    \new_[10585]_ , \new_[10586]_ , \new_[10587]_ , \new_[10588]_ ,
    \new_[10589]_ , \new_[10590]_ , \new_[10591]_ , \new_[10592]_ ,
    \new_[10593]_ , \new_[10594]_ , \new_[10595]_ , \new_[10596]_ ,
    \new_[10597]_ , \new_[10598]_ , \new_[10599]_ , \new_[10600]_ ,
    \new_[10601]_ , \new_[10602]_ , \new_[10603]_ , \new_[10604]_ ,
    \new_[10605]_ , \new_[10606]_ , \new_[10607]_ , \new_[10608]_ ,
    \new_[10609]_ , \new_[10610]_ , \new_[10611]_ , \new_[10612]_ ,
    \new_[10613]_ , \new_[10614]_ , \new_[10615]_ , \new_[10616]_ ,
    \new_[10617]_ , \new_[10618]_ , \new_[10619]_ , \new_[10620]_ ,
    \new_[10621]_ , \new_[10622]_ , \new_[10623]_ , \new_[10624]_ ,
    \new_[10625]_ , \new_[10626]_ , \new_[10627]_ , \new_[10628]_ ,
    \new_[10629]_ , \new_[10630]_ , \new_[10631]_ , \new_[10632]_ ,
    \new_[10633]_ , \new_[10634]_ , \new_[10635]_ , \new_[10636]_ ,
    \new_[10637]_ , \new_[10638]_ , \new_[10639]_ , \new_[10640]_ ,
    \new_[10641]_ , \new_[10642]_ , \new_[10643]_ , \new_[10644]_ ,
    \new_[10645]_ , \new_[10646]_ , \new_[10647]_ , \new_[10648]_ ,
    \new_[10649]_ , \new_[10650]_ , \new_[10651]_ , \new_[10652]_ ,
    \new_[10653]_ , \new_[10654]_ , \new_[10655]_ , \new_[10656]_ ,
    \new_[10657]_ , \new_[10658]_ , \new_[10659]_ , \new_[10660]_ ,
    \new_[10661]_ , \new_[10662]_ , \new_[10663]_ , \new_[10664]_ ,
    \new_[10665]_ , \new_[10666]_ , \new_[10667]_ , \new_[10668]_ ,
    \new_[10669]_ , \new_[10670]_ , \new_[10671]_ , \new_[10672]_ ,
    \new_[10673]_ , \new_[10674]_ , \new_[10675]_ , \new_[10676]_ ,
    \new_[10677]_ , \new_[10678]_ , \new_[10679]_ , \new_[10680]_ ,
    \new_[10681]_ , \new_[10682]_ , \new_[10683]_ , \new_[10684]_ ,
    \new_[10685]_ , \new_[10686]_ , \new_[10687]_ , \new_[10688]_ ,
    \new_[10689]_ , \new_[10690]_ , \new_[10691]_ , \new_[10692]_ ,
    \new_[10693]_ , \new_[10694]_ , \new_[10695]_ , \new_[10696]_ ,
    \new_[10697]_ , \new_[10698]_ , \new_[10699]_ , \new_[10700]_ ,
    \new_[10701]_ , \new_[10702]_ , \new_[10703]_ , \new_[10704]_ ,
    \new_[10705]_ , \new_[10706]_ , \new_[10707]_ , \new_[10708]_ ,
    \new_[10709]_ , \new_[10710]_ , \new_[10711]_ , \new_[10712]_ ,
    \new_[10713]_ , \new_[10714]_ , \new_[10715]_ , \new_[10716]_ ,
    \new_[10717]_ , \new_[10718]_ , \new_[10719]_ , \new_[10720]_ ,
    \new_[10721]_ , \new_[10722]_ , \new_[10723]_ , \new_[10724]_ ,
    \new_[10725]_ , \new_[10726]_ , \new_[10727]_ , \new_[10728]_ ,
    \new_[10729]_ , \new_[10730]_ , \new_[10731]_ , \new_[10732]_ ,
    \new_[10733]_ , \new_[10734]_ , \new_[10735]_ , \new_[10736]_ ,
    \new_[10737]_ , \new_[10738]_ , \new_[10739]_ , \new_[10740]_ ,
    \new_[10741]_ , \new_[10742]_ , \new_[10743]_ , \new_[10744]_ ,
    \new_[10745]_ , \new_[10746]_ , \new_[10747]_ , \new_[10748]_ ,
    \new_[10749]_ , \new_[10750]_ , \new_[10751]_ , \new_[10752]_ ,
    \new_[10753]_ , \new_[10754]_ , \new_[10755]_ , \new_[10756]_ ,
    \new_[10757]_ , \new_[10758]_ , \new_[10759]_ , \new_[10760]_ ,
    \new_[10761]_ , \new_[10762]_ , \new_[10763]_ , \new_[10764]_ ,
    \new_[10765]_ , \new_[10766]_ , \new_[10767]_ , \new_[10768]_ ,
    \new_[10769]_ , \new_[10770]_ , \new_[10771]_ , \new_[10772]_ ,
    \new_[10773]_ , \new_[10774]_ , \new_[10775]_ , \new_[10776]_ ,
    \new_[10777]_ , \new_[10778]_ , \new_[10779]_ , \new_[10780]_ ,
    \new_[10781]_ , \new_[10782]_ , \new_[10783]_ , \new_[10784]_ ,
    \new_[10785]_ , \new_[10786]_ , \new_[10787]_ , \new_[10788]_ ,
    \new_[10789]_ , \new_[10790]_ , \new_[10791]_ , \new_[10792]_ ,
    \new_[10793]_ , \new_[10794]_ , \new_[10795]_ , \new_[10796]_ ,
    \new_[10797]_ , \new_[10798]_ , \new_[10799]_ , \new_[10800]_ ,
    \new_[10801]_ , \new_[10802]_ , \new_[10803]_ , \new_[10804]_ ,
    \new_[10805]_ , \new_[10806]_ , \new_[10807]_ , \new_[10808]_ ,
    \new_[10809]_ , \new_[10810]_ , \new_[10811]_ , \new_[10812]_ ,
    \new_[10813]_ , \new_[10814]_ , \new_[10815]_ , \new_[10816]_ ,
    \new_[10817]_ , \new_[10818]_ , \new_[10819]_ , \new_[10820]_ ,
    \new_[10821]_ , \new_[10822]_ , \new_[10823]_ , \new_[10824]_ ,
    \new_[10825]_ , \new_[10826]_ , \new_[10827]_ , \new_[10828]_ ,
    \new_[10829]_ , \new_[10830]_ , \new_[10831]_ , \new_[10832]_ ,
    \new_[10833]_ , \new_[10834]_ , \new_[10835]_ , \new_[10836]_ ,
    \new_[10837]_ , \new_[10838]_ , \new_[10839]_ , \new_[10840]_ ,
    \new_[10841]_ , \new_[10842]_ , \new_[10843]_ , \new_[10844]_ ,
    \new_[10845]_ , \new_[10846]_ , \new_[10847]_ , \new_[10848]_ ,
    \new_[10849]_ , \new_[10850]_ , \new_[10851]_ , \new_[10852]_ ,
    \new_[10853]_ , \new_[10854]_ , \new_[10855]_ , \new_[10856]_ ,
    \new_[10857]_ , \new_[10858]_ , \new_[10859]_ , \new_[10860]_ ,
    \new_[10861]_ , \new_[10862]_ , \new_[10863]_ , \new_[10864]_ ,
    \new_[10865]_ , \new_[10866]_ , \new_[10867]_ , \new_[10868]_ ,
    \new_[10869]_ , \new_[10870]_ , \new_[10871]_ , \new_[10872]_ ,
    \new_[10873]_ , \new_[10874]_ , \new_[10875]_ , \new_[10876]_ ,
    \new_[10877]_ , \new_[10878]_ , \new_[10879]_ , \new_[10880]_ ,
    \new_[10881]_ , \new_[10882]_ , \new_[10883]_ , \new_[10884]_ ,
    \new_[10885]_ , \new_[10886]_ , \new_[10887]_ , \new_[10888]_ ,
    \new_[10889]_ , \new_[10890]_ , \new_[10891]_ , \new_[10892]_ ,
    \new_[10893]_ , \new_[10894]_ , \new_[10895]_ , \new_[10896]_ ,
    \new_[10897]_ , \new_[10898]_ , \new_[10899]_ , \new_[10900]_ ,
    \new_[10901]_ , \new_[10902]_ , \new_[10903]_ , \new_[10904]_ ,
    \new_[10905]_ , \new_[10906]_ , \new_[10907]_ , \new_[10908]_ ,
    \new_[10909]_ , \new_[10910]_ , \new_[10911]_ , \new_[10912]_ ,
    \new_[10913]_ , \new_[10914]_ , \new_[10915]_ , \new_[10916]_ ,
    \new_[10917]_ , \new_[10918]_ , \new_[10919]_ , \new_[10920]_ ,
    \new_[10921]_ , \new_[10922]_ , \new_[10923]_ , \new_[10924]_ ,
    \new_[10925]_ , \new_[10926]_ , \new_[10927]_ , \new_[10928]_ ,
    \new_[10929]_ , \new_[10930]_ , \new_[10931]_ , \new_[10932]_ ,
    \new_[10933]_ , \new_[10934]_ , \new_[10935]_ , \new_[10936]_ ,
    \new_[10937]_ , \new_[10938]_ , \new_[10939]_ , \new_[10940]_ ,
    \new_[10941]_ , \new_[10942]_ , \new_[10943]_ , \new_[10944]_ ,
    \new_[10945]_ , \new_[10946]_ , \new_[10947]_ , \new_[10948]_ ,
    \new_[10949]_ , \new_[10950]_ , \new_[10951]_ , \new_[10952]_ ,
    \new_[10953]_ , \new_[10954]_ , \new_[10955]_ , \new_[10956]_ ,
    \new_[10957]_ , \new_[10958]_ , \new_[10959]_ , \new_[10960]_ ,
    \new_[10961]_ , \new_[10962]_ , \new_[10963]_ , \new_[10964]_ ,
    \new_[10965]_ , \new_[10966]_ , \new_[10967]_ , \new_[10968]_ ,
    \new_[10969]_ , \new_[10970]_ , \new_[10971]_ , \new_[10972]_ ,
    \new_[10973]_ , \new_[10974]_ , \new_[10975]_ , \new_[10976]_ ,
    \new_[10977]_ , \new_[10978]_ , \new_[10979]_ , \new_[10980]_ ,
    \new_[10981]_ , \new_[10982]_ , \new_[10983]_ , \new_[10984]_ ,
    \new_[10985]_ , \new_[10986]_ , \new_[10987]_ , \new_[10988]_ ,
    \new_[10989]_ , \new_[10990]_ , \new_[10991]_ , \new_[10992]_ ,
    \new_[10993]_ , \new_[10994]_ , \new_[10995]_ , \new_[10996]_ ,
    \new_[10997]_ , \new_[10998]_ , \new_[10999]_ , \new_[11000]_ ,
    \new_[11001]_ , \new_[11002]_ , \new_[11003]_ , \new_[11004]_ ,
    \new_[11005]_ , \new_[11006]_ , \new_[11007]_ , \new_[11008]_ ,
    \new_[11009]_ , \new_[11010]_ , \new_[11011]_ , \new_[11012]_ ,
    \new_[11013]_ , \new_[11014]_ , \new_[11015]_ , \new_[11016]_ ,
    \new_[11017]_ , \new_[11018]_ , \new_[11019]_ , \new_[11020]_ ,
    \new_[11021]_ , \new_[11022]_ , \new_[11023]_ , \new_[11024]_ ,
    \new_[11025]_ , \new_[11026]_ , \new_[11027]_ , \new_[11028]_ ,
    \new_[11029]_ , \new_[11030]_ , \new_[11031]_ , \new_[11032]_ ,
    \new_[11033]_ , \new_[11034]_ , \new_[11035]_ , \new_[11036]_ ,
    \new_[11037]_ , \new_[11038]_ , \new_[11039]_ , \new_[11040]_ ,
    \new_[11041]_ , \new_[11042]_ , \new_[11043]_ , \new_[11044]_ ,
    \new_[11045]_ , \new_[11046]_ , \new_[11047]_ , \new_[11048]_ ,
    \new_[11049]_ , \new_[11050]_ , \new_[11051]_ , \new_[11052]_ ,
    \new_[11053]_ , \new_[11054]_ , \new_[11055]_ , \new_[11056]_ ,
    \new_[11057]_ , \new_[11058]_ , \new_[11059]_ , \new_[11060]_ ,
    \new_[11061]_ , \new_[11062]_ , \new_[11063]_ , \new_[11064]_ ,
    \new_[11065]_ , \new_[11066]_ , \new_[11067]_ , \new_[11068]_ ,
    \new_[11069]_ , \new_[11070]_ , \new_[11071]_ , \new_[11072]_ ,
    \new_[11073]_ , \new_[11074]_ , \new_[11075]_ , \new_[11076]_ ,
    \new_[11077]_ , \new_[11078]_ , \new_[11079]_ , \new_[11080]_ ,
    \new_[11081]_ , \new_[11082]_ , \new_[11083]_ , \new_[11084]_ ,
    \new_[11085]_ , \new_[11086]_ , \new_[11087]_ , \new_[11088]_ ,
    \new_[11089]_ , \new_[11090]_ , \new_[11091]_ , \new_[11092]_ ,
    \new_[11093]_ , \new_[11094]_ , \new_[11095]_ , \new_[11096]_ ,
    \new_[11097]_ , \new_[11098]_ , \new_[11099]_ , \new_[11100]_ ,
    \new_[11101]_ , \new_[11102]_ , \new_[11103]_ , \new_[11104]_ ,
    \new_[11105]_ , \new_[11106]_ , \new_[11107]_ , \new_[11108]_ ,
    \new_[11109]_ , \new_[11110]_ , \new_[11111]_ , \new_[11112]_ ,
    \new_[11113]_ , \new_[11114]_ , \new_[11115]_ , \new_[11116]_ ,
    \new_[11117]_ , \new_[11118]_ , \new_[11119]_ , \new_[11120]_ ,
    \new_[11121]_ , \new_[11122]_ , \new_[11123]_ , \new_[11124]_ ,
    \new_[11125]_ , \new_[11126]_ , \new_[11127]_ , \new_[11128]_ ,
    \new_[11129]_ , \new_[11130]_ , \new_[11131]_ , \new_[11132]_ ,
    \new_[11133]_ , \new_[11134]_ , \new_[11135]_ , \new_[11136]_ ,
    \new_[11137]_ , \new_[11138]_ , \new_[11139]_ , \new_[11140]_ ,
    \new_[11141]_ , \new_[11142]_ , \new_[11143]_ , \new_[11144]_ ,
    \new_[11145]_ , \new_[11146]_ , \new_[11147]_ , \new_[11148]_ ,
    \new_[11149]_ , \new_[11150]_ , \new_[11151]_ , \new_[11152]_ ,
    \new_[11153]_ , \new_[11154]_ , \new_[11155]_ , \new_[11156]_ ,
    \new_[11157]_ , \new_[11158]_ , \new_[11159]_ , \new_[11160]_ ,
    \new_[11161]_ , \new_[11162]_ , \new_[11163]_ , \new_[11164]_ ,
    \new_[11165]_ , \new_[11166]_ , \new_[11167]_ , \new_[11168]_ ,
    \new_[11169]_ , \new_[11170]_ , \new_[11171]_ , \new_[11172]_ ,
    \new_[11173]_ , \new_[11174]_ , \new_[11175]_ , \new_[11176]_ ,
    \new_[11177]_ , \new_[11178]_ , \new_[11179]_ , \new_[11180]_ ,
    \new_[11181]_ , \new_[11182]_ , \new_[11183]_ , \new_[11184]_ ,
    \new_[11185]_ , \new_[11186]_ , \new_[11187]_ , \new_[11188]_ ,
    \new_[11189]_ , \new_[11190]_ , \new_[11191]_ , \new_[11192]_ ,
    \new_[11193]_ , \new_[11194]_ , \new_[11195]_ , \new_[11196]_ ,
    \new_[11197]_ , \new_[11198]_ , \new_[11199]_ , \new_[11200]_ ,
    \new_[11201]_ , \new_[11202]_ , \new_[11203]_ , \new_[11204]_ ,
    \new_[11205]_ , \new_[11206]_ , \new_[11207]_ , \new_[11208]_ ,
    \new_[11209]_ , \new_[11210]_ , \new_[11211]_ , \new_[11212]_ ,
    \new_[11213]_ , \new_[11214]_ , \new_[11215]_ , \new_[11216]_ ,
    \new_[11217]_ , \new_[11218]_ , \new_[11219]_ , \new_[11220]_ ,
    \new_[11221]_ , \new_[11222]_ , \new_[11223]_ , \new_[11224]_ ,
    \new_[11225]_ , \new_[11226]_ , \new_[11227]_ , \new_[11228]_ ,
    \new_[11229]_ , \new_[11230]_ , \new_[11231]_ , \new_[11232]_ ,
    \new_[11233]_ , \new_[11234]_ , \new_[11235]_ , \new_[11236]_ ,
    \new_[11237]_ , \new_[11238]_ , \new_[11239]_ , \new_[11240]_ ,
    \new_[11241]_ , \new_[11242]_ , \new_[11243]_ , \new_[11244]_ ,
    \new_[11245]_ , \new_[11246]_ , \new_[11247]_ , \new_[11248]_ ,
    \new_[11249]_ , \new_[11250]_ , \new_[11251]_ , \new_[11252]_ ,
    \new_[11253]_ , \new_[11254]_ , \new_[11255]_ , \new_[11256]_ ,
    \new_[11257]_ , \new_[11258]_ , \new_[11259]_ , \new_[11260]_ ,
    \new_[11261]_ , \new_[11262]_ , \new_[11263]_ , \new_[11264]_ ,
    \new_[11265]_ , \new_[11266]_ , \new_[11267]_ , \new_[11268]_ ,
    \new_[11269]_ , \new_[11270]_ , \new_[11271]_ , \new_[11272]_ ,
    \new_[11273]_ , \new_[11274]_ , \new_[11275]_ , \new_[11276]_ ,
    \new_[11277]_ , \new_[11278]_ , \new_[11279]_ , \new_[11280]_ ,
    \new_[11281]_ , \new_[11282]_ , \new_[11283]_ , \new_[11284]_ ,
    \new_[11285]_ , \new_[11286]_ , \new_[11287]_ , \new_[11288]_ ,
    \new_[11289]_ , \new_[11290]_ , \new_[11291]_ , \new_[11292]_ ,
    \new_[11293]_ , \new_[11294]_ , \new_[11295]_ , \new_[11296]_ ,
    \new_[11297]_ , \new_[11298]_ , \new_[11299]_ , \new_[11300]_ ,
    \new_[11301]_ , \new_[11302]_ , \new_[11303]_ , \new_[11304]_ ,
    \new_[11305]_ , \new_[11306]_ , \new_[11307]_ , \new_[11308]_ ,
    \new_[11309]_ , \new_[11310]_ , \new_[11311]_ , \new_[11312]_ ,
    \new_[11313]_ , \new_[11314]_ , \new_[11315]_ , \new_[11316]_ ,
    \new_[11317]_ , \new_[11318]_ , \new_[11319]_ , \new_[11320]_ ,
    \new_[11321]_ , \new_[11322]_ , \new_[11323]_ , \new_[11324]_ ,
    \new_[11325]_ , \new_[11326]_ , \new_[11327]_ , \new_[11328]_ ,
    \new_[11329]_ , \new_[11330]_ , \new_[11331]_ , \new_[11332]_ ,
    \new_[11333]_ , \new_[11334]_ , \new_[11335]_ , \new_[11336]_ ,
    \new_[11337]_ , \new_[11338]_ , \new_[11339]_ , \new_[11340]_ ,
    \new_[11341]_ , \new_[11342]_ , \new_[11343]_ , \new_[11344]_ ,
    \new_[11345]_ , \new_[11346]_ , \new_[11347]_ , \new_[11348]_ ,
    \new_[11349]_ , \new_[11350]_ , \new_[11351]_ , \new_[11352]_ ,
    \new_[11353]_ , \new_[11354]_ , \new_[11355]_ , \new_[11356]_ ,
    \new_[11357]_ , \new_[11358]_ , \new_[11359]_ , \new_[11360]_ ,
    \new_[11361]_ , \new_[11362]_ , \new_[11363]_ , \new_[11364]_ ,
    \new_[11365]_ , \new_[11366]_ , \new_[11367]_ , \new_[11368]_ ,
    \new_[11369]_ , \new_[11370]_ , \new_[11371]_ , \new_[11372]_ ,
    \new_[11373]_ , \new_[11374]_ , \new_[11375]_ , \new_[11376]_ ,
    \new_[11377]_ , \new_[11378]_ , \new_[11379]_ , \new_[11380]_ ,
    \new_[11381]_ , \new_[11382]_ , \new_[11383]_ , \new_[11384]_ ,
    \new_[11385]_ , \new_[11386]_ , \new_[11387]_ , \new_[11388]_ ,
    \new_[11389]_ , \new_[11390]_ , \new_[11391]_ , \new_[11392]_ ,
    \new_[11393]_ , \new_[11394]_ , \new_[11395]_ , \new_[11396]_ ,
    \new_[11397]_ , \new_[11398]_ , \new_[11399]_ , \new_[11400]_ ,
    \new_[11401]_ , \new_[11402]_ , \new_[11403]_ , \new_[11404]_ ,
    \new_[11405]_ , \new_[11406]_ , \new_[11407]_ , \new_[11408]_ ,
    \new_[11409]_ , \new_[11410]_ , \new_[11411]_ , \new_[11412]_ ,
    \new_[11413]_ , \new_[11414]_ , \new_[11415]_ , \new_[11416]_ ,
    \new_[11417]_ , \new_[11418]_ , \new_[11419]_ , \new_[11420]_ ,
    \new_[11421]_ , \new_[11422]_ , \new_[11423]_ , \new_[11424]_ ,
    \new_[11425]_ , \new_[11426]_ , \new_[11427]_ , \new_[11428]_ ,
    \new_[11429]_ , \new_[11430]_ , \new_[11431]_ , \new_[11432]_ ,
    \new_[11433]_ , \new_[11434]_ , \new_[11435]_ , \new_[11436]_ ,
    \new_[11437]_ , \new_[11438]_ , \new_[11439]_ , \new_[11440]_ ,
    \new_[11441]_ , \new_[11442]_ , \new_[11443]_ , \new_[11444]_ ,
    \new_[11445]_ , \new_[11446]_ , \new_[11447]_ , \new_[11448]_ ,
    \new_[11449]_ , \new_[11450]_ , \new_[11451]_ , \new_[11452]_ ,
    \new_[11453]_ , \new_[11454]_ , \new_[11455]_ , \new_[11456]_ ,
    \new_[11457]_ , \new_[11458]_ , \new_[11459]_ , \new_[11460]_ ,
    \new_[11461]_ , \new_[11462]_ , \new_[11463]_ , \new_[11464]_ ,
    \new_[11465]_ , \new_[11466]_ , \new_[11467]_ , \new_[11468]_ ,
    \new_[11469]_ , \new_[11470]_ , \new_[11471]_ , \new_[11472]_ ,
    \new_[11473]_ , \new_[11474]_ , \new_[11475]_ , \new_[11476]_ ,
    \new_[11477]_ , \new_[11478]_ , \new_[11479]_ , \new_[11480]_ ,
    \new_[11481]_ , \new_[11482]_ , \new_[11483]_ , \new_[11484]_ ,
    \new_[11485]_ , \new_[11486]_ , \new_[11487]_ , \new_[11488]_ ,
    \new_[11489]_ , \new_[11490]_ , \new_[11491]_ , \new_[11492]_ ,
    \new_[11493]_ , \new_[11494]_ , \new_[11495]_ , \new_[11496]_ ,
    \new_[11497]_ , \new_[11498]_ , \new_[11499]_ , \new_[11500]_ ,
    \new_[11501]_ , \new_[11502]_ , \new_[11503]_ , \new_[11504]_ ,
    \new_[11505]_ , \new_[11506]_ , \new_[11507]_ , \new_[11508]_ ,
    \new_[11509]_ , \new_[11510]_ , \new_[11511]_ , \new_[11512]_ ,
    \new_[11513]_ , \new_[11514]_ , \new_[11515]_ , \new_[11516]_ ,
    \new_[11517]_ , \new_[11518]_ , \new_[11519]_ , \new_[11520]_ ,
    \new_[11521]_ , \new_[11522]_ , \new_[11523]_ , \new_[11524]_ ,
    \new_[11525]_ , \new_[11526]_ , \new_[11527]_ , \new_[11528]_ ,
    \new_[11529]_ , \new_[11530]_ , \new_[11531]_ , \new_[11532]_ ,
    \new_[11533]_ , \new_[11534]_ , \new_[11535]_ , \new_[11536]_ ,
    \new_[11537]_ , \new_[11538]_ , \new_[11539]_ , \new_[11540]_ ,
    \new_[11541]_ , \new_[11542]_ , \new_[11543]_ , \new_[11544]_ ,
    \new_[11545]_ , \new_[11546]_ , \new_[11547]_ , \new_[11548]_ ,
    \new_[11549]_ , \new_[11550]_ , \new_[11551]_ , \new_[11552]_ ,
    \new_[11553]_ , \new_[11554]_ , \new_[11555]_ , \new_[11556]_ ,
    \new_[11557]_ , \new_[11558]_ , \new_[11559]_ , \new_[11560]_ ,
    \new_[11561]_ , \new_[11562]_ , \new_[11563]_ , \new_[11564]_ ,
    \new_[11565]_ , \new_[11566]_ , \new_[11567]_ , \new_[11568]_ ,
    \new_[11569]_ , \new_[11570]_ , \new_[11571]_ , \new_[11572]_ ,
    \new_[11573]_ , \new_[11574]_ , \new_[11575]_ , \new_[11576]_ ,
    \new_[11577]_ , \new_[11578]_ , \new_[11579]_ , \new_[11580]_ ,
    \new_[11581]_ , \new_[11582]_ , \new_[11583]_ , \new_[11584]_ ,
    \new_[11585]_ , \new_[11586]_ , \new_[11587]_ , \new_[11588]_ ,
    \new_[11589]_ , \new_[11590]_ , \new_[11591]_ , \new_[11592]_ ,
    \new_[11593]_ , \new_[11594]_ , \new_[11595]_ , \new_[11596]_ ,
    \new_[11597]_ , \new_[11598]_ , \new_[11599]_ , \new_[11600]_ ,
    \new_[11601]_ , \new_[11602]_ , \new_[11603]_ , \new_[11604]_ ,
    \new_[11605]_ , \new_[11606]_ , \new_[11607]_ , \new_[11608]_ ,
    \new_[11609]_ , \new_[11610]_ , \new_[11611]_ , \new_[11612]_ ,
    \new_[11613]_ , \new_[11614]_ , \new_[11615]_ , \new_[11616]_ ,
    \new_[11617]_ , \new_[11618]_ , \new_[11619]_ , \new_[11620]_ ,
    \new_[11621]_ , \new_[11622]_ , \new_[11623]_ , \new_[11624]_ ,
    \new_[11625]_ , \new_[11626]_ , \new_[11627]_ , \new_[11628]_ ,
    \new_[11629]_ , \new_[11630]_ , \new_[11631]_ , \new_[11632]_ ,
    \new_[11633]_ , \new_[11634]_ , \new_[11635]_ , \new_[11636]_ ,
    \new_[11637]_ , \new_[11638]_ , \new_[11639]_ , \new_[11640]_ ,
    \new_[11641]_ , \new_[11642]_ , \new_[11643]_ , \new_[11644]_ ,
    \new_[11645]_ , \new_[11646]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11649]_ , \new_[11650]_ , \new_[11651]_ , \new_[11652]_ ,
    \new_[11653]_ , \new_[11654]_ , \new_[11655]_ , \new_[11656]_ ,
    \new_[11657]_ , \new_[11658]_ , \new_[11659]_ , \new_[11660]_ ,
    \new_[11661]_ , \new_[11662]_ , \new_[11663]_ , \new_[11664]_ ,
    \new_[11665]_ , \new_[11666]_ , \new_[11667]_ , \new_[11668]_ ,
    \new_[11669]_ , \new_[11670]_ , \new_[11671]_ , \new_[11672]_ ,
    \new_[11673]_ , \new_[11674]_ , \new_[11675]_ , \new_[11676]_ ,
    \new_[11677]_ , \new_[11678]_ , \new_[11679]_ , \new_[11680]_ ,
    \new_[11681]_ , \new_[11682]_ , \new_[11683]_ , \new_[11684]_ ,
    \new_[11685]_ , \new_[11686]_ , \new_[11687]_ , \new_[11688]_ ,
    \new_[11689]_ , \new_[11690]_ , \new_[11691]_ , \new_[11692]_ ,
    \new_[11693]_ , \new_[11694]_ , \new_[11695]_ , \new_[11696]_ ,
    \new_[11697]_ , \new_[11698]_ , \new_[11699]_ , \new_[11700]_ ,
    \new_[11701]_ , \new_[11702]_ , \new_[11703]_ , \new_[11704]_ ,
    \new_[11705]_ , \new_[11706]_ , \new_[11707]_ , \new_[11708]_ ,
    \new_[11709]_ , \new_[11710]_ , \new_[11711]_ , \new_[11712]_ ,
    \new_[11713]_ , \new_[11714]_ , \new_[11715]_ , \new_[11716]_ ,
    \new_[11717]_ , \new_[11718]_ , \new_[11719]_ , \new_[11720]_ ,
    \new_[11721]_ , \new_[11722]_ , \new_[11723]_ , \new_[11724]_ ,
    \new_[11725]_ , \new_[11726]_ , \new_[11727]_ , \new_[11728]_ ,
    \new_[11729]_ , \new_[11730]_ , \new_[11731]_ , \new_[11732]_ ,
    \new_[11733]_ , \new_[11734]_ , \new_[11735]_ , \new_[11736]_ ,
    \new_[11737]_ , \new_[11738]_ , \new_[11739]_ , \new_[11740]_ ,
    \new_[11741]_ , \new_[11742]_ , \new_[11743]_ , \new_[11744]_ ,
    \new_[11745]_ , \new_[11746]_ , \new_[11747]_ , \new_[11748]_ ,
    \new_[11749]_ , \new_[11750]_ , \new_[11751]_ , \new_[11752]_ ,
    \new_[11753]_ , \new_[11754]_ , \new_[11755]_ , \new_[11756]_ ,
    \new_[11757]_ , \new_[11758]_ , \new_[11759]_ , \new_[11760]_ ,
    \new_[11761]_ , \new_[11762]_ , \new_[11763]_ , \new_[11764]_ ,
    \new_[11765]_ , \new_[11766]_ , \new_[11767]_ , \new_[11768]_ ,
    \new_[11769]_ , \new_[11770]_ , \new_[11771]_ , \new_[11772]_ ,
    \new_[11773]_ , \new_[11774]_ , \new_[11775]_ , \new_[11776]_ ,
    \new_[11777]_ , \new_[11778]_ , \new_[11779]_ , \new_[11780]_ ,
    \new_[11781]_ , \new_[11782]_ , \new_[11783]_ , \new_[11784]_ ,
    \new_[11785]_ , \new_[11786]_ , \new_[11787]_ , \new_[11788]_ ,
    \new_[11789]_ , \new_[11790]_ , \new_[11791]_ , \new_[11792]_ ,
    \new_[11793]_ , \new_[11794]_ , \new_[11795]_ , \new_[11796]_ ,
    \new_[11797]_ , \new_[11798]_ , \new_[11799]_ , \new_[11800]_ ,
    \new_[11801]_ , \new_[11802]_ , \new_[11803]_ , \new_[11804]_ ,
    \new_[11805]_ , \new_[11806]_ , \new_[11807]_ , \new_[11808]_ ,
    \new_[11809]_ , \new_[11810]_ , \new_[11811]_ , \new_[11812]_ ,
    \new_[11813]_ , \new_[11814]_ , \new_[11815]_ , \new_[11816]_ ,
    \new_[11817]_ , \new_[11818]_ , \new_[11819]_ , \new_[11820]_ ,
    \new_[11821]_ , \new_[11822]_ , \new_[11823]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11826]_ , \new_[11827]_ , \new_[11828]_ ,
    \new_[11829]_ , \new_[11830]_ , \new_[11831]_ , \new_[11832]_ ,
    \new_[11833]_ , \new_[11834]_ , \new_[11835]_ , \new_[11836]_ ,
    \new_[11837]_ , \new_[11838]_ , \new_[11839]_ , \new_[11840]_ ,
    \new_[11841]_ , \new_[11842]_ , \new_[11843]_ , \new_[11844]_ ,
    \new_[11845]_ , \new_[11846]_ , \new_[11847]_ , \new_[11848]_ ,
    \new_[11849]_ , \new_[11850]_ , \new_[11851]_ , \new_[11852]_ ,
    \new_[11853]_ , \new_[11854]_ , \new_[11855]_ , \new_[11856]_ ,
    \new_[11857]_ , \new_[11858]_ , \new_[11859]_ , \new_[11860]_ ,
    \new_[11861]_ , \new_[11862]_ , \new_[11863]_ , \new_[11864]_ ,
    \new_[11865]_ , \new_[11866]_ , \new_[11867]_ , \new_[11868]_ ,
    \new_[11869]_ , \new_[11870]_ , \new_[11871]_ , \new_[11872]_ ,
    \new_[11873]_ , \new_[11874]_ , \new_[11875]_ , \new_[11876]_ ,
    \new_[11877]_ , \new_[11878]_ , \new_[11879]_ , \new_[11880]_ ,
    \new_[11881]_ , \new_[11882]_ , \new_[11883]_ , \new_[11884]_ ,
    \new_[11885]_ , \new_[11886]_ , \new_[11887]_ , \new_[11888]_ ,
    \new_[11889]_ , \new_[11890]_ , \new_[11891]_ , \new_[11892]_ ,
    \new_[11893]_ , \new_[11894]_ , \new_[11895]_ , \new_[11896]_ ,
    \new_[11897]_ , \new_[11898]_ , \new_[11899]_ , \new_[11900]_ ,
    \new_[11901]_ , \new_[11902]_ , \new_[11903]_ , \new_[11904]_ ,
    \new_[11905]_ , \new_[11906]_ , \new_[11907]_ , \new_[11908]_ ,
    \new_[11909]_ , \new_[11910]_ , \new_[11911]_ , \new_[11912]_ ,
    \new_[11913]_ , \new_[11914]_ , \new_[11915]_ , \new_[11916]_ ,
    \new_[11917]_ , \new_[11918]_ , \new_[11919]_ , \new_[11920]_ ,
    \new_[11921]_ , \new_[11922]_ , \new_[11923]_ , \new_[11924]_ ,
    \new_[11925]_ , \new_[11926]_ , \new_[11927]_ , \new_[11928]_ ,
    \new_[11929]_ , \new_[11930]_ , \new_[11931]_ , \new_[11932]_ ,
    \new_[11933]_ , \new_[11934]_ , \new_[11935]_ , \new_[11936]_ ,
    \new_[11937]_ , \new_[11938]_ , \new_[11939]_ , \new_[11940]_ ,
    \new_[11941]_ , \new_[11942]_ , \new_[11943]_ , \new_[11944]_ ,
    \new_[11945]_ , \new_[11946]_ , \new_[11947]_ , \new_[11948]_ ,
    \new_[11949]_ , \new_[11950]_ , \new_[11951]_ , \new_[11952]_ ,
    \new_[11953]_ , \new_[11954]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11957]_ , \new_[11958]_ , \new_[11959]_ , \new_[11960]_ ,
    \new_[11961]_ , \new_[11962]_ , \new_[11963]_ , \new_[11964]_ ,
    \new_[11965]_ , \new_[11966]_ , \new_[11967]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11971]_ , \new_[11972]_ ,
    \new_[11973]_ , \new_[11974]_ , \new_[11975]_ , \new_[11976]_ ,
    \new_[11977]_ , \new_[11978]_ , \new_[11979]_ , \new_[11980]_ ,
    \new_[11981]_ , \new_[11982]_ , \new_[11983]_ , \new_[11984]_ ,
    \new_[11985]_ , \new_[11986]_ , \new_[11987]_ , \new_[11988]_ ,
    \new_[11989]_ , \new_[11990]_ , \new_[11991]_ , \new_[11992]_ ,
    \new_[11993]_ , \new_[11994]_ , \new_[11995]_ , \new_[11996]_ ,
    \new_[11997]_ , \new_[11998]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12001]_ , \new_[12002]_ , \new_[12003]_ , \new_[12004]_ ,
    \new_[12005]_ , \new_[12006]_ , \new_[12007]_ , \new_[12008]_ ,
    \new_[12009]_ , \new_[12010]_ , \new_[12011]_ , \new_[12012]_ ,
    \new_[12013]_ , \new_[12014]_ , \new_[12015]_ , \new_[12016]_ ,
    \new_[12017]_ , \new_[12018]_ , \new_[12019]_ , \new_[12020]_ ,
    \new_[12021]_ , \new_[12022]_ , \new_[12023]_ , \new_[12024]_ ,
    \new_[12025]_ , \new_[12026]_ , \new_[12027]_ , \new_[12028]_ ,
    \new_[12029]_ , \new_[12030]_ , \new_[12031]_ , \new_[12032]_ ,
    \new_[12033]_ , \new_[12034]_ , \new_[12035]_ , \new_[12036]_ ,
    \new_[12037]_ , \new_[12038]_ , \new_[12039]_ , \new_[12040]_ ,
    \new_[12041]_ , \new_[12042]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12045]_ , \new_[12046]_ , \new_[12047]_ , \new_[12048]_ ,
    \new_[12049]_ , \new_[12050]_ , \new_[12051]_ , \new_[12052]_ ,
    \new_[12053]_ , \new_[12054]_ , \new_[12055]_ , \new_[12056]_ ,
    \new_[12057]_ , \new_[12058]_ , \new_[12059]_ , \new_[12060]_ ,
    \new_[12061]_ , \new_[12062]_ , \new_[12063]_ , \new_[12064]_ ,
    \new_[12065]_ , \new_[12066]_ , \new_[12067]_ , \new_[12068]_ ,
    \new_[12069]_ , \new_[12070]_ , \new_[12071]_ , \new_[12072]_ ,
    \new_[12073]_ , \new_[12074]_ , \new_[12075]_ , \new_[12076]_ ,
    \new_[12077]_ , \new_[12078]_ , \new_[12079]_ , \new_[12080]_ ,
    \new_[12081]_ , \new_[12082]_ , \new_[12083]_ , \new_[12084]_ ,
    \new_[12085]_ , \new_[12086]_ , \new_[12087]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12090]_ , \new_[12091]_ , \new_[12092]_ ,
    \new_[12093]_ , \new_[12094]_ , \new_[12095]_ , \new_[12096]_ ,
    \new_[12097]_ , \new_[12098]_ , \new_[12099]_ , \new_[12100]_ ,
    \new_[12101]_ , \new_[12102]_ , \new_[12103]_ , \new_[12104]_ ,
    \new_[12105]_ , \new_[12106]_ , \new_[12107]_ , \new_[12108]_ ,
    \new_[12109]_ , \new_[12110]_ , \new_[12111]_ , \new_[12112]_ ,
    \new_[12113]_ , \new_[12114]_ , \new_[12115]_ , \new_[12116]_ ,
    \new_[12117]_ , \new_[12118]_ , \new_[12119]_ , \new_[12120]_ ,
    \new_[12121]_ , \new_[12122]_ , \new_[12123]_ , \new_[12124]_ ,
    \new_[12125]_ , \new_[12126]_ , \new_[12127]_ , \new_[12128]_ ,
    \new_[12129]_ , \new_[12130]_ , \new_[12131]_ , \new_[12132]_ ,
    \new_[12133]_ , \new_[12134]_ , \new_[12135]_ , \new_[12136]_ ,
    \new_[12137]_ , \new_[12138]_ , \new_[12139]_ , \new_[12140]_ ,
    \new_[12141]_ , \new_[12142]_ , \new_[12143]_ , \new_[12144]_ ,
    \new_[12145]_ , \new_[12146]_ , \new_[12147]_ , \new_[12148]_ ,
    \new_[12149]_ , \new_[12150]_ , \new_[12151]_ , \new_[12152]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12155]_ , \new_[12156]_ ,
    \new_[12157]_ , \new_[12158]_ , \new_[12159]_ , \new_[12160]_ ,
    \new_[12161]_ , \new_[12162]_ , \new_[12163]_ , \new_[12164]_ ,
    \new_[12165]_ , \new_[12166]_ , \new_[12167]_ , \new_[12168]_ ,
    \new_[12169]_ , \new_[12170]_ , \new_[12171]_ , \new_[12172]_ ,
    \new_[12173]_ , \new_[12174]_ , \new_[12175]_ , \new_[12176]_ ,
    \new_[12177]_ , \new_[12178]_ , \new_[12179]_ , \new_[12180]_ ,
    \new_[12181]_ , \new_[12182]_ , \new_[12183]_ , \new_[12184]_ ,
    \new_[12185]_ , \new_[12186]_ , \new_[12187]_ , \new_[12188]_ ,
    \new_[12189]_ , \new_[12190]_ , \new_[12191]_ , \new_[12192]_ ,
    \new_[12193]_ , \new_[12194]_ , \new_[12195]_ , \new_[12196]_ ,
    \new_[12197]_ , \new_[12198]_ , \new_[12199]_ , \new_[12200]_ ,
    \new_[12201]_ , \new_[12202]_ , \new_[12203]_ , \new_[12204]_ ,
    \new_[12205]_ , \new_[12206]_ , \new_[12207]_ , \new_[12208]_ ,
    \new_[12209]_ , \new_[12210]_ , \new_[12211]_ , \new_[12212]_ ,
    \new_[12213]_ , \new_[12214]_ , \new_[12215]_ , \new_[12216]_ ,
    \new_[12217]_ , \new_[12218]_ , \new_[12219]_ , \new_[12220]_ ,
    \new_[12221]_ , \new_[12222]_ , \new_[12223]_ , \new_[12224]_ ,
    \new_[12225]_ , \new_[12226]_ , \new_[12227]_ , \new_[12228]_ ,
    \new_[12229]_ , \new_[12230]_ , \new_[12231]_ , \new_[12232]_ ,
    \new_[12233]_ , \new_[12234]_ , \new_[12235]_ , \new_[12236]_ ,
    \new_[12237]_ , \new_[12238]_ , \new_[12239]_ , \new_[12240]_ ,
    \new_[12241]_ , \new_[12242]_ , \new_[12243]_ , \new_[12244]_ ,
    \new_[12245]_ , \new_[12246]_ , \new_[12247]_ , \new_[12248]_ ,
    \new_[12249]_ , \new_[12250]_ , \new_[12251]_ , \new_[12252]_ ,
    \new_[12253]_ , \new_[12254]_ , \new_[12255]_ , \new_[12256]_ ,
    \new_[12257]_ , \new_[12258]_ , \new_[12259]_ , \new_[12260]_ ,
    \new_[12261]_ , \new_[12262]_ , \new_[12263]_ , \new_[12264]_ ,
    \new_[12265]_ , \new_[12266]_ , \new_[12267]_ , \new_[12268]_ ,
    \new_[12269]_ , \new_[12270]_ , \new_[12271]_ , \new_[12272]_ ,
    \new_[12273]_ , \new_[12274]_ , \new_[12275]_ , \new_[12276]_ ,
    \new_[12277]_ , \new_[12278]_ , \new_[12279]_ , \new_[12280]_ ,
    \new_[12281]_ , \new_[12282]_ , \new_[12283]_ , \new_[12284]_ ,
    \new_[12285]_ , \new_[12286]_ , \new_[12287]_ , \new_[12288]_ ,
    \new_[12289]_ , \new_[12290]_ , \new_[12291]_ , \new_[12292]_ ,
    \new_[12293]_ , \new_[12294]_ , \new_[12295]_ , \new_[12296]_ ,
    \new_[12297]_ , \new_[12298]_ , \new_[12299]_ , \new_[12300]_ ,
    \new_[12301]_ , \new_[12302]_ , \new_[12303]_ , \new_[12304]_ ,
    \new_[12305]_ , \new_[12306]_ , \new_[12307]_ , \new_[12308]_ ,
    \new_[12309]_ , \new_[12310]_ , \new_[12311]_ , \new_[12312]_ ,
    \new_[12313]_ , \new_[12314]_ , \new_[12315]_ , \new_[12316]_ ,
    \new_[12317]_ , \new_[12318]_ , \new_[12319]_ , \new_[12320]_ ,
    \new_[12321]_ , \new_[12322]_ , \new_[12323]_ , \new_[12324]_ ,
    \new_[12325]_ , \new_[12326]_ , \new_[12327]_ , \new_[12328]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12331]_ , \new_[12332]_ ,
    \new_[12333]_ , \new_[12334]_ , \new_[12335]_ , \new_[12336]_ ,
    \new_[12337]_ , \new_[12338]_ , \new_[12339]_ , \new_[12340]_ ,
    \new_[12341]_ , \new_[12342]_ , \new_[12343]_ , \new_[12344]_ ,
    \new_[12345]_ , \new_[12346]_ , \new_[12347]_ , \new_[12348]_ ,
    \new_[12349]_ , \new_[12350]_ , \new_[12351]_ , \new_[12352]_ ,
    \new_[12353]_ , \new_[12354]_ , \new_[12355]_ , \new_[12356]_ ,
    \new_[12357]_ , \new_[12358]_ , \new_[12359]_ , \new_[12360]_ ,
    \new_[12361]_ , \new_[12362]_ , \new_[12363]_ , \new_[12364]_ ,
    \new_[12365]_ , \new_[12366]_ , \new_[12367]_ , \new_[12368]_ ,
    \new_[12369]_ , \new_[12370]_ , \new_[12371]_ , \new_[12372]_ ,
    \new_[12373]_ , \new_[12374]_ , \new_[12375]_ , \new_[12376]_ ,
    \new_[12377]_ , \new_[12378]_ , \new_[12379]_ , \new_[12380]_ ,
    \new_[12381]_ , \new_[12382]_ , \new_[12383]_ , \new_[12384]_ ,
    \new_[12385]_ , \new_[12386]_ , \new_[12387]_ , \new_[12388]_ ,
    \new_[12389]_ , \new_[12390]_ , \new_[12391]_ , \new_[12392]_ ,
    \new_[12393]_ , \new_[12394]_ , \new_[12395]_ , \new_[12396]_ ,
    \new_[12397]_ , \new_[12398]_ , \new_[12399]_ , \new_[12400]_ ,
    \new_[12401]_ , \new_[12402]_ , \new_[12403]_ , \new_[12404]_ ,
    \new_[12405]_ , \new_[12406]_ , \new_[12407]_ , \new_[12408]_ ,
    \new_[12409]_ , \new_[12410]_ , \new_[12411]_ , \new_[12412]_ ,
    \new_[12413]_ , \new_[12414]_ , \new_[12415]_ , \new_[12416]_ ,
    \new_[12417]_ , \new_[12418]_ , \new_[12419]_ , \new_[12420]_ ,
    \new_[12421]_ , \new_[12422]_ , \new_[12423]_ , \new_[12424]_ ,
    \new_[12425]_ , \new_[12426]_ , \new_[12427]_ , \new_[12428]_ ,
    \new_[12429]_ , \new_[12430]_ , \new_[12431]_ , \new_[12432]_ ,
    \new_[12433]_ , \new_[12434]_ , \new_[12435]_ , \new_[12436]_ ,
    \new_[12437]_ , \new_[12438]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12442]_ , \new_[12443]_ , \new_[12444]_ ,
    \new_[12445]_ , \new_[12446]_ , \new_[12447]_ , \new_[12448]_ ,
    \new_[12449]_ , \new_[12450]_ , \new_[12451]_ , \new_[12452]_ ,
    \new_[12453]_ , \new_[12454]_ , \new_[12455]_ , \new_[12456]_ ,
    \new_[12457]_ , \new_[12458]_ , \new_[12459]_ , \new_[12460]_ ,
    \new_[12461]_ , \new_[12462]_ , \new_[12463]_ , \new_[12464]_ ,
    \new_[12465]_ , \new_[12466]_ , \new_[12467]_ , \new_[12468]_ ,
    \new_[12469]_ , \new_[12470]_ , \new_[12471]_ , \new_[12472]_ ,
    \new_[12473]_ , \new_[12474]_ , \new_[12475]_ , \new_[12476]_ ,
    \new_[12477]_ , \new_[12478]_ , \new_[12479]_ , \new_[12480]_ ,
    \new_[12481]_ , \new_[12482]_ , \new_[12483]_ , \new_[12484]_ ,
    \new_[12485]_ , \new_[12486]_ , \new_[12487]_ , \new_[12488]_ ,
    \new_[12489]_ , \new_[12490]_ , \new_[12491]_ , \new_[12492]_ ,
    \new_[12493]_ , \new_[12494]_ , \new_[12495]_ , \new_[12496]_ ,
    \new_[12497]_ , \new_[12498]_ , \new_[12499]_ , \new_[12500]_ ,
    \new_[12501]_ , \new_[12502]_ , \new_[12503]_ , \new_[12504]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12508]_ ,
    \new_[12509]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12513]_ , \new_[12514]_ , \new_[12515]_ , \new_[12516]_ ,
    \new_[12517]_ , \new_[12518]_ , \new_[12519]_ , \new_[12520]_ ,
    \new_[12521]_ , \new_[12522]_ , \new_[12523]_ , \new_[12524]_ ,
    \new_[12525]_ , \new_[12526]_ , \new_[12527]_ , \new_[12528]_ ,
    \new_[12529]_ , \new_[12530]_ , \new_[12531]_ , \new_[12532]_ ,
    \new_[12533]_ , \new_[12534]_ , \new_[12535]_ , \new_[12536]_ ,
    \new_[12537]_ , \new_[12538]_ , \new_[12539]_ , \new_[12540]_ ,
    \new_[12541]_ , \new_[12542]_ , \new_[12543]_ , \new_[12544]_ ,
    \new_[12545]_ , \new_[12546]_ , \new_[12547]_ , \new_[12548]_ ,
    \new_[12549]_ , \new_[12550]_ , \new_[12551]_ , \new_[12552]_ ,
    \new_[12553]_ , \new_[12554]_ , \new_[12555]_ , \new_[12556]_ ,
    \new_[12557]_ , \new_[12558]_ , \new_[12559]_ , \new_[12560]_ ,
    \new_[12561]_ , \new_[12562]_ , \new_[12563]_ , \new_[12564]_ ,
    \new_[12565]_ , \new_[12566]_ , \new_[12567]_ , \new_[12568]_ ,
    \new_[12569]_ , \new_[12570]_ , \new_[12571]_ , \new_[12572]_ ,
    \new_[12573]_ , \new_[12574]_ , \new_[12575]_ , \new_[12576]_ ,
    \new_[12577]_ , \new_[12578]_ , \new_[12579]_ , \new_[12580]_ ,
    \new_[12581]_ , \new_[12582]_ , \new_[12583]_ , \new_[12584]_ ,
    \new_[12585]_ , \new_[12586]_ , \new_[12587]_ , \new_[12588]_ ,
    \new_[12589]_ , \new_[12590]_ , \new_[12591]_ , \new_[12592]_ ,
    \new_[12593]_ , \new_[12594]_ , \new_[12595]_ , \new_[12596]_ ,
    \new_[12597]_ , \new_[12598]_ , \new_[12599]_ , \new_[12600]_ ,
    \new_[12601]_ , \new_[12602]_ , \new_[12603]_ , \new_[12604]_ ,
    \new_[12605]_ , \new_[12606]_ , \new_[12607]_ , \new_[12608]_ ,
    \new_[12609]_ , \new_[12610]_ , \new_[12611]_ , \new_[12612]_ ,
    \new_[12613]_ , \new_[12614]_ , \new_[12615]_ , \new_[12616]_ ,
    \new_[12617]_ , \new_[12618]_ , \new_[12619]_ , \new_[12620]_ ,
    \new_[12621]_ , \new_[12622]_ , \new_[12623]_ , \new_[12624]_ ,
    \new_[12625]_ , \new_[12626]_ , \new_[12627]_ , \new_[12628]_ ,
    \new_[12629]_ , \new_[12630]_ , \new_[12631]_ , \new_[12632]_ ,
    \new_[12633]_ , \new_[12634]_ , \new_[12635]_ , \new_[12636]_ ,
    \new_[12637]_ , \new_[12638]_ , \new_[12639]_ , \new_[12640]_ ,
    \new_[12641]_ , \new_[12642]_ , \new_[12643]_ , \new_[12644]_ ,
    \new_[12645]_ , \new_[12646]_ , \new_[12647]_ , \new_[12648]_ ,
    \new_[12649]_ , \new_[12650]_ , \new_[12651]_ , \new_[12652]_ ,
    \new_[12653]_ , \new_[12654]_ , \new_[12655]_ , \new_[12656]_ ,
    \new_[12657]_ , \new_[12658]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12661]_ , \new_[12662]_ , \new_[12663]_ , \new_[12664]_ ,
    \new_[12665]_ , \new_[12666]_ , \new_[12667]_ , \new_[12668]_ ,
    \new_[12669]_ , \new_[12670]_ , \new_[12671]_ , \new_[12672]_ ,
    \new_[12673]_ , \new_[12674]_ , \new_[12675]_ , \new_[12676]_ ,
    \new_[12677]_ , \new_[12678]_ , \new_[12679]_ , \new_[12680]_ ,
    \new_[12681]_ , \new_[12682]_ , \new_[12683]_ , \new_[12684]_ ,
    \new_[12685]_ , \new_[12686]_ , \new_[12687]_ , \new_[12688]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12691]_ , \new_[12692]_ ,
    \new_[12693]_ , \new_[12694]_ , \new_[12695]_ , \new_[12696]_ ,
    \new_[12697]_ , \new_[12698]_ , \new_[12699]_ , \new_[12700]_ ,
    \new_[12701]_ , \new_[12702]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12705]_ , \new_[12706]_ , \new_[12707]_ , \new_[12708]_ ,
    \new_[12709]_ , \new_[12710]_ , \new_[12711]_ , \new_[12712]_ ,
    \new_[12713]_ , \new_[12714]_ , \new_[12715]_ , \new_[12716]_ ,
    \new_[12717]_ , \new_[12718]_ , \new_[12719]_ , \new_[12720]_ ,
    \new_[12721]_ , \new_[12722]_ , \new_[12723]_ , \new_[12724]_ ,
    \new_[12725]_ , \new_[12726]_ , \new_[12727]_ , \new_[12728]_ ,
    \new_[12729]_ , \new_[12730]_ , \new_[12731]_ , \new_[12732]_ ,
    \new_[12733]_ , \new_[12734]_ , \new_[12735]_ , \new_[12736]_ ,
    \new_[12737]_ , \new_[12738]_ , \new_[12739]_ , \new_[12740]_ ,
    \new_[12741]_ , \new_[12742]_ , \new_[12743]_ , \new_[12744]_ ,
    \new_[12745]_ , \new_[12746]_ , \new_[12747]_ , \new_[12748]_ ,
    \new_[12749]_ , \new_[12750]_ , \new_[12751]_ , \new_[12752]_ ,
    \new_[12753]_ , \new_[12754]_ , \new_[12755]_ , \new_[12756]_ ,
    \new_[12757]_ , \new_[12758]_ , \new_[12759]_ , \new_[12760]_ ,
    \new_[12761]_ , \new_[12762]_ , \new_[12763]_ , \new_[12764]_ ,
    \new_[12765]_ , \new_[12766]_ , \new_[12767]_ , \new_[12768]_ ,
    \new_[12769]_ , \new_[12770]_ , \new_[12771]_ , \new_[12772]_ ,
    \new_[12773]_ , \new_[12774]_ , \new_[12775]_ , \new_[12776]_ ,
    \new_[12777]_ , \new_[12778]_ , \new_[12779]_ , \new_[12780]_ ,
    \new_[12781]_ , \new_[12782]_ , \new_[12783]_ , \new_[12784]_ ,
    \new_[12785]_ , \new_[12786]_ , \new_[12787]_ , \new_[12788]_ ,
    \new_[12789]_ , \new_[12790]_ , \new_[12791]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12794]_ , \new_[12795]_ , \new_[12796]_ ,
    \new_[12797]_ , \new_[12798]_ , \new_[12799]_ , \new_[12800]_ ,
    \new_[12801]_ , \new_[12802]_ , \new_[12803]_ , \new_[12804]_ ,
    \new_[12805]_ , \new_[12806]_ , \new_[12807]_ , \new_[12808]_ ,
    \new_[12809]_ , \new_[12810]_ , \new_[12811]_ , \new_[12812]_ ,
    \new_[12813]_ , \new_[12814]_ , \new_[12815]_ , \new_[12816]_ ,
    \new_[12817]_ , \new_[12818]_ , \new_[12819]_ , \new_[12820]_ ,
    \new_[12821]_ , \new_[12822]_ , \new_[12823]_ , \new_[12824]_ ,
    \new_[12825]_ , \new_[12826]_ , \new_[12827]_ , \new_[12828]_ ,
    \new_[12829]_ , \new_[12830]_ , \new_[12831]_ , \new_[12832]_ ,
    \new_[12833]_ , \new_[12834]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12837]_ , \new_[12838]_ , \new_[12839]_ , \new_[12840]_ ,
    \new_[12841]_ , \new_[12842]_ , \new_[12843]_ , \new_[12844]_ ,
    \new_[12845]_ , \new_[12846]_ , \new_[12847]_ , \new_[12848]_ ,
    \new_[12849]_ , \new_[12850]_ , \new_[12851]_ , \new_[12852]_ ,
    \new_[12853]_ , \new_[12854]_ , \new_[12855]_ , \new_[12856]_ ,
    \new_[12857]_ , \new_[12858]_ , \new_[12859]_ , \new_[12860]_ ,
    \new_[12861]_ , \new_[12862]_ , \new_[12863]_ , \new_[12864]_ ,
    \new_[12865]_ , \new_[12866]_ , \new_[12867]_ , \new_[12868]_ ,
    \new_[12869]_ , \new_[12870]_ , \new_[12871]_ , \new_[12872]_ ,
    \new_[12873]_ , \new_[12874]_ , \new_[12875]_ , \new_[12876]_ ,
    \new_[12877]_ , \new_[12878]_ , \new_[12879]_ , \new_[12880]_ ,
    \new_[12881]_ , \new_[12882]_ , \new_[12883]_ , \new_[12884]_ ,
    \new_[12885]_ , \new_[12886]_ , \new_[12887]_ , \new_[12888]_ ,
    \new_[12889]_ , \new_[12890]_ , \new_[12891]_ , \new_[12892]_ ,
    \new_[12893]_ , \new_[12894]_ , \new_[12895]_ , \new_[12896]_ ,
    \new_[12897]_ , \new_[12898]_ , \new_[12899]_ , \new_[12900]_ ,
    \new_[12901]_ , \new_[12902]_ , \new_[12903]_ , \new_[12904]_ ,
    \new_[12905]_ , \new_[12906]_ , \new_[12907]_ , \new_[12908]_ ,
    \new_[12909]_ , \new_[12910]_ , \new_[12911]_ , \new_[12912]_ ,
    \new_[12913]_ , \new_[12914]_ , \new_[12915]_ , \new_[12916]_ ,
    \new_[12917]_ , \new_[12918]_ , \new_[12919]_ , \new_[12920]_ ,
    \new_[12921]_ , \new_[12922]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12926]_ , \new_[12927]_ , \new_[12928]_ ,
    \new_[12929]_ , \new_[12930]_ , \new_[12931]_ , \new_[12932]_ ,
    \new_[12933]_ , \new_[12934]_ , \new_[12935]_ , \new_[12936]_ ,
    \new_[12937]_ , \new_[12938]_ , \new_[12939]_ , \new_[12940]_ ,
    \new_[12941]_ , \new_[12942]_ , \new_[12943]_ , \new_[12944]_ ,
    \new_[12945]_ , \new_[12946]_ , \new_[12947]_ , \new_[12948]_ ,
    \new_[12949]_ , \new_[12950]_ , \new_[12951]_ , \new_[12952]_ ,
    \new_[12953]_ , \new_[12954]_ , \new_[12955]_ , \new_[12956]_ ,
    \new_[12957]_ , \new_[12958]_ , \new_[12959]_ , \new_[12960]_ ,
    \new_[12961]_ , \new_[12962]_ , \new_[12963]_ , \new_[12964]_ ,
    \new_[12965]_ , \new_[12966]_ , \new_[12967]_ , \new_[12968]_ ,
    \new_[12969]_ , \new_[12970]_ , \new_[12971]_ , \new_[12972]_ ,
    \new_[12973]_ , \new_[12974]_ , \new_[12975]_ , \new_[12976]_ ,
    \new_[12977]_ , \new_[12978]_ , \new_[12979]_ , \new_[12980]_ ,
    \new_[12981]_ , \new_[12982]_ , \new_[12983]_ , \new_[12984]_ ,
    \new_[12985]_ , \new_[12986]_ , \new_[12987]_ , \new_[12988]_ ,
    \new_[12989]_ , \new_[12990]_ , \new_[12991]_ , \new_[12992]_ ,
    \new_[12993]_ , \new_[12994]_ , \new_[12995]_ , \new_[12996]_ ,
    \new_[12997]_ , \new_[12998]_ , \new_[12999]_ , \new_[13000]_ ,
    \new_[13001]_ , \new_[13002]_ , \new_[13003]_ , \new_[13004]_ ,
    \new_[13005]_ , \new_[13006]_ , \new_[13007]_ , \new_[13008]_ ,
    \new_[13009]_ , \new_[13010]_ , \new_[13011]_ , \new_[13012]_ ,
    \new_[13013]_ , \new_[13014]_ , \new_[13015]_ , \new_[13016]_ ,
    \new_[13017]_ , \new_[13018]_ , \new_[13019]_ , \new_[13020]_ ,
    \new_[13021]_ , \new_[13022]_ , \new_[13023]_ , \new_[13024]_ ,
    \new_[13025]_ , \new_[13026]_ , \new_[13027]_ , \new_[13028]_ ,
    \new_[13029]_ , \new_[13030]_ , \new_[13031]_ , \new_[13032]_ ,
    \new_[13033]_ , \new_[13034]_ , \new_[13035]_ , \new_[13036]_ ,
    \new_[13037]_ , \new_[13038]_ , \new_[13039]_ , \new_[13040]_ ,
    \new_[13041]_ , \new_[13042]_ , \new_[13043]_ , \new_[13044]_ ,
    \new_[13045]_ , \new_[13046]_ , \new_[13047]_ , \new_[13048]_ ,
    \new_[13049]_ , \new_[13050]_ , \new_[13051]_ , \new_[13052]_ ,
    \new_[13053]_ , \new_[13054]_ , \new_[13055]_ , \new_[13056]_ ,
    \new_[13057]_ , \new_[13058]_ , \new_[13059]_ , \new_[13060]_ ,
    \new_[13061]_ , \new_[13062]_ , \new_[13063]_ , \new_[13064]_ ,
    \new_[13065]_ , \new_[13066]_ , \new_[13067]_ , \new_[13068]_ ,
    \new_[13069]_ , \new_[13070]_ , \new_[13071]_ , \new_[13072]_ ,
    \new_[13073]_ , \new_[13074]_ , \new_[13075]_ , \new_[13076]_ ,
    \new_[13077]_ , \new_[13078]_ , \new_[13079]_ , \new_[13080]_ ,
    \new_[13081]_ , \new_[13082]_ , \new_[13083]_ , \new_[13084]_ ,
    \new_[13085]_ , \new_[13086]_ , \new_[13087]_ , \new_[13088]_ ,
    \new_[13089]_ , \new_[13090]_ , \new_[13091]_ , \new_[13092]_ ,
    \new_[13093]_ , \new_[13094]_ , \new_[13095]_ , \new_[13096]_ ,
    \new_[13097]_ , \new_[13098]_ , \new_[13099]_ , \new_[13100]_ ,
    \new_[13101]_ , \new_[13102]_ , \new_[13103]_ , \new_[13104]_ ,
    \new_[13105]_ , \new_[13106]_ , \new_[13107]_ , \new_[13108]_ ,
    \new_[13109]_ , \new_[13110]_ , \new_[13111]_ , \new_[13112]_ ,
    \new_[13113]_ , \new_[13114]_ , \new_[13115]_ , \new_[13116]_ ,
    \new_[13117]_ , \new_[13118]_ , \new_[13119]_ , \new_[13120]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13123]_ , \new_[13124]_ ,
    \new_[13125]_ , \new_[13126]_ , \new_[13127]_ , \new_[13128]_ ,
    \new_[13129]_ , \new_[13130]_ , \new_[13131]_ , \new_[13132]_ ,
    \new_[13133]_ , \new_[13134]_ , \new_[13135]_ , \new_[13136]_ ,
    \new_[13137]_ , \new_[13138]_ , \new_[13139]_ , \new_[13140]_ ,
    \new_[13141]_ , \new_[13142]_ , \new_[13143]_ , \new_[13144]_ ,
    \new_[13145]_ , \new_[13146]_ , \new_[13147]_ , \new_[13148]_ ,
    \new_[13149]_ , \new_[13150]_ , \new_[13151]_ , \new_[13152]_ ,
    \new_[13153]_ , \new_[13154]_ , \new_[13155]_ , \new_[13156]_ ,
    \new_[13157]_ , \new_[13158]_ , \new_[13159]_ , \new_[13160]_ ,
    \new_[13161]_ , \new_[13162]_ , \new_[13163]_ , \new_[13164]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13167]_ , \new_[13168]_ ,
    \new_[13169]_ , \new_[13170]_ , \new_[13171]_ , \new_[13172]_ ,
    \new_[13173]_ , \new_[13174]_ , \new_[13175]_ , \new_[13176]_ ,
    \new_[13177]_ , \new_[13178]_ , \new_[13179]_ , \new_[13180]_ ,
    \new_[13181]_ , \new_[13182]_ , \new_[13183]_ , \new_[13184]_ ,
    \new_[13185]_ , \new_[13186]_ , \new_[13187]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13190]_ , \new_[13191]_ , \new_[13192]_ ,
    \new_[13193]_ , \new_[13194]_ , \new_[13195]_ , \new_[13196]_ ,
    \new_[13197]_ , \new_[13198]_ , \new_[13199]_ , \new_[13200]_ ,
    \new_[13201]_ , \new_[13202]_ , \new_[13203]_ , \new_[13204]_ ,
    \new_[13205]_ , \new_[13206]_ , \new_[13207]_ , \new_[13208]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13211]_ , \new_[13212]_ ,
    \new_[13213]_ , \new_[13214]_ , \new_[13215]_ , \new_[13216]_ ,
    \new_[13217]_ , \new_[13218]_ , \new_[13219]_ , \new_[13220]_ ,
    \new_[13221]_ , \new_[13222]_ , \new_[13223]_ , \new_[13224]_ ,
    \new_[13225]_ , \new_[13226]_ , \new_[13227]_ , \new_[13228]_ ,
    \new_[13229]_ , \new_[13230]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13234]_ , \new_[13235]_ , \new_[13236]_ ,
    \new_[13237]_ , \new_[13238]_ , \new_[13239]_ , \new_[13240]_ ,
    \new_[13241]_ , \new_[13242]_ , \new_[13243]_ , \new_[13244]_ ,
    \new_[13245]_ , \new_[13246]_ , \new_[13247]_ , \new_[13248]_ ,
    \new_[13249]_ , \new_[13250]_ , \new_[13251]_ , \new_[13252]_ ,
    \new_[13253]_ , \new_[13254]_ , \new_[13255]_ , \new_[13256]_ ,
    \new_[13257]_ , \new_[13258]_ , \new_[13259]_ , \new_[13260]_ ,
    \new_[13261]_ , \new_[13262]_ , \new_[13263]_ , \new_[13264]_ ,
    \new_[13265]_ , \new_[13266]_ , \new_[13267]_ , \new_[13268]_ ,
    \new_[13269]_ , \new_[13270]_ , \new_[13271]_ , \new_[13272]_ ,
    \new_[13273]_ , \new_[13274]_ , \new_[13275]_ , \new_[13276]_ ,
    \new_[13277]_ , \new_[13278]_ , \new_[13279]_ , \new_[13280]_ ,
    \new_[13281]_ , \new_[13282]_ , \new_[13283]_ , \new_[13284]_ ,
    \new_[13285]_ , \new_[13286]_ , \new_[13287]_ , \new_[13288]_ ,
    \new_[13289]_ , \new_[13290]_ , \new_[13291]_ , \new_[13292]_ ,
    \new_[13293]_ , \new_[13294]_ , \new_[13295]_ , \new_[13296]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13300]_ ,
    \new_[13301]_ , \new_[13302]_ , \new_[13303]_ , \new_[13304]_ ,
    \new_[13305]_ , \new_[13306]_ , \new_[13307]_ , \new_[13308]_ ,
    \new_[13309]_ , \new_[13310]_ , \new_[13311]_ , \new_[13312]_ ,
    \new_[13313]_ , \new_[13314]_ , \new_[13315]_ , \new_[13316]_ ,
    \new_[13317]_ , \new_[13318]_ , \new_[13319]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13322]_ , \new_[13323]_ , \new_[13324]_ ,
    \new_[13325]_ , \new_[13326]_ , \new_[13327]_ , \new_[13328]_ ,
    \new_[13329]_ , \new_[13330]_ , \new_[13331]_ , \new_[13332]_ ,
    \new_[13333]_ , \new_[13334]_ , \new_[13335]_ , \new_[13336]_ ,
    \new_[13337]_ , \new_[13338]_ , \new_[13339]_ , \new_[13340]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13345]_ , \new_[13346]_ , \new_[13347]_ , \new_[13348]_ ,
    \new_[13349]_ , \new_[13350]_ , \new_[13351]_ , \new_[13352]_ ,
    \new_[13353]_ , \new_[13354]_ , \new_[13355]_ , \new_[13356]_ ,
    \new_[13357]_ , \new_[13358]_ , \new_[13359]_ , \new_[13360]_ ,
    \new_[13361]_ , \new_[13362]_ , \new_[13363]_ , \new_[13364]_ ,
    \new_[13365]_ , \new_[13366]_ , \new_[13367]_ , \new_[13368]_ ,
    \new_[13369]_ , \new_[13370]_ , \new_[13371]_ , \new_[13372]_ ,
    \new_[13373]_ , \new_[13374]_ , \new_[13375]_ , \new_[13376]_ ,
    \new_[13377]_ , \new_[13378]_ , \new_[13379]_ , \new_[13380]_ ,
    \new_[13381]_ , \new_[13382]_ , \new_[13383]_ , \new_[13384]_ ,
    \new_[13385]_ , \new_[13386]_ , \new_[13387]_ , \new_[13388]_ ,
    \new_[13389]_ , \new_[13390]_ , \new_[13391]_ , \new_[13392]_ ,
    \new_[13393]_ , \new_[13394]_ , \new_[13395]_ , \new_[13396]_ ,
    \new_[13397]_ , \new_[13398]_ , \new_[13399]_ , \new_[13400]_ ,
    \new_[13401]_ , \new_[13402]_ , \new_[13403]_ , \new_[13404]_ ,
    \new_[13405]_ , \new_[13406]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13410]_ , \new_[13411]_ , \new_[13412]_ ,
    \new_[13413]_ , \new_[13414]_ , \new_[13415]_ , \new_[13416]_ ,
    \new_[13417]_ , \new_[13418]_ , \new_[13419]_ , \new_[13420]_ ,
    \new_[13421]_ , \new_[13422]_ , \new_[13423]_ , \new_[13424]_ ,
    \new_[13425]_ , \new_[13426]_ , \new_[13427]_ , \new_[13428]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13432]_ ,
    \new_[13433]_ , \new_[13434]_ , \new_[13435]_ , \new_[13436]_ ,
    \new_[13437]_ , \new_[13438]_ , \new_[13439]_ , \new_[13440]_ ,
    \new_[13441]_ , \new_[13442]_ , \new_[13443]_ , \new_[13444]_ ,
    \new_[13445]_ , \new_[13446]_ , \new_[13447]_ , \new_[13448]_ ,
    \new_[13449]_ , \new_[13450]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13453]_ , \new_[13454]_ , \new_[13455]_ , \new_[13456]_ ,
    \new_[13457]_ , \new_[13458]_ , \new_[13459]_ , \new_[13460]_ ,
    \new_[13461]_ , \new_[13462]_ , \new_[13463]_ , \new_[13464]_ ,
    \new_[13465]_ , \new_[13466]_ , \new_[13467]_ , \new_[13468]_ ,
    \new_[13469]_ , \new_[13470]_ , \new_[13471]_ , \new_[13472]_ ,
    \new_[13473]_ , \new_[13474]_ , \new_[13475]_ , \new_[13476]_ ,
    \new_[13477]_ , \new_[13478]_ , \new_[13479]_ , \new_[13480]_ ,
    \new_[13481]_ , \new_[13482]_ , \new_[13483]_ , \new_[13484]_ ,
    \new_[13485]_ , \new_[13486]_ , \new_[13487]_ , \new_[13488]_ ,
    \new_[13489]_ , \new_[13490]_ , \new_[13491]_ , \new_[13492]_ ,
    \new_[13493]_ , \new_[13494]_ , \new_[13495]_ , \new_[13496]_ ,
    \new_[13497]_ , \new_[13498]_ , \new_[13499]_ , \new_[13500]_ ,
    \new_[13501]_ , \new_[13502]_ , \new_[13503]_ , \new_[13504]_ ,
    \new_[13505]_ , \new_[13506]_ , \new_[13507]_ , \new_[13508]_ ,
    \new_[13509]_ , \new_[13510]_ , \new_[13511]_ , \new_[13512]_ ,
    \new_[13513]_ , \new_[13514]_ , \new_[13515]_ , \new_[13516]_ ,
    \new_[13517]_ , \new_[13518]_ , \new_[13519]_ , \new_[13520]_ ,
    \new_[13521]_ , \new_[13522]_ , \new_[13523]_ , \new_[13524]_ ,
    \new_[13525]_ , \new_[13526]_ , \new_[13527]_ , \new_[13528]_ ,
    \new_[13529]_ , \new_[13530]_ , \new_[13531]_ , \new_[13532]_ ,
    \new_[13533]_ , \new_[13534]_ , \new_[13535]_ , \new_[13536]_ ,
    \new_[13537]_ , \new_[13538]_ , \new_[13539]_ , \new_[13540]_ ,
    \new_[13541]_ , \new_[13542]_ , \new_[13543]_ , \new_[13544]_ ,
    \new_[13545]_ , \new_[13546]_ , \new_[13547]_ , \new_[13548]_ ,
    \new_[13549]_ , \new_[13550]_ , \new_[13551]_ , \new_[13552]_ ,
    \new_[13553]_ , \new_[13554]_ , \new_[13555]_ , \new_[13556]_ ,
    \new_[13557]_ , \new_[13558]_ , \new_[13559]_ , \new_[13560]_ ,
    \new_[13561]_ , \new_[13562]_ , \new_[13563]_ , \new_[13564]_ ,
    \new_[13565]_ , \new_[13566]_ , \new_[13567]_ , \new_[13568]_ ,
    \new_[13569]_ , \new_[13570]_ , \new_[13571]_ , \new_[13572]_ ,
    \new_[13573]_ , \new_[13574]_ , \new_[13575]_ , \new_[13576]_ ,
    \new_[13577]_ , \new_[13578]_ , \new_[13579]_ , \new_[13580]_ ,
    \new_[13581]_ , \new_[13582]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13586]_ , \new_[13587]_ , \new_[13588]_ ,
    \new_[13589]_ , \new_[13590]_ , \new_[13591]_ , \new_[13592]_ ,
    \new_[13593]_ , \new_[13594]_ , \new_[13595]_ , \new_[13596]_ ,
    \new_[13597]_ , \new_[13598]_ , \new_[13599]_ , \new_[13600]_ ,
    \new_[13601]_ , \new_[13602]_ , \new_[13603]_ , \new_[13604]_ ,
    \new_[13605]_ , \new_[13606]_ , \new_[13607]_ , \new_[13608]_ ,
    \new_[13609]_ , \new_[13610]_ , \new_[13611]_ , \new_[13612]_ ,
    \new_[13613]_ , \new_[13614]_ , \new_[13615]_ , \new_[13616]_ ,
    \new_[13617]_ , \new_[13618]_ , \new_[13619]_ , \new_[13620]_ ,
    \new_[13621]_ , \new_[13622]_ , \new_[13623]_ , \new_[13624]_ ,
    \new_[13625]_ , \new_[13626]_ , \new_[13627]_ , \new_[13628]_ ,
    \new_[13629]_ , \new_[13630]_ , \new_[13631]_ , \new_[13632]_ ,
    \new_[13633]_ , \new_[13634]_ , \new_[13635]_ , \new_[13636]_ ,
    \new_[13637]_ , \new_[13638]_ , \new_[13639]_ , \new_[13640]_ ,
    \new_[13641]_ , \new_[13642]_ , \new_[13643]_ , \new_[13644]_ ,
    \new_[13645]_ , \new_[13646]_ , \new_[13647]_ , \new_[13648]_ ,
    \new_[13649]_ , \new_[13650]_ , \new_[13651]_ , \new_[13652]_ ,
    \new_[13653]_ , \new_[13654]_ , \new_[13655]_ , \new_[13656]_ ,
    \new_[13657]_ , \new_[13658]_ , \new_[13659]_ , \new_[13660]_ ,
    \new_[13661]_ , \new_[13662]_ , \new_[13663]_ , \new_[13664]_ ,
    \new_[13665]_ , \new_[13666]_ , \new_[13667]_ , \new_[13668]_ ,
    \new_[13669]_ , \new_[13670]_ , \new_[13671]_ , \new_[13672]_ ,
    \new_[13673]_ , \new_[13674]_ , \new_[13675]_ , \new_[13676]_ ,
    \new_[13677]_ , \new_[13678]_ , \new_[13679]_ , \new_[13680]_ ,
    \new_[13681]_ , \new_[13682]_ , \new_[13683]_ , \new_[13684]_ ,
    \new_[13685]_ , \new_[13686]_ , \new_[13687]_ , \new_[13688]_ ,
    \new_[13689]_ , \new_[13690]_ , \new_[13691]_ , \new_[13692]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13695]_ , \new_[13696]_ ,
    \new_[13697]_ , \new_[13698]_ , \new_[13699]_ , \new_[13700]_ ,
    \new_[13701]_ , \new_[13702]_ , \new_[13703]_ , \new_[13704]_ ,
    \new_[13705]_ , \new_[13706]_ , \new_[13707]_ , \new_[13708]_ ,
    \new_[13709]_ , \new_[13710]_ , \new_[13711]_ , \new_[13712]_ ,
    \new_[13713]_ , \new_[13714]_ , \new_[13715]_ , \new_[13716]_ ,
    \new_[13717]_ , \new_[13718]_ , \new_[13719]_ , \new_[13720]_ ,
    \new_[13721]_ , \new_[13722]_ , \new_[13723]_ , \new_[13724]_ ,
    \new_[13725]_ , \new_[13726]_ , \new_[13727]_ , \new_[13728]_ ,
    \new_[13729]_ , \new_[13730]_ , \new_[13731]_ , \new_[13732]_ ,
    \new_[13733]_ , \new_[13734]_ , \new_[13735]_ , \new_[13736]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13739]_ , \new_[13740]_ ,
    \new_[13741]_ , \new_[13742]_ , \new_[13743]_ , \new_[13744]_ ,
    \new_[13745]_ , \new_[13746]_ , \new_[13747]_ , \new_[13748]_ ,
    \new_[13749]_ , \new_[13750]_ , \new_[13751]_ , \new_[13752]_ ,
    \new_[13753]_ , \new_[13754]_ , \new_[13755]_ , \new_[13756]_ ,
    \new_[13757]_ , \new_[13758]_ , \new_[13759]_ , \new_[13760]_ ,
    \new_[13761]_ , \new_[13762]_ , \new_[13763]_ , \new_[13764]_ ,
    \new_[13765]_ , \new_[13766]_ , \new_[13767]_ , \new_[13768]_ ,
    \new_[13769]_ , \new_[13770]_ , \new_[13771]_ , \new_[13772]_ ,
    \new_[13773]_ , \new_[13774]_ , \new_[13775]_ , \new_[13776]_ ,
    \new_[13777]_ , \new_[13778]_ , \new_[13779]_ , \new_[13780]_ ,
    \new_[13781]_ , \new_[13782]_ , \new_[13783]_ , \new_[13784]_ ,
    \new_[13785]_ , \new_[13786]_ , \new_[13787]_ , \new_[13788]_ ,
    \new_[13789]_ , \new_[13790]_ , \new_[13791]_ , \new_[13792]_ ,
    \new_[13793]_ , \new_[13794]_ , \new_[13795]_ , \new_[13796]_ ,
    \new_[13797]_ , \new_[13798]_ , \new_[13799]_ , \new_[13800]_ ,
    \new_[13801]_ , \new_[13802]_ , \new_[13803]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13806]_ , \new_[13807]_ , \new_[13808]_ ,
    \new_[13809]_ , \new_[13810]_ , \new_[13811]_ , \new_[13812]_ ,
    \new_[13813]_ , \new_[13814]_ , \new_[13815]_ , \new_[13816]_ ,
    \new_[13817]_ , \new_[13818]_ , \new_[13819]_ , \new_[13820]_ ,
    \new_[13821]_ , \new_[13822]_ , \new_[13823]_ , \new_[13824]_ ,
    \new_[13825]_ , \new_[13826]_ , \new_[13827]_ , \new_[13828]_ ,
    \new_[13829]_ , \new_[13830]_ , \new_[13831]_ , \new_[13832]_ ,
    \new_[13833]_ , \new_[13834]_ , \new_[13835]_ , \new_[13836]_ ,
    \new_[13837]_ , \new_[13838]_ , \new_[13839]_ , \new_[13840]_ ,
    \new_[13841]_ , \new_[13842]_ , \new_[13843]_ , \new_[13844]_ ,
    \new_[13845]_ , \new_[13846]_ , \new_[13847]_ , \new_[13848]_ ,
    \new_[13849]_ , \new_[13850]_ , \new_[13851]_ , \new_[13852]_ ,
    \new_[13853]_ , \new_[13854]_ , \new_[13855]_ , \new_[13856]_ ,
    \new_[13857]_ , \new_[13858]_ , \new_[13859]_ , \new_[13860]_ ,
    \new_[13861]_ , \new_[13862]_ , \new_[13863]_ , \new_[13864]_ ,
    \new_[13865]_ , \new_[13866]_ , \new_[13867]_ , \new_[13868]_ ,
    \new_[13869]_ , \new_[13870]_ , \new_[13871]_ , \new_[13872]_ ,
    \new_[13873]_ , \new_[13874]_ , \new_[13875]_ , \new_[13876]_ ,
    \new_[13877]_ , \new_[13878]_ , \new_[13879]_ , \new_[13880]_ ,
    \new_[13881]_ , \new_[13882]_ , \new_[13883]_ , \new_[13884]_ ,
    \new_[13885]_ , \new_[13886]_ , \new_[13887]_ , \new_[13888]_ ,
    \new_[13889]_ , \new_[13890]_ , \new_[13891]_ , \new_[13892]_ ,
    \new_[13893]_ , \new_[13894]_ , \new_[13895]_ , \new_[13896]_ ,
    \new_[13897]_ , \new_[13898]_ , \new_[13899]_ , \new_[13900]_ ,
    \new_[13901]_ , \new_[13902]_ , \new_[13903]_ , \new_[13904]_ ,
    \new_[13905]_ , \new_[13906]_ , \new_[13907]_ , \new_[13908]_ ,
    \new_[13909]_ , \new_[13910]_ , \new_[13911]_ , \new_[13912]_ ,
    \new_[13913]_ , \new_[13914]_ , \new_[13915]_ , \new_[13916]_ ,
    \new_[13917]_ , \new_[13918]_ , \new_[13919]_ , \new_[13920]_ ,
    \new_[13921]_ , \new_[13922]_ , \new_[13923]_ , \new_[13924]_ ,
    \new_[13925]_ , \new_[13926]_ , \new_[13927]_ , \new_[13928]_ ,
    \new_[13929]_ , \new_[13930]_ , \new_[13931]_ , \new_[13932]_ ,
    \new_[13933]_ , \new_[13934]_ , \new_[13935]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13938]_ , \new_[13939]_ , \new_[13940]_ ,
    \new_[13941]_ , \new_[13942]_ , \new_[13943]_ , \new_[13944]_ ,
    \new_[13945]_ , \new_[13946]_ , \new_[13947]_ , \new_[13948]_ ,
    \new_[13949]_ , \new_[13950]_ , \new_[13951]_ , \new_[13952]_ ,
    \new_[13953]_ , \new_[13954]_ , \new_[13955]_ , \new_[13956]_ ,
    \new_[13957]_ , \new_[13958]_ , \new_[13959]_ , \new_[13960]_ ,
    \new_[13961]_ , \new_[13962]_ , \new_[13963]_ , \new_[13964]_ ,
    \new_[13965]_ , \new_[13966]_ , \new_[13967]_ , \new_[13968]_ ,
    \new_[13969]_ , \new_[13970]_ , \new_[13971]_ , \new_[13972]_ ,
    \new_[13973]_ , \new_[13974]_ , \new_[13975]_ , \new_[13976]_ ,
    \new_[13977]_ , \new_[13978]_ , \new_[13979]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13982]_ , \new_[13983]_ , \new_[13984]_ ,
    \new_[13985]_ , \new_[13986]_ , \new_[13987]_ , \new_[13988]_ ,
    \new_[13989]_ , \new_[13990]_ , \new_[13991]_ , \new_[13992]_ ,
    \new_[13993]_ , \new_[13994]_ , \new_[13995]_ , \new_[13996]_ ,
    \new_[13997]_ , \new_[13998]_ , \new_[13999]_ , \new_[14000]_ ,
    \new_[14001]_ , \new_[14002]_ , \new_[14003]_ , \new_[14004]_ ,
    \new_[14005]_ , \new_[14006]_ , \new_[14007]_ , \new_[14008]_ ,
    \new_[14009]_ , \new_[14010]_ , \new_[14011]_ , \new_[14012]_ ,
    \new_[14013]_ , \new_[14014]_ , \new_[14015]_ , \new_[14016]_ ,
    \new_[14017]_ , \new_[14018]_ , \new_[14019]_ , \new_[14020]_ ,
    \new_[14021]_ , \new_[14022]_ , \new_[14023]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14026]_ , \new_[14027]_ , \new_[14028]_ ,
    \new_[14029]_ , \new_[14030]_ , \new_[14031]_ , \new_[14032]_ ,
    \new_[14033]_ , \new_[14034]_ , \new_[14035]_ , \new_[14036]_ ,
    \new_[14037]_ , \new_[14038]_ , \new_[14039]_ , \new_[14040]_ ,
    \new_[14041]_ , \new_[14042]_ , \new_[14043]_ , \new_[14044]_ ,
    \new_[14045]_ , \new_[14046]_ , \new_[14047]_ , \new_[14048]_ ,
    \new_[14049]_ , \new_[14050]_ , \new_[14051]_ , \new_[14052]_ ,
    \new_[14053]_ , \new_[14054]_ , \new_[14055]_ , \new_[14056]_ ,
    \new_[14057]_ , \new_[14058]_ , \new_[14059]_ , \new_[14060]_ ,
    \new_[14061]_ , \new_[14062]_ , \new_[14063]_ , \new_[14064]_ ,
    \new_[14065]_ , \new_[14066]_ , \new_[14067]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14070]_ , \new_[14071]_ , \new_[14072]_ ,
    \new_[14073]_ , \new_[14074]_ , \new_[14075]_ , \new_[14076]_ ,
    \new_[14077]_ , \new_[14078]_ , \new_[14079]_ , \new_[14080]_ ,
    \new_[14081]_ , \new_[14082]_ , \new_[14083]_ , \new_[14084]_ ,
    \new_[14085]_ , \new_[14086]_ , \new_[14087]_ , \new_[14088]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14091]_ , \new_[14092]_ ,
    \new_[14093]_ , \new_[14094]_ , \new_[14095]_ , \new_[14096]_ ,
    \new_[14097]_ , \new_[14098]_ , \new_[14099]_ , \new_[14100]_ ,
    \new_[14101]_ , \new_[14102]_ , \new_[14103]_ , \new_[14104]_ ,
    \new_[14105]_ , \new_[14106]_ , \new_[14107]_ , \new_[14108]_ ,
    \new_[14109]_ , \new_[14110]_ , \new_[14111]_ , \new_[14112]_ ,
    \new_[14113]_ , \new_[14114]_ , \new_[14115]_ , \new_[14116]_ ,
    \new_[14117]_ , \new_[14118]_ , \new_[14119]_ , \new_[14120]_ ,
    \new_[14121]_ , \new_[14122]_ , \new_[14123]_ , \new_[14124]_ ,
    \new_[14125]_ , \new_[14126]_ , \new_[14127]_ , \new_[14128]_ ,
    \new_[14129]_ , \new_[14130]_ , \new_[14131]_ , \new_[14132]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14137]_ , \new_[14138]_ , \new_[14139]_ , \new_[14140]_ ,
    \new_[14141]_ , \new_[14142]_ , \new_[14143]_ , \new_[14144]_ ,
    \new_[14145]_ , \new_[14146]_ , \new_[14147]_ , \new_[14148]_ ,
    \new_[14149]_ , \new_[14150]_ , \new_[14151]_ , \new_[14152]_ ,
    \new_[14153]_ , \new_[14154]_ , \new_[14155]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14158]_ , \new_[14159]_ , \new_[14160]_ ,
    \new_[14161]_ , \new_[14162]_ , \new_[14163]_ , \new_[14164]_ ,
    \new_[14165]_ , \new_[14166]_ , \new_[14167]_ , \new_[14168]_ ,
    \new_[14169]_ , \new_[14170]_ , \new_[14171]_ , \new_[14172]_ ,
    \new_[14173]_ , \new_[14174]_ , \new_[14175]_ , \new_[14176]_ ,
    \new_[14177]_ , \new_[14178]_ , \new_[14179]_ , \new_[14180]_ ,
    \new_[14181]_ , \new_[14182]_ , \new_[14183]_ , \new_[14184]_ ,
    \new_[14185]_ , \new_[14186]_ , \new_[14187]_ , \new_[14188]_ ,
    \new_[14189]_ , \new_[14190]_ , \new_[14191]_ , \new_[14192]_ ,
    \new_[14193]_ , \new_[14194]_ , \new_[14195]_ , \new_[14196]_ ,
    \new_[14197]_ , \new_[14198]_ , \new_[14199]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14202]_ , \new_[14203]_ , \new_[14204]_ ,
    \new_[14205]_ , \new_[14206]_ , \new_[14207]_ , \new_[14208]_ ,
    \new_[14209]_ , \new_[14210]_ , \new_[14211]_ , \new_[14212]_ ,
    \new_[14213]_ , \new_[14214]_ , \new_[14215]_ , \new_[14216]_ ,
    \new_[14217]_ , \new_[14218]_ , \new_[14219]_ , \new_[14220]_ ,
    \new_[14221]_ , \new_[14222]_ , \new_[14223]_ , \new_[14224]_ ,
    \new_[14225]_ , \new_[14226]_ , \new_[14227]_ , \new_[14228]_ ,
    \new_[14229]_ , \new_[14230]_ , \new_[14231]_ , \new_[14232]_ ,
    \new_[14233]_ , \new_[14234]_ , \new_[14235]_ , \new_[14236]_ ,
    \new_[14237]_ , \new_[14238]_ , \new_[14239]_ , \new_[14240]_ ,
    \new_[14241]_ , \new_[14242]_ , \new_[14243]_ , \new_[14244]_ ,
    \new_[14245]_ , \new_[14246]_ , \new_[14247]_ , \new_[14248]_ ,
    \new_[14249]_ , \new_[14250]_ , \new_[14251]_ , \new_[14252]_ ,
    \new_[14253]_ , \new_[14254]_ , \new_[14255]_ , \new_[14256]_ ,
    \new_[14257]_ , \new_[14258]_ , \new_[14259]_ , \new_[14260]_ ,
    \new_[14261]_ , \new_[14262]_ , \new_[14263]_ , \new_[14264]_ ,
    \new_[14265]_ , \new_[14266]_ , \new_[14267]_ , \new_[14268]_ ,
    \new_[14269]_ , \new_[14270]_ , \new_[14271]_ , \new_[14272]_ ,
    \new_[14273]_ , \new_[14274]_ , \new_[14275]_ , \new_[14276]_ ,
    \new_[14277]_ , \new_[14278]_ , \new_[14279]_ , \new_[14280]_ ,
    \new_[14281]_ , \new_[14282]_ , \new_[14283]_ , \new_[14284]_ ,
    \new_[14285]_ , \new_[14286]_ , \new_[14287]_ , \new_[14288]_ ,
    \new_[14289]_ , \new_[14290]_ , \new_[14291]_ , \new_[14292]_ ,
    \new_[14293]_ , \new_[14294]_ , \new_[14295]_ , \new_[14296]_ ,
    \new_[14297]_ , \new_[14298]_ , \new_[14299]_ , \new_[14300]_ ,
    \new_[14301]_ , \new_[14302]_ , \new_[14303]_ , \new_[14304]_ ,
    \new_[14305]_ , \new_[14306]_ , \new_[14307]_ , \new_[14308]_ ,
    \new_[14309]_ , \new_[14310]_ , \new_[14311]_ , \new_[14312]_ ,
    \new_[14313]_ , \new_[14314]_ , \new_[14315]_ , \new_[14316]_ ,
    \new_[14317]_ , \new_[14318]_ , \new_[14319]_ , \new_[14320]_ ,
    \new_[14321]_ , \new_[14322]_ , \new_[14323]_ , \new_[14324]_ ,
    \new_[14325]_ , \new_[14326]_ , \new_[14327]_ , \new_[14328]_ ,
    \new_[14329]_ , \new_[14330]_ , \new_[14331]_ , \new_[14332]_ ,
    \new_[14333]_ , \new_[14334]_ , \new_[14335]_ , \new_[14336]_ ,
    \new_[14337]_ , \new_[14338]_ , \new_[14339]_ , \new_[14340]_ ,
    \new_[14341]_ , \new_[14342]_ , \new_[14343]_ , \new_[14344]_ ,
    \new_[14345]_ , \new_[14346]_ , \new_[14347]_ , \new_[14348]_ ,
    \new_[14349]_ , \new_[14350]_ , \new_[14351]_ , \new_[14352]_ ,
    \new_[14353]_ , \new_[14354]_ , \new_[14355]_ , \new_[14356]_ ,
    \new_[14357]_ , \new_[14358]_ , \new_[14359]_ , \new_[14360]_ ,
    \new_[14361]_ , \new_[14362]_ , \new_[14363]_ , \new_[14364]_ ,
    \new_[14365]_ , \new_[14366]_ , \new_[14367]_ , \new_[14368]_ ,
    \new_[14369]_ , \new_[14370]_ , \new_[14371]_ , \new_[14372]_ ,
    \new_[14373]_ , \new_[14374]_ , \new_[14375]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14378]_ , \new_[14379]_ , \new_[14380]_ ,
    \new_[14381]_ , \new_[14382]_ , \new_[14383]_ , \new_[14384]_ ,
    \new_[14385]_ , \new_[14386]_ , \new_[14387]_ , \new_[14388]_ ,
    \new_[14389]_ , \new_[14390]_ , \new_[14391]_ , \new_[14392]_ ,
    \new_[14393]_ , \new_[14394]_ , \new_[14395]_ , \new_[14396]_ ,
    \new_[14397]_ , \new_[14398]_ , \new_[14399]_ , \new_[14400]_ ,
    \new_[14401]_ , \new_[14402]_ , \new_[14403]_ , \new_[14404]_ ,
    \new_[14405]_ , \new_[14406]_ , \new_[14407]_ , \new_[14408]_ ,
    \new_[14409]_ , \new_[14410]_ , \new_[14411]_ , \new_[14412]_ ,
    \new_[14413]_ , \new_[14414]_ , \new_[14415]_ , \new_[14416]_ ,
    \new_[14417]_ , \new_[14418]_ , \new_[14419]_ , \new_[14420]_ ,
    \new_[14421]_ , \new_[14422]_ , \new_[14423]_ , \new_[14424]_ ,
    \new_[14425]_ , \new_[14426]_ , \new_[14427]_ , \new_[14428]_ ,
    \new_[14429]_ , \new_[14430]_ , \new_[14431]_ , \new_[14432]_ ,
    \new_[14433]_ , \new_[14434]_ , \new_[14435]_ , \new_[14436]_ ,
    \new_[14437]_ , \new_[14438]_ , \new_[14439]_ , \new_[14440]_ ,
    \new_[14441]_ , \new_[14442]_ , \new_[14443]_ , \new_[14444]_ ,
    \new_[14445]_ , \new_[14446]_ , \new_[14447]_ , \new_[14448]_ ,
    \new_[14449]_ , \new_[14450]_ , \new_[14451]_ , \new_[14452]_ ,
    \new_[14453]_ , \new_[14454]_ , \new_[14455]_ , \new_[14456]_ ,
    \new_[14457]_ , \new_[14458]_ , \new_[14459]_ , \new_[14460]_ ,
    \new_[14461]_ , \new_[14462]_ , \new_[14463]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14466]_ , \new_[14467]_ , \new_[14468]_ ,
    \new_[14469]_ , \new_[14470]_ , \new_[14471]_ , \new_[14472]_ ,
    \new_[14473]_ , \new_[14474]_ , \new_[14475]_ , \new_[14476]_ ,
    \new_[14477]_ , \new_[14478]_ , \new_[14479]_ , \new_[14480]_ ,
    \new_[14481]_ , \new_[14482]_ , \new_[14483]_ , \new_[14484]_ ,
    \new_[14485]_ , \new_[14486]_ , \new_[14487]_ , \new_[14488]_ ,
    \new_[14489]_ , \new_[14490]_ , \new_[14491]_ , \new_[14492]_ ,
    \new_[14493]_ , \new_[14494]_ , \new_[14495]_ , \new_[14496]_ ,
    \new_[14497]_ , \new_[14498]_ , \new_[14499]_ , \new_[14500]_ ,
    \new_[14501]_ , \new_[14502]_ , \new_[14503]_ , \new_[14504]_ ,
    \new_[14505]_ , \new_[14506]_ , \new_[14507]_ , \new_[14508]_ ,
    \new_[14509]_ , \new_[14510]_ , \new_[14511]_ , \new_[14512]_ ,
    \new_[14513]_ , \new_[14514]_ , \new_[14515]_ , \new_[14516]_ ,
    \new_[14517]_ , \new_[14518]_ , \new_[14519]_ , \new_[14520]_ ,
    \new_[14521]_ , \new_[14522]_ , \new_[14523]_ , \new_[14524]_ ,
    \new_[14525]_ , \new_[14526]_ , \new_[14527]_ , \new_[14528]_ ,
    \new_[14529]_ , \new_[14530]_ , \new_[14531]_ , \new_[14532]_ ,
    \new_[14533]_ , \new_[14534]_ , \new_[14535]_ , \new_[14536]_ ,
    \new_[14537]_ , \new_[14538]_ , \new_[14539]_ , \new_[14540]_ ,
    \new_[14541]_ , \new_[14542]_ , \new_[14543]_ , \new_[14544]_ ,
    \new_[14545]_ , \new_[14546]_ , \new_[14547]_ , \new_[14548]_ ,
    \new_[14549]_ , \new_[14550]_ , \new_[14551]_ , \new_[14552]_ ,
    \new_[14553]_ , \new_[14554]_ , \new_[14555]_ , \new_[14556]_ ,
    \new_[14557]_ , \new_[14558]_ , \new_[14559]_ , \new_[14560]_ ,
    \new_[14561]_ , \new_[14562]_ , \new_[14563]_ , \new_[14564]_ ,
    \new_[14565]_ , \new_[14566]_ , \new_[14567]_ , \new_[14568]_ ,
    \new_[14569]_ , \new_[14570]_ , \new_[14571]_ , \new_[14572]_ ,
    \new_[14573]_ , \new_[14574]_ , \new_[14575]_ , \new_[14576]_ ,
    \new_[14577]_ , \new_[14578]_ , \new_[14579]_ , \new_[14580]_ ,
    \new_[14581]_ , \new_[14582]_ , \new_[14583]_ , \new_[14584]_ ,
    \new_[14585]_ , \new_[14586]_ , \new_[14587]_ , \new_[14588]_ ,
    \new_[14589]_ , \new_[14590]_ , \new_[14591]_ , \new_[14592]_ ,
    \new_[14593]_ , \new_[14594]_ , \new_[14595]_ , \new_[14596]_ ,
    \new_[14597]_ , \new_[14598]_ , \new_[14599]_ , \new_[14600]_ ,
    \new_[14601]_ , \new_[14602]_ , \new_[14603]_ , \new_[14604]_ ,
    \new_[14605]_ , \new_[14606]_ , \new_[14607]_ , \new_[14608]_ ,
    \new_[14609]_ , \new_[14610]_ , \new_[14611]_ , \new_[14612]_ ,
    \new_[14613]_ , \new_[14614]_ , \new_[14615]_ , \new_[14616]_ ,
    \new_[14617]_ , \new_[14618]_ , \new_[14619]_ , \new_[14620]_ ,
    \new_[14621]_ , \new_[14622]_ , \new_[14623]_ , \new_[14624]_ ,
    \new_[14625]_ , \new_[14626]_ , \new_[14627]_ , \new_[14628]_ ,
    \new_[14629]_ , \new_[14630]_ , \new_[14631]_ , \new_[14632]_ ,
    \new_[14633]_ , \new_[14634]_ , \new_[14635]_ , \new_[14636]_ ,
    \new_[14637]_ , \new_[14638]_ , \new_[14639]_ , \new_[14640]_ ,
    \new_[14641]_ , \new_[14642]_ , \new_[14643]_ , \new_[14644]_ ,
    \new_[14645]_ , \new_[14646]_ , \new_[14647]_ , \new_[14648]_ ,
    \new_[14649]_ , \new_[14650]_ , \new_[14651]_ , \new_[14652]_ ,
    \new_[14653]_ , \new_[14654]_ , \new_[14655]_ , \new_[14656]_ ,
    \new_[14657]_ , \new_[14658]_ , \new_[14659]_ , \new_[14660]_ ,
    \new_[14661]_ , \new_[14662]_ , \new_[14663]_ , \new_[14664]_ ,
    \new_[14665]_ , \new_[14666]_ , \new_[14667]_ , \new_[14668]_ ,
    \new_[14669]_ , \new_[14670]_ , \new_[14671]_ , \new_[14672]_ ,
    \new_[14673]_ , \new_[14674]_ , \new_[14675]_ , \new_[14676]_ ,
    \new_[14677]_ , \new_[14678]_ , \new_[14679]_ , \new_[14680]_ ,
    \new_[14681]_ , \new_[14682]_ , \new_[14683]_ , \new_[14684]_ ,
    \new_[14685]_ , \new_[14686]_ , \new_[14687]_ , \new_[14688]_ ,
    \new_[14689]_ , \new_[14690]_ , \new_[14691]_ , \new_[14692]_ ,
    \new_[14693]_ , \new_[14694]_ , \new_[14695]_ , \new_[14696]_ ,
    \new_[14697]_ , \new_[14698]_ , \new_[14699]_ , \new_[14700]_ ,
    \new_[14701]_ , \new_[14702]_ , \new_[14703]_ , \new_[14704]_ ,
    \new_[14705]_ , \new_[14706]_ , \new_[14707]_ , \new_[14708]_ ,
    \new_[14709]_ , \new_[14710]_ , \new_[14711]_ , \new_[14712]_ ,
    \new_[14713]_ , \new_[14714]_ , \new_[14715]_ , \new_[14716]_ ,
    \new_[14717]_ , \new_[14718]_ , \new_[14719]_ , \new_[14720]_ ,
    \new_[14721]_ , \new_[14722]_ , \new_[14723]_ , \new_[14724]_ ,
    \new_[14725]_ , \new_[14726]_ , \new_[14727]_ , \new_[14728]_ ,
    \new_[14729]_ , \new_[14730]_ , \new_[14731]_ , \new_[14732]_ ,
    \new_[14733]_ , \new_[14734]_ , \new_[14735]_ , \new_[14736]_ ,
    \new_[14737]_ , \new_[14738]_ , \new_[14739]_ , \new_[14740]_ ,
    \new_[14741]_ , \new_[14742]_ , \new_[14743]_ , \new_[14744]_ ,
    \new_[14745]_ , \new_[14746]_ , \new_[14747]_ , \new_[14748]_ ,
    \new_[14749]_ , \new_[14750]_ , \new_[14751]_ , \new_[14752]_ ,
    \new_[14753]_ , \new_[14754]_ , \new_[14755]_ , \new_[14756]_ ,
    \new_[14757]_ , \new_[14758]_ , \new_[14759]_ , \new_[14760]_ ,
    \new_[14761]_ , \new_[14762]_ , \new_[14763]_ , \new_[14764]_ ,
    \new_[14765]_ , \new_[14766]_ , \new_[14767]_ , \new_[14768]_ ,
    \new_[14769]_ , \new_[14770]_ , \new_[14771]_ , \new_[14772]_ ,
    \new_[14773]_ , \new_[14774]_ , \new_[14775]_ , \new_[14776]_ ,
    \new_[14777]_ , \new_[14778]_ , \new_[14779]_ , \new_[14780]_ ,
    \new_[14781]_ , \new_[14782]_ , \new_[14783]_ , \new_[14784]_ ,
    \new_[14785]_ , \new_[14786]_ , \new_[14787]_ , \new_[14788]_ ,
    \new_[14789]_ , \new_[14790]_ , \new_[14791]_ , \new_[14792]_ ,
    \new_[14793]_ , \new_[14794]_ , \new_[14795]_ , \new_[14796]_ ,
    \new_[14797]_ , \new_[14798]_ , \new_[14799]_ , \new_[14800]_ ,
    \new_[14801]_ , \new_[14802]_ , \new_[14803]_ , \new_[14804]_ ,
    \new_[14805]_ , \new_[14806]_ , \new_[14807]_ , \new_[14808]_ ,
    \new_[14809]_ , \new_[14810]_ , \new_[14811]_ , \new_[14812]_ ,
    \new_[14813]_ , \new_[14814]_ , \new_[14815]_ , \new_[14816]_ ,
    \new_[14817]_ , \new_[14818]_ , \new_[14819]_ , \new_[14820]_ ,
    \new_[14821]_ , \new_[14822]_ , \new_[14823]_ , \new_[14824]_ ,
    \new_[14825]_ , \new_[14826]_ , \new_[14827]_ , \new_[14828]_ ,
    \new_[14829]_ , \new_[14830]_ , \new_[14831]_ , \new_[14832]_ ,
    \new_[14833]_ , \new_[14834]_ , \new_[14835]_ , \new_[14836]_ ,
    \new_[14837]_ , \new_[14838]_ , \new_[14839]_ , \new_[14840]_ ,
    \new_[14841]_ , \new_[14842]_ , \new_[14843]_ , \new_[14844]_ ,
    \new_[14845]_ , \new_[14846]_ , \new_[14847]_ , \new_[14848]_ ,
    \new_[14849]_ , \new_[14850]_ , \new_[14851]_ , \new_[14852]_ ,
    \new_[14853]_ , \new_[14854]_ , \new_[14855]_ , \new_[14856]_ ,
    \new_[14857]_ , \new_[14858]_ , \new_[14859]_ , \new_[14860]_ ,
    \new_[14861]_ , \new_[14862]_ , \new_[14863]_ , \new_[14864]_ ,
    \new_[14865]_ , \new_[14866]_ , \new_[14867]_ , \new_[14868]_ ,
    \new_[14869]_ , \new_[14870]_ , \new_[14871]_ , \new_[14872]_ ,
    \new_[14873]_ , \new_[14874]_ , \new_[14875]_ , \new_[14876]_ ,
    \new_[14877]_ , \new_[14878]_ , \new_[14879]_ , \new_[14880]_ ,
    \new_[14881]_ , \new_[14882]_ , \new_[14883]_ , \new_[14884]_ ,
    \new_[14885]_ , \new_[14886]_ , \new_[14887]_ , \new_[14888]_ ,
    \new_[14889]_ , \new_[14890]_ , \new_[14891]_ , \new_[14892]_ ,
    \new_[14893]_ , \new_[14894]_ , \new_[14895]_ , \new_[14896]_ ,
    \new_[14897]_ , \new_[14898]_ , \new_[14899]_ , \new_[14900]_ ,
    \new_[14901]_ , \new_[14902]_ , \new_[14903]_ , \new_[14904]_ ,
    \new_[14905]_ , \new_[14906]_ , \new_[14907]_ , \new_[14908]_ ,
    \new_[14909]_ , \new_[14910]_ , \new_[14911]_ , \new_[14912]_ ,
    \new_[14913]_ , \new_[14914]_ , \new_[14915]_ , \new_[14916]_ ,
    \new_[14917]_ , \new_[14918]_ , \new_[14919]_ , \new_[14920]_ ,
    \new_[14921]_ , \new_[14922]_ , \new_[14923]_ , \new_[14924]_ ,
    \new_[14925]_ , \new_[14926]_ , \new_[14927]_ , \new_[14928]_ ,
    \new_[14929]_ , \new_[14930]_ , \new_[14931]_ , \new_[14932]_ ,
    \new_[14933]_ , \new_[14934]_ , \new_[14935]_ , \new_[14936]_ ,
    \new_[14937]_ , \new_[14938]_ , \new_[14939]_ , \new_[14940]_ ,
    \new_[14941]_ , \new_[14942]_ , \new_[14943]_ , \new_[14944]_ ,
    \new_[14945]_ , \new_[14946]_ , \new_[14947]_ , \new_[14948]_ ,
    \new_[14949]_ , \new_[14950]_ , \new_[14951]_ , \new_[14952]_ ,
    \new_[14953]_ , \new_[14954]_ , \new_[14955]_ , \new_[14956]_ ,
    \new_[14957]_ , \new_[14958]_ , \new_[14959]_ , \new_[14960]_ ,
    \new_[14961]_ , \new_[14962]_ , \new_[14963]_ , \new_[14964]_ ,
    \new_[14965]_ , \new_[14966]_ , \new_[14967]_ , \new_[14968]_ ,
    \new_[14969]_ , \new_[14970]_ , \new_[14971]_ , \new_[14972]_ ,
    \new_[14973]_ , \new_[14974]_ , \new_[14975]_ , \new_[14976]_ ,
    \new_[14977]_ , \new_[14978]_ , \new_[14979]_ , \new_[14980]_ ,
    \new_[14981]_ , \new_[14982]_ , \new_[14983]_ , \new_[14984]_ ,
    \new_[14985]_ , \new_[14986]_ , \new_[14987]_ , \new_[14988]_ ,
    \new_[14989]_ , \new_[14990]_ , \new_[14991]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14994]_ , \new_[14995]_ , \new_[14996]_ ,
    \new_[14997]_ , \new_[14998]_ , \new_[14999]_ , \new_[15000]_ ,
    \new_[15001]_ , \new_[15002]_ , \new_[15003]_ , \new_[15004]_ ,
    \new_[15005]_ , \new_[15006]_ , \new_[15007]_ , \new_[15008]_ ,
    \new_[15009]_ , \new_[15010]_ , \new_[15011]_ , \new_[15012]_ ,
    \new_[15013]_ , \new_[15014]_ , \new_[15015]_ , \new_[15016]_ ,
    \new_[15017]_ , \new_[15018]_ , \new_[15019]_ , \new_[15020]_ ,
    \new_[15021]_ , \new_[15022]_ , \new_[15023]_ , \new_[15024]_ ,
    \new_[15025]_ , \new_[15026]_ , \new_[15027]_ , \new_[15028]_ ,
    \new_[15029]_ , \new_[15030]_ , \new_[15031]_ , \new_[15032]_ ,
    \new_[15033]_ , \new_[15034]_ , \new_[15035]_ , \new_[15036]_ ,
    \new_[15037]_ , \new_[15038]_ , \new_[15039]_ , \new_[15040]_ ,
    \new_[15041]_ , \new_[15042]_ , \new_[15043]_ , \new_[15044]_ ,
    \new_[15045]_ , \new_[15046]_ , \new_[15047]_ , \new_[15048]_ ,
    \new_[15049]_ , \new_[15050]_ , \new_[15051]_ , \new_[15052]_ ,
    \new_[15053]_ , \new_[15054]_ , \new_[15055]_ , \new_[15056]_ ,
    \new_[15057]_ , \new_[15058]_ , \new_[15059]_ , \new_[15060]_ ,
    \new_[15061]_ , \new_[15062]_ , \new_[15063]_ , \new_[15064]_ ,
    \new_[15065]_ , \new_[15066]_ , \new_[15067]_ , \new_[15068]_ ,
    \new_[15069]_ , \new_[15070]_ , \new_[15071]_ , \new_[15072]_ ,
    \new_[15073]_ , \new_[15074]_ , \new_[15075]_ , \new_[15076]_ ,
    \new_[15077]_ , \new_[15078]_ , \new_[15079]_ , \new_[15080]_ ,
    \new_[15081]_ , \new_[15082]_ , \new_[15083]_ , \new_[15084]_ ,
    \new_[15085]_ , \new_[15086]_ , \new_[15087]_ , \new_[15088]_ ,
    \new_[15089]_ , \new_[15090]_ , \new_[15091]_ , \new_[15092]_ ,
    \new_[15093]_ , \new_[15094]_ , \new_[15095]_ , \new_[15096]_ ,
    \new_[15097]_ , \new_[15098]_ , \new_[15099]_ , \new_[15100]_ ,
    \new_[15101]_ , \new_[15102]_ , \new_[15103]_ , \new_[15104]_ ,
    \new_[15105]_ , \new_[15106]_ , \new_[15107]_ , \new_[15108]_ ,
    \new_[15109]_ , \new_[15110]_ , \new_[15111]_ , \new_[15112]_ ,
    \new_[15113]_ , \new_[15114]_ , \new_[15115]_ , \new_[15116]_ ,
    \new_[15117]_ , \new_[15118]_ , \new_[15119]_ , \new_[15120]_ ,
    \new_[15121]_ , \new_[15122]_ , \new_[15123]_ , \new_[15124]_ ,
    \new_[15125]_ , \new_[15126]_ , \new_[15127]_ , \new_[15128]_ ,
    \new_[15129]_ , \new_[15130]_ , \new_[15131]_ , \new_[15132]_ ,
    \new_[15133]_ , \new_[15134]_ , \new_[15135]_ , \new_[15136]_ ,
    \new_[15137]_ , \new_[15138]_ , \new_[15139]_ , \new_[15140]_ ,
    \new_[15141]_ , \new_[15142]_ , \new_[15143]_ , \new_[15144]_ ,
    \new_[15145]_ , \new_[15146]_ , \new_[15147]_ , \new_[15148]_ ,
    \new_[15149]_ , \new_[15150]_ , \new_[15151]_ , \new_[15152]_ ,
    \new_[15153]_ , \new_[15154]_ , \new_[15155]_ , \new_[15156]_ ,
    \new_[15157]_ , \new_[15158]_ , \new_[15159]_ , \new_[15160]_ ,
    \new_[15161]_ , \new_[15162]_ , \new_[15163]_ , \new_[15164]_ ,
    \new_[15165]_ , \new_[15166]_ , \new_[15167]_ , \new_[15168]_ ,
    \new_[15169]_ , \new_[15170]_ , \new_[15171]_ , \new_[15172]_ ,
    \new_[15173]_ , \new_[15174]_ , \new_[15175]_ , \new_[15176]_ ,
    \new_[15177]_ , \new_[15178]_ , \new_[15179]_ , \new_[15180]_ ,
    \new_[15181]_ , \new_[15182]_ , \new_[15183]_ , \new_[15184]_ ,
    \new_[15185]_ , \new_[15186]_ , \new_[15187]_ , \new_[15188]_ ,
    \new_[15189]_ , \new_[15190]_ , \new_[15191]_ , \new_[15192]_ ,
    \new_[15193]_ , \new_[15194]_ , \new_[15195]_ , \new_[15196]_ ,
    \new_[15197]_ , \new_[15198]_ , \new_[15199]_ , \new_[15200]_ ,
    \new_[15201]_ , \new_[15202]_ , \new_[15203]_ , \new_[15204]_ ,
    \new_[15205]_ , \new_[15206]_ , \new_[15207]_ , \new_[15208]_ ,
    \new_[15209]_ , \new_[15210]_ , \new_[15211]_ , \new_[15212]_ ,
    \new_[15213]_ , \new_[15214]_ , \new_[15215]_ , \new_[15216]_ ,
    \new_[15217]_ , \new_[15218]_ , \new_[15219]_ , \new_[15220]_ ,
    \new_[15221]_ , \new_[15222]_ , \new_[15223]_ , \new_[15224]_ ,
    \new_[15225]_ , \new_[15226]_ , \new_[15227]_ , \new_[15228]_ ,
    \new_[15229]_ , \new_[15230]_ , \new_[15231]_ , \new_[15232]_ ,
    \new_[15233]_ , \new_[15234]_ , \new_[15235]_ , \new_[15236]_ ,
    \new_[15237]_ , \new_[15238]_ , \new_[15239]_ , \new_[15240]_ ,
    \new_[15241]_ , \new_[15242]_ , \new_[15243]_ , \new_[15244]_ ,
    \new_[15245]_ , \new_[15246]_ , \new_[15247]_ , \new_[15248]_ ,
    \new_[15249]_ , \new_[15250]_ , \new_[15251]_ , \new_[15252]_ ,
    \new_[15253]_ , \new_[15254]_ , \new_[15255]_ , \new_[15256]_ ,
    \new_[15257]_ , \new_[15258]_ , \new_[15259]_ , \new_[15260]_ ,
    \new_[15261]_ , \new_[15262]_ , \new_[15263]_ , \new_[15264]_ ,
    \new_[15265]_ , \new_[15266]_ , \new_[15267]_ , \new_[15268]_ ,
    \new_[15269]_ , \new_[15270]_ , \new_[15271]_ , \new_[15272]_ ,
    \new_[15273]_ , \new_[15274]_ , \new_[15275]_ , \new_[15276]_ ,
    \new_[15277]_ , \new_[15278]_ , \new_[15279]_ , \new_[15280]_ ,
    \new_[15281]_ , \new_[15282]_ , \new_[15283]_ , \new_[15284]_ ,
    \new_[15285]_ , \new_[15286]_ , \new_[15287]_ , \new_[15288]_ ,
    \new_[15289]_ , \new_[15290]_ , \new_[15291]_ , \new_[15292]_ ,
    \new_[15293]_ , \new_[15294]_ , \new_[15295]_ , \new_[15296]_ ,
    \new_[15297]_ , \new_[15298]_ , \new_[15299]_ , \new_[15300]_ ,
    \new_[15301]_ , \new_[15302]_ , \new_[15303]_ , \new_[15304]_ ,
    \new_[15305]_ , \new_[15306]_ , \new_[15307]_ , \new_[15308]_ ,
    \new_[15309]_ , \new_[15310]_ , \new_[15311]_ , \new_[15312]_ ,
    \new_[15313]_ , \new_[15314]_ , \new_[15315]_ , \new_[15316]_ ,
    \new_[15317]_ , \new_[15318]_ , \new_[15319]_ , \new_[15320]_ ,
    \new_[15321]_ , \new_[15322]_ , \new_[15323]_ , \new_[15324]_ ,
    \new_[15325]_ , \new_[15326]_ , \new_[15327]_ , \new_[15328]_ ,
    \new_[15329]_ , \new_[15330]_ , \new_[15331]_ , \new_[15332]_ ,
    \new_[15333]_ , \new_[15334]_ , \new_[15335]_ , \new_[15336]_ ,
    \new_[15337]_ , \new_[15338]_ , \new_[15339]_ , \new_[15340]_ ,
    \new_[15341]_ , \new_[15342]_ , \new_[15343]_ , \new_[15344]_ ,
    \new_[15345]_ , \new_[15346]_ , \new_[15347]_ , \new_[15348]_ ,
    \new_[15349]_ , \new_[15350]_ , \new_[15351]_ , \new_[15352]_ ,
    \new_[15353]_ , \new_[15354]_ , \new_[15355]_ , \new_[15356]_ ,
    \new_[15357]_ , \new_[15358]_ , \new_[15359]_ , \new_[15360]_ ,
    \new_[15361]_ , \new_[15362]_ , \new_[15363]_ , \new_[15364]_ ,
    \new_[15365]_ , \new_[15366]_ , \new_[15367]_ , \new_[15368]_ ,
    \new_[15369]_ , \new_[15370]_ , \new_[15371]_ , \new_[15372]_ ,
    \new_[15373]_ , \new_[15374]_ , \new_[15375]_ , \new_[15376]_ ,
    \new_[15377]_ , \new_[15378]_ , \new_[15379]_ , \new_[15380]_ ,
    \new_[15381]_ , \new_[15382]_ , \new_[15383]_ , \new_[15384]_ ,
    \new_[15385]_ , \new_[15386]_ , \new_[15387]_ , \new_[15388]_ ,
    \new_[15389]_ , \new_[15390]_ , \new_[15391]_ , \new_[15392]_ ,
    \new_[15393]_ , \new_[15394]_ , \new_[15395]_ , \new_[15396]_ ,
    \new_[15397]_ , \new_[15398]_ , \new_[15399]_ , \new_[15400]_ ,
    \new_[15401]_ , \new_[15402]_ , \new_[15403]_ , \new_[15404]_ ,
    \new_[15405]_ , \new_[15406]_ , \new_[15407]_ , \new_[15408]_ ,
    \new_[15409]_ , \new_[15410]_ , \new_[15411]_ , \new_[15412]_ ,
    \new_[15413]_ , \new_[15414]_ , \new_[15415]_ , \new_[15416]_ ,
    \new_[15417]_ , \new_[15418]_ , \new_[15419]_ , \new_[15420]_ ,
    \new_[15421]_ , \new_[15422]_ , \new_[15423]_ , \new_[15424]_ ,
    \new_[15425]_ , \new_[15426]_ , \new_[15427]_ , \new_[15428]_ ,
    \new_[15429]_ , \new_[15430]_ , \new_[15431]_ , \new_[15432]_ ,
    \new_[15433]_ , \new_[15434]_ , \new_[15435]_ , \new_[15436]_ ,
    \new_[15437]_ , \new_[15438]_ , \new_[15439]_ , \new_[15440]_ ,
    \new_[15441]_ , \new_[15442]_ , \new_[15443]_ , \new_[15444]_ ,
    \new_[15445]_ , \new_[15446]_ , \new_[15447]_ , \new_[15448]_ ,
    \new_[15449]_ , \new_[15450]_ , \new_[15451]_ , \new_[15452]_ ,
    \new_[15453]_ , \new_[15454]_ , \new_[15455]_ , \new_[15456]_ ,
    \new_[15457]_ , \new_[15458]_ , \new_[15459]_ , \new_[15460]_ ,
    \new_[15461]_ , \new_[15462]_ , \new_[15463]_ , \new_[15464]_ ,
    \new_[15465]_ , \new_[15466]_ , \new_[15467]_ , \new_[15468]_ ,
    \new_[15469]_ , \new_[15470]_ , \new_[15471]_ , \new_[15472]_ ,
    \new_[15473]_ , \new_[15474]_ , \new_[15475]_ , \new_[15476]_ ,
    \new_[15477]_ , \new_[15478]_ , \new_[15479]_ , \new_[15480]_ ,
    \new_[15481]_ , \new_[15482]_ , \new_[15483]_ , \new_[15484]_ ,
    \new_[15485]_ , \new_[15486]_ , \new_[15487]_ , \new_[15488]_ ,
    \new_[15489]_ , \new_[15490]_ , \new_[15491]_ , \new_[15492]_ ,
    \new_[15493]_ , \new_[15494]_ , \new_[15495]_ , \new_[15496]_ ,
    \new_[15497]_ , \new_[15498]_ , \new_[15499]_ , \new_[15500]_ ,
    \new_[15501]_ , \new_[15502]_ , \new_[15503]_ , \new_[15504]_ ,
    \new_[15505]_ , \new_[15506]_ , \new_[15507]_ , \new_[15508]_ ,
    \new_[15509]_ , \new_[15510]_ , \new_[15511]_ , \new_[15512]_ ,
    \new_[15513]_ , \new_[15514]_ , \new_[15515]_ , \new_[15516]_ ,
    \new_[15517]_ , \new_[15518]_ , \new_[15519]_ , \new_[15520]_ ,
    \new_[15521]_ , \new_[15522]_ , \new_[15523]_ , \new_[15524]_ ,
    \new_[15525]_ , \new_[15526]_ , \new_[15527]_ , \new_[15528]_ ,
    \new_[15529]_ , \new_[15530]_ , \new_[15531]_ , \new_[15532]_ ,
    \new_[15533]_ , \new_[15534]_ , \new_[15535]_ , \new_[15536]_ ,
    \new_[15537]_ , \new_[15538]_ , \new_[15539]_ , \new_[15540]_ ,
    \new_[15541]_ , \new_[15542]_ , \new_[15543]_ , \new_[15544]_ ,
    \new_[15545]_ , \new_[15546]_ , \new_[15547]_ , \new_[15548]_ ,
    \new_[15549]_ , \new_[15550]_ , \new_[15551]_ , \new_[15552]_ ,
    \new_[15553]_ , \new_[15554]_ , \new_[15555]_ , \new_[15556]_ ,
    \new_[15557]_ , \new_[15558]_ , \new_[15559]_ , \new_[15560]_ ,
    \new_[15561]_ , \new_[15562]_ , \new_[15563]_ , \new_[15564]_ ,
    \new_[15565]_ , \new_[15566]_ , \new_[15567]_ , \new_[15568]_ ,
    \new_[15569]_ , \new_[15570]_ , \new_[15571]_ , \new_[15572]_ ,
    \new_[15573]_ , \new_[15574]_ , \new_[15575]_ , \new_[15576]_ ,
    \new_[15577]_ , \new_[15578]_ , \new_[15579]_ , \new_[15580]_ ,
    \new_[15581]_ , \new_[15582]_ , \new_[15583]_ , \new_[15584]_ ,
    \new_[15585]_ , \new_[15586]_ , \new_[15587]_ , \new_[15588]_ ,
    \new_[15589]_ , \new_[15590]_ , \new_[15591]_ , \new_[15592]_ ,
    \new_[15593]_ , \new_[15594]_ , \new_[15595]_ , \new_[15596]_ ,
    \new_[15597]_ , \new_[15598]_ , \new_[15599]_ , \new_[15600]_ ,
    \new_[15601]_ , \new_[15602]_ , \new_[15603]_ , \new_[15604]_ ,
    \new_[15605]_ , \new_[15606]_ , \new_[15607]_ , \new_[15608]_ ,
    \new_[15609]_ , \new_[15610]_ , \new_[15611]_ , \new_[15612]_ ,
    \new_[15613]_ , \new_[15614]_ , \new_[15615]_ , \new_[15616]_ ,
    \new_[15617]_ , \new_[15618]_ , \new_[15619]_ , \new_[15620]_ ,
    \new_[15621]_ , \new_[15622]_ , \new_[15623]_ , \new_[15624]_ ,
    \new_[15625]_ , \new_[15626]_ , \new_[15627]_ , \new_[15628]_ ,
    \new_[15629]_ , \new_[15630]_ , \new_[15631]_ , \new_[15632]_ ,
    \new_[15633]_ , \new_[15634]_ , \new_[15635]_ , \new_[15636]_ ,
    \new_[15637]_ , \new_[15638]_ , \new_[15639]_ , \new_[15640]_ ,
    \new_[15641]_ , \new_[15642]_ , \new_[15643]_ , \new_[15644]_ ,
    \new_[15645]_ , \new_[15646]_ , \new_[15647]_ , \new_[15648]_ ,
    \new_[15649]_ , \new_[15650]_ , \new_[15651]_ , \new_[15652]_ ,
    \new_[15653]_ , \new_[15654]_ , \new_[15655]_ , \new_[15656]_ ,
    \new_[15657]_ , \new_[15658]_ , \new_[15659]_ , \new_[15660]_ ,
    \new_[15661]_ , \new_[15662]_ , \new_[15663]_ , \new_[15664]_ ,
    \new_[15665]_ , \new_[15666]_ , \new_[15667]_ , \new_[15668]_ ,
    \new_[15669]_ , \new_[15670]_ , \new_[15671]_ , \new_[15672]_ ,
    \new_[15673]_ , \new_[15674]_ , \new_[15675]_ , \new_[15676]_ ,
    \new_[15677]_ , \new_[15678]_ , \new_[15679]_ , \new_[15680]_ ,
    \new_[15681]_ , \new_[15682]_ , \new_[15683]_ , \new_[15684]_ ,
    \new_[15685]_ , \new_[15686]_ , \new_[15687]_ , \new_[15688]_ ,
    \new_[15689]_ , \new_[15690]_ , \new_[15691]_ , \new_[15692]_ ,
    \new_[15693]_ , \new_[15694]_ , \new_[15695]_ , \new_[15696]_ ,
    \new_[15697]_ , \new_[15698]_ , \new_[15699]_ , \new_[15700]_ ,
    \new_[15701]_ , \new_[15702]_ , \new_[15703]_ , \new_[15704]_ ,
    \new_[15705]_ , \new_[15706]_ , \new_[15707]_ , \new_[15708]_ ,
    \new_[15709]_ , \new_[15710]_ , \new_[15711]_ , \new_[15712]_ ,
    \new_[15713]_ , \new_[15714]_ , \new_[15715]_ , \new_[15716]_ ,
    \new_[15717]_ , \new_[15718]_ , \new_[15719]_ , \new_[15720]_ ,
    \new_[15721]_ , \new_[15722]_ , \new_[15723]_ , \new_[15724]_ ,
    \new_[15725]_ , \new_[15726]_ , \new_[15727]_ , \new_[15728]_ ,
    \new_[15729]_ , \new_[15730]_ , \new_[15731]_ , \new_[15732]_ ,
    \new_[15733]_ , \new_[15734]_ , \new_[15735]_ , \new_[15736]_ ,
    \new_[15737]_ , \new_[15738]_ , \new_[15739]_ , \new_[15740]_ ,
    \new_[15741]_ , \new_[15742]_ , \new_[15743]_ , \new_[15744]_ ,
    \new_[15745]_ , \new_[15746]_ , \new_[15747]_ , \new_[15748]_ ,
    \new_[15749]_ , \new_[15750]_ , \new_[15751]_ , \new_[15752]_ ,
    \new_[15753]_ , \new_[15754]_ , \new_[15755]_ , \new_[15756]_ ,
    \new_[15757]_ , \new_[15758]_ , \new_[15759]_ , \new_[15760]_ ,
    \new_[15761]_ , \new_[15762]_ , \new_[15763]_ , \new_[15764]_ ,
    \new_[15765]_ , \new_[15766]_ , \new_[15767]_ , \new_[15768]_ ,
    \new_[15769]_ , \new_[15770]_ , \new_[15771]_ , \new_[15772]_ ,
    \new_[15773]_ , \new_[15774]_ , \new_[15775]_ , \new_[15776]_ ,
    \new_[15777]_ , \new_[15778]_ , \new_[15779]_ , \new_[15780]_ ,
    \new_[15781]_ , \new_[15782]_ , \new_[15783]_ , \new_[15784]_ ,
    \new_[15785]_ , \new_[15786]_ , \new_[15787]_ , \new_[15788]_ ,
    \new_[15789]_ , \new_[15790]_ , \new_[15791]_ , \new_[15792]_ ,
    \new_[15793]_ , \new_[15794]_ , \new_[15795]_ , \new_[15796]_ ,
    \new_[15797]_ , \new_[15798]_ , \new_[15799]_ , \new_[15800]_ ,
    \new_[15801]_ , \new_[15802]_ , \new_[15803]_ , \new_[15804]_ ,
    \new_[15805]_ , \new_[15806]_ , \new_[15807]_ , \new_[15808]_ ,
    \new_[15809]_ , \new_[15810]_ , \new_[15811]_ , \new_[15812]_ ,
    \new_[15813]_ , \new_[15814]_ , \new_[15815]_ , \new_[15816]_ ,
    \new_[15817]_ , \new_[15818]_ , \new_[15819]_ , \new_[15820]_ ,
    \new_[15821]_ , \new_[15822]_ , \new_[15823]_ , \new_[15824]_ ,
    \new_[15825]_ , \new_[15826]_ , \new_[15827]_ , \new_[15828]_ ,
    \new_[15829]_ , \new_[15830]_ , \new_[15831]_ , \new_[15832]_ ,
    \new_[15833]_ , \new_[15834]_ , \new_[15835]_ , \new_[15836]_ ,
    \new_[15837]_ , \new_[15838]_ , \new_[15839]_ , \new_[15840]_ ,
    \new_[15841]_ , \new_[15842]_ , \new_[15843]_ , \new_[15844]_ ,
    \new_[15845]_ , \new_[15846]_ , \new_[15847]_ , \new_[15848]_ ,
    \new_[15849]_ , \new_[15850]_ , \new_[15851]_ , \new_[15852]_ ,
    \new_[15853]_ , \new_[15854]_ , \new_[15855]_ , \new_[15856]_ ,
    \new_[15857]_ , \new_[15858]_ , \new_[15859]_ , \new_[15860]_ ,
    \new_[15861]_ , \new_[15862]_ , \new_[15863]_ , \new_[15864]_ ,
    \new_[15865]_ , \new_[15866]_ , \new_[15867]_ , \new_[15868]_ ,
    \new_[15869]_ , \new_[15870]_ , \new_[15871]_ , \new_[15872]_ ,
    \new_[15873]_ , \new_[15874]_ , \new_[15875]_ , \new_[15876]_ ,
    \new_[15877]_ , \new_[15878]_ , \new_[15879]_ , \new_[15880]_ ,
    \new_[15881]_ , \new_[15882]_ , \new_[15883]_ , \new_[15884]_ ,
    \new_[15885]_ , \new_[15886]_ , \new_[15887]_ , \new_[15888]_ ,
    \new_[15889]_ , \new_[15890]_ , \new_[15891]_ , \new_[15892]_ ,
    \new_[15893]_ , \new_[15894]_ , \new_[15895]_ , \new_[15896]_ ,
    \new_[15897]_ , \new_[15898]_ , \new_[15899]_ , \new_[15900]_ ,
    \new_[15901]_ , \new_[15902]_ , \new_[15903]_ , \new_[15904]_ ,
    \new_[15905]_ , \new_[15906]_ , \new_[15907]_ , \new_[15908]_ ,
    \new_[15909]_ , \new_[15910]_ , \new_[15911]_ , \new_[15912]_ ,
    \new_[15913]_ , \new_[15914]_ , \new_[15915]_ , \new_[15916]_ ,
    \new_[15917]_ , \new_[15918]_ , \new_[15919]_ , \new_[15920]_ ,
    \new_[15921]_ , \new_[15922]_ , \new_[15923]_ , \new_[15924]_ ,
    \new_[15925]_ , \new_[15926]_ , \new_[15927]_ , \new_[15928]_ ,
    \new_[15929]_ , \new_[15930]_ , \new_[15931]_ , \new_[15932]_ ,
    \new_[15933]_ , \new_[15934]_ , \new_[15935]_ , \new_[15936]_ ,
    \new_[15937]_ , \new_[15938]_ , \new_[15939]_ , \new_[15940]_ ,
    \new_[15941]_ , \new_[15942]_ , \new_[15943]_ , \new_[15944]_ ,
    \new_[15945]_ , \new_[15946]_ , \new_[15947]_ , \new_[15948]_ ,
    \new_[15949]_ , \new_[15950]_ , \new_[15951]_ , \new_[15952]_ ,
    \new_[15953]_ , \new_[15954]_ , \new_[15955]_ , \new_[15956]_ ,
    \new_[15957]_ , \new_[15958]_ , \new_[15959]_ , \new_[15960]_ ,
    \new_[15961]_ , \new_[15962]_ , \new_[15963]_ , \new_[15964]_ ,
    \new_[15965]_ , \new_[15966]_ , \new_[15967]_ , \new_[15968]_ ,
    \new_[15969]_ , \new_[15970]_ , \new_[15971]_ , \new_[15972]_ ,
    \new_[15973]_ , \new_[15974]_ , \new_[15975]_ , \new_[15976]_ ,
    \new_[15977]_ , \new_[15978]_ , \new_[15979]_ , \new_[15980]_ ,
    \new_[15981]_ , \new_[15982]_ , \new_[15983]_ , \new_[15984]_ ,
    \new_[15985]_ , \new_[15986]_ , \new_[15987]_ , \new_[15988]_ ,
    \new_[15989]_ , \new_[15990]_ , \new_[15991]_ , \new_[15992]_ ,
    \new_[15993]_ , \new_[15994]_ , \new_[15995]_ , \new_[15996]_ ,
    \new_[15997]_ , \new_[15998]_ , \new_[15999]_ , \new_[16000]_ ,
    \new_[16001]_ , \new_[16002]_ , \new_[16003]_ , \new_[16004]_ ,
    \new_[16005]_ , \new_[16006]_ , \new_[16007]_ , \new_[16008]_ ,
    \new_[16009]_ , \new_[16010]_ , \new_[16011]_ , \new_[16012]_ ,
    \new_[16013]_ , \new_[16014]_ , \new_[16015]_ , \new_[16016]_ ,
    \new_[16017]_ , \new_[16018]_ , \new_[16019]_ , \new_[16020]_ ,
    \new_[16021]_ , \new_[16022]_ , \new_[16023]_ , \new_[16024]_ ,
    \new_[16025]_ , \new_[16026]_ , \new_[16027]_ , \new_[16028]_ ,
    \new_[16029]_ , \new_[16030]_ , \new_[16031]_ , \new_[16032]_ ,
    \new_[16033]_ , \new_[16034]_ , \new_[16035]_ , \new_[16036]_ ,
    \new_[16037]_ , \new_[16038]_ , \new_[16039]_ , \new_[16040]_ ,
    \new_[16041]_ , \new_[16042]_ , \new_[16043]_ , \new_[16044]_ ,
    \new_[16045]_ , \new_[16046]_ , \new_[16047]_ , \new_[16048]_ ,
    \new_[16049]_ , \new_[16050]_ , \new_[16051]_ , \new_[16052]_ ,
    \new_[16053]_ , \new_[16054]_ , \new_[16055]_ , \new_[16056]_ ,
    \new_[16057]_ , \new_[16058]_ , \new_[16059]_ , \new_[16060]_ ,
    \new_[16061]_ , \new_[16062]_ , \new_[16063]_ , \new_[16064]_ ,
    \new_[16065]_ , \new_[16066]_ , \new_[16067]_ , \new_[16068]_ ,
    \new_[16069]_ , \new_[16070]_ , \new_[16071]_ , \new_[16072]_ ,
    \new_[16073]_ , \new_[16074]_ , \new_[16075]_ , \new_[16076]_ ,
    \new_[16077]_ , \new_[16078]_ , \new_[16079]_ , \new_[16080]_ ,
    \new_[16081]_ , \new_[16082]_ , \new_[16083]_ , \new_[16084]_ ,
    \new_[16085]_ , \new_[16086]_ , \new_[16087]_ , \new_[16088]_ ,
    \new_[16089]_ , \new_[16090]_ , \new_[16091]_ , \new_[16092]_ ,
    \new_[16093]_ , \new_[16094]_ , \new_[16095]_ , \new_[16096]_ ,
    \new_[16097]_ , \new_[16098]_ , \new_[16099]_ , \new_[16100]_ ,
    \new_[16101]_ , \new_[16102]_ , \new_[16103]_ , \new_[16104]_ ,
    \new_[16105]_ , \new_[16106]_ , \new_[16107]_ , \new_[16108]_ ,
    \new_[16109]_ , \new_[16110]_ , \new_[16111]_ , \new_[16112]_ ,
    \new_[16113]_ , \new_[16114]_ , \new_[16115]_ , \new_[16116]_ ,
    \new_[16117]_ , \new_[16118]_ , \new_[16119]_ , \new_[16120]_ ,
    \new_[16121]_ , \new_[16122]_ , \new_[16123]_ , \new_[16124]_ ,
    \new_[16125]_ , \new_[16126]_ , \new_[16127]_ , \new_[16128]_ ,
    \new_[16129]_ , \new_[16130]_ , \new_[16131]_ , \new_[16132]_ ,
    \new_[16133]_ , \new_[16134]_ , \new_[16135]_ , \new_[16136]_ ,
    \new_[16137]_ , \new_[16138]_ , \new_[16139]_ , \new_[16140]_ ,
    \new_[16141]_ , \new_[16142]_ , \new_[16143]_ , \new_[16144]_ ,
    \new_[16145]_ , \new_[16146]_ , \new_[16147]_ , \new_[16148]_ ,
    \new_[16149]_ , \new_[16150]_ , \new_[16151]_ , \new_[16152]_ ,
    \new_[16153]_ , \new_[16154]_ , \new_[16155]_ , \new_[16156]_ ,
    \new_[16157]_ , \new_[16158]_ , \new_[16159]_ , \new_[16160]_ ,
    \new_[16161]_ , \new_[16162]_ , \new_[16163]_ , \new_[16164]_ ,
    \new_[16165]_ , \new_[16166]_ , \new_[16167]_ , \new_[16168]_ ,
    \new_[16169]_ , \new_[16170]_ , \new_[16171]_ , \new_[16172]_ ,
    \new_[16173]_ , \new_[16174]_ , \new_[16175]_ , \new_[16176]_ ,
    \new_[16177]_ , \new_[16178]_ , \new_[16179]_ , \new_[16180]_ ,
    \new_[16181]_ , \new_[16182]_ , \new_[16183]_ , \new_[16184]_ ,
    \new_[16185]_ , \new_[16186]_ , \new_[16187]_ , \new_[16188]_ ,
    \new_[16189]_ , \new_[16190]_ , \new_[16191]_ , \new_[16192]_ ,
    \new_[16193]_ , \new_[16194]_ , \new_[16195]_ , \new_[16196]_ ,
    \new_[16197]_ , \new_[16198]_ , \new_[16199]_ , \new_[16200]_ ,
    \new_[16201]_ , \new_[16202]_ , \new_[16203]_ , \new_[16204]_ ,
    \new_[16205]_ , \new_[16206]_ , \new_[16207]_ , \new_[16208]_ ,
    \new_[16209]_ , \new_[16210]_ , \new_[16211]_ , \new_[16212]_ ,
    \new_[16213]_ , \new_[16214]_ , \new_[16215]_ , \new_[16216]_ ,
    \new_[16217]_ , \new_[16218]_ , \new_[16219]_ , \new_[16220]_ ,
    \new_[16221]_ , \new_[16222]_ , \new_[16223]_ , \new_[16224]_ ,
    \new_[16225]_ , \new_[16226]_ , \new_[16227]_ , \new_[16228]_ ,
    \new_[16229]_ , \new_[16230]_ , \new_[16231]_ , \new_[16232]_ ,
    \new_[16233]_ , \new_[16234]_ , \new_[16235]_ , \new_[16236]_ ,
    \new_[16237]_ , \new_[16238]_ , \new_[16239]_ , \new_[16240]_ ,
    \new_[16241]_ , \new_[16242]_ , \new_[16243]_ , \new_[16244]_ ,
    \new_[16245]_ , \new_[16246]_ , \new_[16247]_ , \new_[16248]_ ,
    \new_[16249]_ , \new_[16250]_ , \new_[16251]_ , \new_[16252]_ ,
    \new_[16253]_ , \new_[16254]_ , \new_[16255]_ , \new_[16256]_ ,
    \new_[16257]_ , \new_[16258]_ , \new_[16259]_ , \new_[16260]_ ,
    \new_[16261]_ , \new_[16262]_ , \new_[16263]_ , \new_[16264]_ ,
    \new_[16265]_ , \new_[16266]_ , \new_[16267]_ , \new_[16268]_ ,
    \new_[16269]_ , \new_[16270]_ , \new_[16271]_ , \new_[16272]_ ,
    \new_[16273]_ , \new_[16274]_ , \new_[16275]_ , \new_[16276]_ ,
    \new_[16277]_ , \new_[16278]_ , \new_[16279]_ , \new_[16280]_ ,
    \new_[16281]_ , \new_[16282]_ , \new_[16283]_ , \new_[16284]_ ,
    \new_[16285]_ , \new_[16286]_ , \new_[16287]_ , \new_[16288]_ ,
    \new_[16289]_ , \new_[16290]_ , \new_[16291]_ , \new_[16292]_ ,
    \new_[16293]_ , \new_[16294]_ , \new_[16295]_ , \new_[16296]_ ,
    \new_[16297]_ , \new_[16298]_ , \new_[16299]_ , \new_[16300]_ ,
    \new_[16301]_ , \new_[16302]_ , \new_[16303]_ , \new_[16304]_ ,
    \new_[16305]_ , \new_[16306]_ , \new_[16307]_ , \new_[16308]_ ,
    \new_[16309]_ , \new_[16310]_ , \new_[16311]_ , \new_[16312]_ ,
    \new_[16313]_ , \new_[16314]_ , \new_[16315]_ , \new_[16316]_ ,
    \new_[16317]_ , \new_[16318]_ , \new_[16319]_ , \new_[16320]_ ,
    \new_[16321]_ , \new_[16322]_ , \new_[16323]_ , \new_[16324]_ ,
    \new_[16325]_ , \new_[16326]_ , \new_[16327]_ , \new_[16328]_ ,
    \new_[16329]_ , \new_[16330]_ , \new_[16331]_ , \new_[16332]_ ,
    \new_[16333]_ , \new_[16334]_ , \new_[16335]_ , \new_[16336]_ ,
    \new_[16337]_ , \new_[16338]_ , \new_[16339]_ , \new_[16340]_ ,
    \new_[16341]_ , \new_[16343]_ , \new_[16344]_ , \new_[16345]_ ,
    \new_[16346]_ , \new_[16347]_ , \new_[16348]_ , \new_[16349]_ ,
    \new_[16350]_ , \new_[16351]_ , \new_[16352]_ , \new_[16353]_ ,
    \new_[16354]_ , \new_[16355]_ , \new_[16356]_ , \new_[16357]_ ,
    \new_[16358]_ , \new_[16359]_ , \new_[16360]_ , \new_[16361]_ ,
    \new_[16362]_ , \new_[16363]_ , \new_[16364]_ , \new_[16365]_ ,
    \new_[16366]_ , \new_[16367]_ , \new_[16368]_ , \new_[16369]_ ,
    \new_[16370]_ , \new_[16371]_ , \new_[16372]_ , \new_[16373]_ ,
    \new_[16374]_ , \new_[16375]_ , \new_[16376]_ , \new_[16377]_ ,
    \new_[16378]_ , \new_[16379]_ , \new_[16380]_ , \new_[16381]_ ,
    \new_[16382]_ , \new_[16383]_ , \new_[16384]_ , \new_[16385]_ ,
    \new_[16386]_ , \new_[16387]_ , \new_[16388]_ , \new_[16389]_ ,
    \new_[16390]_ , \new_[16391]_ , \new_[16392]_ , \new_[16393]_ ,
    \new_[16394]_ , \new_[16395]_ , \new_[16396]_ , \new_[16397]_ ,
    \new_[16398]_ , \new_[16399]_ , \new_[16400]_ , \new_[16401]_ ,
    \new_[16402]_ , \new_[16403]_ , \new_[16404]_ , \new_[16405]_ ,
    \new_[16406]_ , \new_[16407]_ , \new_[16408]_ , \new_[16409]_ ,
    \new_[16410]_ , \new_[16411]_ , \new_[16412]_ , \new_[16413]_ ,
    \new_[16414]_ , \new_[16415]_ , \new_[16416]_ , \new_[16417]_ ,
    \new_[16418]_ , \new_[16419]_ , \new_[16420]_ , \new_[16421]_ ,
    \new_[16422]_ , \new_[16423]_ , \new_[16424]_ , \new_[16425]_ ,
    \new_[16426]_ , \new_[16427]_ , \new_[16428]_ , \new_[16429]_ ,
    \new_[16430]_ , \new_[16431]_ , \new_[16432]_ , \new_[16433]_ ,
    \new_[16434]_ , \new_[16435]_ , \new_[16436]_ , \new_[16437]_ ,
    \new_[16438]_ , \new_[16439]_ , \new_[16440]_ , \new_[16441]_ ,
    \new_[16442]_ , \new_[16443]_ , \new_[16444]_ , \new_[16445]_ ,
    \new_[16446]_ , \new_[16447]_ , \new_[16448]_ , \new_[16449]_ ,
    \new_[16450]_ , \new_[16451]_ , \new_[16452]_ , \new_[16453]_ ,
    \new_[16454]_ , \new_[16455]_ , \new_[16456]_ , \new_[16457]_ ,
    \new_[16458]_ , \new_[16459]_ , \new_[16460]_ , \new_[16461]_ ,
    \new_[16462]_ , \new_[16463]_ , \new_[16464]_ , \new_[16465]_ ,
    \new_[16466]_ , \new_[16467]_ , \new_[16468]_ , \new_[16469]_ ,
    \new_[16470]_ , \new_[16471]_ , \new_[16472]_ , \new_[16473]_ ,
    \new_[16474]_ , \new_[16475]_ , \new_[16476]_ , \new_[16477]_ ,
    \new_[16478]_ , \new_[16479]_ , \new_[16480]_ , \new_[16481]_ ,
    \new_[16482]_ , \new_[16483]_ , \new_[16484]_ , \new_[16485]_ ,
    \new_[16486]_ , \new_[16487]_ , \new_[16488]_ , \new_[16489]_ ,
    \new_[16490]_ , \new_[16491]_ , \new_[16492]_ , \new_[16493]_ ,
    \new_[16494]_ , \new_[16495]_ , \new_[16496]_ , \new_[16497]_ ,
    \new_[16498]_ , \new_[16499]_ , \new_[16500]_ , \new_[16501]_ ,
    \new_[16502]_ , \new_[16503]_ , \new_[16504]_ , \new_[16505]_ ,
    \new_[16506]_ , \new_[16507]_ , \new_[16508]_ , \new_[16509]_ ,
    \new_[16510]_ , \new_[16511]_ , \new_[16512]_ , \new_[16513]_ ,
    \new_[16514]_ , \new_[16515]_ , \new_[16516]_ , \new_[16517]_ ,
    \new_[16518]_ , \new_[16519]_ , \new_[16520]_ , \new_[16521]_ ,
    \new_[16522]_ , \new_[16523]_ , \new_[16524]_ , \new_[16525]_ ,
    \new_[16526]_ , \new_[16527]_ , \new_[16528]_ , \new_[16529]_ ,
    \new_[16530]_ , \new_[16531]_ , \new_[16532]_ , \new_[16533]_ ,
    \new_[16534]_ , \new_[16535]_ , \new_[16536]_ , \new_[16537]_ ,
    \new_[16538]_ , \new_[16539]_ , \new_[16540]_ , \new_[16541]_ ,
    \new_[16542]_ , \new_[16543]_ , \new_[16544]_ , \new_[16545]_ ,
    \new_[16546]_ , \new_[16547]_ , \new_[16548]_ , \new_[16549]_ ,
    \new_[16550]_ , \new_[16551]_ , \new_[16552]_ , \new_[16553]_ ,
    \new_[16554]_ , \new_[16555]_ , \new_[16556]_ , \new_[16557]_ ,
    \new_[16558]_ , \new_[16559]_ , \new_[16560]_ , \new_[16561]_ ,
    \new_[16562]_ , \new_[16563]_ , \new_[16564]_ , \new_[16565]_ ,
    \new_[16566]_ , \new_[16567]_ , \new_[16568]_ , \new_[16569]_ ,
    \new_[16570]_ , \new_[16571]_ , \new_[16572]_ , \new_[16573]_ ,
    \new_[16574]_ , \new_[16575]_ , \new_[16576]_ , \new_[16577]_ ,
    \new_[16578]_ , \new_[16579]_ , \new_[16580]_ , \new_[16581]_ ,
    \new_[16582]_ , \new_[16583]_ , \new_[16584]_ , \new_[16585]_ ,
    \new_[16586]_ , \new_[16587]_ , \new_[16588]_ , \new_[16589]_ ,
    \new_[16590]_ , \new_[16591]_ , \new_[16592]_ , \new_[16593]_ ,
    \new_[16594]_ , \new_[16595]_ , \new_[16596]_ , \new_[16597]_ ,
    \new_[16598]_ , \new_[16599]_ , \new_[16600]_ , \new_[16601]_ ,
    \new_[16602]_ , \new_[16603]_ , \new_[16604]_ , \new_[16605]_ ,
    \new_[16606]_ , \new_[16607]_ , \new_[16608]_ , \new_[16609]_ ,
    \new_[16610]_ , \new_[16611]_ , \new_[16612]_ , \new_[16613]_ ,
    \new_[16614]_ , \new_[16615]_ , \new_[16616]_ , \new_[16617]_ ,
    \new_[16618]_ , \new_[16619]_ , \new_[16620]_ , \new_[16621]_ ,
    \new_[16622]_ , \new_[16623]_ , \new_[16624]_ , \new_[16625]_ ,
    \new_[16626]_ , \new_[16627]_ , \new_[16628]_ , \new_[16629]_ ,
    \new_[16630]_ , \new_[16631]_ , \new_[16632]_ , \new_[16633]_ ,
    \new_[16634]_ , \new_[16635]_ , \new_[16636]_ , \new_[16637]_ ,
    \new_[16638]_ , \new_[16639]_ , \new_[16640]_ , \new_[16641]_ ,
    \new_[16642]_ , \new_[16643]_ , \new_[16644]_ , \new_[16645]_ ,
    \new_[16646]_ , \new_[16647]_ , \new_[16648]_ , \new_[16649]_ ,
    \new_[16650]_ , \new_[16651]_ , \new_[16652]_ , \new_[16653]_ ,
    \new_[16654]_ , \new_[16655]_ , \new_[16656]_ , \new_[16657]_ ,
    \new_[16658]_ , \new_[16659]_ , \new_[16660]_ , \new_[16661]_ ,
    \new_[16662]_ , \new_[16663]_ , \new_[16664]_ , \new_[16665]_ ,
    \new_[16666]_ , \new_[16667]_ , \new_[16668]_ , \new_[16669]_ ,
    \new_[16670]_ , \new_[16671]_ , \new_[16672]_ , \new_[16673]_ ,
    \new_[16674]_ , \new_[16675]_ , \new_[16676]_ , \new_[16677]_ ,
    \new_[16678]_ , \new_[16679]_ , \new_[16680]_ , \new_[16681]_ ,
    \new_[16682]_ , \new_[16683]_ , \new_[16684]_ , \new_[16685]_ ,
    \new_[16686]_ , \new_[16687]_ , \new_[16688]_ , \new_[16689]_ ,
    \new_[16690]_ , \new_[16691]_ , \new_[16692]_ , \new_[16693]_ ,
    \new_[16694]_ , \new_[16695]_ , \new_[16696]_ , \new_[16697]_ ,
    \new_[16698]_ , \new_[16699]_ , \new_[16700]_ , \new_[16701]_ ,
    \new_[16702]_ , \new_[16703]_ , \new_[16704]_ , \new_[16705]_ ,
    \new_[16706]_ , \new_[16707]_ , \new_[16708]_ , \new_[16709]_ ,
    \new_[16710]_ , \new_[16711]_ , \new_[16712]_ , \new_[16713]_ ,
    \new_[16714]_ , \new_[16715]_ , \new_[16716]_ , \new_[16717]_ ,
    \new_[16718]_ , \new_[16719]_ , \new_[16720]_ , \new_[16721]_ ,
    \new_[16722]_ , \new_[16723]_ , \new_[16724]_ , \new_[16725]_ ,
    \new_[16726]_ , \new_[16731]_ , \new_[16732]_ , \new_[16733]_ ,
    \new_[16734]_ , \new_[16735]_ , \new_[16736]_ , \new_[16737]_ ,
    \new_[16738]_ , \new_[16739]_ , \new_[16740]_ , \new_[16741]_ ,
    \new_[16742]_ , \new_[16743]_ , \new_[16744]_ , \new_[16745]_ ,
    \new_[16746]_ , \new_[16747]_ , \new_[16748]_ , \new_[16749]_ ,
    \new_[16750]_ , \new_[16751]_ , \new_[16752]_ , \new_[16753]_ ,
    \new_[16754]_ , \new_[16755]_ , \new_[16756]_ , \new_[16757]_ ,
    \new_[16758]_ , \new_[16759]_ , \new_[16760]_ , \new_[16761]_ ,
    \new_[16762]_ , \new_[16763]_ , \new_[16764]_ , \new_[16765]_ ,
    \new_[16766]_ , \new_[16767]_ , \new_[16768]_ , \new_[16769]_ ,
    \new_[16770]_ , \new_[16771]_ , \new_[16772]_ , \new_[16773]_ ,
    \new_[16774]_ , \new_[16775]_ , \new_[16776]_ , \new_[16777]_ ,
    \new_[16778]_ , \new_[16779]_ , \new_[16780]_ , \new_[16781]_ ,
    \new_[16782]_ , \new_[16783]_ , \new_[16784]_ , \new_[16785]_ ,
    \new_[16786]_ , \new_[16787]_ , \new_[16788]_ , \new_[16789]_ ,
    \new_[16790]_ , \new_[16791]_ , \new_[16792]_ , \new_[16793]_ ,
    \new_[16794]_ , \new_[16795]_ , \new_[16796]_ , \new_[16797]_ ,
    \new_[16798]_ , \new_[16799]_ , \new_[16800]_ , \new_[16801]_ ,
    \new_[16802]_ , \new_[16803]_ , \new_[16804]_ , \new_[16805]_ ,
    \new_[16806]_ , \new_[16807]_ , \new_[16808]_ , \new_[16809]_ ,
    \new_[16810]_ , \new_[16811]_ , \new_[16812]_ , \new_[16813]_ ,
    \new_[16814]_ , \new_[16815]_ , \new_[16816]_ , \new_[16817]_ ,
    \new_[16818]_ , \new_[16819]_ , \new_[16820]_ , \new_[16821]_ ,
    \new_[16822]_ , \new_[16823]_ , \new_[16824]_ , \new_[16825]_ ,
    \new_[16826]_ , \new_[16827]_ , \new_[16828]_ , \new_[16829]_ ,
    \new_[16830]_ , \new_[16831]_ , \new_[16832]_ , \new_[16833]_ ,
    \new_[16834]_ , \new_[16835]_ , \new_[16836]_ , \new_[16837]_ ,
    \new_[16838]_ , \new_[16839]_ , \new_[16840]_ , \new_[16841]_ ,
    \new_[16842]_ , \new_[16843]_ , \new_[16844]_ , \new_[16845]_ ,
    \new_[16846]_ , \new_[16847]_ , \new_[16848]_ , \new_[16849]_ ,
    \new_[16850]_ , \new_[16851]_ , \new_[16852]_ , \new_[16853]_ ,
    \new_[16854]_ , \new_[16855]_ , \new_[16856]_ , \new_[16857]_ ,
    \new_[16858]_ , \new_[16859]_ , \new_[16860]_ , \new_[16861]_ ,
    \new_[16862]_ , \new_[16863]_ , \new_[16864]_ , \new_[16865]_ ,
    \new_[16866]_ , \new_[16867]_ , \new_[16868]_ , \new_[16869]_ ,
    \new_[16870]_ , \new_[16871]_ , \new_[16872]_ , \new_[16873]_ ,
    \new_[16874]_ , \new_[16875]_ , \new_[16876]_ , \new_[16877]_ ,
    \new_[16878]_ , \new_[16879]_ , \new_[16880]_ , \new_[16881]_ ,
    \new_[16882]_ , \new_[16883]_ , \new_[16884]_ , \new_[16885]_ ,
    \new_[16886]_ , \new_[16887]_ , \new_[16888]_ , \new_[16889]_ ,
    \new_[16890]_ , \new_[16891]_ , \new_[16892]_ , \new_[16893]_ ,
    \new_[16894]_ , \new_[16895]_ , \new_[16896]_ , \new_[16897]_ ,
    \new_[16898]_ , \new_[16899]_ , \new_[16900]_ , \new_[16901]_ ,
    \new_[16902]_ , \new_[16903]_ , \new_[16904]_ , \new_[16905]_ ,
    \new_[16906]_ , \new_[16907]_ , \new_[16908]_ , \new_[16909]_ ,
    \new_[16910]_ , \new_[16911]_ , \new_[16912]_ , \new_[16913]_ ,
    \new_[16914]_ , \new_[16915]_ , \new_[16916]_ , \new_[16917]_ ,
    \new_[16918]_ , \new_[16919]_ , \new_[16920]_ , \new_[16921]_ ,
    \new_[16922]_ , \new_[16923]_ , \new_[16924]_ , \new_[16925]_ ,
    \new_[16926]_ , \new_[16927]_ , \new_[16928]_ , \new_[16929]_ ,
    \new_[16930]_ , \new_[16931]_ , \new_[16932]_ , \new_[16933]_ ,
    \new_[16934]_ , \new_[16935]_ , \new_[16936]_ , \new_[16937]_ ,
    \new_[16938]_ , \new_[16939]_ , \new_[16940]_ , \new_[16941]_ ,
    \new_[16942]_ , \new_[16943]_ , \new_[16944]_ , \new_[16945]_ ,
    \new_[16946]_ , \new_[16947]_ , \new_[16948]_ , \new_[16949]_ ,
    \new_[16950]_ , \new_[16951]_ , \new_[16952]_ , \new_[16953]_ ,
    \new_[16954]_ , \new_[16955]_ , \new_[16956]_ , \new_[16957]_ ,
    \new_[16958]_ , \new_[16959]_ , \new_[16960]_ , \new_[16961]_ ,
    \new_[16962]_ , \new_[16963]_ , \new_[16964]_ , \new_[16965]_ ,
    \new_[16966]_ , \new_[16967]_ , \new_[16968]_ , \new_[16969]_ ,
    \new_[16970]_ , \new_[16971]_ , \new_[16972]_ , \new_[16973]_ ,
    \new_[16974]_ , \new_[16975]_ , \new_[16976]_ , \new_[16977]_ ,
    \new_[16978]_ , \new_[16979]_ , \new_[16980]_ , \new_[16981]_ ,
    \new_[16982]_ , \new_[16983]_ , \new_[16984]_ , \new_[16985]_ ,
    \new_[16986]_ , \new_[16987]_ , \new_[16988]_ , \new_[16989]_ ,
    \new_[16990]_ , \new_[16991]_ , \new_[16992]_ , \new_[16993]_ ,
    \new_[16994]_ , \new_[16995]_ , \new_[16996]_ , \new_[16997]_ ,
    \new_[16998]_ , \new_[16999]_ , \new_[17000]_ , \new_[17001]_ ,
    \new_[17002]_ , \new_[17003]_ , \new_[17004]_ , \new_[17005]_ ,
    \new_[17006]_ , \new_[17007]_ , \new_[17008]_ , \new_[17009]_ ,
    \new_[17010]_ , \new_[17011]_ , \new_[17012]_ , \new_[17013]_ ,
    \new_[17014]_ , \new_[17015]_ , \new_[17016]_ , \new_[17017]_ ,
    \new_[17018]_ , \new_[17019]_ , \new_[17020]_ , \new_[17021]_ ,
    \new_[17022]_ , \new_[17023]_ , \new_[17024]_ , \new_[17025]_ ,
    \new_[17026]_ , \new_[17027]_ , \new_[17028]_ , \new_[17029]_ ,
    \new_[17030]_ , \new_[17031]_ , \new_[17032]_ , \new_[17033]_ ,
    \new_[17034]_ , \new_[17035]_ , \new_[17036]_ , \new_[17037]_ ,
    \new_[17038]_ , \new_[17039]_ , \new_[17040]_ , \new_[17041]_ ,
    \new_[17042]_ , \new_[17043]_ , \new_[17044]_ , \new_[17045]_ ,
    \new_[17046]_ , \new_[17047]_ , \new_[17048]_ , \new_[17049]_ ,
    \new_[17050]_ , \new_[17051]_ , \new_[17052]_ , \new_[17053]_ ,
    \new_[17054]_ , \new_[17055]_ , \new_[17056]_ , \new_[17057]_ ,
    \new_[17058]_ , \new_[17059]_ , \new_[17060]_ , \new_[17061]_ ,
    \new_[17062]_ , \new_[17063]_ , \new_[17064]_ , \new_[17065]_ ,
    \new_[17066]_ , \new_[17067]_ , \new_[17068]_ , \new_[17069]_ ,
    \new_[17070]_ , \new_[17071]_ , \new_[17072]_ , \new_[17073]_ ,
    \new_[17074]_ , \new_[17075]_ , \new_[17076]_ , \new_[17077]_ ,
    \new_[17078]_ , \new_[17079]_ , \new_[17080]_ , \new_[17081]_ ,
    \new_[17082]_ , \new_[17083]_ , \new_[17084]_ , \new_[17085]_ ,
    \new_[17086]_ , \new_[17087]_ , \new_[17088]_ , \new_[17089]_ ,
    \new_[17090]_ , \new_[17091]_ , \new_[17092]_ , \new_[17093]_ ,
    \new_[17094]_ , \new_[17095]_ , \new_[17096]_ , \new_[17097]_ ,
    \new_[17098]_ , \new_[17099]_ , \new_[17100]_ , \new_[17101]_ ,
    \new_[17102]_ , \new_[17103]_ , \new_[17104]_ , \new_[17105]_ ,
    \new_[17106]_ , \new_[17107]_ , \new_[17108]_ , \new_[17109]_ ,
    \new_[17110]_ , \new_[17111]_ , \new_[17112]_ , \new_[17113]_ ,
    \new_[17114]_ , \new_[17115]_ , \new_[17116]_ , \new_[17117]_ ,
    \new_[17118]_ , \new_[17119]_ , \new_[17120]_ , \new_[17121]_ ,
    \new_[17122]_ , \new_[17123]_ , \new_[17124]_ , \new_[17125]_ ,
    \new_[17126]_ , \new_[17127]_ , \new_[17128]_ , \new_[17129]_ ,
    \new_[17130]_ , \new_[17131]_ , \new_[17132]_ , \new_[17133]_ ,
    \new_[17134]_ , \new_[17135]_ , \new_[17136]_ , \new_[17137]_ ,
    \new_[17138]_ , \new_[17139]_ , \new_[17140]_ , \new_[17141]_ ,
    \new_[17142]_ , \new_[17143]_ , \new_[17144]_ , \new_[17145]_ ,
    \new_[17146]_ , \new_[17147]_ , \new_[17148]_ , \new_[17149]_ ,
    \new_[17150]_ , \new_[17151]_ , \new_[17152]_ , \new_[17153]_ ,
    \new_[17154]_ , \new_[17155]_ , \new_[17156]_ , \new_[17157]_ ,
    \new_[17158]_ , \new_[17159]_ , \new_[17160]_ , \new_[17161]_ ,
    \new_[17162]_ , \new_[17163]_ , \new_[17164]_ , \new_[17165]_ ,
    \new_[17166]_ , \new_[17167]_ , \new_[17168]_ , \new_[17169]_ ,
    \new_[17170]_ , \new_[17171]_ , \new_[17172]_ , \new_[17173]_ ,
    \new_[17174]_ , \new_[17175]_ , \new_[17176]_ , \new_[17177]_ ,
    \new_[17178]_ , \new_[17179]_ , \new_[17180]_ , \new_[17181]_ ,
    \new_[17182]_ , \new_[17183]_ , \new_[17184]_ , \new_[17185]_ ,
    \new_[17186]_ , \new_[17187]_ , \new_[17188]_ , \new_[17189]_ ,
    \new_[17190]_ , \new_[17191]_ , \new_[17192]_ , \new_[17193]_ ,
    \new_[17194]_ , \new_[17195]_ , \new_[17196]_ , \new_[17197]_ ,
    \new_[17198]_ , \new_[17199]_ , \new_[17200]_ , \new_[17201]_ ,
    \new_[17202]_ , \new_[17203]_ , \new_[17204]_ , \new_[17205]_ ,
    \new_[17206]_ , \new_[17207]_ , \new_[17208]_ , \new_[17209]_ ,
    \new_[17210]_ , \new_[17211]_ , \new_[17212]_ , \new_[17213]_ ,
    \new_[17214]_ , \new_[17215]_ , \new_[17216]_ , \new_[17217]_ ,
    \new_[17218]_ , \new_[17219]_ , \new_[17220]_ , \new_[17221]_ ,
    \new_[17222]_ , \new_[17223]_ , \new_[17224]_ , \new_[17225]_ ,
    \new_[17226]_ , \new_[17227]_ , \new_[17228]_ , \new_[17229]_ ,
    \new_[17230]_ , \new_[17231]_ , \new_[17232]_ , \new_[17233]_ ,
    \new_[17234]_ , \new_[17235]_ , \new_[17236]_ , \new_[17237]_ ,
    \new_[17238]_ , \new_[17239]_ , \new_[17240]_ , \new_[17241]_ ,
    \new_[17242]_ , \new_[17243]_ , \new_[17244]_ , \new_[17245]_ ,
    \new_[17246]_ , \new_[17247]_ , \new_[17248]_ , \new_[17249]_ ,
    \new_[17250]_ , \new_[17251]_ , \new_[17252]_ , \new_[17253]_ ,
    \new_[17254]_ , \new_[17255]_ , \new_[17256]_ , \new_[17257]_ ,
    \new_[17258]_ , \new_[17259]_ , \new_[17260]_ , \new_[17261]_ ,
    \new_[17262]_ , \new_[17263]_ , \new_[17264]_ , \new_[17265]_ ,
    \new_[17266]_ , \new_[17267]_ , \new_[17268]_ , \new_[17269]_ ,
    \new_[17270]_ , \new_[17271]_ , \new_[17272]_ , \new_[17273]_ ,
    \new_[17274]_ , \new_[17275]_ , \new_[17276]_ , \new_[17277]_ ,
    \new_[17278]_ , \new_[17279]_ , \new_[17280]_ , \new_[17281]_ ,
    \new_[17282]_ , \new_[17283]_ , \new_[17284]_ , \new_[17285]_ ,
    \new_[17286]_ , \new_[17287]_ , \new_[17288]_ , \new_[17289]_ ,
    \new_[17290]_ , \new_[17291]_ , \new_[17292]_ , \new_[17293]_ ,
    \new_[17294]_ , \new_[17295]_ , \new_[17296]_ , \new_[17297]_ ,
    \new_[17298]_ , \new_[17299]_ , \new_[17300]_ , \new_[17301]_ ,
    \new_[17302]_ , \new_[17303]_ , \new_[17304]_ , \new_[17305]_ ,
    \new_[17306]_ , \new_[17307]_ , \new_[17308]_ , \new_[17309]_ ,
    \new_[17310]_ , \new_[17311]_ , \new_[17312]_ , \new_[17313]_ ,
    \new_[17314]_ , \new_[17315]_ , \new_[17316]_ , \new_[17317]_ ,
    \new_[17318]_ , \new_[17319]_ , \new_[17320]_ , \new_[17321]_ ,
    \new_[17322]_ , \new_[17323]_ , \new_[17324]_ , \new_[17325]_ ,
    \new_[17326]_ , \new_[17327]_ , \new_[17328]_ , \new_[17329]_ ,
    \new_[17330]_ , \new_[17331]_ , \new_[17332]_ , \new_[17333]_ ,
    \new_[17334]_ , \new_[17335]_ , \new_[17336]_ , \new_[17337]_ ,
    \new_[17338]_ , \new_[17339]_ , \new_[17340]_ , \new_[17341]_ ,
    \new_[17342]_ , \new_[17343]_ , \new_[17344]_ , \new_[17345]_ ,
    \new_[17346]_ , \new_[17347]_ , \new_[17348]_ , \new_[17349]_ ,
    \new_[17350]_ , \new_[17351]_ , \new_[17352]_ , \new_[17353]_ ,
    \new_[17354]_ , \new_[17355]_ , \new_[17356]_ , \new_[17357]_ ,
    \new_[17358]_ , \new_[17359]_ , \new_[17360]_ , \new_[17361]_ ,
    \new_[17362]_ , \new_[17363]_ , \new_[17364]_ , \new_[17365]_ ,
    \new_[17366]_ , \new_[17367]_ , \new_[17368]_ , \new_[17369]_ ,
    \new_[17370]_ , \new_[17371]_ , \new_[17372]_ , \new_[17373]_ ,
    \new_[17377]_ , \new_[17378]_ , \new_[17379]_ , \new_[17380]_ ,
    \new_[17381]_ , \new_[17382]_ , \new_[17383]_ , \new_[17384]_ ,
    \new_[17385]_ , \new_[17386]_ , \new_[17387]_ , \new_[17388]_ ,
    \new_[17389]_ , \new_[17390]_ , \new_[17391]_ , \new_[17392]_ ,
    \new_[17393]_ , \new_[17394]_ , \new_[17395]_ , \new_[17396]_ ,
    \new_[17397]_ , \new_[17398]_ , \new_[17399]_ , \new_[17400]_ ,
    \new_[17401]_ , \new_[17402]_ , \new_[17403]_ , \new_[17404]_ ,
    \new_[17405]_ , \new_[17406]_ , \new_[17407]_ , \new_[17408]_ ,
    \new_[17409]_ , \new_[17410]_ , \new_[17411]_ , \new_[17412]_ ,
    \new_[17413]_ , \new_[17414]_ , \new_[17415]_ , \new_[17416]_ ,
    \new_[17417]_ , \new_[17418]_ , \new_[17419]_ , \new_[17420]_ ,
    \new_[17421]_ , \new_[17422]_ , \new_[17423]_ , \new_[17424]_ ,
    \new_[17425]_ , \new_[17426]_ , \new_[17427]_ , \new_[17428]_ ,
    \new_[17429]_ , \new_[17430]_ , \new_[17431]_ , \new_[17432]_ ,
    \new_[17433]_ , \new_[17434]_ , \new_[17435]_ , \new_[17436]_ ,
    \new_[17437]_ , \new_[17438]_ , \new_[17439]_ , \new_[17440]_ ,
    \new_[17441]_ , \new_[17442]_ , \new_[17443]_ , \new_[17444]_ ,
    \new_[17445]_ , \new_[17446]_ , \new_[17447]_ , \new_[17448]_ ,
    \new_[17449]_ , \new_[17450]_ , \new_[17451]_ , \new_[17452]_ ,
    \new_[17453]_ , \new_[17454]_ , \new_[17455]_ , \new_[17456]_ ,
    \new_[17457]_ , \new_[17458]_ , \new_[17459]_ , \new_[17460]_ ,
    \new_[17461]_ , \new_[17462]_ , \new_[17463]_ , \new_[17464]_ ,
    \new_[17465]_ , \new_[17466]_ , \new_[17467]_ , \new_[17468]_ ,
    \new_[17469]_ , \new_[17470]_ , \new_[17471]_ , \new_[17472]_ ,
    \new_[17473]_ , \new_[17474]_ , \new_[17475]_ , \new_[17476]_ ,
    \new_[17477]_ , \new_[17478]_ , \new_[17479]_ , \new_[17480]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17483]_ , \new_[17484]_ ,
    \new_[17485]_ , \new_[17486]_ , \new_[17487]_ , \new_[17488]_ ,
    \new_[17489]_ , \new_[17490]_ , \new_[17491]_ , \new_[17492]_ ,
    \new_[17493]_ , \new_[17494]_ , \new_[17495]_ , \new_[17496]_ ,
    \new_[17497]_ , \new_[17498]_ , \new_[17499]_ , \new_[17500]_ ,
    \new_[17501]_ , \new_[17502]_ , \new_[17503]_ , \new_[17504]_ ,
    \new_[17505]_ , \new_[17506]_ , \new_[17507]_ , \new_[17508]_ ,
    \new_[17509]_ , \new_[17510]_ , \new_[17511]_ , \new_[17512]_ ,
    \new_[17513]_ , \new_[17514]_ , \new_[17515]_ , \new_[17516]_ ,
    \new_[17517]_ , \new_[17518]_ , \new_[17519]_ , \new_[17520]_ ,
    \new_[17521]_ , \new_[17522]_ , \new_[17523]_ , \new_[17524]_ ,
    \new_[17525]_ , \new_[17526]_ , \new_[17527]_ , \new_[17528]_ ,
    \new_[17529]_ , \new_[17530]_ , \new_[17531]_ , \new_[17532]_ ,
    \new_[17533]_ , \new_[17534]_ , \new_[17535]_ , \new_[17536]_ ,
    \new_[17537]_ , \new_[17538]_ , \new_[17539]_ , \new_[17540]_ ,
    \new_[17541]_ , \new_[17542]_ , \new_[17543]_ , \new_[17544]_ ,
    \new_[17545]_ , \new_[17546]_ , \new_[17547]_ , \new_[17548]_ ,
    \new_[17549]_ , \new_[17550]_ , \new_[17551]_ , \new_[17552]_ ,
    \new_[17553]_ , \new_[17554]_ , \new_[17555]_ , \new_[17556]_ ,
    \new_[17557]_ , \new_[17558]_ , \new_[17559]_ , \new_[17560]_ ,
    \new_[17561]_ , \new_[17562]_ , \new_[17563]_ , \new_[17564]_ ,
    \new_[17565]_ , \new_[17566]_ , \new_[17567]_ , \new_[17568]_ ,
    \new_[17569]_ , \new_[17570]_ , \new_[17571]_ , \new_[17572]_ ,
    \new_[17573]_ , \new_[17574]_ , \new_[17575]_ , \new_[17582]_ ,
    \new_[17583]_ , \new_[17584]_ , \new_[17585]_ , \new_[17586]_ ,
    \new_[17587]_ , \new_[17588]_ , \new_[17589]_ , \new_[17590]_ ,
    \new_[17591]_ , \new_[17592]_ , \new_[17593]_ , \new_[17594]_ ,
    \new_[17595]_ , \new_[17596]_ , \new_[17597]_ , \new_[17598]_ ,
    \new_[17599]_ , \new_[17600]_ , \new_[17601]_ , \new_[17602]_ ,
    \new_[17603]_ , \new_[17604]_ , \new_[17605]_ , \new_[17606]_ ,
    \new_[17607]_ , \new_[17608]_ , \new_[17609]_ , \new_[17610]_ ,
    \new_[17611]_ , \new_[17612]_ , \new_[17613]_ , \new_[17614]_ ,
    \new_[17615]_ , \new_[17616]_ , \new_[17617]_ , \new_[17618]_ ,
    \new_[17619]_ , \new_[17620]_ , \new_[17621]_ , \new_[17622]_ ,
    \new_[17623]_ , \new_[17624]_ , \new_[17625]_ , \new_[17626]_ ,
    \new_[17627]_ , \new_[17628]_ , \new_[17629]_ , \new_[17630]_ ,
    \new_[17631]_ , \new_[17632]_ , \new_[17633]_ , \new_[17634]_ ,
    \new_[17635]_ , \new_[17636]_ , \new_[17637]_ , \new_[17638]_ ,
    \new_[17639]_ , \new_[17640]_ , \new_[17641]_ , \new_[17642]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17645]_ , \new_[17646]_ ,
    \new_[17647]_ , \new_[17648]_ , \new_[17649]_ , \new_[17650]_ ,
    \new_[17651]_ , \new_[17652]_ , \new_[17653]_ , \new_[17654]_ ,
    \new_[17655]_ , \new_[17656]_ , \new_[17657]_ , \new_[17658]_ ,
    \new_[17659]_ , \new_[17660]_ , \new_[17661]_ , \new_[17662]_ ,
    \new_[17663]_ , \new_[17664]_ , \new_[17665]_ , \new_[17666]_ ,
    \new_[17667]_ , \new_[17668]_ , \new_[17669]_ , \new_[17670]_ ,
    \new_[17671]_ , \new_[17672]_ , \new_[17673]_ , \new_[17674]_ ,
    \new_[17675]_ , \new_[17676]_ , \new_[17677]_ , \new_[17678]_ ,
    \new_[17679]_ , \new_[17680]_ , \new_[17681]_ , \new_[17682]_ ,
    \new_[17683]_ , \new_[17684]_ , \new_[17685]_ , \new_[17686]_ ,
    \new_[17687]_ , \new_[17688]_ , \new_[17689]_ , \new_[17690]_ ,
    \new_[17691]_ , \new_[17692]_ , \new_[17693]_ , \new_[17694]_ ,
    \new_[17695]_ , \new_[17696]_ , \new_[17697]_ , \new_[17698]_ ,
    \new_[17699]_ , \new_[17700]_ , \new_[17701]_ , \new_[17702]_ ,
    \new_[17703]_ , \new_[17704]_ , \new_[17705]_ , \new_[17706]_ ,
    \new_[17707]_ , \new_[17708]_ , \new_[17709]_ , \new_[17710]_ ,
    \new_[17711]_ , \new_[17712]_ , \new_[17713]_ , \new_[17714]_ ,
    \new_[17715]_ , \new_[17716]_ , \new_[17717]_ , \new_[17718]_ ,
    \new_[17719]_ , \new_[17720]_ , \new_[17721]_ , \new_[17722]_ ,
    \new_[17723]_ , \new_[17724]_ , \new_[17725]_ , \new_[17726]_ ,
    \new_[17727]_ , \new_[17728]_ , \new_[17729]_ , \new_[17730]_ ,
    \new_[17731]_ , \new_[17732]_ , \new_[17733]_ , \new_[17734]_ ,
    \new_[17735]_ , \new_[17736]_ , \new_[17737]_ , \new_[17738]_ ,
    \new_[17739]_ , \new_[17740]_ , \new_[17741]_ , \new_[17742]_ ,
    \new_[17743]_ , \new_[17744]_ , \new_[17745]_ , \new_[17746]_ ,
    \new_[17747]_ , \new_[17748]_ , \new_[17749]_ , \new_[17750]_ ,
    \new_[17751]_ , \new_[17752]_ , \new_[17753]_ , \new_[17754]_ ,
    \new_[17755]_ , \new_[17756]_ , \new_[17757]_ , \new_[17758]_ ,
    \new_[17759]_ , \new_[17760]_ , \new_[17761]_ , \new_[17762]_ ,
    \new_[17763]_ , \new_[17764]_ , \new_[17765]_ , \new_[17766]_ ,
    \new_[17767]_ , \new_[17768]_ , \new_[17769]_ , \new_[17770]_ ,
    \new_[17771]_ , \new_[17772]_ , \new_[17773]_ , \new_[17774]_ ,
    \new_[17775]_ , \new_[17776]_ , \new_[17777]_ , \new_[17778]_ ,
    \new_[17779]_ , \new_[17780]_ , \new_[17781]_ , \new_[17782]_ ,
    \new_[17783]_ , \new_[17784]_ , \new_[17785]_ , \new_[17786]_ ,
    \new_[17787]_ , \new_[17788]_ , \new_[17789]_ , \new_[17790]_ ,
    \new_[17791]_ , \new_[17792]_ , \new_[17793]_ , \new_[17794]_ ,
    \new_[17795]_ , \new_[17796]_ , \new_[17797]_ , \new_[17798]_ ,
    \new_[17799]_ , \new_[17800]_ , \new_[17801]_ , \new_[17802]_ ,
    \new_[17803]_ , \new_[17804]_ , \new_[17805]_ , \new_[17806]_ ,
    \new_[17807]_ , \new_[17808]_ , \new_[17809]_ , \new_[17810]_ ,
    \new_[17811]_ , \new_[17812]_ , \new_[17813]_ , \new_[17814]_ ,
    \new_[17815]_ , \new_[17816]_ , \new_[17817]_ , \new_[17818]_ ,
    \new_[17819]_ , \new_[17820]_ , \new_[17821]_ , \new_[17822]_ ,
    \new_[17823]_ , \new_[17824]_ , \new_[17825]_ , \new_[17826]_ ,
    \new_[17827]_ , \new_[17828]_ , \new_[17829]_ , \new_[17830]_ ,
    \new_[17831]_ , \new_[17832]_ , \new_[17833]_ , \new_[17834]_ ,
    \new_[17835]_ , \new_[17836]_ , \new_[17837]_ , \new_[17838]_ ,
    \new_[17839]_ , \new_[17840]_ , \new_[17841]_ , \new_[17842]_ ,
    \new_[17843]_ , \new_[17844]_ , \new_[17845]_ , \new_[17846]_ ,
    \new_[17847]_ , \new_[17848]_ , \new_[17849]_ , \new_[17850]_ ,
    \new_[17851]_ , \new_[17852]_ , \new_[17853]_ , \new_[17854]_ ,
    \new_[17855]_ , \new_[17856]_ , \new_[17857]_ , \new_[17858]_ ,
    \new_[17859]_ , \new_[17860]_ , \new_[17861]_ , \new_[17862]_ ,
    \new_[17863]_ , \new_[17864]_ , \new_[17865]_ , \new_[17866]_ ,
    \new_[17867]_ , \new_[17868]_ , \new_[17869]_ , \new_[17870]_ ,
    \new_[17871]_ , \new_[17872]_ , \new_[17873]_ , \new_[17874]_ ,
    \new_[17875]_ , \new_[17876]_ , \new_[17877]_ , \new_[17878]_ ,
    \new_[17879]_ , \new_[17880]_ , \new_[17881]_ , \new_[17882]_ ,
    \new_[17883]_ , \new_[17884]_ , \new_[17885]_ , \new_[17886]_ ,
    \new_[17887]_ , \new_[17888]_ , \new_[17889]_ , \new_[17890]_ ,
    \new_[17891]_ , \new_[17892]_ , \new_[17893]_ , \new_[17894]_ ,
    \new_[17895]_ , \new_[17896]_ , \new_[17897]_ , \new_[17898]_ ,
    \new_[17899]_ , \new_[17900]_ , \new_[17901]_ , \new_[17902]_ ,
    \new_[17903]_ , \new_[17904]_ , \new_[17905]_ , \new_[17906]_ ,
    \new_[17907]_ , \new_[17908]_ , \new_[17909]_ , \new_[17910]_ ,
    \new_[17911]_ , \new_[17912]_ , \new_[17913]_ , \new_[17914]_ ,
    \new_[17915]_ , \new_[17916]_ , \new_[17917]_ , \new_[17918]_ ,
    \new_[17919]_ , \new_[17920]_ , \new_[17921]_ , \new_[17922]_ ,
    \new_[17923]_ , \new_[17924]_ , \new_[17925]_ , \new_[17926]_ ,
    \new_[17927]_ , \new_[17928]_ , \new_[17929]_ , \new_[17930]_ ,
    \new_[17931]_ , \new_[17932]_ , \new_[17933]_ , \new_[17934]_ ,
    \new_[17935]_ , \new_[17936]_ , \new_[17937]_ , \new_[17938]_ ,
    \new_[17939]_ , \new_[17940]_ , \new_[17941]_ , \new_[17942]_ ,
    \new_[17943]_ , \new_[17944]_ , \new_[17945]_ , \new_[17946]_ ,
    \new_[17947]_ , \new_[17948]_ , \new_[17949]_ , \new_[17950]_ ,
    \new_[17951]_ , \new_[17952]_ , \new_[17953]_ , \new_[17954]_ ,
    \new_[17955]_ , \new_[17956]_ , \new_[17957]_ , \new_[17958]_ ,
    \new_[17959]_ , \new_[17960]_ , \new_[17961]_ , \new_[17962]_ ,
    \new_[17963]_ , \new_[17964]_ , \new_[17965]_ , \new_[17966]_ ,
    \new_[17967]_ , \new_[17968]_ , \new_[17969]_ , \new_[17970]_ ,
    \new_[17971]_ , \new_[17972]_ , \new_[17973]_ , \new_[17974]_ ,
    \new_[17975]_ , \new_[17976]_ , \new_[17977]_ , \new_[17978]_ ,
    \new_[17979]_ , \new_[17980]_ , \new_[17981]_ , \new_[17982]_ ,
    \new_[17983]_ , \new_[17984]_ , \new_[17985]_ , \new_[17986]_ ,
    \new_[17987]_ , \new_[17988]_ , \new_[17989]_ , \new_[17990]_ ,
    \new_[17991]_ , \new_[17992]_ , \new_[17993]_ , \new_[17994]_ ,
    \new_[17995]_ , \new_[17996]_ , \new_[17997]_ , \new_[17998]_ ,
    \new_[17999]_ , \new_[18000]_ , \new_[18001]_ , \new_[18002]_ ,
    \new_[18003]_ , \new_[18004]_ , \new_[18005]_ , \new_[18006]_ ,
    \new_[18007]_ , \new_[18008]_ , \new_[18009]_ , \new_[18010]_ ,
    \new_[18011]_ , \new_[18012]_ , \new_[18013]_ , \new_[18014]_ ,
    \new_[18015]_ , \new_[18016]_ , \new_[18017]_ , \new_[18018]_ ,
    \new_[18019]_ , \new_[18020]_ , \new_[18021]_ , \new_[18022]_ ,
    \new_[18023]_ , \new_[18024]_ , \new_[18025]_ , \new_[18026]_ ,
    \new_[18027]_ , \new_[18028]_ , \new_[18029]_ , \new_[18030]_ ,
    \new_[18031]_ , \new_[18032]_ , \new_[18033]_ , \new_[18034]_ ,
    \new_[18035]_ , \new_[18036]_ , \new_[18037]_ , \new_[18038]_ ,
    \new_[18039]_ , \new_[18040]_ , \new_[18041]_ , \new_[18042]_ ,
    \new_[18043]_ , \new_[18044]_ , \new_[18045]_ , \new_[18046]_ ,
    \new_[18047]_ , \new_[18048]_ , \new_[18049]_ , \new_[18050]_ ,
    \new_[18051]_ , \new_[18052]_ , \new_[18053]_ , \new_[18054]_ ,
    \new_[18055]_ , \new_[18056]_ , \new_[18057]_ , \new_[18058]_ ,
    \new_[18059]_ , \new_[18060]_ , \new_[18061]_ , \new_[18062]_ ,
    \new_[18063]_ , \new_[18064]_ , \new_[18065]_ , \new_[18066]_ ,
    \new_[18067]_ , \new_[18068]_ , \new_[18069]_ , \new_[18070]_ ,
    \new_[18071]_ , \new_[18072]_ , \new_[18073]_ , \new_[18074]_ ,
    \new_[18075]_ , \new_[18076]_ , \new_[18077]_ , \new_[18078]_ ,
    \new_[18079]_ , \new_[18080]_ , \new_[18081]_ , \new_[18082]_ ,
    \new_[18083]_ , \new_[18084]_ , \new_[18085]_ , \new_[18086]_ ,
    \new_[18087]_ , \new_[18088]_ , \new_[18089]_ , \new_[18090]_ ,
    \new_[18091]_ , \new_[18092]_ , \new_[18093]_ , \new_[18094]_ ,
    \new_[18095]_ , \new_[18096]_ , \new_[18097]_ , \new_[18098]_ ,
    \new_[18099]_ , \new_[18100]_ , \new_[18101]_ , \new_[18102]_ ,
    \new_[18103]_ , \new_[18104]_ , \new_[18105]_ , \new_[18106]_ ,
    \new_[18107]_ , \new_[18108]_ , \new_[18109]_ , \new_[18110]_ ,
    \new_[18111]_ , \new_[18112]_ , \new_[18113]_ , \new_[18114]_ ,
    \new_[18115]_ , \new_[18116]_ , \new_[18117]_ , \new_[18118]_ ,
    \new_[18119]_ , \new_[18120]_ , \new_[18121]_ , \new_[18122]_ ,
    \new_[18123]_ , \new_[18124]_ , \new_[18125]_ , \new_[18126]_ ,
    \new_[18127]_ , \new_[18128]_ , \new_[18129]_ , \new_[18130]_ ,
    \new_[18131]_ , \new_[18132]_ , \new_[18133]_ , \new_[18134]_ ,
    \new_[18135]_ , \new_[18136]_ , \new_[18137]_ , \new_[18138]_ ,
    \new_[18139]_ , \new_[18140]_ , \new_[18141]_ , \new_[18142]_ ,
    \new_[18143]_ , \new_[18144]_ , \new_[18145]_ , \new_[18146]_ ,
    \new_[18147]_ , \new_[18148]_ , \new_[18149]_ , \new_[18150]_ ,
    \new_[18151]_ , \new_[18152]_ , \new_[18153]_ , \new_[18154]_ ,
    \new_[18155]_ , \new_[18156]_ , \new_[18157]_ , \new_[18158]_ ,
    \new_[18159]_ , \new_[18160]_ , \new_[18161]_ , \new_[18162]_ ,
    \new_[18163]_ , \new_[18164]_ , \new_[18165]_ , \new_[18166]_ ,
    \new_[18167]_ , \new_[18168]_ , \new_[18169]_ , \new_[18170]_ ,
    \new_[18171]_ , \new_[18172]_ , \new_[18173]_ , \new_[18174]_ ,
    \new_[18175]_ , \new_[18176]_ , \new_[18177]_ , \new_[18178]_ ,
    \new_[18179]_ , \new_[18180]_ , \new_[18181]_ , \new_[18182]_ ,
    \new_[18183]_ , \new_[18184]_ , \new_[18185]_ , \new_[18186]_ ,
    \new_[18187]_ , \new_[18188]_ , \new_[18189]_ , \new_[18190]_ ,
    \new_[18191]_ , \new_[18192]_ , \new_[18193]_ , \new_[18194]_ ,
    \new_[18195]_ , \new_[18196]_ , \new_[18197]_ , \new_[18198]_ ,
    \new_[18199]_ , \new_[18200]_ , \new_[18201]_ , \new_[18202]_ ,
    \new_[18203]_ , \new_[18204]_ , \new_[18205]_ , \new_[18206]_ ,
    \new_[18207]_ , \new_[18208]_ , \new_[18209]_ , \new_[18210]_ ,
    \new_[18211]_ , \new_[18212]_ , \new_[18213]_ , \new_[18214]_ ,
    \new_[18215]_ , \new_[18216]_ , \new_[18217]_ , \new_[18218]_ ,
    \new_[18219]_ , \new_[18220]_ , \new_[18221]_ , \new_[18222]_ ,
    \new_[18223]_ , \new_[18224]_ , \new_[18225]_ , \new_[18226]_ ,
    \new_[18227]_ , \new_[18228]_ , \new_[18229]_ , \new_[18230]_ ,
    \new_[18231]_ , \new_[18232]_ , \new_[18233]_ , \new_[18234]_ ,
    \new_[18235]_ , \new_[18236]_ , \new_[18237]_ , \new_[18238]_ ,
    \new_[18239]_ , \new_[18240]_ , \new_[18241]_ , \new_[18242]_ ,
    \new_[18243]_ , \new_[18244]_ , \new_[18245]_ , \new_[18246]_ ,
    \new_[18247]_ , \new_[18248]_ , \new_[18249]_ , \new_[18250]_ ,
    \new_[18251]_ , \new_[18252]_ , \new_[18253]_ , \new_[18254]_ ,
    \new_[18255]_ , \new_[18256]_ , \new_[18257]_ , \new_[18258]_ ,
    \new_[18259]_ , \new_[18260]_ , \new_[18261]_ , \new_[18262]_ ,
    \new_[18263]_ , \new_[18264]_ , \new_[18265]_ , \new_[18266]_ ,
    \new_[18267]_ , \new_[18268]_ , \new_[18269]_ , \new_[18270]_ ,
    \new_[18271]_ , \new_[18272]_ , \new_[18273]_ , \new_[18274]_ ,
    \new_[18275]_ , \new_[18276]_ , \new_[18277]_ , \new_[18278]_ ,
    \new_[18279]_ , \new_[18280]_ , \new_[18281]_ , \new_[18282]_ ,
    \new_[18283]_ , \new_[18284]_ , \new_[18285]_ , \new_[18286]_ ,
    \new_[18287]_ , \new_[18288]_ , \new_[18289]_ , \new_[18290]_ ,
    \new_[18291]_ , \new_[18292]_ , \new_[18293]_ , \new_[18294]_ ,
    \new_[18295]_ , \new_[18296]_ , \new_[18297]_ , \new_[18298]_ ,
    \new_[18299]_ , \new_[18300]_ , \new_[18301]_ , \new_[18302]_ ,
    \new_[18303]_ , \new_[18304]_ , \new_[18305]_ , \new_[18306]_ ,
    \new_[18307]_ , \new_[18308]_ , \new_[18309]_ , \new_[18310]_ ,
    \new_[18311]_ , \new_[18312]_ , \new_[18313]_ , \new_[18315]_ ,
    \new_[18316]_ , \new_[18317]_ , \new_[18318]_ , \new_[18319]_ ,
    \new_[18320]_ , \new_[18321]_ , \new_[18322]_ , \new_[18323]_ ,
    \new_[18324]_ , \new_[18325]_ , \new_[18326]_ , \new_[18327]_ ,
    \new_[18328]_ , \new_[18329]_ , \new_[18330]_ , \new_[18331]_ ,
    \new_[18332]_ , \new_[18333]_ , \new_[18334]_ , \new_[18335]_ ,
    \new_[18336]_ , \new_[18337]_ , \new_[18338]_ , \new_[18339]_ ,
    \new_[18340]_ , \new_[18341]_ , \new_[18342]_ , \new_[18343]_ ,
    \new_[18344]_ , \new_[18345]_ , \new_[18346]_ , \new_[18347]_ ,
    \new_[18348]_ , \new_[18349]_ , \new_[18350]_ , \new_[18351]_ ,
    \new_[18352]_ , \new_[18353]_ , \new_[18354]_ , \new_[18355]_ ,
    \new_[18356]_ , \new_[18357]_ , \new_[18358]_ , \new_[18359]_ ,
    \new_[18360]_ , \new_[18361]_ , \new_[18362]_ , \new_[18363]_ ,
    \new_[18364]_ , \new_[18365]_ , \new_[18366]_ , \new_[18367]_ ,
    \new_[18368]_ , \new_[18369]_ , \new_[18370]_ , \new_[18371]_ ,
    \new_[18372]_ , \new_[18373]_ , \new_[18374]_ , \new_[18375]_ ,
    \new_[18376]_ , \new_[18380]_ , \new_[18381]_ , \new_[18382]_ ,
    \new_[18383]_ , \new_[18384]_ , \new_[18385]_ , \new_[18386]_ ,
    \new_[18387]_ , \new_[18389]_ , \new_[18390]_ , \new_[18392]_ ,
    \new_[18396]_ , \new_[18397]_ , \new_[18398]_ , \new_[18399]_ ,
    \new_[18400]_ , \new_[18401]_ , \new_[18402]_ , \new_[18403]_ ,
    \new_[18404]_ , \new_[18405]_ , \new_[18406]_ , \new_[18407]_ ,
    \new_[18408]_ , \new_[18409]_ , \new_[18410]_ , \new_[18411]_ ,
    \new_[18412]_ , \new_[18413]_ , \new_[18414]_ , \new_[18415]_ ,
    \new_[18416]_ , \new_[18417]_ , \new_[18418]_ , \new_[18419]_ ,
    \new_[18420]_ , \new_[18421]_ , \new_[18422]_ , \new_[18423]_ ,
    \new_[18424]_ , \new_[18425]_ , \new_[18426]_ , \new_[18427]_ ,
    \new_[18428]_ , \new_[18429]_ , \new_[18430]_ , \new_[18431]_ ,
    \new_[18432]_ , \new_[18433]_ , \new_[18434]_ , \new_[18435]_ ,
    \new_[18436]_ , \new_[18437]_ , \new_[18438]_ , \new_[18439]_ ,
    \new_[18440]_ , \new_[18441]_ , \new_[18442]_ , \new_[18443]_ ,
    \new_[18444]_ , \new_[18445]_ , \new_[18446]_ , \new_[18447]_ ,
    \new_[18448]_ , \new_[18449]_ , \new_[18450]_ , \new_[18451]_ ,
    \new_[18452]_ , \new_[18453]_ , \new_[18454]_ , \new_[18455]_ ,
    \new_[18456]_ , \new_[18457]_ , \new_[18458]_ , \new_[18459]_ ,
    \new_[18460]_ , \new_[18461]_ , \new_[18462]_ , \new_[18463]_ ,
    \new_[18464]_ , \new_[18465]_ , \new_[18466]_ , \new_[18467]_ ,
    \new_[18468]_ , \new_[18469]_ , \new_[18470]_ , \new_[18471]_ ,
    \new_[18472]_ , \new_[18473]_ , \new_[18474]_ , \new_[18475]_ ,
    \new_[18476]_ , \new_[18477]_ , \new_[18483]_ , \new_[18484]_ ,
    \new_[18485]_ , \new_[18486]_ , \new_[18487]_ , \new_[18488]_ ,
    \new_[18489]_ , \new_[18490]_ , \new_[18491]_ , \new_[18492]_ ,
    \new_[18493]_ , \new_[18494]_ , \new_[18495]_ , \new_[18496]_ ,
    \new_[18497]_ , \new_[18498]_ , \new_[18499]_ , \new_[18500]_ ,
    \new_[18501]_ , \new_[18502]_ , \new_[18503]_ , \new_[18504]_ ,
    \new_[18505]_ , \new_[18506]_ , \new_[18507]_ , \new_[18508]_ ,
    \new_[18509]_ , \new_[18510]_ , \new_[18511]_ , \new_[18512]_ ,
    \new_[18513]_ , \new_[18514]_ , \new_[18515]_ , \new_[18516]_ ,
    \new_[18517]_ , \new_[18518]_ , \new_[18519]_ , \new_[18520]_ ,
    \new_[18521]_ , \new_[18522]_ , \new_[18523]_ , \new_[18524]_ ,
    \new_[18525]_ , \new_[18526]_ , \new_[18527]_ , \new_[18528]_ ,
    \new_[18529]_ , \new_[18530]_ , \new_[18531]_ , \new_[18532]_ ,
    \new_[18533]_ , \new_[18534]_ , \new_[18535]_ , \new_[18536]_ ,
    \new_[18537]_ , \new_[18538]_ , \new_[18539]_ , \new_[18540]_ ,
    \new_[18541]_ , \new_[18542]_ , \new_[18543]_ , \new_[18544]_ ,
    \new_[18545]_ , \new_[18546]_ , \new_[18547]_ , \new_[18548]_ ,
    \new_[18549]_ , \new_[18550]_ , \new_[18551]_ , \new_[18552]_ ,
    \new_[18553]_ , \new_[18554]_ , \new_[18555]_ , \new_[18556]_ ,
    \new_[18557]_ , \new_[18558]_ , \new_[18559]_ , \new_[18560]_ ,
    \new_[18561]_ , \new_[18562]_ , \new_[18563]_ , \new_[18564]_ ,
    \new_[18565]_ , \new_[18566]_ , \new_[18567]_ , \new_[18568]_ ,
    \new_[18569]_ , \new_[18570]_ , \new_[18571]_ , \new_[18572]_ ,
    \new_[18573]_ , \new_[18574]_ , \new_[18575]_ , \new_[18576]_ ,
    \new_[18577]_ , \new_[18578]_ , \new_[18579]_ , \new_[18580]_ ,
    \new_[18581]_ , \new_[18582]_ , \new_[18583]_ , \new_[18584]_ ,
    \new_[18585]_ , \new_[18586]_ , \new_[18587]_ , \new_[18588]_ ,
    \new_[18589]_ , \new_[18590]_ , \new_[18591]_ , \new_[18592]_ ,
    \new_[18593]_ , \new_[18594]_ , \new_[18595]_ , \new_[18596]_ ,
    \new_[18597]_ , \new_[18598]_ , \new_[18599]_ , \new_[18600]_ ,
    \new_[18601]_ , \new_[18602]_ , \new_[18603]_ , \new_[18604]_ ,
    \new_[18605]_ , \new_[18606]_ , \new_[18607]_ , \new_[18608]_ ,
    \new_[18609]_ , \new_[18610]_ , \new_[18611]_ , \new_[18612]_ ,
    \new_[18613]_ , \new_[18614]_ , \new_[18615]_ , \new_[18616]_ ,
    \new_[18617]_ , \new_[18618]_ , \new_[18619]_ , \new_[18620]_ ,
    \new_[18621]_ , \new_[18622]_ , \new_[18623]_ , \new_[18624]_ ,
    \new_[18625]_ , \new_[18626]_ , \new_[18627]_ , \new_[18628]_ ,
    \new_[18629]_ , \new_[18630]_ , \new_[18631]_ , \new_[18632]_ ,
    \new_[18633]_ , \new_[18634]_ , \new_[18635]_ , \new_[18636]_ ,
    \new_[18637]_ , \new_[18638]_ , \new_[18639]_ , \new_[18640]_ ,
    \new_[18641]_ , \new_[18642]_ , \new_[18643]_ , \new_[18644]_ ,
    \new_[18645]_ , \new_[18646]_ , \new_[18647]_ , \new_[18648]_ ,
    \new_[18649]_ , \new_[18650]_ , \new_[18651]_ , \new_[18652]_ ,
    \new_[18653]_ , \new_[18654]_ , \new_[18655]_ , \new_[18656]_ ,
    \new_[18657]_ , \new_[18658]_ , \new_[18659]_ , \new_[18660]_ ,
    \new_[18661]_ , \new_[18662]_ , \new_[18663]_ , \new_[18664]_ ,
    \new_[18665]_ , \new_[18666]_ , \new_[18667]_ , \new_[18668]_ ,
    \new_[18669]_ , \new_[18670]_ , \new_[18671]_ , \new_[18672]_ ,
    \new_[18673]_ , \new_[18674]_ , \new_[18675]_ , \new_[18676]_ ,
    \new_[18677]_ , \new_[18678]_ , \new_[18679]_ , \new_[18680]_ ,
    \new_[18681]_ , \new_[18682]_ , \new_[18683]_ , \new_[18684]_ ,
    \new_[18685]_ , \new_[18686]_ , \new_[18687]_ , \new_[18688]_ ,
    \new_[18689]_ , \new_[18690]_ , \new_[18691]_ , \new_[18692]_ ,
    \new_[18693]_ , \new_[18694]_ , \new_[18695]_ , \new_[18696]_ ,
    \new_[18697]_ , \new_[18698]_ , \new_[18699]_ , \new_[18700]_ ,
    \new_[18701]_ , \new_[18702]_ , \new_[18703]_ , \new_[18704]_ ,
    \new_[18705]_ , \new_[18706]_ , \new_[18707]_ , \new_[18708]_ ,
    \new_[18709]_ , \new_[18710]_ , \new_[18711]_ , \new_[18712]_ ,
    \new_[18713]_ , \new_[18714]_ , \new_[18715]_ , \new_[18716]_ ,
    \new_[18717]_ , \new_[18718]_ , \new_[18719]_ , \new_[18720]_ ,
    \new_[18721]_ , \new_[18722]_ , \new_[18723]_ , \new_[18724]_ ,
    \new_[18725]_ , \new_[18726]_ , \new_[18727]_ , \new_[18728]_ ,
    \new_[18729]_ , \new_[18730]_ , \new_[18731]_ , \new_[18732]_ ,
    \new_[18733]_ , \new_[18734]_ , \new_[18735]_ , \new_[18736]_ ,
    \new_[18737]_ , \new_[18738]_ , \new_[18739]_ , \new_[18740]_ ,
    \new_[18741]_ , \new_[18742]_ , \new_[18743]_ , \new_[18744]_ ,
    \new_[18745]_ , \new_[18746]_ , \new_[18747]_ , \new_[18748]_ ,
    \new_[18749]_ , \new_[18750]_ , \new_[18751]_ , \new_[18752]_ ,
    \new_[18753]_ , \new_[18754]_ , \new_[18755]_ , \new_[18756]_ ,
    \new_[18757]_ , \new_[18758]_ , \new_[18759]_ , \new_[18760]_ ,
    \new_[18761]_ , \new_[18762]_ , \new_[18763]_ , \new_[18764]_ ,
    \new_[18765]_ , \new_[18766]_ , \new_[18767]_ , \new_[18768]_ ,
    \new_[18769]_ , \new_[18770]_ , \new_[18771]_ , \new_[18772]_ ,
    \new_[18773]_ , \new_[18774]_ , \new_[18775]_ , \new_[18776]_ ,
    \new_[18777]_ , \new_[18778]_ , \new_[18779]_ , \new_[18780]_ ,
    \new_[18781]_ , \new_[18782]_ , \new_[18783]_ , \new_[18784]_ ,
    \new_[18785]_ , \new_[18786]_ , \new_[18787]_ , \new_[18788]_ ,
    \new_[18789]_ , \new_[18790]_ , \new_[18791]_ , \new_[18792]_ ,
    \new_[18793]_ , \new_[18794]_ , \new_[18795]_ , \new_[18796]_ ,
    \new_[18797]_ , \new_[18798]_ , \new_[18799]_ , \new_[18800]_ ,
    \new_[18801]_ , \new_[18802]_ , \new_[18803]_ , \new_[18804]_ ,
    \new_[18805]_ , \new_[18806]_ , \new_[18807]_ , \new_[18808]_ ,
    \new_[18809]_ , \new_[18810]_ , \new_[18811]_ , \new_[18812]_ ,
    \new_[18813]_ , \new_[18814]_ , \new_[18815]_ , \new_[18816]_ ,
    \new_[18817]_ , \new_[18818]_ , \new_[18819]_ , \new_[18820]_ ,
    \new_[18821]_ , \new_[18822]_ , \new_[18823]_ , \new_[18824]_ ,
    \new_[18825]_ , \new_[18826]_ , \new_[18827]_ , \new_[18828]_ ,
    \new_[18829]_ , \new_[18830]_ , \new_[18831]_ , \new_[18832]_ ,
    \new_[18833]_ , \new_[18834]_ , \new_[18835]_ , \new_[18836]_ ,
    \new_[18837]_ , \new_[18838]_ , \new_[18839]_ , \new_[18840]_ ,
    \new_[18841]_ , \new_[18842]_ , \new_[18843]_ , \new_[18844]_ ,
    \new_[18845]_ , \new_[18846]_ , \new_[18847]_ , \new_[18848]_ ,
    \new_[18849]_ , \new_[18850]_ , \new_[18851]_ , \new_[18852]_ ,
    \new_[18853]_ , \new_[18854]_ , \new_[18855]_ , \new_[18856]_ ,
    \new_[18857]_ , \new_[18858]_ , \new_[18859]_ , \new_[18860]_ ,
    \new_[18861]_ , \new_[18862]_ , \new_[18863]_ , \new_[18864]_ ,
    \new_[18865]_ , \new_[18866]_ , \new_[18867]_ , \new_[18868]_ ,
    \new_[18869]_ , \new_[18870]_ , \new_[18871]_ , \new_[18872]_ ,
    \new_[18873]_ , \new_[18874]_ , \new_[18875]_ , \new_[18876]_ ,
    \new_[18877]_ , \new_[18878]_ , \new_[18879]_ , \new_[18880]_ ,
    \new_[18881]_ , \new_[18882]_ , \new_[18883]_ , \new_[18884]_ ,
    \new_[18885]_ , \new_[18886]_ , \new_[18887]_ , \new_[18888]_ ,
    \new_[18889]_ , \new_[18890]_ , \new_[18891]_ , \new_[18892]_ ,
    \new_[18893]_ , \new_[18894]_ , \new_[18895]_ , \new_[18896]_ ,
    \new_[18897]_ , \new_[18898]_ , \new_[18899]_ , \new_[18900]_ ,
    \new_[18901]_ , \new_[18902]_ , \new_[18903]_ , \new_[18904]_ ,
    \new_[18905]_ , \new_[18906]_ , \new_[18907]_ , \new_[18908]_ ,
    \new_[18909]_ , \new_[18910]_ , \new_[18911]_ , \new_[18912]_ ,
    \new_[18913]_ , \new_[18914]_ , \new_[18915]_ , \new_[18916]_ ,
    \new_[18917]_ , \new_[18918]_ , \new_[18919]_ , \new_[18920]_ ,
    \new_[18921]_ , \new_[18922]_ , \new_[18923]_ , \new_[18924]_ ,
    \new_[18925]_ , \new_[18926]_ , \new_[18927]_ , \new_[18928]_ ,
    \new_[18929]_ , \new_[18930]_ , \new_[18931]_ , \new_[18932]_ ,
    \new_[18933]_ , \new_[18934]_ , \new_[18935]_ , \new_[18936]_ ,
    \new_[18937]_ , \new_[18938]_ , \new_[18939]_ , \new_[18940]_ ,
    \new_[18941]_ , \new_[18942]_ , \new_[18943]_ , \new_[18944]_ ,
    \new_[18945]_ , \new_[18946]_ , \new_[18947]_ , \new_[18948]_ ,
    \new_[18949]_ , \new_[18950]_ , \new_[18951]_ , \new_[18952]_ ,
    \new_[18953]_ , \new_[18954]_ , \new_[18955]_ , \new_[18956]_ ,
    \new_[18957]_ , \new_[18958]_ , \new_[18959]_ , \new_[18960]_ ,
    \new_[18961]_ , \new_[18962]_ , \new_[18963]_ , \new_[18964]_ ,
    \new_[18965]_ , \new_[18966]_ , \new_[18967]_ , \new_[18968]_ ,
    \new_[18969]_ , \new_[18970]_ , \new_[18971]_ , \new_[18972]_ ,
    \new_[18973]_ , \new_[18974]_ , \new_[18975]_ , \new_[18976]_ ,
    \new_[18977]_ , \new_[18978]_ , \new_[18979]_ , \new_[18980]_ ,
    \new_[18981]_ , \new_[18982]_ , \new_[18983]_ , \new_[18984]_ ,
    \new_[18985]_ , \new_[18986]_ , \new_[18987]_ , \new_[18988]_ ,
    \new_[18989]_ , \new_[18990]_ , \new_[18991]_ , \new_[18992]_ ,
    \new_[18993]_ , \new_[18994]_ , \new_[18995]_ , \new_[18996]_ ,
    \new_[18997]_ , \new_[18998]_ , \new_[18999]_ , \new_[19000]_ ,
    \new_[19001]_ , \new_[19002]_ , \new_[19003]_ , \new_[19004]_ ,
    \new_[19005]_ , \new_[19006]_ , \new_[19007]_ , \new_[19008]_ ,
    \new_[19009]_ , \new_[19010]_ , \new_[19011]_ , \new_[19012]_ ,
    \new_[19013]_ , \new_[19014]_ , \new_[19015]_ , \new_[19016]_ ,
    \new_[19017]_ , \new_[19018]_ , \new_[19019]_ , \new_[19020]_ ,
    \new_[19021]_ , \new_[19022]_ , \new_[19023]_ , \new_[19024]_ ,
    \new_[19025]_ , \new_[19026]_ , \new_[19027]_ , \new_[19028]_ ,
    \new_[19029]_ , \new_[19030]_ , \new_[19031]_ , \new_[19032]_ ,
    \new_[19033]_ , \new_[19034]_ , \new_[19035]_ , \new_[19036]_ ,
    \new_[19037]_ , \new_[19038]_ , \new_[19039]_ , \new_[19040]_ ,
    \new_[19041]_ , \new_[19042]_ , \new_[19043]_ , \new_[19044]_ ,
    \new_[19045]_ , \new_[19046]_ , \new_[19047]_ , \new_[19048]_ ,
    \new_[19049]_ , \new_[19050]_ , \new_[19051]_ , \new_[19052]_ ,
    \new_[19053]_ , \new_[19054]_ , \new_[19055]_ , \new_[19056]_ ,
    \new_[19057]_ , \new_[19058]_ , \new_[19059]_ , \new_[19060]_ ,
    \new_[19061]_ , \new_[19062]_ , \new_[19063]_ , \new_[19064]_ ,
    \new_[19065]_ , \new_[19066]_ , \new_[19067]_ , \new_[19068]_ ,
    \new_[19069]_ , \new_[19070]_ , \new_[19071]_ , \new_[19072]_ ,
    \new_[19073]_ , \new_[19074]_ , \new_[19075]_ , \new_[19076]_ ,
    \new_[19077]_ , \new_[19079]_ , \new_[19080]_ , \new_[19081]_ ,
    \new_[19088]_ , \new_[19089]_ , \new_[19090]_ , \new_[19091]_ ,
    \new_[19092]_ , \new_[19093]_ , \new_[19094]_ , \new_[19095]_ ,
    \new_[19096]_ , \new_[19097]_ , \new_[19098]_ , \new_[19099]_ ,
    \new_[19100]_ , \new_[19101]_ , \new_[19102]_ , \new_[19103]_ ,
    \new_[19104]_ , \new_[19105]_ , \new_[19106]_ , \new_[19107]_ ,
    \new_[19108]_ , \new_[19109]_ , \new_[19110]_ , \new_[19111]_ ,
    \new_[19112]_ , \new_[19113]_ , \new_[19114]_ , \new_[19115]_ ,
    \new_[19116]_ , \new_[19117]_ , \new_[19118]_ , \new_[19119]_ ,
    \new_[19120]_ , \new_[19121]_ , \new_[19122]_ , \new_[19123]_ ,
    \new_[19124]_ , \new_[19125]_ , \new_[19126]_ , \new_[19127]_ ,
    \new_[19128]_ , \new_[19129]_ , \new_[19130]_ , \new_[19131]_ ,
    \new_[19132]_ , \new_[19133]_ , \new_[19134]_ , \new_[19135]_ ,
    \new_[19136]_ , \new_[19137]_ , \new_[19138]_ , \new_[19139]_ ,
    \new_[19140]_ , \new_[19141]_ , \new_[19142]_ , \new_[19143]_ ,
    \new_[19144]_ , \new_[19145]_ , \new_[19146]_ , \new_[19147]_ ,
    \new_[19148]_ , \new_[19149]_ , \new_[19150]_ , \new_[19151]_ ,
    \new_[19152]_ , \new_[19153]_ , \new_[19154]_ , \new_[19155]_ ,
    \new_[19156]_ , \new_[19157]_ , \new_[19158]_ , \new_[19159]_ ,
    \new_[19160]_ , \new_[19161]_ , \new_[19162]_ , \new_[19163]_ ,
    \new_[19164]_ , \new_[19165]_ , \new_[19166]_ , \new_[19167]_ ,
    \new_[19168]_ , \new_[19169]_ , \new_[19170]_ , \new_[19171]_ ,
    \new_[19172]_ , \new_[19173]_ , \new_[19174]_ , \new_[19175]_ ,
    \new_[19176]_ , \new_[19177]_ , \new_[19178]_ , \new_[19179]_ ,
    \new_[19180]_ , \new_[19181]_ , \new_[19182]_ , \new_[19183]_ ,
    \new_[19184]_ , \new_[19185]_ , \new_[19186]_ , \new_[19187]_ ,
    \new_[19188]_ , \new_[19189]_ , \new_[19190]_ , \new_[19191]_ ,
    \new_[19192]_ , \new_[19193]_ , \new_[19194]_ , \new_[19195]_ ,
    \new_[19196]_ , \new_[19197]_ , \new_[19198]_ , \new_[19199]_ ,
    \new_[19200]_ , \new_[19201]_ , \new_[19202]_ , \new_[19203]_ ,
    \new_[19204]_ , \new_[19205]_ , \new_[19206]_ , \new_[19207]_ ,
    \new_[19208]_ , \new_[19209]_ , \new_[19210]_ , \new_[19211]_ ,
    \new_[19212]_ , \new_[19213]_ , \new_[19214]_ , \new_[19215]_ ,
    \new_[19216]_ , \new_[19217]_ , \new_[19218]_ , \new_[19219]_ ,
    \new_[19220]_ , \new_[19221]_ , \new_[19222]_ , \new_[19223]_ ,
    \new_[19224]_ , \new_[19225]_ , \new_[19226]_ , \new_[19227]_ ,
    \new_[19228]_ , \new_[19229]_ , \new_[19230]_ , \new_[19231]_ ,
    \new_[19232]_ , \new_[19233]_ , \new_[19234]_ , \new_[19235]_ ,
    \new_[19236]_ , \new_[19237]_ , \new_[19238]_ , \new_[19239]_ ,
    \new_[19240]_ , \new_[19241]_ , \new_[19242]_ , \new_[19243]_ ,
    \new_[19244]_ , \new_[19245]_ , \new_[19246]_ , \new_[19247]_ ,
    \new_[19248]_ , \new_[19250]_ , \new_[19251]_ , \new_[19252]_ ,
    \new_[19253]_ , \new_[19254]_ , \new_[19255]_ , \new_[19256]_ ,
    \new_[19257]_ , \new_[19258]_ , \new_[19259]_ , \new_[19260]_ ,
    \new_[19261]_ , \new_[19262]_ , \new_[19263]_ , \new_[19264]_ ,
    \new_[19265]_ , \new_[19266]_ , \new_[19267]_ , \new_[19268]_ ,
    \new_[19269]_ , \new_[19270]_ , \new_[19271]_ , \new_[19272]_ ,
    \new_[19273]_ , \new_[19274]_ , \new_[19275]_ , \new_[19276]_ ,
    \new_[19277]_ , \new_[19278]_ , \new_[19279]_ , \new_[19280]_ ,
    \new_[19281]_ , \new_[19283]_ , \new_[19284]_ , \new_[19286]_ ,
    \new_[19287]_ , \new_[19288]_ , \new_[19289]_ , \new_[19290]_ ,
    \new_[19291]_ , \new_[19292]_ , \new_[19293]_ , \new_[19294]_ ,
    \new_[19295]_ , \new_[19296]_ , \new_[19297]_ , \new_[19298]_ ,
    \new_[19299]_ , \new_[19300]_ , \new_[19301]_ , \new_[19302]_ ,
    \new_[19303]_ , \new_[19304]_ , \new_[19305]_ , \new_[19306]_ ,
    \new_[19307]_ , \new_[19308]_ , \new_[19310]_ , \new_[19311]_ ,
    \new_[19312]_ , \new_[19313]_ , \new_[19314]_ , \new_[19315]_ ,
    \new_[19316]_ , \new_[19317]_ , \new_[19318]_ , \new_[19319]_ ,
    \new_[19320]_ , \new_[19321]_ , \new_[19322]_ , \new_[19323]_ ,
    \new_[19324]_ , \new_[19325]_ , \new_[19326]_ , \new_[19327]_ ,
    \new_[19328]_ , \new_[19329]_ , \new_[19330]_ , \new_[19331]_ ,
    \new_[19332]_ , \new_[19333]_ , \new_[19334]_ , \new_[19335]_ ,
    \new_[19336]_ , \new_[19337]_ , \new_[19338]_ , \new_[19339]_ ,
    \new_[19340]_ , \new_[19341]_ , \new_[19342]_ , \new_[19345]_ ,
    \new_[19346]_ , \new_[19347]_ , \new_[19348]_ , \new_[19349]_ ,
    \new_[19350]_ , \new_[19351]_ , \new_[19352]_ , \new_[19353]_ ,
    \new_[19354]_ , \new_[19355]_ , \new_[19356]_ , \new_[19357]_ ,
    \new_[19358]_ , \new_[19360]_ , \new_[19361]_ , \new_[19362]_ ,
    \new_[19363]_ , \new_[19364]_ , \new_[19365]_ , \new_[19366]_ ,
    \new_[19367]_ , \new_[19368]_ , \new_[19369]_ , \new_[19370]_ ,
    \new_[19371]_ , \new_[19372]_ , \new_[19373]_ , \new_[19374]_ ,
    \new_[19375]_ , \new_[19376]_ , \new_[19377]_ , \new_[19378]_ ,
    \new_[19379]_ , \new_[19380]_ , \new_[19381]_ , \new_[19382]_ ,
    \new_[19383]_ , \new_[19384]_ , \new_[19385]_ , \new_[19386]_ ,
    \new_[19387]_ , \new_[19388]_ , \new_[19389]_ , \new_[19390]_ ,
    \new_[19391]_ , \new_[19392]_ , \new_[19393]_ , \new_[19394]_ ,
    \new_[19395]_ , \new_[19396]_ , \new_[19397]_ , \new_[19398]_ ,
    \new_[19399]_ , \new_[19400]_ , \new_[19401]_ , \new_[19402]_ ,
    \new_[19403]_ , \new_[19404]_ , \new_[19405]_ , \new_[19406]_ ,
    \new_[19407]_ , \new_[19408]_ , \new_[19409]_ , \new_[19410]_ ,
    \new_[19411]_ , \new_[19412]_ , \new_[19413]_ , \new_[19414]_ ,
    \new_[19415]_ , \new_[19416]_ , \new_[19417]_ , \new_[19418]_ ,
    \new_[19419]_ , \new_[19420]_ , \new_[19421]_ , \new_[19422]_ ,
    \new_[19423]_ , \new_[19424]_ , \new_[19425]_ , \new_[19426]_ ,
    \new_[19427]_ , \new_[19428]_ , \new_[19429]_ , \new_[19430]_ ,
    \new_[19431]_ , \new_[19432]_ , \new_[19433]_ , \new_[19434]_ ,
    \new_[19435]_ , \new_[19436]_ , \new_[19437]_ , \new_[19438]_ ,
    \new_[19439]_ , \new_[19440]_ , \new_[19441]_ , \new_[19442]_ ,
    \new_[19443]_ , \new_[19444]_ , \new_[19445]_ , \new_[19446]_ ,
    \new_[19447]_ , \new_[19448]_ , \new_[19449]_ , \new_[19450]_ ,
    \new_[19468]_ , \new_[19469]_ , \new_[19470]_ , \new_[19471]_ ,
    \new_[19472]_ , \new_[19473]_ , \new_[19474]_ , \new_[19475]_ ,
    \new_[19476]_ , \new_[19477]_ , \new_[19478]_ , \new_[19479]_ ,
    \new_[19480]_ , \new_[19481]_ , \new_[19482]_ , \new_[19483]_ ,
    \new_[19484]_ , \new_[19485]_ , \new_[19486]_ , \new_[19487]_ ,
    \new_[19488]_ , \new_[19489]_ , \new_[19490]_ , \new_[19491]_ ,
    \new_[19492]_ , \new_[19493]_ , \new_[19494]_ , \new_[19495]_ ,
    \new_[19496]_ , \new_[19497]_ , \new_[19498]_ , \new_[19499]_ ,
    \new_[19500]_ , \new_[19501]_ , \new_[19502]_ , \new_[19503]_ ,
    \new_[19504]_ , \new_[19505]_ , \new_[19506]_ , \new_[19507]_ ,
    \new_[19508]_ , \new_[19509]_ , \new_[19510]_ , \new_[19511]_ ,
    \new_[19512]_ , \new_[19513]_ , \new_[19514]_ , \new_[19515]_ ,
    \new_[19516]_ , \new_[19517]_ , \new_[19518]_ , \new_[19519]_ ,
    \new_[19520]_ , \new_[19521]_ , \new_[19522]_ , \new_[19523]_ ,
    \new_[19524]_ , \new_[19525]_ , \new_[19526]_ , \new_[19527]_ ,
    \new_[19528]_ , \new_[19529]_ , \new_[19530]_ , \new_[19531]_ ,
    \new_[19532]_ , \new_[19533]_ , \new_[19534]_ , \new_[19535]_ ,
    \new_[19536]_ , \new_[19537]_ , \new_[19538]_ , \new_[19539]_ ,
    \new_[19540]_ , \new_[19541]_ , \new_[19542]_ , \new_[19543]_ ,
    \new_[19544]_ , \new_[19545]_ , \new_[19546]_ , \new_[19547]_ ,
    \new_[19548]_ , \new_[19549]_ , \new_[19550]_ , \new_[19551]_ ,
    \new_[19552]_ , \new_[19553]_ , \new_[19554]_ , \new_[19555]_ ,
    \new_[19556]_ , \new_[19557]_ , \new_[19558]_ , \new_[19559]_ ,
    \new_[19560]_ , \new_[19561]_ , \new_[19562]_ , \new_[19563]_ ,
    \new_[19564]_ , \new_[19565]_ , \new_[19566]_ , \new_[19567]_ ,
    \new_[19568]_ , \new_[19569]_ , \new_[19570]_ , \new_[19571]_ ,
    \new_[19572]_ , \new_[19573]_ , \new_[19574]_ , \new_[19575]_ ,
    \new_[19576]_ , \new_[19577]_ , \new_[19578]_ , \new_[19579]_ ,
    \new_[19580]_ , \new_[19581]_ , \new_[19582]_ , \new_[19583]_ ,
    \new_[19584]_ , \new_[19585]_ , \new_[19586]_ , \new_[19587]_ ,
    \new_[19588]_ , \new_[19589]_ , \new_[19590]_ , \new_[19591]_ ,
    \new_[19592]_ , \new_[19593]_ , \new_[19594]_ , \new_[19595]_ ,
    \new_[19596]_ , \new_[19597]_ , \new_[19598]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19601]_ , \new_[19602]_ , \new_[19603]_ ,
    \new_[19604]_ , \new_[19605]_ , \new_[19606]_ , \new_[19607]_ ,
    \new_[19608]_ , \new_[19609]_ , \new_[19610]_ , \new_[19611]_ ,
    \new_[19612]_ , \new_[19613]_ , \new_[19614]_ , \new_[19615]_ ,
    \new_[19616]_ , \new_[19617]_ , \new_[19618]_ , \new_[19619]_ ,
    \new_[19620]_ , \new_[19621]_ , \new_[19622]_ , \new_[19623]_ ,
    \new_[19624]_ , \new_[19625]_ , \new_[19626]_ , \new_[19627]_ ,
    \new_[19628]_ , \new_[19629]_ , \new_[19630]_ , \new_[19631]_ ,
    \new_[19632]_ , \new_[19633]_ , \new_[19634]_ , \new_[19635]_ ,
    \new_[19636]_ , \new_[19637]_ , \new_[19638]_ , \new_[19639]_ ,
    \new_[19640]_ , \new_[19641]_ , \new_[19642]_ , \new_[19643]_ ,
    \new_[19644]_ , \new_[19645]_ , \new_[19646]_ , \new_[19647]_ ,
    \new_[19648]_ , \new_[19649]_ , \new_[19650]_ , \new_[19651]_ ,
    \new_[19652]_ , \new_[19653]_ , \new_[19654]_ , \new_[19655]_ ,
    \new_[19656]_ , \new_[19657]_ , \new_[19658]_ , \new_[19659]_ ,
    \new_[19660]_ , \new_[19661]_ , \new_[19662]_ , \new_[19663]_ ,
    \new_[19664]_ , \new_[19665]_ , \new_[19666]_ , \new_[19667]_ ,
    \new_[19668]_ , \new_[19669]_ , \new_[19670]_ , \new_[19671]_ ,
    \new_[19672]_ , \new_[19673]_ , \new_[19674]_ , \new_[19675]_ ,
    \new_[19676]_ , \new_[19677]_ , \new_[19678]_ , \new_[19679]_ ,
    \new_[19680]_ , \new_[19681]_ , \new_[19682]_ , \new_[19683]_ ,
    \new_[19684]_ , \new_[19685]_ , \new_[19686]_ , \new_[19687]_ ,
    \new_[19688]_ , \new_[19689]_ , \new_[19690]_ , \new_[19691]_ ,
    \new_[19692]_ , \new_[19693]_ , \new_[19694]_ , \new_[19695]_ ,
    \new_[19696]_ , \new_[19697]_ , \new_[19698]_ , \new_[19699]_ ,
    \new_[19700]_ , \new_[19701]_ , \new_[19702]_ , \new_[19703]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19706]_ , \new_[19707]_ ,
    \new_[19708]_ , \new_[19709]_ , \new_[19710]_ , \new_[19711]_ ,
    \new_[19712]_ , \new_[19713]_ , \new_[19714]_ , \new_[19715]_ ,
    \new_[19716]_ , \new_[19717]_ , \new_[19718]_ , \new_[19719]_ ,
    \new_[19720]_ , \new_[19721]_ , \new_[19722]_ , \new_[19723]_ ,
    \new_[19724]_ , \new_[19725]_ , \new_[19726]_ , \new_[19727]_ ,
    \new_[19728]_ , \new_[19729]_ , \new_[19730]_ , \new_[19731]_ ,
    \new_[19732]_ , \new_[19733]_ , \new_[19734]_ , \new_[19735]_ ,
    \new_[19736]_ , \new_[19737]_ , \new_[19738]_ , \new_[19739]_ ,
    \new_[19740]_ , \new_[19748]_ , \new_[19749]_ , \new_[19750]_ ,
    \new_[19751]_ , \new_[19752]_ , \new_[19753]_ , \new_[19754]_ ,
    \new_[19755]_ , \new_[19756]_ , \new_[19757]_ , \new_[19758]_ ,
    \new_[19759]_ , \new_[19760]_ , \new_[19761]_ , \new_[19762]_ ,
    \new_[19763]_ , \new_[19764]_ , \new_[19765]_ , \new_[19766]_ ,
    \new_[19767]_ , \new_[19768]_ , \new_[19769]_ , \new_[19770]_ ,
    \new_[19771]_ , \new_[19772]_ , \new_[19773]_ , \new_[19774]_ ,
    \new_[19775]_ , \new_[19776]_ , \new_[19777]_ , \new_[19778]_ ,
    \new_[19779]_ , \new_[19780]_ , \new_[19781]_ , \new_[19782]_ ,
    \new_[19783]_ , \new_[19784]_ , \new_[19785]_ , \new_[19786]_ ,
    \new_[19787]_ , \new_[19788]_ , \new_[19789]_ , \new_[19790]_ ,
    \new_[19791]_ , \new_[19792]_ , \new_[19793]_ , \new_[19794]_ ,
    \new_[19795]_ , \new_[19796]_ , \new_[19797]_ , \new_[19798]_ ,
    \new_[19799]_ , \new_[19800]_ , \new_[19801]_ , \new_[19802]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19805]_ , \new_[19806]_ ,
    \new_[19807]_ , \new_[19808]_ , \new_[19809]_ , \new_[19810]_ ,
    \new_[19811]_ , \new_[19812]_ , \new_[19813]_ , \new_[19814]_ ,
    \new_[19815]_ , \new_[19816]_ , \new_[19817]_ , \new_[19818]_ ,
    \new_[19819]_ , \new_[19820]_ , \new_[19821]_ , \new_[19822]_ ,
    \new_[19823]_ , \new_[19824]_ , \new_[19825]_ , \new_[19826]_ ,
    \new_[19827]_ , \new_[19828]_ , \new_[19829]_ , \new_[19830]_ ,
    \new_[19831]_ , \new_[19832]_ , \new_[19833]_ , \new_[19834]_ ,
    \new_[19835]_ , \new_[19836]_ , \new_[19837]_ , \new_[19838]_ ,
    \new_[19839]_ , \new_[19840]_ , \new_[19841]_ , \new_[19842]_ ,
    \new_[19843]_ , \new_[19844]_ , \new_[19845]_ , \new_[19846]_ ,
    \new_[19847]_ , \new_[19848]_ , \new_[19849]_ , \new_[19850]_ ,
    \new_[19851]_ , \new_[19852]_ , \new_[19853]_ , \new_[19854]_ ,
    \new_[19855]_ , \new_[19856]_ , \new_[19857]_ , \new_[19858]_ ,
    \new_[19859]_ , \new_[19860]_ , \new_[19861]_ , \new_[19862]_ ,
    \new_[19863]_ , \new_[19864]_ , \new_[19865]_ , \new_[19866]_ ,
    \new_[19867]_ , \new_[19868]_ , \new_[19869]_ , \new_[19870]_ ,
    \new_[19871]_ , \new_[19872]_ , \new_[19873]_ , \new_[19874]_ ,
    \new_[19875]_ , \new_[19876]_ , \new_[19877]_ , \new_[19878]_ ,
    \new_[19879]_ , \new_[19880]_ , \new_[19881]_ , \new_[19882]_ ,
    \new_[19883]_ , \new_[19884]_ , \new_[19885]_ , \new_[19886]_ ,
    \new_[19887]_ , \new_[19888]_ , \new_[19889]_ , \new_[19890]_ ,
    \new_[19891]_ , \new_[19892]_ , \new_[19893]_ , \new_[19894]_ ,
    \new_[19895]_ , \new_[19896]_ , \new_[19897]_ , \new_[19898]_ ,
    \new_[19899]_ , \new_[19900]_ , \new_[19901]_ , \new_[19902]_ ,
    \new_[19903]_ , \new_[19904]_ , \new_[19905]_ , \new_[19906]_ ,
    \new_[19907]_ , \new_[19908]_ , \new_[19909]_ , \new_[19910]_ ,
    \new_[19911]_ , \new_[19912]_ , \new_[19913]_ , \new_[19914]_ ,
    \new_[19915]_ , \new_[19916]_ , \new_[19917]_ , \new_[19918]_ ,
    \new_[19919]_ , \new_[19920]_ , \new_[19921]_ , \new_[19922]_ ,
    \new_[19923]_ , \new_[19924]_ , \new_[19925]_ , \new_[19926]_ ,
    \new_[19927]_ , \new_[19928]_ , \new_[19929]_ , \new_[19930]_ ,
    \new_[19931]_ , \new_[19932]_ , \new_[19933]_ , \new_[19934]_ ,
    \new_[19935]_ , \new_[19936]_ , \new_[19937]_ , \new_[19938]_ ,
    \new_[19939]_ , \new_[19940]_ , \new_[19941]_ , \new_[19942]_ ,
    \new_[19943]_ , \new_[19944]_ , \new_[19945]_ , \new_[19946]_ ,
    \new_[19947]_ , \new_[19948]_ , \new_[19949]_ , \new_[19950]_ ,
    \new_[19951]_ , \new_[19952]_ , \new_[19953]_ , \new_[19954]_ ,
    \new_[19955]_ , \new_[19956]_ , \new_[19957]_ , \new_[19958]_ ,
    \new_[19959]_ , \new_[19960]_ , \new_[19961]_ , \new_[19962]_ ,
    \new_[19963]_ , \new_[19964]_ , \new_[19965]_ , \new_[19966]_ ,
    \new_[19967]_ , \new_[19968]_ , \new_[19969]_ , \new_[19970]_ ,
    \new_[19971]_ , \new_[19972]_ , \new_[19973]_ , \new_[19974]_ ,
    \new_[19975]_ , \new_[19976]_ , \new_[19977]_ , \new_[19978]_ ,
    \new_[19979]_ , \new_[19980]_ , \new_[19981]_ , \new_[19982]_ ,
    \new_[19983]_ , \new_[19984]_ , \new_[19985]_ , \new_[19986]_ ,
    \new_[19987]_ , \new_[19988]_ , \new_[19989]_ , \new_[19990]_ ,
    \new_[19991]_ , \new_[19992]_ , \new_[19993]_ , \new_[19994]_ ,
    \new_[19995]_ , \new_[19996]_ , \new_[19997]_ , \new_[19998]_ ,
    \new_[19999]_ , \new_[20000]_ , \new_[20001]_ , \new_[20002]_ ,
    \new_[20003]_ , \new_[20004]_ , \new_[20005]_ , \new_[20006]_ ,
    \new_[20007]_ , \new_[20008]_ , \new_[20009]_ , \new_[20010]_ ,
    \new_[20011]_ , \new_[20012]_ , \new_[20013]_ , \new_[20014]_ ,
    \new_[20015]_ , \new_[20016]_ , \new_[20017]_ , \new_[20018]_ ,
    \new_[20019]_ , \new_[20020]_ , \new_[20021]_ , \new_[20022]_ ,
    \new_[20023]_ , \new_[20024]_ , \new_[20025]_ , \new_[20026]_ ,
    \new_[20027]_ , \new_[20028]_ , \new_[20029]_ , \new_[20030]_ ,
    \new_[20031]_ , \new_[20032]_ , \new_[20033]_ , \new_[20034]_ ,
    \new_[20035]_ , \new_[20036]_ , \new_[20037]_ , \new_[20038]_ ,
    \new_[20039]_ , \new_[20040]_ , \new_[20041]_ , \new_[20042]_ ,
    \new_[20043]_ , \new_[20044]_ , \new_[20045]_ , \new_[20046]_ ,
    \new_[20047]_ , \new_[20048]_ , \new_[20049]_ , \new_[20050]_ ,
    \new_[20051]_ , \new_[20052]_ , \new_[20053]_ , \new_[20054]_ ,
    \new_[20055]_ , \new_[20056]_ , \new_[20057]_ , \new_[20058]_ ,
    \new_[20059]_ , \new_[20060]_ , \new_[20061]_ , \new_[20062]_ ,
    \new_[20063]_ , \new_[20064]_ , \new_[20065]_ , \new_[20066]_ ,
    \new_[20067]_ , \new_[20068]_ , \new_[20069]_ , \new_[20070]_ ,
    \new_[20071]_ , \new_[20072]_ , \new_[20073]_ , \new_[20074]_ ,
    \new_[20075]_ , \new_[20076]_ , \new_[20077]_ , \new_[20078]_ ,
    \new_[20079]_ , \new_[20080]_ , \new_[20081]_ , \new_[20082]_ ,
    \new_[20083]_ , \new_[20084]_ , \new_[20085]_ , \new_[20086]_ ,
    \new_[20087]_ , \new_[20088]_ , \new_[20089]_ , \new_[20090]_ ,
    \new_[20091]_ , \new_[20092]_ , \new_[20093]_ , \new_[20094]_ ,
    \new_[20095]_ , \new_[20096]_ , \new_[20097]_ , \new_[20098]_ ,
    \new_[20099]_ , \new_[20100]_ , \new_[20101]_ , \new_[20102]_ ,
    \new_[20103]_ , \new_[20104]_ , \new_[20105]_ , \new_[20106]_ ,
    \new_[20107]_ , \new_[20108]_ , \new_[20109]_ , \new_[20110]_ ,
    \new_[20111]_ , \new_[20112]_ , \new_[20113]_ , \new_[20114]_ ,
    \new_[20115]_ , \new_[20116]_ , \new_[20117]_ , \new_[20118]_ ,
    \new_[20119]_ , \new_[20120]_ , \new_[20121]_ , \new_[20122]_ ,
    \new_[20123]_ , \new_[20124]_ , \new_[20125]_ , \new_[20126]_ ,
    \new_[20127]_ , \new_[20128]_ , \new_[20129]_ , \new_[20130]_ ,
    \new_[20131]_ , \new_[20132]_ , \new_[20133]_ , \new_[20134]_ ,
    \new_[20135]_ , \new_[20136]_ , \new_[20137]_ , \new_[20138]_ ,
    \new_[20139]_ , \new_[20140]_ , \new_[20141]_ , \new_[20142]_ ,
    \new_[20143]_ , \new_[20144]_ , \new_[20145]_ , \new_[20146]_ ,
    \new_[20147]_ , \new_[20148]_ , \new_[20149]_ , \new_[20150]_ ,
    \new_[20151]_ , \new_[20152]_ , \new_[20153]_ , \new_[20154]_ ,
    \new_[20155]_ , \new_[20156]_ , \new_[20157]_ , \new_[20158]_ ,
    \new_[20159]_ , \new_[20160]_ , \new_[20161]_ , \new_[20162]_ ,
    \new_[20163]_ , \new_[20164]_ , \new_[20165]_ , \new_[20166]_ ,
    \new_[20167]_ , \new_[20168]_ , \new_[20169]_ , \new_[20170]_ ,
    \new_[20171]_ , \new_[20172]_ , \new_[20173]_ , \new_[20174]_ ,
    \new_[20175]_ , \new_[20176]_ , \new_[20178]_ , \new_[20179]_ ,
    \new_[20180]_ , \new_[20181]_ , \new_[20182]_ , \new_[20183]_ ,
    \new_[20185]_ , \new_[20191]_ , \new_[20199]_ , \new_[20200]_ ,
    \new_[20201]_ , \new_[20202]_ , \new_[20203]_ , \new_[20204]_ ,
    \new_[20205]_ , \new_[20207]_ , \new_[20208]_ , \new_[20209]_ ,
    \new_[20210]_ , \new_[20211]_ , \new_[20212]_ , \new_[20213]_ ,
    \new_[20214]_ , \new_[20215]_ , \new_[20216]_ , \new_[20217]_ ,
    \new_[20218]_ , \new_[20219]_ , \new_[20220]_ , \new_[20221]_ ,
    \new_[20222]_ , \new_[20223]_ , \new_[20224]_ , \new_[20226]_ ,
    \new_[20227]_ , \new_[20228]_ , \new_[20229]_ , \new_[20230]_ ,
    \new_[20231]_ , \new_[20232]_ , \new_[20233]_ , \new_[20234]_ ,
    \new_[20235]_ , \new_[20236]_ , \new_[20237]_ , \new_[20238]_ ,
    \new_[20239]_ , \new_[20240]_ , \new_[20241]_ , \new_[20242]_ ,
    \new_[20243]_ , \new_[20244]_ , \new_[20245]_ , \new_[20246]_ ,
    \new_[20247]_ , \new_[20248]_ , \new_[20249]_ , \new_[20250]_ ,
    \new_[20251]_ , \new_[20252]_ , \new_[20253]_ , \new_[20254]_ ,
    \new_[20255]_ , \new_[20256]_ , \new_[20257]_ , \new_[20258]_ ,
    \new_[20259]_ , \new_[20260]_ , \new_[20262]_ , \new_[20263]_ ,
    \new_[20265]_ , \new_[20266]_ , \new_[20267]_ , \new_[20268]_ ,
    \new_[20269]_ , \new_[20270]_ , \new_[20271]_ , \new_[20272]_ ,
    \new_[20273]_ , \new_[20274]_ , \new_[20275]_ , \new_[20276]_ ,
    \new_[20277]_ , \new_[20278]_ , \new_[20279]_ , \new_[20280]_ ,
    \new_[20281]_ , \new_[20282]_ , \new_[20285]_ , \new_[20286]_ ,
    \new_[20287]_ , \new_[20288]_ , \new_[20289]_ , \new_[20294]_ ,
    \new_[20295]_ , \new_[20296]_ , \new_[20297]_ , \new_[20298]_ ,
    \new_[20301]_ , \new_[20302]_ , \new_[20303]_ , \new_[20304]_ ,
    \new_[20306]_ , \new_[20309]_ , \new_[20310]_ , \new_[20311]_ ,
    \new_[20312]_ , \new_[20314]_ , \new_[20316]_ , \new_[20317]_ ,
    \new_[20319]_ , \new_[20323]_ , \new_[20324]_ , \new_[20325]_ ,
    \new_[20326]_ , \new_[20327]_ , \new_[20328]_ , \new_[20329]_ ,
    \new_[20330]_ , \new_[20331]_ , \new_[20332]_ , \new_[20333]_ ,
    \new_[20334]_ , \new_[20335]_ , \new_[20336]_ , \new_[20337]_ ,
    \new_[20338]_ , \new_[20339]_ , \new_[20340]_ , \new_[20341]_ ,
    \new_[20342]_ , \new_[20343]_ , \new_[20344]_ , \new_[20345]_ ,
    \new_[20346]_ , \new_[20347]_ , \new_[20348]_ , \new_[20349]_ ,
    \new_[20350]_ , \new_[20351]_ , \new_[20352]_ , \new_[20353]_ ,
    \new_[20354]_ , \new_[20355]_ , \new_[20356]_ , \new_[20357]_ ,
    \new_[20358]_ , \new_[20359]_ , \new_[20360]_ , \new_[20361]_ ,
    \new_[20362]_ , \new_[20363]_ , \new_[20364]_ , \new_[20365]_ ,
    \new_[20366]_ , \new_[20367]_ , \new_[20368]_ , \new_[20369]_ ,
    \new_[20370]_ , \new_[20371]_ , \new_[20372]_ , \new_[20373]_ ,
    \new_[20374]_ , \new_[20375]_ , \new_[20376]_ , \new_[20377]_ ,
    \new_[20378]_ , \new_[20379]_ , \new_[20380]_ , \new_[20381]_ ,
    \new_[20382]_ , \new_[20383]_ , \new_[20384]_ , \new_[20385]_ ,
    \new_[20386]_ , \new_[20387]_ , \new_[20388]_ , \new_[20389]_ ,
    \new_[20390]_ , \new_[20391]_ , \new_[20392]_ , \new_[20393]_ ,
    \new_[20394]_ , \new_[20395]_ , \new_[20396]_ , \new_[20397]_ ,
    \new_[20398]_ , \new_[20399]_ , \new_[20400]_ , \new_[20401]_ ,
    \new_[20402]_ , \new_[20403]_ , \new_[20404]_ , \new_[20405]_ ,
    \new_[20406]_ , \new_[20407]_ , \new_[20408]_ , \new_[20409]_ ,
    \new_[20410]_ , \new_[20411]_ , \new_[20412]_ , \new_[20413]_ ,
    \new_[20414]_ , \new_[20415]_ , \new_[20416]_ , \new_[20417]_ ,
    \new_[20418]_ , \new_[20419]_ , \new_[20420]_ , \new_[20421]_ ,
    \new_[20422]_ , \new_[20423]_ , \new_[20424]_ , \new_[20425]_ ,
    \new_[20426]_ , \new_[20427]_ , \new_[20428]_ , \new_[20429]_ ,
    \new_[20430]_ , \new_[20431]_ , \new_[20432]_ , \new_[20433]_ ,
    \new_[20434]_ , \new_[20435]_ , \new_[20436]_ , \new_[20437]_ ,
    \new_[20438]_ , \new_[20439]_ , \new_[20440]_ , \new_[20441]_ ,
    \new_[20442]_ , \new_[20443]_ , \new_[20444]_ , \new_[20445]_ ,
    \new_[20446]_ , \new_[20447]_ , \new_[20448]_ , \new_[20449]_ ,
    \new_[20450]_ , \new_[20451]_ , \new_[20452]_ , \new_[20453]_ ,
    \new_[20454]_ , \new_[20455]_ , \new_[20456]_ , \new_[20457]_ ,
    \new_[20458]_ , \new_[20459]_ , \new_[20460]_ , \new_[20461]_ ,
    \new_[20462]_ , \new_[20463]_ , \new_[20464]_ , \new_[20465]_ ,
    \new_[20466]_ , \new_[20467]_ , \new_[20468]_ , \new_[20469]_ ,
    \new_[20470]_ , \new_[20471]_ , \new_[20472]_ , \new_[20473]_ ,
    \new_[20474]_ , \new_[20475]_ , \new_[20476]_ , \new_[20477]_ ,
    \new_[20478]_ , \new_[20479]_ , \new_[20480]_ , \new_[20481]_ ,
    \new_[20482]_ , \new_[20483]_ , \new_[20484]_ , \new_[20485]_ ,
    \new_[20486]_ , \new_[20487]_ , \new_[20488]_ , \new_[20489]_ ,
    \new_[20490]_ , \new_[20491]_ , \new_[20492]_ , \new_[20493]_ ,
    \new_[20494]_ , \new_[20495]_ , \new_[20496]_ , \new_[20497]_ ,
    \new_[20498]_ , \new_[20499]_ , \new_[20500]_ , \new_[20501]_ ,
    \new_[20502]_ , \new_[20503]_ , \new_[20504]_ , \new_[20505]_ ,
    \new_[20506]_ , \new_[20507]_ , \new_[20508]_ , \new_[20509]_ ,
    \new_[20510]_ , \new_[20511]_ , \new_[20512]_ , \new_[20520]_ ,
    \new_[20521]_ , \new_[20522]_ , \new_[20523]_ , \new_[20524]_ ,
    \new_[20525]_ , \new_[20526]_ , \new_[20527]_ , \new_[20528]_ ,
    \new_[20529]_ , \new_[20530]_ , \new_[20531]_ , \new_[20532]_ ,
    \new_[20533]_ , \new_[20534]_ , \new_[20535]_ , \new_[20536]_ ,
    \new_[20537]_ , \new_[20538]_ , \new_[20539]_ , \new_[20540]_ ,
    \new_[20541]_ , \new_[20542]_ , \new_[20543]_ , \new_[20544]_ ,
    \new_[20545]_ , \new_[20546]_ , \new_[20547]_ , \new_[20548]_ ,
    \new_[20549]_ , \new_[20550]_ , \new_[20551]_ , \new_[20552]_ ,
    \new_[20553]_ , \new_[20554]_ , \new_[20555]_ , \new_[20556]_ ,
    \new_[20557]_ , \new_[20558]_ , \new_[20559]_ , \new_[20560]_ ,
    \new_[20561]_ , \new_[20562]_ , \new_[20563]_ , \new_[20564]_ ,
    \new_[20565]_ , \new_[20566]_ , \new_[20567]_ , \new_[20568]_ ,
    \new_[20569]_ , \new_[20570]_ , \new_[20571]_ , \new_[20572]_ ,
    \new_[20573]_ , \new_[20574]_ , \new_[20575]_ , \new_[20576]_ ,
    \new_[20577]_ , \new_[20578]_ , \new_[20579]_ , \new_[20580]_ ,
    \new_[20581]_ , \new_[20582]_ , \new_[20583]_ , \new_[20584]_ ,
    \new_[20585]_ , \new_[20586]_ , \new_[20587]_ , \new_[20588]_ ,
    \new_[20589]_ , \new_[20590]_ , \new_[20591]_ , \new_[20592]_ ,
    \new_[20593]_ , \new_[20594]_ , \new_[20595]_ , \new_[20596]_ ,
    \new_[20597]_ , \new_[20598]_ , \new_[20599]_ , \new_[20600]_ ,
    \new_[20601]_ , \new_[20602]_ , \new_[20603]_ , \new_[20604]_ ,
    \new_[20605]_ , \new_[20606]_ , \new_[20607]_ , \new_[20608]_ ,
    \new_[20609]_ , \new_[20610]_ , \new_[20611]_ , \new_[20612]_ ,
    \new_[20613]_ , \new_[20614]_ , \new_[20615]_ , \new_[20616]_ ,
    \new_[20617]_ , \new_[20618]_ , \new_[20619]_ , \new_[20620]_ ,
    \new_[20621]_ , \new_[20622]_ , \new_[20623]_ , \new_[20624]_ ,
    \new_[20625]_ , \new_[20626]_ , \new_[20627]_ , \new_[20628]_ ,
    \new_[20629]_ , \new_[20631]_ , \new_[20632]_ , \new_[20633]_ ,
    \new_[20634]_ , \new_[20635]_ , \new_[20636]_ , \new_[20637]_ ,
    \new_[20638]_ , \new_[20639]_ , \new_[20640]_ , \new_[20641]_ ,
    \new_[20642]_ , \new_[20643]_ , \new_[20644]_ , \new_[20645]_ ,
    \new_[20646]_ , \new_[20647]_ , \new_[20648]_ , \new_[20649]_ ,
    \new_[20650]_ , \new_[20651]_ , \new_[20652]_ , \new_[20653]_ ,
    \new_[20654]_ , \new_[20655]_ , \new_[20656]_ , \new_[20657]_ ,
    \new_[20658]_ , \new_[20659]_ , \new_[20660]_ , \new_[20661]_ ,
    \new_[20662]_ , \new_[20663]_ , \new_[20664]_ , \new_[20665]_ ,
    \new_[20666]_ , \new_[20667]_ , \new_[20668]_ , \new_[20669]_ ,
    \new_[20670]_ , \new_[20671]_ , \new_[20672]_ , \new_[20673]_ ,
    \new_[20674]_ , \new_[20675]_ , \new_[20676]_ , \new_[20677]_ ,
    \new_[20678]_ , \new_[20679]_ , \new_[20680]_ , \new_[20681]_ ,
    \new_[20682]_ , \new_[20683]_ , \new_[20684]_ , \new_[20685]_ ,
    \new_[20686]_ , \new_[20687]_ , \new_[20688]_ , \new_[20689]_ ,
    \new_[20690]_ , \new_[20691]_ , \new_[20692]_ , \new_[20693]_ ,
    \new_[20694]_ , \new_[20695]_ , \new_[20696]_ , \new_[20697]_ ,
    \new_[20698]_ , \new_[20699]_ , \new_[20700]_ , \new_[20701]_ ,
    \new_[20702]_ , \new_[20703]_ , \new_[20704]_ , \new_[20705]_ ,
    \new_[20706]_ , \new_[20707]_ , \new_[20708]_ , \new_[20709]_ ,
    \new_[20710]_ , \new_[20711]_ , \new_[20712]_ , \new_[20713]_ ,
    \new_[20714]_ , \new_[20715]_ , \new_[20716]_ , \new_[20717]_ ,
    \new_[20718]_ , \new_[20719]_ , \new_[20720]_ , \new_[20721]_ ,
    \new_[20722]_ , \new_[20723]_ , \new_[20724]_ , \new_[20725]_ ,
    \new_[20726]_ , \new_[20727]_ , \new_[20728]_ , \new_[20729]_ ,
    \new_[20730]_ , \new_[20731]_ , \new_[20732]_ , \new_[20733]_ ,
    \new_[20734]_ , \new_[20735]_ , \new_[20736]_ , \new_[20737]_ ,
    \new_[20738]_ , \new_[20739]_ , \new_[20740]_ , \new_[20741]_ ,
    \new_[20742]_ , \new_[20743]_ , \new_[20744]_ , \new_[20745]_ ,
    \new_[20746]_ , \new_[20747]_ , \new_[20748]_ , \new_[20749]_ ,
    \new_[20750]_ , \new_[20751]_ , \new_[20752]_ , \new_[20753]_ ,
    \new_[20754]_ , \new_[20755]_ , \new_[20756]_ , \new_[20757]_ ,
    \new_[20758]_ , \new_[20759]_ , \new_[20760]_ , \new_[20761]_ ,
    \new_[20762]_ , \new_[20763]_ , \new_[20764]_ , \new_[20765]_ ,
    \new_[20766]_ , \new_[20767]_ , \new_[20768]_ , \new_[20769]_ ,
    \new_[20770]_ , \new_[20771]_ , \new_[20772]_ , \new_[20773]_ ,
    \new_[20774]_ , \new_[20775]_ , \new_[20776]_ , \new_[20777]_ ,
    \new_[20778]_ , \new_[20779]_ , \new_[20780]_ , \new_[20781]_ ,
    \new_[20782]_ , \new_[20783]_ , \new_[20784]_ , \new_[20785]_ ,
    \new_[20786]_ , \new_[20787]_ , \new_[20788]_ , \new_[20789]_ ,
    \new_[20790]_ , \new_[20791]_ , \new_[20792]_ , \new_[20793]_ ,
    \new_[20794]_ , \new_[20795]_ , \new_[20796]_ , \new_[20797]_ ,
    \new_[20798]_ , \new_[20799]_ , \new_[20800]_ , \new_[20801]_ ,
    \new_[20802]_ , \new_[20803]_ , \new_[20804]_ , \new_[20805]_ ,
    \new_[20806]_ , \new_[20807]_ , \new_[20808]_ , \new_[20809]_ ,
    \new_[20810]_ , \new_[20811]_ , \new_[20812]_ , \new_[20813]_ ,
    \new_[20814]_ , \new_[20815]_ , \new_[20816]_ , \new_[20817]_ ,
    \new_[20818]_ , \new_[20819]_ , \new_[20820]_ , \new_[20821]_ ,
    \new_[20822]_ , \new_[20823]_ , \new_[20824]_ , \new_[20825]_ ,
    \new_[20826]_ , \new_[20827]_ , \new_[20828]_ , \new_[20829]_ ,
    \new_[20830]_ , \new_[20831]_ , \new_[20832]_ , \new_[20833]_ ,
    \new_[20834]_ , \new_[20835]_ , \new_[20836]_ , \new_[20837]_ ,
    \new_[20838]_ , \new_[20839]_ , \new_[20840]_ , \new_[20841]_ ,
    \new_[20842]_ , \new_[20843]_ , \new_[20844]_ , \new_[20845]_ ,
    \new_[20846]_ , \new_[20847]_ , \new_[20848]_ , \new_[20849]_ ,
    \new_[20850]_ , \new_[20851]_ , \new_[20852]_ , \new_[20853]_ ,
    \new_[20854]_ , \new_[20855]_ , \new_[20856]_ , \new_[20857]_ ,
    \new_[20858]_ , \new_[20859]_ , \new_[20860]_ , \new_[20861]_ ,
    \new_[20862]_ , \new_[20863]_ , \new_[20864]_ , \new_[20865]_ ,
    \new_[20866]_ , \new_[20867]_ , \new_[20868]_ , \new_[20869]_ ,
    \new_[20870]_ , \new_[20871]_ , \new_[20872]_ , \new_[20873]_ ,
    \new_[20874]_ , \new_[20875]_ , \new_[20876]_ , \new_[20877]_ ,
    \new_[20878]_ , \new_[20879]_ , \new_[20880]_ , \new_[20881]_ ,
    \new_[20882]_ , \new_[20883]_ , \new_[20884]_ , \new_[20885]_ ,
    \new_[20886]_ , \new_[20887]_ , \new_[20888]_ , \new_[20889]_ ,
    \new_[20890]_ , \new_[20891]_ , \new_[20892]_ , \new_[20893]_ ,
    \new_[20894]_ , \new_[20895]_ , \new_[20896]_ , \new_[20897]_ ,
    \new_[20898]_ , \new_[20899]_ , \new_[20900]_ , \new_[20901]_ ,
    \new_[20902]_ , \new_[20903]_ , \new_[20904]_ , \new_[20905]_ ,
    \new_[20906]_ , \new_[20907]_ , \new_[20908]_ , \new_[20909]_ ,
    \new_[20910]_ , \new_[20911]_ , \new_[20912]_ , \new_[20913]_ ,
    \new_[20914]_ , \new_[20915]_ , \new_[20916]_ , \new_[20917]_ ,
    \new_[20918]_ , \new_[20919]_ , \new_[20920]_ , \new_[20921]_ ,
    \new_[20922]_ , \new_[20923]_ , \new_[20924]_ , \new_[20925]_ ,
    \new_[20926]_ , \new_[20927]_ , \new_[20928]_ , \new_[20929]_ ,
    \new_[20930]_ , \new_[20931]_ , \new_[20932]_ , \new_[20933]_ ,
    \new_[20934]_ , \new_[20935]_ , \new_[20936]_ , \new_[20937]_ ,
    \new_[20938]_ , \new_[20939]_ , \new_[20940]_ , \new_[20941]_ ,
    \new_[20942]_ , \new_[20943]_ , \new_[20944]_ , \new_[20945]_ ,
    \new_[20946]_ , \new_[20947]_ , \new_[20948]_ , \new_[20949]_ ,
    \new_[20950]_ , \new_[20951]_ , \new_[20952]_ , \new_[20953]_ ,
    \new_[20954]_ , \new_[20955]_ , \new_[20956]_ , \new_[20957]_ ,
    \new_[20958]_ , \new_[20959]_ , \new_[20960]_ , \new_[20961]_ ,
    \new_[20962]_ , \new_[20963]_ , \new_[20964]_ , \new_[20965]_ ,
    \new_[20966]_ , \new_[20967]_ , \new_[20968]_ , \new_[20969]_ ,
    \new_[20970]_ , \new_[20971]_ , \new_[20972]_ , \new_[20973]_ ,
    \new_[20974]_ , \new_[20975]_ , \new_[20976]_ , \new_[20977]_ ,
    \new_[20978]_ , \new_[20979]_ , \new_[20980]_ , \new_[20981]_ ,
    \new_[20982]_ , \new_[20983]_ , \new_[20984]_ , \new_[20985]_ ,
    \new_[20986]_ , \new_[20987]_ , \new_[20988]_ , \new_[20989]_ ,
    \new_[20990]_ , \new_[20991]_ , \new_[20992]_ , \new_[20993]_ ,
    \new_[20994]_ , \new_[20995]_ , \new_[20996]_ , \new_[20997]_ ,
    \new_[20998]_ , \new_[20999]_ , \new_[21000]_ , \new_[21001]_ ,
    \new_[21002]_ , \new_[21003]_ , \new_[21004]_ , \new_[21005]_ ,
    \new_[21006]_ , \new_[21007]_ , \new_[21008]_ , \new_[21009]_ ,
    \new_[21010]_ , \new_[21011]_ , \new_[21012]_ , \new_[21013]_ ,
    \new_[21014]_ , \new_[21015]_ , \new_[21017]_ , \new_[21018]_ ,
    \new_[21019]_ , \new_[21020]_ , \new_[21021]_ , \new_[21022]_ ,
    \new_[21023]_ , \new_[21028]_ , \new_[21030]_ , \new_[21031]_ ,
    \new_[21035]_ , \new_[21038]_ , \new_[21044]_ , \new_[21046]_ ,
    \new_[21048]_ , \new_[21049]_ , \new_[21053]_ , \new_[21054]_ ,
    \new_[21055]_ , \new_[21056]_ , \new_[21057]_ , \new_[21059]_ ,
    \new_[21060]_ , \new_[21061]_ , \new_[21062]_ , \new_[21063]_ ,
    \new_[21064]_ , \new_[21067]_ , \new_[21068]_ , \new_[21069]_ ,
    \new_[21070]_ , \new_[21071]_ , \new_[21072]_ , \new_[21073]_ ,
    \new_[21075]_ , \new_[21076]_ , \new_[21077]_ , \new_[21078]_ ,
    \new_[21080]_ , \new_[21081]_ , \new_[21082]_ , \new_[21083]_ ,
    \new_[21084]_ , \new_[21085]_ , \new_[21086]_ , \new_[21087]_ ,
    \new_[21088]_ , \new_[21090]_ , \new_[21091]_ , \new_[21092]_ ,
    \new_[21093]_ , \new_[21094]_ , \new_[21095]_ , \new_[21097]_ ,
    \new_[21098]_ , \new_[21099]_ , \new_[21100]_ , \new_[21101]_ ,
    \new_[21102]_ , \new_[21103]_ , \new_[21104]_ , \new_[21105]_ ,
    \new_[21106]_ , \new_[21107]_ , \new_[21108]_ , \new_[21109]_ ,
    \new_[21110]_ , \new_[21111]_ , \new_[21112]_ , \new_[21113]_ ,
    \new_[21114]_ , \new_[21115]_ , \new_[21118]_ , \new_[21119]_ ,
    \new_[21121]_ , \new_[21122]_ , \new_[21124]_ , \new_[21126]_ ,
    \new_[21128]_ , \new_[21129]_ , \new_[21130]_ , \new_[21131]_ ,
    \new_[21134]_ , \new_[21136]_ , \new_[21137]_ , \new_[21138]_ ,
    \new_[21139]_ , \new_[21140]_ , \new_[21142]_ , \new_[21145]_ ,
    \new_[21148]_ , \new_[21149]_ , \new_[21150]_ , \new_[21152]_ ,
    \new_[21153]_ , \new_[21154]_ , \new_[21155]_ , \new_[21157]_ ,
    \new_[21158]_ , \new_[21159]_ , \new_[21160]_ , \new_[21162]_ ,
    \new_[21163]_ , \new_[21164]_ , \new_[21166]_ , \new_[21168]_ ,
    \new_[21169]_ , \new_[21170]_ , \new_[21171]_ , \new_[21172]_ ,
    \new_[21173]_ , \new_[21174]_ , \new_[21176]_ , \new_[21177]_ ,
    \new_[21178]_ , \new_[21179]_ , \new_[21180]_ , \new_[21181]_ ,
    \new_[21182]_ , \new_[21183]_ , \new_[21184]_ , \new_[21185]_ ,
    \new_[21186]_ , \new_[21187]_ , \new_[21188]_ , \new_[21189]_ ,
    \new_[21190]_ , \new_[21191]_ , \new_[21192]_ , \new_[21193]_ ,
    \new_[21194]_ , \new_[21195]_ , \new_[21196]_ , \new_[21197]_ ,
    \new_[21198]_ , \new_[21199]_ , \new_[21200]_ , \new_[21201]_ ,
    \new_[21202]_ , \new_[21203]_ , \new_[21204]_ , \new_[21205]_ ,
    \new_[21206]_ , \new_[21207]_ , \new_[21208]_ , \new_[21209]_ ,
    \new_[21210]_ , \new_[21211]_ , \new_[21212]_ , \new_[21213]_ ,
    \new_[21214]_ , \new_[21215]_ , \new_[21216]_ , \new_[21217]_ ,
    \new_[21218]_ , \new_[21219]_ , \new_[21220]_ , \new_[21221]_ ,
    \new_[21222]_ , \new_[21223]_ , \new_[21224]_ , \new_[21225]_ ,
    \new_[21226]_ , \new_[21227]_ , \new_[21228]_ , \new_[21229]_ ,
    \new_[21230]_ , \new_[21231]_ , \new_[21232]_ , \new_[21233]_ ,
    \new_[21234]_ , \new_[21235]_ , \new_[21236]_ , \new_[21237]_ ,
    \new_[21238]_ , \new_[21239]_ , \new_[21240]_ , \new_[21241]_ ,
    \new_[21242]_ , \new_[21243]_ , \new_[21244]_ , \new_[21245]_ ,
    \new_[21246]_ , \new_[21247]_ , \new_[21248]_ , \new_[21249]_ ,
    \new_[21250]_ , \new_[21251]_ , \new_[21252]_ , \new_[21253]_ ,
    \new_[21254]_ , \new_[21255]_ , \new_[21256]_ , \new_[21257]_ ,
    \new_[21258]_ , \new_[21259]_ , \new_[21260]_ , \new_[21261]_ ,
    \new_[21262]_ , \new_[21263]_ , \new_[21264]_ , \new_[21265]_ ,
    \new_[21266]_ , \new_[21267]_ , \new_[21268]_ , \new_[21269]_ ,
    \new_[21270]_ , \new_[21271]_ , \new_[21272]_ , \new_[21273]_ ,
    \new_[21274]_ , \new_[21275]_ , \new_[21276]_ , \new_[21277]_ ,
    \new_[21278]_ , \new_[21279]_ , \new_[21280]_ , \new_[21281]_ ,
    \new_[21282]_ , \new_[21283]_ , \new_[21284]_ , \new_[21285]_ ,
    \new_[21286]_ , \new_[21287]_ , \new_[21288]_ , \new_[21289]_ ,
    \new_[21290]_ , \new_[21291]_ , \new_[21292]_ , \new_[21293]_ ,
    \new_[21294]_ , \new_[21295]_ , \new_[21296]_ , \new_[21297]_ ,
    \new_[21298]_ , \new_[21299]_ , \new_[21300]_ , \new_[21301]_ ,
    \new_[21302]_ , \new_[21303]_ , \new_[21304]_ , \new_[21305]_ ,
    \new_[21306]_ , \new_[21307]_ , \new_[21308]_ , \new_[21309]_ ,
    \new_[21310]_ , \new_[21311]_ , \new_[21312]_ , \new_[21313]_ ,
    \new_[21314]_ , \new_[21315]_ , \new_[21316]_ , \new_[21317]_ ,
    \new_[21318]_ , \new_[21319]_ , \new_[21320]_ , \new_[21321]_ ,
    \new_[21322]_ , \new_[21323]_ , \new_[21324]_ , \new_[21325]_ ,
    \new_[21326]_ , \new_[21327]_ , \new_[21328]_ , \new_[21329]_ ,
    \new_[21330]_ , \new_[21331]_ , \new_[21332]_ , \new_[21333]_ ,
    \new_[21334]_ , \new_[21335]_ , \new_[21336]_ , \new_[21337]_ ,
    \new_[21338]_ , \new_[21339]_ , \new_[21340]_ , \new_[21341]_ ,
    \new_[21342]_ , \new_[21343]_ , \new_[21344]_ , \new_[21345]_ ,
    \new_[21346]_ , \new_[21347]_ , \new_[21348]_ , \new_[21349]_ ,
    \new_[21350]_ , \new_[21351]_ , \new_[21352]_ , \new_[21353]_ ,
    \new_[21354]_ , \new_[21355]_ , \new_[21356]_ , \new_[21357]_ ,
    \new_[21358]_ , \new_[21359]_ , \new_[21360]_ , \new_[21361]_ ,
    \new_[21362]_ , \new_[21363]_ , \new_[21364]_ , \new_[21365]_ ,
    \new_[21366]_ , \new_[21367]_ , \new_[21368]_ , \new_[21369]_ ,
    \new_[21370]_ , \new_[21371]_ , \new_[21372]_ , \new_[21373]_ ,
    \new_[21374]_ , \new_[21375]_ , \new_[21376]_ , \new_[21377]_ ,
    \new_[21378]_ , \new_[21379]_ , \new_[21380]_ , \new_[21381]_ ,
    \new_[21382]_ , \new_[21383]_ , \new_[21384]_ , \new_[21385]_ ,
    \new_[21386]_ , \new_[21387]_ , \new_[21388]_ , \new_[21389]_ ,
    \new_[21390]_ , \new_[21391]_ , \new_[21392]_ , \new_[21393]_ ,
    \new_[21394]_ , \new_[21395]_ , \new_[21396]_ , \new_[21397]_ ,
    \new_[21398]_ , \new_[21399]_ , \new_[21400]_ , \new_[21401]_ ,
    \new_[21402]_ , \new_[21403]_ , \new_[21404]_ , \new_[21405]_ ,
    \new_[21406]_ , \new_[21407]_ , \new_[21408]_ , \new_[21409]_ ,
    \new_[21410]_ , \new_[21411]_ , \new_[21412]_ , \new_[21413]_ ,
    \new_[21414]_ , \new_[21415]_ , \new_[21416]_ , \new_[21417]_ ,
    \new_[21418]_ , \new_[21419]_ , \new_[21420]_ , \new_[21421]_ ,
    \new_[21422]_ , \new_[21423]_ , \new_[21424]_ , \new_[21425]_ ,
    \new_[21426]_ , \new_[21427]_ , \new_[21428]_ , \new_[21429]_ ,
    \new_[21430]_ , \new_[21431]_ , \new_[21432]_ , \new_[21433]_ ,
    \new_[21434]_ , \new_[21435]_ , \new_[21436]_ , \new_[21437]_ ,
    \new_[21438]_ , \new_[21439]_ , \new_[21440]_ , \new_[21441]_ ,
    \new_[21442]_ , \new_[21443]_ , \new_[21444]_ , \new_[21445]_ ,
    \new_[21446]_ , \new_[21447]_ , \new_[21448]_ , \new_[21449]_ ,
    \new_[21450]_ , \new_[21451]_ , \new_[21452]_ , \new_[21453]_ ,
    \new_[21454]_ , \new_[21455]_ , \new_[21456]_ , \new_[21457]_ ,
    \new_[21458]_ , \new_[21459]_ , \new_[21460]_ , \new_[21461]_ ,
    \new_[21462]_ , \new_[21463]_ , \new_[21464]_ , \new_[21465]_ ,
    \new_[21466]_ , \new_[21467]_ , \new_[21468]_ , \new_[21469]_ ,
    \new_[21470]_ , \new_[21471]_ , \new_[21472]_ , \new_[21473]_ ,
    \new_[21474]_ , \new_[21475]_ , \new_[21476]_ , \new_[21477]_ ,
    \new_[21478]_ , \new_[21479]_ , \new_[21480]_ , \new_[21481]_ ,
    \new_[21482]_ , \new_[21483]_ , \new_[21484]_ , \new_[21485]_ ,
    \new_[21486]_ , \new_[21487]_ , \new_[21488]_ , \new_[21489]_ ,
    \new_[21490]_ , \new_[21491]_ , \new_[21492]_ , \new_[21493]_ ,
    \new_[21494]_ , \new_[21495]_ , \new_[21496]_ , \new_[21497]_ ,
    \new_[21498]_ , \new_[21499]_ , \new_[21500]_ , \new_[21501]_ ,
    \new_[21502]_ , \new_[21503]_ , \new_[21504]_ , \new_[21505]_ ,
    \new_[21506]_ , \new_[21507]_ , \new_[21508]_ , \new_[21509]_ ,
    \new_[21510]_ , \new_[21511]_ , \new_[21512]_ , \new_[21513]_ ,
    \new_[21514]_ , \new_[21515]_ , \new_[21516]_ , \new_[21517]_ ,
    \new_[21518]_ , \new_[21519]_ , \new_[21520]_ , \new_[21521]_ ,
    \new_[21522]_ , \new_[21523]_ , \new_[21524]_ , \new_[21525]_ ,
    \new_[21526]_ , \new_[21527]_ , \new_[21528]_ , \new_[21529]_ ,
    \new_[21530]_ , \new_[21531]_ , \new_[21532]_ , \new_[21533]_ ,
    \new_[21534]_ , \new_[21535]_ , \new_[21536]_ , \new_[21537]_ ,
    \new_[21538]_ , \new_[21539]_ , \new_[21540]_ , \new_[21541]_ ,
    \new_[21542]_ , \new_[21543]_ , \new_[21544]_ , \new_[21545]_ ,
    \new_[21546]_ , \new_[21547]_ , \new_[21548]_ , \new_[21549]_ ,
    \new_[21550]_ , \new_[21551]_ , \new_[21552]_ , \new_[21553]_ ,
    \new_[21554]_ , \new_[21555]_ , \new_[21556]_ , \new_[21557]_ ,
    \new_[21558]_ , \new_[21559]_ , \new_[21560]_ , \new_[21561]_ ,
    \new_[21562]_ , \new_[21563]_ , \new_[21564]_ , \new_[21565]_ ,
    \new_[21566]_ , \new_[21567]_ , \new_[21568]_ , \new_[21569]_ ,
    \new_[21570]_ , \new_[21571]_ , \new_[21572]_ , \new_[21573]_ ,
    \new_[21574]_ , \new_[21575]_ , \new_[21576]_ , \new_[21577]_ ,
    \new_[21578]_ , \new_[21579]_ , \new_[21580]_ , \new_[21581]_ ,
    \new_[21582]_ , \new_[21583]_ , \new_[21584]_ , \new_[21585]_ ,
    \new_[21586]_ , \new_[21587]_ , \new_[21588]_ , \new_[21589]_ ,
    \new_[21590]_ , \new_[21591]_ , \new_[21592]_ , \new_[21593]_ ,
    \new_[21594]_ , \new_[21595]_ , \new_[21596]_ , \new_[21597]_ ,
    \new_[21598]_ , \new_[21599]_ , \new_[21600]_ , \new_[21601]_ ,
    \new_[21602]_ , \new_[21603]_ , \new_[21604]_ , \new_[21605]_ ,
    \new_[21606]_ , \new_[21607]_ , \new_[21608]_ , \new_[21609]_ ,
    \new_[21610]_ , \new_[21611]_ , \new_[21612]_ , \new_[21613]_ ,
    \new_[21614]_ , \new_[21615]_ , \new_[21616]_ , \new_[21617]_ ,
    \new_[21618]_ , \new_[21620]_ , \new_[21621]_ , \new_[21622]_ ,
    \new_[21623]_ , \new_[21624]_ , \new_[21625]_ , \new_[21626]_ ,
    \new_[21627]_ , \new_[21628]_ , \new_[21629]_ , \new_[21630]_ ,
    \new_[21631]_ , \new_[21632]_ , \new_[21633]_ , \new_[21634]_ ,
    \new_[21635]_ , \new_[21636]_ , \new_[21637]_ , \new_[21638]_ ,
    \new_[21639]_ , \new_[21640]_ , \new_[21641]_ , \new_[21642]_ ,
    \new_[21643]_ , \new_[21644]_ , \new_[21645]_ , \new_[21646]_ ,
    \new_[21647]_ , \new_[21648]_ , \new_[21649]_ , \new_[21650]_ ,
    \new_[21651]_ , \new_[21652]_ , \new_[21653]_ , \new_[21654]_ ,
    \new_[21655]_ , \new_[21656]_ , \new_[21657]_ , \new_[21658]_ ,
    \new_[21659]_ , \new_[21660]_ , \new_[21661]_ , \new_[21662]_ ,
    \new_[21663]_ , \new_[21664]_ , \new_[21665]_ , \new_[21666]_ ,
    \new_[21667]_ , \new_[21668]_ , \new_[21669]_ , \new_[21670]_ ,
    \new_[21671]_ , \new_[21672]_ , \new_[21673]_ , \new_[21674]_ ,
    \new_[21675]_ , \new_[21676]_ , \new_[21677]_ , \new_[21678]_ ,
    \new_[21679]_ , \new_[21680]_ , \new_[21681]_ , \new_[21682]_ ,
    \new_[21683]_ , \new_[21684]_ , \new_[21685]_ , \new_[21686]_ ,
    \new_[21687]_ , \new_[21688]_ , \new_[21689]_ , \new_[21690]_ ,
    \new_[21691]_ , \new_[21692]_ , \new_[21693]_ , \new_[21694]_ ,
    \new_[21695]_ , \new_[21696]_ , \new_[21697]_ , \new_[21698]_ ,
    \new_[21699]_ , \new_[21700]_ , \new_[21701]_ , \new_[21702]_ ,
    \new_[21703]_ , \new_[21704]_ , \new_[21705]_ , \new_[21706]_ ,
    \new_[21707]_ , \new_[21708]_ , \new_[21709]_ , \new_[21710]_ ,
    \new_[21711]_ , \new_[21712]_ , \new_[21713]_ , \new_[21714]_ ,
    \new_[21715]_ , \new_[21716]_ , \new_[21717]_ , \new_[21718]_ ,
    \new_[21719]_ , \new_[21720]_ , \new_[21721]_ , \new_[21722]_ ,
    \new_[21723]_ , \new_[21724]_ , \new_[21725]_ , \new_[21726]_ ,
    \new_[21727]_ , \new_[21728]_ , \new_[21729]_ , \new_[21730]_ ,
    \new_[21731]_ , \new_[21732]_ , \new_[21733]_ , \new_[21734]_ ,
    \new_[21735]_ , \new_[21736]_ , \new_[21737]_ , \new_[21738]_ ,
    \new_[21739]_ , \new_[21740]_ , \new_[21741]_ , \new_[21742]_ ,
    \new_[21743]_ , \new_[21744]_ , \new_[21745]_ , \new_[21746]_ ,
    \new_[21747]_ , \new_[21748]_ , \new_[21749]_ , \new_[21750]_ ,
    \new_[21751]_ , \new_[21752]_ , \new_[21753]_ , \new_[21754]_ ,
    \new_[21755]_ , \new_[21756]_ , \new_[21757]_ , \new_[21758]_ ,
    \new_[21759]_ , \new_[21760]_ , \new_[21761]_ , \new_[21762]_ ,
    \new_[21763]_ , \new_[21764]_ , \new_[21765]_ , \new_[21766]_ ,
    \new_[21767]_ , \new_[21768]_ , \new_[21769]_ , \new_[21770]_ ,
    \new_[21771]_ , \new_[21772]_ , \new_[21773]_ , \new_[21774]_ ,
    \new_[21775]_ , \new_[21776]_ , \new_[21777]_ , \new_[21778]_ ,
    \new_[21779]_ , \new_[21780]_ , \new_[21781]_ , \new_[21782]_ ,
    \new_[21783]_ , \new_[21784]_ , \new_[21785]_ , \new_[21786]_ ,
    \new_[21787]_ , \new_[21788]_ , \new_[21789]_ , \new_[21790]_ ,
    \new_[21791]_ , \new_[21792]_ , \new_[21793]_ , \new_[21794]_ ,
    \new_[21795]_ , \new_[21796]_ , \new_[21797]_ , \new_[21798]_ ,
    \new_[21799]_ , \new_[21800]_ , \new_[21801]_ , \new_[21802]_ ,
    \new_[21803]_ , \new_[21804]_ , \new_[21805]_ , \new_[21806]_ ,
    \new_[21807]_ , \new_[21808]_ , \new_[21809]_ , \new_[21810]_ ,
    \new_[21811]_ , \new_[21812]_ , \new_[21813]_ , \new_[21814]_ ,
    \new_[21815]_ , \new_[21816]_ , \new_[21817]_ , \new_[21818]_ ,
    \new_[21819]_ , \new_[21820]_ , \new_[21821]_ , \new_[21822]_ ,
    \new_[21823]_ , \new_[21824]_ , \new_[21825]_ , \new_[21826]_ ,
    \new_[21827]_ , \new_[21828]_ , \new_[21829]_ , \new_[21830]_ ,
    \new_[21831]_ , \new_[21832]_ , \new_[21833]_ , \new_[21834]_ ,
    \new_[21835]_ , \new_[21836]_ , \new_[21837]_ , \new_[21838]_ ,
    \new_[21839]_ , \new_[21840]_ , \new_[21841]_ , \new_[21842]_ ,
    \new_[21843]_ , \new_[21844]_ , \new_[21845]_ , \new_[21846]_ ,
    \new_[21847]_ , \new_[21848]_ , \new_[21849]_ , \new_[21850]_ ,
    \new_[21851]_ , \new_[21852]_ , \new_[21853]_ , \new_[21854]_ ,
    \new_[21855]_ , \new_[21856]_ , \new_[21857]_ , \new_[21858]_ ,
    \new_[21859]_ , \new_[21860]_ , \new_[21861]_ , \new_[21862]_ ,
    \new_[21863]_ , \new_[21864]_ , \new_[21865]_ , \new_[21866]_ ,
    \new_[21867]_ , \new_[21868]_ , \new_[21869]_ , \new_[21870]_ ,
    \new_[21871]_ , \new_[21872]_ , \new_[21873]_ , \new_[21874]_ ,
    \new_[21875]_ , \new_[21876]_ , \new_[21877]_ , \new_[21878]_ ,
    \new_[21879]_ , \new_[21880]_ , \new_[21881]_ , \new_[21882]_ ,
    \new_[21883]_ , \new_[21884]_ , \new_[21885]_ , \new_[21886]_ ,
    \new_[21887]_ , \new_[21888]_ , \new_[21889]_ , \new_[21890]_ ,
    \new_[21891]_ , \new_[21892]_ , \new_[21893]_ , \new_[21894]_ ,
    \new_[21895]_ , \new_[21896]_ , \new_[21897]_ , \new_[21898]_ ,
    \new_[21899]_ , \new_[21900]_ , \new_[21901]_ , \new_[21902]_ ,
    \new_[21903]_ , \new_[21904]_ , \new_[21905]_ , \new_[21906]_ ,
    \new_[21907]_ , \new_[21908]_ , \new_[21909]_ , \new_[21910]_ ,
    \new_[21911]_ , \new_[21912]_ , \new_[21913]_ , \new_[21914]_ ,
    \new_[21915]_ , \new_[21916]_ , \new_[21917]_ , \new_[21918]_ ,
    \new_[21919]_ , \new_[21920]_ , \new_[21921]_ , \new_[21922]_ ,
    \new_[21923]_ , \new_[21924]_ , \new_[21925]_ , \new_[21926]_ ,
    \new_[21927]_ , \new_[21928]_ , \new_[21929]_ , \new_[21930]_ ,
    \new_[21931]_ , \new_[21932]_ , \new_[21933]_ , \new_[21934]_ ,
    \new_[21935]_ , \new_[21936]_ , \new_[21937]_ , \new_[21938]_ ,
    \new_[21939]_ , \new_[21940]_ , \new_[21941]_ , \new_[21942]_ ,
    \new_[21943]_ , \new_[21944]_ , \new_[21945]_ , \new_[21946]_ ,
    \new_[21947]_ , \new_[21948]_ , \new_[21949]_ , \new_[21950]_ ,
    \new_[21951]_ , \new_[21952]_ , \new_[21953]_ , \new_[21954]_ ,
    \new_[21955]_ , \new_[21956]_ , \new_[21957]_ , \new_[21958]_ ,
    \new_[21959]_ , \new_[21960]_ , \new_[21961]_ , \new_[21962]_ ,
    \new_[21963]_ , \new_[21964]_ , \new_[21965]_ , \new_[21966]_ ,
    \new_[21967]_ , \new_[21968]_ , \new_[21969]_ , \new_[21970]_ ,
    \new_[21971]_ , \new_[21972]_ , \new_[21973]_ , \new_[21974]_ ,
    \new_[21975]_ , \new_[21976]_ , \new_[21977]_ , \new_[21978]_ ,
    \new_[21979]_ , \new_[21980]_ , \new_[21981]_ , \new_[21982]_ ,
    \new_[21983]_ , \new_[21984]_ , \new_[21985]_ , \new_[21986]_ ,
    \new_[21987]_ , \new_[21988]_ , \new_[21989]_ , \new_[21990]_ ,
    \new_[21991]_ , \new_[21992]_ , \new_[21993]_ , \new_[21994]_ ,
    \new_[21995]_ , \new_[21996]_ , \new_[21998]_ , \new_[21999]_ ,
    \new_[22000]_ , \new_[22001]_ , \new_[22002]_ , \new_[22003]_ ,
    \new_[22004]_ , \new_[22005]_ , \new_[22006]_ , \new_[22007]_ ,
    \new_[22008]_ , \new_[22009]_ , \new_[22010]_ , \new_[22011]_ ,
    \new_[22012]_ , \new_[22013]_ , \new_[22014]_ , \new_[22015]_ ,
    \new_[22016]_ , \new_[22017]_ , \new_[22018]_ , \new_[22019]_ ,
    \new_[22025]_ , \new_[22029]_ , \new_[22037]_ , \new_[22043]_ ,
    \new_[22047]_ , \new_[22053]_ , \new_[22062]_ , \new_[22067]_ ,
    \new_[22069]_ , \new_[22071]_ , \new_[22075]_ , \new_[22076]_ ,
    \new_[22077]_ , \new_[22078]_ , \new_[22079]_ , \new_[22080]_ ,
    \new_[22081]_ , \new_[22082]_ , \new_[22083]_ , \new_[22084]_ ,
    \new_[22085]_ , \new_[22086]_ , \new_[22087]_ , \new_[22088]_ ,
    \new_[22089]_ , \new_[22090]_ , \new_[22092]_ , \new_[22093]_ ,
    \new_[22094]_ , \new_[22095]_ , \new_[22096]_ , \new_[22097]_ ,
    \new_[22098]_ , \new_[22099]_ , \new_[22100]_ , \new_[22101]_ ,
    \new_[22102]_ , \new_[22103]_ , \new_[22104]_ , \new_[22105]_ ,
    \new_[22106]_ , \new_[22107]_ , \new_[22108]_ , \new_[22109]_ ,
    \new_[22110]_ , \new_[22111]_ , \new_[22112]_ , \new_[22113]_ ,
    \new_[22114]_ , \new_[22115]_ , \new_[22116]_ , \new_[22117]_ ,
    \new_[22118]_ , \new_[22119]_ , \new_[22120]_ , \new_[22121]_ ,
    \new_[22122]_ , \new_[22123]_ , \new_[22124]_ , \new_[22125]_ ,
    \new_[22126]_ , \new_[22127]_ , \new_[22128]_ , \new_[22129]_ ,
    \new_[22130]_ , \new_[22131]_ , \new_[22132]_ , \new_[22133]_ ,
    \new_[22134]_ , \new_[22135]_ , \new_[22136]_ , \new_[22137]_ ,
    \new_[22138]_ , \new_[22139]_ , \new_[22140]_ , \new_[22142]_ ,
    \new_[22143]_ , \new_[22144]_ , \new_[22145]_ , \new_[22146]_ ,
    \new_[22147]_ , \new_[22148]_ , \new_[22149]_ , \new_[22150]_ ,
    \new_[22151]_ , \new_[22152]_ , \new_[22153]_ , \new_[22155]_ ,
    \new_[22156]_ , \new_[22157]_ , \new_[22158]_ , \new_[22159]_ ,
    \new_[22160]_ , \new_[22161]_ , \new_[22162]_ , \new_[22163]_ ,
    \new_[22164]_ , \new_[22165]_ , \new_[22166]_ , \new_[22167]_ ,
    \new_[22168]_ , \new_[22169]_ , \new_[22170]_ , \new_[22171]_ ,
    \new_[22172]_ , \new_[22173]_ , \new_[22174]_ , \new_[22175]_ ,
    \new_[22176]_ , \new_[22177]_ , \new_[22178]_ , \new_[22179]_ ,
    \new_[22180]_ , \new_[22181]_ , \new_[22182]_ , \new_[22183]_ ,
    \new_[22184]_ , \new_[22185]_ , \new_[22186]_ , \new_[22187]_ ,
    \new_[22188]_ , \new_[22189]_ , \new_[22190]_ , \new_[22191]_ ,
    \new_[22192]_ , \new_[22193]_ , \new_[22194]_ , \new_[22195]_ ,
    \new_[22196]_ , \new_[22197]_ , \new_[22198]_ , \new_[22199]_ ,
    \new_[22200]_ , \new_[22201]_ , \new_[22202]_ , \new_[22203]_ ,
    \new_[22204]_ , \new_[22205]_ , \new_[22206]_ , \new_[22207]_ ,
    \new_[22208]_ , \new_[22209]_ , \new_[22210]_ , \new_[22211]_ ,
    \new_[22212]_ , \new_[22213]_ , \new_[22214]_ , \new_[22215]_ ,
    \new_[22216]_ , \new_[22217]_ , \new_[22218]_ , \new_[22219]_ ,
    \new_[22220]_ , \new_[22221]_ , \new_[22222]_ , \new_[22223]_ ,
    \new_[22224]_ , \new_[22225]_ , \new_[22226]_ , \new_[22227]_ ,
    \new_[22228]_ , \new_[22229]_ , \new_[22230]_ , \new_[22231]_ ,
    \new_[22232]_ , \new_[22233]_ , \new_[22234]_ , \new_[22235]_ ,
    \new_[22236]_ , \new_[22237]_ , \new_[22238]_ , \new_[22239]_ ,
    \new_[22240]_ , \new_[22241]_ , \new_[22242]_ , \new_[22243]_ ,
    \new_[22244]_ , \new_[22245]_ , \new_[22246]_ , \new_[22247]_ ,
    \new_[22248]_ , \new_[22249]_ , \new_[22250]_ , \new_[22251]_ ,
    \new_[22252]_ , \new_[22253]_ , \new_[22254]_ , \new_[22255]_ ,
    \new_[22256]_ , \new_[22257]_ , \new_[22258]_ , \new_[22259]_ ,
    \new_[22260]_ , \new_[22261]_ , \new_[22262]_ , \new_[22263]_ ,
    \new_[22264]_ , \new_[22265]_ , \new_[22266]_ , \new_[22267]_ ,
    \new_[22268]_ , \new_[22269]_ , \new_[22270]_ , \new_[22271]_ ,
    \new_[22272]_ , \new_[22273]_ , \new_[22274]_ , \new_[22275]_ ,
    \new_[22276]_ , \new_[22277]_ , \new_[22278]_ , \new_[22279]_ ,
    \new_[22280]_ , \new_[22281]_ , \new_[22282]_ , \new_[22283]_ ,
    \new_[22284]_ , \new_[22285]_ , \new_[22286]_ , \new_[22287]_ ,
    \new_[22288]_ , \new_[22289]_ , \new_[22290]_ , \new_[22291]_ ,
    \new_[22292]_ , \new_[22293]_ , \new_[22294]_ , \new_[22295]_ ,
    \new_[22296]_ , \new_[22297]_ , \new_[22298]_ , \new_[22299]_ ,
    \new_[22300]_ , \new_[22301]_ , \new_[22302]_ , \new_[22303]_ ,
    \new_[22304]_ , \new_[22305]_ , \new_[22306]_ , \new_[22307]_ ,
    \new_[22308]_ , \new_[22309]_ , \new_[22310]_ , \new_[22311]_ ,
    \new_[22312]_ , \new_[22313]_ , \new_[22314]_ , \new_[22315]_ ,
    \new_[22316]_ , \new_[22317]_ , \new_[22318]_ , \new_[22319]_ ,
    \new_[22320]_ , \new_[22321]_ , \new_[22322]_ , \new_[22323]_ ,
    \new_[22324]_ , \new_[22325]_ , \new_[22326]_ , \new_[22327]_ ,
    \new_[22328]_ , \new_[22329]_ , \new_[22330]_ , \new_[22331]_ ,
    \new_[22332]_ , \new_[22333]_ , \new_[22334]_ , \new_[22335]_ ,
    \new_[22336]_ , \new_[22337]_ , \new_[22338]_ , \new_[22339]_ ,
    \new_[22340]_ , \new_[22341]_ , \new_[22342]_ , \new_[22343]_ ,
    \new_[22344]_ , \new_[22345]_ , \new_[22346]_ , \new_[22347]_ ,
    \new_[22348]_ , \new_[22349]_ , \new_[22350]_ , \new_[22351]_ ,
    \new_[22352]_ , \new_[22353]_ , \new_[22354]_ , \new_[22355]_ ,
    \new_[22356]_ , \new_[22357]_ , \new_[22358]_ , \new_[22359]_ ,
    \new_[22360]_ , \new_[22361]_ , \new_[22362]_ , \new_[22363]_ ,
    \new_[22364]_ , \new_[22365]_ , \new_[22366]_ , \new_[22367]_ ,
    \new_[22368]_ , \new_[22369]_ , \new_[22370]_ , \new_[22371]_ ,
    \new_[22372]_ , \new_[22373]_ , \new_[22374]_ , \new_[22375]_ ,
    \new_[22376]_ , \new_[22377]_ , \new_[22378]_ , \new_[22379]_ ,
    \new_[22380]_ , \new_[22381]_ , \new_[22382]_ , \new_[22383]_ ,
    \new_[22384]_ , \new_[22385]_ , \new_[22386]_ , \new_[22387]_ ,
    \new_[22388]_ , \new_[22389]_ , \new_[22390]_ , \new_[22391]_ ,
    \new_[22392]_ , \new_[22393]_ , \new_[22394]_ , \new_[22395]_ ,
    \new_[22396]_ , \new_[22397]_ , \new_[22398]_ , \new_[22399]_ ,
    \new_[22400]_ , \new_[22401]_ , \new_[22402]_ , \new_[22403]_ ,
    \new_[22404]_ , \new_[22405]_ , \new_[22406]_ , \new_[22407]_ ,
    \new_[22408]_ , \new_[22409]_ , \new_[22410]_ , \new_[22411]_ ,
    \new_[22412]_ , \new_[22413]_ , \new_[22414]_ , \new_[22415]_ ,
    \new_[22416]_ , \new_[22417]_ , \new_[22418]_ , \new_[22419]_ ,
    \new_[22420]_ , \new_[22421]_ , \new_[22422]_ , \new_[22423]_ ,
    \new_[22424]_ , \new_[22425]_ , \new_[22426]_ , \new_[22427]_ ,
    \new_[22428]_ , \new_[22429]_ , \new_[22430]_ , \new_[22431]_ ,
    \new_[22432]_ , \new_[22433]_ , \new_[22434]_ , \new_[22435]_ ,
    \new_[22436]_ , \new_[22437]_ , \new_[22438]_ , \new_[22439]_ ,
    \new_[22440]_ , \new_[22441]_ , \new_[22442]_ , \new_[22443]_ ,
    \new_[22444]_ , \new_[22445]_ , \new_[22446]_ , \new_[22447]_ ,
    \new_[22448]_ , \new_[22449]_ , \new_[22450]_ , \new_[22451]_ ,
    \new_[22452]_ , \new_[22453]_ , \new_[22454]_ , \new_[22455]_ ,
    \new_[22456]_ , \new_[22457]_ , \new_[22458]_ , \new_[22459]_ ,
    \new_[22460]_ , \new_[22461]_ , \new_[22462]_ , \new_[22463]_ ,
    \new_[22464]_ , \new_[22465]_ , \new_[22466]_ , \new_[22467]_ ,
    \new_[22468]_ , \new_[22469]_ , \new_[22470]_ , \new_[22471]_ ,
    \new_[22472]_ , \new_[22473]_ , \new_[22474]_ , \new_[22475]_ ,
    \new_[22476]_ , \new_[22477]_ , \new_[22478]_ , \new_[22479]_ ,
    \new_[22480]_ , \new_[22481]_ , \new_[22482]_ , \new_[22483]_ ,
    \new_[22484]_ , \new_[22485]_ , \new_[22486]_ , \new_[22487]_ ,
    \new_[22488]_ , \new_[22489]_ , \new_[22490]_ , \new_[22491]_ ,
    \new_[22492]_ , \new_[22493]_ , \new_[22494]_ , \new_[22495]_ ,
    \new_[22496]_ , \new_[22497]_ , \new_[22498]_ , \new_[22499]_ ,
    \new_[22500]_ , \new_[22501]_ , \new_[22502]_ , \new_[22503]_ ,
    \new_[22504]_ , \new_[22505]_ , \new_[22506]_ , \new_[22507]_ ,
    \new_[22508]_ , \new_[22509]_ , \new_[22510]_ , \new_[22511]_ ,
    \new_[22512]_ , \new_[22513]_ , \new_[22514]_ , \new_[22515]_ ,
    \new_[22516]_ , \new_[22517]_ , \new_[22518]_ , \new_[22519]_ ,
    \new_[22520]_ , \new_[22521]_ , \new_[22522]_ , \new_[22523]_ ,
    \new_[22524]_ , \new_[22525]_ , \new_[22526]_ , \new_[22527]_ ,
    \new_[22528]_ , \new_[22529]_ , \new_[22530]_ , \new_[22531]_ ,
    \new_[22532]_ , \new_[22533]_ , \new_[22534]_ , \new_[22535]_ ,
    \new_[22536]_ , \new_[22537]_ , \new_[22538]_ , \new_[22539]_ ,
    \new_[22540]_ , \new_[22541]_ , \new_[22542]_ , \new_[22543]_ ,
    \new_[22544]_ , \new_[22545]_ , \new_[22546]_ , \new_[22547]_ ,
    \new_[22548]_ , \new_[22549]_ , \new_[22550]_ , \new_[22551]_ ,
    \new_[22552]_ , \new_[22553]_ , \new_[22554]_ , \new_[22555]_ ,
    \new_[22556]_ , \new_[22557]_ , \new_[22558]_ , \new_[22559]_ ,
    \new_[22560]_ , \new_[22561]_ , \new_[22562]_ , \new_[22563]_ ,
    \new_[22564]_ , \new_[22565]_ , \new_[22566]_ , \new_[22567]_ ,
    \new_[22568]_ , \new_[22569]_ , \new_[22570]_ , \new_[22571]_ ,
    \new_[22572]_ , \new_[22573]_ , \new_[22574]_ , \new_[22575]_ ,
    \new_[22576]_ , \new_[22577]_ , \new_[22578]_ , \new_[22579]_ ,
    \new_[22580]_ , \new_[22581]_ , \new_[22582]_ , \new_[22583]_ ,
    \new_[22584]_ , \new_[22585]_ , \new_[22586]_ , \new_[22587]_ ,
    \new_[22588]_ , \new_[22589]_ , \new_[22590]_ , \new_[22591]_ ,
    \new_[22592]_ , \new_[22593]_ , \new_[22594]_ , \new_[22595]_ ,
    \new_[22596]_ , \new_[22597]_ , \new_[22598]_ , \new_[22599]_ ,
    \new_[22600]_ , \new_[22601]_ , \new_[22602]_ , \new_[22603]_ ,
    \new_[22604]_ , \new_[22605]_ , \new_[22606]_ , \new_[22607]_ ,
    \new_[22608]_ , \new_[22609]_ , \new_[22610]_ , \new_[22611]_ ,
    \new_[22612]_ , \new_[22613]_ , \new_[22614]_ , \new_[22615]_ ,
    \new_[22616]_ , \new_[22617]_ , \new_[22618]_ , \new_[22619]_ ,
    \new_[22620]_ , \new_[22621]_ , \new_[22622]_ , \new_[22623]_ ,
    \new_[22624]_ , \new_[22625]_ , \new_[22626]_ , \new_[22627]_ ,
    \new_[22628]_ , \new_[22629]_ , \new_[22630]_ , \new_[22631]_ ,
    \new_[22632]_ , \new_[22633]_ , \new_[22634]_ , \new_[22635]_ ,
    \new_[22636]_ , \new_[22637]_ , \new_[22638]_ , \new_[22639]_ ,
    \new_[22640]_ , \new_[22641]_ , \new_[22642]_ , \new_[22643]_ ,
    \new_[22644]_ , \new_[22645]_ , \new_[22646]_ , \new_[22647]_ ,
    \new_[22648]_ , \new_[22649]_ , \new_[22650]_ , \new_[22651]_ ,
    \new_[22652]_ , \new_[22653]_ , \new_[22654]_ , \new_[22655]_ ,
    \new_[22656]_ , \new_[22657]_ , \new_[22658]_ , \new_[22659]_ ,
    \new_[22660]_ , \new_[22661]_ , \new_[22662]_ , \new_[22663]_ ,
    \new_[22664]_ , \new_[22665]_ , \new_[22666]_ , \new_[22667]_ ,
    \new_[22668]_ , \new_[22669]_ , \new_[22670]_ , \new_[22671]_ ,
    \new_[22672]_ , \new_[22673]_ , \new_[22674]_ , \new_[22675]_ ,
    \new_[22676]_ , \new_[22677]_ , \new_[22678]_ , \new_[22679]_ ,
    \new_[22680]_ , \new_[22681]_ , \new_[22682]_ , \new_[22683]_ ,
    \new_[22684]_ , \new_[22685]_ , \new_[22686]_ , \new_[22687]_ ,
    \new_[22688]_ , \new_[22689]_ , \new_[22690]_ , \new_[22691]_ ,
    \new_[22692]_ , \new_[22693]_ , \new_[22694]_ , \new_[22695]_ ,
    \new_[22696]_ , \new_[22697]_ , \new_[22698]_ , \new_[22699]_ ,
    \new_[22700]_ , \new_[22701]_ , \new_[22702]_ , \new_[22703]_ ,
    \new_[22704]_ , \new_[22705]_ , \new_[22706]_ , \new_[22707]_ ,
    \new_[22708]_ , \new_[22709]_ , \new_[22710]_ , \new_[22711]_ ,
    \new_[22712]_ , \new_[22713]_ , \new_[22714]_ , \new_[22715]_ ,
    \new_[22716]_ , \new_[22717]_ , \new_[22718]_ , \new_[22719]_ ,
    \new_[22720]_ , \new_[22721]_ , \new_[22722]_ , \new_[22723]_ ,
    \new_[22724]_ , \new_[22725]_ , \new_[22726]_ , \new_[22727]_ ,
    \new_[22728]_ , \new_[22729]_ , \new_[22730]_ , \new_[22731]_ ,
    \new_[22732]_ , \new_[22733]_ , \new_[22734]_ , \new_[22735]_ ,
    \new_[22736]_ , \new_[22737]_ , \new_[22738]_ , \new_[22739]_ ,
    \new_[22740]_ , \new_[22741]_ , \new_[22742]_ , \new_[22743]_ ,
    \new_[22744]_ , \new_[22745]_ , \new_[22746]_ , \new_[22747]_ ,
    \new_[22748]_ , \new_[22749]_ , \new_[22750]_ , \new_[22751]_ ,
    \new_[22752]_ , \new_[22753]_ , \new_[22754]_ , \new_[22755]_ ,
    \new_[22756]_ , \new_[22757]_ , \new_[22758]_ , \new_[22759]_ ,
    \new_[22760]_ , \new_[22761]_ , \new_[22762]_ , \new_[22763]_ ,
    \new_[22764]_ , \new_[22765]_ , \new_[22766]_ , \new_[22767]_ ,
    \new_[22768]_ , \new_[22769]_ , \new_[22770]_ , \new_[22771]_ ,
    \new_[22772]_ , \new_[22773]_ , \new_[22774]_ , \new_[22775]_ ,
    \new_[22776]_ , \new_[22777]_ , \new_[22778]_ , \new_[22779]_ ,
    \new_[22780]_ , \new_[22781]_ , \new_[22782]_ , \new_[22783]_ ,
    \new_[22784]_ , \new_[22785]_ , \new_[22786]_ , \new_[22787]_ ,
    \new_[22788]_ , \new_[22789]_ , \new_[22790]_ , \new_[22791]_ ,
    \new_[22792]_ , \new_[22793]_ , \new_[22794]_ , \new_[22795]_ ,
    \new_[22796]_ , \new_[22797]_ , \new_[22798]_ , \new_[22799]_ ,
    \new_[22800]_ , \new_[22801]_ , \new_[22802]_ , \new_[22803]_ ,
    \new_[22804]_ , \new_[22805]_ , \new_[22806]_ , \new_[22807]_ ,
    \new_[22808]_ , \new_[22809]_ , \new_[22810]_ , \new_[22811]_ ,
    \new_[22812]_ , \new_[22813]_ , \new_[22814]_ , \new_[22815]_ ,
    \new_[22816]_ , \new_[22817]_ , \new_[22818]_ , \new_[22819]_ ,
    \new_[22820]_ , \new_[22821]_ , \new_[22822]_ , \new_[22823]_ ,
    \new_[22824]_ , \new_[22825]_ , \new_[22826]_ , \new_[22827]_ ,
    \new_[22828]_ , \new_[22829]_ , \new_[22830]_ , \new_[22831]_ ,
    \new_[22832]_ , \new_[22833]_ , \new_[22834]_ , \new_[22835]_ ,
    \new_[22836]_ , \new_[22837]_ , \new_[22838]_ , \new_[22839]_ ,
    \new_[22840]_ , \new_[22841]_ , \new_[22842]_ , \new_[22843]_ ,
    \new_[22844]_ , \new_[22845]_ , \new_[22846]_ , \new_[22847]_ ,
    \new_[22848]_ , \new_[22849]_ , \new_[22850]_ , \new_[22851]_ ,
    \new_[22852]_ , \new_[22853]_ , \new_[22854]_ , \new_[22855]_ ,
    \new_[22856]_ , \new_[22857]_ , \new_[22858]_ , \new_[22859]_ ,
    \new_[22860]_ , \new_[22861]_ , \new_[22862]_ , \new_[22863]_ ,
    \new_[22864]_ , \new_[22865]_ , \new_[22866]_ , \new_[22867]_ ,
    \new_[22868]_ , \new_[22869]_ , \new_[22870]_ , \new_[22871]_ ,
    \new_[22872]_ , \new_[22873]_ , \new_[22874]_ , \new_[22875]_ ,
    \new_[22876]_ , \new_[22877]_ , \new_[22878]_ , \new_[22879]_ ,
    \new_[22880]_ , \new_[22881]_ , \new_[22882]_ , \new_[22883]_ ,
    \new_[22884]_ , \new_[22885]_ , \new_[22886]_ , \new_[22887]_ ,
    \new_[22888]_ , \new_[22889]_ , \new_[22890]_ , \new_[22891]_ ,
    \new_[22892]_ , \new_[22893]_ , \new_[22894]_ , \new_[22895]_ ,
    \new_[22896]_ , \new_[22897]_ , \new_[22898]_ , \new_[22899]_ ,
    \new_[22900]_ , \new_[22901]_ , \new_[22902]_ , \new_[22903]_ ,
    \new_[22904]_ , \new_[22905]_ , \new_[22906]_ , \new_[22907]_ ,
    \new_[22908]_ , \new_[22909]_ , \new_[22910]_ , \new_[22911]_ ,
    \new_[22912]_ , \new_[22913]_ , \new_[22914]_ , \new_[22915]_ ,
    \new_[22916]_ , \new_[22917]_ , \new_[22918]_ , \new_[22919]_ ,
    \new_[22920]_ , \new_[22921]_ , \new_[22922]_ , \new_[22923]_ ,
    \new_[22924]_ , \new_[22925]_ , \new_[22926]_ , \new_[22927]_ ,
    \new_[22928]_ , \new_[22929]_ , \new_[22930]_ , \new_[22931]_ ,
    \new_[22932]_ , \new_[22933]_ , \new_[22934]_ , \new_[22935]_ ,
    \new_[22936]_ , \new_[22937]_ , \new_[22938]_ , \new_[22939]_ ,
    \new_[22940]_ , \new_[22941]_ , \new_[22942]_ , \new_[22943]_ ,
    \new_[22944]_ , \new_[22945]_ , \new_[22946]_ , \new_[22947]_ ,
    \new_[22948]_ , \new_[22949]_ , \new_[22950]_ , \new_[22951]_ ,
    \new_[22952]_ , \new_[22953]_ , \new_[22954]_ , \new_[22955]_ ,
    \new_[22956]_ , \new_[22957]_ , \new_[22958]_ , \new_[22959]_ ,
    \new_[22960]_ , \new_[22961]_ , \new_[22962]_ , \new_[22963]_ ,
    \new_[22964]_ , \new_[22965]_ , \new_[22966]_ , \new_[22967]_ ,
    \new_[22968]_ , \new_[22969]_ , \new_[22970]_ , \new_[22971]_ ,
    \new_[22972]_ , \new_[22973]_ , \new_[22974]_ , \new_[22975]_ ,
    \new_[22976]_ , \new_[22977]_ , \new_[22978]_ , \new_[22979]_ ,
    \new_[22980]_ , \new_[22981]_ , \new_[22982]_ , \new_[22983]_ ,
    \new_[22984]_ , \new_[22985]_ , \new_[22986]_ , \new_[22987]_ ,
    \new_[22988]_ , \new_[22989]_ , \new_[22990]_ , \new_[22991]_ ,
    \new_[22992]_ , \new_[22993]_ , \new_[22994]_ , \new_[22995]_ ,
    \new_[22996]_ , \new_[22997]_ , \new_[22998]_ , \new_[22999]_ ,
    \new_[23000]_ , \new_[23001]_ , \new_[23002]_ , \new_[23003]_ ,
    \new_[23004]_ , \new_[23005]_ , \new_[23006]_ , \new_[23007]_ ,
    \new_[23008]_ , \new_[23009]_ , \new_[23010]_ , \new_[23011]_ ,
    \new_[23012]_ , \new_[23013]_ , \new_[23014]_ , \new_[23015]_ ,
    \new_[23016]_ , \new_[23017]_ , \new_[23018]_ , \new_[23019]_ ,
    \new_[23020]_ , \new_[23021]_ , \new_[23022]_ , \new_[23023]_ ,
    \new_[23024]_ , \new_[23025]_ , \new_[23026]_ , \new_[23027]_ ,
    \new_[23028]_ , \new_[23029]_ , \new_[23030]_ , \new_[23031]_ ,
    \new_[23032]_ , \new_[23033]_ , \new_[23034]_ , \new_[23035]_ ,
    \new_[23036]_ , \new_[23037]_ , \new_[23038]_ , \new_[23039]_ ,
    \new_[23040]_ , \new_[23041]_ , \new_[23042]_ , \new_[23043]_ ,
    \new_[23044]_ , \new_[23045]_ , \new_[23046]_ , \new_[23047]_ ,
    \new_[23048]_ , \new_[23049]_ , \new_[23050]_ , \new_[23051]_ ,
    \new_[23052]_ , \new_[23053]_ , \new_[23054]_ , \new_[23055]_ ,
    \new_[23056]_ , \new_[23057]_ , \new_[23058]_ , \new_[23059]_ ,
    \new_[23060]_ , \new_[23061]_ , \new_[23062]_ , \new_[23063]_ ,
    \new_[23064]_ , \new_[23065]_ , \new_[23066]_ , \new_[23067]_ ,
    \new_[23068]_ , \new_[23069]_ , \new_[23070]_ , \new_[23071]_ ,
    \new_[23072]_ , \new_[23073]_ , \new_[23074]_ , \new_[23075]_ ,
    \new_[23076]_ , \new_[23077]_ , \new_[23078]_ , \new_[23079]_ ,
    \new_[23080]_ , \new_[23081]_ , \new_[23082]_ , \new_[23083]_ ,
    \new_[23084]_ , \new_[23085]_ , \new_[23086]_ , \new_[23087]_ ,
    \new_[23088]_ , \new_[23089]_ , \new_[23090]_ , \new_[23091]_ ,
    \new_[23092]_ , \new_[23093]_ , \new_[23094]_ , \new_[23095]_ ,
    \new_[23096]_ , \new_[23097]_ , \new_[23098]_ , \new_[23099]_ ,
    \new_[23100]_ , \new_[23101]_ , \new_[23102]_ , \new_[23103]_ ,
    \new_[23104]_ , \new_[23105]_ , \new_[23106]_ , \new_[23107]_ ,
    \new_[23108]_ , \new_[23109]_ , \new_[23110]_ , \new_[23111]_ ,
    \new_[23112]_ , \new_[23113]_ , \new_[23114]_ , \new_[23115]_ ,
    \new_[23116]_ , \new_[23117]_ , \new_[23118]_ , \new_[23119]_ ,
    \new_[23120]_ , \new_[23121]_ , \new_[23122]_ , \new_[23123]_ ,
    \new_[23124]_ , \new_[23125]_ , \new_[23126]_ , \new_[23127]_ ,
    \new_[23128]_ , \new_[23129]_ , \new_[23130]_ , \new_[23131]_ ,
    \new_[23132]_ , \new_[23133]_ , \new_[23134]_ , \new_[23135]_ ,
    \new_[23136]_ , \new_[23137]_ , \new_[23138]_ , \new_[23139]_ ,
    \new_[23140]_ , \new_[23141]_ , \new_[23142]_ , \new_[23143]_ ,
    \new_[23144]_ , \new_[23145]_ , \new_[23146]_ , \new_[23147]_ ,
    \new_[23148]_ , \new_[23149]_ , \new_[23150]_ , \new_[23152]_ ,
    \new_[23153]_ , \new_[23154]_ , \new_[23155]_ , \new_[23156]_ ,
    \new_[23157]_ , \new_[23158]_ , \new_[23160]_ , \new_[23162]_ ,
    \new_[23163]_ , \new_[23164]_ , \new_[23165]_ , \new_[23166]_ ,
    \new_[23167]_ , \new_[23168]_ , \new_[23169]_ , \new_[23170]_ ,
    \new_[23171]_ , \new_[23172]_ , \new_[23173]_ , \new_[23174]_ ,
    \new_[23175]_ , \new_[23176]_ , \new_[23177]_ , \new_[23178]_ ,
    \new_[23179]_ , \new_[23180]_ , \new_[23181]_ , \new_[23182]_ ,
    \new_[23183]_ , \new_[23184]_ , \new_[23185]_ , \new_[23186]_ ,
    \new_[23187]_ , \new_[23188]_ , \new_[23189]_ , \new_[23190]_ ,
    \new_[23191]_ , \new_[23192]_ , \new_[23193]_ , \new_[23194]_ ,
    \new_[23195]_ , \new_[23196]_ , \new_[23197]_ , \new_[23198]_ ,
    \new_[23199]_ , \new_[23200]_ , \new_[23201]_ , \new_[23202]_ ,
    \new_[23203]_ , \new_[23204]_ , \new_[23205]_ , \new_[23206]_ ,
    \new_[23207]_ , \new_[23208]_ , \new_[23209]_ , \new_[23210]_ ,
    \new_[23211]_ , \new_[23212]_ , \new_[23213]_ , \new_[23214]_ ,
    \new_[23215]_ , \new_[23216]_ , \new_[23217]_ , \new_[23218]_ ,
    \new_[23219]_ , \new_[23220]_ , \new_[23221]_ , \new_[23222]_ ,
    \new_[23223]_ , \new_[23224]_ , \new_[23225]_ , \new_[23226]_ ,
    \new_[23227]_ , \new_[23228]_ , \new_[23229]_ , \new_[23230]_ ,
    \new_[23231]_ , \new_[23232]_ , \new_[23233]_ , \new_[23234]_ ,
    \new_[23235]_ , \new_[23236]_ , \new_[23237]_ , \new_[23238]_ ,
    \new_[23239]_ , \new_[23240]_ , \new_[23241]_ , \new_[23242]_ ,
    \new_[23243]_ , \new_[23244]_ , \new_[23245]_ , \new_[23246]_ ,
    \new_[23247]_ , \new_[23248]_ , \new_[23249]_ , \new_[23250]_ ,
    \new_[23251]_ , \new_[23252]_ , \new_[23253]_ , \new_[23254]_ ,
    \new_[23255]_ , \new_[23256]_ , \new_[23257]_ , \new_[23258]_ ,
    \new_[23259]_ , \new_[23260]_ , \new_[23261]_ , \new_[23262]_ ,
    \new_[23263]_ , \new_[23264]_ , \new_[23265]_ , \new_[23266]_ ,
    \new_[23267]_ , \new_[23268]_ , \new_[23269]_ , \new_[23270]_ ,
    \new_[23271]_ , \new_[23272]_ , \new_[23273]_ , \new_[23274]_ ,
    \new_[23275]_ , \new_[23276]_ , \new_[23277]_ , \new_[23278]_ ,
    \new_[23279]_ , \new_[23280]_ , \new_[23281]_ , \new_[23302]_ ,
    \new_[23306]_ , \new_[23321]_ , \new_[23326]_ , \new_[23327]_ ,
    \new_[23328]_ , \new_[23329]_ , \new_[23330]_ , \new_[23331]_ ,
    \new_[23332]_ , \new_[23333]_ , \new_[23334]_ , \new_[23335]_ ,
    \new_[23336]_ , \new_[23337]_ , \new_[23338]_ , \new_[23339]_ ,
    \new_[23340]_ , \new_[23341]_ , \new_[23342]_ , \new_[23343]_ ,
    \new_[23344]_ , \new_[23345]_ , \new_[23346]_ , \new_[23347]_ ,
    \new_[23348]_ , \new_[23349]_ , \new_[23350]_ , \new_[23351]_ ,
    \new_[23352]_ , \new_[23353]_ , \new_[23354]_ , \new_[23355]_ ,
    \new_[23356]_ , \new_[23357]_ , \new_[23358]_ , \new_[23359]_ ,
    \new_[23360]_ , \new_[23361]_ , \new_[23362]_ , \new_[23363]_ ,
    \new_[23364]_ , \new_[23365]_ , \new_[23366]_ , \new_[23367]_ ,
    \new_[23368]_ , \new_[23369]_ , \new_[23370]_ , \new_[23371]_ ,
    \new_[23372]_ , \new_[23373]_ , \new_[23374]_ , \new_[23375]_ ,
    \new_[23376]_ , \new_[23377]_ , \new_[23378]_ , \new_[23379]_ ,
    \new_[23380]_ , \new_[23381]_ , \new_[23382]_ , \new_[23383]_ ,
    \new_[23384]_ , \new_[23385]_ , \new_[23386]_ , \new_[23387]_ ,
    \new_[23388]_ , \new_[23389]_ , \new_[23390]_ , \new_[23391]_ ,
    \new_[23392]_ , \new_[23393]_ , \new_[23394]_ , \new_[23395]_ ,
    \new_[23396]_ , \new_[23397]_ , \new_[23398]_ , \new_[23399]_ ,
    \new_[23400]_ , \new_[23401]_ , \new_[23402]_ , \new_[23403]_ ,
    \new_[23404]_ , \new_[23405]_ , \new_[23406]_ , \new_[23407]_ ,
    \new_[23408]_ , \new_[23409]_ , \new_[23410]_ , \new_[23411]_ ,
    \new_[23412]_ , \new_[23413]_ , \new_[23414]_ , \new_[23415]_ ,
    \new_[23416]_ , \new_[23417]_ , \new_[23418]_ , \new_[23419]_ ,
    \new_[23420]_ , \new_[23421]_ , \new_[23422]_ , \new_[23423]_ ,
    \new_[23424]_ , \new_[23425]_ , \new_[23426]_ , \new_[23427]_ ,
    \new_[23428]_ , \new_[23429]_ , \new_[23430]_ , \new_[23431]_ ,
    \new_[23432]_ , \new_[23433]_ , \new_[23434]_ , \new_[23435]_ ,
    \new_[23436]_ , \new_[23437]_ , \new_[23438]_ , \new_[23439]_ ,
    \new_[23440]_ , \new_[23441]_ , \new_[23442]_ , \new_[23443]_ ,
    \new_[23444]_ , \new_[23445]_ , \new_[23446]_ , \new_[23447]_ ,
    \new_[23448]_ , \new_[23449]_ , \new_[23450]_ , \new_[23451]_ ,
    \new_[23452]_ , \new_[23453]_ , \new_[23454]_ , \new_[23455]_ ,
    \new_[23456]_ , \new_[23457]_ , \new_[23458]_ , \new_[23459]_ ,
    \new_[23460]_ , \new_[23461]_ , \new_[23462]_ , \new_[23463]_ ,
    \new_[23464]_ , \new_[23465]_ , \new_[23466]_ , \new_[23467]_ ,
    \new_[23468]_ , \new_[23469]_ , \new_[23470]_ , \new_[23471]_ ,
    \new_[23472]_ , \new_[23473]_ , \new_[23474]_ , \new_[23475]_ ,
    \new_[23476]_ , \new_[23477]_ , \new_[23478]_ , \new_[23479]_ ,
    \new_[23480]_ , \new_[23481]_ , \new_[23482]_ , \new_[23483]_ ,
    \new_[23484]_ , \new_[23485]_ , \new_[23486]_ , \new_[23487]_ ,
    \new_[23488]_ , \new_[23489]_ , \new_[23490]_ , \new_[23491]_ ,
    \new_[23492]_ , \new_[23493]_ , \new_[23494]_ , \new_[23495]_ ,
    \new_[23496]_ , \new_[23497]_ , \new_[23498]_ , \new_[23499]_ ,
    \new_[23500]_ , \new_[23501]_ , \new_[23502]_ , \new_[23503]_ ,
    \new_[23504]_ , \new_[23505]_ , \new_[23506]_ , \new_[23507]_ ,
    \new_[23508]_ , \new_[23509]_ , \new_[23510]_ , \new_[23511]_ ,
    \new_[23512]_ , \new_[23513]_ , \new_[23514]_ , \new_[23515]_ ,
    \new_[23516]_ , \new_[23517]_ , \new_[23518]_ , \new_[23519]_ ,
    \new_[23520]_ , \new_[23521]_ , \new_[23522]_ , \new_[23523]_ ,
    \new_[23524]_ , \new_[23525]_ , \new_[23526]_ , \new_[23527]_ ,
    \new_[23528]_ , \new_[23529]_ , \new_[23530]_ , \new_[23531]_ ,
    \new_[23532]_ , \new_[23533]_ , \new_[23534]_ , \new_[23535]_ ,
    \new_[23536]_ , \new_[23537]_ , \new_[23538]_ , \new_[23539]_ ,
    \new_[23540]_ , \new_[23541]_ , \new_[23542]_ , \new_[23543]_ ,
    \new_[23544]_ , \new_[23545]_ , \new_[23546]_ , \new_[23547]_ ,
    \new_[23548]_ , \new_[23549]_ , \new_[23550]_ , \new_[23551]_ ,
    \new_[23552]_ , \new_[23553]_ , \new_[23554]_ , \new_[23555]_ ,
    \new_[23556]_ , \new_[23557]_ , \new_[23558]_ , \new_[23559]_ ,
    \new_[23560]_ , \new_[23561]_ , \new_[23562]_ , \new_[23563]_ ,
    \new_[23564]_ , \new_[23565]_ , \new_[23566]_ , \new_[23567]_ ,
    \new_[23568]_ , \new_[23569]_ , \new_[23570]_ , \new_[23571]_ ,
    \new_[23572]_ , \new_[23573]_ , \new_[23574]_ , \new_[23575]_ ,
    \new_[23576]_ , \new_[23577]_ , \new_[23578]_ , \new_[23579]_ ,
    \new_[23580]_ , \new_[23581]_ , \new_[23582]_ , \new_[23583]_ ,
    \new_[23584]_ , \new_[23585]_ , \new_[23586]_ , \new_[23587]_ ,
    \new_[23588]_ , \new_[23589]_ , \new_[23590]_ , \new_[23591]_ ,
    \new_[23592]_ , \new_[23593]_ , \new_[23594]_ , \new_[23595]_ ,
    \new_[23596]_ , \new_[23597]_ , \new_[23598]_ , \new_[23599]_ ,
    \new_[23600]_ , \new_[23601]_ , \new_[23602]_ , \new_[23603]_ ,
    \new_[23604]_ , \new_[23605]_ , \new_[23606]_ , \new_[23607]_ ,
    \new_[23608]_ , \new_[23609]_ , \new_[23610]_ , \new_[23611]_ ,
    \new_[23612]_ , \new_[23613]_ , \new_[23614]_ , \new_[23615]_ ,
    \new_[23616]_ , \new_[23617]_ , \new_[23618]_ , \new_[23619]_ ,
    \new_[23620]_ , \new_[23621]_ , \new_[23622]_ , \new_[23623]_ ,
    \new_[23624]_ , \new_[23625]_ , \new_[23626]_ , \new_[23627]_ ,
    \new_[23628]_ , \new_[23629]_ , \new_[23630]_ , \new_[23631]_ ,
    \new_[23632]_ , \new_[23633]_ , \new_[23634]_ , \new_[23635]_ ,
    \new_[23636]_ , \new_[23637]_ , \new_[23638]_ , \new_[23639]_ ,
    \new_[23640]_ , \new_[23641]_ , \new_[23642]_ , \new_[23643]_ ,
    \new_[23644]_ , \new_[23645]_ , \new_[23646]_ , \new_[23647]_ ,
    \new_[23648]_ , \new_[23649]_ , \new_[23650]_ , \new_[23651]_ ,
    \new_[23652]_ , \new_[23653]_ , \new_[23654]_ , \new_[23655]_ ,
    \new_[23656]_ , \new_[23657]_ , \new_[23658]_ , \new_[23659]_ ,
    \new_[23660]_ , \new_[23661]_ , \new_[23662]_ , \new_[23663]_ ,
    \new_[23664]_ , \new_[23665]_ , \new_[23666]_ , \new_[23667]_ ,
    \new_[23668]_ , \new_[23669]_ , \new_[23670]_ , \new_[23671]_ ,
    \new_[23672]_ , \new_[23673]_ , \new_[23674]_ , \new_[23675]_ ,
    \new_[23676]_ , \new_[23677]_ , \new_[23678]_ , \new_[23679]_ ,
    \new_[23680]_ , \new_[23681]_ , \new_[23682]_ , \new_[23683]_ ,
    \new_[23684]_ , \new_[23685]_ , \new_[23686]_ , \new_[23687]_ ,
    \new_[23688]_ , \new_[23689]_ , \new_[23690]_ , \new_[23691]_ ,
    \new_[23692]_ , \new_[23693]_ , \new_[23694]_ , \new_[23695]_ ,
    \new_[23696]_ , \new_[23697]_ , \new_[23698]_ , \new_[23699]_ ,
    \new_[23700]_ , \new_[23701]_ , \new_[23702]_ , \new_[23703]_ ,
    \new_[23704]_ , \new_[23705]_ , \new_[23706]_ , \new_[23707]_ ,
    \new_[23708]_ , \new_[23709]_ , \new_[23710]_ , \new_[23711]_ ,
    \new_[23712]_ , \new_[23713]_ , \new_[23714]_ , \new_[23715]_ ,
    \new_[23716]_ , \new_[23717]_ , \new_[23718]_ , \new_[23719]_ ,
    \new_[23720]_ , \new_[23721]_ , \new_[23722]_ , \new_[23723]_ ,
    \new_[23724]_ , \new_[23725]_ , \new_[23726]_ , \new_[23727]_ ,
    \new_[23728]_ , \new_[23729]_ , \new_[23730]_ , \new_[23731]_ ,
    \new_[23732]_ , \new_[23733]_ , \new_[23734]_ , \new_[23735]_ ,
    \new_[23736]_ , \new_[23737]_ , \new_[23738]_ , \new_[23739]_ ,
    \new_[23740]_ , \new_[23741]_ , \new_[23742]_ , \new_[23743]_ ,
    \new_[23744]_ , \new_[23745]_ , \new_[23746]_ , \new_[23747]_ ,
    \new_[23748]_ , \new_[23749]_ , \new_[23750]_ , \new_[23751]_ ,
    \new_[23752]_ , \new_[23753]_ , \new_[23754]_ , \new_[23755]_ ,
    \new_[23756]_ , \new_[23757]_ , \new_[23758]_ , \new_[23759]_ ,
    \new_[23760]_ , \new_[23761]_ , \new_[23762]_ , \new_[23763]_ ,
    \new_[23764]_ , \new_[23765]_ , \new_[23766]_ , \new_[23767]_ ,
    \new_[23768]_ , \new_[23769]_ , \new_[23770]_ , \new_[23771]_ ,
    \new_[23772]_ , \new_[23773]_ , \new_[23774]_ , \new_[23775]_ ,
    \new_[23776]_ , \new_[23777]_ , \new_[23778]_ , \new_[23779]_ ,
    \new_[23780]_ , \new_[23781]_ , \new_[23782]_ , \new_[23783]_ ,
    \new_[23784]_ , \new_[23785]_ , \new_[23786]_ , \new_[23787]_ ,
    \new_[23788]_ , \new_[23789]_ , \new_[23790]_ , \new_[23791]_ ,
    \new_[23792]_ , \new_[23793]_ , \new_[23794]_ , \new_[23795]_ ,
    \new_[23796]_ , \new_[23797]_ , \new_[23798]_ , \new_[23799]_ ,
    \new_[23800]_ , \new_[23801]_ , \new_[23802]_ , \new_[23803]_ ,
    \new_[23804]_ , \new_[23805]_ , \new_[23806]_ , \new_[23807]_ ,
    \new_[23808]_ , \new_[23809]_ , \new_[23810]_ , \new_[23811]_ ,
    \new_[23812]_ , \new_[23813]_ , \new_[23814]_ , \new_[23815]_ ,
    \new_[23816]_ , \new_[23817]_ , \new_[23818]_ , \new_[23819]_ ,
    \new_[23820]_ , \new_[23821]_ , \new_[23822]_ , \new_[23823]_ ,
    \new_[23824]_ , \new_[23825]_ , \new_[23826]_ , \new_[23827]_ ,
    \new_[23828]_ , \new_[23829]_ , \new_[23830]_ , \new_[23831]_ ,
    \new_[23832]_ , \new_[23833]_ , \new_[23834]_ , \new_[23835]_ ,
    \new_[23836]_ , \new_[23837]_ , \new_[23838]_ , \new_[23839]_ ,
    \new_[23840]_ , \new_[23841]_ , \new_[23842]_ , \new_[23843]_ ,
    \new_[23844]_ , \new_[23845]_ , \new_[23846]_ , \new_[23847]_ ,
    \new_[23848]_ , \new_[23849]_ , \new_[23850]_ , \new_[23851]_ ,
    \new_[23852]_ , \new_[23853]_ , \new_[23854]_ , \new_[23855]_ ,
    \new_[23856]_ , \new_[23857]_ , \new_[23858]_ , \new_[23859]_ ,
    \new_[23860]_ , \new_[23861]_ , \new_[23862]_ , \new_[23863]_ ,
    \new_[23864]_ , \new_[23865]_ , \new_[23866]_ , \new_[23867]_ ,
    \new_[23868]_ , \new_[23869]_ , \new_[23870]_ , \new_[23871]_ ,
    \new_[23872]_ , \new_[23873]_ , \new_[23874]_ , \new_[23875]_ ,
    \new_[23876]_ , \new_[23877]_ , \new_[23878]_ , \new_[23879]_ ,
    \new_[23880]_ , \new_[23881]_ , \new_[23882]_ , \new_[23883]_ ,
    \new_[23884]_ , \new_[23885]_ , \new_[23886]_ , \new_[23887]_ ,
    \new_[23888]_ , \new_[23889]_ , \new_[23890]_ , \new_[23891]_ ,
    \new_[23892]_ , \new_[23893]_ , \new_[23894]_ , \new_[23895]_ ,
    \new_[23896]_ , \new_[23897]_ , \new_[23898]_ , \new_[23899]_ ,
    \new_[23900]_ , \new_[23901]_ , \new_[23902]_ , \new_[23903]_ ,
    \new_[23904]_ , \new_[23905]_ , \new_[23906]_ , \new_[23907]_ ,
    \new_[23908]_ , \new_[23909]_ , \new_[23910]_ , \new_[23911]_ ,
    \new_[23912]_ , \new_[23913]_ , \new_[23914]_ , \new_[23915]_ ,
    \new_[23916]_ , \new_[23917]_ , \new_[23918]_ , \new_[23919]_ ,
    \new_[23920]_ , \new_[23921]_ , \new_[23922]_ , \new_[23923]_ ,
    \new_[23924]_ , \new_[23925]_ , \new_[23926]_ , \new_[23927]_ ,
    \new_[23928]_ , \new_[23929]_ , \new_[23930]_ , \new_[23931]_ ,
    \new_[23932]_ , \new_[23933]_ , \new_[23934]_ , \new_[23935]_ ,
    \new_[23936]_ , \new_[23937]_ , \new_[23938]_ , \new_[23939]_ ,
    \new_[23940]_ , \new_[23941]_ , \new_[23942]_ , \new_[23943]_ ,
    \new_[23944]_ , \new_[23945]_ , \new_[23946]_ , \new_[23947]_ ,
    \new_[23948]_ , \new_[23949]_ , \new_[23950]_ , \new_[23951]_ ,
    \new_[23952]_ , \new_[23953]_ , \new_[23954]_ , \new_[23955]_ ,
    \new_[23956]_ , \new_[23957]_ , \new_[23958]_ , \new_[23959]_ ,
    \new_[23960]_ , \new_[23961]_ , \new_[23962]_ , \new_[23963]_ ,
    \new_[23964]_ , \new_[23965]_ , \new_[23966]_ , \new_[23967]_ ,
    \new_[23968]_ , \new_[23969]_ , \new_[23970]_ , \new_[23971]_ ,
    \new_[23972]_ , \new_[23973]_ , \new_[23974]_ , \new_[23975]_ ,
    \new_[23976]_ , \new_[23977]_ , \new_[23978]_ , \new_[23979]_ ,
    \new_[23980]_ , \new_[23981]_ , \new_[23982]_ , \new_[23983]_ ,
    \new_[23984]_ , \new_[23985]_ , \new_[23986]_ , \new_[23987]_ ,
    \new_[23988]_ , \new_[23989]_ , \new_[23990]_ , \new_[23991]_ ,
    \new_[23992]_ , \new_[23993]_ , \new_[23994]_ , \new_[23995]_ ,
    \new_[23996]_ , \new_[23997]_ , \new_[23998]_ , \new_[23999]_ ,
    \new_[24000]_ , \new_[24001]_ , \new_[24002]_ , \new_[24003]_ ,
    \new_[24004]_ , \new_[24005]_ , \new_[24006]_ , \new_[24007]_ ,
    \new_[24008]_ , \new_[24009]_ , \new_[24010]_ , \new_[24011]_ ,
    \new_[24012]_ , \new_[24013]_ , \new_[24014]_ , \new_[24015]_ ,
    \new_[24016]_ , \new_[24017]_ , \new_[24018]_ , \new_[24019]_ ,
    \new_[24020]_ , \new_[24021]_ , \new_[24022]_ , \new_[24023]_ ,
    \new_[24024]_ , \new_[24025]_ , \new_[24026]_ , \new_[24027]_ ,
    \new_[24028]_ , \new_[24029]_ , \new_[24030]_ , \new_[24031]_ ,
    \new_[24032]_ , \new_[24033]_ , \new_[24034]_ , \new_[24035]_ ,
    \new_[24036]_ , \new_[24037]_ , \new_[24038]_ , \new_[24039]_ ,
    \new_[24040]_ , \new_[24041]_ , \new_[24042]_ , \new_[24043]_ ,
    \new_[24044]_ , \new_[24045]_ , \new_[24046]_ , \new_[24047]_ ,
    \new_[24048]_ , \new_[24049]_ , \new_[24050]_ , \new_[24051]_ ,
    \new_[24052]_ , \new_[24053]_ , \new_[24054]_ , \new_[24055]_ ,
    \new_[24056]_ , \new_[24057]_ , \new_[24058]_ , \new_[24059]_ ,
    \new_[24060]_ , \new_[24061]_ , \new_[24062]_ , \new_[24063]_ ,
    \new_[24064]_ , \new_[24065]_ , \new_[24066]_ , \new_[24067]_ ,
    \new_[24068]_ , \new_[24069]_ , \new_[24070]_ , \new_[24071]_ ,
    \new_[24072]_ , \new_[24073]_ , \new_[24074]_ , \new_[24075]_ ,
    \new_[24076]_ , \new_[24077]_ , \new_[24078]_ , \new_[24079]_ ,
    \new_[24080]_ , \new_[24081]_ , \new_[24082]_ , \new_[24083]_ ,
    \new_[24084]_ , \new_[24085]_ , \new_[24086]_ , \new_[24087]_ ,
    \new_[24088]_ , \new_[24089]_ , \new_[24090]_ , \new_[24091]_ ,
    \new_[24092]_ , \new_[24093]_ , \new_[24094]_ , \new_[24095]_ ,
    \new_[24096]_ , \new_[24097]_ , \new_[24098]_ , \new_[24099]_ ,
    \new_[24100]_ , \new_[24101]_ , \new_[24102]_ , \new_[24103]_ ,
    \new_[24104]_ , \new_[24105]_ , \new_[24106]_ , \new_[24107]_ ,
    \new_[24108]_ , \new_[24109]_ , \new_[24110]_ , \new_[24111]_ ,
    \new_[24112]_ , \new_[24113]_ , \new_[24114]_ , \new_[24115]_ ,
    \new_[24116]_ , \new_[24117]_ , \new_[24118]_ , \new_[24119]_ ,
    \new_[24120]_ , \new_[24121]_ , \new_[24122]_ , \new_[24123]_ ,
    \new_[24124]_ , \new_[24125]_ , \new_[24126]_ , \new_[24127]_ ,
    \new_[24128]_ , \new_[24129]_ , \new_[24130]_ , \new_[24131]_ ,
    \new_[24132]_ , \new_[24133]_ , \new_[24134]_ , \new_[24135]_ ,
    \new_[24136]_ , \new_[24137]_ , \new_[24138]_ , \new_[24139]_ ,
    \new_[24140]_ , \new_[24141]_ , \new_[24142]_ , \new_[24143]_ ,
    \new_[24144]_ , \new_[24145]_ , \new_[24146]_ , \new_[24147]_ ,
    \new_[24148]_ , \new_[24149]_ , \new_[24150]_ , \new_[24151]_ ,
    \new_[24152]_ , \new_[24153]_ , \new_[24154]_ , \new_[24155]_ ,
    \new_[24156]_ , \new_[24157]_ , \new_[24158]_ , \new_[24159]_ ,
    \new_[24160]_ , \new_[24161]_ , \new_[24162]_ , \new_[24163]_ ,
    \new_[24164]_ , \new_[24165]_ , \new_[24166]_ , \new_[24167]_ ,
    \new_[24168]_ , \new_[24169]_ , \new_[24170]_ , \new_[24171]_ ,
    \new_[24172]_ , \new_[24173]_ , \new_[24174]_ , \new_[24175]_ ,
    \new_[24176]_ , \new_[24177]_ , \new_[24178]_ , \new_[24179]_ ,
    \new_[24180]_ , \new_[24181]_ , \new_[24182]_ , \new_[24183]_ ,
    \new_[24184]_ , \new_[24185]_ , \new_[24186]_ , \new_[24187]_ ,
    \new_[24188]_ , \new_[24189]_ , \new_[24190]_ , \new_[24191]_ ,
    \new_[24192]_ , \new_[24193]_ , \new_[24194]_ , \new_[24195]_ ,
    \new_[24196]_ , \new_[24197]_ , \new_[24198]_ , \new_[24199]_ ,
    \new_[24200]_ , \new_[24201]_ , \new_[24202]_ , \new_[24203]_ ,
    \new_[24204]_ , \new_[24205]_ , \new_[24206]_ , \new_[24207]_ ,
    \new_[24208]_ , \new_[24209]_ , \new_[24210]_ , \new_[24211]_ ,
    \new_[24212]_ , \new_[24213]_ , \new_[24214]_ , \new_[24215]_ ,
    \new_[24216]_ , \new_[24217]_ , \new_[24218]_ , \new_[24219]_ ,
    \new_[24220]_ , \new_[24221]_ , \new_[24222]_ , \new_[24223]_ ,
    \new_[24224]_ , \new_[24225]_ , \new_[24226]_ , \new_[24227]_ ,
    \new_[24228]_ , \new_[24229]_ , \new_[24230]_ , \new_[24231]_ ,
    \new_[24232]_ , \new_[24233]_ , \new_[24234]_ , \new_[24235]_ ,
    \new_[24236]_ , \new_[24237]_ , \new_[24238]_ , \new_[24239]_ ,
    \new_[24240]_ , \new_[24241]_ , \new_[24242]_ , \new_[24243]_ ,
    \new_[24244]_ , \new_[24245]_ , \new_[24246]_ , \new_[24247]_ ,
    \new_[24248]_ , \new_[24249]_ , \new_[24250]_ , \new_[24251]_ ,
    \new_[24252]_ , \new_[24253]_ , \new_[24254]_ , \new_[24255]_ ,
    \new_[24256]_ , \new_[24257]_ , \new_[24258]_ , \new_[24259]_ ,
    \new_[24260]_ , \new_[24261]_ , \new_[24262]_ , \new_[24263]_ ,
    \new_[24264]_ , \new_[24265]_ , \new_[24266]_ , \new_[24267]_ ,
    \new_[24268]_ , \new_[24269]_ , \new_[24270]_ , \new_[24271]_ ,
    \new_[24272]_ , \new_[24273]_ , \new_[24274]_ , \new_[24275]_ ,
    \new_[24276]_ , \new_[24277]_ , \new_[24278]_ , \new_[24279]_ ,
    \new_[24280]_ , \new_[24281]_ , \new_[24282]_ , \new_[24283]_ ,
    \new_[24284]_ , \new_[24285]_ , \new_[24286]_ , \new_[24287]_ ,
    \new_[24288]_ , \new_[24289]_ , \new_[24290]_ , \new_[24291]_ ,
    \new_[24292]_ , \new_[24293]_ , \new_[24294]_ , \new_[24295]_ ,
    \new_[24296]_ , \new_[24297]_ , \new_[24298]_ , \new_[24299]_ ,
    \new_[24300]_ , \new_[24301]_ , \new_[24302]_ , \new_[24303]_ ,
    \new_[24304]_ , \new_[24305]_ , \new_[24306]_ , \new_[24307]_ ,
    \new_[24308]_ , \new_[24309]_ , \new_[24310]_ , \new_[24311]_ ,
    \new_[24312]_ , \new_[24313]_ , \new_[24314]_ , \new_[24315]_ ,
    \new_[24316]_ , \new_[24317]_ , \new_[24318]_ , \new_[24319]_ ,
    \new_[24320]_ , \new_[24321]_ , \new_[24322]_ , \new_[24323]_ ,
    \new_[24324]_ , \new_[24325]_ , \new_[24326]_ , \new_[24327]_ ,
    \new_[24328]_ , \new_[24329]_ , \new_[24330]_ , \new_[24331]_ ,
    \new_[24332]_ , \new_[24333]_ , \new_[24334]_ , \new_[24335]_ ,
    \new_[24336]_ , \new_[24337]_ , \new_[24338]_ , \new_[24339]_ ,
    \new_[24340]_ , \new_[24341]_ , \new_[24342]_ , \new_[24343]_ ,
    \new_[24344]_ , \new_[24345]_ , \new_[24346]_ , \new_[24347]_ ,
    \new_[24348]_ , \new_[24349]_ , \new_[24350]_ , \new_[24351]_ ,
    \new_[24352]_ , \new_[24353]_ , \new_[24354]_ , \new_[24355]_ ,
    \new_[24356]_ , \new_[24357]_ , \new_[24358]_ , \new_[24359]_ ,
    \new_[24360]_ , \new_[24361]_ , \new_[24362]_ , \new_[24363]_ ,
    \new_[24364]_ , \new_[24365]_ , \new_[24366]_ , \new_[24367]_ ,
    \new_[24368]_ , \new_[24369]_ , \new_[24370]_ , \new_[24371]_ ,
    \new_[24372]_ , \new_[24373]_ , \new_[24374]_ , \new_[24375]_ ,
    \new_[24376]_ , \new_[24377]_ , \new_[24378]_ , \new_[24379]_ ,
    \new_[24380]_ , \new_[24381]_ , \new_[24382]_ , \new_[24383]_ ,
    \new_[24384]_ , \new_[24385]_ , \new_[24386]_ , \new_[24387]_ ,
    \new_[24388]_ , \new_[24389]_ , \new_[24390]_ , \new_[24391]_ ,
    \new_[24392]_ , \new_[24393]_ , \new_[24394]_ , \new_[24395]_ ,
    \new_[24396]_ , \new_[24397]_ , \new_[24398]_ , \new_[24399]_ ,
    \new_[24400]_ , \new_[24401]_ , \new_[24402]_ , \new_[24403]_ ,
    \new_[24404]_ , \new_[24405]_ , \new_[24406]_ , \new_[24407]_ ,
    \new_[24408]_ , \new_[24409]_ , \new_[24410]_ , \new_[24411]_ ,
    \new_[24412]_ , \new_[24413]_ , \new_[24414]_ , \new_[24415]_ ,
    \new_[24416]_ , \new_[24417]_ , \new_[24418]_ , \new_[24419]_ ,
    \new_[24420]_ , \new_[24421]_ , \new_[24422]_ , \new_[24423]_ ,
    \new_[24424]_ , \new_[24425]_ , \new_[24426]_ , \new_[24427]_ ,
    \new_[24428]_ , \new_[24429]_ , \new_[24430]_ , \new_[24431]_ ,
    \new_[24432]_ , \new_[24433]_ , \new_[24434]_ , \new_[24435]_ ,
    \new_[24436]_ , \new_[24437]_ , \new_[24438]_ , \new_[24439]_ ,
    \new_[24440]_ , \new_[24441]_ , \new_[24442]_ , \new_[24443]_ ,
    \new_[24444]_ , \new_[24445]_ , \new_[24446]_ , \new_[24447]_ ,
    \new_[24448]_ , \new_[24449]_ , \new_[24450]_ , \new_[24451]_ ,
    \new_[24452]_ , \new_[24453]_ , \new_[24454]_ , \new_[24455]_ ,
    \new_[24456]_ , \new_[24457]_ , \new_[24458]_ , \new_[24459]_ ,
    \new_[24460]_ , \new_[24461]_ , \new_[24462]_ , \new_[24463]_ ,
    \new_[24464]_ , \new_[24465]_ , \new_[24466]_ , \new_[24467]_ ,
    \new_[24468]_ , \new_[24469]_ , \new_[24470]_ , \new_[24471]_ ,
    \new_[24472]_ , \new_[24473]_ , \new_[24474]_ , \new_[24475]_ ,
    \new_[24476]_ , \new_[24477]_ , \new_[24478]_ , \new_[24479]_ ,
    \new_[24480]_ , \new_[24481]_ , \new_[24482]_ , \new_[24483]_ ,
    \new_[24484]_ , \new_[24485]_ , \new_[24486]_ , \new_[24487]_ ,
    \new_[24488]_ , \new_[24489]_ , \new_[24490]_ , \new_[24491]_ ,
    \new_[24492]_ , \new_[24493]_ , \new_[24494]_ , \new_[24495]_ ,
    \new_[24496]_ , \new_[24497]_ , \new_[24498]_ , \new_[24499]_ ,
    \new_[24500]_ , \new_[24501]_ , \new_[24502]_ , \new_[24503]_ ,
    \new_[24504]_ , \new_[24505]_ , \new_[24506]_ , \new_[24507]_ ,
    \new_[24508]_ , \new_[24509]_ , \new_[24510]_ , \new_[24511]_ ,
    \new_[24512]_ , \new_[24513]_ , \new_[24514]_ , \new_[24515]_ ,
    \new_[24516]_ , \new_[24517]_ , \new_[24518]_ , \new_[24519]_ ,
    \new_[24520]_ , \new_[24521]_ , \new_[24522]_ , \new_[24523]_ ,
    \new_[24524]_ , \new_[24525]_ , \new_[24526]_ , \new_[24527]_ ,
    \new_[24528]_ , \new_[24529]_ , \new_[24530]_ , \new_[24531]_ ,
    \new_[24532]_ , \new_[24533]_ , \new_[24534]_ , \new_[24535]_ ,
    \new_[24536]_ , \new_[24537]_ , \new_[24538]_ , \new_[24539]_ ,
    \new_[24540]_ , \new_[24541]_ , \new_[24542]_ , \new_[24543]_ ,
    \new_[24544]_ , \new_[24545]_ , \new_[24546]_ , \new_[24547]_ ,
    \new_[24548]_ , \new_[24549]_ , \new_[24550]_ , \new_[24551]_ ,
    \new_[24552]_ , \new_[24553]_ , \new_[24554]_ , \new_[24555]_ ,
    \new_[24556]_ , \new_[24557]_ , \new_[24558]_ , \new_[24559]_ ,
    \new_[24560]_ , \new_[24561]_ , \new_[24562]_ , \new_[24563]_ ,
    \new_[24564]_ , \new_[24565]_ , \new_[24566]_ , \new_[24567]_ ,
    \new_[24568]_ , \new_[24569]_ , \new_[24570]_ , \new_[24571]_ ,
    \new_[24572]_ , \new_[24573]_ , \new_[24574]_ , \new_[24575]_ ,
    \new_[24576]_ , \new_[24577]_ , \new_[24578]_ , \new_[24579]_ ,
    \new_[24580]_ , \new_[24581]_ , \new_[24582]_ , \new_[24583]_ ,
    \new_[24584]_ , \new_[24585]_ , \new_[24586]_ , \new_[24587]_ ,
    \new_[24588]_ , \new_[24589]_ , \new_[24590]_ , \new_[24591]_ ,
    \new_[24592]_ , \new_[24593]_ , \new_[24594]_ , \new_[24595]_ ,
    \new_[24596]_ , \new_[24597]_ , \new_[24598]_ , \new_[24599]_ ,
    \new_[24600]_ , \new_[24601]_ , \new_[24602]_ , \new_[24603]_ ,
    \new_[24604]_ , \new_[24605]_ , \new_[24606]_ , \new_[24607]_ ,
    \new_[24608]_ , \new_[24609]_ , \new_[24610]_ , \new_[24611]_ ,
    \new_[24612]_ , \new_[24613]_ , \new_[24614]_ , \new_[24615]_ ,
    \new_[24616]_ , \new_[24617]_ , \new_[24618]_ , \new_[24619]_ ,
    \new_[24620]_ , \new_[24621]_ , \new_[24622]_ , \new_[24623]_ ,
    \new_[24624]_ , \new_[24625]_ , \new_[24626]_ , \new_[24627]_ ,
    \new_[24628]_ , \new_[24629]_ , \new_[24630]_ , \new_[24631]_ ,
    \new_[24632]_ , \new_[24633]_ , \new_[24634]_ , \new_[24635]_ ,
    \new_[24636]_ , \new_[24637]_ , \new_[24638]_ , \new_[24639]_ ,
    \new_[24640]_ , \new_[24641]_ , \new_[24642]_ , \new_[24643]_ ,
    \new_[24644]_ , \new_[24645]_ , \new_[24646]_ , \new_[24647]_ ,
    \new_[24648]_ , \new_[24649]_ , \new_[24650]_ , \new_[24651]_ ,
    \new_[24652]_ , \new_[24653]_ , \new_[24654]_ , \new_[24655]_ ,
    \new_[24656]_ , \new_[24657]_ , \new_[24658]_ , \new_[24659]_ ,
    \new_[24660]_ , \new_[24661]_ , \new_[24662]_ , \new_[24663]_ ,
    \new_[24664]_ , \new_[24665]_ , \new_[24666]_ , \new_[24667]_ ,
    \new_[24668]_ , \new_[24669]_ , \new_[24670]_ , \new_[24671]_ ,
    \new_[24672]_ , \new_[24673]_ , \new_[24674]_ , \new_[24675]_ ,
    \new_[24676]_ , \new_[24677]_ , \new_[24678]_ , \new_[24679]_ ,
    \new_[24680]_ , \new_[24681]_ , \new_[24682]_ , \new_[24683]_ ,
    \new_[24684]_ , \new_[24685]_ , \new_[24686]_ , \new_[24687]_ ,
    \new_[24688]_ , \new_[24689]_ , \new_[24690]_ , \new_[24691]_ ,
    \new_[24692]_ , \new_[24693]_ , \new_[24694]_ , \new_[24695]_ ,
    \new_[24696]_ , \new_[24697]_ , \new_[24699]_ , \new_[24700]_ ,
    \new_[24701]_ , \new_[24702]_ , \new_[24703]_ , \new_[24704]_ ,
    \new_[24705]_ , \new_[24706]_ , \new_[24707]_ , \new_[24708]_ ,
    \new_[24709]_ , \new_[24710]_ , \new_[24711]_ , \new_[24712]_ ,
    \new_[24713]_ , \new_[24714]_ , \new_[24715]_ , \new_[24716]_ ,
    \new_[24717]_ , \new_[24718]_ , \new_[24719]_ , \new_[24720]_ ,
    \new_[24721]_ , \new_[24722]_ , \new_[24723]_ , \new_[24724]_ ,
    \new_[24725]_ , \new_[24726]_ , \new_[24727]_ , \new_[24728]_ ,
    \new_[24729]_ , \new_[24730]_ , \new_[24731]_ , \new_[24732]_ ,
    \new_[24733]_ , \new_[24734]_ , \new_[24735]_ , \new_[24736]_ ,
    \new_[24737]_ , \new_[24738]_ , \new_[24739]_ , \new_[24740]_ ,
    \new_[24741]_ , \new_[24742]_ , \new_[24743]_ , \new_[24744]_ ,
    \new_[24745]_ , \new_[24746]_ , \new_[24747]_ , \new_[24748]_ ,
    \new_[24749]_ , \new_[24750]_ , \new_[24751]_ , \new_[24752]_ ,
    \new_[24753]_ , \new_[24754]_ , \new_[24755]_ , \new_[24756]_ ,
    \new_[24757]_ , \new_[24758]_ , \new_[24759]_ , \new_[24760]_ ,
    \new_[24761]_ , \new_[24762]_ , \new_[24763]_ , \new_[24764]_ ,
    \new_[24765]_ , \new_[24766]_ , \new_[24767]_ , \new_[24768]_ ,
    \new_[24769]_ , \new_[24770]_ , \new_[24771]_ , \new_[24772]_ ,
    \new_[24773]_ , \new_[24774]_ , \new_[24775]_ , \new_[24776]_ ,
    \new_[24777]_ , \new_[24778]_ , \new_[24779]_ , \new_[24780]_ ,
    \new_[24782]_ , \new_[24783]_ , \new_[24785]_ , \new_[24787]_ ,
    \new_[24788]_ , \new_[24790]_ , \new_[24791]_ , \new_[24792]_ ,
    \new_[24793]_ , \new_[24794]_ , \new_[24795]_ , \new_[24796]_ ,
    \new_[24797]_ , \new_[24798]_ , \new_[24799]_ , \new_[24800]_ ,
    \new_[24801]_ , \new_[24802]_ , \new_[24803]_ , \new_[24804]_ ,
    \new_[24805]_ , \new_[24806]_ , \new_[24807]_ , \new_[24808]_ ,
    \new_[24809]_ , \new_[24810]_ , \new_[24811]_ , \new_[24812]_ ,
    \new_[24813]_ , \new_[24814]_ , \new_[24815]_ , \new_[24816]_ ,
    \new_[24817]_ , \new_[24818]_ , \new_[24819]_ , \new_[24820]_ ,
    \new_[24821]_ , \new_[24822]_ , \new_[24823]_ , \new_[24824]_ ,
    \new_[24825]_ , \new_[24826]_ , \new_[24827]_ , \new_[24828]_ ,
    \new_[24829]_ , \new_[24830]_ , \new_[24831]_ , \new_[24832]_ ,
    \new_[24833]_ , \new_[24834]_ , \new_[24835]_ , \new_[24836]_ ,
    \new_[24837]_ , \new_[24838]_ , \new_[24839]_ , \new_[24840]_ ,
    \new_[24841]_ , \new_[24842]_ , \new_[24843]_ , \new_[24844]_ ,
    \new_[24845]_ , \new_[24846]_ , \new_[24847]_ , \new_[24848]_ ,
    \new_[24849]_ , \new_[24850]_ , \new_[24851]_ , \new_[24852]_ ,
    \new_[24853]_ , \new_[24854]_ , \new_[24855]_ , \new_[24856]_ ,
    \new_[24857]_ , \new_[24858]_ , \new_[24859]_ , \new_[24860]_ ,
    \new_[24861]_ , \new_[24862]_ , \new_[24863]_ , \new_[24864]_ ,
    \new_[24865]_ , \new_[24866]_ , \new_[24867]_ , \new_[24868]_ ,
    \new_[24869]_ , \new_[24870]_ , \new_[24871]_ , \new_[24872]_ ,
    \new_[24873]_ , \new_[24874]_ , \new_[24875]_ , \new_[24876]_ ,
    \new_[24877]_ , \new_[24878]_ , \new_[24879]_ , \new_[24880]_ ,
    \new_[24881]_ , \new_[24882]_ , \new_[24883]_ , \new_[24884]_ ,
    \new_[24885]_ , \new_[24886]_ , \new_[24887]_ , \new_[24888]_ ,
    \new_[24889]_ , \new_[24890]_ , \new_[24891]_ , \new_[24892]_ ,
    \new_[24893]_ , \new_[24894]_ , \new_[24895]_ , \new_[24896]_ ,
    \new_[24897]_ , \new_[24898]_ , \new_[24899]_ , \new_[24900]_ ,
    \new_[24901]_ , \new_[24902]_ , \new_[24903]_ , \new_[24904]_ ,
    \new_[24905]_ , \new_[24906]_ , \new_[24907]_ , \new_[24908]_ ,
    \new_[24909]_ , \new_[24910]_ , \new_[24911]_ , \new_[24912]_ ,
    \new_[24913]_ , \new_[24914]_ , \new_[24915]_ , \new_[24916]_ ,
    \new_[24917]_ , \new_[24918]_ , \new_[24919]_ , \new_[24920]_ ,
    \new_[24921]_ , \new_[24922]_ , \new_[24923]_ , \new_[24924]_ ,
    \new_[24925]_ , \new_[24926]_ , \new_[24927]_ , \new_[24928]_ ,
    \new_[24929]_ , \new_[24930]_ , \new_[24931]_ , \new_[24932]_ ,
    \new_[24933]_ , \new_[24934]_ , \new_[24935]_ , \new_[24936]_ ,
    \new_[24937]_ , \new_[24938]_ , \new_[24939]_ , \new_[24940]_ ,
    \new_[24941]_ , \new_[24942]_ , \new_[24943]_ , \new_[24944]_ ,
    \new_[24945]_ , \new_[24946]_ , \new_[24947]_ , \new_[24948]_ ,
    \new_[24949]_ , \new_[24950]_ , \new_[24951]_ , \new_[24952]_ ,
    \new_[24953]_ , \new_[24954]_ , \new_[24955]_ , \new_[24956]_ ,
    \new_[24957]_ , \new_[24958]_ , \new_[24959]_ , \new_[24960]_ ,
    \new_[24961]_ , \new_[24962]_ , \new_[24963]_ , \new_[24964]_ ,
    \new_[24965]_ , \new_[24966]_ , \new_[24967]_ , \new_[24968]_ ,
    \new_[24969]_ , \new_[24970]_ , \new_[24971]_ , \new_[24972]_ ,
    \new_[24973]_ , \new_[24974]_ , \new_[24975]_ , \new_[24976]_ ,
    \new_[24977]_ , \new_[24978]_ , \new_[24979]_ , \new_[24980]_ ,
    \new_[24981]_ , \new_[24982]_ , \new_[24983]_ , \new_[24984]_ ,
    \new_[24985]_ , \new_[24986]_ , \new_[24987]_ , \new_[24988]_ ,
    \new_[24989]_ , \new_[24990]_ , \new_[24991]_ , \new_[24992]_ ,
    \new_[24993]_ , \new_[24994]_ , \new_[24995]_ , \new_[24996]_ ,
    \new_[24997]_ , \new_[24998]_ , \new_[24999]_ , \new_[25000]_ ,
    \new_[25001]_ , \new_[25002]_ , \new_[25003]_ , \new_[25004]_ ,
    \new_[25005]_ , \new_[25006]_ , \new_[25007]_ , \new_[25008]_ ,
    \new_[25009]_ , \new_[25010]_ , \new_[25011]_ , \new_[25012]_ ,
    \new_[25013]_ , \new_[25014]_ , \new_[25015]_ , \new_[25016]_ ,
    \new_[25017]_ , \new_[25018]_ , \new_[25019]_ , \new_[25020]_ ,
    \new_[25021]_ , \new_[25022]_ , \new_[25023]_ , \new_[25024]_ ,
    \new_[25025]_ , \new_[25026]_ , \new_[25027]_ , \new_[25028]_ ,
    \new_[25029]_ , \new_[25030]_ , \new_[25031]_ , \new_[25032]_ ,
    \new_[25033]_ , \new_[25034]_ , \new_[25035]_ , \new_[25036]_ ,
    \new_[25037]_ , \new_[25038]_ , \new_[25039]_ , \new_[25040]_ ,
    \new_[25041]_ , \new_[25042]_ , \new_[25043]_ , \new_[25044]_ ,
    \new_[25045]_ , \new_[25046]_ , \new_[25047]_ , \new_[25048]_ ,
    \new_[25049]_ , \new_[25050]_ , \new_[25051]_ , \new_[25052]_ ,
    \new_[25053]_ , \new_[25054]_ , \new_[25055]_ , \new_[25056]_ ,
    \new_[25057]_ , \new_[25058]_ , \new_[25059]_ , \new_[25060]_ ,
    \new_[25061]_ , \new_[25062]_ , \new_[25063]_ , \new_[25064]_ ,
    \new_[25065]_ , \new_[25066]_ , \new_[25067]_ , \new_[25068]_ ,
    \new_[25069]_ , \new_[25070]_ , \new_[25071]_ , \new_[25072]_ ,
    \new_[25073]_ , \new_[25074]_ , \new_[25075]_ , \new_[25076]_ ,
    \new_[25077]_ , \new_[25078]_ , \new_[25079]_ , \new_[25080]_ ,
    \new_[25081]_ , \new_[25082]_ , \new_[25083]_ , \new_[25084]_ ,
    \new_[25085]_ , \new_[25086]_ , \new_[25087]_ , \new_[25088]_ ,
    \new_[25089]_ , \new_[25090]_ , \new_[25091]_ , \new_[25092]_ ,
    \new_[25093]_ , \new_[25094]_ , \new_[25095]_ , \new_[25096]_ ,
    \new_[25097]_ , \new_[25098]_ , \new_[25099]_ , \new_[25100]_ ,
    \new_[25101]_ , \new_[25102]_ , \new_[25103]_ , \new_[25104]_ ,
    \new_[25105]_ , \new_[25106]_ , \new_[25107]_ , \new_[25108]_ ,
    \new_[25109]_ , \new_[25110]_ , \new_[25111]_ , \new_[25112]_ ,
    \new_[25113]_ , \new_[25114]_ , \new_[25115]_ , \new_[25116]_ ,
    \new_[25117]_ , \new_[25118]_ , \new_[25119]_ , \new_[25120]_ ,
    \new_[25121]_ , \new_[25122]_ , \new_[25123]_ , \new_[25124]_ ,
    \new_[25125]_ , \new_[25126]_ , \new_[25127]_ , \new_[25128]_ ,
    \new_[25129]_ , \new_[25130]_ , \new_[25131]_ , \new_[25132]_ ,
    \new_[25133]_ , \new_[25134]_ , \new_[25135]_ , \new_[25136]_ ,
    \new_[25137]_ , \new_[25138]_ , \new_[25139]_ , \new_[25140]_ ,
    \new_[25141]_ , \new_[25142]_ , \new_[25143]_ , \new_[25144]_ ,
    \new_[25145]_ , \new_[25146]_ , \new_[25147]_ , \new_[25148]_ ,
    \new_[25149]_ , \new_[25150]_ , \new_[25151]_ , \new_[25152]_ ,
    \new_[25153]_ , \new_[25154]_ , \new_[25155]_ , \new_[25156]_ ,
    \new_[25157]_ , \new_[25158]_ , \new_[25159]_ , \new_[25160]_ ,
    \new_[25161]_ , \new_[25162]_ , \new_[25163]_ , \new_[25164]_ ,
    \new_[25165]_ , \new_[25166]_ , \new_[25167]_ , \new_[25168]_ ,
    \new_[25169]_ , \new_[25170]_ , \new_[25171]_ , \new_[25172]_ ,
    \new_[25173]_ , \new_[25174]_ , \new_[25175]_ , \new_[25176]_ ,
    \new_[25177]_ , \new_[25178]_ , \new_[25179]_ , \new_[25180]_ ,
    \new_[25181]_ , \new_[25182]_ , \new_[25183]_ , \new_[25184]_ ,
    \new_[25185]_ , \new_[25186]_ , \new_[25187]_ , \new_[25188]_ ,
    \new_[25189]_ , \new_[25190]_ , \new_[25191]_ , \new_[25192]_ ,
    \new_[25193]_ , \new_[25194]_ , \new_[25195]_ , \new_[25196]_ ,
    \new_[25197]_ , \new_[25198]_ , \new_[25199]_ , \new_[25200]_ ,
    \new_[25201]_ , \new_[25202]_ , \new_[25203]_ , \new_[25204]_ ,
    \new_[25205]_ , \new_[25206]_ , \new_[25207]_ , \new_[25208]_ ,
    \new_[25209]_ , \new_[25210]_ , \new_[25211]_ , \new_[25212]_ ,
    \new_[25213]_ , \new_[25214]_ , \new_[25215]_ , \new_[25216]_ ,
    \new_[25217]_ , \new_[25218]_ , \new_[25219]_ , \new_[25220]_ ,
    \new_[25221]_ , \new_[25222]_ , \new_[25223]_ , \new_[25224]_ ,
    \new_[25225]_ , \new_[25226]_ , \new_[25227]_ , \new_[25228]_ ,
    \new_[25229]_ , \new_[25230]_ , \new_[25231]_ , \new_[25232]_ ,
    \new_[25233]_ , \new_[25234]_ , \new_[25235]_ , \new_[25236]_ ,
    \new_[25237]_ , \new_[25238]_ , \new_[25239]_ , \new_[25240]_ ,
    \new_[25241]_ , \new_[25242]_ , \new_[25243]_ , \new_[25244]_ ,
    \new_[25245]_ , \new_[25246]_ , \new_[25247]_ , \new_[25248]_ ,
    \new_[25249]_ , \new_[25250]_ , \new_[25251]_ , \new_[25252]_ ,
    \new_[25253]_ , \new_[25254]_ , \new_[25255]_ , \new_[25256]_ ,
    \new_[25257]_ , \new_[25258]_ , \new_[25259]_ , \new_[25260]_ ,
    \new_[25261]_ , \new_[25262]_ , \new_[25263]_ , \new_[25264]_ ,
    \new_[25265]_ , \new_[25266]_ , \new_[25267]_ , \new_[25268]_ ,
    \new_[25269]_ , \new_[25270]_ , \new_[25271]_ , \new_[25272]_ ,
    \new_[25273]_ , \new_[25274]_ , \new_[25275]_ , \new_[25276]_ ,
    \new_[25277]_ , \new_[25278]_ , \new_[25279]_ , \new_[25280]_ ,
    \new_[25281]_ , \new_[25282]_ , \new_[25283]_ , \new_[25284]_ ,
    \new_[25285]_ , \new_[25286]_ , \new_[25287]_ , \new_[25288]_ ,
    \new_[25289]_ , \new_[25290]_ , \new_[25291]_ , \new_[25292]_ ,
    \new_[25293]_ , \new_[25294]_ , \new_[25295]_ , \new_[25296]_ ,
    \new_[25297]_ , \new_[25298]_ , \new_[25299]_ , \new_[25300]_ ,
    \new_[25301]_ , \new_[25302]_ , \new_[25303]_ , \new_[25304]_ ,
    \new_[25305]_ , \new_[25306]_ , \new_[25307]_ , \new_[25308]_ ,
    \new_[25309]_ , \new_[25310]_ , \new_[25311]_ , \new_[25312]_ ,
    \new_[25313]_ , \new_[25314]_ , \new_[25315]_ , \new_[25316]_ ,
    \new_[25317]_ , \new_[25318]_ , \new_[25319]_ , \new_[25320]_ ,
    \new_[25321]_ , \new_[25322]_ , \new_[25323]_ , \new_[25324]_ ,
    \new_[25325]_ , \new_[25326]_ , \new_[25327]_ , \new_[25328]_ ,
    \new_[25329]_ , \new_[25330]_ , \new_[25331]_ , \new_[25332]_ ,
    \new_[25333]_ , \new_[25334]_ , \new_[25335]_ , \new_[25336]_ ,
    \new_[25337]_ , \new_[25338]_ , \new_[25339]_ , \new_[25340]_ ,
    \new_[25341]_ , \new_[25342]_ , \new_[25343]_ , \new_[25344]_ ,
    \new_[25345]_ , \new_[25346]_ , \new_[25347]_ , \new_[25348]_ ,
    \new_[25349]_ , \new_[25350]_ , \new_[25351]_ , \new_[25352]_ ,
    \new_[25353]_ , \new_[25354]_ , \new_[25355]_ , \new_[25356]_ ,
    \new_[25357]_ , \new_[25358]_ , \new_[25359]_ , \new_[25360]_ ,
    \new_[25361]_ , \new_[25362]_ , \new_[25363]_ , \new_[25364]_ ,
    \new_[25365]_ , \new_[25366]_ , \new_[25367]_ , \new_[25368]_ ,
    \new_[25369]_ , \new_[25370]_ , \new_[25371]_ , \new_[25372]_ ,
    \new_[25373]_ , \new_[25374]_ , \new_[25375]_ , \new_[25376]_ ,
    \new_[25377]_ , \new_[25378]_ , \new_[25379]_ , \new_[25380]_ ,
    \new_[25381]_ , \new_[25382]_ , \new_[25383]_ , \new_[25384]_ ,
    \new_[25385]_ , \new_[25386]_ , \new_[25387]_ , \new_[25388]_ ,
    \new_[25389]_ , \new_[25390]_ , \new_[25391]_ , \new_[25392]_ ,
    \new_[25393]_ , \new_[25394]_ , \new_[25395]_ , \new_[25396]_ ,
    \new_[25397]_ , \new_[25398]_ , \new_[25399]_ , \new_[25400]_ ,
    \new_[25401]_ , \new_[25402]_ , \new_[25403]_ , \new_[25404]_ ,
    \new_[25405]_ , \new_[25406]_ , \new_[25407]_ , \new_[25408]_ ,
    \new_[25409]_ , \new_[25410]_ , \new_[25411]_ , \new_[25412]_ ,
    \new_[25413]_ , \new_[25414]_ , \new_[25415]_ , \new_[25416]_ ,
    \new_[25417]_ , \new_[25418]_ , \new_[25419]_ , \new_[25420]_ ,
    \new_[25421]_ , \new_[25422]_ , \new_[25423]_ , \new_[25424]_ ,
    \new_[25425]_ , \new_[25426]_ , \new_[25427]_ , \new_[25428]_ ,
    \new_[25429]_ , \new_[25430]_ , \new_[25431]_ , \new_[25432]_ ,
    \new_[25433]_ , \new_[25434]_ , \new_[25435]_ , \new_[25436]_ ,
    \new_[25437]_ , \new_[25438]_ , \new_[25439]_ , \new_[25440]_ ,
    \new_[25441]_ , \new_[25442]_ , \new_[25443]_ , \new_[25444]_ ,
    \new_[25445]_ , \new_[25446]_ , \new_[25447]_ , \new_[25448]_ ,
    \new_[25449]_ , \new_[25450]_ , \new_[25451]_ , \new_[25452]_ ,
    \new_[25453]_ , \new_[25454]_ , \new_[25455]_ , \new_[25456]_ ,
    \new_[25457]_ , \new_[25458]_ , \new_[25459]_ , \new_[25460]_ ,
    \new_[25461]_ , \new_[25462]_ , \new_[25463]_ , \new_[25464]_ ,
    \new_[25465]_ , \new_[25466]_ , \new_[25467]_ , \new_[25468]_ ,
    \new_[25469]_ , \new_[25470]_ , \new_[25471]_ , \new_[25472]_ ,
    \new_[25473]_ , \new_[25474]_ , \new_[25475]_ , \new_[25476]_ ,
    \new_[25477]_ , \new_[25478]_ , \new_[25479]_ , \new_[25480]_ ,
    \new_[25481]_ , \new_[25482]_ , \new_[25483]_ , \new_[25484]_ ,
    \new_[25485]_ , \new_[25486]_ , \new_[25487]_ , \new_[25488]_ ,
    \new_[25489]_ , \new_[25490]_ , \new_[25491]_ , \new_[25492]_ ,
    \new_[25493]_ , \new_[25494]_ , \new_[25495]_ , \new_[25496]_ ,
    \new_[25497]_ , \new_[25498]_ , \new_[25499]_ , \new_[25500]_ ,
    \new_[25501]_ , \new_[25502]_ , \new_[25503]_ , \new_[25504]_ ,
    \new_[25505]_ , \new_[25506]_ , \new_[25507]_ , \new_[25508]_ ,
    \new_[25509]_ , \new_[25510]_ , \new_[25511]_ , \new_[25512]_ ,
    \new_[25513]_ , \new_[25514]_ , \new_[25515]_ , \new_[25516]_ ,
    \new_[25517]_ , \new_[25518]_ , \new_[25519]_ , \new_[25520]_ ,
    \new_[25521]_ , \new_[25522]_ , \new_[25523]_ , \new_[25524]_ ,
    \new_[25525]_ , \new_[25526]_ , \new_[25527]_ , \new_[25528]_ ,
    \new_[25529]_ , \new_[25530]_ , \new_[25531]_ , \new_[25532]_ ,
    \new_[25533]_ , \new_[25534]_ , \new_[25535]_ , \new_[25536]_ ,
    \new_[25537]_ , \new_[25538]_ , \new_[25539]_ , \new_[25540]_ ,
    \new_[25541]_ , \new_[25542]_ , \new_[25543]_ , \new_[25544]_ ,
    \new_[25545]_ , \new_[25546]_ , \new_[25547]_ , \new_[25548]_ ,
    \new_[25549]_ , \new_[25550]_ , \new_[25551]_ , \new_[25552]_ ,
    \new_[25553]_ , \new_[25554]_ , \new_[25555]_ , \new_[25556]_ ,
    \new_[25557]_ , \new_[25558]_ , \new_[25559]_ , \new_[25560]_ ,
    \new_[25561]_ , \new_[25562]_ , \new_[25563]_ , \new_[25564]_ ,
    \new_[25565]_ , \new_[25566]_ , \new_[25567]_ , \new_[25568]_ ,
    \new_[25569]_ , \new_[25570]_ , \new_[25571]_ , \new_[25572]_ ,
    \new_[25573]_ , \new_[25574]_ , \new_[25575]_ , \new_[25576]_ ,
    \new_[25577]_ , \new_[25578]_ , \new_[25579]_ , \new_[25580]_ ,
    \new_[25581]_ , \new_[25582]_ , \new_[25583]_ , \new_[25584]_ ,
    \new_[25585]_ , \new_[25586]_ , \new_[25587]_ , \new_[25588]_ ,
    \new_[25589]_ , \new_[25590]_ , \new_[25591]_ , \new_[25592]_ ,
    \new_[25593]_ , \new_[25594]_ , \new_[25595]_ , \new_[25596]_ ,
    \new_[25597]_ , \new_[25598]_ , \new_[25599]_ , \new_[25600]_ ,
    \new_[25601]_ , \new_[25602]_ , \new_[25603]_ , \new_[25604]_ ,
    \new_[25605]_ , \new_[25606]_ , \new_[25607]_ , \new_[25608]_ ,
    \new_[25609]_ , \new_[25610]_ , \new_[25611]_ , \new_[25612]_ ,
    \new_[25613]_ , \new_[25614]_ , \new_[25615]_ , \new_[25616]_ ,
    \new_[25617]_ , \new_[25618]_ , \new_[25619]_ , \new_[25620]_ ,
    \new_[25621]_ , \new_[25622]_ , \new_[25623]_ , \new_[25624]_ ,
    \new_[25625]_ , \new_[25626]_ , \new_[25627]_ , \new_[25628]_ ,
    \new_[25629]_ , \new_[25630]_ , \new_[25631]_ , \new_[25632]_ ,
    \new_[25633]_ , \new_[25634]_ , \new_[25635]_ , \new_[25636]_ ,
    \new_[25637]_ , \new_[25638]_ , \new_[25639]_ , \new_[25640]_ ,
    \new_[25641]_ , \new_[25642]_ , \new_[25643]_ , \new_[25644]_ ,
    \new_[25645]_ , \new_[25646]_ , \new_[25647]_ , \new_[25648]_ ,
    \new_[25649]_ , \new_[25650]_ , \new_[25651]_ , \new_[25652]_ ,
    \new_[25653]_ , \new_[25654]_ , \new_[25655]_ , \new_[25656]_ ,
    \new_[25657]_ , \new_[25658]_ , \new_[25659]_ , \new_[25660]_ ,
    \new_[25661]_ , \new_[25662]_ , \new_[25663]_ , \new_[25664]_ ,
    \new_[25665]_ , \new_[25666]_ , \new_[25667]_ , \new_[25668]_ ,
    \new_[25669]_ , \new_[25670]_ , \new_[25671]_ , \new_[25672]_ ,
    \new_[25673]_ , \new_[25674]_ , \new_[25675]_ , \new_[25676]_ ,
    \new_[25677]_ , \new_[25678]_ , \new_[25679]_ , \new_[25680]_ ,
    \new_[25681]_ , \new_[25682]_ , \new_[25683]_ , \new_[25684]_ ,
    \new_[25685]_ , \new_[25686]_ , \new_[25687]_ , \new_[25688]_ ,
    \new_[25689]_ , \new_[25690]_ , \new_[25691]_ , \new_[25692]_ ,
    \new_[25693]_ , \new_[25694]_ , \new_[25695]_ , \new_[25696]_ ,
    \new_[25697]_ , \new_[25698]_ , \new_[25699]_ , \new_[25700]_ ,
    \new_[25701]_ , \new_[25702]_ , \new_[25703]_ , \new_[25704]_ ,
    \new_[25705]_ , \new_[25706]_ , \new_[25707]_ , \new_[25708]_ ,
    \new_[25709]_ , \new_[25710]_ , \new_[25711]_ , \new_[25712]_ ,
    \new_[25713]_ , \new_[25714]_ , \new_[25715]_ , \new_[25716]_ ,
    \new_[25717]_ , \new_[25718]_ , \new_[25719]_ , \new_[25720]_ ,
    \new_[25721]_ , \new_[25722]_ , \new_[25723]_ , \new_[25724]_ ,
    \new_[25725]_ , \new_[25726]_ , \new_[25727]_ , \new_[25728]_ ,
    \new_[25729]_ , \new_[25730]_ , \new_[25731]_ , \new_[25732]_ ,
    \new_[25733]_ , \new_[25734]_ , \new_[25735]_ , \new_[25736]_ ,
    \new_[25737]_ , \new_[25738]_ , \new_[25739]_ , \new_[25740]_ ,
    \new_[25741]_ , \new_[25742]_ , \new_[25743]_ , \new_[25744]_ ,
    \new_[25745]_ , \new_[25746]_ , \new_[25747]_ , \new_[25748]_ ,
    \new_[25749]_ , \new_[25750]_ , \new_[25751]_ , \new_[25752]_ ,
    \new_[25753]_ , \new_[25754]_ , \new_[25755]_ , \new_[25756]_ ,
    \new_[25757]_ , \new_[25758]_ , \new_[25759]_ , \new_[25760]_ ,
    \new_[25761]_ , \new_[25762]_ , \new_[25763]_ , \new_[25764]_ ,
    \new_[25765]_ , \new_[25766]_ , \new_[25767]_ , \new_[25768]_ ,
    \new_[25769]_ , \new_[25770]_ , \new_[25771]_ , \new_[25772]_ ,
    \new_[25773]_ , \new_[25774]_ , \new_[25775]_ , \new_[25776]_ ,
    \new_[25777]_ , \new_[25778]_ , \new_[25779]_ , \new_[25780]_ ,
    \new_[25781]_ , \new_[25782]_ , \new_[25783]_ , \new_[25784]_ ,
    \new_[25785]_ , \new_[25786]_ , \new_[25787]_ , \new_[25788]_ ,
    \new_[25789]_ , \new_[25790]_ , \new_[25791]_ , \new_[25792]_ ,
    \new_[25793]_ , \new_[25794]_ , \new_[25795]_ , \new_[25796]_ ,
    \new_[25797]_ , \new_[25798]_ , \new_[25799]_ , \new_[25800]_ ,
    \new_[25801]_ , \new_[25802]_ , \new_[25803]_ , \new_[25804]_ ,
    \new_[25805]_ , \new_[25806]_ , \new_[25807]_ , \new_[25808]_ ,
    \new_[25809]_ , \new_[25810]_ , \new_[25811]_ , \new_[25812]_ ,
    \new_[25813]_ , \new_[25814]_ , \new_[25815]_ , \new_[25816]_ ,
    \new_[25817]_ , \new_[25818]_ , \new_[25819]_ , \new_[25820]_ ,
    \new_[25821]_ , \new_[25822]_ , \new_[25823]_ , \new_[25824]_ ,
    \new_[25825]_ , \new_[25826]_ , \new_[25827]_ , \new_[25828]_ ,
    \new_[25829]_ , \new_[25830]_ , \new_[25831]_ , \new_[25832]_ ,
    \new_[25833]_ , \new_[25834]_ , \new_[25835]_ , \new_[25836]_ ,
    \new_[25837]_ , \new_[25838]_ , \new_[25839]_ , \new_[25840]_ ,
    \new_[25841]_ , \new_[25842]_ , \new_[25843]_ , \new_[25844]_ ,
    \new_[25845]_ , \new_[25846]_ , \new_[25847]_ , \new_[25848]_ ,
    \new_[25849]_ , \new_[25850]_ , \new_[25851]_ , \new_[25852]_ ,
    \new_[25853]_ , \new_[25854]_ , \new_[25855]_ , \new_[25856]_ ,
    \new_[25857]_ , \new_[25858]_ , \new_[25859]_ , \new_[25860]_ ,
    \new_[25861]_ , \new_[25862]_ , \new_[25863]_ , \new_[25864]_ ,
    \new_[25865]_ , \new_[25866]_ , \new_[25867]_ , \new_[25868]_ ,
    \new_[25869]_ , \new_[25870]_ , \new_[25871]_ , \new_[25872]_ ,
    \new_[25873]_ , \new_[25874]_ , \new_[25875]_ , \new_[25876]_ ,
    \new_[25877]_ , \new_[25878]_ , \new_[25879]_ , \new_[25880]_ ,
    \new_[25881]_ , \new_[25882]_ , \new_[25883]_ , \new_[25884]_ ,
    \new_[25885]_ , \new_[25886]_ , \new_[25887]_ , \new_[25888]_ ,
    \new_[25889]_ , \new_[25890]_ , \new_[25891]_ , \new_[25892]_ ,
    \new_[25893]_ , \new_[25894]_ , \new_[25895]_ , \new_[25896]_ ,
    \new_[25897]_ , \new_[25898]_ , \new_[25899]_ , \new_[25900]_ ,
    \new_[25901]_ , \new_[25902]_ , \new_[25903]_ , \new_[25904]_ ,
    \new_[25905]_ , \new_[25906]_ , \new_[25907]_ , \new_[25908]_ ,
    \new_[25909]_ , \new_[25910]_ , \new_[25911]_ , \new_[25912]_ ,
    \new_[25913]_ , \new_[25914]_ , \new_[25915]_ , \new_[25916]_ ,
    \new_[25917]_ , \new_[25918]_ , \new_[25919]_ , \new_[25920]_ ,
    \new_[25921]_ , \new_[25922]_ , \new_[25923]_ , \new_[25924]_ ,
    \new_[25925]_ , \new_[25926]_ , \new_[25927]_ , \new_[25928]_ ,
    \new_[25929]_ , \new_[25930]_ , \new_[25931]_ , \new_[25932]_ ,
    \new_[25933]_ , \new_[25934]_ , \new_[25935]_ , \new_[25936]_ ,
    \new_[25937]_ , \new_[25938]_ , \new_[25939]_ , \new_[25940]_ ,
    \new_[25941]_ , \new_[25942]_ , \new_[25943]_ , \new_[25944]_ ,
    \new_[25945]_ , \new_[25946]_ , \new_[25947]_ , \new_[25948]_ ,
    \new_[25949]_ , \new_[25950]_ , \new_[25951]_ , \new_[25952]_ ,
    \new_[25953]_ , \new_[25954]_ , \new_[25955]_ , \new_[25956]_ ,
    \new_[25957]_ , \new_[25958]_ , \new_[25959]_ , \new_[25960]_ ,
    \new_[25961]_ , \new_[25962]_ , \new_[25963]_ , \new_[25964]_ ,
    \new_[25965]_ , \new_[25966]_ , \new_[25967]_ , \new_[25968]_ ,
    \new_[25969]_ , \new_[25970]_ , \new_[25971]_ , \new_[25972]_ ,
    \new_[25973]_ , \new_[25974]_ , \new_[25975]_ , \new_[25976]_ ,
    \new_[25977]_ , \new_[25978]_ , \new_[25979]_ , \new_[25980]_ ,
    \new_[25981]_ , \new_[25982]_ , \new_[25983]_ , \new_[25984]_ ,
    \new_[25985]_ , \new_[25986]_ , \new_[25987]_ , \new_[25988]_ ,
    \new_[25989]_ , \new_[25990]_ , \new_[25991]_ , \new_[25992]_ ,
    \new_[25993]_ , \new_[25994]_ , \new_[25995]_ , \new_[25996]_ ,
    \new_[25997]_ , \new_[25998]_ , \new_[25999]_ , \new_[26000]_ ,
    \new_[26001]_ , \new_[26002]_ , \new_[26003]_ , \new_[26004]_ ,
    \new_[26005]_ , \new_[26006]_ , \new_[26007]_ , \new_[26008]_ ,
    \new_[26009]_ , \new_[26010]_ , \new_[26011]_ , \new_[26012]_ ,
    \new_[26013]_ , \new_[26014]_ , \new_[26015]_ , \new_[26016]_ ,
    \new_[26017]_ , \new_[26018]_ , \new_[26019]_ , \new_[26020]_ ,
    \new_[26021]_ , \new_[26022]_ , \new_[26023]_ , \new_[26024]_ ,
    \new_[26025]_ , \new_[26026]_ , \new_[26027]_ , \new_[26028]_ ,
    \new_[26029]_ , \new_[26030]_ , \new_[26031]_ , \new_[26032]_ ,
    \new_[26033]_ , \new_[26034]_ , \new_[26035]_ , \new_[26036]_ ,
    \new_[26037]_ , \new_[26038]_ , \new_[26039]_ , \new_[26040]_ ,
    \new_[26041]_ , \new_[26042]_ , \new_[26043]_ , \new_[26044]_ ,
    \new_[26045]_ , \new_[26046]_ , \new_[26047]_ , \new_[26048]_ ,
    \new_[26049]_ , \new_[26050]_ , \new_[26051]_ , \new_[26052]_ ,
    \new_[26053]_ , \new_[26054]_ , \new_[26055]_ , \new_[26056]_ ,
    \new_[26057]_ , \new_[26058]_ , \new_[26059]_ , \new_[26060]_ ,
    \new_[26061]_ , \new_[26062]_ , \new_[26063]_ , \new_[26064]_ ,
    \new_[26065]_ , \new_[26066]_ , \new_[26067]_ , \new_[26068]_ ,
    \new_[26069]_ , \new_[26070]_ , \new_[26071]_ , \new_[26072]_ ,
    \new_[26073]_ , \new_[26074]_ , \new_[26075]_ , \new_[26076]_ ,
    \new_[26077]_ , \new_[26078]_ , \new_[26079]_ , \new_[26080]_ ,
    \new_[26081]_ , \new_[26082]_ , \new_[26083]_ , \new_[26084]_ ,
    \new_[26085]_ , \new_[26086]_ , \new_[26087]_ , \new_[26088]_ ,
    \new_[26089]_ , \new_[26090]_ , \new_[26091]_ , \new_[26092]_ ,
    \new_[26093]_ , \new_[26094]_ , \new_[26095]_ , \new_[26096]_ ,
    \new_[26097]_ , \new_[26098]_ , \new_[26099]_ , \new_[26100]_ ,
    \new_[26101]_ , \new_[26102]_ , \new_[26103]_ , \new_[26104]_ ,
    \new_[26105]_ , \new_[26106]_ , \new_[26107]_ , \new_[26108]_ ,
    \new_[26109]_ , \new_[26110]_ , \new_[26111]_ , \new_[26112]_ ,
    \new_[26113]_ , \new_[26114]_ , \new_[26115]_ , \new_[26116]_ ,
    \new_[26117]_ , \new_[26118]_ , \new_[26119]_ , \new_[26120]_ ,
    \new_[26121]_ , \new_[26122]_ , \new_[26123]_ , \new_[26124]_ ,
    \new_[26125]_ , \new_[26126]_ , \new_[26127]_ , \new_[26128]_ ,
    \new_[26129]_ , \new_[26130]_ , \new_[26131]_ , \new_[26132]_ ,
    \new_[26133]_ , \new_[26134]_ , \new_[26135]_ , \new_[26136]_ ,
    \new_[26137]_ , \new_[26138]_ , \new_[26139]_ , \new_[26140]_ ,
    \new_[26141]_ , \new_[26142]_ , \new_[26143]_ , \new_[26144]_ ,
    \new_[26145]_ , \new_[26146]_ , \new_[26147]_ , \new_[26148]_ ,
    \new_[26149]_ , \new_[26150]_ , \new_[26151]_ , \new_[26152]_ ,
    \new_[26153]_ , \new_[26154]_ , \new_[26155]_ , \new_[26156]_ ,
    \new_[26157]_ , \new_[26158]_ , \new_[26159]_ , \new_[26160]_ ,
    \new_[26161]_ , \new_[26162]_ , \new_[26163]_ , \new_[26164]_ ,
    \new_[26165]_ , \new_[26166]_ , \new_[26167]_ , \new_[26168]_ ,
    \new_[26169]_ , \new_[26170]_ , \new_[26171]_ , \new_[26172]_ ,
    \new_[26173]_ , \new_[26174]_ , \new_[26175]_ , \new_[26176]_ ,
    \new_[26177]_ , \new_[26178]_ , \new_[26179]_ , \new_[26180]_ ,
    \new_[26181]_ , \new_[26182]_ , \new_[26183]_ , \new_[26184]_ ,
    \new_[26185]_ , \new_[26186]_ , \new_[26187]_ , \new_[26188]_ ,
    \new_[26189]_ , \new_[26190]_ , \new_[26191]_ , \new_[26192]_ ,
    \new_[26193]_ , \new_[26194]_ , \new_[26195]_ , \new_[26196]_ ,
    \new_[26197]_ , \new_[26198]_ , \new_[26199]_ , \new_[26200]_ ,
    \new_[26201]_ , \new_[26202]_ , \new_[26203]_ , \new_[26204]_ ,
    \new_[26205]_ , \new_[26206]_ , \new_[26207]_ , \new_[26208]_ ,
    \new_[26209]_ , \new_[26210]_ , \new_[26211]_ , \new_[26212]_ ,
    \new_[26213]_ , \new_[26214]_ , \new_[26215]_ , \new_[26216]_ ,
    \new_[26217]_ , \new_[26218]_ , \new_[26219]_ , \new_[26220]_ ,
    \new_[26221]_ , \new_[26222]_ , \new_[26223]_ , \new_[26224]_ ,
    \new_[26225]_ , \new_[26226]_ , \new_[26227]_ , \new_[26228]_ ,
    \new_[26229]_ , \new_[26230]_ , \new_[26231]_ , \new_[26232]_ ,
    \new_[26233]_ , \new_[26234]_ , \new_[26235]_ , \new_[26236]_ ,
    \new_[26237]_ , \new_[26238]_ , \new_[26239]_ , \new_[26240]_ ,
    \new_[26241]_ , \new_[26242]_ , \new_[26243]_ , \new_[26244]_ ,
    \new_[26245]_ , \new_[26246]_ , \new_[26247]_ , \new_[26248]_ ,
    \new_[26249]_ , \new_[26250]_ , \new_[26251]_ , \new_[26252]_ ,
    \new_[26253]_ , \new_[26254]_ , \new_[26255]_ , \new_[26256]_ ,
    \new_[26257]_ , \new_[26258]_ , \new_[26259]_ , \new_[26260]_ ,
    \new_[26261]_ , \new_[26262]_ , \new_[26263]_ , \new_[26264]_ ,
    \new_[26265]_ , \new_[26266]_ , \new_[26267]_ , \new_[26268]_ ,
    \new_[26269]_ , \new_[26270]_ , \new_[26271]_ , \new_[26272]_ ,
    \new_[26273]_ , \new_[26274]_ , \new_[26275]_ , \new_[26276]_ ,
    \new_[26277]_ , \new_[26278]_ , \new_[26279]_ , \new_[26280]_ ,
    \new_[26281]_ , \new_[26282]_ , \new_[26283]_ , \new_[26284]_ ,
    \new_[26285]_ , \new_[26286]_ , \new_[26287]_ , \new_[26288]_ ,
    \new_[26289]_ , \new_[26290]_ , \new_[26291]_ , \new_[26292]_ ,
    \new_[26293]_ , \new_[26294]_ , \new_[26295]_ , \new_[26296]_ ,
    \new_[26297]_ , \new_[26298]_ , \new_[26299]_ , \new_[26300]_ ,
    \new_[26301]_ , \new_[26302]_ , \new_[26303]_ , \new_[26304]_ ,
    \new_[26305]_ , \new_[26306]_ , \new_[26307]_ , \new_[26308]_ ,
    \new_[26309]_ , \new_[26310]_ , \new_[26311]_ , \new_[26312]_ ,
    \new_[26313]_ , \new_[26314]_ , \new_[26315]_ , \new_[26316]_ ,
    \new_[26317]_ , \new_[26318]_ , \new_[26319]_ , \new_[26320]_ ,
    \new_[26321]_ , \new_[26322]_ , \new_[26323]_ , \new_[26324]_ ,
    \new_[26325]_ , \new_[26326]_ , \new_[26327]_ , \new_[26328]_ ,
    \new_[26329]_ , \new_[26330]_ , \new_[26331]_ , \new_[26332]_ ,
    \new_[26333]_ , \new_[26334]_ , \new_[26335]_ , \new_[26336]_ ,
    \new_[26337]_ , \new_[26338]_ , \new_[26339]_ , \new_[26340]_ ,
    \new_[26341]_ , \new_[26342]_ , \new_[26343]_ , \new_[26344]_ ,
    \new_[26345]_ , \new_[26346]_ , \new_[26347]_ , \new_[26348]_ ,
    \new_[26349]_ , \new_[26350]_ , \new_[26351]_ , \new_[26352]_ ,
    \new_[26353]_ , \new_[26354]_ , \new_[26355]_ , \new_[26356]_ ,
    \new_[26357]_ , \new_[26358]_ , \new_[26359]_ , \new_[26360]_ ,
    \new_[26361]_ , \new_[26362]_ , \new_[26363]_ , \new_[26364]_ ,
    \new_[26365]_ , \new_[26366]_ , \new_[26367]_ , \new_[26368]_ ,
    \new_[26369]_ , \new_[26370]_ , \new_[26371]_ , \new_[26372]_ ,
    \new_[26373]_ , \new_[26374]_ , \new_[26375]_ , \new_[26376]_ ,
    \new_[26377]_ , \new_[26378]_ , \new_[26379]_ , \new_[26380]_ ,
    \new_[26381]_ , \new_[26382]_ , \new_[26383]_ , \new_[26384]_ ,
    \new_[26385]_ , \new_[26386]_ , \new_[26387]_ , \new_[26388]_ ,
    \new_[26389]_ , \new_[26390]_ , \new_[26391]_ , \new_[26392]_ ,
    \new_[26393]_ , \new_[26394]_ , \new_[26395]_ , \new_[26396]_ ,
    \new_[26397]_ , \new_[26398]_ , \new_[26399]_ , \new_[26400]_ ,
    \new_[26401]_ , \new_[26402]_ , \new_[26403]_ , \new_[26404]_ ,
    \new_[26405]_ , \new_[26406]_ , \new_[26407]_ , \new_[26408]_ ,
    \new_[26409]_ , \new_[26410]_ , \new_[26411]_ , \new_[26412]_ ,
    \new_[26413]_ , \new_[26414]_ , \new_[26415]_ , \new_[26416]_ ,
    \new_[26417]_ , \new_[26418]_ , \new_[26419]_ , \new_[26420]_ ,
    \new_[26421]_ , \new_[26422]_ , \new_[26423]_ , \new_[26424]_ ,
    \new_[26425]_ , \new_[26426]_ , \new_[26427]_ , \new_[26428]_ ,
    \new_[26429]_ , \new_[26430]_ , \new_[26431]_ , \new_[26432]_ ,
    \new_[26433]_ , \new_[26434]_ , \new_[26435]_ , \new_[26436]_ ,
    \new_[26437]_ , \new_[26438]_ , \new_[26439]_ , \new_[26440]_ ,
    \new_[26441]_ , \new_[26442]_ , \new_[26443]_ , \new_[26444]_ ,
    \new_[26445]_ , \new_[26446]_ , \new_[26447]_ , \new_[26448]_ ,
    \new_[26449]_ , \new_[26450]_ , \new_[26451]_ , \new_[26452]_ ,
    \new_[26453]_ , \new_[26454]_ , \new_[26455]_ , \new_[26456]_ ,
    \new_[26457]_ , \new_[26458]_ , \new_[26459]_ , \new_[26460]_ ,
    \new_[26461]_ , \new_[26462]_ , \new_[26463]_ , \new_[26464]_ ,
    \new_[26465]_ , \new_[26466]_ , \new_[26467]_ , \new_[26468]_ ,
    \new_[26469]_ , \new_[26470]_ , \new_[26471]_ , \new_[26472]_ ,
    \new_[26473]_ , \new_[26474]_ , \new_[26475]_ , \new_[26476]_ ,
    \new_[26477]_ , \new_[26478]_ , \new_[26479]_ , \new_[26480]_ ,
    \new_[26481]_ , \new_[26482]_ , \new_[26483]_ , \new_[26484]_ ,
    \new_[26485]_ , \new_[26486]_ , \new_[26487]_ , \new_[26488]_ ,
    \new_[26489]_ , \new_[26490]_ , \new_[26491]_ , \new_[26492]_ ,
    \new_[26493]_ , \new_[26494]_ , \new_[26495]_ , \new_[26496]_ ,
    \new_[26497]_ , \new_[26498]_ , \new_[26499]_ , \new_[26500]_ ,
    \new_[26501]_ , \new_[26502]_ , \new_[26503]_ , \new_[26504]_ ,
    \new_[26505]_ , \new_[26506]_ , \new_[26507]_ , \new_[26508]_ ,
    \new_[26509]_ , \new_[26510]_ , \new_[26511]_ , \new_[26512]_ ,
    \new_[26513]_ , \new_[26514]_ , \new_[26515]_ , \new_[26516]_ ,
    \new_[26517]_ , \new_[26518]_ , \new_[26519]_ , \new_[26520]_ ,
    \new_[26521]_ , \new_[26522]_ , \new_[26523]_ , \new_[26524]_ ,
    \new_[26525]_ , \new_[26526]_ , \new_[26527]_ , \new_[26528]_ ,
    \new_[26529]_ , \new_[26530]_ , \new_[26531]_ , \new_[26532]_ ,
    \new_[26533]_ , \new_[26534]_ , \new_[26535]_ , \new_[26536]_ ,
    \new_[26537]_ , \new_[26538]_ , \new_[26539]_ , \new_[26540]_ ,
    \new_[26541]_ , \new_[26542]_ , \new_[26543]_ , \new_[26544]_ ,
    \new_[26545]_ , \new_[26546]_ , \new_[26547]_ , \new_[26548]_ ,
    \new_[26549]_ , \new_[26550]_ , \new_[26551]_ , \new_[26552]_ ,
    \new_[26553]_ , \new_[26554]_ , \new_[26555]_ , \new_[26556]_ ,
    \new_[26557]_ , \new_[26558]_ , \new_[26559]_ , \new_[26560]_ ,
    \new_[26561]_ , \new_[26562]_ , \new_[26563]_ , \new_[26564]_ ,
    \new_[26565]_ , \new_[26566]_ , \new_[26567]_ , \new_[26568]_ ,
    \new_[26569]_ , \new_[26570]_ , \new_[26571]_ , \new_[26572]_ ,
    \new_[26573]_ , \new_[26574]_ , \new_[26575]_ , \new_[26576]_ ,
    \new_[26577]_ , \new_[26578]_ , \new_[26579]_ , \new_[26580]_ ,
    \new_[26581]_ , \new_[26582]_ , \new_[26583]_ , \new_[26584]_ ,
    \new_[26585]_ , \new_[26586]_ , \new_[26587]_ , \new_[26588]_ ,
    \new_[26589]_ , \new_[26590]_ , \new_[26591]_ , \new_[26592]_ ,
    \new_[26593]_ , \new_[26594]_ , \new_[26595]_ , \new_[26596]_ ,
    \new_[26597]_ , \new_[26598]_ , \new_[26599]_ , \new_[26600]_ ,
    \new_[26601]_ , \new_[26602]_ , \new_[26603]_ , \new_[26604]_ ,
    \new_[26605]_ , \new_[26606]_ , \new_[26607]_ , \new_[26608]_ ,
    \new_[26609]_ , \new_[26610]_ , \new_[26611]_ , \new_[26612]_ ,
    \new_[26613]_ , \new_[26614]_ , \new_[26615]_ , \new_[26616]_ ,
    \new_[26617]_ , \new_[26618]_ , \new_[26619]_ , \new_[26620]_ ,
    \new_[26621]_ , \new_[26622]_ , \new_[26623]_ , \new_[26624]_ ,
    \new_[26625]_ , \new_[26626]_ , \new_[26627]_ , \new_[26628]_ ,
    \new_[26629]_ , \new_[26630]_ , \new_[26631]_ , \new_[26632]_ ,
    \new_[26633]_ , \new_[26634]_ , \new_[26635]_ , \new_[26636]_ ,
    \new_[26637]_ , \new_[26638]_ , \new_[26639]_ , \new_[26640]_ ,
    \new_[26641]_ , \new_[26642]_ , \new_[26643]_ , \new_[26644]_ ,
    \new_[26645]_ , \new_[26646]_ , \new_[26647]_ , \new_[26648]_ ,
    \new_[26649]_ , \new_[26650]_ , \new_[26651]_ , \new_[26652]_ ,
    \new_[26653]_ , \new_[26654]_ , \new_[26655]_ , \new_[26656]_ ,
    \new_[26657]_ , \new_[26658]_ , \new_[26659]_ , \new_[26660]_ ,
    \new_[26661]_ , \new_[26662]_ , \new_[26663]_ , \new_[26664]_ ,
    \new_[26665]_ , \new_[26666]_ , \new_[26667]_ , \new_[26668]_ ,
    \new_[26669]_ , \new_[26670]_ , \new_[26671]_ , \new_[26672]_ ,
    \new_[26673]_ , \new_[26674]_ , \new_[26675]_ , \new_[26676]_ ,
    \new_[26677]_ , \new_[26678]_ , \new_[26679]_ , \new_[26680]_ ,
    \new_[26681]_ , \new_[26682]_ , \new_[26683]_ , \new_[26684]_ ,
    \new_[26685]_ , \new_[26686]_ , \new_[26687]_ , \new_[26688]_ ,
    \new_[26689]_ , \new_[26690]_ , \new_[26691]_ , \new_[26692]_ ,
    \new_[26693]_ , \new_[26694]_ , \new_[26695]_ , \new_[26696]_ ,
    \new_[26697]_ , \new_[26698]_ , \new_[26699]_ , \new_[26700]_ ,
    \new_[26701]_ , \new_[26702]_ , \new_[26703]_ , \new_[26704]_ ,
    \new_[26705]_ , \new_[26706]_ , \new_[26707]_ , \new_[26708]_ ,
    \new_[26709]_ , \new_[26710]_ , \new_[26711]_ , \new_[26712]_ ,
    \new_[26713]_ , \new_[26714]_ , \new_[26715]_ , \new_[26716]_ ,
    \new_[26717]_ , \new_[26718]_ , \new_[26719]_ , \new_[26720]_ ,
    \new_[26721]_ , \new_[26722]_ , \new_[26723]_ , \new_[26724]_ ,
    \new_[26725]_ , \new_[26726]_ , \new_[26727]_ , \new_[26728]_ ,
    \new_[26729]_ , \new_[26730]_ , \new_[26731]_ , \new_[26732]_ ,
    \new_[26733]_ , \new_[26734]_ , \new_[26735]_ , \new_[26736]_ ,
    \new_[26737]_ , \new_[26738]_ , \new_[26739]_ , \new_[26740]_ ,
    \new_[26741]_ , \new_[26742]_ , \new_[26743]_ , \new_[26744]_ ,
    \new_[26745]_ , \new_[26746]_ , \new_[26747]_ , \new_[26748]_ ,
    \new_[26749]_ , \new_[26750]_ , \new_[26751]_ , \new_[26752]_ ,
    \new_[26753]_ , \new_[26754]_ , \new_[26755]_ , \new_[26756]_ ,
    \new_[26757]_ , \new_[26758]_ , \new_[26759]_ , \new_[26760]_ ,
    \new_[26761]_ , \new_[26762]_ , \new_[26763]_ , \new_[26764]_ ,
    \new_[26765]_ , \new_[26766]_ , \new_[26767]_ , \new_[26768]_ ,
    \new_[26769]_ , \new_[26770]_ , \new_[26771]_ , \new_[26772]_ ,
    \new_[26773]_ , \new_[26774]_ , \new_[26775]_ , \new_[26776]_ ,
    \new_[26777]_ , \new_[26778]_ , \new_[26779]_ , \new_[26780]_ ,
    \new_[26781]_ , \new_[26782]_ , \new_[26783]_ , \new_[26784]_ ,
    \new_[26785]_ , \new_[26786]_ , \new_[26787]_ , \new_[26788]_ ,
    \new_[26789]_ , \new_[26790]_ , \new_[26791]_ , \new_[26792]_ ,
    \new_[26793]_ , \new_[26794]_ , \new_[26795]_ , \new_[26796]_ ,
    \new_[26797]_ , \new_[26798]_ , \new_[26799]_ , \new_[26800]_ ,
    \new_[26801]_ , \new_[26802]_ , \new_[26803]_ , \new_[26804]_ ,
    \new_[26805]_ , \new_[26806]_ , \new_[26807]_ , \new_[26808]_ ,
    \new_[26809]_ , \new_[26810]_ , \new_[26811]_ , \new_[26812]_ ,
    \new_[26813]_ , \new_[26814]_ , \new_[26815]_ , \new_[26816]_ ,
    \new_[26817]_ , \new_[26818]_ , \new_[26819]_ , \new_[26820]_ ,
    \new_[26821]_ , \new_[26822]_ , \new_[26823]_ , \new_[26824]_ ,
    \new_[26825]_ , \new_[26826]_ , \new_[26827]_ , \new_[26828]_ ,
    \new_[26829]_ , \new_[26830]_ , \new_[26831]_ , \new_[26832]_ ,
    \new_[26833]_ , \new_[26834]_ , \new_[26835]_ , \new_[26836]_ ,
    \new_[26837]_ , \new_[26838]_ , \new_[26839]_ , \new_[26840]_ ,
    \new_[26841]_ , \new_[26842]_ , \new_[26843]_ , \new_[26844]_ ,
    \new_[26845]_ , \new_[26846]_ , \new_[26847]_ , \new_[26848]_ ,
    \new_[26849]_ , \new_[26850]_ , \new_[26851]_ , \new_[26852]_ ,
    \new_[26853]_ , \new_[26854]_ , \new_[26855]_ , \new_[26856]_ ,
    \new_[26857]_ , \new_[26858]_ , \new_[26859]_ , \new_[26860]_ ,
    \new_[26861]_ , \new_[26862]_ , \new_[26863]_ , \new_[26864]_ ,
    \new_[26865]_ , \new_[26866]_ , \new_[26867]_ , \new_[26868]_ ,
    \new_[26869]_ , \new_[26870]_ , \new_[26871]_ , \new_[26872]_ ,
    \new_[26873]_ , \new_[26874]_ , \new_[26875]_ , \new_[26876]_ ,
    \new_[26877]_ , \new_[26878]_ , \new_[26879]_ , \new_[26880]_ ,
    \new_[26881]_ , \new_[26882]_ , \new_[26883]_ , \new_[26884]_ ,
    \new_[26885]_ , \new_[26886]_ , \new_[26887]_ , \new_[26888]_ ,
    \new_[26889]_ , \new_[26890]_ , \new_[26891]_ , \new_[26892]_ ,
    \new_[26893]_ , \new_[26894]_ , \new_[26895]_ , \new_[26896]_ ,
    \new_[26897]_ , \new_[26898]_ , \new_[26899]_ , \new_[26900]_ ,
    \new_[26901]_ , \new_[26902]_ , \new_[26903]_ , \new_[26904]_ ,
    \new_[26905]_ , \new_[26906]_ , \new_[26907]_ , \new_[26908]_ ,
    \new_[26909]_ , \new_[26910]_ , \new_[26911]_ , \new_[26912]_ ,
    \new_[26913]_ , \new_[26914]_ , \new_[26915]_ , \new_[26916]_ ,
    \new_[26917]_ , \new_[26918]_ , \new_[26919]_ , \new_[26920]_ ,
    \new_[26921]_ , \new_[26922]_ , \new_[26923]_ , \new_[26924]_ ,
    \new_[26925]_ , \new_[26926]_ , \new_[26927]_ , \new_[26928]_ ,
    \new_[26929]_ , \new_[26930]_ , \new_[26931]_ , \new_[26932]_ ,
    \new_[26933]_ , \new_[26934]_ , \new_[26935]_ , \new_[26936]_ ,
    \new_[26937]_ , \new_[26938]_ , \new_[26939]_ , \new_[26940]_ ,
    \new_[26941]_ , \new_[26942]_ , \new_[26943]_ , \new_[26944]_ ,
    \new_[26945]_ , \new_[26946]_ , \new_[26947]_ , \new_[26948]_ ,
    \new_[26949]_ , \new_[26950]_ , \new_[26951]_ , \new_[26952]_ ,
    \new_[26953]_ , \new_[26954]_ , \new_[26955]_ , \new_[26956]_ ,
    \new_[26957]_ , \new_[26958]_ , \new_[26959]_ , \new_[26960]_ ,
    \new_[26961]_ , \new_[26962]_ , \new_[26963]_ , \new_[26964]_ ,
    \new_[26965]_ , \new_[26966]_ , \new_[26967]_ , \new_[26968]_ ,
    \new_[26969]_ , \new_[26970]_ , \new_[26971]_ , \new_[26972]_ ,
    \new_[26973]_ , \new_[26974]_ , \new_[26975]_ , \new_[26976]_ ,
    \new_[26977]_ , \new_[26978]_ , \new_[26979]_ , \new_[26980]_ ,
    \new_[26981]_ , \new_[26982]_ , \new_[26983]_ , \new_[26984]_ ,
    \new_[26985]_ , \new_[26986]_ , \new_[26987]_ , \new_[26988]_ ,
    \new_[26989]_ , \new_[26990]_ , \new_[26991]_ , \new_[26992]_ ,
    \new_[26993]_ , \new_[26994]_ , \new_[26995]_ , \new_[26996]_ ,
    \new_[26997]_ , \new_[26998]_ , \new_[26999]_ , \new_[27000]_ ,
    \new_[27001]_ , \new_[27002]_ , \new_[27003]_ , \new_[27004]_ ,
    \new_[27005]_ , \new_[27006]_ , \new_[27007]_ , \new_[27008]_ ,
    \new_[27009]_ , \new_[27010]_ , \new_[27011]_ , \new_[27012]_ ,
    \new_[27013]_ , \new_[27014]_ , \new_[27015]_ , \new_[27016]_ ,
    \new_[27017]_ , \new_[27018]_ , \new_[27019]_ , \new_[27020]_ ,
    \new_[27021]_ , \new_[27022]_ , \new_[27023]_ , \new_[27024]_ ,
    \new_[27025]_ , \new_[27026]_ , \new_[27027]_ , \new_[27028]_ ,
    \new_[27029]_ , \new_[27030]_ , \new_[27031]_ , \new_[27032]_ ,
    \new_[27033]_ , \new_[27034]_ , \new_[27035]_ , \new_[27036]_ ,
    \new_[27037]_ , \new_[27038]_ , \new_[27039]_ , \new_[27040]_ ,
    \new_[27041]_ , \new_[27042]_ , \new_[27043]_ , \new_[27044]_ ,
    \new_[27045]_ , \new_[27046]_ , \new_[27047]_ , \new_[27048]_ ,
    \new_[27049]_ , \new_[27050]_ , \new_[27051]_ , \new_[27052]_ ,
    \new_[27053]_ , \new_[27054]_ , \new_[27055]_ , \new_[27056]_ ,
    \new_[27057]_ , \new_[27058]_ , \new_[27059]_ , \new_[27060]_ ,
    \new_[27061]_ , \new_[27062]_ , \new_[27063]_ , \new_[27064]_ ,
    \new_[27065]_ , \new_[27066]_ , \new_[27067]_ , \new_[27068]_ ,
    \new_[27069]_ , \new_[27070]_ , \new_[27071]_ , \new_[27072]_ ,
    \new_[27073]_ , \new_[27074]_ , \new_[27075]_ , \new_[27076]_ ,
    \new_[27077]_ , \new_[27078]_ , \new_[27079]_ , \new_[27080]_ ,
    \new_[27081]_ , \new_[27082]_ , \new_[27083]_ , \new_[27084]_ ,
    \new_[27085]_ , \new_[27086]_ , \new_[27087]_ , \new_[27088]_ ,
    \new_[27089]_ , \new_[27090]_ , \new_[27091]_ , \new_[27092]_ ,
    \new_[27093]_ , \new_[27094]_ , \new_[27095]_ , \new_[27096]_ ,
    \new_[27097]_ , \new_[27098]_ , \new_[27099]_ , \new_[27100]_ ,
    \new_[27101]_ , \new_[27102]_ , \new_[27103]_ , \new_[27104]_ ,
    \new_[27105]_ , \new_[27106]_ , \new_[27107]_ , \new_[27108]_ ,
    \new_[27109]_ , \new_[27110]_ , \new_[27111]_ , \new_[27112]_ ,
    \new_[27113]_ , \new_[27114]_ , \new_[27115]_ , \new_[27116]_ ,
    \new_[27117]_ , \new_[27118]_ , \new_[27119]_ , \new_[27120]_ ,
    \new_[27121]_ , \new_[27122]_ , \new_[27123]_ , \new_[27124]_ ,
    \new_[27125]_ , \new_[27126]_ , \new_[27127]_ , \new_[27128]_ ,
    \new_[27129]_ , \new_[27130]_ , \new_[27131]_ , \new_[27132]_ ,
    \new_[27133]_ , \new_[27134]_ , \new_[27135]_ , \new_[27136]_ ,
    \new_[27137]_ , \new_[27138]_ , \new_[27139]_ , \new_[27140]_ ,
    \new_[27141]_ , \new_[27142]_ , \new_[27143]_ , \new_[27144]_ ,
    \new_[27145]_ , \new_[27146]_ , \new_[27147]_ , \new_[27148]_ ,
    \new_[27149]_ , \new_[27150]_ , \new_[27151]_ , \new_[27152]_ ,
    \new_[27153]_ , \new_[27154]_ , \new_[27155]_ , \new_[27156]_ ,
    \new_[27157]_ , \new_[27158]_ , \new_[27159]_ , \new_[27160]_ ,
    \new_[27161]_ , \new_[27162]_ , \new_[27163]_ , \new_[27164]_ ,
    \new_[27165]_ , \new_[27166]_ , \new_[27167]_ , \new_[27168]_ ,
    \new_[27169]_ , \new_[27170]_ , \new_[27171]_ , \new_[27172]_ ,
    \new_[27173]_ , \new_[27174]_ , \new_[27175]_ , \new_[27176]_ ,
    \new_[27177]_ , \new_[27178]_ , \new_[27179]_ , \new_[27180]_ ,
    \new_[27181]_ , \new_[27182]_ , \new_[27183]_ , \new_[27184]_ ,
    \new_[27185]_ , \new_[27186]_ , \new_[27187]_ , \new_[27188]_ ,
    \new_[27189]_ , \new_[27190]_ , \new_[27191]_ , \new_[27192]_ ,
    \new_[27193]_ , \new_[27194]_ , \new_[27195]_ , \new_[27196]_ ,
    \new_[27197]_ , \new_[27198]_ , \new_[27199]_ , \new_[27200]_ ,
    \new_[27201]_ , \new_[27202]_ , \new_[27203]_ , \new_[27204]_ ,
    \new_[27205]_ , \new_[27206]_ , \new_[27207]_ , \new_[27208]_ ,
    \new_[27209]_ , \new_[27210]_ , \new_[27211]_ , \new_[27212]_ ,
    \new_[27213]_ , \new_[27214]_ , \new_[27215]_ , \new_[27216]_ ,
    \new_[27217]_ , \new_[27218]_ , \new_[27219]_ , \new_[27220]_ ,
    \new_[27221]_ , \new_[27222]_ , \new_[27223]_ , \new_[27224]_ ,
    \new_[27225]_ , \new_[27226]_ , \new_[27227]_ , \new_[27228]_ ,
    \new_[27229]_ , \new_[27230]_ , \new_[27231]_ , \new_[27232]_ ,
    \new_[27233]_ , \new_[27234]_ , \new_[27235]_ , \new_[27236]_ ,
    \new_[27237]_ , \new_[27238]_ , \new_[27239]_ , \new_[27240]_ ,
    \new_[27241]_ , \new_[27242]_ , \new_[27243]_ , \new_[27244]_ ,
    \new_[27245]_ , \new_[27246]_ , \new_[27247]_ , \new_[27248]_ ,
    \new_[27249]_ , \new_[27250]_ , \new_[27251]_ , \new_[27252]_ ,
    \new_[27253]_ , \new_[27254]_ , \new_[27255]_ , \new_[27256]_ ,
    \new_[27257]_ , \new_[27258]_ , \new_[27259]_ , \new_[27260]_ ,
    \new_[27261]_ , \new_[27262]_ , \new_[27263]_ , \new_[27264]_ ,
    \new_[27265]_ , \new_[27266]_ , \new_[27267]_ , \new_[27268]_ ,
    \new_[27269]_ , \new_[27270]_ , \new_[27271]_ , \new_[27272]_ ,
    \new_[27273]_ , \new_[27274]_ , \new_[27275]_ , \new_[27276]_ ,
    \new_[27277]_ , \new_[27278]_ , \new_[27279]_ , \new_[27280]_ ,
    \new_[27281]_ , \new_[27282]_ , \new_[27283]_ , \new_[27284]_ ,
    \new_[27285]_ , \new_[27286]_ , \new_[27287]_ , \new_[27288]_ ,
    \new_[27289]_ , \new_[27290]_ , \new_[27291]_ , \new_[27292]_ ,
    \new_[27293]_ , \new_[27294]_ , \new_[27295]_ , \new_[27296]_ ,
    \new_[27297]_ , \new_[27298]_ , \new_[27299]_ , \new_[27300]_ ,
    \new_[27301]_ , \new_[27302]_ , \new_[27303]_ , \new_[27304]_ ,
    \new_[27305]_ , \new_[27306]_ , \new_[27307]_ , \new_[27308]_ ,
    \new_[27309]_ , \new_[27310]_ , \new_[27311]_ , \new_[27312]_ ,
    \new_[27313]_ , \new_[27314]_ , \new_[27315]_ , \new_[27316]_ ,
    \new_[27317]_ , \new_[27318]_ , \new_[27319]_ , \new_[27320]_ ,
    \new_[27321]_ , \new_[27322]_ , \new_[27323]_ , \new_[27324]_ ,
    \new_[27325]_ , \new_[27326]_ , \new_[27327]_ , \new_[27328]_ ,
    \new_[27329]_ , \new_[27330]_ , \new_[27331]_ , \new_[27332]_ ,
    \new_[27333]_ , \new_[27334]_ , \new_[27335]_ , \new_[27336]_ ,
    \new_[27337]_ , \new_[27338]_ , \new_[27339]_ , \new_[27340]_ ,
    \new_[27341]_ , \new_[27342]_ , \new_[27343]_ , \new_[27344]_ ,
    \new_[27345]_ , \new_[27346]_ , \new_[27347]_ , \new_[27348]_ ,
    \new_[27349]_ , \new_[27350]_ , \new_[27351]_ , \new_[27352]_ ,
    \new_[27353]_ , \new_[27354]_ , \new_[27355]_ , \new_[27356]_ ,
    \new_[27357]_ , \new_[27358]_ , \new_[27359]_ , \new_[27360]_ ,
    \new_[27361]_ , \new_[27362]_ , \new_[27363]_ , \new_[27364]_ ,
    \new_[27365]_ , \new_[27366]_ , \new_[27367]_ , \new_[27368]_ ,
    \new_[27369]_ , \new_[27370]_ , \new_[27371]_ , \new_[27372]_ ,
    \new_[27373]_ , \new_[27374]_ , \new_[27375]_ , \new_[27376]_ ,
    \new_[27377]_ , \new_[27378]_ , \new_[27379]_ , \new_[27380]_ ,
    \new_[27381]_ , \new_[27382]_ , \new_[27383]_ , \new_[27384]_ ,
    \new_[27385]_ , \new_[27386]_ , \new_[27387]_ , \new_[27388]_ ,
    \new_[27389]_ , \new_[27390]_ , \new_[27391]_ , \new_[27392]_ ,
    \new_[27393]_ , \new_[27394]_ , \new_[27395]_ , \new_[27396]_ ,
    \new_[27397]_ , \new_[27398]_ , \new_[27399]_ , \new_[27400]_ ,
    \new_[27401]_ , \new_[27402]_ , \new_[27403]_ , \new_[27404]_ ,
    \new_[27405]_ , \new_[27406]_ , \new_[27407]_ , \new_[27408]_ ,
    \new_[27409]_ , \new_[27410]_ , \new_[27411]_ , \new_[27412]_ ,
    \new_[27413]_ , \new_[27414]_ , \new_[27415]_ , \new_[27416]_ ,
    \new_[27417]_ , \new_[27418]_ , \new_[27419]_ , \new_[27420]_ ,
    \new_[27421]_ , \new_[27422]_ , \new_[27423]_ , \new_[27424]_ ,
    \new_[27425]_ , \new_[27426]_ , \new_[27427]_ , \new_[27428]_ ,
    \new_[27429]_ , \new_[27430]_ , \new_[27431]_ , \new_[27432]_ ,
    \new_[27433]_ , \new_[27434]_ , \new_[27435]_ , \new_[27436]_ ,
    \new_[27437]_ , \new_[27438]_ , \new_[27439]_ , \new_[27440]_ ,
    \new_[27441]_ , \new_[27442]_ , \new_[27443]_ , \new_[27444]_ ,
    \new_[27445]_ , \new_[27446]_ , \new_[27447]_ , \new_[27448]_ ,
    \new_[27449]_ , \new_[27450]_ , \new_[27451]_ , \new_[27452]_ ,
    \new_[27453]_ , \new_[27454]_ , \new_[27455]_ , \new_[27456]_ ,
    \new_[27457]_ , \new_[27458]_ , \new_[27459]_ , \new_[27460]_ ,
    \new_[27461]_ , \new_[27462]_ , \new_[27463]_ , \new_[27464]_ ,
    \new_[27465]_ , \new_[27466]_ , \new_[27467]_ , \new_[27468]_ ,
    \new_[27469]_ , \new_[27470]_ , \new_[27471]_ , \new_[27472]_ ,
    \new_[27473]_ , \new_[27474]_ , \new_[27475]_ , \new_[27476]_ ,
    \new_[27477]_ , \new_[27478]_ , \new_[27479]_ , \new_[27480]_ ,
    \new_[27481]_ , \new_[27482]_ , \new_[27483]_ , \new_[27484]_ ,
    \new_[27485]_ , \new_[27486]_ , \new_[27487]_ , \new_[27488]_ ,
    \new_[27489]_ , \new_[27490]_ , \new_[27491]_ , \new_[27492]_ ,
    \new_[27493]_ , \new_[27494]_ , \new_[27495]_ , \new_[27496]_ ,
    \new_[27497]_ , \new_[27498]_ , \new_[27499]_ , \new_[27500]_ ,
    \new_[27501]_ , \new_[27502]_ , \new_[27503]_ , \new_[27504]_ ,
    \new_[27505]_ , \new_[27506]_ , \new_[27507]_ , \new_[27508]_ ,
    \new_[27509]_ , \new_[27510]_ , \new_[27511]_ , \new_[27512]_ ,
    \new_[27513]_ , \new_[27514]_ , \new_[27515]_ , \new_[27516]_ ,
    \new_[27517]_ , \new_[27518]_ , \new_[27519]_ , \new_[27520]_ ,
    \new_[27521]_ , \new_[27522]_ , \new_[27523]_ , \new_[27524]_ ,
    \new_[27525]_ , \new_[27526]_ , \new_[27527]_ , \new_[27528]_ ,
    \new_[27529]_ , \new_[27530]_ , \new_[27531]_ , \new_[27532]_ ,
    \new_[27533]_ , \new_[27534]_ , \new_[27535]_ , \new_[27536]_ ,
    \new_[27537]_ , \new_[27538]_ , \new_[27539]_ , \new_[27540]_ ,
    \new_[27541]_ , \new_[27542]_ , \new_[27543]_ , \new_[27544]_ ,
    \new_[27545]_ , \new_[27546]_ , \new_[27547]_ , \new_[27548]_ ,
    \new_[27549]_ , \new_[27550]_ , \new_[27551]_ , \new_[27552]_ ,
    \new_[27553]_ , \new_[27554]_ , \new_[27555]_ , \new_[27556]_ ,
    \new_[27557]_ , \new_[27558]_ , \new_[27559]_ , \new_[27560]_ ,
    \new_[27561]_ , \new_[27562]_ , \new_[27563]_ , \new_[27564]_ ,
    \new_[27565]_ , \new_[27566]_ , \new_[27567]_ , \new_[27568]_ ,
    \new_[27569]_ , \new_[27570]_ , \new_[27571]_ , \new_[27572]_ ,
    \new_[27573]_ , \new_[27574]_ , \new_[27575]_ , \new_[27576]_ ,
    \new_[27577]_ , \new_[27578]_ , \new_[27579]_ , \new_[27580]_ ,
    \new_[27581]_ , \new_[27582]_ , \new_[27583]_ , \new_[27584]_ ,
    \new_[27585]_ , \new_[27586]_ , \new_[27587]_ , \new_[27588]_ ,
    \new_[27589]_ , \new_[27590]_ , \new_[27591]_ , \new_[27592]_ ,
    \new_[27593]_ , \new_[27594]_ , \new_[27595]_ , \new_[27596]_ ,
    \new_[27597]_ , \new_[27598]_ , \new_[27599]_ , \new_[27600]_ ,
    \new_[27601]_ , \new_[27602]_ , \new_[27603]_ , \new_[27604]_ ,
    \new_[27605]_ , \new_[27606]_ , \new_[27607]_ , \new_[27608]_ ,
    \new_[27609]_ , \new_[27610]_ , \new_[27611]_ , \new_[27612]_ ,
    \new_[27613]_ , \new_[27614]_ , \new_[27615]_ , \new_[27616]_ ,
    \new_[27617]_ , \new_[27618]_ , \new_[27619]_ , \new_[27620]_ ,
    \new_[27621]_ , \new_[27622]_ , \new_[27623]_ , \new_[27624]_ ,
    \new_[27625]_ , \new_[27626]_ , \new_[27627]_ , \new_[27628]_ ,
    \new_[27629]_ , \new_[27630]_ , \new_[27631]_ , \new_[27632]_ ,
    \new_[27633]_ , \new_[27634]_ , \new_[27635]_ , \new_[27636]_ ,
    \new_[27637]_ , \new_[27638]_ , \new_[27639]_ , \new_[27640]_ ,
    \new_[27641]_ , \new_[27642]_ , \new_[27643]_ , \new_[27644]_ ,
    \new_[27645]_ , \new_[27646]_ , \new_[27647]_ , \new_[27648]_ ,
    \new_[27649]_ , \new_[27650]_ , \new_[27651]_ , \new_[27652]_ ,
    \new_[27653]_ , \new_[27654]_ , \new_[27655]_ , \new_[27656]_ ,
    \new_[27657]_ , \new_[27658]_ , \new_[27659]_ , \new_[27660]_ ,
    \new_[27661]_ , \new_[27662]_ , \new_[27663]_ , \new_[27664]_ ,
    \new_[27665]_ , \new_[27666]_ , \new_[27667]_ , \new_[27668]_ ,
    \new_[27669]_ , \new_[27670]_ , \new_[27671]_ , \new_[27672]_ ,
    \new_[27673]_ , \new_[27674]_ , \new_[27675]_ , \new_[27676]_ ,
    \new_[27677]_ , \new_[27678]_ , \new_[27679]_ , \new_[27680]_ ,
    \new_[27681]_ , \new_[27682]_ , \new_[27683]_ , \new_[27684]_ ,
    \new_[27685]_ , \new_[27686]_ , \new_[27687]_ , \new_[27688]_ ,
    \new_[27689]_ , \new_[27690]_ , \new_[27691]_ , \new_[27692]_ ,
    \new_[27693]_ , \new_[27694]_ , \new_[27695]_ , \new_[27696]_ ,
    \new_[27697]_ , \new_[27698]_ , \new_[27699]_ , \new_[27700]_ ,
    \new_[27701]_ , \new_[27702]_ , \new_[27703]_ , \new_[27704]_ ,
    \new_[27705]_ , \new_[27706]_ , \new_[27707]_ , \new_[27708]_ ,
    \new_[27709]_ , \new_[27710]_ , \new_[27711]_ , \new_[27712]_ ,
    \new_[27713]_ , \new_[27714]_ , \new_[27715]_ , \new_[27716]_ ,
    \new_[27717]_ , \new_[27718]_ , \new_[27719]_ , \new_[27720]_ ,
    \new_[27721]_ , \new_[27722]_ , \new_[27723]_ , \new_[27724]_ ,
    \new_[27725]_ , \new_[27726]_ , \new_[27727]_ , \new_[27728]_ ,
    \new_[27729]_ , \new_[27730]_ , \new_[27731]_ , \new_[27732]_ ,
    \new_[27733]_ , \new_[27734]_ , \new_[27735]_ , \new_[27736]_ ,
    \new_[27737]_ , \new_[27738]_ , \new_[27739]_ , \new_[27740]_ ,
    \new_[27741]_ , \new_[27742]_ , \new_[27743]_ , \new_[27744]_ ,
    \new_[27745]_ , \new_[27746]_ , \new_[27747]_ , \new_[27748]_ ,
    \new_[27749]_ , \new_[27750]_ , \new_[27751]_ , \new_[27752]_ ,
    \new_[27753]_ , \new_[27754]_ , \new_[27755]_ , \new_[27756]_ ,
    \new_[27757]_ , \new_[27758]_ , \new_[27759]_ , \new_[27760]_ ,
    \new_[27761]_ , \new_[27762]_ , \new_[27763]_ , \new_[27764]_ ,
    \new_[27765]_ , \new_[27766]_ , \new_[27767]_ , \new_[27768]_ ,
    \new_[27769]_ , \new_[27770]_ , \new_[27771]_ , \new_[27772]_ ,
    \new_[27773]_ , \new_[27774]_ , \new_[27775]_ , \new_[27776]_ ,
    \new_[27777]_ , \new_[27778]_ , \new_[27779]_ , \new_[27780]_ ,
    \new_[27781]_ , \new_[27782]_ , \new_[27783]_ , \new_[27784]_ ,
    \new_[27785]_ , \new_[27786]_ , \new_[27787]_ , \new_[27788]_ ,
    \new_[27789]_ , \new_[27790]_ , \new_[27791]_ , \new_[27792]_ ,
    \new_[27793]_ , \new_[27794]_ , \new_[27795]_ , \new_[27796]_ ,
    \new_[27797]_ , \new_[27798]_ , \new_[27799]_ , \new_[27800]_ ,
    \new_[27801]_ , \new_[27802]_ , \new_[27803]_ , \new_[27804]_ ,
    \new_[27805]_ , \new_[27806]_ , \new_[27807]_ , \new_[27808]_ ,
    \new_[27809]_ , \new_[27810]_ , \new_[27811]_ , \new_[27812]_ ,
    \new_[27813]_ , \new_[27814]_ , \new_[27815]_ , \new_[27816]_ ,
    \new_[27817]_ , \new_[27818]_ , \new_[27819]_ , \new_[27820]_ ,
    \new_[27821]_ , \new_[27822]_ , \new_[27823]_ , \new_[27824]_ ,
    \new_[27825]_ , \new_[27826]_ , \new_[27827]_ , \new_[27828]_ ,
    \new_[27829]_ , \new_[27830]_ , \new_[27831]_ , \new_[27832]_ ,
    \new_[27833]_ , \new_[27834]_ , \new_[27835]_ , \new_[27836]_ ,
    \new_[27837]_ , \new_[27838]_ , \new_[27839]_ , \new_[27840]_ ,
    \new_[27841]_ , \new_[27842]_ , \new_[27843]_ , \new_[27844]_ ,
    \new_[27845]_ , \new_[27846]_ , \new_[27847]_ , \new_[27848]_ ,
    \new_[27849]_ , \new_[27850]_ , \new_[27851]_ , \new_[27852]_ ,
    \new_[27853]_ , \new_[27854]_ , \new_[27855]_ , \new_[27856]_ ,
    \new_[27857]_ , \new_[27858]_ , \new_[27859]_ , \new_[27860]_ ,
    \new_[27861]_ , \new_[27862]_ , \new_[27863]_ , \new_[27864]_ ,
    \new_[27865]_ , \new_[27866]_ , \new_[27867]_ , \new_[27868]_ ,
    \new_[27869]_ , \new_[27870]_ , \new_[27871]_ , \new_[27872]_ ,
    \new_[27873]_ , \new_[27874]_ , \new_[27875]_ , \new_[27876]_ ,
    \new_[27877]_ , \new_[27878]_ , \new_[27879]_ , \new_[27880]_ ,
    \new_[27881]_ , \new_[27882]_ , \new_[27883]_ , \new_[27884]_ ,
    \new_[27885]_ , \new_[27886]_ , \new_[27887]_ , \new_[27888]_ ,
    \new_[27889]_ , \new_[27890]_ , \new_[27891]_ , \new_[27892]_ ,
    \new_[27893]_ , \new_[27894]_ , \new_[27895]_ , \new_[27896]_ ,
    \new_[27897]_ , \new_[27898]_ , \new_[27899]_ , \new_[27900]_ ,
    \new_[27901]_ , \new_[27902]_ , \new_[27903]_ , \new_[27904]_ ,
    \new_[27905]_ , \new_[27906]_ , \new_[27907]_ , \new_[27908]_ ,
    \new_[27909]_ , \new_[27910]_ , \new_[27911]_ , \new_[27912]_ ,
    \new_[27913]_ , \new_[27914]_ , \new_[27915]_ , \new_[27916]_ ,
    \new_[27917]_ , \new_[27918]_ , \new_[27919]_ , \new_[27920]_ ,
    \new_[27921]_ , \new_[27922]_ , \new_[27923]_ , \new_[27924]_ ,
    \new_[27925]_ , \new_[27926]_ , \new_[27927]_ , \new_[27928]_ ,
    \new_[27929]_ , \new_[27930]_ , \new_[27931]_ , \new_[27932]_ ,
    \new_[27933]_ , \new_[27934]_ , \new_[27935]_ , \new_[27936]_ ,
    \new_[27937]_ , \new_[27938]_ , \new_[27939]_ , \new_[27940]_ ,
    \new_[27941]_ , \new_[27942]_ , \new_[27943]_ , \new_[27944]_ ,
    \new_[27945]_ , \new_[27946]_ , \new_[27947]_ , \new_[27948]_ ,
    \new_[27949]_ , \new_[27950]_ , \new_[27951]_ , \new_[27952]_ ,
    \new_[27953]_ , \new_[27954]_ , \new_[27955]_ , \new_[27956]_ ,
    \new_[27957]_ , \new_[27958]_ , \new_[27959]_ , \new_[27960]_ ,
    \new_[27961]_ , \new_[27962]_ , \new_[27963]_ , \new_[27964]_ ,
    \new_[27965]_ , \new_[27966]_ , \new_[27967]_ , \new_[27968]_ ,
    \new_[27969]_ , \new_[27970]_ , \new_[27971]_ , \new_[27972]_ ,
    \new_[27973]_ , \new_[27974]_ , \new_[27975]_ , \new_[27976]_ ,
    \new_[27977]_ , \new_[27978]_ , \new_[27979]_ , \new_[27980]_ ,
    \new_[27981]_ , \new_[27982]_ , \new_[27983]_ , \new_[27984]_ ,
    \new_[27985]_ , \new_[27986]_ , \new_[27987]_ , \new_[27988]_ ,
    \new_[27989]_ , \new_[27990]_ , \new_[27991]_ , \new_[27992]_ ,
    \new_[27993]_ , \new_[27994]_ , \new_[27995]_ , \new_[27996]_ ,
    \new_[27997]_ , \new_[27998]_ , \new_[27999]_ , \new_[28000]_ ,
    \new_[28001]_ , \new_[28002]_ , \new_[28003]_ , \new_[28004]_ ,
    \new_[28005]_ , \new_[28006]_ , \new_[28007]_ , \new_[28008]_ ,
    \new_[28009]_ , \new_[28010]_ , \new_[28011]_ , \new_[28012]_ ,
    \new_[28013]_ , \new_[28014]_ , \new_[28015]_ , \new_[28016]_ ,
    \new_[28017]_ , \new_[28018]_ , \new_[28019]_ , \new_[28020]_ ,
    \new_[28021]_ , \new_[28022]_ , \new_[28023]_ , \new_[28024]_ ,
    \new_[28025]_ , \new_[28026]_ , \new_[28027]_ , \new_[28028]_ ,
    \new_[28029]_ , \new_[28030]_ , \new_[28031]_ , \new_[28032]_ ,
    \new_[28033]_ , \new_[28034]_ , \new_[28035]_ , \new_[28036]_ ,
    \new_[28037]_ , \new_[28038]_ , \new_[28039]_ , \new_[28040]_ ,
    \new_[28041]_ , \new_[28042]_ , \new_[28043]_ , \new_[28044]_ ,
    \new_[28045]_ , \new_[28046]_ , \new_[28047]_ , \new_[28048]_ ,
    \new_[28049]_ , \new_[28050]_ , \new_[28051]_ , \new_[28052]_ ,
    \new_[28053]_ , \new_[28054]_ , \new_[28055]_ , \new_[28056]_ ,
    \new_[28057]_ , \new_[28058]_ , \new_[28059]_ , \new_[28060]_ ,
    \new_[28061]_ , \new_[28062]_ , \new_[28063]_ , \new_[28064]_ ,
    \new_[28065]_ , \new_[28066]_ , \new_[28067]_ , \new_[28068]_ ,
    \new_[28069]_ , \new_[28070]_ , \new_[28071]_ , \new_[28072]_ ,
    \new_[28073]_ , \new_[28074]_ , \new_[28075]_ , \new_[28076]_ ,
    \new_[28077]_ , \new_[28078]_ , \new_[28079]_ , \new_[28080]_ ,
    \new_[28081]_ , \new_[28082]_ , \new_[28083]_ , \new_[28084]_ ,
    \new_[28085]_ , \new_[28086]_ , \new_[28087]_ , \new_[28088]_ ,
    \new_[28089]_ , \new_[28090]_ , \new_[28091]_ , \new_[28092]_ ,
    \new_[28093]_ , \new_[28094]_ , \new_[28095]_ , \new_[28096]_ ,
    \new_[28097]_ , \new_[28098]_ , \new_[28099]_ , \new_[28100]_ ,
    \new_[28101]_ , \new_[28102]_ , \new_[28103]_ , \new_[28104]_ ,
    \new_[28105]_ , \new_[28106]_ , \new_[28107]_ , \new_[28108]_ ,
    \new_[28109]_ , \new_[28110]_ , \new_[28111]_ , \new_[28112]_ ,
    \new_[28113]_ , \new_[28114]_ , \new_[28115]_ , \new_[28116]_ ,
    \new_[28117]_ , \new_[28118]_ , \new_[28119]_ , \new_[28120]_ ,
    \new_[28121]_ , \new_[28122]_ , \new_[28123]_ , \new_[28124]_ ,
    \new_[28125]_ , \new_[28126]_ , \new_[28127]_ , \new_[28128]_ ,
    \new_[28129]_ , \new_[28130]_ , \new_[28131]_ , \new_[28132]_ ,
    \new_[28133]_ , \new_[28134]_ , \new_[28135]_ , \new_[28136]_ ,
    \new_[28137]_ , \new_[28138]_ , \new_[28139]_ , \new_[28140]_ ,
    \new_[28141]_ , \new_[28142]_ , \new_[28143]_ , \new_[28144]_ ,
    \new_[28145]_ , \new_[28146]_ , \new_[28147]_ , \new_[28148]_ ,
    \new_[28149]_ , \new_[28150]_ , \new_[28151]_ , \new_[28152]_ ,
    \new_[28153]_ , \new_[28154]_ , \new_[28155]_ , \new_[28156]_ ,
    \new_[28157]_ , \new_[28158]_ , \new_[28159]_ , \new_[28160]_ ,
    \new_[28161]_ , \new_[28162]_ , \new_[28163]_ , \new_[28164]_ ,
    \new_[28165]_ , \new_[28166]_ , \new_[28167]_ , \new_[28168]_ ,
    \new_[28169]_ , \new_[28170]_ , \new_[28171]_ , \new_[28172]_ ,
    \new_[28173]_ , \new_[28174]_ , \new_[28175]_ , \new_[28176]_ ,
    \new_[28177]_ , \new_[28178]_ , \new_[28179]_ , \new_[28180]_ ,
    \new_[28181]_ , \new_[28182]_ , \new_[28183]_ , \new_[28184]_ ,
    \new_[28185]_ , \new_[28186]_ , \new_[28187]_ , \new_[28188]_ ,
    \new_[28189]_ , \new_[28190]_ , \new_[28191]_ , \new_[28192]_ ,
    \new_[28193]_ , \new_[28194]_ , \new_[28195]_ , \new_[28196]_ ,
    \new_[28197]_ , \new_[28198]_ , \new_[28199]_ , \new_[28200]_ ,
    \new_[28201]_ , \new_[28202]_ , \new_[28203]_ , \new_[28204]_ ,
    \new_[28205]_ , \new_[28206]_ , \new_[28207]_ , \new_[28208]_ ,
    \new_[28209]_ , \new_[28210]_ , \new_[28211]_ , \new_[28212]_ ,
    \new_[28213]_ , \new_[28214]_ , \new_[28215]_ , \new_[28216]_ ,
    \new_[28217]_ , \new_[28218]_ , \new_[28219]_ , \new_[28220]_ ,
    \new_[28221]_ , \new_[28222]_ , \new_[28223]_ , \new_[28224]_ ,
    \new_[28225]_ , \new_[28226]_ , \new_[28227]_ , \new_[28228]_ ,
    \new_[28229]_ , \new_[28230]_ , \new_[28231]_ , \new_[28232]_ ,
    \new_[28233]_ , \new_[28234]_ , \new_[28235]_ , \new_[28236]_ ,
    \new_[28237]_ , \new_[28238]_ , \new_[28239]_ , \new_[28240]_ ,
    \new_[28241]_ , \new_[28242]_ , \new_[28243]_ , \new_[28244]_ ,
    \new_[28245]_ , \new_[28246]_ , \new_[28247]_ , \new_[28248]_ ,
    \new_[28249]_ , \new_[28250]_ , \new_[28251]_ , \new_[28252]_ ,
    \new_[28253]_ , \new_[28254]_ , \new_[28255]_ , \new_[28256]_ ,
    \new_[28257]_ , \new_[28258]_ , \new_[28259]_ , \new_[28260]_ ,
    \new_[28261]_ , \new_[28262]_ , \new_[28263]_ , \new_[28264]_ ,
    \new_[28265]_ , \new_[28266]_ , \new_[28267]_ , \new_[28268]_ ,
    \new_[28269]_ , \new_[28270]_ , \new_[28271]_ , \new_[28272]_ ,
    \new_[28273]_ , \new_[28274]_ , \new_[28275]_ , \new_[28276]_ ,
    \new_[28277]_ , \new_[28278]_ , \new_[28279]_ , \new_[28280]_ ,
    \new_[28281]_ , \new_[28282]_ , \new_[28283]_ , \new_[28284]_ ,
    \new_[28285]_ , \new_[28286]_ , \new_[28287]_ , \new_[28288]_ ,
    \new_[28289]_ , \new_[28290]_ , \new_[28291]_ , \new_[28292]_ ,
    \new_[28293]_ , \new_[28294]_ , \new_[28295]_ , \new_[28296]_ ,
    \new_[28297]_ , \new_[28298]_ , \new_[28299]_ , \new_[28300]_ ,
    \new_[28301]_ , \new_[28302]_ , \new_[28303]_ , \new_[28304]_ ,
    \new_[28305]_ , \new_[28306]_ , \new_[28307]_ , \new_[28308]_ ,
    \new_[28309]_ , \new_[28310]_ , \new_[28311]_ , \new_[28312]_ ,
    \new_[28313]_ , \new_[28314]_ , \new_[28315]_ , \new_[28316]_ ,
    \new_[28317]_ , \new_[28318]_ , \new_[28319]_ , \new_[28320]_ ,
    \new_[28321]_ , \new_[28322]_ , \new_[28323]_ , \new_[28324]_ ,
    \new_[28325]_ , \new_[28326]_ , \new_[28327]_ , \new_[28328]_ ,
    \new_[28329]_ , \new_[28330]_ , \new_[28331]_ , \new_[28332]_ ,
    \new_[28333]_ , \new_[28334]_ , \new_[28335]_ , \new_[28336]_ ,
    \new_[28337]_ , \new_[28338]_ , \new_[28339]_ , \new_[28340]_ ,
    \new_[28341]_ , \new_[28342]_ , \new_[28343]_ , \new_[28344]_ ,
    \new_[28345]_ , \new_[28346]_ , \new_[28347]_ , \new_[28348]_ ,
    \new_[28349]_ , \new_[28350]_ , \new_[28351]_ , \new_[28352]_ ,
    \new_[28353]_ , \new_[28354]_ , \new_[28355]_ , \new_[28356]_ ,
    \new_[28357]_ , \new_[28358]_ , \new_[28359]_ , \new_[28360]_ ,
    \new_[28361]_ , \new_[28362]_ , \new_[28363]_ , \new_[28364]_ ,
    \new_[28365]_ , \new_[28366]_ , \new_[28367]_ , \new_[28368]_ ,
    \new_[28369]_ , \new_[28370]_ , \new_[28371]_ , \new_[28372]_ ,
    \new_[28373]_ , \new_[28374]_ , \new_[28375]_ , \new_[28376]_ ,
    \new_[28377]_ , \new_[28378]_ , \new_[28379]_ , \new_[28380]_ ,
    \new_[28381]_ , \new_[28382]_ , \new_[28383]_ , \new_[28384]_ ,
    \new_[28385]_ , \new_[28386]_ , \new_[28387]_ , \new_[28388]_ ,
    \new_[28389]_ , \new_[28390]_ , \new_[28391]_ , \new_[28392]_ ,
    \new_[28393]_ , \new_[28394]_ , \new_[28395]_ , \new_[28396]_ ,
    \new_[28397]_ , \new_[28398]_ , \new_[28399]_ , \new_[28400]_ ,
    \new_[28401]_ , \new_[28402]_ , \new_[28403]_ , \new_[28404]_ ,
    \new_[28405]_ , \new_[28406]_ , \new_[28407]_ , \new_[28408]_ ,
    \new_[28409]_ , \new_[28410]_ , \new_[28411]_ , \new_[28412]_ ,
    \new_[28413]_ , \new_[28414]_ , \new_[28415]_ , \new_[28416]_ ,
    \new_[28417]_ , \new_[28418]_ , \new_[28419]_ , \new_[28420]_ ,
    \new_[28421]_ , \new_[28422]_ , \new_[28423]_ , \new_[28424]_ ,
    \new_[28425]_ , \new_[28426]_ , \new_[28427]_ , \new_[28428]_ ,
    \new_[28429]_ , \new_[28430]_ , \new_[28431]_ , \new_[28432]_ ,
    \new_[28433]_ , \new_[28434]_ , \new_[28435]_ , \new_[28436]_ ,
    \new_[28437]_ , \new_[28438]_ , \new_[28439]_ , \new_[28440]_ ,
    \new_[28441]_ , \new_[28442]_ , \new_[28443]_ , \new_[28444]_ ,
    \new_[28445]_ , \new_[28446]_ , \new_[28447]_ , \new_[28448]_ ,
    \new_[28449]_ , \new_[28450]_ , \new_[28451]_ , \new_[28452]_ ,
    \new_[28453]_ , \new_[28454]_ , \new_[28455]_ , \new_[28456]_ ,
    \new_[28457]_ , \new_[28458]_ , \new_[28459]_ , \new_[28460]_ ,
    \new_[28461]_ , \new_[28462]_ , \new_[28463]_ , \new_[28464]_ ,
    \new_[28465]_ , \new_[28466]_ , \new_[28467]_ , \new_[28468]_ ,
    \new_[28469]_ , \new_[28470]_ , \new_[28471]_ , \new_[28472]_ ,
    \new_[28473]_ , \new_[28474]_ , \new_[28475]_ , \new_[28476]_ ,
    \new_[28477]_ , \new_[28478]_ , \new_[28479]_ , \new_[28480]_ ,
    \new_[28481]_ , \new_[28482]_ , \new_[28483]_ , \new_[28484]_ ,
    \new_[28485]_ , \new_[28486]_ , \new_[28487]_ , \new_[28488]_ ,
    \new_[28489]_ , \new_[28490]_ , \new_[28491]_ , \new_[28492]_ ,
    \new_[28493]_ , \new_[28494]_ , \new_[28495]_ , \new_[28496]_ ,
    \new_[28497]_ , \new_[28498]_ , \new_[28499]_ , \new_[28500]_ ,
    \new_[28501]_ , \new_[28502]_ , \new_[28503]_ , \new_[28504]_ ,
    \new_[28505]_ , \new_[28506]_ , \new_[28507]_ , \new_[28508]_ ,
    \new_[28509]_ , \new_[28510]_ , \new_[28511]_ , \new_[28512]_ ,
    \new_[28513]_ , \new_[28514]_ , \new_[28515]_ , \new_[28516]_ ,
    \new_[28517]_ , \new_[28518]_ , \new_[28519]_ , \new_[28520]_ ,
    \new_[28521]_ , \new_[28522]_ , \new_[28523]_ , \new_[28524]_ ,
    \new_[28525]_ , \new_[28526]_ , \new_[28527]_ , \new_[28528]_ ,
    \new_[28529]_ , \new_[28530]_ , \new_[28531]_ , \new_[28532]_ ,
    \new_[28533]_ , \new_[28534]_ , \new_[28535]_ , \new_[28536]_ ,
    \new_[28537]_ , \new_[28538]_ , \new_[28539]_ , \new_[28540]_ ,
    \new_[28541]_ , \new_[28542]_ , \new_[28543]_ , \new_[28544]_ ,
    \new_[28545]_ , \new_[28546]_ , \new_[28547]_ , \new_[28548]_ ,
    \new_[28549]_ , \new_[28550]_ , \new_[28551]_ , \new_[28552]_ ,
    \new_[28553]_ , \new_[28554]_ , \new_[28555]_ , \new_[28556]_ ,
    \new_[28557]_ , \new_[28558]_ , \new_[28559]_ , \new_[28560]_ ,
    \new_[28561]_ , \new_[28562]_ , \new_[28563]_ , \new_[28564]_ ,
    \new_[28565]_ , \new_[28566]_ , \new_[28567]_ , \new_[28568]_ ,
    \new_[28569]_ , \new_[28570]_ , \new_[28571]_ , \new_[28572]_ ,
    \new_[28573]_ , \new_[28574]_ , \new_[28575]_ , \new_[28576]_ ,
    \new_[28577]_ , \new_[28578]_ , \new_[28579]_ , \new_[28580]_ ,
    \new_[28581]_ , \new_[28582]_ , \new_[28583]_ , \new_[28584]_ ,
    \new_[28585]_ , \new_[28586]_ , \new_[28587]_ , \new_[28588]_ ,
    \new_[28589]_ , \new_[28590]_ , \new_[28591]_ , \new_[28592]_ ,
    \new_[28593]_ , \new_[28594]_ , \new_[28595]_ , \new_[28596]_ ,
    \new_[28597]_ , \new_[28598]_ , \new_[28599]_ , \new_[28600]_ ,
    \new_[28601]_ , \new_[28602]_ , \new_[28603]_ , \new_[28604]_ ,
    \new_[28605]_ , \new_[28606]_ , \new_[28607]_ , \new_[28608]_ ,
    \new_[28609]_ , \new_[28610]_ , \new_[28611]_ , \new_[28612]_ ,
    \new_[28613]_ , \new_[28614]_ , \new_[28615]_ , \new_[28616]_ ,
    \new_[28617]_ , \new_[28618]_ , \new_[28619]_ , \new_[28620]_ ,
    \new_[28621]_ , \new_[28622]_ , \new_[28623]_ , \new_[28624]_ ,
    \new_[28625]_ , \new_[28626]_ , \new_[28627]_ , \new_[28628]_ ,
    \new_[28629]_ , \new_[28630]_ , \new_[28631]_ , \new_[28632]_ ,
    \new_[28633]_ , \new_[28634]_ , \new_[28635]_ , \new_[28636]_ ,
    \new_[28637]_ , \new_[28638]_ , \new_[28639]_ , \new_[28640]_ ,
    \new_[28641]_ , \new_[28642]_ , \new_[28643]_ , \new_[28644]_ ,
    \new_[28645]_ , \new_[28646]_ , \new_[28647]_ , \new_[28648]_ ,
    \new_[28649]_ , \new_[28650]_ , \new_[28651]_ , \new_[28652]_ ,
    \new_[28653]_ , \new_[28654]_ , \new_[28655]_ , \new_[28656]_ ,
    \new_[28657]_ , \new_[28658]_ , \new_[28659]_ , \new_[28660]_ ,
    \new_[28661]_ , \new_[28662]_ , \new_[28663]_ , \new_[28664]_ ,
    \new_[28665]_ , \new_[28666]_ , \new_[28667]_ , \new_[28668]_ ,
    \new_[28669]_ , \new_[28670]_ , \new_[28671]_ , \new_[28672]_ ,
    \new_[28673]_ , \new_[28674]_ , \new_[28675]_ , \new_[28676]_ ,
    \new_[28677]_ , \new_[28678]_ , \new_[28679]_ , \new_[28680]_ ,
    \new_[28681]_ , \new_[28682]_ , \new_[28683]_ , \new_[28684]_ ,
    \new_[28685]_ , \new_[28686]_ , \new_[28687]_ , \new_[28688]_ ,
    \new_[28689]_ , \new_[28690]_ , \new_[28691]_ , \new_[28692]_ ,
    \new_[28693]_ , \new_[28694]_ , \new_[28695]_ , \new_[28696]_ ,
    \new_[28697]_ , \new_[28698]_ , \new_[28699]_ , \new_[28700]_ ,
    \new_[28701]_ , \new_[28702]_ , \new_[28703]_ , \new_[28704]_ ,
    \new_[28705]_ , \new_[28706]_ , \new_[28707]_ , \new_[28708]_ ,
    \new_[28709]_ , \new_[28710]_ , \new_[28711]_ , \new_[28712]_ ,
    \new_[28713]_ , \new_[28714]_ , \new_[28715]_ , \new_[28716]_ ,
    \new_[28717]_ , \new_[28718]_ , \new_[28719]_ , \new_[28720]_ ,
    \new_[28721]_ , \new_[28722]_ , \new_[28723]_ , \new_[28724]_ ,
    \new_[28725]_ , \new_[28726]_ , \new_[28727]_ , \new_[28728]_ ,
    \new_[28729]_ , \new_[28730]_ , \new_[28731]_ , \new_[28732]_ ,
    \new_[28733]_ , \new_[28734]_ , \new_[28735]_ , \new_[28736]_ ,
    \new_[28737]_ , \new_[28738]_ , \new_[28739]_ , \new_[28740]_ ,
    \new_[28741]_ , \new_[28742]_ , \new_[28743]_ , \new_[28744]_ ,
    \new_[28745]_ , \new_[28746]_ , \new_[28747]_ , \new_[28748]_ ,
    \new_[28749]_ , \new_[28750]_ , \new_[28751]_ , \new_[28752]_ ,
    \new_[28753]_ , \new_[28754]_ , \new_[28755]_ , \new_[28756]_ ,
    \new_[28757]_ , \new_[28758]_ , \new_[28759]_ , \new_[28760]_ ,
    \new_[28761]_ , \new_[28762]_ , \new_[28763]_ , \new_[28764]_ ,
    \new_[28765]_ , \new_[28766]_ , \new_[28767]_ , \new_[28768]_ ,
    \new_[28769]_ , \new_[28770]_ , \new_[28771]_ , \new_[28772]_ ,
    \new_[28773]_ , \new_[28774]_ , \new_[28775]_ , \new_[28776]_ ,
    \new_[28777]_ , \new_[28778]_ , \new_[28779]_ , \new_[28780]_ ,
    \new_[28781]_ , \new_[28782]_ , \new_[28783]_ , \new_[28784]_ ,
    \new_[28785]_ , \new_[28786]_ , \new_[28787]_ , \new_[28788]_ ,
    \new_[28789]_ , \new_[28790]_ , \new_[28791]_ , \new_[28792]_ ,
    \new_[28793]_ , \new_[28794]_ , \new_[28795]_ , \new_[28796]_ ,
    \new_[28797]_ , \new_[28798]_ , \new_[28799]_ , \new_[28800]_ ,
    \new_[28801]_ , \new_[28802]_ , \new_[28803]_ , \new_[28804]_ ,
    \new_[28805]_ , \new_[28806]_ , \new_[28807]_ , \new_[28808]_ ,
    \new_[28809]_ , \new_[28810]_ , \new_[28811]_ , \new_[28812]_ ,
    \new_[28813]_ , \new_[28814]_ , \new_[28815]_ , \new_[28816]_ ,
    \new_[28817]_ , \new_[28818]_ , \new_[28819]_ , \new_[28820]_ ,
    \new_[28821]_ , \new_[28822]_ , \new_[28823]_ , \new_[28824]_ ,
    \new_[28825]_ , \new_[28826]_ , \new_[28827]_ , \new_[28828]_ ,
    \new_[28829]_ , \new_[28830]_ , \new_[28831]_ , \new_[28832]_ ,
    \new_[28833]_ , \new_[28834]_ , \new_[28835]_ , \new_[28836]_ ,
    \new_[28837]_ , \new_[28838]_ , \new_[28839]_ , \new_[28840]_ ,
    \new_[28841]_ , \new_[28842]_ , \new_[28843]_ , \new_[28844]_ ,
    \new_[28845]_ , \new_[28846]_ , \new_[28847]_ , \new_[28848]_ ,
    \new_[28849]_ , \new_[28850]_ , \new_[28851]_ , \new_[28852]_ ,
    \new_[28853]_ , \new_[28854]_ , \new_[28855]_ , \new_[28856]_ ,
    \new_[28857]_ , \new_[28858]_ , \new_[28859]_ , \new_[28860]_ ,
    \new_[28861]_ , \new_[28862]_ , \new_[28863]_ , \new_[28864]_ ,
    \new_[28865]_ , \new_[28866]_ , \new_[28867]_ , \new_[28868]_ ,
    \new_[28869]_ , \new_[28870]_ , \new_[28871]_ , \new_[28872]_ ,
    \new_[28873]_ , \new_[28874]_ , \new_[28875]_ , \new_[28876]_ ,
    \new_[28877]_ , \new_[28878]_ , \new_[28879]_ , \new_[28880]_ ,
    \new_[28881]_ , \new_[28882]_ , \new_[28883]_ , \new_[28884]_ ,
    \new_[28885]_ , \new_[28886]_ , \new_[28887]_ , \new_[28888]_ ,
    \new_[28889]_ , \new_[28890]_ , \new_[28891]_ , \new_[28892]_ ,
    \new_[28893]_ , \new_[28894]_ , \new_[28895]_ , \new_[28896]_ ,
    \new_[28897]_ , \new_[28898]_ , \new_[28899]_ , \new_[28900]_ ,
    \new_[28901]_ , \new_[28902]_ , \new_[28903]_ , \new_[28904]_ ,
    \new_[28905]_ , \new_[28906]_ , \new_[28907]_ , \new_[28908]_ ,
    \new_[28909]_ , \new_[28910]_ , \new_[28911]_ , \new_[28912]_ ,
    \new_[28913]_ , \new_[28914]_ , \new_[28915]_ , \new_[28916]_ ,
    \new_[28917]_ , \new_[28918]_ , \new_[28919]_ , \new_[28920]_ ,
    \new_[28921]_ , \new_[28922]_ , \new_[28923]_ , \new_[28924]_ ,
    \new_[28925]_ , \new_[28926]_ , \new_[28927]_ , \new_[28928]_ ,
    \new_[28929]_ , \new_[28930]_ , \new_[28931]_ , \new_[28932]_ ,
    \new_[28933]_ , \new_[28934]_ , \new_[28935]_ , \new_[28936]_ ,
    \new_[28937]_ , \new_[28938]_ , \new_[28939]_ , \new_[28940]_ ,
    \new_[28941]_ , \new_[28942]_ , \new_[28943]_ , \new_[28944]_ ,
    \new_[28945]_ , \new_[28946]_ , \new_[28947]_ , \new_[28948]_ ,
    \new_[28949]_ , \new_[28950]_ , \new_[28951]_ , \new_[28952]_ ,
    \new_[28953]_ , \new_[28954]_ , \new_[28955]_ , \new_[28956]_ ,
    \new_[28957]_ , \new_[28958]_ , \new_[28959]_ , \new_[28960]_ ,
    \new_[28961]_ , \new_[28962]_ , \new_[28963]_ , \new_[28964]_ ,
    \new_[28965]_ , \new_[28966]_ , \new_[28967]_ , \new_[28968]_ ,
    \new_[28969]_ , \new_[28970]_ , \new_[28971]_ , \new_[28972]_ ,
    \new_[28973]_ , \new_[28974]_ , \new_[28975]_ , \new_[28976]_ ,
    \new_[28977]_ , \new_[28978]_ , \new_[28979]_ , \new_[28980]_ ,
    \new_[28981]_ , \new_[28982]_ , \new_[28983]_ , \new_[28984]_ ,
    \new_[28985]_ , \new_[28986]_ , \new_[28987]_ , \new_[28988]_ ,
    \new_[28989]_ , \new_[28990]_ , \new_[28991]_ , \new_[28992]_ ,
    \new_[28993]_ , \new_[28994]_ , \new_[28995]_ , \new_[28996]_ ,
    \new_[28997]_ , \new_[28998]_ , \new_[28999]_ , \new_[29000]_ ,
    \new_[29001]_ , \new_[29002]_ , \new_[29003]_ , \new_[29004]_ ,
    \new_[29005]_ , \new_[29006]_ , \new_[29007]_ , \new_[29008]_ ,
    \new_[29009]_ , \new_[29010]_ , \new_[29011]_ , \new_[29012]_ ,
    \new_[29013]_ , \new_[29014]_ , \new_[29015]_ , \new_[29016]_ ,
    \new_[29017]_ , \new_[29018]_ , \new_[29019]_ , \new_[29020]_ ,
    \new_[29021]_ , \new_[29022]_ , \new_[29023]_ , \new_[29024]_ ,
    \new_[29025]_ , \new_[29026]_ , \new_[29027]_ , \new_[29028]_ ,
    \new_[29029]_ , \new_[29030]_ , \new_[29031]_ , \new_[29032]_ ,
    \new_[29033]_ , \new_[29034]_ , \new_[29035]_ , \new_[29036]_ ,
    \new_[29037]_ , \new_[29038]_ , \new_[29039]_ , \new_[29040]_ ,
    \new_[29041]_ , \new_[29042]_ , \new_[29043]_ , \new_[29044]_ ,
    \new_[29045]_ , \new_[29046]_ , \new_[29047]_ , \new_[29048]_ ,
    \new_[29049]_ , \new_[29050]_ , \new_[29051]_ , \new_[29052]_ ,
    \new_[29053]_ , \new_[29054]_ , \new_[29055]_ , \new_[29056]_ ,
    \new_[29057]_ , \new_[29058]_ , \new_[29059]_ , \new_[29060]_ ,
    \new_[29061]_ , \new_[29062]_ , \new_[29063]_ , \new_[29064]_ ,
    \new_[29065]_ , \new_[29066]_ , \new_[29067]_ , \new_[29068]_ ,
    \new_[29069]_ , \new_[29070]_ , \new_[29071]_ , \new_[29072]_ ,
    \new_[29073]_ , \new_[29074]_ , \new_[29075]_ , \new_[29076]_ ,
    \new_[29077]_ , \new_[29078]_ , \new_[29079]_ , \new_[29080]_ ,
    \new_[29081]_ , \new_[29082]_ , \new_[29083]_ , \new_[29084]_ ,
    \new_[29085]_ , \new_[29086]_ , \new_[29087]_ , \new_[29088]_ ,
    \new_[29089]_ , \new_[29090]_ , \new_[29091]_ , \new_[29092]_ ,
    \new_[29093]_ , \new_[29094]_ , \new_[29095]_ , \new_[29096]_ ,
    \new_[29097]_ , \new_[29098]_ , \new_[29099]_ , \new_[29100]_ ,
    \new_[29101]_ , \new_[29102]_ , \new_[29103]_ , \new_[29104]_ ,
    \new_[29105]_ , \new_[29106]_ , \new_[29107]_ , \new_[29108]_ ,
    \new_[29109]_ , \new_[29110]_ , \new_[29111]_ , \new_[29112]_ ,
    \new_[29113]_ , \new_[29114]_ , \new_[29115]_ , \new_[29116]_ ,
    \new_[29117]_ , \new_[29118]_ , \new_[29119]_ , \new_[29120]_ ,
    \new_[29121]_ , \new_[29122]_ , \new_[29123]_ , \new_[29124]_ ,
    \new_[29125]_ , \new_[29126]_ , \new_[29127]_ , \new_[29128]_ ,
    \new_[29129]_ , \new_[29130]_ , \new_[29131]_ , \new_[29132]_ ,
    \new_[29133]_ , \new_[29134]_ , \new_[29135]_ , \new_[29136]_ ,
    \new_[29137]_ , \new_[29138]_ , \new_[29139]_ , \new_[29140]_ ,
    \new_[29141]_ , \new_[29142]_ , \new_[29143]_ , \new_[29144]_ ,
    \new_[29145]_ , \new_[29146]_ , \new_[29147]_ , \new_[29148]_ ,
    \new_[29149]_ , \new_[29150]_ , \new_[29151]_ , \new_[29152]_ ,
    \new_[29153]_ , \new_[29154]_ , \new_[29155]_ , \new_[29156]_ ,
    \new_[29157]_ , \new_[29158]_ , \new_[29159]_ , \new_[29160]_ ,
    \new_[29161]_ , \new_[29162]_ , \new_[29163]_ , \new_[29164]_ ,
    \new_[29165]_ , \new_[29166]_ , \new_[29167]_ , \new_[29168]_ ,
    \new_[29169]_ , \new_[29170]_ , \new_[29171]_ , \new_[29172]_ ,
    \new_[29173]_ , \new_[29174]_ , \new_[29175]_ , \new_[29176]_ ,
    \new_[29177]_ , \new_[29178]_ , \new_[29179]_ , \new_[29180]_ ,
    \new_[29181]_ , \new_[29182]_ , \new_[29183]_ , \new_[29184]_ ,
    \new_[29185]_ , \new_[29186]_ , \new_[29187]_ , \new_[29188]_ ,
    \new_[29189]_ , \new_[29190]_ , \new_[29191]_ , \new_[29192]_ ,
    \new_[29193]_ , \new_[29194]_ , \new_[29195]_ , \new_[29196]_ ,
    \new_[29197]_ , \new_[29198]_ , \new_[29199]_ , \new_[29200]_ ,
    \new_[29201]_ , \new_[29202]_ , \new_[29203]_ , \new_[29204]_ ,
    \new_[29205]_ , \new_[29206]_ , \new_[29207]_ , \new_[29208]_ ,
    \new_[29209]_ , \new_[29210]_ , \new_[29211]_ , \new_[29212]_ ,
    \new_[29213]_ , \new_[29214]_ , \new_[29215]_ , \new_[29216]_ ,
    \new_[29217]_ , \new_[29218]_ , \new_[29219]_ , \new_[29220]_ ,
    \new_[29221]_ , \new_[29222]_ , \new_[29223]_ , \new_[29224]_ ,
    \new_[29225]_ , \new_[29226]_ , \new_[29227]_ , \new_[29228]_ ,
    \new_[29229]_ , \new_[29230]_ , \new_[29231]_ , \new_[29232]_ ,
    \new_[29233]_ , \new_[29234]_ , \new_[29235]_ , \new_[29236]_ ,
    \new_[29237]_ , \new_[29238]_ , \new_[29239]_ , \new_[29240]_ ,
    \new_[29241]_ , \new_[29242]_ , \new_[29243]_ , \new_[29244]_ ,
    \new_[29245]_ , \new_[29246]_ , \new_[29247]_ , \new_[29248]_ ,
    \new_[29249]_ , \new_[29250]_ , \new_[29251]_ , \new_[29252]_ ,
    \new_[29253]_ , \new_[29254]_ , \new_[29255]_ , \new_[29256]_ ,
    \new_[29257]_ , \new_[29258]_ , \new_[29259]_ , \new_[29260]_ ,
    \new_[29261]_ , \new_[29262]_ , \new_[29263]_ , \new_[29264]_ ,
    \new_[29265]_ , \new_[29266]_ , \new_[29267]_ , \new_[29268]_ ,
    \new_[29269]_ , \new_[29270]_ , \new_[29271]_ , \new_[29272]_ ,
    \new_[29273]_ , \new_[29274]_ , \new_[29275]_ , \new_[29276]_ ,
    \new_[29277]_ , \new_[29278]_ , \new_[29279]_ , \new_[29280]_ ,
    \new_[29281]_ , \new_[29282]_ , \new_[29283]_ , \new_[29284]_ ,
    \new_[29285]_ , \new_[29286]_ , \new_[29287]_ , \new_[29288]_ ,
    \new_[29289]_ , \new_[29290]_ , \new_[29291]_ , \new_[29292]_ ,
    \new_[29293]_ , \new_[29294]_ , \new_[29295]_ , \new_[29296]_ ,
    \new_[29297]_ , \new_[29298]_ , \new_[29299]_ , \new_[29300]_ ,
    \new_[29301]_ , \new_[29302]_ , \new_[29303]_ , \new_[29304]_ ,
    \new_[29305]_ , \new_[29306]_ , \new_[29307]_ , \new_[29308]_ ,
    \new_[29309]_ , \new_[29310]_ , \new_[29311]_ , \new_[29312]_ ,
    \new_[29313]_ , \new_[29314]_ , \new_[29315]_ , \new_[29316]_ ,
    \new_[29317]_ , \new_[29318]_ , \new_[29319]_ , \new_[29320]_ ,
    \new_[29321]_ , \new_[29322]_ , \new_[29323]_ , \new_[29324]_ ,
    \new_[29325]_ , \new_[29326]_ , \new_[29327]_ , \new_[29328]_ ,
    \new_[29329]_ , \new_[29330]_ , \new_[29331]_ , \new_[29332]_ ,
    \new_[29333]_ , \new_[29334]_ , \new_[29335]_ , \new_[29336]_ ,
    \new_[29337]_ , \new_[29338]_ , \new_[29339]_ , \new_[29340]_ ,
    \new_[29341]_ , \new_[29342]_ , \new_[29343]_ , \new_[29344]_ ,
    \new_[29345]_ , \new_[29346]_ , \new_[29347]_ , \new_[29348]_ ,
    \new_[29349]_ , \new_[29350]_ , \new_[29351]_ , \new_[29352]_ ,
    \new_[29353]_ , \new_[29354]_ , \new_[29355]_ , \new_[29356]_ ,
    \new_[29357]_ , \new_[29358]_ , \new_[29359]_ , \new_[29360]_ ,
    \new_[29361]_ , \new_[29362]_ , \new_[29363]_ , \new_[29364]_ ,
    \new_[29365]_ , \new_[29366]_ , \new_[29367]_ , \new_[29368]_ ,
    \new_[29369]_ , \new_[29370]_ , \new_[29371]_ , \new_[29372]_ ,
    \new_[29373]_ , \new_[29374]_ , \new_[29375]_ , \new_[29376]_ ,
    \new_[29377]_ , \new_[29378]_ , \new_[29379]_ , \new_[29380]_ ,
    \new_[29381]_ , \new_[29382]_ , \new_[29383]_ , \new_[29384]_ ,
    \new_[29385]_ , \new_[29386]_ , \new_[29387]_ , \new_[29388]_ ,
    \new_[29389]_ , \new_[29390]_ , \new_[29391]_ , \new_[29392]_ ,
    \new_[29393]_ , \new_[29394]_ , \new_[29395]_ , \new_[29396]_ ,
    \new_[29397]_ , \new_[29398]_ , \new_[29399]_ , \new_[29400]_ ,
    \new_[29401]_ , \new_[29402]_ , \new_[29403]_ , \new_[29404]_ ,
    \new_[29405]_ , \new_[29406]_ , \new_[29407]_ , \new_[29408]_ ,
    \new_[29409]_ , \new_[29410]_ , \new_[29411]_ , \new_[29412]_ ,
    \new_[29413]_ , \new_[29414]_ , \new_[29415]_ , \new_[29416]_ ,
    \new_[29417]_ , \new_[29418]_ , \new_[29419]_ , \new_[29420]_ ,
    \new_[29421]_ , \new_[29422]_ , \new_[29423]_ , \new_[29424]_ ,
    \new_[29425]_ , \new_[29426]_ , \new_[29427]_ , \new_[29428]_ ,
    \new_[29429]_ , \new_[29430]_ , \new_[29431]_ , \new_[29432]_ ,
    \new_[29433]_ , \new_[29434]_ , \new_[29435]_ , \new_[29436]_ ,
    \new_[29437]_ , \new_[29438]_ , \new_[29439]_ , \new_[29440]_ ,
    \new_[29441]_ , \new_[29442]_ , \new_[29443]_ , \new_[29444]_ ,
    \new_[29445]_ , \new_[29446]_ , \new_[29447]_ , \new_[29448]_ ,
    \new_[29449]_ , \new_[29450]_ , \new_[29451]_ , \new_[29452]_ ,
    \new_[29453]_ , \new_[29454]_ , \new_[29455]_ , \new_[29456]_ ,
    \new_[29457]_ , \new_[29458]_ , \new_[29459]_ , \new_[29460]_ ,
    \new_[29461]_ , \new_[29462]_ , \new_[29463]_ , \new_[29464]_ ,
    \new_[29465]_ , \new_[29466]_ , \new_[29467]_ , \new_[29468]_ ,
    \new_[29469]_ , \new_[29470]_ , \new_[29471]_ , \new_[29472]_ ,
    \new_[29473]_ , \new_[29474]_ , \new_[29475]_ , \new_[29476]_ ,
    \new_[29477]_ , \new_[29478]_ , \new_[29479]_ , \new_[29480]_ ,
    \new_[29481]_ , \new_[29482]_ , \new_[29483]_ , \new_[29484]_ ,
    \new_[29485]_ , \new_[29486]_ , \new_[29487]_ , \new_[29488]_ ,
    \new_[29489]_ , \new_[29490]_ , \new_[29491]_ , \new_[29492]_ ,
    \new_[29493]_ , \new_[29494]_ , \new_[29495]_ , \new_[29496]_ ,
    \new_[29497]_ , \new_[29498]_ , \new_[29499]_ , \new_[29500]_ ,
    \new_[29501]_ , \new_[29502]_ , \new_[29503]_ , \new_[29504]_ ,
    \new_[29505]_ , \new_[29506]_ , \new_[29507]_ , \new_[29508]_ ,
    \new_[29509]_ , \new_[29510]_ , \new_[29511]_ , \new_[29512]_ ,
    \new_[29513]_ , \new_[29514]_ , \new_[29515]_ , \new_[29516]_ ,
    \new_[29517]_ , \new_[29518]_ , \new_[29519]_ , \new_[29520]_ ,
    \new_[29521]_ , \new_[29522]_ , \new_[29523]_ , \new_[29524]_ ,
    \new_[29525]_ , \new_[29526]_ , \new_[29527]_ , \new_[29528]_ ,
    \new_[29529]_ , \new_[29530]_ , \new_[29531]_ , \new_[29532]_ ,
    \new_[29533]_ , \new_[29534]_ , \new_[29535]_ , \new_[29536]_ ,
    \new_[29537]_ , \new_[29538]_ , \new_[29539]_ , \new_[29540]_ ,
    \new_[29541]_ , \new_[29542]_ , \new_[29543]_ , \new_[29544]_ ,
    \new_[29545]_ , \new_[29546]_ , \new_[29547]_ , \new_[29548]_ ,
    \new_[29549]_ , \new_[29550]_ , \new_[29551]_ , \new_[29552]_ ,
    \new_[29553]_ , \new_[29554]_ , \new_[29555]_ , \new_[29556]_ ,
    \new_[29557]_ , \new_[29558]_ , \new_[29559]_ , \new_[29560]_ ,
    \new_[29561]_ , \new_[29562]_ , \new_[29563]_ , \new_[29564]_ ,
    \new_[29565]_ , \new_[29566]_ , \new_[29567]_ , \new_[29568]_ ,
    \new_[29569]_ , \new_[29570]_ , \new_[29571]_ , \new_[29572]_ ,
    \new_[29573]_ , \new_[29574]_ , \new_[29575]_ , \new_[29576]_ ,
    \new_[29577]_ , \new_[29578]_ , \new_[29579]_ , \new_[29580]_ ,
    \new_[29581]_ , \new_[29582]_ , \new_[29583]_ , \new_[29584]_ ,
    \new_[29585]_ , \new_[29586]_ , \new_[29587]_ , \new_[29588]_ ,
    \new_[29589]_ , \new_[29590]_ , \new_[29591]_ , \new_[29592]_ ,
    \new_[29593]_ , \new_[29594]_ , \new_[29595]_ , \new_[29596]_ ,
    \new_[29597]_ , \new_[29598]_ , \new_[29599]_ , \new_[29600]_ ,
    \new_[29601]_ , \new_[29602]_ , \new_[29603]_ , \new_[29604]_ ,
    \new_[29605]_ , \new_[29606]_ , \new_[29607]_ , \new_[29608]_ ,
    \new_[29609]_ , \new_[29610]_ , \new_[29611]_ , \new_[29612]_ ,
    \new_[29613]_ , \new_[29614]_ , \new_[29615]_ , \new_[29616]_ ,
    \new_[29617]_ , \new_[29618]_ , \new_[29619]_ , \new_[29620]_ ,
    \new_[29621]_ , \new_[29622]_ , \new_[29623]_ , \new_[29624]_ ,
    \new_[29625]_ , \new_[29626]_ , \new_[29627]_ , \new_[29628]_ ,
    \new_[29629]_ , \new_[29630]_ , \new_[29631]_ , \new_[29632]_ ,
    \new_[29633]_ , \new_[29634]_ , \new_[29635]_ , \new_[29636]_ ,
    \new_[29637]_ , \new_[29638]_ , \new_[29639]_ , \new_[29640]_ ,
    \new_[29641]_ , \new_[29642]_ , \new_[29643]_ , \new_[29644]_ ,
    \new_[29645]_ , \new_[29646]_ , \new_[29647]_ , \new_[29648]_ ,
    \new_[29649]_ , \new_[29650]_ , \new_[29651]_ , \new_[29652]_ ,
    \new_[29653]_ , \new_[29654]_ , \new_[29655]_ , \new_[29656]_ ,
    \new_[29657]_ , \new_[29658]_ , \new_[29659]_ , \new_[29660]_ ,
    \new_[29661]_ , \new_[29662]_ , \new_[29663]_ , \new_[29664]_ ,
    \new_[29665]_ , \new_[29666]_ , \new_[29667]_ , \new_[29668]_ ,
    \new_[29669]_ , \new_[29670]_ , \new_[29671]_ , \new_[29672]_ ,
    \new_[29673]_ , \new_[29674]_ , \new_[29675]_ , \new_[29676]_ ,
    \new_[29677]_ , \new_[29678]_ , \new_[29679]_ , \new_[29680]_ ,
    \new_[29681]_ , \new_[29682]_ , \new_[29683]_ , \new_[29684]_ ,
    \new_[29685]_ , \new_[29686]_ , \new_[29687]_ , \new_[29688]_ ,
    \new_[29689]_ , \new_[29690]_ , \new_[29691]_ , \new_[29692]_ ,
    \new_[29693]_ , \new_[29694]_ , \new_[29695]_ , \new_[29696]_ ,
    \new_[29697]_ , \new_[29698]_ , \new_[29699]_ , \new_[29700]_ ,
    \new_[29701]_ , \new_[29702]_ , \new_[29703]_ , \new_[29704]_ ,
    \new_[29705]_ , \new_[29706]_ , \new_[29707]_ , \new_[29708]_ ,
    \new_[29709]_ , \new_[29710]_ , \new_[29711]_ , \new_[29712]_ ,
    \new_[29713]_ , \new_[29714]_ , \new_[29715]_ , \new_[29716]_ ,
    \new_[29717]_ , \new_[29718]_ , \new_[29719]_ , \new_[29720]_ ,
    \new_[29721]_ , \new_[29722]_ , \new_[29723]_ , \new_[29724]_ ,
    \new_[29725]_ , \new_[29726]_ , \new_[29727]_ , \new_[29728]_ ,
    \new_[29729]_ , \new_[29730]_ , \new_[29731]_ , \new_[29732]_ ,
    \new_[29733]_ , \new_[29734]_ , \new_[29735]_ , \new_[29736]_ ,
    \new_[29737]_ , \new_[29738]_ , \new_[29739]_ , \new_[29740]_ ,
    \new_[29741]_ , \new_[29742]_ , \new_[29743]_ , \new_[29744]_ ,
    \new_[29745]_ , \new_[29746]_ , \new_[29747]_ , \new_[29748]_ ,
    \new_[29749]_ , \new_[29750]_ , \new_[29751]_ , \new_[29752]_ ,
    \new_[29753]_ , \new_[29754]_ , \new_[29755]_ , \new_[29756]_ ,
    \new_[29757]_ , \new_[29758]_ , \new_[29759]_ , \new_[29760]_ ,
    \new_[29761]_ , \new_[29762]_ , \new_[29763]_ , \new_[29764]_ ,
    \new_[29765]_ , \new_[29766]_ , \new_[29767]_ , \new_[29768]_ ,
    \new_[29769]_ , \new_[29770]_ , \new_[29771]_ , \new_[29772]_ ,
    \new_[29773]_ , \new_[29774]_ , \new_[29775]_ , \new_[29776]_ ,
    \new_[29777]_ , \new_[29778]_ , \new_[29779]_ , \new_[29780]_ ,
    \new_[29781]_ , \new_[29782]_ , \new_[29783]_ , \new_[29784]_ ,
    \new_[29785]_ , \new_[29786]_ , \new_[29787]_ , \new_[29788]_ ,
    \new_[29789]_ , \new_[29790]_ , \new_[29791]_ , \new_[29792]_ ,
    \new_[29793]_ , \new_[29794]_ , \new_[29795]_ , \new_[29796]_ ,
    \new_[29797]_ , \new_[29798]_ , \new_[29799]_ , \new_[29800]_ ,
    \new_[29801]_ , \new_[29802]_ , \new_[29803]_ , \new_[29804]_ ,
    \new_[29805]_ , \new_[29806]_ , \new_[29807]_ , \new_[29808]_ ,
    \new_[29809]_ , \new_[29810]_ , \new_[29811]_ , \new_[29812]_ ,
    \new_[29813]_ , \new_[29814]_ , \new_[29815]_ , \new_[29816]_ ,
    \new_[29817]_ , \new_[29818]_ , \new_[29819]_ , \new_[29820]_ ,
    \new_[29821]_ , \new_[29822]_ , \new_[29823]_ , \new_[29824]_ ,
    \new_[29825]_ , \new_[29826]_ , \new_[29827]_ , \new_[29828]_ ,
    \new_[29829]_ , \new_[29830]_ , \new_[29831]_ , \new_[29832]_ ,
    \new_[29833]_ , \new_[29834]_ , \new_[29835]_ , \new_[29836]_ ,
    \new_[29837]_ , \new_[29838]_ , \new_[29839]_ , \new_[29840]_ ,
    \new_[29841]_ , \new_[29842]_ , \new_[29843]_ , \new_[29844]_ ,
    \new_[29845]_ , \new_[29846]_ , \new_[29847]_ , \new_[29848]_ ,
    \new_[29849]_ , \new_[29850]_ , \new_[29851]_ , \new_[29852]_ ,
    \new_[29853]_ , \new_[29854]_ , \new_[29855]_ , \new_[29856]_ ,
    \new_[29857]_ , \new_[29858]_ , \new_[29859]_ , \new_[29860]_ ,
    \new_[29861]_ , \new_[29862]_ , \new_[29863]_ , \new_[29864]_ ,
    \new_[29865]_ , \new_[29866]_ , \new_[29867]_ , \new_[29868]_ ,
    \new_[29869]_ , \new_[29870]_ , \new_[29871]_ , \new_[29872]_ ,
    \new_[29873]_ , \new_[29874]_ , \new_[29875]_ , \new_[29876]_ ,
    \new_[29877]_ , \new_[29878]_ , \new_[29879]_ , \new_[29880]_ ,
    \new_[29881]_ , \new_[29882]_ , \new_[29883]_ , \new_[29884]_ ,
    \new_[29885]_ , \new_[29886]_ , \new_[29887]_ , \new_[29888]_ ,
    \new_[29889]_ , \new_[29890]_ , \new_[29891]_ , \new_[29892]_ ,
    \new_[29893]_ , \new_[29894]_ , \new_[29895]_ , \new_[29896]_ ,
    \new_[29897]_ , \new_[29898]_ , \new_[29899]_ , \new_[29900]_ ,
    \new_[29901]_ , \new_[29902]_ , \new_[29903]_ , \new_[29904]_ ,
    \new_[29905]_ , \new_[29906]_ , \new_[29907]_ , \new_[29908]_ ,
    \new_[29909]_ , \new_[29910]_ , \new_[29911]_ , \new_[29912]_ ,
    \new_[29913]_ , \new_[29914]_ , \new_[29915]_ , \new_[29916]_ ,
    \new_[29917]_ , \new_[29918]_ , \new_[29919]_ , \new_[29920]_ ,
    \new_[29921]_ , \new_[29922]_ , \new_[29923]_ , \new_[29924]_ ,
    \new_[29925]_ , \new_[29926]_ , \new_[29927]_ , \new_[29928]_ ,
    \new_[29929]_ , \new_[29930]_ , \new_[29931]_ , \new_[29932]_ ,
    \new_[29933]_ , \new_[29934]_ , \new_[29935]_ , \new_[29936]_ ,
    \new_[29937]_ , \new_[29938]_ , \new_[29939]_ , \new_[29940]_ ,
    \new_[29941]_ , \new_[29942]_ , \new_[29943]_ , \new_[29944]_ ,
    \new_[29945]_ , \new_[29946]_ , \new_[29947]_ , \new_[29948]_ ,
    \new_[29949]_ , \new_[29950]_ , \new_[29951]_ , \new_[29952]_ ,
    \new_[29953]_ , \new_[29954]_ , \new_[29955]_ , \new_[29956]_ ,
    \new_[29957]_ , \new_[29958]_ , \new_[29959]_ , \new_[29960]_ ,
    \new_[29961]_ , \new_[29962]_ , \new_[29963]_ , \new_[29964]_ ,
    \new_[29965]_ , \new_[29966]_ , \new_[29967]_ , \new_[29968]_ ,
    \new_[29969]_ , \new_[29970]_ , \new_[29971]_ , \new_[29972]_ ,
    \new_[29973]_ , \new_[29974]_ , \new_[29975]_ , \new_[29976]_ ,
    \new_[29977]_ , \new_[29978]_ , \new_[29979]_ , \new_[29980]_ ,
    \new_[29981]_ , \new_[29982]_ , \new_[29983]_ , \new_[29984]_ ,
    \new_[29985]_ , \new_[29986]_ , \new_[29987]_ , \new_[29988]_ ,
    \new_[29989]_ , \new_[29990]_ , \new_[29991]_ , \new_[29992]_ ,
    \new_[29993]_ , \new_[29994]_ , \new_[29995]_ , \new_[29996]_ ,
    \new_[29997]_ , \new_[29998]_ , \new_[29999]_ , \new_[30000]_ ,
    \new_[30001]_ , \new_[30002]_ , \new_[30003]_ , \new_[30004]_ ,
    \new_[30005]_ , \new_[30006]_ , \new_[30007]_ , \new_[30008]_ ,
    \new_[30009]_ , \new_[30010]_ , \new_[30011]_ , \new_[30012]_ ,
    \new_[30013]_ , \new_[30014]_ , \new_[30015]_ , \new_[30016]_ ,
    \new_[30017]_ , \new_[30018]_ , \new_[30019]_ , \new_[30020]_ ,
    \new_[30021]_ , \new_[30022]_ , \new_[30023]_ , \new_[30024]_ ,
    \new_[30025]_ , \new_[30026]_ , \new_[30027]_ , \new_[30028]_ ,
    \new_[30029]_ , \new_[30030]_ , \new_[30031]_ , \new_[30032]_ ,
    \new_[30033]_ , \new_[30034]_ , \new_[30035]_ , \new_[30036]_ ,
    \new_[30037]_ , \new_[30038]_ , \new_[30039]_ , \new_[30040]_ ,
    \new_[30041]_ , \new_[30042]_ , \new_[30043]_ , \new_[30044]_ ,
    \new_[30045]_ , \new_[30046]_ , \new_[30047]_ , \new_[30048]_ ,
    \new_[30049]_ , \new_[30050]_ , \new_[30051]_ , \new_[30052]_ ,
    \new_[30053]_ , \new_[30054]_ , \new_[30055]_ , \new_[30056]_ ,
    \new_[30057]_ , \new_[30058]_ , \new_[30059]_ , \new_[30060]_ ,
    \new_[30061]_ , \new_[30062]_ , \new_[30063]_ , \new_[30064]_ ,
    \new_[30065]_ , \new_[30066]_ , \new_[30067]_ , \new_[30068]_ ,
    \new_[30069]_ , \new_[30070]_ , \new_[30071]_ , \new_[30072]_ ,
    \new_[30073]_ , \new_[30074]_ , \new_[30075]_ , \new_[30076]_ ,
    \new_[30077]_ , \new_[30078]_ , \new_[30079]_ , \new_[30080]_ ,
    \new_[30081]_ , \new_[30082]_ , \new_[30083]_ , \new_[30084]_ ,
    \new_[30085]_ , \new_[30086]_ , \new_[30087]_ , \new_[30088]_ ,
    \new_[30089]_ , \new_[30090]_ , \new_[30091]_ , \new_[30092]_ ,
    \new_[30093]_ , \new_[30094]_ , \new_[30095]_ , \new_[30096]_ ,
    \new_[30097]_ , \new_[30098]_ , \new_[30099]_ , \new_[30100]_ ,
    \new_[30101]_ , \new_[30102]_ , \new_[30103]_ , \new_[30104]_ ,
    \new_[30105]_ , \new_[30106]_ , \new_[30107]_ , \new_[30108]_ ,
    \new_[30109]_ , \new_[30110]_ , \new_[30111]_ , \new_[30112]_ ,
    \new_[30113]_ , \new_[30114]_ , \new_[30115]_ , \new_[30116]_ ,
    \new_[30117]_ , \new_[30118]_ , \new_[30119]_ , \new_[30120]_ ,
    \new_[30121]_ , \new_[30122]_ , \new_[30123]_ , \new_[30124]_ ,
    \new_[30125]_ , \new_[30126]_ , \new_[30127]_ , \new_[30128]_ ,
    \new_[30129]_ , \new_[30130]_ , \new_[30131]_ , \new_[30132]_ ,
    \new_[30133]_ , \new_[30134]_ , \new_[30135]_ , \new_[30136]_ ,
    \new_[30137]_ , \new_[30138]_ , \new_[30139]_ , \new_[30140]_ ,
    \new_[30141]_ , \new_[30142]_ , \new_[30143]_ , \new_[30144]_ ,
    \new_[30145]_ , \new_[30146]_ , \new_[30147]_ , \new_[30148]_ ,
    \new_[30149]_ , \new_[30150]_ , \new_[30151]_ , \new_[30152]_ ,
    \new_[30153]_ , \new_[30154]_ , \new_[30155]_ , \new_[30156]_ ,
    \new_[30157]_ , \new_[30158]_ , \new_[30159]_ , \new_[30160]_ ,
    \new_[30161]_ , \new_[30162]_ , \new_[30163]_ , \new_[30164]_ ,
    \new_[30165]_ , \new_[30166]_ , \new_[30167]_ , \new_[30168]_ ,
    \new_[30169]_ , \new_[30170]_ , \new_[30171]_ , \new_[30172]_ ,
    \new_[30173]_ , \new_[30174]_ , \new_[30175]_ , \new_[30176]_ ,
    \new_[30177]_ , \new_[30178]_ , \new_[30179]_ , \new_[30180]_ ,
    \new_[30181]_ , \new_[30182]_ , \new_[30183]_ , \new_[30184]_ ,
    \new_[30185]_ , \new_[30186]_ , \new_[30187]_ , \new_[30188]_ ,
    \new_[30189]_ , \new_[30190]_ , \new_[30191]_ , \new_[30192]_ ,
    \new_[30193]_ , \new_[30194]_ , \new_[30195]_ , \new_[30196]_ ,
    \new_[30197]_ , \new_[30198]_ , \new_[30199]_ , \new_[30200]_ ,
    \new_[30201]_ , \new_[30202]_ , \new_[30203]_ , \new_[30204]_ ,
    \new_[30205]_ , \new_[30206]_ , \new_[30207]_ , \new_[30208]_ ,
    \new_[30209]_ , \new_[30210]_ , \new_[30211]_ , \new_[30212]_ ,
    \new_[30213]_ , \new_[30214]_ , \new_[30215]_ , \new_[30216]_ ,
    \new_[30217]_ , \new_[30218]_ , \new_[30219]_ , \new_[30220]_ ,
    \new_[30221]_ , \new_[30222]_ , \new_[30223]_ , \new_[30224]_ ,
    \new_[30225]_ , \new_[30226]_ , \new_[30227]_ , \new_[30228]_ ,
    \new_[30229]_ , \new_[30230]_ , \new_[30231]_ , \new_[30232]_ ,
    \new_[30233]_ , \new_[30234]_ , \new_[30235]_ , \new_[30236]_ ,
    \new_[30237]_ , \new_[30238]_ , \new_[30239]_ , \new_[30240]_ ,
    \new_[30241]_ , \new_[30242]_ , \new_[30243]_ , \new_[30244]_ ,
    \new_[30245]_ , \new_[30246]_ , \new_[30247]_ , \new_[30248]_ ,
    \new_[30249]_ , \new_[30250]_ , \new_[30251]_ , \new_[30252]_ ,
    \new_[30253]_ , \new_[30254]_ , \new_[30255]_ , \new_[30256]_ ,
    \new_[30257]_ , \new_[30258]_ , \new_[30259]_ , \new_[30260]_ ,
    \new_[30261]_ , \new_[30262]_ , \new_[30263]_ , \new_[30264]_ ,
    \new_[30265]_ , \new_[30266]_ , \new_[30267]_ , \new_[30268]_ ,
    \new_[30269]_ , \new_[30270]_ , \new_[30271]_ , \new_[30272]_ ,
    \new_[30273]_ , \new_[30274]_ , \new_[30275]_ , \new_[30276]_ ,
    \new_[30277]_ , \new_[30278]_ , \new_[30279]_ , \new_[30280]_ ,
    \new_[30281]_ , \new_[30282]_ , \new_[30283]_ , \new_[30284]_ ,
    \new_[30285]_ , \new_[30286]_ , \new_[30287]_ , \new_[30288]_ ,
    \new_[30289]_ , \new_[30290]_ , \new_[30291]_ , \new_[30292]_ ,
    \new_[30293]_ , \new_[30294]_ , \new_[30295]_ , \new_[30296]_ ,
    \new_[30297]_ , \new_[30298]_ , \new_[30299]_ , \new_[30300]_ ,
    \new_[30301]_ , \new_[30302]_ , \new_[30303]_ , \new_[30304]_ ,
    \new_[30305]_ , \new_[30306]_ , \new_[30307]_ , \new_[30308]_ ,
    \new_[30309]_ , \new_[30310]_ , \new_[30311]_ , \new_[30312]_ ,
    \new_[30313]_ , \new_[30314]_ , \new_[30315]_ , \new_[30316]_ ,
    \new_[30317]_ , \new_[30318]_ , \new_[30319]_ , \new_[30320]_ ,
    \new_[30321]_ , \new_[30322]_ , \new_[30323]_ , \new_[30324]_ ,
    \new_[30325]_ , \new_[30326]_ , \new_[30327]_ , \new_[30328]_ ,
    \new_[30329]_ , \new_[30330]_ , \new_[30331]_ , \new_[30332]_ ,
    \new_[30333]_ , \new_[30334]_ , \new_[30335]_ , \new_[30336]_ ,
    \new_[30337]_ , \new_[30338]_ , \new_[30339]_ , \new_[30340]_ ,
    \new_[30341]_ , \new_[30342]_ , \new_[30343]_ , \new_[30344]_ ,
    \new_[30345]_ , \new_[30346]_ , \new_[30347]_ , \new_[30348]_ ,
    \new_[30349]_ , \new_[30350]_ , \new_[30351]_ , \new_[30352]_ ,
    \new_[30353]_ , \new_[30354]_ , \new_[30355]_ , \new_[30356]_ ,
    \new_[30357]_ , \new_[30358]_ , \new_[30359]_ , \new_[30360]_ ,
    \new_[30361]_ , \new_[30362]_ , \new_[30363]_ , \new_[30364]_ ,
    \new_[30365]_ , \new_[30366]_ , \new_[30367]_ , \new_[30368]_ ,
    \new_[30369]_ , \new_[30370]_ , \new_[30371]_ , \new_[30372]_ ,
    \new_[30373]_ , \new_[30374]_ , \new_[30375]_ , \new_[30376]_ ,
    \new_[30377]_ , \new_[30378]_ , \new_[30379]_ , \new_[30380]_ ,
    \new_[30381]_ , \new_[30382]_ , \new_[30383]_ , \new_[30384]_ ,
    \new_[30385]_ , \new_[30386]_ , \new_[30387]_ , \new_[30388]_ ,
    \new_[30389]_ , \new_[30390]_ , \new_[30391]_ , \new_[30392]_ ,
    \new_[30393]_ , \new_[30394]_ , \new_[30395]_ , \new_[30396]_ ,
    \new_[30397]_ , \new_[30398]_ , \new_[30399]_ , \new_[30400]_ ,
    \new_[30401]_ , \new_[30402]_ , \new_[30403]_ , \new_[30404]_ ,
    \new_[30405]_ , \new_[30406]_ , \new_[30407]_ , \new_[30408]_ ,
    \new_[30409]_ , \new_[30410]_ , \new_[30411]_ , \new_[30412]_ ,
    \new_[30413]_ , \new_[30414]_ , \new_[30415]_ , \new_[30416]_ ,
    \new_[30417]_ , \new_[30418]_ , \new_[30419]_ , \new_[30420]_ ,
    \new_[30421]_ , \new_[30422]_ , \new_[30423]_ , \new_[30424]_ ,
    \new_[30425]_ , \new_[30426]_ , \new_[30427]_ , \new_[30428]_ ,
    \new_[30429]_ , \new_[30430]_ , \new_[30431]_ , \new_[30432]_ ,
    \new_[30433]_ , \new_[30434]_ , \new_[30435]_ , \new_[30436]_ ,
    \new_[30437]_ , \new_[30438]_ , \new_[30439]_ , \new_[30440]_ ,
    \new_[30441]_ , \new_[30442]_ , \new_[30443]_ , \new_[30444]_ ,
    \new_[30445]_ , \new_[30446]_ , \new_[30447]_ , \new_[30448]_ ,
    \new_[30449]_ , \new_[30450]_ , \new_[30451]_ , \new_[30452]_ ,
    \new_[30453]_ , \new_[30454]_ , \new_[30455]_ , \new_[30456]_ ,
    \new_[30457]_ , \new_[30458]_ , \new_[30459]_ , \new_[30460]_ ,
    \new_[30461]_ , \new_[30462]_ , \new_[30463]_ , \new_[30464]_ ,
    \new_[30465]_ , \new_[30466]_ , \new_[30467]_ , \new_[30468]_ ,
    \new_[30469]_ , \new_[30470]_ , \new_[30471]_ , \new_[30472]_ ,
    \new_[30473]_ , \new_[30474]_ , \new_[30475]_ , \new_[30476]_ ,
    \new_[30477]_ , \new_[30478]_ , \new_[30479]_ , \new_[30480]_ ,
    \new_[30481]_ , \new_[30482]_ , \new_[30483]_ , \new_[30484]_ ,
    \new_[30485]_ , \new_[30486]_ , \new_[30487]_ , \new_[30488]_ ,
    \new_[30489]_ , \new_[30490]_ , \new_[30491]_ , \new_[30492]_ ,
    \new_[30493]_ , \new_[30494]_ , \new_[30495]_ , \new_[30496]_ ,
    \new_[30497]_ , \new_[30498]_ , \new_[30499]_ , \new_[30500]_ ,
    \new_[30501]_ , \new_[30502]_ , \new_[30503]_ , \new_[30504]_ ,
    \new_[30505]_ , \new_[30506]_ , \new_[30507]_ , \new_[30508]_ ,
    \new_[30509]_ , \new_[30510]_ , \new_[30511]_ , \new_[30512]_ ,
    \new_[30513]_ , \new_[30514]_ , \new_[30515]_ , \new_[30516]_ ,
    \new_[30517]_ , \new_[30518]_ , \new_[30519]_ , \new_[30520]_ ,
    \new_[30521]_ , \new_[30522]_ , \new_[30523]_ , \new_[30524]_ ,
    \new_[30525]_ , \new_[30526]_ , \new_[30527]_ , \new_[30528]_ ,
    \new_[30529]_ , \new_[30530]_ , \new_[30531]_ , \new_[30532]_ ,
    \new_[30533]_ , \new_[30534]_ , \new_[30535]_ , \new_[30536]_ ,
    \new_[30537]_ , \new_[30538]_ , \new_[30539]_ , \new_[30540]_ ,
    \new_[30541]_ , \new_[30542]_ , \new_[30543]_ , \new_[30544]_ ,
    \new_[30545]_ , \new_[30546]_ , \new_[30547]_ , \new_[30548]_ ,
    \new_[30549]_ , \new_[30550]_ , \new_[30551]_ , \new_[30552]_ ,
    \new_[30553]_ , \new_[30554]_ , \new_[30555]_ , \new_[30556]_ ,
    \new_[30557]_ , \new_[30558]_ , \new_[30559]_ , \new_[30560]_ ,
    \new_[30561]_ , \new_[30562]_ , \new_[30563]_ , \new_[30564]_ ,
    \new_[30565]_ , \new_[30566]_ , \new_[30567]_ , \new_[30568]_ ,
    \new_[30569]_ , \new_[30570]_ , \new_[30571]_ , \new_[30572]_ ,
    \new_[30573]_ , \new_[30574]_ , \new_[30575]_ , \new_[30576]_ ,
    \new_[30577]_ , \new_[30578]_ , \new_[30579]_ , \new_[30580]_ ,
    \new_[30581]_ , \new_[30582]_ , \new_[30583]_ , \new_[30584]_ ,
    \new_[30585]_ , \new_[30586]_ , \new_[30587]_ , \new_[30588]_ ,
    \new_[30589]_ , \new_[30590]_ , \new_[30591]_ , \new_[30592]_ ,
    \new_[30593]_ , \new_[30594]_ , \new_[30595]_ , \new_[30596]_ ,
    \new_[30597]_ , \new_[30598]_ , \new_[30599]_ , \new_[30600]_ ,
    \new_[30601]_ , \new_[30602]_ , \new_[30603]_ , \new_[30604]_ ,
    \new_[30605]_ , \new_[30606]_ , \new_[30607]_ , \new_[30608]_ ,
    \new_[30609]_ , \new_[30610]_ , \new_[30611]_ , \new_[30612]_ ,
    \new_[30613]_ , \new_[30614]_ , \new_[30615]_ , \new_[30616]_ ,
    \new_[30617]_ , \new_[30618]_ , \new_[30619]_ , \new_[30620]_ ,
    \new_[30621]_ , \new_[30622]_ , \new_[30623]_ , \new_[30624]_ ,
    \new_[30625]_ , \new_[30626]_ , \new_[30627]_ , \new_[30628]_ ,
    \new_[30629]_ , \new_[30630]_ , \new_[30631]_ , \new_[30632]_ ,
    \new_[30633]_ , \new_[30634]_ , \new_[30635]_ , \new_[30636]_ ,
    \new_[30637]_ , \new_[30638]_ , \new_[30639]_ , \new_[30640]_ ,
    \new_[30641]_ , \new_[30642]_ , \new_[30643]_ , \new_[30644]_ ,
    \new_[30645]_ , \new_[30646]_ , \new_[30647]_ , \new_[30648]_ ,
    \new_[30649]_ , \new_[30650]_ , \new_[30651]_ , \new_[30652]_ ,
    \new_[30653]_ , \new_[30654]_ , \new_[30655]_ , \new_[30656]_ ,
    \new_[30657]_ , \new_[30658]_ , \new_[30659]_ , \new_[30660]_ ,
    \new_[30661]_ , \new_[30662]_ , \new_[30663]_ , \new_[30664]_ ,
    \new_[30665]_ , \new_[30666]_ , \new_[30667]_ , \new_[30668]_ ,
    \new_[30669]_ , \new_[30670]_ , \new_[30671]_ , \new_[30672]_ ,
    \new_[30673]_ , \new_[30674]_ , \new_[30675]_ , \new_[30676]_ ,
    \new_[30677]_ , \new_[30678]_ , \new_[30679]_ , \new_[30680]_ ,
    \new_[30681]_ , \new_[30682]_ , \new_[30683]_ , \new_[30684]_ ,
    \new_[30685]_ , \new_[30686]_ , \new_[30687]_ , \new_[30688]_ ,
    \new_[30689]_ , \new_[30690]_ , \new_[30691]_ , \new_[30692]_ ,
    \new_[30693]_ , \new_[30694]_ , \new_[30695]_ , \new_[30696]_ ,
    \new_[30697]_ , \new_[30698]_ , \new_[30699]_ , \new_[30700]_ ,
    \new_[30701]_ , \new_[30702]_ , \new_[30703]_ , \new_[30704]_ ,
    \new_[30705]_ , \new_[30706]_ , \new_[30707]_ , \new_[30708]_ ,
    \new_[30709]_ , \new_[30710]_ , \new_[30711]_ , \new_[30712]_ ,
    \new_[30713]_ , \new_[30714]_ , \new_[30715]_ , \new_[30716]_ ,
    \new_[30717]_ , \new_[30718]_ , \new_[30719]_ , \new_[30720]_ ,
    \new_[30721]_ , \new_[30722]_ , \new_[30723]_ , \new_[30724]_ ,
    \new_[30725]_ , \new_[30726]_ , \new_[30727]_ , \new_[30728]_ ,
    \new_[30729]_ , \new_[30730]_ , \new_[30731]_ , \new_[30732]_ ,
    \new_[30733]_ , \new_[30734]_ , \new_[30735]_ , \new_[30736]_ ,
    \new_[30737]_ , \new_[30738]_ , \new_[30739]_ , \new_[30740]_ ,
    \new_[30741]_ , \new_[30742]_ , \new_[30743]_ , \new_[30744]_ ,
    \new_[30745]_ , \new_[30746]_ , \new_[30747]_ , \new_[30748]_ ,
    \new_[30749]_ , \new_[30750]_ , \new_[30751]_ , \new_[30752]_ ,
    \new_[30753]_ , \new_[30754]_ , \new_[30755]_ , \new_[30756]_ ,
    \new_[30757]_ , \new_[30758]_ , \new_[30759]_ , \new_[30760]_ ,
    \new_[30761]_ , \new_[30762]_ , \new_[30763]_ , \new_[30764]_ ,
    \new_[30765]_ , \new_[30766]_ , \new_[30767]_ , \new_[30768]_ ,
    \new_[30769]_ , \new_[30770]_ , \new_[30771]_ , \new_[30772]_ ,
    \new_[30773]_ , \new_[30774]_ , \new_[30775]_ , \new_[30776]_ ,
    \new_[30777]_ , \new_[30778]_ , \new_[30779]_ , \new_[30780]_ ,
    \new_[30781]_ , \new_[30782]_ , \new_[30783]_ , \new_[30784]_ ,
    \new_[30785]_ , \new_[30786]_ , \new_[30787]_ , \new_[30788]_ ,
    \new_[30789]_ , \new_[30790]_ , \new_[30791]_ , \new_[30792]_ ,
    \new_[30793]_ , \new_[30794]_ , \new_[30795]_ , \new_[30796]_ ,
    \new_[30797]_ , \new_[30798]_ , \new_[30799]_ , \new_[30800]_ ,
    \new_[30801]_ , \new_[30802]_ , \new_[30803]_ , \new_[30804]_ ,
    \new_[30805]_ , \new_[30806]_ , \new_[30807]_ , \new_[30808]_ ,
    \new_[30809]_ , \new_[30810]_ , \new_[30811]_ , \new_[30812]_ ,
    \new_[30813]_ , \new_[30814]_ , \new_[30815]_ , \new_[30816]_ ,
    \new_[30817]_ , \new_[30818]_ , \new_[30819]_ , \new_[30820]_ ,
    \new_[30821]_ , \new_[30822]_ , \new_[30823]_ , \new_[30824]_ ,
    \new_[30825]_ , \new_[30826]_ , \new_[30827]_ , \new_[30828]_ ,
    \new_[30829]_ , \new_[30830]_ , \new_[30831]_ , \new_[30832]_ ,
    \new_[30833]_ , \new_[30834]_ , \new_[30835]_ , \new_[30836]_ ,
    \new_[30837]_ , \new_[30838]_ , \new_[30839]_ , \new_[30840]_ ,
    \new_[30841]_ , \new_[30842]_ , \new_[30843]_ , \new_[30844]_ ,
    \new_[30845]_ , \new_[30846]_ , \new_[30847]_ , \new_[30848]_ ,
    \new_[30849]_ , \new_[30850]_ , \new_[30851]_ , \new_[30852]_ ,
    \new_[30853]_ , \new_[30854]_ , \new_[30855]_ , \new_[30856]_ ,
    \new_[30857]_ , \new_[30858]_ , \new_[30859]_ , \new_[30860]_ ,
    \new_[30861]_ , \new_[30862]_ , \new_[30863]_ , \new_[30864]_ ,
    \new_[30865]_ , \new_[30866]_ , \new_[30867]_ , \new_[30868]_ ,
    \new_[30869]_ , \new_[30870]_ , \new_[30871]_ , \new_[30872]_ ,
    \new_[30873]_ , \new_[30874]_ , \new_[30875]_ , \new_[30876]_ ,
    \new_[30877]_ , \new_[30878]_ , \new_[30879]_ , \new_[30880]_ ,
    \new_[30881]_ , \new_[30882]_ , \new_[30883]_ , \new_[30884]_ ,
    \new_[30885]_ , \new_[30886]_ , \new_[30887]_ , \new_[30888]_ ,
    \new_[30889]_ , \new_[30890]_ , \new_[30891]_ , \new_[30892]_ ,
    \new_[30893]_ , \new_[30894]_ , \new_[30895]_ , \new_[30896]_ ,
    \new_[30897]_ , \new_[30898]_ , \new_[30899]_ , \new_[30900]_ ,
    \new_[30901]_ , \new_[30902]_ , \new_[30903]_ , \new_[30904]_ ,
    \new_[30905]_ , \new_[30906]_ , \new_[30907]_ , \new_[30908]_ ,
    \new_[30909]_ , \new_[30910]_ , \new_[30911]_ , \new_[30912]_ ,
    \new_[30913]_ , \new_[30914]_ , \new_[30915]_ , \new_[30916]_ ,
    \new_[30917]_ , \new_[30918]_ , \new_[30919]_ , \new_[30920]_ ,
    \new_[30921]_ , \new_[30922]_ , \new_[30923]_ , \new_[30924]_ ,
    \new_[30925]_ , \new_[30926]_ , \new_[30927]_ , \new_[30928]_ ,
    \new_[30929]_ , \new_[30930]_ , \new_[30931]_ , \new_[30932]_ ,
    \new_[30933]_ , \new_[30934]_ , \new_[30935]_ , \new_[30936]_ ,
    \new_[30937]_ , \new_[30938]_ , \new_[30939]_ , \new_[30940]_ ,
    \new_[30941]_ , \new_[30942]_ , \new_[30943]_ , \new_[30944]_ ,
    \new_[30945]_ , \new_[30946]_ , \new_[30947]_ , \new_[30948]_ ,
    \new_[30949]_ , \new_[30950]_ , \new_[30951]_ , \new_[30952]_ ,
    \new_[30953]_ , \new_[30954]_ , \new_[30955]_ , \new_[30956]_ ,
    \new_[30957]_ , \new_[30958]_ , \new_[30959]_ , \new_[30960]_ ,
    \new_[30961]_ , \new_[30962]_ , \new_[30963]_ , \new_[30964]_ ,
    \new_[30965]_ , \new_[30966]_ , \new_[30967]_ , \new_[30968]_ ,
    \new_[30969]_ , \new_[30970]_ , \new_[30971]_ , \new_[30972]_ ,
    \new_[30973]_ , \new_[30974]_ , \new_[30975]_ , \new_[30976]_ ,
    \new_[30977]_ , \new_[30978]_ , \new_[30979]_ , \new_[30980]_ ,
    \new_[30981]_ , \new_[30982]_ , \new_[30983]_ , \new_[30984]_ ,
    \new_[30985]_ , \new_[30986]_ , \new_[30987]_ , \new_[30988]_ ,
    \new_[30989]_ , \new_[30990]_ , \new_[30991]_ , \new_[30992]_ ,
    \new_[30993]_ , \new_[30994]_ , \new_[30995]_ , \new_[30996]_ ,
    \new_[30997]_ , \new_[30998]_ , \new_[30999]_ , \new_[31000]_ ,
    \new_[31001]_ , \new_[31002]_ , \new_[31003]_ , \new_[31004]_ ,
    \new_[31005]_ , \new_[31006]_ , \new_[31007]_ , \new_[31008]_ ,
    \new_[31009]_ , \new_[31010]_ , \new_[31011]_ , \new_[31012]_ ,
    \new_[31013]_ , \new_[31014]_ , \new_[31015]_ , \new_[31016]_ ,
    \new_[31017]_ , \new_[31018]_ , \new_[31019]_ , \new_[31020]_ ,
    \new_[31021]_ , \new_[31022]_ , \new_[31023]_ , \new_[31024]_ ,
    \new_[31025]_ , \new_[31026]_ , \new_[31027]_ , \new_[31028]_ ,
    \new_[31029]_ , \new_[31030]_ , \new_[31031]_ , \new_[31032]_ ,
    \new_[31033]_ , \new_[31034]_ , \new_[31035]_ , \new_[31036]_ ,
    \new_[31037]_ , \new_[31038]_ , \new_[31039]_ , \new_[31040]_ ,
    \new_[31041]_ , \new_[31042]_ , \new_[31043]_ , \new_[31044]_ ,
    \new_[31045]_ , \new_[31046]_ , \new_[31047]_ , \new_[31048]_ ,
    \new_[31049]_ , \new_[31050]_ , \new_[31051]_ , \new_[31052]_ ,
    \new_[31053]_ , \new_[31054]_ , \new_[31055]_ , \new_[31056]_ ,
    \new_[31057]_ , \new_[31058]_ , \new_[31059]_ , \new_[31060]_ ,
    \new_[31061]_ , \new_[31062]_ , \new_[31063]_ , \new_[31064]_ ,
    \new_[31065]_ , \new_[31066]_ , \new_[31067]_ , \new_[31068]_ ,
    \new_[31069]_ , \new_[31070]_ , \new_[31071]_ , \new_[31072]_ ,
    \new_[31073]_ , \new_[31074]_ , \new_[31075]_ , \new_[31076]_ ,
    \new_[31077]_ , \new_[31078]_ , \new_[31079]_ , \new_[31080]_ ,
    \new_[31081]_ , \new_[31082]_ , \new_[31083]_ , \new_[31084]_ ,
    \new_[31085]_ , \new_[31086]_ , \new_[31087]_ , \new_[31088]_ ,
    \new_[31089]_ , \new_[31090]_ , \new_[31091]_ , \new_[31092]_ ,
    \new_[31093]_ , \new_[31094]_ , \new_[31095]_ , \new_[31096]_ ,
    \new_[31097]_ , \new_[31098]_ , \new_[31099]_ , \new_[31100]_ ,
    \new_[31101]_ , \new_[31102]_ , \new_[31103]_ , \new_[31104]_ ,
    \new_[31105]_ , \new_[31106]_ , \new_[31107]_ , \new_[31108]_ ,
    \new_[31109]_ , \new_[31110]_ , \new_[31111]_ , \new_[31112]_ ,
    \new_[31113]_ , \new_[31114]_ , \new_[31115]_ , \new_[31116]_ ,
    \new_[31117]_ , \new_[31118]_ , \new_[31119]_ , \new_[31120]_ ,
    \new_[31121]_ , \new_[31122]_ , \new_[31123]_ , \new_[31124]_ ,
    \new_[31125]_ , \new_[31126]_ , \new_[31127]_ , \new_[31128]_ ,
    \new_[31129]_ , \new_[31130]_ , \new_[31131]_ , \new_[31132]_ ,
    \new_[31133]_ , \new_[31134]_ , \new_[31135]_ , \new_[31136]_ ,
    \new_[31137]_ , \new_[31138]_ , \new_[31139]_ , \new_[31140]_ ,
    \new_[31141]_ , \new_[31142]_ , \new_[31143]_ , \new_[31144]_ ,
    \new_[31145]_ , \new_[31146]_ , \new_[31147]_ , \new_[31148]_ ,
    \new_[31149]_ , \new_[31150]_ , \new_[31151]_ , \new_[31152]_ ,
    \new_[31153]_ , \new_[31154]_ , \new_[31155]_ , \new_[31156]_ ,
    \new_[31157]_ , \new_[31158]_ , \new_[31159]_ , \new_[31160]_ ,
    \new_[31161]_ , \new_[31162]_ , \new_[31163]_ , \new_[31164]_ ,
    \new_[31165]_ , \new_[31166]_ , \new_[31167]_ , \new_[31168]_ ,
    \new_[31169]_ , \new_[31170]_ , \new_[31171]_ , \new_[31172]_ ,
    \new_[31173]_ , \new_[31174]_ , \new_[31175]_ , \new_[31176]_ ,
    \new_[31177]_ , \new_[31178]_ , \new_[31179]_ , \new_[31180]_ ,
    \new_[31181]_ , \new_[31182]_ , \new_[31183]_ , \new_[31184]_ ,
    \new_[31185]_ , \new_[31186]_ , \new_[31187]_ , \new_[31188]_ ,
    \new_[31189]_ , \new_[31190]_ , \new_[31191]_ , \new_[31192]_ ,
    \new_[31193]_ , \new_[31194]_ , \new_[31195]_ , \new_[31196]_ ,
    \new_[31197]_ , \new_[31198]_ , \new_[31199]_ , \new_[31200]_ ,
    \new_[31201]_ , \new_[31202]_ , \new_[31203]_ , \new_[31204]_ ,
    \new_[31205]_ , \new_[31206]_ , \new_[31207]_ , \new_[31208]_ ,
    \new_[31209]_ , \new_[31210]_ , \new_[31211]_ , \new_[31212]_ ,
    \new_[31213]_ , \new_[31214]_ , \new_[31215]_ , \new_[31216]_ ,
    \new_[31217]_ , \new_[31218]_ , \new_[31219]_ , \new_[31220]_ ,
    \new_[31221]_ , \new_[31222]_ , \new_[31223]_ , \new_[31224]_ ,
    \new_[31225]_ , \new_[31226]_ , \new_[31227]_ , \new_[31228]_ ,
    \new_[31229]_ , \new_[31230]_ , \new_[31231]_ , \new_[31232]_ ,
    \new_[31233]_ , \new_[31234]_ , \new_[31235]_ , \new_[31236]_ ,
    \new_[31237]_ , \new_[31238]_ , \new_[31239]_ , \new_[31240]_ ,
    \new_[31241]_ , \new_[31242]_ , \new_[31243]_ , \new_[31244]_ ,
    \new_[31245]_ , \new_[31246]_ , \new_[31247]_ , \new_[31248]_ ,
    \new_[31249]_ , \new_[31250]_ , \new_[31251]_ , \new_[31252]_ ,
    \new_[31253]_ , \new_[31254]_ , \new_[31255]_ , \new_[31256]_ ,
    \new_[31257]_ , \new_[31258]_ , \new_[31259]_ , \new_[31260]_ ,
    \new_[31261]_ , \new_[31262]_ , \new_[31263]_ , \new_[31264]_ ,
    \new_[31265]_ , \new_[31266]_ , \new_[31267]_ , \new_[31268]_ ,
    \new_[31269]_ , \new_[31270]_ , \new_[31271]_ , \new_[31272]_ ,
    \new_[31273]_ , \new_[31274]_ , \new_[31275]_ , \new_[31276]_ ,
    \new_[31277]_ , \new_[31278]_ , \new_[31279]_ , \new_[31280]_ ,
    \new_[31281]_ , \new_[31282]_ , \new_[31283]_ , \new_[31284]_ ,
    \new_[31285]_ , \new_[31286]_ , \new_[31287]_ , \new_[31288]_ ,
    \new_[31289]_ , \new_[31290]_ , \new_[31291]_ , \new_[31292]_ ,
    \new_[31293]_ , \new_[31294]_ , \new_[31295]_ , \new_[31296]_ ,
    \new_[31297]_ , \new_[31298]_ , \new_[31299]_ , \new_[31300]_ ,
    \new_[31301]_ , \new_[31302]_ , \new_[31303]_ , \new_[31304]_ ,
    \new_[31305]_ , \new_[31306]_ , \new_[31307]_ , \new_[31308]_ ,
    \new_[31309]_ , \new_[31310]_ , \new_[31311]_ , \new_[31312]_ ,
    \new_[31313]_ , \new_[31314]_ , \new_[31315]_ , \new_[31316]_ ,
    \new_[31317]_ , \new_[31318]_ , \new_[31319]_ , \new_[31320]_ ,
    \new_[31321]_ , \new_[31322]_ , \new_[31323]_ , \new_[31324]_ ,
    \new_[31325]_ , \new_[31326]_ , \new_[31327]_ , \new_[31328]_ ,
    \new_[31329]_ , \new_[31330]_ , \new_[31331]_ , \new_[31332]_ ,
    \new_[31333]_ , \new_[31334]_ , \new_[31335]_ , \new_[31336]_ ,
    \new_[31337]_ , \new_[31338]_ , \new_[31339]_ , \new_[31340]_ ,
    \new_[31341]_ , \new_[31342]_ , \new_[31343]_ , \new_[31344]_ ,
    \new_[31345]_ , \new_[31346]_ , \new_[31347]_ , \new_[31348]_ ,
    \new_[31349]_ , \new_[31350]_ , \new_[31351]_ , \new_[31352]_ ,
    \new_[31353]_ , \new_[31354]_ , \new_[31355]_ , \new_[31356]_ ,
    \new_[31357]_ , \new_[31358]_ , \new_[31359]_ , \new_[31360]_ ,
    \new_[31361]_ , \new_[31362]_ , \new_[31363]_ , \new_[31364]_ ,
    \new_[31365]_ , \new_[31366]_ , \new_[31367]_ , \new_[31368]_ ,
    \new_[31369]_ , \new_[31370]_ , \new_[31371]_ , \new_[31372]_ ,
    \new_[31373]_ , \new_[31374]_ , \new_[31375]_ , \new_[31376]_ ,
    \new_[31377]_ , \new_[31378]_ , \new_[31379]_ , \new_[31380]_ ,
    \new_[31381]_ , \new_[31382]_ , \new_[31383]_ , \new_[31384]_ ,
    \new_[31385]_ , \new_[31386]_ , \new_[31387]_ , \new_[31388]_ ,
    \new_[31389]_ , \new_[31390]_ , \new_[31391]_ , \new_[31392]_ ,
    \new_[31393]_ , \new_[31394]_ , \new_[31395]_ , \new_[31396]_ ,
    \new_[31397]_ , \new_[31398]_ , \new_[31399]_ , \new_[31400]_ ,
    \new_[31401]_ , \new_[31402]_ , \new_[31403]_ , \new_[31404]_ ,
    \new_[31405]_ , \new_[31406]_ , \new_[31407]_ , \new_[31408]_ ,
    \new_[31409]_ , \new_[31410]_ , \new_[31411]_ , \new_[31412]_ ,
    \new_[31413]_ , \new_[31414]_ , \new_[31415]_ , \new_[31416]_ ,
    \new_[31417]_ , \new_[31418]_ , \new_[31419]_ , \new_[31420]_ ,
    \new_[31421]_ , \new_[31422]_ , \new_[31423]_ , \new_[31424]_ ,
    \new_[31425]_ , \new_[31426]_ , \new_[31427]_ , \new_[31428]_ ,
    \new_[31429]_ , \new_[31430]_ , \new_[31431]_ , \new_[31432]_ ,
    \new_[31433]_ , \new_[31434]_ , \new_[31435]_ , \new_[31436]_ ,
    \new_[31437]_ , \new_[31438]_ , \new_[31439]_ , \new_[31440]_ ,
    \new_[31441]_ , \new_[31442]_ , \new_[31443]_ , \new_[31444]_ ,
    \new_[31445]_ , \new_[31446]_ , \new_[31447]_ , \new_[31448]_ ,
    \new_[31449]_ , \new_[31450]_ , \new_[31451]_ , \new_[31452]_ ,
    \new_[31453]_ , \new_[31454]_ , \new_[31455]_ , \new_[31456]_ ,
    \new_[31457]_ , \new_[31458]_ , \new_[31459]_ , \new_[31460]_ ,
    \new_[31461]_ , \new_[31462]_ , \new_[31463]_ , \new_[31464]_ ,
    \new_[31465]_ , \new_[31466]_ , \new_[31467]_ , \new_[31468]_ ,
    \new_[31469]_ , \new_[31470]_ , \new_[31471]_ , \new_[31472]_ ,
    \new_[31473]_ , \new_[31474]_ , \new_[31475]_ , \new_[31476]_ ,
    \new_[31477]_ , \new_[31478]_ , \new_[31479]_ , \new_[31480]_ ,
    \new_[31481]_ , \new_[31482]_ , \new_[31483]_ , \new_[31484]_ ,
    \new_[31485]_ , \new_[31486]_ , \new_[31487]_ , \new_[31488]_ ,
    \new_[31489]_ , \new_[31490]_ , \new_[31491]_ , \new_[31492]_ ,
    \new_[31493]_ , \new_[31494]_ , \new_[31495]_ , \new_[31496]_ ,
    \new_[31497]_ , \new_[31498]_ , \new_[31499]_ , \new_[31500]_ ,
    \new_[31501]_ , \new_[31502]_ , \new_[31503]_ , \new_[31504]_ ,
    \new_[31505]_ , \new_[31506]_ , \new_[31507]_ , \new_[31508]_ ,
    \new_[31509]_ , \new_[31510]_ , \new_[31511]_ , \new_[31512]_ ,
    \new_[31513]_ , \new_[31514]_ , \new_[31515]_ , \new_[31516]_ ,
    \new_[31517]_ , \new_[31518]_ , \new_[31519]_ , \new_[31520]_ ,
    \new_[31521]_ , \new_[31522]_ , \new_[31523]_ , \new_[31524]_ ,
    \new_[31525]_ , \new_[31526]_ , \new_[31527]_ , \new_[31528]_ ,
    \new_[31529]_ , \new_[31530]_ , \new_[31531]_ , \new_[31532]_ ,
    \new_[31533]_ , \new_[31534]_ , \new_[31535]_ , \new_[31536]_ ,
    \new_[31537]_ , \new_[31538]_ , \new_[31539]_ , \new_[31540]_ ,
    \new_[31541]_ , \new_[31542]_ , \new_[31543]_ , \new_[31544]_ ,
    \new_[31545]_ , \new_[31546]_ , \new_[31547]_ , \new_[31548]_ ,
    \new_[31549]_ , \new_[31550]_ , \new_[31551]_ , \new_[31552]_ ,
    \new_[31553]_ , \new_[31554]_ , \new_[31555]_ , \new_[31556]_ ,
    \new_[31557]_ , \new_[31558]_ , \new_[31559]_ , \new_[31560]_ ,
    \new_[31561]_ , \new_[31562]_ , \new_[31563]_ , \new_[31564]_ ,
    \new_[31565]_ , \new_[31566]_ , \new_[31567]_ , \new_[31568]_ ,
    \new_[31569]_ , \new_[31570]_ , \new_[31571]_ , \new_[31572]_ ,
    \new_[31573]_ , \new_[31574]_ , \new_[31575]_ , \new_[31576]_ ,
    \new_[31577]_ , \new_[31578]_ , \new_[31579]_ , \new_[31580]_ ,
    \new_[31581]_ , \new_[31582]_ , \new_[31583]_ , \new_[31584]_ ,
    \new_[31585]_ , \new_[31586]_ , \new_[31587]_ , \new_[31588]_ ,
    \new_[31589]_ , \new_[31590]_ , \new_[31591]_ , \new_[31592]_ ,
    \new_[31593]_ , \new_[31594]_ , \new_[31595]_ , \new_[31596]_ ,
    \new_[31597]_ , \new_[31598]_ , \new_[31599]_ , \new_[31600]_ ,
    \new_[31601]_ , \new_[31602]_ , \new_[31603]_ , \new_[31604]_ ,
    \new_[31605]_ , \new_[31606]_ , \new_[31607]_ , \new_[31608]_ ,
    \new_[31609]_ , \new_[31610]_ , \new_[31611]_ , \new_[31612]_ ,
    \new_[31613]_ , \new_[31614]_ , \new_[31615]_ , \new_[31616]_ ,
    \new_[31617]_ , \new_[31618]_ , \new_[31619]_ , \new_[31620]_ ,
    \new_[31621]_ , \new_[31622]_ , \new_[31623]_ , \new_[31624]_ ,
    \new_[31625]_ , \new_[31626]_ , \new_[31627]_ , \new_[31628]_ ,
    \new_[31629]_ , \new_[31630]_ , \new_[31631]_ , \new_[31632]_ ,
    \new_[31633]_ , \new_[31634]_ , \new_[31635]_ , \new_[31636]_ ,
    \new_[31637]_ , \new_[31638]_ , \new_[31639]_ , \new_[31640]_ ,
    \new_[31641]_ , \new_[31642]_ , \new_[31643]_ , \new_[31644]_ ,
    \new_[31645]_ , \new_[31646]_ , \new_[31647]_ , \new_[31648]_ ,
    \new_[31649]_ , \new_[31650]_ , \new_[31651]_ , \new_[31652]_ ,
    \new_[31653]_ , \new_[31654]_ , \new_[31655]_ , \new_[31656]_ ,
    \new_[31657]_ , \new_[31658]_ , \new_[31659]_ , \new_[31660]_ ,
    \new_[31661]_ , \new_[31662]_ , \new_[31663]_ , \new_[31664]_ ,
    \new_[31665]_ , \new_[31666]_ , \new_[31667]_ , \new_[31668]_ ,
    \new_[31669]_ , \new_[31670]_ , \new_[31671]_ , \new_[31672]_ ,
    \new_[31673]_ , \new_[31674]_ , \new_[31675]_ , \new_[31676]_ ,
    \new_[31677]_ , \new_[31678]_ , \new_[31679]_ , \new_[31680]_ ,
    \new_[31681]_ , \new_[31682]_ , \new_[31683]_ , \new_[31684]_ ,
    \new_[31685]_ , \new_[31686]_ , \new_[31687]_ , \new_[31688]_ ,
    \new_[31689]_ , \new_[31690]_ , \new_[31691]_ , \new_[31692]_ ,
    \new_[31693]_ , \new_[31694]_ , \new_[31695]_ , \new_[31696]_ ,
    \new_[31697]_ , \new_[31698]_ , \new_[31699]_ , \new_[31700]_ ,
    \new_[31701]_ , \new_[31702]_ , \new_[31703]_ , \new_[31704]_ ,
    \new_[31705]_ , \new_[31706]_ , \new_[31707]_ , \new_[31708]_ ,
    \new_[31709]_ , \new_[31710]_ , \new_[31711]_ , \new_[31712]_ ,
    \new_[31713]_ , \new_[31714]_ , \new_[31715]_ , \new_[31716]_ ,
    \new_[31717]_ , \new_[31718]_ , \new_[31719]_ , \new_[31720]_ ,
    \new_[31721]_ , \new_[31722]_ , \new_[31723]_ , \new_[31724]_ ,
    \new_[31725]_ , \new_[31726]_ , \new_[31727]_ , \new_[31728]_ ,
    \new_[31729]_ , \new_[31730]_ , \new_[31731]_ , \new_[31732]_ ,
    \new_[31733]_ , \new_[31734]_ , \new_[31735]_ , \new_[31736]_ ,
    \new_[31737]_ , \new_[31738]_ , \new_[31739]_ , \new_[31740]_ ,
    \new_[31741]_ , \new_[31742]_ , \new_[31743]_ , \new_[31744]_ ,
    \new_[31745]_ , \new_[31746]_ , \new_[31747]_ , \new_[31748]_ ,
    \new_[31749]_ , \new_[31750]_ , \new_[31751]_ , \new_[31752]_ ,
    \new_[31753]_ , \new_[31754]_ , \new_[31755]_ , \new_[31756]_ ,
    \new_[31757]_ , \new_[31758]_ , \new_[31759]_ , \new_[31760]_ ,
    \new_[31761]_ , \new_[31762]_ , \new_[31763]_ , \new_[31764]_ ,
    \new_[31765]_ , \new_[31766]_ , \new_[31767]_ , \new_[31768]_ ,
    \new_[31769]_ , \new_[31770]_ , \new_[31771]_ , \new_[31772]_ ,
    \new_[31773]_ , \new_[31774]_ , \new_[31775]_ , \new_[31776]_ ,
    \new_[31777]_ , \new_[31778]_ , \new_[31779]_ , \new_[31780]_ ,
    \new_[31781]_ , \new_[31782]_ , \new_[31783]_ , \new_[31784]_ ,
    \new_[31785]_ , \new_[31786]_ , \new_[31787]_ , \new_[31788]_ ,
    \new_[31789]_ , \new_[31790]_ , \new_[31791]_ , \new_[31792]_ ,
    \new_[31793]_ , \new_[31794]_ , \new_[31795]_ , \new_[31796]_ ,
    \new_[31797]_ , \new_[31798]_ , \new_[31799]_ , \new_[31800]_ ,
    \new_[31801]_ , \new_[31802]_ , \new_[31803]_ , \new_[31804]_ ,
    \new_[31805]_ , \new_[31806]_ , \new_[31807]_ , \new_[31808]_ ,
    \new_[31809]_ , \new_[31810]_ , \new_[31811]_ , \new_[31812]_ ,
    \new_[31813]_ , \new_[31814]_ , \new_[31815]_ , \new_[31816]_ ,
    \new_[31817]_ , \new_[31818]_ , \new_[31819]_ , \new_[31820]_ ,
    \new_[31821]_ , \new_[31822]_ , \new_[31823]_ , \new_[31824]_ ,
    \new_[31825]_ , \new_[31826]_ , \new_[31827]_ , \new_[31828]_ ,
    \new_[31829]_ , \new_[31830]_ , \new_[31831]_ , \new_[31832]_ ,
    \new_[31833]_ , \new_[31834]_ , \new_[31835]_ , \new_[31836]_ ,
    \new_[31837]_ , \new_[31838]_ , \new_[31839]_ , \new_[31840]_ ,
    \new_[31841]_ , \new_[31842]_ , \new_[31843]_ , \new_[31844]_ ,
    \new_[31845]_ , \new_[31846]_ , \new_[31847]_ , \new_[31848]_ ,
    \new_[31849]_ , \new_[31850]_ , \new_[31851]_ , \new_[31852]_ ,
    \new_[31853]_ , \new_[31854]_ , \new_[31855]_ , \new_[31856]_ ,
    \new_[31857]_ , \new_[31858]_ , \new_[31859]_ , \new_[31860]_ ,
    \new_[31861]_ , \new_[31862]_ , \new_[31863]_ , \new_[31864]_ ,
    \new_[31865]_ , \new_[31866]_ , \new_[31867]_ , \new_[31868]_ ,
    \new_[31869]_ , \new_[31870]_ , \new_[31871]_ , \new_[31872]_ ,
    \new_[31873]_ , \new_[31874]_ , \new_[31875]_ , \new_[31876]_ ,
    \new_[31877]_ , \new_[31878]_ , \new_[31879]_ , \new_[31880]_ ,
    \new_[31881]_ , \new_[31882]_ , \new_[31883]_ , \new_[31884]_ ,
    \new_[31885]_ , \new_[31886]_ , \new_[31887]_ , \new_[31888]_ ,
    \new_[31889]_ , \new_[31890]_ , \new_[31891]_ , \new_[31892]_ ,
    \new_[31893]_ , \new_[31894]_ , \new_[31895]_ , \new_[31896]_ ,
    \new_[31897]_ , \new_[31898]_ , \new_[31899]_ , \new_[31900]_ ,
    \new_[31901]_ , \new_[31902]_ , \new_[31903]_ , \new_[31904]_ ,
    \new_[31905]_ , \new_[31906]_ , \new_[31907]_ , \new_[31908]_ ,
    \new_[31909]_ , \new_[31910]_ , \new_[31911]_ , \new_[31912]_ ,
    \new_[31913]_ , \new_[31914]_ , \new_[31915]_ , \new_[31916]_ ,
    \new_[31917]_ , \new_[31918]_ , \new_[31919]_ , \new_[31920]_ ,
    \new_[31921]_ , \new_[31922]_ , \new_[31923]_ , \new_[31924]_ ,
    \new_[31925]_ , \new_[31926]_ , \new_[31927]_ , \new_[31928]_ ,
    \new_[31929]_ , \new_[31930]_ , \new_[31931]_ , \new_[31932]_ ,
    \new_[31933]_ , \new_[31934]_ , \new_[31935]_ , \new_[31936]_ ,
    \new_[31937]_ , \new_[31938]_ , \new_[31939]_ , \new_[31940]_ ,
    \new_[31941]_ , \new_[31943]_ , \new_[31944]_ , \new_[31945]_ ,
    \new_[31946]_ , \new_[31947]_ , \new_[31948]_ , \new_[31949]_ ,
    \new_[31950]_ , \new_[31951]_ , \new_[31952]_ , \new_[31953]_ ,
    \new_[31954]_ , \new_[31955]_ , \new_[31956]_ , \new_[31957]_ ,
    \new_[31958]_ , \new_[31959]_ , \new_[31960]_ , \new_[31961]_ ,
    \new_[31962]_ , \new_[31963]_ , \new_[31964]_ , \new_[31965]_ ,
    \new_[31966]_ , \new_[31967]_ , \new_[31968]_ , \new_[31969]_ ,
    \new_[31970]_ , \new_[31971]_ , \new_[31972]_ , \new_[31973]_ ,
    \new_[31974]_ , \new_[31975]_ , \new_[31976]_ , \new_[31977]_ ,
    \new_[31978]_ , \new_[31979]_ , \new_[31980]_ , \new_[31981]_ ,
    \new_[31982]_ , \new_[31983]_ , \new_[31984]_ , \new_[31985]_ ,
    \new_[31986]_ , \new_[31987]_ , \new_[31988]_ , \new_[31989]_ ,
    \new_[31990]_ , \new_[31991]_ , \new_[31992]_ , \new_[31993]_ ,
    \new_[31994]_ , \new_[31995]_ , \new_[31996]_ , \new_[31997]_ ,
    \new_[31998]_ , \new_[31999]_ , \new_[32000]_ , \new_[32001]_ ,
    \new_[32002]_ , \new_[32003]_ , \new_[32004]_ , \new_[32005]_ ,
    \new_[32006]_ , \new_[32007]_ , \new_[32008]_ , \new_[32009]_ ,
    \new_[32010]_ , \new_[32011]_ , \new_[32012]_ , \new_[32014]_ ,
    \new_[32015]_ , \new_[32016]_ , \new_[32017]_ , \new_[32018]_ ,
    \new_[32019]_ , \new_[32020]_ , \new_[32021]_ , \new_[32022]_ ,
    \new_[32023]_ , \new_[32025]_ , \new_[32026]_ , \new_[32027]_ ,
    \new_[32028]_ , \new_[32029]_ , \new_[32030]_ , \new_[32031]_ ,
    \new_[32032]_ , \new_[32033]_ , \new_[32034]_ , \new_[32036]_ ,
    \new_[32037]_ , \new_[32038]_ , \new_[32039]_ , \new_[32040]_ ,
    \new_[32041]_ , \new_[32042]_ , \new_[32043]_ , \new_[32044]_ ,
    \new_[32045]_ , \new_[32046]_ , \new_[32047]_ , \new_[32048]_ ,
    \new_[32049]_ , \new_[32050]_ , \new_[32051]_ , \new_[32052]_ ,
    \new_[32053]_ , \new_[32054]_ , \new_[32055]_ , \new_[32056]_ ,
    \new_[32057]_ , \new_[32058]_ , \new_[32059]_ , \new_[32060]_ ,
    \new_[32061]_ , \new_[32062]_ , \new_[32063]_ , \new_[32064]_ ,
    \new_[32065]_ , \new_[32066]_ , \new_[32067]_ , \new_[32068]_ ,
    \new_[32069]_ , \new_[32070]_ , \new_[32072]_ , \new_[32073]_ ,
    \new_[32074]_ , \new_[32075]_ , \new_[32076]_ , \new_[32077]_ ,
    \new_[32078]_ , \new_[32079]_ , \new_[32080]_ , \new_[32081]_ ,
    \new_[32082]_ , \new_[32083]_ , \new_[32084]_ , \new_[32085]_ ,
    \new_[32086]_ , \new_[32087]_ , \new_[32088]_ , \new_[32089]_ ,
    \new_[32090]_ , \new_[32092]_ , \new_[32093]_ , \new_[32094]_ ,
    \new_[32095]_ , \new_[32096]_ , \new_[32097]_ , \new_[32098]_ ,
    \new_[32099]_ , \new_[32100]_ , \new_[32101]_ , \new_[32103]_ ,
    \new_[32104]_ , \new_[32105]_ , \new_[32106]_ , \new_[32107]_ ,
    \new_[32108]_ , \new_[32109]_ , \new_[32110]_ , \new_[32111]_ ,
    \new_[32112]_ , \new_[32114]_ , \new_[32115]_ , \new_[32116]_ ,
    \new_[32117]_ , \new_[32118]_ , \new_[32119]_ , \new_[32120]_ ,
    \new_[32121]_ , \new_[32122]_ , \new_[32123]_ , \new_[32124]_ ,
    \new_[32125]_ , \new_[32126]_ , \new_[32127]_ , \new_[32128]_ ,
    \new_[32129]_ , \new_[32130]_ , \new_[32131]_ , \new_[32132]_ ,
    \new_[32133]_ , \new_[32134]_ , \new_[32135]_ , \new_[32137]_ ,
    \new_[32138]_ , \new_[32139]_ , \new_[32140]_ , \new_[32141]_ ,
    \new_[32142]_ , \new_[32143]_ , \new_[32144]_ , \new_[32145]_ ,
    \new_[32146]_ , \new_[32148]_ , \new_[32149]_ , \new_[32150]_ ,
    \new_[32151]_ , \new_[32152]_ , \new_[32153]_ , \new_[32154]_ ,
    \new_[32155]_ , \new_[32156]_ , \new_[32157]_ , \new_[32158]_ ,
    \new_[32159]_ , \new_[32160]_ , \new_[32161]_ , \new_[32162]_ ,
    \new_[32163]_ , \new_[32164]_ , \new_[32165]_ , \new_[32166]_ ,
    \new_[32167]_ , \new_[32168]_ , \new_[32169]_ , \new_[32170]_ ,
    \new_[32171]_ , \new_[32172]_ , \new_[32173]_ , \new_[32174]_ ,
    \new_[32175]_ , \new_[32176]_ , \new_[32177]_ , \new_[32178]_ ,
    \new_[32179]_ , \new_[32180]_ , \new_[32181]_ , \new_[32182]_ ,
    \new_[32183]_ , \new_[32184]_ , \new_[32185]_ , \new_[32186]_ ,
    \new_[32187]_ , \new_[32188]_ , \new_[32189]_ , \new_[32190]_ ,
    \new_[32191]_ , \new_[32192]_ , \new_[32193]_ , \new_[32195]_ ,
    \new_[32196]_ , \new_[32197]_ , \new_[32198]_ , \new_[32199]_ ,
    \new_[32200]_ , \new_[32201]_ , \new_[32202]_ , \new_[32203]_ ,
    \new_[32204]_ , \new_[32206]_ , \new_[32207]_ , \new_[32208]_ ,
    \new_[32209]_ , \new_[32210]_ , \new_[32211]_ , \new_[32212]_ ,
    \new_[32213]_ , \new_[32214]_ , \new_[32215]_ , \new_[32216]_ ,
    \new_[32217]_ , \new_[32218]_ , \new_[32219]_ , \new_[32220]_ ,
    \new_[32221]_ , \new_[32222]_ , \new_[32223]_ , \new_[32225]_ ,
    \new_[32226]_ , \new_[32227]_ , \new_[32228]_ , \new_[32229]_ ,
    \new_[32230]_ , \new_[32231]_ , \new_[32232]_ , \new_[32233]_ ,
    \new_[32234]_ , \new_[32236]_ , \new_[32237]_ , \new_[32238]_ ,
    \new_[32239]_ , \new_[32240]_ , \new_[32241]_ , \new_[32242]_ ,
    \new_[32243]_ , \new_[32244]_ , \new_[32245]_ , \new_[32247]_ ,
    \new_[32248]_ , \new_[32249]_ , \new_[32250]_ , \new_[32251]_ ,
    \new_[32252]_ , \new_[32253]_ , \new_[32254]_ , \new_[32255]_ ,
    \new_[32256]_ , \new_[32257]_ , \new_[32258]_ , \new_[32259]_ ,
    \new_[32260]_ , \new_[32261]_ , \new_[32262]_ , \new_[32263]_ ,
    \new_[32264]_ , \new_[32265]_ , \new_[32266]_ , \new_[32267]_ ,
    \new_[32268]_ , \new_[32269]_ , \new_[32270]_ , \new_[32271]_ ,
    \new_[32272]_ , \new_[32273]_ , \new_[32274]_ , \new_[32275]_ ,
    \new_[32276]_ , \new_[32277]_ , \new_[32278]_ , \new_[32279]_ ,
    \new_[32280]_ , \new_[32281]_ , \new_[32282]_ , \new_[32283]_ ,
    \new_[32284]_ , \new_[32285]_ , \new_[32286]_ , \new_[32287]_ ,
    \new_[32288]_ , \new_[32289]_ , \new_[32291]_ , \new_[32293]_ ,
    \new_[32294]_ , \new_[32295]_ , \new_[32296]_ , \new_[32297]_ ,
    \new_[32298]_ , \new_[32299]_ , \new_[32300]_ , \new_[32301]_ ,
    \new_[32302]_ , \new_[32303]_ , \new_[32304]_ , \new_[32305]_ ,
    \new_[32306]_ , \new_[32307]_ , \new_[32308]_ , \new_[32309]_ ,
    \new_[32310]_ , \new_[32311]_ , \new_[32312]_ , \new_[32313]_ ,
    \new_[32314]_ , \new_[32315]_ , \new_[32316]_ , \new_[32317]_ ,
    \new_[32318]_ , \new_[32319]_ , \new_[32320]_ , \new_[32321]_ ,
    \new_[32322]_ , \new_[32323]_ , \new_[32324]_ , \new_[32325]_ ,
    \new_[32326]_ , \new_[32327]_ , \new_[32328]_ , \new_[32329]_ ,
    \new_[32330]_ , \new_[32331]_ , \new_[32333]_ , \new_[32335]_ ,
    \new_[32336]_ , \new_[32337]_ , \new_[32338]_ , \new_[32339]_ ,
    \new_[32340]_ , \new_[32341]_ , \new_[32342]_ , \new_[32343]_ ,
    \new_[32344]_ , \new_[32345]_ , \new_[32346]_ , \new_[32347]_ ,
    \new_[32348]_ , \new_[32349]_ , \new_[32350]_ , \new_[32351]_ , n5094,
    n5099, n5104, n5109, n5114, n5119, n5124, n5129, n5134, n5139, n5144,
    n5149, n5154, n5159, n5164, n5169, n5174, n5179, n5184, n5189, n5194,
    n5199, n5204, n5209, n5214, n5219, n5224, n5229, n5234, n5239, n5244,
    n5249, n5254, n5259, n5264, n5269, n5274, n5279, n5284, n5289, n5294,
    n5299, n5304, n5309, n5314, n5319, n5324, n5329, n5334, n5339, n5344,
    n5349, n5354, n5359, n5364, n5369, n5374, n5379, n5384, n5389, n5394,
    n5399, n5404, n5409, n5414, n5419, n5424, n5429, n5434, n5439, n5444,
    n5449, n5454, n5459, n5464, n5469, n5474, n5479, n5484, n5489, n5494,
    n5499, n5504, n5509, n5514, n5519, n5524, n5529, n5534, n5539, n5544,
    n5549, n5554, n5559, n5564, n5569, n5574, n5579, n5584, n5589, n5594,
    n5599, n5604, n5609, n5614, n5619, n5624, n5629, n5634, n5639, n5644,
    n5649, n5654, n5659, n5664, n5669, n5674, n5679, n5684, n5689, n5694,
    n5699, n5704, n5709, n5714, n5719, n5724, n5729, n5734, n5739, n5744,
    n5749, n5754, n5759, n5764, n5769, n5774, n5779, n5784, n5789, n5794,
    n5799, n5804, n5809, n5814, n5819, n5824, n5829, n5834, n5839, n5844,
    n5849, n5854, n5859, n5864, n5869, n5874, n5879, n5884, n5889, n5894,
    n5899, n5904, n5909, n5914, n5919, n5924, n5929, n5934, n5939, n5944,
    n5949, n5954, n5959, n5964, n5969, n5974, n5979, n5984, n5989, n5994,
    n5999, n6004, n6009, n6014, n6019, n6024, n6029, n6034, n6039, n6044,
    n6049, n6054, n6059, n6064, n6069, n6074, n6079, n6084, n6089, n6094,
    n6099, n6104, n6109, n6114, n6119, n6124, n6129, n6134, n6139, n6144,
    n6149, n6154, n6159, n6164, n6169, n6174, n6179, n6184, n6189, n6194,
    n6199, n6204, n6209, n6214, n6219, n6224, n6229, n6234, n6239, n6244,
    n6249, n6254, n6259, n6264, n6269, n6274, n6279, n6284, n6289, n6294,
    n6299, n6304, n6309, n6314, n6319, n6324, n6329, n6334, n6339, n6344,
    n6349, n6354, n6359, n6364, n6369, n6374, n6379, n6384, n6389, n6394,
    n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444,
    n6449, n6454, n6459, n6464, n6469, n6474, n6479, n6484, n6489, n6494,
    n6499, n6504, n6509, n6514, n6519, n6524, n6529, n6534, n6539, n6544,
    n6549, n6554, n6559, n6564, n6569, n6574, n6579, n6584, n6589, n6594,
    n6599, n6604, n6609, n6614, n6619, n6624, n6629, n6634, n6639, n6644,
    n6649, n6654, n6659, n6664, n6669, n6674, n6679, n6684, n6689, n6694,
    n6699, n6704, n6709, n6714, n6719, n6724, n6729, n6734, n6739, n6744,
    n6749, n6754, n6759, n6764, n6769, n6774, n6779, n6784, n6789, n6794,
    n6799, n6804, n6809, n6814, n6819, n6824, n6829, n6834, n6839, n6844,
    n6849, n6854, n6859, n6864, n6869, n6874, n6879, n6884, n6889, n6894,
    n6899, n6904, n6909, n6914, n6919, n6924, n6929, n6934, n6939, n6944,
    n6949, n6954, n6959, n6964, n6969, n6974, n6979, n6984, n6989, n6994,
    n6999, n7004, n7009, n7014, n7019, n7024, n7029, n7034, n7039, n7044,
    n7049, n7054, n7059, n7064, n7069, n7074, n7079, n7084, n7089, n7094,
    n7099, n7104, n7109, n7114, n7119, n7124, n7129, n7134, n7139, n7144,
    n7149, n7154, n7159, n7164, n7169, n7174, n7179, n7184, n7189, n7194,
    n7199, n7204, n7209, n7214, n7219, n7224, n7229, n7234, n7239, n7244,
    n7249, n7254, n7259, n7264, n7269, n7274, n7279, n7284, n7289, n7294,
    n7299, n7304, n7309, n7314, n7319, n7324, n7329, n7334, n7339, n7344,
    n7349, n7354, n7359, n7364, n7369, n7374, n7379, n7384, n7389, n7394,
    n7399, n7404, n7409, n7414, n7419, n7424, n7429, n7434, n7439, n7444,
    n7449, n7454, n7459, n7464, n7469, n7474, n7479, n7484, n7489, n7494,
    n7499, n7504, n7509, n7514, n7519, n7524, n7529, n7534, n7539, n7544,
    n7549, n7554, n7559, n7564, n7569, n7574, n7579, n7584, n7589, n7594,
    n7599, n7604, n7609, n7614, n7619, n7624, n7629, n7634, n7639, n7644,
    n7649, n7654, n7659, n7664, n7669, n7674, n7679, n7684, n7689, n7694,
    n7699, n7704, n7709, n7714, n7719, n7724, n7729, n7734, n7739, n7744,
    n7749, n7754, n7759, n7764, n7769, n7774, n7779, n7784, n7789, n7794,
    n7799, n7804, n7809, n7814, n7819, n7824, n7829, n7834, n7839, n7844,
    n7849, n7854, n7859, n7864, n7869, n7874, n7879, n7884, n7889, n7894,
    n7899, n7904, n7909, n7914, n7919, n7924, n7929, n7934, n7939, n7944,
    n7949, n7954, n7959, n7964, n7969, n7974, n7979, n7984, n7989, n7994,
    n7999, n8004, n8009, n8014, n8019, n8024, n8029, n8034, n8039, n8044,
    n8049, n8054, n8059, n8064, n8069, n8074, n8079, n8084, n8089, n8094,
    n8099, n8104, n8109, n8114, n8119, n8124, n8129, n8134, n8139, n8144,
    n8149, n8154, n8159, n8164, n8169, n8174, n8179, n8184, n8189, n8194,
    n8199, n8204, n8209, n8214, n8219, n8224, n8229, n8234, n8239, n8244,
    n8249, n8254, n8259, n8264, n8269, n8274, n8279, n8284, n8289, n8294,
    n8299, n8304, n8309, n8314, n8319, n8324, n8329, n8334, n8339, n8344,
    n8349, n8354, n8359, n8364, n8369, n8374, n8379, n8384, n8389, n8394,
    n8399, n8404, n8409, n8414, n8419, n8424, n8429, n8434, n8439, n8444,
    n8449, n8454, n8459, n8464, n8469, n8474, n8479, n8484, n8489, n8494,
    n8499, n8504, n8509, n8514, n8519, n8524, n8529, n8534, n8539, n8544,
    n8549, n8554, n8559, n8564, n8569, n8574, n8579, n8584, n8589, n8594,
    n8599, n8604, n8609, n8614, n8619, n8624, n8629, n8634, n8639, n8644,
    n8649, n8654, n8659, n8664, n8669, n8674, n8679, n8684, n8689, n8694,
    n8699, n8704, n8709, n8714, n8719, n8724, n8729, n8734, n8739, n8744,
    n8749, n8754, n8759, n8764, n8769, n8774, n8779, n8784, n8789, n8794,
    n8799, n8804, n8809, n8814, n8819, n8824, n8829, n8834, n8839, n8844,
    n8849, n8854, n8859, n8864, n8869, n8874, n8879, n8884, n8889, n8894,
    n8899, n8904, n8909, n8914, n8919, n8924, n8929, n8934, n8939;
  assign \m1_data_o[14]  = ~\new_[25644]_  | ~\new_[25836]_  | ~\new_[3436]_  | ~\new_[25638]_ ;
  assign \m1_data_o[12]  = ~\new_[25600]_  | ~\new_[25862]_  | ~\new_[3439]_  | ~\new_[25864]_ ;
  assign \m1_data_o[9]  = ~\new_[25896]_  | ~\new_[25526]_  | ~\new_[3441]_  | ~\new_[26458]_ ;
  assign \m1_data_o[6]  = ~\new_[25932]_  | ~\new_[25937]_  | ~\new_[3443]_  | ~\new_[24747]_ ;
  assign \m1_data_o[4]  = ~\new_[25979]_  | ~\new_[24708]_  | ~\new_[3446]_  | ~\new_[25289]_ ;
  assign \m1_data_o[2]  = ~\new_[26011]_  | ~\new_[26055]_  | ~\new_[3447]_  | ~\new_[26012]_ ;
  assign \m1_data_o[1]  = ~\new_[26018]_  | ~\new_[25961]_  | ~\new_[3448]_  | ~\new_[24651]_ ;
  assign \m2_data_o[12]  = ~\new_[27107]_  | ~\new_[27109]_  | ~\new_[3467]_  | ~\new_[23133]_ ;
  assign \m2_data_o[11]  = ~\new_[27116]_  | ~\new_[27211]_  | ~\new_[3442]_  | ~\new_[23989]_ ;
  assign \m2_data_o[6]  = ~\new_[27144]_  | ~\new_[27128]_  | ~\new_[3445]_  | ~\new_[24000]_ ;
  assign \m2_data_o[5]  = ~\new_[27179]_  | ~\new_[27927]_  | ~\new_[3454]_  | ~\new_[24055]_ ;
  assign \m2_data_o[2]  = ~\new_[27262]_  | ~\new_[27252]_  | ~\new_[3472]_  | ~\new_[24009]_ ;
  assign \m2_data_o[1]  = ~\new_[27159]_  | ~\new_[27342]_  | ~\new_[3435]_  | ~\new_[24125]_ ;
  assign \m3_data_o[14]  = ~\new_[24540]_  | ~\new_[26656]_  | ~\new_[3462]_  | ~\new_[27260]_ ;
  assign \m3_data_o[12]  = ~\new_[25680]_  | ~\new_[27296]_  | ~\new_[3463]_  | ~\new_[27486]_ ;
  assign \m3_data_o[11]  = ~\new_[25636]_  | ~\new_[27477]_  | ~\new_[3464]_  | ~\new_[27044]_ ;
  assign \m3_data_o[6]  = ~\new_[25768]_  | ~\new_[27157]_  | ~\new_[3470]_  | ~\new_[27121]_ ;
  assign \m3_data_o[5]  = ~\new_[25626]_  | ~\new_[27303]_  | ~\new_[3471]_  | ~\new_[27386]_ ;
  assign \m3_data_o[4]  = ~\new_[25619]_  | ~\new_[27381]_  | ~\new_[3473]_  | ~\new_[27308]_ ;
  assign \m3_data_o[2]  = ~\new_[26090]_  | ~\new_[27238]_  | ~\new_[3417]_  | ~\new_[26997]_ ;
  assign \m3_data_o[1]  = ~\new_[25204]_  | ~\new_[27295]_  | ~\new_[3419]_  | ~\new_[27712]_ ;
  assign \m5_data_o[14]  = ~\new_[25348]_  | ~\new_[25340]_  | ~\new_[3450]_  | ~\new_[23974]_ ;
  assign \m5_data_o[12]  = ~\new_[26475]_  | ~\new_[26221]_  | ~\new_[3451]_  | ~\new_[23961]_ ;
  assign \m5_data_o[9]  = ~\new_[25995]_  | ~\new_[25927]_  | ~\new_[3452]_  | ~\new_[24151]_ ;
  assign \m5_data_o[6]  = ~\new_[26135]_  | ~\new_[25986]_  | ~\new_[3456]_  | ~\new_[23957]_ ;
  assign \m5_data_o[5]  = ~\new_[26102]_  | ~\new_[25275]_  | ~\new_[3440]_  | ~\new_[24519]_ ;
  assign \m5_data_o[4]  = ~\new_[25694]_  | ~\new_[26063]_  | ~\new_[3418]_  | ~\new_[24168]_ ;
  assign \m5_data_o[2]  = ~\new_[25292]_  | ~\new_[26519]_  | ~\new_[3460]_  | ~\new_[24502]_ ;
  assign \m5_data_o[1]  = ~\new_[25287]_  | ~\new_[25297]_  | ~\new_[3437]_  | ~\new_[23964]_ ;
  assign \m6_data_o[12]  = ~\new_[26000]_  | ~\new_[25392]_  | ~\new_[3466]_  | ~\new_[25659]_ ;
  assign \m6_data_o[11]  = ~\new_[25451]_  | ~\new_[25758]_  | ~\new_[3469]_  | ~\new_[25345]_ ;
  assign \m6_data_o[6]  = ~\new_[25454]_  | ~\new_[25367]_  | ~\new_[3455]_  | ~\new_[25585]_ ;
  assign \m6_data_o[5]  = ~\new_[25490]_  | ~\new_[25491]_  | ~\new_[3459]_  | ~\new_[25591]_ ;
  assign \m6_data_o[2]  = ~\new_[25445]_  | ~\new_[25514]_  | ~\new_[3465]_  | ~\new_[25806]_ ;
  assign \m6_data_o[1]  = ~\new_[25517]_  | ~\new_[25125]_  | ~\new_[3468]_  | ~\new_[25519]_ ;
  assign \m7_data_o[14]  = ~\new_[22574]_  | ~\new_[22650]_  | ~\new_[3438]_  | ~\new_[25799]_ ;
  assign \m7_data_o[12]  = ~\new_[22690]_  | ~\new_[22662]_  | ~\new_[3444]_  | ~\new_[26448]_ ;
  assign \m7_data_o[9]  = ~\new_[22623]_  | ~\new_[22617]_  | ~\new_[3449]_  | ~\new_[25647]_ ;
  assign \m7_data_o[6]  = ~\new_[22636]_  | ~\new_[22589]_  | ~\new_[3453]_  | ~\new_[25279]_ ;
  assign \m7_data_o[4]  = ~\new_[22579]_  | ~\new_[22578]_  | ~\new_[3457]_  | ~\new_[25653]_ ;
  assign \m7_data_o[2]  = ~\new_[22620]_  | ~\new_[22647]_  | ~\new_[3458]_  | ~\new_[25776]_ ;
  assign \m7_data_o[1]  = ~\new_[22640]_  | ~\new_[22566]_  | ~\new_[3461]_  | ~\new_[25780]_ ;
  assign \m0_data_o[9]  = ~\new_[21710]_  | ~\new_[24753]_  | ~\new_[3515]_  | ~\new_[25485]_ ;
  assign \m0_data_o[4]  = ~\new_[21767]_  | ~\new_[25874]_  | ~\new_[3528]_  | ~\new_[25863]_ ;
  assign \m0_data_o[2]  = ~\new_[21902]_  | ~\new_[24711]_  | ~\new_[3484]_  | ~\new_[24736]_ ;
  assign \m0_data_o[1]  = ~\new_[21923]_  | ~\new_[24772]_  | ~\new_[3494]_  | ~\new_[26060]_ ;
  assign \m0_data_o[11]  = ~\new_[21780]_  | ~\new_[25579]_  | ~\new_[3506]_  | ~\new_[25718]_ ;
  assign \m0_data_o[6]  = ~\new_[21848]_  | ~\new_[25807]_  | ~\new_[3525]_  | ~\new_[25747]_ ;
  assign \m1_data_o[13]  = ~\new_[25847]_  | ~\new_[25849]_  | ~\new_[3483]_  | ~\new_[25850]_ ;
  assign \m0_data_o[5]  = ~\new_[21868]_  | ~\new_[25673]_  | ~\new_[3526]_  | ~\new_[24728]_ ;
  assign \m1_data_o[10]  = ~\new_[25549]_  | ~\new_[24723]_  | ~\new_[3486]_  | ~\new_[25546]_ ;
  assign \m1_data_o[15]  = ~\new_[26037]_  | ~\new_[25808]_  | ~\new_[3480]_  | ~\new_[25678]_ ;
  assign \m0_data_o[14]  = ~\new_[21669]_  | ~\new_[25709]_  | ~\new_[3523]_  | ~\new_[25377]_ ;
  assign \m1_data_o[7]  = ~\new_[25920]_  | ~\new_[24775]_  | ~\new_[3493]_  | ~\new_[25922]_ ;
  assign \m0_data_o[12]  = ~\new_[21763]_  | ~\new_[25576]_  | ~\new_[3503]_  | ~\new_[25698]_ ;
  assign \m1_data_o[8]  = ~\new_[25305]_  | ~\new_[24865]_  | ~\new_[3490]_  | ~\new_[25910]_ ;
  assign \m1_data_o[3]  = ~\new_[25994]_  | ~\new_[25997]_  | ~\new_[3496]_  | ~\new_[25998]_ ;
  assign \m1_data_o[0]  = ~\new_[25895]_  | ~\new_[25883]_  | ~\new_[3500]_  | ~\new_[24779]_ ;
  assign \m2_data_o[14]  = ~\new_[23205]_  | ~\new_[23981]_  | ~\new_[3520]_  | ~\new_[27293]_ ;
  assign \m2_data_o[13]  = ~\new_[27266]_  | ~\new_[27104]_  | ~\new_[3516]_  | ~\new_[24048]_ ;
  assign \m2_data_o[10]  = ~\new_[27175]_  | ~\new_[26935]_  | ~\new_[3478]_  | ~\new_[24011]_ ;
  assign \m2_data_o[8]  = ~\new_[27865]_  | ~\new_[27164]_  | ~\new_[3518]_  | ~\new_[24049]_ ;
  assign \m2_data_o[3]  = ~\new_[27331]_  | ~\new_[27169]_  | ~\new_[3527]_  | ~\new_[24007]_ ;
  assign \m3_data_o[13]  = ~\new_[25684]_  | ~\new_[27066]_  | ~\new_[3519]_  | ~\new_[27912]_ ;
  assign \m3_data_o[8]  = ~\new_[25981]_  | ~\new_[27245]_  | ~\new_[3524]_  | ~\new_[27047]_ ;
  assign \m3_data_o[10]  = ~\new_[25611]_  | ~\new_[27391]_  | ~\new_[3522]_  | ~\new_[27301]_ ;
  assign \m3_data_o[15]  = ~\new_[25317]_  | ~\new_[27340]_  | ~\new_[3517]_  | ~\new_[27059]_ ;
  assign \m3_data_o[3]  = ~\new_[25559]_  | ~\new_[27457]_  | ~\new_[3530]_  | ~\new_[27456]_ ;
  assign \m3_data_o[0]  = ~\new_[26512]_  | ~\new_[26870]_  | ~\new_[3477]_  | ~\new_[26606]_ ;
  assign \m4_data_o[14]  = ~\new_[21747]_  | ~\new_[24014]_  | ~\new_[3475]_  | ~\new_[26957]_ ;
  assign \m4_data_o[12]  = ~\new_[21887]_  | ~\new_[23525]_  | ~\new_[3479]_  | ~\new_[26938]_ ;
  assign \m4_data_o[9]  = ~\new_[21893]_  | ~\new_[23275]_  | ~\new_[3482]_  | ~\new_[26749]_ ;
  assign \m4_data_o[6]  = ~\new_[21900]_  | ~\new_[25945]_  | ~\new_[3485]_  | ~\new_[23979]_ ;
  assign \m4_data_o[5]  = ~\new_[21901]_  | ~\new_[23971]_  | ~\new_[3488]_  | ~\new_[27412]_ ;
  assign \m4_data_o[4]  = ~\new_[21905]_  | ~\new_[24142]_  | ~\new_[3489]_  | ~\new_[27416]_ ;
  assign \m4_data_o[2]  = ~\new_[21908]_  | ~\new_[24150]_  | ~\new_[3492]_  | ~\new_[27422]_ ;
  assign \m4_data_o[1]  = ~\new_[21911]_  | ~\new_[24154]_  | ~\new_[3495]_  | ~\new_[26773]_ ;
  assign \m5_data_o[15]  = ~\new_[26116]_  | ~\new_[24666]_  | ~\new_[3502]_  | ~\new_[24182]_ ;
  assign \m5_data_o[13]  = ~\new_[25302]_  | ~\new_[26492]_  | ~\new_[3507]_  | ~\new_[23965]_ ;
  assign \m5_data_o[10]  = ~\new_[26137]_  | ~\new_[25946]_  | ~\new_[3509]_  | ~\new_[24185]_ ;
  assign \m4_data_o[11]  = ~\new_[21891]_  | ~\new_[24127]_  | ~\new_[3481]_  | ~\new_[27162]_ ;
  assign \m5_data_o[8]  = ~\new_[24731]_  | ~\new_[26376]_  | ~\new_[3510]_  | ~\new_[23980]_ ;
  assign \m5_data_o[7]  = ~\new_[26343]_  | ~\new_[25726]_  | ~\new_[3511]_  | ~\new_[24385]_ ;
  assign \m5_data_o[3]  = ~\new_[25819]_  | ~\new_[25286]_  | ~\new_[3497]_  | ~\new_[23175]_ ;
  assign \m6_data_o[15]  = ~\new_[25033]_  | ~\new_[25426]_  | ~\new_[3501]_  | ~\new_[25756]_ ;
  assign \m6_data_o[14]  = ~\new_[21711]_  | ~\new_[25481]_  | ~\new_[3529]_  | ~\new_[27126]_ ;
  assign \m5_data_o[0]  = ~\new_[25300]_  | ~\new_[25952]_  | ~\new_[3504]_  | ~\new_[24138]_ ;
  assign \m6_data_o[13]  = ~\new_[25435]_  | ~\new_[25444]_  | ~\new_[3513]_  | ~\new_[25436]_ ;
  assign \m6_data_o[10]  = ~\new_[25118]_  | ~\new_[25461]_  | ~\new_[3476]_  | ~\new_[25462]_ ;
  assign \m6_data_o[8]  = ~\new_[25474]_  | ~\new_[25643]_  | ~\new_[3499]_  | ~\new_[25608]_ ;
  assign \m6_data_o[3]  = ~\new_[25217]_  | ~\new_[25507]_  | ~\new_[3521]_  | ~\new_[25205]_ ;
  assign \m6_data_o[0]  = ~\new_[26084]_  | ~\new_[25186]_  | ~\new_[3474]_  | ~\new_[25686]_ ;
  assign \m7_data_o[15]  = ~\new_[22629]_  | ~\new_[22610]_  | ~\new_[3491]_  | ~\new_[25730]_ ;
  assign \m7_data_o[13]  = ~\new_[22612]_  | ~\new_[23070]_  | ~\new_[3487]_  | ~\new_[24702]_ ;
  assign \m7_data_o[10]  = ~\new_[22616]_  | ~\new_[22622]_  | ~\new_[3498]_  | ~\new_[25603]_ ;
  assign \m7_data_o[8]  = ~\new_[21583]_  | ~\new_[22619]_  | ~\new_[3505]_  | ~\new_[25615]_ ;
  assign \m7_data_o[7]  = ~\new_[22664]_  | ~\new_[21586]_  | ~\new_[3508]_  | ~\new_[24671]_ ;
  assign \m7_data_o[3]  = ~\new_[22569]_  | ~\new_[22567]_  | ~\new_[3512]_  | ~\new_[25568]_ ;
  assign \m7_data_o[0]  = ~\new_[22691]_  | ~\new_[21579]_  | ~\new_[3514]_  | ~\new_[25630]_ ;
  assign \new_[3417]_  = ~\new_[26103]_  & ~\new_[3594]_ ;
  assign \new_[3418]_  = ~\new_[25675]_  & ~\new_[3575]_ ;
  assign \new_[3419]_  = ~\new_[24595]_  & ~\new_[3596]_ ;
  assign \m0_data_o[15]  = ~\new_[21681]_  | ~\new_[25667]_  | ~\new_[3585]_  | ~\new_[25745]_ ;
  assign \m0_data_o[13]  = ~\new_[21741]_  | ~\new_[25128]_  | ~\new_[3537]_  | ~\new_[25369]_ ;
  assign \m0_data_o[10]  = ~\new_[21861]_  | ~\new_[25649]_  | ~\new_[3571]_  | ~\new_[25639]_ ;
  assign \m0_data_o[8]  = ~\new_[21865]_  | ~\new_[25704]_  | ~\new_[3584]_  | ~\new_[25277]_ ;
  assign \m0_data_o[7]  = ~\new_[21926]_  | ~\new_[25552]_  | ~\new_[3592]_  | ~\new_[26041]_ ;
  assign \m0_data_o[3]  = ~\new_[21890]_  | ~\new_[25465]_  | ~\new_[3603]_  | ~\new_[25901]_ ;
  assign \m0_data_o[0]  = ~\new_[21930]_  | ~\new_[26043]_  | ~\new_[3558]_  | ~\new_[25646]_ ;
  assign \m2_data_o[15]  = ~\new_[23232]_  | ~\new_[27523]_  | ~\new_[3583]_  | ~\new_[23978]_ ;
  assign \m4_data_o[15]  = ~\new_[21883]_  | ~\new_[24119]_  | ~\new_[3531]_  | ~\new_[27385]_ ;
  assign \m4_data_o[13]  = ~\new_[21885]_  | ~\new_[24122]_  | ~\new_[3536]_  | ~\new_[27100]_ ;
  assign \m4_data_o[8]  = ~\new_[21895]_  | ~\new_[23986]_  | ~\new_[3542]_  | ~\new_[26848]_ ;
  assign \m4_data_o[7]  = ~\new_[21896]_  | ~\new_[24134]_  | ~\new_[3546]_  | ~\new_[26926]_ ;
  assign \m4_data_o[10]  = ~\new_[21722]_  | ~\new_[24128]_  | ~\new_[3540]_  | ~\new_[27142]_ ;
  assign \m4_data_o[3]  = ~\new_[21907]_  | ~\new_[24146]_  | ~\new_[3553]_  | ~\new_[27420]_ ;
  assign \m4_data_o[0]  = ~\new_[21916]_  | ~\new_[24176]_  | ~\new_[3559]_  | ~\new_[26758]_ ;
  assign \new_[3435]_  = ~\new_[32046]_  & ~\new_[25580]_ ;
  assign \new_[3436]_  = ~\new_[25834]_  & ~\new_[3599]_ ;
  assign \new_[3437]_  = ~\new_[25765]_  & ~\new_[3581]_ ;
  assign \new_[3438]_  = ~\new_[25870]_  & ~\new_[3572]_ ;
  assign \new_[3439]_  = ~\new_[25857]_  & ~\new_[3602]_ ;
  assign \new_[3440]_  = ~\new_[32257]_  & ~\new_[25273]_ ;
  assign \new_[3441]_  = ~\new_[24908]_  & ~\new_[3535]_ ;
  assign \new_[3442]_  = ~\new_[3595]_  & ~\new_[25409]_ ;
  assign \new_[3443]_  = ~\new_[25931]_  & ~\new_[3545]_ ;
  assign \new_[3444]_  = ~\new_[25596]_  & ~\new_[3573]_ ;
  assign \new_[3445]_  = ~\new_[3543]_  & ~\new_[25560]_ ;
  assign \new_[3446]_  = ~\new_[25976]_  & ~\new_[3552]_ ;
  assign \new_[3447]_  = ~\new_[26069]_  & ~\new_[3560]_ ;
  assign \new_[3448]_  = ~\new_[24741]_  & ~\new_[3561]_ ;
  assign \new_[3449]_  = ~\new_[25607]_  & ~\new_[3574]_ ;
  assign \new_[3450]_  = ~\new_[26280]_  & ~\new_[3564]_ ;
  assign \new_[3451]_  = ~\new_[26128]_  & ~\new_[3566]_ ;
  assign \new_[3452]_  = ~\new_[26434]_  & ~\new_[3567]_ ;
  assign \new_[3453]_  = ~\new_[25544]_  & ~\new_[3576]_ ;
  assign \new_[3454]_  = ~\new_[3548]_  & ~\new_[25484]_ ;
  assign \new_[3455]_  = ~\new_[3551]_  & ~\new_[25494]_ ;
  assign \new_[3456]_  = ~\new_[26139]_  & ~\new_[3568]_ ;
  assign \new_[3457]_  = ~\new_[25453]_  & ~\new_[3577]_ ;
  assign \new_[3458]_  = ~\new_[25627]_  & ~\new_[3579]_ ;
  assign \new_[3459]_  = ~\new_[3554]_  & ~\new_[25487]_ ;
  assign \new_[3460]_  = ~\new_[26003]_  & ~\new_[3578]_ ;
  assign \new_[3461]_  = ~\new_[25571]_  & ~\new_[3580]_ ;
  assign \new_[3462]_  = ~\new_[32082]_  & ~\new_[25728]_ ;
  assign \new_[3463]_  = ~\new_[3586]_  & ~\new_[25691]_ ;
  assign \new_[3464]_  = ~\new_[3587]_  & ~\new_[25735]_ ;
  assign \new_[3465]_  = ~\new_[25687]_  & ~\new_[3562]_ ;
  assign \new_[3466]_  = ~\new_[3532]_  & ~\new_[25443]_ ;
  assign \new_[3467]_  = ~\new_[3590]_  & ~\new_[24634]_ ;
  assign \new_[3468]_  = ~\new_[24725]_  & ~\new_[3563]_ ;
  assign \new_[3469]_  = ~\new_[3534]_  & ~\new_[26142]_ ;
  assign \new_[3470]_  = ~\new_[3589]_  & ~\new_[25558]_ ;
  assign \new_[3471]_  = ~\new_[3591]_  & ~\new_[25753]_ ;
  assign \new_[3472]_  = ~\new_[24915]_  & ~\new_[3565]_ ;
  assign \new_[3473]_  = ~\new_[32158]_  & ~\new_[25176]_ ;
  assign \new_[3474]_  = ~\new_[32124]_  & ~\new_[26545]_ ;
  assign \new_[3475]_  = ~\new_[3533]_ ;
  assign \new_[3476]_  = ~\new_[3609]_  & ~\new_[25459]_ ;
  assign \new_[3477]_  = ~\new_[25880]_  & ~\new_[3644]_ ;
  assign \new_[3478]_  = ~\new_[3645]_  & ~\new_[25362]_ ;
  assign \new_[3479]_  = ~\new_[3538]_ ;
  assign \new_[3480]_  = ~\new_[26053]_  & ~\new_[3647]_ ;
  assign \new_[3481]_  = ~\new_[3539]_ ;
  assign \new_[3482]_  = ~\new_[3541]_ ;
  assign \new_[3483]_  = ~\new_[25844]_  & ~\new_[3648]_ ;
  assign \new_[3484]_  = ~\new_[3544]_ ;
  assign \new_[3485]_  = ~\new_[3547]_ ;
  assign \new_[3486]_  = ~\new_[25881]_  & ~\new_[3652]_ ;
  assign \new_[3487]_  = ~\new_[25771]_  & ~\new_[3627]_ ;
  assign \new_[3488]_  = ~\new_[3549]_ ;
  assign \new_[3489]_  = ~\new_[3550]_ ;
  assign \new_[3490]_  = ~\new_[25907]_  & ~\new_[3606]_ ;
  assign \new_[3491]_  = ~\new_[25822]_  & ~\new_[3626]_ ;
  assign \new_[3492]_  = ~\new_[3555]_ ;
  assign \new_[3493]_  = ~\new_[25916]_  & ~\new_[3610]_ ;
  assign \new_[3494]_  = ~\new_[3556]_ ;
  assign \new_[3495]_  = ~\new_[3557]_ ;
  assign \new_[3496]_  = ~\new_[32318]_  & ~\new_[25987]_ ;
  assign \new_[3497]_  = ~\new_[3631]_  & ~\new_[26035]_ ;
  assign \new_[3498]_  = ~\new_[25695]_  & ~\new_[3628]_ ;
  assign \new_[3499]_  = ~\new_[3612]_  & ~\new_[24697]_ ;
  assign \new_[3500]_  = ~\new_[24959]_  & ~\new_[3619]_ ;
  assign \new_[3501]_  = ~\new_[25774]_  & ~\new_[3646]_ ;
  assign \new_[3502]_  = ~\new_[25410]_  & ~\new_[3620]_ ;
  assign \new_[3503]_  = ~\new_[3569]_ ;
  assign \new_[3504]_  = ~\new_[25299]_  & ~\new_[3633]_ ;
  assign \new_[3505]_  = ~\new_[24645]_  & ~\new_[3629]_ ;
  assign \new_[3506]_  = ~\new_[3570]_ ;
  assign \new_[3507]_  = ~\new_[26123]_  & ~\new_[3621]_ ;
  assign \new_[3508]_  = ~\new_[25670]_  & ~\new_[3630]_ ;
  assign \new_[3509]_  = ~\new_[26136]_  & ~\new_[3622]_ ;
  assign \new_[3510]_  = ~\new_[25955]_  & ~\new_[3623]_ ;
  assign \new_[3511]_  = ~\new_[26150]_  & ~\new_[3624]_ ;
  assign \new_[3512]_  = ~\new_[32216]_  & ~\new_[26025]_ ;
  assign \new_[3513]_  = ~\new_[25456]_  & ~\new_[3649]_ ;
  assign \new_[3514]_  = ~\new_[25418]_  & ~\new_[3632]_ ;
  assign \new_[3515]_  = ~\new_[3582]_ ;
  assign \new_[3516]_  = ~\new_[25676]_  & ~\new_[3641]_ ;
  assign \new_[3517]_  = ~\new_[25818]_  & ~\new_[3634]_ ;
  assign \new_[3518]_  = ~\new_[3651]_  & ~\new_[24543]_ ;
  assign \new_[3519]_  = ~\new_[25447]_  & ~\new_[3636]_ ;
  assign \new_[3520]_  = ~\new_[3588]_ ;
  assign \new_[3521]_  = ~\new_[3615]_  & ~\new_[26147]_ ;
  assign \new_[3522]_  = ~\new_[3639]_  & ~\new_[25783]_ ;
  assign \new_[3523]_  = ~\new_[3593]_ ;
  assign \new_[3524]_  = ~\new_[3640]_  & ~\new_[25341]_ ;
  assign \new_[3525]_  = ~\new_[3597]_ ;
  assign \new_[3526]_  = ~\new_[3598]_ ;
  assign \new_[3527]_  = ~\new_[3618]_  & ~\new_[24690]_ ;
  assign \new_[3528]_  = ~\new_[3600]_ ;
  assign \new_[3529]_  = ~\new_[3601]_ ;
  assign \new_[3530]_  = ~\new_[3643]_  & ~\new_[26108]_ ;
  assign \new_[3531]_  = ~\new_[3604]_ ;
  assign \new_[3532]_  = ~\new_[27184]_  | ~\new_[25441]_  | ~\new_[3677]_  | ~\new_[25437]_ ;
  assign \new_[3533]_  = ~\new_[24120]_  | ~\new_[24017]_  | ~\new_[3714]_  | ~\new_[25884]_ ;
  assign \new_[3534]_  = ~\new_[27305]_  | ~\new_[25450]_  | ~\new_[3678]_  | ~\new_[25373]_ ;
  assign \new_[3535]_  = ~\new_[25888]_  | ~\new_[25890]_  | ~\new_[3715]_  | ~\new_[25886]_ ;
  assign \new_[3536]_  = ~\new_[3605]_ ;
  assign \new_[3537]_  = ~\new_[3607]_ ;
  assign \new_[3538]_  = ~\new_[24003]_  | ~\new_[25898]_  | ~\new_[3716]_  | ~\new_[24124]_ ;
  assign \new_[3539]_  = ~\new_[23996]_  | ~\new_[26523]_  | ~\new_[3717]_  | ~\new_[23506]_ ;
  assign \new_[3540]_  = ~\new_[3608]_ ;
  assign \new_[3541]_  = ~\new_[24129]_  | ~\new_[25448]_  | ~\new_[3718]_  | ~\new_[23995]_ ;
  assign \new_[3542]_  = ~\new_[3611]_ ;
  assign \new_[3543]_  = ~\new_[25584]_  | ~\new_[26495]_  | ~\new_[3680]_  | ~\new_[27140]_ ;
  assign \new_[3544]_  = ~\new_[23983]_  | ~\new_[25941]_  | ~\new_[3719]_  | ~\new_[25934]_ ;
  assign \new_[3545]_  = ~\new_[25954]_  | ~\new_[24755]_  | ~\new_[3720]_  | ~\new_[24765]_ ;
  assign \new_[3546]_  = ~\new_[3613]_ ;
  assign \new_[3547]_  = ~\new_[24137]_  | ~\new_[25939]_  | ~\new_[3653]_  | ~\new_[24136]_ ;
  assign \new_[3548]_  = ~\new_[25388]_  | ~\new_[25787]_  | ~\new_[3681]_  | ~\new_[27747]_ ;
  assign \new_[3549]_  = ~\new_[24139]_  | ~\new_[25951]_  | ~\new_[3655]_  | ~\new_[23973]_ ;
  assign \new_[3550]_  = ~\new_[24141]_  | ~\new_[25963]_  | ~\new_[3656]_  | ~\new_[24140]_ ;
  assign \new_[3551]_  = ~\new_[27150]_  | ~\new_[25344]_  | ~\new_[3682]_  | ~\new_[25482]_ ;
  assign \new_[3552]_  = ~\new_[25973]_  | ~\new_[25974]_  | ~\new_[3657]_  | ~\new_[25969]_ ;
  assign \new_[3553]_  = ~\new_[3614]_ ;
  assign \new_[3554]_  = ~\new_[27154]_  | ~\new_[25731]_  | ~\new_[3683]_  | ~\new_[25773]_ ;
  assign \new_[3555]_  = ~\new_[23156]_  | ~\new_[25982]_  | ~\new_[3658]_  | ~\new_[24147]_ ;
  assign \new_[3556]_  = ~\new_[24156]_  | ~\new_[26088]_  | ~\new_[3659]_  | ~\new_[25992]_ ;
  assign \new_[3557]_  = ~\new_[23153]_  | ~\new_[25989]_  | ~\new_[3660]_  | ~\new_[24152]_ ;
  assign \new_[3558]_  = ~\new_[3616]_ ;
  assign \new_[3559]_  = ~\new_[3617]_ ;
  assign \new_[3560]_  = ~\new_[26093]_  | ~\new_[24663]_  | ~\new_[3661]_  | ~\new_[26006]_ ;
  assign \new_[3561]_  = ~\new_[24659]_  | ~\new_[26016]_  | ~\new_[3662]_  | ~\new_[24643]_ ;
  assign \new_[3562]_  = ~\new_[27163]_  | ~\new_[26045]_  | ~\new_[3686]_  | ~\new_[25503]_ ;
  assign \new_[3563]_  = ~\new_[27520]_  | ~\new_[25817]_  | ~\new_[3687]_  | ~\new_[25796]_ ;
  assign \new_[3564]_  = ~\new_[25358]_  | ~\new_[25349]_  | ~\new_[3663]_  | ~\new_[25368]_ ;
  assign \new_[3565]_  = ~\new_[25705]_  | ~\new_[25699]_  | ~\new_[3688]_  | ~\new_[27294]_ ;
  assign \new_[3566]_  = ~\new_[25281]_  | ~\new_[26478]_  | ~\new_[3664]_  | ~\new_[25284]_ ;
  assign \new_[3567]_  = ~\new_[25929]_  | ~\new_[26566]_  | ~\new_[3666]_  | ~\new_[24750]_ ;
  assign \new_[3568]_  = ~\new_[25272]_  | ~\new_[26145]_  | ~\new_[3667]_  | ~\new_[25618]_ ;
  assign \new_[3569]_  = ~\new_[24042]_  | ~\new_[24579]_  | ~\new_[3689]_  | ~\new_[24638]_ ;
  assign \new_[3570]_  = ~\new_[24083]_  | ~\new_[25742]_  | ~\new_[3690]_  | ~\new_[25587]_ ;
  assign \new_[3571]_  = ~\new_[3625]_ ;
  assign \new_[3572]_  = ~\new_[24029]_  | ~\new_[27314]_  | ~\new_[3691]_  | ~\new_[22666]_ ;
  assign \new_[3573]_  = ~\new_[23977]_  | ~\new_[27313]_  | ~\new_[3692]_  | ~\new_[22638]_ ;
  assign \new_[3574]_  = ~\new_[24032]_  | ~\new_[27255]_  | ~\new_[3694]_  | ~\new_[22625]_ ;
  assign \new_[3575]_  = ~\new_[25280]_  | ~\new_[24556]_  | ~\new_[3668]_  | ~\new_[25278]_ ;
  assign \new_[3576]_  = ~\new_[24090]_  | ~\new_[27421]_  | ~\new_[3695]_  | ~\new_[22683]_ ;
  assign \new_[3577]_  = ~\new_[24033]_  | ~\new_[27111]_  | ~\new_[3697]_  | ~\new_[22585]_ ;
  assign \new_[3578]_  = ~\new_[26526]_  | ~\new_[25290]_  | ~\new_[3669]_  | ~\new_[24672]_ ;
  assign \new_[3579]_  = ~\new_[24503]_  | ~\new_[27430]_  | ~\new_[3698]_  | ~\new_[22673]_ ;
  assign \new_[3580]_  = ~\new_[24001]_  | ~\new_[27173]_  | ~\new_[3699]_  | ~\new_[22621]_ ;
  assign \new_[3581]_  = ~\new_[25295]_  | ~\new_[25296]_  | ~\new_[3670]_  | ~\new_[25928]_ ;
  assign \new_[3582]_  = ~\new_[23982]_  | ~\new_[26140]_  | ~\new_[3700]_  | ~\new_[25748]_ ;
  assign \new_[3583]_  = ~\new_[3635]_ ;
  assign \new_[3584]_  = ~\new_[3637]_ ;
  assign \new_[3585]_  = ~\new_[3638]_ ;
  assign \new_[3586]_  = ~\new_[27471]_  | ~\new_[25688]_  | ~\new_[3701]_  | ~\new_[27043]_ ;
  assign \new_[3587]_  = ~\new_[27124]_  | ~\new_[26544]_  | ~\new_[3702]_  | ~\new_[27321]_ ;
  assign \new_[3588]_  = ~\new_[27297]_  | ~\new_[26112]_  | ~\new_[3671]_  | ~\new_[26505]_ ;
  assign \new_[3589]_  = ~\new_[27147]_  | ~\new_[25489]_  | ~\new_[3704]_  | ~\new_[27333]_ ;
  assign \new_[3590]_  = ~\new_[25393]_  | ~\new_[25395]_  | ~\new_[3672]_  | ~\new_[27259]_ ;
  assign \new_[3591]_  = ~\new_[27312]_  | ~\new_[25784]_  | ~\new_[3705]_  | ~\new_[27810]_ ;
  assign \new_[3592]_  = ~\new_[3642]_ ;
  assign \new_[3593]_  = ~\new_[24078]_  | ~\new_[25428]_  | ~\new_[3673]_  | ~\new_[25417]_ ;
  assign \new_[3594]_  = ~\new_[27076]_  | ~\new_[26182]_  | ~\new_[3706]_  | ~\new_[27452]_ ;
  assign \new_[3595]_  = ~\new_[25407]_  | ~\new_[25595]_  | ~\new_[3674]_  | ~\new_[27112]_ ;
  assign \new_[3596]_  = ~\new_[27223]_  | ~\new_[24546]_  | ~\new_[3707]_  | ~\new_[27215]_ ;
  assign \new_[3597]_  = ~\new_[24050]_  | ~\new_[26080]_  | ~\new_[3708]_  | ~\new_[25812]_ ;
  assign \new_[3598]_  = ~\new_[24077]_  | ~\new_[25366]_  | ~\new_[3709]_  | ~\new_[25404]_ ;
  assign \new_[3599]_  = ~\new_[25830]_  | ~\new_[25832]_  | ~\new_[3710]_  | ~\new_[25828]_ ;
  assign \new_[3600]_  = ~\new_[24107]_  | ~\new_[25858]_  | ~\new_[3711]_  | ~\new_[25629]_ ;
  assign \new_[3601]_  = ~\new_[25762]_  | ~\new_[25215]_  | ~\new_[3676]_  | ~\new_[27125]_ ;
  assign \new_[3602]_  = ~\new_[25486]_  | ~\new_[25855]_  | ~\new_[3712]_  | ~\new_[25614]_ ;
  assign \new_[3603]_  = ~\new_[3650]_ ;
  assign \new_[3604]_  = ~\new_[24118]_  | ~\new_[25184]_  | ~\new_[3766]_  | ~\new_[24024]_ ;
  assign \new_[3605]_  = ~\new_[24012]_  | ~\new_[25893]_  | ~\new_[3767]_  | ~\new_[24013]_ ;
  assign \new_[3606]_  = ~\new_[25515]_  | ~\new_[25511]_  | ~\new_[3768]_  | ~\new_[25905]_ ;
  assign \new_[3607]_  = ~\new_[24085]_  | ~\new_[25520]_  | ~\new_[3743]_  | ~\new_[26133]_ ;
  assign \new_[3608]_  = ~\new_[23369]_  | ~\new_[25477]_  | ~\new_[3769]_  | ~\new_[23397]_ ;
  assign \new_[3609]_  = ~\new_[27248]_  | ~\new_[25321]_  | ~\new_[3740]_  | ~\new_[24548]_ ;
  assign \new_[3610]_  = ~\new_[24791]_  | ~\new_[25452]_  | ~\new_[3770]_  | ~\new_[24793]_ ;
  assign \new_[3611]_  = ~\new_[23257]_  | ~\new_[25923]_  | ~\new_[3771]_  | ~\new_[24131]_ ;
  assign \new_[3612]_  = ~\new_[27789]_  | ~\new_[26490]_  | ~\new_[3741]_  | ~\new_[25455]_ ;
  assign \new_[3613]_  = ~\new_[24133]_  | ~\new_[26306]_  | ~\new_[3721]_  | ~\new_[24132]_ ;
  assign \new_[3614]_  = ~\new_[24145]_  | ~\new_[24715]_  | ~\new_[3722]_  | ~\new_[24144]_ ;
  assign \new_[3615]_  = ~\new_[27222]_  | ~\new_[26146]_  | ~\new_[3744]_  | ~\new_[25251]_ ;
  assign \new_[3616]_  = ~\new_[24114]_  | ~\new_[25492]_  | ~\new_[3724]_  | ~\new_[24762]_ ;
  assign \new_[3617]_  = ~\new_[24504]_  | ~\new_[26001]_  | ~\new_[3723]_  | ~\new_[23147]_ ;
  assign \new_[3618]_  = ~\new_[25512]_  | ~\new_[26027]_  | ~\new_[3745]_  | ~\new_[26737]_ ;
  assign \new_[3619]_  = ~\new_[26019]_  | ~\new_[25906]_  | ~\new_[3725]_  | ~\new_[24648]_ ;
  assign \new_[3620]_  = ~\new_[25415]_  | ~\new_[26115]_  | ~\new_[3726]_  | ~\new_[25422]_ ;
  assign \new_[3621]_  = ~\new_[26143]_  | ~\new_[26500]_  | ~\new_[3727]_  | ~\new_[26122]_ ;
  assign \new_[3622]_  = ~\new_[26461]_  | ~\new_[25968]_  | ~\new_[3728]_  | ~\new_[24713]_ ;
  assign \new_[3623]_  = ~\new_[26144]_  | ~\new_[25964]_  | ~\new_[3729]_  | ~\new_[25971]_ ;
  assign \new_[3624]_  = ~\new_[26417]_  | ~\new_[25570]_  | ~\new_[3730]_  | ~\new_[26149]_ ;
  assign \new_[3625]_  = ~\new_[23987]_  | ~\new_[25325]_  | ~\new_[3751]_  | ~\new_[25304]_ ;
  assign \new_[3626]_  = ~\new_[24101]_  | ~\new_[27278]_  | ~\new_[3747]_  | ~\new_[22624]_ ;
  assign \new_[3627]_  = ~\new_[24082]_  | ~\new_[27316]_  | ~\new_[3748]_  | ~\new_[22641]_ ;
  assign \new_[3628]_  = ~\new_[24059]_  | ~\new_[27282]_  | ~\new_[3749]_  | ~\new_[22630]_ ;
  assign \new_[3629]_  = ~\new_[24038]_  | ~\new_[27247]_  | ~\new_[3750]_  | ~\new_[21577]_ ;
  assign \new_[3630]_  = ~\new_[24075]_  | ~\new_[27068]_  | ~\new_[3752]_  | ~\new_[22614]_ ;
  assign \new_[3631]_  = ~\new_[25786]_  | ~\new_[25283]_  | ~\new_[3732]_  | ~\new_[25759]_ ;
  assign \new_[3632]_  = ~\new_[24037]_  | ~\new_[27045]_  | ~\new_[3753]_  | ~\new_[22609]_ ;
  assign \new_[3633]_  = ~\new_[25962]_  | ~\new_[25298]_  | ~\new_[3733]_  | ~\new_[25972]_ ;
  assign \new_[3634]_  = ~\new_[27227]_  | ~\new_[25327]_  | ~\new_[32004]_  | ~\new_[27268]_ ;
  assign \new_[3635]_  = ~\new_[27091]_  | ~\new_[25356]_  | ~\new_[3734]_  | ~\new_[26340]_ ;
  assign \new_[3636]_  = ~\new_[27178]_  | ~\new_[25504]_  | ~\new_[3754]_  | ~\new_[27790]_ ;
  assign \new_[3637]_  = ~\new_[24062]_  | ~\new_[26429]_  | ~\new_[3755]_  | ~\new_[25383]_ ;
  assign \new_[3638]_  = ~\new_[23975]_  | ~\new_[25856]_  | ~\new_[3731]_  | ~\new_[25814]_ ;
  assign \new_[3639]_  = ~\new_[27825]_  | ~\new_[24680]_  | ~\new_[3756]_  | ~\new_[26588]_ ;
  assign \new_[3640]_  = ~\new_[27603]_  | ~\new_[25729]_  | ~\new_[3757]_  | ~\new_[27349]_ ;
  assign \new_[3641]_  = ~\new_[24773]_  | ~\new_[25682]_  | ~\new_[3735]_  | ~\new_[27276]_ ;
  assign \new_[3642]_  = ~\new_[24071]_  | ~\new_[26067]_  | ~\new_[3759]_  | ~\new_[25744]_ ;
  assign \new_[3643]_  = ~\new_[27253]_  | ~\new_[25763]_  | ~\new_[3760]_  | ~\new_[26963]_ ;
  assign \new_[3644]_  = ~\new_[27374]_  | ~\new_[25875]_  | ~\new_[3761]_  | ~\new_[27436]_ ;
  assign \new_[3645]_  = ~\new_[25557]_  | ~\new_[25551]_  | ~\new_[3736]_  | ~\new_[27119]_ ;
  assign \new_[3646]_  = ~\new_[27122]_  | ~\new_[25423]_  | ~\new_[3737]_  | ~\new_[25421]_ ;
  assign \new_[3647]_  = ~\new_[25288]_  | ~\new_[25985]_  | ~\new_[3762]_  | ~\new_[24719]_ ;
  assign \new_[3648]_  = ~\new_[25589]_  | ~\new_[25843]_  | ~\new_[3763]_  | ~\new_[25641]_ ;
  assign \new_[3649]_  = ~\new_[27217]_  | ~\new_[25432]_  | ~\new_[32008]_  | ~\new_[25470]_ ;
  assign \new_[3650]_  = ~\new_[24121]_  | ~\new_[25522]_  | ~\new_[3765]_  | ~\new_[25885]_ ;
  assign \new_[3651]_  = ~\new_[25442]_  | ~\new_[26190]_  | ~\new_[3738]_  | ~\new_[27131]_ ;
  assign \new_[3652]_  = ~\new_[24658]_  | ~\new_[24664]_  | ~\new_[3764]_  | ~\new_[25878]_ ;
  assign \new_[3653]_  = (~\new_[3775]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[6] );
  assign \new_[3654]_  = (~\new_[32259]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[5] );
  assign \new_[3655]_  = (~\new_[32259]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[5] );
  assign \new_[3656]_  = (~\new_[32160]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[4] );
  assign \new_[3657]_  = (~\new_[32160]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[4] );
  assign \new_[3658]_  = (~\new_[3776]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[2] );
  assign \new_[3659]_  = (~\new_[32048]_  | ~\new_[26491]_ ) & (~\s13_data_i[1]  | ~\new_[28726]_ );
  assign \new_[3660]_  = (~\new_[32048]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[1] );
  assign \new_[3661]_  = (~\new_[3776]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[2] );
  assign \new_[3662]_  = (~\new_[32048]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[1] );
  assign \new_[3663]_  = (~\new_[32084]_  | ~\new_[32260]_ ) & (~\new_[32267]_  | ~\s13_data_i[14] );
  assign \new_[3664]_  = (~\new_[3772]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[12] );
  assign \new_[3665]_  = (~\new_[3773]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[11] );
  assign \new_[3666]_  = (~\new_[3774]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[9] );
  assign \new_[3667]_  = (~\new_[3775]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[6] );
  assign \new_[3668]_  = (~\new_[32160]_  | ~\new_[32260]_ ) & (~\new_[32267]_  | ~\s13_data_i[4] );
  assign \new_[3669]_  = (~\new_[3776]_  | ~\new_[32260]_ ) & (~\new_[32267]_  | ~\s13_data_i[2] );
  assign \new_[3670]_  = (~\new_[32048]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[1] );
  assign \new_[3671]_  = (~\new_[32084]_  | ~\new_[32049]_ ) & (~\new_[32056]_  | ~\s13_data_i[14] );
  assign \new_[3672]_  = (~\new_[3772]_  | ~\new_[32049]_ ) & (~\new_[32056]_  | ~\s13_data_i[12] );
  assign \new_[3673]_  = (~\new_[32084]_  | ~\new_[26491]_ ) & (~\s13_data_i[14]  | ~\new_[28726]_ );
  assign \new_[3674]_  = (~\new_[3773]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[11] );
  assign \new_[3675]_  = (~\new_[3774]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[9] );
  assign \new_[3676]_  = (~\new_[32084]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[14] );
  assign \new_[3677]_  = (~\new_[3772]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[12] );
  assign \new_[3678]_  = (~\new_[3773]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[11] );
  assign \new_[3679]_  = (~\new_[3774]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[9] );
  assign \new_[3680]_  = (~\new_[3775]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[6] );
  assign \new_[3681]_  = (~\new_[32259]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[5] );
  assign \new_[3682]_  = (~\new_[3775]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[6] );
  assign \new_[3683]_  = (~\new_[32259]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[5] );
  assign \new_[3684]_  = (~\new_[32160]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[4] );
  assign \new_[3685]_  = (~\new_[32160]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[4] );
  assign \new_[3686]_  = (~\new_[3776]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[2] );
  assign \new_[3687]_  = (~\new_[32048]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[1] );
  assign \new_[3688]_  = (~\new_[3776]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[2] );
  assign \new_[3689]_  = (~\new_[3772]_  | ~\new_[29043]_ ) & (~\s13_data_i[12]  | ~\new_[28726]_ );
  assign \new_[3690]_  = (~\new_[3773]_  | ~\new_[26491]_ ) & (~\s13_data_i[11]  | ~\new_[28726]_ );
  assign \new_[3691]_  = (~\new_[32084]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[14] );
  assign \new_[3692]_  = (~\new_[3772]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[12] );
  assign \new_[3693]_  = (~\new_[3773]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[11] );
  assign \new_[3694]_  = (~\new_[3774]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[9] );
  assign \new_[3695]_  = (~\new_[3775]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[6] );
  assign \new_[3696]_  = (~\new_[32259]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[5] );
  assign \new_[3697]_  = (~\new_[32160]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[4] );
  assign \new_[3698]_  = (~\new_[3776]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[2] );
  assign \new_[3699]_  = (~\new_[32048]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[1] );
  assign \new_[3700]_  = (~\new_[3774]_  | ~\new_[29043]_ ) & (~\s13_data_i[9]  | ~\new_[28726]_ );
  assign \new_[3701]_  = (~\new_[3772]_  | ~\new_[32161]_ ) & (~\new_[32168]_  | ~\s13_data_i[12] );
  assign \new_[3702]_  = (~\new_[3773]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[11] );
  assign \new_[3703]_  = (~\new_[3774]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[9] );
  assign \new_[3704]_  = (~\new_[3775]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[6] );
  assign \new_[3705]_  = (~\new_[32259]_  | ~\new_[32161]_ ) & (~\new_[32168]_  | ~\s13_data_i[5] );
  assign \new_[3706]_  = (~\new_[3776]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[2] );
  assign \new_[3707]_  = (~\new_[32048]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[1] );
  assign \new_[3708]_  = (~\new_[3775]_  | ~\new_[29043]_ ) & (~\s13_data_i[6]  | ~\new_[28726]_ );
  assign \new_[3709]_  = (~\new_[32259]_  | ~\new_[26491]_ ) & (~\s13_data_i[5]  | ~\new_[28726]_ );
  assign \new_[3710]_  = (~\new_[32084]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[14] );
  assign \new_[3711]_  = (~\new_[32160]_  | ~\new_[29043]_ ) & (~\s13_data_i[4]  | ~\new_[28726]_ );
  assign \new_[3712]_  = (~\new_[3772]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[12] );
  assign \new_[3713]_  = (~\new_[3773]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[11] );
  assign \new_[3714]_  = (~\new_[32084]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[14] );
  assign \new_[3715]_  = (~\new_[3774]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[9] );
  assign \new_[3716]_  = (~\new_[3772]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[12] );
  assign \new_[3717]_  = (~\new_[3773]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[11] );
  assign \new_[3718]_  = (~\new_[3774]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[9] );
  assign \new_[3719]_  = (~\new_[3776]_  | ~\new_[26491]_ ) & (~\s13_data_i[2]  | ~\new_[28726]_ );
  assign \new_[3720]_  = (~\new_[3775]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[6] );
  assign \new_[3721]_  = (~\new_[3781]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[7] );
  assign \new_[3722]_  = (~\new_[32320]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[3] );
  assign \new_[3723]_  = (~\new_[32126]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[0] );
  assign \new_[3724]_  = (~\new_[32126]_  | ~\new_[29043]_ ) & (~\s13_data_i[0]  | ~\new_[28726]_ );
  assign \new_[3725]_  = (~\new_[32126]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[0] );
  assign \new_[3726]_  = (~\new_[32006]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[15] );
  assign \new_[3727]_  = (~\new_[32010]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[13] );
  assign \new_[3728]_  = (~\new_[3779]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[10] );
  assign \new_[3729]_  = (~\new_[3780]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[8] );
  assign \new_[3730]_  = (~\new_[3781]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[7] );
  assign \new_[3731]_  = (~\new_[32006]_  | ~\new_[26491]_ ) & (~\s13_data_i[15]  | ~\new_[28726]_ );
  assign \new_[3732]_  = (~\new_[32320]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[3] );
  assign \new_[3733]_  = (~\new_[32126]_  | ~\new_[28712]_ ) & (~\new_[32267]_  | ~\s13_data_i[0] );
  assign \new_[3734]_  = (~\new_[32006]_  | ~\new_[32049]_ ) & (~\new_[32056]_  | ~\s13_data_i[15] );
  assign \new_[3735]_  = (~\new_[32010]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[13] );
  assign \new_[3736]_  = (~\new_[3779]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[10] );
  assign \new_[3737]_  = (~\new_[32006]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[15] );
  assign \new_[3738]_  = (~\new_[3780]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[8] );
  assign \new_[3739]_  = (~\new_[3781]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[7] );
  assign \new_[3740]_  = (~\new_[3779]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[10] );
  assign \new_[3741]_  = (~\new_[3780]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[8] );
  assign \new_[3742]_  = (~\new_[3781]_  | ~\new_[32127]_ ) & (~\new_[32134]_  | ~\s13_data_i[7] );
  assign \new_[3743]_  = (~\new_[32010]_  | ~\new_[29043]_ ) & (~\s13_data_i[13]  | ~\new_[28726]_ );
  assign \new_[3744]_  = (~\new_[32320]_  | ~\new_[24630]_ ) & (~\new_[32134]_  | ~\s13_data_i[3] );
  assign \new_[3745]_  = (~\new_[32320]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[3] );
  assign \new_[3746]_  = (~\new_[32126]_  | ~\new_[24571]_ ) & (~\new_[32056]_  | ~\s13_data_i[0] );
  assign \new_[3747]_  = (~\new_[32006]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[15] );
  assign \new_[3748]_  = (~\new_[32010]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[13] );
  assign \new_[3749]_  = (~\new_[3779]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[10] );
  assign \new_[3750]_  = (~\new_[3780]_  | ~\new_[32343]_ ) & (~\new_[32338]_  | ~\s13_data_i[8] );
  assign \new_[3751]_  = (~\new_[3779]_  | ~\new_[29043]_ ) & (~\s13_data_i[10]  | ~\new_[28726]_ );
  assign \new_[3752]_  = (~\new_[3781]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[7] );
  assign \new_[3753]_  = (~\new_[32126]_  | ~\new_[26525]_ ) & (~\new_[32338]_  | ~\s13_data_i[0] );
  assign \new_[3754]_  = (~\new_[32010]_  | ~\new_[32161]_ ) & (~\new_[32168]_  | ~\s13_data_i[13] );
  assign \new_[3755]_  = (~\new_[3780]_  | ~\new_[29043]_ ) & (~\s13_data_i[8]  | ~\new_[28726]_ );
  assign \new_[3756]_  = (~\new_[3779]_  | ~\new_[32161]_ ) & (~\new_[32168]_  | ~\s13_data_i[10] );
  assign \new_[3757]_  = (~\new_[3780]_  | ~\new_[32161]_ ) & (~\new_[32168]_  | ~\s13_data_i[8] );
  assign \new_[3758]_  = (~\new_[3781]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[7] );
  assign \new_[3759]_  = (~\new_[3781]_  | ~\new_[26491]_ ) & (~\s13_data_i[7]  | ~\new_[28726]_ );
  assign \new_[3760]_  = (~\new_[32320]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[3] );
  assign \new_[3761]_  = (~\new_[32126]_  | ~\new_[26641]_ ) & (~\new_[32168]_  | ~\s13_data_i[0] );
  assign \new_[3762]_  = (~\new_[32006]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[15] );
  assign \new_[3763]_  = (~\new_[32010]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[13] );
  assign \new_[3764]_  = (~\new_[3779]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[10] );
  assign \new_[3765]_  = (~\new_[32320]_  | ~\new_[29043]_ ) & (~\s13_data_i[3]  | ~\new_[28726]_ );
  assign \new_[3766]_  = (~\new_[32006]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[15] );
  assign \new_[3767]_  = (~\new_[32010]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[13] );
  assign \new_[3768]_  = (~\new_[3780]_  | ~\new_[32321]_ ) & (~\new_[32327]_  | ~\s13_data_i[8] );
  assign \new_[3769]_  = (~\new_[3779]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[10] );
  assign \new_[3770]_  = (~\new_[3781]_  | ~\new_[28695]_ ) & (~\new_[32327]_  | ~\s13_data_i[7] );
  assign \new_[3771]_  = (~\new_[3780]_  | ~\new_[27781]_ ) & (~\new_[28851]_  | ~\s13_data_i[8] );
  assign \new_[3772]_  = \new_[3805]_  ? \new_[5881]_  : \s15_data_i[12] ;
  assign \new_[3773]_  = \new_[3806]_  ? \new_[5882]_  : \s15_data_i[11] ;
  assign \new_[3774]_  = \new_[3807]_  ? \new_[5883]_  : \s15_data_i[9] ;
  assign \new_[3775]_  = \new_[3808]_  ? \new_[5881]_  : \s15_data_i[6] ;
  assign \new_[3776]_  = \new_[3811]_  ? \new_[32340]_  : \s15_data_i[2] ;
  assign m6_ack_o = \new_[8521]_  | \new_[3802]_ ;
  assign m7_ack_o = \new_[8535]_  | \new_[3803]_ ;
  assign \new_[3779]_  = \new_[3821]_  ? \new_[5881]_  : \s15_data_i[10] ;
  assign \new_[3780]_  = \new_[3822]_  ? \new_[5881]_  : \s15_data_i[8] ;
  assign \new_[3781]_  = \new_[3823]_  ? \new_[5883]_  : \s15_data_i[7] ;
  assign m0_ack_o = \new_[11004]_  | \new_[3813]_ ;
  assign m1_ack_o = \new_[12907]_  | \new_[3818]_ ;
  assign m2_ack_o = \new_[8524]_  | \new_[3815]_ ;
  assign m3_ack_o = \new_[9449]_  | \new_[3816]_ ;
  assign m4_ack_o = \new_[8545]_  | \new_[3817]_ ;
  assign m5_ack_o = \new_[8514]_  | \new_[3814]_ ;
  assign m1_err_o = \new_[11001]_  | \new_[3837]_ ;
  assign m1_rty_o = \new_[12910]_  | \new_[3838]_ ;
  assign m2_err_o = \new_[8003]_  | \new_[3831]_ ;
  assign m2_rty_o = \new_[8525]_  | \new_[3832]_ ;
  assign m3_err_o = \new_[9450]_  | \new_[3835]_ ;
  assign m3_rty_o = \new_[9453]_  | \new_[3836]_ ;
  assign m4_err_o = \new_[8546]_  | \new_[31943]_ ;
  assign m4_rty_o = \new_[9460]_  | \new_[31955]_ ;
  assign m5_err_o = \new_[8518]_  | \new_[31966]_ ;
  assign m5_rty_o = \new_[9413]_  | \new_[3828]_ ;
  assign m6_err_o = \new_[8000]_  | \new_[3829]_ ;
  assign m6_rty_o = \new_[8523]_  | \new_[3830]_ ;
  assign m7_err_o = \new_[9439]_  | \new_[3833]_ ;
  assign m7_rty_o = \new_[7306]_  | \new_[3834]_ ;
  assign \new_[3802]_  = ~\new_[16053]_  | ~\new_[14637]_  | ~\new_[11082]_  | ~\new_[3848]_ ;
  assign \new_[3803]_  = ~\new_[14786]_  | ~\new_[16169]_  | ~\new_[11087]_  | ~\new_[3849]_ ;
  assign \new_[3804]_  = \\rf_rf_dout_reg[14] ;
  assign \new_[3805]_  = \\rf_rf_dout_reg[12] ;
  assign \new_[3806]_  = \\rf_rf_dout_reg[11] ;
  assign \new_[3807]_  = \\rf_rf_dout_reg[9] ;
  assign \new_[3808]_  = \\rf_rf_dout_reg[6] ;
  assign \new_[3809]_  = \\rf_rf_dout_reg[5] ;
  assign \new_[3810]_  = \\rf_rf_dout_reg[4] ;
  assign \new_[3811]_  = \\rf_rf_dout_reg[2] ;
  assign \new_[3812]_  = \\rf_rf_dout_reg[1] ;
  assign \new_[3813]_  = ~\new_[17041]_  | ~\new_[16159]_  | ~\new_[14369]_  | ~\new_[3865]_ ;
  assign \new_[3814]_  = ~\new_[14749]_  | ~\new_[13353]_  | ~\new_[12954]_  | ~\new_[3864]_ ;
  assign \new_[3815]_  = ~\new_[9728]_  | ~\new_[16062]_  | ~\new_[12984]_  | ~\new_[3866]_ ;
  assign \new_[3816]_  = ~\new_[13396]_  | ~\new_[17076]_  | ~\new_[13029]_  | ~\new_[3867]_ ;
  assign \new_[3817]_  = ~\new_[16115]_  | ~\new_[13315]_  | ~\new_[13026]_  | ~\new_[3868]_ ;
  assign \new_[3818]_  = ~\new_[17082]_  | ~\new_[17083]_  | ~\new_[14434]_  | ~\new_[3869]_ ;
  assign \new_[3819]_  = \\rf_rf_dout_reg[15] ;
  assign \new_[3820]_  = \\rf_rf_dout_reg[13] ;
  assign \new_[3821]_  = \\rf_rf_dout_reg[10] ;
  assign \new_[3822]_  = \\rf_rf_dout_reg[8] ;
  assign \new_[3823]_  = \\rf_rf_dout_reg[7] ;
  assign \new_[3824]_  = \\rf_rf_dout_reg[3] ;
  assign \new_[3825]_  = \\rf_rf_dout_reg[0] ;
  assign m0_err_o = ~\new_[4186]_  | ~\new_[15664]_  | ~\new_[15661]_  | ~\new_[12868]_ ;
  assign m0_rty_o = ~\new_[4187]_  | ~\new_[15667]_  | ~\new_[15665]_  | ~\new_[12876]_ ;
  assign \new_[3828]_  = ~\new_[13366]_  | ~\new_[14758]_  | ~\new_[4018]_  | ~\new_[14373]_ ;
  assign \new_[3829]_  = ~\new_[13254]_  | ~\new_[16854]_  | ~\new_[4019]_  | ~\new_[14390]_ ;
  assign \new_[3830]_  = ~\new_[13260]_  | ~\new_[16857]_  | ~\new_[4020]_  | ~\new_[11083]_ ;
  assign \new_[3831]_  = ~\new_[9729]_  | ~\new_[16067]_  | ~\new_[4021]_  | ~\new_[11084]_ ;
  assign \new_[3832]_  = ~\new_[9730]_  | ~\new_[16070]_  | ~\new_[4022]_  | ~\new_[11085]_ ;
  assign \new_[3833]_  = ~\new_[9787]_  | ~\new_[11435]_  | ~\new_[4023]_  | ~\new_[11088]_ ;
  assign \new_[3834]_  = ~\new_[16178]_  | ~\new_[16177]_  | ~\new_[4024]_  | ~\new_[11089]_ ;
  assign \new_[3835]_  = ~\new_[16189]_  | ~\new_[14816]_  | ~\new_[4025]_  | ~\new_[14423]_ ;
  assign \new_[3836]_  = ~\new_[16223]_  | ~\new_[14812]_  | ~\new_[4026]_  | ~\new_[14424]_ ;
  assign \new_[3837]_  = ~\new_[17878]_  | ~\new_[16213]_  | ~\new_[4027]_  | ~\new_[15802]_ ;
  assign \new_[3838]_  = ~\new_[17102]_  | ~\new_[17104]_  | ~\new_[4028]_  | ~\new_[14435]_ ;
  assign n5104 = ~\new_[32269]_ ;
  assign n5099 = ~\new_[3852]_ ;
  assign n5094 = ~\new_[3854]_ ;
  assign n5134 = ~\new_[3856]_ ;
  assign n5129 = ~\new_[5629]_  & (~\new_[3903]_  | ~\new_[4688]_ );
  assign n5124 = ~\new_[3858]_ ;
  assign n5119 = ~\new_[3859]_ ;
  assign n5114 = ~\new_[3860]_ ;
  assign n5109 = ~\new_[3863]_ ;
  assign \new_[3848]_  = ~\new_[10947]_  & ~\new_[4030]_ ;
  assign \new_[3849]_  = ~\new_[10965]_  & ~\new_[4029]_ ;
  assign n5169 = ~\new_[5629]_  & (~\new_[4031]_  | ~\new_[4681]_ );
  assign n5149 = ~\new_[5629]_  & (~\new_[4032]_  | ~\new_[4683]_ );
  assign \new_[3852]_  = ~\new_[32275]_  | (~\new_[4033]_  & ~\new_[4684]_ );
  assign n5144 = ~\new_[5629]_  & (~\new_[4034]_  | ~\new_[4388]_ );
  assign \new_[3854]_  = ~\new_[32275]_  | (~\new_[4035]_  & ~\new_[32000]_ );
  assign n5139 = ~\new_[5629]_  & (~\new_[4100]_  | ~\new_[4686]_ );
  assign \new_[3856]_  = ~\new_[32275]_  | (~\new_[4165]_  & ~\new_[4687]_ );
  assign n5164 = ~\new_[3870]_ ;
  assign \new_[3858]_  = ~\new_[32275]_  | (~\new_[4183]_  & ~\new_[4691]_ );
  assign \new_[3859]_  = ~\new_[32275]_  | (~\new_[4184]_  & ~\new_[4692]_ );
  assign \new_[3860]_  = ~\new_[32275]_  | (~\new_[32175]_  & ~\new_[32183]_ );
  assign n5159 = ~\new_[3871]_ ;
  assign n5154 = ~\new_[3872]_ ;
  assign \new_[3863]_  = ~\new_[32275]_  | (~\new_[4185]_  & ~\new_[4695]_ );
  assign \new_[3864]_  = ~\new_[4189]_  & ~\new_[10930]_ ;
  assign \new_[3865]_  = ~\new_[4188]_  & ~\new_[10942]_ ;
  assign \new_[3866]_  = ~\new_[4190]_  & ~\new_[12862]_ ;
  assign \new_[3867]_  = ~\new_[4191]_  & ~\new_[12894]_ ;
  assign \new_[3868]_  = ~\new_[4192]_  & ~\new_[9459]_ ;
  assign \new_[3869]_  = ~\new_[4193]_  & ~\new_[10999]_ ;
  assign \new_[3870]_  = ~\new_[32275]_  | (~\new_[4281]_  & ~\new_[4689]_ );
  assign \new_[3871]_  = ~\new_[32275]_  | (~\new_[4282]_  & ~\new_[4847]_ );
  assign \new_[3872]_  = ~\new_[32275]_  | (~\new_[4283]_  & ~\new_[4694]_ );
  assign \new_[3873]_  = \\rf_conf15_reg[0] ;
  assign \new_[3874]_  = \\rf_conf15_reg[10] ;
  assign \new_[3875]_  = \\rf_conf15_reg[11] ;
  assign \new_[3876]_  = \\rf_conf15_reg[12] ;
  assign \new_[3877]_  = \\rf_conf15_reg[13] ;
  assign \new_[3878]_  = \\rf_conf15_reg[14] ;
  assign \new_[3879]_  = \\rf_conf15_reg[15] ;
  assign \new_[3880]_  = \\rf_conf15_reg[1] ;
  assign \new_[3881]_  = \\rf_conf15_reg[2] ;
  assign \new_[3882]_  = \\rf_conf15_reg[3] ;
  assign \new_[3883]_  = \\rf_conf15_reg[4] ;
  assign \new_[3884]_  = \\rf_conf15_reg[5] ;
  assign \new_[3885]_  = \\rf_conf15_reg[6] ;
  assign \new_[3886]_  = \\rf_conf15_reg[7] ;
  assign \new_[3887]_  = \\rf_conf15_reg[8] ;
  assign \new_[3888]_  = \\rf_conf15_reg[9] ;
  assign \m0_data_o[31]  = ~\new_[21778]_  | ~\new_[25648]_  | ~\new_[4380]_  | ~\new_[25917]_ ;
  assign \m0_data_o[30]  = ~\new_[21942]_  | ~\new_[25390]_  | ~\new_[4364]_  | ~\new_[25531]_ ;
  assign \m0_data_o[29]  = ~\new_[21888]_  | ~\new_[25938]_  | ~\new_[4384]_  | ~\new_[25561]_ ;
  assign \m0_data_o[28]  = ~\new_[22661]_  | ~\new_[26098]_  | ~\new_[4407]_  | ~\new_[26047]_ ;
  assign \m0_data_o[26]  = ~\new_[21718]_  | ~\new_[25471]_  | ~\new_[4308]_  | ~\new_[25547]_ ;
  assign \m0_data_o[25]  = ~\new_[21754]_  | ~\new_[25567]_  | ~\new_[4328]_  | ~\new_[25766]_ ;
  assign \m0_data_o[24]  = ~\new_[21684]_  | ~\new_[25732]_  | ~\new_[4347]_  | ~\new_[25495]_ ;
  assign \m0_data_o[23]  = ~\new_[21814]_  | ~\new_[25661]_  | ~\new_[4366]_  | ~\new_[25291]_ ;
  assign \m0_data_o[22]  = ~\new_[21931]_  | ~\new_[25622]_  | ~\new_[4372]_  | ~\new_[26058]_ ;
  assign \m0_data_o[21]  = ~\new_[21873]_  | ~\new_[25852]_  | ~\new_[4387]_  | ~\new_[25825]_ ;
  assign \m0_data_o[20]  = ~\new_[21892]_  | ~\new_[24769]_  | ~\new_[4403]_  | ~\new_[25002]_ ;
  assign \m0_data_o[19]  = ~\new_[21922]_  | ~\new_[25900]_  | ~\new_[4406]_  | ~\new_[26009]_ ;
  assign \m0_data_o[18]  = ~\new_[21949]_  | ~\new_[25634]_  | ~\new_[4408]_  | ~\new_[26527]_ ;
  assign \m0_data_o[17]  = ~\new_[21910]_  | ~\new_[26425]_  | ~\new_[4426]_  | ~\new_[26124]_ ;
  assign \new_[3903]_  = ~\new_[4182]_ ;
  assign \m0_data_o[16]  = ~\new_[21647]_  | ~\new_[24847]_  | ~\new_[4196]_  | ~\new_[25294]_ ;
  assign \m0_data_o[27]  = ~\new_[21646]_  | ~\new_[25319]_  | ~\new_[4425]_  | ~\new_[25840]_ ;
  assign \m1_data_o[31]  = ~\new_[21869]_  | ~\new_[25752]_  | ~\new_[4358]_  | ~\new_[27645]_ ;
  assign \m1_data_o[30]  = ~\new_[21799]_  | ~\new_[25318]_  | ~\new_[4363]_  | ~\new_[26791]_ ;
  assign \m1_data_o[29]  = ~\new_[21805]_  | ~\new_[25538]_  | ~\new_[4368]_  | ~\new_[27279]_ ;
  assign \m1_data_o[28]  = ~\new_[21726]_  | ~\new_[26049]_  | ~\new_[4369]_  | ~\new_[26605]_ ;
  assign \m1_data_o[27]  = ~\new_[21665]_  | ~\new_[26483]_  | ~\new_[4370]_  | ~\new_[27872]_ ;
  assign \m1_data_o[26]  = ~\new_[21702]_  | ~\new_[25809]_  | ~\new_[4371]_  | ~\new_[27049]_ ;
  assign \m1_data_o[25]  = ~\new_[21818]_  | ~\new_[26056]_  | ~\new_[4373]_  | ~\new_[27433]_ ;
  assign \m1_data_o[24]  = ~\new_[21842]_  | ~\new_[26472]_  | ~\new_[4374]_  | ~\new_[27065]_ ;
  assign \m1_data_o[23]  = ~\new_[21863]_  | ~\new_[25586]_  | ~\new_[4375]_  | ~\new_[27432]_ ;
  assign \m1_data_o[22]  = ~\new_[21954]_  | ~\new_[26207]_  | ~\new_[4376]_  | ~\new_[26584]_ ;
  assign \m1_data_o[21]  = ~\new_[21947]_  | ~\new_[26020]_  | ~\new_[4377]_  | ~\new_[27443]_ ;
  assign \m1_data_o[20]  = ~\new_[21853]_  | ~\new_[25772]_  | ~\new_[4378]_  | ~\new_[27435]_ ;
  assign \m1_data_o[17]  = ~\new_[21832]_  | ~\new_[25837]_  | ~\new_[4389]_  | ~\new_[27351]_ ;
  assign \m1_data_o[19]  = ~\new_[21755]_  | ~\new_[24575]_  | ~\new_[4381]_  | ~\new_[27250]_ ;
  assign \m1_data_o[18]  = ~\new_[21849]_  | ~\new_[25815]_  | ~\new_[4385]_  | ~\new_[27344]_ ;
  assign \m1_data_o[16]  = ~\new_[21859]_  | ~\new_[25940]_  | ~\new_[4392]_  | ~\new_[26854]_ ;
  assign \m2_data_o[31]  = ~\new_[23216]_  | ~\new_[24175]_  | ~\new_[4421]_  | ~\new_[27226]_ ;
  assign \m2_data_o[29]  = ~\new_[23259]_  | ~\new_[24181]_  | ~\new_[4429]_  | ~\new_[27221]_ ;
  assign \m2_data_o[28]  = ~\new_[23260]_  | ~\new_[24183]_  | ~\new_[4432]_  | ~\new_[27468]_ ;
  assign \m2_data_o[27]  = ~\new_[23188]_  | ~\new_[24488]_  | ~\new_[4433]_  | ~\new_[27475]_ ;
  assign \m2_data_o[26]  = ~\new_[23263]_  | ~\new_[24285]_  | ~\new_[4434]_  | ~\new_[27785]_ ;
  assign \m2_data_o[25]  = ~\new_[23264]_  | ~\new_[24188]_  | ~\new_[4194]_  | ~\new_[26691]_ ;
  assign \m2_data_o[24]  = ~\new_[23191]_  | ~\new_[23958]_  | ~\new_[4195]_  | ~\new_[27478]_ ;
  assign \m2_data_o[23]  = ~\new_[23193]_  | ~\new_[23116]_  | ~\new_[4303]_  | ~\new_[26646]_ ;
  assign \m2_data_o[22]  = ~\new_[24530]_  | ~\new_[23963]_  | ~\new_[4304]_  | ~\new_[27052]_ ;
  assign \m2_data_o[21]  = ~\new_[23196]_  | ~\new_[23966]_  | ~\new_[4305]_  | ~\new_[27413]_ ;
  assign \m2_data_o[20]  = ~\new_[23197]_  | ~\new_[23994]_  | ~\new_[4306]_  | ~\new_[27399]_ ;
  assign \m2_data_o[18]  = ~\new_[23199]_  | ~\new_[24041]_  | ~\new_[4309]_  | ~\new_[27069]_ ;
  assign \m2_data_o[19]  = ~\new_[24522]_  | ~\new_[23960]_  | ~\new_[4307]_  | ~\new_[27186]_ ;
  assign \m2_data_o[17]  = ~\new_[23240]_  | ~\new_[24463]_  | ~\new_[4311]_  | ~\new_[27075]_ ;
  assign \m2_data_o[16]  = ~\new_[23201]_  | ~\new_[27089]_  | ~\new_[4314]_  | ~\new_[23976]_ ;
  assign \m2_data_o[30]  = ~\new_[23242]_  | ~\new_[24178]_  | ~\new_[4427]_  | ~\new_[26808]_ ;
  assign \m3_data_o[31]  = ~\new_[21765]_  | ~\new_[27202]_  | ~\new_[4341]_  | ~\new_[26787]_ ;
  assign \m3_data_o[30]  = ~\new_[21770]_  | ~\new_[27209]_  | ~\new_[4346]_  | ~\new_[27207]_ ;
  assign \m3_data_o[29]  = ~\new_[21866]_  | ~\new_[26796]_  | ~\new_[4350]_  | ~\new_[27361]_ ;
  assign \m3_data_o[28]  = ~\new_[21773]_  | ~\new_[27318]_  | ~\new_[4351]_  | ~\new_[27345]_ ;
  assign \m3_data_o[27]  = ~\new_[21776]_  | ~\new_[27287]_  | ~\new_[4352]_  | ~\new_[27800]_ ;
  assign \m3_data_o[26]  = ~\new_[21800]_  | ~\new_[27256]_  | ~\new_[4353]_  | ~\new_[27283]_ ;
  assign \m3_data_o[25]  = ~\new_[21783]_  | ~\new_[27239]_  | ~\new_[4354]_  | ~\new_[26778]_ ;
  assign \m3_data_o[24]  = ~\new_[21786]_  | ~\new_[27243]_  | ~\new_[4355]_  | ~\new_[27168]_ ;
  assign \m3_data_o[23]  = ~\new_[21788]_  | ~\new_[27387]_  | ~\new_[4356]_  | ~\new_[27300]_ ;
  assign \m3_data_o[22]  = ~\new_[21790]_  | ~\new_[27446]_  | ~\new_[4357]_  | ~\new_[27236]_ ;
  assign \m3_data_o[18]  = ~\new_[21756]_  | ~\new_[27411]_  | ~\new_[4362]_  | ~\new_[27598]_ ;
  assign \m3_data_o[17]  = ~\new_[21809]_  | ~\new_[27064]_  | ~\new_[4365]_  | ~\new_[27118]_ ;
  assign \m3_data_o[16]  = ~\new_[21803]_  | ~\new_[27327]_  | ~\new_[4367]_  | ~\new_[27263]_ ;
  assign \m3_data_o[19]  = ~\new_[21796]_  | ~\new_[27257]_  | ~\new_[4361]_  | ~\new_[27607]_ ;
  assign \m3_data_o[20]  = ~\new_[21877]_  | ~\new_[27357]_  | ~\new_[4360]_  | ~\new_[27390]_ ;
  assign \m3_data_o[21]  = ~\new_[21819]_  | ~\new_[27332]_  | ~\new_[4359]_  | ~\new_[27453]_ ;
  assign \m4_data_o[31]  = ~\new_[21839]_  | ~\new_[24158]_  | ~\new_[4383]_  | ~\new_[27428]_ ;
  assign \m4_data_o[30]  = ~\new_[21851]_  | ~\new_[24058]_  | ~\new_[4386]_  | ~\new_[26792]_ ;
  assign \m4_data_o[29]  = ~\new_[21856]_  | ~\new_[23990]_  | ~\new_[4390]_  | ~\new_[27077]_ ;
  assign \m4_data_o[28]  = ~\new_[21927]_  | ~\new_[24010]_  | ~\new_[4391]_  | ~\new_[26872]_ ;
  assign \m4_data_o[27]  = ~\new_[21860]_  | ~\new_[24070]_  | ~\new_[4393]_  | ~\new_[27350]_ ;
  assign \m4_data_o[26]  = ~\new_[21862]_  | ~\new_[23972]_  | ~\new_[4394]_  | ~\new_[26830]_ ;
  assign \m4_data_o[25]  = ~\new_[21903]_  | ~\new_[24084]_  | ~\new_[4395]_  | ~\new_[27149]_ ;
  assign \m4_data_o[24]  = ~\new_[21870]_  | ~\new_[24051]_  | ~\new_[4396]_  | ~\new_[27269]_ ;
  assign \m4_data_o[23]  = ~\new_[22675]_  | ~\new_[24047]_  | ~\new_[4397]_  | ~\new_[27362]_ ;
  assign \m4_data_o[21]  = ~\new_[21791]_  | ~\new_[24104]_  | ~\new_[4399]_  | ~\new_[27370]_ ;
  assign \m4_data_o[20]  = ~\new_[22582]_  | ~\new_[23143]_  | ~\new_[4400]_  | ~\new_[27171]_ ;
  assign \m4_data_o[19]  = ~\new_[21876]_  | ~\new_[23991]_  | ~\new_[4401]_  | ~\new_[26772]_ ;
  assign \m4_data_o[18]  = ~\new_[21772]_  | ~\new_[24115]_  | ~\new_[4402]_  | ~\new_[27376]_ ;
  assign \m4_data_o[17]  = ~\new_[21878]_  | ~\new_[23953]_  | ~\new_[4404]_  | ~\new_[27380]_ ;
  assign \m4_data_o[16]  = ~\new_[21880]_  | ~\new_[24025]_  | ~\new_[4405]_  | ~\new_[27192]_ ;
  assign \m4_data_o[22]  = ~\new_[21874]_  | ~\new_[24098]_  | ~\new_[4398]_  | ~\new_[27366]_ ;
  assign \m5_data_o[31]  = ~\new_[21875]_  | ~\new_[24161]_  | ~\new_[4409]_  | ~\new_[27434]_ ;
  assign \m5_data_o[30]  = ~\new_[22344]_  | ~\new_[24057]_  | ~\new_[4410]_  | ~\new_[27358]_ ;
  assign \m5_data_o[29]  = ~\new_[21857]_  | ~\new_[24163]_  | ~\new_[4411]_  | ~\new_[27346]_ ;
  assign \m5_data_o[28]  = ~\new_[21935]_  | ~\new_[24165]_  | ~\new_[4412]_  | ~\new_[27328]_ ;
  assign \m5_data_o[27]  = ~\new_[21938]_  | ~\new_[24073]_  | ~\new_[4413]_  | ~\new_[27317]_ ;
  assign \m5_data_o[26]  = ~\new_[21940]_  | ~\new_[24069]_  | ~\new_[4415]_  | ~\new_[27440]_ ;
  assign \m5_data_o[25]  = ~\new_[21943]_  | ~\new_[24169]_  | ~\new_[4416]_  | ~\new_[27292]_ ;
  assign \m5_data_o[24]  = ~\new_[21948]_  | ~\new_[24056]_  | ~\new_[4417]_  | ~\new_[27275]_ ;
  assign \m5_data_o[21]  = ~\new_[21957]_  | ~\new_[24173]_  | ~\new_[4422]_  | ~\new_[27454]_ ;
  assign \m5_data_o[20]  = ~\new_[21960]_  | ~\new_[24174]_  | ~\new_[4423]_  | ~\new_[27455]_ ;
  assign \m5_data_o[19]  = ~\new_[21758]_  | ~\new_[24177]_  | ~\new_[4424]_  | ~\new_[27963]_ ;
  assign \m5_data_o[18]  = ~\new_[21965]_  | ~\new_[24518]_  | ~\new_[4428]_  | ~\new_[27936]_ ;
  assign \m5_data_o[16]  = ~\new_[21971]_  | ~\new_[24180]_  | ~\new_[4431]_  | ~\new_[27138]_ ;
  assign \m5_data_o[23]  = ~\new_[21951]_  | ~\new_[24045]_  | ~\new_[4419]_  | ~\new_[27445]_ ;
  assign \m5_data_o[17]  = ~\new_[21966]_  | ~\new_[24179]_  | ~\new_[4430]_  | ~\new_[27166]_ ;
  assign \m5_data_o[22]  = ~\new_[21955]_  | ~\new_[24086]_  | ~\new_[4420]_  | ~\new_[27450]_ ;
  assign \m6_data_o[31]  = ~\new_[21658]_  | ~\new_[25835]_  | ~\new_[4310]_  | ~\new_[27070]_ ;
  assign \m6_data_o[30]  = ~\new_[21661]_  | ~\new_[25702]_  | ~\new_[4312]_  | ~\new_[27074]_ ;
  assign \m6_data_o[29]  = ~\new_[21664]_  | ~\new_[25737]_  | ~\new_[4313]_  | ~\new_[27079]_ ;
  assign \m6_data_o[28]  = ~\new_[21668]_  | ~\new_[25782]_  | ~\new_[4315]_  | ~\new_[27330]_ ;
  assign \m6_data_o[27]  = ~\new_[21673]_  | ~\new_[25757]_  | ~\new_[4316]_  | ~\new_[27087]_ ;
  assign \m6_data_o[26]  = ~\new_[21676]_  | ~\new_[26407]_  | ~\new_[4317]_  | ~\new_[27315]_ ;
  assign \m6_data_o[25]  = ~\new_[21678]_  | ~\new_[25365]_  | ~\new_[4318]_  | ~\new_[27096]_ ;
  assign \m6_data_o[23]  = ~\new_[21682]_  | ~\new_[27280]_  | ~\new_[4320]_  | ~\new_[25703]_ ;
  assign \m6_data_o[22]  = ~\new_[21685]_  | ~\new_[25382]_  | ~\new_[4321]_  | ~\new_[27271]_ ;
  assign \m6_data_o[21]  = ~\new_[21688]_  | ~\new_[25655]_  | ~\new_[4322]_  | ~\new_[27106]_ ;
  assign \m6_data_o[20]  = ~\new_[21691]_  | ~\new_[25398]_  | ~\new_[4323]_  | ~\new_[26810]_ ;
  assign \m6_data_o[19]  = ~\new_[21694]_  | ~\new_[25403]_  | ~\new_[4324]_  | ~\new_[27110]_ ;
  assign \m6_data_o[17]  = ~\new_[21700]_  | ~\new_[24735]_  | ~\new_[4326]_  | ~\new_[27204]_ ;
  assign \m6_data_o[24]  = ~\new_[21680]_  | ~\new_[25713]_  | ~\new_[4319]_  | ~\new_[27299]_ ;
  assign \m6_data_o[16]  = ~\new_[21704]_  | ~\new_[25419]_  | ~\new_[4327]_  | ~\new_[27182]_ ;
  assign \m6_data_o[18]  = ~\new_[21697]_  | ~\new_[25440]_  | ~\new_[4325]_  | ~\new_[26780]_ ;
  assign \m7_data_o[31]  = ~\new_[20063]_  | ~\new_[25537]_  | ~\new_[4329]_  | ~\new_[27397]_ ;
  assign \m7_data_o[30]  = ~\new_[20043]_  | ~\new_[25540]_  | ~\new_[4330]_  | ~\new_[27176]_ ;
  assign \m7_data_o[29]  = ~\new_[20044]_  | ~\new_[25637]_  | ~\new_[4331]_  | ~\new_[27129]_ ;
  assign \m7_data_o[28]  = ~\new_[20094]_  | ~\new_[25740]_  | ~\new_[4332]_  | ~\new_[27183]_ ;
  assign \m7_data_o[27]  = ~\new_[20051]_  | ~\new_[25554]_  | ~\new_[4333]_  | ~\new_[27868]_ ;
  assign \m7_data_o[26]  = ~\new_[20113]_  | ~\new_[25769]_  | ~\new_[4335]_  | ~\new_[27404]_ ;
  assign \m7_data_o[25]  = ~\new_[19992]_  | ~\new_[25516]_  | ~\new_[4336]_  | ~\new_[27244]_ ;
  assign \m7_data_o[23]  = ~\new_[20050]_  | ~\new_[25472]_  | ~\new_[4339]_  | ~\new_[27067]_ ;
  assign \m7_data_o[22]  = ~\new_[20130]_  | ~\new_[25306]_  | ~\new_[4340]_  | ~\new_[27483]_ ;
  assign \m7_data_o[21]  = ~\new_[20055]_  | ~\new_[25572]_  | ~\new_[4342]_  | ~\new_[27448]_ ;
  assign \m7_data_o[20]  = ~\new_[20128]_  | ~\new_[24733]_  | ~\new_[4343]_  | ~\new_[27438]_ ;
  assign \m7_data_o[24]  = ~\new_[20114]_  | ~\new_[25562]_  | ~\new_[4337]_  | ~\new_[27053]_ ;
  assign \m7_data_o[18]  = ~\new_[20056]_  | ~\new_[25510]_  | ~\new_[4345]_  | ~\new_[27203]_ ;
  assign \m7_data_o[19]  = ~\new_[20123]_  | ~\new_[25936]_  | ~\new_[4344]_  | ~\new_[27200]_ ;
  assign \m7_data_o[16]  = ~\new_[20059]_  | ~\new_[25532]_  | ~\new_[4349]_  | ~\new_[27148]_ ;
  assign \m7_data_o[17]  = ~\new_[20058]_  | ~\new_[25581]_  | ~\new_[4348]_  | ~\new_[27185]_ ;
  assign \new_[4018]_  = ~\new_[31978]_  & ~\new_[10937]_ ;
  assign \new_[4019]_  = ~\new_[4301]_  & ~\new_[9418]_ ;
  assign \new_[4020]_  = ~\new_[4302]_  & ~\new_[9421]_ ;
  assign \new_[4021]_  = ~\new_[12863]_  & ~\new_[4334]_ ;
  assign \new_[4022]_  = ~\new_[12865]_  & ~\new_[4338]_ ;
  assign \new_[4023]_  = ~\new_[31986]_  & ~\new_[12886]_ ;
  assign \new_[4024]_  = ~\new_[4300]_  & ~\new_[9442]_ ;
  assign \new_[4025]_  = ~\new_[4379]_  & ~\new_[12896]_ ;
  assign \new_[4026]_  = ~\new_[4382]_  & ~\new_[9454]_ ;
  assign \new_[4027]_  = ~\new_[11005]_  & ~\new_[4414]_ ;
  assign \new_[4028]_  = ~\new_[12912]_  & ~\new_[4418]_ ;
  assign \new_[4029]_  = ~\new_[16152]_  | ~\new_[4846]_  | ~\new_[17068]_  | ~\new_[17050]_ ;
  assign \new_[4030]_  = ~\new_[17709]_  | ~\new_[4845]_  | ~\new_[17708]_  | ~\new_[14636]_ ;
  assign \new_[4031]_  = ~\new_[4197]_ ;
  assign \new_[4032]_  = ~\new_[4198]_ ;
  assign \new_[4033]_  = ~\new_[4740]_  | ~\new_[5557]_  | ~\new_[4888]_ ;
  assign \new_[4034]_  = ~\new_[4199]_ ;
  assign \new_[4035]_  = ~\new_[5564]_  | ~\new_[5565]_  | ~\new_[5566]_  | ~\new_[4742]_ ;
  assign \new_[4036]_  = \\rf_conf0_reg[0] ;
  assign \new_[4037]_  = \\rf_conf0_reg[10] ;
  assign \new_[4038]_  = \\rf_conf0_reg[11] ;
  assign \new_[4039]_  = \\rf_conf0_reg[12] ;
  assign \new_[4040]_  = \\rf_conf0_reg[13] ;
  assign \new_[4041]_  = \\rf_conf0_reg[14] ;
  assign \new_[4042]_  = \\rf_conf0_reg[15] ;
  assign \new_[4043]_  = \\rf_conf0_reg[1] ;
  assign \new_[4044]_  = \\rf_conf0_reg[2] ;
  assign \new_[4045]_  = \\rf_conf0_reg[3] ;
  assign \new_[4046]_  = \\rf_conf0_reg[4] ;
  assign \new_[4047]_  = \\rf_conf0_reg[5] ;
  assign \new_[4048]_  = \\rf_conf0_reg[6] ;
  assign \new_[4049]_  = \\rf_conf0_reg[7] ;
  assign \new_[4050]_  = \\rf_conf0_reg[8] ;
  assign \new_[4051]_  = \\rf_conf0_reg[9] ;
  assign \new_[4052]_  = \\rf_conf12_reg[0] ;
  assign \new_[4053]_  = \\rf_conf12_reg[10] ;
  assign \new_[4054]_  = \\rf_conf12_reg[11] ;
  assign \new_[4055]_  = \\rf_conf12_reg[12] ;
  assign \new_[4056]_  = \\rf_conf12_reg[13] ;
  assign \new_[4057]_  = \\rf_conf12_reg[14] ;
  assign \new_[4058]_  = \\rf_conf12_reg[15] ;
  assign \new_[4059]_  = \\rf_conf12_reg[1] ;
  assign \new_[4060]_  = \\rf_conf12_reg[2] ;
  assign \new_[4061]_  = \\rf_conf12_reg[3] ;
  assign \new_[4062]_  = \\rf_conf12_reg[4] ;
  assign \new_[4063]_  = \\rf_conf12_reg[5] ;
  assign \new_[4064]_  = \\rf_conf12_reg[6] ;
  assign \new_[4065]_  = \\rf_conf12_reg[7] ;
  assign \new_[4066]_  = \\rf_conf12_reg[8] ;
  assign \new_[4067]_  = \\rf_conf12_reg[9] ;
  assign \new_[4068]_  = \\rf_conf13_reg[0] ;
  assign \new_[4069]_  = \\rf_conf13_reg[10] ;
  assign \new_[4070]_  = \\rf_conf13_reg[11] ;
  assign \new_[4071]_  = \\rf_conf13_reg[12] ;
  assign \new_[4072]_  = \\rf_conf13_reg[13] ;
  assign \new_[4073]_  = \\rf_conf13_reg[14] ;
  assign \new_[4074]_  = \\rf_conf13_reg[15] ;
  assign \new_[4075]_  = \\rf_conf13_reg[1] ;
  assign \new_[4076]_  = \\rf_conf13_reg[4] ;
  assign \new_[4077]_  = \\rf_conf13_reg[5] ;
  assign \new_[4078]_  = \\rf_conf13_reg[6] ;
  assign \new_[4079]_  = \\rf_conf13_reg[7] ;
  assign \new_[4080]_  = \\rf_conf13_reg[8] ;
  assign \new_[4081]_  = \\rf_conf13_reg[9] ;
  assign \new_[4082]_  = \\rf_conf14_reg[0] ;
  assign \new_[4083]_  = \\rf_conf14_reg[10] ;
  assign \new_[4084]_  = \\rf_conf14_reg[11] ;
  assign \new_[4085]_  = \\rf_conf14_reg[12] ;
  assign \new_[4086]_  = \\rf_conf14_reg[13] ;
  assign \new_[4087]_  = \\rf_conf14_reg[14] ;
  assign \new_[4088]_  = \\rf_conf14_reg[15] ;
  assign \new_[4089]_  = \\rf_conf14_reg[1] ;
  assign \new_[4090]_  = \\rf_conf14_reg[3] ;
  assign \new_[4091]_  = \\rf_conf14_reg[4] ;
  assign \new_[4092]_  = \\rf_conf14_reg[5] ;
  assign \new_[4093]_  = \\rf_conf14_reg[6] ;
  assign \new_[4094]_  = \\rf_conf14_reg[7] ;
  assign \new_[4095]_  = \\rf_conf14_reg[8] ;
  assign \new_[4096]_  = \\rf_conf14_reg[9] ;
  assign \new_[4097]_  = \\rf_conf13_reg[2] ;
  assign \new_[4098]_  = \\rf_conf13_reg[3] ;
  assign \new_[4099]_  = \\rf_conf14_reg[2] ;
  assign \new_[4100]_  = ~\new_[4232]_ ;
  assign \new_[4101]_  = \\rf_conf1_reg[0] ;
  assign \new_[4102]_  = \\rf_conf1_reg[10] ;
  assign \new_[4103]_  = \\rf_conf1_reg[11] ;
  assign \new_[4104]_  = \\rf_conf1_reg[12] ;
  assign \new_[4105]_  = \\rf_conf1_reg[13] ;
  assign \new_[4106]_  = \\rf_conf1_reg[14] ;
  assign \new_[4107]_  = \\rf_conf1_reg[15] ;
  assign \new_[4108]_  = \\rf_conf1_reg[1] ;
  assign \new_[4109]_  = \\rf_conf1_reg[2] ;
  assign \new_[4110]_  = \\rf_conf1_reg[3] ;
  assign \new_[4111]_  = \\rf_conf1_reg[4] ;
  assign \new_[4112]_  = \\rf_conf1_reg[5] ;
  assign \new_[4113]_  = \\rf_conf1_reg[6] ;
  assign \new_[4114]_  = \\rf_conf1_reg[7] ;
  assign \new_[4115]_  = \\rf_conf1_reg[8] ;
  assign \new_[4116]_  = \\rf_conf1_reg[9] ;
  assign \new_[4117]_  = \\rf_conf2_reg[0] ;
  assign \new_[4118]_  = \\rf_conf2_reg[10] ;
  assign \new_[4119]_  = \\rf_conf2_reg[11] ;
  assign \new_[4120]_  = \\rf_conf2_reg[12] ;
  assign \new_[4121]_  = \\rf_conf2_reg[13] ;
  assign \new_[4122]_  = \\rf_conf2_reg[14] ;
  assign \new_[4123]_  = \\rf_conf2_reg[15] ;
  assign \new_[4124]_  = \\rf_conf2_reg[1] ;
  assign \new_[4125]_  = \\rf_conf2_reg[2] ;
  assign \new_[4126]_  = \\rf_conf2_reg[3] ;
  assign \new_[4127]_  = \\rf_conf2_reg[4] ;
  assign \new_[4128]_  = \\rf_conf2_reg[5] ;
  assign \new_[4129]_  = \\rf_conf2_reg[6] ;
  assign \new_[4130]_  = \\rf_conf2_reg[7] ;
  assign \new_[4131]_  = \\rf_conf2_reg[8] ;
  assign \new_[4132]_  = \\rf_conf2_reg[9] ;
  assign \new_[4133]_  = \\rf_conf3_reg[0] ;
  assign \new_[4134]_  = \\rf_conf3_reg[10] ;
  assign \new_[4135]_  = \\rf_conf3_reg[11] ;
  assign \new_[4136]_  = \\rf_conf3_reg[12] ;
  assign \new_[4137]_  = \\rf_conf3_reg[13] ;
  assign \new_[4138]_  = \\rf_conf3_reg[14] ;
  assign \new_[4139]_  = \\rf_conf3_reg[15] ;
  assign \new_[4140]_  = \\rf_conf3_reg[1] ;
  assign \new_[4141]_  = \\rf_conf3_reg[2] ;
  assign \new_[4142]_  = \\rf_conf3_reg[3] ;
  assign \new_[4143]_  = \\rf_conf3_reg[4] ;
  assign \new_[4144]_  = \\rf_conf3_reg[5] ;
  assign \new_[4145]_  = \\rf_conf3_reg[6] ;
  assign \new_[4146]_  = \\rf_conf3_reg[7] ;
  assign \new_[4147]_  = \\rf_conf3_reg[8] ;
  assign \new_[4148]_  = \\rf_conf3_reg[9] ;
  assign \new_[4149]_  = \\rf_conf5_reg[0] ;
  assign \new_[4150]_  = \\rf_conf5_reg[10] ;
  assign \new_[4151]_  = \\rf_conf5_reg[11] ;
  assign \new_[4152]_  = \\rf_conf5_reg[12] ;
  assign \new_[4153]_  = \\rf_conf5_reg[13] ;
  assign \new_[4154]_  = \\rf_conf5_reg[14] ;
  assign \new_[4155]_  = \\rf_conf5_reg[15] ;
  assign \new_[4156]_  = \\rf_conf5_reg[1] ;
  assign \new_[4157]_  = \\rf_conf5_reg[2] ;
  assign \new_[4158]_  = \\rf_conf5_reg[3] ;
  assign \new_[4159]_  = \\rf_conf5_reg[4] ;
  assign \new_[4160]_  = \\rf_conf5_reg[5] ;
  assign \new_[4161]_  = \\rf_conf5_reg[6] ;
  assign \new_[4162]_  = \\rf_conf5_reg[7] ;
  assign \new_[4163]_  = \\rf_conf5_reg[8] ;
  assign \new_[4164]_  = \\rf_conf5_reg[9] ;
  assign \new_[4165]_  = ~\new_[4743]_  | ~\new_[5572]_  | ~\new_[4894]_ ;
  assign \new_[4166]_  = \\rf_conf7_reg[0] ;
  assign \new_[4167]_  = \\rf_conf7_reg[10] ;
  assign \new_[4168]_  = \\rf_conf7_reg[11] ;
  assign \new_[4169]_  = \\rf_conf7_reg[12] ;
  assign \new_[4170]_  = \\rf_conf7_reg[13] ;
  assign \new_[4171]_  = \\rf_conf7_reg[14] ;
  assign \new_[4172]_  = \\rf_conf7_reg[15] ;
  assign \new_[4173]_  = \\rf_conf7_reg[1] ;
  assign \new_[4174]_  = \\rf_conf7_reg[2] ;
  assign \new_[4175]_  = \\rf_conf7_reg[3] ;
  assign \new_[4176]_  = \\rf_conf7_reg[4] ;
  assign \new_[4177]_  = \\rf_conf7_reg[5] ;
  assign \new_[4178]_  = \\rf_conf7_reg[6] ;
  assign \new_[4179]_  = \\rf_conf7_reg[7] ;
  assign \new_[4180]_  = \\rf_conf7_reg[8] ;
  assign \new_[4181]_  = \\rf_conf7_reg[9] ;
  assign \new_[4182]_  = ~\new_[4895]_  | ~\new_[5577]_  | ~\new_[4744]_ ;
  assign \new_[4183]_  = ~\new_[5584]_  | ~\new_[5438]_  | ~\new_[5669]_  | ~\new_[4745]_ ;
  assign \new_[4184]_  = ~\new_[5588]_  | ~\new_[5441]_  | ~\new_[5670]_  | ~\new_[4746]_ ;
  assign \new_[4185]_  = ~\new_[5604]_  | ~\new_[5448]_  | ~\new_[5605]_  | ~\new_[4747]_ ;
  assign \new_[4186]_  = ~\new_[14333]_  & ~\new_[4649]_ ;
  assign \new_[4187]_  = ~\new_[14336]_  & ~\new_[4652]_ ;
  assign \new_[4188]_  = ~\new_[13368]_  | ~\new_[16150]_  | ~\new_[16144]_  | ~\new_[4844]_ ;
  assign \new_[4189]_  = ~\new_[17015]_  | ~\new_[18652]_  | ~\new_[14746]_  | ~\new_[4848]_ ;
  assign \new_[4190]_  = ~\new_[16861]_  | ~\new_[18560]_  | ~\new_[16059]_  | ~\new_[4849]_ ;
  assign \new_[4191]_  = ~\new_[17059]_  | ~\new_[16187]_  | ~\new_[17043]_  | ~\new_[4850]_ ;
  assign \new_[4192]_  = ~\new_[16950]_  | ~\new_[14709]_  | ~\new_[14707]_  | ~\new_[4851]_ ;
  assign \new_[4193]_  = ~\new_[17079]_  | ~\new_[18665]_  | ~\new_[17078]_  | ~\new_[4852]_ ;
  assign \new_[4194]_  = ~\new_[4435]_ ;
  assign \new_[4195]_  = ~\new_[4436]_ ;
  assign \new_[4196]_  = ~\new_[4437]_ ;
  assign \new_[4197]_  = ~\new_[5421]_  | ~\new_[5420]_  | ~\new_[5422]_  | ~\new_[4883]_ ;
  assign \new_[4198]_  = ~\new_[4885]_  | ~\new_[5423]_  | ~\new_[4884]_ ;
  assign \new_[4199]_  = ~\new_[4889]_  | ~\new_[5562]_  | ~\new_[4890]_ ;
  assign \new_[4200]_  = \\rf_conf10_reg[0] ;
  assign \new_[4201]_  = \\rf_conf10_reg[10] ;
  assign \new_[4202]_  = \\rf_conf10_reg[11] ;
  assign \new_[4203]_  = \\rf_conf10_reg[12] ;
  assign \new_[4204]_  = \\rf_conf10_reg[13] ;
  assign \new_[4205]_  = \\rf_conf10_reg[14] ;
  assign \new_[4206]_  = \\rf_conf10_reg[15] ;
  assign \new_[4207]_  = \\rf_conf10_reg[1] ;
  assign \new_[4208]_  = \\rf_conf10_reg[2] ;
  assign \new_[4209]_  = \\rf_conf10_reg[3] ;
  assign \new_[4210]_  = \\rf_conf10_reg[4] ;
  assign \new_[4211]_  = \\rf_conf10_reg[5] ;
  assign \new_[4212]_  = \\rf_conf10_reg[6] ;
  assign \new_[4213]_  = \\rf_conf10_reg[7] ;
  assign \new_[4214]_  = \\rf_conf10_reg[8] ;
  assign \new_[4215]_  = \\rf_conf10_reg[9] ;
  assign \new_[4216]_  = \\rf_conf11_reg[0] ;
  assign \new_[4217]_  = \\rf_conf11_reg[10] ;
  assign \new_[4218]_  = \\rf_conf11_reg[11] ;
  assign \new_[4219]_  = \\rf_conf11_reg[12] ;
  assign \new_[4220]_  = \\rf_conf11_reg[13] ;
  assign \new_[4221]_  = \\rf_conf11_reg[14] ;
  assign \new_[4222]_  = \\rf_conf11_reg[15] ;
  assign \new_[4223]_  = \\rf_conf11_reg[1] ;
  assign \new_[4224]_  = \\rf_conf11_reg[4] ;
  assign \new_[4225]_  = \\rf_conf11_reg[5] ;
  assign \new_[4226]_  = \\rf_conf11_reg[6] ;
  assign \new_[4227]_  = \\rf_conf11_reg[7] ;
  assign \new_[4228]_  = \\rf_conf11_reg[8] ;
  assign \new_[4229]_  = \\rf_conf11_reg[9] ;
  assign \new_[4230]_  = \\rf_conf11_reg[2] ;
  assign \new_[4231]_  = \\rf_conf11_reg[3] ;
  assign \new_[4232]_  = ~\new_[4893]_  | ~\new_[5430]_  | ~\new_[4891]_ ;
  assign \new_[4233]_  = \\rf_conf4_reg[0] ;
  assign \new_[4234]_  = \\rf_conf4_reg[10] ;
  assign \new_[4235]_  = \\rf_conf4_reg[11] ;
  assign \new_[4236]_  = \\rf_conf4_reg[12] ;
  assign \new_[4237]_  = \\rf_conf4_reg[13] ;
  assign \new_[4238]_  = \\rf_conf4_reg[14] ;
  assign \new_[4239]_  = \\rf_conf4_reg[15] ;
  assign \new_[4240]_  = \\rf_conf4_reg[1] ;
  assign \new_[4241]_  = \\rf_conf4_reg[4] ;
  assign \new_[4242]_  = \\rf_conf4_reg[5] ;
  assign \new_[4243]_  = \\rf_conf4_reg[6] ;
  assign \new_[4244]_  = \\rf_conf4_reg[7] ;
  assign \new_[4245]_  = \\rf_conf4_reg[8] ;
  assign \new_[4246]_  = \\rf_conf4_reg[9] ;
  assign \new_[4247]_  = \\rf_conf4_reg[2] ;
  assign \new_[4248]_  = \\rf_conf4_reg[3] ;
  assign \new_[4249]_  = \\rf_conf6_reg[0] ;
  assign \new_[4250]_  = \\rf_conf6_reg[10] ;
  assign \new_[4251]_  = \\rf_conf6_reg[11] ;
  assign \new_[4252]_  = \\rf_conf6_reg[12] ;
  assign \new_[4253]_  = \\rf_conf6_reg[13] ;
  assign \new_[4254]_  = \\rf_conf6_reg[14] ;
  assign \new_[4255]_  = \\rf_conf6_reg[15] ;
  assign \new_[4256]_  = \\rf_conf6_reg[1] ;
  assign \new_[4257]_  = \\rf_conf6_reg[4] ;
  assign \new_[4258]_  = \\rf_conf6_reg[5] ;
  assign \new_[4259]_  = \\rf_conf6_reg[6] ;
  assign \new_[4260]_  = \\rf_conf6_reg[7] ;
  assign \new_[4261]_  = \\rf_conf6_reg[8] ;
  assign \new_[4262]_  = \\rf_conf6_reg[9] ;
  assign \new_[4263]_  = \\rf_conf6_reg[2] ;
  assign \new_[4264]_  = \\rf_conf6_reg[3] ;
  assign \new_[4265]_  = \\rf_conf9_reg[0] ;
  assign \new_[4266]_  = \\rf_conf9_reg[10] ;
  assign \new_[4267]_  = \\rf_conf9_reg[11] ;
  assign \new_[4268]_  = \\rf_conf9_reg[12] ;
  assign \new_[4269]_  = \\rf_conf9_reg[13] ;
  assign \new_[4270]_  = \\rf_conf9_reg[14] ;
  assign \new_[4271]_  = \\rf_conf9_reg[15] ;
  assign \new_[4272]_  = \\rf_conf9_reg[1] ;
  assign \new_[4273]_  = \\rf_conf9_reg[2] ;
  assign \new_[4274]_  = \\rf_conf9_reg[3] ;
  assign \new_[4275]_  = \\rf_conf9_reg[4] ;
  assign \new_[4276]_  = \\rf_conf9_reg[5] ;
  assign \new_[4277]_  = \\rf_conf9_reg[6] ;
  assign \new_[4278]_  = \\rf_conf9_reg[7] ;
  assign \new_[4279]_  = \\rf_conf9_reg[8] ;
  assign \new_[4280]_  = \\rf_conf9_reg[9] ;
  assign \new_[4281]_  = ~\new_[4897]_  | ~\new_[5083]_  | ~\new_[4898]_ ;
  assign \new_[4282]_  = ~\new_[5443]_  | ~\new_[5444]_  | ~\new_[5084]_  | ~\new_[4899]_ ;
  assign \new_[4283]_  = ~\new_[4901]_  | ~\new_[5085]_  | ~\new_[4900]_ ;
  assign n5174 = ~\new_[5046]_  | ~\new_[4828]_ ;
  assign n5179 = ~\new_[5047]_  | ~\new_[4829]_ ;
  assign n5184 = ~\new_[5048]_  | ~\new_[4830]_ ;
  assign n5189 = ~\new_[5049]_  | ~\new_[4831]_ ;
  assign n5194 = ~\new_[5050]_  | ~\new_[4832]_ ;
  assign n5199 = ~\new_[5051]_  | ~\new_[4833]_ ;
  assign n5204 = ~\new_[5052]_  | ~\new_[4834]_ ;
  assign n5209 = ~\new_[5053]_  | ~\new_[4835]_ ;
  assign n5214 = ~\new_[5054]_  | ~\new_[4836]_ ;
  assign n5219 = ~\new_[5055]_  | ~\new_[4837]_ ;
  assign n5224 = ~\new_[5056]_  | ~\new_[4838]_ ;
  assign n5229 = ~\new_[5057]_  | ~\new_[4839]_ ;
  assign n5234 = ~\new_[5058]_  | ~\new_[4840]_ ;
  assign n5244 = ~\new_[5060]_  | ~\new_[4842]_ ;
  assign n5239 = ~\new_[5059]_  | ~\new_[4841]_ ;
  assign n5249 = ~\new_[5061]_  | ~\new_[4843]_ ;
  assign \new_[4300]_  = ~\new_[17053]_  | ~\new_[17054]_  | ~\new_[5088]_  | ~\new_[16175]_ ;
  assign \new_[4301]_  = ~\new_[17716]_  | ~\new_[14641]_  | ~\new_[5092]_  | ~\new_[17713]_ ;
  assign \new_[4302]_  = ~\new_[17662]_  | ~\new_[18557]_  | ~\new_[5093]_  | ~\new_[17720]_ ;
  assign \new_[4303]_  = ~\new_[4600]_ ;
  assign \new_[4304]_  = ~\new_[4601]_ ;
  assign \new_[4305]_  = ~\new_[4602]_ ;
  assign \new_[4306]_  = ~\new_[4603]_ ;
  assign \new_[4307]_  = ~\new_[4604]_ ;
  assign \new_[4308]_  = ~\new_[4605]_ ;
  assign \new_[4309]_  = ~\new_[4606]_ ;
  assign \new_[4310]_  = ~\new_[4607]_ ;
  assign \new_[4311]_  = ~\new_[4608]_ ;
  assign \new_[4312]_  = ~\new_[4609]_ ;
  assign \new_[4313]_  = ~\new_[4610]_ ;
  assign \new_[4314]_  = ~\new_[4611]_ ;
  assign \new_[4315]_  = ~\new_[4612]_ ;
  assign \new_[4316]_  = ~\new_[4613]_ ;
  assign \new_[4317]_  = ~\new_[4614]_ ;
  assign \new_[4318]_  = ~\new_[4615]_ ;
  assign \new_[4319]_  = ~\new_[4616]_ ;
  assign \new_[4320]_  = ~\new_[4617]_ ;
  assign \new_[4321]_  = ~\new_[4618]_ ;
  assign \new_[4322]_  = ~\new_[4619]_ ;
  assign \new_[4323]_  = ~\new_[4620]_ ;
  assign \new_[4324]_  = ~\new_[4621]_ ;
  assign \new_[4325]_  = ~\new_[4622]_ ;
  assign \new_[4326]_  = ~\new_[4623]_ ;
  assign \new_[4327]_  = ~\new_[4624]_ ;
  assign \new_[4328]_  = ~\new_[4625]_ ;
  assign \new_[4329]_  = ~\new_[4626]_ ;
  assign \new_[4330]_  = ~\new_[4627]_ ;
  assign \new_[4331]_  = ~\new_[4628]_ ;
  assign \new_[4332]_  = ~\new_[4629]_ ;
  assign \new_[4333]_  = ~\new_[4630]_ ;
  assign \new_[4334]_  = ~\new_[16872]_  | ~\new_[18564]_  | ~\new_[5086]_  | ~\new_[14659]_ ;
  assign \new_[4335]_  = ~\new_[4631]_ ;
  assign \new_[4336]_  = ~\new_[4632]_ ;
  assign \new_[4337]_  = ~\new_[4633]_ ;
  assign \new_[4338]_  = ~\new_[16878]_  | ~\new_[17738]_  | ~\new_[5087]_  | ~\new_[16071]_ ;
  assign \new_[4339]_  = ~\new_[4634]_ ;
  assign \new_[4340]_  = ~\new_[4635]_ ;
  assign \new_[4341]_  = ~\new_[4636]_ ;
  assign \new_[4342]_  = ~\new_[4637]_ ;
  assign \new_[4343]_  = ~\new_[4638]_ ;
  assign \new_[4344]_  = ~\new_[4639]_ ;
  assign \new_[4345]_  = ~\new_[4640]_ ;
  assign \new_[4346]_  = ~\new_[4641]_ ;
  assign \new_[4347]_  = ~\new_[4642]_ ;
  assign \new_[4348]_  = ~\new_[4643]_ ;
  assign \new_[4349]_  = ~\new_[4644]_ ;
  assign \new_[4350]_  = ~\new_[4645]_ ;
  assign \new_[4351]_  = ~\new_[4646]_ ;
  assign \new_[4352]_  = ~\new_[4647]_ ;
  assign \new_[4353]_  = ~\new_[4648]_ ;
  assign \new_[4354]_  = ~\new_[4650]_ ;
  assign \new_[4355]_  = ~\new_[4651]_ ;
  assign \new_[4356]_  = ~\new_[4653]_ ;
  assign \new_[4357]_  = ~\new_[4654]_ ;
  assign \new_[4358]_  = ~\new_[4655]_ ;
  assign \new_[4359]_  = ~\new_[4656]_ ;
  assign \new_[4360]_  = ~\new_[4657]_ ;
  assign \new_[4361]_  = ~\new_[4658]_ ;
  assign \new_[4362]_  = ~\new_[4659]_ ;
  assign \new_[4363]_  = ~\new_[4660]_ ;
  assign \new_[4364]_  = ~\new_[4661]_ ;
  assign \new_[4365]_  = ~\new_[4662]_ ;
  assign \new_[4366]_  = ~\new_[4663]_ ;
  assign \new_[4367]_  = ~\new_[4664]_ ;
  assign \new_[4368]_  = ~\new_[4665]_ ;
  assign \new_[4369]_  = ~\new_[4666]_ ;
  assign \new_[4370]_  = ~\new_[4667]_ ;
  assign \new_[4371]_  = ~\new_[4668]_ ;
  assign \new_[4372]_  = ~\new_[4669]_ ;
  assign \new_[4373]_  = ~\new_[4670]_ ;
  assign \new_[4374]_  = ~\new_[4671]_ ;
  assign \new_[4375]_  = ~\new_[4672]_ ;
  assign \new_[4376]_  = ~\new_[4673]_ ;
  assign \new_[4377]_  = ~\new_[4674]_ ;
  assign \new_[4378]_  = ~\new_[4675]_ ;
  assign \new_[4379]_  = ~\new_[17107]_  | ~\new_[16196]_  | ~\new_[5094]_  | ~\new_[17061]_ ;
  assign \new_[4380]_  = ~\new_[4676]_ ;
  assign \new_[4381]_  = ~\new_[4677]_ ;
  assign \new_[4382]_  = ~\new_[17045]_  | ~\new_[16195]_  | ~\new_[5095]_  | ~\new_[17065]_ ;
  assign \new_[4383]_  = ~\new_[4678]_ ;
  assign \new_[4384]_  = ~\new_[4679]_ ;
  assign \new_[4385]_  = ~\new_[4680]_ ;
  assign \new_[4386]_  = ~\new_[4682]_ ;
  assign \new_[4387]_  = ~\new_[4685]_ ;
  assign \new_[4388]_  = ~\new_[4741]_  & ~\new_[5081]_ ;
  assign \new_[4389]_  = ~\new_[4690]_ ;
  assign \new_[4390]_  = ~\new_[4693]_ ;
  assign \new_[4391]_  = ~\new_[4696]_ ;
  assign \new_[4392]_  = ~\new_[4697]_ ;
  assign \new_[4393]_  = ~\new_[4698]_ ;
  assign \new_[4394]_  = ~\new_[4699]_ ;
  assign \new_[4395]_  = ~\new_[4700]_ ;
  assign \new_[4396]_  = ~\new_[4701]_ ;
  assign \new_[4397]_  = ~\new_[4702]_ ;
  assign \new_[4398]_  = ~\new_[4703]_ ;
  assign \new_[4399]_  = ~\new_[4704]_ ;
  assign \new_[4400]_  = ~\new_[4705]_ ;
  assign \new_[4401]_  = ~\new_[4706]_ ;
  assign \new_[4402]_  = ~\new_[4707]_ ;
  assign \new_[4403]_  = ~\new_[4708]_ ;
  assign \new_[4404]_  = ~\new_[4709]_ ;
  assign \new_[4405]_  = ~\new_[4710]_ ;
  assign \new_[4406]_  = ~\new_[4711]_ ;
  assign \new_[4407]_  = ~\new_[4712]_ ;
  assign \new_[4408]_  = ~\new_[4713]_ ;
  assign \new_[4409]_  = ~\new_[4714]_ ;
  assign \new_[4410]_  = ~\new_[4715]_ ;
  assign \new_[4411]_  = ~\new_[4716]_ ;
  assign \new_[4412]_  = ~\new_[4717]_ ;
  assign \new_[4413]_  = ~\new_[4718]_ ;
  assign \new_[4414]_  = ~\new_[17090]_  | ~\new_[17091]_  | ~\new_[5096]_  | ~\new_[17089]_ ;
  assign \new_[4415]_  = ~\new_[4719]_ ;
  assign \new_[4416]_  = ~\new_[4720]_ ;
  assign \new_[4417]_  = ~\new_[4721]_ ;
  assign \new_[4418]_  = ~\new_[16220]_  | ~\new_[17888]_  | ~\new_[5097]_  | ~\new_[17098]_ ;
  assign \new_[4419]_  = ~\new_[4722]_ ;
  assign \new_[4420]_  = ~\new_[4723]_ ;
  assign \new_[4421]_  = ~\new_[4724]_ ;
  assign \new_[4422]_  = ~\new_[4725]_ ;
  assign \new_[4423]_  = ~\new_[4726]_ ;
  assign \new_[4424]_  = ~\new_[4727]_ ;
  assign \new_[4425]_  = ~\new_[4728]_ ;
  assign \new_[4426]_  = ~\new_[4729]_ ;
  assign \new_[4427]_  = ~\new_[4730]_ ;
  assign \new_[4428]_  = ~\new_[4731]_ ;
  assign \new_[4429]_  = ~\new_[4732]_ ;
  assign \new_[4430]_  = ~\new_[4733]_ ;
  assign \new_[4431]_  = ~\new_[4734]_ ;
  assign \new_[4432]_  = ~\new_[4735]_ ;
  assign \new_[4433]_  = ~\new_[4736]_ ;
  assign \new_[4434]_  = ~\new_[4737]_ ;
  assign \new_[4435]_  = ~\new_[25314]_  | ~\new_[25965]_  | ~\new_[4880]_  | ~\new_[27423]_ ;
  assign \new_[4436]_  = ~\new_[26148]_  | ~\new_[26436]_  | ~\new_[4882]_  | ~\new_[27102]_ ;
  assign \new_[4437]_  = ~\new_[23959]_  | ~\new_[25293]_  | ~\new_[5101]_  | ~\new_[25274]_ ;
  assign \new_[4438]_  = \\rf_conf8_reg[0] ;
  assign \new_[4439]_  = \\rf_conf8_reg[10] ;
  assign \new_[4440]_  = \\rf_conf8_reg[11] ;
  assign \new_[4441]_  = \\rf_conf8_reg[12] ;
  assign \new_[4442]_  = \\rf_conf8_reg[13] ;
  assign \new_[4443]_  = \\rf_conf8_reg[14] ;
  assign \new_[4444]_  = \\rf_conf8_reg[15] ;
  assign \new_[4445]_  = \\rf_conf8_reg[1] ;
  assign \new_[4446]_  = \\rf_conf8_reg[4] ;
  assign \new_[4447]_  = \\rf_conf8_reg[5] ;
  assign \new_[4448]_  = \\rf_conf8_reg[6] ;
  assign \new_[4449]_  = \\rf_conf8_reg[7] ;
  assign \new_[4450]_  = \\rf_conf8_reg[8] ;
  assign \new_[4451]_  = \\rf_conf8_reg[9] ;
  assign \new_[4452]_  = \\rf_conf8_reg[2] ;
  assign \new_[4453]_  = \\rf_conf8_reg[3] ;
  assign \new_[4454]_  = rf_rf_we_reg;
  assign \new_[4455]_  = ~rf_rf_ack_reg;
  assign n5254 = ~\new_[4982]_  | ~\new_[5276]_ ;
  assign n5259 = ~\new_[4983]_  | ~\new_[5277]_ ;
  assign n5264 = ~\new_[4984]_  | ~\new_[5278]_ ;
  assign n5269 = ~\new_[4985]_  | ~\new_[5279]_ ;
  assign n5274 = ~\new_[4986]_  | ~\new_[5280]_ ;
  assign n5279 = ~\new_[4987]_  | ~\new_[5281]_ ;
  assign n5284 = ~\new_[4988]_  | ~\new_[5282]_ ;
  assign n5289 = ~\new_[4989]_  | ~\new_[5283]_ ;
  assign n5294 = ~\new_[4990]_  | ~\new_[5284]_ ;
  assign n5299 = ~\new_[4991]_  | ~\new_[5285]_ ;
  assign n5304 = ~\new_[4992]_  | ~\new_[5286]_ ;
  assign n5309 = ~\new_[4993]_  | ~\new_[5287]_ ;
  assign n5314 = ~\new_[4994]_  | ~\new_[5288]_ ;
  assign n5319 = ~\new_[4995]_  | ~\new_[5289]_ ;
  assign n5324 = ~\new_[4996]_  | ~\new_[5290]_ ;
  assign n5329 = ~\new_[4997]_  | ~\new_[5291]_ ;
  assign n5334 = ~\new_[4998]_  | ~\new_[5212]_ ;
  assign n5339 = ~\new_[4999]_  | ~\new_[5213]_ ;
  assign n5344 = ~\new_[5000]_  | ~\new_[5214]_ ;
  assign n5349 = ~\new_[5001]_  | ~\new_[5215]_ ;
  assign n5354 = ~\new_[5002]_  | ~\new_[5216]_ ;
  assign n5359 = ~\new_[5003]_  | ~\new_[5217]_ ;
  assign n5364 = ~\new_[5004]_  | ~\new_[5218]_ ;
  assign n5369 = ~\new_[5005]_  | ~\new_[5219]_ ;
  assign n5374 = ~\new_[5006]_  | ~\new_[5220]_ ;
  assign n5379 = ~\new_[5007]_  | ~\new_[5221]_ ;
  assign n5384 = ~\new_[5008]_  | ~\new_[5223]_ ;
  assign n5389 = ~\new_[5009]_  | ~\new_[5222]_ ;
  assign n5394 = ~\new_[5010]_  | ~\new_[5224]_ ;
  assign n5399 = ~\new_[5011]_  | ~\new_[5225]_ ;
  assign n5404 = ~\new_[5012]_  | ~\new_[5226]_ ;
  assign n5409 = ~\new_[5013]_  | ~\new_[5227]_ ;
  assign n5414 = ~\new_[5228]_  | ~\new_[5014]_ ;
  assign n5424 = ~\new_[5230]_  | ~\new_[5016]_ ;
  assign n5419 = ~\new_[5229]_  | ~\new_[5015]_ ;
  assign n5429 = ~\new_[5017]_  | ~\new_[5231]_ ;
  assign n5434 = ~\new_[5232]_  | ~\new_[5018]_ ;
  assign n5439 = ~\new_[5233]_  | ~\new_[5019]_ ;
  assign n5444 = ~\new_[5020]_  | ~\new_[5234]_ ;
  assign n5449 = ~\new_[5021]_  | ~\new_[5235]_ ;
  assign n5559 = ~\new_[5236]_  | ~\new_[5022]_ ;
  assign n5564 = ~\new_[5237]_  | ~\new_[5023]_ ;
  assign n5454 = ~\new_[5238]_  | ~\new_[5024]_ ;
  assign n5459 = ~\new_[5239]_  | ~\new_[5025]_ ;
  assign n5464 = ~\new_[5240]_  | ~\new_[5026]_ ;
  assign n5469 = ~\new_[5241]_  | ~\new_[5027]_ ;
  assign n5474 = ~\new_[5242]_  | ~\new_[5028]_ ;
  assign n5479 = ~\new_[5029]_  | ~\new_[5243]_ ;
  assign n5484 = ~\new_[5030]_  | ~\new_[5244]_ ;
  assign n5489 = ~\new_[5031]_  | ~\new_[5245]_ ;
  assign n5494 = ~\new_[5032]_  | ~\new_[5246]_ ;
  assign n5504 = ~\new_[5034]_  | ~\new_[5248]_ ;
  assign n5509 = ~\new_[5035]_  | ~\new_[5249]_ ;
  assign n5499 = ~\new_[5033]_  | ~\new_[5247]_ ;
  assign n5514 = ~\new_[5036]_  | ~\new_[5250]_ ;
  assign n5519 = ~\new_[5037]_  | ~\new_[5251]_ ;
  assign n5569 = ~\new_[5038]_  | ~\new_[5252]_ ;
  assign n5524 = ~\new_[5040]_  | ~\new_[5253]_ ;
  assign n5534 = ~\new_[5041]_  | ~\new_[5255]_ ;
  assign n5529 = ~\new_[5039]_  | ~\new_[5254]_ ;
  assign n5539 = ~\new_[5042]_  | ~\new_[5256]_ ;
  assign n5544 = ~\new_[5043]_  | ~\new_[5257]_ ;
  assign n5549 = ~\new_[5044]_  | ~\new_[5258]_ ;
  assign n5554 = ~\new_[5045]_  | ~\new_[5259]_ ;
  assign n5574 = ~\new_[4918]_  | ~\new_[5308]_ ;
  assign n5579 = ~\new_[4919]_  | ~\new_[5309]_ ;
  assign n5584 = ~\new_[4920]_  | ~\new_[5310]_ ;
  assign n5594 = ~\new_[4922]_  | ~\new_[5312]_ ;
  assign n5589 = ~\new_[4921]_  | ~\new_[5311]_ ;
  assign n5599 = ~\new_[4923]_  | ~\new_[5313]_ ;
  assign n5604 = ~\new_[4924]_  | ~\new_[5314]_ ;
  assign n5609 = ~\new_[4925]_  | ~\new_[5315]_ ;
  assign n5614 = ~\new_[4926]_  | ~\new_[5316]_ ;
  assign n5619 = ~\new_[4927]_  | ~\new_[5317]_ ;
  assign n5624 = ~\new_[4928]_  | ~\new_[5318]_ ;
  assign n5629 = ~\new_[4929]_  | ~\new_[5319]_ ;
  assign n5634 = ~\new_[4930]_  | ~\new_[5320]_ ;
  assign n5639 = ~\new_[4931]_  | ~\new_[5321]_ ;
  assign n5644 = ~\new_[4932]_  | ~\new_[5322]_ ;
  assign n5649 = ~\new_[4933]_  | ~\new_[5323]_ ;
  assign n5654 = ~\new_[4934]_  | ~\new_[5324]_ ;
  assign n5659 = ~\new_[4935]_  | ~\new_[5325]_ ;
  assign n5664 = ~\new_[4936]_  | ~\new_[5326]_ ;
  assign n5669 = ~\new_[4937]_  | ~\new_[5327]_ ;
  assign n5674 = ~\new_[4938]_  | ~\new_[5328]_ ;
  assign n5679 = ~\new_[4939]_  | ~\new_[5329]_ ;
  assign n5689 = ~\new_[4941]_  | ~\new_[5331]_ ;
  assign n5684 = ~\new_[4940]_  | ~\new_[5330]_ ;
  assign n5694 = ~\new_[4942]_  | ~\new_[5332]_ ;
  assign n5699 = ~\new_[4943]_  | ~\new_[5333]_ ;
  assign n5704 = ~\new_[4944]_  | ~\new_[5334]_ ;
  assign n5709 = ~\new_[4945]_  | ~\new_[5335]_ ;
  assign n5714 = ~\new_[4946]_  | ~\new_[5336]_ ;
  assign n5719 = ~\new_[4947]_  | ~\new_[5337]_ ;
  assign n5724 = ~\new_[4948]_  | ~\new_[5338]_ ;
  assign n5729 = ~\new_[4949]_  | ~\new_[5339]_ ;
  assign n5734 = ~\new_[4950]_  | ~\new_[5340]_ ;
  assign n5739 = ~\new_[4951]_  | ~\new_[5341]_ ;
  assign n5744 = ~\new_[4952]_  | ~\new_[5342]_ ;
  assign n5749 = ~\new_[4953]_  | ~\new_[5343]_ ;
  assign n5754 = ~\new_[4954]_  | ~\new_[5344]_ ;
  assign n5759 = ~\new_[4955]_  | ~\new_[5345]_ ;
  assign n5764 = ~\new_[4956]_  | ~\new_[5346]_ ;
  assign n5769 = ~\new_[4957]_  | ~\new_[5347]_ ;
  assign n5774 = ~\new_[4958]_  | ~\new_[5348]_ ;
  assign n5784 = ~\new_[4960]_  | ~\new_[5350]_ ;
  assign n5779 = ~\new_[4959]_  | ~\new_[5349]_ ;
  assign n5789 = ~\new_[4961]_  | ~\new_[5351]_ ;
  assign n5794 = ~\new_[4962]_  | ~\new_[5352]_ ;
  assign n5799 = ~\new_[4963]_  | ~\new_[5353]_ ;
  assign n5804 = ~\new_[4964]_  | ~\new_[5354]_ ;
  assign n5809 = ~\new_[4965]_  | ~\new_[5355]_ ;
  assign n5814 = ~\new_[5062]_  | ~\new_[5260]_ ;
  assign n5819 = ~\new_[5063]_  | ~\new_[5261]_ ;
  assign n5824 = ~\new_[5064]_  | ~\new_[5262]_ ;
  assign n5829 = ~\new_[5065]_  | ~\new_[5263]_ ;
  assign n5834 = ~\new_[5066]_  | ~\new_[5264]_ ;
  assign n5839 = ~\new_[5067]_  | ~\new_[5265]_ ;
  assign n5844 = ~\new_[5068]_  | ~\new_[5266]_ ;
  assign n5849 = ~\new_[5070]_  | ~\new_[5267]_ ;
  assign n5859 = ~\new_[5071]_  | ~\new_[5269]_ ;
  assign n5854 = ~\new_[5069]_  | ~\new_[5268]_ ;
  assign n5864 = ~\new_[5072]_  | ~\new_[5270]_ ;
  assign n5869 = ~\new_[5073]_  | ~\new_[5271]_ ;
  assign n5874 = ~\new_[5074]_  | ~\new_[5272]_ ;
  assign n5879 = ~\new_[5075]_  | ~\new_[5273]_ ;
  assign n5884 = ~\new_[5076]_  | ~\new_[5274]_ ;
  assign n5889 = ~\new_[5077]_  | ~\new_[5275]_ ;
  assign n5894 = ~\new_[5388]_  | ~\new_[4966]_ ;
  assign n5904 = ~\new_[5390]_  | ~\new_[4968]_ ;
  assign n5899 = ~\new_[5389]_  | ~\new_[4967]_ ;
  assign n5909 = ~\new_[5391]_  | ~\new_[4969]_ ;
  assign n5914 = ~\new_[5392]_  | ~\new_[4970]_ ;
  assign n5919 = ~\new_[5393]_  | ~\new_[4971]_ ;
  assign n5924 = ~\new_[5394]_  | ~\new_[4972]_ ;
  assign n5929 = ~\new_[5395]_  | ~\new_[4973]_ ;
  assign n5934 = ~\new_[5396]_  | ~\new_[4974]_ ;
  assign n5939 = ~\new_[5397]_  | ~\new_[4975]_ ;
  assign n5944 = ~\new_[5398]_  | ~\new_[4976]_ ;
  assign n5949 = ~\new_[5399]_  | ~\new_[4977]_ ;
  assign n5954 = ~\new_[5400]_  | ~\new_[4978]_ ;
  assign n5959 = ~\new_[5401]_  | ~\new_[4979]_ ;
  assign n5964 = ~\new_[5402]_  | ~\new_[4980]_ ;
  assign n5969 = ~\new_[5403]_  | ~\new_[4981]_ ;
  assign \new_[4600]_  = ~\new_[24545]_  | ~\new_[24559]_  | ~\new_[5100]_  | ~\new_[27970]_ ;
  assign \new_[4601]_  = ~\new_[26014]_  | ~\new_[25566]_  | ~\new_[5102]_  | ~\new_[27880]_ ;
  assign \new_[4602]_  = ~\new_[25967]_  | ~\new_[24734]_  | ~\new_[5103]_  | ~\new_[27419]_ ;
  assign \new_[4603]_  = ~\new_[25918]_  | ~\new_[25458]_  | ~\new_[5104]_  | ~\new_[27063]_ ;
  assign \new_[4604]_  = ~\new_[25542]_  | ~\new_[25877]_  | ~\new_[5105]_  | ~\new_[27389]_ ;
  assign \new_[4605]_  = ~\new_[24053]_  | ~\new_[26002]_  | ~\new_[5113]_  | ~\new_[25723]_ ;
  assign \new_[4606]_  = ~\new_[26441]_  | ~\new_[25323]_  | ~\new_[5106]_  | ~\new_[27319]_ ;
  assign \new_[4607]_  = ~\new_[26747]_  | ~\new_[25324]_  | ~\new_[5107]_  | ~\new_[25322]_ ;
  assign \new_[4608]_  = ~\new_[25333]_  | ~\new_[25693]_  | ~\new_[5108]_  | ~\new_[27354]_ ;
  assign \new_[4609]_  = ~\new_[27786]_  | ~\new_[25792]_  | ~\new_[5109]_  | ~\new_[24567]_ ;
  assign \new_[4610]_  = ~\new_[27304]_  | ~\new_[25339]_  | ~\new_[5110]_  | ~\new_[25725]_ ;
  assign \new_[4611]_  = ~\new_[25789]_  | ~\new_[25805]_  | ~\new_[5111]_  | ~\new_[27143]_ ;
  assign \new_[4612]_  = ~\new_[27336]_  | ~\new_[25777]_  | ~\new_[5112]_  | ~\new_[25803]_ ;
  assign \new_[4613]_  = ~\new_[27324]_  | ~\new_[25350]_  | ~\new_[5114]_  | ~\new_[25778]_ ;
  assign \new_[4614]_  = ~\new_[27090]_  | ~\new_[25750]_  | ~\new_[5115]_  | ~\new_[25352]_ ;
  assign \new_[4615]_  = ~\new_[27092]_  | ~\new_[25739]_  | ~\new_[5116]_  | ~\new_[25361]_ ;
  assign \new_[4616]_  = ~\new_[27522]_  | ~\new_[25727]_  | ~\new_[5117]_  | ~\new_[26481]_ ;
  assign \new_[4617]_  = ~\new_[27286]_  | ~\new_[25374]_  | ~\new_[5118]_  | ~\new_[25371]_ ;
  assign \new_[4618]_  = ~\new_[26154]_  | ~\new_[25685]_  | ~\new_[5119]_  | ~\new_[27101]_ ;
  assign \new_[4619]_  = ~\new_[27265]_  | ~\new_[25389]_  | ~\new_[5120]_  | ~\new_[25385]_ ;
  assign \new_[4620]_  = ~\new_[27335]_  | ~\new_[25575]_  | ~\new_[5121]_  | ~\new_[25651]_ ;
  assign \new_[4621]_  = ~\new_[27108]_  | ~\new_[25628]_  | ~\new_[5122]_  | ~\new_[25399]_ ;
  assign \new_[4622]_  = ~\new_[27229]_  | ~\new_[24686]_  | ~\new_[5123]_  | ~\new_[25406]_ ;
  assign \new_[4623]_  = ~\new_[27117]_  | ~\new_[24603]_  | ~\new_[5124]_  | ~\new_[25412]_ ;
  assign \new_[4624]_  = ~\new_[27190]_  | ~\new_[24536]_  | ~\new_[5125]_  | ~\new_[25563]_ ;
  assign \new_[4625]_  = ~\new_[24034]_  | ~\new_[26445]_  | ~\new_[5126]_  | ~\new_[25521]_ ;
  assign \new_[4626]_  = ~\new_[24015]_  | ~\new_[27174]_  | ~\new_[32337]_  | ~\new_[22665]_ ;
  assign \new_[4627]_  = ~\new_[24061]_  | ~\new_[26619]_  | ~\new_[5127]_  | ~\new_[22637]_ ;
  assign \new_[4628]_  = ~\new_[24064]_  | ~\new_[27061]_  | ~\new_[5128]_  | ~\new_[22584]_ ;
  assign \new_[4629]_  = ~\new_[24019]_  | ~\new_[27220]_  | ~\new_[5129]_  | ~\new_[22644]_ ;
  assign \new_[4630]_  = ~\new_[24022]_  | ~\new_[27273]_  | ~\new_[5130]_  | ~\new_[22604]_ ;
  assign \new_[4631]_  = ~\new_[24023]_  | ~\new_[27187]_  | ~\new_[5131]_  | ~\new_[22568]_ ;
  assign \new_[4632]_  = ~\new_[24046]_  | ~\new_[26722]_  | ~\new_[5132]_  | ~\new_[22599]_ ;
  assign \new_[4633]_  = ~\new_[23969]_  | ~\new_[26671]_  | ~\new_[5133]_  | ~\new_[22564]_ ;
  assign \new_[4634]_  = ~\new_[24040]_  | ~\new_[27235]_  | ~\new_[5134]_  | ~\new_[22626]_ ;
  assign \new_[4635]_  = ~\new_[24190]_  | ~\new_[27484]_  | ~\new_[5135]_  | ~\new_[22603]_ ;
  assign \new_[4636]_  = ~\new_[27197]_  | ~\new_[24637]_  | ~\new_[5136]_  | ~\new_[27684]_ ;
  assign \new_[4637]_  = ~\new_[23967]_  | ~\new_[27195]_  | ~\new_[5137]_  | ~\new_[22684]_ ;
  assign \new_[4638]_  = ~\new_[23130]_  | ~\new_[27234]_  | ~\new_[5138]_  | ~\new_[21581]_ ;
  assign \new_[4639]_  = ~\new_[24143]_  | ~\new_[27417]_  | ~\new_[5139]_  | ~\new_[22674]_ ;
  assign \new_[4640]_  = ~\new_[24130]_  | ~\new_[27134]_  | ~\new_[5140]_  | ~\new_[22668]_ ;
  assign \new_[4641]_  = ~\new_[27205]_  | ~\new_[25899]_  | ~\new_[5141]_  | ~\new_[27225]_ ;
  assign \new_[4642]_  = ~\new_[24031]_  | ~\new_[25496]_  | ~\new_[5145]_  | ~\new_[25816]_ ;
  assign \new_[4643]_  = ~\new_[23813]_  | ~\new_[27208]_  | ~\new_[5142]_  | ~\new_[22660]_ ;
  assign \new_[4644]_  = ~\new_[23150]_  | ~\new_[27201]_  | ~\new_[5143]_  | ~\new_[22576]_ ;
  assign \new_[4645]_  = ~\new_[27214]_  | ~\new_[24717]_  | ~\new_[5144]_  | ~\new_[27212]_ ;
  assign \new_[4646]_  = ~\new_[27219]_  | ~\new_[25788]_  | ~\new_[5146]_  | ~\new_[27338]_ ;
  assign \new_[4647]_  = ~\new_[26802]_  | ~\new_[25597]_  | ~\new_[5147]_  | ~\new_[27078]_ ;
  assign \new_[4648]_  = ~\new_[27230]_  | ~\new_[25604]_  | ~\new_[5148]_  | ~\new_[26579]_ ;
  assign \new_[4649]_  = ~\new_[12870]_  | ~\new_[12872]_  | ~\new_[5098]_  | ~\new_[14335]_ ;
  assign \new_[4650]_  = ~\new_[27237]_  | ~\new_[25609]_  | ~\new_[5149]_  | ~\new_[27146]_ ;
  assign \new_[4651]_  = ~\new_[27242]_  | ~\new_[25529]_  | ~\new_[5150]_  | ~\new_[27113]_ ;
  assign \new_[4652]_  = ~\new_[14337]_  | ~\new_[12883]_  | ~\new_[5099]_  | ~\new_[12879]_ ;
  assign \new_[4653]_  = ~\new_[27097]_  | ~\new_[25624]_  | ~\new_[5151]_  | ~\new_[27193]_ ;
  assign \new_[4654]_  = ~\new_[27355]_  | ~\new_[25743]_  | ~\new_[5152]_  | ~\new_[27469]_ ;
  assign \new_[4655]_  = ~\new_[25337]_  | ~\new_[25942]_  | ~\new_[5153]_  | ~\new_[25633]_ ;
  assign \new_[4656]_  = ~\new_[27424]_  | ~\new_[25632]_  | ~\new_[5154]_  | ~\new_[27768]_ ;
  assign \new_[4657]_  = ~\new_[26944]_  | ~\new_[25391]_  | ~\new_[5155]_  | ~\new_[27398]_ ;
  assign \new_[4658]_  = ~\new_[27480]_  | ~\new_[25810]_  | ~\new_[5156]_  | ~\new_[27307]_ ;
  assign \new_[4659]_  = ~\new_[27153]_  | ~\new_[25666]_  | ~\new_[5157]_  | ~\new_[27258]_ ;
  assign \new_[4660]_  = ~\new_[25347]_  | ~\new_[25565]_  | ~\new_[5158]_  | ~\new_[26126]_ ;
  assign \new_[4661]_  = ~\new_[24159]_  | ~\new_[25414]_  | ~\new_[5167]_  | ~\new_[25535]_ ;
  assign \new_[4662]_  = ~\new_[27274]_  | ~\new_[24602]_  | ~\new_[5159]_  | ~\new_[27228]_ ;
  assign \new_[4663]_  = ~\new_[24486]_  | ~\new_[25379]_  | ~\new_[5160]_  | ~\new_[25958]_ ;
  assign \new_[4664]_  = ~\new_[27306]_  | ~\new_[25635]_  | ~\new_[5161]_  | ~\new_[27050]_ ;
  assign \new_[4665]_  = ~\new_[26141]_  | ~\new_[25672]_  | ~\new_[32276]_  | ~\new_[25523]_ ;
  assign \new_[4666]_  = ~\new_[24576]_  | ~\new_[24681]_  | ~\new_[31998]_  | ~\new_[26017]_ ;
  assign \new_[4667]_  = ~\new_[25692]_  | ~\new_[25736]_  | ~\new_[5163]_  | ~\new_[25690]_ ;
  assign \new_[4668]_  = ~\new_[25813]_  | ~\new_[25668]_  | ~\new_[5164]_  | ~\new_[25411]_ ;
  assign \new_[4669]_  = ~\new_[24172]_  | ~\new_[25754]_  | ~\new_[5168]_  | ~\new_[25376]_ ;
  assign \new_[4670]_  = ~\new_[25712]_  | ~\new_[25476]_  | ~\new_[5165]_  | ~\new_[25930]_ ;
  assign \new_[4671]_  = ~\new_[24729]_  | ~\new_[25983]_  | ~\new_[5166]_  | ~\new_[26301]_ ;
  assign \new_[4672]_  = ~\new_[26558]_  | ~\new_[25311]_  | ~\new_[5169]_  | ~\new_[24706]_ ;
  assign \new_[4673]_  = ~\new_[25332]_  | ~\new_[25548]_  | ~\new_[5170]_  | ~\new_[25746]_ ;
  assign \new_[4674]_  = ~\new_[25601]_  | ~\new_[26070]_  | ~\new_[5171]_  | ~\new_[26075]_ ;
  assign \new_[4675]_  = ~\new_[25764]_  | ~\new_[26048]_  | ~\new_[5172]_  | ~\new_[26062]_ ;
  assign \new_[4676]_  = ~\new_[23651]_  | ~\new_[25593]_  | ~\new_[5162]_  | ~\new_[25467]_ ;
  assign \new_[4677]_  = ~\new_[25797]_  | ~\new_[25779]_  | ~\new_[5173]_  | ~\new_[25307]_ ;
  assign \new_[4678]_  = ~\new_[24103]_  | ~\new_[25594]_  | ~\new_[5174]_  | ~\new_[23111]_ ;
  assign \new_[4679]_  = ~\new_[24110]_  | ~\new_[25276]_  | ~\new_[5192]_  | ~\new_[25663]_ ;
  assign \new_[4680]_  = ~\new_[25820]_  | ~\new_[25338]_  | ~\new_[5175]_  | ~\new_[26032]_ ;
  assign \new_[4681]_  = ~\new_[5195]_  & ~\new_[5080]_ ;
  assign \new_[4682]_  = ~\new_[24167]_  | ~\new_[25359]_  | ~\new_[5176]_  | ~\new_[23970]_ ;
  assign \new_[4683]_  = ~\new_[4886]_  & ~\new_[5424]_ ;
  assign \new_[4684]_  = ~\new_[5428]_  | ~\new_[5663]_  | ~\new_[5427]_ ;
  assign \new_[4685]_  = ~\new_[24087]_  | ~\new_[25897]_  | ~\new_[5179]_  | ~\new_[25716]_ ;
  assign \new_[4686]_  = ~\new_[4892]_  & ~\new_[5082]_ ;
  assign \new_[4687]_  = ~\new_[5433]_  | ~\new_[5432]_  | ~\new_[5574]_ ;
  assign \new_[4688]_  = ~\new_[4896]_  & ~\new_[5435]_ ;
  assign \new_[4689]_  = ~\new_[5581]_  | ~\new_[5582]_  | ~\new_[5436]_ ;
  assign \new_[4690]_  = ~\new_[25556]_  | ~\new_[25527]_  | ~\new_[5177]_  | ~\new_[25707]_ ;
  assign \new_[4691]_  = ~\new_[5439]_  | ~\new_[5586]_  | ~\new_[32065]_ ;
  assign \new_[4692]_  = ~\new_[5442]_  | ~\new_[5591]_  | ~\new_[5589]_ ;
  assign \new_[4693]_  = ~\new_[23177]_  | ~\new_[25500]_  | ~\new_[5178]_  | ~\new_[24533]_ ;
  assign \new_[4694]_  = ~\new_[5601]_  | ~\new_[5602]_  | ~\new_[5446]_ ;
  assign \new_[4695]_  = ~\new_[5449]_  | ~\new_[5673]_  | ~\new_[5606]_ ;
  assign \new_[4696]_  = ~\new_[24089]_  | ~\new_[25384]_  | ~\new_[5180]_  | ~\new_[24072]_ ;
  assign \new_[4697]_  = ~\new_[25960]_  | ~\new_[25650]_  | ~\new_[5181]_  | ~\new_[25438]_ ;
  assign \new_[4698]_  = ~\new_[24076]_  | ~\new_[25430]_  | ~\new_[5182]_  | ~\new_[24067]_ ;
  assign \new_[4699]_  = ~\new_[23998]_  | ~\new_[25631]_  | ~\new_[5183]_  | ~\new_[24171]_ ;
  assign \new_[4700]_  = ~\new_[23100]_  | ~\new_[25599]_  | ~\new_[5184]_  | ~\new_[23519]_ ;
  assign \new_[4701]_  = ~\new_[24093]_  | ~\new_[25677]_  | ~\new_[5185]_  | ~\new_[24092]_ ;
  assign \new_[4702]_  = ~\new_[24095]_  | ~\new_[25833]_  | ~\new_[5186]_  | ~\new_[24066]_ ;
  assign \new_[4703]_  = ~\new_[24096]_  | ~\new_[24618]_  | ~\new_[5187]_  | ~\new_[24036]_ ;
  assign \new_[4704]_  = ~\new_[24102]_  | ~\new_[25845]_  | ~\new_[5188]_  | ~\new_[24100]_ ;
  assign \new_[4705]_  = ~\new_[23993]_  | ~\new_[25524]_  | ~\new_[5189]_  | ~\new_[24105]_ ;
  assign \new_[4706]_  = ~\new_[24109]_  | ~\new_[25446]_  | ~\new_[5190]_  | ~\new_[24108]_ ;
  assign \new_[4707]_  = ~\new_[24112]_  | ~\new_[25360]_  | ~\new_[5191]_  | ~\new_[24030]_ ;
  assign \new_[4708]_  = ~\new_[24018]_  | ~\new_[25887]_  | ~\new_[4853]_  | ~\new_[25876]_ ;
  assign \new_[4709]_  = ~\new_[24027]_  | ~\new_[25285]_  | ~\new_[5193]_  | ~\new_[24116]_ ;
  assign \new_[4710]_  = ~\new_[24026]_  | ~\new_[25233]_  | ~\new_[5194]_  | ~\new_[23179]_ ;
  assign \new_[4711]_  = ~\new_[24148]_  | ~\new_[25988]_  | ~\new_[4854]_  | ~\new_[24714]_ ;
  assign \new_[4712]_  = ~\new_[23612]_  | ~\new_[26023]_  | ~\new_[4876]_  | ~\new_[26026]_ ;
  assign \new_[4713]_  = ~\new_[24164]_  | ~\new_[24606]_  | ~\new_[4856]_  | ~\new_[26034]_ ;
  assign \new_[4714]_  = ~\new_[26473]_  | ~\new_[25865]_  | ~\new_[4855]_  | ~\new_[25577]_ ;
  assign \new_[4715]_  = ~\new_[25652]_  | ~\new_[26029]_  | ~\new_[4857]_  | ~\new_[26028]_ ;
  assign \new_[4716]_  = ~\new_[25721]_  | ~\new_[24626]_  | ~\new_[4858]_  | ~\new_[24629]_ ;
  assign \new_[4717]_  = ~\new_[26044]_  | ~\new_[25785]_  | ~\new_[4859]_  | ~\new_[25794]_ ;
  assign \new_[4718]_  = ~\new_[26335]_  | ~\new_[26052]_  | ~\new_[4860]_  | ~\new_[26050]_ ;
  assign \new_[4719]_  = ~\new_[26177]_  | ~\new_[26057]_  | ~\new_[4861]_  | ~\new_[25741]_ ;
  assign \new_[4720]_  = ~\new_[24587]_  | ~\new_[26040]_  | ~\new_[4862]_  | ~\new_[24588]_ ;
  assign \new_[4721]_  = ~\new_[26066]_  | ~\new_[25689]_  | ~\new_[4863]_  | ~\new_[26064]_ ;
  assign \new_[4722]_  = ~\new_[25671]_  | ~\new_[26072]_  | ~\new_[4864]_  | ~\new_[26071]_ ;
  assign \new_[4723]_  = ~\new_[24551]_  | ~\new_[26079]_  | ~\new_[4865]_  | ~\new_[26078]_ ;
  assign \new_[4724]_  = ~\new_[26086]_  | ~\new_[26095]_  | ~\new_[4866]_  | ~\new_[27451]_ ;
  assign \new_[4725]_  = ~\new_[26087]_  | ~\new_[25623]_  | ~\new_[4867]_  | ~\new_[24539]_ ;
  assign \new_[4726]_  = ~\new_[26094]_  | ~\new_[25588]_  | ~\new_[4868]_  | ~\new_[26092]_ ;
  assign \new_[4727]_  = ~\new_[25569]_  | ~\new_[26099]_  | ~\new_[4869]_  | ~\new_[25574]_ ;
  assign \new_[4728]_  = ~\new_[24187]_  | ~\new_[26559]_  | ~\new_[4881]_  | ~\new_[26129]_ ;
  assign \new_[4729]_  = ~\new_[24516]_  | ~\new_[26516]_  | ~\new_[4871]_  | ~\new_[26107]_ ;
  assign \new_[4730]_  = ~\new_[26101]_  | ~\new_[26104]_  | ~\new_[4870]_  | ~\new_[27955]_ ;
  assign \new_[4731]_  = ~\new_[25539]_  | ~\new_[26555]_  | ~\new_[4872]_  | ~\new_[25545]_ ;
  assign \new_[4732]_  = ~\new_[25473]_  | ~\new_[26113]_  | ~\new_[4874]_  | ~\new_[26805]_ ;
  assign \new_[4733]_  = ~\new_[26539]_  | ~\new_[26109]_  | ~\new_[4873]_  | ~\new_[26106]_ ;
  assign \new_[4734]_  = ~\new_[25468]_  | ~\new_[25534]_  | ~\new_[4875]_  | ~\new_[25479]_ ;
  assign \new_[4735]_  = ~\new_[26125]_  | ~\new_[26119]_  | ~\new_[4877]_  | ~\new_[27859]_ ;
  assign \new_[4736]_  = ~\new_[26127]_  | ~\new_[26004]_  | ~\new_[4878]_  | ~\new_[27473]_ ;
  assign \new_[4737]_  = ~\new_[26134]_  | ~\new_[25921]_  | ~\new_[4879]_  | ~\new_[27479]_ ;
  assign s15_cyc_o = ~\new_[5450]_  & ~n7424;
  assign \new_[4739]_  = ~\new_[5661]_  & ~\new_[5425]_ ;
  assign \new_[4740]_  = ~\new_[5555]_  & ~\new_[5426]_ ;
  assign \new_[4741]_  = ~\new_[5705]_  | ~\new_[5794]_  | ~\new_[5792]_  | ~\new_[5793]_ ;
  assign \new_[4742]_  = ~\new_[5563]_  & ~\new_[5429]_ ;
  assign \new_[4743]_  = ~\new_[5666]_  & ~\new_[5431]_ ;
  assign \new_[4744]_  = ~\new_[5575]_  & ~\new_[5434]_ ;
  assign \new_[4745]_  = ~\new_[5583]_  & ~\new_[5437]_ ;
  assign \new_[4746]_  = ~\new_[5587]_  & ~\new_[5440]_ ;
  assign \new_[4747]_  = ~\new_[5603]_  & ~\new_[5447]_ ;
  assign n5974 = ~\new_[5292]_  | ~\new_[5452]_ ;
  assign n5979 = ~\new_[5293]_  | ~\new_[5453]_ ;
  assign n5984 = ~\new_[5294]_  | ~\new_[5454]_ ;
  assign n5989 = ~\new_[5295]_  | ~\new_[5455]_ ;
  assign n5994 = ~\new_[5296]_  | ~\new_[5456]_ ;
  assign n6004 = ~\new_[5298]_  | ~\new_[5458]_ ;
  assign n6009 = ~\new_[5299]_  | ~\new_[5459]_ ;
  assign n5999 = ~\new_[5297]_  | ~\new_[5457]_ ;
  assign n6014 = ~\new_[5300]_  | ~\new_[5460]_ ;
  assign n6019 = ~\new_[5301]_  | ~\new_[5461]_ ;
  assign n6024 = ~\new_[5302]_  | ~\new_[5462]_ ;
  assign n6029 = ~\new_[5303]_  | ~\new_[5463]_ ;
  assign n6034 = ~\new_[5304]_  | ~\new_[5464]_ ;
  assign n6039 = ~\new_[5305]_  | ~\new_[5465]_ ;
  assign n6044 = ~\new_[5306]_  | ~\new_[5467]_ ;
  assign n6049 = ~\new_[5307]_  | ~\new_[5466]_ ;
  assign n6054 = ~\new_[5516]_  | ~\new_[5196]_ ;
  assign n6059 = ~\new_[5518]_  | ~\new_[5197]_ ;
  assign n6069 = ~\new_[5519]_  | ~\new_[5199]_ ;
  assign n6064 = ~\new_[5517]_  | ~\new_[5198]_ ;
  assign n6074 = ~\new_[5520]_  | ~\new_[5200]_ ;
  assign n6079 = ~\new_[5521]_  | ~\new_[5201]_ ;
  assign n6084 = ~\new_[5522]_  | ~\new_[5202]_ ;
  assign n6089 = ~\new_[5523]_  | ~\new_[5203]_ ;
  assign n6124 = ~\new_[5524]_  | ~\new_[5204]_ ;
  assign n6129 = ~\new_[5525]_  | ~\new_[5205]_ ;
  assign n6094 = ~\new_[5526]_  | ~\new_[5206]_ ;
  assign n6099 = ~\new_[5527]_  | ~\new_[5207]_ ;
  assign n6104 = ~\new_[5528]_  | ~\new_[5208]_ ;
  assign n6109 = ~\new_[5529]_  | ~\new_[5209]_ ;
  assign n6114 = ~\new_[5530]_  | ~\new_[5210]_ ;
  assign n6119 = ~\new_[5531]_  | ~\new_[5211]_ ;
  assign n6134 = ~\new_[5356]_  | ~\new_[5468]_ ;
  assign n6139 = ~\new_[5357]_  | ~\new_[5469]_ ;
  assign n6144 = ~\new_[5358]_  | ~\new_[5470]_ ;
  assign n6149 = ~\new_[5359]_  | ~\new_[5471]_ ;
  assign n6154 = ~\new_[5360]_  | ~\new_[5472]_ ;
  assign n6159 = ~\new_[5361]_  | ~\new_[5473]_ ;
  assign n6164 = ~\new_[5362]_  | ~\new_[5474]_ ;
  assign n6169 = ~\new_[5363]_  | ~\new_[5475]_ ;
  assign n6204 = ~\new_[5364]_  | ~\new_[5476]_ ;
  assign n6209 = ~\new_[5365]_  | ~\new_[5477]_ ;
  assign n6174 = ~\new_[5366]_  | ~\new_[5478]_ ;
  assign n6179 = ~\new_[5367]_  | ~\new_[5479]_ ;
  assign n6184 = ~\new_[5368]_  | ~\new_[5480]_ ;
  assign n6189 = ~\new_[5369]_  | ~\new_[5481]_ ;
  assign n6194 = ~\new_[5370]_  | ~\new_[5482]_ ;
  assign n6199 = ~\new_[5371]_  | ~\new_[5483]_ ;
  assign n6214 = ~\new_[5372]_  | ~\new_[5484]_ ;
  assign n6219 = ~\new_[5373]_  | ~\new_[5485]_ ;
  assign n6224 = ~\new_[5374]_  | ~\new_[5486]_ ;
  assign n6229 = ~\new_[5375]_  | ~\new_[5487]_ ;
  assign n6234 = ~\new_[5376]_  | ~\new_[5488]_ ;
  assign n6239 = ~\new_[5377]_  | ~\new_[5489]_ ;
  assign n6244 = ~\new_[5378]_  | ~\new_[5490]_ ;
  assign n6249 = ~\new_[5379]_  | ~\new_[5491]_ ;
  assign n6284 = ~\new_[5380]_  | ~\new_[5492]_ ;
  assign n6289 = ~\new_[5381]_  | ~\new_[5493]_ ;
  assign n6254 = ~\new_[5382]_  | ~\new_[5494]_ ;
  assign n6259 = ~\new_[5383]_  | ~\new_[5495]_ ;
  assign n6264 = ~\new_[5384]_  | ~\new_[5496]_ ;
  assign n6269 = ~\new_[5385]_  | ~\new_[5497]_ ;
  assign n6274 = ~\new_[5386]_  | ~\new_[5498]_ ;
  assign n6279 = ~\new_[5387]_  | ~\new_[5499]_ ;
  assign n6294 = ~\new_[5404]_  | ~\new_[5500]_ ;
  assign n6299 = ~\new_[5405]_  | ~\new_[5501]_ ;
  assign n6304 = ~\new_[5406]_  | ~\new_[5502]_ ;
  assign n6309 = ~\new_[5407]_  | ~\new_[5503]_ ;
  assign n6314 = ~\new_[5408]_  | ~\new_[5504]_ ;
  assign n6319 = ~\new_[5409]_  | ~\new_[5505]_ ;
  assign n6324 = ~\new_[5410]_  | ~\new_[5506]_ ;
  assign n6329 = ~\new_[5411]_  | ~\new_[5507]_ ;
  assign n6334 = ~\new_[5412]_  | ~\new_[5508]_ ;
  assign n6339 = ~\new_[5413]_  | ~\new_[5509]_ ;
  assign n6344 = ~\new_[5414]_  | ~\new_[5510]_ ;
  assign n6349 = ~\new_[5415]_  | ~\new_[5511]_ ;
  assign n6354 = ~\new_[5416]_  | ~\new_[5512]_ ;
  assign n6359 = ~\new_[5417]_  | ~\new_[5513]_ ;
  assign n6364 = ~\new_[5418]_  | ~\new_[5514]_ ;
  assign n6369 = ~\new_[5419]_  | ~\new_[5515]_ ;
  assign \new_[4828]_  = ~\s15_data_o[0]  | ~\new_[5619]_ ;
  assign \new_[4829]_  = ~\s15_data_o[10]  | ~\new_[5619]_ ;
  assign \new_[4830]_  = ~\s15_data_o[11]  | ~\new_[5619]_ ;
  assign \new_[4831]_  = ~\s15_data_o[12]  | ~\new_[5619]_ ;
  assign \new_[4832]_  = ~\s15_data_o[13]  | ~\new_[5619]_ ;
  assign \new_[4833]_  = ~\s15_data_o[14]  | ~\new_[5619]_ ;
  assign \new_[4834]_  = ~\s15_data_o[15]  | ~\new_[5619]_ ;
  assign \new_[4835]_  = ~\s15_data_o[1]  | ~\new_[5619]_ ;
  assign \new_[4836]_  = ~\s15_data_o[2]  | ~\new_[5619]_ ;
  assign \new_[4837]_  = ~\s15_data_o[3]  | ~\new_[5619]_ ;
  assign \new_[4838]_  = ~\s15_data_o[4]  | ~\new_[5619]_ ;
  assign \new_[4839]_  = ~\s15_data_o[5]  | ~\new_[5619]_ ;
  assign \new_[4840]_  = ~\s15_data_o[6]  | ~\new_[5619]_ ;
  assign \new_[4841]_  = ~\s15_data_o[7]  | ~\new_[5619]_ ;
  assign \new_[4842]_  = ~\s15_data_o[8]  | ~\new_[5619]_ ;
  assign \new_[4843]_  = ~\s15_data_o[9]  | ~\new_[5619]_ ;
  assign \new_[4844]_  = ~\new_[11326]_  | ~\new_[5451]_ ;
  assign \new_[4845]_  = ~\new_[32127]_  | ~\new_[5451]_  | ~\new_[13527]_ ;
  assign \new_[4846]_  = ~\new_[32343]_  | ~\new_[5451]_  | ~\new_[8851]_ ;
  assign \new_[4847]_  = ~\new_[5597]_  | ~\new_[5445]_  | ~\new_[5596]_ ;
  assign \new_[4848]_  = ~\new_[32260]_  | ~\new_[5451]_  | ~\new_[31981]_ ;
  assign \new_[4849]_  = ~\new_[32049]_  | ~\new_[5451]_  | ~\new_[14838]_ ;
  assign \new_[4850]_  = ~\new_[32161]_  | ~\new_[5451]_  | ~\new_[14844]_ ;
  assign \new_[4851]_  = ~\new_[27781]_  | ~\new_[5451]_  | ~\new_[14856]_ ;
  assign \new_[4852]_  = ~\new_[32321]_  | ~\new_[5451]_  | ~\new_[14861]_ ;
  assign \new_[4853]_  = (~\new_[5654]_  | ~\new_[26491]_ ) & (~\s13_data_i[20]  | ~\new_[28726]_ );
  assign \new_[4854]_  = (~\new_[5655]_  | ~\new_[29043]_ ) & (~\s13_data_i[19]  | ~\new_[28726]_ );
  assign \new_[4855]_  = (~\new_[32267]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[32260]_ );
  assign \new_[4856]_  = (~\new_[5656]_  | ~\new_[26491]_ ) & (~\s13_data_i[18]  | ~\new_[28726]_ );
  assign \new_[4857]_  = (~\new_[32267]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[32260]_ );
  assign \new_[4858]_  = (~\new_[32267]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[32260]_ );
  assign \new_[4859]_  = (~\new_[32267]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[32260]_ );
  assign \new_[4860]_  = (~\new_[32267]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[32260]_ );
  assign \new_[4861]_  = (~\new_[32267]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[28712]_ );
  assign \new_[4862]_  = (~\new_[32267]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[32260]_ );
  assign \new_[4863]_  = (~\new_[32267]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[32260]_ );
  assign \new_[4864]_  = (~\new_[32267]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[28712]_ );
  assign \new_[4865]_  = (~\new_[32267]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[28712]_ );
  assign \new_[4866]_  = (~\new_[32056]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[24571]_ );
  assign \new_[4867]_  = (~\new_[32267]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[32260]_ );
  assign \new_[4868]_  = (~\new_[32267]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[28712]_ );
  assign \new_[4869]_  = (~\new_[32267]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[32260]_ );
  assign \new_[4870]_  = (~\new_[32056]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[24571]_ );
  assign \new_[4871]_  = (~\new_[5657]_  | ~\new_[29043]_ ) & (~\s13_data_i[17]  | ~\new_[28726]_ );
  assign \new_[4872]_  = (~\new_[32267]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[32260]_ );
  assign \new_[4873]_  = (~\new_[32267]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[32260]_ );
  assign \new_[4874]_  = (~\new_[32056]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[32049]_ );
  assign \new_[4875]_  = (~\new_[32267]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[32260]_ );
  assign \new_[4876]_  = (~\new_[31999]_  | ~\new_[26491]_ ) & (~\s13_data_i[28]  | ~\new_[28726]_ );
  assign \new_[4877]_  = (~\new_[32056]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[24571]_ );
  assign \new_[4878]_  = (~\new_[32056]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[32049]_ );
  assign \new_[4879]_  = (~\new_[32056]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[24571]_ );
  assign \new_[4880]_  = (~\new_[32056]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[32049]_ );
  assign \new_[4881]_  = (~\new_[5658]_  | ~\new_[29043]_ ) & (~\s13_data_i[27]  | ~\new_[28726]_ );
  assign \new_[4882]_  = (~\new_[32056]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[32049]_ );
  assign \new_[4883]_  = ~\new_[5659]_  & ~\new_[5548]_ ;
  assign \new_[4884]_  = ~\new_[5549]_  & ~\new_[5660]_ ;
  assign \new_[4885]_  = ~\new_[5550]_  & ~\new_[5551]_ ;
  assign \new_[4886]_  = ~\new_[5726]_  | ~\new_[5837]_  | ~\new_[5701]_  | ~\new_[5782]_ ;
  assign \new_[4887]_  = ~\new_[5552]_  & ~\new_[5553]_ ;
  assign \new_[4888]_  = ~\new_[5662]_  & ~\new_[5556]_ ;
  assign \new_[4889]_  = ~\new_[5560]_  & ~\new_[5561]_ ;
  assign \new_[4890]_  = ~\new_[5559]_  & ~\new_[5664]_ ;
  assign \new_[4891]_  = ~\new_[5567]_  & ~\new_[5665]_ ;
  assign \new_[4892]_  = ~\new_[5738]_  | ~\new_[5842]_  | ~\new_[5709]_  | ~\new_[5866]_ ;
  assign \new_[4893]_  = ~\new_[5568]_  & ~\new_[5569]_ ;
  assign \new_[4894]_  = ~\new_[5570]_  & ~\new_[5571]_ ;
  assign \new_[4895]_  = ~\new_[5576]_  & ~\new_[5667]_ ;
  assign \new_[4896]_  = ~\new_[5743]_  | ~\new_[5744]_  | ~\new_[5844]_  | ~\new_[5872]_ ;
  assign \new_[4897]_  = ~\new_[5579]_  & ~\new_[5580]_ ;
  assign \new_[4898]_  = ~\new_[5578]_  & ~\new_[5668]_ ;
  assign \new_[4899]_  = ~\new_[5671]_  & ~\new_[5594]_ ;
  assign \new_[4900]_  = ~\new_[5598]_  & ~\new_[5672]_ ;
  assign \new_[4901]_  = ~\new_[5599]_  & ~\new_[5600]_ ;
  assign n6374 = ~\new_[5532]_  | ~\new_[5630]_ ;
  assign n6379 = ~\new_[5533]_  | ~\new_[5631]_ ;
  assign n6384 = ~\new_[5534]_  | ~\new_[5632]_ ;
  assign n6389 = ~\new_[5535]_  | ~\new_[5633]_ ;
  assign n6394 = ~\new_[5536]_  | ~\new_[5634]_ ;
  assign n6399 = ~\new_[5537]_  | ~\new_[5635]_ ;
  assign n6404 = ~\new_[5538]_  | ~\new_[5636]_ ;
  assign n6409 = ~\new_[5539]_  | ~\new_[5637]_ ;
  assign n6444 = ~\new_[5540]_  | ~\new_[5638]_ ;
  assign n6449 = ~\new_[5542]_  | ~\new_[5639]_ ;
  assign n6419 = ~\new_[5543]_  | ~\new_[5641]_ ;
  assign n6414 = ~\new_[5541]_  | ~\new_[5640]_ ;
  assign n6424 = ~\new_[5544]_  | ~\new_[5642]_ ;
  assign n6429 = ~\new_[5545]_  | ~\new_[5643]_ ;
  assign n6434 = ~\new_[5546]_  | ~\new_[5644]_ ;
  assign n6439 = ~\new_[5547]_  | ~\new_[5645]_ ;
  assign \new_[4918]_  = ~\new_[5620]_  | ~\new_[4101]_ ;
  assign \new_[4919]_  = ~\new_[5620]_  | ~\new_[4102]_ ;
  assign \new_[4920]_  = ~\new_[5620]_  | ~\new_[4103]_ ;
  assign \new_[4921]_  = ~\new_[5620]_  | ~\new_[4104]_ ;
  assign \new_[4922]_  = ~\new_[5620]_  | ~\new_[4105]_ ;
  assign \new_[4923]_  = ~\new_[5620]_  | ~\new_[4106]_ ;
  assign \new_[4924]_  = ~\new_[5620]_  | ~\new_[4107]_ ;
  assign \new_[4925]_  = ~\new_[5620]_  | ~\new_[4108]_ ;
  assign \new_[4926]_  = ~\new_[5620]_  | ~\new_[4109]_ ;
  assign \new_[4927]_  = ~\new_[5620]_  | ~\new_[4110]_ ;
  assign \new_[4928]_  = ~\new_[5620]_  | ~\new_[4111]_ ;
  assign \new_[4929]_  = ~\new_[5620]_  | ~\new_[4112]_ ;
  assign \new_[4930]_  = ~\new_[5620]_  | ~\new_[4113]_ ;
  assign \new_[4931]_  = ~\new_[5620]_  | ~\new_[4114]_ ;
  assign \new_[4932]_  = ~\new_[5620]_  | ~\new_[4115]_ ;
  assign \new_[4933]_  = ~\new_[5620]_  | ~\new_[4116]_ ;
  assign \new_[4934]_  = ~\new_[5621]_  | ~\new_[4117]_ ;
  assign \new_[4935]_  = ~\new_[5621]_  | ~\new_[4118]_ ;
  assign \new_[4936]_  = ~\new_[5621]_  | ~\new_[4119]_ ;
  assign \new_[4937]_  = ~\new_[5621]_  | ~\new_[4120]_ ;
  assign \new_[4938]_  = ~\new_[5621]_  | ~\new_[4121]_ ;
  assign \new_[4939]_  = ~\new_[5621]_  | ~\new_[4122]_ ;
  assign \new_[4940]_  = ~\new_[5621]_  | ~\new_[4123]_ ;
  assign \new_[4941]_  = ~\new_[5621]_  | ~\new_[4124]_ ;
  assign \new_[4942]_  = ~\new_[5621]_  | ~\new_[4125]_ ;
  assign \new_[4943]_  = ~\new_[5621]_  | ~\new_[4126]_ ;
  assign \new_[4944]_  = ~\new_[5621]_  | ~\new_[4127]_ ;
  assign \new_[4945]_  = ~\new_[5621]_  | ~\new_[4128]_ ;
  assign \new_[4946]_  = ~\new_[5621]_  | ~\new_[4129]_ ;
  assign \new_[4947]_  = ~\new_[5621]_  | ~\new_[4130]_ ;
  assign \new_[4948]_  = ~\new_[5621]_  | ~\new_[4131]_ ;
  assign \new_[4949]_  = ~\new_[5621]_  | ~\new_[4132]_ ;
  assign \new_[4950]_  = ~\new_[5622]_  | ~\new_[4133]_ ;
  assign \new_[4951]_  = ~\new_[5622]_  | ~\new_[4134]_ ;
  assign \new_[4952]_  = ~\new_[5622]_  | ~\new_[4135]_ ;
  assign \new_[4953]_  = ~\new_[5622]_  | ~\new_[4136]_ ;
  assign \new_[4954]_  = ~\new_[5622]_  | ~\new_[4137]_ ;
  assign \new_[4955]_  = ~\new_[5622]_  | ~\new_[4138]_ ;
  assign \new_[4956]_  = ~\new_[5622]_  | ~\new_[4139]_ ;
  assign \new_[4957]_  = ~\new_[5622]_  | ~\new_[4140]_ ;
  assign \new_[4958]_  = ~\new_[5622]_  | ~\new_[4141]_ ;
  assign \new_[4959]_  = ~\new_[5622]_  | ~\new_[4142]_ ;
  assign \new_[4960]_  = ~\new_[5622]_  | ~\new_[4143]_ ;
  assign \new_[4961]_  = ~\new_[5622]_  | ~\new_[4144]_ ;
  assign \new_[4962]_  = ~\new_[5622]_  | ~\new_[4145]_ ;
  assign \new_[4963]_  = ~\new_[5622]_  | ~\new_[4146]_ ;
  assign \new_[4964]_  = ~\new_[5622]_  | ~\new_[4147]_ ;
  assign \new_[4965]_  = ~\new_[5622]_  | ~\new_[4148]_ ;
  assign \new_[4966]_  = ~\s15_data_o[0]  | ~\new_[5624]_ ;
  assign \new_[4967]_  = ~\s15_data_o[10]  | ~\new_[5624]_ ;
  assign \new_[4968]_  = ~\s15_data_o[11]  | ~\new_[5624]_ ;
  assign \new_[4969]_  = ~\s15_data_o[12]  | ~\new_[5624]_ ;
  assign \new_[4970]_  = ~\s15_data_o[13]  | ~\new_[5624]_ ;
  assign \new_[4971]_  = ~\s15_data_o[14]  | ~\new_[5624]_ ;
  assign \new_[4972]_  = ~\s15_data_o[15]  | ~\new_[5624]_ ;
  assign \new_[4973]_  = ~\s15_data_o[1]  | ~\new_[5624]_ ;
  assign \new_[4974]_  = ~\s15_data_o[2]  | ~\new_[5624]_ ;
  assign \new_[4975]_  = ~\s15_data_o[3]  | ~\new_[5624]_ ;
  assign \new_[4976]_  = ~\s15_data_o[4]  | ~\new_[5624]_ ;
  assign \new_[4977]_  = ~\s15_data_o[5]  | ~\new_[5624]_ ;
  assign \new_[4978]_  = ~\s15_data_o[6]  | ~\new_[5624]_ ;
  assign \new_[4979]_  = ~\s15_data_o[7]  | ~\new_[5624]_ ;
  assign \new_[4980]_  = ~\s15_data_o[8]  | ~\new_[5624]_ ;
  assign \new_[4981]_  = ~\s15_data_o[9]  | ~\new_[5624]_ ;
  assign \new_[4982]_  = ~\new_[5610]_  | ~\new_[4036]_ ;
  assign \new_[4983]_  = ~\new_[5610]_  | ~\new_[4037]_ ;
  assign \new_[4984]_  = ~\new_[5610]_  | ~\new_[4038]_ ;
  assign \new_[4985]_  = ~\new_[5610]_  | ~\new_[4039]_ ;
  assign \new_[4986]_  = ~\new_[5610]_  | ~\new_[4040]_ ;
  assign \new_[4987]_  = ~\new_[5610]_  | ~\new_[4041]_ ;
  assign \new_[4988]_  = ~\new_[5610]_  | ~\new_[4042]_ ;
  assign \new_[4989]_  = ~\new_[5610]_  | ~\new_[4043]_ ;
  assign \new_[4990]_  = ~\new_[5610]_  | ~\new_[4044]_ ;
  assign \new_[4991]_  = ~\new_[5610]_  | ~\new_[4045]_ ;
  assign \new_[4992]_  = ~\new_[5610]_  | ~\new_[4046]_ ;
  assign \new_[4993]_  = ~\new_[5610]_  | ~\new_[4047]_ ;
  assign \new_[4994]_  = ~\new_[5610]_  | ~\new_[4048]_ ;
  assign \new_[4995]_  = ~\new_[5610]_  | ~\new_[4049]_ ;
  assign \new_[4996]_  = ~\new_[5610]_  | ~\new_[4050]_ ;
  assign \new_[4997]_  = ~\new_[5610]_  | ~\new_[4051]_ ;
  assign \new_[4998]_  = ~\new_[5612]_  | ~\new_[4052]_ ;
  assign \new_[4999]_  = ~\new_[5611]_  | ~\new_[4053]_ ;
  assign \new_[5000]_  = ~\new_[5612]_  | ~\new_[4054]_ ;
  assign \new_[5001]_  = ~\new_[5611]_  | ~\new_[4055]_ ;
  assign \new_[5002]_  = ~\new_[5612]_  | ~\new_[4056]_ ;
  assign \new_[5003]_  = ~\new_[5611]_  | ~\new_[4057]_ ;
  assign \new_[5004]_  = ~\new_[5612]_  | ~\new_[4058]_ ;
  assign \new_[5005]_  = ~\new_[5613]_  | ~\new_[4059]_ ;
  assign \new_[5006]_  = ~\new_[5611]_  | ~\new_[4060]_ ;
  assign \new_[5007]_  = ~\new_[5613]_  | ~\new_[4061]_ ;
  assign \new_[5008]_  = ~\new_[5613]_  | ~\new_[4062]_ ;
  assign \new_[5009]_  = ~\new_[5612]_  | ~\new_[4063]_ ;
  assign \new_[5010]_  = ~\new_[5613]_  | ~\new_[4064]_ ;
  assign \new_[5011]_  = ~\new_[5613]_  | ~\new_[4065]_ ;
  assign \new_[5012]_  = ~\new_[5613]_  | ~\new_[4066]_ ;
  assign \new_[5013]_  = ~\new_[5612]_  | ~\new_[4067]_ ;
  assign \new_[5014]_  = ~\new_[5614]_  | ~\new_[4068]_ ;
  assign \new_[5015]_  = ~\new_[5614]_  | ~\new_[4069]_ ;
  assign \new_[5016]_  = ~\new_[5614]_  | ~\new_[4070]_ ;
  assign \new_[5017]_  = ~\new_[5614]_  | ~\new_[4071]_ ;
  assign \new_[5018]_  = ~\new_[5614]_  | ~\new_[4072]_ ;
  assign \new_[5019]_  = ~\new_[5614]_  | ~\new_[4073]_ ;
  assign \new_[5020]_  = ~\new_[5614]_  | ~\new_[4074]_ ;
  assign \new_[5021]_  = ~\new_[5614]_  | ~\new_[4075]_ ;
  assign \new_[5022]_  = ~\new_[5614]_  | ~\new_[4097]_ ;
  assign \new_[5023]_  = ~\new_[5614]_  | ~\new_[4098]_ ;
  assign \new_[5024]_  = ~\new_[5614]_  | ~\new_[4076]_ ;
  assign \new_[5025]_  = ~\new_[5614]_  | ~\new_[4077]_ ;
  assign \new_[5026]_  = ~\new_[5614]_  | ~\new_[4078]_ ;
  assign \new_[5027]_  = ~\new_[5614]_  | ~\new_[4079]_ ;
  assign \new_[5028]_  = ~\new_[5614]_  | ~\new_[4080]_ ;
  assign \new_[5029]_  = ~\new_[5614]_  | ~\new_[4081]_ ;
  assign \new_[5030]_  = ~\new_[5616]_  | ~\new_[4082]_ ;
  assign \new_[5031]_  = ~\new_[5615]_  | ~\new_[4083]_ ;
  assign \new_[5032]_  = ~\new_[5616]_  | ~\new_[4084]_ ;
  assign \new_[5033]_  = ~\new_[5615]_  | ~\new_[4085]_ ;
  assign \new_[5034]_  = ~\new_[5616]_  | ~\new_[4086]_ ;
  assign \new_[5035]_  = ~\new_[5615]_  | ~\new_[4087]_ ;
  assign \new_[5036]_  = ~\new_[5616]_  | ~\new_[4088]_ ;
  assign \new_[5037]_  = ~\new_[5617]_  | ~\new_[4089]_ ;
  assign \new_[5038]_  = ~\new_[5615]_  | ~\new_[4099]_ ;
  assign \new_[5039]_  = ~\new_[5617]_  | ~\new_[4091]_ ;
  assign \new_[5040]_  = ~\new_[5617]_  | ~\new_[4090]_ ;
  assign \new_[5041]_  = ~\new_[5616]_  | ~\new_[4092]_ ;
  assign \new_[5042]_  = ~\new_[5617]_  | ~\new_[4093]_ ;
  assign \new_[5043]_  = ~\new_[5617]_  | ~\new_[4094]_ ;
  assign \new_[5044]_  = ~\new_[5617]_  | ~\new_[4095]_ ;
  assign \new_[5045]_  = ~\new_[5616]_  | ~\new_[4096]_ ;
  assign \new_[5046]_  = ~\new_[5618]_  | ~\new_[3873]_ ;
  assign \new_[5047]_  = ~\new_[5618]_  | ~\new_[3874]_ ;
  assign \new_[5048]_  = ~\new_[5618]_  | ~\new_[3875]_ ;
  assign \new_[5049]_  = ~\new_[5618]_  | ~\new_[3876]_ ;
  assign \new_[5050]_  = ~\new_[5618]_  | ~\new_[3877]_ ;
  assign \new_[5051]_  = ~\new_[5618]_  | ~\new_[3878]_ ;
  assign \new_[5052]_  = ~\new_[5618]_  | ~\new_[3879]_ ;
  assign \new_[5053]_  = ~\new_[5618]_  | ~\new_[3880]_ ;
  assign \new_[5054]_  = ~\new_[5618]_  | ~\new_[3881]_ ;
  assign \new_[5055]_  = ~\new_[5618]_  | ~\new_[3882]_ ;
  assign \new_[5056]_  = ~\new_[5618]_  | ~\new_[3883]_ ;
  assign \new_[5057]_  = ~\new_[5618]_  | ~\new_[3884]_ ;
  assign \new_[5058]_  = ~\new_[5618]_  | ~\new_[3885]_ ;
  assign \new_[5059]_  = ~\new_[5618]_  | ~\new_[3886]_ ;
  assign \new_[5060]_  = ~\new_[5618]_  | ~\new_[3887]_ ;
  assign \new_[5061]_  = ~\new_[5618]_  | ~\new_[3888]_ ;
  assign \new_[5062]_  = ~\new_[5623]_  | ~\new_[4149]_ ;
  assign \new_[5063]_  = ~\new_[5623]_  | ~\new_[4150]_ ;
  assign \new_[5064]_  = ~\new_[5623]_  | ~\new_[4151]_ ;
  assign \new_[5065]_  = ~\new_[5623]_  | ~\new_[4152]_ ;
  assign \new_[5066]_  = ~\new_[5623]_  | ~\new_[4153]_ ;
  assign \new_[5067]_  = ~\new_[5623]_  | ~\new_[4154]_ ;
  assign \new_[5068]_  = ~\new_[5623]_  | ~\new_[4155]_ ;
  assign \new_[5069]_  = ~\new_[5623]_  | ~\new_[4157]_ ;
  assign \new_[5070]_  = ~\new_[5623]_  | ~\new_[4156]_ ;
  assign \new_[5071]_  = ~\new_[5623]_  | ~\new_[4158]_ ;
  assign \new_[5072]_  = ~\new_[5623]_  | ~\new_[4159]_ ;
  assign \new_[5073]_  = ~\new_[5623]_  | ~\new_[4160]_ ;
  assign \new_[5074]_  = ~\new_[5623]_  | ~\new_[4161]_ ;
  assign \new_[5075]_  = ~\new_[5623]_  | ~\new_[4162]_ ;
  assign \new_[5076]_  = ~\new_[5623]_  | ~\new_[4163]_ ;
  assign \new_[5077]_  = ~\new_[5623]_  | ~\new_[4164]_ ;
  assign n6459 = ~\new_[5629]_  & ~\new_[31781]_ ;
  assign n6454 = ~\new_[6201]_  & ~\new_[5629]_ ;
  assign \new_[5080]_  = ~\new_[5608]_  | ~\new_[5834]_ ;
  assign \new_[5081]_  = ~\new_[5609]_  | ~\new_[5840]_ ;
  assign \new_[5082]_  = ~\new_[5708]_  | ~\new_[5625]_ ;
  assign \new_[5083]_  = ~\new_[5626]_  & (~\new_[5941]_  | ~\new_[4098]_ );
  assign \new_[5084]_  = ~\new_[5627]_  & (~\new_[5941]_  | ~\new_[4079]_ );
  assign \new_[5085]_  = ~\new_[5628]_  & (~\new_[5941]_  | ~\new_[4080]_ );
  assign \new_[5086]_  = ~\new_[32049]_  | ~\new_[14838]_  | ~\new_[31988]_ ;
  assign \new_[5087]_  = ~\new_[32049]_  | ~\new_[14838]_  | ~\new_[31980]_ ;
  assign \new_[5088]_  = ~\new_[32343]_  | ~\new_[31989]_  | ~\new_[31980]_ ;
  assign \new_[5089]_  = ~\new_[27781]_  | ~\new_[14856]_  | ~\new_[31997]_ ;
  assign \new_[5090]_  = ~\new_[27781]_  | ~\new_[14856]_  | ~\new_[31985]_ ;
  assign \new_[5091]_  = ~\new_[32260]_  | ~\new_[31981]_  | ~\new_[31997]_ ;
  assign \new_[5092]_  = ~\new_[32127]_  | ~\new_[13527]_  | ~\new_[31988]_ ;
  assign \new_[5093]_  = ~\new_[32127]_  | ~\new_[13527]_  | ~\new_[31980]_ ;
  assign \new_[5094]_  = ~\new_[32161]_  | ~\new_[14844]_  | ~\new_[31988]_ ;
  assign \new_[5095]_  = ~\new_[32161]_  | ~\new_[14844]_  | ~\new_[31980]_ ;
  assign \new_[5096]_  = ~\new_[32321]_  | ~\new_[14861]_  | ~\new_[31988]_ ;
  assign \new_[5097]_  = ~\new_[32321]_  | ~\new_[14861]_  | ~\new_[31980]_ ;
  assign \new_[5098]_  = (~\new_[11326]_  | ~\new_[31988]_ ) & (~\new_[17757]_  | ~s13_err_i);
  assign \new_[5099]_  = (~\new_[11326]_  | ~\new_[31985]_ ) & (~\new_[17757]_  | ~s13_rty_i);
  assign \new_[5100]_  = (~\new_[32056]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[32049]_ );
  assign \new_[5101]_  = (~\new_[5646]_  | ~\new_[26491]_ ) & (~\s13_data_i[16]  | ~\new_[28726]_ );
  assign \new_[5102]_  = (~\new_[32056]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[32049]_ );
  assign \new_[5103]_  = (~\new_[32056]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[32049]_ );
  assign \new_[5104]_  = (~\new_[32056]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[32049]_ );
  assign \new_[5105]_  = (~\new_[32056]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[24571]_ );
  assign \new_[5106]_  = (~\new_[32056]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[24571]_ );
  assign \new_[5107]_  = (~\new_[32134]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[32127]_ );
  assign \new_[5108]_  = (~\new_[32056]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[24571]_ );
  assign \new_[5109]_  = (~\new_[32134]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[24630]_ );
  assign \new_[5110]_  = (~\new_[32134]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[24630]_ );
  assign \new_[5111]_  = (~\new_[32056]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[24571]_ );
  assign \new_[5112]_  = (~\new_[32134]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[24630]_ );
  assign \new_[5113]_  = (~\new_[5647]_  | ~\new_[26491]_ ) & (~\s13_data_i[26]  | ~\new_[28726]_ );
  assign \new_[5114]_  = (~\new_[32134]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[24630]_ );
  assign \new_[5115]_  = (~\new_[32134]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[32127]_ );
  assign \new_[5116]_  = (~\new_[32134]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[24630]_ );
  assign \new_[5117]_  = (~\new_[32134]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[24630]_ );
  assign \new_[5118]_  = (~\new_[32134]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[32127]_ );
  assign \new_[5119]_  = (~\new_[32134]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[24630]_ );
  assign \new_[5120]_  = (~\new_[32134]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[24630]_ );
  assign \new_[5121]_  = (~\new_[32134]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[24630]_ );
  assign \new_[5122]_  = (~\new_[32134]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[24630]_ );
  assign \new_[5123]_  = (~\new_[32134]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[24630]_ );
  assign \new_[5124]_  = (~\new_[32134]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[32127]_ );
  assign \new_[5125]_  = (~\new_[32134]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[24630]_ );
  assign \new_[5126]_  = (~\new_[5648]_  | ~\new_[29043]_ ) & (~\s13_data_i[25]  | ~\new_[28726]_ );
  assign \new_[5127]_  = (~\new_[32338]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[32343]_ );
  assign \new_[5128]_  = (~\new_[32338]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[26525]_ );
  assign \new_[5129]_  = (~\new_[32338]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[26525]_ );
  assign \new_[5130]_  = (~\new_[32338]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[32343]_ );
  assign \new_[5131]_  = (~\new_[32338]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[26525]_ );
  assign \new_[5132]_  = (~\new_[32338]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[26525]_ );
  assign \new_[5133]_  = (~\new_[32338]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[26525]_ );
  assign \new_[5134]_  = (~\new_[32338]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[26525]_ );
  assign \new_[5135]_  = (~\new_[32338]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[26525]_ );
  assign \new_[5136]_  = (~\new_[32168]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[32161]_ );
  assign \new_[5137]_  = (~\new_[32338]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[26525]_ );
  assign \new_[5138]_  = (~\new_[32338]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[26525]_ );
  assign \new_[5139]_  = (~\new_[32338]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[26525]_ );
  assign \new_[5140]_  = (~\new_[32338]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[32343]_ );
  assign \new_[5141]_  = (~\new_[32168]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[32161]_ );
  assign \new_[5142]_  = (~\new_[32338]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[26525]_ );
  assign \new_[5143]_  = (~\new_[32338]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[26525]_ );
  assign \new_[5144]_  = (~\new_[32168]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[26641]_ );
  assign \new_[5145]_  = (~\new_[5649]_  | ~\new_[26491]_ ) & (~\s13_data_i[24]  | ~\new_[28726]_ );
  assign \new_[5146]_  = (~\new_[32168]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[26641]_ );
  assign \new_[5147]_  = (~\new_[32168]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[32161]_ );
  assign \new_[5148]_  = (~\new_[32168]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[26641]_ );
  assign \new_[5149]_  = (~\new_[32168]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[26641]_ );
  assign \new_[5150]_  = (~\new_[32168]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[26641]_ );
  assign \new_[5151]_  = (~\new_[32168]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[26641]_ );
  assign \new_[5152]_  = (~\new_[32168]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[26641]_ );
  assign \new_[5153]_  = (~\new_[32327]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[32321]_ );
  assign \new_[5154]_  = (~\new_[32168]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[26641]_ );
  assign \new_[5155]_  = (~\new_[32168]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[26641]_ );
  assign \new_[5156]_  = (~\new_[32168]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[26641]_ );
  assign \new_[5157]_  = (~\new_[32168]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[32161]_ );
  assign \new_[5158]_  = (~\new_[32327]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[32321]_ );
  assign \new_[5159]_  = (~\new_[32168]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[26641]_ );
  assign \new_[5160]_  = (~\new_[5650]_  | ~\new_[29043]_ ) & (~\s13_data_i[23]  | ~\new_[28726]_ );
  assign \new_[5161]_  = (~\new_[32168]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[26641]_ );
  assign \new_[5162]_  = (~\new_[32339]_  | ~\new_[26491]_ ) & (~\new_[28726]_  | ~\s13_data_i[31] );
  assign \new_[5163]_  = (~\new_[32327]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[28695]_ );
  assign \new_[5164]_  = (~\new_[32327]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[28695]_ );
  assign \new_[5165]_  = (~\new_[32327]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[28695]_ );
  assign \new_[5166]_  = (~\new_[32327]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[28695]_ );
  assign \new_[5167]_  = (~\new_[5651]_  | ~\new_[29043]_ ) & (~\s13_data_i[30]  | ~\new_[28726]_ );
  assign \new_[5168]_  = (~\new_[5652]_  | ~\new_[26491]_ ) & (~\s13_data_i[22]  | ~\new_[28726]_ );
  assign \new_[5169]_  = (~\new_[32327]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[28695]_ );
  assign \new_[5170]_  = (~\new_[32327]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[28695]_ );
  assign \new_[5171]_  = (~\new_[32327]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[32321]_ );
  assign \new_[5172]_  = (~\new_[32327]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[28695]_ );
  assign \new_[5173]_  = (~\new_[32327]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[28695]_ );
  assign \new_[5174]_  = (~\new_[28851]_  | ~\s13_data_i[31] ) & (~\new_[32339]_  | ~\new_[29472]_ );
  assign \new_[5175]_  = (~\new_[32327]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[32321]_ );
  assign \new_[5176]_  = (~\new_[28851]_  | ~\s13_data_i[30] ) & (~\new_[5651]_  | ~\new_[29472]_ );
  assign \new_[5177]_  = (~\new_[32327]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[32321]_ );
  assign \new_[5178]_  = (~\new_[28851]_  | ~\s13_data_i[29] ) & (~\new_[32277]_  | ~\new_[29472]_ );
  assign \new_[5179]_  = (~\new_[5653]_  | ~\new_[26491]_ ) & (~\s13_data_i[21]  | ~\new_[28726]_ );
  assign \new_[5180]_  = (~\new_[28851]_  | ~\s13_data_i[28] ) & (~\new_[31999]_  | ~\new_[29472]_ );
  assign \new_[5181]_  = (~\new_[32327]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[32321]_ );
  assign \new_[5182]_  = (~\new_[28851]_  | ~\s13_data_i[27] ) & (~\new_[5658]_  | ~\new_[29472]_ );
  assign \new_[5183]_  = (~\new_[28851]_  | ~\s13_data_i[26] ) & (~\new_[5647]_  | ~\new_[29472]_ );
  assign \new_[5184]_  = (~\new_[28851]_  | ~\s13_data_i[25] ) & (~\new_[5648]_  | ~\new_[29472]_ );
  assign \new_[5185]_  = (~\new_[28851]_  | ~\s13_data_i[24] ) & (~\new_[5649]_  | ~\new_[29472]_ );
  assign \new_[5186]_  = (~\new_[28851]_  | ~\s13_data_i[23] ) & (~\new_[5650]_  | ~\new_[29472]_ );
  assign \new_[5187]_  = (~\new_[28851]_  | ~\s13_data_i[22] ) & (~\new_[5652]_  | ~\new_[29472]_ );
  assign \new_[5188]_  = (~\new_[28851]_  | ~\s13_data_i[21] ) & (~\new_[5653]_  | ~\new_[29472]_ );
  assign \new_[5189]_  = (~\new_[28851]_  | ~\s13_data_i[20] ) & (~\new_[5654]_  | ~\new_[29472]_ );
  assign \new_[5190]_  = (~\new_[28851]_  | ~\s13_data_i[19] ) & (~\new_[5655]_  | ~\new_[29472]_ );
  assign \new_[5191]_  = (~\new_[28851]_  | ~\s13_data_i[18] ) & (~\new_[5656]_  | ~\new_[29472]_ );
  assign \new_[5192]_  = (~\new_[32277]_  | ~\new_[29043]_ ) & (~\s13_data_i[29]  | ~\new_[28726]_ );
  assign \new_[5193]_  = (~\new_[28851]_  | ~\s13_data_i[17] ) & (~\new_[5657]_  | ~\new_[29472]_ );
  assign \new_[5194]_  = (~\new_[28851]_  | ~\s13_data_i[16] ) & (~\new_[5646]_  | ~\new_[29472]_ );
  assign \new_[5195]_  = ~\new_[5853]_  | ~\new_[5852]_  | ~\new_[5699]_  | ~\new_[5778]_ ;
  assign \new_[5196]_  = ~\s15_data_o[0]  | ~\new_[5681]_ ;
  assign \new_[5197]_  = ~\s15_data_o[10]  | ~\new_[5681]_ ;
  assign \new_[5198]_  = ~\s15_data_o[11]  | ~\new_[5682]_ ;
  assign \new_[5199]_  = ~\s15_data_o[12]  | ~\new_[5681]_ ;
  assign \new_[5200]_  = ~\s15_data_o[13]  | ~\new_[5681]_ ;
  assign \new_[5201]_  = ~\s15_data_o[14]  | ~\new_[5682]_ ;
  assign \new_[5202]_  = ~\s15_data_o[15]  | ~\new_[5682]_ ;
  assign \new_[5203]_  = ~\s15_data_o[1]  | ~\new_[5681]_ ;
  assign \new_[5204]_  = ~\s15_data_o[2]  | ~\new_[5681]_ ;
  assign \new_[5205]_  = ~\s15_data_o[3]  | ~\new_[5681]_ ;
  assign \new_[5206]_  = ~\s15_data_o[4]  | ~\new_[5681]_ ;
  assign \new_[5207]_  = ~\s15_data_o[5]  | ~\new_[5682]_ ;
  assign \new_[5208]_  = ~\s15_data_o[6]  | ~\new_[5682]_ ;
  assign \new_[5209]_  = ~\s15_data_o[7]  | ~\new_[5682]_ ;
  assign \new_[5210]_  = ~\s15_data_o[8]  | ~\new_[5682]_ ;
  assign \new_[5211]_  = ~\s15_data_o[9]  | ~\new_[5682]_ ;
  assign \new_[5212]_  = ~\s15_data_o[0]  | ~\new_[5683]_ ;
  assign \new_[5213]_  = ~\s15_data_o[10]  | ~\new_[5683]_ ;
  assign \new_[5214]_  = ~\s15_data_o[11]  | ~\new_[5683]_ ;
  assign \new_[5215]_  = ~\s15_data_o[12]  | ~\new_[5683]_ ;
  assign \new_[5216]_  = ~\s15_data_o[13]  | ~\new_[5683]_ ;
  assign \new_[5217]_  = ~\s15_data_o[14]  | ~\new_[5683]_ ;
  assign \new_[5218]_  = ~\s15_data_o[15]  | ~\new_[5683]_ ;
  assign \new_[5219]_  = ~\s15_data_o[1]  | ~\new_[5683]_ ;
  assign \new_[5220]_  = ~\s15_data_o[2]  | ~\new_[5683]_ ;
  assign \new_[5221]_  = ~\s15_data_o[3]  | ~\new_[5683]_ ;
  assign \new_[5222]_  = ~\s15_data_o[5]  | ~\new_[5683]_ ;
  assign \new_[5223]_  = ~\s15_data_o[4]  | ~\new_[5683]_ ;
  assign \new_[5224]_  = ~\s15_data_o[6]  | ~\new_[5683]_ ;
  assign \new_[5225]_  = ~\s15_data_o[7]  | ~\new_[5683]_ ;
  assign \new_[5226]_  = ~\s15_data_o[8]  | ~\new_[5683]_ ;
  assign \new_[5227]_  = ~\s15_data_o[9]  | ~\new_[5683]_ ;
  assign \new_[5228]_  = ~\s15_data_o[0]  | ~\new_[5685]_ ;
  assign \new_[5229]_  = ~\s15_data_o[10]  | ~\new_[5685]_ ;
  assign \new_[5230]_  = ~\s15_data_o[11]  | ~\new_[5686]_ ;
  assign \new_[5231]_  = ~\s15_data_o[12]  | ~\new_[5684]_ ;
  assign \new_[5232]_  = ~\s15_data_o[13]  | ~\new_[5686]_ ;
  assign \new_[5233]_  = ~\s15_data_o[14]  | ~\new_[5686]_ ;
  assign \new_[5234]_  = ~\s15_data_o[15]  | ~\new_[5684]_ ;
  assign \new_[5235]_  = ~\s15_data_o[1]  | ~\new_[5684]_ ;
  assign \new_[5236]_  = ~\s15_data_o[2]  | ~\new_[5685]_ ;
  assign \new_[5237]_  = ~\s15_data_o[3]  | ~\new_[5686]_ ;
  assign \new_[5238]_  = ~\s15_data_o[4]  | ~\new_[5686]_ ;
  assign \new_[5239]_  = ~\s15_data_o[5]  | ~\new_[5685]_ ;
  assign \new_[5240]_  = ~\s15_data_o[6]  | ~\new_[5685]_ ;
  assign \new_[5241]_  = ~\s15_data_o[7]  | ~\new_[5685]_ ;
  assign \new_[5242]_  = ~\s15_data_o[8]  | ~\new_[5686]_ ;
  assign \new_[5243]_  = ~\s15_data_o[9]  | ~\new_[5684]_ ;
  assign \new_[5244]_  = ~\s15_data_o[0]  | ~\new_[5687]_ ;
  assign \new_[5245]_  = ~\s15_data_o[10]  | ~\new_[5687]_ ;
  assign \new_[5246]_  = ~\s15_data_o[11]  | ~\new_[5687]_ ;
  assign \new_[5247]_  = ~\s15_data_o[12]  | ~\new_[5687]_ ;
  assign \new_[5248]_  = ~\s15_data_o[13]  | ~\new_[5687]_ ;
  assign \new_[5249]_  = ~\s15_data_o[14]  | ~\new_[5687]_ ;
  assign \new_[5250]_  = ~\s15_data_o[15]  | ~\new_[5687]_ ;
  assign \new_[5251]_  = ~\s15_data_o[1]  | ~\new_[5687]_ ;
  assign \new_[5252]_  = ~\s15_data_o[2]  | ~\new_[5687]_ ;
  assign \new_[5253]_  = ~\s15_data_o[3]  | ~\new_[5687]_ ;
  assign \new_[5254]_  = ~\s15_data_o[4]  | ~\new_[5687]_ ;
  assign \new_[5255]_  = ~\s15_data_o[5]  | ~\new_[5687]_ ;
  assign \new_[5256]_  = ~\s15_data_o[6]  | ~\new_[5687]_ ;
  assign \new_[5257]_  = ~\s15_data_o[7]  | ~\new_[5687]_ ;
  assign \new_[5258]_  = ~\s15_data_o[8]  | ~\new_[5687]_ ;
  assign \new_[5259]_  = ~\s15_data_o[9]  | ~\new_[5687]_ ;
  assign \new_[5260]_  = ~\s15_data_o[0]  | ~\new_[5692]_ ;
  assign \new_[5261]_  = ~\s15_data_o[10]  | ~\new_[5692]_ ;
  assign \new_[5262]_  = ~\s15_data_o[11]  | ~\new_[5692]_ ;
  assign \new_[5263]_  = ~\s15_data_o[12]  | ~\new_[5692]_ ;
  assign \new_[5264]_  = ~\s15_data_o[13]  | ~\new_[5692]_ ;
  assign \new_[5265]_  = ~\s15_data_o[14]  | ~\new_[5692]_ ;
  assign \new_[5266]_  = ~\s15_data_o[15]  | ~\new_[5692]_ ;
  assign \new_[5267]_  = ~\s15_data_o[1]  | ~\new_[5692]_ ;
  assign \new_[5268]_  = ~\s15_data_o[2]  | ~\new_[5692]_ ;
  assign \new_[5269]_  = ~\s15_data_o[3]  | ~\new_[5692]_ ;
  assign \new_[5270]_  = ~\s15_data_o[4]  | ~\new_[5692]_ ;
  assign \new_[5271]_  = ~\s15_data_o[5]  | ~\new_[5692]_ ;
  assign \new_[5272]_  = ~\s15_data_o[6]  | ~\new_[5692]_ ;
  assign \new_[5273]_  = ~\s15_data_o[7]  | ~\new_[5692]_ ;
  assign \new_[5274]_  = ~\s15_data_o[8]  | ~\new_[5692]_ ;
  assign \new_[5275]_  = ~\s15_data_o[9]  | ~\new_[5692]_ ;
  assign \new_[5276]_  = ~\s15_data_o[0]  | ~\new_[5679]_ ;
  assign \new_[5277]_  = ~\s15_data_o[10]  | ~\new_[5679]_ ;
  assign \new_[5278]_  = ~\s15_data_o[11]  | ~\new_[5679]_ ;
  assign \new_[5279]_  = ~\s15_data_o[12]  | ~\new_[5679]_ ;
  assign \new_[5280]_  = ~\s15_data_o[13]  | ~\new_[5679]_ ;
  assign \new_[5281]_  = ~\s15_data_o[14]  | ~\new_[5679]_ ;
  assign \new_[5282]_  = ~\s15_data_o[15]  | ~\new_[5679]_ ;
  assign \new_[5283]_  = ~\s15_data_o[1]  | ~\new_[5679]_ ;
  assign \new_[5284]_  = ~\s15_data_o[2]  | ~\new_[5679]_ ;
  assign \new_[5285]_  = ~\s15_data_o[3]  | ~\new_[5679]_ ;
  assign \new_[5286]_  = ~\s15_data_o[4]  | ~\new_[5679]_ ;
  assign \new_[5287]_  = ~\s15_data_o[5]  | ~\new_[5679]_ ;
  assign \new_[5288]_  = ~\s15_data_o[6]  | ~\new_[5679]_ ;
  assign \new_[5289]_  = ~\s15_data_o[7]  | ~\new_[5679]_ ;
  assign \new_[5290]_  = ~\s15_data_o[8]  | ~\new_[5679]_ ;
  assign \new_[5291]_  = ~\s15_data_o[9]  | ~\new_[5679]_ ;
  assign \new_[5292]_  = ~\new_[5680]_  | ~\new_[4200]_ ;
  assign \new_[5293]_  = ~\new_[5680]_  | ~\new_[4201]_ ;
  assign \new_[5294]_  = ~\new_[5680]_  | ~\new_[4202]_ ;
  assign \new_[5295]_  = ~\new_[5680]_  | ~\new_[4203]_ ;
  assign \new_[5296]_  = ~\new_[5680]_  | ~\new_[4204]_ ;
  assign \new_[5297]_  = ~\new_[5680]_  | ~\new_[4205]_ ;
  assign \new_[5298]_  = ~\new_[5680]_  | ~\new_[4206]_ ;
  assign \new_[5299]_  = ~\new_[5680]_  | ~\new_[4207]_ ;
  assign \new_[5300]_  = ~\new_[5680]_  | ~\new_[4208]_ ;
  assign \new_[5301]_  = ~\new_[5680]_  | ~\new_[4209]_ ;
  assign \new_[5302]_  = ~\new_[5680]_  | ~\new_[4210]_ ;
  assign \new_[5303]_  = ~\new_[5680]_  | ~\new_[4211]_ ;
  assign \new_[5304]_  = ~\new_[5680]_  | ~\new_[4212]_ ;
  assign \new_[5305]_  = ~\new_[5680]_  | ~\new_[4213]_ ;
  assign \new_[5306]_  = ~\new_[5680]_  | ~\new_[4214]_ ;
  assign \new_[5307]_  = ~\new_[5680]_  | ~\new_[4215]_ ;
  assign \new_[5308]_  = ~\s15_data_o[0]  | ~\new_[5689]_ ;
  assign \new_[5309]_  = ~\s15_data_o[10]  | ~\new_[5689]_ ;
  assign \new_[5310]_  = ~\s15_data_o[11]  | ~\new_[5689]_ ;
  assign \new_[5311]_  = ~\s15_data_o[12]  | ~\new_[5689]_ ;
  assign \new_[5312]_  = ~\s15_data_o[13]  | ~\new_[5689]_ ;
  assign \new_[5313]_  = ~\s15_data_o[14]  | ~\new_[5689]_ ;
  assign \new_[5314]_  = ~\s15_data_o[15]  | ~\new_[5689]_ ;
  assign \new_[5315]_  = ~\s15_data_o[1]  | ~\new_[5689]_ ;
  assign \new_[5316]_  = ~\s15_data_o[2]  | ~\new_[5689]_ ;
  assign \new_[5317]_  = ~\s15_data_o[3]  | ~\new_[5689]_ ;
  assign \new_[5318]_  = ~\s15_data_o[4]  | ~\new_[5689]_ ;
  assign \new_[5319]_  = ~\s15_data_o[5]  | ~\new_[5689]_ ;
  assign \new_[5320]_  = ~\s15_data_o[6]  | ~\new_[5689]_ ;
  assign \new_[5321]_  = ~\s15_data_o[7]  | ~\new_[5689]_ ;
  assign \new_[5322]_  = ~\s15_data_o[8]  | ~\new_[5689]_ ;
  assign \new_[5323]_  = ~\s15_data_o[9]  | ~\new_[5689]_ ;
  assign \new_[5324]_  = ~\s15_data_o[0]  | ~\new_[5690]_ ;
  assign \new_[5325]_  = ~\s15_data_o[10]  | ~\new_[5690]_ ;
  assign \new_[5326]_  = ~\s15_data_o[11]  | ~\new_[5690]_ ;
  assign \new_[5327]_  = ~\s15_data_o[12]  | ~\new_[5690]_ ;
  assign \new_[5328]_  = ~\s15_data_o[13]  | ~\new_[5690]_ ;
  assign \new_[5329]_  = ~\s15_data_o[14]  | ~\new_[5690]_ ;
  assign \new_[5330]_  = ~\s15_data_o[15]  | ~\new_[5690]_ ;
  assign \new_[5331]_  = ~\s15_data_o[1]  | ~\new_[5690]_ ;
  assign \new_[5332]_  = ~\s15_data_o[2]  | ~\new_[5690]_ ;
  assign \new_[5333]_  = ~\s15_data_o[3]  | ~\new_[5690]_ ;
  assign \new_[5334]_  = ~\s15_data_o[4]  | ~\new_[5690]_ ;
  assign \new_[5335]_  = ~\s15_data_o[5]  | ~\new_[5690]_ ;
  assign \new_[5336]_  = ~\s15_data_o[6]  | ~\new_[5690]_ ;
  assign \new_[5337]_  = ~\s15_data_o[7]  | ~\new_[5690]_ ;
  assign \new_[5338]_  = ~\s15_data_o[8]  | ~\new_[5690]_ ;
  assign \new_[5339]_  = ~\s15_data_o[9]  | ~\new_[5690]_ ;
  assign \new_[5340]_  = ~\s15_data_o[0]  | ~\new_[5691]_ ;
  assign \new_[5341]_  = ~\s15_data_o[10]  | ~\new_[5691]_ ;
  assign \new_[5342]_  = ~\s15_data_o[11]  | ~\new_[5691]_ ;
  assign \new_[5343]_  = ~\s15_data_o[12]  | ~\new_[5691]_ ;
  assign \new_[5344]_  = ~\s15_data_o[13]  | ~\new_[5691]_ ;
  assign \new_[5345]_  = ~\s15_data_o[14]  | ~\new_[5691]_ ;
  assign \new_[5346]_  = ~\s15_data_o[15]  | ~\new_[5691]_ ;
  assign \new_[5347]_  = ~\s15_data_o[1]  | ~\new_[5691]_ ;
  assign \new_[5348]_  = ~\s15_data_o[2]  | ~\new_[5691]_ ;
  assign \new_[5349]_  = ~\s15_data_o[3]  | ~\new_[5691]_ ;
  assign \new_[5350]_  = ~\s15_data_o[4]  | ~\new_[5691]_ ;
  assign \new_[5351]_  = ~\s15_data_o[5]  | ~\new_[5691]_ ;
  assign \new_[5352]_  = ~\s15_data_o[6]  | ~\new_[5691]_ ;
  assign \new_[5353]_  = ~\s15_data_o[7]  | ~\new_[5691]_ ;
  assign \new_[5354]_  = ~\s15_data_o[8]  | ~\new_[5691]_ ;
  assign \new_[5355]_  = ~\s15_data_o[9]  | ~\new_[5691]_ ;
  assign \new_[5356]_  = ~\new_[5674]_  | ~\new_[4233]_ ;
  assign \new_[5357]_  = ~\new_[5674]_  | ~\new_[4234]_ ;
  assign \new_[5358]_  = ~\new_[5674]_  | ~\new_[4235]_ ;
  assign \new_[5359]_  = ~\new_[5674]_  | ~\new_[4236]_ ;
  assign \new_[5360]_  = ~\new_[5674]_  | ~\new_[4237]_ ;
  assign \new_[5361]_  = ~\new_[5674]_  | ~\new_[4238]_ ;
  assign \new_[5362]_  = ~\new_[5674]_  | ~\new_[4239]_ ;
  assign \new_[5363]_  = ~\new_[5674]_  | ~\new_[4240]_ ;
  assign \new_[5364]_  = ~\new_[5674]_  | ~\new_[4247]_ ;
  assign \new_[5365]_  = ~\new_[5674]_  | ~\new_[4248]_ ;
  assign \new_[5366]_  = ~\new_[5674]_  | ~\new_[4241]_ ;
  assign \new_[5367]_  = ~\new_[5674]_  | ~\new_[4242]_ ;
  assign \new_[5368]_  = ~\new_[5674]_  | ~\new_[4243]_ ;
  assign \new_[5369]_  = ~\new_[5674]_  | ~\new_[4244]_ ;
  assign \new_[5370]_  = ~\new_[5674]_  | ~\new_[4245]_ ;
  assign \new_[5371]_  = ~\new_[5674]_  | ~\new_[4246]_ ;
  assign \new_[5372]_  = ~\new_[5693]_  | ~\new_[4249]_ ;
  assign \new_[5373]_  = ~\new_[5848]_  | ~\new_[4250]_ ;
  assign \new_[5374]_  = ~\new_[5693]_  | ~\new_[4251]_ ;
  assign \new_[5375]_  = ~\new_[5848]_  | ~\new_[4252]_ ;
  assign \new_[5376]_  = ~\new_[5693]_  | ~\new_[4253]_ ;
  assign \new_[5377]_  = ~\new_[5848]_  | ~\new_[4254]_ ;
  assign \new_[5378]_  = ~\new_[5693]_  | ~\new_[4255]_ ;
  assign \new_[5379]_  = ~\new_[5693]_  | ~\new_[4256]_ ;
  assign \new_[5380]_  = ~\new_[5848]_  | ~\new_[4263]_ ;
  assign \new_[5381]_  = ~\new_[5693]_  | ~\new_[4264]_ ;
  assign \new_[5382]_  = ~\new_[5693]_  | ~\new_[4257]_ ;
  assign \new_[5383]_  = ~\new_[5693]_  | ~\new_[4258]_ ;
  assign \new_[5384]_  = ~\new_[5693]_  | ~\new_[4259]_ ;
  assign \new_[5385]_  = ~\new_[5693]_  | ~\new_[4260]_ ;
  assign \new_[5386]_  = ~\new_[5693]_  | ~\new_[4261]_ ;
  assign \new_[5387]_  = ~\new_[5693]_  | ~\new_[4262]_ ;
  assign \new_[5388]_  = ~\new_[5694]_  | ~\new_[4166]_ ;
  assign \new_[5389]_  = ~\new_[5694]_  | ~\new_[4167]_ ;
  assign \new_[5390]_  = ~\new_[5694]_  | ~\new_[4168]_ ;
  assign \new_[5391]_  = ~\new_[5694]_  | ~\new_[4169]_ ;
  assign \new_[5392]_  = ~\new_[5694]_  | ~\new_[4170]_ ;
  assign \new_[5393]_  = ~\new_[5694]_  | ~\new_[4171]_ ;
  assign \new_[5394]_  = ~\new_[5694]_  | ~\new_[4172]_ ;
  assign \new_[5395]_  = ~\new_[5694]_  | ~\new_[4173]_ ;
  assign \new_[5396]_  = ~\new_[5694]_  | ~\new_[4174]_ ;
  assign \new_[5397]_  = ~\new_[5694]_  | ~\new_[4175]_ ;
  assign \new_[5398]_  = ~\new_[5694]_  | ~\new_[4176]_ ;
  assign \new_[5399]_  = ~\new_[5694]_  | ~\new_[4177]_ ;
  assign \new_[5400]_  = ~\new_[5694]_  | ~\new_[4178]_ ;
  assign \new_[5401]_  = ~\new_[5694]_  | ~\new_[4179]_ ;
  assign \new_[5402]_  = ~\new_[5694]_  | ~\new_[4180]_ ;
  assign \new_[5403]_  = ~\new_[5694]_  | ~\new_[4181]_ ;
  assign \new_[5404]_  = ~\new_[5696]_  | ~\new_[4265]_ ;
  assign \new_[5405]_  = ~\new_[5849]_  | ~\new_[4266]_ ;
  assign \new_[5406]_  = ~\new_[5696]_  | ~\new_[4267]_ ;
  assign \new_[5407]_  = ~\new_[5849]_  | ~\new_[4268]_ ;
  assign \new_[5408]_  = ~\new_[5696]_  | ~\new_[4269]_ ;
  assign \new_[5409]_  = ~\new_[5849]_  | ~\new_[4270]_ ;
  assign \new_[5410]_  = ~\new_[5696]_  | ~\new_[4271]_ ;
  assign \new_[5411]_  = ~\new_[5696]_  | ~\new_[4272]_ ;
  assign \new_[5412]_  = ~\new_[5849]_  | ~\new_[4273]_ ;
  assign \new_[5413]_  = ~\new_[5696]_  | ~\new_[4274]_ ;
  assign \new_[5414]_  = ~\new_[5696]_  | ~\new_[4275]_ ;
  assign \new_[5415]_  = ~\new_[5696]_  | ~\new_[4276]_ ;
  assign \new_[5416]_  = ~\new_[5696]_  | ~\new_[4277]_ ;
  assign \new_[5417]_  = ~\new_[5696]_  | ~\new_[4278]_ ;
  assign \new_[5418]_  = ~\new_[5696]_  | ~\new_[4279]_ ;
  assign \new_[5419]_  = ~\new_[5696]_  | ~\new_[4280]_ ;
  assign \new_[5420]_  = ~\new_[5675]_  & (~\new_[5953]_  | ~\new_[4117]_ );
  assign \new_[5421]_  = ~\new_[5697]_  & (~\new_[32068]_  | ~\new_[4149]_ );
  assign \new_[5422]_  = ~\new_[5698]_  & (~\new_[5960]_  | ~\new_[4249]_ );
  assign \new_[5423]_  = ~\new_[5700]_  & (~\new_[5960]_  | ~\new_[4250]_ );
  assign \new_[5424]_  = ~\new_[5702]_  | ~\new_[5856]_ ;
  assign \new_[5425]_  = ~\new_[5703]_  | (~\new_[5885]_  & ~\new_[31446]_ );
  assign \new_[5426]_  = ~\new_[5704]_  | (~\new_[5885]_  & ~\new_[31734]_ );
  assign \new_[5427]_  = ~\new_[32170]_  & (~\new_[32068]_  | ~\new_[4152]_ );
  assign \new_[5428]_  = ~\new_[5558]_ ;
  assign \new_[5429]_  = ~\new_[5706]_  | (~\new_[5885]_  & ~\new_[31642]_ );
  assign \new_[5430]_  = ~\new_[5707]_  & (~\new_[5960]_  | ~\new_[4255]_ );
  assign \new_[5431]_  = ~\new_[5710]_  | (~\new_[5885]_  & ~\new_[31823]_ );
  assign \new_[5432]_  = ~\new_[5711]_  & (~\new_[32192]_  | ~\new_[4089]_ );
  assign \new_[5433]_  = ~\new_[5573]_ ;
  assign \new_[5434]_  = ~\new_[5712]_  | ~\new_[5804]_ ;
  assign \new_[5435]_  = ~\new_[5713]_  | ~\new_[5807]_ ;
  assign \new_[5436]_  = ~\new_[5714]_  & (~\new_[6029]_  | ~\new_[4264]_ );
  assign \new_[5437]_  = ~\new_[5715]_  | (~\new_[5885]_  & ~\new_[31786]_ );
  assign \new_[5438]_  = ~\new_[5676]_  & (~\new_[6017]_  | ~\new_[4241]_ );
  assign \new_[5439]_  = ~\new_[5585]_ ;
  assign \new_[5440]_  = ~\new_[5716]_  | (~\new_[5885]_  & ~\new_[31792]_ );
  assign \new_[5441]_  = ~\new_[5677]_  & (~\new_[6017]_  | ~\new_[4242]_ );
  assign \new_[5442]_  = ~\new_[5590]_ ;
  assign \new_[5443]_  = ~\new_[5718]_  & (~\new_[32068]_  | ~\new_[4162]_ );
  assign \new_[5444]_  = ~\new_[5595]_ ;
  assign \new_[5445]_  = ~\new_[5719]_  & (~\new_[6029]_  | ~\new_[4260]_ );
  assign \new_[5446]_  = ~\new_[5720]_  & (~\new_[6029]_  | ~\new_[4261]_ );
  assign \new_[5447]_  = ~\new_[5721]_  | (~\new_[5885]_  & ~\new_[31802]_ );
  assign \new_[5448]_  = ~\new_[5678]_  & (~\new_[6017]_  | ~\new_[4246]_ );
  assign \new_[5449]_  = ~\new_[5607]_ ;
  assign \new_[5450]_  = ~\new_[5629]_ ;
  assign \new_[5451]_  = \new_[31781]_  ? \new_[5880]_  : s15_ack_i;
  assign \new_[5452]_  = ~\s15_data_o[0]  | ~\new_[5763]_ ;
  assign \new_[5453]_  = ~\s15_data_o[10]  | ~\new_[5763]_ ;
  assign \new_[5454]_  = ~\s15_data_o[11]  | ~\new_[5763]_ ;
  assign \new_[5455]_  = ~\s15_data_o[12]  | ~\new_[5763]_ ;
  assign \new_[5456]_  = ~\s15_data_o[13]  | ~\new_[5763]_ ;
  assign \new_[5457]_  = ~\s15_data_o[14]  | ~\new_[5763]_ ;
  assign \new_[5458]_  = ~\s15_data_o[15]  | ~\new_[5763]_ ;
  assign \new_[5459]_  = ~\s15_data_o[1]  | ~\new_[5763]_ ;
  assign \new_[5460]_  = ~\s15_data_o[2]  | ~\new_[5763]_ ;
  assign \new_[5461]_  = ~\s15_data_o[3]  | ~\new_[5763]_ ;
  assign \new_[5462]_  = ~\s15_data_o[4]  | ~\new_[5763]_ ;
  assign \new_[5463]_  = ~\s15_data_o[5]  | ~\new_[5763]_ ;
  assign \new_[5464]_  = ~\s15_data_o[6]  | ~\new_[5763]_ ;
  assign \new_[5465]_  = ~\s15_data_o[7]  | ~\new_[5763]_ ;
  assign \new_[5466]_  = ~\s15_data_o[9]  | ~\new_[5763]_ ;
  assign \new_[5467]_  = ~\s15_data_o[8]  | ~\new_[5763]_ ;
  assign \new_[5468]_  = ~\s15_data_o[0]  | ~\new_[5722]_ ;
  assign \new_[5469]_  = ~\s15_data_o[10]  | ~\new_[5722]_ ;
  assign \new_[5470]_  = ~\s15_data_o[11]  | ~\new_[5722]_ ;
  assign \new_[5471]_  = ~\s15_data_o[12]  | ~\new_[5722]_ ;
  assign \new_[5472]_  = ~\s15_data_o[13]  | ~\new_[5722]_ ;
  assign \new_[5473]_  = ~\s15_data_o[14]  | ~\new_[5722]_ ;
  assign \new_[5474]_  = ~\s15_data_o[15]  | ~\new_[5722]_ ;
  assign \new_[5475]_  = ~\s15_data_o[1]  | ~\new_[5722]_ ;
  assign \new_[5476]_  = ~\s15_data_o[2]  | ~\new_[5722]_ ;
  assign \new_[5477]_  = ~\s15_data_o[3]  | ~\new_[5722]_ ;
  assign \new_[5478]_  = ~\s15_data_o[4]  | ~\new_[5722]_ ;
  assign \new_[5479]_  = ~\s15_data_o[5]  | ~\new_[5722]_ ;
  assign \new_[5480]_  = ~\s15_data_o[6]  | ~\new_[5722]_ ;
  assign \new_[5481]_  = ~\s15_data_o[7]  | ~\new_[5722]_ ;
  assign \new_[5482]_  = ~\s15_data_o[8]  | ~\new_[5722]_ ;
  assign \new_[5483]_  = ~\s15_data_o[9]  | ~\new_[5722]_ ;
  assign \new_[5484]_  = ~\s15_data_o[0]  | ~\new_[5773]_ ;
  assign \new_[5485]_  = ~\s15_data_o[10]  | ~\new_[5773]_ ;
  assign \new_[5486]_  = ~\s15_data_o[11]  | ~\new_[5774]_ ;
  assign \new_[5487]_  = ~\s15_data_o[12]  | ~\new_[5772]_ ;
  assign \new_[5488]_  = ~\s15_data_o[13]  | ~\new_[5774]_ ;
  assign \new_[5489]_  = ~\s15_data_o[14]  | ~\new_[5774]_ ;
  assign \new_[5490]_  = ~\s15_data_o[15]  | ~\new_[5772]_ ;
  assign \new_[5491]_  = ~\s15_data_o[1]  | ~\new_[5772]_ ;
  assign \new_[5492]_  = ~\s15_data_o[2]  | ~\new_[5773]_ ;
  assign \new_[5493]_  = ~\s15_data_o[3]  | ~\new_[5774]_ ;
  assign \new_[5494]_  = ~\s15_data_o[4]  | ~\new_[5774]_ ;
  assign \new_[5495]_  = ~\s15_data_o[5]  | ~\new_[5773]_ ;
  assign \new_[5496]_  = ~\s15_data_o[6]  | ~\new_[5773]_ ;
  assign \new_[5497]_  = ~\s15_data_o[7]  | ~\new_[5773]_ ;
  assign \new_[5498]_  = ~\s15_data_o[8]  | ~\new_[5774]_ ;
  assign \new_[5499]_  = ~\s15_data_o[9]  | ~\new_[5772]_ ;
  assign \new_[5500]_  = ~\s15_data_o[0]  | ~\new_[5776]_ ;
  assign \new_[5501]_  = ~\s15_data_o[10]  | ~\new_[5776]_ ;
  assign \new_[5502]_  = ~\s15_data_o[11]  | ~\new_[5776]_ ;
  assign \new_[5503]_  = ~\s15_data_o[12]  | ~\new_[5776]_ ;
  assign \new_[5504]_  = ~\s15_data_o[13]  | ~\new_[5776]_ ;
  assign \new_[5505]_  = ~\s15_data_o[14]  | ~\new_[5776]_ ;
  assign \new_[5506]_  = ~\s15_data_o[15]  | ~\new_[5776]_ ;
  assign \new_[5507]_  = ~\s15_data_o[1]  | ~\new_[5776]_ ;
  assign \new_[5508]_  = ~\s15_data_o[2]  | ~\new_[5776]_ ;
  assign \new_[5509]_  = ~\s15_data_o[3]  | ~\new_[5776]_ ;
  assign \new_[5510]_  = ~\s15_data_o[4]  | ~\new_[5776]_ ;
  assign \new_[5511]_  = ~\s15_data_o[5]  | ~\new_[5776]_ ;
  assign \new_[5512]_  = ~\s15_data_o[6]  | ~\new_[5776]_ ;
  assign \new_[5513]_  = ~\s15_data_o[7]  | ~\new_[5776]_ ;
  assign \new_[5514]_  = ~\s15_data_o[8]  | ~\new_[5776]_ ;
  assign \new_[5515]_  = ~\s15_data_o[9]  | ~\new_[5776]_ ;
  assign \new_[5516]_  = ~\new_[5764]_  | ~\new_[4216]_ ;
  assign \new_[5517]_  = ~\new_[5764]_  | ~\new_[4218]_ ;
  assign \new_[5518]_  = ~\new_[5764]_  | ~\new_[4217]_ ;
  assign \new_[5519]_  = ~\new_[5764]_  | ~\new_[4219]_ ;
  assign \new_[5520]_  = ~\new_[5764]_  | ~\new_[4220]_ ;
  assign \new_[5521]_  = ~\new_[5764]_  | ~\new_[4221]_ ;
  assign \new_[5522]_  = ~\new_[5764]_  | ~\new_[4222]_ ;
  assign \new_[5523]_  = ~\new_[5764]_  | ~\new_[4223]_ ;
  assign \new_[5524]_  = ~\new_[5764]_  | ~\new_[4230]_ ;
  assign \new_[5525]_  = ~\new_[5764]_  | ~\new_[4231]_ ;
  assign \new_[5526]_  = ~\new_[5764]_  | ~\new_[4224]_ ;
  assign \new_[5527]_  = ~\new_[5764]_  | ~\new_[4225]_ ;
  assign \new_[5528]_  = ~\new_[5764]_  | ~\new_[4226]_ ;
  assign \new_[5529]_  = ~\new_[5764]_  | ~\new_[4227]_ ;
  assign \new_[5530]_  = ~\new_[5764]_  | ~\new_[4228]_ ;
  assign \new_[5531]_  = ~\new_[5764]_  | ~\new_[4229]_ ;
  assign \new_[5532]_  = ~\new_[5723]_  | ~\new_[4438]_ ;
  assign \new_[5533]_  = ~\new_[5723]_  | ~\new_[4439]_ ;
  assign \new_[5534]_  = ~\new_[5723]_  | ~\new_[4440]_ ;
  assign \new_[5535]_  = ~\new_[5723]_  | ~\new_[4441]_ ;
  assign \new_[5536]_  = ~\new_[5723]_  | ~\new_[4442]_ ;
  assign \new_[5537]_  = ~\new_[5723]_  | ~\new_[4443]_ ;
  assign \new_[5538]_  = ~\new_[5723]_  | ~\new_[4444]_ ;
  assign \new_[5539]_  = ~\new_[5723]_  | ~\new_[4445]_ ;
  assign \new_[5540]_  = ~\new_[5723]_  | ~\new_[4452]_ ;
  assign \new_[5541]_  = ~\new_[5723]_  | ~\new_[4446]_ ;
  assign \new_[5542]_  = ~\new_[5723]_  | ~\new_[4453]_ ;
  assign \new_[5543]_  = ~\new_[5723]_  | ~\new_[4447]_ ;
  assign \new_[5544]_  = ~\new_[5723]_  | ~\new_[4448]_ ;
  assign \new_[5545]_  = ~\new_[5723]_  | ~\new_[4449]_ ;
  assign \new_[5546]_  = ~\new_[5723]_  | ~\new_[4450]_ ;
  assign \new_[5547]_  = ~\new_[5723]_  | ~\new_[4451]_ ;
  assign \new_[5548]_  = ~\new_[5777]_  | ~\new_[5851]_ ;
  assign \new_[5549]_  = ~\new_[5779]_  | ~\new_[5780]_ ;
  assign \new_[5550]_  = ~\new_[5781]_  | ~\new_[5855]_ ;
  assign \new_[5551]_  = ~\new_[5724]_  | ~\new_[5725]_ ;
  assign \new_[5552]_  = ~\new_[5783]_  | (~\new_[32316]_  & ~\new_[31299]_ );
  assign \new_[5553]_  = ~\new_[5836]_  | (~\new_[5892]_  & ~\new_[31702]_ );
  assign \new_[5554]_  = ~\new_[5784]_  & (~\new_[5889]_  | ~\new_[4440]_ );
  assign \new_[5555]_  = ~\new_[5786]_  | (~\new_[5958]_  & ~\new_[31805]_ );
  assign \new_[5556]_  = ~\new_[5838]_  | (~\new_[5892]_  & ~\new_[31912]_ );
  assign \new_[5557]_  = ~\new_[5787]_  & (~\new_[5943]_  | ~\new_[4085]_ );
  assign \new_[5558]_  = ~\new_[5729]_  | ~\new_[5730]_ ;
  assign \new_[5559]_  = ~\new_[5789]_  | ~\new_[5788]_ ;
  assign \new_[5560]_  = ~\new_[5790]_  | ~\new_[5863]_ ;
  assign \new_[5561]_  = ~\new_[5731]_  | ~\new_[5732]_ ;
  assign \new_[5562]_  = ~\new_[5791]_  & (~\new_[6026]_  | ~\new_[4204]_ );
  assign \new_[5563]_  = ~\new_[5795]_  | (~\new_[32316]_  & ~\new_[31762]_ );
  assign \new_[5564]_  = ~\new_[5733]_  & (~\new_[6017]_  | ~\new_[4238]_ );
  assign \new_[5565]_  = ~\new_[5796]_  & (~\new_[6026]_  | ~\new_[4205]_ );
  assign \new_[5566]_  = ~\new_[5797]_  & (~\new_[5889]_  | ~\new_[4443]_ );
  assign \new_[5567]_  = ~\new_[5798]_  | ~\new_[5799]_ ;
  assign \new_[5568]_  = ~\new_[5800]_  | ~\new_[5865]_ ;
  assign \new_[5569]_  = ~\new_[5736]_  | ~\new_[5737]_ ;
  assign \new_[5570]_  = ~\new_[5739]_  | (~\new_[5945]_  & ~\new_[31916]_ );
  assign \new_[5571]_  = ~\new_[5801]_  | (~\new_[5958]_  & ~\new_[31649]_ );
  assign \new_[5572]_  = ~\new_[5802]_  & (~\new_[5889]_  | ~\new_[4445]_ );
  assign \new_[5573]_  = ~\new_[5740]_  | ~\new_[5741]_ ;
  assign \new_[5574]_  = ~\new_[5803]_  & (~\new_[6027]_  | ~\new_[4156]_ );
  assign \new_[5575]_  = ~\new_[5742]_  | ~\new_[5843]_ ;
  assign \new_[5576]_  = ~\new_[5869]_  | ~\new_[5805]_ ;
  assign \new_[5577]_  = ~\new_[5806]_  & (~\new_[6027]_  | ~\new_[4157]_ );
  assign \new_[5578]_  = ~\new_[5808]_  | (~\new_[5957]_  & ~\new_[31774]_ );
  assign \new_[5579]_  = ~\new_[5809]_  | (~\new_[5942]_  & ~\new_[31731]_ );
  assign \new_[5580]_  = ~\new_[5745]_  | ~\new_[5746]_ ;
  assign \new_[5581]_  = ~\new_[5747]_  & (~\new_[6187]_  | ~\new_[4248]_ );
  assign \new_[5582]_  = ~\new_[5810]_  & (~\new_[6026]_  | ~\new_[4209]_ );
  assign \new_[5583]_  = ~\new_[5811]_  | (~\new_[5959]_  & ~\new_[31701]_ );
  assign \new_[5584]_  = ~\new_[5812]_  & (~\new_[6025]_  | ~\new_[4210]_ );
  assign \new_[5585]_  = ~\new_[5748]_  | ~\new_[5749]_ ;
  assign \new_[5586]_  = ~\new_[5813]_  & (~\new_[5943]_  | ~\new_[4091]_ );
  assign \new_[5587]_  = ~\new_[5814]_  | (~\new_[5959]_  & ~\new_[31748]_ );
  assign \new_[5588]_  = ~\new_[5815]_  & (~\new_[6025]_  | ~\new_[4211]_ );
  assign \new_[5589]_  = ~\new_[5816]_  & (~\new_[6027]_  | ~\new_[4160]_ );
  assign \new_[5590]_  = ~\new_[5750]_  | ~\new_[5751]_ ;
  assign \new_[5591]_  = ~\new_[5817]_  & (~\new_[5943]_  | ~\new_[4092]_ );
  assign \new_[5592]_  = ~\new_[5818]_  | (~\new_[5958]_  & ~\new_[31879]_ );
  assign \new_[5593]_  = ~\new_[5845]_  | (~\new_[5892]_  & ~\new_[31663]_ );
  assign \new_[5594]_  = ~\new_[5820]_  | (~\new_[5942]_  & ~\new_[31657]_ );
  assign \new_[5595]_  = ~\new_[5754]_  | ~\new_[5755]_ ;
  assign \new_[5596]_  = ~\new_[5821]_  & (~\new_[6026]_  | ~\new_[4213]_ );
  assign \new_[5597]_  = ~\new_[5756]_  & (~\new_[6187]_  | ~\new_[4244]_ );
  assign \new_[5598]_  = ~\new_[5822]_  | (~\new_[5942]_  & ~\new_[31926]_ );
  assign \new_[5599]_  = ~\new_[5823]_  | (~\new_[5957]_  & ~\new_[31630]_ );
  assign \new_[5600]_  = ~\new_[5757]_  | ~\new_[5759]_ ;
  assign \new_[5601]_  = ~\new_[5758]_  & (~\new_[6187]_  | ~\new_[4245]_ );
  assign \new_[5602]_  = ~\new_[5824]_  & (~\new_[6026]_  | ~\new_[4214]_ );
  assign \new_[5603]_  = ~\new_[5825]_  | (~\new_[32316]_  & ~\new_[31754]_ );
  assign \new_[5604]_  = ~\new_[5826]_  & (~\new_[6025]_  | ~\new_[4215]_ );
  assign \new_[5605]_  = ~\new_[5827]_  & (~\new_[5943]_  | ~\new_[4096]_ );
  assign \new_[5606]_  = ~\new_[5828]_  & (~\new_[6027]_  | ~\new_[4164]_ );
  assign \new_[5607]_  = ~\new_[5760]_  | ~\new_[5761]_ ;
  assign \new_[5608]_  = ~\new_[5954]_  | ~\new_[4036]_ ;
  assign \new_[5609]_  = ~\new_[5954]_  | ~\new_[4040]_ ;
  assign \new_[5610]_  = ~\new_[5679]_ ;
  assign \new_[5611]_  = ~\new_[5683]_ ;
  assign \new_[5612]_  = ~\new_[5683]_ ;
  assign \new_[5613]_  = ~\new_[5683]_ ;
  assign \new_[5614]_  = ~\new_[5684]_ ;
  assign \new_[5615]_  = ~\new_[5687]_ ;
  assign \new_[5616]_  = ~\new_[5687]_ ;
  assign \new_[5617]_  = ~\new_[5687]_ ;
  assign \new_[5618]_  = \new_[5688]_ ;
  assign \new_[5619]_  = ~\new_[5688]_ ;
  assign \new_[5620]_  = ~\new_[5689]_ ;
  assign \new_[5621]_  = ~\new_[5690]_ ;
  assign \new_[5622]_  = ~\new_[5691]_ ;
  assign \new_[5623]_  = ~\new_[5692]_ ;
  assign \new_[5624]_  = \new_[5695]_ ;
  assign \new_[5625]_  = ~\new_[5941]_  | ~\new_[4074]_ ;
  assign \new_[5626]_  = ~\new_[5829]_  & ~\new_[31896]_ ;
  assign \new_[5627]_  = ~\new_[5829]_  & ~\new_[31613]_ ;
  assign \new_[5628]_  = ~\new_[5829]_  & ~\new_[31606]_ ;
  assign \new_[5629]_  = \new_[32274]_ ;
  assign \new_[5630]_  = ~\s15_data_o[0]  | ~\new_[5832]_ ;
  assign \new_[5631]_  = ~\s15_data_o[10]  | ~\new_[5832]_ ;
  assign \new_[5632]_  = ~\s15_data_o[11]  | ~\new_[5832]_ ;
  assign \new_[5633]_  = ~\s15_data_o[12]  | ~\new_[5832]_ ;
  assign \new_[5634]_  = ~\s15_data_o[13]  | ~\new_[5832]_ ;
  assign \new_[5635]_  = ~\s15_data_o[14]  | ~\new_[5832]_ ;
  assign \new_[5636]_  = ~\s15_data_o[15]  | ~\new_[5832]_ ;
  assign \new_[5637]_  = ~\s15_data_o[1]  | ~\new_[5832]_ ;
  assign \new_[5638]_  = ~\s15_data_o[2]  | ~\new_[5832]_ ;
  assign \new_[5639]_  = ~\s15_data_o[3]  | ~\new_[5832]_ ;
  assign \new_[5640]_  = ~\s15_data_o[4]  | ~\new_[5832]_ ;
  assign \new_[5641]_  = ~\s15_data_o[5]  | ~\new_[5832]_ ;
  assign \new_[5642]_  = ~\s15_data_o[6]  | ~\new_[5832]_ ;
  assign \new_[5643]_  = ~\s15_data_o[7]  | ~\new_[5832]_ ;
  assign \new_[5644]_  = ~\s15_data_o[8]  | ~\new_[5832]_ ;
  assign \new_[5645]_  = ~\s15_data_o[9]  | ~\new_[5832]_ ;
  assign \new_[5646]_  = \new_[32278]_  & \s15_data_i[16] ;
  assign \new_[5647]_  = \new_[32340]_  & \s15_data_i[26] ;
  assign \new_[5648]_  = \new_[32340]_  & \s15_data_i[25] ;
  assign \new_[5649]_  = \new_[32340]_  & \s15_data_i[24] ;
  assign \new_[5650]_  = \new_[32340]_  & \s15_data_i[23] ;
  assign \new_[5651]_  = \new_[32278]_  & \s15_data_i[30] ;
  assign \new_[5652]_  = \new_[32278]_  & \s15_data_i[22] ;
  assign \new_[5653]_  = \new_[32340]_  & \s15_data_i[21] ;
  assign \new_[5654]_  = \new_[32340]_  & \s15_data_i[20] ;
  assign \new_[5655]_  = \new_[32340]_  & \s15_data_i[19] ;
  assign \new_[5656]_  = \new_[32278]_  & \s15_data_i[18] ;
  assign \new_[5657]_  = \new_[32278]_  & \s15_data_i[17] ;
  assign \new_[5658]_  = \new_[32340]_  & \s15_data_i[27] ;
  assign \new_[5659]_  = ~\new_[5833]_  | ~\new_[5850]_ ;
  assign \new_[5660]_  = ~\new_[5835]_  | ~\new_[5854]_ ;
  assign \new_[5661]_  = ~\new_[5857]_  | ~\new_[5858]_ ;
  assign \new_[5662]_  = ~\new_[5860]_  | ~\new_[5859]_ ;
  assign \new_[5663]_  = ~\new_[5861]_  & (~\new_[6020]_  | ~\new_[4441]_ );
  assign \new_[5664]_  = ~\new_[5839]_  | ~\new_[5862]_ ;
  assign \new_[5665]_  = ~\new_[5841]_  | ~\new_[5864]_ ;
  assign \new_[5666]_  = ~\new_[5867]_  | ~\new_[5868]_ ;
  assign \new_[5667]_  = ~\new_[5870]_  | ~\new_[5871]_ ;
  assign \new_[5668]_  = ~\new_[5873]_  | (~\new_[5949]_  & ~\new_[31682]_ );
  assign \new_[5669]_  = ~\new_[5874]_  & (~\new_[6020]_  | ~\new_[4446]_ );
  assign \new_[5670]_  = ~\new_[5875]_  & (~\new_[6020]_  | ~\new_[4447]_ );
  assign \new_[5671]_  = ~\new_[5846]_  | ~\new_[5877]_ ;
  assign \new_[5672]_  = ~\new_[5878]_  | (~\new_[5949]_  & ~\new_[31829]_ );
  assign \new_[5673]_  = ~\new_[5879]_  & (~\new_[6020]_  | ~\new_[4451]_ );
  assign \new_[5674]_  = ~\new_[5722]_ ;
  assign \new_[5675]_  = ~\new_[6022]_  & ~\new_[31785]_ ;
  assign \new_[5676]_  = ~\new_[5892]_  & ~\new_[31557]_ ;
  assign \new_[5677]_  = ~\new_[5892]_  & ~\new_[31816]_ ;
  assign \new_[5678]_  = ~\new_[5892]_  & ~\new_[31620]_ ;
  assign \new_[5679]_  = ~\new_[5762]_ ;
  assign \new_[5680]_  = ~\new_[5763]_ ;
  assign \new_[5681]_  = \new_[5765]_ ;
  assign \new_[5682]_  = \new_[5765]_ ;
  assign \new_[5683]_  = ~\new_[5766]_ ;
  assign \new_[5684]_  = ~\new_[5767]_ ;
  assign \new_[5685]_  = ~\new_[5767]_ ;
  assign \new_[5686]_  = ~\new_[5767]_ ;
  assign \new_[5687]_  = ~\new_[32191]_ ;
  assign \new_[5688]_  = ~\new_[6016]_  | ~\new_[4454]_ ;
  assign \new_[5689]_  = ~\new_[5768]_ ;
  assign \new_[5690]_  = ~\new_[5769]_ ;
  assign \new_[5691]_  = ~\new_[5770]_ ;
  assign \new_[5692]_  = ~\new_[5771]_ ;
  assign \new_[5693]_  = ~\new_[5772]_ ;
  assign \new_[5694]_  = \new_[5775]_ ;
  assign \new_[5695]_  = ~\new_[5775]_ ;
  assign \new_[5696]_  = ~\new_[5776]_ ;
  assign \new_[5697]_  = ~\new_[5890]_  & ~\new_[31807]_ ;
  assign \new_[5698]_  = ~\new_[5888]_  & ~\new_[31693]_ ;
  assign \new_[5699]_  = ~\new_[5886]_  | ~\new_[3873]_ ;
  assign \new_[5700]_  = ~\new_[5888]_  & ~\new_[31917]_ ;
  assign \new_[5701]_  = ~\new_[5886]_  | ~\new_[3874]_ ;
  assign \new_[5702]_  = ~\new_[5893]_  | ~\new_[4266]_ ;
  assign \new_[5703]_  = ~\new_[5887]_  | ~\new_[3875]_ ;
  assign \new_[5704]_  = ~\new_[5887]_  | ~\new_[3876]_ ;
  assign \new_[5705]_  = ~\new_[5886]_  | ~\new_[3877]_ ;
  assign \new_[5706]_  = ~\new_[5887]_  | ~\new_[3878]_ ;
  assign \new_[5707]_  = ~\new_[5888]_  & ~\new_[31727]_ ;
  assign \new_[5708]_  = ~\new_[5886]_  | ~\new_[3879]_ ;
  assign \new_[5709]_  = ~\new_[5893]_  | ~\new_[4271]_ ;
  assign \new_[5710]_  = ~\new_[5887]_  | ~\new_[3880]_ ;
  assign \new_[5711]_  = ~\new_[5884]_  & ~\new_[31646]_ ;
  assign \new_[5712]_  = ~\new_[5887]_  | ~\new_[3881]_ ;
  assign \new_[5713]_  = ~\new_[32188]_  | ~\new_[4060]_ ;
  assign \new_[5714]_  = ~\new_[5888]_  & ~\new_[31558]_ ;
  assign \new_[5715]_  = ~\new_[5887]_  | ~\new_[3883]_ ;
  assign \new_[5716]_  = ~\new_[5887]_  | ~\new_[3884]_ ;
  assign \new_[5717]_  = ~\new_[5886]_  | ~\new_[3885]_ ;
  assign \new_[5718]_  = ~\new_[5890]_  & ~\new_[31904]_ ;
  assign \new_[5719]_  = ~\new_[5888]_  & ~\new_[31601]_ ;
  assign \new_[5720]_  = ~\new_[5888]_  & ~\new_[31680]_ ;
  assign \new_[5721]_  = ~\new_[5887]_  | ~\new_[3888]_ ;
  assign \new_[5722]_  = \new_[5831]_ ;
  assign \new_[5723]_  = ~\new_[5934]_ ;
  assign \new_[5724]_  = ~\new_[5952]_  | ~\new_[4102]_ ;
  assign \new_[5725]_  = ~\new_[5953]_  | ~\new_[4118]_ ;
  assign \new_[5726]_  = ~\new_[5954]_  | ~\new_[4037]_ ;
  assign \new_[5727]_  = ~\new_[5952]_  | ~\new_[4103]_ ;
  assign \new_[5728]_  = ~\new_[5953]_  | ~\new_[4119]_ ;
  assign \new_[5729]_  = ~\new_[5952]_  | ~\new_[4104]_ ;
  assign \new_[5730]_  = ~\new_[5953]_  | ~\new_[4120]_ ;
  assign \new_[5731]_  = ~\new_[5952]_  | ~\new_[4105]_ ;
  assign \new_[5732]_  = ~\new_[5953]_  | ~\new_[4121]_ ;
  assign \new_[5733]_  = ~\new_[5955]_  & ~\new_[31653]_ ;
  assign \new_[5734]_  = ~\new_[5952]_  | ~\new_[4106]_ ;
  assign \new_[5735]_  = ~\new_[5953]_  | ~\new_[4122]_ ;
  assign \new_[5736]_  = ~\new_[5952]_  | ~\new_[4107]_ ;
  assign \new_[5737]_  = ~\new_[5953]_  | ~\new_[4123]_ ;
  assign \new_[5738]_  = ~\new_[5954]_  | ~\new_[4042]_ ;
  assign \new_[5739]_  = ~\new_[5954]_  | ~\new_[4043]_ ;
  assign \new_[5740]_  = ~\new_[5952]_  | ~\new_[4108]_ ;
  assign \new_[5741]_  = ~\new_[5953]_  | ~\new_[4124]_ ;
  assign \new_[5742]_  = ~\new_[5954]_  | ~\new_[4044]_ ;
  assign \new_[5743]_  = ~\new_[5952]_  | ~\new_[4109]_ ;
  assign \new_[5744]_  = ~\new_[5953]_  | ~\new_[4125]_ ;
  assign \new_[5745]_  = ~\new_[5952]_  | ~\new_[4110]_ ;
  assign \new_[5746]_  = ~\new_[5953]_  | ~\new_[4126]_ ;
  assign \new_[5747]_  = ~\new_[5955]_  & ~\new_[31768]_ ;
  assign \new_[5748]_  = ~\new_[5952]_  | ~\new_[4111]_ ;
  assign \new_[5749]_  = ~\new_[5953]_  | ~\new_[4127]_ ;
  assign \new_[5750]_  = ~\new_[5952]_  | ~\new_[4112]_ ;
  assign \new_[5751]_  = ~\new_[5953]_  | ~\new_[4128]_ ;
  assign \new_[5752]_  = ~\new_[5952]_  | ~\new_[4113]_ ;
  assign \new_[5753]_  = ~\new_[5953]_  | ~\new_[4129]_ ;
  assign \new_[5754]_  = ~\new_[5952]_  | ~\new_[4114]_ ;
  assign \new_[5755]_  = ~\new_[5953]_  | ~\new_[4130]_ ;
  assign \new_[5756]_  = ~\new_[5955]_  & ~\new_[31886]_ ;
  assign \new_[5757]_  = ~\new_[5952]_  | ~\new_[4115]_ ;
  assign \new_[5758]_  = ~\new_[5955]_  & ~\new_[31858]_ ;
  assign \new_[5759]_  = ~\new_[5953]_  | ~\new_[4131]_ ;
  assign \new_[5760]_  = ~\new_[5952]_  | ~\new_[4116]_ ;
  assign \new_[5761]_  = ~\new_[5953]_  | ~\new_[4132]_ ;
  assign \new_[5762]_  = ~\new_[5935]_  | ~\new_[6389]_ ;
  assign \new_[5763]_  = ~\new_[32284]_ ;
  assign \new_[5764]_  = \new_[5847]_ ;
  assign \new_[5765]_  = ~\new_[5847]_ ;
  assign \new_[5766]_  = ~\new_[5937]_  | ~\new_[4454]_ ;
  assign \new_[5767]_  = ~\new_[5941]_  | ~\new_[4454]_ ;
  assign \new_[5768]_  = ~\new_[5935]_  | ~\new_[6373]_ ;
  assign \new_[5769]_  = ~\new_[5935]_  | ~\new_[32287]_ ;
  assign \new_[5770]_  = ~\new_[5935]_  | ~\new_[32330]_ ;
  assign \new_[5771]_  = ~\new_[32070]_  | ~\new_[4454]_ ;
  assign \new_[5772]_  = ~\new_[5848]_ ;
  assign \new_[5773]_  = ~\new_[5848]_ ;
  assign \new_[5774]_  = ~\new_[5848]_ ;
  assign \new_[5775]_  = ~\new_[5947]_  | ~\new_[4454]_ ;
  assign \new_[5776]_  = ~\new_[5849]_ ;
  assign \new_[5777]_  = ~\new_[5937]_  | ~\new_[4052]_ ;
  assign \new_[5778]_  = ~\new_[5941]_  | ~\new_[4068]_ ;
  assign \new_[5779]_  = ~\new_[5937]_  | ~\new_[4053]_ ;
  assign \new_[5780]_  = ~\new_[32192]_  | ~\new_[4083]_ ;
  assign \new_[5781]_  = ~\new_[32171]_  | ~\new_[4134]_ ;
  assign \new_[5782]_  = ~\new_[5941]_  | ~\new_[4069]_ ;
  assign \new_[5783]_  = ~\new_[5946]_  | ~\new_[4168]_ ;
  assign \new_[5784]_  = ~\new_[5936]_  & ~\new_[31413]_ ;
  assign \new_[5785]_  = ~\new_[5938]_  & ~\new_[31412]_ ;
  assign \new_[5786]_  = ~\new_[5946]_  | ~\new_[4169]_ ;
  assign \new_[5787]_  = ~\new_[5940]_  & ~\new_[31572]_ ;
  assign \new_[5788]_  = ~\new_[32192]_  | ~\new_[4086]_ ;
  assign \new_[5789]_  = ~\new_[5937]_  | ~\new_[4056]_ ;
  assign \new_[5790]_  = ~\new_[32171]_  | ~\new_[4137]_ ;
  assign \new_[5791]_  = ~\new_[5961]_  & ~\new_[31755]_ ;
  assign \new_[5792]_  = ~\new_[5960]_  | ~\new_[4253]_ ;
  assign \new_[5793]_  = ~\new_[5946]_  | ~\new_[4170]_ ;
  assign \new_[5794]_  = ~\new_[5941]_  | ~\new_[4072]_ ;
  assign \new_[5795]_  = ~\new_[5946]_  | ~\new_[4171]_ ;
  assign \new_[5796]_  = ~\new_[5962]_  & ~\new_[31662]_ ;
  assign \new_[5797]_  = ~\new_[5936]_  & ~\new_[31700]_ ;
  assign \new_[5798]_  = ~\new_[5937]_  | ~\new_[4058]_ ;
  assign \new_[5799]_  = ~\new_[32192]_  | ~\new_[4088]_ ;
  assign \new_[5800]_  = ~\new_[32171]_  | ~\new_[4139]_ ;
  assign \new_[5801]_  = ~\new_[5946]_  | ~\new_[4173]_ ;
  assign \new_[5802]_  = ~\new_[5936]_  & ~\new_[31580]_ ;
  assign \new_[5803]_  = ~\new_[5951]_  & ~\new_[31659]_ ;
  assign \new_[5804]_  = ~\new_[5941]_  | ~\new_[4097]_ ;
  assign \new_[5805]_  = ~\new_[5946]_  | ~\new_[4174]_ ;
  assign \new_[5806]_  = ~\new_[5951]_  & ~\new_[31929]_ ;
  assign \new_[5807]_  = ~\new_[5943]_  | ~\new_[4099]_ ;
  assign \new_[5808]_  = ~\new_[32171]_  | ~\new_[4142]_ ;
  assign \new_[5809]_  = ~\new_[4061]_  | ~\new_[5939]_ ;
  assign \new_[5810]_  = ~\new_[5962]_  & ~\new_[31811]_ ;
  assign \new_[5811]_  = ~\new_[5948]_  | ~\new_[4176]_ ;
  assign \new_[5812]_  = ~\new_[5962]_  & ~\new_[31670]_ ;
  assign \new_[5813]_  = ~\new_[5938]_  & ~\new_[31600]_ ;
  assign \new_[5814]_  = ~\new_[5946]_  | ~\new_[4177]_ ;
  assign \new_[5815]_  = ~\new_[5962]_  & ~\new_[31801]_ ;
  assign \new_[5816]_  = ~\new_[5951]_  & ~\new_[31708]_ ;
  assign \new_[5817]_  = ~\new_[5938]_  & ~\new_[31891]_ ;
  assign \new_[5818]_  = ~\new_[5946]_  | ~\new_[4178]_ ;
  assign \new_[5819]_  = ~\new_[5936]_  & ~\new_[31851]_ ;
  assign \new_[5820]_  = ~\new_[5939]_  | ~\new_[4065]_ ;
  assign \new_[5821]_  = ~\new_[5962]_  & ~\new_[31909]_ ;
  assign \new_[5822]_  = ~\new_[5939]_  | ~\new_[4066]_ ;
  assign \new_[5823]_  = ~\new_[5950]_  | ~\new_[4147]_ ;
  assign \new_[5824]_  = ~\new_[5961]_  & ~\new_[31761]_ ;
  assign \new_[5825]_  = ~\new_[5946]_  | ~\new_[4181]_ ;
  assign \new_[5826]_  = ~\new_[5962]_  & ~\new_[31627]_ ;
  assign \new_[5827]_  = ~\new_[5940]_  & ~\new_[31632]_ ;
  assign \new_[5828]_  = ~\new_[5951]_  & ~\new_[31771]_ ;
  assign \new_[5829]_  = ~\new_[5886]_ ;
  assign \new_[5830]_  = \\s14_msel_arb2_state_reg[0] ;
  assign \new_[5831]_  = ~\new_[6272]_  & ~\new_[31931]_ ;
  assign \new_[5832]_  = \new_[5934]_ ;
  assign \new_[5833]_  = ~\new_[6021]_  | ~\new_[4438]_ ;
  assign \new_[5834]_  = ~\new_[6017]_  | ~\new_[4233]_ ;
  assign \new_[5835]_  = ~\new_[6020]_  | ~\new_[4439]_ ;
  assign \new_[5836]_  = ~\new_[6018]_  | ~\new_[4235]_ ;
  assign \new_[5837]_  = ~\new_[6017]_  | ~\new_[4234]_ ;
  assign \new_[5838]_  = ~\new_[6187]_  | ~\new_[4236]_ ;
  assign \new_[5839]_  = ~\new_[6020]_  | ~\new_[4442]_ ;
  assign \new_[5840]_  = ~\new_[6017]_  | ~\new_[4237]_ ;
  assign \new_[5841]_  = ~\new_[6020]_  | ~\new_[4444]_ ;
  assign \new_[5842]_  = ~\new_[6017]_  | ~\new_[4239]_ ;
  assign \new_[5843]_  = ~\new_[6018]_  | ~\new_[4247]_ ;
  assign \new_[5844]_  = ~\new_[6020]_  | ~\new_[4452]_ ;
  assign \new_[5845]_  = ~\new_[6018]_  | ~\new_[4243]_ ;
  assign \new_[5846]_  = ~\new_[6021]_  | ~\new_[4449]_ ;
  assign \new_[5847]_  = ~\new_[6011]_  | ~\new_[4454]_ ;
  assign \new_[5848]_  = ~\new_[6029]_  | ~\new_[4454]_ ;
  assign \new_[5849]_  = ~\new_[6030]_  | ~\new_[4454]_ ;
  assign \new_[5850]_  = ~\new_[6012]_  | ~\new_[4216]_ ;
  assign \new_[5851]_  = ~\new_[32192]_  | ~\new_[4082]_ ;
  assign \new_[5852]_  = ~\new_[6026]_  | ~\new_[4200]_ ;
  assign \new_[5853]_  = ~\new_[6030]_  | ~\new_[4265]_ ;
  assign \new_[5854]_  = ~\new_[6010]_  | ~\new_[4217]_ ;
  assign \new_[5855]_  = ~\new_[6027]_  | ~\new_[4150]_ ;
  assign \new_[5856]_  = ~\new_[6026]_  | ~\new_[4201]_ ;
  assign \new_[5857]_  = ~\new_[6030]_  | ~\new_[4267]_ ;
  assign \new_[5858]_  = ~\new_[32288]_  | ~\new_[4202]_ ;
  assign \new_[5859]_  = ~\new_[32288]_  | ~\new_[4203]_ ;
  assign \new_[5860]_  = ~\new_[6030]_  | ~\new_[4268]_ ;
  assign \new_[5861]_  = ~\new_[6013]_  & ~\new_[31635]_ ;
  assign \new_[5862]_  = ~\new_[6010]_  | ~\new_[4220]_ ;
  assign \new_[5863]_  = ~\new_[6027]_  | ~\new_[4153]_ ;
  assign \new_[5864]_  = ~\new_[6010]_  | ~\new_[4222]_ ;
  assign \new_[5865]_  = ~\new_[6027]_  | ~\new_[4155]_ ;
  assign \new_[5866]_  = ~\new_[6026]_  | ~\new_[4206]_ ;
  assign \new_[5867]_  = ~\new_[6030]_  | ~\new_[4272]_ ;
  assign \new_[5868]_  = ~\new_[32285]_  | ~\new_[4207]_ ;
  assign \new_[5869]_  = ~\new_[6028]_  | ~\new_[4263]_ ;
  assign \new_[5870]_  = ~\new_[6030]_  | ~\new_[4273]_ ;
  assign \new_[5871]_  = ~\new_[32288]_  | ~\new_[4208]_ ;
  assign \new_[5872]_  = ~\new_[6010]_  | ~\new_[4230]_ ;
  assign \new_[5873]_  = ~\new_[6010]_  | ~\new_[4231]_ ;
  assign \new_[5874]_  = ~\new_[6013]_  & ~\new_[31555]_ ;
  assign \new_[5875]_  = ~\new_[6013]_  & ~\new_[31717]_ ;
  assign \new_[5876]_  = ~\new_[6030]_  | ~\new_[4277]_ ;
  assign \new_[5877]_  = ~\new_[6012]_  | ~\new_[4227]_ ;
  assign \new_[5878]_  = ~\new_[6010]_  | ~\new_[4228]_ ;
  assign \new_[5879]_  = ~\new_[6013]_  & ~\new_[31918]_ ;
  assign \new_[5880]_  = ~\new_[32282]_ ;
  assign \new_[5881]_  = ~\new_[32282]_ ;
  assign \new_[5882]_  = ~\new_[32315]_ ;
  assign \new_[5883]_  = ~\new_[32341]_ ;
  assign \new_[5884]_  = ~\new_[5939]_ ;
  assign \new_[5885]_  = ~\new_[5941]_ ;
  assign \new_[5886]_  = ~\new_[5944]_ ;
  assign \new_[5887]_  = ~\new_[5944]_ ;
  assign \new_[5888]_  = ~\new_[5948]_ ;
  assign \new_[5889]_  = ~\new_[5949]_ ;
  assign \new_[5890]_  = ~\new_[5950]_ ;
  assign \new_[5891]_  = ~\new_[32171]_ ;
  assign \new_[5892]_  = ~\new_[5954]_ ;
  assign \new_[5893]_  = ~\new_[5961]_ ;
  assign \new_[5894]_  = \\s10_msel_arb0_state_reg[1] ;
  assign \new_[5895]_  = \\s11_msel_arb0_state_reg[1] ;
  assign \new_[5896]_  = \\s12_msel_arb0_state_reg[1] ;
  assign \new_[5897]_  = \\s13_msel_arb0_state_reg[1] ;
  assign \new_[5898]_  = \\s14_msel_arb0_state_reg[1] ;
  assign \new_[5899]_  = \\s15_msel_arb0_state_reg[1] ;
  assign \new_[5900]_  = \\s1_msel_arb0_state_reg[1] ;
  assign \new_[5901]_  = \\s2_msel_arb0_state_reg[1] ;
  assign \new_[5902]_  = \\s3_msel_arb0_state_reg[1] ;
  assign \new_[5903]_  = \\s4_msel_arb0_state_reg[1] ;
  assign \new_[5904]_  = \\s5_msel_arb0_state_reg[1] ;
  assign \new_[5905]_  = \\s6_msel_arb0_state_reg[1] ;
  assign \new_[5906]_  = \\s8_msel_arb0_state_reg[1] ;
  assign \new_[5907]_  = \\s9_msel_arb0_state_reg[1] ;
  assign \new_[5908]_  = \\s0_msel_arb0_state_reg[1] ;
  assign \new_[5909]_  = \\s11_msel_arb0_state_reg[0] ;
  assign \new_[5910]_  = \\s11_msel_arb1_state_reg[1] ;
  assign \new_[5911]_  = \\s12_msel_arb0_state_reg[0] ;
  assign \new_[5912]_  = \\s13_msel_arb0_state_reg[0] ;
  assign \new_[5913]_  = \\s13_msel_arb2_state_reg[0] ;
  assign \new_[5914]_  = \\s14_msel_arb0_state_reg[0] ;
  assign \new_[5915]_  = \\s15_msel_arb2_state_reg[0] ;
  assign \new_[5916]_  = \\s15_msel_arb3_state_reg[1] ;
  assign \new_[5917]_  = \\s3_msel_arb0_state_reg[0] ;
  assign \new_[5918]_  = \\s4_msel_arb0_state_reg[0] ;
  assign \new_[5919]_  = \\s4_msel_arb2_state_reg[0] ;
  assign \new_[5920]_  = \\s4_msel_arb2_state_reg[1] ;
  assign \new_[5921]_  = \\s5_msel_arb0_state_reg[0] ;
  assign \new_[5922]_  = \\s5_msel_arb3_state_reg[1] ;
  assign \new_[5923]_  = \\s6_msel_arb0_state_reg[0] ;
  assign \new_[5924]_  = \\s6_msel_arb1_state_reg[0] ;
  assign \new_[5925]_  = \\s6_msel_arb1_state_reg[1] ;
  assign \new_[5926]_  = \\s7_msel_arb0_state_reg[0] ;
  assign \new_[5927]_  = \\s8_msel_arb0_state_reg[0] ;
  assign \new_[5928]_  = \\s8_msel_arb1_state_reg[1] ;
  assign \new_[5929]_  = \\s8_msel_arb3_state_reg[1] ;
  assign \new_[5930]_  = \\s9_msel_arb3_state_reg[0] ;
  assign \new_[5931]_  = \\s9_msel_arb2_state_reg[0] ;
  assign \new_[5932]_  = \\s0_msel_arb2_state_reg[0] ;
  assign \new_[5933]_  = \\s7_msel_arb0_state_reg[1] ;
  assign \new_[5934]_  = ~\new_[6188]_  & ~\new_[31931]_ ;
  assign \new_[5935]_  = ~\new_[6009]_ ;
  assign \new_[5936]_  = ~\new_[6012]_ ;
  assign \new_[5937]_  = ~\new_[6014]_ ;
  assign \new_[5938]_  = \new_[6014]_ ;
  assign \new_[5939]_  = ~\new_[6014]_ ;
  assign \new_[5940]_  = \new_[6014]_ ;
  assign \new_[5941]_  = ~\new_[6015]_ ;
  assign \new_[5942]_  = ~\new_[32192]_ ;
  assign \new_[5943]_  = \new_[32192]_ ;
  assign \new_[5944]_  = ~\new_[6016]_ ;
  assign \new_[5945]_  = ~\new_[6018]_ ;
  assign \new_[5946]_  = ~\new_[6019]_ ;
  assign \new_[5947]_  = ~\new_[6019]_ ;
  assign \new_[5948]_  = ~\new_[6019]_ ;
  assign \new_[5949]_  = ~\new_[6021]_ ;
  assign \new_[5950]_  = ~\new_[32172]_ ;
  assign \new_[5951]_  = \new_[32172]_ ;
  assign \new_[5952]_  = ~\new_[6022]_ ;
  assign \new_[5953]_  = ~\new_[6023]_ ;
  assign \new_[5954]_  = ~\new_[6024]_ ;
  assign \new_[5955]_  = \new_[6024]_ ;
  assign \new_[5956]_  = ~\new_[6025]_ ;
  assign \new_[5957]_  = ~\new_[6027]_ ;
  assign \new_[5958]_  = ~\new_[6028]_ ;
  assign \new_[5959]_  = ~\new_[6029]_ ;
  assign \new_[5960]_  = \new_[6029]_ ;
  assign \new_[5961]_  = ~\new_[6030]_ ;
  assign \new_[5962]_  = ~\new_[6030]_ ;
  assign \new_[5963]_  = \\s10_msel_arb2_state_reg[1] ;
  assign \new_[5964]_  = \\s10_msel_arb2_state_reg[0] ;
  assign \new_[5965]_  = \\s11_msel_arb2_state_reg[1] ;
  assign \new_[5966]_  = \\s11_msel_arb3_state_reg[1] ;
  assign \new_[5967]_  = \\s12_msel_arb1_state_reg[1] ;
  assign \new_[5968]_  = \\s12_msel_arb2_state_reg[0] ;
  assign \new_[5969]_  = \\s12_msel_arb2_state_reg[1] ;
  assign \new_[5970]_  = \\s13_msel_arb1_state_reg[1] ;
  assign \new_[5971]_  = \\s13_msel_arb2_state_reg[1] ;
  assign \new_[5972]_  = \\s14_msel_arb2_state_reg[1] ;
  assign \new_[5973]_  = \\s14_msel_arb2_state_reg[2] ;
  assign \new_[5974]_  = \\s15_msel_arb0_state_reg[0] ;
  assign \new_[5975]_  = \\s15_msel_arb1_state_reg[1] ;
  assign \new_[5976]_  = \\s15_msel_arb2_state_reg[1] ;
  assign \new_[5977]_  = \\s15_msel_arb2_state_reg[2] ;
  assign \new_[5978]_  = \\s1_msel_arb0_state_reg[0] ;
  assign \new_[5979]_  = \\s1_msel_arb2_state_reg[0] ;
  assign \new_[5980]_  = \\s1_msel_arb2_state_reg[1] ;
  assign \new_[5981]_  = \\s2_msel_arb2_state_reg[0] ;
  assign \new_[5982]_  = \\s2_msel_arb2_state_reg[1] ;
  assign \new_[5983]_  = \\s2_msel_arb0_state_reg[0] ;
  assign \new_[5984]_  = \\s3_msel_arb1_state_reg[1] ;
  assign \new_[5985]_  = \\s3_msel_arb2_state_reg[0] ;
  assign \new_[5986]_  = \\s3_msel_arb2_state_reg[1] ;
  assign \new_[5987]_  = \\s3_msel_arb3_state_reg[1] ;
  assign \new_[5988]_  = \\s4_msel_arb2_state_reg[2] ;
  assign \new_[5989]_  = \\s5_msel_arb1_state_reg[1] ;
  assign \new_[5990]_  = \\s5_msel_arb2_state_reg[1] ;
  assign \new_[5991]_  = \\s5_msel_arb3_state_reg[0] ;
  assign \new_[5992]_  = \\s5_msel_arb3_state_reg[2] ;
  assign \new_[5993]_  = \\s6_msel_arb2_state_reg[1] ;
  assign \new_[5994]_  = \\s6_msel_arb2_state_reg[0] ;
  assign \new_[5995]_  = \\s6_msel_arb3_state_reg[1] ;
  assign \new_[5996]_  = \\s6_msel_arb3_state_reg[0] ;
  assign \new_[5997]_  = \\s7_msel_arb2_state_reg[0] ;
  assign \new_[5998]_  = \\s7_msel_arb2_state_reg[1] ;
  assign \new_[5999]_  = \\s8_msel_arb2_state_reg[0] ;
  assign \new_[6000]_  = \\s8_msel_arb2_state_reg[1] ;
  assign \new_[6001]_  = \\s8_msel_arb3_state_reg[0] ;
  assign \new_[6002]_  = \\s9_msel_arb0_state_reg[0] ;
  assign \new_[6003]_  = \\s9_msel_arb2_state_reg[2] ;
  assign \new_[6004]_  = \\s0_msel_arb0_state_reg[0] ;
  assign \new_[6005]_  = \\s0_msel_arb2_state_reg[1] ;
  assign \new_[6006]_  = \\s0_msel_arb2_state_reg[2] ;
  assign \new_[6007]_  = \\s0_msel_arb3_state_reg[0] ;
  assign n6464 = ~\new_[9837]_  | ~\new_[9838]_  | ~\new_[7298]_  | ~\new_[6357]_ ;
  assign \new_[6009]_  = ~\new_[32173]_  | ~\new_[4454]_ ;
  assign \new_[6010]_  = ~\new_[32329]_ ;
  assign \new_[6011]_  = ~\new_[32329]_ ;
  assign \new_[6012]_  = ~\new_[32329]_ ;
  assign \new_[6013]_  = \new_[32329]_ ;
  assign \new_[6014]_  = ~\new_[6223]_  | ~\new_[6390]_ ;
  assign \new_[6015]_  = ~\new_[6223]_  | ~\new_[6373]_ ;
  assign \new_[6016]_  = ~\new_[6222]_  & ~\new_[6287]_ ;
  assign \new_[6017]_  = \new_[6187]_ ;
  assign \new_[6018]_  = \new_[6187]_ ;
  assign \new_[6019]_  = ~\new_[6374]_  | ~\new_[6221]_ ;
  assign \new_[6020]_  = ~\new_[6188]_ ;
  assign \new_[6021]_  = ~\new_[6188]_ ;
  assign \new_[6022]_  = ~\new_[32173]_  | ~\new_[6373]_ ;
  assign \new_[6023]_  = ~\new_[32287]_  | ~\new_[32173]_ ;
  assign \new_[6024]_  = ~\new_[6390]_  | ~\new_[32173]_ ;
  assign \new_[6025]_  = ~\new_[32286]_ ;
  assign \new_[6026]_  = ~\new_[32286]_ ;
  assign \new_[6027]_  = \new_[32070]_ ;
  assign \new_[6028]_  = ~\new_[32316]_ ;
  assign \new_[6029]_  = ~\new_[32317]_ ;
  assign \new_[6030]_  = ~\new_[6198]_ ;
  assign \new_[6031]_  = \\s14_msel_arb3_state_reg[0] ;
  assign \new_[6032]_  = \\s12_msel_arb1_state_reg[0] ;
  assign \new_[6033]_  = \\s10_msel_arb1_state_reg[0] ;
  assign \new_[6034]_  = \\s10_msel_arb1_state_reg[1] ;
  assign \new_[6035]_  = \\s10_msel_arb2_state_reg[2] ;
  assign \new_[6036]_  = \\s11_msel_arb0_state_reg[2] ;
  assign \new_[6037]_  = \\s11_msel_arb1_state_reg[2] ;
  assign \new_[6038]_  = \\s11_msel_arb2_state_reg[0] ;
  assign \new_[6039]_  = \\s11_msel_arb2_state_reg[2] ;
  assign \new_[6040]_  = \\s11_msel_arb1_state_reg[0] ;
  assign \new_[6041]_  = \\s11_msel_arb3_state_reg[2] ;
  assign \new_[6042]_  = \\s12_msel_arb0_state_reg[2] ;
  assign \new_[6043]_  = \\s12_msel_arb1_state_reg[2] ;
  assign \new_[6044]_  = \\s12_msel_arb2_state_reg[2] ;
  assign \new_[6045]_  = \\s13_msel_arb0_state_reg[2] ;
  assign \new_[6046]_  = \\s12_msel_arb3_state_reg[1] ;
  assign \new_[6047]_  = \\s13_msel_arb2_state_reg[2] ;
  assign \new_[6048]_  = \\s13_msel_arb3_state_reg[1] ;
  assign \new_[6049]_  = \\s14_msel_arb1_state_reg[2] ;
  assign \new_[6050]_  = \\s14_msel_arb1_state_reg[1] ;
  assign \new_[6051]_  = \\s14_msel_arb0_state_reg[2] ;
  assign \new_[6052]_  = \\s14_msel_arb3_state_reg[1] ;
  assign \new_[6053]_  = \\s14_msel_arb3_state_reg[2] ;
  assign \new_[6054]_  = \\s15_msel_arb1_state_reg[0] ;
  assign \new_[6055]_  = \\s15_msel_arb3_state_reg[0] ;
  assign \new_[6056]_  = \\s1_msel_arb0_state_reg[2] ;
  assign \new_[6057]_  = \\s1_msel_arb1_state_reg[1] ;
  assign \new_[6058]_  = \\s1_msel_arb2_state_reg[2] ;
  assign \new_[6059]_  = \\s1_msel_arb3_state_reg[0] ;
  assign \new_[6060]_  = \\s1_msel_arb3_state_reg[1] ;
  assign \new_[6061]_  = \\s2_msel_arb1_state_reg[1] ;
  assign \new_[6062]_  = \\s2_msel_arb0_state_reg[2] ;
  assign \new_[6063]_  = \\s2_msel_arb2_state_reg[2] ;
  assign \new_[6064]_  = \\s2_msel_arb3_state_reg[0] ;
  assign \new_[6065]_  = \\s2_msel_arb3_state_reg[1] ;
  assign \new_[6066]_  = \\s3_msel_arb1_state_reg[0] ;
  assign \new_[6067]_  = \\s3_msel_arb0_state_reg[2] ;
  assign \new_[6068]_  = \\s3_msel_arb2_state_reg[2] ;
  assign \new_[6069]_  = \\s4_msel_arb1_state_reg[0] ;
  assign \new_[6070]_  = \\s4_msel_arb1_state_reg[1] ;
  assign \new_[6071]_  = \\s4_msel_arb3_state_reg[0] ;
  assign \new_[6072]_  = \\s5_msel_arb1_state_reg[0] ;
  assign \new_[6073]_  = \\s5_msel_arb1_state_reg[2] ;
  assign \new_[6074]_  = \\s5_msel_arb0_state_reg[2] ;
  assign \new_[6075]_  = \\s6_msel_arb0_state_reg[2] ;
  assign \new_[6076]_  = \\s6_msel_arb1_state_reg[2] ;
  assign \new_[6077]_  = \\s6_msel_arb2_state_reg[2] ;
  assign \new_[6078]_  = \\s7_msel_arb1_state_reg[0] ;
  assign \new_[6079]_  = \\s7_msel_arb1_state_reg[2] ;
  assign \new_[6080]_  = \\s7_msel_arb0_state_reg[2] ;
  assign \new_[6081]_  = \\s7_msel_arb2_state_reg[2] ;
  assign \new_[6082]_  = \\s7_msel_arb3_state_reg[2] ;
  assign \new_[6083]_  = \\s8_msel_arb0_state_reg[2] ;
  assign \new_[6084]_  = \\s8_msel_arb1_state_reg[0] ;
  assign \new_[6085]_  = \\s7_msel_arb3_state_reg[1] ;
  assign \new_[6086]_  = \\s8_msel_arb3_state_reg[2] ;
  assign \new_[6087]_  = \\s9_msel_arb0_state_reg[2] ;
  assign \new_[6088]_  = \\s9_msel_arb2_state_reg[1] ;
  assign \new_[6089]_  = \\s9_msel_arb1_state_reg[2] ;
  assign \new_[6090]_  = \\s9_msel_arb3_state_reg[1] ;
  assign \new_[6091]_  = \\s0_msel_arb0_state_reg[2] ;
  assign \new_[6092]_  = \\s0_msel_arb1_state_reg[1] ;
  assign \new_[6093]_  = \\s0_msel_arb1_state_reg[2] ;
  assign \new_[6094]_  = \\s10_msel_arb0_state_reg[0] ;
  assign \new_[6095]_  = \\s0_msel_arb3_state_reg[2] ;
  assign \new_[6096]_  = \\s13_msel_arb1_state_reg[0] ;
  assign n6474 = \new_[8362]_  | \new_[8363]_  | \new_[6364]_  | \new_[9871]_ ;
  assign n6479 = \new_[8364]_  | \new_[8365]_  | \new_[6365]_  | \new_[11564]_ ;
  assign n6484 = \new_[8367]_  | \new_[8368]_  | \new_[6366]_  | \new_[9880]_ ;
  assign n6489 = \new_[8371]_  | \new_[7902]_  | \new_[6367]_  | \new_[8858]_ ;
  assign n6494 = ~\new_[6599]_  | ~\new_[7899]_  | ~\new_[6601]_  | ~\new_[8796]_ ;
  assign n6509 = \new_[8375]_  | \new_[7904]_  | \new_[6368]_  | \new_[8865]_ ;
  assign n6514 = \new_[8377]_  | \new_[8378]_  | \new_[6369]_  | \new_[8869]_ ;
  assign n6519 = \new_[8379]_  | \new_[8380]_  | \new_[6370]_  | \new_[11633]_ ;
  assign n6524 = \new_[8383]_  | \new_[8384]_  | \new_[6371]_  | \new_[8875]_ ;
  assign n6529 = \new_[8386]_  | \new_[8387]_  | \new_[6372]_  | \new_[9931]_ ;
  assign \s15_data_o[31]  = ~\new_[6646]_  | ~\new_[7348]_  | ~\new_[6644]_  | ~\new_[6645]_ ;
  assign \s15_data_o[30]  = ~\new_[6649]_  | ~\new_[7349]_  | ~\new_[6647]_  | ~\new_[6648]_ ;
  assign \s15_data_o[29]  = ~\new_[8039]_  | ~\new_[6651]_  | ~\new_[6650]_  | ~\new_[7350]_ ;
  assign \s15_data_o[28]  = ~\new_[6654]_  | ~\new_[7351]_  | ~\new_[6652]_  | ~\new_[6653]_ ;
  assign \s15_data_o[27]  = ~\new_[6657]_  | ~\new_[7352]_  | ~\new_[6655]_  | ~\new_[6656]_ ;
  assign \s15_data_o[26]  = ~\new_[6660]_  | ~\new_[7353]_  | ~\new_[6658]_  | ~\new_[6659]_ ;
  assign \s15_data_o[25]  = ~\new_[6663]_  | ~\new_[7354]_  | ~\new_[6661]_  | ~\new_[6662]_ ;
  assign \s15_data_o[24]  = ~\new_[6666]_  | ~\new_[7356]_  | ~\new_[6664]_  | ~\new_[6665]_ ;
  assign \s15_data_o[23]  = ~\new_[6669]_  | ~\new_[7358]_  | ~\new_[6667]_  | ~\new_[6668]_ ;
  assign \s15_data_o[22]  = ~\new_[6672]_  | ~\new_[8044]_  | ~\new_[6670]_  | ~\new_[6671]_ ;
  assign \s15_data_o[21]  = ~\new_[8046]_  | ~\new_[6675]_  | ~\new_[6673]_  | ~\new_[6674]_ ;
  assign \s15_data_o[20]  = ~\new_[6678]_  | ~\new_[7360]_  | ~\new_[6676]_  | ~\new_[6677]_ ;
  assign \s15_data_o[19]  = ~\new_[8049]_  | ~\new_[6681]_  | ~\new_[6679]_  | ~\new_[6680]_ ;
  assign \s15_data_o[18]  = ~\new_[6684]_  | ~\new_[7364]_  | ~\new_[6683]_  | ~\new_[6682]_ ;
  assign \s15_data_o[17]  = ~\new_[6687]_  | ~\new_[7368]_  | ~\new_[6685]_  | ~\new_[6686]_ ;
  assign \s15_data_o[16]  = ~\new_[6690]_  | ~\new_[7371]_  | ~\new_[6688]_  | ~\new_[6689]_ ;
  assign \s15_addr_o[31]  = ~\new_[6700]_  | ~\new_[7393]_  | ~\new_[6431]_  | ~\new_[6699]_ ;
  assign \s15_addr_o[30]  = ~\new_[6702]_  | ~\new_[7394]_  | ~\new_[6432]_  | ~\new_[6701]_ ;
  assign \s15_addr_o[29]  = ~\new_[7395]_  | ~\new_[6705]_  | ~\new_[6703]_  | ~\new_[6704]_ ;
  assign \s15_addr_o[28]  = ~\new_[6707]_  | ~\new_[7396]_  | ~\new_[6433]_  | ~\new_[6706]_ ;
  assign \s15_addr_o[23]  = ~\new_[6710]_  | ~\new_[7397]_  | ~\new_[6708]_  | ~\new_[6709]_ ;
  assign \s15_addr_o[22]  = ~\new_[6713]_  | ~\new_[7398]_  | ~\new_[6711]_  | ~\new_[6712]_ ;
  assign \s15_addr_o[21]  = ~\new_[6716]_  | ~\new_[7399]_  | ~\new_[6714]_  | ~\new_[6715]_ ;
  assign \s15_addr_o[20]  = ~\new_[6719]_  | ~\new_[7401]_  | ~\new_[6717]_  | ~\new_[6718]_ ;
  assign \s15_addr_o[19]  = ~\new_[6722]_  | ~\new_[7402]_  | ~\new_[6720]_  | ~\new_[6721]_ ;
  assign \s15_addr_o[18]  = ~\new_[6726]_  | ~\new_[7403]_  | ~\new_[6723]_  | ~\new_[6725]_ ;
  assign \s15_addr_o[17]  = ~\new_[8088]_  | ~\new_[6729]_  | ~\new_[6727]_  | ~\new_[6728]_ ;
  assign \s15_addr_o[16]  = ~\new_[6732]_  | ~\new_[7404]_  | ~\new_[6730]_  | ~\new_[6731]_ ;
  assign \s15_addr_o[15]  = ~\new_[6735]_  | ~\new_[7405]_  | ~\new_[6733]_  | ~\new_[6734]_ ;
  assign \s15_addr_o[14]  = ~\new_[6738]_  | ~\new_[8091]_  | ~\new_[6736]_  | ~\new_[6737]_ ;
  assign \s15_addr_o[13]  = ~\new_[6741]_  | ~\new_[8092]_  | ~\new_[6739]_  | ~\new_[6740]_ ;
  assign \s15_addr_o[12]  = ~\new_[6744]_  | ~\new_[8093]_  | ~\new_[6742]_  | ~\new_[6743]_ ;
  assign \s15_addr_o[11]  = ~\new_[6747]_  | ~\new_[7407]_  | ~\new_[6745]_  | ~\new_[6746]_ ;
  assign \s15_addr_o[10]  = ~\new_[6750]_  | ~\new_[7408]_  | ~\new_[6748]_  | ~\new_[6749]_ ;
  assign \s15_addr_o[9]  = ~\new_[6753]_  | ~\new_[7409]_  | ~\new_[6751]_  | ~\new_[6752]_ ;
  assign \s15_addr_o[8]  = ~\new_[6756]_  | ~\new_[7410]_  | ~\new_[6754]_  | ~\new_[6755]_ ;
  assign \s15_addr_o[7]  = ~\new_[6759]_  | ~\new_[7411]_  | ~\new_[6757]_  | ~\new_[6758]_ ;
  assign \s15_addr_o[6]  = ~\new_[6762]_  | ~\new_[7412]_  | ~\new_[6760]_  | ~\new_[6761]_ ;
  assign \s15_addr_o[1]  = ~\new_[6765]_  | ~\new_[7415]_  | ~\new_[6763]_  | ~\new_[6764]_ ;
  assign \s15_addr_o[0]  = ~\new_[6768]_  | ~\new_[7417]_  | ~\new_[6766]_  | ~\new_[6767]_ ;
  assign \s15_sel_o[3]  = ~\new_[6771]_  | ~\new_[7418]_  | ~\new_[6769]_  | ~\new_[6770]_ ;
  assign \s15_sel_o[2]  = ~\new_[6774]_  | ~\new_[7420]_  | ~\new_[6772]_  | ~\new_[6773]_ ;
  assign \s15_sel_o[1]  = ~\new_[6776]_  | ~\new_[7422]_  | ~\new_[7421]_  | ~\new_[6775]_ ;
  assign n6499 = ~\new_[18389]_  | ~\new_[10252]_  | ~\new_[6358]_  | ~\new_[7304]_ ;
  assign \s15_sel_o[0]  = ~\new_[6778]_  | ~\new_[7424]_  | ~\new_[7423]_  | ~\new_[6777]_ ;
  assign n6504 = ~\new_[18390]_  | ~\new_[10265]_  | ~\new_[6359]_  | ~\new_[7309]_ ;
  assign n6664 = ~\new_[18401]_  | ~\new_[11955]_  | ~\new_[6360]_  | ~\new_[7337]_ ;
  assign n6534 = ~\new_[18396]_  | ~\new_[10346]_  | ~\new_[6361]_  | ~\new_[7345]_ ;
  assign n6539 = ~\new_[18403]_  | ~\new_[10358]_  | ~\new_[6362]_  | ~\new_[7357]_ ;
  assign n6469 = ~\new_[18385]_  | ~\new_[11906]_  | ~\new_[6363]_  | ~\new_[7279]_ ;
  assign n6544 = ~\new_[7380]_  | ~\new_[6620]_  | ~\new_[7282]_  | ~\new_[6631]_ ;
  assign n6554 = ~\new_[7381]_  | ~\new_[6621]_  | ~\new_[7286]_  | ~\new_[6634]_ ;
  assign n6559 = ~\new_[7383]_  | ~\new_[6622]_  | ~\new_[7291]_  | ~\new_[6635]_ ;
  assign n6564 = ~\new_[9835]_  | ~\new_[8836]_  | ~\new_[8515]_  | ~\new_[6425]_ ;
  assign n6569 = ~\new_[7385]_  | ~\new_[6623]_  | ~\new_[7297]_  | ~\new_[6636]_ ;
  assign n6574 = ~\new_[6426]_  | ~\new_[8007]_  | ~\new_[7300]_ ;
  assign n6584 = ~\new_[7387]_  | ~\new_[6624]_  | ~\new_[7312]_  | ~\new_[6638]_ ;
  assign n6589 = ~\new_[7388]_  | ~\new_[6625]_  | ~\new_[7318]_  | ~\new_[6639]_ ;
  assign n6594 = ~\new_[9849]_  | ~\new_[9850]_  | ~\new_[8551]_  | ~\new_[6427]_ ;
  assign n6604 = ~\new_[7389]_  | ~\new_[6626]_  | ~\new_[7320]_  | ~\new_[6640]_ ;
  assign n6614 = ~\new_[7391]_  | ~\new_[6627]_  | ~\new_[7328]_  | ~\new_[6641]_ ;
  assign n6619 = ~\new_[6695]_  | ~\new_[7330]_  | ~\new_[7331]_  | ~\new_[7329]_ ;
  assign n6629 = ~\new_[6697]_  | ~\new_[7952]_  | ~\new_[7336]_  | ~\new_[7335]_ ;
  assign n6634 = ~\new_[7392]_  | ~\new_[6628]_  | ~\new_[7339]_  | ~\new_[6642]_ ;
  assign n6654 = ~\new_[9858]_  | ~\new_[8850]_  | ~\new_[8567]_  | ~\new_[6428]_ ;
  assign n6649 = ~\new_[11541]_  | ~\new_[9860]_  | ~\new_[8038]_  | ~\new_[6429]_ ;
  assign n6659 = ~\new_[9861]_  | ~\new_[11544]_  | ~\new_[8047]_  | ~\new_[6430]_ ;
  assign \new_[6174]_  = \\s10_msel_arb1_state_reg[2] ;
  assign n6579 = ~\new_[6629]_  | ~\new_[8504]_  | ~\new_[8534]_  | ~\new_[8533]_ ;
  assign \new_[6176]_  = \\s11_msel_arb3_state_reg[0] ;
  assign n6599 = ~\new_[7276]_  | ~\new_[6691]_  | ~\new_[8027]_  | ~\new_[8491]_ ;
  assign n6609 = ~\new_[7277]_  | ~\new_[6692]_  | ~\new_[7327]_  | ~\new_[8493]_ ;
  assign n6644 = ~\new_[6693]_  | ~\new_[6630]_  | ~\new_[6643]_  | ~\new_[7968]_ ;
  assign n6549 = ~\new_[6632]_  | ~\new_[6694]_  | ~\new_[7284]_  | ~\new_[6633]_ ;
  assign n6624 = ~\new_[8030]_  | ~\new_[6696]_  | ~\new_[7332]_  | ~\new_[8031]_ ;
  assign n6639 = ~\new_[7341]_  | ~\new_[6698]_  | ~\new_[7343]_  | ~\new_[7342]_ ;
  assign \new_[6183]_  = \\s9_msel_arb3_state_reg[2] ;
  assign \new_[6184]_  = \\s9_msel_arb1_state_reg[0] ;
  assign \new_[6185]_  = \\s8_msel_arb2_state_reg[2] ;
  assign \new_[6186]_  = \\s8_msel_arb1_state_reg[2] ;
  assign \new_[6187]_  = ~\new_[6272]_ ;
  assign \new_[6188]_  = ~\new_[6389]_  | ~\new_[32333]_ ;
  assign \new_[6189]_  = \\s5_msel_arb2_state_reg[2] ;
  assign \new_[6190]_  = \\s5_msel_arb2_state_reg[0] ;
  assign \new_[6191]_  = \\s4_msel_arb1_state_reg[2] ;
  assign \new_[6192]_  = \\s4_msel_arb3_state_reg[1] ;
  assign \new_[6193]_  = \\s4_msel_arb0_state_reg[2] ;
  assign \new_[6194]_  = \\s3_msel_arb1_state_reg[2] ;
  assign \new_[6195]_  = \\s1_msel_arb3_state_reg[2] ;
  assign \new_[6196]_  = \\s1_msel_arb1_state_reg[0] ;
  assign \new_[6197]_  = \\s1_msel_arb1_state_reg[2] ;
  assign \new_[6198]_  = ~\new_[32333]_  | ~\new_[6373]_ ;
  assign \new_[6199]_  = \\s13_msel_arb1_state_reg[2] ;
  assign \new_[6200]_  = \\s13_msel_arb3_state_reg[2] ;
  assign \new_[6201]_  = ~s15_we_o | ~\new_[31931]_ ;
  assign \new_[6202]_  = \\s10_msel_arb0_state_reg[2] ;
  assign \new_[6203]_  = \\s10_msel_arb3_state_reg[2] ;
  assign \new_[6204]_  = \\s12_msel_arb3_state_reg[0] ;
  assign \new_[6205]_  = \\s12_msel_arb3_state_reg[2] ;
  assign \new_[6206]_  = \\s13_msel_arb3_state_reg[0] ;
  assign \new_[6207]_  = \\s14_msel_arb1_state_reg[0] ;
  assign \new_[6208]_  = \\s15_msel_arb1_state_reg[2] ;
  assign \new_[6209]_  = \\s15_msel_arb3_state_reg[2] ;
  assign \new_[6210]_  = \\s2_msel_arb1_state_reg[0] ;
  assign \new_[6211]_  = \\s2_msel_arb1_state_reg[2] ;
  assign \new_[6212]_  = \\s3_msel_arb3_state_reg[0] ;
  assign \new_[6213]_  = \\s3_msel_arb3_state_reg[2] ;
  assign \new_[6214]_  = \\s4_msel_arb3_state_reg[2] ;
  assign \new_[6215]_  = \\s9_msel_arb1_state_reg[1] ;
  assign \new_[6216]_  = \\s0_msel_arb1_state_reg[0] ;
  assign \new_[6217]_  = \\s0_msel_arb3_state_reg[1] ;
  assign n6719 = ~\new_[7873]_  | ~\new_[7453]_  | ~\new_[8311]_  | ~\new_[6615]_ ;
  assign n6884 = ~\new_[7881]_  | ~\new_[7205]_  | ~\new_[8351]_  | ~\new_[6619]_ ;
  assign n6814 = ~\new_[7216]_  | ~\new_[8220]_  | ~\new_[8746]_  | ~\new_[7245]_ ;
  assign \new_[6221]_  = ~\new_[6287]_ ;
  assign \new_[6222]_  = ~\new_[32289]_ ;
  assign \new_[6223]_  = \new_[32289]_ ;
  assign n6674 = ~\new_[9827]_  | ~\new_[8834]_  | ~\new_[8510]_  | ~\new_[6602]_ ;
  assign n6694 = ~\new_[11499]_  | ~\new_[9834]_  | ~\new_[9404]_  | ~\new_[6603]_ ;
  assign n6739 = ~\new_[8675]_  | ~\new_[7428]_  | ~\new_[8727]_  | ~\new_[6616]_ ;
  assign n6744 = ~\new_[8066]_  | ~\new_[7266]_  | ~\new_[8010]_  | ~\new_[7303]_ ;
  assign n6749 = ~\new_[9841]_  | ~\new_[9842]_  | ~\new_[9448]_  | ~\new_[6605]_ ;
  assign n6769 = ~\new_[8069]_  | ~\new_[7267]_  | ~\new_[8015]_  | ~\new_[7308]_ ;
  assign n6759 = ~\new_[8839]_  | ~\new_[8840]_  | ~\new_[9458]_  | ~\new_[6606]_ ;
  assign n6779 = ~\new_[9846]_  | ~\new_[9847]_  | ~\new_[9461]_  | ~\new_[6607]_ ;
  assign n6809 = ~\new_[8843]_  | ~\new_[9853]_  | ~\new_[8552]_  | ~\new_[6608]_ ;
  assign n6824 = ~\new_[9854]_  | ~\new_[8844]_  | ~\new_[9481]_  | ~\new_[6609]_ ;
  assign n6834 = ~\new_[8845]_  | ~\new_[8846]_  | ~\new_[8553]_  | ~\new_[6610]_ ;
  assign n6839 = ~\new_[9855]_  | ~\new_[9856]_  | ~\new_[8558]_  | ~\new_[6611]_ ;
  assign n6849 = ~\new_[8848]_  | ~\new_[8847]_  | ~\new_[8560]_  | ~\new_[6612]_ ;
  assign n6859 = ~\new_[8849]_  | ~\new_[9857]_  | ~\new_[8561]_  | ~\new_[6613]_ ;
  assign n6864 = ~\new_[8077]_  | ~\new_[7268]_  | ~\new_[8041]_  | ~\new_[7344]_ ;
  assign n6874 = ~\new_[8079]_  | ~\new_[7269]_  | ~\new_[8040]_  | ~\new_[7355]_ ;
  assign n6889 = ~\new_[13464]_  | ~\new_[9863]_  | ~\new_[8571]_  | ~\new_[6614]_ ;
  assign n6794 = ~\new_[8188]_  | ~\new_[7215]_  | ~\new_[7890]_  | ~\new_[6617]_ ;
  assign n6869 = ~\new_[8700]_  | ~\new_[7880]_  | ~\new_[8347]_  | ~\new_[6618]_ ;
  assign n6724 = ~\new_[6604]_  | ~\new_[8004]_  | ~\new_[8002]_ ;
  assign n6734 = ~\new_[7951]_  | ~\new_[7273]_  | ~\new_[8008]_  | ~\new_[7302]_ ;
  assign \new_[6245]_  = \\s10_msel_arb3_state_reg[1] ;
  assign \new_[6246]_  = \\s10_msel_arb3_state_reg[0] ;
  assign n6669 = ~\new_[7362]_  | ~\new_[8498]_  | ~\new_[7281]_  | ~\new_[9389]_ ;
  assign n6679 = ~\new_[7363]_  | ~\new_[7971]_  | ~\new_[7991]_  | ~\new_[8477]_ ;
  assign n6684 = ~\new_[7365]_  | ~\new_[7270]_  | ~\new_[7285]_  | ~\new_[8478]_ ;
  assign n6699 = ~\new_[7366]_  | ~\new_[7972]_  | ~\new_[7994]_  | ~\new_[8479]_ ;
  assign n6709 = ~\new_[7271]_  | ~\new_[7367]_  | ~\new_[7295]_  | ~\new_[8481]_ ;
  assign n6714 = ~\new_[7272]_  | ~\new_[7369]_  | ~\new_[6637]_  | ~\new_[8483]_ ;
  assign n6754 = ~\new_[7370]_  | ~\new_[7975]_  | ~\new_[8014]_  | ~\new_[8485]_ ;
  assign n6764 = ~\new_[7274]_  | ~\new_[7372]_  | ~\new_[7311]_  | ~\new_[8487]_ ;
  assign n6784 = ~\new_[7373]_  | ~\new_[7978]_  | ~\new_[8024]_  | ~\new_[8489]_ ;
  assign n6789 = ~\new_[8575]_  | ~\new_[7275]_  | ~\new_[7317]_  | ~\new_[8490]_ ;
  assign n6804 = ~\new_[7374]_  | ~\new_[7979]_  | ~\new_[7326]_  | ~\new_[8492]_ ;
  assign n6819 = ~\new_[7375]_  | ~\new_[7980]_  | ~\new_[7333]_  | ~\new_[8494]_ ;
  assign n6829 = ~\new_[7981]_  | ~\new_[7376]_  | ~\new_[7334]_  | ~\new_[7964]_ ;
  assign n6844 = ~\new_[7377]_  | ~\new_[7982]_  | ~\new_[8033]_  | ~\new_[8495]_ ;
  assign n6854 = ~\new_[7378]_  | ~\new_[7278]_  | ~\new_[8036]_  | ~\new_[7967]_ ;
  assign n6879 = ~\new_[7379]_  | ~\new_[7985]_  | ~\new_[7359]_  | ~\new_[8497]_ ;
  assign n6689 = ~\new_[8511]_  | ~\new_[7382]_  | ~\new_[7289]_  | ~\new_[8512]_ ;
  assign n6704 = ~\new_[7384]_  | ~\new_[7293]_  | ~\new_[7294]_  | ~\new_[7996]_ ;
  assign n6729 = ~\new_[7386]_  | ~\new_[8528]_  | ~\new_[8529]_  | ~\new_[7299]_ ;
  assign n6774 = ~\new_[8071]_  | ~\new_[7315]_  | ~\new_[7316]_  | ~\new_[8022]_ ;
  assign n6799 = ~\new_[7323]_  | ~\new_[7390]_  | ~\new_[7325]_  | ~\new_[7324]_ ;
  assign \new_[6268]_  = \\s6_msel_arb3_state_reg[2] ;
  assign \new_[6269]_  = \\s7_msel_arb3_state_reg[0] ;
  assign \new_[6270]_  = \\s7_msel_arb1_state_reg[1] ;
  assign \new_[6271]_  = \\s15_msel_arb0_state_reg[2] ;
  assign \new_[6272]_  = ~\new_[6391]_  | ~\new_[6374]_ ;
  assign \new_[6273]_  = \\s2_msel_arb3_state_reg[2] ;
  assign \new_[6274]_  = s15_next_reg;
  assign n6924 = ~\new_[9628]_  | ~\new_[7431]_  | ~\new_[8296]_  | ~\new_[7254]_ ;
  assign n7079 = ~\new_[7876]_  | ~\new_[8176]_  | ~\new_[8324]_  | ~\new_[7243]_ ;
  assign n7124 = ~\new_[7877]_  | ~\new_[7798]_  | ~\new_[8335]_  | ~\new_[7246]_ ;
  assign n7244 = ~\new_[7879]_  | ~\new_[7822]_  | ~\new_[7896]_  | ~\new_[7249]_ ;
  assign n6934 = ~\new_[7448]_  | ~\new_[7432]_  | ~\new_[8298]_  | ~\new_[7236]_ ;
  assign n6944 = ~\new_[7870]_  | ~\new_[8133]_  | ~\new_[9692]_  | ~\new_[7940]_ ;
  assign n7004 = ~\new_[8283]_  | ~\new_[8140]_  | ~\new_[8721]_  | ~\new_[7239]_ ;
  assign n7029 = ~\new_[7874]_  | ~\new_[8156]_  | ~\new_[8315]_  | ~\new_[7240]_ ;
  assign n7284 = ~\new_[8284]_  | ~\new_[8161]_  | ~\new_[8731]_  | ~\new_[7241]_ ;
  assign n7254 = ~\new_[8288]_  | ~\new_[7734]_  | ~\new_[7892]_  | ~\new_[7244]_ ;
  assign n7149 = ~\new_[8289]_  | ~\new_[8225]_  | ~\new_[9739]_  | ~\new_[7248]_ ;
  assign n7169 = ~\new_[8290]_  | ~\new_[8259]_  | ~\new_[8760]_  | ~\new_[7250]_ ;
  assign \new_[6287]_  = ~\new_[32331]_ ;
  assign n7214 = ~\new_[8704]_  | ~\new_[8469]_  | ~\new_[9753]_  | ~\new_[7252]_ ;
  assign n7224 = ~\new_[8706]_  | ~\new_[9823]_  | ~\new_[9681]_  | ~\new_[7253]_ ;
  assign n6954 = ~\new_[8712]_  | ~\new_[9636]_  | ~\new_[8713]_  | ~\new_[7255]_ ;
  assign n6984 = ~\new_[9649]_  | ~\new_[8672]_  | ~\new_[9703]_  | ~\new_[7256]_ ;
  assign n7294 = ~\new_[9657]_  | ~\new_[8677]_  | ~\new_[9710]_  | ~\new_[7257]_ ;
  assign n7279 = ~\new_[8969]_  | ~\new_[8449]_  | ~\new_[8322]_  | ~\new_[7258]_ ;
  assign n7264 = ~\new_[9663]_  | ~\new_[8682]_  | ~\new_[9722]_  | ~\new_[7259]_ ;
  assign n7104 = ~\new_[8327]_  | ~\new_[9665]_  | ~\new_[8744]_  | ~\new_[7260]_ ;
  assign n7119 = ~\new_[8749]_  | ~\new_[8223]_  | ~\new_[8332]_  | ~\new_[7261]_ ;
  assign n7134 = ~\new_[8755]_  | ~\new_[9667]_  | ~\new_[9734]_  | ~\new_[7262]_ ;
  assign n7249 = ~\new_[8341]_  | ~\new_[8692]_  | ~\new_[8758]_  | ~\new_[7263]_ ;
  assign n7184 = ~\new_[9746]_  | ~\new_[9669]_  | ~\new_[9747]_  | ~\new_[7264]_ ;
  assign n7204 = ~\new_[8766]_  | ~\new_[8747]_  | ~\new_[9750]_  | ~\new_[7265]_ ;
  assign n6904 = ~\new_[8060]_  | ~\new_[7986]_  | ~\new_[9395]_  | ~\new_[7280]_ ;
  assign n6939 = ~\new_[8061]_  | ~\new_[7989]_  | ~\new_[7990]_  | ~\new_[7283]_ ;
  assign n6929 = ~\new_[11495]_  | ~\new_[9832]_  | ~\new_[9397]_  | ~\new_[7227]_ ;
  assign n7229 = ~\new_[9833]_  | ~\new_[11497]_  | ~\new_[9398]_  | ~\new_[7228]_ ;
  assign n6899 = ~\new_[8062]_  | ~\new_[7993]_  | ~\new_[7288]_  | ~\new_[7287]_ ;
  assign n7219 = ~\new_[8063]_  | ~\new_[7995]_  | ~\new_[7292]_  | ~\new_[8513]_ ;
  assign n6894 = ~\new_[8838]_  | ~\new_[9840]_  | ~\new_[9420]_  | ~\new_[7229]_ ;
  assign n7009 = ~\new_[8065]_  | ~\new_[8526]_  | ~\new_[8527]_  | ~\new_[8005]_ ;
  assign n7014 = ~\new_[7230]_  | ~\new_[9434]_  | ~\new_[8530]_ ;
  assign n7289 = ~\new_[8067]_  | ~\new_[8011]_  | ~\new_[8536]_  | ~\new_[7305]_ ;
  assign n7034 = ~\new_[9843]_  | ~\new_[9844]_  | ~\new_[9452]_  | ~\new_[7231]_ ;
  assign n7059 = ~\new_[8841]_  | ~\new_[9845]_  | ~\new_[10991]_  | ~\new_[7232]_ ;
  assign n7069 = ~\new_[8070]_  | ~\new_[8021]_  | ~\new_[7314]_  | ~\new_[7313]_ ;
  assign n7084 = ~\new_[8072]_  | ~\new_[8025]_  | ~\new_[8548]_  | ~\new_[7319]_ ;
  assign n7094 = ~\new_[11521]_  | ~\new_[9851]_  | ~\new_[9471]_  | ~\new_[7233]_ ;
  assign n7099 = ~\new_[8074]_  | ~\new_[8029]_  | ~\new_[7322]_  | ~\new_[7321]_ ;
  assign n7259 = ~\new_[9852]_  | ~\new_[8842]_  | ~\new_[9475]_  | ~\new_[7234]_ ;
  assign n7129 = ~\new_[8075]_  | ~\new_[8032]_  | ~\new_[8554]_  | ~\new_[7338]_ ;
  assign n7159 = ~\new_[8076]_  | ~\new_[8034]_  | ~\new_[8035]_  | ~\new_[7340]_ ;
  assign n7239 = ~\new_[8078]_  | ~\new_[8562]_  | ~\new_[8563]_  | ~\new_[8037]_ ;
  assign n7209 = ~\new_[8081]_  | ~\new_[7953]_  | ~\new_[8050]_  | ~\new_[7361]_ ;
  assign n6914 = ~\new_[8664]_  | ~\new_[7445]_  | ~\new_[8294]_  | ~\new_[7235]_ ;
  assign n6959 = ~\new_[8668]_  | ~\new_[7871]_  | ~\new_[8302]_  | ~\new_[7237]_ ;
  assign n6974 = ~\new_[8671]_  | ~\new_[7872]_  | ~\new_[8308]_  | ~\new_[7238]_ ;
  assign n7054 = ~\new_[8681]_  | ~\new_[7875]_  | ~\new_[8320]_  | ~\new_[7242]_ ;
  assign n7144 = ~\new_[8685]_  | ~\new_[7878]_  | ~\new_[8339]_  | ~\new_[7247]_ ;
  assign n7234 = ~\new_[9671]_  | ~\new_[8291]_  | ~\new_[9748]_  | ~\new_[7251]_ ;
  assign n6919 = ~\new_[8132]_  | ~\new_[7954]_  | ~\new_[7430]_  | ~\new_[7429]_ ;
  assign n6949 = ~\new_[8134]_  | ~\new_[7955]_  | ~\new_[7441]_  | ~\new_[7438]_ ;
  assign n6964 = ~\new_[8137]_  | ~\new_[7956]_  | ~\new_[7447]_  | ~\new_[7446]_ ;
  assign n6994 = ~\new_[7450]_  | ~\new_[7957]_  | ~\new_[7451]_  | ~\new_[7449]_ ;
  assign n7019 = ~\new_[8146]_  | ~\new_[7958]_  | ~\new_[8676]_  | ~\new_[9334]_ ;
  assign n7049 = ~\new_[8172]_  | ~\new_[7959]_  | ~\new_[9659]_  | ~\new_[8679]_ ;
  assign n7074 = ~\new_[7599]_  | ~\new_[7960]_  | ~\new_[7603]_  | ~\new_[7595]_ ;
  assign n7274 = ~\new_[7653]_  | ~\new_[7961]_  | ~\new_[7656]_  | ~\new_[7646]_ ;
  assign n7109 = ~\new_[8219]_  | ~\new_[7962]_  | ~\new_[7715]_  | ~\new_[7699]_ ;
  assign n7114 = ~\new_[7777]_  | ~\new_[7963]_  | ~\new_[7780]_  | ~\new_[7769]_ ;
  assign n7139 = ~\new_[7800]_  | ~\new_[7965]_  | ~\new_[8670]_  | ~\new_[8684]_ ;
  assign n7154 = ~\new_[8235]_  | ~\new_[7966]_  | ~\new_[7807]_  | ~\new_[7802]_ ;
  assign n7174 = ~\new_[8268]_  | ~\new_[7969]_  | ~\new_[8699]_  | ~\new_[8698]_ ;
  assign n7194 = ~\new_[8279]_  | ~\new_[7970]_  | ~\new_[9673]_  | ~\new_[8701]_ ;
  assign n6969 = ~\new_[7973]_  | ~\new_[8051]_  | ~\new_[7290]_  | ~\new_[8480]_ ;
  assign n6979 = ~\new_[8501]_  | ~\new_[8052]_  | ~\new_[7296]_  | ~\new_[8482]_ ;
  assign n6999 = ~\new_[8053]_  | ~\new_[7974]_  | ~\new_[8001]_  | ~\new_[8484]_ ;
  assign n7039 = ~\new_[8054]_  | ~\new_[7976]_  | ~\new_[8541]_  | ~\new_[8486]_ ;
  assign n7064 = ~\new_[7977]_  | ~\new_[8055]_  | ~\new_[8020]_  | ~\new_[8488]_ ;
  assign n7269 = ~\new_[8056]_  | ~\new_[8505]_  | ~\new_[8028]_  | ~\new_[9391]_ ;
  assign n7164 = ~\new_[8506]_  | ~\new_[8057]_  | ~\new_[8559]_  | ~\new_[9392]_ ;
  assign n7179 = ~\new_[8058]_  | ~\new_[7983]_  | ~\new_[7346]_  | ~\new_[8496]_ ;
  assign n7189 = ~\new_[7984]_  | ~\new_[8059]_  | ~\new_[7347]_  | ~\new_[9393]_ ;
  assign n6909 = ~\new_[8587]_  | ~\new_[7987]_  | ~\new_[8509]_  | ~\new_[8508]_ ;
  assign n6989 = ~\new_[8064]_  | ~\new_[7998]_  | ~\new_[8522]_  | ~\new_[7999]_ ;
  assign n7024 = ~\new_[8068]_  | ~\new_[8537]_  | ~\new_[8538]_  | ~\new_[8013]_ ;
  assign n7044 = ~\new_[9523]_  | ~\new_[8017]_  | ~\new_[8544]_  | ~\new_[9457]_ ;
  assign n7089 = ~\new_[8073]_  | ~\new_[8549]_  | ~\new_[8550]_  | ~\new_[8026]_ ;
  assign n7199 = ~\new_[8043]_  | ~\new_[8080]_  | ~\new_[8570]_  | ~\new_[8045]_ ;
  assign \new_[6357]_  = ~\new_[8086]_  & ~\new_[6724]_ ;
  assign \new_[6358]_  = ~\new_[6584]_  & ~\new_[8404]_ ;
  assign \new_[6359]_  = ~\new_[6585]_  & ~\new_[8405]_ ;
  assign \new_[6360]_  = ~\new_[6586]_  & ~\new_[11650]_ ;
  assign \new_[6361]_  = ~\new_[6587]_  & ~\new_[8424]_ ;
  assign \new_[6362]_  = ~\new_[6588]_  & ~\new_[8427]_ ;
  assign \new_[6363]_  = ~\new_[6589]_  & ~\new_[9864]_ ;
  assign \new_[6364]_  = ~\new_[20287]_  | ~\new_[11912]_  | ~\new_[6590]_  | ~\new_[8808]_ ;
  assign \new_[6365]_  = ~\new_[20294]_  | ~\new_[11916]_  | ~\new_[6591]_  | ~\new_[8809]_ ;
  assign \new_[6366]_  = ~\new_[20304]_  | ~\new_[11922]_  | ~\new_[6592]_  | ~\new_[8810]_ ;
  assign \new_[6367]_  = ~\new_[18386]_  | ~\new_[9109]_  | ~\new_[6593]_  | ~\new_[8370]_ ;
  assign \new_[6368]_  = ~\new_[18392]_  | ~\new_[9135]_  | ~\new_[6594]_  | ~\new_[8374]_ ;
  assign \new_[6369]_  = ~\new_[19340]_  | ~\new_[9142]_  | ~\new_[6595]_  | ~\new_[8821]_ ;
  assign \new_[6370]_  = ~\new_[20345]_  | ~\new_[11946]_  | ~\new_[6596]_  | ~\new_[8823]_ ;
  assign \new_[6371]_  = ~\new_[20314]_  | ~\new_[9157]_  | ~\new_[6597]_  | ~\new_[8824]_ ;
  assign \new_[6372]_  = ~\new_[20319]_  | ~\new_[11960]_  | ~\new_[6598]_  | ~\new_[8827]_ ;
  assign \new_[6373]_  = ~\new_[6434]_ ;
  assign \new_[6374]_  = ~\new_[6435]_ ;
  assign \new_[6375]_  = \\s13_msel_pri_out_reg[0] ;
  assign \new_[6376]_  = \\s3_msel_pri_out_reg[0] ;
  assign n7344 = ~\new_[8660]_  | ~\new_[8145]_  | ~\new_[9709]_  | ~\new_[7944]_ ;
  assign n7339 = ~\new_[9655]_  | ~\new_[8144]_  | ~\new_[8725]_  | ~\new_[7943]_ ;
  assign s0_stb_o = \new_[8471]_  | \new_[7220]_ ;
  assign n7304 = ~\new_[8282]_  | ~\new_[9644]_  | ~\new_[9700]_  | ~\new_[7942]_ ;
  assign n7419 = ~\new_[8285]_  | ~\new_[8173]_  | ~\new_[8736]_  | ~\new_[7945]_ ;
  assign n7369 = ~\new_[8287]_  | ~\new_[8197]_  | ~\new_[9724]_  | ~\new_[7947]_ ;
  assign n7314 = ~\new_[9674]_  | ~\new_[8131]_  | ~\new_[9684]_  | ~\new_[7939]_ ;
  assign n7324 = ~\new_[8281]_  | ~\new_[8136]_  | ~\new_[9697]_  | ~\new_[7941]_ ;
  assign s9_stb_o = \new_[7307]_  | \new_[8012]_ ;
  assign n7364 = ~\new_[8286]_  | ~\new_[8177]_  | ~\new_[9719]_  | ~\new_[7946]_ ;
  assign n7399 = ~\new_[8703]_  | ~\new_[8224]_  | ~\new_[8336]_  | ~\new_[7948]_ ;
  assign s12_stb_o = \new_[10978]_  | \new_[7310]_ ;
  assign \new_[6389]_  = ~\new_[6578]_ ;
  assign \new_[6390]_  = ~\new_[6578]_ ;
  assign \new_[6391]_  = ~\new_[6578]_ ;
  assign n7299 = ~\new_[8304]_  | ~\new_[8138]_  | ~\new_[8305]_  | ~\new_[7949]_ ;
  assign n7354 = ~\new_[8733]_  | ~\new_[8680]_  | ~\new_[9714]_  | ~\new_[7950]_ ;
  assign n7394 = ~\new_[9829]_  | ~\new_[9831]_  | ~\new_[10904]_  | ~\new_[7933]_ ;
  assign n7319 = ~\new_[8835]_  | ~\new_[11502]_  | ~\new_[10922]_  | ~\new_[7934]_ ;
  assign n7329 = ~\new_[8837]_  | ~\new_[9836]_  | ~\new_[10933]_  | ~\new_[7935]_ ;
  assign n7334 = ~\new_[8592]_  | ~\new_[8519]_  | ~\new_[8520]_  | ~\new_[7997]_ ;
  assign n7349 = ~\new_[8598]_  | ~\new_[8542]_  | ~\new_[9456]_  | ~\new_[8016]_ ;
  assign n7359 = ~\new_[9848]_  | ~\new_[11516]_  | ~\new_[11011]_  | ~\new_[7937]_ ;
  assign n7404 = ~\new_[11530]_  | ~\new_[11533]_  | ~\new_[11052]_  | ~\new_[7938]_ ;
  assign n7379 = ~\new_[8612]_  | ~\new_[8568]_  | ~\new_[8569]_  | ~\new_[8042]_ ;
  assign n7309 = ~\new_[8662]_  | ~\new_[8476]_  | ~\new_[8663]_  | ~\new_[8661]_ ;
  assign n7414 = ~\new_[8143]_  | ~\new_[8502]_  | ~\new_[8674]_  | ~\new_[8673]_ ;
  assign n7389 = ~\new_[8499]_  | ~\new_[8572]_  | ~\new_[7988]_  | ~\new_[9390]_ ;
  assign n7384 = ~\new_[8507]_  | ~\new_[8584]_  | ~\new_[8048]_  | ~\new_[9394]_ ;
  assign n7409 = ~\new_[8607]_  | ~\new_[8555]_  | ~\new_[8557]_  | ~\new_[8556]_ ;
  assign n7374 = ~\new_[8564]_  | ~\new_[8611]_  | ~\new_[8566]_  | ~\new_[8565]_ ;
  assign \s15_data_o[15]  = ~\new_[8574]_  | ~\new_[9502]_  | ~\new_[8573]_  | ~\new_[9501]_ ;
  assign \s15_data_o[14]  = ~\new_[8577]_  | ~\new_[9505]_  | ~\new_[9503]_  | ~\new_[8576]_ ;
  assign \s15_data_o[13]  = ~\new_[8579]_  | ~\new_[9507]_  | ~\new_[9506]_  | ~\new_[8578]_ ;
  assign \s15_data_o[12]  = ~\new_[8581]_  | ~\new_[9509]_  | ~\new_[9508]_  | ~\new_[8580]_ ;
  assign \s15_data_o[11]  = ~\new_[8583]_  | ~\new_[9511]_  | ~\new_[9510]_  | ~\new_[8582]_ ;
  assign \s15_data_o[10]  = ~\new_[8586]_  | ~\new_[9513]_  | ~\new_[9512]_  | ~\new_[8585]_ ;
  assign \s15_data_o[9]  = ~\new_[9515]_  | ~\new_[8589]_  | ~\new_[8588]_  | ~\new_[9514]_ ;
  assign \s15_data_o[8]  = ~\new_[8591]_  | ~\new_[9517]_  | ~\new_[8590]_  | ~\new_[9516]_ ;
  assign \s15_data_o[7]  = ~\new_[8594]_  | ~\new_[9519]_  | ~\new_[9518]_  | ~\new_[8593]_ ;
  assign \s15_data_o[6]  = ~\new_[8596]_  | ~\new_[9521]_  | ~\new_[9520]_  | ~\new_[8595]_ ;
  assign \s15_data_o[5]  = ~\new_[8599]_  | ~\new_[9524]_  | ~\new_[8597]_  | ~\new_[9522]_ ;
  assign \s15_data_o[4]  = ~\new_[8601]_  | ~\new_[9526]_  | ~\new_[9525]_  | ~\new_[8600]_ ;
  assign \s15_data_o[3]  = ~\new_[8603]_  | ~\new_[9528]_  | ~\new_[9527]_  | ~\new_[8602]_ ;
  assign \s15_data_o[2]  = ~\new_[8605]_  | ~\new_[9530]_  | ~\new_[9529]_  | ~\new_[8604]_ ;
  assign \s15_data_o[1]  = ~\new_[8608]_  | ~\new_[9532]_  | ~\new_[8606]_  | ~\new_[9531]_ ;
  assign \s15_data_o[0]  = ~\new_[8610]_  | ~\new_[9534]_  | ~\new_[8609]_  | ~\new_[9533]_ ;
  assign s15_we_o = ~\new_[8642]_  | ~\new_[9550]_  | ~\new_[9549]_  | ~\new_[8641]_ ;
  assign \new_[6425]_  = ~\new_[7400]_  & ~\new_[8617]_ ;
  assign \new_[6426]_  = ~\new_[7419]_  & ~\new_[7301]_ ;
  assign \new_[6427]_  = ~\new_[7406]_  & ~\new_[8627]_ ;
  assign \new_[6428]_  = ~\new_[7413]_  & ~\new_[8102]_ ;
  assign \new_[6429]_  = ~\new_[8634]_  & ~\new_[7414]_ ;
  assign \new_[6430]_  = ~\new_[8635]_  & ~\new_[7416]_ ;
  assign \new_[6431]_  = (~\new_[8851]_  | ~\m7_addr_i[31] ) & (~\new_[32346]_  | ~\m0_addr_i[31] );
  assign \new_[6432]_  = (~\new_[8851]_  | ~\new_[31885]_ ) & (~\new_[32346]_  | ~\new_[31292]_ );
  assign \new_[6433]_  = (~\new_[8851]_  | ~\new_[30577]_ ) & (~\new_[32346]_  | ~\new_[30957]_ );
  assign \new_[6434]_  = ~\s15_addr_o[2]  | ~\new_[7923]_ ;
  assign \new_[6435]_  = ~\s15_addr_o[4]  | ~\new_[32304]_ ;
  assign \new_[6436]_  = \\s11_msel_pri_out_reg[0] ;
  assign \new_[6437]_  = \\s12_msel_pri_out_reg[0] ;
  assign \new_[6438]_  = \\s5_msel_pri_out_reg[0] ;
  assign \new_[6439]_  = \\s6_msel_pri_out_reg[0] ;
  assign \new_[6440]_  = \\s8_msel_pri_out_reg[0] ;
  assign \new_[6441]_  = ~s12_next_reg;
  assign \new_[6442]_  = ~s13_next_reg;
  assign \new_[6443]_  = ~s14_next_reg;
  assign \new_[6444]_  = ~s3_next_reg;
  assign \new_[6445]_  = ~s6_next_reg;
  assign \new_[6446]_  = ~s9_next_reg;
  assign \new_[6447]_  = ~s8_next_reg;
  assign \new_[6448]_  = ~s0_next_reg;
  assign \new_[6449]_  = \\s8_msel_pri_out_reg[1] ;
  assign \s0_data_o[30]  = ~\new_[11992]_  | ~\new_[9214]_  | ~\new_[10374]_  | ~\new_[11986]_ ;
  assign \s0_data_o[25]  = ~\new_[9251]_  | ~\new_[12054]_  | ~\new_[12041]_  | ~\new_[12044]_ ;
  assign \s0_data_o[24]  = ~\new_[9255]_  | ~\new_[12060]_  | ~\new_[12055]_  | ~\new_[10439]_ ;
  assign \s0_data_o[19]  = ~\new_[13696]_  | ~\new_[9282]_  | ~\new_[10472]_  | ~\new_[10473]_ ;
  assign \s0_data_o[18]  = ~\new_[12099]_  | ~\new_[9284]_  | ~\new_[12096]_  | ~\new_[10474]_ ;
  assign \s0_data_o[17]  = ~\new_[13711]_  | ~\new_[9288]_  | ~\new_[12102]_  | ~\new_[10478]_ ;
  assign \s0_data_o[16]  = ~\new_[9290]_  | ~\new_[12118]_  | ~\new_[10480]_  | ~\new_[12116]_ ;
  assign \s0_data_o[15]  = ~\new_[12123]_  | ~\new_[9291]_  | ~\new_[10483]_  | ~\new_[12120]_ ;
  assign \s0_addr_o[31]  = ~\new_[12273]_  | ~\new_[9311]_  | ~\new_[13817]_  | ~\new_[12272]_ ;
  assign \s0_addr_o[30]  = ~\new_[10539]_  | ~\new_[9504]_  | ~\new_[12277]_  | ~\new_[13142]_ ;
  assign \s0_addr_o[27]  = ~\new_[12294]_  | ~\new_[9315]_  | ~\new_[12292]_  | ~\new_[13839]_ ;
  assign \s0_addr_o[26]  = ~\new_[12297]_  | ~\new_[9316]_  | ~\new_[13840]_  | ~\new_[12296]_ ;
  assign \s0_addr_o[23]  = ~\new_[11822]_  | ~\new_[9319]_  | ~\new_[12314]_  | ~\new_[10550]_ ;
  assign \s0_addr_o[21]  = ~\new_[11670]_  | ~\new_[9320]_  | ~\new_[12337]_  | ~\new_[12339]_ ;
  assign \s0_addr_o[18]  = ~\new_[13892]_  | ~\new_[9321]_  | ~\new_[9967]_  | ~\new_[12360]_ ;
  assign \s0_addr_o[17]  = ~\new_[12368]_  | ~\new_[9322]_  | ~\new_[10574]_  | ~\new_[12366]_ ;
  assign \s0_addr_o[16]  = ~\new_[9323]_  | ~\new_[12377]_  | ~\new_[10578]_  | ~\new_[12375]_ ;
  assign \s0_addr_o[15]  = ~\new_[13922]_  | ~\new_[8678]_  | ~\new_[12379]_  | ~\new_[10583]_ ;
  assign \s0_addr_o[10]  = ~\new_[13963]_  | ~\new_[9333]_  | ~\new_[12423]_  | ~\new_[9629]_ ;
  assign \s0_addr_o[7]  = ~\new_[13980]_  | ~\new_[9335]_  | ~\new_[12447]_  | ~\new_[10606]_ ;
  assign \s0_addr_o[6]  = ~\new_[13984]_  | ~\new_[9336]_  | ~\new_[12456]_  | ~\new_[10614]_ ;
  assign \s0_addr_o[5]  = ~\new_[12469]_  | ~\new_[8659]_  | ~\new_[10616]_  | ~\new_[10617]_ ;
  assign \s0_addr_o[4]  = ~\new_[12481]_  | ~\new_[9337]_  | ~\new_[10620]_  | ~\new_[12479]_ ;
  assign \s0_addr_o[0]  = ~\new_[14007]_  | ~\new_[9340]_  | ~\new_[10052]_  | ~\new_[10637]_ ;
  assign \s0_sel_o[3]  = ~\new_[13459]_  | ~\new_[9344]_  | ~\new_[10641]_  | ~\new_[10642]_ ;
  assign \s0_sel_o[2]  = ~\new_[14017]_  | ~\new_[9346]_  | ~\new_[10645]_  | ~\new_[10647]_ ;
  assign \s0_sel_o[0]  = ~\new_[14029]_  | ~\new_[9350]_  | ~\new_[9991]_  | ~\new_[10660]_ ;
  assign s0_we_o = ~\new_[14034]_  | ~\new_[9355]_  | ~\new_[10663]_  | ~\new_[10666]_ ;
  assign s3_stb_o = \new_[8023]_  | \new_[9462]_ ;
  assign s7_stb_o = \new_[9425]_  | \new_[8006]_ ;
  assign \s8_data_o[31]  = ~\new_[8958]_  | ~\new_[11809]_  | ~\new_[10054]_  | ~\new_[8956]_ ;
  assign \s8_data_o[30]  = ~\new_[8963]_  | ~\new_[10056]_  | ~\new_[10055]_  | ~\new_[8961]_ ;
  assign \s8_data_o[28]  = ~\new_[8966]_  | ~\new_[10065]_  | ~\new_[11811]_  | ~\new_[10064]_ ;
  assign \s8_data_o[26]  = ~\new_[8971]_  | ~\new_[11813]_  | ~\new_[10071]_  | ~\new_[8970]_ ;
  assign \s8_data_o[24]  = ~\new_[8976]_  | ~\new_[11815]_  | ~\new_[8974]_  | ~\new_[8975]_ ;
  assign \s8_data_o[22]  = ~\new_[8979]_  | ~\new_[10084]_  | ~\new_[11818]_  | ~\new_[8978]_ ;
  assign \s8_data_o[21]  = ~\new_[8981]_  | ~\new_[10086]_  | ~\new_[10085]_  | ~\new_[8980]_ ;
  assign \s8_data_o[20]  = ~\new_[8983]_  | ~\new_[10090]_  | ~\new_[10089]_  | ~\new_[8982]_ ;
  assign \s8_data_o[19]  = ~\new_[8985]_  | ~\new_[10092]_  | ~\new_[11829]_  | ~\new_[8984]_ ;
  assign \s8_data_o[18]  = ~\new_[8989]_  | ~\new_[11832]_  | ~\new_[8987]_  | ~\new_[8988]_ ;
  assign \s8_data_o[14]  = ~\new_[9000]_  | ~\new_[10104]_  | ~\new_[11837]_  | ~\new_[10103]_ ;
  assign \s8_data_o[8]  = ~\new_[9008]_  | ~\new_[11855]_  | ~\new_[9007]_  | ~\new_[10126]_ ;
  assign \s8_data_o[4]  = ~\new_[9018]_  | ~\new_[11864]_  | ~\new_[9016]_  | ~\new_[9017]_ ;
  assign \s8_data_o[3]  = ~\new_[9021]_  | ~\new_[10143]_  | ~\new_[11866]_  | ~\new_[9020]_ ;
  assign \s8_data_o[1]  = ~\new_[9025]_  | ~\new_[11873]_  | ~\new_[9023]_  | ~\new_[9024]_ ;
  assign \s8_data_o[0]  = ~\new_[9032]_  | ~\new_[10148]_  | ~\new_[9028]_  | ~\new_[9029]_ ;
  assign \s8_addr_o[31]  = ~\new_[9033]_  | ~\new_[9035]_  | ~\new_[11874]_  | ~\new_[9034]_ ;
  assign \s8_addr_o[30]  = ~\new_[11877]_  | ~\new_[9039]_  | ~\new_[10149]_  | ~\new_[9038]_ ;
  assign \s8_addr_o[29]  = ~\new_[9042]_  | ~\new_[10152]_  | ~\new_[10151]_  | ~\new_[9041]_ ;
  assign \s8_addr_o[28]  = ~\new_[11882]_  | ~\new_[9046]_  | ~\new_[10153]_  | ~\new_[9043]_ ;
  assign \s8_addr_o[27]  = ~\new_[11883]_  | ~\new_[9050]_  | ~\new_[10154]_  | ~\new_[10155]_ ;
  assign \s8_addr_o[26]  = ~\new_[9053]_  | ~\new_[9051]_  | ~\new_[11886]_  | ~\new_[10156]_ ;
  assign \s8_addr_o[25]  = ~\new_[11888]_  | ~\new_[9057]_  | ~\new_[10157]_  | ~\new_[10158]_ ;
  assign \s8_addr_o[24]  = ~\new_[9060]_  | ~\new_[10162]_  | ~\new_[9058]_  | ~\new_[9059]_ ;
  assign \s8_addr_o[23]  = ~\new_[9064]_  | ~\new_[10163]_  | ~\new_[11891]_  | ~\new_[9062]_ ;
  assign \s8_addr_o[22]  = ~\new_[9066]_  | ~\new_[10165]_  | ~\new_[10164]_  | ~\new_[9065]_ ;
  assign \s8_addr_o[20]  = ~\new_[9072]_  | ~\new_[9073]_  | ~\new_[10171]_  | ~\new_[10173]_ ;
  assign \s8_addr_o[19]  = ~\new_[9076]_  | ~\new_[10179]_  | ~\new_[10175]_  | ~\new_[9075]_ ;
  assign \s8_addr_o[17]  = ~\new_[9080]_  | ~\new_[10190]_  | ~\new_[11899]_  | ~\new_[9079]_ ;
  assign \s8_addr_o[15]  = ~\new_[9083]_  | ~\new_[10198]_  | ~\new_[11903]_  | ~\new_[9082]_ ;
  assign \s8_addr_o[12]  = ~\new_[9088]_  | ~\new_[11910]_  | ~\new_[10209]_  | ~\new_[9087]_ ;
  assign \s8_addr_o[8]  = ~\new_[10221]_  | ~\new_[9097]_  | ~\new_[10184]_  | ~\new_[10219]_ ;
  assign \s8_addr_o[4]  = ~\new_[9104]_  | ~\new_[10233]_  | ~\new_[11920]_  | ~\new_[10232]_ ;
  assign \s8_addr_o[2]  = ~\new_[11926]_  | ~\new_[9107]_  | ~\new_[10239]_  | ~\new_[10240]_ ;
  assign \s8_addr_o[0]  = ~\new_[9112]_  | ~\new_[10246]_  | ~\new_[11927]_  | ~\new_[9111]_ ;
  assign \s8_sel_o[3]  = ~\new_[9115]_  | ~\new_[11930]_  | ~\new_[9114]_  | ~\new_[10247]_ ;
  assign \s8_sel_o[2]  = ~\new_[9119]_  | ~\new_[11931]_  | ~\new_[9117]_  | ~\new_[9118]_ ;
  assign \s8_sel_o[0]  = ~\new_[9125]_  | ~\new_[10254]_  | ~\new_[11933]_  | ~\new_[9124]_ ;
  assign s8_stb_o = \new_[8532]_  | \new_[8009]_ ;
  assign \s9_data_o[31]  = ~\new_[9128]_  | ~\new_[10259]_  | ~\new_[8754]_  | ~\new_[10258]_ ;
  assign \s9_data_o[30]  = ~\new_[10263]_  | ~\new_[9130]_  | ~\new_[10260]_  | ~\new_[10261]_ ;
  assign \s9_data_o[26]  = ~\new_[11938]_  | ~\new_[9136]_  | ~\new_[10279]_  | ~\new_[9134]_ ;
  assign \s9_data_o[25]  = ~\new_[9139]_  | ~\new_[10283]_  | ~\new_[10281]_  | ~\new_[9138]_ ;
  assign \s9_data_o[24]  = ~\new_[9140]_  | ~\new_[10287]_  | ~\new_[10285]_  | ~\new_[10284]_ ;
  assign \s9_data_o[22]  = ~\new_[9141]_  | ~\new_[10293]_  | ~\new_[10291]_  | ~\new_[10292]_ ;
  assign \s9_data_o[20]  = ~\new_[9147]_  | ~\new_[10297]_  | ~\new_[9146]_  | ~\new_[10296]_ ;
  assign \s9_data_o[18]  = ~\new_[10303]_  | ~\new_[9151]_  | ~\new_[9149]_  | ~\new_[10302]_ ;
  assign \s9_data_o[17]  = ~\new_[10307]_  | ~\new_[9152]_  | ~\new_[10304]_  | ~\new_[10305]_ ;
  assign \s9_data_o[14]  = ~\new_[9156]_  | ~\new_[10317]_  | ~\new_[10315]_  | ~\new_[10316]_ ;
  assign \s9_data_o[6]  = ~\new_[10339]_  | ~\new_[9172]_  | ~\new_[9171]_  | ~\new_[10337]_ ;
  assign \s9_data_o[5]  = ~\new_[10342]_  | ~\new_[9175]_  | ~\new_[9173]_  | ~\new_[9174]_ ;
  assign \s9_data_o[3]  = ~\new_[9182]_  | ~\new_[9183]_  | ~\new_[10345]_  | ~\new_[9179]_ ;
  assign \s9_data_o[1]  = ~\new_[9187]_  | ~\new_[10350]_  | ~\new_[9186]_  | ~\new_[10665]_ ;
  assign \s9_addr_o[30]  = ~\new_[9193]_  | ~\new_[9194]_  | ~\new_[10363]_  | ~\new_[9192]_ ;
  assign \s9_addr_o[28]  = ~\new_[11970]_  | ~\new_[9200]_  | ~\new_[10367]_  | ~\new_[10369]_ ;
  assign \s9_addr_o[27]  = ~\new_[10371]_  | ~\new_[9204]_  | ~\new_[9201]_  | ~\new_[9202]_ ;
  assign \s9_addr_o[25]  = ~\new_[9208]_  | ~\new_[10375]_  | ~\new_[9207]_  | ~\new_[10373]_ ;
  assign \s9_addr_o[24]  = ~\new_[9210]_  | ~\new_[13657]_  | ~\new_[9209]_  | ~\new_[10376]_ ;
  assign \s9_addr_o[21]  = ~\new_[10387]_  | ~\new_[9223]_  | ~\new_[10385]_  | ~\new_[10386]_ ;
  assign \s9_addr_o[19]  = ~\new_[9226]_  | ~\new_[9227]_  | ~\new_[10391]_  | ~\new_[10393]_ ;
  assign \s9_addr_o[15]  = ~\new_[12021]_  | ~\new_[9234]_  | ~\new_[10408]_  | ~\new_[9233]_ ;
  assign \s9_addr_o[14]  = ~\new_[10411]_  | ~\new_[9236]_  | ~\new_[10409]_  | ~\new_[9235]_ ;
  assign \s9_addr_o[13]  = ~\new_[9238]_  | ~\new_[12029]_  | ~\new_[9237]_  | ~\new_[10415]_ ;
  assign \s9_addr_o[12]  = ~\new_[14960]_  | ~\new_[9241]_  | ~\new_[10419]_  | ~\new_[9239]_ ;
  assign \s9_addr_o[10]  = ~\new_[9246]_  | ~\new_[12039]_  | ~\new_[9245]_  | ~\new_[10428]_ ;
  assign \s9_addr_o[9]  = ~\new_[9248]_  | ~\new_[10432]_  | ~\new_[10430]_  | ~\new_[9247]_ ;
  assign \s9_addr_o[5]  = ~\new_[10445]_  | ~\new_[9256]_  | ~\new_[10443]_  | ~\new_[10444]_ ;
  assign \s9_addr_o[2]  = ~\new_[9259]_  | ~\new_[10455]_  | ~\new_[10453]_  | ~\new_[10454]_ ;
  assign \s9_addr_o[1]  = ~\new_[9263]_  | ~\new_[9261]_  | ~\new_[9260]_  | ~\new_[10456]_ ;
  assign \s9_addr_o[0]  = ~\new_[9265]_  | ~\new_[9266]_  | ~\new_[10458]_  | ~\new_[10459]_ ;
  assign \s9_sel_o[2]  = ~\new_[9268]_  | ~\new_[10465]_  | ~\new_[10462]_  | ~\new_[9269]_ ;
  assign \s9_sel_o[0]  = ~\new_[12081]_  | ~\new_[9276]_  | ~\new_[10468]_  | ~\new_[9275]_ ;
  assign s9_we_o = ~\new_[9278]_  | ~\new_[10471]_  | ~\new_[9277]_  | ~\new_[10470]_ ;
  assign \s11_addr_o[28]  = ~\new_[13163]_  | ~\new_[9327]_  | ~\new_[12394]_  | ~\new_[15216]_ ;
  assign \s11_addr_o[27]  = ~\new_[13938]_  | ~\new_[9328]_  | ~\new_[15217]_  | ~\new_[12399]_ ;
  assign \s11_addr_o[26]  = ~\new_[13944]_  | ~\new_[9330]_  | ~\new_[12401]_  | ~\new_[15223]_ ;
  assign \s12_data_o[28]  = ~\new_[15010]_  | ~\new_[9341]_  | ~\new_[10640]_  | ~\new_[12494]_ ;
  assign \s12_data_o[15]  = ~\new_[9351]_  | ~\new_[9352]_  | ~\new_[11185]_  | ~\new_[15329]_ ;
  assign \s12_data_o[14]  = ~\new_[15332]_  | ~\new_[9353]_  | ~\new_[10667]_  | ~\new_[12519]_ ;
  assign \s12_data_o[12]  = ~\new_[9572]_  | ~\new_[14037]_  | ~\new_[8658]_  | ~\new_[15335]_ ;
  assign \s12_data_o[10]  = ~\new_[9358]_  | ~\new_[14038]_  | ~\new_[9573]_  | ~\new_[15341]_ ;
  assign \s12_data_o[6]  = ~\new_[15350]_  | ~\new_[8933]_  | ~\new_[12535]_  | ~\new_[10087]_ ;
  assign \s12_addr_o[19]  = ~\new_[10696]_  | ~\new_[9371]_  | ~\new_[11833]_  | ~\new_[15404]_ ;
  assign \s12_addr_o[16]  = ~\new_[15412]_  | ~\new_[9244]_  | ~\new_[10702]_  | ~\new_[14085]_ ;
  assign \s12_addr_o[15]  = ~\new_[15415]_  | ~\new_[9375]_  | ~\new_[10703]_  | ~\new_[14088]_ ;
  assign \s12_addr_o[14]  = ~\new_[15417]_  | ~\new_[9376]_  | ~\new_[10704]_  | ~\new_[13347]_ ;
  assign \s12_addr_o[13]  = ~\new_[15421]_  | ~\new_[9377]_  | ~\new_[10705]_  | ~\new_[11561]_ ;
  assign \s12_addr_o[12]  = ~\new_[10706]_  | ~\new_[9379]_  | ~\new_[14885]_  | ~\new_[14093]_ ;
  assign \s12_addr_o[11]  = ~\new_[14095]_  | ~\new_[9380]_  | ~\new_[15433]_  | ~\new_[10708]_ ;
  assign \s12_addr_o[8]  = ~\new_[10711]_  | ~\new_[9382]_  | ~\new_[15436]_  | ~\new_[12490]_ ;
  assign \s12_addr_o[7]  = ~\new_[12580]_  | ~\new_[8867]_  | ~\new_[10713]_  | ~\new_[15439]_ ;
  assign \s12_addr_o[6]  = ~\new_[15442]_  | ~\new_[9383]_  | ~\new_[10714]_  | ~\new_[12582]_ ;
  assign \s12_addr_o[2]  = ~\new_[14689]_  | ~\new_[8828]_  | ~\new_[10722]_  | ~\new_[12591]_ ;
  assign \s12_addr_o[1]  = ~\new_[15456]_  | ~\new_[9388]_  | ~\new_[10724]_  | ~\new_[12609]_ ;
  assign \s12_addr_o[0]  = ~\new_[15626]_  | ~\new_[9384]_  | ~\new_[11097]_  | ~\new_[12962]_ ;
  assign \s12_sel_o[3]  = ~\new_[14978]_  | ~\new_[9385]_  | ~\new_[10482]_  | ~\new_[12593]_ ;
  assign \s12_sel_o[2]  = ~\new_[15460]_  | ~\new_[9386]_  | ~\new_[10208]_  | ~\new_[11515]_ ;
  assign \s12_sel_o[1]  = ~\new_[15862]_  | ~\new_[9387]_  | ~\new_[10725]_  | ~\new_[12599]_ ;
  assign \new_[6578]_  = ~\new_[32294]_  | ~\new_[7923]_ ;
  assign \s14_data_o[21]  = ~\new_[9411]_  | ~\new_[12850]_  | ~\new_[10927]_  | ~\new_[10928]_ ;
  assign \s14_addr_o[14]  = ~\new_[9476]_  | ~\new_[12931]_  | ~\new_[11032]_  | ~\new_[11033]_ ;
  assign \s14_addr_o[10]  = ~\new_[9482]_  | ~\new_[12937]_  | ~\new_[11040]_  | ~\new_[11041]_ ;
  assign \s14_sel_o[3]  = ~\new_[9495]_  | ~\new_[12964]_  | ~\new_[11067]_  | ~\new_[11068]_ ;
  assign s14_stb_o = \new_[8018]_  | \new_[8019]_ ;
  assign \new_[6584]_  = \new_[8775]_  | \new_[9558]_  | \new_[9798]_  | \new_[8637]_ ;
  assign \new_[6585]_  = \new_[8777]_  | \new_[9559]_  | \new_[9803]_  | \new_[8638]_ ;
  assign \new_[6586]_  = \new_[8784]_  | \new_[11141]_  | \new_[9815]_  | \new_[8639]_ ;
  assign \new_[6587]_  = \new_[8786]_  | \new_[9565]_  | \new_[9822]_  | \new_[8640]_ ;
  assign \new_[6588]_  = \new_[8787]_  | \new_[9566]_  | \new_[9826]_  | \new_[8643]_ ;
  assign \new_[6589]_  = \new_[8789]_  | \new_[9553]_  | \new_[9773]_  | \new_[8644]_ ;
  assign \new_[6590]_  = ~\new_[7924]_  & (~\new_[8666]_  | ~\new_[28424]_ );
  assign \new_[6591]_  = ~\new_[7925]_  & (~\new_[9287]_  | ~\new_[28151]_ );
  assign \new_[6592]_  = ~\new_[7926]_  & (~\new_[8669]_  | ~\new_[28744]_ );
  assign \new_[6593]_  = ~\new_[7927]_  & (~\new_[8139]_  | ~\new_[30263]_ );
  assign \new_[6594]_  = ~\new_[7928]_  & (~\new_[8175]_  | ~\new_[28143]_ );
  assign \new_[6595]_  = ~\new_[7929]_  & (~\new_[8178]_  | ~\new_[28109]_ );
  assign \new_[6596]_  = ~\new_[7930]_  & (~\new_[8683]_  | ~\new_[28690]_ );
  assign \new_[6597]_  = ~\new_[7931]_  & (~\new_[8221]_  | ~\new_[28736]_ );
  assign \new_[6598]_  = ~\new_[7932]_  & (~\new_[8686]_  | ~\new_[28330]_ );
  assign \new_[6599]_  = ~\new_[7936]_  & (~\new_[8142]_  | ~\new_[23176]_ );
  assign \new_[6600]_  = ~\s15_addr_o[5] ;
  assign \new_[6601]_  = ~\new_[8104]_  & ~\new_[9893]_ ;
  assign \new_[6602]_  = ~\new_[8613]_  & ~\new_[8083]_ ;
  assign \new_[6603]_  = ~\new_[8085]_  & ~\new_[8616]_ ;
  assign \new_[6604]_  = ~\new_[8082]_  & ~\new_[8475]_ ;
  assign \new_[6605]_  = ~\new_[8087]_  & ~\new_[8620]_ ;
  assign \new_[6606]_  = ~\new_[8089]_  & ~\new_[8623]_ ;
  assign \new_[6607]_  = ~\new_[8090]_  & ~\new_[8626]_ ;
  assign \new_[6608]_  = ~\new_[8094]_  & ~\new_[9545]_ ;
  assign \new_[6609]_  = ~\new_[8095]_  & ~\new_[8631]_ ;
  assign \new_[6610]_  = ~\new_[8632]_  & ~\new_[8096]_ ;
  assign \new_[6611]_  = ~\new_[8097]_  & ~\new_[8098]_ ;
  assign \new_[6612]_  = ~\new_[8099]_  & ~\new_[8100]_ ;
  assign \new_[6613]_  = ~\new_[8101]_  & ~\new_[8633]_ ;
  assign \new_[6614]_  = ~\new_[9548]_  & ~\new_[8103]_ ;
  assign \new_[6615]_  = ~\new_[8106]_  & (~\new_[13428]_  | ~\new_[30237]_ );
  assign \new_[6616]_  = ~\new_[8105]_  & (~\new_[16233]_  | ~\new_[28332]_ );
  assign \new_[6617]_  = ~\new_[7425]_  & (~\new_[16238]_  | ~\new_[30281]_ );
  assign \new_[6618]_  = ~\new_[7426]_  & (~\new_[16229]_  | ~\new_[28986]_ );
  assign \new_[6619]_  = ~\new_[7427]_  & (~\new_[17156]_  | ~\new_[26759]_ );
  assign \new_[6620]_  = ~\new_[7882]_  & ~\new_[8926]_ ;
  assign \new_[6621]_  = ~\new_[7883]_  & ~\new_[8929]_ ;
  assign \new_[6622]_  = ~\new_[7884]_  & ~\new_[8932]_ ;
  assign \new_[6623]_  = ~\new_[7885]_  & ~\new_[8934]_ ;
  assign \new_[6624]_  = ~\new_[7887]_  & ~\new_[8940]_ ;
  assign \new_[6625]_  = ~\new_[7888]_  & ~\new_[8943]_ ;
  assign \new_[6626]_  = ~\new_[7891]_  & ~\new_[8946]_ ;
  assign \new_[6627]_  = ~\new_[7894]_  & ~\new_[8948]_ ;
  assign \new_[6628]_  = ~\new_[7895]_  & ~\new_[8957]_ ;
  assign \new_[6629]_  = ~\new_[8358]_  & ~\new_[7903]_ ;
  assign \new_[6630]_  = ~\new_[9935]_  & ~\new_[7912]_ ;
  assign \new_[6631]_  = ~\new_[8295]_  & (~\new_[8450]_  | ~\new_[28424]_ );
  assign \new_[6632]_  = ~\new_[7900]_  & ~\new_[8853]_ ;
  assign \new_[6633]_  = ~\new_[9782]_  & (~\new_[8451]_  | ~\new_[27980]_ );
  assign \new_[6634]_  = ~\new_[8300]_  & (~\new_[8452]_  | ~\new_[28151]_ );
  assign \new_[6635]_  = ~\new_[8303]_  & (~\new_[8453]_  | ~\new_[28744]_ );
  assign \new_[6636]_  = ~\new_[8309]_  & (~\new_[8454]_  | ~\new_[30263]_ );
  assign \new_[6637]_  = ~\new_[8719]_  & ~\new_[7907]_ ;
  assign \new_[6638]_  = ~\new_[8321]_  & (~\new_[8455]_  | ~\new_[28143]_ );
  assign \new_[6639]_  = ~\new_[8325]_  & (~\new_[8456]_  | ~\new_[28109]_ );
  assign \new_[6640]_  = ~\new_[8326]_  & (~\new_[8457]_  | ~\new_[28690]_ );
  assign \new_[6641]_  = ~\new_[8330]_  & (~\new_[8458]_  | ~\new_[28736]_ );
  assign \new_[6642]_  = ~\new_[8340]_  & (~\new_[8459]_  | ~\new_[28330]_ );
  assign \new_[6643]_  = ~\new_[8343]_  & ~\new_[7910]_ ;
  assign \new_[6644]_  = (~\new_[32346]_  | ~\m0_data_i[31] ) & (~\new_[9929]_  | ~\m1_data_i[31] );
  assign \new_[6645]_  = (~\new_[13530]_  | ~\m2_data_i[31] ) & (~\new_[8408]_  | ~\m3_data_i[31] );
  assign \new_[6646]_  = (~\new_[11773]_  | ~\m6_data_i[31] ) & (~\new_[8391]_  | ~\m7_data_i[31] );
  assign \new_[6647]_  = (~\new_[32346]_  | ~\m0_data_i[30] ) & (~\new_[9929]_  | ~\m1_data_i[30] );
  assign \new_[6648]_  = (~\new_[8447]_  | ~\m6_data_i[30] ) & (~\new_[8851]_  | ~\m7_data_i[30] );
  assign \new_[6649]_  = (~\new_[13530]_  | ~\m2_data_i[30] ) & (~\new_[8407]_  | ~\m3_data_i[30] );
  assign \new_[6650]_  = (~\new_[8447]_  | ~\m6_data_i[29] ) & (~\new_[8851]_  | ~\m7_data_i[29] );
  assign \new_[6651]_  = (~\new_[8921]_  | ~\m2_data_i[29] ) & (~\new_[8407]_  | ~\m3_data_i[29] );
  assign \new_[6652]_  = (~\new_[32346]_  | ~\m0_data_i[28] ) & (~\new_[9929]_  | ~\m1_data_i[28] );
  assign \new_[6653]_  = (~\new_[8921]_  | ~\m2_data_i[28] ) & (~\new_[8407]_  | ~\m3_data_i[28] );
  assign \new_[6654]_  = (~\new_[11773]_  | ~\m6_data_i[28] ) & (~\new_[31989]_  | ~\m7_data_i[28] );
  assign \new_[6655]_  = (~\new_[32346]_  | ~\m0_data_i[27] ) & (~\new_[9929]_  | ~\m1_data_i[27] );
  assign \new_[6656]_  = (~\new_[13530]_  | ~\m2_data_i[27] ) & (~\new_[8407]_  | ~\m3_data_i[27] );
  assign \new_[6657]_  = (~\new_[11773]_  | ~\m6_data_i[27] ) & (~\new_[8391]_  | ~\m7_data_i[27] );
  assign \new_[6658]_  = (~\new_[32346]_  | ~\m0_data_i[26] ) & (~\new_[9929]_  | ~\m1_data_i[26] );
  assign \new_[6659]_  = (~\new_[8921]_  | ~\m2_data_i[26] ) & (~\new_[8408]_  | ~\m3_data_i[26] );
  assign \new_[6660]_  = (~\new_[8447]_  | ~\m6_data_i[26] ) & (~\new_[8391]_  | ~\m7_data_i[26] );
  assign \new_[6661]_  = (~\new_[32346]_  | ~\m0_data_i[25] ) & (~\new_[9929]_  | ~\m1_data_i[25] );
  assign \new_[6662]_  = (~\new_[8921]_  | ~\m2_data_i[25] ) & (~\new_[8408]_  | ~\m3_data_i[25] );
  assign \new_[6663]_  = (~\new_[8447]_  | ~\m6_data_i[25] ) & (~\new_[31989]_  | ~\m7_data_i[25] );
  assign \new_[6664]_  = (~\new_[32346]_  | ~\m0_data_i[24] ) & (~\new_[9929]_  | ~\m1_data_i[24] );
  assign \new_[6665]_  = (~\new_[8921]_  | ~\m2_data_i[24] ) & (~\new_[8407]_  | ~\m3_data_i[24] );
  assign \new_[6666]_  = (~\new_[8447]_  | ~\m6_data_i[24] ) & (~\new_[31989]_  | ~\m7_data_i[24] );
  assign \new_[6667]_  = (~\new_[32346]_  | ~\m0_data_i[23] ) & (~\new_[9929]_  | ~\m1_data_i[23] );
  assign \new_[6668]_  = (~\new_[8921]_  | ~\m2_data_i[23] ) & (~\new_[8408]_  | ~\m3_data_i[23] );
  assign \new_[6669]_  = (~\new_[11773]_  | ~\m6_data_i[23] ) & (~\new_[8391]_  | ~\m7_data_i[23] );
  assign \new_[6670]_  = (~\new_[32346]_  | ~\m0_data_i[22] ) & (~\new_[9929]_  | ~\m1_data_i[22] );
  assign \new_[6671]_  = (~\new_[8921]_  | ~\m2_data_i[22] ) & (~\new_[8407]_  | ~\m3_data_i[22] );
  assign \new_[6672]_  = (~\new_[8447]_  | ~\m6_data_i[22] ) & (~\new_[31989]_  | ~\m7_data_i[22] );
  assign \new_[6673]_  = (~\new_[32346]_  | ~\m0_data_i[21] ) & (~\new_[9929]_  | ~\m1_data_i[21] );
  assign \new_[6674]_  = (~\new_[13530]_  | ~\m2_data_i[21] ) & (~\new_[8407]_  | ~\m3_data_i[21] );
  assign \new_[6675]_  = (~\new_[8447]_  | ~\m6_data_i[21] ) & (~\new_[8851]_  | ~\m7_data_i[21] );
  assign \new_[6676]_  = (~\new_[32346]_  | ~\m0_data_i[20] ) & (~\new_[9929]_  | ~\m1_data_i[20] );
  assign \new_[6677]_  = (~\new_[13530]_  | ~\m2_data_i[20] ) & (~\new_[8408]_  | ~\m3_data_i[20] );
  assign \new_[6678]_  = (~\new_[8447]_  | ~\m6_data_i[20] ) & (~\new_[8851]_  | ~\m7_data_i[20] );
  assign \new_[6679]_  = (~\new_[32346]_  | ~\m0_data_i[19] ) & (~\new_[9929]_  | ~\m1_data_i[19] );
  assign \new_[6680]_  = (~\new_[13530]_  | ~\m2_data_i[19] ) & (~\new_[8408]_  | ~\m3_data_i[19] );
  assign \new_[6681]_  = (~\new_[8447]_  | ~\m6_data_i[19] ) & (~\new_[8851]_  | ~\m7_data_i[19] );
  assign \new_[6682]_  = (~\new_[8921]_  | ~\m2_data_i[18] ) & (~\new_[8408]_  | ~\m3_data_i[18] );
  assign \new_[6683]_  = (~\new_[32346]_  | ~\m0_data_i[18] ) & (~\new_[9929]_  | ~\m1_data_i[18] );
  assign \new_[6684]_  = (~\new_[11773]_  | ~\m6_data_i[18] ) & (~\new_[8391]_  | ~\m7_data_i[18] );
  assign \new_[6685]_  = (~\new_[13530]_  | ~\m2_data_i[17] ) & (~\new_[8407]_  | ~\m3_data_i[17] );
  assign \new_[6686]_  = (~\new_[32346]_  | ~\m0_data_i[17] ) & (~\new_[13487]_  | ~\m1_data_i[17] );
  assign \new_[6687]_  = (~\new_[11773]_  | ~\m6_data_i[17] ) & (~\new_[8391]_  | ~\m7_data_i[17] );
  assign \new_[6688]_  = (~\new_[32346]_  | ~\m0_data_i[16] ) & (~\new_[9929]_  | ~\m1_data_i[16] );
  assign \new_[6689]_  = (~\new_[8921]_  | ~\m2_data_i[16] ) & (~\new_[8407]_  | ~\m3_data_i[16] );
  assign \new_[6690]_  = (~\new_[8447]_  | ~\m6_data_i[16] ) & (~\new_[8391]_  | ~\m7_data_i[16] );
  assign \new_[6691]_  = ~\new_[7889]_  & ~\new_[8903]_ ;
  assign \new_[6692]_  = ~\new_[7893]_  & ~\new_[8906]_ ;
  assign \new_[6693]_  = ~\new_[8444]_  & ~\new_[7897]_ ;
  assign \new_[6694]_  = ~\new_[7898]_  & ~\new_[7901]_ ;
  assign \new_[6695]_  = ~\new_[7913]_  & ~\new_[8949]_ ;
  assign \new_[6696]_  = ~\new_[8782]_  & ~\new_[7905]_ ;
  assign \new_[6697]_  = ~\new_[8468]_  & ~\new_[7909]_ ;
  assign \new_[6698]_  = ~\new_[8356]_  & ~\new_[7906]_ ;
  assign \new_[6699]_  = (~\new_[8447]_  | ~\m6_addr_i[31] ) & (~\new_[14850]_  | ~\new_[31001]_ );
  assign \new_[6700]_  = (~\new_[11613]_  | ~\m3_addr_i[31] ) & (~\new_[13526]_  | ~\m4_addr_i[31] );
  assign \new_[6701]_  = (~\new_[8447]_  | ~\m6_addr_i[30] ) & (~\new_[14850]_  | ~\new_[31147]_ );
  assign \new_[6702]_  = (~\new_[11613]_  | ~\m3_addr_i[30] ) & (~\new_[13526]_  | ~\m4_addr_i[30] );
  assign \new_[6703]_  = (~\new_[8447]_  | ~\m6_addr_i[29] ) & (~\new_[14850]_  | ~\new_[31407]_ );
  assign \new_[6704]_  = (~\new_[11613]_  | ~\m3_addr_i[29] ) & (~\new_[13526]_  | ~\m4_addr_i[29] );
  assign \new_[6705]_  = (~\new_[8851]_  | ~\new_[31531]_ ) & (~\new_[32346]_  | ~\new_[31481]_ );
  assign \new_[6706]_  = (~\new_[8447]_  | ~\m6_addr_i[28] ) & (~\new_[14850]_  | ~\new_[31276]_ );
  assign \new_[6707]_  = (~\new_[11613]_  | ~\m3_addr_i[28] ) & (~\new_[13526]_  | ~\m4_addr_i[28] );
  assign \new_[6708]_  = (~\new_[32346]_  | ~\m0_addr_i[23] ) & (~\new_[9929]_  | ~\m1_addr_i[23] );
  assign \new_[6709]_  = (~\new_[8921]_  | ~\m2_addr_i[23] ) & (~\new_[8408]_  | ~\m3_addr_i[23] );
  assign \new_[6710]_  = (~\new_[8447]_  | ~\m6_addr_i[23] ) & (~\new_[31989]_  | ~\m7_addr_i[23] );
  assign \new_[6711]_  = (~\new_[32346]_  | ~\m0_addr_i[22] ) & (~\new_[9929]_  | ~\m1_addr_i[22] );
  assign \new_[6712]_  = (~\new_[8921]_  | ~\m2_addr_i[22] ) & (~\new_[8408]_  | ~\m3_addr_i[22] );
  assign \new_[6713]_  = (~\new_[8447]_  | ~\m6_addr_i[22] ) & (~\new_[31989]_  | ~\m7_addr_i[22] );
  assign \new_[6714]_  = (~\new_[8447]_  | ~\m6_addr_i[21] ) & (~\new_[8851]_  | ~\m7_addr_i[21] );
  assign \new_[6715]_  = (~\new_[32346]_  | ~\m0_addr_i[21] ) & (~\new_[13487]_  | ~\m1_addr_i[21] );
  assign \new_[6716]_  = (~\new_[13530]_  | ~\m2_addr_i[21] ) & (~\new_[8407]_  | ~\m3_addr_i[21] );
  assign \new_[6717]_  = (~\new_[32346]_  | ~\m0_addr_i[20] ) & (~\new_[9929]_  | ~\m1_addr_i[20] );
  assign \new_[6718]_  = (~\new_[8921]_  | ~\m2_addr_i[20] ) & (~\new_[8407]_  | ~\m3_addr_i[20] );
  assign \new_[6719]_  = (~\new_[8447]_  | ~\m6_addr_i[20] ) & (~\new_[31989]_  | ~\m7_addr_i[20] );
  assign \new_[6720]_  = (~\new_[32346]_  | ~\m0_addr_i[19] ) & (~\new_[9929]_  | ~\m1_addr_i[19] );
  assign \new_[6721]_  = (~\new_[8921]_  | ~\m2_addr_i[19] ) & (~\new_[8407]_  | ~\m3_addr_i[19] );
  assign \new_[6722]_  = (~\new_[8447]_  | ~\m6_addr_i[19] ) & (~\new_[8391]_  | ~\m7_addr_i[19] );
  assign \new_[6723]_  = (~\new_[32346]_  | ~\m0_addr_i[18] ) & (~\new_[9929]_  | ~\m1_addr_i[18] );
  assign \new_[6724]_  = ~\new_[7911]_  | ~\new_[10028]_ ;
  assign \new_[6725]_  = (~\new_[8921]_  | ~\m2_addr_i[18] ) & (~\new_[8407]_  | ~\m3_addr_i[18] );
  assign \new_[6726]_  = (~\new_[8447]_  | ~\m6_addr_i[18] ) & (~\new_[8391]_  | ~\m7_addr_i[18] );
  assign \new_[6727]_  = (~\new_[32346]_  | ~\m0_addr_i[17] ) & (~\new_[9929]_  | ~\m1_addr_i[17] );
  assign \new_[6728]_  = (~\new_[8921]_  | ~\m2_addr_i[17] ) & (~\new_[8407]_  | ~\m3_addr_i[17] );
  assign \new_[6729]_  = (~\new_[8447]_  | ~\m6_addr_i[17] ) & (~\new_[8851]_  | ~\m7_addr_i[17] );
  assign \new_[6730]_  = (~\new_[32346]_  | ~\m0_addr_i[16] ) & (~\new_[9929]_  | ~\m1_addr_i[16] );
  assign \new_[6731]_  = (~\new_[8921]_  | ~\m2_addr_i[16] ) & (~\new_[8407]_  | ~\m3_addr_i[16] );
  assign \new_[6732]_  = (~\new_[8447]_  | ~\m6_addr_i[16] ) & (~\new_[31989]_  | ~\m7_addr_i[16] );
  assign \new_[6733]_  = (~\new_[8447]_  | ~\m6_addr_i[15] ) & (~\new_[8851]_  | ~\m7_addr_i[15] );
  assign \new_[6734]_  = (~\new_[32346]_  | ~\m0_addr_i[15] ) & (~\new_[13487]_  | ~\m1_addr_i[15] );
  assign \new_[6735]_  = (~\new_[13530]_  | ~\m2_addr_i[15] ) & (~\new_[8407]_  | ~\m3_addr_i[15] );
  assign \new_[6736]_  = (~\new_[32346]_  | ~\m0_addr_i[14] ) & (~\new_[9929]_  | ~\m1_addr_i[14] );
  assign \new_[6737]_  = (~\new_[8921]_  | ~\m2_addr_i[14] ) & (~\new_[8407]_  | ~\m3_addr_i[14] );
  assign \new_[6738]_  = (~\new_[11773]_  | ~\m6_addr_i[14] ) & (~\new_[8391]_  | ~\m7_addr_i[14] );
  assign \new_[6739]_  = (~\new_[32346]_  | ~\m0_addr_i[13] ) & (~\new_[9929]_  | ~\m1_addr_i[13] );
  assign \new_[6740]_  = (~\new_[8921]_  | ~\m2_addr_i[13] ) & (~\new_[8408]_  | ~\m3_addr_i[13] );
  assign \new_[6741]_  = (~\new_[8447]_  | ~\m6_addr_i[13] ) & (~\new_[8391]_  | ~\m7_addr_i[13] );
  assign \new_[6742]_  = (~\new_[32346]_  | ~\m0_addr_i[12] ) & (~\new_[9929]_  | ~\m1_addr_i[12] );
  assign \new_[6743]_  = (~\new_[8921]_  | ~\m2_addr_i[12] ) & (~\new_[8408]_  | ~\m3_addr_i[12] );
  assign \new_[6744]_  = (~\new_[8447]_  | ~\m6_addr_i[12] ) & (~\new_[8391]_  | ~\m7_addr_i[12] );
  assign \new_[6745]_  = (~\new_[32346]_  | ~\m0_addr_i[11] ) & (~\new_[9929]_  | ~\m1_addr_i[11] );
  assign \new_[6746]_  = (~\new_[8921]_  | ~\m2_addr_i[11] ) & (~\new_[8407]_  | ~\m3_addr_i[11] );
  assign \new_[6747]_  = (~\new_[11773]_  | ~\m6_addr_i[11] ) & (~\new_[8851]_  | ~\m7_addr_i[11] );
  assign \new_[6748]_  = (~\new_[32346]_  | ~\m0_addr_i[10] ) & (~\new_[9929]_  | ~\m1_addr_i[10] );
  assign \new_[6749]_  = (~\new_[8921]_  | ~\m2_addr_i[10] ) & (~\new_[8408]_  | ~\m3_addr_i[10] );
  assign \new_[6750]_  = (~\new_[11773]_  | ~\m6_addr_i[10] ) & (~\new_[8851]_  | ~\m7_addr_i[10] );
  assign \new_[6751]_  = (~\new_[8447]_  | ~\m6_addr_i[9] ) & (~\new_[8851]_  | ~\m7_addr_i[9] );
  assign \new_[6752]_  = (~\new_[32346]_  | ~\m0_addr_i[9] ) & (~\new_[13487]_  | ~\m1_addr_i[9] );
  assign \new_[6753]_  = (~\new_[8921]_  | ~\m2_addr_i[9] ) & (~\new_[11613]_  | ~\m3_addr_i[9] );
  assign \new_[6754]_  = (~\new_[32346]_  | ~\m0_addr_i[8] ) & (~\new_[9929]_  | ~\m1_addr_i[8] );
  assign \new_[6755]_  = (~\new_[8921]_  | ~\m2_addr_i[8] ) & (~\new_[8407]_  | ~\m3_addr_i[8] );
  assign \new_[6756]_  = (~\new_[8447]_  | ~\m6_addr_i[8] ) & (~\new_[8391]_  | ~\m7_addr_i[8] );
  assign \new_[6757]_  = (~\new_[32346]_  | ~\m0_addr_i[7] ) & (~\new_[9929]_  | ~\m1_addr_i[7] );
  assign \new_[6758]_  = (~\new_[13530]_  | ~\m2_addr_i[7] ) & (~\new_[8407]_  | ~\m3_addr_i[7] );
  assign \new_[6759]_  = (~\new_[11773]_  | ~\m6_addr_i[7] ) & (~\new_[8391]_  | ~\m7_addr_i[7] );
  assign \new_[6760]_  = (~\new_[32346]_  | ~\m0_addr_i[6] ) & (~\new_[9929]_  | ~\m1_addr_i[6] );
  assign \new_[6761]_  = (~\new_[8921]_  | ~\m2_addr_i[6] ) & (~\new_[8407]_  | ~\m3_addr_i[6] );
  assign \new_[6762]_  = (~\new_[11773]_  | ~\m6_addr_i[6] ) & (~\new_[8391]_  | ~\m7_addr_i[6] );
  assign \new_[6763]_  = (~\new_[32346]_  | ~\m0_addr_i[1] ) & (~\new_[9929]_  | ~\m1_addr_i[1] );
  assign \new_[6764]_  = (~\new_[13530]_  | ~\m2_addr_i[1] ) & (~\new_[8408]_  | ~\m3_addr_i[1] );
  assign \new_[6765]_  = (~\new_[11773]_  | ~\m6_addr_i[1] ) & (~\new_[8851]_  | ~\m7_addr_i[1] );
  assign \new_[6766]_  = (~\new_[32346]_  | ~\m0_addr_i[0] ) & (~\new_[9929]_  | ~\m1_addr_i[0] );
  assign \new_[6767]_  = (~\new_[8921]_  | ~\m2_addr_i[0] ) & (~\new_[8407]_  | ~\m3_addr_i[0] );
  assign \new_[6768]_  = (~\new_[11773]_  | ~\m6_addr_i[0] ) & (~\new_[8851]_  | ~\m7_addr_i[0] );
  assign \new_[6769]_  = (~\new_[8447]_  | ~\m6_sel_i[3] ) & (~\new_[8851]_  | ~\m7_sel_i[3] );
  assign \new_[6770]_  = (~\new_[32346]_  | ~\m0_sel_i[3] ) & (~\new_[13487]_  | ~\m1_sel_i[3] );
  assign \new_[6771]_  = (~\new_[13530]_  | ~\m2_sel_i[3] ) & (~\new_[8407]_  | ~\m3_sel_i[3] );
  assign \new_[6772]_  = (~\new_[32346]_  | ~\m0_sel_i[2] ) & (~\new_[9929]_  | ~\m1_sel_i[2] );
  assign \new_[6773]_  = (~\new_[8921]_  | ~\m2_sel_i[2] ) & (~\new_[8408]_  | ~\m3_sel_i[2] );
  assign \new_[6774]_  = (~\new_[8447]_  | ~\m6_sel_i[2] ) & (~\new_[8851]_  | ~\m7_sel_i[2] );
  assign \new_[6775]_  = (~\new_[8921]_  | ~\m2_sel_i[1] ) & (~\new_[8408]_  | ~\m3_sel_i[1] );
  assign \new_[6776]_  = (~\new_[11773]_  | ~\m6_sel_i[1] ) & (~\new_[8391]_  | ~\m7_sel_i[1] );
  assign \new_[6777]_  = (~\new_[8921]_  | ~\m2_sel_i[0] ) & (~\new_[8408]_  | ~\m3_sel_i[0] );
  assign \new_[6778]_  = (~\new_[11773]_  | ~\m6_sel_i[0] ) & (~\new_[8851]_  | ~\m7_sel_i[0] );
  assign \new_[6779]_  = \\s15_msel_pri_out_reg[0] ;
  assign \new_[6780]_  = \\s2_msel_pri_out_reg[0] ;
  assign \new_[6781]_  = \\s1_msel_pri_out_reg[0] ;
  assign \new_[6782]_  = \\s7_msel_pri_out_reg[0] ;
  assign \new_[6783]_  = \\s9_msel_pri_out_reg[0] ;
  assign \new_[6784]_  = \\s0_msel_pri_out_reg[0] ;
  assign \new_[6785]_  = ~s11_next_reg;
  assign \new_[6786]_  = ~s2_next_reg;
  assign \new_[6787]_  = ~s4_next_reg;
  assign \new_[6788]_  = ~s7_next_reg;
  assign \new_[6789]_  = \\s11_msel_pri_out_reg[1] ;
  assign \new_[6790]_  = \\s12_msel_pri_out_reg[1] ;
  assign \new_[6791]_  = \\s13_msel_pri_out_reg[1] ;
  assign \new_[6792]_  = \\s3_msel_pri_out_reg[1] ;
  assign \new_[6793]_  = \\s5_msel_pri_out_reg[1] ;
  assign \new_[6794]_  = \\s6_msel_pri_out_reg[1] ;
  assign n7429 = (~\new_[9310]_  & ~rst_i) | (~\new_[31183]_  & ~\new_[31810]_ );
  assign s6_cyc_o = ~n7484;
  assign \s0_data_o[29]  = ~\new_[10388]_  | ~\new_[12003]_  | ~\new_[9218]_  | ~\new_[11998]_ ;
  assign \s0_data_o[26]  = ~\new_[10422]_  | ~\new_[12037]_  | ~\new_[12030]_  | ~\new_[10420]_ ;
  assign \s0_data_o[14]  = ~\new_[13725]_  | ~\new_[10486]_  | ~\new_[10484]_  | ~\new_[10485]_ ;
  assign \s0_data_o[13]  = ~\new_[10490]_  | ~\new_[13731]_  | ~\new_[10488]_  | ~\new_[10489]_ ;
  assign \s0_data_o[12]  = ~\new_[10493]_  | ~\new_[12150]_  | ~\new_[12142]_  | ~\new_[12146]_ ;
  assign \s0_data_o[11]  = ~\new_[13745]_  | ~\new_[10499]_  | ~\new_[10495]_  | ~\new_[10496]_ ;
  assign \s0_data_o[10]  = ~\new_[10505]_  | ~\new_[10506]_  | ~\new_[10502]_  | ~\new_[13750]_ ;
  assign \s0_data_o[9]  = ~\new_[10508]_  | ~\new_[12179]_  | ~\new_[12130]_  | ~\new_[9180]_ ;
  assign \s0_data_o[8]  = ~\new_[10513]_  | ~\new_[12189]_  | ~\new_[12180]_  | ~\new_[9301]_ ;
  assign \s0_data_o[7]  = ~\new_[10519]_  | ~\new_[12203]_  | ~\new_[12192]_  | ~\new_[10516]_ ;
  assign \s0_data_o[6]  = ~\new_[12215]_  | ~\new_[10524]_  | ~\new_[10595]_  | ~\new_[10523]_ ;
  assign \s0_data_o[5]  = ~\new_[10527]_  | ~\new_[12224]_  | ~\new_[9307]_  | ~\new_[12219]_ ;
  assign \s0_data_o[4]  = ~\new_[13783]_  | ~\new_[12235]_  | ~\new_[12227]_  | ~\new_[9308]_ ;
  assign \s0_data_o[3]  = ~\new_[10532]_  | ~\new_[12245]_  | ~\new_[12386]_  | ~\new_[12243]_ ;
  assign \s0_data_o[2]  = ~\new_[9916]_  | ~\new_[13800]_  | ~\new_[10533]_  | ~\new_[10534]_ ;
  assign \s0_data_o[1]  = ~\new_[12259]_  | ~\new_[10537]_  | ~\new_[12255]_  | ~\new_[9309]_ ;
  assign \s0_data_o[0]  = ~\new_[10538]_  | ~\new_[12266]_  | ~\new_[12260]_  | ~\new_[12265]_ ;
  assign \s0_addr_o[25]  = ~\new_[10545]_  | ~\new_[12303]_  | ~\new_[13843]_  | ~\new_[12298]_ ;
  assign \s0_addr_o[24]  = ~\new_[10548]_  | ~\new_[12312]_  | ~\new_[13848]_  | ~\new_[12308]_ ;
  assign \s0_addr_o[22]  = ~\new_[12331]_  | ~\new_[13859]_  | ~\new_[12326]_  | ~\new_[8832]_ ;
  assign \s0_addr_o[13]  = ~\new_[12398]_  | ~\new_[12400]_  | ~\new_[12390]_  | ~\new_[9326]_ ;
  assign \s0_addr_o[9]  = ~\new_[10600]_  | ~\new_[11173]_  | ~\new_[12432]_  | ~\new_[13016]_ ;
  assign \s0_addr_o[8]  = ~\new_[10602]_  | ~\new_[10603]_  | ~\new_[9604]_  | ~\new_[12439]_ ;
  assign \s0_addr_o[3]  = ~\new_[12487]_  | ~\new_[10629]_  | ~\new_[10625]_  | ~\new_[12485]_ ;
  assign \s0_addr_o[1]  = ~\new_[10634]_  | ~\new_[10231]_  | ~\new_[12500]_  | ~\new_[12689]_ ;
  assign \s0_addr_o[2]  = ~\new_[13999]_  | ~\new_[10633]_  | ~\new_[10632]_  | ~\new_[12495]_ ;
  assign \s0_sel_o[1]  = ~\new_[10655]_  | ~\new_[10657]_  | ~\new_[10653]_  | ~\new_[12513]_ ;
  assign s1_stb_o = \new_[8472]_  | \new_[8473]_ ;
  assign \s2_data_o[31]  = ~\new_[10972]_  | ~\new_[14338]_  | ~\new_[12895]_  | ~\new_[15668]_ ;
  assign \s2_data_o[30]  = ~\new_[10982]_  | ~\new_[12900]_  | ~\new_[15669]_  | ~\new_[14339]_ ;
  assign \s2_data_o[28]  = ~\new_[10998]_  | ~\new_[14342]_  | ~\new_[15670]_  | ~\new_[15671]_ ;
  assign \s2_data_o[26]  = ~\new_[15678]_  | ~\new_[11014]_  | ~\new_[15674]_  | ~\new_[15676]_ ;
  assign s8_cyc_o = ~n7494;
  assign s2_stb_o = \new_[10994]_  | \new_[8547]_ ;
  assign \s3_data_o[30]  = ~\new_[11145]_  | ~\new_[14488]_  | ~\new_[13093]_  | ~\new_[11144]_ ;
  assign \s3_data_o[29]  = ~\new_[11148]_  | ~\new_[15886]_  | ~\new_[13094]_  | ~\new_[11147]_ ;
  assign \s3_data_o[17]  = ~\new_[9581]_  | ~\new_[13115]_  | ~\new_[11164]_  | ~\new_[9580]_ ;
  assign \s3_data_o[15]  = ~\new_[9584]_  | ~\new_[13119]_  | ~\new_[11166]_  | ~\new_[9583]_ ;
  assign \s3_data_o[14]  = ~\new_[9587]_  | ~\new_[13121]_  | ~\new_[13120]_  | ~\new_[9585]_ ;
  assign \s3_data_o[13]  = ~\new_[9589]_  | ~\new_[13123]_  | ~\new_[13122]_  | ~\new_[9588]_ ;
  assign \s3_data_o[12]  = ~\new_[9591]_  | ~\new_[13125]_  | ~\new_[13124]_  | ~\new_[9590]_ ;
  assign \s3_data_o[10]  = ~\new_[9594]_  | ~\new_[13130]_  | ~\new_[13128]_  | ~\new_[9593]_ ;
  assign \s3_data_o[9]  = ~\new_[9596]_  | ~\new_[13132]_  | ~\new_[13131]_  | ~\new_[9595]_ ;
  assign \s3_data_o[8]  = ~\new_[9598]_  | ~\new_[13134]_  | ~\new_[11169]_  | ~\new_[9597]_ ;
  assign \s3_data_o[7]  = ~\new_[9600]_  | ~\new_[13135]_  | ~\new_[11170]_  | ~\new_[9599]_ ;
  assign \s3_data_o[6]  = ~\new_[9603]_  | ~\new_[13137]_  | ~\new_[11171]_  | ~\new_[9601]_ ;
  assign \s3_data_o[5]  = ~\new_[9606]_  | ~\new_[13138]_  | ~\new_[11172]_  | ~\new_[9605]_ ;
  assign \s3_data_o[4]  = ~\new_[9608]_  | ~\new_[13140]_  | ~\new_[13139]_  | ~\new_[9607]_ ;
  assign \s3_data_o[3]  = ~\new_[9611]_  | ~\new_[13141]_  | ~\new_[11175]_  | ~\new_[9610]_ ;
  assign \s3_data_o[2]  = ~\new_[9613]_  | ~\new_[13144]_  | ~\new_[13143]_  | ~\new_[9612]_ ;
  assign \s3_data_o[1]  = ~\new_[9615]_  | ~\new_[13146]_  | ~\new_[13145]_  | ~\new_[9614]_ ;
  assign \s3_data_o[0]  = ~\new_[9617]_  | ~\new_[13147]_  | ~\new_[11176]_  | ~\new_[9616]_ ;
  assign \s3_addr_o[28]  = ~\new_[9620]_  | ~\new_[13158]_  | ~\new_[13156]_  | ~\new_[11184]_ ;
  assign \s3_addr_o[27]  = ~\new_[9621]_  | ~\new_[13162]_  | ~\new_[13160]_  | ~\new_[11186]_ ;
  assign \s3_addr_o[26]  = ~\new_[10201]_  | ~\new_[13441]_  | ~\new_[13164]_  | ~\new_[11187]_ ;
  assign \s3_addr_o[25]  = ~\new_[11112]_  | ~\new_[13166]_  | ~\new_[13159]_  | ~\new_[13081]_ ;
  assign \s3_addr_o[24]  = ~\new_[9624]_  | ~\new_[13939]_  | ~\new_[13167]_  | ~\new_[11188]_ ;
  assign \s3_addr_o[15]  = ~\new_[9641]_  | ~\new_[14483]_  | ~\new_[11210]_  | ~\new_[9640]_ ;
  assign \s3_addr_o[14]  = ~\new_[9643]_  | ~\new_[13186]_  | ~\new_[11215]_  | ~\new_[9642]_ ;
  assign \s3_addr_o[8]  = ~\new_[9654]_  | ~\new_[13202]_  | ~\new_[11228]_  | ~\new_[9653]_ ;
  assign \s3_addr_o[5]  = ~\new_[9656]_  | ~\new_[13650]_  | ~\new_[12560]_  | ~\new_[10006]_ ;
  assign \s3_addr_o[4]  = ~\new_[9658]_  | ~\new_[13595]_  | ~\new_[13615]_  | ~\new_[10195]_ ;
  assign \s3_addr_o[3]  = ~\new_[10076]_  | ~\new_[13545]_  | ~\new_[11870]_  | ~\new_[10091]_ ;
  assign \s3_addr_o[2]  = ~\new_[9989]_  | ~\new_[13506]_  | ~\new_[11751]_  | ~\new_[10009]_ ;
  assign \s3_addr_o[0]  = ~\new_[11018]_  | ~\new_[14157]_  | ~\new_[13043]_  | ~\new_[14405]_ ;
  assign s3_we_o = ~\new_[9632]_  | ~\new_[14022]_  | ~\new_[11695]_  | ~\new_[9943]_ ;
  assign \s3_sel_o[1]  = ~\new_[10081]_  | ~\new_[13546]_  | ~\new_[11853]_  | ~\new_[10095]_ ;
  assign \s4_data_o[31]  = ~\new_[15425]_  | ~\new_[10669]_  | ~\new_[12880]_  | ~\new_[12544]_ ;
  assign \s4_data_o[30]  = ~\new_[16333]_  | ~\new_[10181]_  | ~\new_[12351]_  | ~\new_[11958]_ ;
  assign \s4_data_o[28]  = ~\new_[16319]_  | ~\new_[9992]_  | ~\new_[11778]_  | ~\new_[11755]_ ;
  assign \s4_data_o[24]  = ~\new_[14974]_  | ~\new_[10024]_  | ~\new_[12404]_  | ~\new_[12233]_ ;
  assign \s4_data_o[23]  = ~\new_[15020]_  | ~\new_[9666]_  | ~\new_[11741]_  | ~\new_[11233]_ ;
  assign \s4_data_o[22]  = ~\new_[15129]_  | ~\new_[9626]_  | ~\new_[11190]_  | ~\new_[11197]_ ;
  assign \s4_data_o[19]  = ~\new_[14537]_  | ~\new_[9638]_  | ~\new_[11217]_  | ~\new_[11211]_ ;
  assign n7434 = (~\new_[9312]_  & ~rst_i) | (~\new_[30812]_  & ~\new_[31718]_ );
  assign \s4_data_o[18]  = ~\new_[14871]_  | ~\new_[10005]_  | ~\new_[11194]_  | ~\new_[11865]_ ;
  assign \s4_data_o[13]  = ~\new_[15561]_  | ~\new_[10382]_  | ~\new_[12493]_  | ~\new_[11246]_ ;
  assign \s4_data_o[12]  = ~\new_[14904]_  | ~\new_[11121]_  | ~\new_[11953]_  | ~\new_[11247]_ ;
  assign \s4_data_o[11]  = ~\new_[15303]_  | ~\new_[10220]_  | ~\new_[12902]_  | ~\new_[12756]_ ;
  assign \s4_data_o[10]  = ~\new_[15818]_  | ~\new_[9586]_  | ~\new_[11997]_  | ~\new_[11340]_ ;
  assign \s4_data_o[8]  = ~\new_[14947]_  | ~\new_[9672]_  | ~\new_[11860]_  | ~\new_[11249]_ ;
  assign \s4_data_o[7]  = ~\new_[14903]_  | ~\new_[9908]_  | ~\new_[12412]_  | ~\new_[12112]_ ;
  assign \s4_data_o[4]  = ~\new_[15779]_  | ~\new_[10813]_  | ~\new_[11309]_  | ~\new_[11640]_ ;
  assign \s4_data_o[1]  = ~\new_[14527]_  | ~\new_[9676]_  | ~\new_[11947]_  | ~\new_[11659]_ ;
  assign \s4_addr_o[22]  = ~\new_[14529]_  | ~\new_[10413]_  | ~\new_[11199]_  | ~\new_[11195]_ ;
  assign \s4_addr_o[20]  = ~\new_[14912]_  | ~\new_[9668]_  | ~\new_[11872]_  | ~\new_[11244]_ ;
  assign \s4_addr_o[19]  = ~\new_[14787]_  | ~\new_[10865]_  | ~\new_[11446]_  | ~\new_[11225]_ ;
  assign \s4_addr_o[17]  = ~\new_[15017]_  | ~\new_[9670]_  | ~\new_[13025]_  | ~\new_[11248]_ ;
  assign \s4_addr_o[14]  = ~\new_[14674]_  | ~\new_[10959]_  | ~\new_[12942]_  | ~\new_[11559]_ ;
  assign \s4_addr_o[12]  = ~\new_[15923]_  | ~\new_[10608]_  | ~\new_[11251]_  | ~\new_[11587]_ ;
  assign \s4_addr_o[11]  = ~\new_[14541]_  | ~\new_[9675]_  | ~\new_[11300]_  | ~\new_[11213]_ ;
  assign \s4_addr_o[9]  = ~\new_[14559]_  | ~\new_[9677]_  | ~\new_[11261]_  | ~\new_[11263]_ ;
  assign \s4_addr_o[8]  = ~\new_[14562]_  | ~\new_[9679]_  | ~\new_[11266]_  | ~\new_[11268]_ ;
  assign \s4_addr_o[6]  = ~\new_[14568]_  | ~\new_[9680]_  | ~\new_[11272]_  | ~\new_[11273]_ ;
  assign \s4_addr_o[4]  = ~\new_[14574]_  | ~\new_[9683]_  | ~\new_[11278]_  | ~\new_[11279]_ ;
  assign \s4_addr_o[3]  = ~\new_[14577]_  | ~\new_[9687]_  | ~\new_[11280]_  | ~\new_[14576]_ ;
  assign \s4_addr_o[2]  = ~\new_[14578]_  | ~\new_[9689]_  | ~\new_[11281]_  | ~\new_[11282]_ ;
  assign \s4_addr_o[1]  = ~\new_[14580]_  | ~\new_[9691]_  | ~\new_[11283]_  | ~\new_[11284]_ ;
  assign \s4_addr_o[0]  = ~\new_[14582]_  | ~\new_[9693]_  | ~\new_[11285]_  | ~\new_[11286]_ ;
  assign \s4_sel_o[2]  = ~\new_[15986]_  | ~\new_[9695]_  | ~\new_[11291]_  | ~\new_[11292]_ ;
  assign s4_stb_o = \new_[8516]_  | \new_[8517]_ ;
  assign s9_cyc_o = ~n7489;
  assign \s6_data_o[30]  = ~\new_[9781]_  | ~\new_[13395]_  | ~\new_[11424]_  | ~\new_[9778]_ ;
  assign \s6_data_o[25]  = ~\new_[9791]_  | ~\new_[11438]_  | ~\new_[11437]_  | ~\new_[9790]_ ;
  assign \s6_data_o[24]  = ~\new_[9793]_  | ~\new_[11440]_  | ~\new_[11439]_  | ~\new_[9792]_ ;
  assign \s6_data_o[22]  = ~\new_[9797]_  | ~\new_[11447]_  | ~\new_[11445]_  | ~\new_[9796]_ ;
  assign \s6_data_o[21]  = ~\new_[9800]_  | ~\new_[13415]_  | ~\new_[11448]_  | ~\new_[9799]_ ;
  assign \s6_data_o[20]  = ~\new_[9804]_  | ~\new_[13416]_  | ~\new_[11449]_  | ~\new_[9802]_ ;
  assign \s6_data_o[19]  = ~\new_[9806]_  | ~\new_[11455]_  | ~\new_[11451]_  | ~\new_[9805]_ ;
  assign \s6_addr_o[18]  = ~\new_[9868]_  | ~\new_[11553]_  | ~\new_[11551]_  | ~\new_[9867]_ ;
  assign \s6_addr_o[17]  = ~\new_[9870]_  | ~\new_[11557]_  | ~\new_[11555]_  | ~\new_[9869]_ ;
  assign \s6_addr_o[13]  = ~\new_[9879]_  | ~\new_[11569]_  | ~\new_[11568]_  | ~\new_[9877]_ ;
  assign \s6_addr_o[11]  = ~\new_[9883]_  | ~\new_[11575]_  | ~\new_[11574]_  | ~\new_[9881]_ ;
  assign \s6_addr_o[8]  = ~\new_[9887]_  | ~\new_[11588]_  | ~\new_[11584]_  | ~\new_[9886]_ ;
  assign \s6_addr_o[7]  = ~\new_[9892]_  | ~\new_[11590]_  | ~\new_[11589]_  | ~\new_[9890]_ ;
  assign \s6_addr_o[6]  = ~\new_[9895]_  | ~\new_[11593]_  | ~\new_[11591]_  | ~\new_[11592]_ ;
  assign \s6_addr_o[1]  = ~\new_[9906]_  | ~\new_[13476]_  | ~\new_[11606]_  | ~\new_[11608]_ ;
  assign \s6_sel_o[0]  = ~\new_[9913]_  | ~\new_[11623]_  | ~\new_[11621]_  | ~\new_[11622]_ ;
  assign \s7_data_o[29]  = ~\new_[14842]_  | ~\new_[9918]_  | ~\new_[11637]_  | ~\new_[11639]_ ;
  assign \s7_data_o[19]  = ~\new_[14857]_  | ~\new_[9938]_  | ~\new_[11664]_  | ~\new_[11665]_ ;
  assign \s7_data_o[18]  = ~\new_[9941]_  | ~\new_[11667]_  | ~\new_[11666]_  | ~\new_[13494]_ ;
  assign \s7_data_o[11]  = ~\new_[11679]_  | ~\new_[9959]_  | ~\new_[11678]_  | ~\new_[13507]_ ;
  assign \s7_data_o[10]  = ~\new_[14863]_  | ~\new_[9961]_  | ~\new_[11680]_  | ~\new_[9960]_ ;
  assign \s7_data_o[9]  = ~\new_[11682]_  | ~\new_[9963]_  | ~\new_[11681]_  | ~\new_[13509]_ ;
  assign \s7_data_o[8]  = ~\new_[14864]_  | ~\new_[9964]_  | ~\new_[11683]_  | ~\new_[11685]_ ;
  assign \s7_data_o[6]  = ~\new_[11688]_  | ~\new_[9969]_  | ~\new_[13512]_  | ~\new_[13511]_ ;
  assign \s7_data_o[3]  = ~\new_[9974]_  | ~\new_[11693]_  | ~\new_[11692]_  | ~\new_[13516]_ ;
  assign \s7_data_o[0]  = ~\new_[9981]_  | ~\new_[11700]_  | ~\new_[11698]_  | ~\new_[13519]_ ;
  assign \s7_addr_o[31]  = ~\new_[9982]_  | ~\new_[11702]_  | ~\new_[11701]_  | ~\new_[13520]_ ;
  assign \s7_addr_o[30]  = ~\new_[14870]_  | ~\new_[9984]_  | ~\new_[11703]_  | ~\new_[11704]_ ;
  assign \s7_addr_o[27]  = ~\new_[9995]_  | ~\new_[11711]_  | ~\new_[14874]_  | ~\new_[11710]_ ;
  assign \s7_addr_o[26]  = ~\new_[14875]_  | ~\new_[9996]_  | ~\new_[11713]_  | ~\new_[11714]_ ;
  assign \s7_addr_o[25]  = ~\new_[9997]_  | ~\new_[11716]_  | ~\new_[11715]_  | ~\new_[13524]_ ;
  assign \s7_addr_o[23]  = ~\new_[14879]_  | ~\new_[10003]_  | ~\new_[11719]_  | ~\new_[10000]_ ;
  assign \s7_addr_o[22]  = ~\new_[14881]_  | ~\new_[10004]_  | ~\new_[11720]_  | ~\new_[11721]_ ;
  assign \s7_addr_o[20]  = ~\new_[11727]_  | ~\new_[10010]_  | ~\new_[11726]_  | ~\new_[14883]_ ;
  assign \s7_addr_o[18]  = ~\new_[14886]_  | ~\new_[10011]_  | ~\new_[11732]_  | ~\new_[11733]_ ;
  assign \s7_addr_o[17]  = ~\new_[14887]_  | ~\new_[10012]_  | ~\new_[11734]_  | ~\new_[11735]_ ;
  assign \s7_addr_o[8]  = ~\new_[10023]_  | ~\new_[11770]_  | ~\new_[11768]_  | ~\new_[13537]_ ;
  assign \s7_addr_o[5]  = ~\new_[10031]_  | ~\new_[11777]_  | ~\new_[11776]_  | ~\new_[13541]_ ;
  assign \s7_addr_o[4]  = ~\new_[10034]_  | ~\new_[11780]_  | ~\new_[11779]_  | ~\new_[13542]_ ;
  assign \s7_addr_o[3]  = ~\new_[10039]_  | ~\new_[11782]_  | ~\new_[11781]_  | ~\new_[13543]_ ;
  assign \s7_addr_o[2]  = ~\new_[10041]_  | ~\new_[11784]_  | ~\new_[13544]_  | ~\new_[11783]_ ;
  assign \s7_addr_o[0]  = ~\new_[11789]_  | ~\new_[10046]_  | ~\new_[14896]_  | ~\new_[10044]_ ;
  assign \s8_data_o[29]  = ~\new_[10059]_  | ~\new_[10061]_  | ~\new_[10058]_  | ~\new_[8964]_ ;
  assign \s8_data_o[27]  = ~\new_[10068]_  | ~\new_[10070]_  | ~\new_[10066]_  | ~\new_[8968]_ ;
  assign \s8_data_o[25]  = ~\new_[10074]_  | ~\new_[10075]_  | ~\new_[10073]_  | ~\new_[8973]_ ;
  assign \s8_data_o[23]  = ~\new_[10079]_  | ~\new_[10082]_  | ~\new_[10078]_  | ~\new_[8977]_ ;
  assign \s8_data_o[17]  = ~\new_[10094]_  | ~\new_[10096]_  | ~\new_[10093]_  | ~\new_[8991]_ ;
  assign \s8_data_o[16]  = ~\new_[10099]_  | ~\new_[10100]_  | ~\new_[10098]_  | ~\new_[8994]_ ;
  assign \s8_data_o[15]  = ~\new_[11836]_  | ~\new_[10102]_  | ~\new_[10101]_  | ~\new_[8995]_ ;
  assign \s8_data_o[13]  = ~\new_[10106]_  | ~\new_[10107]_  | ~\new_[10105]_  | ~\new_[9001]_ ;
  assign \s8_data_o[12]  = ~\new_[10111]_  | ~\new_[10112]_  | ~\new_[10108]_  | ~\new_[10109]_ ;
  assign \s8_data_o[11]  = ~\new_[10115]_  | ~\new_[10116]_  | ~\new_[10113]_  | ~\new_[10114]_ ;
  assign \s8_data_o[10]  = ~\new_[11846]_  | ~\new_[10121]_  | ~\new_[10117]_  | ~\new_[10118]_ ;
  assign \s8_data_o[9]  = ~\new_[11850]_  | ~\new_[10124]_  | ~\new_[10122]_  | ~\new_[10123]_ ;
  assign \s8_data_o[7]  = ~\new_[11858]_  | ~\new_[10129]_  | ~\new_[10127]_  | ~\new_[9010]_ ;
  assign \s8_data_o[6]  = ~\new_[10133]_  | ~\new_[10134]_  | ~\new_[10132]_  | ~\new_[9012]_ ;
  assign \s8_data_o[5]  = ~\new_[11861]_  | ~\new_[10139]_  | ~\new_[10135]_  | ~\new_[9014]_ ;
  assign \s8_data_o[2]  = ~\new_[11868]_  | ~\new_[10146]_  | ~\new_[10145]_  | ~\new_[9022]_ ;
  assign \s8_addr_o[21]  = ~\new_[10167]_  | ~\new_[10170]_  | ~\new_[10166]_  | ~\new_[9069]_ ;
  assign \s8_addr_o[18]  = ~\new_[10186]_  | ~\new_[10185]_  | ~\new_[10183]_  | ~\new_[9077]_ ;
  assign \s8_addr_o[16]  = ~\new_[10193]_  | ~\new_[10194]_  | ~\new_[10192]_  | ~\new_[9081]_ ;
  assign \s8_addr_o[14]  = ~\new_[10200]_  | ~\new_[10202]_  | ~\new_[10199]_  | ~\new_[9084]_ ;
  assign \s8_addr_o[13]  = ~\new_[10206]_  | ~\new_[10207]_  | ~\new_[10205]_  | ~\new_[9085]_ ;
  assign \s8_addr_o[11]  = ~\new_[10211]_  | ~\new_[10213]_  | ~\new_[10210]_  | ~\new_[9090]_ ;
  assign \s8_addr_o[9]  = ~\new_[11913]_  | ~\new_[10218]_  | ~\new_[10217]_  | ~\new_[9094]_ ;
  assign \s8_addr_o[10]  = ~\new_[10215]_  | ~\new_[10216]_  | ~\new_[10214]_  | ~\new_[9093]_ ;
  assign \s8_addr_o[7]  = ~\new_[10223]_  | ~\new_[10225]_  | ~\new_[10222]_  | ~\new_[9099]_ ;
  assign \s8_addr_o[6]  = ~\new_[11918]_  | ~\new_[10227]_  | ~\new_[10226]_  | ~\new_[9101]_ ;
  assign \s8_addr_o[5]  = ~\new_[11919]_  | ~\new_[10230]_  | ~\new_[10228]_  | ~\new_[9103]_ ;
  assign \s8_addr_o[3]  = ~\new_[11924]_  | ~\new_[10237]_  | ~\new_[10235]_  | ~\new_[9106]_ ;
  assign \s8_addr_o[1]  = ~\new_[10242]_  | ~\new_[10244]_  | ~\new_[10241]_  | ~\new_[9108]_ ;
  assign \s8_sel_o[1]  = ~\new_[10250]_  | ~\new_[10251]_  | ~\new_[10249]_  | ~\new_[9121]_ ;
  assign s8_we_o = ~\new_[10256]_  | ~\new_[10257]_  | ~\new_[9821]_  | ~\new_[9126]_ ;
  assign \s9_data_o[29]  = ~\new_[11936]_  | ~\new_[10269]_  | ~\new_[10264]_  | ~\new_[10266]_ ;
  assign \s9_data_o[28]  = ~\new_[10272]_  | ~\new_[10273]_  | ~\new_[10270]_  | ~\new_[10271]_ ;
  assign \s9_data_o[27]  = ~\new_[10276]_  | ~\new_[10278]_  | ~\new_[10274]_  | ~\new_[10275]_ ;
  assign \s9_data_o[23]  = ~\new_[10290]_  | ~\new_[9817]_  | ~\new_[10288]_  | ~\new_[10289]_ ;
  assign \s9_data_o[21]  = ~\new_[14948]_  | ~\new_[10295]_  | ~\new_[9144]_  | ~\new_[10294]_ ;
  assign \s9_data_o[19]  = ~\new_[10299]_  | ~\new_[10300]_  | ~\new_[10298]_  | ~\new_[9148]_ ;
  assign \s9_data_o[16]  = ~\new_[11948]_  | ~\new_[10310]_  | ~\new_[10309]_  | ~\new_[9154]_ ;
  assign \s9_data_o[15]  = ~\new_[10313]_  | ~\new_[10314]_  | ~\new_[9155]_  | ~\new_[10312]_ ;
  assign \s9_data_o[13]  = ~\new_[10319]_  | ~\new_[10320]_  | ~\new_[9158]_  | ~\new_[10318]_ ;
  assign \s9_data_o[12]  = ~\new_[10322]_  | ~\new_[10323]_  | ~\new_[9160]_  | ~\new_[10321]_ ;
  assign \s9_data_o[11]  = ~\new_[13643]_  | ~\new_[10324]_  | ~\new_[9162]_  | ~\new_[9163]_ ;
  assign \s9_data_o[10]  = ~\new_[10326]_  | ~\new_[14951]_  | ~\new_[9164]_  | ~\new_[10325]_ ;
  assign \s9_data_o[9]  = ~\new_[10329]_  | ~\new_[10328]_  | ~\new_[9166]_  | ~\new_[10327]_ ;
  assign \s9_data_o[8]  = ~\new_[10332]_  | ~\new_[10333]_  | ~\new_[10331]_  | ~\new_[10330]_ ;
  assign \s9_data_o[7]  = ~\new_[10336]_  | ~\new_[14954]_  | ~\new_[9169]_  | ~\new_[10335]_ ;
  assign \s9_data_o[4]  = ~\new_[13646]_  | ~\new_[10343]_  | ~\new_[9177]_  | ~\new_[9178]_ ;
  assign \s9_data_o[2]  = ~\new_[14955]_  | ~\new_[10349]_  | ~\new_[9184]_  | ~\new_[10348]_ ;
  assign \s9_data_o[0]  = ~\new_[10355]_  | ~\new_[10356]_  | ~\new_[9188]_  | ~\new_[10353]_ ;
  assign \s9_addr_o[31]  = ~\new_[10360]_  | ~\new_[10362]_  | ~\new_[10357]_  | ~\new_[9191]_ ;
  assign \s9_addr_o[29]  = ~\new_[10365]_  | ~\new_[10366]_  | ~\new_[9195]_  | ~\new_[9196]_ ;
  assign \s9_addr_o[26]  = ~\new_[14992]_  | ~\new_[10372]_  | ~\new_[9205]_  | ~\new_[9206]_ ;
  assign \s9_addr_o[23]  = ~\new_[10380]_  | ~\new_[10381]_  | ~\new_[10378]_  | ~\new_[9211]_ ;
  assign \s9_addr_o[22]  = ~\new_[11994]_  | ~\new_[10384]_  | ~\new_[9215]_  | ~\new_[10383]_ ;
  assign \s9_addr_o[20]  = ~\new_[10390]_  | ~\new_[12001]_  | ~\new_[9225]_  | ~\new_[10389]_ ;
  assign \s9_addr_o[18]  = ~\new_[10396]_  | ~\new_[13665]_  | ~\new_[9228]_  | ~\new_[9229]_ ;
  assign \s9_addr_o[17]  = ~\new_[12013]_  | ~\new_[10401]_  | ~\new_[9230]_  | ~\new_[10399]_ ;
  assign \s9_addr_o[16]  = ~\new_[12016]_  | ~\new_[10405]_  | ~\new_[9231]_  | ~\new_[10403]_ ;
  assign \s9_addr_o[11]  = ~\new_[10423]_  | ~\new_[10424]_  | ~\new_[9242]_  | ~\new_[10421]_ ;
  assign \s9_addr_o[8]  = ~\new_[12050]_  | ~\new_[10434]_  | ~\new_[10433]_  | ~\new_[9250]_ ;
  assign \s9_addr_o[7]  = ~\new_[10436]_  | ~\new_[12053]_  | ~\new_[9252]_  | ~\new_[9253]_ ;
  assign \s9_addr_o[6]  = ~\new_[12057]_  | ~\new_[10442]_  | ~\new_[10438]_  | ~\new_[9254]_ ;
  assign \s9_addr_o[4]  = ~\new_[10448]_  | ~\new_[10449]_  | ~\new_[9257]_  | ~\new_[10447]_ ;
  assign \s9_addr_o[3]  = ~\new_[10450]_  | ~\new_[10452]_  | ~\new_[9357]_  | ~\new_[13683]_ ;
  assign \s9_sel_o[3]  = ~\new_[12074]_  | ~\new_[10461]_  | ~\new_[10460]_  | ~\new_[9267]_ ;
  assign \s9_sel_o[1]  = ~\new_[12078]_  | ~\new_[10466]_  | ~\new_[9270]_  | ~\new_[9272]_ ;
  assign s0_cyc_o = ~n7499;
  assign s10_stb_o = \new_[10970]_  | \new_[8539]_ ;
  assign \s11_data_o[31]  = ~\new_[15122]_  | ~\new_[10546]_  | ~\new_[13845]_  | ~\new_[12564]_ ;
  assign \s11_data_o[27]  = ~\new_[10551]_  | ~\new_[15130]_  | ~\new_[11934]_  | ~\new_[12316]_ ;
  assign \s11_data_o[25]  = ~\new_[14831]_  | ~\new_[10553]_  | ~\new_[12323]_  | ~\new_[12325]_ ;
  assign \s11_data_o[23]  = ~\new_[15142]_  | ~\new_[10556]_  | ~\new_[12330]_  | ~\new_[12332]_ ;
  assign \s11_data_o[22]  = ~\new_[14825]_  | ~\new_[10558]_  | ~\new_[12333]_  | ~\new_[12335]_ ;
  assign \s11_data_o[21]  = ~\new_[15146]_  | ~\new_[10559]_  | ~\new_[12569]_  | ~\new_[12338]_ ;
  assign \s11_data_o[20]  = ~\new_[15149]_  | ~\new_[10560]_  | ~\new_[12340]_  | ~\new_[12341]_ ;
  assign \s11_data_o[19]  = ~\new_[15152]_  | ~\new_[10561]_  | ~\new_[12343]_  | ~\new_[12578]_ ;
  assign \s11_data_o[17]  = ~\new_[10563]_  | ~\new_[10564]_  | ~\new_[13873]_  | ~\new_[15157]_ ;
  assign \s11_data_o[16]  = ~\new_[15160]_  | ~\new_[10565]_  | ~\new_[12353]_  | ~\new_[12354]_ ;
  assign \s11_data_o[14]  = ~\new_[15165]_  | ~\new_[10570]_  | ~\new_[13882]_  | ~\new_[10569]_ ;
  assign \s11_data_o[13]  = ~\new_[15166]_  | ~\new_[10571]_  | ~\new_[13887]_  | ~\new_[10917]_ ;
  assign \s11_data_o[12]  = ~\new_[15171]_  | ~\new_[10572]_  | ~\new_[12358]_  | ~\new_[12359]_ ;
  assign \s11_data_o[11]  = ~\new_[13894]_  | ~\new_[10573]_  | ~\new_[12436]_  | ~\new_[15174]_ ;
  assign \s11_data_o[9]  = ~\new_[15641]_  | ~\new_[10576]_  | ~\new_[13899]_  | ~\new_[10575]_ ;
  assign \s11_data_o[7]  = ~\new_[13908]_  | ~\new_[10577]_  | ~\new_[12370]_  | ~\new_[15183]_ ;
  assign \s11_data_o[4]  = ~\new_[15193]_  | ~\new_[10368]_  | ~\new_[10581]_  | ~\new_[12378]_ ;
  assign \s11_data_o[3]  = ~\new_[10584]_  | ~\new_[15198]_  | ~\new_[12380]_  | ~\new_[10582]_ ;
  assign \s11_data_o[1]  = ~\new_[13925]_  | ~\new_[10586]_  | ~\new_[10047]_  | ~\new_[15201]_ ;
  assign \s11_data_o[0]  = ~\new_[10587]_  | ~\new_[9650]_  | ~\new_[14402]_  | ~\new_[15204]_ ;
  assign \s11_addr_o[30]  = ~\new_[15210]_  | ~\new_[10589]_  | ~\new_[13930]_  | ~\new_[9325]_ ;
  assign \s11_addr_o[29]  = ~\new_[10590]_  | ~\new_[12393]_  | ~\new_[12392]_  | ~\new_[15213]_ ;
  assign \s11_addr_o[31]  = ~\new_[12389]_  | ~\new_[15207]_  | ~\new_[13929]_  | ~\new_[9324]_ ;
  assign \s11_addr_o[25]  = ~\new_[12406]_  | ~\new_[15226]_  | ~\new_[13946]_  | ~\new_[9331]_ ;
  assign \s11_addr_o[22]  = ~\new_[10592]_  | ~\new_[10594]_  | ~\new_[13955]_  | ~\new_[15234]_ ;
  assign \s11_addr_o[19]  = ~\new_[12427]_  | ~\new_[10597]_  | ~\new_[15242]_  | ~\new_[12426]_ ;
  assign \s11_addr_o[18]  = ~\new_[12429]_  | ~\new_[10598]_  | ~\new_[15245]_  | ~\new_[12428]_ ;
  assign \s11_addr_o[17]  = ~\new_[12433]_  | ~\new_[10599]_  | ~\new_[13690]_  | ~\new_[15248]_ ;
  assign \s11_addr_o[16]  = ~\new_[10601]_  | ~\new_[9619]_  | ~\new_[15252]_  | ~\new_[12434]_ ;
  assign \s11_addr_o[12]  = ~\new_[10604]_  | ~\new_[10605]_  | ~\new_[15262]_  | ~\new_[12444]_ ;
  assign \s11_addr_o[10]  = ~\new_[15268]_  | ~\new_[10607]_  | ~\new_[12449]_  | ~\new_[12450]_ ;
  assign \s11_addr_o[8]  = ~\new_[11537]_  | ~\new_[10612]_  | ~\new_[14567]_  | ~\new_[12455]_ ;
  assign \s11_addr_o[7]  = ~\new_[13983]_  | ~\new_[10613]_  | ~\new_[12457]_  | ~\new_[15272]_ ;
  assign \s11_addr_o[4]  = ~\new_[15279]_  | ~\new_[10618]_  | ~\new_[12467]_  | ~\new_[12468]_ ;
  assign \s11_addr_o[3]  = ~\new_[10619]_  | ~\new_[14522]_  | ~\new_[13056]_  | ~\new_[12472]_ ;
  assign \s11_addr_o[2]  = ~\new_[13988]_  | ~\new_[10621]_  | ~\new_[15282]_  | ~\new_[9618]_ ;
  assign \s11_addr_o[1]  = ~\new_[12478]_  | ~\new_[10623]_  | ~\new_[15284]_  | ~\new_[12477]_ ;
  assign \s11_addr_o[0]  = ~\new_[15286]_  | ~\new_[10624]_  | ~\new_[12480]_  | ~\new_[11168]_ ;
  assign \s11_sel_o[2]  = ~\new_[13992]_  | ~\new_[10626]_  | ~\new_[12484]_  | ~\new_[14505]_ ;
  assign \s11_sel_o[1]  = ~\new_[10628]_  | ~\new_[15291]_  | ~\new_[13101]_  | ~\new_[12488]_ ;
  assign \s11_sel_o[0]  = ~\new_[12491]_  | ~\new_[10631]_  | ~\new_[15294]_  | ~\new_[12489]_ ;
  assign s11_stb_o = \new_[8540]_  | \new_[10974]_ ;
  assign \s12_data_o[31]  = ~\new_[13577]_  | ~\new_[10635]_  | ~\new_[9338]_  | ~\new_[15299]_ ;
  assign \s12_data_o[30]  = ~\new_[15300]_  | ~\new_[10636]_  | ~\new_[12501]_  | ~\new_[9339]_ ;
  assign \s12_data_o[29]  = ~\new_[10638]_  | ~\new_[10639]_  | ~\new_[15301]_  | ~\new_[12502]_ ;
  assign s12_cyc_o = ~n7464;
  assign \s12_data_o[26]  = ~\new_[12506]_  | ~\new_[10644]_  | ~\new_[15308]_  | ~\new_[9343]_ ;
  assign \s12_data_o[25]  = ~\new_[15311]_  | ~\new_[10514]_  | ~\new_[9345]_  | ~\new_[14013]_ ;
  assign \s12_data_o[24]  = ~\new_[10648]_  | ~\new_[14016]_  | ~\new_[15312]_  | ~\new_[10646]_ ;
  assign \s12_data_o[23]  = ~\new_[10649]_  | ~\new_[10650]_  | ~\new_[15316]_  | ~\new_[12509]_ ;
  assign \s12_data_o[22]  = ~\new_[10182]_  | ~\new_[15317]_  | ~\new_[10547]_  | ~\new_[13660]_ ;
  assign \s12_data_o[21]  = ~\new_[14733]_  | ~\new_[14021]_  | ~\new_[10651]_  | ~\new_[9347]_ ;
  assign \s12_data_o[20]  = ~\new_[10552]_  | ~\new_[10656]_  | ~\new_[12514]_  | ~\new_[15319]_ ;
  assign \s12_data_o[19]  = ~\new_[14023]_  | ~\new_[10658]_  | ~\new_[9348]_  | ~\new_[15323]_ ;
  assign \s12_data_o[18]  = ~\new_[14024]_  | ~\new_[10659]_  | ~\new_[14868]_  | ~\new_[8702]_ ;
  assign \s12_data_o[17]  = ~\new_[14027]_  | ~\new_[10661]_  | ~\new_[15324]_  | ~\new_[9349]_ ;
  assign \s12_data_o[16]  = ~\new_[9622]_  | ~\new_[15328]_  | ~\new_[12518]_  | ~\new_[10662]_ ;
  assign \s12_data_o[11]  = ~\new_[12526]_  | ~\new_[12527]_  | ~\new_[15337]_  | ~\new_[9356]_ ;
  assign \s12_data_o[4]  = ~\new_[13218]_  | ~\new_[10672]_  | ~\new_[8769]_  | ~\new_[15354]_ ;
  assign \s12_data_o[3]  = ~\new_[10673]_  | ~\new_[14045]_  | ~\new_[10557]_  | ~\new_[15357]_ ;
  assign \s12_data_o[2]  = ~\new_[14047]_  | ~\new_[12785]_  | ~\new_[15361]_  | ~\new_[9362]_ ;
  assign \s12_data_o[0]  = ~\new_[11820]_  | ~\new_[12543]_  | ~\new_[14956]_  | ~\new_[9363]_ ;
  assign \s12_addr_o[31]  = ~\new_[10678]_  | ~\new_[14053]_  | ~\new_[15368]_  | ~\new_[10677]_ ;
  assign \s12_addr_o[30]  = ~\new_[14054]_  | ~\new_[10680]_  | ~\new_[9725]_  | ~\new_[15372]_ ;
  assign \s12_addr_o[29]  = ~\new_[15715]_  | ~\new_[10683]_  | ~\new_[10681]_  | ~\new_[11212]_ ;
  assign \s12_addr_o[27]  = ~\new_[15384]_  | ~\new_[10204]_  | ~\new_[12274]_  | ~\new_[10686]_ ;
  assign \s12_addr_o[25]  = ~\new_[10036]_  | ~\new_[15390]_  | ~\new_[12549]_  | ~\new_[10689]_ ;
  assign \s12_addr_o[23]  = ~\new_[10693]_  | ~\new_[15395]_  | ~\new_[12551]_  | ~\new_[10692]_ ;
  assign \s12_addr_o[22]  = ~\new_[10694]_  | ~\new_[15397]_  | ~\new_[9364]_  | ~\new_[14074]_ ;
  assign \s12_addr_o[21]  = ~\new_[10819]_  | ~\new_[13242]_  | ~\new_[9396]_  | ~\new_[15399]_ ;
  assign s13_cyc_o = ~n7469;
  assign \s12_addr_o[20]  = ~\new_[10695]_  | ~\new_[14076]_  | ~\new_[10593]_  | ~\new_[15402]_ ;
  assign \s12_addr_o[17]  = ~\new_[15408]_  | ~\new_[10701]_  | ~\new_[10699]_  | ~\new_[14081]_ ;
  assign \s12_addr_o[18]  = ~\new_[13185]_  | ~\new_[10698]_  | ~\new_[15405]_  | ~\new_[10697]_ ;
  assign \s12_addr_o[9]  = ~\new_[11095]_  | ~\new_[10710]_  | ~\new_[12574]_  | ~\new_[15434]_ ;
  assign \s12_addr_o[10]  = ~\new_[15431]_  | ~\new_[14490]_  | ~\new_[10709]_  | ~\new_[9381]_ ;
  assign \s12_addr_o[5]  = ~\new_[15446]_  | ~\new_[11079]_  | ~\new_[10716]_  | ~\new_[12586]_ ;
  assign \s12_addr_o[3]  = ~\new_[14937]_  | ~\new_[10721]_  | ~\new_[10720]_  | ~\new_[12588]_ ;
  assign \s12_addr_o[4]  = ~\new_[15449]_  | ~\new_[10718]_  | ~\new_[10929]_  | ~\new_[14104]_ ;
  assign \s12_sel_o[0]  = ~\new_[15463]_  | ~\new_[10726]_  | ~\new_[10954]_  | ~\new_[12601]_ ;
  assign s12_we_o = ~\new_[15466]_  | ~\new_[10728]_  | ~\new_[10727]_  | ~\new_[14117]_ ;
  assign \s13_data_o[31]  = ~\new_[10730]_  | ~\new_[10731]_  | ~\new_[11914]_  | ~\new_[10729]_ ;
  assign \s13_data_o[30]  = ~\new_[10733]_  | ~\new_[10735]_  | ~\new_[11503]_  | ~\new_[10732]_ ;
  assign \s13_data_o[29]  = ~\new_[10737]_  | ~\new_[10736]_  | ~\new_[12826]_  | ~\new_[11130]_ ;
  assign s14_cyc_o = ~n7474;
  assign \s13_data_o[28]  = ~\new_[10136]_  | ~\new_[10739]_  | ~\new_[12614]_  | ~\new_[12615]_ ;
  assign \s13_data_o[27]  = ~\new_[10168]_  | ~\new_[10742]_  | ~\new_[12202]_  | ~\new_[10740]_ ;
  assign \s13_data_o[26]  = ~\new_[10745]_  | ~\new_[10746]_  | ~\new_[12620]_  | ~\new_[10743]_ ;
  assign \s13_data_o[25]  = ~\new_[10747]_  | ~\new_[10748]_  | ~\new_[12623]_  | ~\new_[12624]_ ;
  assign \s13_data_o[24]  = ~\new_[10750]_  | ~\new_[10751]_  | ~\new_[12626]_  | ~\new_[10749]_ ;
  assign \s13_data_o[19]  = ~\new_[10761]_  | ~\new_[10762]_  | ~\new_[12650]_  | ~\new_[10760]_ ;
  assign \s13_data_o[18]  = ~\new_[10763]_  | ~\new_[10764]_  | ~\new_[12656]_  | ~\new_[12657]_ ;
  assign \s13_data_o[17]  = ~\new_[10765]_  | ~\new_[10766]_  | ~\new_[12661]_  | ~\new_[12663]_ ;
  assign \s13_data_o[16]  = ~\new_[10768]_  | ~\new_[10769]_  | ~\new_[12664]_  | ~\new_[12666]_ ;
  assign \s13_data_o[15]  = ~\new_[10771]_  | ~\new_[10772]_  | ~\new_[12668]_  | ~\new_[10770]_ ;
  assign \s13_data_o[14]  = ~\new_[10774]_  | ~\new_[10775]_  | ~\new_[12670]_  | ~\new_[10773]_ ;
  assign \s13_data_o[13]  = ~\new_[10776]_  | ~\new_[14163]_  | ~\new_[12674]_  | ~\new_[12675]_ ;
  assign \s13_data_o[12]  = ~\new_[10779]_  | ~\new_[14165]_  | ~\new_[10777]_  | ~\new_[12678]_ ;
  assign \s13_data_o[10]  = ~\new_[14172]_  | ~\new_[10783]_  | ~\new_[10781]_  | ~\new_[10782]_ ;
  assign \s13_data_o[9]  = ~\new_[10785]_  | ~\new_[12683]_  | ~\new_[10784]_  | ~\new_[14175]_ ;
  assign \s13_data_o[7]  = ~\new_[10788]_  | ~\new_[10789]_  | ~\new_[12691]_  | ~\new_[10787]_ ;
  assign \s13_data_o[6]  = ~\new_[10791]_  | ~\new_[14181]_  | ~\new_[10790]_  | ~\new_[12694]_ ;
  assign \s13_data_o[4]  = ~\new_[10793]_  | ~\new_[12707]_  | ~\new_[12704]_  | ~\new_[10792]_ ;
  assign \s13_data_o[3]  = ~\new_[12709]_  | ~\new_[10794]_  | ~\new_[12708]_  | ~\new_[14187]_ ;
  assign \s13_data_o[0]  = ~\new_[10799]_  | ~\new_[10800]_  | ~\new_[12717]_  | ~\new_[10797]_ ;
  assign \s13_addr_o[31]  = ~\new_[10801]_  | ~\new_[10803]_  | ~\new_[12718]_  | ~\new_[12719]_ ;
  assign \s13_addr_o[30]  = ~\new_[10805]_  | ~\new_[14204]_  | ~\new_[12722]_  | ~\new_[10804]_ ;
  assign \s13_addr_o[28]  = ~\new_[10812]_  | ~\new_[12729]_  | ~\new_[12727]_  | ~\new_[10810]_ ;
  assign \s13_addr_o[26]  = ~\new_[10815]_  | ~\new_[12736]_  | ~\new_[12734]_  | ~\new_[12735]_ ;
  assign \s13_addr_o[25]  = ~\new_[10818]_  | ~\new_[12740]_  | ~\new_[12737]_  | ~\new_[12738]_ ;
  assign \s13_addr_o[24]  = ~\new_[10821]_  | ~\new_[12744]_  | ~\new_[12741]_  | ~\new_[12742]_ ;
  assign \s13_addr_o[23]  = ~\new_[10824]_  | ~\new_[10825]_  | ~\new_[12745]_  | ~\new_[10823]_ ;
  assign \s13_addr_o[22]  = ~\new_[10829]_  | ~\new_[10830]_  | ~\new_[12746]_  | ~\new_[10828]_ ;
  assign \s13_addr_o[21]  = ~\new_[10833]_  | ~\new_[10834]_  | ~\new_[12749]_  | ~\new_[10832]_ ;
  assign \s13_addr_o[20]  = ~\new_[10836]_  | ~\new_[10837]_  | ~\new_[12752]_  | ~\new_[12753]_ ;
  assign \s13_addr_o[19]  = ~\new_[10839]_  | ~\new_[10840]_  | ~\new_[12754]_  | ~\new_[12755]_ ;
  assign \s13_addr_o[18]  = ~\new_[10842]_  | ~\new_[10843]_  | ~\new_[12758]_  | ~\new_[12759]_ ;
  assign \s13_addr_o[17]  = ~\new_[10844]_  | ~\new_[10845]_  | ~\new_[12763]_  | ~\new_[12764]_ ;
  assign \s13_addr_o[16]  = ~\new_[10847]_  | ~\new_[10848]_  | ~\new_[12766]_  | ~\new_[10846]_ ;
  assign \s13_addr_o[15]  = ~\new_[10850]_  | ~\new_[10851]_  | ~\new_[12768]_  | ~\new_[10849]_ ;
  assign \s13_addr_o[14]  = ~\new_[10853]_  | ~\new_[10854]_  | ~\new_[12769]_  | ~\new_[10852]_ ;
  assign \s13_addr_o[13]  = ~\new_[10856]_  | ~\new_[10857]_  | ~\new_[12772]_  | ~\new_[10855]_ ;
  assign \s13_addr_o[12]  = ~\new_[10859]_  | ~\new_[10860]_  | ~\new_[12773]_  | ~\new_[10858]_ ;
  assign \s13_addr_o[11]  = ~\new_[10862]_  | ~\new_[10863]_  | ~\new_[12775]_  | ~\new_[10861]_ ;
  assign \s13_addr_o[10]  = ~\new_[10866]_  | ~\new_[10867]_  | ~\new_[12778]_  | ~\new_[10864]_ ;
  assign \s13_addr_o[9]  = ~\new_[10869]_  | ~\new_[10870]_  | ~\new_[12780]_  | ~\new_[10868]_ ;
  assign \s13_addr_o[8]  = ~\new_[10872]_  | ~\new_[14259]_  | ~\new_[12782]_  | ~\new_[10871]_ ;
  assign \s13_addr_o[7]  = ~\new_[10873]_  | ~\new_[10874]_  | ~\new_[12786]_  | ~\new_[12788]_ ;
  assign \s13_addr_o[6]  = ~\new_[12792]_  | ~\new_[10876]_  | ~\new_[12790]_  | ~\new_[10875]_ ;
  assign \s13_addr_o[5]  = ~\new_[10878]_  | ~\new_[10879]_  | ~\new_[12794]_  | ~\new_[10877]_ ;
  assign \s13_addr_o[4]  = ~\new_[10881]_  | ~\new_[10882]_  | ~\new_[12798]_  | ~\new_[12799]_ ;
  assign \s13_addr_o[3]  = ~\new_[10884]_  | ~\new_[10885]_  | ~\new_[12800]_  | ~\new_[10883]_ ;
  assign \s13_addr_o[2]  = ~\new_[12805]_  | ~\new_[10886]_  | ~\new_[12803]_  | ~\new_[12804]_ ;
  assign \s13_addr_o[1]  = ~\new_[10888]_  | ~\new_[10889]_  | ~\new_[12807]_  | ~\new_[12808]_ ;
  assign \s13_addr_o[0]  = ~\new_[10891]_  | ~\new_[14275]_  | ~\new_[12810]_  | ~\new_[10890]_ ;
  assign \s13_sel_o[3]  = ~\new_[10893]_  | ~\new_[14278]_  | ~\new_[12812]_  | ~\new_[10892]_ ;
  assign \s13_sel_o[2]  = ~\new_[10895]_  | ~\new_[14283]_  | ~\new_[12816]_  | ~\new_[10894]_ ;
  assign \s13_sel_o[1]  = ~\new_[10898]_  | ~\new_[10897]_  | ~\new_[12818]_  | ~\new_[10896]_ ;
  assign \s13_sel_o[0]  = ~\new_[10900]_  | ~\new_[10901]_  | ~\new_[12819]_  | ~\new_[10899]_ ;
  assign s13_we_o = ~\new_[12823]_  | ~\new_[10903]_  | ~\new_[12821]_  | ~\new_[10902]_ ;
  assign s13_stb_o = \new_[9455]_  | \new_[8543]_ ;
  assign \s14_data_o[31]  = ~\new_[10907]_  | ~\new_[12830]_  | ~\new_[10905]_  | ~\new_[10906]_ ;
  assign \s14_data_o[30]  = ~\new_[10909]_  | ~\new_[10910]_  | ~\new_[10908]_  | ~\new_[12831]_ ;
  assign \s14_data_o[29]  = ~\new_[10912]_  | ~\new_[10913]_  | ~\new_[10911]_  | ~\new_[12833]_ ;
  assign \s14_data_o[28]  = ~\new_[10914]_  | ~\new_[12836]_  | ~\new_[9399]_  | ~\new_[9400]_ ;
  assign \s14_data_o[27]  = ~\new_[10916]_  | ~\new_[12838]_  | ~\new_[9401]_  | ~\new_[10915]_ ;
  assign \s14_data_o[25]  = ~\new_[10921]_  | ~\new_[12842]_  | ~\new_[10920]_  | ~\new_[9403]_ ;
  assign \s14_data_o[24]  = ~\new_[10923]_  | ~\new_[12845]_  | ~\new_[9405]_  | ~\new_[9406]_ ;
  assign \s14_data_o[26]  = ~\new_[10919]_  | ~\new_[12841]_  | ~\new_[9402]_  | ~\new_[10918]_ ;
  assign \s14_data_o[23]  = ~\new_[10924]_  | ~\new_[12847]_  | ~\new_[9407]_  | ~\new_[9408]_ ;
  assign \s14_data_o[22]  = ~\new_[10925]_  | ~\new_[12849]_  | ~\new_[9409]_  | ~\new_[9410]_ ;
  assign \s14_data_o[20]  = ~\new_[10932]_  | ~\new_[12852]_  | ~\new_[9412]_  | ~\new_[10931]_ ;
  assign \s14_data_o[19]  = ~\new_[12854]_  | ~\new_[10936]_  | ~\new_[10934]_  | ~\new_[10935]_ ;
  assign \s14_data_o[18]  = ~\new_[10940]_  | ~\new_[12857]_  | ~\new_[9414]_  | ~\new_[10938]_ ;
  assign \s14_data_o[17]  = ~\new_[10945]_  | ~\new_[12858]_  | ~\new_[10941]_  | ~\new_[10943]_ ;
  assign \s14_data_o[16]  = ~\new_[10948]_  | ~\new_[12859]_  | ~\new_[10946]_  | ~\new_[9417]_ ;
  assign \s14_data_o[15]  = ~\new_[10950]_  | ~\new_[12861]_  | ~\new_[10949]_  | ~\new_[9419]_ ;
  assign \s14_data_o[14]  = ~\new_[10952]_  | ~\new_[12864]_  | ~\new_[10951]_  | ~\new_[9422]_ ;
  assign \s14_data_o[13]  = ~\new_[10953]_  | ~\new_[12866]_  | ~\new_[9423]_  | ~\new_[9424]_ ;
  assign s3_cyc_o = ~n7479;
  assign \s14_data_o[12]  = ~\new_[10955]_  | ~\new_[12869]_  | ~\new_[9426]_  | ~\new_[9427]_ ;
  assign \s14_data_o[11]  = ~\new_[10956]_  | ~\new_[12871]_  | ~\new_[9428]_  | ~\new_[9429]_ ;
  assign \s14_data_o[8]  = ~\new_[10960]_  | ~\new_[12881]_  | ~\new_[9432]_  | ~\new_[9433]_ ;
  assign \s14_data_o[7]  = ~\new_[12882]_  | ~\new_[10962]_  | ~\new_[9435]_  | ~\new_[10961]_ ;
  assign \s14_data_o[6]  = ~\new_[10964]_  | ~\new_[12884]_  | ~\new_[9436]_  | ~\new_[10963]_ ;
  assign \s14_data_o[5]  = ~\new_[10966]_  | ~\new_[12885]_  | ~\new_[9437]_  | ~\new_[9438]_ ;
  assign \s14_data_o[4]  = ~\new_[12887]_  | ~\new_[10968]_  | ~\new_[10967]_  | ~\new_[9440]_ ;
  assign \s14_data_o[3]  = ~\new_[12889]_  | ~\new_[12890]_  | ~\new_[9441]_  | ~\new_[9443]_ ;
  assign \s14_data_o[2]  = ~\new_[10969]_  | ~\new_[12891]_  | ~\new_[9444]_  | ~\new_[9445]_ ;
  assign \s14_data_o[1]  = ~\new_[12892]_  | ~\new_[12893]_  | ~\new_[9446]_  | ~\new_[9447]_ ;
  assign \s14_data_o[0]  = ~\new_[10973]_  | ~\new_[12897]_  | ~\new_[10971]_  | ~\new_[9451]_ ;
  assign \s14_addr_o[31]  = ~\new_[10977]_  | ~\new_[12898]_  | ~\new_[10975]_  | ~\new_[10976]_ ;
  assign \s14_addr_o[30]  = ~\new_[10981]_  | ~\new_[12899]_  | ~\new_[10979]_  | ~\new_[10980]_ ;
  assign \s14_addr_o[29]  = ~\new_[10985]_  | ~\new_[12901]_  | ~\new_[10983]_  | ~\new_[10984]_ ;
  assign \s14_addr_o[28]  = ~\new_[10989]_  | ~\new_[12904]_  | ~\new_[10987]_  | ~\new_[10988]_ ;
  assign \s14_addr_o[27]  = ~\new_[10993]_  | ~\new_[12905]_  | ~\new_[10990]_  | ~\new_[10992]_ ;
  assign \s14_addr_o[26]  = ~\new_[10997]_  | ~\new_[12908]_  | ~\new_[10995]_  | ~\new_[10996]_ ;
  assign \s14_addr_o[25]  = ~\new_[11003]_  | ~\new_[12909]_  | ~\new_[11000]_  | ~\new_[11002]_ ;
  assign \s14_addr_o[24]  = ~\new_[11008]_  | ~\new_[12913]_  | ~\new_[11006]_  | ~\new_[11007]_ ;
  assign \s14_addr_o[23]  = ~\new_[11010]_  | ~\new_[12914]_  | ~\new_[11009]_  | ~\new_[9463]_ ;
  assign \s14_addr_o[22]  = ~\new_[11013]_  | ~\new_[12915]_  | ~\new_[11012]_  | ~\new_[9464]_ ;
  assign \s14_addr_o[21]  = ~\new_[11015]_  | ~\new_[12917]_  | ~\new_[9465]_  | ~\new_[9466]_ ;
  assign \s14_addr_o[20]  = ~\new_[11017]_  | ~\new_[12918]_  | ~\new_[9467]_  | ~\new_[9468]_ ;
  assign \s14_addr_o[19]  = ~\new_[11019]_  | ~\new_[12920]_  | ~\new_[9469]_  | ~\new_[9470]_ ;
  assign \s14_addr_o[18]  = ~\new_[11023]_  | ~\new_[12922]_  | ~\new_[11020]_  | ~\new_[11021]_ ;
  assign \s14_addr_o[17]  = ~\new_[11025]_  | ~\new_[12924]_  | ~\new_[9472]_  | ~\new_[11024]_ ;
  assign \s14_addr_o[16]  = ~\new_[11028]_  | ~\new_[12927]_  | ~\new_[9473]_  | ~\new_[11027]_ ;
  assign \s14_addr_o[15]  = ~\new_[12928]_  | ~\new_[11030]_  | ~\new_[9474]_  | ~\new_[11029]_ ;
  assign \s14_addr_o[13]  = ~\new_[11035]_  | ~\new_[12932]_  | ~\new_[11034]_  | ~\new_[9477]_ ;
  assign \s14_addr_o[12]  = ~\new_[11037]_  | ~\new_[12935]_  | ~\new_[11036]_  | ~\new_[9478]_ ;
  assign \s14_addr_o[11]  = ~\new_[11039]_  | ~\new_[12936]_  | ~\new_[9479]_  | ~\new_[9480]_ ;
  assign \s14_addr_o[9]  = ~\new_[11044]_  | ~\new_[12940]_  | ~\new_[9483]_  | ~\new_[11043]_ ;
  assign \s14_addr_o[8]  = ~\new_[11047]_  | ~\new_[12943]_  | ~\new_[9484]_  | ~\new_[11046]_ ;
  assign \s14_addr_o[7]  = ~\new_[11049]_  | ~\new_[12945]_  | ~\new_[9485]_  | ~\new_[11048]_ ;
  assign \s14_addr_o[6]  = ~\new_[11051]_  | ~\new_[12946]_  | ~\new_[9486]_  | ~\new_[9487]_ ;
  assign \s14_addr_o[5]  = ~\new_[12947]_  | ~\new_[12948]_  | ~\new_[9488]_  | ~\new_[9489]_ ;
  assign \new_[7205]_  = ~\new_[12553]_  & ~\new_[8470]_ ;
  assign \s14_addr_o[4]  = ~\new_[12950]_  | ~\new_[11055]_  | ~\new_[9490]_  | ~\new_[11054]_ ;
  assign \s14_addr_o[3]  = ~\new_[11057]_  | ~\new_[12952]_  | ~\new_[9491]_  | ~\new_[9492]_ ;
  assign \s14_addr_o[2]  = ~\new_[12955]_  | ~\new_[11060]_  | ~\new_[9493]_  | ~\new_[11058]_ ;
  assign \s14_addr_o[1]  = ~\new_[11062]_  | ~\new_[12958]_  | ~\new_[9494]_  | ~\new_[11061]_ ;
  assign \s14_addr_o[0]  = ~\new_[11066]_  | ~\new_[12961]_  | ~\new_[11064]_  | ~\new_[11065]_ ;
  assign \s14_sel_o[2]  = ~\new_[12965]_  | ~\new_[11071]_  | ~\new_[11069]_  | ~\new_[9496]_ ;
  assign \s14_sel_o[1]  = ~\new_[11072]_  | ~\new_[12967]_  | ~\new_[9497]_  | ~\new_[9498]_ ;
  assign \s14_sel_o[0]  = ~\new_[11074]_  | ~\new_[12970]_  | ~\new_[9499]_  | ~\new_[11073]_ ;
  assign s14_we_o = ~\new_[11077]_  | ~\new_[12972]_  | ~\new_[11076]_  | ~\new_[9500]_ ;
  assign \new_[7215]_  = ~\new_[8464]_  & ~\new_[9300]_ ;
  assign \new_[7216]_  = ~\new_[13697]_  & ~\new_[8465]_ ;
  assign s15_stb_o = ~\new_[11143]_  | ~\new_[11122]_  | ~\new_[11104]_  | ~\new_[11132]_ ;
  assign \new_[7218]_  = ~\new_[11146]_  | ~\new_[11106]_  | ~\new_[11138]_  | ~\new_[11125]_ ;
  assign \s15_addr_o[24]  = ~\new_[9717]_  | ~\new_[9828]_  | ~\new_[9744]_  | ~\new_[9776]_ ;
  assign \new_[7220]_  = ~\new_[15791]_  | ~\new_[11101]_  | ~\new_[9535]_  | ~\new_[13021]_ ;
  assign \new_[7221]_  = ~s5_next_reg;
  assign \new_[7222]_  = \\s14_msel_pri_out_reg[0] ;
  assign \s15_addr_o[27]  = ~\new_[9602]_  | ~\new_[9609]_  | ~\new_[11113]_  | ~\new_[11154]_ ;
  assign \new_[7224]_  = \\s4_msel_pri_out_reg[0] ;
  assign \s15_addr_o[25]  = ~\new_[10017]_  | ~\new_[9575]_  | ~\new_[9678]_  | ~\new_[9631]_ ;
  assign \s15_addr_o[26]  = ~\new_[9664]_  | ~\new_[9685]_  | ~\new_[11056]_  | ~\new_[9625]_ ;
  assign \new_[7227]_  = ~\new_[8614]_  & ~\new_[9537]_ ;
  assign \new_[7228]_  = ~\new_[8615]_  & ~\new_[11107]_ ;
  assign \new_[7229]_  = ~\new_[8618]_  & ~\new_[8619]_ ;
  assign \new_[7230]_  = ~\new_[8636]_  & ~\new_[8531]_ ;
  assign \new_[7231]_  = ~\new_[8621]_  & ~\new_[8622]_ ;
  assign \new_[7232]_  = ~\new_[8624]_  & ~\new_[8625]_ ;
  assign \new_[7233]_  = ~\new_[8628]_  & ~\new_[8629]_ ;
  assign \new_[7234]_  = ~\new_[8630]_  & ~\new_[9544]_ ;
  assign \new_[7235]_  = ~\new_[8646]_  & (~\new_[17138]_  | ~\new_[28064]_ );
  assign \new_[7236]_  = ~\new_[8648]_  & (~\new_[16227]_  | ~\new_[26672]_ );
  assign \new_[7237]_  = ~\new_[8650]_  & (~\new_[16230]_  | ~\new_[28971]_ );
  assign \new_[7238]_  = ~\new_[8651]_  & (~\new_[17143]_  | ~\new_[28629]_ );
  assign \new_[7239]_  = ~\new_[8107]_  & (~\new_[16228]_  | ~\new_[28827]_ );
  assign \new_[7240]_  = ~\new_[8109]_  & (~\new_[16236]_  | ~\new_[29362]_ );
  assign \new_[7241]_  = ~\new_[8110]_  & (~\new_[17147]_  | ~\new_[28662]_ );
  assign \new_[7242]_  = ~\new_[8111]_  & (~\new_[17145]_  | ~\new_[28156]_ );
  assign \new_[7243]_  = ~\new_[8113]_  & (~\new_[17150]_  | ~\new_[29348]_ );
  assign \new_[7244]_  = ~\new_[8116]_  & (~\new_[14819]_  | ~\new_[27999]_ );
  assign \new_[7245]_  = ~\new_[8117]_  & (~\new_[16239]_  | ~\new_[29085]_ );
  assign \new_[7246]_  = ~\new_[8119]_  & (~\new_[17142]_  | ~\new_[29265]_ );
  assign \new_[7247]_  = ~\new_[8121]_  & (~\new_[17141]_  | ~\new_[26977]_ );
  assign \new_[7248]_  = ~\new_[8122]_  & (~\new_[17948]_  | ~\new_[29353]_ );
  assign \new_[7249]_  = ~\new_[8124]_  & (~\new_[17154]_  | ~\new_[29373]_ );
  assign \new_[7250]_  = ~\new_[8125]_  & (~\new_[11483]_  | ~\new_[28970]_ );
  assign \new_[7251]_  = ~\new_[8126]_  & (~\new_[17155]_  | ~\new_[29542]_ );
  assign \new_[7252]_  = ~\new_[8129]_  & (~\new_[16242]_  | ~\new_[29155]_ );
  assign \new_[7253]_  = ~\new_[8645]_  & (~\new_[17013]_  | ~\new_[29090]_ );
  assign \new_[7254]_  = ~\new_[8647]_  & (~\new_[14759]_  | ~\new_[26786]_ );
  assign \new_[7255]_  = ~\new_[8649]_  & (~\new_[14762]_  | ~\new_[27085]_ );
  assign \new_[7256]_  = ~\new_[8652]_  & (~\new_[17056]_  | ~\new_[27852]_ );
  assign \new_[7257]_  = ~\new_[8108]_  & (~\new_[14779]_  | ~\new_[27814]_ );
  assign \new_[7258]_  = ~\new_[8112]_  & (~\new_[11419]_  | ~\new_[26455]_ );
  assign \new_[7259]_  = ~\new_[8114]_  & (~\new_[14769]_  | ~\new_[29283]_ );
  assign \new_[7260]_  = ~\new_[8115]_  & (~\new_[14793]_  | ~\new_[29073]_ );
  assign \new_[7261]_  = ~\new_[8118]_  & (~\new_[14767]_  | ~\new_[28117]_ );
  assign \new_[7262]_  = ~\new_[8120]_  & (~\new_[14768]_  | ~\new_[27939]_ );
  assign \new_[7263]_  = ~\new_[8123]_  & (~\new_[14813]_  | ~\new_[26711]_ );
  assign \new_[7264]_  = ~\new_[8127]_  & (~\new_[17114]_  | ~\new_[28058]_ );
  assign \new_[7265]_  = ~\new_[8128]_  & (~\new_[17112]_  | ~\new_[26259]_ );
  assign \new_[7266]_  = ~\new_[8313]_  & ~\new_[8936]_ ;
  assign \new_[7267]_  = ~\new_[8317]_  & ~\new_[8939]_ ;
  assign \new_[7268]_  = ~\new_[8345]_  & ~\new_[8965]_ ;
  assign \new_[7269]_  = ~\new_[8349]_  & ~\new_[8967]_ ;
  assign \new_[7270]_  = ~\new_[9875]_  & ~\new_[8431]_ ;
  assign \new_[7271]_  = ~\new_[8433]_  & ~\new_[9884]_ ;
  assign \new_[7272]_  = ~\new_[8434]_  & ~\new_[9889]_ ;
  assign \new_[7273]_  = ~\new_[8814]_  & ~\new_[8436]_ ;
  assign \new_[7274]_  = ~\new_[8437]_  & ~\new_[9909]_ ;
  assign \new_[7275]_  = ~\new_[11618]_  & ~\new_[8439]_ ;
  assign \new_[7276]_  = ~\new_[8440]_  & ~\new_[8870]_ ;
  assign \new_[7277]_  = ~\new_[8441]_  & ~\new_[8874]_ ;
  assign \new_[7278]_  = ~\new_[8879]_  & ~\new_[8443]_ ;
  assign \new_[7279]_  = ~\new_[9774]_  & ~\new_[8361]_ ;
  assign \new_[7280]_  = ~\new_[8705]_  & (~\new_[8986]_  | ~\new_[27903]_ );
  assign \new_[7281]_  = ~\new_[8293]_  & ~\new_[8392]_ ;
  assign \new_[7282]_  = ~\new_[9686]_  & (~\new_[8992]_  | ~\new_[27876]_ );
  assign \new_[7283]_  = ~\new_[8708]_  & (~\new_[8993]_  | ~\new_[27980]_ );
  assign \new_[7284]_  = ~\new_[8770]_  & ~\new_[8394]_ ;
  assign \new_[7285]_  = ~\new_[8709]_  & ~\new_[8395]_ ;
  assign \new_[7286]_  = ~\new_[9694]_  & (~\new_[8997]_  | ~\new_[27933]_ );
  assign \new_[7287]_  = ~\new_[8710]_  & (~\new_[8998]_  | ~\new_[24582]_ );
  assign \new_[7288]_  = ~\new_[8711]_  & (~\new_[8999]_  | ~\new_[27919]_ );
  assign \new_[7289]_  = ~\new_[8772]_  & ~\new_[8397]_ ;
  assign \new_[7290]_  = ~\new_[8715]_  & ~\new_[8398]_ ;
  assign \new_[7291]_  = ~\new_[9698]_  & (~\new_[9003]_  | ~\new_[26748]_ );
  assign \new_[7292]_  = ~\new_[8716]_  & (~\new_[9004]_  | ~\new_[28761]_ );
  assign \new_[7293]_  = ~\new_[9882]_  & ~\new_[8369]_ ;
  assign \new_[7294]_  = ~\new_[8773]_  & ~\new_[8400]_ ;
  assign \new_[7295]_  = ~\new_[8307]_  & ~\new_[8401]_ ;
  assign \new_[7296]_  = ~\new_[8718]_  & ~\new_[8402]_ ;
  assign \new_[7297]_  = ~\new_[9701]_  & (~\new_[9006]_  | ~\new_[29066]_ );
  assign \new_[7298]_  = (~\new_[11929]_  | ~\new_[28683]_ ) & (~\new_[9113]_  | ~\new_[29416]_ );
  assign \new_[7299]_  = ~\new_[11405]_  & (~\new_[9011]_  | ~\new_[23094]_ );
  assign \new_[7300]_  = ~\new_[8353]_  & (~\new_[11932]_  | ~\new_[26507]_ );
  assign \new_[7301]_  = ~\new_[22488]_  | ~\new_[10080]_  | ~\new_[19352]_  | ~\new_[10131]_ ;
  assign \new_[7302]_  = ~\new_[8359]_  & (~\new_[14919]_  | ~\new_[26507]_ );
  assign \new_[7303]_  = ~\new_[8312]_  & (~\new_[9013]_  | ~\new_[27837]_ );
  assign \new_[7304]_  = ~\new_[8816]_  & ~\new_[8372]_ ;
  assign \new_[7305]_  = ~\new_[8729]_  & (~\new_[9015]_  | ~\new_[23092]_ );
  assign \new_[7306]_  = ~\new_[9777]_  | ~\new_[11421]_  | ~\new_[14802]_  | ~\new_[16173]_ ;
  assign \new_[7307]_  = ~\new_[9780]_  | ~\new_[14791]_  | ~\new_[9742]_  | ~\new_[9779]_ ;
  assign \new_[7308]_  = ~\new_[8316]_  & (~\new_[9019]_  | ~\new_[29033]_ );
  assign \new_[7309]_  = ~\new_[8818]_  & ~\new_[8373]_ ;
  assign \new_[7310]_  = ~\new_[14683]_  | ~\new_[9788]_  | ~\new_[16109]_  | ~\new_[11436]_ ;
  assign \new_[7311]_  = ~\new_[8319]_  & ~\new_[8406]_ ;
  assign \new_[7312]_  = ~\new_[9715]_  & (~\new_[9027]_  | ~\new_[29196]_ );
  assign \new_[7313]_  = ~\new_[8737]_  & (~\new_[9030]_  | ~\new_[26946]_ );
  assign \new_[7314]_  = ~\new_[8738]_  & (~\new_[9031]_  | ~\new_[24628]_ );
  assign \new_[7315]_  = ~\new_[11616]_  & ~\new_[8376]_ ;
  assign \new_[7316]_  = ~\new_[8779]_  & ~\new_[8410]_ ;
  assign \new_[7317]_  = ~\new_[8739]_  & ~\new_[8411]_ ;
  assign \new_[7318]_  = ~\new_[9720]_  & (~\new_[9037]_  | ~\new_[26589]_ );
  assign \new_[7319]_  = ~\new_[8740]_  & (~\new_[9040]_  | ~\new_[29637]_ );
  assign \new_[7320]_  = ~\new_[9726]_  & (~\new_[9045]_  | ~\new_[26823]_ );
  assign \new_[7321]_  = ~\new_[9727]_  & (~\new_[9047]_  | ~\new_[27847]_ );
  assign \new_[7322]_  = ~\new_[8743]_  & (~\new_[9048]_  | ~\new_[28694]_ );
  assign \new_[7323]_  = ~\new_[8381]_  & ~\new_[9917]_ ;
  assign \new_[7324]_  = ~\new_[9813]_  & (~\new_[9049]_  | ~\new_[27847]_ );
  assign \new_[7325]_  = ~\new_[8781]_  & ~\new_[8414]_ ;
  assign \new_[7326]_  = ~\new_[8329]_  & ~\new_[8415]_ ;
  assign \new_[7327]_  = ~\new_[8745]_  & ~\new_[8416]_ ;
  assign \new_[7328]_  = ~\new_[9731]_  & (~\new_[9054]_  | ~\new_[27767]_ );
  assign \new_[7329]_  = ~\new_[8748]_  & (~\new_[9055]_  | ~\new_[29102]_ );
  assign \new_[7330]_  = ~\new_[8950]_  & ~\new_[8418]_ ;
  assign \new_[7331]_  = ~\new_[8331]_  & (~\new_[9056]_  | ~\new_[28047]_ );
  assign \new_[7332]_  = ~\new_[8783]_  & ~\new_[8419]_ ;
  assign \new_[7333]_  = ~\new_[8334]_  & ~\new_[8420]_ ;
  assign \new_[7334]_  = ~\new_[8750]_  & ~\new_[8421]_ ;
  assign \new_[7335]_  = ~\new_[8337]_  & (~\new_[10161]_  | ~\new_[26827]_ );
  assign \new_[7336]_  = ~\new_[8752]_  & (~\new_[9061]_  | ~\new_[28003]_ );
  assign \new_[7337]_  = ~\new_[9816]_  & ~\new_[8385]_ ;
  assign \new_[7338]_  = ~\new_[8753]_  & (~\new_[9063]_  | ~\new_[28101]_ );
  assign \new_[7339]_  = ~\new_[9740]_  & (~\new_[9068]_  | ~\new_[27819]_ );
  assign \new_[7340]_  = ~\new_[8757]_  & (~\new_[9070]_  | ~\new_[24501]_ );
  assign \new_[7341]_  = ~\new_[8388]_  & ~\new_[9933]_ ;
  assign \new_[7342]_  = ~\new_[9820]_  & (~\new_[9071]_  | ~\new_[24501]_ );
  assign \new_[7343]_  = ~\new_[8785]_  & ~\new_[8423]_ ;
  assign \new_[7344]_  = ~\new_[8344]_  & (~\new_[9074]_  | ~\new_[27924]_ );
  assign \new_[7345]_  = ~\new_[8829]_  & ~\new_[8389]_ ;
  assign \new_[7346]_  = ~\new_[8346]_  & ~\new_[8425]_ ;
  assign \new_[7347]_  = ~\new_[8764]_  & ~\new_[8426]_ ;
  assign \new_[7348]_  = (~\new_[8910]_  | ~\m4_data_i[31] ) & (~\new_[9923]_  | ~\m5_data_i[31] );
  assign \new_[7349]_  = (~\new_[8910]_  | ~\m4_data_i[30] ) & (~\new_[9923]_  | ~\m5_data_i[30] );
  assign \new_[7350]_  = (~\new_[32346]_  | ~\m0_data_i[29] ) & (~\new_[13487]_  | ~\m1_data_i[29] );
  assign \new_[7351]_  = (~\new_[8910]_  | ~\m4_data_i[28] ) & (~\new_[14850]_  | ~\m5_data_i[28] );
  assign \new_[7352]_  = (~\new_[8910]_  | ~\m4_data_i[27] ) & (~\new_[9923]_  | ~\m5_data_i[27] );
  assign \new_[7353]_  = (~\new_[8910]_  | ~\m4_data_i[26] ) & (~\new_[9923]_  | ~\m5_data_i[26] );
  assign \new_[7354]_  = (~\new_[13526]_  | ~\m4_data_i[25] ) & (~\new_[14850]_  | ~\m5_data_i[25] );
  assign \new_[7355]_  = ~\new_[8348]_  & (~\new_[9078]_  | ~\new_[28157]_ );
  assign \new_[7356]_  = (~\new_[8910]_  | ~\m4_data_i[24] ) & (~\new_[9923]_  | ~\m5_data_i[24] );
  assign \new_[7357]_  = ~\new_[8830]_  & ~\new_[8390]_ ;
  assign \new_[7358]_  = (~\new_[8910]_  | ~\m4_data_i[23] ) & (~\new_[9923]_  | ~\m5_data_i[23] );
  assign \new_[7359]_  = ~\new_[9751]_  & ~\new_[8428]_ ;
  assign \new_[7360]_  = (~\new_[8910]_  | ~\m4_data_i[20] ) & (~\new_[9923]_  | ~\m5_data_i[20] );
  assign \new_[7361]_  = ~\new_[8352]_  & (~\new_[10196]_  | ~\new_[28553]_ );
  assign \new_[7362]_  = ~\new_[8429]_  & ~\new_[8292]_ ;
  assign \new_[7363]_  = ~\new_[8886]_  & ~\new_[8297]_ ;
  assign \new_[7364]_  = (~\new_[8910]_  | ~\m4_data_i[18] ) & (~\new_[9923]_  | ~\m5_data_i[18] );
  assign \new_[7365]_  = ~\new_[8430]_  & ~\new_[8299]_ ;
  assign \new_[7366]_  = ~\new_[8432]_  & ~\new_[8301]_ ;
  assign \new_[7367]_  = ~\new_[8306]_  & ~\new_[8891]_ ;
  assign \new_[7368]_  = (~\new_[13526]_  | ~\m4_data_i[17] ) & (~\new_[14850]_  | ~\m5_data_i[17] );
  assign \new_[7369]_  = ~\new_[8310]_  & ~\new_[8435]_ ;
  assign \new_[7370]_  = ~\new_[8895]_  & ~\new_[8314]_ ;
  assign \new_[7371]_  = (~\new_[13526]_  | ~\m4_data_i[16] ) & (~\new_[14850]_  | ~\m5_data_i[16] );
  assign \new_[7372]_  = ~\new_[8318]_  & ~\new_[8899]_ ;
  assign \new_[7373]_  = ~\new_[8438]_  & ~\new_[8323]_ ;
  assign \new_[7374]_  = ~\new_[8904]_  & ~\new_[8328]_ ;
  assign \new_[7375]_  = ~\new_[8907]_  & ~\new_[8333]_ ;
  assign \new_[7376]_  = ~\new_[9732]_  & ~\new_[8442]_ ;
  assign \new_[7377]_  = ~\new_[8912]_  & ~\new_[8338]_ ;
  assign \new_[7378]_  = ~\new_[8915]_  & ~\new_[8342]_ ;
  assign \new_[7379]_  = ~\new_[8920]_  & ~\new_[8350]_ ;
  assign \new_[7380]_  = ~\new_[11911]_  & ~\new_[8393]_ ;
  assign \new_[7381]_  = ~\new_[11915]_  & ~\new_[8396]_ ;
  assign \new_[7382]_  = ~\new_[8771]_  & ~\new_[8366]_ ;
  assign \new_[7383]_  = ~\new_[11921]_  & ~\new_[8399]_ ;
  assign \new_[7384]_  = ~\new_[8811]_  & ~\new_[8354]_ ;
  assign \new_[7385]_  = ~\new_[10243]_  & ~\new_[8403]_ ;
  assign \new_[7386]_  = ~\new_[8357]_  & ~\new_[8360]_ ;
  assign \new_[7387]_  = ~\new_[10280]_  & ~\new_[8409]_ ;
  assign \new_[7388]_  = ~\new_[11941]_  & ~\new_[8412]_ ;
  assign \new_[7389]_  = ~\new_[11945]_  & ~\new_[8413]_ ;
  assign \new_[7390]_  = ~\new_[8355]_  & ~\new_[8382]_ ;
  assign \new_[7391]_  = ~\new_[11950]_  & ~\new_[8417]_ ;
  assign \new_[7392]_  = ~\new_[11959]_  & ~\new_[8422]_ ;
  assign \new_[7393]_  = (~\new_[13530]_  | ~\new_[31537]_ ) & (~\new_[13487]_  | ~\m1_addr_i[31] );
  assign \new_[7394]_  = (~\new_[13530]_  | ~\new_[31486]_ ) & (~\new_[13487]_  | ~\new_[31308]_ );
  assign \new_[7395]_  = (~\new_[8921]_  | ~\new_[31000]_ ) & (~\new_[13487]_  | ~\new_[31538]_ );
  assign \new_[7396]_  = (~\new_[13530]_  | ~\new_[31547]_ ) & (~\new_[13487]_  | ~\new_[31458]_ );
  assign \new_[7397]_  = (~\new_[8910]_  | ~\m4_addr_i[23] ) & (~\new_[9923]_  | ~\m5_addr_i[23] );
  assign \new_[7398]_  = (~\new_[8910]_  | ~\m4_addr_i[22] ) & (~\new_[9923]_  | ~\m5_addr_i[22] );
  assign \new_[7399]_  = (~\new_[8910]_  | ~\m4_addr_i[21] ) & (~\new_[9923]_  | ~\m5_addr_i[21] );
  assign \new_[7400]_  = ~\new_[18404]_  | ~\new_[10077]_  | ~\new_[21263]_  | ~\new_[14255]_ ;
  assign \new_[7401]_  = (~\new_[8910]_  | ~\m4_addr_i[20] ) & (~\new_[9923]_  | ~\m5_addr_i[20] );
  assign \new_[7402]_  = (~\new_[8910]_  | ~\m4_addr_i[19] ) & (~\new_[9923]_  | ~\m5_addr_i[19] );
  assign \new_[7403]_  = (~\new_[8910]_  | ~\m4_addr_i[18] ) & (~\new_[9923]_  | ~\m5_addr_i[18] );
  assign \new_[7404]_  = (~\new_[8910]_  | ~\m4_addr_i[16] ) & (~\new_[9923]_  | ~\m5_addr_i[16] );
  assign \new_[7405]_  = (~\new_[8910]_  | ~\m4_addr_i[15] ) & (~\new_[9923]_  | ~\m5_addr_i[15] );
  assign \new_[7406]_  = ~\new_[17378]_  | ~\new_[10083]_  | ~\new_[21293]_  | ~\new_[14289]_ ;
  assign \new_[7407]_  = (~\new_[8910]_  | ~\m4_addr_i[11] ) & (~\new_[9923]_  | ~\m5_addr_i[11] );
  assign \new_[7408]_  = (~\new_[8910]_  | ~\m4_addr_i[10] ) & (~\new_[9923]_  | ~\m5_addr_i[10] );
  assign \new_[7409]_  = (~\new_[8910]_  | ~\m4_addr_i[9] ) & (~\new_[9923]_  | ~\m5_addr_i[9] );
  assign \new_[7410]_  = (~\new_[8910]_  | ~\m4_addr_i[8] ) & (~\new_[9923]_  | ~\m5_addr_i[8] );
  assign \new_[7411]_  = (~\new_[8910]_  | ~\m4_addr_i[7] ) & (~\new_[9923]_  | ~\m5_addr_i[7] );
  assign \new_[7412]_  = (~\new_[8910]_  | ~\m4_addr_i[6] ) & (~\new_[9923]_  | ~\m5_addr_i[6] );
  assign \new_[7413]_  = ~\new_[18419]_  | ~\new_[10088]_  | ~\new_[20364]_  | ~\new_[14324]_ ;
  assign \new_[7414]_  = ~\new_[8445]_  | ~\new_[13552]_ ;
  assign \new_[7415]_  = (~\new_[8910]_  | ~\m4_addr_i[1] ) & (~\new_[9923]_  | ~\m5_addr_i[1] );
  assign \new_[7416]_  = ~\new_[8446]_  | ~\new_[11812]_ ;
  assign \new_[7417]_  = (~\new_[8910]_  | ~\m4_addr_i[0] ) & (~\new_[9923]_  | ~\m5_addr_i[0] );
  assign \new_[7418]_  = (~\new_[8910]_  | ~\m4_sel_i[3] ) & (~\new_[9923]_  | ~\m5_sel_i[3] );
  assign \new_[7419]_  = ~\new_[20285]_  | ~\new_[10130]_  | ~\new_[20386]_  | ~\new_[12796]_ ;
  assign \new_[7420]_  = (~\new_[8910]_  | ~\m4_sel_i[2] ) & (~\new_[9923]_  | ~\m5_sel_i[2] );
  assign \new_[7421]_  = (~\new_[32346]_  | ~\m0_sel_i[1] ) & (~\new_[13487]_  | ~\m1_sel_i[1] );
  assign \new_[7422]_  = (~\new_[8910]_  | ~\m4_sel_i[1] ) & (~\new_[9923]_  | ~\m5_sel_i[1] );
  assign \new_[7423]_  = (~\new_[32346]_  | ~\m0_sel_i[0] ) & (~\new_[13487]_  | ~\m1_sel_i[0] );
  assign \new_[7424]_  = (~\new_[13526]_  | ~\m4_sel_i[0] ) & (~\new_[9923]_  | ~\m5_sel_i[0] );
  assign \new_[7425]_  = ~\new_[19362]_  | (~\new_[10510]_  & ~\new_[28036]_ );
  assign \new_[7426]_  = ~\new_[19365]_  | (~\new_[10521]_  & ~\new_[28711]_ );
  assign \new_[7427]_  = ~\new_[20361]_  | (~\new_[10525]_  & ~\new_[27972]_ );
  assign \new_[7428]_  = ~\new_[10440]_  & ~\new_[9203]_ ;
  assign \new_[7429]_  = ~\new_[12005]_  & (~\new_[10798]_  | ~\new_[24493]_ );
  assign \new_[7430]_  = ~\new_[9365]_  & ~\new_[9212]_ ;
  assign \new_[7431]_  = ~\new_[9092]_  & ~\new_[12143]_ ;
  assign \new_[7432]_  = ~\new_[12458]_  & ~\new_[9294]_ ;
  assign n7439 = (~\new_[10535]_  & ~rst_i) | (~\new_[30931]_  & ~\new_[31564]_ );
  assign \new_[7434]_  = \\s15_msel_pri_out_reg[1] ;
  assign \new_[7435]_  = \\s10_msel_pri_out_reg[0] ;
  assign \new_[7436]_  = \\s2_msel_pri_out_reg[1] ;
  assign \new_[7437]_  = \\s1_msel_pri_out_reg[1] ;
  assign \new_[7438]_  = ~\new_[12008]_  & (~\new_[10802]_  | ~\new_[24481]_ );
  assign \new_[7439]_  = \\s7_msel_pri_out_reg[1] ;
  assign \new_[7440]_  = \\s0_msel_pri_out_reg[1] ;
  assign \new_[7441]_  = ~\new_[9366]_  & ~\new_[9213]_ ;
  assign s5_cyc_o = ~n7589;
  assign n7444 = (~\new_[10536]_  & ~rst_i) | (~\new_[31209]_  & ~\new_[31846]_ );
  assign \s12_data_o[5]  = ~\new_[15351]_  | ~\new_[12537]_  | ~\new_[9361]_  | ~\new_[14043]_ ;
  assign \new_[7445]_  = ~\new_[9293]_  & ~\new_[9086]_ ;
  assign \new_[7446]_  = ~\new_[12012]_  & (~\new_[10806]_  | ~\new_[24477]_ );
  assign \new_[7447]_  = ~\new_[9367]_  & ~\new_[9216]_ ;
  assign \new_[7448]_  = ~\new_[12061]_  & ~\new_[9095]_ ;
  assign \new_[7449]_  = ~\new_[12015]_  & (~\new_[10809]_  | ~\new_[27967]_ );
  assign \new_[7450]_  = ~\new_[12784]_  & ~\new_[9110]_ ;
  assign \new_[7451]_  = ~\new_[9368]_  & ~\new_[9217]_ ;
  assign n7484 = ~\new_[9262]_  & ~\new_[10457]_ ;
  assign \new_[7453]_  = ~\new_[9116]_  & ~\new_[12492]_ ;
  assign \s0_data_o[31]  = ~\new_[11976]_  | ~\new_[11977]_  | ~\new_[9199]_  | ~\new_[11973]_ ;
  assign \s0_data_o[28]  = ~\new_[12011]_  | ~\new_[12014]_  | ~\new_[12006]_  | ~\new_[10397]_ ;
  assign \s0_data_o[27]  = ~\new_[12024]_  | ~\new_[12027]_  | ~\new_[9232]_  | ~\new_[12019]_ ;
  assign \s0_data_o[23]  = ~\new_[12066]_  | ~\new_[12069]_  | ~\new_[9258]_  | ~\new_[12063]_ ;
  assign \s0_data_o[22]  = ~\new_[12077]_  | ~\new_[12075]_  | ~\new_[9264]_  | ~\new_[12072]_ ;
  assign \s0_data_o[21]  = ~\new_[12080]_  | ~\new_[13692]_  | ~\new_[9271]_  | ~\new_[10467]_ ;
  assign \s0_data_o[20]  = ~\new_[12086]_  | ~\new_[13693]_  | ~\new_[9280]_  | ~\new_[12084]_ ;
  assign \s0_addr_o[28]  = ~\new_[12288]_  | ~\new_[13836]_  | ~\new_[9313]_  | ~\new_[12286]_ ;
  assign \s0_addr_o[20]  = ~\new_[12348]_  | ~\new_[12350]_  | ~\new_[12344]_  | ~\new_[10562]_ ;
  assign \s0_addr_o[19]  = ~\new_[13883]_  | ~\new_[12357]_  | ~\new_[10566]_  | ~\new_[10567]_ ;
  assign s7_cyc_o = ~n7554;
  assign \s0_addr_o[14]  = ~\new_[12388]_  | ~\new_[11209]_  | ~\new_[11231]_  | ~\new_[10588]_ ;
  assign \s0_addr_o[12]  = ~\new_[12407]_  | ~\new_[12409]_  | ~\new_[9329]_  | ~\new_[12403]_ ;
  assign \s0_addr_o[11]  = ~\new_[13956]_  | ~\new_[12419]_  | ~\new_[9577]_  | ~\new_[10591]_ ;
  assign \s1_data_o[28]  = ~\new_[14059]_  | ~\new_[14062]_  | ~\new_[15381]_  | ~\new_[10685]_ ;
  assign \s1_data_o[26]  = ~\new_[14072]_  | ~\new_[14540]_  | ~\new_[14069]_  | ~\new_[11081]_ ;
  assign \s1_data_o[25]  = ~\new_[12042]_  | ~\new_[14075]_  | ~\new_[15400]_  | ~\new_[15401]_ ;
  assign \s1_data_o[24]  = ~\new_[13551]_  | ~\new_[12557]_  | ~\new_[14077]_  | ~\new_[15403]_ ;
  assign \s1_data_o[23]  = ~\new_[14083]_  | ~\new_[14084]_  | ~\new_[15406]_  | ~\new_[10700]_ ;
  assign \s1_data_o[22]  = ~\new_[15414]_  | ~\new_[12566]_  | ~\new_[14087]_  | ~\new_[15413]_ ;
  assign \s1_data_o[21]  = ~\new_[12607]_  | ~\new_[14092]_  | ~\new_[15419]_  | ~\new_[15420]_ ;
  assign \s1_data_o[20]  = ~\new_[15428]_  | ~\new_[14097]_  | ~\new_[14486]_  | ~\new_[10707]_ ;
  assign \s1_data_o[19]  = ~\new_[15435]_  | ~\new_[12941]_  | ~\new_[14197]_  | ~\new_[15432]_ ;
  assign \s1_data_o[16]  = ~\new_[13497]_  | ~\new_[14106]_  | ~\new_[15453]_  | ~\new_[10719]_ ;
  assign \s1_data_o[14]  = ~\new_[12595]_  | ~\new_[14111]_  | ~\new_[14110]_  | ~\new_[15459]_ ;
  assign \s1_data_o[12]  = ~\new_[14118]_  | ~\new_[12605]_  | ~\new_[15464]_  | ~\new_[15465]_ ;
  assign \s1_data_o[11]  = ~\new_[11707]_  | ~\new_[15468]_  | ~\new_[14119]_  | ~\new_[14120]_ ;
  assign \s1_data_o[10]  = ~\new_[12610]_  | ~\new_[13623]_  | ~\new_[14380]_  | ~\new_[15469]_ ;
  assign \s1_data_o[9]  = ~\new_[12979]_  | ~\new_[14125]_  | ~\new_[15470]_  | ~\new_[14123]_ ;
  assign \s1_data_o[8]  = ~\new_[12618]_  | ~\new_[15473]_  | ~\new_[15472]_  | ~\new_[14127]_ ;
  assign \s1_data_o[7]  = ~\new_[12621]_  | ~\new_[15477]_  | ~\new_[14129]_  | ~\new_[14130]_ ;
  assign \s1_data_o[5]  = ~\new_[12637]_  | ~\new_[14143]_  | ~\new_[15482]_  | ~\new_[15483]_ ;
  assign \s1_data_o[2]  = ~\new_[12667]_  | ~\new_[15491]_  | ~\new_[15489]_  | ~\new_[14155]_ ;
  assign \s1_addr_o[31]  = ~\new_[12682]_  | ~\new_[14173]_  | ~\new_[14168]_  | ~\new_[15504]_ ;
  assign \s1_addr_o[29]  = ~\new_[15515]_  | ~\new_[12696]_  | ~\new_[15512]_  | ~\new_[15514]_ ;
  assign \s1_addr_o[24]  = ~\new_[12728]_  | ~\new_[14211]_  | ~\new_[15535]_  | ~\new_[14207]_ ;
  assign \s1_addr_o[23]  = ~\new_[14214]_  | ~\new_[15546]_  | ~\new_[15538]_  | ~\new_[10814]_ ;
  assign \s1_addr_o[21]  = ~\new_[15551]_  | ~\new_[14225]_  | ~\new_[15550]_  | ~\new_[10827]_ ;
  assign \s1_addr_o[19]  = ~\new_[15558]_  | ~\new_[12761]_  | ~\new_[14232]_  | ~\new_[15557]_ ;
  assign \s1_addr_o[18]  = ~\new_[15566]_  | ~\new_[12767]_  | ~\new_[14236]_  | ~\new_[15563]_ ;
  assign \s1_addr_o[17]  = ~\new_[12771]_  | ~\new_[14244]_  | ~\new_[15568]_  | ~\new_[15569]_ ;
  assign \s1_addr_o[16]  = ~\new_[14247]_  | ~\new_[12776]_  | ~\new_[15574]_  | ~\new_[14245]_ ;
  assign \s1_addr_o[15]  = ~\new_[15580]_  | ~\new_[12781]_  | ~\new_[14251]_  | ~\new_[15579]_ ;
  assign \s1_addr_o[14]  = ~\new_[15586]_  | ~\new_[12787]_  | ~\new_[14254]_  | ~\new_[15584]_ ;
  assign \s1_addr_o[13]  = ~\new_[15592]_  | ~\new_[12793]_  | ~\new_[15589]_  | ~\new_[14261]_ ;
  assign \s1_addr_o[11]  = ~\new_[14270]_  | ~\new_[12806]_  | ~\new_[15600]_  | ~\new_[15601]_ ;
  assign \s1_addr_o[10]  = ~\new_[15608]_  | ~\new_[12813]_  | ~\new_[14273]_  | ~\new_[15606]_ ;
  assign \s1_addr_o[9]  = ~\new_[15614]_  | ~\new_[12817]_  | ~\new_[14277]_  | ~\new_[14280]_ ;
  assign \s1_addr_o[8]  = ~\new_[15616]_  | ~\new_[12822]_  | ~\new_[14290]_  | ~\new_[14285]_ ;
  assign \s1_addr_o[7]  = ~\new_[15620]_  | ~\new_[12825]_  | ~\new_[14291]_  | ~\new_[15619]_ ;
  assign \s1_addr_o[6]  = ~\new_[15623]_  | ~\new_[12827]_  | ~\new_[14295]_  | ~\new_[14296]_ ;
  assign \s1_addr_o[5]  = ~\new_[15629]_  | ~\new_[12829]_  | ~\new_[14297]_  | ~\new_[14298]_ ;
  assign \s1_addr_o[4]  = ~\new_[15631]_  | ~\new_[12835]_  | ~\new_[14304]_  | ~\new_[14305]_ ;
  assign \s1_addr_o[3]  = ~\new_[15635]_  | ~\new_[12839]_  | ~\new_[14311]_  | ~\new_[14312]_ ;
  assign \s1_addr_o[2]  = ~\new_[15637]_  | ~\new_[12844]_  | ~\new_[14317]_  | ~\new_[14319]_ ;
  assign \s1_addr_o[1]  = ~\new_[15645]_  | ~\new_[12846]_  | ~\new_[14323]_  | ~\new_[15643]_ ;
  assign \s1_addr_o[0]  = ~\new_[15652]_  | ~\new_[12851]_  | ~\new_[14326]_  | ~\new_[15649]_ ;
  assign \s1_sel_o[3]  = ~\new_[15654]_  | ~\new_[12855]_  | ~\new_[14328]_  | ~\new_[15653]_ ;
  assign \s1_sel_o[1]  = ~\new_[15658]_  | ~\new_[12860]_  | ~\new_[15656]_  | ~\new_[15657]_ ;
  assign \s1_sel_o[0]  = ~\new_[15660]_  | ~\new_[12867]_  | ~\new_[14331]_  | ~\new_[15659]_ ;
  assign s1_we_o = ~\new_[15663]_  | ~\new_[12873]_  | ~\new_[14332]_  | ~\new_[14334]_ ;
  assign \s2_data_o[29]  = ~\new_[12903]_  | ~\new_[14341]_  | ~\new_[10986]_  | ~\new_[14340]_ ;
  assign \s2_data_o[27]  = ~\new_[12911]_  | ~\new_[14344]_  | ~\new_[15672]_  | ~\new_[14343]_ ;
  assign \s2_data_o[25]  = ~\new_[12919]_  | ~\new_[15684]_  | ~\new_[12916]_  | ~\new_[11016]_ ;
  assign \s2_data_o[24]  = ~\new_[12923]_  | ~\new_[15688]_  | ~\new_[12921]_  | ~\new_[11022]_ ;
  assign \s2_data_o[23]  = ~\new_[12926]_  | ~\new_[14354]_  | ~\new_[12925]_  | ~\new_[11026]_ ;
  assign \s2_data_o[22]  = ~\new_[12930]_  | ~\new_[14355]_  | ~\new_[12929]_  | ~\new_[11031]_ ;
  assign \s2_data_o[21]  = ~\new_[12934]_  | ~\new_[14361]_  | ~\new_[12933]_  | ~\new_[11038]_ ;
  assign \s2_data_o[20]  = ~\new_[12938]_  | ~\new_[15706]_  | ~\new_[14362]_  | ~\new_[11042]_ ;
  assign \s2_data_o[19]  = ~\new_[15710]_  | ~\new_[14368]_  | ~\new_[14367]_  | ~\new_[11045]_ ;
  assign \s2_data_o[18]  = ~\new_[15713]_  | ~\new_[15714]_  | ~\new_[12944]_  | ~\new_[11050]_ ;
  assign \s2_data_o[17]  = ~\new_[12951]_  | ~\new_[15716]_  | ~\new_[12949]_  | ~\new_[11053]_ ;
  assign \s2_data_o[16]  = ~\new_[12956]_  | ~\new_[14372]_  | ~\new_[12953]_  | ~\new_[11059]_ ;
  assign \s2_data_o[15]  = ~\new_[12960]_  | ~\new_[14378]_  | ~\new_[12959]_  | ~\new_[11063]_ ;
  assign \s2_data_o[14]  = ~\new_[12966]_  | ~\new_[14381]_  | ~\new_[12963]_  | ~\new_[11070]_ ;
  assign \s2_data_o[13]  = ~\new_[12969]_  | ~\new_[15729]_  | ~\new_[12968]_  | ~\new_[11075]_ ;
  assign \s2_data_o[12]  = ~\new_[12974]_  | ~\new_[15733]_  | ~\new_[12971]_  | ~\new_[12973]_ ;
  assign \s2_data_o[11]  = ~\new_[12976]_  | ~\new_[15735]_  | ~\new_[12975]_  | ~\new_[11078]_ ;
  assign \s2_data_o[10]  = ~\new_[12978]_  | ~\new_[15738]_  | ~\new_[12977]_  | ~\new_[11080]_ ;
  assign \s2_data_o[9]  = ~\new_[12982]_  | ~\new_[14392]_  | ~\new_[12980]_  | ~\new_[12981]_ ;
  assign \s2_data_o[8]  = ~\new_[12986]_  | ~\new_[14393]_  | ~\new_[12983]_  | ~\new_[12985]_ ;
  assign \s2_data_o[7]  = ~\new_[12989]_  | ~\new_[14395]_  | ~\new_[12987]_  | ~\new_[12988]_ ;
  assign \s2_data_o[6]  = ~\new_[12992]_  | ~\new_[15750]_  | ~\new_[12990]_  | ~\new_[12991]_ ;
  assign \s2_data_o[5]  = ~\new_[12995]_  | ~\new_[14397]_  | ~\new_[12993]_  | ~\new_[12994]_ ;
  assign \s2_data_o[4]  = ~\new_[12998]_  | ~\new_[15756]_  | ~\new_[12996]_  | ~\new_[12997]_ ;
  assign \s2_data_o[3]  = ~\new_[13000]_  | ~\new_[14403]_  | ~\new_[12999]_  | ~\new_[11086]_ ;
  assign \s2_data_o[2]  = ~\new_[13003]_  | ~\new_[14406]_  | ~\new_[13001]_  | ~\new_[13002]_ ;
  assign \s2_data_o[1]  = ~\new_[13005]_  | ~\new_[15765]_  | ~\new_[13004]_  | ~\new_[11090]_ ;
  assign \s2_data_o[0]  = ~\new_[13008]_  | ~\new_[14410]_  | ~\new_[13007]_  | ~\new_[11091]_ ;
  assign \s2_addr_o[31]  = ~\new_[13010]_  | ~\new_[14412]_  | ~\new_[13009]_  | ~\new_[11092]_ ;
  assign \s2_addr_o[30]  = ~\new_[13013]_  | ~\new_[14415]_  | ~\new_[13012]_  | ~\new_[11093]_ ;
  assign \s2_addr_o[29]  = ~\new_[13015]_  | ~\new_[14419]_  | ~\new_[13014]_  | ~\new_[11094]_ ;
  assign \s2_addr_o[28]  = ~\new_[15781]_  | ~\new_[14422]_  | ~\new_[13017]_  | ~\new_[11096]_ ;
  assign \s2_addr_o[27]  = ~\new_[15786]_  | ~\new_[14425]_  | ~\new_[13018]_  | ~\new_[11098]_ ;
  assign \s2_addr_o[26]  = ~\new_[15790]_  | ~\new_[14430]_  | ~\new_[13019]_  | ~\new_[11099]_ ;
  assign \s2_addr_o[25]  = ~\new_[15795]_  | ~\new_[14431]_  | ~\new_[13022]_  | ~\new_[11102]_ ;
  assign \s2_addr_o[24]  = ~\new_[13027]_  | ~\new_[14433]_  | ~\new_[13024]_  | ~\new_[11105]_ ;
  assign n7494 = ~\new_[9273]_  & ~\new_[9274]_ ;
  assign \s2_addr_o[23]  = ~\new_[13030]_  | ~\new_[15805]_  | ~\new_[13028]_  | ~\new_[11108]_ ;
  assign \s2_addr_o[22]  = ~\new_[13032]_  | ~\new_[15807]_  | ~\new_[13031]_  | ~\new_[11109]_ ;
  assign \s2_addr_o[21]  = ~\new_[13035]_  | ~\new_[14440]_  | ~\new_[13034]_  | ~\new_[11110]_ ;
  assign \s2_addr_o[20]  = ~\new_[15816]_  | ~\new_[15819]_  | ~\new_[13037]_  | ~\new_[11111]_ ;
  assign \s2_addr_o[19]  = ~\new_[15826]_  | ~\new_[15829]_  | ~\new_[13039]_  | ~\new_[11114]_ ;
  assign \s2_addr_o[18]  = ~\new_[15835]_  | ~\new_[14447]_  | ~\new_[13040]_  | ~\new_[11115]_ ;
  assign \s2_addr_o[17]  = ~\new_[13042]_  | ~\new_[14450]_  | ~\new_[13041]_  | ~\new_[11116]_ ;
  assign \s2_addr_o[16]  = ~\new_[13044]_  | ~\new_[15856]_  | ~\new_[14451]_  | ~\new_[11117]_ ;
  assign \s2_addr_o[15]  = ~\new_[13045]_  | ~\new_[15857]_  | ~\new_[14454]_  | ~\new_[11118]_ ;
  assign \s2_addr_o[14]  = ~\new_[13046]_  | ~\new_[15858]_  | ~\new_[14458]_  | ~\new_[11119]_ ;
  assign \s2_addr_o[13]  = ~\new_[13050]_  | ~\new_[14463]_  | ~\new_[13047]_  | ~\new_[11120]_ ;
  assign \s2_addr_o[12]  = ~\new_[13052]_  | ~\new_[14465]_  | ~\new_[13051]_  | ~\new_[11123]_ ;
  assign \s2_addr_o[11]  = ~\new_[15863]_  | ~\new_[14467]_  | ~\new_[14466]_  | ~\new_[11124]_ ;
  assign \s2_addr_o[10]  = ~\new_[15865]_  | ~\new_[14470]_  | ~\new_[13055]_  | ~\new_[11126]_ ;
  assign \s2_addr_o[9]  = ~\new_[13057]_  | ~\new_[15868]_  | ~\new_[14471]_  | ~\new_[11127]_ ;
  assign \s2_addr_o[8]  = ~\new_[13059]_  | ~\new_[14472]_  | ~\new_[13058]_  | ~\new_[11128]_ ;
  assign \s2_addr_o[7]  = ~\new_[15869]_  | ~\new_[15870]_  | ~\new_[13060]_  | ~\new_[11129]_ ;
  assign \s2_addr_o[6]  = ~\new_[13061]_  | ~\new_[14474]_  | ~\new_[14473]_  | ~\new_[11131]_ ;
  assign \s2_addr_o[5]  = ~\new_[13064]_  | ~\new_[15872]_  | ~\new_[13062]_  | ~\new_[13063]_ ;
  assign \s2_addr_o[4]  = ~\new_[13067]_  | ~\new_[14476]_  | ~\new_[13065]_  | ~\new_[13066]_ ;
  assign \s2_addr_o[3]  = ~\new_[13069]_  | ~\new_[15875]_  | ~\new_[13068]_  | ~\new_[11133]_ ;
  assign \s2_addr_o[2]  = ~\new_[13072]_  | ~\new_[14479]_  | ~\new_[13070]_  | ~\new_[13071]_ ;
  assign \s2_addr_o[1]  = ~\new_[13074]_  | ~\new_[15876]_  | ~\new_[13073]_  | ~\new_[11134]_ ;
  assign \s2_addr_o[0]  = ~\new_[13077]_  | ~\new_[14480]_  | ~\new_[13076]_  | ~\new_[11135]_ ;
  assign \s2_sel_o[3]  = ~\new_[13079]_  | ~\new_[15879]_  | ~\new_[13078]_  | ~\new_[11136]_ ;
  assign \s2_sel_o[2]  = ~\new_[13082]_  | ~\new_[15882]_  | ~\new_[13080]_  | ~\new_[11137]_ ;
  assign \s2_sel_o[1]  = ~\new_[13084]_  | ~\new_[14482]_  | ~\new_[13083]_  | ~\new_[11139]_ ;
  assign \s2_sel_o[0]  = ~\new_[13086]_  | ~\new_[14484]_  | ~\new_[13085]_  | ~\new_[11140]_ ;
  assign s2_we_o = ~\new_[13090]_  | ~\new_[14485]_  | ~\new_[13088]_  | ~\new_[13089]_ ;
  assign \s3_data_o[31]  = ~\new_[14487]_  | ~\new_[15885]_  | ~\new_[13092]_  | ~\new_[11142]_ ;
  assign \s3_data_o[28]  = ~\new_[14492]_  | ~\new_[14493]_  | ~\new_[13096]_  | ~\new_[11149]_ ;
  assign \s3_data_o[27]  = ~\new_[13098]_  | ~\new_[14494]_  | ~\new_[13097]_  | ~\new_[11150]_ ;
  assign \s3_data_o[26]  = ~\new_[14495]_  | ~\new_[15888]_  | ~\new_[13099]_  | ~\new_[11151]_ ;
  assign \s3_data_o[25]  = ~\new_[14497]_  | ~\new_[14498]_  | ~\new_[14496]_  | ~\new_[11152]_ ;
  assign \s3_data_o[24]  = ~\new_[14499]_  | ~\new_[15890]_  | ~\new_[13100]_  | ~\new_[11153]_ ;
  assign \s3_data_o[23]  = ~\new_[14500]_  | ~\new_[14501]_  | ~\new_[13102]_  | ~\new_[11156]_ ;
  assign \s3_data_o[22]  = ~\new_[14502]_  | ~\new_[13104]_  | ~\new_[13103]_  | ~\new_[11157]_ ;
  assign \s3_data_o[21]  = ~\new_[13105]_  | ~\new_[13106]_  | ~\new_[11158]_  | ~\new_[9574]_ ;
  assign \s3_data_o[20]  = ~\new_[11160]_  | ~\new_[13107]_  | ~\new_[11159]_  | ~\new_[9576]_ ;
  assign \s3_data_o[19]  = ~\new_[13108]_  | ~\new_[14508]_  | ~\new_[11161]_  | ~\new_[9578]_ ;
  assign \s3_data_o[18]  = ~\new_[13110]_  | ~\new_[13111]_  | ~\new_[13109]_  | ~\new_[9579]_ ;
  assign \s3_data_o[16]  = ~\new_[13116]_  | ~\new_[13117]_  | ~\new_[11165]_  | ~\new_[9582]_ ;
  assign \s3_data_o[11]  = ~\new_[13126]_  | ~\new_[13127]_  | ~\new_[11167]_  | ~\new_[9592]_ ;
  assign \new_[7595]_  = ~\new_[12028]_  & (~\new_[10820]_  | ~\new_[27776]_ );
  assign \s3_addr_o[31]  = ~\new_[11178]_  | ~\new_[13150]_  | ~\new_[13148]_  | ~\new_[11177]_ ;
  assign \s3_addr_o[30]  = ~\new_[11180]_  | ~\new_[13152]_  | ~\new_[13151]_  | ~\new_[11179]_ ;
  assign \s3_addr_o[29]  = ~\new_[11182]_  | ~\new_[13155]_  | ~\new_[13153]_  | ~\new_[11181]_ ;
  assign \new_[7599]_  = ~\new_[12815]_  & ~\new_[9137]_ ;
  assign \s3_addr_o[23]  = ~\new_[13168]_  | ~\new_[13169]_  | ~\new_[11192]_  | ~\new_[10554]_ ;
  assign \s3_addr_o[22]  = ~\new_[13796]_  | ~\new_[13171]_  | ~\new_[11198]_  | ~\new_[9627]_ ;
  assign \s3_addr_o[21]  = ~\new_[13172]_  | ~\new_[13760]_  | ~\new_[11200]_  | ~\new_[9630]_ ;
  assign \new_[7603]_  = ~\new_[9369]_  & ~\new_[9219]_ ;
  assign \s3_addr_o[20]  = ~\new_[13724]_  | ~\new_[13718]_  | ~\new_[11203]_  | ~\new_[9633]_ ;
  assign \s3_addr_o[19]  = ~\new_[13176]_  | ~\new_[13177]_  | ~\new_[11204]_  | ~\new_[9634]_ ;
  assign \s3_addr_o[18]  = ~\new_[13179]_  | ~\new_[13180]_  | ~\new_[11205]_  | ~\new_[9635]_ ;
  assign \s3_addr_o[17]  = ~\new_[13181]_  | ~\new_[13182]_  | ~\new_[11901]_  | ~\new_[9637]_ ;
  assign \s3_addr_o[16]  = ~\new_[13183]_  | ~\new_[13444]_  | ~\new_[11207]_  | ~\new_[9639]_ ;
  assign \s3_addr_o[13]  = ~\new_[13187]_  | ~\new_[13188]_  | ~\new_[11216]_  | ~\new_[9645]_ ;
  assign \s3_addr_o[12]  = ~\new_[13191]_  | ~\new_[13192]_  | ~\new_[11219]_  | ~\new_[9646]_ ;
  assign \s3_addr_o[11]  = ~\new_[13194]_  | ~\new_[14544]_  | ~\new_[11222]_  | ~\new_[9648]_ ;
  assign \s3_addr_o[9]  = ~\new_[13199]_  | ~\new_[13200]_  | ~\new_[11227]_  | ~\new_[9652]_ ;
  assign \s3_addr_o[10]  = ~\new_[13196]_  | ~\new_[14918]_  | ~\new_[11223]_  | ~\new_[9651]_ ;
  assign \s3_addr_o[7]  = ~\new_[13133]_  | ~\new_[14448]_  | ~\new_[11235]_  | ~\new_[9623]_ ;
  assign \s3_addr_o[6]  = ~\new_[12802]_  | ~\new_[14137]_  | ~\new_[12888]_  | ~\new_[10926]_ ;
  assign \s3_addr_o[1]  = ~\new_[13204]_  | ~\new_[13149]_  | ~\new_[13490]_  | ~\new_[9660]_ ;
  assign \s3_sel_o[2]  = ~\new_[13601]_  | ~\new_[13592]_  | ~\new_[11923]_  | ~\new_[10180]_ ;
  assign \s3_sel_o[3]  = ~\new_[13682]_  | ~\new_[13759]_  | ~\new_[12512]_  | ~\new_[9661]_ ;
  assign \s3_sel_o[0]  = ~\new_[13528]_  | ~\new_[14869]_  | ~\new_[11763]_  | ~\new_[9662]_ ;
  assign \s4_data_o[29]  = ~\new_[14902]_  | ~\new_[11238]_  | ~\new_[11825]_  | ~\new_[11842]_ ;
  assign \s4_data_o[27]  = ~\new_[14551]_  | ~\new_[11240]_  | ~\new_[11239]_  | ~\new_[11218]_ ;
  assign \s4_data_o[26]  = ~\new_[15133]_  | ~\new_[11241]_  | ~\new_[11196]_  | ~\new_[12416]_ ;
  assign \s4_data_o[25]  = ~\new_[15542]_  | ~\new_[11243]_  | ~\new_[12957]_  | ~\new_[12853]_ ;
  assign \s4_data_o[21]  = ~\new_[14894]_  | ~\new_[11696]_  | ~\new_[11761]_  | ~\new_[11189]_ ;
  assign \s4_data_o[20]  = ~\new_[14545]_  | ~\new_[11220]_  | ~\new_[11230]_  | ~\new_[11224]_ ;
  assign \s4_data_o[17]  = ~\new_[14835]_  | ~\new_[11847]_  | ~\new_[11193]_  | ~\new_[11556]_ ;
  assign \s4_data_o[16]  = ~\new_[14827]_  | ~\new_[11657]_  | ~\new_[11796]_  | ~\new_[11675]_ ;
  assign \s4_data_o[15]  = ~\new_[14710]_  | ~\new_[11245]_  | ~\new_[11208]_  | ~\new_[11425]_ ;
  assign \s4_data_o[14]  = ~\new_[14655]_  | ~\new_[13049]_  | ~\new_[12431]_  | ~\new_[11881]_ ;
  assign \s4_data_o[9]  = ~\new_[15259]_  | ~\new_[12134]_  | ~\new_[12777]_  | ~\new_[15517]_ ;
  assign \s4_data_o[6]  = ~\new_[15801]_  | ~\new_[12757]_  | ~\new_[11287]_  | ~\new_[14552]_ ;
  assign \s4_data_o[5]  = ~\new_[14914]_  | ~\new_[11518]_  | ~\new_[12459]_  | ~\new_[14963]_ ;
  assign \s4_data_o[3]  = ~\new_[14889]_  | ~\new_[11480]_  | ~\new_[12287]_  | ~\new_[14923]_ ;
  assign \s4_data_o[2]  = ~\new_[15560]_  | ~\new_[12139]_  | ~\new_[11391]_  | ~\new_[15778]_ ;
  assign \s4_data_o[0]  = ~\new_[14959]_  | ~\new_[11401]_  | ~\new_[11214]_  | ~\new_[15344]_ ;
  assign \s4_addr_o[31]  = ~\new_[14533]_  | ~\new_[11252]_  | ~\new_[11232]_  | ~\new_[14901]_ ;
  assign \s4_addr_o[30]  = ~\new_[14535]_  | ~\new_[11253]_  | ~\new_[11234]_  | ~\new_[14548]_ ;
  assign \s4_addr_o[29]  = ~\new_[14554]_  | ~\new_[11257]_  | ~\new_[11255]_  | ~\new_[14553]_ ;
  assign \s4_addr_o[28]  = ~\new_[14556]_  | ~\new_[11260]_  | ~\new_[11258]_  | ~\new_[14555]_ ;
  assign \s4_addr_o[27]  = ~\new_[14558]_  | ~\new_[11264]_  | ~\new_[11262]_  | ~\new_[14557]_ ;
  assign \s4_addr_o[25]  = ~\new_[14534]_  | ~\new_[11201]_  | ~\new_[11748]_  | ~\new_[14872]_ ;
  assign \s4_addr_o[24]  = ~\new_[16518]_  | ~\new_[11242]_  | ~\new_[11191]_  | ~\new_[15836]_ ;
  assign \s4_addr_o[26]  = ~\new_[14561]_  | ~\new_[11267]_  | ~\new_[11265]_  | ~\new_[14560]_ ;
  assign \s4_addr_o[23]  = ~\new_[14520]_  | ~\new_[11202]_  | ~\new_[11183]_  | ~\new_[11810]_ ;
  assign \s4_addr_o[21]  = ~\new_[14538]_  | ~\new_[11206]_  | ~\new_[11221]_  | ~\new_[11226]_ ;
  assign \new_[7646]_  = ~\new_[12031]_  & (~\new_[10822]_  | ~\new_[24480]_ );
  assign \s4_addr_o[18]  = ~\new_[15056]_  | ~\new_[11322]_  | ~\new_[13023]_  | ~\new_[12706]_ ;
  assign \s4_addr_o[16]  = ~\new_[14962]_  | ~\new_[11250]_  | ~\new_[13020]_  | ~\new_[12575]_ ;
  assign \s4_addr_o[15]  = ~\new_[14897]_  | ~\new_[11394]_  | ~\new_[12906]_  | ~\new_[12473]_ ;
  assign \s4_addr_o[13]  = ~\new_[16033]_  | ~\new_[12939]_  | ~\new_[12232]_  | ~\new_[11585]_ ;
  assign \s4_addr_o[10]  = ~\new_[15939]_  | ~\new_[11259]_  | ~\new_[11254]_  | ~\new_[11256]_ ;
  assign \s4_addr_o[7]  = ~\new_[14564]_  | ~\new_[11271]_  | ~\new_[11269]_  | ~\new_[11270]_ ;
  assign \new_[7653]_  = ~\new_[12820]_  & ~\new_[9143]_ ;
  assign \s4_addr_o[5]  = ~\new_[14571]_  | ~\new_[11277]_  | ~\new_[11275]_  | ~\new_[11276]_ ;
  assign \s4_sel_o[3]  = ~\new_[14583]_  | ~\new_[11290]_  | ~\new_[11288]_  | ~\new_[11289]_ ;
  assign \new_[7656]_  = ~\new_[9370]_  & ~\new_[9220]_ ;
  assign \s4_sel_o[1]  = ~\new_[15987]_  | ~\new_[11295]_  | ~\new_[11294]_  | ~\new_[11293]_ ;
  assign \s4_sel_o[0]  = ~\new_[14590]_  | ~\new_[11298]_  | ~\new_[11296]_  | ~\new_[11297]_ ;
  assign s4_we_o = ~\new_[14598]_  | ~\new_[11301]_  | ~\new_[11299]_  | ~\new_[14597]_ ;
  assign \s5_data_o[31]  = ~\new_[13219]_  | ~\new_[11304]_  | ~\new_[11303]_  | ~\new_[14599]_ ;
  assign \s5_data_o[29]  = ~\new_[13222]_  | ~\new_[11307]_  | ~\new_[11306]_  | ~\new_[14601]_ ;
  assign \s5_data_o[28]  = ~\new_[13223]_  | ~\new_[11311]_  | ~\new_[11310]_  | ~\new_[14602]_ ;
  assign \s5_data_o[27]  = ~\new_[13224]_  | ~\new_[11313]_  | ~\new_[11312]_  | ~\new_[14603]_ ;
  assign \s5_data_o[26]  = ~\new_[13225]_  | ~\new_[11317]_  | ~\new_[11315]_  | ~\new_[14605]_ ;
  assign \s5_data_o[25]  = ~\new_[13228]_  | ~\new_[11319]_  | ~\new_[11318]_  | ~\new_[14606]_ ;
  assign \s5_data_o[24]  = ~\new_[13229]_  | ~\new_[11321]_  | ~\new_[11320]_  | ~\new_[14607]_ ;
  assign \s5_data_o[22]  = ~\new_[13233]_  | ~\new_[11325]_  | ~\new_[11323]_  | ~\new_[14610]_ ;
  assign \s5_data_o[19]  = ~\new_[13239]_  | ~\new_[11330]_  | ~\new_[11329]_  | ~\new_[14617]_ ;
  assign \s5_data_o[17]  = ~\new_[13243]_  | ~\new_[11334]_  | ~\new_[11333]_  | ~\new_[14621]_ ;
  assign \s5_data_o[16]  = ~\new_[13244]_  | ~\new_[11336]_  | ~\new_[11335]_  | ~\new_[14623]_ ;
  assign \s5_data_o[15]  = ~\new_[13246]_  | ~\new_[11338]_  | ~\new_[11337]_  | ~\new_[14626]_ ;
  assign \s5_data_o[14]  = ~\new_[13248]_  | ~\new_[11341]_  | ~\new_[11339]_  | ~\new_[14630]_ ;
  assign \s5_data_o[13]  = ~\new_[13251]_  | ~\new_[11343]_  | ~\new_[11342]_  | ~\new_[14635]_ ;
  assign n7489 = ~\new_[9279]_  & ~\new_[9281]_ ;
  assign \s5_data_o[12]  = ~\new_[13253]_  | ~\new_[11346]_  | ~\new_[14639]_  | ~\new_[14640]_ ;
  assign \s5_data_o[11]  = ~\new_[13255]_  | ~\new_[11347]_  | ~\new_[14642]_  | ~\new_[14644]_ ;
  assign \s5_data_o[10]  = ~\new_[13259]_  | ~\new_[11348]_  | ~\new_[14647]_  | ~\new_[14648]_ ;
  assign \s5_data_o[9]  = ~\new_[13262]_  | ~\new_[11350]_  | ~\new_[11349]_  | ~\new_[14651]_ ;
  assign \s5_data_o[8]  = ~\new_[13263]_  | ~\new_[11352]_  | ~\new_[11351]_  | ~\new_[14654]_ ;
  assign \s5_data_o[7]  = ~\new_[13264]_  | ~\new_[11355]_  | ~\new_[14656]_  | ~\new_[14658]_ ;
  assign \s5_data_o[6]  = ~\new_[13266]_  | ~\new_[11357]_  | ~\new_[11356]_  | ~\new_[14660]_ ;
  assign \s5_data_o[5]  = ~\new_[13268]_  | ~\new_[11360]_  | ~\new_[11359]_  | ~\new_[14662]_ ;
  assign \s5_data_o[1]  = ~\new_[14667]_  | ~\new_[11365]_  | ~\new_[13278]_  | ~\new_[13279]_ ;
  assign \s5_addr_o[23]  = ~\new_[13303]_  | ~\new_[11370]_  | ~\new_[11368]_  | ~\new_[14698]_ ;
  assign \s5_addr_o[22]  = ~\new_[14700]_  | ~\new_[11371]_  | ~\new_[13304]_  | ~\new_[14699]_ ;
  assign \s5_addr_o[21]  = ~\new_[13305]_  | ~\new_[11375]_  | ~\new_[11373]_  | ~\new_[14702]_ ;
  assign \s5_addr_o[18]  = ~\new_[13318]_  | ~\new_[11382]_  | ~\new_[11380]_  | ~\new_[14712]_ ;
  assign \s5_addr_o[11]  = ~\new_[13336]_  | ~\new_[11392]_  | ~\new_[11389]_  | ~\new_[14735]_ ;
  assign \s5_addr_o[10]  = ~\new_[13338]_  | ~\new_[11395]_  | ~\new_[11393]_  | ~\new_[14736]_ ;
  assign \s5_addr_o[1]  = ~\new_[13370]_  | ~\new_[11410]_  | ~\new_[11407]_  | ~\new_[14763]_ ;
  assign \s5_addr_o[0]  = ~\new_[13373]_  | ~\new_[11412]_  | ~\new_[14765]_  | ~\new_[14766]_ ;
  assign \s5_sel_o[3]  = ~\new_[13378]_  | ~\new_[11413]_  | ~\new_[13376]_  | ~\new_[14771]_ ;
  assign \s6_data_o[31]  = ~\new_[11422]_  | ~\new_[11423]_  | ~\new_[13391]_  | ~\new_[13392]_ ;
  assign s5_stb_o = \new_[12856]_  | \new_[9415]_ ;
  assign \s6_data_o[29]  = ~\new_[11428]_  | ~\new_[11429]_  | ~\new_[11426]_  | ~\new_[11427]_ ;
  assign \s6_data_o[28]  = ~\new_[14798]_  | ~\new_[11431]_  | ~\new_[13397]_  | ~\new_[13398]_ ;
  assign \s6_data_o[27]  = ~\new_[11433]_  | ~\new_[13402]_  | ~\new_[11432]_  | ~\new_[9784]_ ;
  assign \s6_data_o[26]  = ~\new_[13403]_  | ~\new_[13405]_  | ~\new_[11434]_  | ~\new_[9786]_ ;
  assign \new_[7699]_  = ~\new_[12033]_  & (~\new_[10826]_  | ~\new_[23101]_ );
  assign \s6_data_o[23]  = ~\new_[11443]_  | ~\new_[11444]_  | ~\new_[11442]_  | ~\new_[13412]_ ;
  assign \s6_data_o[18]  = ~\new_[11458]_  | ~\new_[11459]_  | ~\new_[11456]_  | ~\new_[11457]_ ;
  assign \s6_data_o[17]  = ~\new_[13419]_  | ~\new_[13420]_  | ~\new_[11460]_  | ~\new_[9807]_ ;
  assign \s6_data_o[16]  = ~\new_[13421]_  | ~\new_[11462]_  | ~\new_[11461]_  | ~\new_[9809]_ ;
  assign \s6_data_o[15]  = ~\new_[11465]_  | ~\new_[11466]_  | ~\new_[11463]_  | ~\new_[9811]_ ;
  assign \s6_data_o[14]  = ~\new_[11468]_  | ~\new_[11469]_  | ~\new_[11467]_  | ~\new_[9812]_ ;
  assign \s6_data_o[13]  = ~\new_[11471]_  | ~\new_[11472]_  | ~\new_[11470]_  | ~\new_[13422]_ ;
  assign \s6_data_o[12]  = ~\new_[11474]_  | ~\new_[13423]_  | ~\new_[11473]_  | ~\new_[9814]_ ;
  assign \s6_data_o[11]  = ~\new_[11477]_  | ~\new_[13425]_  | ~\new_[11476]_  | ~\new_[11475]_ ;
  assign \s6_data_o[10]  = ~\new_[11478]_  | ~\new_[13429]_  | ~\new_[13426]_  | ~\new_[13427]_ ;
  assign \s6_data_o[9]  = ~\new_[14817]_  | ~\new_[11481]_  | ~\new_[13430]_  | ~\new_[13431]_ ;
  assign \s6_data_o[8]  = ~\new_[14820]_  | ~\new_[11482]_  | ~\new_[13432]_  | ~\new_[13433]_ ;
  assign \s6_data_o[7]  = ~\new_[11486]_  | ~\new_[11487]_  | ~\new_[11484]_  | ~\new_[11485]_ ;
  assign \s6_data_o[6]  = ~\new_[11489]_  | ~\new_[11490]_  | ~\new_[13435]_  | ~\new_[13436]_ ;
  assign \s6_data_o[5]  = ~\new_[11492]_  | ~\new_[11493]_  | ~\new_[13438]_  | ~\new_[13439]_ ;
  assign \new_[7715]_  = ~\new_[9372]_  & ~\new_[9221]_ ;
  assign \s6_data_o[4]  = ~\new_[11496]_  | ~\new_[11494]_  | ~\new_[13440]_  | ~\new_[9830]_ ;
  assign \s6_data_o[3]  = ~\new_[14824]_  | ~\new_[11498]_  | ~\new_[13443]_  | ~\new_[13442]_ ;
  assign \s6_data_o[2]  = ~\new_[11500]_  | ~\new_[11501]_  | ~\new_[13445]_  | ~\new_[13446]_ ;
  assign \s6_data_o[1]  = ~\new_[14826]_  | ~\new_[11504]_  | ~\new_[13447]_  | ~\new_[13448]_ ;
  assign \s6_data_o[0]  = ~\new_[11506]_  | ~\new_[11507]_  | ~\new_[11505]_  | ~\new_[9839]_ ;
  assign \s6_addr_o[31]  = ~\new_[11508]_  | ~\new_[13451]_  | ~\new_[13449]_  | ~\new_[13450]_ ;
  assign \s6_addr_o[30]  = ~\new_[11510]_  | ~\new_[11511]_  | ~\new_[11509]_  | ~\new_[13452]_ ;
  assign \s6_addr_o[29]  = ~\new_[11513]_  | ~\new_[14828]_  | ~\new_[11512]_  | ~\new_[13453]_ ;
  assign \s6_addr_o[28]  = ~\new_[11517]_  | ~\new_[11519]_  | ~\new_[11514]_  | ~\new_[13454]_ ;
  assign \s6_addr_o[27]  = ~\new_[11522]_  | ~\new_[11523]_  | ~\new_[11520]_  | ~\new_[13455]_ ;
  assign \s6_addr_o[26]  = ~\new_[13458]_  | ~\new_[11524]_  | ~\new_[13456]_  | ~\new_[13457]_ ;
  assign \s6_addr_o[25]  = ~\new_[11526]_  | ~\new_[11527]_  | ~\new_[11525]_  | ~\new_[13460]_ ;
  assign \s6_addr_o[24]  = ~\new_[13461]_  | ~\new_[11531]_  | ~\new_[11528]_  | ~\new_[11529]_ ;
  assign \s6_addr_o[23]  = ~\new_[11534]_  | ~\new_[11535]_  | ~\new_[11532]_  | ~\new_[13462]_ ;
  assign \s6_addr_o[22]  = ~\new_[14829]_  | ~\new_[11538]_  | ~\new_[11536]_  | ~\new_[13463]_ ;
  assign \s6_addr_o[21]  = ~\new_[11542]_  | ~\new_[11543]_  | ~\new_[11540]_  | ~\new_[9859]_ ;
  assign \s6_addr_o[20]  = ~\new_[11546]_  | ~\new_[11547]_  | ~\new_[11545]_  | ~\new_[9862]_ ;
  assign \s6_addr_o[19]  = ~\new_[11550]_  | ~\new_[13466]_  | ~\new_[11548]_  | ~\new_[9865]_ ;
  assign \new_[7734]_  = ~\new_[9302]_  & ~\new_[10668]_ ;
  assign \s6_addr_o[16]  = ~\new_[11560]_  | ~\new_[13467]_  | ~\new_[11558]_  | ~\new_[9873]_ ;
  assign \s6_addr_o[15]  = ~\new_[14832]_  | ~\new_[11563]_  | ~\new_[13468]_  | ~\new_[11562]_ ;
  assign \s6_addr_o[14]  = ~\new_[11566]_  | ~\new_[13469]_  | ~\new_[11565]_  | ~\new_[9876]_ ;
  assign \s6_addr_o[12]  = ~\new_[11573]_  | ~\new_[13470]_  | ~\new_[11571]_  | ~\new_[11572]_ ;
  assign \s6_addr_o[10]  = ~\new_[11578]_  | ~\new_[11580]_  | ~\new_[11576]_  | ~\new_[11577]_ ;
  assign \s6_addr_o[9]  = ~\new_[11582]_  | ~\new_[13471]_  | ~\new_[11581]_  | ~\new_[9885]_ ;
  assign \s6_addr_o[5]  = ~\new_[11595]_  | ~\new_[13472]_  | ~\new_[11594]_  | ~\new_[9898]_ ;
  assign \s6_addr_o[4]  = ~\new_[13473]_  | ~\new_[11599]_  | ~\new_[11596]_  | ~\new_[9900]_ ;
  assign \s6_addr_o[3]  = ~\new_[11601]_  | ~\new_[11602]_  | ~\new_[11600]_  | ~\new_[9902]_ ;
  assign n7449 = (~\new_[10541]_  & ~rst_i) | (~\new_[30982]_  & ~\new_[31597]_ );
  assign \s6_addr_o[2]  = ~\new_[11604]_  | ~\new_[11605]_  | ~\new_[11603]_  | ~\new_[13474]_ ;
  assign \s6_addr_o[0]  = ~\new_[11612]_  | ~\new_[13477]_  | ~\new_[11609]_  | ~\new_[11610]_ ;
  assign \s6_sel_o[3]  = ~\new_[11614]_  | ~\new_[11615]_  | ~\new_[13478]_  | ~\new_[9911]_ ;
  assign \s6_sel_o[2]  = ~\new_[14840]_  | ~\new_[11617]_  | ~\new_[13479]_  | ~\new_[13480]_ ;
  assign \s6_sel_o[1]  = ~\new_[11619]_  | ~\new_[11620]_  | ~\new_[13481]_  | ~\new_[13482]_ ;
  assign s6_we_o = ~\new_[11627]_  | ~\new_[11628]_  | ~\new_[11625]_  | ~\new_[11626]_ ;
  assign s6_stb_o = \new_[10944]_  | \new_[9416]_ ;
  assign \s7_data_o[31]  = ~\new_[11632]_  | ~\new_[11631]_  | ~\new_[11630]_  | ~\new_[13483]_ ;
  assign \s7_data_o[30]  = ~\new_[11635]_  | ~\new_[11636]_  | ~\new_[14841]_  | ~\new_[11634]_ ;
  assign \s7_data_o[28]  = ~\new_[11642]_  | ~\new_[11643]_  | ~\new_[14843]_  | ~\new_[11641]_ ;
  assign \s7_data_o[27]  = ~\new_[14845]_  | ~\new_[11646]_  | ~\new_[9919]_  | ~\new_[11645]_ ;
  assign \s7_data_o[26]  = ~\new_[14846]_  | ~\new_[11648]_  | ~\new_[9921]_  | ~\new_[11647]_ ;
  assign \s7_data_o[25]  = ~\new_[14847]_  | ~\new_[13484]_  | ~\new_[11649]_  | ~\new_[9922]_ ;
  assign \s7_data_o[24]  = ~\new_[14851]_  | ~\new_[13486]_  | ~\new_[11652]_  | ~\new_[9925]_ ;
  assign \s7_data_o[23]  = ~\new_[11655]_  | ~\new_[14853]_  | ~\new_[11653]_  | ~\new_[9928]_ ;
  assign \s7_data_o[22]  = ~\new_[11658]_  | ~\new_[11660]_  | ~\new_[11656]_  | ~\new_[13488]_ ;
  assign \s7_data_o[21]  = ~\new_[11662]_  | ~\new_[14854]_  | ~\new_[11661]_  | ~\new_[9934]_ ;
  assign \s7_data_o[20]  = ~\new_[14855]_  | ~\new_[13489]_  | ~\new_[11663]_  | ~\new_[9936]_ ;
  assign \s7_data_o[17]  = ~\new_[14858]_  | ~\new_[11669]_  | ~\new_[9942]_  | ~\new_[11668]_ ;
  assign \s7_data_o[16]  = ~\new_[11673]_  | ~\new_[13496]_  | ~\new_[14859]_  | ~\new_[9944]_ ;
  assign \s7_data_o[15]  = ~\new_[13498]_  | ~\new_[13499]_  | ~\new_[9947]_  | ~\new_[9948]_ ;
  assign \s7_data_o[14]  = ~\new_[13500]_  | ~\new_[13501]_  | ~\new_[9949]_  | ~\new_[9951]_ ;
  assign \s7_data_o[13]  = ~\new_[13502]_  | ~\new_[13503]_  | ~\new_[9953]_  | ~\new_[9954]_ ;
  assign \s7_data_o[12]  = ~\new_[14862]_  | ~\new_[13505]_  | ~\new_[11676]_  | ~\new_[9956]_ ;
  assign \new_[7769]_  = ~\new_[12036]_  & (~\new_[10831]_  | ~\new_[24495]_ );
  assign \s7_data_o[7]  = ~\new_[14865]_  | ~\new_[11686]_  | ~\new_[9965]_  | ~\new_[13510]_ ;
  assign \s7_data_o[5]  = ~\new_[13513]_  | ~\new_[13514]_  | ~\new_[11689]_  | ~\new_[9970]_ ;
  assign \s7_data_o[4]  = ~\new_[13515]_  | ~\new_[11691]_  | ~\new_[9971]_  | ~\new_[11690]_ ;
  assign \s7_data_o[1]  = ~\new_[11697]_  | ~\new_[14867]_  | ~\new_[9977]_  | ~\new_[9979]_ ;
  assign \s7_data_o[2]  = ~\new_[13517]_  | ~\new_[13518]_  | ~\new_[9976]_  | ~\new_[9975]_ ;
  assign \s7_addr_o[29]  = ~\new_[13521]_  | ~\new_[13522]_  | ~\new_[11706]_  | ~\new_[9985]_ ;
  assign \s7_addr_o[28]  = ~\new_[14873]_  | ~\new_[11709]_  | ~\new_[9988]_  | ~\new_[11708]_ ;
  assign \new_[7777]_  = ~\new_[9159]_  & ~\new_[12828]_ ;
  assign \s7_addr_o[24]  = ~\new_[14877]_  | ~\new_[11718]_  | ~\new_[11717]_  | ~\new_[9999]_ ;
  assign \s7_addr_o[21]  = ~\new_[11724]_  | ~\new_[11725]_  | ~\new_[14882]_  | ~\new_[11723]_ ;
  assign \new_[7780]_  = ~\new_[9373]_  & ~\new_[9222]_ ;
  assign \s7_addr_o[19]  = ~\new_[11731]_  | ~\new_[11730]_  | ~\new_[14884]_  | ~\new_[11729]_ ;
  assign \s7_addr_o[16]  = ~\new_[11737]_  | ~\new_[11738]_  | ~\new_[11736]_  | ~\new_[13529]_ ;
  assign \s7_addr_o[15]  = ~\new_[11740]_  | ~\new_[11742]_  | ~\new_[11739]_  | ~\new_[13532]_ ;
  assign \s7_addr_o[14]  = ~\new_[11744]_  | ~\new_[11745]_  | ~\new_[11743]_  | ~\new_[13533]_ ;
  assign \s7_addr_o[13]  = ~\new_[11749]_  | ~\new_[11750]_  | ~\new_[11747]_  | ~\new_[13534]_ ;
  assign \s7_addr_o[12]  = ~\new_[14890]_  | ~\new_[11754]_  | ~\new_[10018]_  | ~\new_[11752]_ ;
  assign \s7_addr_o[11]  = ~\new_[14891]_  | ~\new_[11757]_  | ~\new_[10019]_  | ~\new_[11756]_ ;
  assign \s7_addr_o[10]  = ~\new_[11760]_  | ~\new_[11762]_  | ~\new_[14892]_  | ~\new_[11758]_ ;
  assign \s7_addr_o[9]  = ~\new_[14893]_  | ~\new_[11766]_  | ~\new_[10020]_  | ~\new_[11765]_ ;
  assign \s7_addr_o[7]  = ~\new_[13538]_  | ~\new_[11772]_  | ~\new_[11771]_  | ~\new_[10025]_ ;
  assign \s7_addr_o[6]  = ~\new_[13540]_  | ~\new_[11775]_  | ~\new_[10029]_  | ~\new_[11774]_ ;
  assign \s7_addr_o[1]  = ~\new_[11787]_  | ~\new_[11788]_  | ~\new_[11785]_  | ~\new_[13547]_ ;
  assign \s7_sel_o[3]  = ~\new_[11792]_  | ~\new_[11793]_  | ~\new_[11790]_  | ~\new_[14898]_ ;
  assign \s7_sel_o[2]  = ~\new_[11795]_  | ~\new_[11798]_  | ~\new_[11794]_  | ~\new_[14899]_ ;
  assign \s7_sel_o[1]  = ~\new_[14900]_  | ~\new_[11801]_  | ~\new_[10049]_  | ~\new_[11800]_ ;
  assign \s7_sel_o[0]  = ~\new_[11803]_  | ~\new_[11804]_  | ~\new_[11802]_  | ~\new_[13548]_ ;
  assign s7_we_o = ~\new_[13550]_  | ~\new_[11805]_  | ~\new_[10051]_  | ~\new_[13549]_ ;
  assign \new_[7798]_  = ~\new_[12533]_  & ~\new_[9161]_ ;
  assign n7454 = (~\new_[10542]_  & ~rst_i) | (~\new_[30904]_  & ~\new_[31575]_ );
  assign \new_[7800]_  = ~\new_[9165]_  & ~\new_[12834]_ ;
  assign s11_cyc_o = ~n7539;
  assign \new_[7802]_  = ~\new_[12045]_  & (~\new_[10838]_  | ~\new_[24489]_ );
  assign \s10_data_o[31]  = ~\new_[14970]_  | ~\new_[12090]_  | ~\new_[13698]_  | ~\new_[12088]_ ;
  assign \s10_data_o[26]  = ~\new_[12104]_  | ~\new_[12105]_  | ~\new_[16346]_  | ~\new_[13708]_ ;
  assign \s10_data_o[25]  = ~\new_[12106]_  | ~\new_[12108]_  | ~\new_[13709]_  | ~\new_[14980]_ ;
  assign \s10_data_o[22]  = ~\new_[13715]_  | ~\new_[12115]_  | ~\new_[14984]_  | ~\new_[12114]_ ;
  assign \new_[7807]_  = ~\new_[9374]_  & ~\new_[9224]_ ;
  assign \s10_data_o[15]  = ~\new_[12128]_  | ~\new_[16348]_  | ~\new_[12127]_  | ~\new_[13726]_ ;
  assign \s10_data_o[14]  = ~\new_[13727]_  | ~\new_[12131]_  | ~\new_[12471]_  | ~\new_[15141]_ ;
  assign \s10_data_o[6]  = ~\new_[12157]_  | ~\new_[15011]_  | ~\new_[12155]_  | ~\new_[13743]_ ;
  assign \s10_data_o[2]  = ~\new_[12168]_  | ~\new_[15015]_  | ~\new_[15359]_  | ~\new_[13754]_ ;
  assign \s10_data_o[1]  = ~\new_[12172]_  | ~\new_[15016]_  | ~\new_[12169]_  | ~\new_[13756]_ ;
  assign \s10_data_o[0]  = ~\new_[12175]_  | ~\new_[16362]_  | ~\new_[12174]_  | ~\new_[13758]_ ;
  assign \s10_addr_o[30]  = ~\new_[16365]_  | ~\new_[12184]_  | ~\new_[12182]_  | ~\new_[13763]_ ;
  assign n7499 = ~\new_[10476]_  & ~\new_[9283]_ ;
  assign \s10_addr_o[28]  = ~\new_[12191]_  | ~\new_[15023]_  | ~\new_[16366]_  | ~\new_[12572]_ ;
  assign \s10_addr_o[27]  = ~\new_[12196]_  | ~\new_[15024]_  | ~\new_[13766]_  | ~\new_[12194]_ ;
  assign \s10_addr_o[26]  = ~\new_[11302]_  | ~\new_[15025]_  | ~\new_[12198]_  | ~\new_[16367]_ ;
  assign \s10_addr_o[25]  = ~\new_[12205]_  | ~\new_[15026]_  | ~\new_[13768]_  | ~\new_[11808]_ ;
  assign \s10_addr_o[24]  = ~\new_[12208]_  | ~\new_[13770]_  | ~\new_[16368]_  | ~\new_[12207]_ ;
  assign \s10_addr_o[23]  = ~\new_[16369]_  | ~\new_[12212]_  | ~\new_[13771]_  | ~\new_[13772]_ ;
  assign \new_[7822]_  = ~\new_[10679]_  & ~\new_[9176]_ ;
  assign \s10_addr_o[14]  = ~\new_[12242]_  | ~\new_[15046]_  | ~\new_[12241]_  | ~\new_[13789]_ ;
  assign \s10_addr_o[12]  = ~\new_[14926]_  | ~\new_[12247]_  | ~\new_[13794]_  | ~\new_[12246]_ ;
  assign \s10_addr_o[11]  = ~\new_[13799]_  | ~\new_[12249]_  | ~\new_[13798]_  | ~\new_[15054]_ ;
  assign \s10_addr_o[6]  = ~\new_[15076]_  | ~\new_[12262]_  | ~\new_[13807]_  | ~\new_[15073]_ ;
  assign n7459 = (~\new_[10544]_  & ~rst_i) | (~\new_[30916]_  & ~\new_[31935]_ );
  assign \s10_sel_o[0]  = ~\new_[15113]_  | ~\new_[12289]_  | ~\new_[13833]_  | ~\new_[16388]_ ;
  assign s10_we_o = ~\new_[13838]_  | ~\new_[12293]_  | ~\new_[15114]_  | ~\new_[12290]_ ;
  assign \s11_data_o[30]  = ~\new_[15195]_  | ~\new_[12305]_  | ~\new_[12300]_  | ~\new_[12301]_ ;
  assign \s11_data_o[29]  = ~\new_[15125]_  | ~\new_[12309]_  | ~\new_[12306]_  | ~\new_[12307]_ ;
  assign \s11_data_o[28]  = ~\new_[15128]_  | ~\new_[12315]_  | ~\new_[12310]_  | ~\new_[12313]_ ;
  assign \s11_data_o[26]  = ~\new_[12321]_  | ~\new_[15134]_  | ~\new_[12319]_  | ~\new_[12320]_ ;
  assign \s11_data_o[24]  = ~\new_[12329]_  | ~\new_[15138]_  | ~\new_[12327]_  | ~\new_[12328]_ ;
  assign \s11_data_o[15]  = ~\new_[13880]_  | ~\new_[15163]_  | ~\new_[11453]_  | ~\new_[10568]_ ;
  assign \s11_data_o[10]  = ~\new_[15175]_  | ~\new_[12365]_  | ~\new_[11229]_  | ~\new_[12363]_ ;
  assign \s11_data_o[6]  = ~\new_[13910]_  | ~\new_[15186]_  | ~\new_[12371]_  | ~\new_[10579]_ ;
  assign \s11_data_o[5]  = ~\new_[15189]_  | ~\new_[12376]_  | ~\new_[12373]_  | ~\new_[10580]_ ;
  assign \s11_data_o[2]  = ~\new_[15200]_  | ~\new_[12384]_  | ~\new_[12382]_  | ~\new_[10585]_ ;
  assign \s11_addr_o[24]  = ~\new_[15228]_  | ~\new_[12410]_  | ~\new_[9332]_  | ~\new_[12408]_ ;
  assign \s11_addr_o[15]  = ~\new_[12437]_  | ~\new_[13974]_  | ~\new_[12435]_  | ~\new_[15254]_ ;
  assign \s11_addr_o[14]  = ~\new_[14513]_  | ~\new_[12440]_  | ~\new_[12438]_  | ~\new_[11174]_ ;
  assign \s11_addr_o[5]  = ~\new_[13986]_  | ~\new_[12466]_  | ~\new_[14566]_  | ~\new_[10615]_ ;
  assign n7464 = ~\new_[9285]_  & ~\new_[10479]_ ;
  assign s11_we_o = ~\new_[12497]_  | ~\new_[13998]_  | ~\new_[15295]_  | ~\new_[12496]_ ;
  assign \s12_data_o[27]  = ~\new_[12505]_  | ~\new_[15307]_  | ~\new_[9342]_  | ~\new_[10643]_ ;
  assign \s12_data_o[8]  = ~\new_[11966]_  | ~\new_[12532]_  | ~\new_[9360]_  | ~\new_[15346]_ ;
  assign \s12_data_o[7]  = ~\new_[15349]_  | ~\new_[12534]_  | ~\new_[9098]_  | ~\new_[14041]_ ;
  assign \s12_data_o[1]  = ~\new_[15364]_  | ~\new_[14049]_  | ~\new_[9378]_  | ~\new_[10674]_ ;
  assign \s12_addr_o[28]  = ~\new_[14082]_  | ~\new_[15378]_  | ~\new_[10887]_  | ~\new_[10684]_ ;
  assign n7469 = ~\new_[12107]_  & ~\new_[9286]_ ;
  assign \s12_addr_o[26]  = ~\new_[14063]_  | ~\new_[15385]_  | ~\new_[10042]_  | ~\new_[10687]_ ;
  assign \s12_addr_o[24]  = ~\new_[15394]_  | ~\new_[14070]_  | ~\new_[10690]_  | ~\new_[10691]_ ;
  assign n7474 = ~\new_[9289]_  & ~\new_[10481]_ ;
  assign \s13_data_o[23]  = ~\new_[12633]_  | ~\new_[14139]_  | ~\new_[12632]_  | ~\new_[10752]_ ;
  assign \s13_data_o[22]  = ~\new_[12639]_  | ~\new_[14142]_  | ~\new_[10754]_  | ~\new_[12636]_ ;
  assign \s13_data_o[21]  = ~\new_[12643]_  | ~\new_[14146]_  | ~\new_[12641]_  | ~\new_[10756]_ ;
  assign \s13_data_o[20]  = ~\new_[12649]_  | ~\new_[14148]_  | ~\new_[12647]_  | ~\new_[10759]_ ;
  assign s2_cyc_o = ~n7544;
  assign \s13_data_o[11]  = ~\new_[14169]_  | ~\new_[12681]_  | ~\new_[12680]_  | ~\new_[10780]_ ;
  assign \s13_data_o[8]  = ~\new_[14177]_  | ~\new_[12688]_  | ~\new_[12685]_  | ~\new_[10786]_ ;
  assign \s13_data_o[5]  = ~\new_[12701]_  | ~\new_[12703]_  | ~\new_[12698]_  | ~\new_[14182]_ ;
  assign \s13_data_o[2]  = ~\new_[14192]_  | ~\new_[12712]_  | ~\new_[10795]_  | ~\new_[12711]_ ;
  assign \s13_data_o[1]  = ~\new_[12715]_  | ~\new_[14196]_  | ~\new_[10796]_  | ~\new_[12713]_ ;
  assign \s13_addr_o[29]  = ~\new_[14206]_  | ~\new_[12725]_  | ~\new_[10807]_  | ~\new_[10808]_ ;
  assign \s13_addr_o[27]  = ~\new_[12732]_  | ~\new_[12733]_  | ~\new_[12730]_  | ~\new_[12731]_ ;
  assign n7479 = ~\new_[9292]_  & ~\new_[12133]_ ;
  assign \s14_data_o[9]  = ~\new_[12877]_  | ~\new_[12878]_  | ~\new_[9431]_  | ~\new_[10958]_ ;
  assign \s14_data_o[10]  = ~\new_[12874]_  | ~\new_[12875]_  | ~\new_[9430]_  | ~\new_[10957]_ ;
  assign \new_[7870]_  = ~\new_[12062]_  & ~\new_[9096]_ ;
  assign \new_[7871]_  = ~\new_[9102]_  & ~\new_[9295]_ ;
  assign \new_[7872]_  = ~\new_[10238]_  & ~\new_[9296]_ ;
  assign \new_[7873]_  = ~\new_[12070]_  & ~\new_[9297]_ ;
  assign \new_[7874]_  = ~\new_[13688]_  & ~\new_[9127]_ ;
  assign \new_[7875]_  = ~\new_[9132]_  & ~\new_[9298]_ ;
  assign \new_[7876]_  = ~\new_[12083]_  & ~\new_[9299]_ ;
  assign \new_[7877]_  = ~\new_[12093]_  & ~\new_[9303]_ ;
  assign \new_[7878]_  = ~\new_[10517]_  & ~\new_[9168]_ ;
  assign \new_[7879]_  = ~\new_[12101]_  & ~\new_[9304]_ ;
  assign \new_[7880]_  = ~\new_[10351]_  & ~\new_[9305]_ ;
  assign \new_[7881]_  = ~\new_[12135]_  & ~\new_[9306]_ ;
  assign \new_[7882]_  = ~\new_[24718]_  | ~\new_[8990]_ ;
  assign \new_[7883]_  = ~\new_[25160]_  | ~\new_[8996]_ ;
  assign \new_[7884]_  = ~\new_[25165]_  | ~\new_[9002]_ ;
  assign \new_[7885]_  = ~\new_[19385]_  | ~\new_[9005]_ ;
  assign \s12_data_o[9]  = ~\new_[12530]_  | ~\new_[12531]_  | ~\new_[9359]_  | ~\new_[15342]_ ;
  assign \new_[7887]_  = ~\new_[19391]_  | ~\new_[9026]_ ;
  assign \new_[7888]_  = ~\new_[19392]_  | ~\new_[9036]_ ;
  assign \new_[7889]_  = ~\new_[29114]_  & (~\new_[10529]_  | ~\new_[22807]_ );
  assign \new_[7890]_  = ~\new_[9240]_  & (~\new_[11236]_  | ~\new_[30175]_ );
  assign \new_[7891]_  = ~\new_[25196]_  | ~\new_[9044]_ ;
  assign \new_[7892]_  = ~\new_[9243]_  & (~\new_[11237]_  | ~\new_[29358]_ );
  assign \new_[7893]_  = ~\new_[28653]_  & (~\new_[10530]_  | ~\new_[22707]_ );
  assign \new_[7894]_  = ~\new_[19393]_  | ~\new_[9052]_ ;
  assign \new_[7895]_  = ~\new_[25203]_  | ~\new_[9067]_ ;
  assign \new_[7896]_  = ~\new_[9249]_  & (~\new_[11965]_  | ~\new_[29337]_ );
  assign \new_[7897]_  = ~\new_[28260]_  & (~\new_[10531]_  | ~\new_[21422]_ );
  assign \new_[7898]_  = ~\new_[29424]_  & (~\new_[10555]_  | ~\new_[22949]_ );
  assign \new_[7899]_  = \new_[9009]_  | \new_[23103]_ ;
  assign \new_[7900]_  = ~\new_[28252]_  & (~\new_[10609]_  | ~\new_[22853]_ );
  assign \new_[7901]_  = ~\new_[26677]_  & (~\new_[10610]_  | ~\new_[29382]_ );
  assign \new_[7902]_  = ~\new_[28810]_  & (~\new_[10627]_  | ~\new_[23034]_ );
  assign \new_[7903]_  = ~\new_[27840]_  & (~\new_[10528]_  | ~\new_[27491]_ );
  assign \new_[7904]_  = ~\new_[28374]_  & (~\new_[10652]_  | ~\new_[22925]_ );
  assign \new_[7905]_  = ~\new_[28628]_  & (~\new_[10670]_  | ~\new_[29493]_ );
  assign \new_[7906]_  = ~\new_[27910]_  & (~\new_[10676]_  | ~\new_[27713]_ );
  assign \new_[7907]_  = ~\new_[28869]_  & (~\new_[10811]_  | ~\new_[21449]_ );
  assign \s12_data_o[13]  = ~\new_[14036]_  | ~\new_[12525]_  | ~\new_[9354]_  | ~\new_[15333]_ ;
  assign \new_[7909]_  = ~\new_[27916]_  & (~\new_[10717]_  | ~\new_[23041]_ );
  assign \new_[7910]_  = ~\new_[28145]_  & (~\new_[10841]_  | ~\new_[20428]_ );
  assign \new_[7911]_  = (~\new_[10630]_  | ~\new_[30408]_ ) & (~\new_[22713]_  | ~\new_[30408]_ );
  assign \new_[7912]_  = ~\new_[28131]_  & (~\new_[10596]_  | ~\new_[21431]_ );
  assign \new_[7913]_  = ~\new_[18414]_  | ~\new_[9314]_ ;
  assign n7504 = (~\new_[11155]_  & ~rst_i) | (~\new_[30453]_  & ~\new_[31935]_ );
  assign \new_[7915]_  = \\s9_msel_pri_out_reg[1] ;
  assign \new_[7916]_  = \\s4_msel_pri_out_reg[1] ;
  assign \new_[7917]_  = \\s14_msel_pri_out_reg[1] ;
  assign \new_[7918]_  = \\s10_msel_pri_out_reg[1] ;
  assign \new_[7919]_  = ~s1_next_reg;
  assign \new_[7920]_  = ~s10_next_reg;
  assign \new_[7921]_  = ~\s15_addr_o[4] ;
  assign \new_[7922]_  = ~\s15_addr_o[4] ;
  assign \new_[7923]_  = ~\new_[9317]_  & ~\new_[10549]_ ;
  assign \new_[7924]_  = \new_[9757]_  | \new_[9554]_ ;
  assign \new_[7925]_  = \new_[9758]_  | \new_[9555]_ ;
  assign \new_[7926]_  = \new_[9759]_  | \new_[9556]_ ;
  assign \new_[7927]_  = \new_[9760]_  | \new_[9557]_ ;
  assign \new_[7928]_  = \new_[9762]_  | \new_[9560]_ ;
  assign \new_[7929]_  = \new_[9763]_  | \new_[9561]_ ;
  assign \new_[7930]_  = \new_[9764]_  | \new_[9562]_ ;
  assign \new_[7931]_  = \new_[9765]_  | \new_[9563]_ ;
  assign \new_[7932]_  = \new_[9767]_  | \new_[9564]_ ;
  assign \new_[7933]_  = ~\new_[9536]_  & ~\new_[11103]_ ;
  assign \new_[7934]_  = ~\new_[9538]_  & ~\new_[9539]_ ;
  assign \new_[7935]_  = ~\new_[9540]_  & ~\new_[9541]_ ;
  assign \new_[7936]_  = ~\new_[21179]_  | ~\new_[11381]_  | ~\new_[19351]_  | ~\new_[10370]_ ;
  assign \new_[7937]_  = ~\new_[9542]_  & ~\new_[9543]_ ;
  assign \new_[7938]_  = ~\new_[9546]_  & ~\new_[9547]_ ;
  assign \new_[7939]_  = ~\new_[9567]_  & (~\new_[17139]_  | ~\new_[29547]_ );
  assign \new_[7940]_  = ~\new_[9568]_  & (~\new_[13424]_  | ~\new_[28034]_ );
  assign \new_[7941]_  = ~\new_[9569]_  & (~\new_[16231]_  | ~\new_[30182]_ );
  assign \new_[7942]_  = ~\new_[9571]_  & (~\new_[16234]_  | ~\new_[29760]_ );
  assign \new_[7943]_  = ~\new_[9551]_  & (~\new_[14773]_  | ~\new_[27894]_ );
  assign \new_[7944]_  = ~\new_[9552]_  & (~\new_[17146]_  | ~\new_[26484]_ );
  assign \new_[7945]_  = ~\new_[8654]_  & (~\new_[17148]_  | ~\new_[29110]_ );
  assign \new_[7946]_  = ~\new_[8655]_  & (~\new_[14818]_  | ~\new_[29160]_ );
  assign \new_[7947]_  = ~\new_[8656]_  & (~\new_[17153]_  | ~\new_[29538]_ );
  assign \new_[7948]_  = ~\new_[8657]_  & (~\new_[13434]_  | ~\new_[29143]_ );
  assign \new_[7949]_  = ~\new_[9570]_  & (~\new_[11411]_  | ~\new_[28367]_ );
  assign \new_[7950]_  = ~\new_[8653]_  & (~\new_[16162]_  | ~\new_[28100]_ );
  assign \new_[7951]_  = ~\new_[8790]_  & ~\new_[9897]_ ;
  assign \new_[7952]_  = ~\new_[8751]_  & ~\new_[8953]_ ;
  assign \new_[7953]_  = ~\new_[8768]_  & ~\new_[8972]_ ;
  assign \new_[7954]_  = ~\new_[8792]_  & ~\new_[11978]_ ;
  assign \new_[7955]_  = ~\new_[8793]_  & ~\new_[11979]_ ;
  assign \new_[7956]_  = ~\new_[8794]_  & ~\new_[11980]_ ;
  assign \new_[7957]_  = ~\new_[8795]_  & ~\new_[11981]_ ;
  assign \new_[7958]_  = ~\new_[8797]_  & ~\new_[11982]_ ;
  assign \new_[7959]_  = ~\new_[8798]_  & ~\new_[11983]_ ;
  assign \new_[7960]_  = ~\new_[8799]_  & ~\new_[11984]_ ;
  assign \new_[7961]_  = ~\new_[8800]_  & ~\new_[11985]_ ;
  assign \new_[7962]_  = ~\new_[8801]_  & ~\new_[11987]_ ;
  assign \new_[7963]_  = ~\new_[8802]_  & ~\new_[11988]_ ;
  assign \new_[7964]_  = (~\new_[10160]_  | ~\new_[29144]_ ) & (~\new_[14927]_  | ~\new_[29730]_ );
  assign \new_[7965]_  = ~\new_[8803]_  & ~\new_[13656]_ ;
  assign \new_[7966]_  = ~\new_[8804]_  & ~\new_[11989]_ ;
  assign \new_[7967]_  = (~\new_[10172]_  | ~\new_[28822]_ ) & (~\new_[13607]_  | ~\new_[28771]_ );
  assign \new_[7968]_  = (~\new_[10174]_  | ~\new_[28854]_ ) & (~\new_[11895]_  | ~\new_[28025]_ );
  assign \new_[7969]_  = ~\new_[8805]_  & ~\new_[11990]_ ;
  assign \new_[7970]_  = ~\new_[8806]_  & ~\new_[11991]_ ;
  assign \new_[7971]_  = ~\new_[9874]_  & ~\new_[8887]_ ;
  assign \new_[7972]_  = ~\new_[9878]_  & ~\new_[8888]_ ;
  assign \new_[7973]_  = ~\new_[8889]_  & ~\new_[11570]_ ;
  assign \new_[7974]_  = ~\new_[9891]_  & ~\new_[8894]_ ;
  assign \new_[7975]_  = ~\new_[9903]_  & ~\new_[8896]_ ;
  assign \new_[7976]_  = ~\new_[9904]_  & ~\new_[8898]_ ;
  assign \new_[7977]_  = ~\new_[8900]_  & ~\new_[9910]_ ;
  assign \new_[7978]_  = ~\new_[9912]_  & ~\new_[8902]_ ;
  assign \new_[7979]_  = ~\new_[11638]_  & ~\new_[8905]_ ;
  assign \new_[7980]_  = ~\new_[9920]_  & ~\new_[8908]_ ;
  assign \new_[7981]_  = ~\new_[10001]_  & ~\new_[8876]_ ;
  assign \new_[7982]_  = ~\new_[9927]_  & ~\new_[8913]_ ;
  assign \new_[7983]_  = ~\new_[9940]_  & ~\new_[8918]_ ;
  assign \new_[7984]_  = ~\new_[8919]_  & ~\new_[13495]_ ;
  assign \new_[7985]_  = ~\new_[9946]_  & ~\new_[8922]_ ;
  assign \new_[7986]_  = ~\new_[8925]_  & ~\new_[11549]_ ;
  assign \new_[7987]_  = ~\new_[13465]_  & ~\new_[8807]_ ;
  assign \new_[7988]_  = ~\new_[8707]_  & ~\new_[8852]_ ;
  assign \new_[7989]_  = ~\new_[8928]_  & ~\new_[9872]_ ;
  assign \new_[7990]_  = ~\new_[9688]_  & (~\new_[10097]_  | ~\new_[27838]_ );
  assign \new_[7991]_  = ~\new_[9690]_  & ~\new_[8854]_ ;
  assign \s0_addr_o[29]  = ~\new_[12282]_  | ~\new_[12283]_  | ~\new_[13828]_  | ~\new_[10540]_ ;
  assign \new_[7993]_  = ~\new_[8930]_  & ~\new_[8855]_ ;
  assign \new_[7994]_  = ~\new_[9696]_  & ~\new_[8856]_ ;
  assign \new_[7995]_  = ~\new_[11767]_  & ~\new_[8857]_ ;
  assign \new_[7996]_  = ~\new_[9789]_  & (~\new_[10110]_  | ~\new_[26635]_ );
  assign \new_[7997]_  = ~\new_[9702]_  & (~\new_[10119]_  | ~\new_[23138]_ );
  assign \new_[7998]_  = ~\new_[11586]_  & ~\new_[8813]_ ;
  assign \new_[7999]_  = ~\new_[11441]_  & (~\new_[10120]_  | ~\new_[23138]_ );
  assign \new_[8000]_  = ~\new_[11344]_  | ~\new_[11345]_  | ~\new_[14638]_  | ~\new_[13252]_ ;
  assign \new_[8001]_  = ~\new_[8720]_  & ~\new_[8859]_ ;
  assign \new_[8002]_  = ~\new_[8722]_  & (~\new_[10125]_  | ~\new_[23176]_ );
  assign \new_[8003]_  = ~\new_[14657]_  | ~\new_[11354]_  | ~\new_[11353]_  | ~\new_[16063]_ ;
  assign \new_[8004]_  = ~\new_[8724]_  & ~\new_[8723]_ ;
  assign \new_[8005]_  = ~\new_[9706]_  & (~\new_[10128]_  | ~\new_[23094]_ );
  assign \new_[8006]_  = ~\new_[11363]_  | ~\new_[17867]_  | ~\new_[13272]_  | ~\new_[14778]_ ;
  assign \new_[8007]_  = ~\new_[8791]_  & (~\new_[11905]_  | ~\new_[28332]_ );
  assign \new_[8008]_  = ~\new_[8726]_  & ~\new_[8815]_ ;
  assign \new_[8009]_  = ~\new_[13282]_  | ~\new_[14783]_  | ~\new_[9736]_  | ~\new_[9771]_ ;
  assign \new_[8010]_  = ~\new_[8728]_  & (~\new_[10138]_  | ~\new_[28666]_ );
  assign \new_[8011]_  = ~\new_[8938]_  & ~\new_[11597]_ ;
  assign \new_[8012]_  = ~\new_[11367]_  | ~\new_[14792]_  | ~\new_[16101]_  | ~\new_[13393]_ ;
  assign \new_[8013]_  = ~\new_[11450]_  & (~\new_[10140]_  | ~\new_[23092]_ );
  assign \new_[8014]_  = ~\new_[8730]_  & ~\new_[8861]_ ;
  assign \new_[8015]_  = ~\new_[8732]_  & (~\new_[10142]_  | ~\new_[28660]_ );
  assign \new_[8016]_  = ~\new_[9713]_  & (~\new_[10144]_  | ~\new_[26586]_ );
  assign \new_[8017]_  = ~\new_[13475]_  & ~\new_[8819]_ ;
  assign \new_[8018]_  = ~\new_[13307]_  | ~\new_[11409]_  | ~\new_[16205]_  | ~\new_[16206]_ ;
  assign \new_[8019]_  = ~\new_[11377]_  | ~\new_[14808]_  | ~\new_[11376]_  | ~\new_[14807]_ ;
  assign \new_[8020]_  = ~\new_[8735]_  & ~\new_[8864]_ ;
  assign \new_[8021]_  = ~\new_[8942]_  & ~\new_[8866]_ ;
  assign \new_[8022]_  = ~\new_[9808]_  & (~\new_[10147]_  | ~\new_[26946]_ );
  assign \new_[8023]_  = ~\new_[11385]_  | ~\new_[13418]_  | ~\new_[14731]_  | ~\new_[14814]_ ;
  assign \new_[8024]_  = ~\new_[9716]_  & ~\new_[8868]_ ;
  assign \new_[8025]_  = ~\new_[8945]_  & ~\new_[9914]_ ;
  assign \new_[8026]_  = ~\new_[11464]_  & (~\new_[10150]_  | ~\new_[29637]_ );
  assign \new_[8027]_  = ~\new_[9723]_  & ~\new_[8871]_ ;
  assign \new_[8028]_  = ~\new_[8742]_  & ~\new_[8872]_ ;
  assign \new_[8029]_  = ~\new_[10048]_  & ~\new_[8873]_ ;
  assign \new_[8030]_  = ~\new_[8825]_  & ~\new_[11644]_ ;
  assign \new_[8031]_  = ~\new_[8826]_  & (~\new_[10159]_  | ~\new_[29102]_ );
  assign \new_[8032]_  = ~\new_[8955]_  & ~\new_[9924]_ ;
  assign \new_[8033]_  = ~\new_[9737]_  & ~\new_[8878]_ ;
  assign \new_[8034]_  = ~\new_[8960]_  & ~\new_[9932]_ ;
  assign \new_[8035]_  = ~\new_[9741]_  & (~\new_[10169]_  | ~\new_[24569]_ );
  assign \new_[8036]_  = ~\new_[8759]_  & ~\new_[8880]_ ;
  assign \new_[8037]_  = ~\new_[9743]_  & (~\new_[10178]_  | ~\new_[27956]_ );
  assign \new_[8038]_  = (~\new_[13649]_  | ~\new_[28698]_ ) & (~\new_[10352]_  | ~\new_[28689]_ );
  assign \new_[8039]_  = (~\new_[13526]_  | ~\m4_data_i[29] ) & (~\new_[14850]_  | ~\m5_data_i[29] );
  assign \new_[8040]_  = ~\new_[8765]_  & (~\new_[10188]_  | ~\new_[29017]_ );
  assign \new_[8041]_  = ~\new_[8761]_  & (~\new_[10177]_  | ~\new_[28206]_ );
  assign \new_[8042]_  = ~\new_[9749]_  & (~\new_[10189]_  | ~\new_[24509]_ );
  assign \new_[8043]_  = ~\new_[8831]_  & ~\new_[11672]_ ;
  assign \new_[8044]_  = (~\new_[13526]_  | ~\m4_data_i[22] ) & (~\new_[9923]_  | ~\m5_data_i[22] );
  assign \new_[8045]_  = ~\new_[11491]_  & (~\new_[10191]_  | ~\new_[24509]_ );
  assign \new_[8046]_  = (~\new_[13526]_  | ~\m4_data_i[21] ) & (~\new_[14850]_  | ~\m5_data_i[21] );
  assign \new_[8047]_  = (~\new_[13651]_  | ~\new_[27759]_ ) & (~\new_[10364]_  | ~\new_[28320]_ );
  assign \new_[8048]_  = ~\new_[8767]_  & ~\new_[8883]_ ;
  assign \new_[8049]_  = (~\new_[13526]_  | ~\m4_data_i[19] ) & (~\new_[14850]_  | ~\m5_data_i[19] );
  assign \new_[8050]_  = ~\new_[9754]_  & (~\new_[10197]_  | ~\new_[29567]_ );
  assign \new_[8051]_  = ~\new_[8714]_  & ~\new_[8890]_ ;
  assign \new_[8052]_  = ~\new_[8717]_  & ~\new_[8892]_ ;
  assign \new_[8053]_  = ~\new_[8893]_  & ~\new_[9704]_ ;
  assign \new_[8054]_  = ~\new_[8897]_  & ~\new_[9711]_ ;
  assign \new_[8055]_  = ~\new_[8734]_  & ~\new_[8901]_ ;
  assign \new_[8056]_  = ~\new_[9993]_  & ~\new_[8741]_ ;
  assign \new_[8057]_  = ~\new_[8756]_  & ~\new_[10008]_ ;
  assign \new_[8058]_  = ~\new_[8917]_  & ~\new_[8762]_ ;
  assign \new_[8059]_  = ~\new_[8763]_  & ~\new_[10013]_ ;
  assign \new_[8060]_  = ~\new_[10203]_  & ~\new_[8924]_ ;
  assign \new_[8061]_  = ~\new_[9091]_  & ~\new_[8927]_ ;
  assign \new_[8062]_  = ~\new_[9100]_  & ~\new_[8931]_ ;
  assign \new_[8063]_  = ~\new_[9105]_  & ~\new_[10021]_ ;
  assign \new_[8064]_  = ~\new_[8812]_  & ~\new_[8774]_ ;
  assign \new_[8065]_  = ~\new_[9122]_  & ~\new_[9950]_ ;
  assign \new_[8066]_  = ~\new_[9123]_  & ~\new_[8860]_ ;
  assign \new_[8067]_  = ~\new_[10255]_  & ~\new_[8937]_ ;
  assign \new_[8068]_  = ~\new_[8817]_  & ~\new_[8776]_ ;
  assign \new_[8069]_  = ~\new_[9131]_  & ~\new_[8862]_ ;
  assign \new_[8070]_  = ~\new_[10282]_  & ~\new_[8941]_ ;
  assign \new_[8071]_  = ~\new_[8820]_  & ~\new_[8778]_ ;
  assign \new_[8072]_  = ~\new_[9145]_  & ~\new_[8944]_ ;
  assign \new_[8073]_  = ~\new_[8822]_  & ~\new_[8780]_ ;
  assign \new_[8074]_  = ~\new_[9153]_  & ~\new_[8947]_ ;
  assign \new_[8075]_  = ~\new_[9167]_  & ~\new_[8954]_ ;
  assign \new_[8076]_  = ~\new_[10340]_  & ~\new_[8959]_ ;
  assign \new_[8077]_  = ~\new_[9181]_  & ~\new_[8881]_ ;
  assign \new_[8078]_  = ~\new_[9185]_  & ~\new_[10060]_ ;
  assign \new_[8079]_  = ~\new_[9190]_  & ~\new_[8882]_ ;
  assign \new_[8080]_  = ~\new_[8788]_  & ~\new_[8833]_ ;
  assign \new_[8081]_  = ~\new_[9198]_  & ~\new_[8884]_ ;
  assign \new_[8082]_  = ~\new_[20316]_  | ~\new_[11852]_  | ~\new_[20377]_  | ~\new_[13809]_ ;
  assign \new_[8083]_  = ~\new_[8885]_  | ~\new_[11746]_ ;
  assign s4_cyc_o = ~n7549;
  assign \new_[8085]_  = ~\new_[18412]_  | ~\new_[11814]_  | ~\new_[20376]_  | ~\new_[15576]_ ;
  assign \new_[8086]_  = ~\new_[18409]_  | ~\new_[11816]_  | ~\new_[18408]_  | ~\new_[14260]_ ;
  assign \new_[8087]_  = ~\new_[19389]_  | ~\new_[11817]_  | ~\new_[21282]_  | ~\new_[14269]_ ;
  assign \new_[8088]_  = (~\new_[13526]_  | ~\m4_addr_i[17] ) & (~\new_[14850]_  | ~\m5_addr_i[17] );
  assign \new_[8089]_  = ~\new_[18411]_  | ~\new_[11819]_  | ~\new_[21288]_  | ~\new_[14274]_ ;
  assign \new_[8090]_  = ~\new_[18413]_  | ~\new_[11821]_  | ~\new_[21296]_  | ~\new_[14282]_ ;
  assign \new_[8091]_  = (~\new_[13526]_  | ~\m4_addr_i[14] ) & (~\new_[9923]_  | ~\m5_addr_i[14] );
  assign \new_[8092]_  = (~\new_[13526]_  | ~\m4_addr_i[13] ) & (~\new_[9923]_  | ~\m5_addr_i[13] );
  assign \new_[8093]_  = (~\new_[13526]_  | ~\m4_addr_i[12] ) & (~\new_[9923]_  | ~\m5_addr_i[12] );
  assign \new_[8094]_  = ~\new_[21306]_  | ~\new_[11823]_  | ~\new_[20381]_  | ~\new_[15627]_ ;
  assign \new_[8095]_  = ~\new_[19394]_  | ~\new_[11824]_  | ~\new_[21303]_  | ~\new_[14303]_ ;
  assign \new_[8096]_  = ~\new_[8909]_  | ~\new_[8952]_ ;
  assign \new_[8097]_  = ~\new_[19395]_  | ~\new_[11826]_  | ~\new_[21320]_  | ~\new_[14310]_ ;
  assign \new_[8098]_  = ~\new_[8911]_  | ~\new_[10053]_ ;
  assign \new_[8099]_  = ~\new_[18416]_  | ~\new_[11827]_  | ~\new_[21319]_  | ~\new_[12840]_ ;
  assign \new_[8100]_  = ~\new_[8914]_  | ~\new_[8962]_ ;
  assign \new_[8101]_  = ~\new_[21318]_  | ~\new_[11828]_  | ~\new_[17377]_  | ~\new_[14320]_ ;
  assign \new_[8102]_  = ~\new_[8916]_  | ~\new_[10063]_ ;
  assign \new_[8103]_  = ~\new_[8923]_  | ~\new_[13553]_ ;
  assign \new_[8104]_  = ~\new_[22486]_  | ~\new_[11830]_  | ~\new_[20326]_  | ~\new_[11856]_ ;
  assign \new_[8105]_  = ~\new_[18398]_  | (~\new_[10501]_  & ~\new_[26630]_ );
  assign \new_[8106]_  = ~\new_[17373]_  | (~\new_[10498]_  & ~\new_[27995]_ );
  assign \new_[8107]_  = ~\new_[19374]_  | (~\new_[12158]_  & ~\new_[29005]_ );
  assign \new_[8108]_  = ~\new_[19356]_  | (~\new_[12161]_  & ~\new_[26332]_ );
  assign \new_[8109]_  = ~\new_[20324]_  | (~\new_[12163]_  & ~\new_[26719]_ );
  assign \new_[8110]_  = ~\new_[19357]_  | (~\new_[12164]_  & ~\new_[27850]_ );
  assign \new_[8111]_  = ~\new_[19350]_  | (~\new_[12167]_  & ~\new_[28931]_ );
  assign \new_[8112]_  = ~\new_[19360]_  | (~\new_[12170]_  & ~\new_[26877]_ );
  assign \new_[8113]_  = ~\new_[20331]_  | (~\new_[12173]_  & ~\new_[26683]_ );
  assign \new_[8114]_  = ~\new_[19353]_  | (~\new_[12176]_  & ~\new_[30007]_ );
  assign \new_[8115]_  = ~\new_[20340]_  | (~\new_[12181]_  & ~\new_[28290]_ );
  assign \new_[8116]_  = ~\new_[20341]_  | (~\new_[12183]_  & ~\new_[27843]_ );
  assign \new_[8117]_  = ~\new_[21212]_  | (~\new_[12185]_  & ~\new_[27891]_ );
  assign \new_[8118]_  = ~\new_[19363]_  | (~\new_[12186]_  & ~\new_[28973]_ );
  assign \new_[8119]_  = ~\new_[21231]_  | (~\new_[12190]_  & ~\new_[28254]_ );
  assign \new_[8120]_  = ~\new_[19364]_  | (~\new_[12193]_  & ~\new_[28032]_ );
  assign \new_[8121]_  = ~\new_[21195]_  | (~\new_[12195]_  & ~\new_[26654]_ );
  assign \new_[8122]_  = ~\new_[20354]_  | (~\new_[12197]_  & ~\new_[27885]_ );
  assign \new_[8123]_  = ~\new_[19358]_  | (~\new_[12199]_  & ~\new_[26501]_ );
  assign \new_[8124]_  = ~\new_[21249]_  | (~\new_[12201]_  & ~\new_[27869]_ );
  assign \new_[8125]_  = ~\new_[20333]_  | (~\new_[12204]_  & ~\new_[27858]_ );
  assign \new_[8126]_  = ~\new_[18399]_  | (~\new_[12209]_  & ~\new_[28752]_ );
  assign \new_[8127]_  = ~\new_[20350]_  | (~\new_[12206]_  & ~\new_[28264]_ );
  assign \new_[8128]_  = ~\new_[20360]_  | (~\new_[12210]_  & ~\new_[24742]_ );
  assign \new_[8129]_  = ~\new_[19379]_  | (~\new_[12214]_  & ~\new_[27889]_ );
  assign n7549 = ~\new_[12059]_  & ~\new_[10446]_ ;
  assign \new_[8131]_  = ~\new_[15269]_  & ~\new_[10491]_ ;
  assign \new_[8132]_  = ~\new_[10212]_  & ~\new_[12770]_ ;
  assign \new_[8133]_  = ~\new_[10492]_  & ~\new_[12462]_ ;
  assign \new_[8134]_  = ~\new_[12774]_  & ~\new_[10224]_ ;
  assign n7589 = ~\new_[10451]_  & ~\new_[12064]_ ;
  assign \new_[8136]_  = ~\new_[15283]_  & ~\new_[10494]_ ;
  assign \new_[8137]_  = ~\new_[10234]_  & ~\new_[12779]_ ;
  assign \new_[8138]_  = ~\new_[10622]_  & ~\new_[12152]_ ;
  assign \new_[8139]_  = ~\new_[10404]_  | ~\new_[28510]_ ;
  assign \new_[8140]_  = ~\new_[13997]_  & ~\new_[10500]_ ;
  assign n7594 = (~\new_[12261]_  & ~rst_i) | (~\new_[31076]_  & ~\new_[31888]_ );
  assign \new_[8142]_  = ~\new_[10407]_  | ~\new_[26769]_ ;
  assign \new_[8143]_  = ~\new_[14262]_  & ~\new_[10377]_ ;
  assign \new_[8144]_  = ~\new_[10379]_  & ~\new_[14966]_ ;
  assign \new_[8145]_  = ~\new_[14005]_  & ~\new_[10441]_ ;
  assign \new_[8146]_  = ~\new_[10253]_  & ~\new_[12801]_ ;
  assign \s1_data_o[31]  = ~\new_[14048]_  | ~\new_[14050]_  | ~\new_[10816]_  | ~\new_[15363]_ ;
  assign \s1_data_o[30]  = ~\new_[13298]_  | ~\new_[15370]_  | ~\new_[10675]_  | ~\new_[15367]_ ;
  assign \s1_data_o[29]  = ~\new_[14055]_  | ~\new_[15376]_  | ~\new_[9647]_  | ~\new_[15374]_ ;
  assign \s1_data_o[27]  = ~\new_[15389]_  | ~\new_[15391]_  | ~\new_[10688]_  | ~\new_[15387]_ ;
  assign \s1_data_o[17]  = ~\new_[15447]_  | ~\new_[14256]_  | ~\new_[10715]_  | ~\new_[15444]_ ;
  assign \s1_data_o[18]  = ~\new_[15440]_  | ~\new_[14102]_  | ~\new_[10712]_  | ~\new_[14942]_ ;
  assign \s1_data_o[15]  = ~\new_[15457]_  | ~\new_[14108]_  | ~\new_[10723]_  | ~\new_[13414]_ ;
  assign \s1_data_o[13]  = ~\new_[15462]_  | ~\new_[14113]_  | ~\new_[15461]_  | ~\new_[12600]_ ;
  assign \s1_data_o[6]  = ~\new_[15479]_  | ~\new_[15480]_  | ~\new_[14135]_  | ~\new_[12629]_ ;
  assign \new_[8156]_  = ~\new_[10503]_  & ~\new_[12504]_ ;
  assign \s1_data_o[4]  = ~\new_[15485]_  | ~\new_[14150]_  | ~\new_[14145]_  | ~\new_[12645]_ ;
  assign \s1_data_o[3]  = ~\new_[15487]_  | ~\new_[14153]_  | ~\new_[15486]_  | ~\new_[12655]_ ;
  assign \s1_data_o[1]  = ~\new_[15495]_  | ~\new_[14162]_  | ~\new_[14159]_  | ~\new_[12671]_ ;
  assign \s1_data_o[0]  = ~\new_[15499]_  | ~\new_[15501]_  | ~\new_[10778]_  | ~\new_[15497]_ ;
  assign \new_[8161]_  = ~\new_[14011]_  & ~\new_[10504]_ ;
  assign \s1_addr_o[30]  = ~\new_[15508]_  | ~\new_[14179]_  | ~\new_[15506]_  | ~\new_[12684]_ ;
  assign \s1_addr_o[28]  = ~\new_[14184]_  | ~\new_[14186]_  | ~\new_[12699]_  | ~\new_[15518]_ ;
  assign \s1_addr_o[27]  = ~\new_[14191]_  | ~\new_[14193]_  | ~\new_[15523]_  | ~\new_[12710]_ ;
  assign \s1_addr_o[26]  = ~\new_[15528]_  | ~\new_[14200]_  | ~\new_[12714]_  | ~\new_[14198]_ ;
  assign \s1_addr_o[25]  = ~\new_[14205]_  | ~\new_[14203]_  | ~\new_[12720]_  | ~\new_[15532]_ ;
  assign \s1_addr_o[22]  = ~\new_[14220]_  | ~\new_[15549]_  | ~\new_[10817]_  | ~\new_[14218]_ ;
  assign \s1_addr_o[20]  = ~\new_[14230]_  | ~\new_[15555]_  | ~\new_[10835]_  | ~\new_[14227]_ ;
  assign n7519 = (~\new_[12270]_  & ~rst_i) | (~\new_[30878]_  & ~\new_[31576]_ );
  assign \s1_addr_o[12]  = ~\new_[14263]_  | ~\new_[14264]_  | ~\new_[10880]_  | ~\new_[15595]_ ;
  assign \s1_sel_o[2]  = ~\new_[14329]_  | ~\new_[15655]_  | ~\new_[10939]_  | ~\new_[14330]_ ;
  assign \new_[8172]_  = ~\new_[10267]_  & ~\new_[12809]_ ;
  assign \new_[8173]_  = ~\new_[14018]_  & ~\new_[10277]_ ;
  assign n7514 = (~\new_[12275]_  & ~rst_i) | (~\new_[31091]_  & ~\new_[31759]_ );
  assign \new_[8175]_  = ~\new_[10414]_  | ~\new_[28554]_ ;
  assign \new_[8176]_  = ~\new_[10286]_  & ~\new_[12515]_ ;
  assign \new_[8177]_  = ~\new_[14025]_  & ~\new_[10509]_ ;
  assign \new_[8178]_  = ~\new_[10418]_  | ~\new_[28186]_ ;
  assign \s5_data_o[30]  = ~\new_[13220]_  | ~\new_[13221]_  | ~\new_[11305]_  | ~\new_[14600]_ ;
  assign \s5_data_o[23]  = ~\new_[13231]_  | ~\new_[13232]_  | ~\new_[14609]_  | ~\new_[13230]_ ;
  assign \s5_data_o[21]  = ~\new_[13234]_  | ~\new_[13235]_  | ~\new_[11327]_  | ~\new_[14613]_ ;
  assign \s5_data_o[20]  = ~\new_[13237]_  | ~\new_[13238]_  | ~\new_[11328]_  | ~\new_[14614]_ ;
  assign \s5_data_o[18]  = ~\new_[13240]_  | ~\new_[13241]_  | ~\new_[11331]_  | ~\new_[14619]_ ;
  assign \s5_data_o[4]  = ~\new_[13270]_  | ~\new_[14663]_  | ~\new_[11361]_  | ~\new_[13269]_ ;
  assign \s5_data_o[3]  = ~\new_[13274]_  | ~\new_[14664]_  | ~\new_[11362]_  | ~\new_[13273]_ ;
  assign \s5_data_o[2]  = ~\new_[13276]_  | ~\new_[13277]_  | ~\new_[14665]_  | ~\new_[11364]_ ;
  assign \s5_data_o[0]  = ~\new_[13280]_  | ~\new_[13281]_  | ~\new_[14668]_  | ~\new_[11366]_ ;
  assign \new_[8188]_  = ~\new_[12085]_  & ~\new_[10664]_ ;
  assign \s5_addr_o[31]  = ~\new_[13284]_  | ~\new_[13285]_  | ~\new_[14669]_  | ~\new_[14670]_ ;
  assign \s5_addr_o[30]  = ~\new_[13287]_  | ~\new_[14675]_  | ~\new_[14672]_  | ~\new_[13286]_ ;
  assign \s5_addr_o[29]  = ~\new_[13290]_  | ~\new_[13289]_  | ~\new_[14676]_  | ~\new_[13288]_ ;
  assign \s5_addr_o[28]  = ~\new_[13292]_  | ~\new_[14681]_  | ~\new_[13291]_  | ~\new_[14680]_ ;
  assign \s5_addr_o[27]  = ~\new_[13295]_  | ~\new_[14684]_  | ~\new_[14682]_  | ~\new_[13294]_ ;
  assign \s5_addr_o[26]  = ~\new_[13297]_  | ~\new_[14690]_  | ~\new_[14686]_  | ~\new_[13296]_ ;
  assign \s5_addr_o[25]  = ~\new_[13300]_  | ~\new_[14694]_  | ~\new_[14692]_  | ~\new_[13299]_ ;
  assign \s5_addr_o[24]  = ~\new_[13302]_  | ~\new_[13301]_  | ~\new_[14695]_  | ~\new_[14696]_ ;
  assign \new_[8197]_  = ~\new_[15331]_  & ~\new_[10301]_ ;
  assign \s5_addr_o[20]  = ~\new_[13309]_  | ~\new_[13310]_  | ~\new_[11378]_  | ~\new_[14703]_ ;
  assign \s5_addr_o[19]  = ~\new_[13312]_  | ~\new_[13314]_  | ~\new_[11379]_  | ~\new_[14708]_ ;
  assign \s5_addr_o[17]  = ~\new_[13322]_  | ~\new_[14720]_  | ~\new_[14716]_  | ~\new_[13319]_ ;
  assign \s5_addr_o[16]  = ~\new_[13325]_  | ~\new_[13326]_  | ~\new_[14723]_  | ~\new_[14724]_ ;
  assign n7599 = (~\new_[12280]_  & ~rst_i) | (~\new_[30496]_  & ~\new_[31830]_ );
  assign \s5_addr_o[15]  = ~\new_[13327]_  | ~\new_[13328]_  | ~\new_[14726]_  | ~\new_[14727]_ ;
  assign \s5_addr_o[14]  = ~\new_[13329]_  | ~\new_[13330]_  | ~\new_[14728]_  | ~\new_[14729]_ ;
  assign \s5_addr_o[13]  = ~\new_[13333]_  | ~\new_[13332]_  | ~\new_[14730]_  | ~\new_[13331]_ ;
  assign \s5_addr_o[12]  = ~\new_[13335]_  | ~\new_[14734]_  | ~\new_[11386]_  | ~\new_[13334]_ ;
  assign \s5_addr_o[9]  = ~\new_[13340]_  | ~\new_[13341]_  | ~\new_[14737]_  | ~\new_[13339]_ ;
  assign \s5_addr_o[8]  = ~\new_[14739]_  | ~\new_[13342]_  | ~\new_[14738]_  | ~\new_[11397]_ ;
  assign \s5_addr_o[7]  = ~\new_[13343]_  | ~\new_[14740]_  | ~\new_[11398]_  | ~\new_[11399]_ ;
  assign \s5_addr_o[6]  = ~\new_[13346]_  | ~\new_[13348]_  | ~\new_[14741]_  | ~\new_[13344]_ ;
  assign \s5_addr_o[5]  = ~\new_[13352]_  | ~\new_[14748]_  | ~\new_[14747]_  | ~\new_[13351]_ ;
  assign \s5_addr_o[4]  = ~\new_[13356]_  | ~\new_[13358]_  | ~\new_[14753]_  | ~\new_[13354]_ ;
  assign \s5_addr_o[3]  = ~\new_[14757]_  | ~\new_[13362]_  | ~\new_[11404]_  | ~\new_[13361]_ ;
  assign \s5_addr_o[2]  = ~\new_[14760]_  | ~\new_[14761]_  | ~\new_[13365]_  | ~\new_[11406]_ ;
  assign \s5_sel_o[2]  = ~\new_[14776]_  | ~\new_[13381]_  | ~\new_[11414]_  | ~\new_[13380]_ ;
  assign \s5_sel_o[1]  = ~\new_[14781]_  | ~\new_[13382]_  | ~\new_[11415]_  | ~\new_[14780]_ ;
  assign \s5_sel_o[0]  = ~\new_[14782]_  | ~\new_[13385]_  | ~\new_[11416]_  | ~\new_[13383]_ ;
  assign s5_we_o = ~\new_[14789]_  | ~\new_[13389]_  | ~\new_[11418]_  | ~\new_[13387]_ ;
  assign \new_[8219]_  = ~\new_[10306]_  & ~\new_[12824]_ ;
  assign \new_[8220]_  = ~\new_[15340]_  & ~\new_[10512]_ ;
  assign \new_[8221]_  = ~\new_[10425]_  | ~\new_[28291]_ ;
  assign s10_cyc_o = ~n7659;
  assign \new_[8223]_  = ~\new_[10671]_  & ~\new_[12188]_ ;
  assign \new_[8224]_  = ~\new_[10515]_  & ~\new_[12536]_ ;
  assign \new_[8225]_  = ~\new_[15366]_  & ~\new_[10518]_ ;
  assign n7524 = (~\new_[12295]_  & ~rst_i) | (~\new_[30669]_  & ~\new_[31698]_ );
  assign n7539 = ~\new_[13704]_  & ~\new_[10475]_ ;
  assign \s10_data_o[30]  = ~\new_[13700]_  | ~\new_[14971]_  | ~\new_[16343]_  | ~\new_[12092]_ ;
  assign \s10_data_o[29]  = ~\new_[14973]_  | ~\new_[14975]_  | ~\new_[13701]_  | ~\new_[12095]_ ;
  assign \s10_data_o[28]  = ~\new_[13706]_  | ~\new_[14976]_  | ~\new_[16344]_  | ~\new_[12097]_ ;
  assign \s10_data_o[27]  = ~\new_[16345]_  | ~\new_[14977]_  | ~\new_[13707]_  | ~\new_[12100]_ ;
  assign \s10_data_o[24]  = ~\new_[13713]_  | ~\new_[14981]_  | ~\new_[12109]_  | ~\new_[13712]_ ;
  assign \s10_data_o[23]  = ~\new_[14982]_  | ~\new_[14983]_  | ~\new_[13714]_  | ~\new_[12113]_ ;
  assign \s10_data_o[21]  = ~\new_[15946]_  | ~\new_[14985]_  | ~\new_[13716]_  | ~\new_[12117]_ ;
  assign \new_[8235]_  = ~\new_[10338]_  & ~\new_[12837]_ ;
  assign \s10_data_o[20]  = ~\new_[14986]_  | ~\new_[14987]_  | ~\new_[13717]_  | ~\new_[12119]_ ;
  assign \s10_data_o[19]  = ~\new_[14988]_  | ~\new_[14989]_  | ~\new_[12121]_  | ~\new_[12122]_ ;
  assign \s10_data_o[17]  = ~\new_[13721]_  | ~\new_[14821]_  | ~\new_[12124]_  | ~\new_[12125]_ ;
  assign \s10_data_o[16]  = ~\new_[13723]_  | ~\new_[14994]_  | ~\new_[12126]_  | ~\new_[13722]_ ;
  assign \s10_data_o[13]  = ~\new_[14995]_  | ~\new_[13728]_  | ~\new_[12132]_  | ~\new_[14996]_ ;
  assign \s10_data_o[12]  = ~\new_[16351]_  | ~\new_[14998]_  | ~\new_[13729]_  | ~\new_[12136]_ ;
  assign \s10_data_o[11]  = ~\new_[15000]_  | ~\new_[15001]_  | ~\new_[13733]_  | ~\new_[12140]_ ;
  assign \s10_data_o[10]  = ~\new_[15002]_  | ~\new_[15003]_  | ~\new_[13735]_  | ~\new_[12144]_ ;
  assign \s10_data_o[8]  = ~\new_[15006]_  | ~\new_[15007]_  | ~\new_[13740]_  | ~\new_[12151]_ ;
  assign \s10_data_o[5]  = ~\new_[13747]_  | ~\new_[15012]_  | ~\new_[12159]_  | ~\new_[12160]_ ;
  assign \s10_addr_o[31]  = ~\new_[15018]_  | ~\new_[15019]_  | ~\new_[16363]_  | ~\new_[12178]_ ;
  assign \s10_addr_o[29]  = ~\new_[15021]_  | ~\new_[15022]_  | ~\new_[13764]_  | ~\new_[12187]_ ;
  assign \s10_addr_o[22]  = ~\new_[15027]_  | ~\new_[15029]_  | ~\new_[13658]_  | ~\new_[12213]_ ;
  assign \s10_addr_o[21]  = ~\new_[13211]_  | ~\new_[15031]_  | ~\new_[13773]_  | ~\new_[12217]_ ;
  assign \s10_addr_o[20]  = ~\new_[15032]_  | ~\new_[15033]_  | ~\new_[13774]_  | ~\new_[12222]_ ;
  assign \s10_addr_o[19]  = ~\new_[13777]_  | ~\new_[15035]_  | ~\new_[16370]_  | ~\new_[12226]_ ;
  assign \s10_addr_o[18]  = ~\new_[13780]_  | ~\new_[15037]_  | ~\new_[11314]_  | ~\new_[13779]_ ;
  assign \s10_addr_o[17]  = ~\new_[15038]_  | ~\new_[15040]_  | ~\new_[13782]_  | ~\new_[12231]_ ;
  assign \s10_addr_o[16]  = ~\new_[13785]_  | ~\new_[15042]_  | ~\new_[15041]_  | ~\new_[12236]_ ;
  assign \s10_addr_o[15]  = ~\new_[15044]_  | ~\new_[15045]_  | ~\new_[13786]_  | ~\new_[12239]_ ;
  assign \s10_addr_o[13]  = ~\new_[13791]_  | ~\new_[15050]_  | ~\new_[15048]_  | ~\new_[13792]_ ;
  assign \s10_addr_o[10]  = ~\new_[15058]_  | ~\new_[15060]_  | ~\new_[12250]_  | ~\new_[12251]_ ;
  assign \s10_addr_o[9]  = ~\new_[15061]_  | ~\new_[15063]_  | ~\new_[12253]_  | ~\new_[12254]_ ;
  assign \new_[8259]_  = ~\new_[10520]_  & ~\new_[10682]_ ;
  assign \s10_addr_o[5]  = ~\new_[15078]_  | ~\new_[15110]_  | ~\new_[13811]_  | ~\new_[12263]_ ;
  assign \s10_addr_o[4]  = ~\new_[16380]_  | ~\new_[15080]_  | ~\new_[13813]_  | ~\new_[12268]_ ;
  assign \s10_addr_o[3]  = ~\new_[13816]_  | ~\new_[15085]_  | ~\new_[12269]_  | ~\new_[15082]_ ;
  assign \s10_addr_o[0]  = ~\new_[15097]_  | ~\new_[15098]_  | ~\new_[13824]_  | ~\new_[12278]_ ;
  assign \s10_sel_o[2]  = ~\new_[15105]_  | ~\new_[15106]_  | ~\new_[13829]_  | ~\new_[12281]_ ;
  assign \s10_sel_o[1]  = ~\new_[15108]_  | ~\new_[14866]_  | ~\new_[13831]_  | ~\new_[12285]_ ;
  assign \s11_data_o[18]  = ~\new_[15383]_  | ~\new_[13872]_  | ~\new_[12345]_  | ~\new_[12346]_ ;
  assign \s11_data_o[8]  = ~\new_[13904]_  | ~\new_[15180]_  | ~\new_[12367]_  | ~\new_[12369]_ ;
  assign \new_[8268]_  = ~\new_[12843]_  & ~\new_[10347]_ ;
  assign \s11_addr_o[23]  = ~\new_[13953]_  | ~\new_[15232]_  | ~\new_[11163]_  | ~\new_[12411]_ ;
  assign \s11_addr_o[20]  = ~\new_[15241]_  | ~\new_[13962]_  | ~\new_[12417]_  | ~\new_[12420]_ ;
  assign \s11_addr_o[13]  = ~\new_[13129]_  | ~\new_[15260]_  | ~\new_[12441]_  | ~\new_[12442]_ ;
  assign \s11_addr_o[11]  = ~\new_[14503]_  | ~\new_[13979]_  | ~\new_[12445]_  | ~\new_[12446]_ ;
  assign \s11_addr_o[9]  = ~\new_[15270]_  | ~\new_[13981]_  | ~\new_[12451]_  | ~\new_[12452]_ ;
  assign \s11_addr_o[6]  = ~\new_[13985]_  | ~\new_[15274]_  | ~\new_[12460]_  | ~\new_[12461]_ ;
  assign \s11_sel_o[3]  = ~\new_[13112]_  | ~\new_[15288]_  | ~\new_[11162]_  | ~\new_[12483]_ ;
  assign n7529 = (~\new_[12304]_  & ~rst_i) | (~\new_[31151]_  & ~\new_[31678]_ );
  assign s1_cyc_o = ~n7654;
  assign n7544 = ~\new_[12129]_  & ~\new_[10487]_ ;
  assign \new_[8279]_  = ~\new_[10359]_  & ~\new_[12848]_ ;
  assign n7534 = (~\new_[12317]_  & ~rst_i) | (~\new_[31028]_  & ~\new_[31804]_ );
  assign \new_[8281]_  = ~\new_[13685]_  & ~\new_[10229]_ ;
  assign \new_[8282]_  = ~\new_[13686]_  & ~\new_[10497]_ ;
  assign \new_[8283]_  = ~\new_[12071]_  & ~\new_[10248]_ ;
  assign \new_[8284]_  = ~\new_[13689]_  & ~\new_[10262]_ ;
  assign \new_[8285]_  = ~\new_[13691]_  & ~\new_[10507]_ ;
  assign \new_[8286]_  = ~\new_[10469]_  & ~\new_[11940]_ ;
  assign \new_[8287]_  = ~\new_[13694]_  & ~\new_[10511]_ ;
  assign \new_[8288]_  = ~\new_[12087]_  & ~\new_[10311]_ ;
  assign \new_[8289]_  = ~\new_[13703]_  & ~\new_[10334]_ ;
  assign \new_[8290]_  = ~\new_[10477]_  & ~\new_[10344]_ ;
  assign \new_[8291]_  = ~\new_[10354]_  & ~\new_[10522]_ ;
  assign \new_[8292]_  = ~\new_[28310]_  & (~\new_[12216]_  | ~\new_[21360]_ );
  assign \new_[8293]_  = ~\new_[27797]_  & (~\new_[12324]_  | ~\new_[22698]_ );
  assign \new_[8294]_  = ~\new_[10392]_  & (~\new_[13190]_  | ~\new_[29549]_ );
  assign \new_[8295]_  = ~\new_[28327]_  & (~\new_[12612]_  | ~\new_[26822]_ );
  assign \new_[8296]_  = ~\new_[10394]_  & (~\new_[14542]_  | ~\new_[26466]_ );
  assign \new_[8297]_  = ~\new_[28038]_  & (~\new_[12218]_  | ~\new_[22711]_ );
  assign \new_[8298]_  = ~\new_[10395]_  & (~\new_[13193]_  | ~\new_[27816]_ );
  assign \new_[8299]_  = ~\new_[28068]_  & (~\new_[12220]_  | ~\new_[24236]_ );
  assign \new_[8300]_  = ~\new_[28354]_  & (~\new_[12616]_  | ~\new_[27758]_ );
  assign \new_[8301]_  = ~\new_[28729]_  & (~\new_[12221]_  | ~\new_[22796]_ );
  assign \new_[8302]_  = ~\new_[10398]_  & (~\new_[13195]_  | ~\new_[29084]_ );
  assign \new_[8303]_  = ~\new_[28603]_  & (~\new_[12619]_  | ~\new_[26735]_ );
  assign \new_[8304]_  = ~\new_[12067]_  & ~\new_[10236]_ ;
  assign \new_[8305]_  = ~\new_[10400]_  & (~\new_[13197]_  | ~\new_[28623]_ );
  assign \new_[8306]_  = ~\new_[28617]_  & (~\new_[12223]_  | ~\new_[22797]_ );
  assign \new_[8307]_  = ~\new_[27938]_  & (~\new_[12352]_  | ~\new_[21452]_ );
  assign \new_[8308]_  = ~\new_[10402]_  & (~\new_[13198]_  | ~\new_[29161]_ );
  assign \new_[8309]_  = ~\new_[29847]_  & (~\new_[12622]_  | ~\new_[27608]_ );
  assign \new_[8310]_  = ~\new_[28925]_  & (~\new_[12225]_  | ~\new_[22655]_ );
  assign \new_[8311]_  = ~\new_[10406]_  & (~\new_[13201]_  | ~\new_[29993]_ );
  assign \new_[8312]_  = ~\new_[28613]_  & (~\new_[12627]_  | ~\new_[27950]_ );
  assign \new_[8313]_  = ~\new_[20391]_  | ~\new_[10137]_ ;
  assign \new_[8314]_  = ~\new_[28018]_  & (~\new_[12228]_  | ~\new_[22563]_ );
  assign \new_[8315]_  = ~\new_[10410]_  & (~\new_[13203]_  | ~\new_[29580]_ );
  assign \new_[8316]_  = ~\new_[28607]_  & (~\new_[12631]_  | ~\new_[26741]_ );
  assign \new_[8317]_  = ~\new_[20379]_  | ~\new_[10141]_ ;
  assign \new_[8318]_  = ~\new_[29321]_  & (~\new_[12229]_  | ~\new_[20425]_ );
  assign \new_[8319]_  = ~\new_[27784]_  & (~\new_[12374]_  | ~\new_[20421]_ );
  assign \new_[8320]_  = ~\new_[10412]_  & (~\new_[13687]_  | ~\new_[28843]_ );
  assign \new_[8321]_  = ~\new_[30056]_  & (~\new_[12634]_  | ~\new_[27621]_ );
  assign \new_[8322]_  = ~\new_[10416]_  & (~\new_[13613]_  | ~\new_[24482]_ );
  assign \new_[8323]_  = ~\new_[28387]_  & (~\new_[12230]_  | ~\new_[22809]_ );
  assign \new_[8324]_  = ~\new_[10417]_  & (~\new_[13600]_  | ~\new_[29731]_ );
  assign \new_[8325]_  = ~\new_[28325]_  & (~\new_[12638]_  | ~\new_[27613]_ );
  assign \new_[8326]_  = ~\new_[28316]_  & (~\new_[12642]_  | ~\new_[27641]_ );
  assign \new_[8327]_  = ~\new_[13695]_  & ~\new_[10308]_ ;
  assign \new_[8328]_  = ~\new_[28292]_  & (~\new_[12234]_  | ~\new_[21403]_ );
  assign \new_[8329]_  = ~\new_[27804]_  & (~\new_[12395]_  | ~\new_[21342]_ );
  assign \new_[8330]_  = ~\new_[28060]_  & (~\new_[12646]_  | ~\new_[27632]_ );
  assign \new_[8331]_  = ~\new_[27788]_  & (~\new_[12700]_  | ~\new_[28139]_ );
  assign \new_[8332]_  = ~\new_[10426]_  & (~\new_[14550]_  | ~\new_[27809]_ );
  assign \new_[8333]_  = ~\new_[29343]_  & (~\new_[12237]_  | ~\new_[22700]_ );
  assign \new_[8334]_  = ~\new_[28608]_  & (~\new_[12402]_  | ~\new_[22524]_ );
  assign \new_[8335]_  = ~\new_[10427]_  & (~\new_[14468]_  | ~\new_[30288]_ );
  assign \new_[8336]_  = ~\new_[10429]_  & (~\new_[15749]_  | ~\new_[29310]_ );
  assign \new_[8337]_  = ~\new_[28087]_  & (~\new_[12651]_  | ~\new_[28429]_ );
  assign \new_[8338]_  = ~\new_[28657]_  & (~\new_[12238]_  | ~\new_[22079]_ );
  assign \new_[8339]_  = ~\new_[10431]_  & (~\new_[14208]_  | ~\new_[27798]_ );
  assign \new_[8340]_  = ~\new_[28620]_  & (~\new_[12653]_  | ~\new_[27644]_ );
  assign \new_[8341]_  = ~\new_[13705]_  & ~\new_[10341]_ ;
  assign \new_[8342]_  = ~\new_[28805]_  & (~\new_[12240]_  | ~\new_[21443]_ );
  assign \new_[8343]_  = ~\new_[28019]_  & (~\new_[12425]_  | ~\new_[21439]_ );
  assign \new_[8344]_  = ~\new_[28599]_  & (~\new_[12659]_  | ~\new_[26874]_ );
  assign \new_[8345]_  = ~\new_[20371]_  | ~\new_[10176]_ ;
  assign \new_[8346]_  = ~\new_[28625]_  & (~\new_[12430]_  | ~\new_[20439]_ );
  assign \new_[8347]_  = ~\new_[10435]_  & (~\new_[13575]_  | ~\new_[30190]_ );
  assign \new_[8348]_  = ~\new_[30165]_  & (~\new_[12662]_  | ~\new_[26704]_ );
  assign \new_[8349]_  = ~\new_[20387]_  | ~\new_[10187]_ ;
  assign \new_[8350]_  = ~\new_[28755]_  & (~\new_[12244]_  | ~\new_[22840]_ );
  assign \new_[8351]_  = ~\new_[10437]_  & (~\new_[13531]_  | ~\new_[27777]_ );
  assign \new_[8352]_  = ~\new_[29533]_  & (~\new_[12665]_  | ~\new_[28074]_ );
  assign \new_[8353]_  = ~\new_[28022]_  & (~\new_[12795]_  | ~\new_[26795]_ );
  assign \new_[8354]_  = ~\new_[29982]_  & (~\new_[12347]_  | ~\new_[22862]_ );
  assign \new_[8355]_  = ~\new_[30119]_  & (~\new_[12391]_  | ~\new_[22984]_ );
  assign \new_[8356]_  = ~\new_[28720]_  & (~\new_[12414]_  | ~\new_[23098]_ );
  assign \new_[8357]_  = ~\new_[27873]_  & (~\new_[12498]_  | ~\new_[23261]_ );
  assign \new_[8358]_  = ~\new_[26533]_  & (~\new_[12364]_  | ~\new_[20429]_ );
  assign \new_[8359]_  = ~\new_[27363]_  & (~\new_[12797]_  | ~\new_[26362]_ );
  assign \new_[8360]_  = ~\new_[27866]_  & (~\new_[12361]_  | ~\new_[23025]_ );
  assign \new_[8361]_  = ~\new_[28841]_  & (~\new_[12443]_  | ~\new_[23228]_ );
  assign \new_[8362]_  = ~\new_[27823]_  & (~\new_[12453]_  | ~\new_[21491]_ );
  assign \new_[8363]_  = ~\new_[26482]_  & (~\new_[12454]_  | ~\new_[21616]_ );
  assign \new_[8364]_  = ~\new_[27890]_  & (~\new_[12463]_  | ~\new_[21594]_ );
  assign \new_[8365]_  = ~\new_[26460]_  & (~\new_[12464]_  | ~\new_[22986]_ );
  assign \new_[8366]_  = ~\new_[27977]_  & (~\new_[12465]_  | ~\new_[27982]_ );
  assign \new_[8367]_  = ~\new_[27906]_  & (~\new_[12474]_  | ~\new_[21113]_ );
  assign \new_[8368]_  = ~\new_[26452]_  & (~\new_[12475]_  | ~\new_[22946]_ );
  assign \new_[8369]_  = ~\new_[28922]_  & (~\new_[12476]_  | ~\new_[29352]_ );
  assign \new_[8370]_  = ~\new_[29066]_  | (~\new_[12783]_  & ~\new_[24812]_ );
  assign \new_[8371]_  = ~\new_[29599]_  & (~\new_[12486]_  | ~\new_[19425]_ );
  assign \new_[8372]_  = ~\new_[28175]_  & (~\new_[12503]_  | ~\new_[23940]_ );
  assign \new_[8373]_  = ~\new_[28779]_  & (~\new_[12507]_  | ~\new_[23330]_ );
  assign \new_[8374]_  = ~\new_[29196]_  | (~\new_[12814]_  & ~\new_[26204]_ );
  assign \new_[8375]_  = ~\new_[26964]_  & (~\new_[12510]_  | ~\new_[19442]_ );
  assign \new_[8376]_  = ~\new_[24647]_  & (~\new_[12511]_  | ~\new_[28277]_ );
  assign \new_[8377]_  = ~\new_[27839]_  & (~\new_[12516]_  | ~\new_[19438]_ );
  assign \new_[8378]_  = ~\new_[26457]_  & (~\new_[12517]_  | ~\new_[22889]_ );
  assign \new_[8379]_  = ~\new_[27829]_  & (~\new_[12520]_  | ~\new_[19709]_ );
  assign \new_[8380]_  = ~\new_[24598]_  & (~\new_[12521]_  | ~\new_[23003]_ );
  assign \new_[8381]_  = ~\new_[28290]_  & (~\new_[12522]_  | ~\new_[22923]_ );
  assign \new_[8382]_  = ~\new_[29675]_  & (~\new_[12523]_  | ~\new_[29209]_ );
  assign \new_[8383]_  = ~\new_[27502]_  & (~\new_[12528]_  | ~\new_[20447]_ );
  assign \new_[8384]_  = ~\new_[26510]_  & (~\new_[12529]_  | ~\new_[23033]_ );
  assign \new_[8385]_  = ~\new_[28085]_  & (~\new_[12538]_  | ~\new_[24299]_ );
  assign \new_[8386]_  = ~\new_[27931]_  & (~\new_[12540]_  | ~\new_[19449]_ );
  assign \new_[8387]_  = ~\new_[24538]_  & (~\new_[12541]_  | ~\new_[22910]_ );
  assign \new_[8388]_  = ~\new_[26501]_  & (~\new_[12542]_  | ~\new_[22970]_ );
  assign \new_[8389]_  = ~\new_[28084]_  & (~\new_[12546]_  | ~\new_[24277]_ );
  assign \new_[8390]_  = ~\new_[29135]_  & (~\new_[12550]_  | ~\new_[24369]_ );
  assign \new_[8391]_  = ~\new_[31995]_ ;
  assign \new_[8392]_  = ~\new_[28319]_  & (~\new_[12716]_  | ~\new_[21436]_ );
  assign \new_[8393]_  = ~\new_[27823]_  & (~\new_[12559]_  | ~\new_[21766]_ );
  assign \new_[8394]_  = ~\new_[28263]_  & (~\new_[12561]_  | ~\new_[19423]_ );
  assign \new_[8395]_  = ~\new_[28716]_  & (~\new_[12721]_  | ~\new_[20433]_ );
  assign \new_[8396]_  = ~\new_[27890]_  & (~\new_[12562]_  | ~\new_[24326]_ );
  assign \new_[8397]_  = ~\new_[28356]_  & (~\new_[12563]_  | ~\new_[21505]_ );
  assign \new_[8398]_  = ~\new_[29679]_  & (~\new_[12723]_  | ~\new_[21353]_ );
  assign \new_[8399]_  = ~\new_[27906]_  & (~\new_[12565]_  | ~\new_[22893]_ );
  assign \new_[8400]_  = ~\new_[28913]_  & (~\new_[12567]_  | ~\new_[19426]_ );
  assign \new_[8401]_  = ~\new_[28715]_  & (~\new_[12724]_  | ~\new_[21373]_ );
  assign \new_[8402]_  = ~\new_[28056]_  & (~\new_[12726]_  | ~\new_[26167]_ );
  assign \new_[8403]_  = ~\new_[29599]_  & (~\new_[12568]_  | ~\new_[21539]_ );
  assign \new_[8404]_  = ~\new_[27857]_  & (~\new_[12570]_  | ~\new_[20524]_ );
  assign \new_[8405]_  = ~\new_[28975]_  & (~\new_[12571]_  | ~\new_[22924]_ );
  assign \new_[8406]_  = ~\new_[28059]_  & (~\new_[12739]_  | ~\new_[20422]_ );
  assign \new_[8407]_  = ~\new_[8863]_ ;
  assign \new_[8408]_  = ~\new_[8863]_ ;
  assign \new_[8409]_  = ~\new_[26964]_  & (~\new_[12573]_  | ~\new_[21552]_ );
  assign \new_[8410]_  = ~\new_[26634]_  & (~\new_[12576]_  | ~\new_[20472]_ );
  assign \new_[8411]_  = ~\new_[29274]_  & (~\new_[12743]_  | ~\new_[22649]_ );
  assign \new_[8412]_  = ~\new_[27839]_  & (~\new_[12577]_  | ~\new_[21356]_ );
  assign \new_[8413]_  = ~\new_[27829]_  & (~\new_[12579]_  | ~\new_[21759]_ );
  assign \new_[8414]_  = ~\new_[29407]_  & (~\new_[12581]_  | ~\new_[20477]_ );
  assign \new_[8415]_  = ~\new_[28487]_  & (~\new_[12747]_  | ~\new_[22793]_ );
  assign \new_[8416]_  = ~\new_[28557]_  & (~\new_[12748]_  | ~\new_[20415]_ );
  assign \new_[8417]_  = ~\new_[27502]_  & (~\new_[12583]_  | ~\new_[22914]_ );
  assign \new_[8418]_  = ~\new_[28628]_  & (~\new_[12584]_  | ~\new_[29740]_ );
  assign \new_[8419]_  = ~\new_[29313]_  & (~\new_[12585]_  | ~\new_[20503]_ );
  assign \new_[8420]_  = ~\new_[29361]_  & (~\new_[12750]_  | ~\new_[20414]_ );
  assign \new_[8421]_  = ~\new_[28667]_  & (~\new_[12751]_  | ~\new_[23721]_ );
  assign \new_[8422]_  = ~\new_[27931]_  & (~\new_[12587]_  | ~\new_[21534]_ );
  assign \new_[8423]_  = ~\new_[26649]_  & (~\new_[12589]_  | ~\new_[19433]_ );
  assign \new_[8424]_  = ~\new_[28006]_  & (~\new_[12590]_  | ~\new_[21521]_ );
  assign \new_[8425]_  = ~\new_[29148]_  & (~\new_[12760]_  | ~\new_[21416]_ );
  assign \new_[8426]_  = ~\new_[28929]_  & (~\new_[12762]_  | ~\new_[22821]_ );
  assign \new_[8427]_  = ~\new_[29752]_  & (~\new_[12592]_  | ~\new_[22922]_ );
  assign \new_[8428]_  = ~\new_[26503]_  & (~\new_[12765]_  | ~\new_[21352]_ );
  assign \new_[8429]_  = ~\new_[27878]_  & (~\new_[12322]_  | ~\new_[20440]_ );
  assign \new_[8430]_  = ~\new_[26966]_  & (~\new_[12334]_  | ~\new_[22782]_ );
  assign \new_[8431]_  = ~\new_[27975]_  & (~\new_[12336]_  | ~\new_[22779]_ );
  assign \new_[8432]_  = ~\new_[28552]_  & (~\new_[12342]_  | ~\new_[19410]_ );
  assign \new_[8433]_  = ~\new_[27900]_  & (~\new_[12349]_  | ~\new_[19405]_ );
  assign \new_[8434]_  = ~\new_[27995]_  & (~\new_[12355]_  | ~\new_[19412]_ );
  assign \new_[8435]_  = ~\new_[29087]_  & (~\new_[12356]_  | ~\new_[22757]_ );
  assign \new_[8436]_  = ~\new_[26587]_  & (~\new_[12362]_  | ~\new_[24208]_ );
  assign \new_[8437]_  = ~\new_[28931]_  & (~\new_[12372]_  | ~\new_[19414]_ );
  assign \new_[8438]_  = ~\new_[26683]_  & (~\new_[12381]_  | ~\new_[19415]_ );
  assign \new_[8439]_  = ~\new_[29666]_  & (~\new_[12383]_  | ~\new_[24206]_ );
  assign \new_[8440]_  = ~\new_[28036]_  & (~\new_[12385]_  | ~\new_[18422]_ );
  assign \new_[8441]_  = ~\new_[27891]_  & (~\new_[12397]_  | ~\new_[22788]_ );
  assign \new_[8442]_  = ~\new_[28611]_  & (~\new_[12405]_  | ~\new_[21448]_ );
  assign \new_[8443]_  = ~\new_[28635]_  & (~\new_[12418]_  | ~\new_[21441]_ );
  assign \new_[8444]_  = ~\new_[27858]_  & (~\new_[12422]_  | ~\new_[22800]_ );
  assign \new_[8445]_  = (~\new_[12548]_  | ~\new_[29856]_ ) & (~\new_[26157]_  | ~\new_[29856]_ );
  assign \new_[8446]_  = (~\new_[12552]_  | ~\new_[27902]_ ) & (~\new_[22696]_  | ~\new_[27902]_ );
  assign \new_[8447]_  = ~\new_[8935]_ ;
  assign \s11_addr_o[21]  = ~\new_[15239]_  | ~\new_[13437]_  | ~\new_[12413]_  | ~\new_[12415]_ ;
  assign \new_[8449]_  = ~\new_[10654]_  & ~\new_[11939]_ ;
  assign \new_[8450]_  = ~\new_[10734]_  | ~\new_[26839]_ ;
  assign \new_[8451]_  = ~\new_[10611]_  | ~\new_[28532]_ ;
  assign \new_[8452]_  = ~\new_[10738]_  | ~\new_[28541]_ ;
  assign \new_[8453]_  = ~\new_[10741]_  | ~\new_[27602]_ ;
  assign \new_[8454]_  = ~\new_[10744]_  | ~\new_[28510]_ ;
  assign \new_[8455]_  = ~\new_[10753]_  | ~\new_[28554]_ ;
  assign \new_[8456]_  = ~\new_[10755]_  | ~\new_[28186]_ ;
  assign \new_[8457]_  = ~\new_[10757]_  | ~\new_[28384]_ ;
  assign \new_[8458]_  = ~\new_[10758]_  | ~\new_[28291]_ ;
  assign \new_[8459]_  = ~\new_[10767]_  | ~\new_[28294]_ ;
  assign n7559 = (~\new_[13048]_  & ~rst_i) | (~\new_[30917]_  & ~\new_[31564]_ );
  assign n7564 = (~\new_[13053]_  & ~rst_i) | (~\new_[30928]_  & ~\new_[31846]_ );
  assign n7569 = (~\new_[13054]_  & ~rst_i) | (~\new_[30614]_  & ~\new_[31810]_ );
  assign n7574 = (~\new_[13075]_  & ~rst_i) | (~\new_[31040]_  & ~\new_[31718]_ );
  assign \new_[8464]_  = ~\new_[29114]_  & (~\new_[13006]_  | ~\new_[22680]_ );
  assign \new_[8465]_  = ~\new_[28653]_  & (~\new_[13011]_  | ~\new_[22716]_ );
  assign n7579 = (~\new_[13087]_  & ~rst_i) | (~\new_[30880]_  & ~\new_[31597]_ );
  assign n7584 = (~\new_[13095]_  & ~rst_i) | (~\new_[30817]_  & ~\new_[31575]_ );
  assign \new_[8468]_  = ~\new_[21322]_  | ~\new_[10543]_ ;
  assign \new_[8469]_  = ~\new_[10526]_  & ~\new_[15398]_ ;
  assign \new_[8470]_  = ~\new_[28755]_  & (~\new_[13033]_  | ~\new_[22842]_ );
  assign \new_[8471]_  = ~\new_[14391]_  | ~\new_[14429]_  | ~\new_[11100]_  | ~\new_[14427]_ ;
  assign \new_[8472]_  = ~\new_[13114]_  | ~\new_[14510]_  | ~\new_[14509]_  | ~\new_[13113]_ ;
  assign \new_[8473]_  = ~\new_[13118]_  | ~\new_[14511]_  | ~\new_[15901]_  | ~\new_[15902]_ ;
  assign \new_[8474]_  = ~\new_[9317]_ ;
  assign \new_[8475]_  = ~\new_[22505]_  | ~\new_[13565]_  | ~\new_[21258]_  | ~\new_[11854]_ ;
  assign \new_[8476]_  = ~\new_[9770]_  & ~\new_[13654]_ ;
  assign \new_[8477]_  = (~\new_[11834]_  | ~\new_[26766]_ ) & (~\new_[13573]_  | ~\new_[28051]_ );
  assign \new_[8478]_  = (~\new_[11835]_  | ~\new_[28701]_ ) & (~\new_[13574]_  | ~\new_[28314]_ );
  assign \new_[8479]_  = (~\new_[11839]_  | ~\new_[28630]_ ) & (~\new_[13578]_  | ~\new_[28323]_ );
  assign \new_[8480]_  = (~\new_[11840]_  | ~\new_[30077]_ ) & (~\new_[14915]_  | ~\new_[29423]_ );
  assign \new_[8481]_  = (~\new_[11843]_  | ~\new_[28126]_ ) & (~\new_[13580]_  | ~\new_[26608]_ );
  assign \new_[8482]_  = (~\new_[11844]_  | ~\new_[29658]_ ) & (~\new_[14917]_  | ~\new_[28764]_ );
  assign \new_[8483]_  = (~\new_[11849]_  | ~\new_[29273]_ ) & (~\new_[11848]_  | ~\new_[29416]_ );
  assign \new_[8484]_  = (~\new_[11851]_  | ~\new_[28879]_ ) & (~\new_[13582]_  | ~\new_[29713]_ );
  assign \new_[8485]_  = (~\new_[11863]_  | ~\new_[29237]_ ) & (~\new_[13586]_  | ~\new_[28008]_ );
  assign \new_[8486]_  = (~\new_[11867]_  | ~\new_[28758]_ ) & (~\new_[13587]_  | ~\new_[27957]_ );
  assign \new_[8487]_  = (~\new_[11869]_  | ~\new_[29678]_ ) & (~\new_[13591]_  | ~\new_[29140]_ );
  assign \new_[8488]_  = (~\new_[11871]_  | ~\new_[29586]_ ) & (~\new_[14921]_  | ~\new_[29059]_ );
  assign \new_[8489]_  = (~\new_[11875]_  | ~\new_[29279]_ ) & (~\new_[13594]_  | ~\new_[28295]_ );
  assign \new_[8490]_  = (~\new_[11876]_  | ~\new_[29301]_ ) & (~\new_[14922]_  | ~\new_[29345]_ );
  assign \new_[8491]_  = (~\new_[11880]_  | ~\new_[29187]_ ) & (~\new_[11879]_  | ~\new_[29703]_ );
  assign \new_[8492]_  = (~\new_[11884]_  | ~\new_[28261]_ ) & (~\new_[14925]_  | ~\new_[28757]_ );
  assign \new_[8493]_  = (~\new_[11887]_  | ~\new_[28030]_ ) & (~\new_[11885]_  | ~\new_[28237]_ );
  assign \new_[8494]_  = (~\new_[11889]_  | ~\new_[29041]_ ) & (~\new_[13602]_  | ~\new_[29010]_ );
  assign \new_[8495]_  = (~\new_[11894]_  | ~\new_[26639]_ ) & (~\new_[13603]_  | ~\new_[28588]_ );
  assign \new_[8496]_  = (~\new_[11898]_  | ~\new_[28077]_ ) & (~\new_[13610]_  | ~\new_[28364]_ );
  assign \new_[8497]_  = (~\new_[11902]_  | ~\new_[27000]_ ) & (~\new_[13614]_  | ~\new_[28320]_ );
  assign \new_[8498]_  = ~\new_[11552]_  & ~\new_[9955]_ ;
  assign \new_[8499]_  = ~\new_[9957]_  & ~\new_[11554]_ ;
  assign n7509 = ~\new_[30310]_  | (~\new_[12098]_  & ~rst_i);
  assign \new_[8501]_  = ~\new_[9968]_  & ~\new_[11579]_ ;
  assign \new_[8502]_  = ~\new_[9705]_  & ~\new_[13652]_ ;
  assign n7554 = ~\new_[10463]_  & ~\new_[10464]_ ;
  assign \new_[8504]_  = ~\new_[9899]_  & ~\new_[9973]_ ;
  assign \new_[8505]_  = ~\new_[11629]_  & ~\new_[9994]_ ;
  assign \new_[8506]_  = ~\new_[10007]_  & ~\new_[11654]_ ;
  assign \new_[8507]_  = ~\new_[10015]_  & ~\new_[11674]_ ;
  assign \new_[8508]_  = ~\new_[11420]_  & (~\new_[11831]_  | ~\new_[27903]_ );
  assign \new_[8509]_  = ~\new_[11383]_  & ~\new_[9866]_ ;
  assign \new_[8510]_  = (~\new_[13617]_  | ~\new_[26610]_ ) & (~\new_[11909]_  | ~\new_[28723]_ );
  assign \new_[8511]_  = ~\new_[9783]_  & ~\new_[11567]_ ;
  assign \new_[8512]_  = ~\new_[9785]_  & (~\new_[11838]_  | ~\new_[24582]_ );
  assign \new_[8513]_  = ~\new_[9699]_  & (~\new_[11841]_  | ~\new_[26635]_ );
  assign \new_[8514]_  = ~\new_[13345]_  | ~\new_[14744]_  | ~\new_[14742]_  | ~\new_[14743]_ ;
  assign \new_[8515]_  = (~\new_[11925]_  | ~\new_[27884]_ ) & (~\new_[13624]_  | ~\new_[26608]_ );
  assign \new_[8516]_  = ~\new_[13350]_  | ~\new_[16139]_  | ~\new_[13226]_  | ~\new_[16138]_ ;
  assign \new_[8517]_  = ~\new_[13227]_  | ~\new_[17861]_  | ~\new_[16019]_  | ~\new_[17017]_ ;
  assign \new_[8518]_  = ~\new_[13355]_  | ~\new_[14752]_  | ~\new_[14750]_  | ~\new_[14751]_ ;
  assign \new_[8519]_  = ~\new_[10027]_  & ~\new_[11583]_ ;
  assign \new_[8520]_  = ~\new_[11308]_  & (~\new_[11845]_  | ~\new_[23071]_ );
  assign \new_[8521]_  = ~\new_[14631]_  | ~\new_[13249]_  | ~\new_[13247]_  | ~\new_[16846]_ ;
  assign \new_[8522]_  = ~\new_[11384]_  & ~\new_[9888]_ ;
  assign \new_[8523]_  = ~\new_[14646]_  | ~\new_[13256]_  | ~\new_[16055]_  | ~\new_[14645]_ ;
  assign \new_[8524]_  = ~\new_[16058]_  | ~\new_[13261]_  | ~\new_[11316]_  | ~\new_[16057]_ ;
  assign \new_[8525]_  = ~\new_[16069]_  | ~\new_[13267]_  | ~\new_[11358]_  | ~\new_[16068]_ ;
  assign \new_[8526]_  = ~\new_[9952]_  & ~\new_[9894]_ ;
  assign \new_[8527]_  = ~\new_[9707]_  & (~\new_[11857]_  | ~\new_[27894]_ );
  assign \new_[8528]_  = ~\new_[9896]_  & ~\new_[9794]_ ;
  assign \new_[8529]_  = ~\new_[9761]_  & ~\new_[10072]_ ;
  assign \new_[8530]_  = ~\new_[9755]_  & (~\new_[13628]_  | ~\new_[28742]_ );
  assign \new_[8531]_  = ~\new_[22476]_  | ~\new_[13558]_  | ~\new_[18387]_  | ~\new_[13584]_ ;
  assign \new_[8532]_  = ~\new_[16165]_  | ~\new_[16166]_  | ~\new_[9735]_  | ~\new_[16164]_ ;
  assign \new_[8533]_  = ~\new_[9769]_  & (~\new_[11859]_  | ~\new_[28742]_ );
  assign \new_[8534]_  = ~\new_[9708]_  & ~\new_[9795]_ ;
  assign \new_[8535]_  = ~\new_[16215]_  | ~\new_[14784]_  | ~\new_[9772]_  | ~\new_[11417]_ ;
  assign \new_[8536]_  = ~\new_[11324]_  & (~\new_[11862]_  | ~\new_[24580]_ );
  assign \new_[8537]_  = ~\new_[11598]_  & ~\new_[9801]_ ;
  assign \new_[8538]_  = ~\new_[11387]_  & ~\new_[9901]_ ;
  assign \new_[8539]_  = ~\new_[16921]_  | ~\new_[13406]_  | ~\new_[16920]_  | ~\new_[16184]_ ;
  assign \new_[8540]_  = ~\new_[16096]_  | ~\new_[16190]_  | ~\new_[11369]_  | ~\new_[11430]_ ;
  assign \new_[8541]_  = ~\new_[9712]_  & ~\new_[9905]_ ;
  assign \new_[8542]_  = ~\new_[10037]_  & ~\new_[11607]_ ;
  assign \new_[8543]_  = ~\new_[13306]_  | ~\new_[16203]_  | ~\new_[14805]_  | ~\new_[14806]_ ;
  assign \new_[8544]_  = ~\new_[11390]_  & ~\new_[9907]_ ;
  assign \new_[8545]_  = ~\new_[16112]_  | ~\new_[13311]_  | ~\new_[14704]_  | ~\new_[14705]_ ;
  assign \new_[8546]_  = ~\new_[13317]_  | ~\new_[16117]_  | ~\new_[16116]_  | ~\new_[13316]_ ;
  assign \new_[8547]_  = ~\new_[13323]_  | ~\new_[14809]_  | ~\new_[13321]_  | ~\new_[16210]_ ;
  assign \new_[8548]_  = ~\new_[9721]_  & (~\new_[11878]_  | ~\new_[28746]_ );
  assign \new_[8549]_  = ~\new_[11624]_  & ~\new_[9810]_ ;
  assign \new_[8550]_  = ~\new_[11396]_  & ~\new_[9915]_ ;
  assign \new_[8551]_  = (~\new_[11944]_  | ~\new_[28665]_ ) & (~\new_[11943]_  | ~\new_[29703]_ );
  assign \new_[8552]_  = (~\new_[13640]_  | ~\new_[27828]_ ) & (~\new_[11949]_  | ~\new_[28237]_ );
  assign \new_[8553]_  = (~\new_[14950]_  | ~\new_[29339]_ ) & (~\new_[11952]_  | ~\new_[29730]_ );
  assign \new_[8554]_  = ~\new_[9733]_  & (~\new_[11892]_  | ~\new_[27934]_ );
  assign \new_[8555]_  = ~\new_[13485]_  & ~\new_[9819]_ ;
  assign \new_[8556]_  = ~\new_[11479]_  & (~\new_[11893]_  | ~\new_[28101]_ );
  assign \new_[8557]_  = ~\new_[11400]_  & ~\new_[9926]_ ;
  assign \new_[8558]_  = (~\new_[13644]_  | ~\new_[27833]_ ) & (~\new_[11957]_  | ~\new_[28588]_ );
  assign \new_[8559]_  = ~\new_[9738]_  & ~\new_[9930]_ ;
  assign \new_[8560]_  = (~\new_[13645]_  | ~\new_[27449]_ ) & (~\new_[11961]_  | ~\new_[28771]_ );
  assign \new_[8561]_  = (~\new_[13647]_  | ~\new_[27439]_ ) & (~\new_[11962]_  | ~\new_[28025]_ );
  assign \new_[8562]_  = ~\new_[10062]_  & ~\new_[9937]_ ;
  assign \new_[8563]_  = ~\new_[9745]_  & (~\new_[11896]_  | ~\new_[26637]_ );
  assign \new_[8564]_  = ~\new_[9824]_  & ~\new_[13492]_ ;
  assign \new_[8565]_  = ~\new_[11488]_  & (~\new_[11897]_  | ~\new_[27956]_ );
  assign \new_[8566]_  = ~\new_[11402]_  & ~\new_[9939]_ ;
  assign \new_[8567]_  = (~\new_[11964]_  | ~\new_[28041]_ ) & (~\new_[11963]_  | ~\new_[28364]_ );
  assign \new_[8568]_  = ~\new_[10069]_  & ~\new_[11671]_ ;
  assign \new_[8569]_  = ~\new_[11372]_  & (~\new_[11900]_  | ~\new_[26528]_ );
  assign \new_[8570]_  = ~\new_[11403]_  & ~\new_[9945]_ ;
  assign \new_[8571]_  = (~\new_[14957]_  | ~\new_[26662]_ ) & (~\new_[11968]_  | ~\new_[28343]_ );
  assign \new_[8572]_  = ~\new_[9682]_  & ~\new_[9958]_ ;
  assign \new_[8573]_  = (~\new_[13530]_  | ~\m2_data_i[15] ) & (~\new_[11613]_  | ~\m3_data_i[15] );
  assign \new_[8574]_  = (~\new_[11773]_  | ~\m6_data_i[15] ) & (~\new_[31989]_  | ~\m7_data_i[15] );
  assign \new_[8575]_  = ~\new_[9986]_  & ~\new_[9718]_ ;
  assign \new_[8576]_  = (~\new_[13530]_  | ~\m2_data_i[14] ) & (~\new_[11611]_  | ~\m3_data_i[14] );
  assign \new_[8577]_  = (~\new_[11773]_  | ~\m6_data_i[14] ) & (~\new_[11539]_  | ~\m7_data_i[14] );
  assign \new_[8578]_  = (~\new_[13530]_  | ~\m2_data_i[13] ) & (~\new_[11611]_  | ~\m3_data_i[13] );
  assign \new_[8579]_  = (~\new_[11773]_  | ~\m6_data_i[13] ) & (~\new_[31989]_  | ~\m7_data_i[13] );
  assign \new_[8580]_  = (~\new_[13530]_  | ~\m2_data_i[12] ) & (~\new_[11611]_  | ~\m3_data_i[12] );
  assign \new_[8581]_  = (~\new_[11773]_  | ~\m6_data_i[12] ) & (~\new_[11539]_  | ~\m7_data_i[12] );
  assign \new_[8582]_  = (~\new_[13530]_  | ~\m2_data_i[11] ) & (~\new_[11611]_  | ~\m3_data_i[11] );
  assign \new_[8583]_  = (~\new_[11773]_  | ~\m6_data_i[11] ) & (~\new_[31989]_  | ~\m7_data_i[11] );
  assign \new_[8584]_  = ~\new_[9752]_  & ~\new_[10016]_ ;
  assign \new_[8585]_  = (~\new_[13530]_  | ~\m2_data_i[10] ) & (~\new_[11611]_  | ~\m3_data_i[10] );
  assign \new_[8586]_  = (~\new_[11773]_  | ~\m6_data_i[10] ) & (~\new_[11539]_  | ~\m7_data_i[10] );
  assign \new_[8587]_  = ~\new_[9775]_  & ~\new_[9756]_ ;
  assign \new_[8588]_  = (~\new_[13530]_  | ~\m2_data_i[9] ) & (~\new_[11613]_  | ~\m3_data_i[9] );
  assign \new_[8589]_  = (~\new_[11773]_  | ~\m6_data_i[9] ) & (~\new_[31989]_  | ~\m7_data_i[9] );
  assign \new_[8590]_  = (~\new_[13530]_  | ~\m2_data_i[8] ) & (~\new_[11613]_  | ~\m3_data_i[8] );
  assign \new_[8591]_  = (~\new_[11773]_  | ~\m6_data_i[8] ) & (~\new_[11539]_  | ~\m7_data_i[8] );
  assign \new_[8592]_  = ~\new_[10245]_  & ~\new_[10026]_ ;
  assign \new_[8593]_  = (~\new_[13530]_  | ~\m2_data_i[7] ) & (~\new_[11611]_  | ~\m3_data_i[7] );
  assign \new_[8594]_  = (~\new_[11773]_  | ~\m6_data_i[7] ) & (~\new_[11539]_  | ~\m7_data_i[7] );
  assign \new_[8595]_  = (~\new_[13530]_  | ~\m2_data_i[6] ) & (~\new_[11611]_  | ~\m3_data_i[6] );
  assign \new_[8596]_  = (~\new_[11773]_  | ~\m6_data_i[6] ) & (~\new_[11539]_  | ~\m7_data_i[6] );
  assign \new_[8597]_  = (~\new_[11773]_  | ~\m6_data_i[5] ) & (~\new_[31989]_  | ~\m7_data_i[5] );
  assign \new_[8598]_  = ~\new_[10268]_  & ~\new_[10035]_ ;
  assign \new_[8599]_  = (~\new_[13530]_  | ~\m2_data_i[5] ) & (~\new_[11611]_  | ~\m3_data_i[5] );
  assign \new_[8600]_  = (~\new_[13530]_  | ~\m2_data_i[4] ) & (~\new_[11611]_  | ~\m3_data_i[4] );
  assign \new_[8601]_  = (~\new_[11773]_  | ~\m6_data_i[4] ) & (~\new_[31989]_  | ~\m7_data_i[4] );
  assign \new_[8602]_  = (~\new_[13530]_  | ~\m2_data_i[3] ) & (~\new_[11611]_  | ~\m3_data_i[3] );
  assign \new_[8603]_  = (~\new_[11773]_  | ~\m6_data_i[3] ) & (~\new_[11539]_  | ~\m7_data_i[3] );
  assign \new_[8604]_  = (~\new_[13530]_  | ~\m2_data_i[2] ) & (~\new_[11611]_  | ~\m3_data_i[2] );
  assign \new_[8605]_  = (~\new_[11773]_  | ~\m6_data_i[2] ) & (~\new_[31989]_  | ~\m7_data_i[2] );
  assign \new_[8606]_  = (~\new_[13530]_  | ~\m2_data_i[1] ) & (~\new_[11613]_  | ~\m3_data_i[1] );
  assign \new_[8607]_  = ~\new_[9818]_  & ~\new_[9766]_ ;
  assign \new_[8608]_  = (~\new_[11773]_  | ~\m6_data_i[1] ) & (~\new_[11539]_  | ~\m7_data_i[1] );
  assign \new_[8609]_  = (~\new_[13530]_  | ~\m2_data_i[0] ) & (~\new_[11613]_  | ~\m3_data_i[0] );
  assign \new_[8610]_  = (~\new_[11773]_  | ~\m6_data_i[0] ) & (~\new_[31989]_  | ~\m7_data_i[0] );
  assign \new_[8611]_  = ~\new_[9768]_  & ~\new_[9825]_ ;
  assign \new_[8612]_  = ~\new_[10361]_  & ~\new_[10067]_ ;
  assign \new_[8613]_  = ~\new_[19380]_  | ~\new_[13554]_  | ~\new_[21262]_  | ~\new_[15567]_ ;
  assign \new_[8614]_  = ~\new_[20366]_  | ~\new_[13555]_  | ~\new_[19605]_  | ~\new_[15571]_ ;
  assign \new_[8615]_  = ~\new_[21268]_  | ~\new_[13556]_  | ~\new_[18405]_  | ~\new_[16513]_ ;
  assign \new_[8616]_  = ~\new_[9962]_  | ~\new_[11759]_ ;
  assign \new_[8617]_  = ~\new_[9966]_  | ~\new_[10022]_ ;
  assign \new_[8618]_  = ~\new_[21277]_  | ~\new_[13557]_  | ~\new_[20368]_  | ~\new_[12789]_ ;
  assign \new_[8619]_  = ~\new_[9972]_  | ~\new_[10030]_ ;
  assign \new_[8620]_  = ~\new_[11694]_  | ~\new_[10032]_ ;
  assign \new_[8621]_  = ~\new_[21283]_  | ~\new_[13559]_  | ~\new_[21312]_  | ~\new_[14271]_ ;
  assign \new_[8622]_  = ~\new_[9978]_  | ~\new_[10033]_ ;
  assign \new_[8623]_  = ~\new_[9980]_  | ~\new_[10038]_ ;
  assign \new_[8624]_  = ~\new_[19383]_  | ~\new_[14908]_  | ~\new_[21289]_  | ~\new_[12811]_ ;
  assign \new_[8625]_  = ~\new_[11699]_  | ~\new_[10040]_ ;
  assign \new_[8626]_  = ~\new_[9983]_  | ~\new_[10043]_ ;
  assign \new_[8627]_  = ~\new_[9987]_  | ~\new_[10045]_ ;
  assign \new_[8628]_  = ~\new_[19390]_  | ~\new_[13560]_  | ~\new_[21279]_  | ~\new_[15618]_ ;
  assign \new_[8629]_  = ~\new_[9990]_  | ~\new_[11791]_ ;
  assign \new_[8630]_  = ~\new_[18406]_  | ~\new_[13561]_  | ~\new_[21272]_  | ~\new_[15624]_ ;
  assign \new_[8631]_  = ~\new_[9998]_  | ~\new_[10050]_ ;
  assign \new_[8632]_  = ~\new_[21280]_  | ~\new_[13562]_  | ~\new_[18415]_  | ~\new_[12832]_ ;
  assign \new_[8633]_  = ~\new_[11728]_  | ~\new_[10057]_ ;
  assign \new_[8634]_  = ~\new_[21313]_  | ~\new_[13563]_  | ~\new_[21304]_  | ~\new_[15644]_ ;
  assign \new_[8635]_  = ~\new_[19398]_  | ~\new_[13564]_  | ~\new_[21327]_  | ~\new_[15650]_ ;
  assign \new_[8636]_  = ~\new_[19354]_  | ~\new_[13583]_  | ~\new_[20390]_  | ~\new_[15597]_ ;
  assign \new_[8637]_  = ~\new_[28647]_  & (~\new_[12018]_  | ~\new_[28420]_ );
  assign \new_[8638]_  = ~\new_[29942]_  & (~\new_[12023]_  | ~\new_[28574]_ );
  assign \new_[8639]_  = ~\new_[28673]_  & (~\new_[12038]_  | ~\new_[27130]_ );
  assign \new_[8640]_  = ~\new_[28738]_  & (~\new_[12048]_  | ~\new_[28606]_ );
  assign \new_[8641]_  = (~\new_[13530]_  | ~m2_we_i) & (~\new_[11613]_  | ~m3_we_i);
  assign \new_[8642]_  = (~\new_[11773]_  | ~m6_we_i) & (~\new_[31989]_  | ~m7_we_i);
  assign \new_[8643]_  = ~\new_[29076]_  & (~\new_[12051]_  | ~\new_[28346]_ );
  assign \new_[8644]_  = ~\new_[29555]_  & (~\new_[12056]_  | ~\new_[28193]_ );
  assign \new_[8645]_  = ~\new_[19341]_  | (~\new_[12137]_  & ~\new_[28300]_ );
  assign \new_[8646]_  = ~\new_[21122]_  | (~\new_[12138]_  & ~\new_[27878]_ );
  assign \new_[8647]_  = ~\new_[19345]_  | (~\new_[12141]_  & ~\new_[28252]_ );
  assign \new_[8648]_  = ~\new_[21134]_  | (~\new_[12145]_  & ~\new_[27842]_ );
  assign \new_[8649]_  = ~\new_[19347]_  | (~\new_[12148]_  & ~\new_[26801]_ );
  assign \new_[8650]_  = ~\new_[20298]_  | (~\new_[12149]_  & ~\new_[28552]_ );
  assign \new_[8651]_  = ~\new_[20310]_  | (~\new_[12153]_  & ~\new_[27900]_ );
  assign \new_[8652]_  = ~\new_[20312]_  | (~\new_[12156]_  & ~\new_[26508]_ );
  assign \new_[8653]_  = ~\new_[20327]_  | (~\new_[13753]_  & ~\new_[28706]_ );
  assign \new_[8654]_  = ~\new_[20346]_  | (~\new_[13755]_  & ~\new_[29673]_ );
  assign \new_[8655]_  = ~\new_[20332]_  | (~\new_[13757]_  & ~\new_[28195]_ );
  assign \new_[8656]_  = ~\new_[20362]_  | (~\new_[13761]_  & ~\new_[29152]_ );
  assign \new_[8657]_  = ~\new_[19376]_  | (~\new_[13765]_  & ~\new_[29643]_ );
  assign \new_[8658]_  = (~\m5_data_i[12]  | ~\new_[18004]_ ) & (~\m6_data_i[12]  | ~\new_[17241]_ );
  assign \new_[8659]_  = (~\m1_addr_i[5]  | ~\new_[17277]_ ) & (~\m0_addr_i[5]  | ~\new_[16280]_ );
  assign \new_[8660]_  = \new_[12076]_  & \new_[14958]_ ;
  assign \new_[8661]_  = ~\new_[12002]_  & (~\new_[14195]_  | ~\new_[28626]_ );
  assign \new_[8662]_  = ~\new_[15565]_  & ~\new_[11907]_ ;
  assign \new_[8663]_  = ~\new_[12554]_  & ~\new_[11993]_ ;
  assign \new_[8664]_  = ~\new_[12058]_  & ~\new_[12448]_ ;
  assign n7609 = (~\new_[13795]_  & ~rst_i) | (~\new_[31130]_  & ~\new_[31853]_ );
  assign \new_[8666]_  = ~\new_[12004]_  | ~\new_[26839]_ ;
  assign n7659 = ~\new_[12089]_  & ~\new_[12091]_ ;
  assign \new_[8668]_  = ~\new_[12065]_  & ~\new_[12470]_ ;
  assign \new_[8669]_  = ~\new_[12010]_  | ~\new_[27602]_ ;
  assign \new_[8670]_  = ~\new_[14079]_  & ~\new_[11999]_ ;
  assign \new_[8671]_  = ~\new_[12068]_  & ~\new_[12482]_ ;
  assign \new_[8672]_  = ~\new_[15292]_  & ~\new_[11928]_ ;
  assign \new_[8673]_  = ~\new_[11972]_  & (~\new_[14210]_  | ~\new_[26570]_ );
  assign \new_[8674]_  = ~\new_[12555]_  & ~\new_[11995]_ ;
  assign \new_[8675]_  = ~\new_[12073]_  & ~\new_[14004]_ ;
  assign \new_[8676]_  = ~\new_[12556]_  & ~\new_[11996]_ ;
  assign \new_[8677]_  = ~\new_[14010]_  & ~\new_[11935]_ ;
  assign \new_[8678]_  = (~\m1_addr_i[15]  | ~\new_[17277]_ ) & (~\m0_addr_i[15]  | ~\new_[16280]_ );
  assign \new_[8679]_  = ~\new_[12025]_  & (~\new_[14216]_  | ~\new_[27943]_ );
  assign \new_[8680]_  = ~\new_[14015]_  & ~\new_[12166]_ ;
  assign \new_[8681]_  = ~\new_[12079]_  & ~\new_[12508]_ ;
  assign \new_[8682]_  = ~\new_[11942]_  & ~\new_[12177]_ ;
  assign \new_[8683]_  = ~\new_[12032]_  | ~\new_[28384]_ ;
  assign \new_[8684]_  = ~\new_[12040]_  & (~\new_[14228]_  | ~\new_[26688]_ );
  assign \new_[8685]_  = ~\new_[13702]_  & ~\new_[12539]_ ;
  assign \new_[8686]_  = ~\new_[12043]_  | ~\new_[28294]_ ;
  assign \s10_data_o[18]  = ~\new_[14990]_  | ~\new_[14991]_  | ~\new_[13719]_  | ~\new_[13720]_ ;
  assign \s10_data_o[9]  = ~\new_[15004]_  | ~\new_[15005]_  | ~\new_[12147]_  | ~\new_[13737]_ ;
  assign \s10_data_o[7]  = ~\new_[15008]_  | ~\new_[15009]_  | ~\new_[12154]_  | ~\new_[13849]_ ;
  assign \s10_data_o[4]  = ~\new_[16359]_  | ~\new_[15013]_  | ~\new_[12162]_  | ~\new_[13751]_ ;
  assign \s10_data_o[3]  = ~\new_[15014]_  | ~\new_[16361]_  | ~\new_[12165]_  | ~\new_[13752]_ ;
  assign \new_[8692]_  = ~\new_[14051]_  & ~\new_[12200]_ ;
  assign \s10_addr_o[8]  = ~\new_[15067]_  | ~\new_[15069]_  | ~\new_[12256]_  | ~\new_[15066]_ ;
  assign \s10_addr_o[7]  = ~\new_[15070]_  | ~\new_[15071]_  | ~\new_[12258]_  | ~\new_[13803]_ ;
  assign \s10_addr_o[2]  = ~\new_[15089]_  | ~\new_[15091]_  | ~\new_[11806]_  | ~\new_[15086]_ ;
  assign \s10_addr_o[1]  = ~\new_[15093]_  | ~\new_[15095]_  | ~\new_[12276]_  | ~\new_[16381]_ ;
  assign \s10_sel_o[3]  = ~\new_[16384]_  | ~\new_[15101]_  | ~\new_[14116]_  | ~\new_[13826]_ ;
  assign \new_[8698]_  = ~\new_[12049]_  & (~\new_[14234]_  | ~\new_[27796]_ );
  assign \new_[8699]_  = ~\new_[12558]_  & ~\new_[12000]_ ;
  assign \new_[8700]_  = ~\new_[12103]_  & ~\new_[12547]_ ;
  assign \new_[8701]_  = ~\new_[12052]_  & (~\new_[14235]_  | ~\new_[28375]_ );
  assign \new_[8702]_  = (~\m5_data_i[18]  | ~\new_[18004]_ ) & (~\m6_data_i[18]  | ~\new_[17241]_ );
  assign \new_[8703]_  = ~\new_[12094]_  & ~\new_[11954]_ ;
  assign \new_[8704]_  = ~\new_[13730]_  & ~\new_[11969]_ ;
  assign \new_[8705]_  = ~\new_[30134]_  & (~\new_[14124]_  | ~\new_[28298]_ );
  assign \new_[8706]_  = ~\new_[14961]_  & ~\new_[11908]_ ;
  assign \new_[8707]_  = ~\new_[28338]_  & (~\new_[13855]_  | ~\new_[22835]_ );
  assign \new_[8708]_  = ~\new_[29424]_  & (~\new_[14126]_  | ~\new_[26299]_ );
  assign \new_[8709]_  = ~\new_[27799]_  & (~\new_[13863]_  | ~\new_[22777]_ );
  assign \new_[8710]_  = ~\new_[28831]_  & (~\new_[14128]_  | ~\new_[23093]_ );
  assign \new_[8711]_  = ~\new_[24623]_  & (~\new_[14161]_  | ~\new_[28525]_ );
  assign \new_[8712]_  = ~\new_[13684]_  & ~\new_[11917]_ ;
  assign \new_[8713]_  = ~\new_[12009]_  & (~\new_[14546]_  | ~\new_[27806]_ );
  assign \new_[8714]_  = ~\new_[29232]_  & (~\new_[13775]_  | ~\new_[24210]_ );
  assign \new_[8715]_  = ~\new_[29543]_  & (~\new_[13871]_  | ~\new_[21354]_ );
  assign \new_[8716]_  = ~\new_[26858]_  & (~\new_[14164]_  | ~\new_[28551]_ );
  assign \new_[8717]_  = ~\new_[28028]_  & (~\new_[13776]_  | ~\new_[22736]_ );
  assign \new_[8718]_  = ~\new_[28812]_  & (~\new_[13879]_  | ~\new_[22682]_ );
  assign \new_[8719]_  = ~\new_[29363]_  & (~\new_[13886]_  | ~\new_[18424]_ );
  assign \new_[8720]_  = ~\new_[28342]_  & (~\new_[13891]_  | ~\new_[20419]_ );
  assign \new_[8721]_  = ~\new_[12017]_  & (~\new_[15938]_  | ~\new_[29532]_ );
  assign \new_[8722]_  = ~\new_[23109]_  & (~\new_[14133]_  | ~\new_[28570]_ );
  assign \new_[8723]_  = ~\new_[23103]_  & (~\new_[14167]_  | ~\new_[28522]_ );
  assign \new_[8724]_  = ~\new_[27372]_  & (~\new_[14166]_  | ~\new_[26806]_ );
  assign \new_[8725]_  = ~\new_[11974]_  & (~\new_[15932]_  | ~\new_[26451]_ );
  assign \new_[8726]_  = ~\new_[27935]_  & (~\new_[13896]_  | ~\new_[19421]_ );
  assign \new_[8727]_  = ~\new_[11975]_  & (~\new_[14516]_  | ~\new_[27989]_ );
  assign \new_[8728]_  = ~\new_[28777]_  & (~\new_[14170]_  | ~\new_[24751]_ );
  assign \new_[8729]_  = ~\new_[28124]_  & (~\new_[14136]_  | ~\new_[26585]_ );
  assign \new_[8730]_  = ~\new_[28062]_  & (~\new_[13903]_  | ~\new_[21420]_ );
  assign \new_[8731]_  = ~\new_[12022]_  & (~\new_[16475]_  | ~\new_[29131]_ );
  assign \new_[8732]_  = ~\new_[30306]_  & (~\new_[14174]_  | ~\new_[26248]_ );
  assign \new_[8733]_  = ~\new_[14968]_  & ~\new_[11937]_ ;
  assign \new_[8734]_  = ~\new_[30171]_  & (~\new_[13781]_  | ~\new_[21371]_ );
  assign \new_[8735]_  = ~\new_[28605]_  & (~\new_[13916]_  | ~\new_[21425]_ );
  assign \new_[8736]_  = ~\new_[12026]_  & (~\new_[16341]_  | ~\new_[29074]_ );
  assign \new_[8737]_  = ~\new_[28037]_  & (~\new_[14140]_  | ~\new_[23547]_ );
  assign \new_[8738]_  = ~\new_[24479]_  & (~\new_[14178]_  | ~\new_[28743]_ );
  assign \new_[8739]_  = ~\new_[28063]_  & (~\new_[13924]_  | ~\new_[21402]_ );
  assign \new_[8740]_  = ~\new_[30143]_  & (~\new_[14144]_  | ~\new_[26837]_ );
  assign \new_[8741]_  = ~\new_[29843]_  & (~\new_[13784]_  | ~\new_[22727]_ );
  assign \new_[8742]_  = ~\new_[28616]_  & (~\new_[13931]_  | ~\new_[21488]_ );
  assign \new_[8743]_  = ~\new_[28155]_  & (~\new_[14180]_  | ~\new_[24461]_ );
  assign \new_[8744]_  = ~\new_[12034]_  & (~\new_[14876]_  | ~\new_[28615]_ );
  assign \new_[8745]_  = ~\new_[28165]_  & (~\new_[13937]_  | ~\new_[22764]_ );
  assign \new_[8746]_  = ~\new_[12035]_  & (~\new_[14860]_  | ~\new_[29378]_ );
  assign \new_[8747]_  = ~\new_[15393]_  & ~\new_[12211]_ ;
  assign \new_[8748]_  = ~\new_[30358]_  & (~\new_[14147]_  | ~\new_[24621]_ );
  assign \new_[8749]_  = ~\new_[13699]_  & ~\new_[11951]_ ;
  assign \new_[8750]_  = ~\new_[28212]_  & (~\new_[13948]_  | ~\new_[20442]_ );
  assign \new_[8751]_  = ~\new_[25189]_  | ~\new_[11890]_ ;
  assign \new_[8752]_  = ~\new_[28321]_  & (~\new_[14183]_  | ~\new_[24544]_ );
  assign \new_[8753]_  = ~\new_[29236]_  & (~\new_[14151]_  | ~\new_[26712]_ );
  assign \new_[8754]_  = (~\m4_data_i[31]  | ~\new_[16307]_ ) & (~\m3_data_i[31]  | ~\new_[17249]_ );
  assign \new_[8755]_  = ~\new_[14972]_  & ~\new_[11956]_ ;
  assign \new_[8756]_  = ~\new_[28581]_  & (~\new_[13787]_  | ~\new_[22832]_ );
  assign \new_[8757]_  = ~\new_[28720]_  & (~\new_[14152]_  | ~\new_[24633]_ );
  assign \new_[8758]_  = ~\new_[12046]_  & (~\new_[14999]_  | ~\new_[26536]_ );
  assign \new_[8759]_  = ~\new_[28618]_  & (~\new_[13960]_  | ~\new_[22771]_ );
  assign \new_[8760]_  = ~\new_[12047]_  & (~\new_[13606]_  | ~\new_[29535]_ );
  assign \new_[8761]_  = ~\new_[27929]_  & (~\new_[14188]_  | ~\new_[24541]_ );
  assign \new_[8762]_  = ~\new_[28920]_  & (~\new_[13788]_  | ~\new_[22822]_ );
  assign \new_[8763]_  = ~\new_[29243]_  & (~\new_[13790]_  | ~\new_[23845]_ );
  assign \new_[8764]_  = ~\new_[28624]_  & (~\new_[13969]_  | ~\new_[19407]_ );
  assign \new_[8765]_  = ~\new_[28983]_  & (~\new_[14189]_  | ~\new_[26428]_ );
  assign \new_[8766]_  = ~\new_[14997]_  & ~\new_[11967]_ ;
  assign \new_[8767]_  = ~\new_[28600]_  & (~\new_[13976]_  | ~\new_[20444]_ );
  assign \new_[8768]_  = ~\new_[27041]_  | ~\new_[11904]_ ;
  assign \new_[8769]_  = (~\m5_data_i[4]  | ~\new_[18004]_ ) & (~\m6_data_i[4]  | ~\new_[17241]_ );
  assign \new_[8770]_  = ~\new_[26454]_  & (~\new_[13856]_  | ~\new_[20476]_ );
  assign \new_[8771]_  = ~\new_[28831]_  & (~\new_[13864]_  | ~\new_[21939]_ );
  assign \new_[8772]_  = ~\new_[24623]_  & (~\new_[13865]_  | ~\new_[20005]_ );
  assign \new_[8773]_  = ~\new_[26858]_  & (~\new_[13874]_  | ~\new_[23019]_ );
  assign \new_[8774]_  = ~\new_[28735]_  & (~\new_[13881]_  | ~\new_[22976]_ );
  assign \new_[8775]_  = ~\new_[28613]_  & (~\new_[13898]_  | ~\new_[20462]_ );
  assign \new_[8776]_  = ~\new_[28124]_  & (~\new_[13900]_  | ~\new_[24296]_ );
  assign \new_[8777]_  = ~\new_[28607]_  & (~\new_[13909]_  | ~\new_[20483]_ );
  assign \new_[8778]_  = ~\new_[28037]_  & (~\new_[13917]_  | ~\new_[23714]_ );
  assign \new_[8779]_  = ~\new_[24479]_  & (~\new_[13918]_  | ~\new_[20509]_ );
  assign \new_[8780]_  = ~\new_[30143]_  & (~\new_[13926]_  | ~\new_[22156]_ );
  assign \new_[8781]_  = ~\new_[28155]_  & (~\new_[13932]_  | ~\new_[21498]_ );
  assign \new_[8782]_  = ~\new_[30358]_  & (~\new_[13940]_  | ~\new_[20480]_ );
  assign \new_[8783]_  = ~\new_[27788]_  & (~\new_[13941]_  | ~\new_[20491]_ );
  assign \new_[8784]_  = ~\new_[28087]_  & (~\new_[13950]_  | ~\new_[21524]_ );
  assign \new_[8785]_  = ~\new_[26462]_  & (~\new_[13957]_  | ~\new_[19786]_ );
  assign \new_[8786]_  = ~\new_[28599]_  & (~\new_[13964]_  | ~\new_[20486]_ );
  assign \new_[8787]_  = ~\new_[30165]_  & (~\new_[13970]_  | ~\new_[20475]_ );
  assign \new_[8788]_  = ~\new_[28044]_  & (~\new_[13971]_  | ~\new_[21602]_ );
  assign \new_[8789]_  = ~\new_[29533]_  & (~\new_[13852]_  | ~\new_[21481]_ );
  assign \new_[8790]_  = ~\new_[26630]_  & (~\new_[13893]_  | ~\new_[21401]_ );
  assign \new_[8791]_  = ~\new_[27363]_  & (~\new_[14350]_  | ~\new_[26362]_ );
  assign \new_[8792]_  = ~\new_[27823]_  & (~\new_[13797]_  | ~\new_[21567]_ );
  assign \new_[8793]_  = ~\new_[27890]_  & (~\new_[13801]_  | ~\new_[24393]_ );
  assign \new_[8794]_  = ~\new_[27906]_  & (~\new_[13802]_  | ~\new_[23026]_ );
  assign \new_[8795]_  = ~\new_[29599]_  & (~\new_[13806]_  | ~\new_[21543]_ );
  assign \new_[8796]_  = \new_[20369]_  & \new_[11971]_ ;
  assign \new_[8797]_  = ~\new_[27949]_  & (~\new_[13814]_  | ~\new_[22933]_ );
  assign \new_[8798]_  = ~\new_[29147]_  & (~\new_[13818]_  | ~\new_[22993]_ );
  assign \new_[8799]_  = ~\new_[26964]_  & (~\new_[13822]_  | ~\new_[21485]_ );
  assign \new_[8800]_  = ~\new_[27839]_  & (~\new_[13827]_  | ~\new_[21522]_ );
  assign \new_[8801]_  = ~\new_[27829]_  & (~\new_[13830]_  | ~\new_[22898]_ );
  assign \new_[8802]_  = ~\new_[27502]_  & (~\new_[13834]_  | ~\new_[21600]_ );
  assign \new_[8803]_  = ~\new_[27916]_  & (~\new_[13837]_  | ~\new_[23052]_ );
  assign \new_[8804]_  = ~\new_[27931]_  & (~\new_[13841]_  | ~\new_[20512]_ );
  assign \new_[8805]_  = ~\new_[28226]_  & (~\new_[13847]_  | ~\new_[22864]_ );
  assign \new_[8806]_  = ~\new_[29585]_  & (~\new_[13850]_  | ~\new_[22997]_ );
  assign \new_[8807]_  = ~\new_[29126]_  & (~\new_[13977]_  | ~\new_[29318]_ );
  assign \new_[8808]_  = ~\new_[27876]_  | (~\new_[14241]_  & ~\new_[26250]_ );
  assign \new_[8809]_  = ~\new_[27933]_  | (~\new_[14248]_  & ~\new_[25351]_ );
  assign \new_[8810]_  = ~\new_[26748]_  | (~\new_[14253]_  & ~\new_[26206]_ );
  assign \new_[8811]_  = ~\new_[28172]_  & (~\new_[13989]_  | ~\new_[21618]_ );
  assign \new_[8812]_  = ~\new_[26508]_  & (~\new_[13993]_  | ~\new_[22991]_ );
  assign \new_[8813]_  = ~\new_[24492]_  & (~\new_[13994]_  | ~\new_[24730]_ );
  assign \new_[8814]_  = ~\new_[28022]_  & (~\new_[13778]_  | ~\new_[24336]_ );
  assign \new_[8815]_  = ~\new_[26819]_  & (~\new_[14212]_  | ~\new_[20416]_ );
  assign \new_[8816]_  = ~\new_[27949]_  & (~\new_[14006]_  | ~\new_[21574]_ );
  assign \new_[8817]_  = ~\new_[26332]_  & (~\new_[14008]_  | ~\new_[22943]_ );
  assign \new_[8818]_  = ~\new_[29147]_  & (~\new_[14012]_  | ~\new_[23049]_ );
  assign \new_[8819]_  = ~\new_[28173]_  & (~\new_[14014]_  | ~\new_[28956]_ );
  assign \new_[8820]_  = ~\new_[26877]_  & (~\new_[14019]_  | ~\new_[21572]_ );
  assign \new_[8821]_  = ~\new_[26589]_  | (~\new_[14286]_  & ~\new_[26200]_ );
  assign \new_[8822]_  = ~\new_[30007]_  & (~\new_[14026]_  | ~\new_[21604]_ );
  assign \new_[8823]_  = ~\new_[26823]_  | (~\new_[14293]_  & ~\new_[24768]_ );
  assign \new_[8824]_  = ~\new_[27767]_  | (~\new_[14300]_  & ~\new_[26233]_ );
  assign \new_[8825]_  = ~\new_[28973]_  & (~\new_[14039]_  | ~\new_[22994]_ );
  assign \new_[8826]_  = ~\new_[29200]_  & (~\new_[14313]_  | ~\new_[28573]_ );
  assign \new_[8827]_  = ~\new_[27819]_  | (~\new_[14266]_  & ~\new_[26279]_ );
  assign \new_[8828]_  = (~\m5_addr_i[2]  | ~\new_[18004]_ ) & (~\m6_addr_i[2]  | ~\new_[17241]_ );
  assign \new_[8829]_  = ~\new_[28226]_  & (~\new_[14056]_  | ~\new_[22979]_ );
  assign \new_[8830]_  = ~\new_[29585]_  & (~\new_[14065]_  | ~\new_[22929]_ );
  assign \new_[8831]_  = ~\new_[24742]_  & (~\new_[14066]_  | ~\new_[21609]_ );
  assign \new_[8832]_  = (~\m1_addr_i[22]  | ~\new_[17277]_ ) & (~\m0_addr_i[22]  | ~\new_[16279]_ );
  assign \new_[8833]_  = ~\new_[26474]_  & (~\new_[14067]_  | ~\new_[27922]_ );
  assign \new_[8834]_  = ~\new_[28064]_  | (~\new_[14345]_  & ~\new_[27437]_ );
  assign \new_[8835]_  = ~\new_[30077]_  | (~\new_[14346]_  & ~\new_[27615]_ );
  assign \new_[8836]_  = ~\new_[28629]_  | (~\new_[14347]_  & ~\new_[26862]_ );
  assign \new_[8837]_  = ~\new_[29658]_  | (~\new_[14348]_  & ~\new_[26409]_ );
  assign \new_[8838]_  = ~\new_[28879]_  | (~\new_[14349]_  & ~\new_[24744]_ );
  assign \new_[8839]_  = ~\new_[29678]_  | (~\new_[14351]_  & ~\new_[24511]_ );
  assign \new_[8840]_  = ~\new_[28156]_  | (~\new_[14352]_  & ~\new_[27558]_ );
  assign \new_[8841]_  = ~\new_[29586]_  | (~\new_[14353]_  & ~\new_[26393]_ );
  assign \new_[8842]_  = ~\new_[27999]_  | (~\new_[14356]_  & ~\new_[28376]_ );
  assign \new_[8843]_  = ~\new_[28030]_  | (~\new_[14357]_  & ~\new_[26450]_ );
  assign \new_[8844]_  = ~\new_[29265]_  | (~\new_[14358]_  & ~\new_[26733]_ );
  assign \new_[8845]_  = ~\new_[29144]_  | (~\new_[14359]_  & ~\new_[25065]_ );
  assign \new_[8846]_  = ~\new_[29143]_  | (~\new_[14360]_  & ~\new_[28491]_ );
  assign \new_[8847]_  = ~\new_[29373]_  | (~\new_[14364]_  & ~\new_[27289]_ );
  assign \new_[8848]_  = ~\new_[28822]_  | (~\new_[14363]_  & ~\new_[26416]_ );
  assign \new_[8849]_  = ~\new_[28854]_  | (~\new_[14365]_  & ~\new_[25386]_ );
  assign \new_[8850]_  = ~\new_[28986]_  | (~\new_[14366]_  & ~\new_[26433]_ );
  assign \new_[8851]_  = ~\new_[31995]_ ;
  assign \new_[8852]_  = ~\new_[28179]_  & (~\new_[14199]_  | ~\new_[24205]_ );
  assign \new_[8853]_  = ~\new_[28189]_  & (~\new_[14086]_  | ~\new_[19468]_ );
  assign \new_[8854]_  = ~\new_[24553]_  & (~\new_[14201]_  | ~\new_[21405]_ );
  assign \new_[8855]_  = ~\new_[27977]_  & (~\new_[14089]_  | ~\new_[29459]_ );
  assign \new_[8856]_  = ~\new_[28648]_  & (~\new_[14202]_  | ~\new_[20427]_ );
  assign \new_[8857]_  = ~\new_[28922]_  & (~\new_[14090]_  | ~\new_[29044]_ );
  assign \new_[8858]_  = ~\new_[29689]_  & (~\new_[14091]_  | ~\new_[17409]_ );
  assign \new_[8859]_  = ~\new_[28255]_  & (~\new_[14209]_  | ~\new_[22814]_ );
  assign \new_[8860]_  = ~\new_[27949]_  & (~\new_[14094]_  | ~\new_[23036]_ );
  assign \new_[8861]_  = ~\new_[28159]_  & (~\new_[14215]_  | ~\new_[21418]_ );
  assign \new_[8862]_  = ~\new_[29147]_  & (~\new_[14096]_  | ~\new_[23047]_ );
  assign \new_[8863]_  = ~\new_[11613]_ ;
  assign \new_[8864]_  = ~\new_[28267]_  & (~\new_[14217]_  | ~\new_[22724]_ );
  assign \new_[8865]_  = ~\new_[29060]_  & (~\new_[14098]_  | ~\new_[17353]_ );
  assign \new_[8866]_  = ~\new_[24647]_  & (~\new_[14099]_  | ~\new_[29757]_ );
  assign \new_[8867]_  = (~\m5_addr_i[7]  | ~\new_[18004]_ ) & (~\m6_addr_i[7]  | ~\new_[17241]_ );
  assign \new_[8868]_  = ~\new_[27998]_  & (~\new_[14219]_  | ~\new_[21393]_ );
  assign \new_[8869]_  = ~\new_[26582]_  & (~\new_[14100]_  | ~\new_[17406]_ );
  assign \new_[8870]_  = ~\new_[28493]_  & (~\new_[14221]_  | ~\new_[22792]_ );
  assign \new_[8871]_  = ~\new_[29247]_  & (~\new_[14222]_  | ~\new_[20431]_ );
  assign \new_[8872]_  = ~\new_[28312]_  & (~\new_[14223]_  | ~\new_[24111]_ );
  assign \new_[8873]_  = ~\new_[29675]_  & (~\new_[14101]_  | ~\new_[28825]_ );
  assign \new_[8874]_  = ~\new_[27870]_  & (~\new_[14224]_  | ~\new_[21419]_ );
  assign \new_[8875]_  = ~\new_[27701]_  & (~\new_[14103]_  | ~\new_[17414]_ );
  assign \new_[8876]_  = ~\new_[29054]_  & (~\new_[14226]_  | ~\new_[19420]_ );
  assign n7604 = ~\new_[30184]_  | (~\new_[14114]_  & ~rst_i);
  assign \new_[8878]_  = ~\new_[25457]_  & (~\new_[14229]_  | ~\new_[21411]_ );
  assign \new_[8879]_  = ~\new_[26714]_  & (~\new_[14231]_  | ~\new_[22827]_ );
  assign \new_[8880]_  = ~\new_[28190]_  & (~\new_[14233]_  | ~\new_[21409]_ );
  assign \new_[8881]_  = ~\new_[28226]_  & (~\new_[14105]_  | ~\new_[23027]_ );
  assign \new_[8882]_  = ~\new_[29585]_  & (~\new_[14107]_  | ~\new_[22895]_ );
  assign \new_[8883]_  = ~\new_[28205]_  & (~\new_[14237]_  | ~\new_[24243]_ );
  assign \new_[8884]_  = ~\new_[28094]_  & (~\new_[14109]_  | ~\new_[21589]_ );
  assign \new_[8885]_  = (~\new_[13978]_  | ~\new_[29179]_ ) & (~\new_[24246]_  | ~\new_[29179]_ );
  assign \new_[8886]_  = ~\new_[27842]_  & (~\new_[13857]_  | ~\new_[21428]_ );
  assign \new_[8887]_  = ~\new_[26485]_  & (~\new_[13858]_  | ~\new_[22799]_ );
  assign \new_[8888]_  = ~\new_[28795]_  & (~\new_[13867]_  | ~\new_[22720]_ );
  assign \new_[8889]_  = ~\new_[28168]_  & (~\new_[13869]_  | ~\new_[22745]_ );
  assign \new_[8890]_  = ~\new_[28948]_  & (~\new_[13870]_  | ~\new_[22743]_ );
  assign \new_[8891]_  = ~\new_[28622]_  & (~\new_[13876]_  | ~\new_[21377]_ );
  assign \new_[8892]_  = ~\new_[28033]_  & (~\new_[13878]_  | ~\new_[21442]_ );
  assign \new_[8893]_  = ~\new_[29005]_  & (~\new_[13889]_  | ~\new_[22754]_ );
  assign \new_[8894]_  = ~\new_[28602]_  & (~\new_[13890]_  | ~\new_[21394]_ );
  assign \new_[8895]_  = ~\new_[26719]_  & (~\new_[13901]_  | ~\new_[20410]_ );
  assign \new_[8896]_  = ~\new_[28326]_  & (~\new_[13902]_  | ~\new_[21390]_ );
  assign \new_[8897]_  = ~\new_[27850]_  & (~\new_[13906]_  | ~\new_[22581]_ );
  assign \new_[8898]_  = ~\new_[28309]_  & (~\new_[13907]_  | ~\new_[22789]_ );
  assign \new_[8899]_  = ~\new_[28347]_  & (~\new_[13912]_  | ~\new_[21372]_ );
  assign \new_[8900]_  = ~\new_[29673]_  & (~\new_[13914]_  | ~\new_[20418]_ );
  assign \new_[8901]_  = ~\new_[28333]_  & (~\new_[13915]_  | ~\new_[21397]_ );
  assign \new_[8902]_  = ~\new_[28782]_  & (~\new_[13920]_  | ~\new_[22586]_ );
  assign \new_[8903]_  = ~\new_[28997]_  & (~\new_[13928]_  | ~\new_[22594]_ );
  assign \new_[8904]_  = ~\new_[27843]_  & (~\new_[13933]_  | ~\new_[19416]_ );
  assign \new_[8905]_  = ~\new_[28627]_  & (~\new_[13934]_  | ~\new_[21374]_ );
  assign \new_[8906]_  = ~\new_[28140]_  & (~\new_[13936]_  | ~\new_[21445]_ );
  assign \new_[8907]_  = ~\new_[28254]_  & (~\new_[13942]_  | ~\new_[20412]_ );
  assign \new_[8908]_  = ~\new_[29088]_  & (~\new_[13943]_  | ~\new_[21415]_ );
  assign \new_[8909]_  = (~\new_[14042]_  | ~\new_[29677]_ ) & (~\new_[26166]_  | ~\new_[29677]_ );
  assign \new_[8910]_  = ~\new_[10002]_ ;
  assign \new_[8911]_  = (~\new_[14046]_  | ~\new_[27103]_ ) & (~\new_[22833]_  | ~\new_[27103]_ );
  assign \new_[8912]_  = ~\new_[26654]_  & (~\new_[13951]_  | ~\new_[20441]_ );
  assign \new_[8913]_  = ~\new_[24572]_  & (~\new_[13952]_  | ~\new_[22572]_ );
  assign \new_[8914]_  = (~\new_[14052]_  | ~\new_[29188]_ ) & (~\new_[22794]_  | ~\new_[29188]_ );
  assign \new_[8915]_  = ~\new_[27869]_  & (~\new_[13958]_  | ~\new_[19413]_ );
  assign \new_[8916]_  = (~\new_[14060]_  | ~\new_[30155]_ ) & (~\new_[23988]_  | ~\new_[30155]_ );
  assign \new_[8917]_  = ~\new_[28711]_  & (~\new_[13965]_  | ~\new_[19419]_ );
  assign \new_[8918]_  = ~\new_[29556]_  & (~\new_[13966]_  | ~\new_[21365]_ );
  assign \new_[8919]_  = ~\new_[28752]_  & (~\new_[13968]_  | ~\new_[22751]_ );
  assign \new_[8920]_  = ~\new_[27972]_  & (~\new_[13972]_  | ~\new_[20437]_ );
  assign \new_[8921]_  = ~\new_[10014]_ ;
  assign \new_[8922]_  = ~\new_[24694]_  & (~\new_[13973]_  | ~\new_[22732]_ );
  assign \new_[8923]_  = (~\new_[14073]_  | ~\new_[29204]_ ) & (~\new_[26179]_  | ~\new_[29204]_ );
  assign \new_[8924]_  = ~\new_[28300]_  & (~\new_[14238]_  | ~\new_[24304]_ );
  assign \new_[8925]_  = ~\new_[29659]_  & (~\new_[14239]_  | ~\new_[23008]_ );
  assign \new_[8926]_  = ~\new_[26482]_  & (~\new_[14240]_  | ~\new_[22901]_ );
  assign \new_[8927]_  = ~\new_[28252]_  & (~\new_[14242]_  | ~\new_[23013]_ );
  assign \new_[8928]_  = ~\new_[28263]_  & (~\new_[14243]_  | ~\new_[19434]_ );
  assign \new_[8929]_  = ~\new_[26460]_  & (~\new_[14246]_  | ~\new_[22885]_ );
  assign \new_[8930]_  = ~\new_[28356]_  & (~\new_[14250]_  | ~\new_[20521]_ );
  assign \new_[8931]_  = ~\new_[26801]_  & (~\new_[14249]_  | ~\new_[24288]_ );
  assign \new_[8932]_  = ~\new_[26452]_  & (~\new_[14252]_  | ~\new_[22890]_ );
  assign \new_[8933]_  = (~\m5_data_i[6]  | ~\new_[18004]_ ) & (~\m6_data_i[6]  | ~\new_[17241]_ );
  assign \new_[8934]_  = ~\new_[28810]_  & (~\new_[14258]_  | ~\new_[22908]_ );
  assign \new_[8935]_  = ~\new_[11773]_ ;
  assign \new_[8936]_  = ~\new_[28175]_  & (~\new_[14265]_  | ~\new_[23119]_ );
  assign \new_[8937]_  = ~\new_[26332]_  & (~\new_[14267]_  | ~\new_[22859]_ );
  assign \new_[8938]_  = ~\new_[26645]_  & (~\new_[14268]_  | ~\new_[20448]_ );
  assign \new_[8939]_  = ~\new_[28779]_  & (~\new_[14272]_  | ~\new_[24439]_ );
  assign \new_[8940]_  = ~\new_[28374]_  & (~\new_[14276]_  | ~\new_[21835]_ );
  assign \new_[8941]_  = ~\new_[26877]_  & (~\new_[14279]_  | ~\new_[23043]_ );
  assign \new_[8942]_  = ~\new_[26634]_  & (~\new_[14281]_  | ~\new_[20493]_ );
  assign \new_[8943]_  = ~\new_[26457]_  & (~\new_[14284]_  | ~\new_[22907]_ );
  assign \new_[8944]_  = ~\new_[30007]_  & (~\new_[14287]_  | ~\new_[22965]_ );
  assign \new_[8945]_  = ~\new_[28936]_  & (~\new_[14288]_  | ~\new_[21526]_ );
  assign \new_[8946]_  = ~\new_[24598]_  & (~\new_[14292]_  | ~\new_[22871]_ );
  assign \new_[8947]_  = ~\new_[28290]_  & (~\new_[14294]_  | ~\new_[21607]_ );
  assign \new_[8948]_  = ~\new_[26510]_  & (~\new_[14299]_  | ~\new_[22903]_ );
  assign \new_[8949]_  = ~\new_[28973]_  & (~\new_[14301]_  | ~\new_[22881]_ );
  assign \new_[8950]_  = ~\new_[29313]_  & (~\new_[14302]_  | ~\new_[20494]_ );
  assign n7654 = ~\new_[12110]_  & ~\new_[12111]_ ;
  assign \new_[8952]_  = (~\new_[13835]_  | ~\new_[29310]_ ) & (~\new_[22741]_  | ~\new_[29310]_ );
  assign \new_[8953]_  = ~\new_[28085]_  & (~\new_[14307]_  | ~\new_[23306]_ );
  assign \new_[8954]_  = ~\new_[28032]_  & (~\new_[14308]_  | ~\new_[22494]_ );
  assign \new_[8955]_  = ~\new_[28257]_  & (~\new_[14309]_  | ~\new_[22989]_ );
  assign \new_[8956]_  = (~\m7_data_i[31]  | ~\new_[16295]_ ) & (~\m0_data_i[31]  | ~\new_[18203]_ );
  assign \new_[8957]_  = ~\new_[24538]_  & (~\new_[14314]_  | ~\new_[22941]_ );
  assign \new_[8958]_  = (~\m2_data_i[31]  | ~\new_[18080]_ ) & (~\m1_data_i[31]  | ~\new_[18167]_ );
  assign \new_[8959]_  = ~\new_[26501]_  & (~\new_[14315]_  | ~\new_[21620]_ );
  assign \new_[8960]_  = ~\new_[26649]_  & (~\new_[14316]_  | ~\new_[19404]_ );
  assign \new_[8961]_  = (~\m5_data_i[30]  | ~\new_[17204]_ ) & (~\m6_data_i[30]  | ~\new_[16287]_ );
  assign \new_[8962]_  = (~\new_[13844]_  | ~\new_[29337]_ ) & (~\new_[22791]_  | ~\new_[29337]_ );
  assign \new_[8963]_  = (~\m7_data_i[30]  | ~\new_[16295]_ ) & (~\m0_data_i[30]  | ~\new_[18204]_ );
  assign \new_[8964]_  = (~\m2_data_i[29]  | ~\new_[16292]_ ) & (~\m1_data_i[29]  | ~\new_[19621]_ );
  assign \new_[8965]_  = ~\new_[28084]_  & (~\new_[14322]_  | ~\new_[23125]_ );
  assign \new_[8966]_  = (~\m2_data_i[28]  | ~\new_[18080]_ ) & (~\m1_data_i[28]  | ~\new_[18167]_ );
  assign \new_[8967]_  = ~\new_[29135]_  & (~\new_[14325]_  | ~\new_[23158]_ );
  assign \new_[8968]_  = (~\m2_data_i[27]  | ~\new_[16292]_ ) & (~\m1_data_i[27]  | ~\new_[18167]_ );
  assign \new_[8969]_  = ~\new_[12082]_  & ~\new_[12171]_ ;
  assign \new_[8970]_  = (~\m2_data_i[26]  | ~\new_[16292]_ ) & (~\m1_data_i[26]  | ~\new_[18167]_ );
  assign \new_[8971]_  = (~\m7_data_i[26]  | ~\new_[16295]_ ) & (~\m0_data_i[26]  | ~\new_[18204]_ );
  assign \new_[8972]_  = ~\new_[28841]_  & (~\new_[14327]_  | ~\new_[24404]_ );
  assign \new_[8973]_  = (~\m7_data_i[25]  | ~\new_[16295]_ ) & (~\m0_data_i[25]  | ~\new_[18203]_ );
  assign \new_[8974]_  = (~\m5_data_i[24]  | ~\new_[17204]_ ) & (~\m6_data_i[24]  | ~\new_[16287]_ );
  assign \new_[8975]_  = (~\m7_data_i[24]  | ~\new_[16295]_ ) & (~\m0_data_i[24]  | ~\new_[18204]_ );
  assign \new_[8976]_  = (~\m2_data_i[24]  | ~\new_[18080]_ ) & (~\m1_data_i[24]  | ~\new_[18167]_ );
  assign \new_[8977]_  = (~\m2_data_i[23]  | ~\new_[16292]_ ) & (~\m1_data_i[23]  | ~\new_[18167]_ );
  assign \new_[8978]_  = (~\m7_data_i[22]  | ~\new_[16295]_ ) & (~\m0_data_i[22]  | ~\new_[18204]_ );
  assign \new_[8979]_  = (~\m2_data_i[22]  | ~\new_[18080]_ ) & (~\m1_data_i[22]  | ~\new_[18167]_ );
  assign \new_[8980]_  = (~\m7_data_i[21]  | ~\new_[16295]_ ) & (~\m0_data_i[21]  | ~\new_[19643]_ );
  assign \new_[8981]_  = (~\m2_data_i[21]  | ~\new_[16292]_ ) & (~\m1_data_i[21]  | ~\new_[18167]_ );
  assign \new_[8982]_  = (~\m2_data_i[20]  | ~\new_[16292]_ ) & (~\m1_data_i[20]  | ~\new_[18167]_ );
  assign \new_[8983]_  = (~\m7_data_i[20]  | ~\new_[16295]_ ) & (~\m0_data_i[20]  | ~\new_[18204]_ );
  assign \new_[8984]_  = (~\m7_data_i[19]  | ~\new_[16295]_ ) & (~\m0_data_i[19]  | ~\new_[19643]_ );
  assign \new_[8985]_  = (~\m2_data_i[19]  | ~\new_[18080]_ ) & (~\m1_data_i[19]  | ~\new_[18167]_ );
  assign \new_[8986]_  = ~\new_[12611]_  | ~\new_[28555]_ ;
  assign \new_[8987]_  = (~\m5_data_i[18]  | ~\new_[17204]_ ) & (~\m6_data_i[18]  | ~\new_[16287]_ );
  assign \new_[8988]_  = (~\m7_data_i[18]  | ~\new_[16295]_ ) & (~\m0_data_i[18]  | ~\new_[19643]_ );
  assign \new_[8989]_  = (~\m2_data_i[18]  | ~\new_[18080]_ ) & (~\m1_data_i[18]  | ~\new_[18167]_ );
  assign \new_[8990]_  = ~\new_[12594]_  | ~\new_[27898]_ ;
  assign \new_[8991]_  = (~\m7_data_i[17]  | ~\new_[16295]_ ) & (~\m0_data_i[17]  | ~\new_[19643]_ );
  assign \new_[8992]_  = \new_[12669]_  | \new_[26250]_ ;
  assign \new_[8993]_  = ~\new_[12613]_  | ~\new_[28532]_ ;
  assign \new_[8994]_  = (~\m2_data_i[16]  | ~\new_[16292]_ ) & (~\m1_data_i[16]  | ~\new_[18167]_ );
  assign \new_[8995]_  = (~\m2_data_i[15]  | ~\new_[16292]_ ) & (~\m1_data_i[15]  | ~\new_[18890]_ );
  assign \new_[8996]_  = ~\new_[12596]_  | ~\new_[27231]_ ;
  assign \new_[8997]_  = \new_[12672]_  | \new_[25351]_ ;
  assign \new_[8998]_  = ~\new_[12617]_  | ~\new_[28722]_ ;
  assign \new_[8999]_  = ~\new_[12673]_  | ~\new_[28492]_ ;
  assign \new_[9000]_  = (~\m2_data_i[14]  | ~\new_[18080]_ ) & (~\m1_data_i[14]  | ~\new_[18167]_ );
  assign \new_[9001]_  = (~\m2_data_i[13]  | ~\new_[16292]_ ) & (~\m1_data_i[13]  | ~\new_[18167]_ );
  assign \new_[9002]_  = ~\new_[12597]_  | ~\new_[26803]_ ;
  assign \new_[9003]_  = \new_[12676]_  | \new_[26206]_ ;
  assign \new_[9004]_  = ~\new_[12677]_  | ~\new_[28481]_ ;
  assign \new_[9005]_  = ~\new_[12598]_  | ~\new_[26192]_ ;
  assign \new_[9006]_  = \new_[12679]_  | \new_[24812]_ ;
  assign \new_[9007]_  = (~\m5_data_i[8]  | ~\new_[17204]_ ) & (~\m6_data_i[8]  | ~\new_[16287]_ );
  assign \new_[9008]_  = (~\m2_data_i[8]  | ~\new_[18080]_ ) & (~\m1_data_i[8]  | ~\new_[18167]_ );
  assign \new_[9009]_  = \new_[12791]_  & \new_[28522]_ ;
  assign \new_[9010]_  = (~\m2_data_i[7]  | ~\new_[16292]_ ) & (~\m1_data_i[7]  | ~\new_[18167]_ );
  assign \new_[9011]_  = ~\new_[12499]_  | ~\new_[28496]_ ;
  assign \new_[9012]_  = (~\m7_data_i[6]  | ~\new_[16295]_ ) & (~\m0_data_i[6]  | ~\new_[18204]_ );
  assign \new_[9013]_  = ~\new_[12625]_  | ~\new_[28420]_ ;
  assign \new_[9014]_  = (~\m2_data_i[5]  | ~\new_[16292]_ ) & (~\m1_data_i[5]  | ~\new_[18167]_ );
  assign \new_[9015]_  = ~\new_[12628]_  | ~\new_[28494]_ ;
  assign \new_[9016]_  = (~\m5_data_i[4]  | ~\new_[17204]_ ) & (~\m6_data_i[4]  | ~\new_[16287]_ );
  assign \new_[9017]_  = (~\m2_data_i[4]  | ~\new_[16292]_ ) & (~\m1_data_i[4]  | ~\new_[19621]_ );
  assign \new_[9018]_  = (~\m7_data_i[4]  | ~\new_[16295]_ ) & (~\m0_data_i[4]  | ~\new_[18204]_ );
  assign \new_[9019]_  = ~\new_[12630]_  | ~\new_[28574]_ ;
  assign \new_[9020]_  = (~\m7_data_i[3]  | ~\new_[16295]_ ) & (~\m0_data_i[3]  | ~\new_[18203]_ );
  assign \new_[9021]_  = (~\m2_data_i[3]  | ~\new_[18080]_ ) & (~\m1_data_i[3]  | ~\new_[18167]_ );
  assign \new_[9022]_  = (~\m2_data_i[2]  | ~\new_[16292]_ ) & (~\m1_data_i[2]  | ~\new_[18890]_ );
  assign \new_[9023]_  = (~\m5_data_i[1]  | ~\new_[17204]_ ) & (~\m6_data_i[1]  | ~\new_[16287]_ );
  assign \new_[9024]_  = (~\m2_data_i[1]  | ~\new_[16292]_ ) & (~\m1_data_i[1]  | ~\new_[18890]_ );
  assign \new_[9025]_  = (~\m7_data_i[1]  | ~\new_[16295]_ ) & (~\m0_data_i[1]  | ~\new_[18204]_ );
  assign \new_[9026]_  = ~\new_[12602]_  | ~\new_[26247]_ ;
  assign \new_[9027]_  = \new_[12687]_  | \new_[26204]_ ;
  assign \new_[9028]_  = (~\m5_data_i[0]  | ~\new_[17204]_ ) & (~\m6_data_i[0]  | ~\new_[16287]_ );
  assign \new_[9029]_  = (~\m7_data_i[0]  | ~\new_[16295]_ ) & (~\m0_data_i[0]  | ~\new_[18204]_ );
  assign \new_[9030]_  = ~\new_[12635]_  | ~\new_[28674]_ ;
  assign \new_[9031]_  = ~\new_[12686]_  | ~\new_[28556]_ ;
  assign \new_[9032]_  = (~\m2_data_i[0]  | ~\new_[18080]_ ) & (~\m1_data_i[0]  | ~\new_[18167]_ );
  assign \new_[9033]_  = (~\new_[16292]_  | ~\m2_addr_i[31] ) & (~\new_[19621]_  | ~\new_[31447]_ );
  assign \new_[9034]_  = (~\new_[16295]_  | ~\m7_addr_i[31] ) & (~\new_[18204]_  | ~\m0_addr_i[31] );
  assign \new_[9035]_  = (~\new_[16287]_  | ~\m6_addr_i[31] ) & (~\new_[18760]_  | ~\new_[31001]_ );
  assign \new_[9036]_  = ~\new_[12603]_  | ~\new_[26437]_ ;
  assign \new_[9037]_  = \new_[12690]_  | \new_[26200]_ ;
  assign \new_[9038]_  = (~\new_[16295]_  | ~\new_[31885]_ ) & (~\new_[18204]_  | ~\new_[31292]_ );
  assign \new_[9039]_  = (~\new_[16287]_  | ~\m6_addr_i[30] ) & (~\new_[18760]_  | ~\new_[31147]_ );
  assign \new_[9040]_  = ~\new_[12640]_  | ~\new_[28097]_ ;
  assign \new_[9041]_  = (~\new_[16287]_  | ~\m6_addr_i[29] ) & (~\new_[17204]_  | ~\new_[31407]_ );
  assign \new_[9042]_  = (~\new_[16292]_  | ~\new_[31000]_ ) & (~\new_[19621]_  | ~\new_[31538]_ );
  assign \new_[9043]_  = (~\new_[16295]_  | ~\new_[30577]_ ) & (~\new_[18204]_  | ~\new_[30957]_ );
  assign \new_[9044]_  = ~\new_[12604]_  | ~\new_[27609]_ ;
  assign \new_[9045]_  = \new_[12692]_  | \new_[24768]_ ;
  assign \new_[9046]_  = (~\new_[16287]_  | ~\m6_addr_i[28] ) & (~\new_[17204]_  | ~\new_[31276]_ );
  assign \new_[9047]_  = ~\new_[12644]_  | ~\new_[28176]_ ;
  assign \new_[9048]_  = ~\new_[12693]_  | ~\new_[28708]_ ;
  assign \new_[9049]_  = ~\new_[12524]_  | ~\new_[28176]_ ;
  assign \new_[9050]_  = (~\new_[16287]_  | ~\m6_addr_i[27] ) & (~\new_[17204]_  | ~\m5_addr_i[27] );
  assign \new_[9051]_  = (~\new_[16287]_  | ~\m6_addr_i[26] ) & (~\new_[18760]_  | ~\m5_addr_i[26] );
  assign \new_[9052]_  = ~\new_[12606]_  | ~\new_[26211]_ ;
  assign \new_[9053]_  = (~\new_[16295]_  | ~\m7_addr_i[26] ) & (~\new_[19643]_  | ~\m0_addr_i[26] );
  assign \new_[9054]_  = \new_[12695]_  | \new_[26233]_ ;
  assign \new_[9055]_  = ~\new_[12648]_  | ~\new_[28564]_ ;
  assign \new_[9056]_  = ~\new_[12697]_  | ~\new_[28573]_ ;
  assign \new_[9057]_  = (~\new_[16287]_  | ~\m6_addr_i[25] ) & (~\new_[18760]_  | ~\m5_addr_i[25] );
  assign \new_[9058]_  = (~\new_[16287]_  | ~\m6_addr_i[24] ) & (~\new_[18760]_  | ~\m5_addr_i[24] );
  assign \new_[9059]_  = (~\new_[16295]_  | ~\m7_addr_i[24] ) & (~\new_[18204]_  | ~\m0_addr_i[24] );
  assign \new_[9060]_  = (~\new_[16292]_  | ~\m2_addr_i[24] ) & (~\new_[19621]_  | ~\m1_addr_i[24] );
  assign \new_[9061]_  = ~\new_[12702]_  | ~\new_[28305]_ ;
  assign \new_[9062]_  = (~\m7_addr_i[23]  | ~\new_[16295]_ ) & (~\m0_addr_i[23]  | ~\new_[18204]_ );
  assign \new_[9063]_  = ~\new_[12652]_  | ~\new_[28477]_ ;
  assign \new_[9064]_  = (~\m2_addr_i[23]  | ~\new_[18080]_ ) & (~\m1_addr_i[23]  | ~\new_[18167]_ );
  assign \new_[9065]_  = (~\m7_addr_i[22]  | ~\new_[16295]_ ) & (~\m0_addr_i[22]  | ~\new_[19643]_ );
  assign \new_[9066]_  = (~\m2_addr_i[22]  | ~\new_[18080]_ ) & (~\m1_addr_i[22]  | ~\new_[18167]_ );
  assign \new_[9067]_  = ~\new_[12608]_  | ~\new_[27703]_ ;
  assign \new_[9068]_  = \new_[12705]_  | \new_[26279]_ ;
  assign \new_[9069]_  = (~\m2_addr_i[21]  | ~\new_[16292]_ ) & (~\m1_addr_i[21]  | ~\new_[18167]_ );
  assign \new_[9070]_  = ~\new_[12654]_  | ~\new_[28643]_ ;
  assign \new_[9071]_  = ~\new_[12545]_  | ~\new_[28643]_ ;
  assign \new_[9072]_  = (~\m7_addr_i[20]  | ~\new_[16295]_ ) & (~\m0_addr_i[20]  | ~\new_[18204]_ );
  assign \new_[9073]_  = (~\m2_addr_i[20]  | ~\new_[16292]_ ) & (~\m1_addr_i[20]  | ~\new_[19621]_ );
  assign \new_[9074]_  = ~\new_[12658]_  | ~\new_[28606]_ ;
  assign \new_[9075]_  = (~\m7_addr_i[19]  | ~\new_[16295]_ ) & (~\m0_addr_i[19]  | ~\new_[19643]_ );
  assign \new_[9076]_  = (~\m2_addr_i[19]  | ~\new_[18080]_ ) & (~\m1_addr_i[19]  | ~\new_[18167]_ );
  assign \new_[9077]_  = (~\m7_addr_i[18]  | ~\new_[16295]_ ) & (~\m0_addr_i[18]  | ~\new_[18204]_ );
  assign \new_[9078]_  = ~\new_[12660]_  | ~\new_[28346]_ ;
  assign \new_[9079]_  = (~\m2_addr_i[17]  | ~\new_[16292]_ ) & (~\m1_addr_i[17]  | ~\new_[18167]_ );
  assign \new_[9080]_  = (~\m7_addr_i[17]  | ~\new_[16295]_ ) & (~\m0_addr_i[17]  | ~\new_[18204]_ );
  assign \new_[9081]_  = (~\m7_addr_i[16]  | ~\new_[16295]_ ) & (~\m0_addr_i[16]  | ~\new_[19643]_ );
  assign \new_[9082]_  = (~\m7_addr_i[15]  | ~\new_[16295]_ ) & (~\m0_addr_i[15]  | ~\new_[19643]_ );
  assign \new_[9083]_  = (~\m2_addr_i[15]  | ~\new_[18080]_ ) & (~\m1_addr_i[15]  | ~\new_[18167]_ );
  assign \new_[9084]_  = (~\m2_addr_i[14]  | ~\new_[16292]_ ) & (~\m1_addr_i[14]  | ~\new_[18167]_ );
  assign \new_[9085]_  = (~\m2_addr_i[13]  | ~\new_[16292]_ ) & (~\m1_addr_i[13]  | ~\new_[18167]_ );
  assign \new_[9086]_  = ~\new_[28310]_  & (~\new_[14371]_  | ~\new_[21483]_ );
  assign \new_[9087]_  = (~\m7_addr_i[12]  | ~\new_[16295]_ ) & (~\m0_addr_i[12]  | ~\new_[18204]_ );
  assign \new_[9088]_  = (~\m2_addr_i[12]  | ~\new_[18080]_ ) & (~\m1_addr_i[12]  | ~\new_[18167]_ );
  assign n7649 = (~\new_[14462]_  & ~rst_i) | (~\new_[31057]_  & ~\new_[31853]_ );
  assign \new_[9090]_  = (~\m2_addr_i[11]  | ~\new_[16292]_ ) & (~\m1_addr_i[11]  | ~\new_[18167]_ );
  assign \new_[9091]_  = ~\new_[18418]_  | ~\new_[12248]_ ;
  assign \new_[9092]_  = ~\new_[29424]_  & (~\new_[14375]_  | ~\new_[22944]_ );
  assign \new_[9093]_  = (~\m7_addr_i[10]  | ~\new_[16295]_ ) & (~\m0_addr_i[10]  | ~\new_[18204]_ );
  assign \new_[9094]_  = (~\m2_addr_i[9]  | ~\new_[16292]_ ) & (~\m1_addr_i[9]  | ~\new_[18167]_ );
  assign \new_[9095]_  = ~\new_[28038]_  & (~\new_[14376]_  | ~\new_[22712]_ );
  assign \new_[9096]_  = ~\new_[28068]_  & (~\new_[14379]_  | ~\new_[24200]_ );
  assign \new_[9097]_  = (~\m7_addr_i[8]  | ~\new_[16295]_ ) & (~\m0_addr_i[8]  | ~\new_[19643]_ );
  assign \new_[9098]_  = (~\m5_data_i[7]  | ~\new_[18004]_ ) & (~\m6_data_i[7]  | ~\new_[17241]_ );
  assign \new_[9099]_  = (~\m2_addr_i[7]  | ~\new_[16292]_ ) & (~\m1_addr_i[7]  | ~\new_[18167]_ );
  assign \new_[9100]_  = ~\new_[19381]_  | ~\new_[12252]_ ;
  assign \new_[9101]_  = (~\m2_addr_i[6]  | ~\new_[16292]_ ) & (~\m1_addr_i[6]  | ~\new_[18167]_ );
  assign \new_[9102]_  = ~\new_[28729]_  & (~\new_[14382]_  | ~\new_[22753]_ );
  assign \new_[9103]_  = (~\m2_addr_i[5]  | ~\new_[16292]_ ) & (~\m1_addr_i[5]  | ~\new_[18167]_ );
  assign \new_[9104]_  = (~\m2_addr_i[4]  | ~\new_[18080]_ ) & (~\m1_addr_i[4]  | ~\new_[18167]_ );
  assign \new_[9105]_  = ~\new_[18407]_  | ~\new_[12257]_ ;
  assign \new_[9106]_  = (~\new_[31399]_  | ~\new_[16292]_ ) & (~\m1_addr_i[3]  | ~\new_[18890]_ );
  assign \new_[9107]_  = (~\m2_addr_i[2]  | ~\new_[16292]_ ) & (~\m1_addr_i[2]  | ~\new_[19621]_ );
  assign \new_[9108]_  = (~\m7_addr_i[1]  | ~\new_[16295]_ ) & (~\m0_addr_i[1]  | ~\new_[19643]_ );
  assign \new_[9109]_  = ~\new_[30412]_  | (~\new_[14385]_  & ~\new_[24885]_ );
  assign \new_[9110]_  = ~\new_[28868]_  & (~\new_[14386]_  | ~\new_[19382]_ );
  assign \new_[9111]_  = (~\m7_addr_i[0]  | ~\new_[16295]_ ) & (~\m0_addr_i[0]  | ~\new_[19643]_ );
  assign \new_[9112]_  = (~\m2_addr_i[0]  | ~\new_[18080]_ ) & (~\m1_addr_i[0]  | ~\new_[18167]_ );
  assign \new_[9113]_  = ~\new_[14387]_  | ~\new_[28091]_  | ~\new_[22838]_ ;
  assign \new_[9114]_  = (~\m5_sel_i[3]  | ~\new_[17204]_ ) & (~\m6_sel_i[3]  | ~\new_[16287]_ );
  assign \new_[9115]_  = (~\m2_sel_i[3]  | ~\new_[18080]_ ) & (~\m1_sel_i[3]  | ~\new_[18167]_ );
  assign \new_[9116]_  = ~\new_[28925]_  & (~\new_[14389]_  | ~\new_[22746]_ );
  assign \new_[9117]_  = (~\m5_sel_i[2]  | ~\new_[17204]_ ) & (~\m6_sel_i[2]  | ~\new_[16287]_ );
  assign \new_[9118]_  = (~\m2_sel_i[2]  | ~\new_[16292]_ ) & (~\m1_sel_i[2]  | ~\new_[19621]_ );
  assign \new_[9119]_  = (~\m7_sel_i[2]  | ~\new_[16295]_ ) & (~\m0_sel_i[2]  | ~\new_[18204]_ );
  assign n7644 = (~\new_[14469]_  & ~rst_i) | (~\new_[30813]_  & ~\new_[31888]_ );
  assign \new_[9121]_  = (~\m7_sel_i[1]  | ~\new_[16295]_ ) & (~\m0_sel_i[1]  | ~\new_[18204]_ );
  assign \new_[9122]_  = ~\new_[20370]_  | ~\new_[12264]_ ;
  assign \new_[9123]_  = ~\new_[20372]_  | ~\new_[12267]_ ;
  assign \new_[9124]_  = (~\m7_sel_i[0]  | ~\new_[16295]_ ) & (~\m0_sel_i[0]  | ~\new_[19643]_ );
  assign \new_[9125]_  = (~\m2_sel_i[0]  | ~\new_[18080]_ ) & (~\m1_sel_i[0]  | ~\new_[18167]_ );
  assign \new_[9126]_  = (~m2_we_i | ~\new_[16292]_ ) & (~m1_we_i | ~\new_[18890]_ );
  assign \new_[9127]_  = ~\new_[28018]_  & (~\new_[14396]_  | ~\new_[22762]_ );
  assign \new_[9128]_  = (~\m7_data_i[31]  | ~\new_[18111]_ ) & (~\m0_data_i[31]  | ~\new_[18027]_ );
  assign n7619 = (~\new_[14475]_  & ~rst_i) | (~\new_[31173]_  & ~\new_[31576]_ );
  assign \new_[9130]_  = (~\m4_data_i[30]  | ~\new_[16307]_ ) & (~\m3_data_i[30]  | ~\new_[17249]_ );
  assign \new_[9131]_  = ~\new_[21305]_  | ~\new_[12271]_ ;
  assign \new_[9132]_  = ~\new_[29321]_  & (~\new_[14398]_  | ~\new_[20438]_ );
  assign n7614 = (~\new_[14478]_  & ~rst_i) | (~\new_[31117]_  & ~\new_[31759]_ );
  assign \new_[9134]_  = (~\m4_data_i[26]  | ~\new_[16308]_ ) & (~\m3_data_i[26]  | ~\new_[18850]_ );
  assign \new_[9135]_  = ~\new_[30345]_  | (~\new_[14400]_  & ~\new_[24964]_ );
  assign \new_[9136]_  = (~\m7_data_i[26]  | ~\new_[18111]_ ) & (~\m0_data_i[26]  | ~\new_[18027]_ );
  assign \new_[9137]_  = ~\new_[29304]_  & (~\new_[14401]_  | ~\new_[19427]_ );
  assign \new_[9138]_  = (~\m7_data_i[25]  | ~\new_[18111]_ ) & (~\m0_data_i[25]  | ~\new_[18027]_ );
  assign \new_[9139]_  = (~\m4_data_i[25]  | ~\new_[16307]_ ) & (~\m3_data_i[25]  | ~\new_[18850]_ );
  assign \new_[9140]_  = (~\m4_data_i[24]  | ~\new_[16307]_ ) & (~\m3_data_i[24]  | ~\new_[18850]_ );
  assign \new_[9141]_  = (~\m4_data_i[22]  | ~\new_[16307]_ ) & (~\m3_data_i[22]  | ~\new_[18850]_ );
  assign \new_[9142]_  = ~\new_[28656]_  | (~\new_[14407]_  & ~\new_[24989]_ );
  assign \new_[9143]_  = ~\new_[27832]_  & (~\new_[14408]_  | ~\new_[20459]_ );
  assign \new_[9144]_  = (~\m4_data_i[21]  | ~\new_[13493]_ ) & (~\m3_data_i[21]  | ~\new_[17249]_ );
  assign \new_[9145]_  = ~\new_[20378]_  | ~\new_[12279]_ ;
  assign \new_[9146]_  = (~\m7_data_i[20]  | ~\new_[18111]_ ) & (~\m0_data_i[20]  | ~\new_[18027]_ );
  assign \new_[9147]_  = (~\m4_data_i[20]  | ~\new_[16307]_ ) & (~\m3_data_i[20]  | ~\new_[17249]_ );
  assign \new_[9148]_  = (~\m4_data_i[19]  | ~\new_[16308]_ ) & (~\m3_data_i[19]  | ~\new_[17249]_ );
  assign \new_[9149]_  = (~\m7_data_i[18]  | ~\new_[18111]_ ) & (~\m0_data_i[18]  | ~\new_[18027]_ );
  assign n7639 = (~\new_[14481]_  & ~rst_i) | (~\new_[31101]_  & ~\new_[31830]_ );
  assign \new_[9151]_  = (~\m5_data_i[18]  | ~\new_[16278]_ ) & (~\m6_data_i[18]  | ~\new_[18035]_ );
  assign \new_[9152]_  = (~\m7_data_i[17]  | ~\new_[18111]_ ) & (~\m0_data_i[17]  | ~\new_[18027]_ );
  assign \new_[9153]_  = ~\new_[19384]_  | ~\new_[12284]_ ;
  assign \new_[9154]_  = (~\m4_data_i[16]  | ~\new_[16308]_ ) & (~\m3_data_i[16]  | ~\new_[18850]_ );
  assign \new_[9155]_  = (~\m7_data_i[15]  | ~\new_[18111]_ ) & (~\m0_data_i[15]  | ~\new_[18027]_ );
  assign \new_[9156]_  = (~\m4_data_i[14]  | ~\new_[13493]_ ) & (~\m3_data_i[14]  | ~\new_[17249]_ );
  assign \new_[9157]_  = ~\new_[27992]_  | (~\new_[14413]_  & ~\new_[26518]_ );
  assign \new_[9158]_  = (~\m4_data_i[13]  | ~\new_[16308]_ ) & (~\m3_data_i[13]  | ~\new_[18850]_ );
  assign \new_[9159]_  = ~\new_[27862]_  & (~\new_[14414]_  | ~\new_[21137]_ );
  assign \new_[9160]_  = (~\m4_data_i[12]  | ~\new_[16308]_ ) & (~\m3_data_i[12]  | ~\new_[18850]_ );
  assign \new_[9161]_  = ~\new_[29343]_  & (~\new_[14417]_  | ~\new_[22722]_ );
  assign \new_[9162]_  = (~\m7_data_i[11]  | ~\new_[18111]_ ) & (~\m0_data_i[11]  | ~\new_[18027]_ );
  assign \new_[9163]_  = (~\m4_data_i[11]  | ~\new_[16307]_ ) & (~\m3_data_i[11]  | ~\new_[18850]_ );
  assign \new_[9164]_  = (~\m4_data_i[10]  | ~\new_[16308]_ ) & (~\m3_data_i[10]  | ~\new_[18850]_ );
  assign \new_[9165]_  = ~\new_[28321]_  & (~\new_[14420]_  | ~\new_[19432]_ );
  assign \new_[9166]_  = (~\m7_data_i[9]  | ~\new_[18111]_ ) & (~\m0_data_i[9]  | ~\new_[18027]_ );
  assign \new_[9167]_  = ~\new_[20385]_  | ~\new_[12291]_ ;
  assign \new_[9168]_  = ~\new_[28657]_  & (~\new_[14421]_  | ~\new_[22787]_ );
  assign \new_[9169]_  = (~\m4_data_i[7]  | ~\new_[16307]_ ) & (~\m3_data_i[7]  | ~\new_[17249]_ );
  assign n7624 = (~\new_[14491]_  & ~rst_i) | (~\new_[30965]_  & ~\new_[31698]_ );
  assign \new_[9171]_  = (~\m4_data_i[6]  | ~\new_[16307]_ ) & (~\m3_data_i[6]  | ~\new_[17249]_ );
  assign \new_[9172]_  = (~\m7_data_i[6]  | ~\new_[18111]_ ) & (~\m0_data_i[6]  | ~\new_[18027]_ );
  assign \new_[9173]_  = (~\m4_data_i[5]  | ~\new_[16307]_ ) & (~\m3_data_i[5]  | ~\new_[17249]_ );
  assign \new_[9174]_  = (~\m5_data_i[5]  | ~\new_[16278]_ ) & (~\m6_data_i[5]  | ~\new_[18036]_ );
  assign \new_[9175]_  = (~\m7_data_i[5]  | ~\new_[18111]_ ) & (~\m0_data_i[5]  | ~\new_[18027]_ );
  assign \new_[9176]_  = ~\new_[28805]_  & (~\new_[14428]_  | ~\new_[21392]_ );
  assign \new_[9177]_  = (~\m7_data_i[4]  | ~\new_[18111]_ ) & (~\m0_data_i[4]  | ~\new_[18027]_ );
  assign \new_[9178]_  = (~\m4_data_i[4]  | ~\new_[16307]_ ) & (~\m3_data_i[4]  | ~\new_[18850]_ );
  assign \new_[9179]_  = (~\m5_data_i[3]  | ~\new_[16278]_ ) & (~\m6_data_i[3]  | ~\new_[18035]_ );
  assign \new_[9180]_  = (~\m1_data_i[9]  | ~\new_[17277]_ ) & (~\m0_data_i[9]  | ~\new_[16279]_ );
  assign \new_[9181]_  = ~\new_[20380]_  | ~\new_[12299]_ ;
  assign \new_[9182]_  = (~\m7_data_i[3]  | ~\new_[18111]_ ) & (~\m0_data_i[3]  | ~\new_[18027]_ );
  assign \new_[9183]_  = (~\m4_data_i[3]  | ~\new_[16307]_ ) & (~\m3_data_i[3]  | ~\new_[17249]_ );
  assign \new_[9184]_  = (~\m4_data_i[2]  | ~\new_[16307]_ ) & (~\m3_data_i[2]  | ~\new_[17249]_ );
  assign \new_[9185]_  = ~\new_[21298]_  | ~\new_[12302]_ ;
  assign \new_[9186]_  = (~\m7_data_i[1]  | ~\new_[18111]_ ) & (~\m0_data_i[1]  | ~\new_[18027]_ );
  assign \new_[9187]_  = (~\m4_data_i[1]  | ~\new_[13493]_ ) & (~\m3_data_i[1]  | ~\new_[17249]_ );
  assign \new_[9188]_  = (~\m4_data_i[0]  | ~\new_[16308]_ ) & (~\m3_data_i[0]  | ~\new_[18850]_ );
  assign n7634 = (~\new_[14455]_  & ~rst_i) | (~\new_[30830]_  & ~\new_[31678]_ );
  assign \new_[9190]_  = ~\new_[21325]_  | ~\new_[12311]_ ;
  assign \new_[9191]_  = (~\new_[16308]_  | ~\m4_addr_i[31] ) & (~\new_[17249]_  | ~\m3_addr_i[31] );
  assign \new_[9192]_  = (~\new_[19559]_  | ~\m6_addr_i[30] ) & (~\new_[16278]_  | ~\new_[31147]_ );
  assign \new_[9193]_  = (~\new_[18111]_  | ~\new_[31885]_ ) & (~\new_[18027]_  | ~\new_[31292]_ );
  assign \new_[9194]_  = (~\new_[16307]_  | ~\m4_addr_i[30] ) & (~\new_[17249]_  | ~\m3_addr_i[30] );
  assign \new_[9195]_  = (~\new_[13493]_  | ~\m4_addr_i[29] ) & (~\new_[17249]_  | ~\m3_addr_i[29] );
  assign \new_[9196]_  = (~\new_[18111]_  | ~\new_[31531]_ ) & (~\new_[18027]_  | ~\new_[31481]_ );
  assign n7629 = (~\new_[13136]_  & ~rst_i) | (~\new_[30516]_  & ~\new_[31804]_ );
  assign \new_[9198]_  = ~\new_[20393]_  | ~\new_[12318]_ ;
  assign \new_[9199]_  = (~\m1_data_i[31]  | ~\new_[17277]_ ) & (~\m0_data_i[31]  | ~\new_[16280]_ );
  assign \new_[9200]_  = (~\new_[16307]_  | ~\m4_addr_i[28] ) & (~\new_[17249]_  | ~\m3_addr_i[28] );
  assign \new_[9201]_  = (~\new_[19559]_  | ~\m6_addr_i[27] ) & (~\new_[16278]_  | ~\m5_addr_i[27] );
  assign \new_[9202]_  = (~\new_[18111]_  | ~\m7_addr_i[27] ) & (~\new_[18027]_  | ~\m0_addr_i[27] );
  assign \new_[9203]_  = ~\new_[26819]_  & (~\new_[14394]_  | ~\new_[20430]_ );
  assign \new_[9204]_  = (~\new_[16307]_  | ~\m4_addr_i[27] ) & (~\new_[18850]_  | ~\m3_addr_i[27] );
  assign \new_[9205]_  = (~\new_[13493]_  | ~\m4_addr_i[26] ) & (~\new_[17249]_  | ~\m3_addr_i[26] );
  assign \new_[9206]_  = (~\new_[18111]_  | ~\m7_addr_i[26] ) & (~\new_[18027]_  | ~\m0_addr_i[26] );
  assign \new_[9207]_  = (~\new_[13493]_  | ~\m4_addr_i[25] ) & (~\new_[17249]_  | ~\m3_addr_i[25] );
  assign \new_[9208]_  = (~\new_[18111]_  | ~\m7_addr_i[25] ) & (~\new_[18027]_  | ~\m0_addr_i[25] );
  assign \new_[9209]_  = (~\new_[13493]_  | ~\m4_addr_i[24] ) & (~\new_[17249]_  | ~\m3_addr_i[24] );
  assign \new_[9210]_  = (~\new_[18111]_  | ~\m7_addr_i[24] ) & (~\new_[18027]_  | ~\m0_addr_i[24] );
  assign \new_[9211]_  = (~\m7_addr_i[23]  | ~\new_[18111]_ ) & (~\m0_addr_i[23]  | ~\new_[18027]_ );
  assign \new_[9212]_  = ~\new_[27466]_  & (~\new_[13491]_  | ~\new_[20631]_ );
  assign \new_[9213]_  = ~\new_[27844]_  & (~\new_[13189]_  | ~\new_[21489]_ );
  assign \new_[9214]_  = (~\m1_data_i[30]  | ~\new_[17277]_ ) & (~\m0_data_i[30]  | ~\new_[16280]_ );
  assign \new_[9215]_  = (~\m4_addr_i[22]  | ~\new_[16307]_ ) & (~\m3_addr_i[22]  | ~\new_[17249]_ );
  assign \new_[9216]_  = ~\new_[27917]_  & (~\new_[13173]_  | ~\new_[21479]_ );
  assign \new_[9217]_  = ~\new_[29287]_  & (~\new_[14464]_  | ~\new_[24258]_ );
  assign \new_[9218]_  = (~\m1_data_i[29]  | ~\new_[17277]_ ) & (~\m0_data_i[29]  | ~\new_[16280]_ );
  assign \new_[9219]_  = ~\new_[27830]_  & (~\new_[14033]_  | ~\new_[24373]_ );
  assign \new_[9220]_  = ~\new_[27849]_  & (~\new_[13846]_  | ~\new_[24270]_ );
  assign \new_[9221]_  = ~\new_[26601]_  & (~\new_[13655]_  | ~\new_[21549]_ );
  assign \new_[9222]_  = ~\new_[27913]_  & (~\new_[13608]_  | ~\new_[23157]_ );
  assign \new_[9223]_  = (~\m4_addr_i[21]  | ~\new_[16307]_ ) & (~\m3_addr_i[21]  | ~\new_[17249]_ );
  assign \new_[9224]_  = ~\new_[26990]_  & (~\new_[13571]_  | ~\new_[21529]_ );
  assign \new_[9225]_  = (~\m4_addr_i[20]  | ~\new_[16307]_ ) & (~\m3_addr_i[20]  | ~\new_[17249]_ );
  assign \new_[9226]_  = (~\m4_addr_i[19]  | ~\new_[16307]_ ) & (~\m3_addr_i[19]  | ~\new_[17249]_ );
  assign \new_[9227]_  = (~\m7_addr_i[19]  | ~\new_[18111]_ ) & (~\m0_addr_i[19]  | ~\new_[18027]_ );
  assign \new_[9228]_  = (~\m7_addr_i[18]  | ~\new_[18111]_ ) & (~\m0_addr_i[18]  | ~\new_[18027]_ );
  assign \new_[9229]_  = (~\m4_addr_i[18]  | ~\new_[16308]_ ) & (~\m3_addr_i[18]  | ~\new_[18850]_ );
  assign \new_[9230]_  = (~\m4_addr_i[17]  | ~\new_[13493]_ ) & (~\m3_addr_i[17]  | ~\new_[17249]_ );
  assign \new_[9231]_  = (~\m4_addr_i[16]  | ~\new_[13493]_ ) & (~\m3_addr_i[16]  | ~\new_[17249]_ );
  assign \new_[9232]_  = (~\m1_data_i[27]  | ~\new_[17277]_ ) & (~\m0_data_i[27]  | ~\new_[16280]_ );
  assign \new_[9233]_  = (~\m4_addr_i[15]  | ~\new_[16308]_ ) & (~\m3_addr_i[15]  | ~\new_[17249]_ );
  assign \new_[9234]_  = (~\m7_addr_i[15]  | ~\new_[18111]_ ) & (~\m0_addr_i[15]  | ~\new_[18027]_ );
  assign \new_[9235]_  = (~\m7_addr_i[14]  | ~\new_[18111]_ ) & (~\m0_addr_i[14]  | ~\new_[18027]_ );
  assign \new_[9236]_  = (~\m4_addr_i[14]  | ~\new_[16307]_ ) & (~\m3_addr_i[14]  | ~\new_[17249]_ );
  assign \new_[9237]_  = (~\m4_addr_i[13]  | ~\new_[13493]_ ) & (~\m3_addr_i[13]  | ~\new_[17249]_ );
  assign \new_[9238]_  = (~\m7_addr_i[13]  | ~\new_[18111]_ ) & (~\m0_addr_i[13]  | ~\new_[18027]_ );
  assign \new_[9239]_  = (~\m4_addr_i[12]  | ~\new_[16308]_ ) & (~\m3_addr_i[12]  | ~\new_[18850]_ );
  assign \new_[9240]_  = \new_[12387]_  & \new_[29187]_ ;
  assign \new_[9241]_  = (~\m7_addr_i[12]  | ~\new_[18111]_ ) & (~\m0_addr_i[12]  | ~\new_[18027]_ );
  assign \new_[9242]_  = (~\m7_addr_i[11]  | ~\new_[18111]_ ) & (~\m0_addr_i[11]  | ~\new_[18027]_ );
  assign \new_[9243]_  = \new_[12396]_  & \new_[28261]_ ;
  assign \new_[9244]_  = (~\m5_addr_i[16]  | ~\new_[18004]_ ) & (~\m6_addr_i[16]  | ~\new_[17241]_ );
  assign \new_[9245]_  = (~\m7_addr_i[10]  | ~\new_[18111]_ ) & (~\m0_addr_i[10]  | ~\new_[18027]_ );
  assign \new_[9246]_  = (~\m4_addr_i[10]  | ~\new_[16307]_ ) & (~\m3_addr_i[10]  | ~\new_[17249]_ );
  assign \new_[9247]_  = (~\m4_addr_i[9]  | ~\new_[16308]_ ) & (~\m3_addr_i[9]  | ~\new_[17249]_ );
  assign \new_[9248]_  = (~\m7_addr_i[9]  | ~\new_[18111]_ ) & (~\m0_addr_i[9]  | ~\new_[18027]_ );
  assign \new_[9249]_  = \new_[12421]_  & \new_[28822]_ ;
  assign \new_[9250]_  = (~\m7_addr_i[8]  | ~\new_[18111]_ ) & (~\m0_addr_i[8]  | ~\new_[18027]_ );
  assign \new_[9251]_  = (~\m1_data_i[25]  | ~\new_[17277]_ ) & (~\m0_data_i[25]  | ~\new_[16279]_ );
  assign \new_[9252]_  = (~\m7_addr_i[7]  | ~\new_[18111]_ ) & (~\m0_addr_i[7]  | ~\new_[18027]_ );
  assign \new_[9253]_  = (~\m4_addr_i[7]  | ~\new_[16307]_ ) & (~\m3_addr_i[7]  | ~\new_[17249]_ );
  assign \new_[9254]_  = (~\m4_addr_i[6]  | ~\new_[16308]_ ) & (~\m3_addr_i[6]  | ~\new_[18850]_ );
  assign \new_[9255]_  = (~\m1_data_i[24]  | ~\new_[17277]_ ) & (~\m0_data_i[24]  | ~\new_[16279]_ );
  assign \new_[9256]_  = (~\m4_addr_i[5]  | ~\new_[16307]_ ) & (~\m3_addr_i[5]  | ~\new_[17249]_ );
  assign \new_[9257]_  = (~\m7_addr_i[4]  | ~\new_[18111]_ ) & (~\m0_addr_i[4]  | ~\new_[18027]_ );
  assign \new_[9258]_  = (~\m1_data_i[23]  | ~\new_[17277]_ ) & (~\m0_data_i[23]  | ~\new_[16280]_ );
  assign \new_[9259]_  = (~\m4_addr_i[2]  | ~\new_[13493]_ ) & (~\m3_addr_i[2]  | ~\new_[17249]_ );
  assign \new_[9260]_  = (~\m7_addr_i[1]  | ~\new_[18111]_ ) & (~\m0_addr_i[1]  | ~\new_[18027]_ );
  assign \new_[9261]_  = (~\m5_addr_i[1]  | ~\new_[16278]_ ) & (~\m6_addr_i[1]  | ~\new_[18035]_ );
  assign \new_[9262]_  = ~\new_[16652]_  | ~\new_[15864]_  | ~\new_[16650]_  | ~\new_[16651]_ ;
  assign \new_[9263]_  = (~\m4_addr_i[1]  | ~\new_[16307]_ ) & (~\m3_addr_i[1]  | ~\new_[18850]_ );
  assign \new_[9264]_  = (~\m1_data_i[22]  | ~\new_[17277]_ ) & (~\m0_data_i[22]  | ~\new_[16280]_ );
  assign \new_[9265]_  = (~\m4_addr_i[0]  | ~\new_[16307]_ ) & (~\m3_addr_i[0]  | ~\new_[17249]_ );
  assign \new_[9266]_  = (~\m5_addr_i[0]  | ~\new_[16278]_ ) & (~\m6_addr_i[0]  | ~\new_[18035]_ );
  assign \new_[9267]_  = (~\m4_sel_i[3]  | ~\new_[16308]_ ) & (~\m3_sel_i[3]  | ~\new_[18850]_ );
  assign \new_[9268]_  = (~\m7_sel_i[2]  | ~\new_[18111]_ ) & (~\m0_sel_i[2]  | ~\new_[18027]_ );
  assign \new_[9269]_  = (~\m4_sel_i[2]  | ~\new_[16308]_ ) & (~\m3_sel_i[2]  | ~\new_[18850]_ );
  assign \new_[9270]_  = (~\m4_sel_i[1]  | ~\new_[16307]_ ) & (~\m3_sel_i[1]  | ~\new_[17249]_ );
  assign \new_[9271]_  = (~\m1_data_i[21]  | ~\new_[17277]_ ) & (~\m0_data_i[21]  | ~\new_[16280]_ );
  assign \new_[9272]_  = (~\m7_sel_i[1]  | ~\new_[18111]_ ) & (~\m0_sel_i[1]  | ~\new_[18027]_ );
  assign \new_[9273]_  = ~\new_[15873]_  | ~\new_[16664]_  | ~\new_[17542]_  | ~\new_[17543]_ ;
  assign \new_[9274]_  = ~\new_[16665]_  | ~\new_[16666]_  | ~\new_[15874]_  | ~\new_[14477]_ ;
  assign \new_[9275]_  = (~\m4_sel_i[0]  | ~\new_[16308]_ ) & (~\m3_sel_i[0]  | ~\new_[18850]_ );
  assign \new_[9276]_  = (~\m5_sel_i[0]  | ~\new_[16278]_ ) & (~\m6_sel_i[0]  | ~\new_[18038]_ );
  assign \new_[9277]_  = (~m7_we_i | ~\new_[18111]_ ) & (~m0_we_i | ~\new_[18027]_ );
  assign \new_[9278]_  = (~m4_we_i | ~\new_[13493]_ ) & (~m3_we_i | ~\new_[17249]_ );
  assign \new_[9279]_  = ~\new_[15878]_  | ~\new_[16673]_  | ~\new_[16671]_  | ~\new_[16672]_ ;
  assign \new_[9280]_  = (~\m1_data_i[20]  | ~\new_[17277]_ ) & (~\m0_data_i[20]  | ~\new_[16280]_ );
  assign \new_[9281]_  = ~\new_[15881]_  | ~\new_[15883]_  | ~\new_[17545]_  | ~\new_[15880]_ ;
  assign \new_[9282]_  = (~\m1_data_i[19]  | ~\new_[17277]_ ) & (~\m0_data_i[19]  | ~\new_[16280]_ );
  assign \new_[9283]_  = ~\new_[15889]_  | ~\new_[15891]_  | ~\new_[15909]_  | ~\new_[16685]_ ;
  assign \new_[9284]_  = (~\m1_data_i[18]  | ~\new_[17277]_ ) & (~\m0_data_i[18]  | ~\new_[16280]_ );
  assign \new_[9285]_  = ~\new_[16688]_  | ~\new_[15894]_  | ~\new_[17541]_  | ~\new_[17557]_ ;
  assign \new_[9286]_  = ~\new_[15898]_  | ~\new_[14506]_  | ~\new_[15895]_  | ~\new_[15897]_ ;
  assign \new_[9287]_  = ~\new_[12007]_  | ~\new_[28541]_ ;
  assign \new_[9288]_  = (~\m1_data_i[17]  | ~\new_[17277]_ ) & (~\m0_data_i[17]  | ~\new_[16280]_ );
  assign \new_[9289]_  = ~\new_[14512]_  | ~\new_[15903]_  | ~\new_[16697]_  | ~\new_[16698]_ ;
  assign \new_[9290]_  = (~\m1_data_i[16]  | ~\new_[17277]_ ) & (~\m0_data_i[16]  | ~\new_[16279]_ );
  assign \new_[9291]_  = (~\m1_data_i[15]  | ~\new_[17277]_ ) & (~\m0_data_i[15]  | ~\new_[16280]_ );
  assign \new_[9292]_  = ~\new_[15912]_  | ~\new_[14519]_  | ~\new_[14518]_  | ~\new_[15911]_ ;
  assign \new_[9293]_  = ~\new_[28319]_  & (~\new_[14370]_  | ~\new_[22819]_ );
  assign \new_[9294]_  = ~\new_[24553]_  & (~\new_[14377]_  | ~\new_[21412]_ );
  assign \new_[9295]_  = ~\new_[28648]_  & (~\new_[14383]_  | ~\new_[20426]_ );
  assign \new_[9296]_  = ~\new_[28715]_  & (~\new_[14384]_  | ~\new_[21378]_ );
  assign \new_[9297]_  = ~\new_[28869]_  & (~\new_[14388]_  | ~\new_[21387]_ );
  assign \new_[9298]_  = ~\new_[28059]_  & (~\new_[14399]_  | ~\new_[20420]_ );
  assign \new_[9299]_  = ~\new_[27998]_  & (~\new_[14404]_  | ~\new_[22706]_ );
  assign \new_[9300]_  = ~\new_[29247]_  & (~\new_[14409]_  | ~\new_[20417]_ );
  assign \new_[9301]_  = (~\m1_data_i[8]  | ~\new_[17277]_ ) & (~\m0_data_i[8]  | ~\new_[16279]_ );
  assign \new_[9302]_  = ~\new_[28487]_  & (~\new_[14411]_  | ~\new_[24225]_ );
  assign \new_[9303]_  = ~\new_[29361]_  & (~\new_[14416]_  | ~\new_[20435]_ );
  assign \new_[9304]_  = ~\new_[28190]_  & (~\new_[14426]_  | ~\new_[22632]_ );
  assign \new_[9305]_  = ~\new_[29148]_  & (~\new_[14432]_  | ~\new_[21434]_ );
  assign \new_[9306]_  = ~\new_[26503]_  & (~\new_[14436]_  | ~\new_[22697]_ );
  assign \new_[9307]_  = (~\m1_data_i[5]  | ~\new_[17277]_ ) & (~\m0_data_i[5]  | ~\new_[16280]_ );
  assign \new_[9308]_  = (~\m1_data_i[4]  | ~\new_[17277]_ ) & (~\m0_data_i[4]  | ~\new_[16279]_ );
  assign \new_[9309]_  = (~\m1_data_i[1]  | ~\new_[17277]_ ) & (~\m0_data_i[1]  | ~\new_[16279]_ );
  assign \new_[9310]_  = ~\new_[13036]_  & ~\new_[14625]_ ;
  assign \new_[9311]_  = (~\new_[17239]_  | ~\m7_addr_i[31] ) & (~\new_[16280]_  | ~\m0_addr_i[31] );
  assign \new_[9312]_  = ~\new_[13038]_  & ~\new_[14677]_ ;
  assign \new_[9313]_  = (~\new_[17240]_  | ~\new_[30577]_ ) & (~\new_[16280]_  | ~\new_[30957]_ );
  assign \new_[9314]_  = ~\new_[28762]_  | ~\new_[13091]_  | ~\new_[30343]_ ;
  assign \new_[9315]_  = (~\new_[17239]_  | ~\m7_addr_i[27] ) & (~\new_[16280]_  | ~\m0_addr_i[27] );
  assign \new_[9316]_  = (~\new_[17239]_  | ~\m7_addr_i[26] ) & (~\new_[16280]_  | ~\m0_addr_i[26] );
  assign \new_[9317]_  = ~\new_[14586]_  | ~\new_[14594]_  | ~\new_[14596]_  | ~\new_[14593]_ ;
  assign \new_[9318]_  = ~\new_[10549]_ ;
  assign \new_[9319]_  = (~\m1_addr_i[23]  | ~\new_[17277]_ ) & (~\m0_addr_i[23]  | ~\new_[16280]_ );
  assign \new_[9320]_  = (~\m1_addr_i[21]  | ~\new_[17277]_ ) & (~\m0_addr_i[21]  | ~\new_[16280]_ );
  assign \new_[9321]_  = (~\m1_addr_i[18]  | ~\new_[17277]_ ) & (~\m0_addr_i[18]  | ~\new_[16280]_ );
  assign \new_[9322]_  = (~\m1_addr_i[17]  | ~\new_[17277]_ ) & (~\m0_addr_i[17]  | ~\new_[16280]_ );
  assign \new_[9323]_  = (~\m1_addr_i[16]  | ~\new_[18192]_ ) & (~\m0_addr_i[16]  | ~\new_[16279]_ );
  assign \new_[9324]_  = (~\new_[17229]_  | ~\m6_addr_i[31] ) & (~\new_[18015]_  | ~\new_[31001]_ );
  assign \new_[9325]_  = (~\new_[17229]_  | ~\m6_addr_i[30] ) & (~\new_[18015]_  | ~\new_[31147]_ );
  assign \new_[9326]_  = (~\m1_addr_i[13]  | ~\new_[17277]_ ) & (~\m0_addr_i[13]  | ~\new_[16279]_ );
  assign \new_[9327]_  = (~\new_[17229]_  | ~\m6_addr_i[28] ) & (~\new_[19547]_  | ~\new_[31276]_ );
  assign \new_[9328]_  = (~\new_[17229]_  | ~\m6_addr_i[27] ) & (~\new_[19547]_  | ~\m5_addr_i[27] );
  assign \new_[9329]_  = (~\m1_addr_i[12]  | ~\new_[17277]_ ) & (~\m0_addr_i[12]  | ~\new_[16280]_ );
  assign \new_[9330]_  = (~\new_[17229]_  | ~\m6_addr_i[26] ) & (~\new_[19547]_  | ~\m5_addr_i[26] );
  assign \new_[9331]_  = (~\new_[17229]_  | ~\m6_addr_i[25] ) & (~\new_[18015]_  | ~\m5_addr_i[25] );
  assign \new_[9332]_  = (~\new_[17229]_  | ~\m6_addr_i[24] ) & (~\new_[18015]_  | ~\m5_addr_i[24] );
  assign \new_[9333]_  = (~\m1_addr_i[10]  | ~\new_[17277]_ ) & (~\m0_addr_i[10]  | ~\new_[16280]_ );
  assign \new_[9334]_  = ~\new_[12020]_  & (~\new_[14213]_  | ~\new_[26761]_ );
  assign \new_[9335]_  = (~\m1_addr_i[7]  | ~\new_[17277]_ ) & (~\m0_addr_i[7]  | ~\new_[16280]_ );
  assign \new_[9336]_  = (~\m1_addr_i[6]  | ~\new_[17277]_ ) & (~\m0_addr_i[6]  | ~\new_[16280]_ );
  assign \new_[9337]_  = (~\m1_addr_i[4]  | ~\new_[17277]_ ) & (~\m0_addr_i[4]  | ~\new_[16280]_ );
  assign \new_[9338]_  = (~\m5_data_i[31]  | ~\new_[18004]_ ) & (~\m6_data_i[31]  | ~\new_[18836]_ );
  assign \new_[9339]_  = (~\m5_data_i[30]  | ~\new_[18004]_ ) & (~\m6_data_i[30]  | ~\new_[17241]_ );
  assign \new_[9340]_  = (~\m1_addr_i[0]  | ~\new_[17277]_ ) & (~\m0_addr_i[0]  | ~\new_[16280]_ );
  assign \new_[9341]_  = (~\m5_data_i[28]  | ~\new_[18004]_ ) & (~\m6_data_i[28]  | ~\new_[17241]_ );
  assign \new_[9342]_  = (~\m5_data_i[27]  | ~\new_[18004]_ ) & (~\m6_data_i[27]  | ~\new_[18836]_ );
  assign \new_[9343]_  = (~\m5_data_i[26]  | ~\new_[18004]_ ) & (~\m6_data_i[26]  | ~\new_[18836]_ );
  assign \new_[9344]_  = (~\m1_sel_i[3]  | ~\new_[17277]_ ) & (~\m0_sel_i[3]  | ~\new_[16280]_ );
  assign \new_[9345]_  = (~\m5_data_i[25]  | ~\new_[18004]_ ) & (~\m6_data_i[25]  | ~\new_[18836]_ );
  assign \new_[9346]_  = (~\m1_sel_i[2]  | ~\new_[17277]_ ) & (~\m0_sel_i[2]  | ~\new_[16280]_ );
  assign \new_[9347]_  = (~\m5_data_i[21]  | ~\new_[18004]_ ) & (~\m6_data_i[21]  | ~\new_[17241]_ );
  assign \new_[9348]_  = (~\m5_data_i[19]  | ~\new_[18004]_ ) & (~\m6_data_i[19]  | ~\new_[18836]_ );
  assign \new_[9349]_  = (~\m5_data_i[17]  | ~\new_[18004]_ ) & (~\m6_data_i[17]  | ~\new_[17241]_ );
  assign \new_[9350]_  = (~\m1_sel_i[0]  | ~\new_[17277]_ ) & (~\m0_sel_i[0]  | ~\new_[16280]_ );
  assign \new_[9351]_  = (~\m7_data_i[15]  | ~\new_[16296]_ ) & (~\m0_data_i[15]  | ~\new_[20545]_ );
  assign \new_[9352]_  = (~\m5_data_i[15]  | ~\new_[18004]_ ) & (~\m6_data_i[15]  | ~\new_[17241]_ );
  assign \new_[9353]_  = (~\m5_data_i[14]  | ~\new_[18004]_ ) & (~\m6_data_i[14]  | ~\new_[17241]_ );
  assign \new_[9354]_  = (~\m5_data_i[13]  | ~\new_[18004]_ ) & (~\m6_data_i[13]  | ~\new_[17241]_ );
  assign \new_[9355]_  = (~m1_we_i | ~\new_[17277]_ ) & (~m0_we_i | ~\new_[16280]_ );
  assign \new_[9356]_  = (~\m5_data_i[11]  | ~\new_[18004]_ ) & (~\m6_data_i[11]  | ~\new_[17241]_ );
  assign \new_[9357]_  = (~\new_[31726]_  | ~\new_[18111]_ ) & (~\m0_addr_i[3]  | ~\new_[18027]_ );
  assign \new_[9358]_  = (~\m7_data_i[10]  | ~\new_[16296]_ ) & (~\m0_data_i[10]  | ~\new_[20545]_ );
  assign \new_[9359]_  = (~\m5_data_i[9]  | ~\new_[18004]_ ) & (~\m6_data_i[9]  | ~\new_[18836]_ );
  assign \new_[9360]_  = (~\m5_data_i[8]  | ~\new_[18004]_ ) & (~\m6_data_i[8]  | ~\new_[18836]_ );
  assign \new_[9361]_  = (~\m5_data_i[5]  | ~\new_[18004]_ ) & (~\m6_data_i[5]  | ~\new_[18836]_ );
  assign \new_[9362]_  = (~\m5_data_i[2]  | ~\new_[18004]_ ) & (~\m6_data_i[2]  | ~\new_[17241]_ );
  assign \new_[9363]_  = (~\m5_data_i[0]  | ~\new_[18004]_ ) & (~\m6_data_i[0]  | ~\new_[17241]_ );
  assign \new_[9364]_  = (~\m5_addr_i[22]  | ~\new_[18004]_ ) & (~\m6_addr_i[22]  | ~\new_[18836]_ );
  assign \new_[9365]_  = ~\new_[28327]_  & (~\new_[13363]_  | ~\new_[21497]_ );
  assign \new_[9366]_  = ~\new_[28354]_  & (~\new_[13369]_  | ~\new_[21490]_ );
  assign \new_[9367]_  = ~\new_[28603]_  & (~\new_[13371]_  | ~\new_[21476]_ );
  assign \new_[9368]_  = ~\new_[29847]_  & (~\new_[13374]_  | ~\new_[20528]_ );
  assign \new_[9369]_  = ~\new_[30056]_  & (~\new_[13384]_  | ~\new_[21459]_ );
  assign \new_[9370]_  = ~\new_[28325]_  & (~\new_[13379]_  | ~\new_[21551]_ );
  assign \new_[9371]_  = (~\m5_addr_i[19]  | ~\new_[18004]_ ) & (~\m6_addr_i[19]  | ~\new_[17241]_ );
  assign \new_[9372]_  = ~\new_[28316]_  & (~\new_[13394]_  | ~\new_[21519]_ );
  assign \new_[9373]_  = ~\new_[28060]_  & (~\new_[13417]_  | ~\new_[21496]_ );
  assign \new_[9374]_  = ~\new_[28620]_  & (~\new_[13359]_  | ~\new_[21515]_ );
  assign \new_[9375]_  = (~\m5_addr_i[15]  | ~\new_[18004]_ ) & (~\m6_addr_i[15]  | ~\new_[17241]_ );
  assign \new_[9376]_  = (~\m5_addr_i[14]  | ~\new_[18004]_ ) & (~\m6_addr_i[14]  | ~\new_[17241]_ );
  assign \new_[9377]_  = (~\m5_addr_i[13]  | ~\new_[18004]_ ) & (~\m6_addr_i[13]  | ~\new_[17241]_ );
  assign \new_[9378]_  = (~\m5_data_i[1]  | ~\new_[18004]_ ) & (~\m6_data_i[1]  | ~\new_[18836]_ );
  assign \new_[9379]_  = (~\m5_addr_i[12]  | ~\new_[18004]_ ) & (~\m6_addr_i[12]  | ~\new_[17241]_ );
  assign \new_[9380]_  = (~\m5_addr_i[11]  | ~\new_[18004]_ ) & (~\m6_addr_i[11]  | ~\new_[17241]_ );
  assign \new_[9381]_  = (~\m5_addr_i[10]  | ~\new_[18004]_ ) & (~\m6_addr_i[10]  | ~\new_[18836]_ );
  assign \new_[9382]_  = (~\m5_addr_i[8]  | ~\new_[18004]_ ) & (~\m6_addr_i[8]  | ~\new_[17241]_ );
  assign \new_[9383]_  = (~\m5_addr_i[6]  | ~\new_[18004]_ ) & (~\m6_addr_i[6]  | ~\new_[17241]_ );
  assign \new_[9384]_  = (~\m5_addr_i[0]  | ~\new_[18004]_ ) & (~\m6_addr_i[0]  | ~\new_[17241]_ );
  assign \new_[9385]_  = (~\m5_sel_i[3]  | ~\new_[18004]_ ) & (~\m6_sel_i[3]  | ~\new_[17241]_ );
  assign \new_[9386]_  = (~\m5_sel_i[2]  | ~\new_[18004]_ ) & (~\m6_sel_i[2]  | ~\new_[17241]_ );
  assign \new_[9387]_  = (~\m5_sel_i[1]  | ~\new_[18004]_ ) & (~\m6_sel_i[1]  | ~\new_[17241]_ );
  assign \new_[9388]_  = (~\m5_addr_i[1]  | ~\new_[18004]_ ) & (~\m6_addr_i[1]  | ~\new_[17241]_ );
  assign \new_[9389]_  = (~\new_[13569]_  | ~\new_[28418]_ ) & (~\new_[13568]_  | ~\new_[28723]_ );
  assign \new_[9390]_  = (~\new_[13570]_  | ~\new_[28693]_ ) & (~\new_[14913]_  | ~\new_[28645]_ );
  assign \new_[9391]_  = (~\new_[13597]_  | ~\new_[29193]_ ) & (~\new_[14924]_  | ~\new_[29031]_ );
  assign \new_[9392]_  = (~\new_[13604]_  | ~\new_[29630]_ ) & (~\new_[14929]_  | ~\new_[28112]_ );
  assign \new_[9393]_  = (~\new_[14930]_  | ~\new_[28200]_ ) & (~\new_[13611]_  | ~\new_[28689]_ );
  assign \new_[9394]_  = (~\new_[13616]_  | ~\new_[28938]_ ) & (~\new_[14931]_  | ~\new_[28343]_ );
  assign \new_[9395]_  = ~\new_[11274]_  & (~\new_[13567]_  | ~\new_[28734]_ );
  assign \new_[9396]_  = (~\m5_addr_i[21]  | ~\new_[18004]_ ) & (~\m6_addr_i[21]  | ~\new_[18836]_ );
  assign \new_[9397]_  = (~\new_[14935]_  | ~\new_[27853]_ ) & (~\new_[13619]_  | ~\new_[28051]_ );
  assign \new_[9398]_  = (~\new_[14936]_  | ~\new_[27945]_ ) & (~\new_[13620]_  | ~\new_[28314]_ );
  assign \new_[9399]_  = (~\m7_data_i[28]  | ~\new_[16297]_ ) & (~\m0_data_i[28]  | ~\new_[19575]_ );
  assign \new_[9400]_  = (~\m2_data_i[28]  | ~\new_[16290]_ ) & (~\m1_data_i[28]  | ~\new_[18174]_ );
  assign \new_[9401]_  = (~\m7_data_i[27]  | ~\new_[16297]_ ) & (~\m0_data_i[27]  | ~\new_[19575]_ );
  assign \new_[9402]_  = (~\m7_data_i[26]  | ~\new_[16297]_ ) & (~\m0_data_i[26]  | ~\new_[18083]_ );
  assign \new_[9403]_  = (~\m2_data_i[25]  | ~\new_[16290]_ ) & (~\m1_data_i[25]  | ~\new_[18174]_ );
  assign \new_[9404]_  = (~\new_[13622]_  | ~\new_[27908]_ ) & (~\new_[13621]_  | ~\new_[28323]_ );
  assign \new_[9405]_  = (~\m7_data_i[24]  | ~\new_[16297]_ ) & (~\m0_data_i[24]  | ~\new_[19575]_ );
  assign \new_[9406]_  = (~\m2_data_i[24]  | ~\new_[16290]_ ) & (~\m1_data_i[24]  | ~\new_[18171]_ );
  assign \new_[9407]_  = (~\m7_data_i[23]  | ~\new_[16297]_ ) & (~\m0_data_i[23]  | ~\new_[19575]_ );
  assign \new_[9408]_  = (~\m2_data_i[23]  | ~\new_[16290]_ ) & (~\m1_data_i[23]  | ~\new_[18174]_ );
  assign \new_[9409]_  = (~\m7_data_i[22]  | ~\new_[16297]_ ) & (~\m0_data_i[22]  | ~\new_[18811]_ );
  assign \new_[9410]_  = (~\m2_data_i[22]  | ~\new_[16290]_ ) & (~\m1_data_i[22]  | ~\new_[18174]_ );
  assign \new_[9411]_  = (~\m2_data_i[21]  | ~\new_[16290]_ ) & (~\m1_data_i[21]  | ~\new_[18174]_ );
  assign \new_[9412]_  = (~\m7_data_i[20]  | ~\new_[16297]_ ) & (~\m0_data_i[20]  | ~\new_[19575]_ );
  assign \new_[9413]_  = ~\new_[14756]_  | ~\new_[16141]_  | ~\new_[13360]_  | ~\new_[14755]_ ;
  assign \new_[9414]_  = (~\m7_data_i[18]  | ~\new_[16297]_ ) & (~\m0_data_i[18]  | ~\new_[18083]_ );
  assign \new_[9415]_  = ~\new_[16827]_  | ~\new_[14764]_  | ~\new_[16035]_  | ~\new_[17032]_ ;
  assign \new_[9416]_  = ~\new_[14629]_  | ~\new_[14772]_  | ~\new_[14628]_  | ~\new_[13377]_ ;
  assign \new_[9417]_  = (~\m2_data_i[16]  | ~\new_[16290]_ ) & (~\m1_data_i[16]  | ~\new_[19627]_ );
  assign \new_[9418]_  = ~\new_[17718]_  | ~\new_[14643]_  | ~\new_[17717]_  | ~\new_[18555]_ ;
  assign \new_[9419]_  = (~\m2_data_i[15]  | ~\new_[16290]_ ) & (~\m1_data_i[15]  | ~\new_[19627]_ );
  assign \new_[9420]_  = (~\new_[13627]_  | ~\new_[28750]_ ) & (~\new_[13626]_  | ~\new_[29713]_ );
  assign \new_[9421]_  = ~\new_[17722]_  | ~\new_[14650]_  | ~\new_[17721]_  | ~\new_[14649]_ ;
  assign \new_[9422]_  = (~\m2_data_i[14]  | ~\new_[16290]_ ) & (~\m1_data_i[14]  | ~\new_[18168]_ );
  assign \new_[9423]_  = (~\m7_data_i[13]  | ~\new_[16297]_ ) & (~\m0_data_i[13]  | ~\new_[18083]_ );
  assign \new_[9424]_  = (~\m2_data_i[13]  | ~\new_[16290]_ ) & (~\m1_data_i[13]  | ~\new_[19627]_ );
  assign \new_[9425]_  = ~\new_[14777]_  | ~\new_[16161]_  | ~\new_[16073]_  | ~\new_[17044]_ ;
  assign \new_[9426]_  = (~\m7_data_i[12]  | ~\new_[16297]_ ) & (~\m0_data_i[12]  | ~\new_[18083]_ );
  assign \new_[9427]_  = (~\m2_data_i[12]  | ~\new_[16290]_ ) & (~\m1_data_i[12]  | ~\new_[19627]_ );
  assign \new_[9428]_  = (~\m7_data_i[11]  | ~\new_[16297]_ ) & (~\m0_data_i[11]  | ~\new_[18083]_ );
  assign \new_[9429]_  = (~\m2_data_i[11]  | ~\new_[16290]_ ) & (~\m1_data_i[11]  | ~\new_[18174]_ );
  assign \new_[9430]_  = (~\m2_data_i[10]  | ~\new_[16290]_ ) & (~\m1_data_i[10]  | ~\new_[18170]_ );
  assign \new_[9431]_  = (~\m7_data_i[9]  | ~\new_[16297]_ ) & (~\m0_data_i[9]  | ~\new_[18083]_ );
  assign \new_[9432]_  = (~\m7_data_i[8]  | ~\new_[16297]_ ) & (~\m0_data_i[8]  | ~\new_[18083]_ );
  assign \new_[9433]_  = (~\m2_data_i[8]  | ~\new_[16290]_ ) & (~\m1_data_i[8]  | ~\new_[18169]_ );
  assign \new_[9434]_  = ~\new_[11408]_  & (~\new_[14932]_  | ~\new_[26484]_ );
  assign \new_[9435]_  = (~\m2_data_i[7]  | ~\new_[16290]_ ) & (~\m1_data_i[7]  | ~\new_[18170]_ );
  assign \new_[9436]_  = (~\m7_data_i[6]  | ~\new_[16297]_ ) & (~\m0_data_i[6]  | ~\new_[18083]_ );
  assign \new_[9437]_  = (~\m7_data_i[5]  | ~\new_[16297]_ ) & (~\m0_data_i[5]  | ~\new_[18083]_ );
  assign \new_[9438]_  = (~\m2_data_i[5]  | ~\new_[16290]_ ) & (~\m1_data_i[5]  | ~\new_[18168]_ );
  assign \new_[9439]_  = ~\new_[16171]_  | ~\new_[14790]_  | ~\new_[14788]_  | ~\new_[16170]_ ;
  assign \new_[9440]_  = (~\m2_data_i[4]  | ~\new_[16290]_ ) & (~\m1_data_i[4]  | ~\new_[18169]_ );
  assign \new_[9441]_  = (~\m7_data_i[3]  | ~\new_[16297]_ ) & (~\m0_data_i[3]  | ~\new_[18083]_ );
  assign \new_[9442]_  = ~\new_[14796]_  | ~\new_[17877]_  | ~\new_[16176]_  | ~\new_[17874]_ ;
  assign \new_[9443]_  = (~\m2_data_i[3]  | ~\new_[16290]_ ) & (~\m1_data_i[3]  | ~\new_[19627]_ );
  assign \new_[9444]_  = (~\m7_data_i[2]  | ~\new_[16297]_ ) & (~\m0_data_i[2]  | ~\new_[18083]_ );
  assign \new_[9445]_  = (~\m2_data_i[2]  | ~\new_[16290]_ ) & (~\m1_data_i[2]  | ~\new_[19627]_ );
  assign \new_[9446]_  = (~\m7_data_i[1]  | ~\new_[16297]_ ) & (~\m0_data_i[1]  | ~\new_[18083]_ );
  assign \new_[9447]_  = (~\m2_data_i[1]  | ~\new_[16290]_ ) & (~\m1_data_i[1]  | ~\new_[18168]_ );
  assign \new_[9448]_  = (~\new_[13630]_  | ~\new_[26631]_ ) & (~\new_[13629]_  | ~\new_[28008]_ );
  assign \new_[9449]_  = ~\new_[16217]_  | ~\new_[14810]_  | ~\new_[16222]_  | ~\new_[16185]_ ;
  assign \new_[9450]_  = ~\new_[16200]_  | ~\new_[14797]_  | ~\new_[13413]_  | ~\new_[17060]_ ;
  assign \new_[9451]_  = (~\m2_data_i[0]  | ~\new_[16290]_ ) & (~\m1_data_i[0]  | ~\new_[18168]_ );
  assign \new_[9452]_  = (~\new_[13632]_  | ~\new_[27930]_ ) & (~\new_[13631]_  | ~\new_[27957]_ );
  assign \new_[9453]_  = ~\new_[16151]_  | ~\new_[14800]_  | ~\new_[13400]_  | ~\new_[17094]_ ;
  assign \new_[9454]_  = ~\new_[14775]_  | ~\new_[18668]_  | ~\new_[16201]_  | ~\new_[18664]_ ;
  assign \new_[9455]_  = ~\new_[16110]_  | ~\new_[14804]_  | ~\new_[11374]_  | ~\new_[13408]_ ;
  assign \new_[9456]_  = ~\new_[11332]_  & (~\new_[13589]_  | ~\new_[28709]_ );
  assign \new_[9457]_  = ~\new_[11454]_  & (~\new_[13590]_  | ~\new_[26586]_ );
  assign \new_[9458]_  = (~\new_[13634]_  | ~\new_[28273]_ ) & (~\new_[13633]_  | ~\new_[29140]_ );
  assign \new_[9459]_  = ~\new_[14711]_  | ~\new_[17811]_  | ~\new_[13313]_  | ~\new_[16114]_ ;
  assign \new_[9460]_  = ~\new_[14718]_  | ~\new_[16956]_  | ~\new_[16120]_  | ~\new_[13320]_ ;
  assign \new_[9461]_  = (~\new_[13636]_  | ~\new_[26954]_ ) & (~\new_[13635]_  | ~\new_[28295]_ );
  assign \new_[9462]_  = ~\new_[16123]_  | ~\new_[14815]_  | ~\new_[17108]_  | ~\new_[17110]_ ;
  assign \new_[9463]_  = (~\m2_addr_i[23]  | ~\new_[16290]_ ) & (~\m1_addr_i[23]  | ~\new_[18171]_ );
  assign \new_[9464]_  = (~\m2_addr_i[22]  | ~\new_[16290]_ ) & (~\m1_addr_i[22]  | ~\new_[18171]_ );
  assign \new_[9465]_  = (~\m7_addr_i[21]  | ~\new_[16297]_ ) & (~\m0_addr_i[21]  | ~\new_[19575]_ );
  assign \new_[9466]_  = (~\m2_addr_i[21]  | ~\new_[16290]_ ) & (~\m1_addr_i[21]  | ~\new_[18174]_ );
  assign \new_[9467]_  = (~\m7_addr_i[20]  | ~\new_[16297]_ ) & (~\m0_addr_i[20]  | ~\new_[18811]_ );
  assign \new_[9468]_  = (~\m2_addr_i[20]  | ~\new_[16290]_ ) & (~\m1_addr_i[20]  | ~\new_[18174]_ );
  assign \new_[9469]_  = (~\m7_addr_i[19]  | ~\new_[16297]_ ) & (~\m0_addr_i[19]  | ~\new_[18811]_ );
  assign \new_[9470]_  = (~\m2_addr_i[19]  | ~\new_[16290]_ ) & (~\m1_addr_i[19]  | ~\new_[18174]_ );
  assign \new_[9471]_  = (~\new_[14949]_  | ~\new_[28915]_ ) & (~\new_[13637]_  | ~\new_[29031]_ );
  assign \new_[9472]_  = (~\m7_addr_i[17]  | ~\new_[16297]_ ) & (~\m0_addr_i[17]  | ~\new_[19575]_ );
  assign \new_[9473]_  = (~\m2_addr_i[16]  | ~\new_[16290]_ ) & (~\m1_addr_i[16]  | ~\new_[18170]_ );
  assign \new_[9474]_  = (~\m2_addr_i[15]  | ~\new_[16290]_ ) & (~\m1_addr_i[15]  | ~\new_[18170]_ );
  assign \new_[9475]_  = (~\new_[13639]_  | ~\new_[26771]_ ) & (~\new_[13638]_  | ~\new_[28757]_ );
  assign \new_[9476]_  = (~\m2_addr_i[14]  | ~\new_[16290]_ ) & (~\m1_addr_i[14]  | ~\new_[18174]_ );
  assign \new_[9477]_  = (~\m2_addr_i[13]  | ~\new_[16290]_ ) & (~\m1_addr_i[13]  | ~\new_[19627]_ );
  assign \new_[9478]_  = (~\m2_addr_i[12]  | ~\new_[16290]_ ) & (~\m1_addr_i[12]  | ~\new_[18171]_ );
  assign \new_[9479]_  = (~\m7_addr_i[11]  | ~\new_[16297]_ ) & (~\m0_addr_i[11]  | ~\new_[18083]_ );
  assign \new_[9480]_  = (~\m2_addr_i[11]  | ~\new_[16290]_ ) & (~\m1_addr_i[11]  | ~\new_[18174]_ );
  assign \new_[9481]_  = (~\new_[13642]_  | ~\new_[28719]_ ) & (~\new_[13641]_  | ~\new_[29010]_ );
  assign \new_[9482]_  = (~\m2_addr_i[10]  | ~\new_[16290]_ ) & (~\m1_addr_i[10]  | ~\new_[18174]_ );
  assign \new_[9483]_  = (~\m7_addr_i[9]  | ~\new_[16297]_ ) & (~\m0_addr_i[9]  | ~\new_[18083]_ );
  assign \new_[9484]_  = (~\m7_addr_i[8]  | ~\new_[16297]_ ) & (~\m0_addr_i[8]  | ~\new_[18083]_ );
  assign \new_[9485]_  = (~\m7_addr_i[7]  | ~\new_[16297]_ ) & (~\m0_addr_i[7]  | ~\new_[18083]_ );
  assign \new_[9486]_  = (~\m7_addr_i[6]  | ~\new_[16297]_ ) & (~\m0_addr_i[6]  | ~\new_[19575]_ );
  assign \new_[9487]_  = (~\m2_addr_i[6]  | ~\new_[16290]_ ) & (~\m1_addr_i[6]  | ~\new_[18174]_ );
  assign \new_[9488]_  = (~\m7_addr_i[5]  | ~\new_[16297]_ ) & (~\new_[31848]_  | ~\new_[18083]_ );
  assign \new_[9489]_  = (~\new_[31095]_  | ~\new_[16290]_ ) & (~\m1_addr_i[5]  | ~\new_[18169]_ );
  assign \new_[9490]_  = (~\m2_addr_i[4]  | ~\new_[16290]_ ) & (~\m1_addr_i[4]  | ~\new_[18170]_ );
  assign \new_[9491]_  = (~\new_[31726]_  | ~\new_[16297]_ ) & (~\m0_addr_i[3]  | ~\new_[18083]_ );
  assign \new_[9492]_  = (~\new_[31399]_  | ~\new_[16290]_ ) & (~\m1_addr_i[3]  | ~\new_[19627]_ );
  assign \new_[9493]_  = (~\m2_addr_i[2]  | ~\new_[16290]_ ) & (~\new_[31477]_  | ~\new_[18170]_ );
  assign \new_[9494]_  = (~\m7_addr_i[1]  | ~\new_[16297]_ ) & (~\m0_addr_i[1]  | ~\new_[19575]_ );
  assign \new_[9495]_  = (~\m2_sel_i[3]  | ~\new_[16290]_ ) & (~\m1_sel_i[3]  | ~\new_[18174]_ );
  assign \new_[9496]_  = (~\m2_sel_i[2]  | ~\new_[16290]_ ) & (~\m1_sel_i[2]  | ~\new_[18174]_ );
  assign \new_[9497]_  = (~\m7_sel_i[1]  | ~\new_[16297]_ ) & (~\m0_sel_i[1]  | ~\new_[18083]_ );
  assign \new_[9498]_  = (~\m2_sel_i[1]  | ~\new_[16290]_ ) & (~\m1_sel_i[1]  | ~\new_[19627]_ );
  assign \new_[9499]_  = (~\m7_sel_i[0]  | ~\new_[16297]_ ) & (~\m0_sel_i[0]  | ~\new_[19575]_ );
  assign \new_[9500]_  = (~m2_we_i | ~\new_[16290]_ ) & (~m1_we_i | ~\new_[18169]_ );
  assign \new_[9501]_  = (~\new_[32347]_  | ~\m0_data_i[15] ) & (~\new_[13487]_  | ~\m1_data_i[15] );
  assign \new_[9502]_  = (~\new_[13526]_  | ~\m4_data_i[15] ) & (~\new_[14849]_  | ~\m5_data_i[15] );
  assign \new_[9503]_  = (~\new_[32347]_  | ~\m0_data_i[14] ) & (~\new_[13487]_  | ~\m1_data_i[14] );
  assign \new_[9504]_  = (~\new_[17239]_  | ~\new_[31885]_ ) & (~\new_[16280]_  | ~\new_[31292]_ );
  assign \new_[9505]_  = (~\new_[13525]_  | ~\m4_data_i[14] ) & (~\new_[14850]_  | ~\m5_data_i[14] );
  assign \new_[9506]_  = (~\new_[32347]_  | ~\m0_data_i[13] ) & (~\new_[13487]_  | ~\m1_data_i[13] );
  assign \new_[9507]_  = (~\new_[13525]_  | ~\m4_data_i[13] ) & (~\new_[14848]_  | ~\m5_data_i[13] );
  assign \new_[9508]_  = (~\new_[32347]_  | ~\m0_data_i[12] ) & (~\new_[13487]_  | ~\m1_data_i[12] );
  assign \new_[9509]_  = (~\new_[13525]_  | ~\m4_data_i[12] ) & (~\new_[14850]_  | ~\m5_data_i[12] );
  assign \new_[9510]_  = (~\new_[32347]_  | ~\m0_data_i[11] ) & (~\new_[13487]_  | ~\m1_data_i[11] );
  assign \new_[9511]_  = (~\new_[13525]_  | ~\m4_data_i[11] ) & (~\new_[14850]_  | ~\m5_data_i[11] );
  assign \new_[9512]_  = (~\new_[32347]_  | ~\m0_data_i[10] ) & (~\new_[13487]_  | ~\m1_data_i[10] );
  assign \new_[9513]_  = (~\new_[13526]_  | ~\m4_data_i[10] ) & (~\new_[14850]_  | ~\m5_data_i[10] );
  assign \new_[9514]_  = (~\new_[32347]_  | ~\m0_data_i[9] ) & (~\new_[13487]_  | ~\m1_data_i[9] );
  assign \new_[9515]_  = (~\new_[13526]_  | ~\m4_data_i[9] ) & (~\new_[14849]_  | ~\m5_data_i[9] );
  assign \new_[9516]_  = (~\new_[32347]_  | ~\m0_data_i[8] ) & (~\new_[13487]_  | ~\m1_data_i[8] );
  assign \new_[9517]_  = (~\new_[13526]_  | ~\m4_data_i[8] ) & (~\new_[14850]_  | ~\m5_data_i[8] );
  assign \new_[9518]_  = (~\new_[32347]_  | ~\m0_data_i[7] ) & (~\new_[13487]_  | ~\m1_data_i[7] );
  assign \new_[9519]_  = (~\new_[13526]_  | ~\m4_data_i[7] ) & (~\new_[14850]_  | ~\m5_data_i[7] );
  assign \new_[9520]_  = (~\new_[32347]_  | ~\m0_data_i[6] ) & (~\new_[13487]_  | ~\m1_data_i[6] );
  assign \new_[9521]_  = (~\new_[13526]_  | ~\m4_data_i[6] ) & (~\new_[14848]_  | ~\m5_data_i[6] );
  assign \new_[9522]_  = (~\new_[32347]_  | ~\m0_data_i[5] ) & (~\new_[13487]_  | ~\m1_data_i[5] );
  assign \new_[9523]_  = ~\new_[11452]_  & ~\new_[11388]_ ;
  assign \new_[9524]_  = (~\new_[13526]_  | ~\m4_data_i[5] ) & (~\new_[14849]_  | ~\m5_data_i[5] );
  assign \new_[9525]_  = (~\new_[32347]_  | ~\m0_data_i[4] ) & (~\new_[13487]_  | ~\m1_data_i[4] );
  assign \new_[9526]_  = (~\new_[13526]_  | ~\m4_data_i[4] ) & (~\new_[14848]_  | ~\m5_data_i[4] );
  assign \new_[9527]_  = (~\new_[32347]_  | ~\m0_data_i[3] ) & (~\new_[13487]_  | ~\m1_data_i[3] );
  assign \new_[9528]_  = (~\new_[13525]_  | ~\m4_data_i[3] ) & (~\new_[14850]_  | ~\m5_data_i[3] );
  assign \new_[9529]_  = (~\new_[32347]_  | ~\m0_data_i[2] ) & (~\new_[13487]_  | ~\m1_data_i[2] );
  assign \new_[9530]_  = (~\new_[13525]_  | ~\m4_data_i[2] ) & (~\new_[14850]_  | ~\m5_data_i[2] );
  assign \new_[9531]_  = (~\new_[32347]_  | ~\m0_data_i[1] ) & (~\new_[13487]_  | ~\m1_data_i[1] );
  assign \new_[9532]_  = (~\new_[13525]_  | ~\m4_data_i[1] ) & (~\new_[14848]_  | ~\m5_data_i[1] );
  assign \new_[9533]_  = (~\new_[32347]_  | ~\m0_data_i[0] ) & (~\new_[13487]_  | ~\m1_data_i[0] );
  assign \new_[9534]_  = (~\new_[13525]_  | ~\m4_data_i[0] ) & (~\new_[14850]_  | ~\m5_data_i[0] );
  assign \new_[9535]_  = ~m0_stb_i | ~\new_[26156]_  | ~\new_[16280]_ ;
  assign \new_[9536]_  = ~\new_[21265]_  | ~\new_[14905]_  | ~\new_[21264]_  | ~\new_[16511]_ ;
  assign \new_[9537]_  = ~\new_[11677]_  | ~\new_[11753]_ ;
  assign \new_[9538]_  = ~\new_[21281]_  | ~\new_[14906]_  | ~\new_[20367]_  | ~\new_[16514]_ ;
  assign \new_[9539]_  = ~\new_[11684]_  | ~\new_[11764]_ ;
  assign \new_[9540]_  = ~\new_[19387]_  | ~\new_[14907]_  | ~\new_[20365]_  | ~\new_[14257]_ ;
  assign \new_[9541]_  = ~\new_[11687]_  | ~\new_[11769]_ ;
  assign \new_[9542]_  = ~\new_[21299]_  | ~\new_[14909]_  | ~\new_[19397]_  | ~\new_[15613]_ ;
  assign \new_[9543]_  = ~\new_[11705]_  | ~\new_[11786]_ ;
  assign \new_[9544]_  = ~\new_[11712]_  | ~\new_[11797]_ ;
  assign \new_[9545]_  = ~\new_[13523]_  | ~\new_[11799]_ ;
  assign \new_[9546]_  = ~\new_[21307]_  | ~\new_[14910]_  | ~\new_[22499]_  | ~\new_[15634]_ ;
  assign \new_[9547]_  = ~\new_[11722]_  | ~\new_[11807]_ ;
  assign \new_[9548]_  = ~\new_[21328]_  | ~\new_[14911]_  | ~\new_[20392]_  | ~\new_[16530]_ ;
  assign \new_[9549]_  = (~\new_[32346]_  | ~m0_we_i) & (~\new_[13487]_  | ~m1_we_i);
  assign \new_[9550]_  = (~\new_[13526]_  | ~m4_we_i) & (~\new_[14850]_  | ~m5_we_i);
  assign \new_[9551]_  = ~\new_[20342]_  | (~\new_[13746]_  & ~\new_[27873]_ );
  assign \new_[9552]_  = ~\new_[20338]_  | (~\new_[13748]_  & ~\new_[26533]_ );
  assign \new_[9553]_  = ~\new_[30259]_  & (~\new_[13566]_  | ~\new_[28256]_ );
  assign \new_[9554]_  = ~\new_[29027]_  & (~\new_[13572]_  | ~\new_[28517]_ );
  assign \new_[9555]_  = ~\new_[28994]_  & (~\new_[13576]_  | ~\new_[28505]_ );
  assign \new_[9556]_  = ~\new_[29137]_  & (~\new_[13579]_  | ~\new_[28198]_ );
  assign \new_[9557]_  = ~\new_[30447]_  & (~\new_[13581]_  | ~\new_[23057]_ );
  assign \new_[9558]_  = ~\new_[28996]_  & (~\new_[13585]_  | ~\new_[21495]_ );
  assign \new_[9559]_  = ~\new_[28858]_  & (~\new_[13588]_  | ~\new_[21467]_ );
  assign \new_[9560]_  = ~\new_[30742]_  & (~\new_[13593]_  | ~\new_[22985]_ );
  assign \new_[9561]_  = ~\new_[29049]_  & (~\new_[13596]_  | ~\new_[23061]_ );
  assign \new_[9562]_  = ~\new_[29325]_  & (~\new_[13598]_  | ~\new_[28809]_ );
  assign \new_[9563]_  = ~\new_[29282]_  & (~\new_[13599]_  | ~\new_[22849]_ );
  assign \new_[9564]_  = ~\new_[29486]_  & (~\new_[13605]_  | ~\new_[28521]_ );
  assign \new_[9565]_  = ~\new_[29030]_  & (~\new_[13609]_  | ~\new_[20866]_ );
  assign \new_[9566]_  = ~\new_[30100]_  & (~\new_[13612]_  | ~\new_[20526]_ );
  assign \new_[9567]_  = ~\new_[21124]_  | (~\new_[13734]_  & ~\new_[26892]_ );
  assign \new_[9568]_  = ~\new_[21139]_  | (~\new_[13736]_  & ~\new_[26966]_ );
  assign \new_[9569]_  = ~\new_[20303]_  | (~\new_[13739]_  & ~\new_[28168]_ );
  assign \new_[9570]_  = ~\new_[21162]_  | (~\new_[13741]_  & ~\new_[28172]_ );
  assign \new_[9571]_  = ~\new_[21168]_  | (~\new_[13742]_  & ~\new_[27867]_ );
  assign \new_[9572]_  = (~\m7_data_i[12]  | ~\new_[16296]_ ) & (~\m0_data_i[12]  | ~\new_[20545]_ );
  assign \new_[9573]_  = (~\m5_data_i[10]  | ~\new_[18004]_ ) & (~\m6_data_i[10]  | ~\new_[17241]_ );
  assign \new_[9574]_  = (~\m2_data_i[21]  | ~\new_[17193]_ ) & (~\m1_data_i[21]  | ~\new_[19633]_ );
  assign \new_[9575]_  = ~\new_[14589]_  & (~\new_[14878]_  | ~\m4_addr_i[25] );
  assign \new_[9576]_  = (~\m2_data_i[20]  | ~\new_[17193]_ ) & (~\m1_data_i[20]  | ~\new_[19633]_ );
  assign \new_[9577]_  = (~\m5_addr_i[11]  | ~\new_[17203]_ ) & (~\m4_addr_i[11]  | ~\new_[17271]_ );
  assign \new_[9578]_  = (~\m2_data_i[19]  | ~\new_[17193]_ ) & (~\m1_data_i[19]  | ~\new_[19633]_ );
  assign \new_[9579]_  = (~\m2_data_i[18]  | ~\new_[17193]_ ) & (~\m1_data_i[18]  | ~\new_[18917]_ );
  assign \new_[9580]_  = (~\m2_data_i[17]  | ~\new_[17193]_ ) & (~\m1_data_i[17]  | ~\new_[18917]_ );
  assign \new_[9581]_  = (~\m4_data_i[17]  | ~\new_[17260]_ ) & (~\m3_data_i[17]  | ~\new_[18175]_ );
  assign \new_[9582]_  = (~\m2_data_i[16]  | ~\new_[17193]_ ) & (~\m1_data_i[16]  | ~\new_[19633]_ );
  assign \new_[9583]_  = (~\m2_data_i[15]  | ~\new_[17193]_ ) & (~\m1_data_i[15]  | ~\new_[18916]_ );
  assign \new_[9584]_  = (~\m4_data_i[15]  | ~\new_[17260]_ ) & (~\m3_data_i[15]  | ~\new_[18175]_ );
  assign \new_[9585]_  = (~\m2_data_i[14]  | ~\new_[17193]_ ) & (~\m1_data_i[14]  | ~\new_[18917]_ );
  assign \new_[9586]_  = (~\m5_data_i[10]  | ~\new_[20544]_ ) & (~\m6_data_i[10]  | ~\new_[17213]_ );
  assign \new_[9587]_  = (~\m4_data_i[14]  | ~\new_[17260]_ ) & (~\m3_data_i[14]  | ~\new_[18175]_ );
  assign \new_[9588]_  = (~\m2_data_i[13]  | ~\new_[17193]_ ) & (~\m1_data_i[13]  | ~\new_[18917]_ );
  assign \new_[9589]_  = (~\m4_data_i[13]  | ~\new_[17260]_ ) & (~\m3_data_i[13]  | ~\new_[18175]_ );
  assign \new_[9590]_  = (~\m2_data_i[12]  | ~\new_[17193]_ ) & (~\m1_data_i[12]  | ~\new_[18917]_ );
  assign \new_[9591]_  = (~\m4_data_i[12]  | ~\new_[17260]_ ) & (~\m3_data_i[12]  | ~\new_[18175]_ );
  assign \new_[9592]_  = (~\m2_data_i[11]  | ~\new_[17193]_ ) & (~\m1_data_i[11]  | ~\new_[18917]_ );
  assign \new_[9593]_  = (~\m2_data_i[10]  | ~\new_[17193]_ ) & (~\m1_data_i[10]  | ~\new_[18917]_ );
  assign \new_[9594]_  = (~\m4_data_i[10]  | ~\new_[17260]_ ) & (~\m3_data_i[10]  | ~\new_[18175]_ );
  assign \new_[9595]_  = (~\m2_data_i[9]  | ~\new_[17193]_ ) & (~\m1_data_i[9]  | ~\new_[18917]_ );
  assign \new_[9596]_  = (~\m4_data_i[9]  | ~\new_[17260]_ ) & (~\m3_data_i[9]  | ~\new_[18175]_ );
  assign \new_[9597]_  = (~\m2_data_i[8]  | ~\new_[17193]_ ) & (~\m1_data_i[8]  | ~\new_[18193]_ );
  assign \new_[9598]_  = (~\m4_data_i[8]  | ~\new_[17260]_ ) & (~\m3_data_i[8]  | ~\new_[18175]_ );
  assign \new_[9599]_  = (~\m2_data_i[7]  | ~\new_[17193]_ ) & (~\m1_data_i[7]  | ~\new_[18917]_ );
  assign \new_[9600]_  = (~\m4_data_i[7]  | ~\new_[17260]_ ) & (~\m3_data_i[7]  | ~\new_[18175]_ );
  assign \new_[9601]_  = (~\m2_data_i[6]  | ~\new_[17193]_ ) & (~\m1_data_i[6]  | ~\new_[18193]_ );
  assign \new_[9602]_  = ~\new_[13213]_  & (~\new_[32348]_  | ~\m0_addr_i[27] );
  assign \new_[9603]_  = (~\m4_data_i[6]  | ~\new_[17260]_ ) & (~\m3_data_i[6]  | ~\new_[18175]_ );
  assign \new_[9604]_  = (~\m5_addr_i[8]  | ~\new_[17203]_ ) & (~\m4_addr_i[8]  | ~\new_[17271]_ );
  assign \new_[9605]_  = (~\m2_data_i[5]  | ~\new_[17193]_ ) & (~\m1_data_i[5]  | ~\new_[18917]_ );
  assign \new_[9606]_  = (~\m4_data_i[5]  | ~\new_[17260]_ ) & (~\m3_data_i[5]  | ~\new_[18175]_ );
  assign \new_[9607]_  = (~\m2_data_i[4]  | ~\new_[17193]_ ) & (~\m1_data_i[4]  | ~\new_[18917]_ );
  assign \new_[9608]_  = (~\m4_data_i[4]  | ~\new_[17260]_ ) & (~\m3_data_i[4]  | ~\new_[18175]_ );
  assign \new_[9609]_  = ~\new_[13214]_  & (~\new_[14830]_  | ~\m7_addr_i[27] );
  assign \new_[9610]_  = (~\m2_data_i[3]  | ~\new_[17193]_ ) & (~\m1_data_i[3]  | ~\new_[18193]_ );
  assign \new_[9611]_  = (~\m4_data_i[3]  | ~\new_[17260]_ ) & (~\m3_data_i[3]  | ~\new_[18175]_ );
  assign \new_[9612]_  = (~\m2_data_i[2]  | ~\new_[17193]_ ) & (~\m1_data_i[2]  | ~\new_[18917]_ );
  assign \new_[9613]_  = (~\m4_data_i[2]  | ~\new_[17260]_ ) & (~\m3_data_i[2]  | ~\new_[18175]_ );
  assign \new_[9614]_  = (~\m2_data_i[1]  | ~\new_[17193]_ ) & (~\m1_data_i[1]  | ~\new_[18917]_ );
  assign \new_[9615]_  = (~\m4_data_i[1]  | ~\new_[17260]_ ) & (~\m3_data_i[1]  | ~\new_[18175]_ );
  assign \new_[9616]_  = (~\m2_data_i[0]  | ~\new_[17193]_ ) & (~\m1_data_i[0]  | ~\new_[18916]_ );
  assign \new_[9617]_  = (~\m4_data_i[0]  | ~\new_[17260]_ ) & (~\m3_data_i[0]  | ~\new_[18175]_ );
  assign \new_[9618]_  = (~\m5_addr_i[2]  | ~\new_[18015]_ ) & (~\m6_addr_i[2]  | ~\new_[17229]_ );
  assign \new_[9619]_  = (~\m5_addr_i[16]  | ~\new_[18016]_ ) & (~\m6_addr_i[16]  | ~\new_[17229]_ );
  assign \new_[9620]_  = (~\new_[17260]_  | ~\m4_addr_i[28] ) & (~\new_[18175]_  | ~\m3_addr_i[28] );
  assign \new_[9621]_  = (~\new_[17260]_  | ~\m4_addr_i[27] ) & (~\new_[18175]_  | ~\m3_addr_i[27] );
  assign \new_[9622]_  = (~\m5_data_i[16]  | ~\new_[18004]_ ) & (~\m6_data_i[16]  | ~\new_[17241]_ );
  assign \new_[9623]_  = (~\m2_addr_i[7]  | ~\new_[17193]_ ) & (~\m1_addr_i[7]  | ~\new_[18916]_ );
  assign \new_[9624]_  = (~\new_[17260]_  | ~\m4_addr_i[24] ) & (~\new_[18175]_  | ~\m3_addr_i[24] );
  assign \new_[9625]_  = ~\new_[13216]_  & (~\new_[14839]_  | ~\m3_addr_i[26] );
  assign \new_[9626]_  = (~\m5_data_i[22]  | ~\new_[18752]_ ) & (~\m6_data_i[22]  | ~\new_[17213]_ );
  assign \new_[9627]_  = (~\m2_addr_i[22]  | ~\new_[17193]_ ) & (~\m1_addr_i[22]  | ~\new_[19633]_ );
  assign \new_[9628]_  = ~\new_[13681]_  & ~\new_[13982]_ ;
  assign \new_[9629]_  = (~\m5_addr_i[10]  | ~\new_[17203]_ ) & (~\m4_addr_i[10]  | ~\new_[17271]_ );
  assign \new_[9630]_  = (~\m2_addr_i[21]  | ~\new_[17193]_ ) & (~\m1_addr_i[21]  | ~\new_[19633]_ );
  assign \new_[9631]_  = ~\new_[13217]_  & (~\new_[14830]_  | ~\m7_addr_i[25] );
  assign \new_[9632]_  = (~m4_we_i | ~\new_[17260]_ ) & (~m3_we_i | ~\new_[18175]_ );
  assign \new_[9633]_  = (~\m2_addr_i[20]  | ~\new_[17193]_ ) & (~\m1_addr_i[20]  | ~\new_[19633]_ );
  assign \new_[9634]_  = (~\m2_addr_i[19]  | ~\new_[17193]_ ) & (~\m1_addr_i[19]  | ~\new_[19633]_ );
  assign \new_[9635]_  = (~\m2_addr_i[18]  | ~\new_[17193]_ ) & (~\m1_addr_i[18]  | ~\new_[18917]_ );
  assign \new_[9636]_  = ~\new_[13738]_  & ~\new_[13987]_ ;
  assign \new_[9637]_  = (~\m2_addr_i[17]  | ~\new_[17193]_ ) & (~\m1_addr_i[17]  | ~\new_[18916]_ );
  assign \new_[9638]_  = (~\m5_data_i[19]  | ~\new_[18755]_ ) & (~\m6_data_i[19]  | ~\new_[17213]_ );
  assign \new_[9639]_  = (~\m2_addr_i[16]  | ~\new_[17193]_ ) & (~\m1_addr_i[16]  | ~\new_[18916]_ );
  assign \new_[9640]_  = (~\m2_addr_i[15]  | ~\new_[17193]_ ) & (~\m1_addr_i[15]  | ~\new_[18917]_ );
  assign \new_[9641]_  = (~\m4_addr_i[15]  | ~\new_[17260]_ ) & (~\m3_addr_i[15]  | ~\new_[18175]_ );
  assign \new_[9642]_  = (~\m2_addr_i[14]  | ~\new_[17193]_ ) & (~\m1_addr_i[14]  | ~\new_[19633]_ );
  assign \new_[9643]_  = (~\m4_addr_i[14]  | ~\new_[17260]_ ) & (~\m3_addr_i[14]  | ~\new_[18175]_ );
  assign \new_[9644]_  = ~\new_[15289]_  & ~\new_[13625]_ ;
  assign \new_[9645]_  = (~\m2_addr_i[13]  | ~\new_[17193]_ ) & (~\m1_addr_i[13]  | ~\new_[19633]_ );
  assign \new_[9646]_  = (~\m2_addr_i[12]  | ~\new_[17193]_ ) & (~\m1_addr_i[12]  | ~\new_[18917]_ );
  assign \new_[9647]_  = (~\m5_data_i[29]  | ~\new_[18738]_ ) & (~\m6_data_i[29]  | ~\new_[18030]_ );
  assign \new_[9648]_  = (~\m2_addr_i[11]  | ~\new_[17193]_ ) & (~\m1_addr_i[11]  | ~\new_[19633]_ );
  assign \new_[9649]_  = ~\new_[14964]_  & ~\new_[13744]_ ;
  assign \new_[9650]_  = (~\m5_data_i[0]  | ~\new_[18016]_ ) & (~\m6_data_i[0]  | ~\new_[17229]_ );
  assign \new_[9651]_  = (~\m2_addr_i[10]  | ~\new_[17193]_ ) & (~\m1_addr_i[10]  | ~\new_[19633]_ );
  assign \new_[9652]_  = (~\m2_addr_i[9]  | ~\new_[17193]_ ) & (~\m1_addr_i[9]  | ~\new_[19633]_ );
  assign \new_[9653]_  = (~\m2_addr_i[8]  | ~\new_[17193]_ ) & (~\m1_addr_i[8]  | ~\new_[18916]_ );
  assign \new_[9654]_  = (~\m4_addr_i[8]  | ~\new_[17260]_ ) & (~\m3_addr_i[8]  | ~\new_[18175]_ );
  assign \new_[9655]_  = ~\new_[14965]_  & ~\new_[14000]_ ;
  assign \new_[9656]_  = (~\m4_addr_i[5]  | ~\new_[17260]_ ) & (~\m3_addr_i[5]  | ~\new_[18175]_ );
  assign \new_[9657]_  = ~\new_[14967]_  & ~\new_[13749]_ ;
  assign \new_[9658]_  = (~\m4_addr_i[4]  | ~\new_[17260]_ ) & (~\m3_addr_i[4]  | ~\new_[18175]_ );
  assign \new_[9659]_  = ~\new_[14078]_  & ~\new_[13659]_ ;
  assign \new_[9660]_  = (~\m2_addr_i[1]  | ~\new_[17193]_ ) & (~\m1_addr_i[1]  | ~\new_[18917]_ );
  assign \new_[9661]_  = (~\m2_sel_i[3]  | ~\new_[17193]_ ) & (~\m1_sel_i[3]  | ~\new_[19633]_ );
  assign \new_[9662]_  = (~\m2_sel_i[0]  | ~\new_[17193]_ ) & (~\m1_sel_i[0]  | ~\new_[19633]_ );
  assign \new_[9663]_  = ~\new_[14969]_  & ~\new_[14030]_ ;
  assign \new_[9664]_  = ~\new_[13208]_  & (~\new_[32348]_  | ~\m0_addr_i[26] );
  assign \new_[9665]_  = ~\new_[13762]_  & ~\new_[14035]_ ;
  assign \new_[9666]_  = (~\m5_data_i[23]  | ~\new_[18749]_ ) & (~\m6_data_i[23]  | ~\new_[17213]_ );
  assign \new_[9667]_  = ~\new_[13767]_  & ~\new_[14044]_ ;
  assign \new_[9668]_  = (~\m5_addr_i[20]  | ~\new_[18748]_ ) & (~\m6_addr_i[20]  | ~\new_[17213]_ );
  assign \new_[9669]_  = ~\new_[13769]_  & ~\new_[14057]_ ;
  assign \new_[9670]_  = (~\m5_addr_i[17]  | ~\new_[18754]_ ) & (~\m6_addr_i[17]  | ~\new_[17213]_ );
  assign \new_[9671]_  = ~\new_[13710]_  & ~\new_[14064]_ ;
  assign \new_[9672]_  = (~\m5_data_i[8]  | ~\new_[18750]_ ) & (~\m6_data_i[8]  | ~\new_[17213]_ );
  assign \new_[9673]_  = ~\new_[14080]_  & ~\new_[13661]_ ;
  assign \new_[9674]_  = ~\new_[13680]_  & ~\new_[13618]_ ;
  assign \new_[9675]_  = (~\m5_addr_i[11]  | ~\new_[18748]_ ) & (~\m6_addr_i[11]  | ~\new_[17213]_ );
  assign \new_[9676]_  = (~\m5_data_i[1]  | ~\new_[18752]_ ) & (~\m6_data_i[1]  | ~\new_[17213]_ );
  assign \new_[9677]_  = (~\m5_addr_i[9]  | ~\new_[18758]_ ) & (~\m6_addr_i[9]  | ~\new_[17213]_ );
  assign \new_[9678]_  = ~\new_[13207]_  & (~\new_[14839]_  | ~\m3_addr_i[25] );
  assign \new_[9679]_  = (~\m5_addr_i[8]  | ~\new_[18754]_ ) & (~\m6_addr_i[8]  | ~\new_[17213]_ );
  assign \new_[9680]_  = (~\m5_addr_i[6]  | ~\new_[18749]_ ) & (~\m6_addr_i[6]  | ~\new_[17213]_ );
  assign \new_[9681]_  = ~\new_[13662]_  & (~\new_[15934]_  | ~\new_[28756]_ );
  assign \new_[9682]_  = ~\new_[28680]_  & (~\new_[15030]_  | ~\new_[22705]_ );
  assign \new_[9683]_  = (~\m5_addr_i[4]  | ~\new_[20544]_ ) & (~\m6_addr_i[4]  | ~\new_[17213]_ );
  assign \new_[9684]_  = ~\new_[13663]_  & (~\new_[15935]_  | ~\new_[29662]_ );
  assign \new_[9685]_  = ~\new_[14584]_  & (~\new_[14878]_  | ~\m4_addr_i[26] );
  assign \new_[9686]_  = ~\new_[27875]_  & (~\new_[15492]_  | ~\new_[23165]_ );
  assign \new_[9687]_  = (~\m5_addr_i[3]  | ~\new_[18750]_ ) & (~\m6_addr_i[3]  | ~\new_[17213]_ );
  assign \new_[9688]_  = ~\new_[26454]_  & (~\new_[15493]_  | ~\new_[24675]_ );
  assign \new_[9689]_  = (~\m5_addr_i[2]  | ~\new_[18758]_ ) & (~\m6_addr_i[2]  | ~\new_[17213]_ );
  assign \new_[9690]_  = ~\new_[24584]_  & (~\new_[15145]_  | ~\new_[22778]_ );
  assign \new_[9691]_  = (~\m5_addr_i[1]  | ~\new_[18759]_ ) & (~\m6_addr_i[1]  | ~\new_[17213]_ );
  assign \new_[9692]_  = ~\new_[13664]_  & (~\new_[14543]_  | ~\new_[29000]_ );
  assign \new_[9693]_  = (~\m5_addr_i[0]  | ~\new_[18759]_ ) & (~\m6_addr_i[0]  | ~\new_[17213]_ );
  assign \new_[9694]_  = ~\new_[26800]_  & (~\new_[15494]_  | ~\new_[24456]_ );
  assign \new_[9695]_  = (~\m5_sel_i[2]  | ~\new_[18751]_ ) & (~\m6_sel_i[2]  | ~\new_[17213]_ );
  assign \new_[9696]_  = ~\new_[28619]_  & (~\new_[15151]_  | ~\new_[21404]_ );
  assign \new_[9697]_  = ~\new_[13666]_  & (~\new_[14547]_  | ~\new_[29871]_ );
  assign \new_[9698]_  = ~\new_[26628]_  & (~\new_[15496]_  | ~\new_[24281]_ );
  assign \new_[9699]_  = ~\new_[29982]_  & (~\new_[15475]_  | ~\new_[24413]_ );
  assign \new_[9700]_  = ~\new_[13667]_  & (~\new_[14549]_  | ~\new_[28897]_ );
  assign \new_[9701]_  = ~\new_[28868]_  & (~\new_[15498]_  | ~\new_[23268]_ );
  assign \new_[9702]_  = ~\new_[28735]_  & (~\new_[15476]_  | ~\new_[26844]_ );
  assign \new_[9703]_  = ~\new_[13668]_  & (~\new_[16314]_  | ~\new_[23067]_ );
  assign \new_[9704]_  = ~\new_[29638]_  & (~\new_[15034]_  | ~\new_[21346]_ );
  assign \new_[9705]_  = ~\new_[24088]_  & (~\new_[15077]_  | ~\new_[21530]_ );
  assign \new_[9706]_  = ~\new_[27866]_  & (~\new_[15478]_  | ~\new_[26616]_ );
  assign \new_[9707]_  = ~\new_[26499]_  & (~\new_[15502]_  | ~\new_[28772]_ );
  assign \new_[9708]_  = ~\new_[24494]_  & (~\new_[15177]_  | ~\new_[21427]_ );
  assign \new_[9709]_  = ~\new_[13653]_  & (~\new_[15762]_  | ~\new_[24653]_ );
  assign \new_[9710]_  = ~\new_[13669]_  & (~\new_[16528]_  | ~\new_[23091]_ );
  assign \new_[9711]_  = ~\new_[28759]_  & (~\new_[15036]_  | ~\new_[21414]_ );
  assign \new_[9712]_  = ~\new_[27813]_  & (~\new_[15184]_  | ~\new_[20409]_ );
  assign \new_[9713]_  = ~\new_[29805]_  & (~\new_[15481]_  | ~\new_[28196]_ );
  assign \new_[9714]_  = ~\new_[13670]_  & (~\new_[16392]_  | ~\new_[27780]_ );
  assign \new_[9715]_  = ~\new_[29304]_  & (~\new_[15507]_  | ~\new_[23137]_ );
  assign \new_[9716]_  = ~\new_[28365]_  & (~\new_[15197]_  | ~\new_[21407]_ );
  assign \new_[9717]_  = ~\new_[14585]_  & (~\new_[14880]_  | ~\m4_addr_i[24] );
  assign \new_[9718]_  = ~\new_[29364]_  & (~\new_[15039]_  | ~\new_[22774]_ );
  assign \new_[9719]_  = ~\new_[13671]_  & (~\new_[14920]_  | ~\new_[29937]_ );
  assign \new_[9720]_  = ~\new_[27832]_  & (~\new_[15509]_  | ~\new_[23968]_ );
  assign \new_[9721]_  = ~\new_[28005]_  & (~\new_[15511]_  | ~\new_[28604]_ );
  assign \new_[9722]_  = ~\new_[13672]_  & (~\new_[16331]_  | ~\new_[28669]_ );
  assign \new_[9723]_  = ~\new_[29092]_  & (~\new_[15206]_  | ~\new_[20432]_ );
  assign \new_[9724]_  = ~\new_[13673]_  & (~\new_[16317]_  | ~\new_[29334]_ );
  assign \new_[9725]_  = (~\new_[16296]_  | ~\new_[31885]_ ) & (~\new_[18764]_  | ~\new_[31292]_ );
  assign \new_[9726]_  = ~\new_[26705]_  & (~\new_[15513]_  | ~\new_[23166]_ );
  assign \new_[9727]_  = ~\new_[30119]_  & (~\new_[15484]_  | ~\new_[23245]_ );
  assign \new_[9728]_  = ~s8_ack_i | ~\new_[18080]_  | ~\new_[30341]_ ;
  assign \new_[9729]_  = ~s8_err_i | ~\new_[18080]_  | ~\new_[30341]_ ;
  assign \new_[9730]_  = ~s8_rty_i | ~\new_[18080]_  | ~\new_[30341]_ ;
  assign \new_[9731]_  = ~\new_[27862]_  & (~\new_[15516]_  | ~\new_[24307]_ );
  assign \new_[9732]_  = ~\new_[30090]_  & (~\new_[15043]_  | ~\new_[20443]_ );
  assign \new_[9733]_  = ~\new_[25158]_  & (~\new_[15519]_  | ~\new_[28230]_ );
  assign \new_[9734]_  = ~\new_[13674]_  & (~\new_[16524]_  | ~\new_[26464]_ );
  assign \new_[9735]_  = ~m2_stb_i | ~\new_[18080]_  | ~\new_[30341]_ ;
  assign \new_[9736]_  = ~m6_stb_i | ~\new_[16287]_  | ~\new_[29420]_ ;
  assign \new_[9737]_  = ~\new_[26486]_  & (~\new_[15231]_  | ~\new_[22798]_ );
  assign \new_[9738]_  = ~\new_[28636]_  & (~\new_[15236]_  | ~\new_[21410]_ );
  assign \new_[9739]_  = ~\new_[13675]_  & (~\new_[16457]_  | ~\new_[29548]_ );
  assign \new_[9740]_  = ~\new_[27893]_  & (~\new_[15520]_  | ~\new_[23087]_ );
  assign \new_[9741]_  = ~\new_[26462]_  & (~\new_[15521]_  | ~\new_[26757]_ );
  assign \new_[9742]_  = ~m4_stb_i | ~\new_[16307]_  | ~\new_[29185]_ ;
  assign \new_[9743]_  = ~\new_[29838]_  & (~\new_[15488]_  | ~\new_[27717]_ );
  assign \new_[9744]_  = ~\new_[13210]_  & (~\new_[32348]_  | ~\m0_addr_i[24] );
  assign \new_[9745]_  = ~\new_[27042]_  & (~\new_[15524]_  | ~\new_[24615]_ );
  assign \new_[9746]_  = ~\new_[14979]_  & ~\new_[13648]_ ;
  assign \new_[9747]_  = ~\new_[13676]_  & (~\new_[16334]_  | ~\new_[27811]_ );
  assign \new_[9748]_  = ~\new_[13677]_  & (~\new_[17350]_  | ~\new_[30027]_ );
  assign \new_[9749]_  = ~\new_[28044]_  & (~\new_[15490]_  | ~\new_[27198]_ );
  assign \new_[9750]_  = ~\new_[13678]_  & (~\new_[16327]_  | ~\new_[24527]_ );
  assign \new_[9751]_  = ~\new_[26456]_  & (~\new_[15256]_  | ~\new_[21454]_ );
  assign \new_[9752]_  = ~\new_[28066]_  & (~\new_[15047]_  | ~\new_[22823]_ );
  assign \new_[9753]_  = ~\new_[13679]_  & (~\new_[17300]_  | ~\new_[28901]_ );
  assign \new_[9754]_  = ~\new_[27864]_  & (~\new_[15527]_  | ~\new_[24709]_ );
  assign \new_[9755]_  = ~\new_[27840]_  & (~\new_[15596]_  | ~\new_[28370]_ );
  assign \new_[9756]_  = ~\new_[30134]_  & (~\new_[15132]_  | ~\new_[21564]_ );
  assign \new_[9757]_  = ~\new_[28327]_  & (~\new_[15139]_  | ~\new_[24327]_ );
  assign \new_[9758]_  = ~\new_[28354]_  & (~\new_[15147]_  | ~\new_[24353]_ );
  assign \new_[9759]_  = ~\new_[28603]_  & (~\new_[15155]_  | ~\new_[23277]_ );
  assign \new_[9760]_  = ~\new_[29847]_  & (~\new_[15162]_  | ~\new_[24473]_ );
  assign \new_[9761]_  = ~\new_[26480]_  & (~\new_[15172]_  | ~\new_[20511]_ );
  assign \new_[9762]_  = ~\new_[30056]_  & (~\new_[15192]_  | ~\new_[23172]_ );
  assign \new_[9763]_  = ~\new_[28325]_  & (~\new_[15202]_  | ~\new_[23220]_ );
  assign \new_[9764]_  = ~\new_[28316]_  & (~\new_[15211]_  | ~\new_[24267]_ );
  assign \new_[9765]_  = ~\new_[28060]_  & (~\new_[15220]_  | ~\new_[24338]_ );
  assign \new_[9766]_  = ~\new_[29236]_  & (~\new_[15227]_  | ~\new_[22953]_ );
  assign \new_[9767]_  = ~\new_[28620]_  & (~\new_[15237]_  | ~\new_[23233]_ );
  assign \new_[9768]_  = ~\new_[29838]_  & (~\new_[15244]_  | ~\new_[22894]_ );
  assign \new_[9769]_  = ~\new_[26642]_  & (~\new_[15598]_  | ~\new_[27662]_ );
  assign \new_[9770]_  = ~\new_[28094]_  & (~\new_[15049]_  | ~\new_[23042]_ );
  assign \new_[9771]_  = ~m7_stb_i | ~\new_[16295]_  | ~\new_[27337]_ ;
  assign \new_[9772]_  = ~s8_ack_i | ~\new_[16295]_  | ~\new_[27337]_ ;
  assign \new_[9773]_  = ~\new_[30406]_  & (~\new_[15564]_  | ~\new_[28740]_ );
  assign \new_[9774]_  = ~\new_[28094]_  & (~\new_[15261]_  | ~\new_[21854]_ );
  assign \new_[9775]_  = ~\new_[28300]_  & (~\new_[15263]_  | ~\new_[24397]_ );
  assign \new_[9776]_  = ~\new_[13205]_  & (~\new_[16322]_  | ~\m2_addr_i[24] );
  assign \new_[9777]_  = ~s8_rty_i | ~\new_[16295]_  | ~\new_[27337]_ ;
  assign \new_[9778]_  = (~\m2_data_i[30]  | ~\new_[17220]_ ) & (~\m1_data_i[30]  | ~\new_[17275]_ );
  assign \new_[9779]_  = ~m5_stb_i | ~\new_[16278]_  | ~\new_[29951]_ ;
  assign \new_[9780]_  = ~\new_[29034]_  | ~\new_[18027]_  | ~m0_stb_i;
  assign \new_[9781]_  = (~\m4_data_i[30]  | ~\new_[18881]_ ) & (~\m3_data_i[30]  | ~\new_[18207]_ );
  assign \new_[9782]_  = ~\new_[28814]_  & (~\new_[15570]_  | ~\new_[28115]_ );
  assign \new_[9783]_  = ~\new_[26801]_  & (~\new_[15275]_  | ~\new_[24123]_ );
  assign \new_[9784]_  = (~\m2_data_i[27]  | ~\new_[17220]_ ) & (~\m1_data_i[27]  | ~\new_[17275]_ );
  assign \new_[9785]_  = ~\new_[28780]_  & (~\new_[15575]_  | ~\new_[28492]_ );
  assign \new_[9786]_  = (~\m2_data_i[26]  | ~\new_[17220]_ ) & (~\m1_data_i[26]  | ~\new_[17274]_ );
  assign \new_[9787]_  = ~s8_err_i | ~\new_[16295]_  | ~\new_[27337]_ ;
  assign \new_[9788]_  = ~m7_stb_i | ~\new_[16296]_  | ~\new_[27347]_ ;
  assign \new_[9789]_  = ~\new_[29057]_  & (~\new_[15582]_  | ~\new_[28481]_ );
  assign \new_[9790]_  = (~\m2_data_i[25]  | ~\new_[17220]_ ) & (~\m1_data_i[25]  | ~\new_[17275]_ );
  assign \new_[9791]_  = (~\m4_data_i[25]  | ~\new_[17267]_ ) & (~\m3_data_i[25]  | ~\new_[18207]_ );
  assign \new_[9792]_  = (~\m2_data_i[24]  | ~\new_[17220]_ ) & (~\m1_data_i[24]  | ~\new_[17275]_ );
  assign \new_[9793]_  = (~\m4_data_i[24]  | ~\new_[18881]_ ) & (~\m3_data_i[24]  | ~\new_[18207]_ );
  assign \new_[9794]_  = ~\new_[26799]_  & (~\new_[15298]_  | ~\new_[28681]_ );
  assign \new_[9795]_  = ~\new_[26463]_  & (~\new_[15540]_  | ~\new_[19409]_ );
  assign \new_[9796]_  = (~\m2_data_i[22]  | ~\new_[17220]_ ) & (~\m1_data_i[22]  | ~\new_[17275]_ );
  assign \new_[9797]_  = (~\m4_data_i[22]  | ~\new_[18881]_ ) & (~\m3_data_i[22]  | ~\new_[18207]_ );
  assign \new_[9798]_  = ~\new_[29584]_  & (~\new_[15599]_  | ~\new_[28048]_ );
  assign \new_[9799]_  = (~\m2_data_i[21]  | ~\new_[17220]_ ) & (~\m1_data_i[21]  | ~\new_[17275]_ );
  assign \new_[9800]_  = (~\m4_data_i[21]  | ~\new_[17267]_ ) & (~\m3_data_i[21]  | ~\new_[18207]_ );
  assign \new_[9801]_  = ~\new_[26469]_  & (~\new_[15302]_  | ~\new_[27742]_ );
  assign \new_[9802]_  = (~\m2_data_i[20]  | ~\new_[17220]_ ) & (~\m1_data_i[20]  | ~\new_[17275]_ );
  assign \new_[9803]_  = ~\new_[29446]_  & (~\new_[15604]_  | ~\new_[28559]_ );
  assign \new_[9804]_  = (~\m4_data_i[20]  | ~\new_[17267]_ ) & (~\m3_data_i[20]  | ~\new_[18207]_ );
  assign \new_[9805]_  = (~\m2_data_i[19]  | ~\new_[17220]_ ) & (~\m1_data_i[19]  | ~\new_[17275]_ );
  assign \new_[9806]_  = (~\m4_data_i[19]  | ~\new_[17267]_ ) & (~\m3_data_i[19]  | ~\new_[18207]_ );
  assign \new_[9807]_  = (~\m2_data_i[17]  | ~\new_[17220]_ ) & (~\m1_data_i[17]  | ~\new_[17275]_ );
  assign \new_[9808]_  = ~\new_[26723]_  & (~\new_[15611]_  | ~\new_[28556]_ );
  assign \new_[9809]_  = (~\m2_data_i[16]  | ~\new_[17220]_ ) & (~\m1_data_i[16]  | ~\new_[17275]_ );
  assign \new_[9810]_  = ~\new_[29303]_  & (~\new_[15325]_  | ~\new_[28853]_ );
  assign \new_[9811]_  = (~\m2_data_i[15]  | ~\new_[17220]_ ) & (~\m1_data_i[15]  | ~\new_[17275]_ );
  assign \new_[9812]_  = (~\m2_data_i[14]  | ~\new_[17220]_ ) & (~\m1_data_i[14]  | ~\new_[17275]_ );
  assign \new_[9813]_  = ~\new_[29250]_  & (~\new_[15622]_  | ~\new_[28708]_ );
  assign \new_[9814]_  = (~\m2_data_i[12]  | ~\new_[17220]_ ) & (~\m1_data_i[12]  | ~\new_[17275]_ );
  assign \new_[9815]_  = ~\new_[29612]_  & (~\new_[15632]_  | ~\new_[28305]_ );
  assign \new_[9816]_  = ~\new_[27916]_  & (~\new_[15352]_  | ~\new_[23044]_ );
  assign \new_[9817]_  = (~\m5_data_i[23]  | ~\new_[16277]_ ) & (~\m6_data_i[23]  | ~\new_[18037]_ );
  assign \new_[9818]_  = ~\new_[28032]_  & (~\new_[15353]_  | ~\new_[22936]_ );
  assign \new_[9819]_  = ~\new_[27794]_  & (~\new_[15355]_  | ~\new_[29503]_ );
  assign \new_[9820]_  = ~\new_[26640]_  & (~\new_[15636]_  | ~\new_[28154]_ );
  assign \new_[9821]_  = (~m7_we_i | ~\new_[16295]_ ) & (~m0_we_i | ~\new_[18203]_ );
  assign \new_[9822]_  = ~\new_[29138]_  & (~\new_[15638]_  | ~\new_[28501]_ );
  assign \new_[9823]_  = ~\new_[13732]_  & ~\new_[15266]_ ;
  assign \new_[9824]_  = ~\new_[28264]_  & (~\new_[15377]_  | ~\new_[23030]_ );
  assign \new_[9825]_  = ~\new_[28334]_  & (~\new_[15379]_  | ~\new_[29124]_ );
  assign \new_[9826]_  = ~\new_[30073]_  & (~\new_[15646]_  | ~\new_[28475]_ );
  assign \new_[9827]_  = ~\new_[28418]_  | (~\new_[15673]_  & ~\new_[24008]_ );
  assign \new_[9828]_  = ~\new_[13206]_  & (~\new_[14895]_  | ~\m6_addr_i[24] );
  assign \new_[9829]_  = ~\new_[28693]_  | (~\new_[15675]_  & ~\new_[24998]_ );
  assign \new_[9830]_  = (~\m2_data_i[4]  | ~\new_[17220]_ ) & (~\m1_data_i[4]  | ~\new_[17274]_ );
  assign \new_[9831]_  = ~\new_[29547]_  | (~\new_[15677]_  & ~\new_[29211]_ );
  assign \new_[9832]_  = ~\new_[26672]_  | (~\new_[15679]_  & ~\new_[26775]_ );
  assign \new_[9833]_  = ~\new_[28701]_  | (~\new_[15680]_  & ~\new_[27572]_ );
  assign \new_[9834]_  = ~\new_[28971]_  | (~\new_[15681]_  & ~\new_[27530]_ );
  assign \new_[9835]_  = ~\new_[28126]_  | (~\new_[15682]_  & ~\new_[23162]_ );
  assign \new_[9836]_  = ~\new_[29760]_  | (~\new_[15683]_  & ~\new_[29761]_ );
  assign \new_[9837]_  = ~\new_[29273]_  | (~\new_[15685]_  & ~\new_[26405]_ );
  assign \new_[9838]_  = ~\new_[30237]_  | (~\new_[15686]_  & ~\new_[24787]_ );
  assign \new_[9839]_  = (~\m2_data_i[0]  | ~\new_[17220]_ ) & (~\m1_data_i[0]  | ~\new_[17275]_ );
  assign \new_[9840]_  = ~\new_[28827]_  | (~\new_[15687]_  & ~\new_[26743]_ );
  assign \new_[9841]_  = ~\new_[29237]_  | (~\new_[15689]_  & ~\new_[25127]_ );
  assign \new_[9842]_  = ~\new_[29362]_  | (~\new_[15690]_  & ~\new_[26885]_ );
  assign \new_[9843]_  = ~\new_[28758]_  | (~\new_[15691]_  & ~\new_[27581]_ );
  assign \new_[9844]_  = ~\new_[28662]_  | (~\new_[15692]_  & ~\new_[27442]_ );
  assign \new_[9845]_  = ~\new_[29110]_  | (~\new_[15693]_  & ~\new_[28472]_ );
  assign \new_[9846]_  = ~\new_[29279]_  | (~\new_[15694]_  & ~\new_[26561]_ );
  assign \new_[9847]_  = ~\new_[29348]_  | (~\new_[15695]_  & ~\new_[26578]_ );
  assign \new_[9848]_  = ~\new_[29301]_  | (~\new_[15696]_  & ~\new_[27965]_ );
  assign \new_[9849]_  = ~\new_[29187]_  | (~\new_[15697]_  & ~\new_[24550]_ );
  assign \new_[9850]_  = ~\new_[30281]_  | (~\new_[15698]_  & ~\new_[24554]_ );
  assign \new_[9851]_  = ~\new_[29538]_  | (~\new_[15699]_  & ~\new_[28571]_ );
  assign \new_[9852]_  = ~\new_[28261]_  | (~\new_[15700]_  & ~\new_[23997]_ );
  assign \new_[9853]_  = ~\new_[29085]_  | (~\new_[15701]_  & ~\new_[26509]_ );
  assign \new_[9854]_  = ~\new_[29041]_  | (~\new_[15702]_  & ~\new_[23924]_ );
  assign \new_[9855]_  = ~\new_[26639]_  | (~\new_[15708]_  & ~\new_[26829]_ );
  assign \new_[9856]_  = ~\new_[26977]_  | (~\new_[15703]_  & ~\new_[27267]_ );
  assign \new_[9857]_  = ~\new_[28970]_  | (~\new_[15704]_  & ~\new_[26272]_ );
  assign \new_[9858]_  = ~\new_[28077]_  | (~\new_[15705]_  & ~\new_[24337]_ );
  assign \new_[9859]_  = (~\m2_addr_i[21]  | ~\new_[17220]_ ) & (~\m1_addr_i[21]  | ~\new_[17275]_ );
  assign \new_[9860]_  = ~\new_[29542]_  | (~\new_[15707]_  & ~\new_[27649]_ );
  assign \new_[9861]_  = ~\new_[27000]_  | (~\new_[15709]_  & ~\new_[26752]_ );
  assign \new_[9862]_  = (~\m2_addr_i[20]  | ~\new_[17220]_ ) & (~\m1_addr_i[20]  | ~\new_[17274]_ );
  assign \new_[9863]_  = ~\new_[29155]_  | (~\new_[15711]_  & ~\new_[28099]_ );
  assign \new_[9864]_  = ~\new_[29278]_  & (~\new_[15407]_  | ~\new_[21514]_ );
  assign \new_[9865]_  = (~\m2_addr_i[19]  | ~\new_[17220]_ ) & (~\m1_addr_i[19]  | ~\new_[17274]_ );
  assign \new_[9866]_  = ~\new_[29659]_  & (~\new_[15409]_  | ~\new_[23021]_ );
  assign \new_[9867]_  = (~\m2_addr_i[18]  | ~\new_[17220]_ ) & (~\m1_addr_i[18]  | ~\new_[17275]_ );
  assign \new_[9868]_  = (~\m4_addr_i[18]  | ~\new_[17267]_ ) & (~\m3_addr_i[18]  | ~\new_[18207]_ );
  assign \new_[9869]_  = (~\m2_addr_i[17]  | ~\new_[17220]_ ) & (~\m1_addr_i[17]  | ~\new_[17275]_ );
  assign \new_[9870]_  = (~\m4_addr_i[17]  | ~\new_[17267]_ ) & (~\m3_addr_i[17]  | ~\new_[18207]_ );
  assign \new_[9871]_  = ~\new_[27925]_  & (~\new_[15410]_  | ~\new_[17403]_ );
  assign \new_[9872]_  = ~\new_[26677]_  & (~\new_[15411]_  | ~\new_[29419]_ );
  assign \new_[9873]_  = (~\m2_addr_i[16]  | ~\new_[17220]_ ) & (~\m1_addr_i[16]  | ~\new_[17275]_ );
  assign \new_[9874]_  = ~\new_[26652]_  & (~\new_[15529]_  | ~\new_[21368]_ );
  assign \new_[9875]_  = ~\new_[26774]_  & (~\new_[15530]_  | ~\new_[19417]_ );
  assign \new_[9876]_  = (~\m2_addr_i[14]  | ~\new_[17220]_ ) & (~\m1_addr_i[14]  | ~\new_[17275]_ );
  assign \new_[9877]_  = (~\m2_addr_i[13]  | ~\new_[17220]_ ) & (~\m1_addr_i[13]  | ~\new_[17275]_ );
  assign \new_[9878]_  = ~\new_[28304]_  & (~\new_[15531]_  | ~\new_[21429]_ );
  assign \new_[9879]_  = (~\m4_addr_i[13]  | ~\new_[18881]_ ) & (~\m3_addr_i[13]  | ~\new_[18207]_ );
  assign \new_[9880]_  = ~\new_[26925]_  & (~\new_[15416]_  | ~\new_[17405]_ );
  assign \new_[9881]_  = (~\m2_addr_i[11]  | ~\new_[17220]_ ) & (~\m1_addr_i[11]  | ~\new_[17275]_ );
  assign \new_[9882]_  = ~\new_[30144]_  & (~\new_[15418]_  | ~\new_[18425]_ );
  assign \new_[9883]_  = (~\m4_addr_i[11]  | ~\new_[17267]_ ) & (~\m3_addr_i[11]  | ~\new_[18207]_ );
  assign \new_[9884]_  = ~\new_[27395]_  & (~\new_[15533]_  | ~\new_[22695]_ );
  assign \new_[9885]_  = (~\m2_addr_i[9]  | ~\new_[17220]_ ) & (~\m1_addr_i[9]  | ~\new_[17275]_ );
  assign \new_[9886]_  = (~\m2_addr_i[8]  | ~\new_[17220]_ ) & (~\m1_addr_i[8]  | ~\new_[17275]_ );
  assign \new_[9887]_  = (~\m4_addr_i[8]  | ~\new_[18881]_ ) & (~\m3_addr_i[8]  | ~\new_[18207]_ );
  assign \new_[9888]_  = ~\new_[26598]_  & (~\new_[15422]_  | ~\new_[20460]_ );
  assign \new_[9889]_  = ~\new_[28691]_  & (~\new_[15534]_  | ~\new_[19411]_ );
  assign \new_[9890]_  = (~\m2_addr_i[7]  | ~\new_[17220]_ ) & (~\m1_addr_i[7]  | ~\new_[17275]_ );
  assign \new_[9891]_  = ~\new_[28995]_  & (~\new_[15536]_  | ~\new_[21376]_ );
  assign \new_[9892]_  = (~\m4_addr_i[7]  | ~\new_[17267]_ ) & (~\m3_addr_i[7]  | ~\new_[18207]_ );
  assign \new_[9893]_  = ~\new_[28775]_  & (~\new_[15423]_  | ~\new_[20718]_ );
  assign \new_[9894]_  = ~\new_[26799]_  & (~\new_[15424]_  | ~\new_[28537]_ );
  assign \new_[9895]_  = (~\m4_addr_i[6]  | ~\new_[17267]_ ) & (~\m3_addr_i[6]  | ~\new_[18207]_ );
  assign \new_[9896]_  = ~\new_[28754]_  & (~\new_[15426]_  | ~\new_[20451]_ );
  assign \new_[9897]_  = ~\new_[26643]_  & (~\new_[15537]_  | ~\new_[21386]_ );
  assign \new_[9898]_  = (~\new_[31095]_  | ~\new_[17220]_ ) & (~\m1_addr_i[5]  | ~\new_[17274]_ );
  assign \new_[9899]_  = ~\new_[26447]_  & (~\new_[15539]_  | ~\new_[21408]_ );
  assign \new_[9900]_  = (~\m2_addr_i[4]  | ~\new_[17220]_ ) & (~\m1_addr_i[4]  | ~\new_[17274]_ );
  assign \new_[9901]_  = ~\new_[26645]_  & (~\new_[15429]_  | ~\new_[20484]_ );
  assign \new_[9902]_  = (~\new_[31399]_  | ~\new_[17220]_ ) & (~\m1_addr_i[3]  | ~\new_[17274]_ );
  assign \new_[9903]_  = ~\new_[26754]_  & (~\new_[15541]_  | ~\new_[22755]_ );
  assign \new_[9904]_  = ~\new_[26583]_  & (~\new_[15543]_  | ~\new_[22805]_ );
  assign \new_[9905]_  = ~\new_[28088]_  & (~\new_[15544]_  | ~\new_[22790]_ );
  assign \new_[9906]_  = (~\m4_addr_i[1]  | ~\new_[17267]_ ) & (~\m3_addr_i[1]  | ~\new_[18207]_ );
  assign \new_[9907]_  = ~\new_[29646]_  & (~\new_[15430]_  | ~\new_[23178]_ );
  assign \new_[9908]_  = (~\m5_data_i[7]  | ~\new_[20544]_ ) & (~\m6_data_i[7]  | ~\new_[17213]_ );
  assign \new_[9909]_  = ~\new_[28848]_  & (~\new_[15545]_  | ~\new_[22756]_ );
  assign \new_[9910]_  = ~\new_[29154]_  & (~\new_[15547]_  | ~\new_[22651]_ );
  assign \new_[9911]_  = (~\m2_sel_i[3]  | ~\new_[17220]_ ) & (~\m1_sel_i[3]  | ~\new_[17275]_ );
  assign \new_[9912]_  = ~\new_[26644]_  & (~\new_[15548]_  | ~\new_[22783]_ );
  assign \new_[9913]_  = (~\m4_sel_i[0]  | ~\new_[17267]_ ) & (~\m3_sel_i[0]  | ~\new_[18207]_ );
  assign \new_[9914]_  = ~\new_[29303]_  & (~\new_[15437]_  | ~\new_[28940]_ );
  assign \new_[9915]_  = ~\new_[28936]_  & (~\new_[15438]_  | ~\new_[21542]_ );
  assign \new_[9916]_  = (~\m1_data_i[2]  | ~\new_[18192]_ ) & (~\m0_data_i[2]  | ~\new_[14834]_ );
  assign \new_[9917]_  = ~\new_[29932]_  & (~\new_[15441]_  | ~\new_[21458]_ );
  assign \new_[9918]_  = (~\m4_data_i[29]  | ~\new_[17268]_ ) & (~\m3_data_i[29]  | ~\new_[20567]_ );
  assign \new_[9919]_  = (~\m4_data_i[27]  | ~\new_[17268]_ ) & (~\m3_data_i[27]  | ~\new_[18853]_ );
  assign \new_[9920]_  = ~\new_[28053]_  & (~\new_[15552]_  | ~\new_[22802]_ );
  assign \new_[9921]_  = (~\m4_data_i[26]  | ~\new_[17268]_ ) & (~\m3_data_i[26]  | ~\new_[18853]_ );
  assign \new_[9922]_  = (~\m4_data_i[25]  | ~\new_[17268]_ ) & (~\m3_data_i[25]  | ~\new_[20567]_ );
  assign \new_[9923]_  = ~\new_[11651]_ ;
  assign \new_[9924]_  = ~\new_[27794]_  & (~\new_[15445]_  | ~\new_[29136]_ );
  assign \new_[9925]_  = (~\m4_data_i[24]  | ~\new_[17268]_ ) & (~\m3_data_i[24]  | ~\new_[20567]_ );
  assign \new_[9926]_  = ~\new_[28257]_  & (~\new_[15448]_  | ~\new_[22679]_ );
  assign \new_[9927]_  = ~\new_[27240]_  & (~\new_[15553]_  | ~\new_[22421]_ );
  assign \new_[9928]_  = (~\m4_data_i[23]  | ~\new_[17268]_ ) & (~\m3_data_i[23]  | ~\new_[20567]_ );
  assign \new_[9929]_  = ~\new_[14852]_ ;
  assign \new_[9930]_  = ~\new_[28141]_  & (~\new_[15554]_  | ~\new_[22829]_ );
  assign \new_[9931]_  = ~\new_[26765]_  & (~\new_[15450]_  | ~\new_[17411]_ );
  assign \new_[9932]_  = ~\new_[27910]_  & (~\new_[15451]_  | ~\new_[29399]_ );
  assign \new_[9933]_  = ~\new_[28804]_  & (~\new_[15452]_  | ~\new_[20488]_ );
  assign \new_[9934]_  = (~\m4_data_i[21]  | ~\new_[17268]_ ) & (~\m3_data_i[21]  | ~\new_[20567]_ );
  assign \new_[9935]_  = ~\new_[27888]_  & (~\new_[15556]_  | ~\new_[18423]_ );
  assign \new_[9936]_  = (~\m4_data_i[20]  | ~\new_[17268]_ ) & (~\m3_data_i[20]  | ~\new_[18852]_ );
  assign \new_[9937]_  = ~\new_[28334]_  & (~\new_[15454]_  | ~\new_[29336]_ );
  assign \new_[9938]_  = (~\m4_data_i[19]  | ~\new_[17268]_ ) & (~\m3_data_i[19]  | ~\new_[20567]_ );
  assign \new_[9939]_  = ~\new_[29297]_  & (~\new_[15455]_  | ~\new_[23029]_ );
  assign \new_[9940]_  = ~\new_[28426]_  & (~\new_[15559]_  | ~\new_[21369]_ );
  assign \new_[9941]_  = (~\m4_data_i[18]  | ~\new_[17268]_ ) & (~\m3_data_i[18]  | ~\new_[18854]_ );
  assign \new_[9942]_  = (~\m4_data_i[17]  | ~\new_[17268]_ ) & (~\m3_data_i[17]  | ~\new_[18853]_ );
  assign \new_[9943]_  = (~m2_we_i | ~\new_[17193]_ ) & (~m1_we_i | ~\new_[18916]_ );
  assign \new_[9944]_  = (~\m5_data_i[16]  | ~\new_[18743]_ ) & (~\m6_data_i[16]  | ~\new_[16289]_ );
  assign \new_[9945]_  = ~\new_[27874]_  & (~\new_[15458]_  | ~\new_[20452]_ );
  assign \new_[9946]_  = ~\new_[26713]_  & (~\new_[15562]_  | ~\new_[22841]_ );
  assign \new_[9947]_  = (~\m5_data_i[15]  | ~\new_[20542]_ ) & (~\m6_data_i[15]  | ~\new_[16289]_ );
  assign \new_[9948]_  = (~\m4_data_i[15]  | ~\new_[17268]_ ) & (~\m3_data_i[15]  | ~\new_[20567]_ );
  assign \new_[9949]_  = (~\m5_data_i[14]  | ~\new_[20542]_ ) & (~\m6_data_i[14]  | ~\new_[16289]_ );
  assign \new_[9950]_  = ~\new_[27873]_  & (~\new_[15593]_  | ~\new_[23132]_ );
  assign \new_[9951]_  = (~\m4_data_i[14]  | ~\new_[17268]_ ) & (~\m3_data_i[14]  | ~\new_[20567]_ );
  assign \new_[9952]_  = ~\new_[28095]_  & (~\new_[15594]_  | ~\new_[20482]_ );
  assign \new_[9953]_  = (~\m5_data_i[13]  | ~\new_[18743]_ ) & (~\m6_data_i[13]  | ~\new_[16289]_ );
  assign \new_[9954]_  = (~\m4_data_i[13]  | ~\new_[17268]_ ) & (~\m3_data_i[13]  | ~\new_[20567]_ );
  assign \new_[9955]_  = ~\new_[28773]_  & (~\new_[15135]_  | ~\new_[21437]_ );
  assign \new_[9956]_  = (~\m4_data_i[12]  | ~\new_[17268]_ ) & (~\m3_data_i[12]  | ~\new_[20567]_ );
  assign \new_[9957]_  = ~\new_[26892]_  & (~\new_[15136]_  | ~\new_[22526]_ );
  assign \new_[9958]_  = ~\new_[28119]_  & (~\new_[15137]_  | ~\new_[21430]_ );
  assign \new_[9959]_  = (~\m4_data_i[11]  | ~\new_[17268]_ ) & (~\m3_data_i[11]  | ~\new_[18852]_ );
  assign \new_[9960]_  = (~\m5_data_i[10]  | ~\new_[18743]_ ) & (~\m6_data_i[10]  | ~\new_[16289]_ );
  assign \new_[9961]_  = (~\m4_data_i[10]  | ~\new_[17268]_ ) & (~\m3_data_i[10]  | ~\new_[20567]_ );
  assign \new_[9962]_  = (~\new_[15280]_  | ~\new_[29146]_ ) & (~\new_[22719]_  | ~\new_[29146]_ );
  assign \new_[9963]_  = (~\m4_data_i[9]  | ~\new_[17268]_ ) & (~\m3_data_i[9]  | ~\new_[18854]_ );
  assign \new_[9964]_  = (~\m4_data_i[8]  | ~\new_[17268]_ ) & (~\m3_data_i[8]  | ~\new_[18852]_ );
  assign \new_[9965]_  = (~\m4_data_i[7]  | ~\new_[17268]_ ) & (~\m3_data_i[7]  | ~\new_[18853]_ );
  assign \new_[9966]_  = (~\new_[15285]_  | ~\new_[29733]_ ) & (~\new_[23686]_  | ~\new_[29733]_ );
  assign \new_[9967]_  = (~\m7_addr_i[18]  | ~\new_[17240]_ ) & (~\m6_addr_i[18]  | ~\new_[18819]_ );
  assign \new_[9968]_  = ~\new_[27867]_  & (~\new_[15159]_  | ~\new_[20423]_ );
  assign \new_[9969]_  = (~\m4_data_i[6]  | ~\new_[17268]_ ) & (~\m3_data_i[6]  | ~\new_[20567]_ );
  assign \new_[9970]_  = (~\m4_data_i[5]  | ~\new_[17268]_ ) & (~\m3_data_i[5]  | ~\new_[18852]_ );
  assign \new_[9971]_  = (~\m4_data_i[4]  | ~\new_[17268]_ ) & (~\m3_data_i[4]  | ~\new_[18853]_ );
  assign \new_[9972]_  = (~\new_[15296]_  | ~\new_[29011]_ ) & (~\new_[26151]_  | ~\new_[29011]_ );
  assign \new_[9973]_  = ~\new_[23129]_  & (~\new_[15176]_  | ~\new_[26176]_ );
  assign \new_[9974]_  = (~\m4_data_i[3]  | ~\new_[17268]_ ) & (~\m3_data_i[3]  | ~\new_[18854]_ );
  assign \new_[9975]_  = (~\m4_data_i[2]  | ~\new_[17268]_ ) & (~\m3_data_i[2]  | ~\new_[18852]_ );
  assign \new_[9976]_  = (~\m5_data_i[2]  | ~\new_[18743]_ ) & (~\m6_data_i[2]  | ~\new_[16289]_ );
  assign \new_[9977]_  = (~\m5_data_i[1]  | ~\new_[20542]_ ) & (~\m6_data_i[1]  | ~\new_[16289]_ );
  assign \new_[9978]_  = (~\new_[15309]_  | ~\new_[28980]_ ) & (~\new_[25640]_  | ~\new_[28980]_ );
  assign \new_[9979]_  = (~\m4_data_i[1]  | ~\new_[17268]_ ) & (~\m3_data_i[1]  | ~\new_[18852]_ );
  assign \new_[9980]_  = (~\new_[15314]_  | ~\new_[29661]_ ) & (~\new_[22449]_  | ~\new_[29661]_ );
  assign \new_[9981]_  = (~\m4_data_i[0]  | ~\new_[17268]_ ) & (~\m3_data_i[0]  | ~\new_[18854]_ );
  assign \new_[9982]_  = (~\new_[17268]_  | ~\m4_addr_i[31] ) & (~\new_[18854]_  | ~\m3_addr_i[31] );
  assign \new_[9983]_  = (~\new_[15321]_  | ~\new_[29292]_ ) & (~\new_[24221]_  | ~\new_[29292]_ );
  assign \new_[9984]_  = (~\new_[17268]_  | ~\m4_addr_i[30] ) & (~\new_[18854]_  | ~\m3_addr_i[30] );
  assign \new_[9985]_  = (~\new_[17268]_  | ~\m4_addr_i[29] ) & (~\new_[20567]_  | ~\m3_addr_i[29] );
  assign \new_[9986]_  = ~\new_[28195]_  & (~\new_[15199]_  | ~\new_[22571]_ );
  assign \new_[9987]_  = (~\new_[15327]_  | ~\new_[29980]_ ) & (~\new_[21362]_  | ~\new_[29980]_ );
  assign \new_[9988]_  = (~\new_[17268]_  | ~\m4_addr_i[28] ) & (~\new_[18853]_  | ~\m3_addr_i[28] );
  assign \new_[9989]_  = (~\m4_addr_i[2]  | ~\new_[17260]_ ) & (~\m3_addr_i[2]  | ~\new_[18175]_ );
  assign \new_[9990]_  = (~\new_[15330]_  | ~\new_[29106]_ ) & (~\new_[26074]_  | ~\new_[29106]_ );
  assign \new_[9991]_  = (~\m5_sel_i[0]  | ~\new_[17202]_ ) & (~\m4_sel_i[0]  | ~\new_[17271]_ );
  assign \new_[9992]_  = (~\m5_data_i[28]  | ~\new_[18747]_ ) & (~\m6_data_i[28]  | ~\new_[17213]_ );
  assign \new_[9993]_  = ~\new_[29152]_  & (~\new_[15208]_  | ~\new_[20383]_ );
  assign \new_[9994]_  = ~\new_[28638]_  & (~\new_[15209]_  | ~\new_[21348]_ );
  assign \new_[9995]_  = (~\new_[17268]_  | ~\m4_addr_i[27] ) & (~\new_[18854]_  | ~\m3_addr_i[27] );
  assign \new_[9996]_  = (~\new_[17268]_  | ~\m4_addr_i[26] ) & (~\new_[18854]_  | ~\m3_addr_i[26] );
  assign \new_[9997]_  = (~\new_[17268]_  | ~\m4_addr_i[25] ) & (~\new_[18854]_  | ~\m3_addr_i[25] );
  assign \new_[9998]_  = (~\new_[15347]_  | ~\new_[30082]_ ) & (~\new_[22780]_  | ~\new_[30082]_ );
  assign \new_[9999]_  = (~\new_[17268]_  | ~\m4_addr_i[24] ) & (~\new_[20567]_  | ~\m3_addr_i[24] );
  assign \new_[10000]_  = (~\m5_addr_i[23]  | ~\new_[18743]_ ) & (~\m6_addr_i[23]  | ~\new_[16289]_ );
  assign \new_[10001]_  = ~\new_[29643]_  & (~\new_[15225]_  | ~\new_[22837]_ );
  assign \new_[10002]_  = ~\new_[13526]_ ;
  assign \new_[10003]_  = (~\m4_addr_i[23]  | ~\new_[17268]_ ) & (~\m3_addr_i[23]  | ~\new_[20567]_ );
  assign \new_[10004]_  = (~\m4_addr_i[22]  | ~\new_[17268]_ ) & (~\m3_addr_i[22]  | ~\new_[18852]_ );
  assign \new_[10005]_  = (~\m5_data_i[18]  | ~\new_[18750]_ ) & (~\m6_data_i[18]  | ~\new_[17213]_ );
  assign \new_[10006]_  = (~\new_[31095]_  | ~\new_[17193]_ ) & (~\m1_addr_i[5]  | ~\new_[18916]_ );
  assign \new_[10007]_  = ~\new_[27885]_  & (~\new_[15233]_  | ~\new_[22834]_ );
  assign \new_[10008]_  = ~\new_[28790]_  & (~\new_[15235]_  | ~\new_[22781]_ );
  assign \new_[10009]_  = (~\m2_addr_i[2]  | ~\new_[17193]_ ) & (~\new_[31477]_  | ~\new_[18916]_ );
  assign \new_[10010]_  = (~\m4_addr_i[20]  | ~\new_[17268]_ ) & (~\m3_addr_i[20]  | ~\new_[20567]_ );
  assign \new_[10011]_  = (~\m4_addr_i[18]  | ~\new_[17268]_ ) & (~\m3_addr_i[18]  | ~\new_[20567]_ );
  assign \new_[10012]_  = (~\m4_addr_i[17]  | ~\new_[17268]_ ) & (~\m3_addr_i[17]  | ~\new_[18852]_ );
  assign \new_[10013]_  = ~\new_[29095]_  & (~\new_[15250]_  | ~\new_[21385]_ );
  assign \new_[10014]_  = ~\new_[13530]_ ;
  assign \new_[10015]_  = ~\new_[27889]_  & (~\new_[15257]_  | ~\new_[22816]_ );
  assign \new_[10016]_  = ~\new_[28035]_  & (~\new_[15258]_  | ~\new_[21382]_ );
  assign \new_[10017]_  = ~\new_[13209]_  & (~\new_[32348]_  | ~\m0_addr_i[25] );
  assign \new_[10018]_  = (~\m4_addr_i[12]  | ~\new_[17268]_ ) & (~\m3_addr_i[12]  | ~\new_[18853]_ );
  assign \new_[10019]_  = (~\m4_addr_i[11]  | ~\new_[17268]_ ) & (~\m3_addr_i[11]  | ~\new_[18853]_ );
  assign \new_[10020]_  = (~\m4_addr_i[9]  | ~\new_[17268]_ ) & (~\m3_addr_i[9]  | ~\new_[18853]_ );
  assign \new_[10021]_  = ~\new_[28172]_  & (~\new_[15581]_  | ~\new_[22454]_ );
  assign \new_[10022]_  = (~\new_[15068]_  | ~\new_[29161]_ ) & (~\new_[21261]_  | ~\new_[29161]_ );
  assign \new_[10023]_  = (~\m4_addr_i[8]  | ~\new_[17268]_ ) & (~\m3_addr_i[8]  | ~\new_[19597]_ );
  assign \new_[10024]_  = (~\m5_data_i[24]  | ~\new_[18756]_ ) & (~\m6_data_i[24]  | ~\new_[17213]_ );
  assign \new_[10025]_  = (~\m4_addr_i[7]  | ~\new_[17268]_ ) & (~\m3_addr_i[7]  | ~\new_[18852]_ );
  assign \new_[10026]_  = ~\new_[26508]_  & (~\new_[15587]_  | ~\new_[23054]_ );
  assign \new_[10027]_  = ~\new_[26598]_  & (~\new_[15588]_  | ~\new_[20450]_ );
  assign \new_[10028]_  = (~\new_[15074]_  | ~\new_[29993]_ ) & (~\new_[24199]_  | ~\new_[29993]_ );
  assign \new_[10029]_  = (~\m4_addr_i[6]  | ~\new_[17268]_ ) & (~\m3_addr_i[6]  | ~\new_[18853]_ );
  assign \new_[10030]_  = (~\new_[15075]_  | ~\new_[29532]_ ) & (~\new_[22738]_  | ~\new_[29532]_ );
  assign \new_[10031]_  = (~\m4_addr_i[5]  | ~\new_[17268]_ ) & (~\m3_addr_i[5]  | ~\new_[19597]_ );
  assign \new_[10032]_  = (~\new_[15083]_  | ~\new_[29580]_ ) & (~\new_[22708]_  | ~\new_[29580]_ );
  assign \new_[10033]_  = (~\new_[15084]_  | ~\new_[29131]_ ) & (~\new_[22801]_  | ~\new_[29131]_ );
  assign \new_[10034]_  = (~\m4_addr_i[4]  | ~\new_[17268]_ ) & (~\m3_addr_i[4]  | ~\new_[18854]_ );
  assign \new_[10035]_  = ~\new_[28706]_  & (~\new_[15605]_  | ~\new_[21582]_ );
  assign \new_[10036]_  = (~\new_[16296]_  | ~\m7_addr_i[25] ) & (~\new_[18766]_  | ~\m0_addr_i[25] );
  assign \new_[10037]_  = ~\new_[29646]_  & (~\new_[15607]_  | ~\new_[24384]_ );
  assign \new_[10038]_  = (~\new_[15090]_  | ~\new_[28843]_ ) & (~\new_[21389]_  | ~\new_[28843]_ );
  assign \new_[10039]_  = (~\m4_addr_i[3]  | ~\new_[17268]_ ) & (~\m3_addr_i[3]  | ~\new_[18854]_ );
  assign \new_[10040]_  = (~\new_[15092]_  | ~\new_[29074]_ ) & (~\new_[22725]_  | ~\new_[29074]_ );
  assign \new_[10041]_  = (~\m4_addr_i[2]  | ~\new_[17268]_ ) & (~\m3_addr_i[2]  | ~\new_[18854]_ );
  assign \new_[10042]_  = (~\new_[16296]_  | ~\m7_addr_i[26] ) & (~\new_[18764]_  | ~\m0_addr_i[26] );
  assign \new_[10043]_  = (~\new_[15096]_  | ~\new_[29731]_ ) & (~\new_[24223]_  | ~\new_[29731]_ );
  assign \new_[10044]_  = (~\m5_addr_i[0]  | ~\new_[18743]_ ) & (~\m6_addr_i[0]  | ~\new_[16289]_ );
  assign \new_[10045]_  = (~\new_[15102]_  | ~\new_[30175]_ ) & (~\new_[24195]_  | ~\new_[30175]_ );
  assign \new_[10046]_  = (~\m4_addr_i[0]  | ~\new_[17268]_ ) & (~\m3_addr_i[0]  | ~\new_[20567]_ );
  assign \new_[10047]_  = (~\m5_data_i[1]  | ~\new_[18015]_ ) & (~\m6_data_i[1]  | ~\new_[17229]_ );
  assign \new_[10048]_  = ~\new_[29407]_  & (~\new_[15621]_  | ~\new_[20498]_ );
  assign \new_[10049]_  = (~\m4_sel_i[1]  | ~\new_[17268]_ ) & (~\m3_sel_i[1]  | ~\new_[18853]_ );
  assign \new_[10050]_  = (~\new_[15112]_  | ~\new_[30288]_ ) & (~\new_[21417]_  | ~\new_[30288]_ );
  assign \new_[10051]_  = (~m4_we_i | ~\new_[17268]_ ) & (~m3_we_i | ~\new_[18853]_ );
  assign \new_[10052]_  = (~\m5_addr_i[0]  | ~\new_[17202]_ ) & (~\m4_addr_i[0]  | ~\new_[17271]_ );
  assign \new_[10053]_  = (~\new_[15116]_  | ~\new_[27798]_ ) & (~\new_[24235]_  | ~\new_[27798]_ );
  assign \new_[10054]_  = (~\m5_data_i[31]  | ~\new_[17204]_ ) & (~\m6_data_i[31]  | ~\new_[16288]_ );
  assign \new_[10055]_  = (~\m2_data_i[30]  | ~\new_[16292]_ ) & (~\m1_data_i[30]  | ~\new_[18890]_ );
  assign \new_[10056]_  = (~\m4_data_i[30]  | ~\new_[17262]_ ) & (~\m3_data_i[30]  | ~\new_[18125]_ );
  assign \new_[10057]_  = (~\new_[15120]_  | ~\new_[29535]_ ) & (~\new_[22583]_  | ~\new_[29535]_ );
  assign \new_[10058]_  = (~\m7_data_i[29]  | ~\new_[16295]_ ) & (~\m0_data_i[29]  | ~\new_[18204]_ );
  assign \new_[10059]_  = (~\m4_data_i[29]  | ~\new_[17262]_ ) & (~\m3_data_i[29]  | ~\new_[17247]_ );
  assign \new_[10060]_  = ~\new_[28264]_  & (~\new_[15639]_  | ~\new_[22876]_ );
  assign \new_[10061]_  = (~\m5_data_i[29]  | ~\new_[17205]_ ) & (~\m6_data_i[29]  | ~\new_[14836]_ );
  assign \new_[10062]_  = ~\new_[29297]_  & (~\new_[15640]_  | ~\new_[21570]_ );
  assign \new_[10063]_  = (~\new_[15124]_  | ~\new_[30190]_ ) & (~\new_[21395]_  | ~\new_[30190]_ );
  assign \new_[10064]_  = (~\m7_data_i[28]  | ~\new_[16295]_ ) & (~\m0_data_i[28]  | ~\new_[18204]_ );
  assign \new_[10065]_  = (~\m5_data_i[28]  | ~\new_[17205]_ ) & (~\m6_data_i[28]  | ~\new_[14836]_ );
  assign \new_[10066]_  = (~\m7_data_i[27]  | ~\new_[16295]_ ) & (~\m0_data_i[27]  | ~\new_[18204]_ );
  assign \new_[10067]_  = ~\new_[24742]_  & (~\new_[15647]_  | ~\new_[22160]_ );
  assign \new_[10068]_  = (~\m4_data_i[27]  | ~\new_[17262]_ ) & (~\m3_data_i[27]  | ~\new_[17247]_ );
  assign \new_[10069]_  = ~\new_[27874]_  & (~\new_[15648]_  | ~\new_[20465]_ );
  assign \new_[10070]_  = (~\m5_data_i[27]  | ~\new_[17205]_ ) & (~\m6_data_i[27]  | ~\new_[18033]_ );
  assign \new_[10071]_  = (~\m5_data_i[26]  | ~\new_[17204]_ ) & (~\m6_data_i[26]  | ~\new_[16288]_ );
  assign \new_[10072]_  = ~\new_[28095]_  & (~\new_[15427]_  | ~\new_[19511]_ );
  assign \new_[10073]_  = (~\m2_data_i[25]  | ~\new_[16292]_ ) & (~\m1_data_i[25]  | ~\new_[19621]_ );
  assign \new_[10074]_  = (~\m4_data_i[25]  | ~\new_[17262]_ ) & (~\m3_data_i[25]  | ~\new_[17247]_ );
  assign \new_[10075]_  = (~\m5_data_i[25]  | ~\new_[17205]_ ) & (~\m6_data_i[25]  | ~\new_[16288]_ );
  assign \new_[10076]_  = (~\m4_addr_i[3]  | ~\new_[17260]_ ) & (~\m3_addr_i[3]  | ~\new_[18175]_ );
  assign \new_[10077]_  = ~\new_[13991]_  | ~\new_[28093]_ ;
  assign \new_[10078]_  = (~\m7_data_i[23]  | ~\new_[16295]_ ) & (~\m0_data_i[23]  | ~\new_[18204]_ );
  assign \new_[10079]_  = (~\m4_data_i[23]  | ~\new_[17262]_ ) & (~\m3_data_i[23]  | ~\new_[17247]_ );
  assign \new_[10080]_  = ~\new_[13812]_  | ~\new_[27989]_ ;
  assign \new_[10081]_  = (~\m4_sel_i[1]  | ~\new_[17260]_ ) & (~\m3_sel_i[1]  | ~\new_[18175]_ );
  assign \new_[10082]_  = (~\m5_data_i[23]  | ~\new_[17204]_ ) & (~\m6_data_i[23]  | ~\new_[14836]_ );
  assign \new_[10083]_  = ~\new_[14031]_  | ~\new_[28910]_ ;
  assign \new_[10084]_  = (~\m5_data_i[22]  | ~\new_[17205]_ ) & (~\m6_data_i[22]  | ~\new_[18033]_ );
  assign \new_[10085]_  = (~\m5_data_i[21]  | ~\new_[17204]_ ) & (~\m6_data_i[21]  | ~\new_[16288]_ );
  assign \new_[10086]_  = (~\m4_data_i[21]  | ~\new_[17262]_ ) & (~\m3_data_i[21]  | ~\new_[17246]_ );
  assign \new_[10087]_  = (~\m7_data_i[6]  | ~\new_[16296]_ ) & (~\m0_data_i[6]  | ~\new_[20545]_ );
  assign \new_[10088]_  = ~\new_[14058]_  | ~\new_[29686]_ ;
  assign \new_[10089]_  = (~\m5_data_i[20]  | ~\new_[17204]_ ) & (~\m6_data_i[20]  | ~\new_[16288]_ );
  assign \new_[10090]_  = (~\m4_data_i[20]  | ~\new_[17262]_ ) & (~\m3_data_i[20]  | ~\new_[17246]_ );
  assign \new_[10091]_  = (~\new_[31399]_  | ~\new_[17193]_ ) & (~\m1_addr_i[3]  | ~\new_[18916]_ );
  assign \new_[10092]_  = (~\m5_data_i[19]  | ~\new_[17205]_ ) & (~\m6_data_i[19]  | ~\new_[16288]_ );
  assign \new_[10093]_  = (~\m2_data_i[17]  | ~\new_[16292]_ ) & (~\m1_data_i[17]  | ~\new_[19621]_ );
  assign \new_[10094]_  = (~\m4_data_i[17]  | ~\new_[17262]_ ) & (~\m3_data_i[17]  | ~\new_[17247]_ );
  assign \new_[10095]_  = (~\m2_sel_i[1]  | ~\new_[17193]_ ) & (~\m1_sel_i[1]  | ~\new_[18917]_ );
  assign \new_[10096]_  = (~\m5_data_i[17]  | ~\new_[17205]_ ) & (~\m6_data_i[17]  | ~\new_[16288]_ );
  assign \new_[10097]_  = ~\new_[14158]_  | ~\new_[28115]_ ;
  assign \new_[10098]_  = (~\m7_data_i[16]  | ~\new_[16295]_ ) & (~\m0_data_i[16]  | ~\new_[18204]_ );
  assign \new_[10099]_  = (~\m4_data_i[16]  | ~\new_[17262]_ ) & (~\m3_data_i[16]  | ~\new_[17247]_ );
  assign \new_[10100]_  = (~\m5_data_i[16]  | ~\new_[17204]_ ) & (~\m6_data_i[16]  | ~\new_[16288]_ );
  assign \new_[10101]_  = (~\m7_data_i[15]  | ~\new_[16295]_ ) & (~\m0_data_i[15]  | ~\new_[18203]_ );
  assign \new_[10102]_  = (~\m5_data_i[15]  | ~\new_[18760]_ ) & (~\m6_data_i[15]  | ~\new_[14836]_ );
  assign \new_[10103]_  = (~\m7_data_i[14]  | ~\new_[16295]_ ) & (~\m0_data_i[14]  | ~\new_[18203]_ );
  assign \new_[10104]_  = (~\m5_data_i[14]  | ~\new_[18760]_ ) & (~\m6_data_i[14]  | ~\new_[14836]_ );
  assign \new_[10105]_  = (~\m7_data_i[13]  | ~\new_[16295]_ ) & (~\m0_data_i[13]  | ~\new_[18203]_ );
  assign \new_[10106]_  = (~\m4_data_i[13]  | ~\new_[17262]_ ) & (~\m3_data_i[13]  | ~\new_[17245]_ );
  assign \new_[10107]_  = (~\m5_data_i[13]  | ~\new_[17205]_ ) & (~\m6_data_i[13]  | ~\new_[14836]_ );
  assign \new_[10108]_  = (~\m2_data_i[12]  | ~\new_[16292]_ ) & (~\m1_data_i[12]  | ~\new_[19621]_ );
  assign \new_[10109]_  = (~\m7_data_i[12]  | ~\new_[16295]_ ) & (~\m0_data_i[12]  | ~\new_[18203]_ );
  assign \new_[10110]_  = ~\new_[13990]_  | ~\new_[28210]_ ;
  assign \new_[10111]_  = (~\m4_data_i[12]  | ~\new_[17262]_ ) & (~\m3_data_i[12]  | ~\new_[17247]_ );
  assign \new_[10112]_  = (~\m5_data_i[12]  | ~\new_[18760]_ ) & (~\m6_data_i[12]  | ~\new_[14836]_ );
  assign \new_[10113]_  = (~\m2_data_i[11]  | ~\new_[16292]_ ) & (~\m1_data_i[11]  | ~\new_[19621]_ );
  assign \new_[10114]_  = (~\m7_data_i[11]  | ~\new_[16295]_ ) & (~\m0_data_i[11]  | ~\new_[18203]_ );
  assign \new_[10115]_  = (~\m4_data_i[11]  | ~\new_[17262]_ ) & (~\m3_data_i[11]  | ~\new_[18846]_ );
  assign \new_[10116]_  = (~\m5_data_i[11]  | ~\new_[17205]_ ) & (~\m6_data_i[11]  | ~\new_[14836]_ );
  assign \new_[10117]_  = (~\m2_data_i[10]  | ~\new_[16292]_ ) & (~\m1_data_i[10]  | ~\new_[19621]_ );
  assign \new_[10118]_  = (~\m7_data_i[10]  | ~\new_[16295]_ ) & (~\m0_data_i[10]  | ~\new_[18203]_ );
  assign \new_[10119]_  = ~\new_[14131]_  | ~\new_[28231]_ ;
  assign \new_[10120]_  = ~\new_[13995]_  | ~\new_[28231]_ ;
  assign \new_[10121]_  = (~\m5_data_i[10]  | ~\new_[17205]_ ) & (~\m6_data_i[10]  | ~\new_[14836]_ );
  assign \new_[10122]_  = (~\m2_data_i[9]  | ~\new_[16292]_ ) & (~\m1_data_i[9]  | ~\new_[18167]_ );
  assign \new_[10123]_  = (~\m7_data_i[9]  | ~\new_[16295]_ ) & (~\m0_data_i[9]  | ~\new_[18203]_ );
  assign \new_[10124]_  = (~\m5_data_i[9]  | ~\new_[18760]_ ) & (~\m6_data_i[9]  | ~\new_[16288]_ );
  assign \new_[10125]_  = ~\new_[14132]_  | ~\new_[26769]_ ;
  assign \new_[10126]_  = (~\m7_data_i[8]  | ~\new_[16295]_ ) & (~\m0_data_i[8]  | ~\new_[18204]_ );
  assign \new_[10127]_  = (~\m7_data_i[7]  | ~\new_[16295]_ ) & (~\m0_data_i[7]  | ~\new_[18203]_ );
  assign \new_[10128]_  = ~\new_[14134]_  | ~\new_[28496]_ ;
  assign \new_[10129]_  = (~\m5_data_i[7]  | ~\new_[18760]_ ) & (~\m6_data_i[7]  | ~\new_[14836]_ );
  assign \new_[10130]_  = ~\new_[14001]_  | ~\new_[28014]_ ;
  assign \new_[10131]_  = ~\new_[14002]_  | ~\new_[28158]_ ;
  assign \new_[10132]_  = (~\m2_data_i[6]  | ~\new_[16292]_ ) & (~\m1_data_i[6]  | ~\new_[18167]_ );
  assign \new_[10133]_  = (~\m4_data_i[6]  | ~\new_[17262]_ ) & (~\m3_data_i[6]  | ~\new_[18846]_ );
  assign \new_[10134]_  = (~\m5_data_i[6]  | ~\new_[17205]_ ) & (~\m6_data_i[6]  | ~\new_[14836]_ );
  assign \new_[10135]_  = (~\m7_data_i[5]  | ~\new_[16295]_ ) & (~\m0_data_i[5]  | ~\new_[18203]_ );
  assign \new_[10136]_  = (~\m4_data_i[28]  | ~\new_[17264]_ ) & (~\m3_data_i[28]  | ~\new_[18128]_ );
  assign \new_[10137]_  = ~\new_[14112]_  | ~\new_[24256]_ ;
  assign \new_[10138]_  = ~\new_[14171]_  | ~\new_[28048]_ ;
  assign \new_[10139]_  = (~\m5_data_i[5]  | ~\new_[17205]_ ) & (~\m6_data_i[5]  | ~\new_[16288]_ );
  assign \new_[10140]_  = ~\new_[14009]_  | ~\new_[28494]_ ;
  assign \new_[10141]_  = ~\new_[14115]_  | ~\new_[24295]_ ;
  assign \new_[10142]_  = ~\new_[14176]_  | ~\new_[28559]_ ;
  assign \new_[10143]_  = (~\m5_data_i[3]  | ~\new_[18760]_ ) & (~\m6_data_i[3]  | ~\new_[14836]_ );
  assign \new_[10144]_  = ~\new_[14138]_  | ~\new_[28416]_ ;
  assign \new_[10145]_  = (~\m7_data_i[2]  | ~\new_[16295]_ ) & (~\m0_data_i[2]  | ~\new_[18203]_ );
  assign \new_[10146]_  = (~\m5_data_i[2]  | ~\new_[17205]_ ) & (~\m6_data_i[2]  | ~\new_[14836]_ );
  assign \new_[10147]_  = ~\new_[14020]_  | ~\new_[28674]_ ;
  assign \new_[10148]_  = (~\m4_data_i[0]  | ~\new_[17262]_ ) & (~\m3_data_i[0]  | ~\new_[18125]_ );
  assign \new_[10149]_  = (~\new_[16292]_  | ~\new_[31486]_ ) & (~\new_[18890]_  | ~\new_[31308]_ );
  assign \new_[10150]_  = ~\new_[14028]_  | ~\new_[28097]_ ;
  assign \new_[10151]_  = (~\new_[16295]_  | ~\new_[31531]_ ) & (~\new_[18204]_  | ~\new_[31481]_ );
  assign \new_[10152]_  = (~\new_[17262]_  | ~\m4_addr_i[29] ) & (~\new_[17247]_  | ~\m3_addr_i[29] );
  assign \new_[10153]_  = (~\new_[16292]_  | ~\new_[31547]_ ) & (~\new_[18890]_  | ~\new_[31458]_ );
  assign \new_[10154]_  = (~\new_[16295]_  | ~\m7_addr_i[27] ) & (~\new_[18204]_  | ~\m0_addr_i[27] );
  assign \new_[10155]_  = (~\new_[16292]_  | ~\m2_addr_i[27] ) & (~\new_[18167]_  | ~\m1_addr_i[27] );
  assign \new_[10156]_  = (~\new_[16292]_  | ~\m2_addr_i[26] ) & (~\new_[18167]_  | ~\m1_addr_i[26] );
  assign \new_[10157]_  = (~\new_[16295]_  | ~\m7_addr_i[25] ) & (~\new_[18204]_  | ~\m0_addr_i[25] );
  assign \new_[10158]_  = (~\new_[16292]_  | ~\m2_addr_i[25] ) & (~\new_[18167]_  | ~\m1_addr_i[25] );
  assign \new_[10159]_  = ~\new_[14040]_  | ~\new_[28564]_ ;
  assign \new_[10160]_  = \new_[14306]_  | \new_[25065]_ ;
  assign \new_[10161]_  = ~\new_[14149]_  | ~\new_[27130]_ ;
  assign \new_[10162]_  = (~\new_[17262]_  | ~\m4_addr_i[24] ) & (~\new_[17247]_  | ~\m3_addr_i[24] );
  assign \new_[10163]_  = (~\m5_addr_i[23]  | ~\new_[17204]_ ) & (~\m6_addr_i[23]  | ~\new_[16288]_ );
  assign \new_[10164]_  = (~\m5_addr_i[22]  | ~\new_[17204]_ ) & (~\m6_addr_i[22]  | ~\new_[16288]_ );
  assign \new_[10165]_  = (~\m4_addr_i[22]  | ~\new_[17262]_ ) & (~\m3_addr_i[22]  | ~\new_[17247]_ );
  assign \new_[10166]_  = (~\m7_addr_i[21]  | ~\new_[16295]_ ) & (~\m0_addr_i[21]  | ~\new_[18204]_ );
  assign \new_[10167]_  = (~\m4_addr_i[21]  | ~\new_[17262]_ ) & (~\m3_addr_i[21]  | ~\new_[17245]_ );
  assign \new_[10168]_  = (~\m4_data_i[27]  | ~\new_[17265]_ ) & (~\m3_data_i[27]  | ~\new_[17248]_ );
  assign \new_[10169]_  = ~\new_[14185]_  | ~\new_[28154]_ ;
  assign \new_[10170]_  = (~\m5_addr_i[21]  | ~\new_[17205]_ ) & (~\m6_addr_i[21]  | ~\new_[18033]_ );
  assign \new_[10171]_  = (~\m5_addr_i[20]  | ~\new_[17204]_ ) & (~\m6_addr_i[20]  | ~\new_[16288]_ );
  assign \new_[10172]_  = \new_[14318]_  | \new_[26416]_ ;
  assign \new_[10173]_  = (~\m4_addr_i[20]  | ~\new_[17262]_ ) & (~\m3_addr_i[20]  | ~\new_[18846]_ );
  assign \new_[10174]_  = \new_[14321]_  | \new_[25386]_ ;
  assign \new_[10175]_  = (~\m5_addr_i[19]  | ~\new_[17204]_ ) & (~\m6_addr_i[19]  | ~\new_[16288]_ );
  assign \new_[10176]_  = ~\new_[14121]_  | ~\new_[24440]_ ;
  assign \new_[10177]_  = ~\new_[14160]_  | ~\new_[28501]_ ;
  assign \new_[10178]_  = ~\new_[14141]_  | ~\new_[28587]_ ;
  assign \new_[10179]_  = (~\m4_addr_i[19]  | ~\new_[17262]_ ) & (~\m3_addr_i[19]  | ~\new_[17247]_ );
  assign \new_[10180]_  = (~\m2_sel_i[2]  | ~\new_[17193]_ ) & (~\m1_sel_i[2]  | ~\new_[19633]_ );
  assign \new_[10181]_  = (~\m5_data_i[30]  | ~\new_[18749]_ ) & (~\m6_data_i[30]  | ~\new_[17213]_ );
  assign \new_[10182]_  = (~\m5_data_i[22]  | ~\new_[18004]_ ) & (~\m6_data_i[22]  | ~\new_[17241]_ );
  assign \new_[10183]_  = (~\m2_addr_i[18]  | ~\new_[16292]_ ) & (~\m1_addr_i[18]  | ~\new_[19621]_ );
  assign \new_[10184]_  = (~\m2_addr_i[8]  | ~\new_[16292]_ ) & (~\m1_addr_i[8]  | ~\new_[18890]_ );
  assign \new_[10185]_  = (~\m5_addr_i[18]  | ~\new_[17204]_ ) & (~\m6_addr_i[18]  | ~\new_[14836]_ );
  assign \new_[10186]_  = (~\m4_addr_i[18]  | ~\new_[17262]_ ) & (~\m3_addr_i[18]  | ~\new_[17246]_ );
  assign \new_[10187]_  = ~\new_[14122]_  | ~\new_[24316]_ ;
  assign \new_[10188]_  = ~\new_[14190]_  | ~\new_[28475]_ ;
  assign \new_[10189]_  = ~\new_[14154]_  | ~\new_[28368]_ ;
  assign \new_[10190]_  = (~\m5_addr_i[17]  | ~\new_[17205]_ ) & (~\m6_addr_i[17]  | ~\new_[18033]_ );
  assign \new_[10191]_  = ~\new_[14068]_  | ~\new_[28368]_ ;
  assign \new_[10192]_  = (~\m2_addr_i[16]  | ~\new_[16292]_ ) & (~\m1_addr_i[16]  | ~\new_[18890]_ );
  assign \new_[10193]_  = (~\m4_addr_i[16]  | ~\new_[17262]_ ) & (~\m3_addr_i[16]  | ~\new_[17247]_ );
  assign \new_[10194]_  = (~\m5_addr_i[16]  | ~\new_[17205]_ ) & (~\m6_addr_i[16]  | ~\new_[14836]_ );
  assign \new_[10195]_  = (~\m2_addr_i[4]  | ~\new_[17193]_ ) & (~\m1_addr_i[4]  | ~\new_[18917]_ );
  assign \new_[10196]_  = ~\new_[14156]_  | ~\new_[28193]_ ;
  assign \new_[10197]_  = ~\new_[14194]_  | ~\new_[28740]_ ;
  assign \new_[10198]_  = (~\m5_addr_i[15]  | ~\new_[17205]_ ) & (~\m6_addr_i[15]  | ~\new_[18033]_ );
  assign \new_[10199]_  = (~\m7_addr_i[14]  | ~\new_[16295]_ ) & (~\m0_addr_i[14]  | ~\new_[18204]_ );
  assign \new_[10200]_  = (~\m4_addr_i[14]  | ~\new_[17262]_ ) & (~\m3_addr_i[14]  | ~\new_[17246]_ );
  assign \new_[10201]_  = (~\new_[17260]_  | ~\m4_addr_i[26] ) & (~\new_[18175]_  | ~\m3_addr_i[26] );
  assign \new_[10202]_  = (~\m5_addr_i[14]  | ~\new_[17205]_ ) & (~\m6_addr_i[14]  | ~\new_[14836]_ );
  assign \new_[10203]_  = ~\new_[22461]_  | ~\new_[13793]_ ;
  assign \new_[10204]_  = (~\new_[17241]_  | ~\m6_addr_i[27] ) & (~\new_[18004]_  | ~\m5_addr_i[27] );
  assign \new_[10205]_  = (~\m7_addr_i[13]  | ~\new_[16295]_ ) & (~\m0_addr_i[13]  | ~\new_[18204]_ );
  assign \new_[10206]_  = (~\m4_addr_i[13]  | ~\new_[17262]_ ) & (~\m3_addr_i[13]  | ~\new_[17246]_ );
  assign \new_[10207]_  = (~\m5_addr_i[13]  | ~\new_[17205]_ ) & (~\m6_addr_i[13]  | ~\new_[14836]_ );
  assign \new_[10208]_  = (~\m7_sel_i[2]  | ~\new_[16296]_ ) & (~\m0_sel_i[2]  | ~\new_[18764]_ );
  assign \new_[10209]_  = (~\m5_addr_i[12]  | ~\new_[17204]_ ) & (~\m6_addr_i[12]  | ~\new_[16288]_ );
  assign \new_[10210]_  = (~\m7_addr_i[11]  | ~\new_[16295]_ ) & (~\m0_addr_i[11]  | ~\new_[18204]_ );
  assign \new_[10211]_  = (~\m4_addr_i[11]  | ~\new_[17262]_ ) & (~\m3_addr_i[11]  | ~\new_[17246]_ );
  assign \new_[10212]_  = ~\new_[27875]_  & (~\new_[15719]_  | ~\new_[21528]_ );
  assign \new_[10213]_  = (~\m5_addr_i[11]  | ~\new_[17205]_ ) & (~\m6_addr_i[11]  | ~\new_[18033]_ );
  assign \new_[10214]_  = (~\m2_addr_i[10]  | ~\new_[16292]_ ) & (~\m1_addr_i[10]  | ~\new_[19621]_ );
  assign \new_[10215]_  = (~\m4_addr_i[10]  | ~\new_[17262]_ ) & (~\m3_addr_i[10]  | ~\new_[17247]_ );
  assign \new_[10216]_  = (~\m5_addr_i[10]  | ~\new_[17204]_ ) & (~\m6_addr_i[10]  | ~\new_[18033]_ );
  assign \new_[10217]_  = (~\m7_addr_i[9]  | ~\new_[16295]_ ) & (~\m0_addr_i[9]  | ~\new_[18203]_ );
  assign \new_[10218]_  = (~\m5_addr_i[9]  | ~\new_[17205]_ ) & (~\m6_addr_i[9]  | ~\new_[14836]_ );
  assign \new_[10219]_  = (~\m4_addr_i[8]  | ~\new_[17262]_ ) & (~\m3_addr_i[8]  | ~\new_[18846]_ );
  assign \new_[10220]_  = (~\m5_data_i[11]  | ~\new_[18757]_ ) & (~\m6_data_i[11]  | ~\new_[17213]_ );
  assign \new_[10221]_  = (~\m5_addr_i[8]  | ~\new_[18760]_ ) & (~\m6_addr_i[8]  | ~\new_[16288]_ );
  assign \new_[10222]_  = (~\m7_addr_i[7]  | ~\new_[16295]_ ) & (~\m0_addr_i[7]  | ~\new_[18203]_ );
  assign \new_[10223]_  = (~\m4_addr_i[7]  | ~\new_[17262]_ ) & (~\m3_addr_i[7]  | ~\new_[17247]_ );
  assign \new_[10224]_  = ~\new_[26800]_  & (~\new_[15723]_  | ~\new_[21500]_ );
  assign \new_[10225]_  = (~\m5_addr_i[7]  | ~\new_[17205]_ ) & (~\m6_addr_i[7]  | ~\new_[14836]_ );
  assign \new_[10226]_  = (~\m7_addr_i[6]  | ~\new_[16295]_ ) & (~\m0_addr_i[6]  | ~\new_[18203]_ );
  assign \new_[10227]_  = (~\m5_addr_i[6]  | ~\new_[17205]_ ) & (~\m6_addr_i[6]  | ~\new_[18033]_ );
  assign \new_[10228]_  = (~\m7_addr_i[5]  | ~\new_[16295]_ ) & (~\new_[31848]_  | ~\new_[18203]_ );
  assign \new_[10229]_  = ~\new_[29232]_  & (~\new_[15725]_  | ~\new_[24211]_ );
  assign \new_[10230]_  = (~\m5_addr_i[5]  | ~\new_[17205]_ ) & (~\m6_addr_i[5]  | ~\new_[14836]_ );
  assign \new_[10231]_  = (~\m7_addr_i[1]  | ~\new_[17239]_ ) & (~\m6_addr_i[1]  | ~\new_[18089]_ );
  assign \new_[10232]_  = (~\m7_addr_i[4]  | ~\new_[16295]_ ) & (~\m0_addr_i[4]  | ~\new_[18203]_ );
  assign \new_[10233]_  = (~\m5_addr_i[4]  | ~\new_[17205]_ ) & (~\m6_addr_i[4]  | ~\new_[14836]_ );
  assign \new_[10234]_  = ~\new_[26628]_  & (~\new_[15728]_  | ~\new_[21471]_ );
  assign \new_[10235]_  = (~\new_[31726]_  | ~\new_[16295]_ ) & (~\m0_addr_i[3]  | ~\new_[18203]_ );
  assign \new_[10236]_  = ~\new_[29982]_  & (~\new_[15732]_  | ~\new_[22940]_ );
  assign \new_[10237]_  = (~\m5_addr_i[3]  | ~\new_[17205]_ ) & (~\m6_addr_i[3]  | ~\new_[14836]_ );
  assign \new_[10238]_  = ~\new_[28617]_  & (~\new_[15734]_  | ~\new_[22734]_ );
  assign \new_[10239]_  = (~\m7_addr_i[2]  | ~\new_[16295]_ ) & (~\m0_addr_i[2]  | ~\new_[18203]_ );
  assign \new_[10240]_  = (~\m4_addr_i[2]  | ~\new_[17262]_ ) & (~\m3_addr_i[2]  | ~\new_[17247]_ );
  assign \new_[10241]_  = (~\m2_addr_i[1]  | ~\new_[16292]_ ) & (~\m1_addr_i[1]  | ~\new_[18890]_ );
  assign \new_[10242]_  = (~\m4_addr_i[1]  | ~\new_[17262]_ ) & (~\m3_addr_i[1]  | ~\new_[17245]_ );
  assign \new_[10243]_  = ~\new_[16355]_  | ~\new_[13804]_ ;
  assign \new_[10244]_  = (~\m5_addr_i[1]  | ~\new_[17204]_ ) & (~\m6_addr_i[1]  | ~\new_[16288]_ );
  assign \new_[10245]_  = ~\new_[22479]_  | ~\new_[13808]_ ;
  assign \new_[10246]_  = (~\m5_addr_i[0]  | ~\new_[17205]_ ) & (~\m6_addr_i[0]  | ~\new_[16288]_ );
  assign \new_[10247]_  = (~\m7_sel_i[3]  | ~\new_[16295]_ ) & (~\m0_sel_i[3]  | ~\new_[19643]_ );
  assign \new_[10248]_  = ~\new_[29638]_  & (~\new_[15739]_  | ~\new_[21367]_ );
  assign \new_[10249]_  = (~\m2_sel_i[1]  | ~\new_[16292]_ ) & (~\m1_sel_i[1]  | ~\new_[19621]_ );
  assign \new_[10250]_  = (~\m4_sel_i[1]  | ~\new_[17262]_ ) & (~\m3_sel_i[1]  | ~\new_[17247]_ );
  assign \new_[10251]_  = (~\m5_sel_i[1]  | ~\new_[17204]_ ) & (~\m6_sel_i[1]  | ~\new_[16288]_ );
  assign \new_[10252]_  = ~\new_[26904]_  | (~\new_[15747]_  & ~\new_[23526]_ );
  assign \new_[10253]_  = ~\new_[28777]_  & (~\new_[15748]_  | ~\new_[19424]_ );
  assign \new_[10254]_  = (~\m5_sel_i[0]  | ~\new_[17205]_ ) & (~\m6_sel_i[0]  | ~\new_[14836]_ );
  assign \new_[10255]_  = ~\new_[20374]_  | ~\new_[13815]_ ;
  assign \new_[10256]_  = (~m5_we_i | ~\new_[18760]_ ) & (~m6_we_i | ~\new_[16288]_ );
  assign \new_[10257]_  = (~m4_we_i | ~\new_[17262]_ ) & (~m3_we_i | ~\new_[18125]_ );
  assign \new_[10258]_  = (~\m5_data_i[31]  | ~\new_[16276]_ ) & (~\m6_data_i[31]  | ~\new_[18036]_ );
  assign \new_[10259]_  = (~\m2_data_i[31]  | ~\new_[17222]_ ) & (~\m1_data_i[31]  | ~\new_[17273]_ );
  assign \new_[10260]_  = (~\m5_data_i[30]  | ~\new_[16276]_ ) & (~\m6_data_i[30]  | ~\new_[19559]_ );
  assign \new_[10261]_  = (~\m2_data_i[30]  | ~\new_[17222]_ ) & (~\m1_data_i[30]  | ~\new_[18177]_ );
  assign \new_[10262]_  = ~\new_[28759]_  & (~\new_[15752]_  | ~\new_[21345]_ );
  assign \new_[10263]_  = (~\m7_data_i[30]  | ~\new_[18111]_ ) & (~\m0_data_i[30]  | ~\new_[18027]_ );
  assign \new_[10264]_  = (~\m7_data_i[29]  | ~\new_[18111]_ ) & (~\m0_data_i[29]  | ~\new_[18027]_ );
  assign \new_[10265]_  = ~\new_[29330]_  | (~\new_[15754]_  & ~\new_[23566]_ );
  assign \new_[10266]_  = (~\m5_data_i[29]  | ~\new_[16276]_ ) & (~\m6_data_i[29]  | ~\new_[18036]_ );
  assign \new_[10267]_  = ~\new_[30306]_  & (~\new_[15755]_  | ~\new_[19450]_ );
  assign \new_[10268]_  = ~\new_[21287]_  | ~\new_[13819]_ ;
  assign \new_[10269]_  = (~\m4_data_i[29]  | ~\new_[16308]_ ) & (~\m3_data_i[29]  | ~\new_[17249]_ );
  assign \new_[10270]_  = (~\m2_data_i[28]  | ~\new_[17222]_ ) & (~\m1_data_i[28]  | ~\new_[18177]_ );
  assign \new_[10271]_  = (~\m5_data_i[28]  | ~\new_[16277]_ ) & (~\m6_data_i[28]  | ~\new_[18036]_ );
  assign \new_[10272]_  = (~\m4_data_i[28]  | ~\new_[16308]_ ) & (~\m3_data_i[28]  | ~\new_[17249]_ );
  assign \new_[10273]_  = (~\m7_data_i[28]  | ~\new_[18111]_ ) & (~\m0_data_i[28]  | ~\new_[18027]_ );
  assign \new_[10274]_  = (~\m5_data_i[27]  | ~\new_[16276]_ ) & (~\m6_data_i[27]  | ~\new_[19559]_ );
  assign \new_[10275]_  = (~\m2_data_i[27]  | ~\new_[17222]_ ) & (~\m1_data_i[27]  | ~\new_[17273]_ );
  assign \new_[10276]_  = (~\m4_data_i[27]  | ~\new_[16308]_ ) & (~\m3_data_i[27]  | ~\new_[17249]_ );
  assign \new_[10277]_  = ~\new_[30171]_  & (~\new_[15758]_  | ~\new_[21363]_ );
  assign \new_[10278]_  = (~\m7_data_i[27]  | ~\new_[18111]_ ) & (~\m0_data_i[27]  | ~\new_[18027]_ );
  assign \new_[10279]_  = (~\m5_data_i[26]  | ~\new_[16276]_ ) & (~\m6_data_i[26]  | ~\new_[19559]_ );
  assign \new_[10280]_  = ~\new_[16349]_  | ~\new_[13820]_ ;
  assign \new_[10281]_  = (~\m2_data_i[25]  | ~\new_[17222]_ ) & (~\m1_data_i[25]  | ~\new_[18177]_ );
  assign \new_[10282]_  = ~\new_[18417]_  | ~\new_[13823]_ ;
  assign \new_[10283]_  = (~\m5_data_i[25]  | ~\new_[16277]_ ) & (~\m6_data_i[25]  | ~\new_[18037]_ );
  assign \new_[10284]_  = (~\m2_data_i[24]  | ~\new_[17222]_ ) & (~\m1_data_i[24]  | ~\new_[18906]_ );
  assign \new_[10285]_  = (~\m7_data_i[24]  | ~\new_[18111]_ ) & (~\m0_data_i[24]  | ~\new_[18027]_ );
  assign \new_[10286]_  = ~\new_[28387]_  & (~\new_[15761]_  | ~\new_[22704]_ );
  assign \new_[10287]_  = (~\m5_data_i[24]  | ~\new_[16277]_ ) & (~\m6_data_i[24]  | ~\new_[18037]_ );
  assign \new_[10288]_  = (~\m7_data_i[23]  | ~\new_[18111]_ ) & (~\m0_data_i[23]  | ~\new_[18027]_ );
  assign \new_[10289]_  = (~\m2_data_i[23]  | ~\new_[17222]_ ) & (~\m1_data_i[23]  | ~\new_[18906]_ );
  assign \new_[10290]_  = (~\m4_data_i[23]  | ~\new_[16308]_ ) & (~\m3_data_i[23]  | ~\new_[17249]_ );
  assign \new_[10291]_  = (~\m7_data_i[22]  | ~\new_[18111]_ ) & (~\m0_data_i[22]  | ~\new_[18027]_ );
  assign \new_[10292]_  = (~\m2_data_i[22]  | ~\new_[17222]_ ) & (~\m1_data_i[22]  | ~\new_[17273]_ );
  assign \new_[10293]_  = (~\m5_data_i[22]  | ~\new_[16277]_ ) & (~\m6_data_i[22]  | ~\new_[18037]_ );
  assign \new_[10294]_  = (~\m7_data_i[21]  | ~\new_[18111]_ ) & (~\m0_data_i[21]  | ~\new_[18027]_ );
  assign \new_[10295]_  = (~\m5_data_i[21]  | ~\new_[16277]_ ) & (~\m6_data_i[21]  | ~\new_[18038]_ );
  assign \new_[10296]_  = (~\m2_data_i[20]  | ~\new_[17222]_ ) & (~\m1_data_i[20]  | ~\new_[17273]_ );
  assign \new_[10297]_  = (~\m5_data_i[20]  | ~\new_[16277]_ ) & (~\m6_data_i[20]  | ~\new_[18038]_ );
  assign \new_[10298]_  = (~\m5_data_i[19]  | ~\new_[16276]_ ) & (~\m6_data_i[19]  | ~\new_[18035]_ );
  assign \new_[10299]_  = (~\m7_data_i[19]  | ~\new_[18111]_ ) & (~\m0_data_i[19]  | ~\new_[18027]_ );
  assign \new_[10300]_  = (~\m2_data_i[19]  | ~\new_[17222]_ ) & (~\m1_data_i[19]  | ~\new_[17273]_ );
  assign \new_[10301]_  = ~\new_[29843]_  & (~\new_[15767]_  | ~\new_[22726]_ );
  assign \new_[10302]_  = (~\m2_data_i[18]  | ~\new_[17222]_ ) & (~\m1_data_i[18]  | ~\new_[17273]_ );
  assign \new_[10303]_  = (~\m4_data_i[18]  | ~\new_[16307]_ ) & (~\m3_data_i[18]  | ~\new_[17249]_ );
  assign \new_[10304]_  = (~\m2_data_i[17]  | ~\new_[17222]_ ) & (~\m1_data_i[17]  | ~\new_[18177]_ );
  assign \new_[10305]_  = (~\m5_data_i[17]  | ~\new_[16276]_ ) & (~\m6_data_i[17]  | ~\new_[18036]_ );
  assign \new_[10306]_  = ~\new_[26705]_  & (~\new_[15769]_  | ~\new_[21460]_ );
  assign \new_[10307]_  = (~\m4_data_i[17]  | ~\new_[16308]_ ) & (~\m3_data_i[17]  | ~\new_[17249]_ );
  assign \new_[10308]_  = ~\new_[30119]_  & (~\new_[15772]_  | ~\new_[21899]_ );
  assign \new_[10309]_  = (~\m5_data_i[16]  | ~\new_[16276]_ ) & (~\m6_data_i[16]  | ~\new_[18035]_ );
  assign \new_[10310]_  = (~\m7_data_i[16]  | ~\new_[18111]_ ) & (~\m0_data_i[16]  | ~\new_[18027]_ );
  assign \new_[10311]_  = ~\new_[28292]_  & (~\new_[15773]_  | ~\new_[21432]_ );
  assign \new_[10312]_  = (~\m2_data_i[15]  | ~\new_[17222]_ ) & (~\m1_data_i[15]  | ~\new_[17273]_ );
  assign \new_[10313]_  = (~\m5_data_i[15]  | ~\new_[18008]_ ) & (~\m6_data_i[15]  | ~\new_[19559]_ );
  assign \new_[10314]_  = (~\m4_data_i[15]  | ~\new_[16308]_ ) & (~\m3_data_i[15]  | ~\new_[17249]_ );
  assign \new_[10315]_  = (~\m2_data_i[14]  | ~\new_[17222]_ ) & (~\m1_data_i[14]  | ~\new_[18177]_ );
  assign \new_[10316]_  = (~\m7_data_i[14]  | ~\new_[18111]_ ) & (~\m0_data_i[14]  | ~\new_[18027]_ );
  assign \new_[10317]_  = (~\m5_data_i[14]  | ~\new_[16278]_ ) & (~\m6_data_i[14]  | ~\new_[19559]_ );
  assign \new_[10318]_  = (~\m7_data_i[13]  | ~\new_[18111]_ ) & (~\m0_data_i[13]  | ~\new_[18027]_ );
  assign \new_[10319]_  = (~\m2_data_i[13]  | ~\new_[17222]_ ) & (~\m1_data_i[13]  | ~\new_[18177]_ );
  assign \new_[10320]_  = (~\m5_data_i[13]  | ~\new_[16278]_ ) & (~\m6_data_i[13]  | ~\new_[18040]_ );
  assign \new_[10321]_  = (~\m7_data_i[12]  | ~\new_[18111]_ ) & (~\m0_data_i[12]  | ~\new_[18027]_ );
  assign \new_[10322]_  = (~\m2_data_i[12]  | ~\new_[17222]_ ) & (~\m1_data_i[12]  | ~\new_[17273]_ );
  assign \new_[10323]_  = (~\m5_data_i[12]  | ~\new_[16278]_ ) & (~\m6_data_i[12]  | ~\new_[18040]_ );
  assign \new_[10324]_  = (~\m5_data_i[11]  | ~\new_[16277]_ ) & (~\m6_data_i[11]  | ~\new_[19559]_ );
  assign \new_[10325]_  = (~\m7_data_i[10]  | ~\new_[18111]_ ) & (~\m0_data_i[10]  | ~\new_[18027]_ );
  assign \new_[10326]_  = (~\m5_data_i[10]  | ~\new_[18008]_ ) & (~\m6_data_i[10]  | ~\new_[19559]_ );
  assign \new_[10327]_  = (~\m2_data_i[9]  | ~\new_[17222]_ ) & (~\m1_data_i[9]  | ~\new_[17273]_ );
  assign \new_[10328]_  = (~\m5_data_i[9]  | ~\new_[16278]_ ) & (~\m6_data_i[9]  | ~\new_[19559]_ );
  assign \new_[10329]_  = (~\m4_data_i[9]  | ~\new_[16307]_ ) & (~\m3_data_i[9]  | ~\new_[17249]_ );
  assign \new_[10330]_  = (~\m7_data_i[8]  | ~\new_[18111]_ ) & (~\m0_data_i[8]  | ~\new_[18027]_ );
  assign \new_[10331]_  = (~\m2_data_i[8]  | ~\new_[17222]_ ) & (~\m1_data_i[8]  | ~\new_[18177]_ );
  assign \new_[10332]_  = (~\m4_data_i[8]  | ~\new_[16307]_ ) & (~\m3_data_i[8]  | ~\new_[17249]_ );
  assign \new_[10333]_  = (~\m5_data_i[8]  | ~\new_[16277]_ ) & (~\m6_data_i[8]  | ~\new_[18040]_ );
  assign \new_[10334]_  = ~\new_[28581]_  & (~\new_[15782]_  | ~\new_[22763]_ );
  assign \new_[10335]_  = (~\m7_data_i[7]  | ~\new_[18111]_ ) & (~\m0_data_i[7]  | ~\new_[18027]_ );
  assign \new_[10336]_  = (~\m5_data_i[7]  | ~\new_[18008]_ ) & (~\m6_data_i[7]  | ~\new_[19559]_ );
  assign \new_[10337]_  = (~\m2_data_i[6]  | ~\new_[17222]_ ) & (~\m1_data_i[6]  | ~\new_[17273]_ );
  assign \new_[10338]_  = ~\new_[27893]_  & (~\new_[15785]_  | ~\new_[21553]_ );
  assign \new_[10339]_  = (~\m5_data_i[6]  | ~\new_[18008]_ ) & (~\m6_data_i[6]  | ~\new_[19559]_ );
  assign \new_[10340]_  = ~\new_[18410]_  | ~\new_[13842]_ ;
  assign \new_[10341]_  = ~\new_[28720]_  & (~\new_[15789]_  | ~\new_[24532]_ );
  assign \new_[10342]_  = (~\m2_data_i[5]  | ~\new_[17222]_ ) & (~\m1_data_i[5]  | ~\new_[17273]_ );
  assign \new_[10343]_  = (~\m5_data_i[4]  | ~\new_[16278]_ ) & (~\m6_data_i[4]  | ~\new_[19559]_ );
  assign \new_[10344]_  = ~\new_[28260]_  & (~\new_[15792]_  | ~\new_[21444]_ );
  assign \new_[10345]_  = (~\m2_data_i[3]  | ~\new_[17222]_ ) & (~\m1_data_i[3]  | ~\new_[18177]_ );
  assign \new_[10346]_  = ~\new_[28242]_  | (~\new_[15794]_  & ~\new_[23827]_ );
  assign \new_[10347]_  = ~\new_[27929]_  & (~\new_[15796]_  | ~\new_[19441]_ );
  assign \new_[10348]_  = (~\m7_data_i[2]  | ~\new_[18111]_ ) & (~\m0_data_i[2]  | ~\new_[18027]_ );
  assign \new_[10349]_  = (~\m5_data_i[2]  | ~\new_[18008]_ ) & (~\m6_data_i[2]  | ~\new_[18039]_ );
  assign \new_[10350]_  = (~\m5_data_i[1]  | ~\new_[16278]_ ) & (~\m6_data_i[1]  | ~\new_[19559]_ );
  assign \new_[10351]_  = ~\new_[28920]_  & (~\new_[15797]_  | ~\new_[22836]_ );
  assign \new_[10352]_  = ~\new_[15798]_  | ~\new_[29449]_  | ~\new_[26181]_ ;
  assign \new_[10353]_  = (~\m2_data_i[0]  | ~\new_[17222]_ ) & (~\m1_data_i[0]  | ~\new_[18906]_ );
  assign \new_[10354]_  = ~\new_[29243]_  & (~\new_[15799]_  | ~\new_[24254]_ );
  assign \new_[10355]_  = (~\m7_data_i[0]  | ~\new_[18111]_ ) & (~\m0_data_i[0]  | ~\new_[18027]_ );
  assign \new_[10356]_  = (~\m5_data_i[0]  | ~\new_[16278]_ ) & (~\m6_data_i[0]  | ~\new_[18040]_ );
  assign \new_[10357]_  = (~\new_[19559]_  | ~\m6_addr_i[31] ) & (~\new_[18008]_  | ~\new_[31001]_ );
  assign \new_[10358]_  = ~\new_[27974]_  | (~\new_[15803]_  & ~\new_[23842]_ );
  assign \new_[10359]_  = ~\new_[28983]_  & (~\new_[15804]_  | ~\new_[19437]_ );
  assign \new_[10360]_  = (~\new_[17222]_  | ~\new_[31537]_ ) & (~\new_[18177]_  | ~\m1_addr_i[31] );
  assign \new_[10361]_  = ~\new_[20389]_  | ~\new_[13851]_ ;
  assign \new_[10362]_  = (~\new_[18111]_  | ~\m7_addr_i[31] ) & (~\new_[18027]_  | ~\m0_addr_i[31] );
  assign \new_[10363]_  = (~\new_[17222]_  | ~\new_[31486]_ ) & (~\new_[18177]_  | ~\new_[31308]_ );
  assign \new_[10364]_  = ~\new_[15806]_  | ~\new_[28569]_  | ~\new_[24217]_ ;
  assign \new_[10365]_  = (~\new_[17222]_  | ~\m2_addr_i[29] ) & (~\new_[18177]_  | ~\new_[31538]_ );
  assign \new_[10366]_  = (~\new_[19559]_  | ~\m6_addr_i[29] ) & (~\new_[16277]_  | ~\new_[31407]_ );
  assign \new_[10367]_  = (~\new_[18111]_  | ~\new_[30577]_ ) & (~\new_[18027]_  | ~\new_[30957]_ );
  assign \new_[10368]_  = (~\m7_data_i[4]  | ~\new_[17232]_ ) & (~\m0_data_i[4]  | ~\new_[18941]_ );
  assign \new_[10369]_  = (~\new_[17222]_  | ~\new_[31547]_ ) & (~\new_[18177]_  | ~\new_[31458]_ );
  assign \new_[10370]_  = ~\new_[26465]_  | (~\new_[14523]_  & ~\new_[23798]_ );
  assign \new_[10371]_  = (~\new_[17222]_  | ~\m2_addr_i[27] ) & (~\new_[18177]_  | ~\m1_addr_i[27] );
  assign \new_[10372]_  = (~\new_[19559]_  | ~\m6_addr_i[26] ) & (~\new_[16277]_  | ~\m5_addr_i[26] );
  assign \new_[10373]_  = (~\new_[17222]_  | ~\m2_addr_i[25] ) & (~\new_[18177]_  | ~\m1_addr_i[25] );
  assign \new_[10374]_  = (~\m7_data_i[30]  | ~\new_[17240]_ ) & (~\m6_data_i[30]  | ~\new_[18819]_ );
  assign \new_[10375]_  = (~\new_[19559]_  | ~\m6_addr_i[25] ) & (~\new_[16277]_  | ~\m5_addr_i[25] );
  assign \new_[10376]_  = (~\new_[19559]_  | ~\m6_addr_i[24] ) & (~\new_[16277]_  | ~\m5_addr_i[24] );
  assign \new_[10377]_  = ~\new_[27372]_  & (~\new_[15741]_  | ~\new_[21536]_ );
  assign \new_[10378]_  = (~\m2_addr_i[23]  | ~\new_[17222]_ ) & (~\m1_addr_i[23]  | ~\new_[18177]_ );
  assign \new_[10379]_  = ~\new_[27866]_  & (~\new_[15743]_  | ~\new_[22858]_ );
  assign \new_[10380]_  = (~\m5_addr_i[23]  | ~\new_[18008]_ ) & (~\m6_addr_i[23]  | ~\new_[19559]_ );
  assign \new_[10381]_  = (~\m4_addr_i[23]  | ~\new_[16308]_ ) & (~\m3_addr_i[23]  | ~\new_[17249]_ );
  assign \new_[10382]_  = (~\m5_data_i[13]  | ~\new_[20544]_ ) & (~\m6_data_i[13]  | ~\new_[17213]_ );
  assign \new_[10383]_  = (~\m5_addr_i[22]  | ~\new_[16276]_ ) & (~\m6_addr_i[22]  | ~\new_[18036]_ );
  assign \new_[10384]_  = (~\m7_addr_i[22]  | ~\new_[18111]_ ) & (~\m0_addr_i[22]  | ~\new_[18027]_ );
  assign \new_[10385]_  = (~\m7_addr_i[21]  | ~\new_[18111]_ ) & (~\m0_addr_i[21]  | ~\new_[18027]_ );
  assign \new_[10386]_  = (~\m2_addr_i[21]  | ~\new_[17222]_ ) & (~\m1_addr_i[21]  | ~\new_[17273]_ );
  assign \new_[10387]_  = (~\m5_addr_i[21]  | ~\new_[16277]_ ) & (~\m6_addr_i[21]  | ~\new_[18035]_ );
  assign \new_[10388]_  = (~\m7_data_i[29]  | ~\new_[17239]_ ) & (~\m6_data_i[29]  | ~\new_[18090]_ );
  assign \new_[10389]_  = (~\m5_addr_i[20]  | ~\new_[16276]_ ) & (~\m6_addr_i[20]  | ~\new_[18036]_ );
  assign \new_[10390]_  = (~\m7_addr_i[20]  | ~\new_[18111]_ ) & (~\m0_addr_i[20]  | ~\new_[18027]_ );
  assign \new_[10391]_  = (~\m2_addr_i[19]  | ~\new_[17222]_ ) & (~\m1_addr_i[19]  | ~\new_[18177]_ );
  assign \new_[10392]_  = \new_[13854]_  & \new_[28418]_ ;
  assign \new_[10393]_  = (~\m5_addr_i[19]  | ~\new_[16276]_ ) & (~\m6_addr_i[19]  | ~\new_[18036]_ );
  assign \new_[10394]_  = ~\new_[28814]_  & (~\new_[14563]_  | ~\new_[28115]_ );
  assign \new_[10395]_  = \new_[13860]_  & \new_[26766]_ ;
  assign \new_[10396]_  = (~\m5_addr_i[18]  | ~\new_[16277]_ ) & (~\m6_addr_i[18]  | ~\new_[18035]_ );
  assign \new_[10397]_  = (~\m1_data_i[28]  | ~\new_[17277]_ ) & (~\m0_data_i[28]  | ~\new_[16279]_ );
  assign \new_[10398]_  = \new_[13868]_  & \new_[28630]_ ;
  assign \new_[10399]_  = (~\m5_addr_i[17]  | ~\new_[16277]_ ) & (~\m6_addr_i[17]  | ~\new_[18036]_ );
  assign \new_[10400]_  = ~\new_[29057]_  & (~\new_[14565]_  | ~\new_[28481]_ );
  assign \new_[10401]_  = (~\m7_addr_i[17]  | ~\new_[18111]_ ) & (~\m0_addr_i[17]  | ~\new_[18027]_ );
  assign \new_[10402]_  = \new_[13877]_  & \new_[28126]_ ;
  assign \new_[10403]_  = (~\m5_addr_i[16]  | ~\new_[16277]_ ) & (~\m6_addr_i[16]  | ~\new_[18036]_ );
  assign \new_[10404]_  = ~\new_[13805]_  & (~\new_[29058]_  | ~\new_[5898]_ );
  assign \new_[10405]_  = (~\m7_addr_i[16]  | ~\new_[18111]_ ) & (~\m0_addr_i[16]  | ~\new_[18027]_ );
  assign \new_[10406]_  = \new_[13888]_  & \new_[29273]_ ;
  assign \new_[10407]_  = ~\new_[13810]_  & (~\new_[30130]_  | ~\new_[31429]_ );
  assign \new_[10408]_  = (~\m5_addr_i[15]  | ~\new_[16276]_ ) & (~\m6_addr_i[15]  | ~\new_[18035]_ );
  assign \new_[10409]_  = (~\m2_addr_i[14]  | ~\new_[17222]_ ) & (~\m1_addr_i[14]  | ~\new_[18177]_ );
  assign \new_[10410]_  = \new_[13905]_  & \new_[29237]_ ;
  assign \new_[10411]_  = (~\m5_addr_i[14]  | ~\new_[16277]_ ) & (~\m6_addr_i[14]  | ~\new_[18035]_ );
  assign \new_[10412]_  = \new_[13913]_  & \new_[29678]_ ;
  assign \new_[10413]_  = (~\m5_addr_i[22]  | ~\new_[20544]_ ) & (~\m6_addr_i[22]  | ~\new_[17213]_ );
  assign \new_[10414]_  = ~\new_[13821]_  & (~\new_[29254]_  | ~\new_[5902]_ );
  assign \new_[10415]_  = (~\m5_addr_i[13]  | ~\new_[16276]_ ) & (~\m6_addr_i[13]  | ~\new_[18036]_ );
  assign \new_[10416]_  = ~\new_[26723]_  & (~\new_[14569]_  | ~\new_[28556]_ );
  assign \new_[10417]_  = \new_[13921]_  & \new_[29279]_ ;
  assign \new_[10418]_  = ~\new_[13825]_  & (~\new_[29115]_  | ~\new_[5903]_ );
  assign \new_[10419]_  = (~\m5_addr_i[12]  | ~\new_[16276]_ ) & (~\m6_addr_i[12]  | ~\new_[18035]_ );
  assign \new_[10420]_  = (~\m1_data_i[26]  | ~\new_[17277]_ ) & (~\m0_data_i[26]  | ~\new_[16279]_ );
  assign \new_[10421]_  = (~\m5_addr_i[11]  | ~\new_[16276]_ ) & (~\m6_addr_i[11]  | ~\new_[18036]_ );
  assign \new_[10422]_  = (~\m7_data_i[26]  | ~\new_[17239]_ ) & (~\m6_data_i[26]  | ~\new_[19581]_ );
  assign \new_[10423]_  = (~\m4_addr_i[11]  | ~\new_[16307]_ ) & (~\m3_addr_i[11]  | ~\new_[17249]_ );
  assign \new_[10424]_  = (~\m2_addr_i[11]  | ~\new_[17222]_ ) & (~\m1_addr_i[11]  | ~\new_[17273]_ );
  assign \new_[10425]_  = ~\new_[13832]_  & (~\new_[29229]_  | ~\new_[5905]_ );
  assign \new_[10426]_  = ~\new_[29200]_  & (~\new_[14573]_  | ~\new_[28573]_ );
  assign \new_[10427]_  = \new_[13945]_  & \new_[29041]_ ;
  assign \new_[10428]_  = (~\m5_addr_i[10]  | ~\new_[16277]_ ) & (~\m6_addr_i[10]  | ~\new_[18036]_ );
  assign \new_[10429]_  = \new_[13949]_  & \new_[29144]_ ;
  assign \new_[10430]_  = (~\m5_addr_i[9]  | ~\new_[18008]_ ) & (~\m6_addr_i[9]  | ~\new_[18035]_ );
  assign \new_[10431]_  = \new_[13954]_  & \new_[26639]_ ;
  assign \new_[10432]_  = (~\m2_addr_i[9]  | ~\new_[17222]_ ) & (~\m1_addr_i[9]  | ~\new_[17273]_ );
  assign \new_[10433]_  = (~\m5_addr_i[8]  | ~\new_[18008]_ ) & (~\m6_addr_i[8]  | ~\new_[18036]_ );
  assign \new_[10434]_  = (~\m4_addr_i[8]  | ~\new_[16308]_ ) & (~\m3_addr_i[8]  | ~\new_[17249]_ );
  assign \new_[10435]_  = \new_[13967]_  & \new_[28077]_ ;
  assign \new_[10436]_  = (~\m5_addr_i[7]  | ~\new_[16277]_ ) & (~\m6_addr_i[7]  | ~\new_[18035]_ );
  assign \new_[10437]_  = \new_[13975]_  & \new_[27000]_ ;
  assign \new_[10438]_  = (~\m5_addr_i[6]  | ~\new_[18008]_ ) & (~\m6_addr_i[6]  | ~\new_[18036]_ );
  assign \new_[10439]_  = (~\m7_data_i[24]  | ~\new_[17239]_ ) & (~\m6_data_i[24]  | ~\new_[18819]_ );
  assign \new_[10440]_  = ~\new_[28022]_  & (~\new_[15745]_  | ~\new_[24241]_ );
  assign \new_[10441]_  = ~\new_[27840]_  & (~\new_[15746]_  | ~\new_[27402]_ );
  assign \new_[10442]_  = (~\m7_addr_i[6]  | ~\new_[18111]_ ) & (~\m0_addr_i[6]  | ~\new_[18027]_ );
  assign \new_[10443]_  = (~\m5_addr_i[5]  | ~\new_[18008]_ ) & (~\m6_addr_i[5]  | ~\new_[18036]_ );
  assign \new_[10444]_  = (~\m7_addr_i[5]  | ~\new_[18111]_ ) & (~\m0_addr_i[5]  | ~\new_[18027]_ );
  assign \new_[10445]_  = (~\new_[31095]_  | ~\new_[17222]_ ) & (~\m1_addr_i[5]  | ~\new_[18177]_ );
  assign \new_[10446]_  = ~\new_[16640]_  | ~\new_[17530]_  | ~\new_[17529]_  | ~\new_[18466]_ ;
  assign \new_[10447]_  = (~\m2_addr_i[4]  | ~\new_[17222]_ ) & (~\m1_addr_i[4]  | ~\new_[18906]_ );
  assign \new_[10448]_  = (~\m4_addr_i[4]  | ~\new_[16307]_ ) & (~\m3_addr_i[4]  | ~\new_[17249]_ );
  assign \new_[10449]_  = (~\m5_addr_i[4]  | ~\new_[18008]_ ) & (~\m6_addr_i[4]  | ~\new_[18039]_ );
  assign \new_[10450]_  = (~\m4_addr_i[3]  | ~\new_[16307]_ ) & (~\m3_addr_i[3]  | ~\new_[17249]_ );
  assign \new_[10451]_  = ~\new_[17535]_  | ~\new_[16644]_  | ~\new_[17533]_  | ~\new_[17534]_ ;
  assign \new_[10452]_  = (~\m5_addr_i[3]  | ~\new_[16278]_ ) & (~\m6_addr_i[3]  | ~\new_[18039]_ );
  assign \new_[10453]_  = (~\m2_addr_i[2]  | ~\new_[17222]_ ) & (~\new_[31477]_  | ~\new_[18177]_ );
  assign \new_[10454]_  = (~\m7_addr_i[2]  | ~\new_[18111]_ ) & (~\m0_addr_i[2]  | ~\new_[18027]_ );
  assign \new_[10455]_  = (~\m5_addr_i[2]  | ~\new_[16277]_ ) & (~\m6_addr_i[2]  | ~\new_[19559]_ );
  assign \new_[10456]_  = (~\m2_addr_i[1]  | ~\new_[17222]_ ) & (~\m1_addr_i[1]  | ~\new_[17273]_ );
  assign \new_[10457]_  = ~\new_[16654]_  | ~\new_[16655]_  | ~\new_[17537]_  | ~\new_[16653]_ ;
  assign \new_[10458]_  = (~\m7_addr_i[0]  | ~\new_[18111]_ ) & (~\m0_addr_i[0]  | ~\new_[18027]_ );
  assign \new_[10459]_  = (~\m2_addr_i[0]  | ~\new_[17222]_ ) & (~\m1_addr_i[0]  | ~\new_[18906]_ );
  assign \new_[10460]_  = (~\m5_sel_i[3]  | ~\new_[16276]_ ) & (~\m6_sel_i[3]  | ~\new_[19559]_ );
  assign \new_[10461]_  = (~\m7_sel_i[3]  | ~\new_[18111]_ ) & (~\m0_sel_i[3]  | ~\new_[18027]_ );
  assign \new_[10462]_  = (~\m2_sel_i[2]  | ~\new_[17222]_ ) & (~\m1_sel_i[2]  | ~\new_[18177]_ );
  assign \new_[10463]_  = ~\new_[17540]_  | ~\new_[16658]_  | ~\new_[16657]_  | ~\new_[17539]_ ;
  assign \new_[10464]_  = ~\new_[16659]_  | ~\new_[18473]_  | ~\new_[18471]_  | ~\new_[18472]_ ;
  assign \new_[10465]_  = (~\m5_sel_i[2]  | ~\new_[16277]_ ) & (~\m6_sel_i[2]  | ~\new_[18038]_ );
  assign \new_[10466]_  = (~\m5_sel_i[1]  | ~\new_[16277]_ ) & (~\m6_sel_i[1]  | ~\new_[18035]_ );
  assign \new_[10467]_  = (~\m5_data_i[21]  | ~\new_[17203]_ ) & (~\m4_data_i[21]  | ~\new_[17271]_ );
  assign \new_[10468]_  = (~\m7_sel_i[0]  | ~\new_[18111]_ ) & (~\m0_sel_i[0]  | ~\new_[18027]_ );
  assign \new_[10469]_  = ~\new_[28642]_  & (~\new_[14579]_  | ~\new_[24160]_ );
  assign \new_[10470]_  = (~m2_we_i | ~\new_[17222]_ ) & (~m1_we_i | ~\new_[18906]_ );
  assign \new_[10471]_  = (~m5_we_i | ~\new_[16277]_ ) & (~m6_we_i | ~\new_[18039]_ );
  assign \new_[10472]_  = (~\m5_data_i[19]  | ~\new_[17203]_ ) & (~\m4_data_i[19]  | ~\new_[17271]_ );
  assign \new_[10473]_  = (~\m7_data_i[19]  | ~\new_[17239]_ ) & (~\m6_data_i[19]  | ~\new_[18819]_ );
  assign \new_[10474]_  = (~\m7_data_i[18]  | ~\new_[17239]_ ) & (~\m6_data_i[18]  | ~\new_[18819]_ );
  assign \new_[10475]_  = ~\new_[17555]_  | ~\new_[16680]_  | ~\new_[16678]_  | ~\new_[16679]_ ;
  assign \new_[10476]_  = ~\new_[16684]_  | ~\new_[16683]_  | ~\new_[17556]_  | ~\new_[15910]_ ;
  assign \new_[10477]_  = ~\new_[26633]_  & (~\new_[14581]_  | ~\new_[24214]_ );
  assign \new_[10478]_  = (~\m7_data_i[17]  | ~\new_[17239]_ ) & (~\m6_data_i[17]  | ~\new_[18819]_ );
  assign \new_[10479]_  = ~\new_[17564]_  | ~\new_[17558]_  | ~\new_[16689]_  | ~\new_[14504]_ ;
  assign \new_[10480]_  = (~\m7_data_i[16]  | ~\new_[17240]_ ) & (~\m6_data_i[16]  | ~\new_[18819]_ );
  assign \new_[10481]_  = ~\new_[15904]_  | ~\new_[15905]_  | ~\new_[14514]_  | ~\new_[14515]_ ;
  assign \new_[10482]_  = (~\m7_sel_i[3]  | ~\new_[16296]_ ) & (~\m0_sel_i[3]  | ~\new_[18763]_ );
  assign \new_[10483]_  = (~\m5_data_i[15]  | ~\new_[18745]_ ) & (~\m4_data_i[15]  | ~\new_[17271]_ );
  assign \new_[10484]_  = (~\m5_data_i[14]  | ~\new_[18745]_ ) & (~\m4_data_i[14]  | ~\new_[17271]_ );
  assign \new_[10485]_  = (~\m1_data_i[14]  | ~\new_[17277]_ ) & (~\m0_data_i[14]  | ~\new_[16279]_ );
  assign \new_[10486]_  = (~\m7_data_i[14]  | ~\new_[17239]_ ) & (~\m6_data_i[14]  | ~\new_[18089]_ );
  assign \new_[10487]_  = ~\new_[15908]_  | ~\new_[16700]_  | ~\new_[17562]_  | ~\new_[17563]_ ;
  assign \new_[10488]_  = (~\m5_data_i[13]  | ~\new_[18745]_ ) & (~\m4_data_i[13]  | ~\new_[17271]_ );
  assign \new_[10489]_  = (~\m7_data_i[13]  | ~\new_[17239]_ ) & (~\m6_data_i[13]  | ~\new_[18090]_ );
  assign \new_[10490]_  = (~\m1_data_i[13]  | ~\new_[17277]_ ) & (~\m0_data_i[13]  | ~\new_[14834]_ );
  assign \new_[10491]_  = ~\new_[28179]_  & (~\new_[15717]_  | ~\new_[24189]_ );
  assign \new_[10492]_  = ~\new_[28716]_  & (~\new_[15721]_  | ~\new_[21347]_ );
  assign \new_[10493]_  = (~\m1_data_i[12]  | ~\new_[17277]_ ) & (~\m0_data_i[12]  | ~\new_[14834]_ );
  assign \new_[10494]_  = ~\new_[29679]_  & (~\new_[15726]_  | ~\new_[21355]_ );
  assign \new_[10495]_  = (~\m5_data_i[11]  | ~\new_[18745]_ ) & (~\m4_data_i[11]  | ~\new_[17271]_ );
  assign \new_[10496]_  = (~\m1_data_i[11]  | ~\new_[17277]_ ) & (~\m0_data_i[11]  | ~\new_[16279]_ );
  assign \new_[10497]_  = ~\new_[28056]_  & (~\new_[15736]_  | ~\new_[26174]_ );
  assign \new_[10498]_  = ~\new_[13996]_  & (~\new_[30206]_  | ~\new_[5973]_ );
  assign \new_[10499]_  = (~\m7_data_i[11]  | ~\new_[17239]_ ) & (~\m6_data_i[11]  | ~\new_[18089]_ );
  assign \new_[10500]_  = ~\new_[28255]_  & (~\new_[15740]_  | ~\new_[22808]_ );
  assign \new_[10501]_  = ~\new_[14003]_  & (~\new_[29169]_  | ~\new_[31235]_ );
  assign \new_[10502]_  = (~\m5_data_i[10]  | ~\new_[17203]_ ) & (~\m4_data_i[10]  | ~\new_[17271]_ );
  assign \new_[10503]_  = ~\new_[28159]_  & (~\new_[15751]_  | ~\new_[22806]_ );
  assign \new_[10504]_  = ~\new_[28088]_  & (~\new_[15753]_  | ~\new_[22592]_ );
  assign \new_[10505]_  = (~\m1_data_i[10]  | ~\new_[18192]_ ) & (~\m0_data_i[10]  | ~\new_[14834]_ );
  assign \new_[10506]_  = (~\m7_data_i[10]  | ~\new_[17239]_ ) & (~\m6_data_i[10]  | ~\new_[19581]_ );
  assign \new_[10507]_  = ~\new_[28267]_  & (~\new_[15757]_  | ~\new_[22825]_ );
  assign \new_[10508]_  = (~\m7_data_i[9]  | ~\new_[17239]_ ) & (~\m6_data_i[9]  | ~\new_[17227]_ );
  assign \new_[10509]_  = ~\new_[29274]_  & (~\new_[15763]_  | ~\new_[22654]_ );
  assign \new_[10510]_  = ~\new_[14032]_  & (~\new_[29300]_  | ~\new_[5988]_ );
  assign \new_[10511]_  = ~\new_[28312]_  & (~\new_[15766]_  | ~\new_[24197]_ );
  assign \new_[10512]_  = ~\new_[28557]_  & (~\new_[15774]_  | ~\new_[21357]_ );
  assign \new_[10513]_  = (~\m7_data_i[8]  | ~\new_[17239]_ ) & (~\m6_data_i[8]  | ~\new_[17227]_ );
  assign \new_[10514]_  = (~\m7_data_i[25]  | ~\new_[16296]_ ) & (~\m0_data_i[25]  | ~\new_[20545]_ );
  assign \new_[10515]_  = ~\new_[28667]_  & (~\new_[15777]_  | ~\new_[24230]_ );
  assign \new_[10516]_  = (~\m1_data_i[7]  | ~\new_[17277]_ ) & (~\m0_data_i[7]  | ~\new_[16279]_ );
  assign \new_[10517]_  = ~\new_[25457]_  & (~\new_[15780]_  | ~\new_[22658]_ );
  assign \new_[10518]_  = ~\new_[28141]_  & (~\new_[15783]_  | ~\new_[24155]_ );
  assign \new_[10519]_  = (~\m7_data_i[7]  | ~\new_[17239]_ ) & (~\m6_data_i[7]  | ~\new_[17227]_ );
  assign \new_[10520]_  = ~\new_[28145]_  & (~\new_[15793]_  | ~\new_[20434]_ );
  assign \new_[10521]_  = ~\new_[14061]_  & (~\new_[30078]_  | ~\new_[6003]_ );
  assign \new_[10522]_  = ~\new_[28929]_  & (~\new_[15800]_  | ~\new_[22761]_ );
  assign \new_[10523]_  = (~\m1_data_i[6]  | ~\new_[17277]_ ) & (~\m0_data_i[6]  | ~\new_[16279]_ );
  assign \new_[10524]_  = (~\m7_data_i[6]  | ~\new_[17239]_ ) & (~\m6_data_i[6]  | ~\new_[18089]_ );
  assign \new_[10525]_  = ~\new_[14071]_  & (~\new_[30072]_  | ~\new_[6006]_ );
  assign \new_[10526]_  = ~\new_[28205]_  & (~\new_[15809]_  | ~\new_[26240]_ );
  assign \new_[10527]_  = (~\m7_data_i[5]  | ~\new_[17239]_ ) & (~\m6_data_i[5]  | ~\new_[17227]_ );
  assign \new_[10528]_  = ~\new_[23859]_  & (~\new_[14774]_  | ~\new_[30432]_ );
  assign \new_[10529]_  = ~\new_[22340]_  & (~\new_[14799]_  | ~\new_[29355]_ );
  assign \new_[10530]_  = ~\new_[22254]_  & (~\new_[14794]_  | ~\new_[30210]_ );
  assign \new_[10531]_  = ~\new_[20348]_  & (~\new_[14803]_  | ~\new_[29701]_ );
  assign \new_[10532]_  = (~\m1_data_i[3]  | ~\new_[17277]_ ) & (~\m0_data_i[3]  | ~\new_[14834]_ );
  assign \new_[10533]_  = (~\m5_data_i[2]  | ~\new_[18745]_ ) & (~\m4_data_i[2]  | ~\new_[17271]_ );
  assign \new_[10534]_  = (~\m7_data_i[2]  | ~\new_[17239]_ ) & (~\m6_data_i[2]  | ~\new_[18090]_ );
  assign \new_[10535]_  = ~\new_[14438]_  & ~\new_[14611]_ ;
  assign \new_[10536]_  = ~\new_[14439]_  & ~\new_[14618]_ ;
  assign \new_[10537]_  = (~\m7_data_i[1]  | ~\new_[17239]_ ) & (~\m6_data_i[1]  | ~\new_[18089]_ );
  assign \new_[10538]_  = (~\m1_data_i[0]  | ~\new_[18192]_ ) & (~\m0_data_i[0]  | ~\new_[14834]_ );
  assign \new_[10539]_  = (~\new_[17271]_  | ~\m4_addr_i[30] ) & (~\new_[32350]_  | ~\m3_addr_i[30] );
  assign \new_[10540]_  = (~\new_[17239]_  | ~\new_[31531]_ ) & (~\new_[16279]_  | ~\new_[31481]_ );
  assign \new_[10541]_  = ~\new_[14442]_  & ~\new_[14685]_ ;
  assign \new_[10542]_  = ~\new_[14441]_  & ~\new_[14691]_ ;
  assign \new_[10543]_  = ~\new_[28964]_  | ~\new_[14489]_  | ~\new_[30105]_ ;
  assign \new_[10544]_  = ~\new_[14443]_  & ~\new_[13283]_ ;
  assign \new_[10545]_  = (~\new_[17240]_  | ~\m7_addr_i[25] ) & (~\new_[14834]_  | ~\m0_addr_i[25] );
  assign \new_[10546]_  = (~\m7_data_i[31]  | ~\new_[17232]_ ) & (~\m0_data_i[31]  | ~\new_[18941]_ );
  assign \new_[10547]_  = (~\m7_data_i[22]  | ~\new_[16296]_ ) & (~\m0_data_i[22]  | ~\new_[18764]_ );
  assign \new_[10548]_  = (~\new_[17239]_  | ~\m7_addr_i[24] ) & (~\new_[14834]_  | ~\m0_addr_i[24] );
  assign \new_[10549]_  = ~\new_[14595]_  | ~\new_[14461]_  | ~\new_[14587]_ ;
  assign \new_[10550]_  = (~\m7_addr_i[23]  | ~\new_[17239]_ ) & (~\m6_addr_i[23]  | ~\new_[18819]_ );
  assign \new_[10551]_  = (~\m7_data_i[27]  | ~\new_[17232]_ ) & (~\m0_data_i[27]  | ~\new_[18941]_ );
  assign \new_[10552]_  = (~\m5_data_i[20]  | ~\new_[18004]_ ) & (~\m6_data_i[20]  | ~\new_[17241]_ );
  assign \new_[10553]_  = (~\m7_data_i[25]  | ~\new_[17232]_ ) & (~\m0_data_i[25]  | ~\new_[18941]_ );
  assign \new_[10554]_  = (~\m2_addr_i[23]  | ~\new_[17193]_ ) & (~\m1_addr_i[23]  | ~\new_[19633]_ );
  assign \new_[10555]_  = ~\new_[14374]_  & ~\new_[22276]_ ;
  assign \new_[10556]_  = (~\m7_data_i[23]  | ~\new_[17232]_ ) & (~\m0_data_i[23]  | ~\new_[18941]_ );
  assign \new_[10557]_  = (~\m7_data_i[3]  | ~\new_[16296]_ ) & (~\m0_data_i[3]  | ~\new_[18764]_ );
  assign \new_[10558]_  = (~\m7_data_i[22]  | ~\new_[17232]_ ) & (~\m0_data_i[22]  | ~\new_[19648]_ );
  assign \new_[10559]_  = (~\m7_data_i[21]  | ~\new_[17232]_ ) & (~\m0_data_i[21]  | ~\new_[20580]_ );
  assign \new_[10560]_  = (~\m7_data_i[20]  | ~\new_[17232]_ ) & (~\m0_data_i[20]  | ~\new_[19648]_ );
  assign \new_[10561]_  = (~\m7_data_i[19]  | ~\new_[17232]_ ) & (~\m0_data_i[19]  | ~\new_[19648]_ );
  assign \new_[10562]_  = (~\m1_addr_i[20]  | ~\new_[17277]_ ) & (~\m0_addr_i[20]  | ~\new_[16279]_ );
  assign \new_[10563]_  = (~\m7_data_i[17]  | ~\new_[17232]_ ) & (~\m0_data_i[17]  | ~\new_[19648]_ );
  assign \new_[10564]_  = (~\m5_data_i[17]  | ~\new_[18016]_ ) & (~\m6_data_i[17]  | ~\new_[17229]_ );
  assign \new_[10565]_  = (~\m7_data_i[16]  | ~\new_[17232]_ ) & (~\m0_data_i[16]  | ~\new_[18941]_ );
  assign \new_[10566]_  = (~\m7_addr_i[19]  | ~\new_[17240]_ ) & (~\m6_addr_i[19]  | ~\new_[18819]_ );
  assign \new_[10567]_  = (~\m1_addr_i[19]  | ~\new_[17277]_ ) & (~\m0_addr_i[19]  | ~\new_[16279]_ );
  assign \new_[10568]_  = (~\m5_data_i[15]  | ~\new_[18016]_ ) & (~\m6_data_i[15]  | ~\new_[17229]_ );
  assign \new_[10569]_  = (~\m5_data_i[14]  | ~\new_[18016]_ ) & (~\m6_data_i[14]  | ~\new_[17229]_ );
  assign \new_[10570]_  = (~\m7_data_i[14]  | ~\new_[17232]_ ) & (~\m0_data_i[14]  | ~\new_[18941]_ );
  assign \new_[10571]_  = (~\m7_data_i[13]  | ~\new_[17232]_ ) & (~\m0_data_i[13]  | ~\new_[18941]_ );
  assign \new_[10572]_  = (~\m7_data_i[12]  | ~\new_[17232]_ ) & (~\m0_data_i[12]  | ~\new_[18941]_ );
  assign \new_[10573]_  = (~\m7_data_i[11]  | ~\new_[17232]_ ) & (~\m0_data_i[11]  | ~\new_[18941]_ );
  assign \new_[10574]_  = (~\m7_addr_i[17]  | ~\new_[17240]_ ) & (~\m6_addr_i[17]  | ~\new_[18819]_ );
  assign \new_[10575]_  = (~\m5_data_i[9]  | ~\new_[18016]_ ) & (~\m6_data_i[9]  | ~\new_[17229]_ );
  assign \new_[10576]_  = (~\m7_data_i[9]  | ~\new_[17232]_ ) & (~\m0_data_i[9]  | ~\new_[18941]_ );
  assign \new_[10577]_  = (~\m7_data_i[7]  | ~\new_[17232]_ ) & (~\m0_data_i[7]  | ~\new_[18941]_ );
  assign \new_[10578]_  = (~\m7_addr_i[16]  | ~\new_[17240]_ ) & (~\m6_addr_i[16]  | ~\new_[18819]_ );
  assign \new_[10579]_  = (~\m5_data_i[6]  | ~\new_[18016]_ ) & (~\m6_data_i[6]  | ~\new_[17229]_ );
  assign \new_[10580]_  = (~\m5_data_i[5]  | ~\new_[18016]_ ) & (~\m6_data_i[5]  | ~\new_[17229]_ );
  assign \new_[10581]_  = (~\m5_data_i[4]  | ~\new_[18015]_ ) & (~\m6_data_i[4]  | ~\new_[17229]_ );
  assign \new_[10582]_  = (~\m5_data_i[3]  | ~\new_[18015]_ ) & (~\m6_data_i[3]  | ~\new_[17229]_ );
  assign \new_[10583]_  = (~\m7_addr_i[15]  | ~\new_[17239]_ ) & (~\m6_addr_i[15]  | ~\new_[19581]_ );
  assign \new_[10584]_  = (~\m7_data_i[3]  | ~\new_[17232]_ ) & (~\m0_data_i[3]  | ~\new_[19648]_ );
  assign \new_[10585]_  = (~\m5_data_i[2]  | ~\new_[18016]_ ) & (~\m6_data_i[2]  | ~\new_[17229]_ );
  assign \new_[10586]_  = (~\m7_data_i[1]  | ~\new_[17232]_ ) & (~\m0_data_i[1]  | ~\new_[18941]_ );
  assign \new_[10587]_  = (~\m7_data_i[0]  | ~\new_[17232]_ ) & (~\m0_data_i[0]  | ~\new_[19648]_ );
  assign \new_[10588]_  = (~\m1_addr_i[14]  | ~\new_[17277]_ ) & (~\m0_addr_i[14]  | ~\new_[16279]_ );
  assign \new_[10589]_  = (~\new_[17232]_  | ~\new_[31885]_ ) & (~\new_[18941]_  | ~\new_[31292]_ );
  assign \new_[10590]_  = (~\new_[17229]_  | ~\m6_addr_i[29] ) & (~\new_[18014]_  | ~\new_[31407]_ );
  assign \new_[10591]_  = (~\m1_addr_i[11]  | ~\new_[17277]_ ) & (~\m0_addr_i[11]  | ~\new_[16279]_ );
  assign \new_[10592]_  = (~\m7_addr_i[22]  | ~\new_[17232]_ ) & (~\m0_addr_i[22]  | ~\new_[18941]_ );
  assign \new_[10593]_  = (~\m7_addr_i[20]  | ~\new_[16296]_ ) & (~\m0_addr_i[20]  | ~\new_[18764]_ );
  assign \new_[10594]_  = (~\m5_addr_i[22]  | ~\new_[18016]_ ) & (~\m6_addr_i[22]  | ~\new_[17229]_ );
  assign \new_[10595]_  = (~\m5_data_i[6]  | ~\new_[17203]_ ) & (~\m4_data_i[6]  | ~\new_[17271]_ );
  assign \new_[10596]_  = ~\new_[12424]_ ;
  assign \new_[10597]_  = (~\m7_addr_i[19]  | ~\new_[17232]_ ) & (~\m0_addr_i[19]  | ~\new_[18941]_ );
  assign \new_[10598]_  = (~\m7_addr_i[18]  | ~\new_[17232]_ ) & (~\m0_addr_i[18]  | ~\new_[20580]_ );
  assign \new_[10599]_  = (~\m7_addr_i[17]  | ~\new_[17232]_ ) & (~\m0_addr_i[17]  | ~\new_[20580]_ );
  assign \new_[10600]_  = (~\m1_addr_i[9]  | ~\new_[17277]_ ) & (~\m0_addr_i[9]  | ~\new_[14834]_ );
  assign \new_[10601]_  = (~\m7_addr_i[16]  | ~\new_[17232]_ ) & (~\m0_addr_i[16]  | ~\new_[19648]_ );
  assign \new_[10602]_  = (~\m1_addr_i[8]  | ~\new_[18192]_ ) & (~\m0_addr_i[8]  | ~\new_[14834]_ );
  assign \new_[10603]_  = (~\m7_addr_i[8]  | ~\new_[17239]_ ) & (~\m6_addr_i[8]  | ~\new_[18089]_ );
  assign \new_[10604]_  = (~\m7_addr_i[12]  | ~\new_[17232]_ ) & (~\m0_addr_i[12]  | ~\new_[18941]_ );
  assign \new_[10605]_  = (~\m5_addr_i[12]  | ~\new_[18016]_ ) & (~\m6_addr_i[12]  | ~\new_[17229]_ );
  assign \new_[10606]_  = (~\m7_addr_i[7]  | ~\new_[17239]_ ) & (~\m6_addr_i[7]  | ~\new_[19581]_ );
  assign \new_[10607]_  = (~\m5_addr_i[10]  | ~\new_[18016]_ ) & (~\m6_addr_i[10]  | ~\new_[17229]_ );
  assign \new_[10608]_  = (~\m5_addr_i[12]  | ~\new_[18751]_ ) & (~\m6_addr_i[12]  | ~\new_[17213]_ );
  assign \new_[10609]_  = ~\new_[14444]_  | ~\new_[22892]_ ;
  assign \new_[10610]_  = ~\new_[14445]_  | ~\new_[23022]_ ;
  assign \new_[10611]_  = ~\new_[14437]_  & (~\new_[29909]_  | ~\new_[5910]_ );
  assign \new_[10612]_  = (~\m7_addr_i[8]  | ~\new_[17232]_ ) & (~\m0_addr_i[8]  | ~\new_[18941]_ );
  assign \new_[10613]_  = (~\m5_addr_i[7]  | ~\new_[18016]_ ) & (~\m6_addr_i[7]  | ~\new_[17229]_ );
  assign \new_[10614]_  = (~\m7_addr_i[6]  | ~\new_[17239]_ ) & (~\m6_addr_i[6]  | ~\new_[19581]_ );
  assign \new_[10615]_  = (~\m5_addr_i[5]  | ~\new_[18015]_ ) & (~\m6_addr_i[5]  | ~\new_[17229]_ );
  assign \new_[10616]_  = (~\m5_addr_i[5]  | ~\new_[18745]_ ) & (~\m4_addr_i[5]  | ~\new_[17271]_ );
  assign \new_[10617]_  = (~\m7_addr_i[5]  | ~\new_[17239]_ ) & (~\m6_addr_i[5]  | ~\new_[19581]_ );
  assign \new_[10618]_  = (~\m5_addr_i[4]  | ~\new_[18015]_ ) & (~\m6_addr_i[4]  | ~\new_[17229]_ );
  assign \new_[10619]_  = (~\m7_addr_i[3]  | ~\new_[17232]_ ) & (~\new_[31884]_  | ~\new_[19648]_ );
  assign \new_[10620]_  = (~\m5_addr_i[4]  | ~\new_[17203]_ ) & (~\m4_addr_i[4]  | ~\new_[17271]_ );
  assign \new_[10621]_  = (~\m7_addr_i[2]  | ~\new_[17232]_ ) & (~\m0_addr_i[2]  | ~\new_[18941]_ );
  assign \new_[10622]_  = ~\new_[30144]_  & (~\new_[14622]_  | ~\new_[18431]_ );
  assign \new_[10623]_  = (~\m7_addr_i[1]  | ~\new_[17232]_ ) & (~\m0_addr_i[1]  | ~\new_[19648]_ );
  assign \new_[10624]_  = (~\m7_addr_i[0]  | ~\new_[17232]_ ) & (~\m0_addr_i[0]  | ~\new_[20580]_ );
  assign \new_[10625]_  = (~\m5_addr_i[3]  | ~\new_[18745]_ ) & (~\m4_addr_i[3]  | ~\new_[17271]_ );
  assign \new_[10626]_  = (~\m7_sel_i[2]  | ~\new_[17232]_ ) & (~\m0_sel_i[2]  | ~\new_[20580]_ );
  assign \new_[10627]_  = ~\new_[14446]_  | ~\new_[21507]_ ;
  assign \new_[10628]_  = (~\m7_sel_i[1]  | ~\new_[17232]_ ) & (~\m0_sel_i[1]  | ~\new_[18941]_ );
  assign \new_[10629]_  = (~\m1_addr_i[3]  | ~\new_[17277]_ ) & (~\new_[31884]_  | ~\new_[14834]_ );
  assign \new_[10630]_  = ~\new_[27574]_  & (~\new_[14632]_  | ~\new_[29020]_ );
  assign \new_[10631]_  = (~\m7_sel_i[0]  | ~\new_[17232]_ ) & (~\m0_sel_i[0]  | ~\new_[19648]_ );
  assign \new_[10632]_  = (~\m5_addr_i[2]  | ~\new_[18745]_ ) & (~\m4_addr_i[2]  | ~\new_[17271]_ );
  assign \new_[10633]_  = (~\new_[31477]_  | ~\new_[17277]_ ) & (~\m0_addr_i[2]  | ~\new_[14834]_ );
  assign \new_[10634]_  = (~\m1_addr_i[1]  | ~\new_[17277]_ ) & (~\m0_addr_i[1]  | ~\new_[14834]_ );
  assign \new_[10635]_  = (~\m7_data_i[31]  | ~\new_[16296]_ ) & (~\m0_data_i[31]  | ~\new_[18765]_ );
  assign \new_[10636]_  = (~\m7_data_i[30]  | ~\new_[16296]_ ) & (~\m0_data_i[30]  | ~\new_[18766]_ );
  assign \new_[10637]_  = (~\m7_addr_i[0]  | ~\new_[17239]_ ) & (~\m6_addr_i[0]  | ~\new_[18819]_ );
  assign \new_[10638]_  = (~\m5_data_i[29]  | ~\new_[18004]_ ) & (~\m6_data_i[29]  | ~\new_[17241]_ );
  assign \new_[10639]_  = (~\m7_data_i[29]  | ~\new_[16296]_ ) & (~\m0_data_i[29]  | ~\new_[18766]_ );
  assign \new_[10640]_  = (~\m7_data_i[28]  | ~\new_[16296]_ ) & (~\m0_data_i[28]  | ~\new_[18763]_ );
  assign \new_[10641]_  = (~\m5_sel_i[3]  | ~\new_[17203]_ ) & (~\m4_sel_i[3]  | ~\new_[17271]_ );
  assign \new_[10642]_  = (~\m7_sel_i[3]  | ~\new_[17239]_ ) & (~\m6_sel_i[3]  | ~\new_[18819]_ );
  assign \new_[10643]_  = (~\m7_data_i[27]  | ~\new_[16296]_ ) & (~\m0_data_i[27]  | ~\new_[20545]_ );
  assign \new_[10644]_  = (~\m7_data_i[26]  | ~\new_[16296]_ ) & (~\m0_data_i[26]  | ~\new_[20545]_ );
  assign \new_[10645]_  = (~\m7_sel_i[2]  | ~\new_[17240]_ ) & (~\m6_sel_i[2]  | ~\new_[19581]_ );
  assign \new_[10646]_  = (~\m7_data_i[24]  | ~\new_[16296]_ ) & (~\m0_data_i[24]  | ~\new_[20545]_ );
  assign \new_[10647]_  = (~\m5_sel_i[2]  | ~\new_[18745]_ ) & (~\m4_sel_i[2]  | ~\new_[17271]_ );
  assign \new_[10648]_  = (~\m5_data_i[24]  | ~\new_[18004]_ ) & (~\m6_data_i[24]  | ~\new_[17241]_ );
  assign \new_[10649]_  = (~\m5_data_i[23]  | ~\new_[18004]_ ) & (~\m6_data_i[23]  | ~\new_[18836]_ );
  assign \new_[10650]_  = (~\m7_data_i[23]  | ~\new_[16296]_ ) & (~\m0_data_i[23]  | ~\new_[18766]_ );
  assign \new_[10651]_  = (~\m7_data_i[21]  | ~\new_[16296]_ ) & (~\m0_data_i[21]  | ~\new_[18764]_ );
  assign \new_[10652]_  = ~\new_[14449]_  | ~\new_[21508]_ ;
  assign \new_[10653]_  = (~\m5_sel_i[1]  | ~\new_[17203]_ ) & (~\m4_sel_i[1]  | ~\new_[17271]_ );
  assign \new_[10654]_  = ~\new_[28043]_  & (~\new_[14673]_  | ~\new_[18429]_ );
  assign \new_[10655]_  = (~\m1_sel_i[1]  | ~\new_[18192]_ ) & (~\m0_sel_i[1]  | ~\new_[14834]_ );
  assign \new_[10656]_  = (~\m7_data_i[20]  | ~\new_[16296]_ ) & (~\m0_data_i[20]  | ~\new_[18765]_ );
  assign \new_[10657]_  = (~\m7_sel_i[1]  | ~\new_[17239]_ ) & (~\m6_sel_i[1]  | ~\new_[18089]_ );
  assign \new_[10658]_  = (~\m7_data_i[19]  | ~\new_[16296]_ ) & (~\m0_data_i[19]  | ~\new_[20545]_ );
  assign \new_[10659]_  = (~\m7_data_i[18]  | ~\new_[16296]_ ) & (~\m0_data_i[18]  | ~\new_[18765]_ );
  assign \new_[10660]_  = (~\m7_sel_i[0]  | ~\new_[17239]_ ) & (~\m6_sel_i[0]  | ~\new_[18819]_ );
  assign \new_[10661]_  = (~\m7_data_i[17]  | ~\new_[16296]_ ) & (~\m0_data_i[17]  | ~\new_[18765]_ );
  assign \new_[10662]_  = (~\m7_data_i[16]  | ~\new_[16296]_ ) & (~\m0_data_i[16]  | ~\new_[20545]_ );
  assign \new_[10663]_  = (~m5_we_i | ~\new_[18745]_ ) & (~m4_we_i | ~\new_[17271]_ );
  assign \new_[10664]_  = ~\new_[28493]_  & (~\new_[14679]_  | ~\new_[22831]_ );
  assign \new_[10665]_  = (~\m2_data_i[1]  | ~\new_[17222]_ ) & (~\m1_data_i[1]  | ~\new_[18906]_ );
  assign \new_[10666]_  = (~m7_we_i | ~\new_[17239]_ ) & (~m6_we_i | ~\new_[18090]_ );
  assign \new_[10667]_  = (~\m7_data_i[14]  | ~\new_[16296]_ ) & (~\m0_data_i[14]  | ~\new_[18764]_ );
  assign \new_[10668]_  = ~\new_[27881]_  & (~\new_[14693]_  | ~\new_[22613]_ );
  assign \new_[10669]_  = (~\m5_data_i[31]  | ~\new_[18753]_ ) & (~\m6_data_i[31]  | ~\new_[17213]_ );
  assign \new_[10670]_  = ~\new_[14452]_  | ~\new_[22884]_ ;
  assign \new_[10671]_  = ~\new_[29125]_  & (~\new_[14688]_  | ~\new_[20034]_ );
  assign \new_[10672]_  = (~\m7_data_i[4]  | ~\new_[16296]_ ) & (~\m0_data_i[4]  | ~\new_[18767]_ );
  assign \new_[10673]_  = (~\m5_data_i[3]  | ~\new_[18004]_ ) & (~\m6_data_i[3]  | ~\new_[17241]_ );
  assign \new_[10674]_  = (~\m7_data_i[1]  | ~\new_[16296]_ ) & (~\m0_data_i[1]  | ~\new_[20545]_ );
  assign \new_[10675]_  = (~\m5_data_i[30]  | ~\new_[18738]_ ) & (~\m6_data_i[30]  | ~\new_[18030]_ );
  assign \new_[10676]_  = ~\new_[14453]_  | ~\new_[22642]_ ;
  assign \new_[10677]_  = (~\new_[17241]_  | ~\m6_addr_i[31] ) & (~\new_[18004]_  | ~\new_[31001]_ );
  assign \new_[10678]_  = (~\new_[16296]_  | ~\m7_addr_i[31] ) & (~\new_[18766]_  | ~\m0_addr_i[31] );
  assign \new_[10679]_  = ~\new_[26714]_  & (~\new_[14604]_  | ~\new_[22750]_ );
  assign \new_[10680]_  = (~\new_[17241]_  | ~\m6_addr_i[30] ) & (~\new_[18004]_  | ~\new_[31147]_ );
  assign \new_[10681]_  = (~\new_[16296]_  | ~\new_[31531]_ ) & (~\new_[18764]_  | ~\new_[31481]_ );
  assign \new_[10682]_  = ~\new_[27888]_  & (~\new_[14701]_  | ~\new_[18421]_ );
  assign \new_[10683]_  = (~\new_[17241]_  | ~\m6_addr_i[29] ) & (~\new_[18004]_  | ~\new_[31407]_ );
  assign \new_[10684]_  = (~\new_[18095]_  | ~\new_[30577]_ ) & (~\new_[18766]_  | ~\new_[30957]_ );
  assign \new_[10685]_  = (~\m5_data_i[28]  | ~\new_[18738]_ ) & (~\m6_data_i[28]  | ~\new_[18030]_ );
  assign \new_[10686]_  = (~\new_[18095]_  | ~\m7_addr_i[27] ) & (~\new_[18766]_  | ~\m0_addr_i[27] );
  assign \new_[10687]_  = (~\new_[17241]_  | ~\m6_addr_i[26] ) & (~\new_[18004]_  | ~\m5_addr_i[26] );
  assign \new_[10688]_  = (~\m5_data_i[27]  | ~\new_[18738]_ ) & (~\m6_data_i[27]  | ~\new_[18030]_ );
  assign \new_[10689]_  = (~\new_[17241]_  | ~\m6_addr_i[25] ) & (~\new_[18004]_  | ~\m5_addr_i[25] );
  assign \new_[10690]_  = (~\new_[16296]_  | ~\m7_addr_i[24] ) & (~\new_[18764]_  | ~\m0_addr_i[24] );
  assign \new_[10691]_  = (~\new_[17241]_  | ~\m6_addr_i[24] ) & (~\new_[18004]_  | ~\m5_addr_i[24] );
  assign \new_[10692]_  = (~\m7_addr_i[23]  | ~\new_[18095]_ ) & (~\m0_addr_i[23]  | ~\new_[20545]_ );
  assign \new_[10693]_  = (~\m5_addr_i[23]  | ~\new_[18004]_ ) & (~\m6_addr_i[23]  | ~\new_[17241]_ );
  assign \new_[10694]_  = (~\m7_addr_i[22]  | ~\new_[16296]_ ) & (~\m0_addr_i[22]  | ~\new_[18766]_ );
  assign \new_[10695]_  = (~\m5_addr_i[20]  | ~\new_[18004]_ ) & (~\m6_addr_i[20]  | ~\new_[17241]_ );
  assign \new_[10696]_  = (~\m7_addr_i[19]  | ~\new_[16296]_ ) & (~\m0_addr_i[19]  | ~\new_[20545]_ );
  assign \new_[10697]_  = (~\m7_addr_i[18]  | ~\new_[16296]_ ) & (~\m0_addr_i[18]  | ~\new_[20545]_ );
  assign \new_[10698]_  = (~\m5_addr_i[18]  | ~\new_[18004]_ ) & (~\m6_addr_i[18]  | ~\new_[17241]_ );
  assign \new_[10699]_  = (~\m7_addr_i[17]  | ~\new_[16296]_ ) & (~\m0_addr_i[17]  | ~\new_[18764]_ );
  assign \new_[10700]_  = (~\m5_data_i[23]  | ~\new_[18738]_ ) & (~\m6_data_i[23]  | ~\new_[18030]_ );
  assign \new_[10701]_  = (~\m5_addr_i[17]  | ~\new_[18004]_ ) & (~\m6_addr_i[17]  | ~\new_[17241]_ );
  assign \new_[10702]_  = (~\m7_addr_i[16]  | ~\new_[16296]_ ) & (~\m0_addr_i[16]  | ~\new_[18764]_ );
  assign \new_[10703]_  = (~\m7_addr_i[15]  | ~\new_[16296]_ ) & (~\m0_addr_i[15]  | ~\new_[18766]_ );
  assign \new_[10704]_  = (~\m7_addr_i[14]  | ~\new_[16296]_ ) & (~\m0_addr_i[14]  | ~\new_[18766]_ );
  assign \new_[10705]_  = (~\m7_addr_i[13]  | ~\new_[16296]_ ) & (~\m0_addr_i[13]  | ~\new_[18766]_ );
  assign \new_[10706]_  = (~\m7_addr_i[12]  | ~\new_[16296]_ ) & (~\m0_addr_i[12]  | ~\new_[20545]_ );
  assign \new_[10707]_  = (~\m5_data_i[20]  | ~\new_[18738]_ ) & (~\m6_data_i[20]  | ~\new_[18030]_ );
  assign \new_[10708]_  = (~\m7_addr_i[11]  | ~\new_[16296]_ ) & (~\m0_addr_i[11]  | ~\new_[20545]_ );
  assign \new_[10709]_  = (~\m7_addr_i[10]  | ~\new_[16296]_ ) & (~\m0_addr_i[10]  | ~\new_[18766]_ );
  assign \new_[10710]_  = (~\m7_addr_i[9]  | ~\new_[16296]_ ) & (~\m0_addr_i[9]  | ~\new_[18766]_ );
  assign \new_[10711]_  = (~\m7_addr_i[8]  | ~\new_[16296]_ ) & (~\m0_addr_i[8]  | ~\new_[20545]_ );
  assign \new_[10712]_  = (~\m5_data_i[18]  | ~\new_[18738]_ ) & (~\m6_data_i[18]  | ~\new_[18030]_ );
  assign \new_[10713]_  = (~\m7_addr_i[7]  | ~\new_[16296]_ ) & (~\m0_addr_i[7]  | ~\new_[18763]_ );
  assign \new_[10714]_  = (~\m7_addr_i[6]  | ~\new_[16296]_ ) & (~\m0_addr_i[6]  | ~\new_[18763]_ );
  assign \new_[10715]_  = (~\m5_data_i[17]  | ~\new_[18738]_ ) & (~\m6_data_i[17]  | ~\new_[18030]_ );
  assign \new_[10716]_  = (~\m7_addr_i[5]  | ~\new_[16296]_ ) & (~\new_[31848]_  | ~\new_[18764]_ );
  assign \new_[10717]_  = ~\new_[14418]_  | ~\new_[19446]_ ;
  assign \new_[10718]_  = (~\m5_addr_i[4]  | ~\new_[18004]_ ) & (~\m6_addr_i[4]  | ~\new_[17241]_ );
  assign \new_[10719]_  = (~\m5_data_i[16]  | ~\new_[18738]_ ) & (~\m6_data_i[16]  | ~\new_[18030]_ );
  assign \new_[10720]_  = (~\new_[31726]_  | ~\new_[18095]_ ) & (~\m0_addr_i[3]  | ~\new_[18762]_ );
  assign \new_[10721]_  = (~\m5_addr_i[3]  | ~\new_[18004]_ ) & (~\m6_addr_i[3]  | ~\new_[17241]_ );
  assign \new_[10722]_  = (~\m7_addr_i[2]  | ~\new_[18095]_ ) & (~\m0_addr_i[2]  | ~\new_[18762]_ );
  assign \new_[10723]_  = (~\m5_data_i[15]  | ~\new_[18738]_ ) & (~\m6_data_i[15]  | ~\new_[18030]_ );
  assign \new_[10724]_  = (~\m7_addr_i[1]  | ~\new_[18095]_ ) & (~\m0_addr_i[1]  | ~\new_[18762]_ );
  assign \new_[10725]_  = (~\m7_sel_i[1]  | ~\new_[18095]_ ) & (~\m0_sel_i[1]  | ~\new_[18762]_ );
  assign \new_[10726]_  = (~\m5_sel_i[0]  | ~\new_[18004]_ ) & (~\m6_sel_i[0]  | ~\new_[17241]_ );
  assign \new_[10727]_  = (~m7_we_i | ~\new_[18095]_ ) & (~m0_we_i | ~\new_[18762]_ );
  assign \new_[10728]_  = (~m5_we_i | ~\new_[18004]_ ) & (~m6_we_i | ~\new_[17241]_ );
  assign \new_[10729]_  = (~\m2_data_i[31]  | ~\new_[17218]_ ) & (~\m1_data_i[31]  | ~\new_[18905]_ );
  assign \new_[10730]_  = (~\m4_data_i[31]  | ~\new_[17266]_ ) & (~\m3_data_i[31]  | ~\new_[18128]_ );
  assign \new_[10731]_  = (~\m5_data_i[31]  | ~\new_[17196]_ ) & (~\m6_data_i[31]  | ~\new_[18045]_ );
  assign \new_[10732]_  = (~\m2_data_i[30]  | ~\new_[17218]_ ) & (~\m1_data_i[30]  | ~\new_[18905]_ );
  assign \new_[10733]_  = (~\m4_data_i[30]  | ~\new_[17265]_ ) & (~\m3_data_i[30]  | ~\new_[17248]_ );
  assign \new_[10734]_  = ~\new_[13154]_  & (~\new_[28992]_  | ~\new_[5909]_ );
  assign \new_[10735]_  = (~\m5_data_i[30]  | ~\new_[17196]_ ) & (~\m6_data_i[30]  | ~\new_[18043]_ );
  assign \new_[10736]_  = (~\m5_data_i[29]  | ~\new_[17196]_ ) & (~\m6_data_i[29]  | ~\new_[19562]_ );
  assign \new_[10737]_  = (~\m4_data_i[29]  | ~\new_[17266]_ ) & (~\m3_data_i[29]  | ~\new_[18128]_ );
  assign \new_[10738]_  = ~\new_[13157]_  & (~\new_[29541]_  | ~\new_[5911]_ );
  assign \new_[10739]_  = (~\m5_data_i[28]  | ~\new_[17196]_ ) & (~\m6_data_i[28]  | ~\new_[18045]_ );
  assign \new_[10740]_  = (~\m2_data_i[27]  | ~\new_[17218]_ ) & (~\m1_data_i[27]  | ~\new_[18905]_ );
  assign \new_[10741]_  = ~\new_[13161]_  & (~\new_[29217]_  | ~\new_[5912]_ );
  assign \new_[10742]_  = (~\m5_data_i[27]  | ~\new_[17196]_ ) & (~\m6_data_i[27]  | ~\new_[18044]_ );
  assign \new_[10743]_  = (~\m2_data_i[26]  | ~\new_[17218]_ ) & (~\m1_data_i[26]  | ~\new_[18905]_ );
  assign \new_[10744]_  = ~\new_[13165]_  & (~\new_[29058]_  | ~\new_[5914]_ );
  assign \new_[10745]_  = (~\m4_data_i[26]  | ~\new_[17264]_ ) & (~\m3_data_i[26]  | ~\new_[17248]_ );
  assign \new_[10746]_  = (~\m5_data_i[26]  | ~\new_[17195]_ ) & (~\m6_data_i[26]  | ~\new_[19562]_ );
  assign \new_[10747]_  = (~\m4_data_i[25]  | ~\new_[17264]_ ) & (~\m3_data_i[25]  | ~\new_[18128]_ );
  assign \new_[10748]_  = (~\m5_data_i[25]  | ~\new_[17196]_ ) & (~\m6_data_i[25]  | ~\new_[18046]_ );
  assign \new_[10749]_  = (~\m2_data_i[24]  | ~\new_[17218]_ ) & (~\m1_data_i[24]  | ~\new_[18905]_ );
  assign \new_[10750]_  = (~\m4_data_i[24]  | ~\new_[17266]_ ) & (~\m3_data_i[24]  | ~\new_[17248]_ );
  assign \new_[10751]_  = (~\m5_data_i[24]  | ~\new_[17196]_ ) & (~\m6_data_i[24]  | ~\new_[18043]_ );
  assign \new_[10752]_  = (~\m4_data_i[23]  | ~\new_[17264]_ ) & (~\m3_data_i[23]  | ~\new_[18849]_ );
  assign \new_[10753]_  = ~\new_[13170]_  & (~\new_[29254]_  | ~\new_[5917]_ );
  assign \new_[10754]_  = (~\m4_data_i[22]  | ~\new_[17264]_ ) & (~\m3_data_i[22]  | ~\new_[18849]_ );
  assign \new_[10755]_  = ~\new_[13174]_  & (~\new_[29115]_  | ~\new_[5918]_ );
  assign \new_[10756]_  = (~\m4_data_i[21]  | ~\new_[17265]_ ) & (~\m3_data_i[21]  | ~\new_[18849]_ );
  assign \new_[10757]_  = ~\new_[13175]_  & (~\new_[29101]_  | ~\new_[5921]_ );
  assign \new_[10758]_  = ~\new_[13178]_  & (~\new_[29229]_  | ~\new_[5923]_ );
  assign \new_[10759]_  = (~\m4_data_i[20]  | ~\new_[17264]_ ) & (~\m3_data_i[20]  | ~\new_[18849]_ );
  assign \new_[10760]_  = (~\m2_data_i[19]  | ~\new_[17218]_ ) & (~\m1_data_i[19]  | ~\new_[18905]_ );
  assign \new_[10761]_  = (~\m4_data_i[19]  | ~\new_[17265]_ ) & (~\m3_data_i[19]  | ~\new_[17248]_ );
  assign \new_[10762]_  = (~\m5_data_i[19]  | ~\new_[17196]_ ) & (~\m6_data_i[19]  | ~\new_[18047]_ );
  assign \new_[10763]_  = (~\m4_data_i[18]  | ~\new_[17266]_ ) & (~\m3_data_i[18]  | ~\new_[18128]_ );
  assign \new_[10764]_  = (~\m5_data_i[18]  | ~\new_[17195]_ ) & (~\m6_data_i[18]  | ~\new_[18047]_ );
  assign \new_[10765]_  = (~\m4_data_i[17]  | ~\new_[17264]_ ) & (~\m3_data_i[17]  | ~\new_[17248]_ );
  assign \new_[10766]_  = (~\m5_data_i[17]  | ~\new_[17196]_ ) & (~\m6_data_i[17]  | ~\new_[19562]_ );
  assign \new_[10767]_  = ~\new_[13184]_  & (~\new_[29167]_  | ~\new_[5927]_ );
  assign \new_[10768]_  = (~\m4_data_i[16]  | ~\new_[17266]_ ) & (~\m3_data_i[16]  | ~\new_[17248]_ );
  assign \new_[10769]_  = (~\m5_data_i[16]  | ~\new_[17196]_ ) & (~\m6_data_i[16]  | ~\new_[18047]_ );
  assign \new_[10770]_  = (~\m2_data_i[15]  | ~\new_[17218]_ ) & (~\m1_data_i[15]  | ~\new_[18905]_ );
  assign \new_[10771]_  = (~\m4_data_i[15]  | ~\new_[17265]_ ) & (~\m3_data_i[15]  | ~\new_[18849]_ );
  assign \new_[10772]_  = (~\m5_data_i[15]  | ~\new_[17196]_ ) & (~\m6_data_i[15]  | ~\new_[18045]_ );
  assign \new_[10773]_  = (~\m2_data_i[14]  | ~\new_[17218]_ ) & (~\m1_data_i[14]  | ~\new_[18905]_ );
  assign \new_[10774]_  = (~\m4_data_i[14]  | ~\new_[17265]_ ) & (~\m3_data_i[14]  | ~\new_[17248]_ );
  assign \new_[10775]_  = (~\m5_data_i[14]  | ~\new_[17196]_ ) & (~\m6_data_i[14]  | ~\new_[19562]_ );
  assign \new_[10776]_  = (~\m4_data_i[13]  | ~\new_[17264]_ ) & (~\m3_data_i[13]  | ~\new_[17248]_ );
  assign \new_[10777]_  = (~\m2_data_i[12]  | ~\new_[17218]_ ) & (~\m1_data_i[12]  | ~\new_[18905]_ );
  assign \new_[10778]_  = (~\m5_data_i[0]  | ~\new_[18738]_ ) & (~\m6_data_i[0]  | ~\new_[18030]_ );
  assign \new_[10779]_  = (~\m4_data_i[12]  | ~\new_[17265]_ ) & (~\m3_data_i[12]  | ~\new_[17248]_ );
  assign \new_[10780]_  = (~\m4_data_i[11]  | ~\new_[17265]_ ) & (~\m3_data_i[11]  | ~\new_[17248]_ );
  assign \new_[10781]_  = (~\m4_data_i[10]  | ~\new_[17264]_ ) & (~\m3_data_i[10]  | ~\new_[18849]_ );
  assign \new_[10782]_  = (~\m2_data_i[10]  | ~\new_[17218]_ ) & (~\m1_data_i[10]  | ~\new_[18905]_ );
  assign \new_[10783]_  = (~\m5_data_i[10]  | ~\new_[17196]_ ) & (~\m6_data_i[10]  | ~\new_[19562]_ );
  assign \new_[10784]_  = (~\m2_data_i[9]  | ~\new_[17218]_ ) & (~\m1_data_i[9]  | ~\new_[18905]_ );
  assign \new_[10785]_  = (~\m5_data_i[9]  | ~\new_[17195]_ ) & (~\m6_data_i[9]  | ~\new_[18043]_ );
  assign \new_[10786]_  = (~\m4_data_i[8]  | ~\new_[17265]_ ) & (~\m3_data_i[8]  | ~\new_[17248]_ );
  assign \new_[10787]_  = (~\m2_data_i[7]  | ~\new_[17218]_ ) & (~\m1_data_i[7]  | ~\new_[18905]_ );
  assign \new_[10788]_  = (~\m4_data_i[7]  | ~\new_[17265]_ ) & (~\m3_data_i[7]  | ~\new_[17248]_ );
  assign \new_[10789]_  = (~\m5_data_i[7]  | ~\new_[17196]_ ) & (~\m6_data_i[7]  | ~\new_[18047]_ );
  assign \new_[10790]_  = (~\m2_data_i[6]  | ~\new_[17218]_ ) & (~\m1_data_i[6]  | ~\new_[18905]_ );
  assign \new_[10791]_  = (~\m4_data_i[6]  | ~\new_[17265]_ ) & (~\m3_data_i[6]  | ~\new_[17248]_ );
  assign \new_[10792]_  = (~\m4_data_i[4]  | ~\new_[17265]_ ) & (~\m3_data_i[4]  | ~\new_[17248]_ );
  assign \new_[10793]_  = (~\m5_data_i[4]  | ~\new_[17195]_ ) & (~\m6_data_i[4]  | ~\new_[18043]_ );
  assign \new_[10794]_  = (~\m5_data_i[3]  | ~\new_[17195]_ ) & (~\m6_data_i[3]  | ~\new_[19562]_ );
  assign \new_[10795]_  = (~\m4_data_i[2]  | ~\new_[17264]_ ) & (~\m3_data_i[2]  | ~\new_[18849]_ );
  assign \new_[10796]_  = (~\m4_data_i[1]  | ~\new_[17264]_ ) & (~\m3_data_i[1]  | ~\new_[18849]_ );
  assign \new_[10797]_  = (~\m2_data_i[0]  | ~\new_[17218]_ ) & (~\m1_data_i[0]  | ~\new_[18905]_ );
  assign \new_[10798]_  = \new_[14608]_  ? \new_[30245]_  : \new_[6036]_ ;
  assign \new_[10799]_  = (~\m5_data_i[0]  | ~\new_[17195]_ ) & (~\m6_data_i[0]  | ~\new_[18043]_ );
  assign \new_[10800]_  = (~\m4_data_i[0]  | ~\new_[17264]_ ) & (~\m3_data_i[0]  | ~\new_[17248]_ );
  assign \new_[10801]_  = (~\new_[18792]_  | ~\m6_addr_i[31] ) & (~\new_[17195]_  | ~\new_[31001]_ );
  assign \new_[10802]_  = \new_[14612]_  ? \new_[29908]_  : \new_[6042]_ ;
  assign \new_[10803]_  = (~\new_[17264]_  | ~\m4_addr_i[31] ) & (~\new_[17248]_  | ~\m3_addr_i[31] );
  assign \new_[10804]_  = (~\new_[17264]_  | ~\m4_addr_i[30] ) & (~\new_[18849]_  | ~\m3_addr_i[30] );
  assign \new_[10805]_  = (~\new_[18792]_  | ~\m6_addr_i[30] ) & (~\new_[17195]_  | ~\new_[31147]_ );
  assign \new_[10806]_  = \new_[14620]_  ? \new_[29765]_  : \new_[6045]_ ;
  assign \new_[10807]_  = (~\new_[18792]_  | ~\m6_addr_i[29] ) & (~\new_[17195]_  | ~\new_[31407]_ );
  assign \new_[10808]_  = (~\new_[17264]_  | ~\m4_addr_i[29] ) & (~\new_[18849]_  | ~\m3_addr_i[29] );
  assign \new_[10809]_  = \new_[14732]_  ? \new_[30268]_  : \new_[6051]_ ;
  assign \new_[10810]_  = (~\new_[17218]_  | ~\new_[31547]_ ) & (~\new_[18905]_  | ~\new_[31458]_ );
  assign \new_[10811]_  = ~\new_[28120]_  & (~\new_[14823]_  | ~\new_[29397]_ );
  assign \new_[10812]_  = (~\new_[17265]_  | ~\m4_addr_i[28] ) & (~\new_[18849]_  | ~\m3_addr_i[28] );
  assign \new_[10813]_  = (~\m5_data_i[4]  | ~\new_[18755]_ ) & (~\m6_data_i[4]  | ~\new_[17213]_ );
  assign \new_[10814]_  = (~\m5_addr_i[23]  | ~\new_[18738]_ ) & (~\m6_addr_i[23]  | ~\new_[18030]_ );
  assign \new_[10815]_  = (~\new_[17265]_  | ~\m4_addr_i[26] ) & (~\new_[18128]_  | ~\m3_addr_i[26] );
  assign \new_[10816]_  = (~\m5_data_i[31]  | ~\new_[18738]_ ) & (~\m6_data_i[31]  | ~\new_[18030]_ );
  assign \new_[10817]_  = (~\m5_addr_i[22]  | ~\new_[18738]_ ) & (~\m6_addr_i[22]  | ~\new_[18030]_ );
  assign \new_[10818]_  = (~\new_[17265]_  | ~\m4_addr_i[25] ) & (~\new_[18128]_  | ~\m3_addr_i[25] );
  assign \new_[10819]_  = (~\m7_addr_i[21]  | ~\new_[16296]_ ) & (~\m0_addr_i[21]  | ~\new_[20545]_ );
  assign \new_[10820]_  = \new_[14671]_  ? \new_[29914]_  : \new_[6067]_ ;
  assign \new_[10821]_  = (~\new_[17265]_  | ~\m4_addr_i[24] ) & (~\new_[18849]_  | ~\m3_addr_i[24] );
  assign \new_[10822]_  = \new_[14678]_  ? \new_[30304]_  : \new_[6193]_ ;
  assign \new_[10823]_  = (~\m2_addr_i[23]  | ~\new_[17218]_ ) & (~\m1_addr_i[23]  | ~\new_[18905]_ );
  assign \new_[10824]_  = (~\m4_addr_i[23]  | ~\new_[17266]_ ) & (~\m3_addr_i[23]  | ~\new_[17248]_ );
  assign \new_[10825]_  = (~\m5_addr_i[23]  | ~\new_[17196]_ ) & (~\m6_addr_i[23]  | ~\new_[18043]_ );
  assign \new_[10826]_  = \new_[14666]_  ? \new_[30062]_  : \new_[6074]_ ;
  assign \new_[10827]_  = (~\m5_addr_i[21]  | ~\new_[18738]_ ) & (~\m6_addr_i[21]  | ~\new_[18030]_ );
  assign \new_[10828]_  = (~\m2_addr_i[22]  | ~\new_[17218]_ ) & (~\m1_addr_i[22]  | ~\new_[18905]_ );
  assign \new_[10829]_  = (~\m4_addr_i[22]  | ~\new_[17266]_ ) & (~\m3_addr_i[22]  | ~\new_[17248]_ );
  assign \new_[10830]_  = (~\m5_addr_i[22]  | ~\new_[17196]_ ) & (~\m6_addr_i[22]  | ~\new_[19562]_ );
  assign \new_[10831]_  = \new_[14615]_  ? \new_[30267]_  : \new_[6075]_ ;
  assign \new_[10832]_  = (~\m2_addr_i[21]  | ~\new_[17218]_ ) & (~\m1_addr_i[21]  | ~\new_[18905]_ );
  assign \new_[10833]_  = (~\m4_addr_i[21]  | ~\new_[17266]_ ) & (~\m3_addr_i[21]  | ~\new_[18128]_ );
  assign \new_[10834]_  = (~\m5_addr_i[21]  | ~\new_[17196]_ ) & (~\m6_addr_i[21]  | ~\new_[19562]_ );
  assign \new_[10835]_  = (~\m5_addr_i[20]  | ~\new_[18738]_ ) & (~\m6_addr_i[20]  | ~\new_[18030]_ );
  assign \new_[10836]_  = (~\m4_addr_i[20]  | ~\new_[17264]_ ) & (~\m3_addr_i[20]  | ~\new_[18128]_ );
  assign \new_[10837]_  = (~\m5_addr_i[20]  | ~\new_[17196]_ ) & (~\m6_addr_i[20]  | ~\new_[19562]_ );
  assign \new_[10838]_  = \new_[14697]_  ? \new_[30024]_  : \new_[6083]_ ;
  assign \new_[10839]_  = (~\m4_addr_i[19]  | ~\new_[17266]_ ) & (~\m3_addr_i[19]  | ~\new_[18128]_ );
  assign \new_[10840]_  = (~\m5_addr_i[19]  | ~\new_[17196]_ ) & (~\m6_addr_i[19]  | ~\new_[19562]_ );
  assign \new_[10841]_  = ~\new_[27675]_  & (~\new_[14822]_  | ~\new_[29817]_ );
  assign \new_[10842]_  = (~\m4_addr_i[18]  | ~\new_[17266]_ ) & (~\m3_addr_i[18]  | ~\new_[17248]_ );
  assign \new_[10843]_  = (~\m5_addr_i[18]  | ~\new_[17195]_ ) & (~\m6_addr_i[18]  | ~\new_[18043]_ );
  assign \new_[10844]_  = (~\m4_addr_i[17]  | ~\new_[17266]_ ) & (~\m3_addr_i[17]  | ~\new_[17248]_ );
  assign \new_[10845]_  = (~\m5_addr_i[17]  | ~\new_[17196]_ ) & (~\m6_addr_i[17]  | ~\new_[18043]_ );
  assign \new_[10846]_  = (~\m2_addr_i[16]  | ~\new_[17218]_ ) & (~\m1_addr_i[16]  | ~\new_[18905]_ );
  assign \new_[10847]_  = (~\m4_addr_i[16]  | ~\new_[17266]_ ) & (~\m3_addr_i[16]  | ~\new_[17248]_ );
  assign \new_[10848]_  = (~\m5_addr_i[16]  | ~\new_[17196]_ ) & (~\m6_addr_i[16]  | ~\new_[18044]_ );
  assign \new_[10849]_  = (~\m2_addr_i[15]  | ~\new_[17218]_ ) & (~\m1_addr_i[15]  | ~\new_[18905]_ );
  assign \new_[10850]_  = (~\m4_addr_i[15]  | ~\new_[17266]_ ) & (~\m3_addr_i[15]  | ~\new_[18128]_ );
  assign \new_[10851]_  = (~\m5_addr_i[15]  | ~\new_[17196]_ ) & (~\m6_addr_i[15]  | ~\new_[18043]_ );
  assign \new_[10852]_  = (~\m2_addr_i[14]  | ~\new_[17218]_ ) & (~\m1_addr_i[14]  | ~\new_[18905]_ );
  assign \new_[10853]_  = (~\m4_addr_i[14]  | ~\new_[17266]_ ) & (~\m3_addr_i[14]  | ~\new_[17248]_ );
  assign \new_[10854]_  = (~\m5_addr_i[14]  | ~\new_[17196]_ ) & (~\m6_addr_i[14]  | ~\new_[19562]_ );
  assign \new_[10855]_  = (~\m2_addr_i[13]  | ~\new_[17218]_ ) & (~\m1_addr_i[13]  | ~\new_[18905]_ );
  assign \new_[10856]_  = (~\m4_addr_i[13]  | ~\new_[17266]_ ) & (~\m3_addr_i[13]  | ~\new_[18128]_ );
  assign \new_[10857]_  = (~\m5_addr_i[13]  | ~\new_[17196]_ ) & (~\m6_addr_i[13]  | ~\new_[18046]_ );
  assign \new_[10858]_  = (~\m2_addr_i[12]  | ~\new_[17218]_ ) & (~\m1_addr_i[12]  | ~\new_[18905]_ );
  assign \new_[10859]_  = (~\m4_addr_i[12]  | ~\new_[17264]_ ) & (~\m3_addr_i[12]  | ~\new_[18128]_ );
  assign \new_[10860]_  = (~\m5_addr_i[12]  | ~\new_[17195]_ ) & (~\m6_addr_i[12]  | ~\new_[19562]_ );
  assign \new_[10861]_  = (~\m2_addr_i[11]  | ~\new_[17218]_ ) & (~\m1_addr_i[11]  | ~\new_[18905]_ );
  assign \new_[10862]_  = (~\m4_addr_i[11]  | ~\new_[17265]_ ) & (~\m3_addr_i[11]  | ~\new_[18128]_ );
  assign \new_[10863]_  = (~\m5_addr_i[11]  | ~\new_[17195]_ ) & (~\m6_addr_i[11]  | ~\new_[18046]_ );
  assign \new_[10864]_  = (~\m2_addr_i[10]  | ~\new_[17218]_ ) & (~\m1_addr_i[10]  | ~\new_[18905]_ );
  assign \new_[10865]_  = (~\m5_addr_i[19]  | ~\new_[18748]_ ) & (~\m6_addr_i[19]  | ~\new_[17213]_ );
  assign \new_[10866]_  = (~\m4_addr_i[10]  | ~\new_[17265]_ ) & (~\m3_addr_i[10]  | ~\new_[17248]_ );
  assign \new_[10867]_  = (~\m5_addr_i[10]  | ~\new_[17196]_ ) & (~\m6_addr_i[10]  | ~\new_[18043]_ );
  assign \new_[10868]_  = (~\m2_addr_i[9]  | ~\new_[17218]_ ) & (~\m1_addr_i[9]  | ~\new_[18905]_ );
  assign \new_[10869]_  = (~\m4_addr_i[9]  | ~\new_[17266]_ ) & (~\m3_addr_i[9]  | ~\new_[17248]_ );
  assign \new_[10870]_  = (~\m5_addr_i[9]  | ~\new_[17196]_ ) & (~\m6_addr_i[9]  | ~\new_[19562]_ );
  assign \new_[10871]_  = (~\m4_addr_i[8]  | ~\new_[17265]_ ) & (~\m3_addr_i[8]  | ~\new_[18849]_ );
  assign \new_[10872]_  = (~\m5_addr_i[8]  | ~\new_[17195]_ ) & (~\m6_addr_i[8]  | ~\new_[19562]_ );
  assign \new_[10873]_  = (~\m5_addr_i[7]  | ~\new_[17195]_ ) & (~\m6_addr_i[7]  | ~\new_[19562]_ );
  assign \new_[10874]_  = (~\m4_addr_i[7]  | ~\new_[17264]_ ) & (~\m3_addr_i[7]  | ~\new_[17248]_ );
  assign \new_[10875]_  = (~\m4_addr_i[6]  | ~\new_[17265]_ ) & (~\m3_addr_i[6]  | ~\new_[18849]_ );
  assign \new_[10876]_  = (~\m5_addr_i[6]  | ~\new_[17196]_ ) & (~\m6_addr_i[6]  | ~\new_[18045]_ );
  assign \new_[10877]_  = (~\m2_addr_i[5]  | ~\new_[17218]_ ) & (~\m1_addr_i[5]  | ~\new_[18905]_ );
  assign \new_[10878]_  = (~\m4_addr_i[5]  | ~\new_[17265]_ ) & (~\m3_addr_i[5]  | ~\new_[17248]_ );
  assign \new_[10879]_  = (~\m5_addr_i[5]  | ~\new_[17195]_ ) & (~\m6_addr_i[5]  | ~\new_[19562]_ );
  assign \new_[10880]_  = (~\m5_addr_i[12]  | ~\new_[18738]_ ) & (~\m6_addr_i[12]  | ~\new_[18030]_ );
  assign \new_[10881]_  = (~\m4_addr_i[4]  | ~\new_[17265]_ ) & (~\m3_addr_i[4]  | ~\new_[17248]_ );
  assign \new_[10882]_  = (~\m5_addr_i[4]  | ~\new_[17196]_ ) & (~\m6_addr_i[4]  | ~\new_[18044]_ );
  assign \new_[10883]_  = (~\m2_addr_i[3]  | ~\new_[17218]_ ) & (~\m1_addr_i[3]  | ~\new_[18905]_ );
  assign \new_[10884]_  = (~\m4_addr_i[3]  | ~\new_[17265]_ ) & (~\m3_addr_i[3]  | ~\new_[18128]_ );
  assign \new_[10885]_  = (~\m5_addr_i[3]  | ~\new_[17196]_ ) & (~\m6_addr_i[3]  | ~\new_[18044]_ );
  assign \new_[10886]_  = (~\m5_addr_i[2]  | ~\new_[17196]_ ) & (~\m6_addr_i[2]  | ~\new_[19562]_ );
  assign \new_[10887]_  = (~\new_[17241]_  | ~\m6_addr_i[28] ) & (~\new_[18004]_  | ~\new_[31276]_ );
  assign \new_[10888]_  = (~\m4_addr_i[1]  | ~\new_[17265]_ ) & (~\m3_addr_i[1]  | ~\new_[17248]_ );
  assign \new_[10889]_  = (~\m5_addr_i[1]  | ~\new_[17196]_ ) & (~\m6_addr_i[1]  | ~\new_[18043]_ );
  assign \new_[10890]_  = (~\m4_addr_i[0]  | ~\new_[17264]_ ) & (~\m3_addr_i[0]  | ~\new_[18849]_ );
  assign \new_[10891]_  = (~\m5_addr_i[0]  | ~\new_[17195]_ ) & (~\m6_addr_i[0]  | ~\new_[19562]_ );
  assign \new_[10892]_  = (~\m4_sel_i[3]  | ~\new_[17264]_ ) & (~\m3_sel_i[3]  | ~\new_[18849]_ );
  assign \new_[10893]_  = (~\m5_sel_i[3]  | ~\new_[17195]_ ) & (~\m6_sel_i[3]  | ~\new_[19562]_ );
  assign \new_[10894]_  = (~\m4_sel_i[2]  | ~\new_[17264]_ ) & (~\m3_sel_i[2]  | ~\new_[18849]_ );
  assign \new_[10895]_  = (~\m5_sel_i[2]  | ~\new_[17195]_ ) & (~\m6_sel_i[2]  | ~\new_[18043]_ );
  assign \new_[10896]_  = (~\m2_sel_i[1]  | ~\new_[17218]_ ) & (~\m1_sel_i[1]  | ~\new_[18905]_ );
  assign \new_[10897]_  = (~\m5_sel_i[1]  | ~\new_[17195]_ ) & (~\m6_sel_i[1]  | ~\new_[19562]_ );
  assign \new_[10898]_  = (~\m4_sel_i[1]  | ~\new_[17265]_ ) & (~\m3_sel_i[1]  | ~\new_[18128]_ );
  assign \new_[10899]_  = (~\m2_sel_i[0]  | ~\new_[17218]_ ) & (~\m1_sel_i[0]  | ~\new_[18905]_ );
  assign \new_[10900]_  = (~\m4_sel_i[0]  | ~\new_[17265]_ ) & (~\m3_sel_i[0]  | ~\new_[18128]_ );
  assign \new_[10901]_  = (~\m5_sel_i[0]  | ~\new_[17196]_ ) & (~\m6_sel_i[0]  | ~\new_[18043]_ );
  assign \new_[10902]_  = (~m2_we_i | ~\new_[17218]_ ) & (~m1_we_i | ~\new_[18905]_ );
  assign \new_[10903]_  = (~m5_we_i | ~\new_[17195]_ ) & (~m6_we_i | ~\new_[18046]_ );
  assign \new_[10904]_  = (~\new_[14934]_  | ~\new_[27941]_ ) & (~\new_[14933]_  | ~\new_[28645]_ );
  assign \new_[10905]_  = (~\m4_data_i[31]  | ~\new_[17272]_ ) & (~\m3_data_i[31]  | ~\new_[17278]_ );
  assign \new_[10906]_  = (~\m7_data_i[31]  | ~\new_[18096]_ ) & (~\m0_data_i[31]  | ~\new_[18083]_ );
  assign \new_[10907]_  = (~\m2_data_i[31]  | ~\new_[16290]_ ) & (~\m1_data_i[31]  | ~\new_[18174]_ );
  assign \new_[10908]_  = (~\m2_data_i[30]  | ~\new_[18070]_ ) & (~\m1_data_i[30]  | ~\new_[18172]_ );
  assign \new_[10909]_  = (~\m4_data_i[30]  | ~\new_[17272]_ ) & (~\m3_data_i[30]  | ~\new_[17280]_ );
  assign \new_[10910]_  = (~\m7_data_i[30]  | ~\new_[16297]_ ) & (~\m0_data_i[30]  | ~\new_[19575]_ );
  assign \new_[10911]_  = (~\m2_data_i[29]  | ~\new_[18070]_ ) & (~\m1_data_i[29]  | ~\new_[18172]_ );
  assign \new_[10912]_  = (~\m4_data_i[29]  | ~\new_[17272]_ ) & (~\m3_data_i[29]  | ~\new_[17279]_ );
  assign \new_[10913]_  = (~\m7_data_i[29]  | ~\new_[16297]_ ) & (~\m0_data_i[29]  | ~\new_[19575]_ );
  assign \new_[10914]_  = (~\m4_data_i[28]  | ~\new_[17272]_ ) & (~\m3_data_i[28]  | ~\new_[17278]_ );
  assign \new_[10915]_  = (~\m2_data_i[27]  | ~\new_[16290]_ ) & (~\m1_data_i[27]  | ~\new_[18174]_ );
  assign \new_[10916]_  = (~\m4_data_i[27]  | ~\new_[17272]_ ) & (~\m3_data_i[27]  | ~\new_[18927]_ );
  assign \new_[10917]_  = (~\m5_data_i[13]  | ~\new_[18015]_ ) & (~\m6_data_i[13]  | ~\new_[17229]_ );
  assign \new_[10918]_  = (~\m2_data_i[26]  | ~\new_[16290]_ ) & (~\m1_data_i[26]  | ~\new_[19627]_ );
  assign \new_[10919]_  = (~\m4_data_i[26]  | ~\new_[17272]_ ) & (~\m3_data_i[26]  | ~\new_[17278]_ );
  assign \new_[10920]_  = (~\m7_data_i[25]  | ~\new_[18096]_ ) & (~\m0_data_i[25]  | ~\new_[18083]_ );
  assign \new_[10921]_  = (~\m4_data_i[25]  | ~\new_[17272]_ ) & (~\m3_data_i[25]  | ~\new_[18927]_ );
  assign \new_[10922]_  = (~\new_[14939]_  | ~\new_[28699]_ ) & (~\new_[14938]_  | ~\new_[29423]_ );
  assign \new_[10923]_  = (~\m4_data_i[24]  | ~\new_[17272]_ ) & (~\m3_data_i[24]  | ~\new_[18927]_ );
  assign \new_[10924]_  = (~\m4_data_i[23]  | ~\new_[17272]_ ) & (~\m3_data_i[23]  | ~\new_[18927]_ );
  assign \new_[10925]_  = (~\m4_data_i[22]  | ~\new_[17272]_ ) & (~\m3_data_i[22]  | ~\new_[18927]_ );
  assign \new_[10926]_  = (~\m2_addr_i[6]  | ~\new_[17193]_ ) & (~\m1_addr_i[6]  | ~\new_[19633]_ );
  assign \new_[10927]_  = (~\m4_data_i[21]  | ~\new_[17272]_ ) & (~\m3_data_i[21]  | ~\new_[17278]_ );
  assign \new_[10928]_  = (~\m7_data_i[21]  | ~\new_[16297]_ ) & (~\m0_data_i[21]  | ~\new_[19575]_ );
  assign \new_[10929]_  = (~\m7_addr_i[4]  | ~\new_[16296]_ ) & (~\m0_addr_i[4]  | ~\new_[18764]_ );
  assign \new_[10930]_  = ~\new_[17016]_  | ~\new_[18653]_  | ~\new_[13349]_  | ~\new_[17018]_ ;
  assign \new_[10931]_  = (~\m2_data_i[20]  | ~\new_[16290]_ ) & (~\m1_data_i[20]  | ~\new_[19627]_ );
  assign \new_[10932]_  = (~\m4_data_i[20]  | ~\new_[17272]_ ) & (~\m3_data_i[20]  | ~\new_[17280]_ );
  assign \new_[10933]_  = (~\new_[14941]_  | ~\new_[27841]_ ) & (~\new_[14940]_  | ~\new_[28764]_ );
  assign \new_[10934]_  = (~\m2_data_i[19]  | ~\new_[18070]_ ) & (~\m1_data_i[19]  | ~\new_[18172]_ );
  assign \new_[10935]_  = (~\m4_data_i[19]  | ~\new_[17272]_ ) & (~\m3_data_i[19]  | ~\new_[17280]_ );
  assign \new_[10936]_  = (~\m7_data_i[19]  | ~\new_[16297]_ ) & (~\m0_data_i[19]  | ~\new_[19575]_ );
  assign \new_[10937]_  = ~\new_[17026]_  | ~\new_[18656]_  | ~\new_[13364]_  | ~\new_[17025]_ ;
  assign \new_[10938]_  = (~\m2_data_i[18]  | ~\new_[16290]_ ) & (~\m1_data_i[18]  | ~\new_[18174]_ );
  assign \new_[10939]_  = (~\m5_sel_i[2]  | ~\new_[18738]_ ) & (~\m6_sel_i[2]  | ~\new_[18030]_ );
  assign \new_[10940]_  = (~\m4_data_i[18]  | ~\new_[17272]_ ) & (~\m3_data_i[18]  | ~\new_[18927]_ );
  assign \new_[10941]_  = (~\m7_data_i[17]  | ~\new_[16297]_ ) & (~\m0_data_i[17]  | ~\new_[19575]_ );
  assign \new_[10942]_  = ~\new_[16183]_  | ~\new_[16156]_  | ~\new_[13372]_  | ~\new_[18657]_ ;
  assign \new_[10943]_  = (~\m2_data_i[17]  | ~\new_[16290]_ ) & (~\m1_data_i[17]  | ~\new_[18174]_ );
  assign \new_[10944]_  = ~\new_[16051]_  | ~\new_[17038]_  | ~\new_[13375]_  | ~\new_[14770]_ ;
  assign \new_[10945]_  = (~\m4_data_i[17]  | ~\new_[17272]_ ) & (~\m3_data_i[17]  | ~\new_[18927]_ );
  assign \new_[10946]_  = (~\m7_data_i[16]  | ~\new_[18096]_ ) & (~\m0_data_i[16]  | ~\new_[19575]_ );
  assign \new_[10947]_  = ~\new_[17707]_  | ~\new_[18553]_  | ~\new_[17706]_  | ~\new_[14634]_ ;
  assign \new_[10948]_  = (~\m4_data_i[16]  | ~\new_[17272]_ ) & (~\m3_data_i[16]  | ~\new_[18927]_ );
  assign \new_[10949]_  = (~\m7_data_i[15]  | ~\new_[16297]_ ) & (~\m0_data_i[15]  | ~\new_[18083]_ );
  assign \new_[10950]_  = (~\m4_data_i[15]  | ~\new_[17272]_ ) & (~\m3_data_i[15]  | ~\new_[17280]_ );
  assign \new_[10951]_  = (~\m7_data_i[14]  | ~\new_[16297]_ ) & (~\m0_data_i[14]  | ~\new_[18083]_ );
  assign \new_[10952]_  = (~\m4_data_i[14]  | ~\new_[17272]_ ) & (~\m3_data_i[14]  | ~\new_[18927]_ );
  assign \new_[10953]_  = (~\m4_data_i[13]  | ~\new_[17272]_ ) & (~\m3_data_i[13]  | ~\new_[17280]_ );
  assign \new_[10954]_  = (~\m7_sel_i[0]  | ~\new_[16296]_ ) & (~\m0_sel_i[0]  | ~\new_[18764]_ );
  assign \new_[10955]_  = (~\m4_data_i[12]  | ~\new_[17272]_ ) & (~\m3_data_i[12]  | ~\new_[17280]_ );
  assign \new_[10956]_  = (~\m4_data_i[11]  | ~\new_[17272]_ ) & (~\m3_data_i[11]  | ~\new_[18927]_ );
  assign \new_[10957]_  = (~\m7_data_i[10]  | ~\new_[16297]_ ) & (~\m0_data_i[10]  | ~\new_[19575]_ );
  assign \new_[10958]_  = (~\m2_data_i[9]  | ~\new_[16290]_ ) & (~\m1_data_i[9]  | ~\new_[19627]_ );
  assign \new_[10959]_  = (~\m5_addr_i[14]  | ~\new_[18759]_ ) & (~\m6_addr_i[14]  | ~\new_[17213]_ );
  assign \new_[10960]_  = (~\m4_data_i[8]  | ~\new_[17272]_ ) & (~\m3_data_i[8]  | ~\new_[17280]_ );
  assign \new_[10961]_  = (~\m4_data_i[7]  | ~\new_[17272]_ ) & (~\m3_data_i[7]  | ~\new_[17280]_ );
  assign \new_[10962]_  = (~\m7_data_i[7]  | ~\new_[18096]_ ) & (~\m0_data_i[7]  | ~\new_[19575]_ );
  assign \new_[10963]_  = (~\m2_data_i[6]  | ~\new_[16290]_ ) & (~\m1_data_i[6]  | ~\new_[18174]_ );
  assign \new_[10964]_  = (~\m4_data_i[6]  | ~\new_[17272]_ ) & (~\m3_data_i[6]  | ~\new_[17280]_ );
  assign \new_[10965]_  = ~\new_[16168]_  | ~\new_[17872]_  | ~\new_[14785]_  | ~\new_[17884]_ ;
  assign \new_[10966]_  = (~\m4_data_i[5]  | ~\new_[17272]_ ) & (~\m3_data_i[5]  | ~\new_[17280]_ );
  assign \new_[10967]_  = (~\m7_data_i[4]  | ~\new_[18096]_ ) & (~\m0_data_i[4]  | ~\new_[18083]_ );
  assign \new_[10968]_  = (~\m4_data_i[4]  | ~\new_[17272]_ ) & (~\m3_data_i[4]  | ~\new_[17280]_ );
  assign \new_[10969]_  = (~\m4_data_i[2]  | ~\new_[17272]_ ) & (~\m3_data_i[2]  | ~\new_[17280]_ );
  assign \new_[10970]_  = ~\new_[17113]_  | ~\new_[17057]_  | ~\new_[13337]_  | ~\new_[14795]_ ;
  assign \new_[10971]_  = (~\m7_data_i[0]  | ~\new_[16297]_ ) & (~\m0_data_i[0]  | ~\new_[18083]_ );
  assign \new_[10972]_  = (~\m2_data_i[31]  | ~\new_[14837]_ ) & (~\m1_data_i[31]  | ~\new_[18888]_ );
  assign \new_[10973]_  = (~\m4_data_i[0]  | ~\new_[17272]_ ) & (~\m3_data_i[0]  | ~\new_[18927]_ );
  assign \new_[10974]_  = ~\new_[17880]_  | ~\new_[17062]_  | ~\new_[16103]_  | ~\new_[14801]_ ;
  assign \new_[10975]_  = (~\new_[16297]_  | ~\new_[31496]_ ) & (~\new_[18083]_  | ~\m0_addr_i[31] );
  assign \new_[10976]_  = (~\new_[18070]_  | ~\m2_addr_i[31] ) & (~\new_[18173]_  | ~\new_[31447]_ );
  assign \new_[10977]_  = (~\new_[17272]_  | ~\m4_addr_i[31] ) & (~\new_[17280]_  | ~\m3_addr_i[31] );
  assign \new_[10978]_  = ~\new_[17883]_  | ~\new_[17882]_  | ~\new_[13308]_  | ~\new_[16204]_ ;
  assign \new_[10979]_  = (~\new_[16297]_  | ~\new_[31885]_ ) & (~\new_[18811]_  | ~\new_[31292]_ );
  assign \new_[10980]_  = (~\new_[18070]_  | ~\new_[31486]_ ) & (~\new_[18173]_  | ~\new_[31308]_ );
  assign \new_[10981]_  = (~\new_[17272]_  | ~\m4_addr_i[30] ) & (~\new_[17280]_  | ~\m3_addr_i[30] );
  assign \new_[10982]_  = (~\m2_data_i[30]  | ~\new_[14837]_ ) & (~\m1_data_i[30]  | ~\new_[18888]_ );
  assign \new_[10983]_  = (~\new_[16297]_  | ~\new_[31531]_ ) & (~\new_[18811]_  | ~\new_[31481]_ );
  assign \new_[10984]_  = (~\new_[18070]_  | ~\m2_addr_i[29] ) & (~\new_[19627]_  | ~\new_[31538]_ );
  assign \new_[10985]_  = (~\new_[17272]_  | ~\m4_addr_i[29] ) & (~\new_[17280]_  | ~\m3_addr_i[29] );
  assign \new_[10986]_  = (~\m2_data_i[29]  | ~\new_[17215]_ ) & (~\m1_data_i[29]  | ~\new_[20541]_ );
  assign \new_[10987]_  = (~\new_[16297]_  | ~\new_[30577]_ ) & (~\new_[18811]_  | ~\new_[30957]_ );
  assign \new_[10988]_  = (~\new_[16290]_  | ~\new_[31547]_ ) & (~\new_[19627]_  | ~\new_[31458]_ );
  assign \new_[10989]_  = (~\new_[17272]_  | ~\m4_addr_i[28] ) & (~\new_[17280]_  | ~\m3_addr_i[28] );
  assign \new_[10990]_  = (~\new_[16297]_  | ~\m7_addr_i[27] ) & (~\new_[18811]_  | ~\m0_addr_i[27] );
  assign \new_[10991]_  = (~\new_[14944]_  | ~\new_[29314]_ ) & (~\new_[14943]_  | ~\new_[29059]_ );
  assign \new_[10992]_  = (~\new_[18070]_  | ~\m2_addr_i[27] ) & (~\new_[19627]_  | ~\m1_addr_i[27] );
  assign \new_[10993]_  = (~\new_[17272]_  | ~\m4_addr_i[27] ) & (~\new_[17280]_  | ~\m3_addr_i[27] );
  assign \new_[10994]_  = ~\new_[16209]_  | ~\new_[17069]_  | ~\new_[16955]_  | ~\new_[16208]_ ;
  assign \new_[10995]_  = (~\new_[16297]_  | ~\m7_addr_i[26] ) & (~\new_[18811]_  | ~\m0_addr_i[26] );
  assign \new_[10996]_  = (~\new_[16290]_  | ~\m2_addr_i[26] ) & (~\new_[18173]_  | ~\m1_addr_i[26] );
  assign \new_[10997]_  = (~\new_[17272]_  | ~\m4_addr_i[26] ) & (~\new_[17280]_  | ~\m3_addr_i[26] );
  assign \new_[10998]_  = (~\m2_data_i[28]  | ~\new_[14837]_ ) & (~\m1_data_i[28]  | ~\new_[18888]_ );
  assign \new_[10999]_  = ~\new_[16211]_  | ~\new_[17885]_  | ~\new_[17080]_  | ~\new_[17081]_ ;
  assign \new_[11000]_  = (~\new_[16297]_  | ~\m7_addr_i[25] ) & (~\new_[18811]_  | ~\m0_addr_i[25] );
  assign \new_[11001]_  = ~\new_[16212]_  | ~\new_[17087]_  | ~\new_[17084]_  | ~\new_[17085]_ ;
  assign \new_[11002]_  = (~\new_[16290]_  | ~\m2_addr_i[25] ) & (~\new_[19627]_  | ~\m1_addr_i[25] );
  assign \new_[11003]_  = (~\new_[17272]_  | ~\m4_addr_i[25] ) & (~\new_[17280]_  | ~\m3_addr_i[25] );
  assign \new_[11004]_  = ~\new_[16224]_  | ~\new_[17893]_  | ~\new_[17088]_  | ~\new_[17106]_ ;
  assign \new_[11005]_  = ~\new_[16182]_  | ~\new_[17886]_  | ~\new_[16216]_  | ~\new_[18666]_ ;
  assign \new_[11006]_  = (~\new_[16297]_  | ~\m7_addr_i[24] ) & (~\new_[18811]_  | ~\m0_addr_i[24] );
  assign \new_[11007]_  = (~\new_[16290]_  | ~\m2_addr_i[24] ) & (~\new_[19627]_  | ~\m1_addr_i[24] );
  assign \new_[11008]_  = (~\new_[17272]_  | ~\m4_addr_i[24] ) & (~\new_[17280]_  | ~\m3_addr_i[24] );
  assign \new_[11009]_  = (~\m7_addr_i[23]  | ~\new_[16297]_ ) & (~\m0_addr_i[23]  | ~\new_[19575]_ );
  assign \new_[11010]_  = (~\m4_addr_i[23]  | ~\new_[17272]_ ) & (~\m3_addr_i[23]  | ~\new_[17280]_ );
  assign \new_[11011]_  = (~\new_[14946]_  | ~\new_[28396]_ ) & (~\new_[14945]_  | ~\new_[29345]_ );
  assign \new_[11012]_  = (~\m7_addr_i[22]  | ~\new_[16297]_ ) & (~\m0_addr_i[22]  | ~\new_[18811]_ );
  assign \new_[11013]_  = (~\m4_addr_i[22]  | ~\new_[17272]_ ) & (~\m3_addr_i[22]  | ~\new_[17280]_ );
  assign \new_[11014]_  = (~\m2_data_i[26]  | ~\new_[14837]_ ) & (~\m1_data_i[26]  | ~\new_[20541]_ );
  assign \new_[11015]_  = (~\m4_addr_i[21]  | ~\new_[17272]_ ) & (~\m3_addr_i[21]  | ~\new_[18927]_ );
  assign \new_[11016]_  = (~\m2_data_i[25]  | ~\new_[17215]_ ) & (~\m1_data_i[25]  | ~\new_[20541]_ );
  assign \new_[11017]_  = (~\m4_addr_i[20]  | ~\new_[17272]_ ) & (~\m3_addr_i[20]  | ~\new_[17279]_ );
  assign \new_[11018]_  = (~\m2_addr_i[0]  | ~\new_[17193]_ ) & (~\m1_addr_i[0]  | ~\new_[19633]_ );
  assign \new_[11019]_  = (~\m4_addr_i[19]  | ~\new_[17272]_ ) & (~\m3_addr_i[19]  | ~\new_[17279]_ );
  assign \new_[11020]_  = (~\m2_addr_i[18]  | ~\new_[18070]_ ) & (~\m1_addr_i[18]  | ~\new_[18172]_ );
  assign \new_[11021]_  = (~\m7_addr_i[18]  | ~\new_[16297]_ ) & (~\m0_addr_i[18]  | ~\new_[18083]_ );
  assign \new_[11022]_  = (~\m2_data_i[24]  | ~\new_[17215]_ ) & (~\m1_data_i[24]  | ~\new_[20541]_ );
  assign \new_[11023]_  = (~\m4_addr_i[18]  | ~\new_[17272]_ ) & (~\m3_addr_i[18]  | ~\new_[17280]_ );
  assign \new_[11024]_  = (~\m2_addr_i[17]  | ~\new_[16290]_ ) & (~\m1_addr_i[17]  | ~\new_[19627]_ );
  assign \new_[11025]_  = (~\m4_addr_i[17]  | ~\new_[17272]_ ) & (~\m3_addr_i[17]  | ~\new_[17279]_ );
  assign \new_[11026]_  = (~\m2_data_i[23]  | ~\new_[17215]_ ) & (~\m1_data_i[23]  | ~\new_[20541]_ );
  assign \new_[11027]_  = (~\m7_addr_i[16]  | ~\new_[16297]_ ) & (~\m0_addr_i[16]  | ~\new_[18083]_ );
  assign \new_[11028]_  = (~\m4_addr_i[16]  | ~\new_[17272]_ ) & (~\m3_addr_i[16]  | ~\new_[17279]_ );
  assign \new_[11029]_  = (~\m4_addr_i[15]  | ~\new_[17272]_ ) & (~\m3_addr_i[15]  | ~\new_[17280]_ );
  assign \new_[11030]_  = (~\m7_addr_i[15]  | ~\new_[16297]_ ) & (~\m0_addr_i[15]  | ~\new_[19575]_ );
  assign \new_[11031]_  = (~\m2_data_i[22]  | ~\new_[17215]_ ) & (~\m1_data_i[22]  | ~\new_[20541]_ );
  assign \new_[11032]_  = (~\m4_addr_i[14]  | ~\new_[17272]_ ) & (~\m3_addr_i[14]  | ~\new_[17278]_ );
  assign \new_[11033]_  = (~\m7_addr_i[14]  | ~\new_[16297]_ ) & (~\m0_addr_i[14]  | ~\new_[18083]_ );
  assign \new_[11034]_  = (~\m7_addr_i[13]  | ~\new_[16297]_ ) & (~\m0_addr_i[13]  | ~\new_[19575]_ );
  assign \new_[11035]_  = (~\m4_addr_i[13]  | ~\new_[17272]_ ) & (~\m3_addr_i[13]  | ~\new_[17278]_ );
  assign \new_[11036]_  = (~\m7_addr_i[12]  | ~\new_[16297]_ ) & (~\m0_addr_i[12]  | ~\new_[18083]_ );
  assign \new_[11037]_  = (~\m4_addr_i[12]  | ~\new_[17272]_ ) & (~\m3_addr_i[12]  | ~\new_[18927]_ );
  assign \new_[11038]_  = (~\m2_data_i[21]  | ~\new_[17215]_ ) & (~\m1_data_i[21]  | ~\new_[19618]_ );
  assign \new_[11039]_  = (~\m4_addr_i[11]  | ~\new_[17272]_ ) & (~\m3_addr_i[11]  | ~\new_[17279]_ );
  assign \new_[11040]_  = (~\m4_addr_i[10]  | ~\new_[17272]_ ) & (~\m3_addr_i[10]  | ~\new_[17278]_ );
  assign \new_[11041]_  = (~\m7_addr_i[10]  | ~\new_[16297]_ ) & (~\m0_addr_i[10]  | ~\new_[19575]_ );
  assign \new_[11042]_  = (~\m2_data_i[20]  | ~\new_[17215]_ ) & (~\m1_data_i[20]  | ~\new_[19619]_ );
  assign \new_[11043]_  = (~\m2_addr_i[9]  | ~\new_[16290]_ ) & (~\m1_addr_i[9]  | ~\new_[19627]_ );
  assign \new_[11044]_  = (~\m4_addr_i[9]  | ~\new_[17272]_ ) & (~\m3_addr_i[9]  | ~\new_[17280]_ );
  assign \new_[11045]_  = (~\m2_data_i[19]  | ~\new_[14837]_ ) & (~\m1_data_i[19]  | ~\new_[19618]_ );
  assign \new_[11046]_  = (~\m2_addr_i[8]  | ~\new_[16290]_ ) & (~\m1_addr_i[8]  | ~\new_[19627]_ );
  assign \new_[11047]_  = (~\m4_addr_i[8]  | ~\new_[17272]_ ) & (~\m3_addr_i[8]  | ~\new_[17280]_ );
  assign \new_[11048]_  = (~\m2_addr_i[7]  | ~\new_[16290]_ ) & (~\m1_addr_i[7]  | ~\new_[18174]_ );
  assign \new_[11049]_  = (~\m4_addr_i[7]  | ~\new_[17272]_ ) & (~\m3_addr_i[7]  | ~\new_[17278]_ );
  assign \new_[11050]_  = (~\m2_data_i[18]  | ~\new_[17216]_ ) & (~\m1_data_i[18]  | ~\new_[18888]_ );
  assign \new_[11051]_  = (~\m4_addr_i[6]  | ~\new_[17272]_ ) & (~\m3_addr_i[6]  | ~\new_[17279]_ );
  assign \new_[11052]_  = (~\new_[14953]_  | ~\new_[27738]_ ) & (~\new_[14952]_  | ~\new_[28112]_ );
  assign \new_[11053]_  = (~\m2_data_i[17]  | ~\new_[17215]_ ) & (~\m1_data_i[17]  | ~\new_[20541]_ );
  assign \new_[11054]_  = (~\m4_addr_i[4]  | ~\new_[17272]_ ) & (~\m3_addr_i[4]  | ~\new_[17280]_ );
  assign \new_[11055]_  = (~\m7_addr_i[4]  | ~\new_[18096]_ ) & (~\m0_addr_i[4]  | ~\new_[18083]_ );
  assign \new_[11056]_  = ~\new_[13215]_  & (~\new_[14830]_  | ~\m7_addr_i[26] );
  assign \new_[11057]_  = (~\m4_addr_i[3]  | ~\new_[17272]_ ) & (~\m3_addr_i[3]  | ~\new_[17280]_ );
  assign \new_[11058]_  = (~\m4_addr_i[2]  | ~\new_[17272]_ ) & (~\m3_addr_i[2]  | ~\new_[17280]_ );
  assign \new_[11059]_  = (~\m2_data_i[16]  | ~\new_[17216]_ ) & (~\m1_data_i[16]  | ~\new_[20541]_ );
  assign \new_[11060]_  = (~\m7_addr_i[2]  | ~\new_[18096]_ ) & (~\m0_addr_i[2]  | ~\new_[18083]_ );
  assign \new_[11061]_  = (~\m2_addr_i[1]  | ~\new_[16290]_ ) & (~\m1_addr_i[1]  | ~\new_[18174]_ );
  assign \new_[11062]_  = (~\m4_addr_i[1]  | ~\new_[17272]_ ) & (~\m3_addr_i[1]  | ~\new_[18927]_ );
  assign \new_[11063]_  = (~\m2_data_i[15]  | ~\new_[17216]_ ) & (~\m1_data_i[15]  | ~\new_[19619]_ );
  assign \new_[11064]_  = (~\m7_addr_i[0]  | ~\new_[16297]_ ) & (~\m0_addr_i[0]  | ~\new_[19575]_ );
  assign \new_[11065]_  = (~\m2_addr_i[0]  | ~\new_[16290]_ ) & (~\m1_addr_i[0]  | ~\new_[18174]_ );
  assign \new_[11066]_  = (~\m4_addr_i[0]  | ~\new_[17272]_ ) & (~\m3_addr_i[0]  | ~\new_[18927]_ );
  assign \new_[11067]_  = (~\m7_sel_i[3]  | ~\new_[16297]_ ) & (~\m0_sel_i[3]  | ~\new_[19575]_ );
  assign \new_[11068]_  = (~\m4_sel_i[3]  | ~\new_[17272]_ ) & (~\m3_sel_i[3]  | ~\new_[17280]_ );
  assign \new_[11069]_  = (~\m7_sel_i[2]  | ~\new_[16297]_ ) & (~\m0_sel_i[2]  | ~\new_[18083]_ );
  assign \new_[11070]_  = (~\m2_data_i[14]  | ~\new_[17216]_ ) & (~\m1_data_i[14]  | ~\new_[19619]_ );
  assign \new_[11071]_  = (~\m4_sel_i[2]  | ~\new_[17272]_ ) & (~\m3_sel_i[2]  | ~\new_[17280]_ );
  assign \new_[11072]_  = (~\m4_sel_i[1]  | ~\new_[17272]_ ) & (~\m3_sel_i[1]  | ~\new_[17279]_ );
  assign \new_[11073]_  = (~\m2_sel_i[0]  | ~\new_[16290]_ ) & (~\m1_sel_i[0]  | ~\new_[19627]_ );
  assign \new_[11074]_  = (~\m4_sel_i[0]  | ~\new_[17272]_ ) & (~\m3_sel_i[0]  | ~\new_[17280]_ );
  assign \new_[11075]_  = (~\m2_data_i[13]  | ~\new_[17216]_ ) & (~\m1_data_i[13]  | ~\new_[18888]_ );
  assign \new_[11076]_  = (~m7_we_i | ~\new_[16297]_ ) & (~m0_we_i | ~\new_[18083]_ );
  assign \new_[11077]_  = (~m4_we_i | ~\new_[17272]_ ) & (~m3_we_i | ~\new_[18927]_ );
  assign \new_[11078]_  = (~\m2_data_i[11]  | ~\new_[17216]_ ) & (~\m1_data_i[11]  | ~\new_[19618]_ );
  assign \new_[11079]_  = (~\m5_addr_i[5]  | ~\new_[18004]_ ) & (~\m6_addr_i[5]  | ~\new_[17241]_ );
  assign \new_[11080]_  = (~\m2_data_i[10]  | ~\new_[17216]_ ) & (~\m1_data_i[10]  | ~\new_[18888]_ );
  assign \new_[11081]_  = (~\m5_data_i[26]  | ~\new_[18738]_ ) & (~\m6_data_i[26]  | ~\new_[18030]_ );
  assign \new_[11082]_  = \new_[13250]_  & \new_[14633]_ ;
  assign \new_[11083]_  = \new_[13257]_  & \new_[13258]_ ;
  assign \new_[11084]_  = \new_[16064]_  & \new_[13265]_ ;
  assign \new_[11085]_  = \new_[16072]_  & \new_[13271]_ ;
  assign \new_[11086]_  = (~\m2_data_i[3]  | ~\new_[17216]_ ) & (~\m1_data_i[3]  | ~\new_[18888]_ );
  assign \new_[11087]_  = \new_[13386]_  & \new_[13410]_ ;
  assign \new_[11088]_  = \new_[13388]_  & \new_[13390]_ ;
  assign \new_[11089]_  = \new_[13401]_  & \new_[13399]_ ;
  assign \new_[11090]_  = (~\m2_data_i[1]  | ~\new_[17216]_ ) & (~\m1_data_i[1]  | ~\new_[19619]_ );
  assign \new_[11091]_  = (~\m2_data_i[0]  | ~\new_[17216]_ ) & (~\m1_data_i[0]  | ~\new_[19618]_ );
  assign \new_[11092]_  = (~\new_[17215]_  | ~\m2_addr_i[31] ) & (~\new_[20541]_  | ~\new_[31447]_ );
  assign \new_[11093]_  = (~\new_[17215]_  | ~\new_[31486]_ ) & (~\new_[20541]_  | ~\new_[31308]_ );
  assign \new_[11094]_  = (~\new_[17215]_  | ~\new_[31000]_ ) & (~\new_[20541]_  | ~\new_[31538]_ );
  assign \new_[11095]_  = (~\m5_addr_i[9]  | ~\new_[18004]_ ) & (~\m6_addr_i[9]  | ~\new_[17241]_ );
  assign \new_[11096]_  = (~\new_[17215]_  | ~\new_[31547]_ ) & (~\new_[20541]_  | ~\new_[31458]_ );
  assign \new_[11097]_  = (~\m7_addr_i[0]  | ~\new_[16296]_ ) & (~\m0_addr_i[0]  | ~\new_[18764]_ );
  assign \new_[11098]_  = (~\new_[17215]_  | ~\m2_addr_i[27] ) & (~\new_[20541]_  | ~\m1_addr_i[27] );
  assign \new_[11099]_  = (~\new_[17215]_  | ~\m2_addr_i[26] ) & (~\new_[20541]_  | ~\m1_addr_i[26] );
  assign \new_[11100]_  = ~m4_stb_i | ~\new_[26164]_  | ~\new_[17271]_ ;
  assign \new_[11101]_  = ~m7_stb_i | ~\new_[25155]_  | ~\new_[17239]_ ;
  assign \new_[11102]_  = (~\new_[17215]_  | ~\m2_addr_i[25] ) & (~\new_[20541]_  | ~\m1_addr_i[25] );
  assign \new_[11103]_  = ~\new_[13504]_  | ~\new_[13535]_ ;
  assign \new_[11104]_  = ~\new_[13407]_  & ~\new_[13409]_ ;
  assign \new_[11105]_  = (~\new_[17215]_  | ~\m2_addr_i[24] ) & (~\new_[20541]_  | ~\m1_addr_i[24] );
  assign \new_[11106]_  = ~\new_[13411]_  & (~\new_[30700]_  | ~\new_[32348]_ );
  assign \new_[11107]_  = ~\new_[13508]_  | ~\new_[13536]_ ;
  assign \new_[11108]_  = (~\m2_addr_i[23]  | ~\new_[17215]_ ) & (~\m1_addr_i[23]  | ~\new_[20541]_ );
  assign \new_[11109]_  = (~\m2_addr_i[22]  | ~\new_[17216]_ ) & (~\m1_addr_i[22]  | ~\new_[19619]_ );
  assign \new_[11110]_  = (~\m2_addr_i[21]  | ~\new_[17215]_ ) & (~\m1_addr_i[21]  | ~\new_[19619]_ );
  assign \new_[11111]_  = (~\m2_addr_i[20]  | ~\new_[17215]_ ) & (~\m1_addr_i[20]  | ~\new_[20541]_ );
  assign \new_[11112]_  = (~\new_[17260]_  | ~\m4_addr_i[25] ) & (~\new_[18175]_  | ~\m3_addr_i[25] );
  assign \new_[11113]_  = ~\new_[13212]_  & (~\new_[14839]_  | ~\m3_addr_i[27] );
  assign \new_[11114]_  = (~\m2_addr_i[19]  | ~\new_[17215]_ ) & (~\m1_addr_i[19]  | ~\new_[19619]_ );
  assign \new_[11115]_  = (~\m2_addr_i[18]  | ~\new_[17215]_ ) & (~\m1_addr_i[18]  | ~\new_[19619]_ );
  assign \new_[11116]_  = (~\m2_addr_i[17]  | ~\new_[14837]_ ) & (~\m1_addr_i[17]  | ~\new_[19619]_ );
  assign \new_[11117]_  = (~\m2_addr_i[16]  | ~\new_[17215]_ ) & (~\m1_addr_i[16]  | ~\new_[19619]_ );
  assign \new_[11118]_  = (~\m2_addr_i[15]  | ~\new_[14837]_ ) & (~\m1_addr_i[15]  | ~\new_[19619]_ );
  assign \new_[11119]_  = (~\m2_addr_i[14]  | ~\new_[17215]_ ) & (~\m1_addr_i[14]  | ~\new_[19619]_ );
  assign \new_[11120]_  = (~\m2_addr_i[13]  | ~\new_[17215]_ ) & (~\m1_addr_i[13]  | ~\new_[19619]_ );
  assign \new_[11121]_  = (~\m5_data_i[12]  | ~\new_[18750]_ ) & (~\m6_data_i[12]  | ~\new_[17213]_ );
  assign \new_[11122]_  = ~\new_[13236]_  & (~\new_[27535]_  | ~\new_[16322]_ );
  assign \new_[11123]_  = (~\m2_addr_i[12]  | ~\new_[17215]_ ) & (~\m1_addr_i[12]  | ~\new_[19619]_ );
  assign \new_[11124]_  = (~\m2_addr_i[11]  | ~\new_[17215]_ ) & (~\m1_addr_i[11]  | ~\new_[20541]_ );
  assign \new_[11125]_  = ~\new_[13245]_  & (~\new_[30483]_  | ~\new_[17327]_ );
  assign \new_[11126]_  = (~\m2_addr_i[10]  | ~\new_[17215]_ ) & (~\m1_addr_i[10]  | ~\new_[20541]_ );
  assign \new_[11127]_  = (~\m2_addr_i[9]  | ~\new_[17215]_ ) & (~\m1_addr_i[9]  | ~\new_[19618]_ );
  assign \new_[11128]_  = (~\m2_addr_i[8]  | ~\new_[14837]_ ) & (~\m1_addr_i[8]  | ~\new_[19619]_ );
  assign \new_[11129]_  = (~\m2_addr_i[7]  | ~\new_[17216]_ ) & (~\m1_addr_i[7]  | ~\new_[19619]_ );
  assign \new_[11130]_  = (~\m2_data_i[29]  | ~\new_[17218]_ ) & (~\m1_data_i[29]  | ~\new_[18905]_ );
  assign \new_[11131]_  = (~\m2_addr_i[6]  | ~\new_[17215]_ ) & (~\m1_addr_i[6]  | ~\new_[19619]_ );
  assign \new_[11132]_  = ~\new_[13275]_  & (~\new_[27270]_  | ~\new_[14895]_ );
  assign \new_[11133]_  = (~\new_[31399]_  | ~\new_[17216]_ ) & (~\m1_addr_i[3]  | ~\new_[19618]_ );
  assign \new_[11134]_  = (~\m2_addr_i[1]  | ~\new_[17215]_ ) & (~\m1_addr_i[1]  | ~\new_[20541]_ );
  assign \new_[11135]_  = (~\m2_addr_i[0]  | ~\new_[17216]_ ) & (~\m1_addr_i[0]  | ~\new_[19619]_ );
  assign \new_[11136]_  = (~\m2_sel_i[3]  | ~\new_[17215]_ ) & (~\m1_sel_i[3]  | ~\new_[19619]_ );
  assign \new_[11137]_  = (~\m2_sel_i[2]  | ~\new_[17216]_ ) & (~\m1_sel_i[2]  | ~\new_[19619]_ );
  assign \new_[11138]_  = ~\new_[13367]_  & (~\new_[16301]_  | ~\new_[30672]_ );
  assign \new_[11139]_  = (~\m2_sel_i[1]  | ~\new_[17215]_ ) & (~\m1_sel_i[1]  | ~\new_[19619]_ );
  assign \new_[11140]_  = (~\m2_sel_i[0]  | ~\new_[17216]_ ) & (~\m1_sel_i[0]  | ~\new_[20541]_ );
  assign \new_[11141]_  = ~\new_[29453]_  & (~\new_[14928]_  | ~\new_[28530]_ );
  assign \new_[11142]_  = (~\m2_data_i[31]  | ~\new_[17193]_ ) & (~\m1_data_i[31]  | ~\new_[18917]_ );
  assign \new_[11143]_  = ~\new_[14687]_  & ~\new_[13404]_ ;
  assign \new_[11144]_  = (~\m2_data_i[30]  | ~\new_[17193]_ ) & (~\m1_data_i[30]  | ~\new_[18917]_ );
  assign \new_[11145]_  = (~\m4_data_i[30]  | ~\new_[17260]_ ) & (~\m3_data_i[30]  | ~\new_[18175]_ );
  assign \new_[11146]_  = ~\new_[13293]_  & (~\new_[14895]_  | ~\new_[29153]_ );
  assign \new_[11147]_  = (~\m2_data_i[29]  | ~\new_[17193]_ ) & (~\m1_data_i[29]  | ~\new_[18917]_ );
  assign \new_[11148]_  = (~\m4_data_i[29]  | ~\new_[17260]_ ) & (~\m3_data_i[29]  | ~\new_[18175]_ );
  assign \new_[11149]_  = (~\m2_data_i[28]  | ~\new_[17193]_ ) & (~\m1_data_i[28]  | ~\new_[18916]_ );
  assign \new_[11150]_  = (~\m2_data_i[27]  | ~\new_[17193]_ ) & (~\m1_data_i[27]  | ~\new_[19633]_ );
  assign \new_[11151]_  = (~\m2_data_i[26]  | ~\new_[17193]_ ) & (~\m1_data_i[26]  | ~\new_[18917]_ );
  assign \new_[11152]_  = (~\m2_data_i[25]  | ~\new_[17193]_ ) & (~\m1_data_i[25]  | ~\new_[18917]_ );
  assign \new_[11153]_  = (~\m2_data_i[24]  | ~\new_[17193]_ ) & (~\m1_data_i[24]  | ~\new_[19633]_ );
  assign \new_[11154]_  = ~\new_[14588]_  & (~\new_[14880]_  | ~\m4_addr_i[27] );
  assign \new_[11155]_  = ~\new_[13283]_  & (~\new_[16323]_  | ~\new_[31935]_ );
  assign \new_[11156]_  = (~\m2_data_i[23]  | ~\new_[17193]_ ) & (~\m1_data_i[23]  | ~\new_[18916]_ );
  assign \new_[11157]_  = (~\m2_data_i[22]  | ~\new_[17193]_ ) & (~\m1_data_i[22]  | ~\new_[19633]_ );
  assign \new_[11158]_  = (~\m7_data_i[21]  | ~\new_[18116]_ ) & (~\m0_data_i[21]  | ~\new_[19637]_ );
  assign \new_[11159]_  = (~\m7_data_i[20]  | ~\new_[18116]_ ) & (~\m0_data_i[20]  | ~\new_[19637]_ );
  assign \new_[11160]_  = (~\m4_data_i[20]  | ~\new_[17260]_ ) & (~\m3_data_i[20]  | ~\new_[18175]_ );
  assign \new_[11161]_  = (~\m7_data_i[19]  | ~\new_[18115]_ ) & (~\m0_data_i[19]  | ~\new_[19637]_ );
  assign \new_[11162]_  = (~\m7_sel_i[3]  | ~\new_[17232]_ ) & (~\m0_sel_i[3]  | ~\new_[20580]_ );
  assign \new_[11163]_  = (~\m7_addr_i[23]  | ~\new_[17232]_ ) & (~\m0_addr_i[23]  | ~\new_[20580]_ );
  assign \new_[11164]_  = (~\m7_data_i[17]  | ~\new_[18115]_ ) & (~\m0_data_i[17]  | ~\new_[18932]_ );
  assign \new_[11165]_  = (~\m7_data_i[16]  | ~\new_[18115]_ ) & (~\m0_data_i[16]  | ~\new_[18932]_ );
  assign \new_[11166]_  = (~\m7_data_i[15]  | ~\new_[18115]_ ) & (~\m0_data_i[15]  | ~\new_[18932]_ );
  assign \new_[11167]_  = (~\m7_data_i[11]  | ~\new_[18115]_ ) & (~\m0_data_i[11]  | ~\new_[18932]_ );
  assign \new_[11168]_  = (~\m5_addr_i[0]  | ~\new_[18016]_ ) & (~\m6_addr_i[0]  | ~\new_[17229]_ );
  assign \new_[11169]_  = (~\m7_data_i[8]  | ~\new_[18115]_ ) & (~\m0_data_i[8]  | ~\new_[18932]_ );
  assign \new_[11170]_  = (~\m7_data_i[7]  | ~\new_[18115]_ ) & (~\m0_data_i[7]  | ~\new_[18932]_ );
  assign \new_[11171]_  = (~\m7_data_i[6]  | ~\new_[18115]_ ) & (~\m0_data_i[6]  | ~\new_[18932]_ );
  assign \new_[11172]_  = (~\m7_data_i[5]  | ~\new_[18115]_ ) & (~\m0_data_i[5]  | ~\new_[18932]_ );
  assign \new_[11173]_  = (~\m5_addr_i[9]  | ~\new_[17202]_ ) & (~\m4_addr_i[9]  | ~\new_[17270]_ );
  assign \new_[11174]_  = (~\m4_addr_i[14]  | ~\new_[18149]_ ) & (~\m3_addr_i[14]  | ~\new_[18928]_ );
  assign \new_[11175]_  = (~\m7_data_i[3]  | ~\new_[18115]_ ) & (~\m0_data_i[3]  | ~\new_[18932]_ );
  assign \new_[11176]_  = (~\m7_data_i[0]  | ~\new_[18115]_ ) & (~\m0_data_i[0]  | ~\new_[18932]_ );
  assign \new_[11177]_  = (~\new_[17193]_  | ~\m2_addr_i[31] ) & (~\new_[18193]_  | ~\new_[31447]_ );
  assign \new_[11178]_  = (~\new_[17260]_  | ~\m4_addr_i[31] ) & (~\new_[18175]_  | ~\m3_addr_i[31] );
  assign \new_[11179]_  = (~\new_[17193]_  | ~\new_[31486]_ ) & (~\new_[18193]_  | ~\new_[31308]_ );
  assign \new_[11180]_  = (~\new_[17260]_  | ~\m4_addr_i[30] ) & (~\new_[18175]_  | ~\m3_addr_i[30] );
  assign \new_[11181]_  = (~\new_[17193]_  | ~\new_[31000]_ ) & (~\new_[18193]_  | ~\new_[31538]_ );
  assign \new_[11182]_  = (~\new_[17260]_  | ~\m4_addr_i[29] ) & (~\new_[18175]_  | ~\m3_addr_i[29] );
  assign \new_[11183]_  = (~\m7_addr_i[23]  | ~\new_[19584]_ ) & (~\m0_addr_i[23]  | ~\new_[18026]_ );
  assign \new_[11184]_  = (~\new_[17193]_  | ~\new_[31547]_ ) & (~\new_[18193]_  | ~\new_[31458]_ );
  assign \new_[11185]_  = (~\m2_data_i[15]  | ~\new_[18067]_ ) & (~\m1_data_i[15]  | ~\new_[20573]_ );
  assign \new_[11186]_  = (~\new_[17193]_  | ~\m2_addr_i[27] ) & (~\new_[18193]_  | ~\m1_addr_i[27] );
  assign \new_[11187]_  = (~\new_[17193]_  | ~\m2_addr_i[26] ) & (~\new_[18193]_  | ~\m1_addr_i[26] );
  assign \new_[11188]_  = (~\new_[17193]_  | ~\m2_addr_i[24] ) & (~\new_[18193]_  | ~\m1_addr_i[24] );
  assign \new_[11189]_  = (~\m2_data_i[21]  | ~\new_[18077]_ ) & (~\m1_data_i[21]  | ~\new_[18182]_ );
  assign \new_[11190]_  = (~\m7_data_i[22]  | ~\new_[18106]_ ) & (~\m0_data_i[22]  | ~\new_[18026]_ );
  assign \new_[11191]_  = (~\new_[18101]_  | ~\m7_addr_i[24] ) & (~\new_[18026]_  | ~\m0_addr_i[24] );
  assign \new_[11192]_  = (~\m7_addr_i[23]  | ~\new_[18115]_ ) & (~\m0_addr_i[23]  | ~\new_[18932]_ );
  assign \new_[11193]_  = (~\m7_data_i[17]  | ~\new_[18109]_ ) & (~\m0_data_i[17]  | ~\new_[18026]_ );
  assign \new_[11194]_  = (~\m7_data_i[18]  | ~\new_[18109]_ ) & (~\m0_data_i[18]  | ~\new_[18026]_ );
  assign \new_[11195]_  = (~\m2_addr_i[22]  | ~\new_[18077]_ ) & (~\m1_addr_i[22]  | ~\new_[18182]_ );
  assign \new_[11196]_  = (~\m7_data_i[26]  | ~\new_[18102]_ ) & (~\m0_data_i[26]  | ~\new_[18026]_ );
  assign \new_[11197]_  = (~\m2_data_i[22]  | ~\new_[18078]_ ) & (~\m1_data_i[22]  | ~\new_[19632]_ );
  assign \new_[11198]_  = (~\m7_addr_i[22]  | ~\new_[18115]_ ) & (~\m0_addr_i[22]  | ~\new_[18932]_ );
  assign \new_[11199]_  = (~\m7_addr_i[22]  | ~\new_[18103]_ ) & (~\m0_addr_i[22]  | ~\new_[18026]_ );
  assign \new_[11200]_  = (~\m7_addr_i[21]  | ~\new_[18116]_ ) & (~\m0_addr_i[21]  | ~\new_[18932]_ );
  assign \new_[11201]_  = (~\new_[17213]_  | ~\m6_addr_i[25] ) & (~\new_[20544]_  | ~\m5_addr_i[25] );
  assign \new_[11202]_  = (~\m5_addr_i[23]  | ~\new_[20544]_ ) & (~\m6_addr_i[23]  | ~\new_[17213]_ );
  assign \new_[11203]_  = (~\m7_addr_i[20]  | ~\new_[18116]_ ) & (~\m0_addr_i[20]  | ~\new_[19637]_ );
  assign \new_[11204]_  = (~\m7_addr_i[19]  | ~\new_[18115]_ ) & (~\m0_addr_i[19]  | ~\new_[19637]_ );
  assign \new_[11205]_  = (~\m7_addr_i[18]  | ~\new_[18115]_ ) & (~\m0_addr_i[18]  | ~\new_[18932]_ );
  assign \new_[11206]_  = (~\m5_addr_i[21]  | ~\new_[20544]_ ) & (~\m6_addr_i[21]  | ~\new_[18787]_ );
  assign \new_[11207]_  = (~\m7_addr_i[16]  | ~\new_[18116]_ ) & (~\m0_addr_i[16]  | ~\new_[18932]_ );
  assign \new_[11208]_  = (~\m7_data_i[15]  | ~\new_[18110]_ ) & (~\m0_data_i[15]  | ~\new_[18026]_ );
  assign \new_[11209]_  = (~\m7_addr_i[14]  | ~\new_[17240]_ ) & (~\m6_addr_i[14]  | ~\new_[18089]_ );
  assign \new_[11210]_  = (~\m7_addr_i[15]  | ~\new_[18116]_ ) & (~\m0_addr_i[15]  | ~\new_[18932]_ );
  assign \new_[11211]_  = (~\m2_data_i[19]  | ~\new_[18077]_ ) & (~\m1_data_i[19]  | ~\new_[18183]_ );
  assign \new_[11212]_  = (~\new_[18067]_  | ~\m2_addr_i[29] ) & (~\new_[19626]_  | ~\new_[31538]_ );
  assign \new_[11213]_  = (~\m2_addr_i[11]  | ~\new_[18077]_ ) & (~\m1_addr_i[11]  | ~\new_[19632]_ );
  assign \new_[11214]_  = (~\m7_data_i[0]  | ~\new_[19584]_ ) & (~\m0_data_i[0]  | ~\new_[18026]_ );
  assign \new_[11215]_  = (~\m7_addr_i[14]  | ~\new_[18116]_ ) & (~\m0_addr_i[14]  | ~\new_[19637]_ );
  assign \new_[11216]_  = (~\m7_addr_i[13]  | ~\new_[18116]_ ) & (~\m0_addr_i[13]  | ~\new_[19637]_ );
  assign \new_[11217]_  = (~\m7_data_i[19]  | ~\new_[18105]_ ) & (~\m0_data_i[19]  | ~\new_[18026]_ );
  assign \new_[11218]_  = (~\m2_data_i[27]  | ~\new_[18077]_ ) & (~\m1_data_i[27]  | ~\new_[18183]_ );
  assign \new_[11219]_  = (~\m7_addr_i[12]  | ~\new_[18116]_ ) & (~\m0_addr_i[12]  | ~\new_[18932]_ );
  assign \new_[11220]_  = (~\m5_data_i[20]  | ~\new_[18753]_ ) & (~\m6_data_i[20]  | ~\new_[17213]_ );
  assign \new_[11221]_  = (~\m7_addr_i[21]  | ~\new_[18100]_ ) & (~\m0_addr_i[21]  | ~\new_[18026]_ );
  assign \new_[11222]_  = (~\m7_addr_i[11]  | ~\new_[18116]_ ) & (~\m0_addr_i[11]  | ~\new_[18932]_ );
  assign \new_[11223]_  = (~\m7_addr_i[10]  | ~\new_[18116]_ ) & (~\m0_addr_i[10]  | ~\new_[19637]_ );
  assign \new_[11224]_  = (~\m2_data_i[20]  | ~\new_[18077]_ ) & (~\m1_data_i[20]  | ~\new_[18183]_ );
  assign \new_[11225]_  = (~\m2_addr_i[19]  | ~\new_[18077]_ ) & (~\m1_addr_i[19]  | ~\new_[19632]_ );
  assign \new_[11226]_  = (~\m2_addr_i[21]  | ~\new_[18077]_ ) & (~\m1_addr_i[21]  | ~\new_[18181]_ );
  assign \new_[11227]_  = (~\m7_addr_i[9]  | ~\new_[18115]_ ) & (~\m0_addr_i[9]  | ~\new_[18932]_ );
  assign \new_[11228]_  = (~\m7_addr_i[8]  | ~\new_[18116]_ ) & (~\m0_addr_i[8]  | ~\new_[18932]_ );
  assign \new_[11229]_  = (~\m5_data_i[10]  | ~\new_[18015]_ ) & (~\m6_data_i[10]  | ~\new_[17229]_ );
  assign \new_[11230]_  = (~\m7_data_i[20]  | ~\new_[18105]_ ) & (~\m0_data_i[20]  | ~\new_[18026]_ );
  assign \new_[11231]_  = (~\m3_addr_i[14]  | ~\new_[32350]_ ) & (~\m2_addr_i[14]  | ~\new_[17223]_ );
  assign \new_[11232]_  = (~\new_[18098]_  | ~\m7_addr_i[31] ) & (~\new_[18026]_  | ~\m0_addr_i[31] );
  assign \new_[11233]_  = (~\m2_data_i[23]  | ~\new_[18078]_ ) & (~\m1_data_i[23]  | ~\new_[19632]_ );
  assign \new_[11234]_  = (~\new_[18098]_  | ~\new_[31885]_ ) & (~\new_[18026]_  | ~\new_[31292]_ );
  assign \new_[11235]_  = (~\m7_addr_i[7]  | ~\new_[18115]_ ) & (~\m0_addr_i[7]  | ~\new_[18932]_ );
  assign \new_[11236]_  = \new_[5988]_  ? \new_[29681]_  : \new_[16320]_ ;
  assign \new_[11237]_  = \new_[6189]_  ? \new_[29505]_  : \new_[16315]_ ;
  assign \new_[11238]_  = (~\m5_data_i[29]  | ~\new_[18749]_ ) & (~\m6_data_i[29]  | ~\new_[17213]_ );
  assign \new_[11239]_  = (~\m7_data_i[27]  | ~\new_[18105]_ ) & (~\m0_data_i[27]  | ~\new_[18026]_ );
  assign \new_[11240]_  = (~\m5_data_i[27]  | ~\new_[18747]_ ) & (~\m6_data_i[27]  | ~\new_[18787]_ );
  assign \new_[11241]_  = (~\m5_data_i[26]  | ~\new_[18754]_ ) & (~\m6_data_i[26]  | ~\new_[17213]_ );
  assign \new_[11242]_  = (~\new_[17213]_  | ~\m6_addr_i[24] ) & (~\new_[20544]_  | ~\m5_addr_i[24] );
  assign \new_[11243]_  = (~\m5_data_i[25]  | ~\new_[18754]_ ) & (~\m6_data_i[25]  | ~\new_[17213]_ );
  assign \new_[11244]_  = (~\m2_addr_i[20]  | ~\new_[18077]_ ) & (~\m1_addr_i[20]  | ~\new_[18189]_ );
  assign \new_[11245]_  = (~\m5_data_i[15]  | ~\new_[18758]_ ) & (~\m6_data_i[15]  | ~\new_[17213]_ );
  assign \new_[11246]_  = (~\m2_data_i[13]  | ~\new_[18077]_ ) & (~\m1_data_i[13]  | ~\new_[18186]_ );
  assign \new_[11247]_  = (~\m2_data_i[12]  | ~\new_[18077]_ ) & (~\m1_data_i[12]  | ~\new_[18186]_ );
  assign \new_[11248]_  = (~\m2_addr_i[17]  | ~\new_[18077]_ ) & (~\m1_addr_i[17]  | ~\new_[19632]_ );
  assign \new_[11249]_  = (~\m2_data_i[8]  | ~\new_[18077]_ ) & (~\m1_data_i[8]  | ~\new_[18190]_ );
  assign \new_[11250]_  = (~\m5_addr_i[16]  | ~\new_[18747]_ ) & (~\m6_addr_i[16]  | ~\new_[17213]_ );
  assign \new_[11251]_  = (~\m7_addr_i[12]  | ~\new_[19584]_ ) & (~\m0_addr_i[12]  | ~\new_[18026]_ );
  assign \new_[11252]_  = (~\new_[17213]_  | ~\m6_addr_i[31] ) & (~\new_[20544]_  | ~\new_[31001]_ );
  assign \new_[11253]_  = (~\new_[17213]_  | ~\m6_addr_i[30] ) & (~\new_[20544]_  | ~\new_[31147]_ );
  assign \new_[11254]_  = (~\m7_addr_i[10]  | ~\new_[18104]_ ) & (~\m0_addr_i[10]  | ~\new_[18026]_ );
  assign \new_[11255]_  = (~\new_[18098]_  | ~\new_[31531]_ ) & (~\new_[18026]_  | ~\new_[31481]_ );
  assign \new_[11256]_  = (~\m2_addr_i[10]  | ~\new_[18077]_ ) & (~\m1_addr_i[10]  | ~\new_[19632]_ );
  assign \new_[11257]_  = (~\new_[17213]_  | ~\m6_addr_i[29] ) & (~\new_[20544]_  | ~\new_[31407]_ );
  assign \new_[11258]_  = (~\new_[18101]_  | ~\new_[30577]_ ) & (~\new_[18026]_  | ~\new_[30957]_ );
  assign \new_[11259]_  = (~\m5_addr_i[10]  | ~\new_[18753]_ ) & (~\m6_addr_i[10]  | ~\new_[17213]_ );
  assign \new_[11260]_  = (~\new_[17213]_  | ~\m6_addr_i[28] ) & (~\new_[20544]_  | ~\new_[31276]_ );
  assign \new_[11261]_  = (~\m7_addr_i[9]  | ~\new_[19584]_ ) & (~\m0_addr_i[9]  | ~\new_[18026]_ );
  assign \new_[11262]_  = (~\new_[18101]_  | ~\m7_addr_i[27] ) & (~\new_[18026]_  | ~\m0_addr_i[27] );
  assign \new_[11263]_  = (~\m2_addr_i[9]  | ~\new_[18078]_ ) & (~\m1_addr_i[9]  | ~\new_[19632]_ );
  assign \new_[11264]_  = (~\new_[17213]_  | ~\m6_addr_i[27] ) & (~\new_[20544]_  | ~\m5_addr_i[27] );
  assign \new_[11265]_  = (~\new_[18101]_  | ~\m7_addr_i[26] ) & (~\new_[18026]_  | ~\m0_addr_i[26] );
  assign \new_[11266]_  = (~\m7_addr_i[8]  | ~\new_[18102]_ ) & (~\m0_addr_i[8]  | ~\new_[18026]_ );
  assign \new_[11267]_  = (~\new_[17213]_  | ~\m6_addr_i[26] ) & (~\new_[20544]_  | ~\m5_addr_i[26] );
  assign \new_[11268]_  = (~\m2_addr_i[8]  | ~\new_[18077]_ ) & (~\m1_addr_i[8]  | ~\new_[19632]_ );
  assign \new_[11269]_  = (~\m7_addr_i[7]  | ~\new_[18102]_ ) & (~\m0_addr_i[7]  | ~\new_[18026]_ );
  assign \new_[11270]_  = (~\m2_addr_i[7]  | ~\new_[18077]_ ) & (~\m1_addr_i[7]  | ~\new_[19632]_ );
  assign \new_[11271]_  = (~\m5_addr_i[7]  | ~\new_[18756]_ ) & (~\m6_addr_i[7]  | ~\new_[17213]_ );
  assign \new_[11272]_  = (~\m7_addr_i[6]  | ~\new_[18106]_ ) & (~\m0_addr_i[6]  | ~\new_[18026]_ );
  assign \new_[11273]_  = (~\m2_addr_i[6]  | ~\new_[18078]_ ) & (~\m1_addr_i[6]  | ~\new_[19632]_ );
  assign \new_[11274]_  = ~\new_[28170]_  & (~\new_[16494]_  | ~\new_[28644]_ );
  assign \new_[11275]_  = (~\m7_addr_i[5]  | ~\new_[18110]_ ) & (~\new_[31848]_  | ~\new_[18026]_ );
  assign \new_[11276]_  = (~\m2_addr_i[5]  | ~\new_[18077]_ ) & (~\m1_addr_i[5]  | ~\new_[18190]_ );
  assign \new_[11277]_  = (~\m5_addr_i[5]  | ~\new_[18755]_ ) & (~\m6_addr_i[5]  | ~\new_[17213]_ );
  assign \new_[11278]_  = (~\m7_addr_i[4]  | ~\new_[19584]_ ) & (~\m0_addr_i[4]  | ~\new_[18026]_ );
  assign \new_[11279]_  = (~\m2_addr_i[4]  | ~\new_[18077]_ ) & (~\m1_addr_i[4]  | ~\new_[18186]_ );
  assign \new_[11280]_  = (~\new_[31726]_  | ~\new_[18107]_ ) & (~\m0_addr_i[3]  | ~\new_[18026]_ );
  assign \new_[11281]_  = (~\m7_addr_i[2]  | ~\new_[18110]_ ) & (~\m0_addr_i[2]  | ~\new_[18026]_ );
  assign \new_[11282]_  = (~\m2_addr_i[2]  | ~\new_[18077]_ ) & (~\m1_addr_i[2]  | ~\new_[18190]_ );
  assign \new_[11283]_  = (~\m7_addr_i[1]  | ~\new_[18099]_ ) & (~\m0_addr_i[1]  | ~\new_[18026]_ );
  assign \new_[11284]_  = (~\m2_addr_i[1]  | ~\new_[18078]_ ) & (~\m1_addr_i[1]  | ~\new_[18184]_ );
  assign \new_[11285]_  = (~\m7_addr_i[0]  | ~\new_[18109]_ ) & (~\m0_addr_i[0]  | ~\new_[18026]_ );
  assign \new_[11286]_  = (~\m2_addr_i[0]  | ~\new_[18077]_ ) & (~\m1_addr_i[0]  | ~\new_[18189]_ );
  assign \new_[11287]_  = (~\m7_data_i[6]  | ~\new_[19584]_ ) & (~\m0_data_i[6]  | ~\new_[18026]_ );
  assign \new_[11288]_  = (~\m7_sel_i[3]  | ~\new_[18100]_ ) & (~\m0_sel_i[3]  | ~\new_[18026]_ );
  assign \new_[11289]_  = (~\m2_sel_i[3]  | ~\new_[18077]_ ) & (~\m1_sel_i[3]  | ~\new_[18181]_ );
  assign \new_[11290]_  = (~\m5_sel_i[3]  | ~\new_[18751]_ ) & (~\m6_sel_i[3]  | ~\new_[17213]_ );
  assign \new_[11291]_  = (~\m7_sel_i[2]  | ~\new_[19584]_ ) & (~\m0_sel_i[2]  | ~\new_[18026]_ );
  assign \new_[11292]_  = (~\m2_sel_i[2]  | ~\new_[18078]_ ) & (~\m1_sel_i[2]  | ~\new_[18188]_ );
  assign \new_[11293]_  = (~\m2_sel_i[1]  | ~\new_[18078]_ ) & (~\m1_sel_i[1]  | ~\new_[18188]_ );
  assign \new_[11294]_  = (~\m7_sel_i[1]  | ~\new_[19584]_ ) & (~\m0_sel_i[1]  | ~\new_[18026]_ );
  assign \new_[11295]_  = (~\m5_sel_i[1]  | ~\new_[18751]_ ) & (~\m6_sel_i[1]  | ~\new_[18787]_ );
  assign \new_[11296]_  = (~\m7_sel_i[0]  | ~\new_[19584]_ ) & (~\m0_sel_i[0]  | ~\new_[18026]_ );
  assign \new_[11297]_  = (~\m2_sel_i[0]  | ~\new_[18078]_ ) & (~\m1_sel_i[0]  | ~\new_[18188]_ );
  assign \new_[11298]_  = (~\m5_sel_i[0]  | ~\new_[20544]_ ) & (~\m6_sel_i[0]  | ~\new_[18787]_ );
  assign \new_[11299]_  = (~m7_we_i | ~\new_[19584]_ ) & (~m0_we_i | ~\new_[18026]_ );
  assign \new_[11300]_  = (~\m7_addr_i[11]  | ~\new_[18104]_ ) & (~\m0_addr_i[11]  | ~\new_[18026]_ );
  assign \new_[11301]_  = (~m5_we_i | ~\new_[18757]_ ) & (~m6_we_i | ~\new_[17213]_ );
  assign \new_[11302]_  = (~\new_[19606]_  | ~\m7_addr_i[26] ) & (~\new_[20547]_  | ~\m0_addr_i[26] );
  assign \new_[11303]_  = (~\m7_data_i[31]  | ~\new_[18835]_ ) & (~\m0_data_i[31]  | ~\new_[20578]_ );
  assign \new_[11304]_  = (~\m5_data_i[31]  | ~\new_[18871]_ ) & (~\m6_data_i[31]  | ~\new_[18052]_ );
  assign \new_[11305]_  = (~\m7_data_i[30]  | ~\new_[18835]_ ) & (~\m0_data_i[30]  | ~\new_[19642]_ );
  assign \new_[11306]_  = (~\m7_data_i[29]  | ~\new_[18835]_ ) & (~\m0_data_i[29]  | ~\new_[20578]_ );
  assign \new_[11307]_  = (~\m5_data_i[29]  | ~\new_[18871]_ ) & (~\m6_data_i[29]  | ~\new_[20552]_ );
  assign \new_[11308]_  = ~\new_[26477]_  & (~\new_[16495]_  | ~\new_[24705]_ );
  assign \new_[11309]_  = (~\m7_data_i[4]  | ~\new_[18108]_ ) & (~\m0_data_i[4]  | ~\new_[18026]_ );
  assign \new_[11310]_  = (~\m7_data_i[28]  | ~\new_[18835]_ ) & (~\m0_data_i[28]  | ~\new_[20578]_ );
  assign \new_[11311]_  = (~\m5_data_i[28]  | ~\new_[18871]_ ) & (~\m6_data_i[28]  | ~\new_[18794]_ );
  assign \new_[11312]_  = (~\m7_data_i[27]  | ~\new_[18835]_ ) & (~\m0_data_i[27]  | ~\new_[19642]_ );
  assign \new_[11313]_  = (~\m5_data_i[27]  | ~\new_[18871]_ ) & (~\m6_data_i[27]  | ~\new_[18794]_ );
  assign \new_[11314]_  = (~\m7_addr_i[18]  | ~\new_[19606]_ ) & (~\m0_addr_i[18]  | ~\new_[18781]_ );
  assign \new_[11315]_  = (~\m7_data_i[26]  | ~\new_[18835]_ ) & (~\m0_data_i[26]  | ~\new_[20578]_ );
  assign \new_[11316]_  = ~s3_ack_i | ~\new_[17193]_  | ~\new_[30709]_ ;
  assign \new_[11317]_  = (~\m5_data_i[26]  | ~\new_[18871]_ ) & (~\m6_data_i[26]  | ~\new_[18052]_ );
  assign \new_[11318]_  = (~\m7_data_i[25]  | ~\new_[18835]_ ) & (~\m0_data_i[25]  | ~\new_[20578]_ );
  assign \new_[11319]_  = (~\m5_data_i[25]  | ~\new_[18871]_ ) & (~\m6_data_i[25]  | ~\new_[20552]_ );
  assign \new_[11320]_  = (~\m7_data_i[24]  | ~\new_[18835]_ ) & (~\m0_data_i[24]  | ~\new_[20578]_ );
  assign \new_[11321]_  = (~\m5_data_i[24]  | ~\new_[18871]_ ) & (~\m6_data_i[24]  | ~\new_[18794]_ );
  assign \new_[11322]_  = (~\m5_addr_i[18]  | ~\new_[18758]_ ) & (~\m6_addr_i[18]  | ~\new_[17213]_ );
  assign \new_[11323]_  = (~\m7_data_i[22]  | ~\new_[18835]_ ) & (~\m0_data_i[22]  | ~\new_[20578]_ );
  assign \new_[11324]_  = ~\new_[26498]_  & (~\new_[16496]_  | ~\new_[28802]_ );
  assign \new_[11325]_  = (~\m5_data_i[22]  | ~\new_[18871]_ ) & (~\m6_data_i[22]  | ~\new_[18052]_ );
  assign \new_[11326]_  = \new_[14833]_  & \new_[29043]_ ;
  assign \new_[11327]_  = (~\m7_data_i[21]  | ~\new_[18835]_ ) & (~\m0_data_i[21]  | ~\new_[20578]_ );
  assign \new_[11328]_  = (~\m7_data_i[20]  | ~\new_[18835]_ ) & (~\m0_data_i[20]  | ~\new_[19642]_ );
  assign \new_[11329]_  = (~\m7_data_i[19]  | ~\new_[18835]_ ) & (~\m0_data_i[19]  | ~\new_[20578]_ );
  assign \new_[11330]_  = (~\m5_data_i[19]  | ~\new_[18871]_ ) & (~\m6_data_i[19]  | ~\new_[18052]_ );
  assign \new_[11331]_  = (~\m7_data_i[18]  | ~\new_[18835]_ ) & (~\m0_data_i[18]  | ~\new_[18937]_ );
  assign \new_[11332]_  = ~\new_[26698]_  & (~\new_[16498]_  | ~\new_[27633]_ );
  assign \new_[11333]_  = (~\m7_data_i[17]  | ~\new_[18835]_ ) & (~\m0_data_i[17]  | ~\new_[20578]_ );
  assign \new_[11334]_  = (~\m5_data_i[17]  | ~\new_[18871]_ ) & (~\m6_data_i[17]  | ~\new_[18052]_ );
  assign \new_[11335]_  = (~\m7_data_i[16]  | ~\new_[18835]_ ) & (~\m0_data_i[16]  | ~\new_[20578]_ );
  assign \new_[11336]_  = (~\m5_data_i[16]  | ~\new_[18871]_ ) & (~\m6_data_i[16]  | ~\new_[18052]_ );
  assign \new_[11337]_  = (~\m7_data_i[15]  | ~\new_[18835]_ ) & (~\m0_data_i[15]  | ~\new_[18937]_ );
  assign \new_[11338]_  = (~\m5_data_i[15]  | ~\new_[18871]_ ) & (~\m6_data_i[15]  | ~\new_[18052]_ );
  assign \new_[11339]_  = (~\m7_data_i[14]  | ~\new_[18835]_ ) & (~\m0_data_i[14]  | ~\new_[18937]_ );
  assign \new_[11340]_  = (~\m2_data_i[10]  | ~\new_[18078]_ ) & (~\m1_data_i[10]  | ~\new_[19632]_ );
  assign \new_[11341]_  = (~\m5_data_i[14]  | ~\new_[18871]_ ) & (~\m6_data_i[14]  | ~\new_[18052]_ );
  assign \new_[11342]_  = (~\m7_data_i[13]  | ~\new_[18835]_ ) & (~\m0_data_i[13]  | ~\new_[18937]_ );
  assign \new_[11343]_  = (~\m5_data_i[13]  | ~\new_[18871]_ ) & (~\m6_data_i[13]  | ~\new_[18052]_ );
  assign \new_[11344]_  = ~s8_err_i | ~\new_[14836]_  | ~\new_[29420]_ ;
  assign \new_[11345]_  = ~s11_err_i | ~\new_[17229]_  | ~\new_[30284]_ ;
  assign \new_[11346]_  = (~\m5_data_i[12]  | ~\new_[18871]_ ) & (~\m6_data_i[12]  | ~\new_[18052]_ );
  assign \new_[11347]_  = (~\m5_data_i[11]  | ~\new_[18871]_ ) & (~\m6_data_i[11]  | ~\new_[18052]_ );
  assign \new_[11348]_  = (~\m5_data_i[10]  | ~\new_[18871]_ ) & (~\m6_data_i[10]  | ~\new_[18052]_ );
  assign \new_[11349]_  = (~\m7_data_i[9]  | ~\new_[18835]_ ) & (~\m0_data_i[9]  | ~\new_[18937]_ );
  assign \new_[11350]_  = (~\m5_data_i[9]  | ~\new_[18871]_ ) & (~\m6_data_i[9]  | ~\new_[18052]_ );
  assign \new_[11351]_  = (~\m7_data_i[8]  | ~\new_[18835]_ ) & (~\m0_data_i[8]  | ~\new_[18937]_ );
  assign \new_[11352]_  = (~\m5_data_i[8]  | ~\new_[18871]_ ) & (~\m6_data_i[8]  | ~\new_[18052]_ );
  assign \new_[11353]_  = ~s3_err_i | ~\new_[17193]_  | ~\new_[30709]_ ;
  assign \new_[11354]_  = ~s2_err_i | ~\new_[17216]_  | ~\new_[29788]_ ;
  assign \new_[11355]_  = (~\m5_data_i[7]  | ~\new_[18871]_ ) & (~\m6_data_i[7]  | ~\new_[18052]_ );
  assign \new_[11356]_  = (~\m7_data_i[6]  | ~\new_[18835]_ ) & (~\m0_data_i[6]  | ~\new_[18937]_ );
  assign \new_[11357]_  = (~\m5_data_i[6]  | ~\new_[18871]_ ) & (~\m6_data_i[6]  | ~\new_[18052]_ );
  assign \new_[11358]_  = ~s3_rty_i | ~\new_[17193]_  | ~\new_[30709]_ ;
  assign \new_[11359]_  = (~\m7_data_i[5]  | ~\new_[18835]_ ) & (~\m0_data_i[5]  | ~\new_[18937]_ );
  assign \new_[11360]_  = (~\m5_data_i[5]  | ~\new_[18871]_ ) & (~\m6_data_i[5]  | ~\new_[18052]_ );
  assign \new_[11361]_  = (~\m5_data_i[4]  | ~\new_[18871]_ ) & (~\m6_data_i[4]  | ~\new_[18795]_ );
  assign \new_[11362]_  = (~\m5_data_i[3]  | ~\new_[18871]_ ) & (~\m6_data_i[3]  | ~\new_[18795]_ );
  assign \new_[11363]_  = ~m4_stb_i | ~\new_[17268]_  | ~\new_[28223]_ ;
  assign \new_[11364]_  = (~\m5_data_i[2]  | ~\new_[18871]_ ) & (~\m6_data_i[2]  | ~\new_[18795]_ );
  assign \new_[11365]_  = (~\m5_data_i[1]  | ~\new_[18871]_ ) & (~\m6_data_i[1]  | ~\new_[18052]_ );
  assign \new_[11366]_  = (~\m5_data_i[0]  | ~\new_[18871]_ ) & (~\m6_data_i[0]  | ~\new_[18795]_ );
  assign \new_[11367]_  = ~m2_stb_i | ~\new_[17222]_  | ~\new_[29709]_ ;
  assign \new_[11368]_  = (~\m7_addr_i[23]  | ~\new_[18835]_ ) & (~\m0_addr_i[23]  | ~\new_[20578]_ );
  assign \new_[11369]_  = ~m6_stb_i | ~\new_[17229]_  | ~\new_[30284]_ ;
  assign \new_[11370]_  = (~\m5_addr_i[23]  | ~\new_[18871]_ ) & (~\m6_addr_i[23]  | ~\new_[18052]_ );
  assign \new_[11371]_  = (~\m5_addr_i[22]  | ~\new_[18871]_ ) & (~\m6_addr_i[22]  | ~\new_[18052]_ );
  assign \new_[11372]_  = ~\new_[23107]_  & (~\new_[16499]_  | ~\new_[25564]_ );
  assign \new_[11373]_  = (~\m7_addr_i[21]  | ~\new_[18835]_ ) & (~\m0_addr_i[21]  | ~\new_[19642]_ );
  assign \new_[11374]_  = ~m4_stb_i | ~\new_[17264]_  | ~\new_[28851]_ ;
  assign \new_[11375]_  = (~\m5_addr_i[21]  | ~\new_[18871]_ ) & (~\m6_addr_i[21]  | ~\new_[18052]_ );
  assign \new_[11376]_  = ~m4_stb_i | ~\new_[17272]_  | ~\new_[29641]_ ;
  assign \new_[11377]_  = ~m2_stb_i | ~\new_[16290]_  | ~\new_[29807]_ ;
  assign \new_[11378]_  = (~\m7_addr_i[20]  | ~\new_[18835]_ ) & (~\m0_addr_i[20]  | ~\new_[19642]_ );
  assign \new_[11379]_  = (~\m7_addr_i[19]  | ~\new_[18835]_ ) & (~\m0_addr_i[19]  | ~\new_[19642]_ );
  assign \new_[11380]_  = (~\m7_addr_i[18]  | ~\new_[18835]_ ) & (~\m0_addr_i[18]  | ~\new_[19642]_ );
  assign \new_[11381]_  = ~\new_[28266]_  | (~\new_[16483]_  & ~\new_[26366]_ );
  assign \new_[11382]_  = (~\m5_addr_i[18]  | ~\new_[18871]_ ) & (~\m6_addr_i[18]  | ~\new_[20552]_ );
  assign \new_[11383]_  = ~\new_[28170]_  & (~\new_[16393]_  | ~\new_[20233]_ );
  assign \new_[11384]_  = ~\new_[26477]_  & (~\new_[16402]_  | ~\new_[21464]_ );
  assign \new_[11385]_  = ~m2_stb_i | ~\new_[17193]_  | ~\new_[30709]_ ;
  assign \new_[11386]_  = (~\m7_addr_i[12]  | ~\new_[18835]_ ) & (~\m0_addr_i[12]  | ~\new_[20578]_ );
  assign \new_[11387]_  = ~\new_[26498]_  & (~\new_[16404]_  | ~\new_[20495]_ );
  assign \new_[11388]_  = ~\new_[29805]_  & (~\new_[16405]_  | ~\new_[24350]_ );
  assign \new_[11389]_  = (~\m7_addr_i[11]  | ~\new_[18835]_ ) & (~\m0_addr_i[11]  | ~\new_[20578]_ );
  assign \new_[11390]_  = ~\new_[26698]_  & (~\new_[16407]_  | ~\new_[21493]_ );
  assign \new_[11391]_  = (~\m7_data_i[2]  | ~\new_[18107]_ ) & (~\m0_data_i[2]  | ~\new_[18026]_ );
  assign \new_[11392]_  = (~\m5_addr_i[11]  | ~\new_[18871]_ ) & (~\m6_addr_i[11]  | ~\new_[18794]_ );
  assign \new_[11393]_  = (~\m7_addr_i[10]  | ~\new_[18835]_ ) & (~\m0_addr_i[10]  | ~\new_[20578]_ );
  assign \new_[11394]_  = (~\m5_addr_i[15]  | ~\new_[18757]_ ) & (~\m6_addr_i[15]  | ~\new_[18787]_ );
  assign \new_[11395]_  = (~\m5_addr_i[10]  | ~\new_[18871]_ ) & (~\m6_addr_i[10]  | ~\new_[20552]_ );
  assign \new_[11396]_  = ~\new_[28005]_  & (~\new_[16410]_  | ~\new_[20487]_ );
  assign \new_[11397]_  = (~\m5_addr_i[8]  | ~\new_[18871]_ ) & (~\m6_addr_i[8]  | ~\new_[18795]_ );
  assign \new_[11398]_  = (~\m7_addr_i[7]  | ~\new_[18835]_ ) & (~\m0_addr_i[7]  | ~\new_[20578]_ );
  assign \new_[11399]_  = (~\m5_addr_i[7]  | ~\new_[18871]_ ) & (~\m6_addr_i[7]  | ~\new_[18794]_ );
  assign \new_[11400]_  = ~\new_[25158]_  & (~\new_[16415]_  | ~\new_[20505]_ );
  assign \new_[11401]_  = (~\m5_data_i[0]  | ~\new_[18757]_ ) & (~\m6_data_i[0]  | ~\new_[17213]_ );
  assign \new_[11402]_  = ~\new_[27042]_  & (~\new_[16420]_  | ~\new_[21492]_ );
  assign \new_[11403]_  = ~\new_[23107]_  & (~\new_[16422]_  | ~\new_[21457]_ );
  assign \new_[11404]_  = (~\m5_addr_i[3]  | ~\new_[18871]_ ) & (~\m6_addr_i[3]  | ~\new_[18795]_ );
  assign \new_[11405]_  = ~\new_[26499]_  & (~\new_[16517]_  | ~\new_[28772]_ );
  assign \new_[11406]_  = (~\m5_addr_i[2]  | ~\new_[18871]_ ) & (~\m6_addr_i[2]  | ~\new_[18795]_ );
  assign \new_[11407]_  = (~\m7_addr_i[1]  | ~\new_[18835]_ ) & (~\m0_addr_i[1]  | ~\new_[20578]_ );
  assign \new_[11408]_  = ~\new_[26642]_  & (~\new_[16538]_  | ~\new_[27662]_ );
  assign \new_[11409]_  = ~m7_stb_i | ~\new_[18096]_  | ~\new_[30106]_ ;
  assign \new_[11410]_  = (~\m5_addr_i[1]  | ~\new_[18871]_ ) & (~\m6_addr_i[1]  | ~\new_[18052]_ );
  assign \new_[11411]_  = ~\new_[21163]_  & (~\new_[16338]_  | ~\new_[26213]_ );
  assign \new_[11412]_  = (~\m5_addr_i[0]  | ~\new_[18871]_ ) & (~\m6_addr_i[0]  | ~\new_[20552]_ );
  assign \new_[11413]_  = (~\m5_sel_i[3]  | ~\new_[18871]_ ) & (~\m6_sel_i[3]  | ~\new_[20552]_ );
  assign \new_[11414]_  = (~\m5_sel_i[2]  | ~\new_[18871]_ ) & (~\m6_sel_i[2]  | ~\new_[18794]_ );
  assign \new_[11415]_  = (~\m5_sel_i[1]  | ~\new_[18871]_ ) & (~\m6_sel_i[1]  | ~\new_[18795]_ );
  assign \new_[11416]_  = (~\m5_sel_i[0]  | ~\new_[18871]_ ) & (~\m6_sel_i[0]  | ~\new_[18795]_ );
  assign \new_[11417]_  = ~s11_ack_i | ~\new_[17232]_  | ~\new_[29604]_ ;
  assign \new_[11418]_  = (~m5_we_i | ~\new_[18871]_ ) & (~m6_we_i | ~\new_[18795]_ );
  assign \new_[11419]_  = ~\new_[22204]_  & (~\new_[16339]_  | ~\new_[27418]_ );
  assign \new_[11420]_  = ~\new_[28875]_  & (~\new_[16509]_  | ~\new_[28585]_ );
  assign \new_[11421]_  = ~s11_rty_i | ~\new_[17232]_  | ~\new_[29604]_ ;
  assign \new_[11422]_  = (~\m7_data_i[31]  | ~\new_[18829]_ ) & (~\m0_data_i[31]  | ~\new_[16284]_ );
  assign \new_[11423]_  = (~\m2_data_i[31]  | ~\new_[17220]_ ) & (~\m1_data_i[31]  | ~\new_[17274]_ );
  assign \new_[11424]_  = (~\m7_data_i[30]  | ~\new_[18830]_ ) & (~\m0_data_i[30]  | ~\new_[16284]_ );
  assign \new_[11425]_  = (~\m2_data_i[15]  | ~\new_[18077]_ ) & (~\m1_data_i[15]  | ~\new_[18190]_ );
  assign \new_[11426]_  = (~\m2_data_i[29]  | ~\new_[17220]_ ) & (~\m1_data_i[29]  | ~\new_[18910]_ );
  assign \new_[11427]_  = (~\m7_data_i[29]  | ~\new_[18829]_ ) & (~\m0_data_i[29]  | ~\new_[18784]_ );
  assign \new_[11428]_  = (~\m4_data_i[29]  | ~\new_[18881]_ ) & (~\m3_data_i[29]  | ~\new_[18207]_ );
  assign \new_[11429]_  = (~\m5_data_i[29]  | ~\new_[18742]_ ) & (~\m6_data_i[29]  | ~\new_[18086]_ );
  assign \new_[11430]_  = ~m7_stb_i | ~\new_[17232]_  | ~\new_[29604]_ ;
  assign \new_[11431]_  = (~\m7_data_i[28]  | ~\new_[18829]_ ) & (~\m0_data_i[28]  | ~\new_[18784]_ );
  assign \new_[11432]_  = (~\m7_data_i[27]  | ~\new_[18830]_ ) & (~\m0_data_i[27]  | ~\new_[16284]_ );
  assign \new_[11433]_  = (~\m4_data_i[27]  | ~\new_[18881]_ ) & (~\m3_data_i[27]  | ~\new_[18207]_ );
  assign \new_[11434]_  = (~\m7_data_i[26]  | ~\new_[18830]_ ) & (~\m0_data_i[26]  | ~\new_[16284]_ );
  assign \new_[11435]_  = ~s11_err_i | ~\new_[17232]_  | ~\new_[29604]_ ;
  assign \new_[11436]_  = ~m5_stb_i | ~\new_[18004]_  | ~\new_[29640]_ ;
  assign \new_[11437]_  = (~\m7_data_i[25]  | ~\new_[18830]_ ) & (~\m0_data_i[25]  | ~\new_[16284]_ );
  assign \new_[11438]_  = (~\m5_data_i[25]  | ~\new_[16275]_ ) & (~\m6_data_i[25]  | ~\new_[18087]_ );
  assign \new_[11439]_  = (~\m7_data_i[24]  | ~\new_[18830]_ ) & (~\m0_data_i[24]  | ~\new_[16284]_ );
  assign \new_[11440]_  = (~\m5_data_i[24]  | ~\new_[18742]_ ) & (~\m6_data_i[24]  | ~\new_[18086]_ );
  assign \new_[11441]_  = ~\new_[23097]_  & (~\new_[16516]_  | ~\new_[28167]_ );
  assign \new_[11442]_  = (~\m2_data_i[23]  | ~\new_[17220]_ ) & (~\m1_data_i[23]  | ~\new_[18910]_ );
  assign \new_[11443]_  = (~\m7_data_i[23]  | ~\new_[18829]_ ) & (~\m0_data_i[23]  | ~\new_[16284]_ );
  assign \new_[11444]_  = (~\m4_data_i[23]  | ~\new_[17267]_ ) & (~\m3_data_i[23]  | ~\new_[18206]_ );
  assign \new_[11445]_  = (~\m7_data_i[22]  | ~\new_[18830]_ ) & (~\m0_data_i[22]  | ~\new_[16284]_ );
  assign \new_[11446]_  = (~\m7_addr_i[19]  | ~\new_[18104]_ ) & (~\m0_addr_i[19]  | ~\new_[18026]_ );
  assign \new_[11447]_  = (~\m5_data_i[22]  | ~\new_[18742]_ ) & (~\m6_data_i[22]  | ~\new_[18086]_ );
  assign \new_[11448]_  = (~\m7_data_i[21]  | ~\new_[18830]_ ) & (~\m0_data_i[21]  | ~\new_[16284]_ );
  assign \new_[11449]_  = (~\m7_data_i[20]  | ~\new_[18830]_ ) & (~\m0_data_i[20]  | ~\new_[16284]_ );
  assign \new_[11450]_  = ~\new_[26665]_  & (~\new_[16519]_  | ~\new_[28164]_ );
  assign \new_[11451]_  = (~\m7_data_i[19]  | ~\new_[18830]_ ) & (~\m0_data_i[19]  | ~\new_[16284]_ );
  assign \new_[11452]_  = ~\new_[28706]_  & (~\new_[16444]_  | ~\new_[22872]_ );
  assign \new_[11453]_  = (~\m7_data_i[15]  | ~\new_[17232]_ ) & (~\m0_data_i[15]  | ~\new_[20580]_ );
  assign \new_[11454]_  = ~\new_[28991]_  & (~\new_[16520]_  | ~\new_[28550]_ );
  assign \new_[11455]_  = (~\m5_data_i[19]  | ~\new_[18742]_ ) & (~\m6_data_i[19]  | ~\new_[18086]_ );
  assign \new_[11456]_  = (~\m4_data_i[18]  | ~\new_[17267]_ ) & (~\m3_data_i[18]  | ~\new_[16312]_ );
  assign \new_[11457]_  = (~\m7_data_i[18]  | ~\new_[18829]_ ) & (~\m0_data_i[18]  | ~\new_[16284]_ );
  assign \new_[11458]_  = (~\m2_data_i[18]  | ~\new_[17220]_ ) & (~\m1_data_i[18]  | ~\new_[18910]_ );
  assign \new_[11459]_  = (~\m5_data_i[18]  | ~\new_[18742]_ ) & (~\m6_data_i[18]  | ~\new_[18087]_ );
  assign \new_[11460]_  = (~\m7_data_i[17]  | ~\new_[18830]_ ) & (~\m0_data_i[17]  | ~\new_[16284]_ );
  assign \new_[11461]_  = (~\m7_data_i[16]  | ~\new_[18830]_ ) & (~\m0_data_i[16]  | ~\new_[16284]_ );
  assign \new_[11462]_  = (~\m5_data_i[16]  | ~\new_[16275]_ ) & (~\m6_data_i[16]  | ~\new_[18086]_ );
  assign \new_[11463]_  = (~\m7_data_i[15]  | ~\new_[18830]_ ) & (~\m0_data_i[15]  | ~\new_[16284]_ );
  assign \new_[11464]_  = ~\new_[29716]_  & (~\new_[16522]_  | ~\new_[28122]_ );
  assign \new_[11465]_  = (~\m4_data_i[15]  | ~\new_[17267]_ ) & (~\m3_data_i[15]  | ~\new_[16312]_ );
  assign \new_[11466]_  = (~\m5_data_i[15]  | ~\new_[16275]_ ) & (~\m6_data_i[15]  | ~\new_[19577]_ );
  assign \new_[11467]_  = (~\m4_data_i[14]  | ~\new_[17267]_ ) & (~\m3_data_i[14]  | ~\new_[16312]_ );
  assign \new_[11468]_  = (~\m7_data_i[14]  | ~\new_[18829]_ ) & (~\m0_data_i[14]  | ~\new_[18784]_ );
  assign \new_[11469]_  = (~\m5_data_i[14]  | ~\new_[16275]_ ) & (~\m6_data_i[14]  | ~\new_[18087]_ );
  assign \new_[11470]_  = (~\m4_data_i[13]  | ~\new_[17267]_ ) & (~\m3_data_i[13]  | ~\new_[16312]_ );
  assign \new_[11471]_  = (~\m7_data_i[13]  | ~\new_[18829]_ ) & (~\m0_data_i[13]  | ~\new_[18784]_ );
  assign \new_[11472]_  = (~\m5_data_i[13]  | ~\new_[16275]_ ) & (~\m6_data_i[13]  | ~\new_[18087]_ );
  assign \new_[11473]_  = (~\m7_data_i[12]  | ~\new_[18830]_ ) & (~\m0_data_i[12]  | ~\new_[16284]_ );
  assign \new_[11474]_  = (~\m4_data_i[12]  | ~\new_[17267]_ ) & (~\m3_data_i[12]  | ~\new_[16312]_ );
  assign \new_[11475]_  = (~\m7_data_i[11]  | ~\new_[18830]_ ) & (~\m0_data_i[11]  | ~\new_[16284]_ );
  assign \new_[11476]_  = (~\m2_data_i[11]  | ~\new_[17220]_ ) & (~\m1_data_i[11]  | ~\new_[18910]_ );
  assign \new_[11477]_  = (~\m4_data_i[11]  | ~\new_[17267]_ ) & (~\m3_data_i[11]  | ~\new_[16312]_ );
  assign \new_[11478]_  = (~\m7_data_i[10]  | ~\new_[18829]_ ) & (~\m0_data_i[10]  | ~\new_[16284]_ );
  assign \new_[11479]_  = ~\new_[28763]_  & (~\new_[16525]_  | ~\new_[28297]_ );
  assign \new_[11480]_  = (~\m5_data_i[3]  | ~\new_[18747]_ ) & (~\m6_data_i[3]  | ~\new_[18787]_ );
  assign \new_[11481]_  = (~\m7_data_i[9]  | ~\new_[18829]_ ) & (~\m0_data_i[9]  | ~\new_[18784]_ );
  assign \new_[11482]_  = (~\m7_data_i[8]  | ~\new_[18829]_ ) & (~\m0_data_i[8]  | ~\new_[16284]_ );
  assign \new_[11483]_  = ~\new_[22440]_  & (~\new_[16340]_  | ~\new_[26572]_ );
  assign \new_[11484]_  = (~\m2_data_i[7]  | ~\new_[17220]_ ) & (~\m1_data_i[7]  | ~\new_[18910]_ );
  assign \new_[11485]_  = (~\m7_data_i[7]  | ~\new_[18830]_ ) & (~\m0_data_i[7]  | ~\new_[16284]_ );
  assign \new_[11486]_  = (~\m4_data_i[7]  | ~\new_[17267]_ ) & (~\m3_data_i[7]  | ~\new_[16312]_ );
  assign \new_[11487]_  = (~\m5_data_i[7]  | ~\new_[16275]_ ) & (~\m6_data_i[7]  | ~\new_[19577]_ );
  assign \new_[11488]_  = ~\new_[28026]_  & (~\new_[16527]_  | ~\new_[28306]_ );
  assign \new_[11489]_  = (~\m5_data_i[6]  | ~\new_[16275]_ ) & (~\m6_data_i[6]  | ~\new_[18087]_ );
  assign \new_[11490]_  = (~\m7_data_i[6]  | ~\new_[18829]_ ) & (~\m0_data_i[6]  | ~\new_[16284]_ );
  assign \new_[11491]_  = ~\new_[27871]_  & (~\new_[16529]_  | ~\new_[28241]_ );
  assign \new_[11492]_  = (~\m2_data_i[5]  | ~\new_[17220]_ ) & (~\m1_data_i[5]  | ~\new_[18180]_ );
  assign \new_[11493]_  = (~\m7_data_i[5]  | ~\new_[18829]_ ) & (~\m0_data_i[5]  | ~\new_[16284]_ );
  assign \new_[11494]_  = (~\m5_data_i[4]  | ~\new_[16275]_ ) & (~\m6_data_i[4]  | ~\new_[19577]_ );
  assign \new_[11495]_  = ~\new_[26766]_  | (~\new_[16534]_  & ~\new_[25439]_ );
  assign \new_[11496]_  = (~\m7_data_i[4]  | ~\new_[18829]_ ) & (~\m0_data_i[4]  | ~\new_[18784]_ );
  assign \new_[11497]_  = ~\new_[28034]_  | (~\new_[16535]_  & ~\new_[27818]_ );
  assign \new_[11498]_  = (~\m7_data_i[3]  | ~\new_[18829]_ ) & (~\m0_data_i[3]  | ~\new_[18784]_ );
  assign \new_[11499]_  = ~\new_[28630]_  | (~\new_[16536]_  & ~\new_[24761]_ );
  assign \new_[11500]_  = (~\m2_data_i[2]  | ~\new_[17220]_ ) & (~\m1_data_i[2]  | ~\new_[18910]_ );
  assign \new_[11501]_  = (~\m7_data_i[2]  | ~\new_[18829]_ ) & (~\m0_data_i[2]  | ~\new_[16284]_ );
  assign \new_[11502]_  = ~\new_[30182]_  | (~\new_[16537]_  & ~\new_[28308]_ );
  assign \new_[11503]_  = (~\m7_data_i[30]  | ~\new_[18112]_ ) & (~\m0_data_i[30]  | ~\new_[18019]_ );
  assign \new_[11504]_  = (~\m7_data_i[1]  | ~\new_[18829]_ ) & (~\m0_data_i[1]  | ~\new_[18784]_ );
  assign \new_[11505]_  = (~\m4_data_i[0]  | ~\new_[17267]_ ) & (~\m3_data_i[0]  | ~\new_[16312]_ );
  assign \new_[11506]_  = (~\m7_data_i[0]  | ~\new_[18829]_ ) & (~\m0_data_i[0]  | ~\new_[18784]_ );
  assign \new_[11507]_  = (~\m5_data_i[0]  | ~\new_[16275]_ ) & (~\m6_data_i[0]  | ~\new_[18087]_ );
  assign \new_[11508]_  = (~\new_[18829]_  | ~\m7_addr_i[31] ) & (~\new_[16284]_  | ~\m0_addr_i[31] );
  assign \new_[11509]_  = (~\new_[19577]_  | ~\m6_addr_i[30] ) & (~\new_[16275]_  | ~\new_[31147]_ );
  assign \new_[11510]_  = (~\new_[17220]_  | ~\new_[31486]_ ) & (~\new_[17274]_  | ~\new_[31308]_ );
  assign \new_[11511]_  = (~\new_[18829]_  | ~\new_[31885]_ ) & (~\new_[16284]_  | ~\new_[31292]_ );
  assign \new_[11512]_  = (~\new_[17267]_  | ~\m4_addr_i[29] ) & (~\new_[16312]_  | ~\m3_addr_i[29] );
  assign \new_[11513]_  = (~\new_[18829]_  | ~\new_[31531]_ ) & (~\new_[16284]_  | ~\new_[31481]_ );
  assign \new_[11514]_  = (~\new_[17267]_  | ~\m4_addr_i[28] ) & (~\new_[16312]_  | ~\m3_addr_i[28] );
  assign \new_[11515]_  = (~\m2_sel_i[2]  | ~\new_[18069]_ ) & (~\m1_sel_i[2]  | ~\new_[18901]_ );
  assign \new_[11516]_  = ~\new_[29160]_  | (~\new_[16539]_  & ~\new_[28813]_ );
  assign \new_[11517]_  = (~\new_[17220]_  | ~\new_[31547]_ ) & (~\new_[17274]_  | ~\new_[31458]_ );
  assign \new_[11518]_  = (~\m5_data_i[5]  | ~\new_[18753]_ ) & (~\m6_data_i[5]  | ~\new_[17213]_ );
  assign \new_[11519]_  = (~\new_[18830]_  | ~\new_[30577]_ ) & (~\new_[18784]_  | ~\new_[30957]_ );
  assign \new_[11520]_  = (~\new_[17220]_  | ~\m2_addr_i[27] ) & (~\new_[18910]_  | ~\m1_addr_i[27] );
  assign \new_[11521]_  = ~\new_[29193]_  | (~\new_[16540]_  & ~\new_[26426]_ );
  assign \new_[11522]_  = (~\new_[17267]_  | ~\m4_addr_i[27] ) & (~\new_[18207]_  | ~\m3_addr_i[27] );
  assign \new_[11523]_  = (~\new_[18830]_  | ~\m7_addr_i[27] ) & (~\new_[18784]_  | ~\m0_addr_i[27] );
  assign \new_[11524]_  = (~\new_[18829]_  | ~\m7_addr_i[26] ) & (~\new_[16284]_  | ~\m0_addr_i[26] );
  assign \new_[11525]_  = (~\new_[19577]_  | ~\m6_addr_i[25] ) & (~\new_[16275]_  | ~\m5_addr_i[25] );
  assign \new_[11526]_  = (~\new_[17267]_  | ~\m4_addr_i[25] ) & (~\new_[18206]_  | ~\m3_addr_i[25] );
  assign \new_[11527]_  = (~\new_[18829]_  | ~\m7_addr_i[25] ) & (~\new_[18784]_  | ~\m0_addr_i[25] );
  assign \new_[11528]_  = (~\new_[19577]_  | ~\m6_addr_i[24] ) & (~\new_[16275]_  | ~\m5_addr_i[24] );
  assign \new_[11529]_  = (~\new_[18829]_  | ~\m7_addr_i[24] ) & (~\new_[18784]_  | ~\m0_addr_i[24] );
  assign \new_[11530]_  = ~\new_[29630]_  | (~\new_[16541]_  & ~\new_[27677]_ );
  assign \new_[11531]_  = (~\new_[17267]_  | ~\m4_addr_i[24] ) & (~\new_[18206]_  | ~\m3_addr_i[24] );
  assign \new_[11532]_  = (~\m7_addr_i[23]  | ~\new_[18830]_ ) & (~\m0_addr_i[23]  | ~\new_[16284]_ );
  assign \new_[11533]_  = ~\new_[29353]_  | (~\new_[16542]_  & ~\new_[28169]_ );
  assign \new_[11534]_  = (~\m4_addr_i[23]  | ~\new_[17267]_ ) & (~\m3_addr_i[23]  | ~\new_[18207]_ );
  assign \new_[11535]_  = (~\m2_addr_i[23]  | ~\new_[17220]_ ) & (~\m1_addr_i[23]  | ~\new_[17274]_ );
  assign \new_[11536]_  = (~\m7_addr_i[22]  | ~\new_[18830]_ ) & (~\m0_addr_i[22]  | ~\new_[16284]_ );
  assign \new_[11537]_  = (~\m5_addr_i[8]  | ~\new_[18015]_ ) & (~\m6_addr_i[8]  | ~\new_[17229]_ );
  assign \new_[11538]_  = (~\m4_addr_i[22]  | ~\new_[17267]_ ) & (~\m3_addr_i[22]  | ~\new_[18206]_ );
  assign \new_[11539]_  = ~\new_[31990]_ ;
  assign \new_[11540]_  = (~\m7_addr_i[21]  | ~\new_[18830]_ ) & (~\m0_addr_i[21]  | ~\new_[16284]_ );
  assign \new_[11541]_  = ~\new_[28200]_  | (~\new_[16543]_  & ~\new_[24854]_ );
  assign \new_[11542]_  = (~\m4_addr_i[21]  | ~\new_[17267]_ ) & (~\m3_addr_i[21]  | ~\new_[16312]_ );
  assign \new_[11543]_  = (~\m5_addr_i[21]  | ~\new_[18742]_ ) & (~\m6_addr_i[21]  | ~\new_[18086]_ );
  assign \new_[11544]_  = ~\new_[26759]_  | (~\new_[16544]_  & ~\new_[26900]_ );
  assign \new_[11545]_  = (~\m7_addr_i[20]  | ~\new_[18830]_ ) & (~\m0_addr_i[20]  | ~\new_[16284]_ );
  assign \new_[11546]_  = (~\m4_addr_i[20]  | ~\new_[17267]_ ) & (~\m3_addr_i[20]  | ~\new_[16312]_ );
  assign \new_[11547]_  = (~\m5_addr_i[20]  | ~\new_[18742]_ ) & (~\m6_addr_i[20]  | ~\new_[18086]_ );
  assign \new_[11548]_  = (~\m7_addr_i[19]  | ~\new_[18830]_ ) & (~\m0_addr_i[19]  | ~\new_[16284]_ );
  assign \new_[11549]_  = ~\new_[29126]_  & (~\new_[16462]_  | ~\new_[29365]_ );
  assign \new_[11550]_  = (~\m4_addr_i[19]  | ~\new_[18881]_ ) & (~\m3_addr_i[19]  | ~\new_[16312]_ );
  assign \new_[11551]_  = (~\m7_addr_i[18]  | ~\new_[18830]_ ) & (~\m0_addr_i[18]  | ~\new_[16284]_ );
  assign \new_[11552]_  = ~\new_[26626]_  & (~\new_[16500]_  | ~\new_[22820]_ );
  assign \new_[11553]_  = (~\m5_addr_i[18]  | ~\new_[18742]_ ) & (~\m6_addr_i[18]  | ~\new_[18087]_ );
  assign \new_[11554]_  = ~\new_[26650]_  & (~\new_[16501]_  | ~\new_[22475]_ );
  assign \new_[11555]_  = (~\m7_addr_i[17]  | ~\new_[18830]_ ) & (~\m0_addr_i[17]  | ~\new_[16284]_ );
  assign \new_[11556]_  = (~\m2_data_i[17]  | ~\new_[18077]_ ) & (~\m1_data_i[17]  | ~\new_[18189]_ );
  assign \new_[11557]_  = (~\m5_addr_i[17]  | ~\new_[18742]_ ) & (~\m6_addr_i[17]  | ~\new_[18086]_ );
  assign \new_[11558]_  = (~\m7_addr_i[16]  | ~\new_[18830]_ ) & (~\m0_addr_i[16]  | ~\new_[16284]_ );
  assign \new_[11559]_  = (~\m2_addr_i[14]  | ~\new_[18078]_ ) & (~\m1_addr_i[14]  | ~\new_[18184]_ );
  assign \new_[11560]_  = (~\m4_addr_i[16]  | ~\new_[17267]_ ) & (~\m3_addr_i[16]  | ~\new_[18207]_ );
  assign \new_[11561]_  = (~\m2_addr_i[13]  | ~\new_[18069]_ ) & (~\m1_addr_i[13]  | ~\new_[18898]_ );
  assign \new_[11562]_  = (~\m7_addr_i[15]  | ~\new_[18830]_ ) & (~\m0_addr_i[15]  | ~\new_[18784]_ );
  assign \new_[11563]_  = (~\m4_addr_i[15]  | ~\new_[17267]_ ) & (~\m3_addr_i[15]  | ~\new_[18206]_ );
  assign \new_[11564]_  = ~\new_[27940]_  & (~\new_[16463]_  | ~\new_[17413]_ );
  assign \new_[11565]_  = (~\m7_addr_i[14]  | ~\new_[18830]_ ) & (~\m0_addr_i[14]  | ~\new_[16284]_ );
  assign \new_[11566]_  = (~\m4_addr_i[14]  | ~\new_[18881]_ ) & (~\m3_addr_i[14]  | ~\new_[18207]_ );
  assign \new_[11567]_  = ~\new_[29218]_  & (~\new_[16464]_  | ~\new_[21477]_ );
  assign \new_[11568]_  = (~\m7_addr_i[13]  | ~\new_[18830]_ ) & (~\m0_addr_i[13]  | ~\new_[16284]_ );
  assign \new_[11569]_  = (~\m5_addr_i[13]  | ~\new_[18742]_ ) & (~\m6_addr_i[13]  | ~\new_[18087]_ );
  assign \new_[11570]_  = ~\new_[28408]_  & (~\new_[16502]_  | ~\new_[21379]_ );
  assign \new_[11571]_  = (~\m2_addr_i[12]  | ~\new_[17220]_ ) & (~\m1_addr_i[12]  | ~\new_[18910]_ );
  assign \new_[11572]_  = (~\m7_addr_i[12]  | ~\new_[18830]_ ) & (~\m0_addr_i[12]  | ~\new_[16284]_ );
  assign \new_[11573]_  = (~\m4_addr_i[12]  | ~\new_[18881]_ ) & (~\m3_addr_i[12]  | ~\new_[18207]_ );
  assign \new_[11574]_  = (~\m7_addr_i[11]  | ~\new_[18830]_ ) & (~\m0_addr_i[11]  | ~\new_[16284]_ );
  assign \new_[11575]_  = (~\m5_addr_i[11]  | ~\new_[18742]_ ) & (~\m6_addr_i[11]  | ~\new_[18087]_ );
  assign \new_[11576]_  = (~\m7_addr_i[10]  | ~\new_[18830]_ ) & (~\m0_addr_i[10]  | ~\new_[16284]_ );
  assign \new_[11577]_  = (~\m2_addr_i[10]  | ~\new_[17220]_ ) & (~\m1_addr_i[10]  | ~\new_[17275]_ );
  assign \new_[11578]_  = (~\m4_addr_i[10]  | ~\new_[18881]_ ) & (~\m3_addr_i[10]  | ~\new_[18207]_ );
  assign \new_[11579]_  = ~\new_[26615]_  & (~\new_[16503]_  | ~\new_[21370]_ );
  assign \new_[11580]_  = (~\m5_addr_i[10]  | ~\new_[18742]_ ) & (~\m6_addr_i[10]  | ~\new_[18087]_ );
  assign \new_[11581]_  = (~\m7_addr_i[9]  | ~\new_[18830]_ ) & (~\m0_addr_i[9]  | ~\new_[16284]_ );
  assign \new_[11582]_  = (~\m4_addr_i[9]  | ~\new_[17267]_ ) & (~\m3_addr_i[9]  | ~\new_[16312]_ );
  assign \new_[11583]_  = ~\new_[24492]_  & (~\new_[16465]_  | ~\new_[29366]_ );
  assign \new_[11584]_  = (~\m7_addr_i[8]  | ~\new_[18830]_ ) & (~\m0_addr_i[8]  | ~\new_[16284]_ );
  assign \new_[11585]_  = (~\m2_addr_i[13]  | ~\new_[18077]_ ) & (~\m1_addr_i[13]  | ~\new_[18181]_ );
  assign \new_[11586]_  = ~\new_[28651]_  & (~\new_[16466]_  | ~\new_[23005]_ );
  assign \new_[11587]_  = (~\m2_addr_i[12]  | ~\new_[18078]_ ) & (~\m1_addr_i[12]  | ~\new_[18188]_ );
  assign \new_[11588]_  = (~\m5_addr_i[8]  | ~\new_[18742]_ ) & (~\m6_addr_i[8]  | ~\new_[18086]_ );
  assign \new_[11589]_  = (~\m7_addr_i[7]  | ~\new_[18830]_ ) & (~\m0_addr_i[7]  | ~\new_[16284]_ );
  assign \new_[11590]_  = (~\m5_addr_i[7]  | ~\new_[18742]_ ) & (~\m6_addr_i[7]  | ~\new_[18086]_ );
  assign \new_[11591]_  = (~\m7_addr_i[6]  | ~\new_[18830]_ ) & (~\m0_addr_i[6]  | ~\new_[16284]_ );
  assign \new_[11592]_  = (~\m2_addr_i[6]  | ~\new_[17220]_ ) & (~\m1_addr_i[6]  | ~\new_[17275]_ );
  assign \new_[11593]_  = (~\m5_addr_i[6]  | ~\new_[18742]_ ) & (~\m6_addr_i[6]  | ~\new_[18087]_ );
  assign \new_[11594]_  = (~\m7_addr_i[5]  | ~\new_[18829]_ ) & (~\new_[31848]_  | ~\new_[16284]_ );
  assign \new_[11595]_  = (~\m4_addr_i[5]  | ~\new_[17267]_ ) & (~\m3_addr_i[5]  | ~\new_[16312]_ );
  assign \new_[11596]_  = (~\m7_addr_i[4]  | ~\new_[18830]_ ) & (~\m0_addr_i[4]  | ~\new_[16284]_ );
  assign \new_[11597]_  = ~\new_[26469]_  & (~\new_[16467]_  | ~\new_[29302]_ );
  assign \new_[11598]_  = ~\new_[28303]_  & (~\new_[16468]_  | ~\new_[20501]_ );
  assign \new_[11599]_  = (~\m5_addr_i[4]  | ~\new_[16275]_ ) & (~\m6_addr_i[4]  | ~\new_[18087]_ );
  assign \new_[11600]_  = (~\new_[31726]_  | ~\new_[18830]_ ) & (~\m0_addr_i[3]  | ~\new_[16284]_ );
  assign \new_[11601]_  = (~\m4_addr_i[3]  | ~\new_[17267]_ ) & (~\m3_addr_i[3]  | ~\new_[16312]_ );
  assign \new_[11602]_  = (~\m5_addr_i[3]  | ~\new_[16275]_ ) & (~\m6_addr_i[3]  | ~\new_[19577]_ );
  assign \new_[11603]_  = (~\m7_addr_i[2]  | ~\new_[18829]_ ) & (~\m0_addr_i[2]  | ~\new_[16284]_ );
  assign \new_[11604]_  = (~\m4_addr_i[2]  | ~\new_[17267]_ ) & (~\m3_addr_i[2]  | ~\new_[16312]_ );
  assign \new_[11605]_  = (~\m5_addr_i[2]  | ~\new_[16275]_ ) & (~\m6_addr_i[2]  | ~\new_[19577]_ );
  assign \new_[11606]_  = (~\m2_addr_i[1]  | ~\new_[17220]_ ) & (~\m1_addr_i[1]  | ~\new_[18910]_ );
  assign \new_[11607]_  = ~\new_[28173]_  & (~\new_[16469]_  | ~\new_[29322]_ );
  assign \new_[11608]_  = (~\m7_addr_i[1]  | ~\new_[18829]_ ) & (~\m0_addr_i[1]  | ~\new_[18784]_ );
  assign \new_[11609]_  = (~\m4_addr_i[0]  | ~\new_[17267]_ ) & (~\m3_addr_i[0]  | ~\new_[16312]_ );
  assign \new_[11610]_  = (~\m7_addr_i[0]  | ~\new_[18829]_ ) & (~\m0_addr_i[0]  | ~\new_[16284]_ );
  assign \new_[11611]_  = \new_[14839]_ ;
  assign \new_[11612]_  = (~\m2_addr_i[0]  | ~\new_[17220]_ ) & (~\m1_addr_i[0]  | ~\new_[18910]_ );
  assign \new_[11613]_  = \new_[14839]_ ;
  assign \new_[11614]_  = (~\m7_sel_i[3]  | ~\new_[18829]_ ) & (~\m0_sel_i[3]  | ~\new_[16284]_ );
  assign \new_[11615]_  = (~\m4_sel_i[3]  | ~\new_[17267]_ ) & (~\m3_sel_i[3]  | ~\new_[18206]_ );
  assign \new_[11616]_  = ~\new_[28043]_  & (~\new_[16470]_  | ~\new_[18430]_ );
  assign \new_[11617]_  = (~\m7_sel_i[2]  | ~\new_[18830]_ ) & (~\m0_sel_i[2]  | ~\new_[16284]_ );
  assign \new_[11618]_  = ~\new_[27984]_  & (~\new_[16504]_  | ~\new_[20384]_ );
  assign \new_[11619]_  = (~\m2_sel_i[1]  | ~\new_[17220]_ ) & (~\m1_sel_i[1]  | ~\new_[18910]_ );
  assign \new_[11620]_  = (~\m7_sel_i[1]  | ~\new_[18829]_ ) & (~\m0_sel_i[1]  | ~\new_[18784]_ );
  assign \new_[11621]_  = (~\m7_sel_i[0]  | ~\new_[18830]_ ) & (~\m0_sel_i[0]  | ~\new_[16284]_ );
  assign \new_[11622]_  = (~\m2_sel_i[0]  | ~\new_[17220]_ ) & (~\m1_sel_i[0]  | ~\new_[17275]_ );
  assign \new_[11623]_  = (~\m5_sel_i[0]  | ~\new_[18742]_ ) & (~\m6_sel_i[0]  | ~\new_[18086]_ );
  assign \new_[11624]_  = ~\new_[30238]_  & (~\new_[16471]_  | ~\new_[20508]_ );
  assign \new_[11625]_  = (~m2_we_i | ~\new_[17220]_ ) & (~m1_we_i | ~\new_[18910]_ );
  assign \new_[11626]_  = (~m7_we_i | ~\new_[18830]_ ) & (~m0_we_i | ~\new_[16284]_ );
  assign \new_[11627]_  = (~m4_we_i | ~\new_[17267]_ ) & (~m3_we_i | ~\new_[16312]_ );
  assign \new_[11628]_  = (~m5_we_i | ~\new_[16275]_ ) & (~m6_we_i | ~\new_[18087]_ );
  assign \new_[11629]_  = ~\new_[28895]_  & (~\new_[16505]_  | ~\new_[22717]_ );
  assign \new_[11630]_  = (~\m7_data_i[31]  | ~\new_[18832]_ ) & (~\m0_data_i[31]  | ~\new_[18066]_ );
  assign \new_[11631]_  = (~\m5_data_i[31]  | ~\new_[18744]_ ) & (~\m6_data_i[31]  | ~\new_[16289]_ );
  assign \new_[11632]_  = (~\m4_data_i[31]  | ~\new_[17268]_ ) & (~\m3_data_i[31]  | ~\new_[19597]_ );
  assign \new_[11633]_  = ~\new_[26670]_  & (~\new_[16472]_  | ~\new_[17418]_ );
  assign \new_[11634]_  = (~\m7_data_i[30]  | ~\new_[18832]_ ) & (~\m0_data_i[30]  | ~\new_[18066]_ );
  assign \new_[11635]_  = (~\m4_data_i[30]  | ~\new_[17268]_ ) & (~\m3_data_i[30]  | ~\new_[19597]_ );
  assign \new_[11636]_  = (~\m5_data_i[30]  | ~\new_[18744]_ ) & (~\m6_data_i[30]  | ~\new_[16289]_ );
  assign \new_[11637]_  = (~\m5_data_i[29]  | ~\new_[20542]_ ) & (~\m6_data_i[29]  | ~\new_[16289]_ );
  assign \new_[11638]_  = ~\new_[27881]_  & (~\new_[16506]_  | ~\new_[22906]_ );
  assign \new_[11639]_  = (~\m7_data_i[29]  | ~\new_[18832]_ ) & (~\m0_data_i[29]  | ~\new_[18066]_ );
  assign \new_[11640]_  = (~\m2_data_i[4]  | ~\new_[18078]_ ) & (~\m1_data_i[4]  | ~\new_[18185]_ );
  assign \new_[11641]_  = (~\m7_data_i[28]  | ~\new_[18832]_ ) & (~\m0_data_i[28]  | ~\new_[18066]_ );
  assign \new_[11642]_  = (~\m4_data_i[28]  | ~\new_[17268]_ ) & (~\m3_data_i[28]  | ~\new_[19597]_ );
  assign \new_[11643]_  = (~\m5_data_i[28]  | ~\new_[18744]_ ) & (~\m6_data_i[28]  | ~\new_[16289]_ );
  assign \new_[11644]_  = ~\new_[29125]_  & (~\new_[16473]_  | ~\new_[20466]_ );
  assign \new_[11645]_  = (~\m7_data_i[27]  | ~\new_[18832]_ ) & (~\m0_data_i[27]  | ~\new_[18066]_ );
  assign \new_[11646]_  = (~\m5_data_i[27]  | ~\new_[18744]_ ) & (~\m6_data_i[27]  | ~\new_[16289]_ );
  assign \new_[11647]_  = (~\m7_data_i[26]  | ~\new_[18832]_ ) & (~\m0_data_i[26]  | ~\new_[18066]_ );
  assign \new_[11648]_  = (~\m5_data_i[26]  | ~\new_[18744]_ ) & (~\m6_data_i[26]  | ~\new_[16289]_ );
  assign \new_[11649]_  = (~\m5_data_i[25]  | ~\new_[20542]_ ) & (~\m6_data_i[25]  | ~\new_[16289]_ );
  assign \new_[11650]_  = ~\new_[27861]_  & (~\new_[16474]_  | ~\new_[21573]_ );
  assign \new_[11651]_  = ~\new_[14850]_ ;
  assign \new_[11652]_  = (~\m5_data_i[24]  | ~\new_[20542]_ ) & (~\m6_data_i[24]  | ~\new_[16289]_ );
  assign \new_[11653]_  = (~\m7_data_i[23]  | ~\new_[18832]_ ) & (~\m0_data_i[23]  | ~\new_[18066]_ );
  assign \new_[11654]_  = ~\new_[27015]_  & (~\new_[16507]_  | ~\new_[24035]_ );
  assign \new_[11655]_  = (~\m5_data_i[23]  | ~\new_[18743]_ ) & (~\m6_data_i[23]  | ~\new_[16289]_ );
  assign \new_[11656]_  = (~\m7_data_i[22]  | ~\new_[18832]_ ) & (~\m0_data_i[22]  | ~\new_[18066]_ );
  assign \new_[11657]_  = (~\m5_data_i[16]  | ~\new_[20544]_ ) & (~\m6_data_i[16]  | ~\new_[17213]_ );
  assign \new_[11658]_  = (~\m4_data_i[22]  | ~\new_[17268]_ ) & (~\m3_data_i[22]  | ~\new_[18854]_ );
  assign \new_[11659]_  = (~\m2_data_i[1]  | ~\new_[18078]_ ) & (~\m1_data_i[1]  | ~\new_[18185]_ );
  assign \new_[11660]_  = (~\m5_data_i[22]  | ~\new_[18744]_ ) & (~\m6_data_i[22]  | ~\new_[16289]_ );
  assign \new_[11661]_  = (~\m7_data_i[21]  | ~\new_[18832]_ ) & (~\m0_data_i[21]  | ~\new_[18066]_ );
  assign \new_[11662]_  = (~\m5_data_i[21]  | ~\new_[20542]_ ) & (~\m6_data_i[21]  | ~\new_[16289]_ );
  assign \new_[11663]_  = (~\m5_data_i[20]  | ~\new_[20542]_ ) & (~\m6_data_i[20]  | ~\new_[16289]_ );
  assign \new_[11664]_  = (~\m5_data_i[19]  | ~\new_[20542]_ ) & (~\m6_data_i[19]  | ~\new_[16289]_ );
  assign \new_[11665]_  = (~\m7_data_i[19]  | ~\new_[18832]_ ) & (~\m0_data_i[19]  | ~\new_[18066]_ );
  assign \new_[11666]_  = (~\m7_data_i[18]  | ~\new_[18832]_ ) & (~\m0_data_i[18]  | ~\new_[18066]_ );
  assign \new_[11667]_  = (~\m5_data_i[18]  | ~\new_[18744]_ ) & (~\m6_data_i[18]  | ~\new_[16289]_ );
  assign \new_[11668]_  = (~\m7_data_i[17]  | ~\new_[18832]_ ) & (~\m0_data_i[17]  | ~\new_[18066]_ );
  assign \new_[11669]_  = (~\m5_data_i[17]  | ~\new_[18744]_ ) & (~\m6_data_i[17]  | ~\new_[16289]_ );
  assign \new_[11670]_  = (~\m7_addr_i[21]  | ~\new_[17240]_ ) & (~\m6_addr_i[21]  | ~\new_[19581]_ );
  assign \new_[11671]_  = ~\new_[26474]_  & (~\new_[16476]_  | ~\new_[29751]_ );
  assign \new_[11672]_  = ~\new_[28677]_  & (~\new_[16477]_  | ~\new_[23231]_ );
  assign \new_[11673]_  = (~\m4_data_i[16]  | ~\new_[17268]_ ) & (~\m3_data_i[16]  | ~\new_[19597]_ );
  assign \new_[11674]_  = ~\new_[26763]_  & (~\new_[16508]_  | ~\new_[21381]_ );
  assign \new_[11675]_  = (~\m2_data_i[16]  | ~\new_[18078]_ ) & (~\m1_data_i[16]  | ~\new_[18184]_ );
  assign \new_[11676]_  = (~\m5_data_i[12]  | ~\new_[18743]_ ) & (~\m6_data_i[12]  | ~\new_[16289]_ );
  assign \new_[11677]_  = (~\new_[16429]_  | ~\new_[26612]_ ) & (~\new_[22830]_  | ~\new_[26612]_ );
  assign \new_[11678]_  = (~\m7_data_i[11]  | ~\new_[18832]_ ) & (~\m0_data_i[11]  | ~\new_[18066]_ );
  assign \new_[11679]_  = (~\m5_data_i[11]  | ~\new_[20542]_ ) & (~\m6_data_i[11]  | ~\new_[16289]_ );
  assign \new_[11680]_  = (~\m7_data_i[10]  | ~\new_[18832]_ ) & (~\m0_data_i[10]  | ~\new_[18066]_ );
  assign \new_[11681]_  = (~\m5_data_i[9]  | ~\new_[18743]_ ) & (~\m6_data_i[9]  | ~\new_[16289]_ );
  assign \new_[11682]_  = (~\m7_data_i[9]  | ~\new_[18832]_ ) & (~\m0_data_i[9]  | ~\new_[18066]_ );
  assign \new_[11683]_  = (~\m5_data_i[8]  | ~\new_[18743]_ ) & (~\m6_data_i[8]  | ~\new_[16289]_ );
  assign \new_[11684]_  = (~\new_[16432]_  | ~\new_[30403]_ ) & (~\new_[24216]_  | ~\new_[30403]_ );
  assign \new_[11685]_  = (~\m7_data_i[8]  | ~\new_[18832]_ ) & (~\m0_data_i[8]  | ~\new_[18066]_ );
  assign \new_[11686]_  = (~\m5_data_i[7]  | ~\new_[18744]_ ) & (~\m6_data_i[7]  | ~\new_[16289]_ );
  assign \new_[11687]_  = (~\new_[16435]_  | ~\new_[29170]_ ) & (~\new_[27501]_  | ~\new_[29170]_ );
  assign \new_[11688]_  = (~\m5_data_i[6]  | ~\new_[20542]_ ) & (~\m6_data_i[6]  | ~\new_[16289]_ );
  assign \new_[11689]_  = (~\m5_data_i[5]  | ~\new_[18743]_ ) & (~\m6_data_i[5]  | ~\new_[16289]_ );
  assign \new_[11690]_  = (~\m7_data_i[4]  | ~\new_[18832]_ ) & (~\m0_data_i[4]  | ~\new_[18066]_ );
  assign \new_[11691]_  = (~\m5_data_i[4]  | ~\new_[18744]_ ) & (~\m6_data_i[4]  | ~\new_[16289]_ );
  assign \new_[11692]_  = (~\m7_data_i[3]  | ~\new_[18832]_ ) & (~\m0_data_i[3]  | ~\new_[18066]_ );
  assign \new_[11693]_  = (~\m5_data_i[3]  | ~\new_[18744]_ ) & (~\m6_data_i[3]  | ~\new_[16289]_ );
  assign \new_[11694]_  = (~\new_[16442]_  | ~\new_[29257]_ ) & (~\new_[22810]_  | ~\new_[29257]_ );
  assign \new_[11695]_  = (~m7_we_i | ~\new_[18115]_ ) & (~m0_we_i | ~\new_[18932]_ );
  assign \new_[11696]_  = (~\m5_data_i[21]  | ~\new_[18752]_ ) & (~\m6_data_i[21]  | ~\new_[18787]_ );
  assign \new_[11697]_  = (~\m7_data_i[1]  | ~\new_[18832]_ ) & (~\m0_data_i[1]  | ~\new_[18066]_ );
  assign \new_[11698]_  = (~\m7_data_i[0]  | ~\new_[18832]_ ) & (~\m0_data_i[0]  | ~\new_[18066]_ );
  assign \new_[11699]_  = (~\new_[16447]_  | ~\new_[29696]_ ) & (~\new_[24113]_  | ~\new_[29696]_ );
  assign \new_[11700]_  = (~\m5_data_i[0]  | ~\new_[18743]_ ) & (~\m6_data_i[0]  | ~\new_[16289]_ );
  assign \new_[11701]_  = (~\new_[18832]_  | ~\new_[31496]_ ) & (~\new_[18066]_  | ~\m0_addr_i[31] );
  assign \new_[11702]_  = (~\new_[16289]_  | ~\m6_addr_i[31] ) & (~\new_[20542]_  | ~\new_[31001]_ );
  assign \new_[11703]_  = (~\new_[16289]_  | ~\m6_addr_i[30] ) & (~\new_[18743]_  | ~\new_[31147]_ );
  assign \new_[11704]_  = (~\new_[18832]_  | ~\new_[31885]_ ) & (~\new_[18066]_  | ~\new_[31292]_ );
  assign \new_[11705]_  = (~\new_[16449]_  | ~\new_[29958]_ ) & (~\new_[26171]_  | ~\new_[29958]_ );
  assign \new_[11706]_  = (~\new_[16289]_  | ~\m6_addr_i[29] ) & (~\new_[18743]_  | ~\new_[31407]_ );
  assign \new_[11707]_  = (~\m5_data_i[11]  | ~\new_[18738]_ ) & (~\m6_data_i[11]  | ~\new_[18031]_ );
  assign \new_[11708]_  = (~\new_[18832]_  | ~\new_[30577]_ ) & (~\new_[18066]_  | ~\new_[30957]_ );
  assign \new_[11709]_  = (~\new_[16289]_  | ~\m6_addr_i[28] ) & (~\new_[20542]_  | ~\new_[31276]_ );
  assign \new_[11710]_  = (~\new_[18832]_  | ~\m7_addr_i[27] ) & (~\new_[18066]_  | ~\m0_addr_i[27] );
  assign \new_[11711]_  = (~\new_[16289]_  | ~\m6_addr_i[27] ) & (~\new_[20542]_  | ~\m5_addr_i[27] );
  assign \new_[11712]_  = (~\new_[16454]_  | ~\new_[29635]_ ) & (~\new_[25095]_  | ~\new_[29635]_ );
  assign \new_[11713]_  = (~\new_[16289]_  | ~\m6_addr_i[26] ) & (~\new_[18743]_  | ~\m5_addr_i[26] );
  assign \new_[11714]_  = (~\new_[18832]_  | ~\m7_addr_i[26] ) & (~\new_[18066]_  | ~\m0_addr_i[26] );
  assign \new_[11715]_  = (~\new_[18832]_  | ~\m7_addr_i[25] ) & (~\new_[18066]_  | ~\m0_addr_i[25] );
  assign \new_[11716]_  = (~\new_[16289]_  | ~\m6_addr_i[25] ) & (~\new_[20542]_  | ~\m5_addr_i[25] );
  assign \new_[11717]_  = (~\new_[18832]_  | ~\m7_addr_i[24] ) & (~\new_[18066]_  | ~\m0_addr_i[24] );
  assign \new_[11718]_  = (~\new_[16289]_  | ~\m6_addr_i[24] ) & (~\new_[20542]_  | ~\m5_addr_i[24] );
  assign \new_[11719]_  = (~\m7_addr_i[23]  | ~\new_[18832]_ ) & (~\m0_addr_i[23]  | ~\new_[18066]_ );
  assign \new_[11720]_  = (~\m5_addr_i[22]  | ~\new_[20542]_ ) & (~\m6_addr_i[22]  | ~\new_[16289]_ );
  assign \new_[11721]_  = (~\m7_addr_i[22]  | ~\new_[18832]_ ) & (~\m0_addr_i[22]  | ~\new_[18066]_ );
  assign \new_[11722]_  = (~\new_[16458]_  | ~\new_[29570]_ ) & (~\new_[24219]_  | ~\new_[29570]_ );
  assign \new_[11723]_  = (~\m7_addr_i[21]  | ~\new_[18832]_ ) & (~\m0_addr_i[21]  | ~\new_[18066]_ );
  assign \new_[11724]_  = (~\m4_addr_i[21]  | ~\new_[17268]_ ) & (~\m3_addr_i[21]  | ~\new_[19597]_ );
  assign \new_[11725]_  = (~\m5_addr_i[21]  | ~\new_[18744]_ ) & (~\m6_addr_i[21]  | ~\new_[16289]_ );
  assign \new_[11726]_  = (~\m5_addr_i[20]  | ~\new_[20542]_ ) & (~\m6_addr_i[20]  | ~\new_[16289]_ );
  assign \new_[11727]_  = (~\m7_addr_i[20]  | ~\new_[18832]_ ) & (~\m0_addr_i[20]  | ~\new_[18066]_ );
  assign \new_[11728]_  = (~\new_[16459]_  | ~\new_[29379]_ ) & (~\new_[22795]_  | ~\new_[29379]_ );
  assign \new_[11729]_  = (~\m7_addr_i[19]  | ~\new_[18832]_ ) & (~\m0_addr_i[19]  | ~\new_[18066]_ );
  assign \new_[11730]_  = (~\m5_addr_i[19]  | ~\new_[18744]_ ) & (~\m6_addr_i[19]  | ~\new_[16289]_ );
  assign \new_[11731]_  = (~\m4_addr_i[19]  | ~\new_[17268]_ ) & (~\m3_addr_i[19]  | ~\new_[18854]_ );
  assign \new_[11732]_  = (~\m5_addr_i[18]  | ~\new_[20542]_ ) & (~\m6_addr_i[18]  | ~\new_[16289]_ );
  assign \new_[11733]_  = (~\m7_addr_i[18]  | ~\new_[18832]_ ) & (~\m0_addr_i[18]  | ~\new_[18066]_ );
  assign \new_[11734]_  = (~\m5_addr_i[17]  | ~\new_[20542]_ ) & (~\m6_addr_i[17]  | ~\new_[16289]_ );
  assign \new_[11735]_  = (~\m7_addr_i[17]  | ~\new_[18832]_ ) & (~\m0_addr_i[17]  | ~\new_[18066]_ );
  assign \new_[11736]_  = (~\m7_addr_i[16]  | ~\new_[18832]_ ) & (~\m0_addr_i[16]  | ~\new_[18066]_ );
  assign \new_[11737]_  = (~\m4_addr_i[16]  | ~\new_[17268]_ ) & (~\m3_addr_i[16]  | ~\new_[18854]_ );
  assign \new_[11738]_  = (~\m5_addr_i[16]  | ~\new_[18744]_ ) & (~\m6_addr_i[16]  | ~\new_[16289]_ );
  assign \new_[11739]_  = (~\m7_addr_i[15]  | ~\new_[18832]_ ) & (~\m0_addr_i[15]  | ~\new_[18066]_ );
  assign \new_[11740]_  = (~\m4_addr_i[15]  | ~\new_[17268]_ ) & (~\m3_addr_i[15]  | ~\new_[18854]_ );
  assign \new_[11741]_  = (~\m7_data_i[23]  | ~\new_[18106]_ ) & (~\m0_data_i[23]  | ~\new_[18026]_ );
  assign \new_[11742]_  = (~\m5_addr_i[15]  | ~\new_[18744]_ ) & (~\m6_addr_i[15]  | ~\new_[16289]_ );
  assign \new_[11743]_  = (~\m7_addr_i[14]  | ~\new_[18832]_ ) & (~\m0_addr_i[14]  | ~\new_[18066]_ );
  assign \new_[11744]_  = (~\m4_addr_i[14]  | ~\new_[17268]_ ) & (~\m3_addr_i[14]  | ~\new_[18854]_ );
  assign \new_[11745]_  = (~\m5_addr_i[14]  | ~\new_[18744]_ ) & (~\m6_addr_i[14]  | ~\new_[16289]_ );
  assign \new_[11746]_  = (~\new_[16373]_  | ~\new_[29549]_ ) & (~\new_[21438]_  | ~\new_[29549]_ );
  assign \new_[11747]_  = (~\m7_addr_i[13]  | ~\new_[18832]_ ) & (~\m0_addr_i[13]  | ~\new_[18066]_ );
  assign \new_[11748]_  = (~\new_[18098]_  | ~\m7_addr_i[25] ) & (~\new_[18026]_  | ~\m0_addr_i[25] );
  assign \new_[11749]_  = (~\m4_addr_i[13]  | ~\new_[17268]_ ) & (~\m3_addr_i[13]  | ~\new_[19597]_ );
  assign \new_[11750]_  = (~\m5_addr_i[13]  | ~\new_[18744]_ ) & (~\m6_addr_i[13]  | ~\new_[16289]_ );
  assign \new_[11751]_  = (~\m7_addr_i[2]  | ~\new_[18115]_ ) & (~\m0_addr_i[2]  | ~\new_[18932]_ );
  assign \new_[11752]_  = (~\m7_addr_i[12]  | ~\new_[18832]_ ) & (~\m0_addr_i[12]  | ~\new_[18066]_ );
  assign \new_[11753]_  = (~\new_[16374]_  | ~\new_[27816]_ ) & (~\new_[24227]_  | ~\new_[27816]_ );
  assign \new_[11754]_  = (~\m5_addr_i[12]  | ~\new_[18744]_ ) & (~\m6_addr_i[12]  | ~\new_[16289]_ );
  assign \new_[11755]_  = (~\m2_data_i[28]  | ~\new_[18077]_ ) & (~\m1_data_i[28]  | ~\new_[19632]_ );
  assign \new_[11756]_  = (~\m7_addr_i[11]  | ~\new_[18832]_ ) & (~\m0_addr_i[11]  | ~\new_[18066]_ );
  assign \new_[11757]_  = (~\m5_addr_i[11]  | ~\new_[18744]_ ) & (~\m6_addr_i[11]  | ~\new_[16289]_ );
  assign \new_[11758]_  = (~\m7_addr_i[10]  | ~\new_[18832]_ ) & (~\m0_addr_i[10]  | ~\new_[18066]_ );
  assign \new_[11759]_  = (~\new_[16375]_  | ~\new_[29084]_ ) & (~\new_[24202]_  | ~\new_[29084]_ );
  assign \new_[11760]_  = (~\m4_addr_i[10]  | ~\new_[17268]_ ) & (~\m3_addr_i[10]  | ~\new_[19597]_ );
  assign \new_[11761]_  = (~\m7_data_i[21]  | ~\new_[18103]_ ) & (~\m0_data_i[21]  | ~\new_[18026]_ );
  assign \new_[11762]_  = (~\m5_addr_i[10]  | ~\new_[18744]_ ) & (~\m6_addr_i[10]  | ~\new_[16289]_ );
  assign \new_[11763]_  = (~\m7_sel_i[0]  | ~\new_[18115]_ ) & (~\m0_sel_i[0]  | ~\new_[19637]_ );
  assign \new_[11764]_  = (~\new_[16376]_  | ~\new_[29871]_ ) & (~\new_[22803]_  | ~\new_[29871]_ );
  assign \new_[11765]_  = (~\m7_addr_i[9]  | ~\new_[18832]_ ) & (~\m0_addr_i[9]  | ~\new_[18066]_ );
  assign \new_[11766]_  = (~\m5_addr_i[9]  | ~\new_[18744]_ ) & (~\m6_addr_i[9]  | ~\new_[16289]_ );
  assign \new_[11767]_  = ~\new_[28913]_  & (~\new_[16515]_  | ~\new_[19429]_ );
  assign \new_[11768]_  = (~\m7_addr_i[8]  | ~\new_[18832]_ ) & (~\m0_addr_i[8]  | ~\new_[18066]_ );
  assign \new_[11769]_  = (~\new_[16377]_  | ~\new_[28897]_ ) & (~\new_[22577]_  | ~\new_[28897]_ );
  assign \new_[11770]_  = (~\m5_addr_i[8]  | ~\new_[18743]_ ) & (~\m6_addr_i[8]  | ~\new_[16289]_ );
  assign \new_[11771]_  = (~\m7_addr_i[7]  | ~\new_[18832]_ ) & (~\m0_addr_i[7]  | ~\new_[18066]_ );
  assign \new_[11772]_  = (~\m5_addr_i[7]  | ~\new_[18743]_ ) & (~\m6_addr_i[7]  | ~\new_[16289]_ );
  assign \new_[11773]_  = ~\new_[13539]_ ;
  assign \new_[11774]_  = (~\m7_addr_i[6]  | ~\new_[18832]_ ) & (~\m0_addr_i[6]  | ~\new_[18066]_ );
  assign \new_[11775]_  = (~\m5_addr_i[6]  | ~\new_[18744]_ ) & (~\m6_addr_i[6]  | ~\new_[16289]_ );
  assign \new_[11776]_  = (~\m7_addr_i[5]  | ~\new_[18832]_ ) & (~\new_[31848]_  | ~\new_[18066]_ );
  assign \new_[11777]_  = (~\m5_addr_i[5]  | ~\new_[18744]_ ) & (~\m6_addr_i[5]  | ~\new_[16289]_ );
  assign \new_[11778]_  = (~\m7_data_i[28]  | ~\new_[18104]_ ) & (~\m0_data_i[28]  | ~\new_[18026]_ );
  assign \new_[11779]_  = (~\m7_addr_i[4]  | ~\new_[18832]_ ) & (~\m0_addr_i[4]  | ~\new_[18066]_ );
  assign \new_[11780]_  = (~\m5_addr_i[4]  | ~\new_[18744]_ ) & (~\m6_addr_i[4]  | ~\new_[16289]_ );
  assign \new_[11781]_  = (~\new_[31726]_  | ~\new_[18832]_ ) & (~\m0_addr_i[3]  | ~\new_[18066]_ );
  assign \new_[11782]_  = (~\m5_addr_i[3]  | ~\new_[18744]_ ) & (~\m6_addr_i[3]  | ~\new_[16289]_ );
  assign \new_[11783]_  = (~\m7_addr_i[2]  | ~\new_[18832]_ ) & (~\m0_addr_i[2]  | ~\new_[18066]_ );
  assign \new_[11784]_  = (~\m5_addr_i[2]  | ~\new_[18744]_ ) & (~\m6_addr_i[2]  | ~\new_[16289]_ );
  assign \new_[11785]_  = (~\m7_addr_i[1]  | ~\new_[18832]_ ) & (~\m0_addr_i[1]  | ~\new_[18066]_ );
  assign \new_[11786]_  = (~\new_[16383]_  | ~\new_[29937]_ ) & (~\new_[24222]_  | ~\new_[29937]_ );
  assign \new_[11787]_  = (~\m4_addr_i[1]  | ~\new_[17268]_ ) & (~\m3_addr_i[1]  | ~\new_[19597]_ );
  assign \new_[11788]_  = (~\m5_addr_i[1]  | ~\new_[18744]_ ) & (~\m6_addr_i[1]  | ~\new_[16289]_ );
  assign \new_[11789]_  = (~\m7_addr_i[0]  | ~\new_[18832]_ ) & (~\m0_addr_i[0]  | ~\new_[18066]_ );
  assign \new_[11790]_  = (~\m7_sel_i[3]  | ~\new_[18832]_ ) & (~\m0_sel_i[3]  | ~\new_[18066]_ );
  assign \new_[11791]_  = (~\new_[16385]_  | ~\new_[29334]_ ) & (~\new_[22715]_  | ~\new_[29334]_ );
  assign \new_[11792]_  = (~\m4_sel_i[3]  | ~\new_[17268]_ ) & (~\m3_sel_i[3]  | ~\new_[18854]_ );
  assign \new_[11793]_  = (~\m5_sel_i[3]  | ~\new_[18744]_ ) & (~\m6_sel_i[3]  | ~\new_[16289]_ );
  assign \new_[11794]_  = (~\m7_sel_i[2]  | ~\new_[18832]_ ) & (~\m0_sel_i[2]  | ~\new_[18066]_ );
  assign \new_[11795]_  = (~\m4_sel_i[2]  | ~\new_[17268]_ ) & (~\m3_sel_i[2]  | ~\new_[18854]_ );
  assign \new_[11796]_  = (~\m7_data_i[16]  | ~\new_[18099]_ ) & (~\m0_data_i[16]  | ~\new_[18026]_ );
  assign \new_[11797]_  = (~\new_[16386]_  | ~\new_[29358]_ ) & (~\new_[21446]_  | ~\new_[29358]_ );
  assign \new_[11798]_  = (~\m5_sel_i[2]  | ~\new_[18744]_ ) & (~\m6_sel_i[2]  | ~\new_[16289]_ );
  assign \new_[11799]_  = (~\new_[16387]_  | ~\new_[29378]_ ) & (~\new_[22772]_  | ~\new_[29378]_ );
  assign \new_[11800]_  = (~\m7_sel_i[1]  | ~\new_[18832]_ ) & (~\m0_sel_i[1]  | ~\new_[18066]_ );
  assign \new_[11801]_  = (~\m5_sel_i[1]  | ~\new_[18744]_ ) & (~\m6_sel_i[1]  | ~\new_[16289]_ );
  assign \new_[11802]_  = (~\m7_sel_i[0]  | ~\new_[18832]_ ) & (~\m0_sel_i[0]  | ~\new_[18066]_ );
  assign \new_[11803]_  = (~\m4_sel_i[0]  | ~\new_[17268]_ ) & (~\m3_sel_i[0]  | ~\new_[19597]_ );
  assign \new_[11804]_  = (~\m5_sel_i[0]  | ~\new_[18744]_ ) & (~\m6_sel_i[0]  | ~\new_[16289]_ );
  assign \new_[11805]_  = (~m5_we_i | ~\new_[18744]_ ) & (~m6_we_i | ~\new_[16289]_ );
  assign \new_[11806]_  = (~\m4_addr_i[2]  | ~\new_[18155]_ ) & (~\m3_addr_i[2]  | ~\new_[18130]_ );
  assign \new_[11807]_  = (~\new_[16390]_  | ~\new_[29548]_ ) & (~\new_[24060]_  | ~\new_[29548]_ );
  assign \new_[11808]_  = (~\new_[18155]_  | ~\m4_addr_i[25] ) & (~\new_[18130]_  | ~\m3_addr_i[25] );
  assign \new_[11809]_  = (~\m4_data_i[31]  | ~\new_[17263]_ ) & (~\m3_data_i[31]  | ~\new_[17247]_ );
  assign \new_[11810]_  = (~\m2_addr_i[23]  | ~\new_[18078]_ ) & (~\m1_addr_i[23]  | ~\new_[19632]_ );
  assign \new_[11811]_  = (~\m4_data_i[28]  | ~\new_[16306]_ ) & (~\m3_data_i[28]  | ~\new_[18846]_ );
  assign \new_[11812]_  = (~\new_[16391]_  | ~\new_[27777]_ ) & (~\new_[24191]_  | ~\new_[27777]_ );
  assign \new_[11813]_  = (~\m4_data_i[26]  | ~\new_[17263]_ ) & (~\m3_data_i[26]  | ~\new_[18125]_ );
  assign \new_[11814]_  = ~\new_[15278]_  | ~\new_[28961]_ ;
  assign \new_[11815]_  = (~\m4_data_i[24]  | ~\new_[17263]_ ) & (~\m3_data_i[24]  | ~\new_[17247]_ );
  assign \new_[11816]_  = ~\new_[15293]_  | ~\new_[29616]_ ;
  assign \new_[11817]_  = ~\new_[15305]_  | ~\new_[28246]_ ;
  assign \new_[11818]_  = (~\m4_data_i[22]  | ~\new_[16306]_ ) & (~\m3_data_i[22]  | ~\new_[18846]_ );
  assign \new_[11819]_  = ~\new_[15313]_  | ~\new_[29858]_ ;
  assign \new_[11820]_  = (~\m2_data_i[0]  | ~\new_[18068]_ ) & (~\m1_data_i[0]  | ~\new_[18901]_ );
  assign \new_[11821]_  = ~\new_[15320]_  | ~\new_[28082]_ ;
  assign \new_[11822]_  = (~\m5_addr_i[23]  | ~\new_[17202]_ ) & (~\m4_addr_i[23]  | ~\new_[17270]_ );
  assign \new_[11823]_  = ~\new_[15338]_  | ~\new_[28243]_ ;
  assign \new_[11824]_  = ~\new_[15345]_  | ~\new_[29001]_ ;
  assign \new_[11825]_  = (~\m7_data_i[29]  | ~\new_[18100]_ ) & (~\m0_data_i[29]  | ~\new_[18026]_ );
  assign \new_[11826]_  = ~\new_[15360]_  | ~\new_[28728]_ ;
  assign \new_[11827]_  = ~\new_[15388]_  | ~\new_[28224]_ ;
  assign \new_[11828]_  = ~\new_[15373]_  | ~\new_[27996]_ ;
  assign \new_[11829]_  = (~\m4_data_i[19]  | ~\new_[16306]_ ) & (~\m3_data_i[19]  | ~\new_[17247]_ );
  assign \new_[11830]_  = ~\new_[21516]_  | ~\new_[26570]_  | ~\new_[16627]_ ;
  assign \new_[11831]_  = ~\new_[15264]_  | ~\new_[28555]_ ;
  assign \new_[11832]_  = (~\m4_data_i[18]  | ~\new_[17263]_ ) & (~\m3_data_i[18]  | ~\new_[17246]_ );
  assign \new_[11833]_  = (~\m2_addr_i[19]  | ~\new_[18067]_ ) & (~\m1_addr_i[19]  | ~\new_[20573]_ );
  assign \new_[11834]_  = \new_[15572]_  | \new_[25439]_ ;
  assign \new_[11835]_  = \new_[15573]_  | \new_[27572]_ ;
  assign \new_[11836]_  = (~\m4_data_i[15]  | ~\new_[16306]_ ) & (~\m3_data_i[15]  | ~\new_[17245]_ );
  assign \new_[11837]_  = (~\m4_data_i[14]  | ~\new_[16306]_ ) & (~\m3_data_i[14]  | ~\new_[17247]_ );
  assign \new_[11838]_  = ~\new_[15276]_  | ~\new_[28722]_ ;
  assign \new_[11839]_  = \new_[15577]_  | \new_[24761]_ ;
  assign \new_[11840]_  = \new_[15578]_  | \new_[27615]_ ;
  assign \new_[11841]_  = ~\new_[15474]_  | ~\new_[28210]_ ;
  assign \new_[11842]_  = (~\m2_data_i[29]  | ~\new_[18077]_ ) & (~\m1_data_i[29]  | ~\new_[18181]_ );
  assign \new_[11843]_  = \new_[15583]_  | \new_[23162]_ ;
  assign \new_[11844]_  = \new_[15585]_  | \new_[26409]_ ;
  assign \new_[11845]_  = ~\new_[15500]_  | ~\new_[28167]_ ;
  assign \new_[11846]_  = (~\m4_data_i[10]  | ~\new_[16306]_ ) & (~\m3_data_i[10]  | ~\new_[17247]_ );
  assign \new_[11847]_  = (~\m5_data_i[17]  | ~\new_[18756]_ ) & (~\m6_data_i[17]  | ~\new_[17213]_ );
  assign \new_[11848]_  = ~\new_[15915]_  | ~\new_[28091]_  | ~\new_[22657]_ ;
  assign \new_[11849]_  = \new_[15590]_  | \new_[26405]_ ;
  assign \new_[11850]_  = (~\m4_data_i[9]  | ~\new_[16306]_ ) & (~\m3_data_i[9]  | ~\new_[17247]_ );
  assign \new_[11851]_  = \new_[15591]_  | \new_[24744]_ ;
  assign \new_[11852]_  = ~\new_[20612]_  | ~\new_[26549]_  | ~\new_[16562]_ ;
  assign \new_[11853]_  = (~\m7_sel_i[1]  | ~\new_[18115]_ ) & (~\m0_sel_i[1]  | ~\new_[18932]_ );
  assign \new_[11854]_  = ~\new_[28266]_  | ~\new_[26375]_  | ~\new_[16563]_ ;
  assign \new_[11855]_  = (~\m4_data_i[8]  | ~\new_[17263]_ ) & (~\m3_data_i[8]  | ~\new_[17246]_ );
  assign \new_[11856]_  = ~\new_[20612]_  | ~\new_[26549]_  | ~\new_[16626]_ ;
  assign \new_[11857]_  = ~\new_[15503]_  | ~\new_[26607]_ ;
  assign \new_[11858]_  = (~\m4_data_i[7]  | ~\new_[16306]_ ) & (~\m3_data_i[7]  | ~\new_[18846]_ );
  assign \new_[11859]_  = ~\new_[15916]_  | ~\new_[28144]_  | ~\new_[22735]_ ;
  assign \new_[11860]_  = (~\m7_data_i[8]  | ~\new_[18110]_ ) & (~\m0_data_i[8]  | ~\new_[18026]_ );
  assign \new_[11861]_  = (~\m4_data_i[5]  | ~\new_[17263]_ ) & (~\m3_data_i[5]  | ~\new_[17245]_ );
  assign \new_[11862]_  = ~\new_[15505]_  | ~\new_[28164]_ ;
  assign \new_[11863]_  = \new_[15602]_  | \new_[25127]_ ;
  assign \new_[11864]_  = (~\m4_data_i[4]  | ~\new_[17263]_ ) & (~\m3_data_i[4]  | ~\new_[18125]_ );
  assign \new_[11865]_  = (~\m2_data_i[18]  | ~\new_[18077]_ ) & (~\m1_data_i[18]  | ~\new_[18189]_ );
  assign \new_[11866]_  = (~\m4_data_i[3]  | ~\new_[16306]_ ) & (~\m3_data_i[3]  | ~\new_[17247]_ );
  assign \new_[11867]_  = \new_[15603]_  | \new_[27581]_ ;
  assign \new_[11868]_  = (~\m4_data_i[2]  | ~\new_[17263]_ ) & (~\m3_data_i[2]  | ~\new_[17247]_ );
  assign \new_[11869]_  = \new_[15609]_  | \new_[24511]_ ;
  assign \new_[11870]_  = (~\new_[31726]_  | ~\new_[18115]_ ) & (~\m0_addr_i[3]  | ~\new_[18932]_ );
  assign \new_[11871]_  = \new_[15610]_  | \new_[26393]_ ;
  assign \new_[11872]_  = (~\m7_addr_i[20]  | ~\new_[18109]_ ) & (~\m0_addr_i[20]  | ~\new_[18026]_ );
  assign \new_[11873]_  = (~\m4_data_i[1]  | ~\new_[17263]_ ) & (~\m3_data_i[1]  | ~\new_[17245]_ );
  assign \new_[11874]_  = (~\new_[16306]_  | ~\m4_addr_i[31] ) & (~\new_[18846]_  | ~\m3_addr_i[31] );
  assign \new_[11875]_  = \new_[15612]_  | \new_[26561]_ ;
  assign \new_[11876]_  = \new_[15615]_  | \new_[27965]_ ;
  assign \new_[11877]_  = (~\new_[17263]_  | ~\m4_addr_i[30] ) & (~\new_[17245]_  | ~\m3_addr_i[30] );
  assign \new_[11878]_  = ~\new_[15510]_  | ~\new_[28122]_ ;
  assign \new_[11879]_  = ~\new_[15917]_  | ~\new_[27951]_  | ~\new_[22775]_ ;
  assign \new_[11880]_  = \new_[15617]_  | \new_[24550]_ ;
  assign \new_[11881]_  = (~\m2_data_i[14]  | ~\new_[18078]_ ) & (~\m1_data_i[14]  | ~\new_[18185]_ );
  assign \new_[11882]_  = (~\new_[17263]_  | ~\m4_addr_i[28] ) & (~\new_[17245]_  | ~\m3_addr_i[28] );
  assign \new_[11883]_  = (~\new_[17263]_  | ~\m4_addr_i[27] ) & (~\new_[17245]_  | ~\m3_addr_i[27] );
  assign \new_[11884]_  = \new_[15625]_  | \new_[23997]_ ;
  assign \new_[11885]_  = ~\new_[15918]_  | ~\new_[29460]_  | ~\new_[23941]_ ;
  assign \new_[11886]_  = (~\new_[16306]_  | ~\m4_addr_i[26] ) & (~\new_[18846]_  | ~\m3_addr_i[26] );
  assign \new_[11887]_  = \new_[15628]_  | \new_[26450]_ ;
  assign \new_[11888]_  = (~\new_[17263]_  | ~\m4_addr_i[25] ) & (~\new_[17245]_  | ~\m3_addr_i[25] );
  assign \new_[11889]_  = \new_[15630]_  | \new_[23924]_ ;
  assign \new_[11890]_  = ~\new_[15467]_  | ~\new_[24330]_ ;
  assign \new_[11891]_  = (~\m4_addr_i[23]  | ~\new_[16306]_ ) & (~\m3_addr_i[23]  | ~\new_[18846]_ );
  assign \new_[11892]_  = ~\new_[15525]_  | ~\new_[28297]_ ;
  assign \new_[11893]_  = ~\new_[15356]_  | ~\new_[28477]_ ;
  assign \new_[11894]_  = \new_[15633]_  | \new_[26829]_ ;
  assign \new_[11895]_  = ~\new_[15919]_  | ~\new_[29284]_  | ~\new_[24249]_ ;
  assign \new_[11896]_  = ~\new_[15522]_  | ~\new_[28306]_ ;
  assign \new_[11897]_  = ~\new_[15380]_  | ~\new_[28587]_ ;
  assign \new_[11898]_  = \new_[15642]_  | \new_[24337]_ ;
  assign \new_[11899]_  = (~\m4_addr_i[17]  | ~\new_[16306]_ ) & (~\m3_addr_i[17]  | ~\new_[17247]_ );
  assign \new_[11900]_  = ~\new_[15526]_  | ~\new_[28241]_ ;
  assign \new_[11901]_  = (~\m7_addr_i[17]  | ~\new_[18116]_ ) & (~\m0_addr_i[17]  | ~\new_[18932]_ );
  assign \new_[11902]_  = \new_[15651]_  | \new_[26752]_ ;
  assign \new_[11903]_  = (~\m4_addr_i[15]  | ~\new_[16306]_ ) & (~\m3_addr_i[15]  | ~\new_[17247]_ );
  assign \new_[11904]_  = ~\new_[15471]_  | ~\new_[27544]_ ;
  assign \new_[11905]_  = ~\new_[16567]_  | ~\new_[27620]_  | ~\new_[19403]_ ;
  assign \new_[11906]_  = ~\new_[28271]_  | (~\new_[16546]_  & ~\new_[23170]_ );
  assign \new_[11907]_  = ~\new_[27864]_  & (~\new_[16547]_  | ~\new_[19436]_ );
  assign \new_[11908]_  = ~\new_[30134]_  & (~\new_[16549]_  | ~\new_[23073]_ );
  assign \new_[11909]_  = ~\new_[16550]_  | ~\new_[28527]_  | ~\new_[22824]_ ;
  assign \new_[11910]_  = (~\m4_addr_i[12]  | ~\new_[17263]_ ) & (~\m3_addr_i[12]  | ~\new_[17245]_ );
  assign \new_[11911]_  = ~\new_[16350]_  | ~\new_[15051]_ ;
  assign \new_[11912]_  = ~\new_[28265]_  | (~\new_[16551]_  & ~\new_[24820]_ );
  assign \new_[11913]_  = (~\m4_addr_i[9]  | ~\new_[17263]_ ) & (~\m3_addr_i[9]  | ~\new_[17247]_ );
  assign \new_[11914]_  = (~\m7_data_i[31]  | ~\new_[18112]_ ) & (~\m0_data_i[31]  | ~\new_[18019]_ );
  assign \new_[11915]_  = ~\new_[16353]_  | ~\new_[15055]_ ;
  assign \new_[11916]_  = ~\new_[28209]_  | (~\new_[16553]_  & ~\new_[24839]_ );
  assign \new_[11917]_  = ~\new_[28831]_  & (~\new_[16556]_  | ~\new_[23010]_ );
  assign \new_[11918]_  = (~\m4_addr_i[6]  | ~\new_[17263]_ ) & (~\m3_addr_i[6]  | ~\new_[17247]_ );
  assign \new_[11919]_  = (~\m4_addr_i[5]  | ~\new_[17263]_ ) & (~\m3_addr_i[5]  | ~\new_[17245]_ );
  assign \new_[11920]_  = (~\m4_addr_i[4]  | ~\new_[16306]_ ) & (~\m3_addr_i[4]  | ~\new_[17247]_ );
  assign \new_[11921]_  = ~\new_[16356]_  | ~\new_[15062]_ ;
  assign \new_[11922]_  = ~\new_[28688]_  | (~\new_[16557]_  & ~\new_[24881]_ );
  assign \new_[11923]_  = (~\m7_sel_i[2]  | ~\new_[18116]_ ) & (~\m0_sel_i[2]  | ~\new_[19637]_ );
  assign \new_[11924]_  = (~\m4_addr_i[3]  | ~\new_[17263]_ ) & (~\m3_addr_i[3]  | ~\new_[18846]_ );
  assign \new_[11925]_  = ~\new_[16558]_  | ~\new_[26180]_  | ~\new_[22826]_ ;
  assign \new_[11926]_  = (~\m5_addr_i[2]  | ~\new_[18760]_ ) & (~\m6_addr_i[2]  | ~\new_[16287]_ );
  assign \new_[11927]_  = (~\m4_addr_i[0]  | ~\new_[16306]_ ) & (~\m3_addr_i[0]  | ~\new_[18846]_ );
  assign \new_[11928]_  = ~\new_[28735]_  & (~\new_[16560]_  | ~\new_[23069]_ );
  assign \new_[11929]_  = ~\new_[16561]_  | ~\new_[26298]_  | ~\new_[22645]_ ;
  assign \new_[11930]_  = (~\m4_sel_i[3]  | ~\new_[17263]_ ) & (~\m3_sel_i[3]  | ~\new_[18125]_ );
  assign \new_[11931]_  = (~\m4_sel_i[2]  | ~\new_[17263]_ ) & (~\m3_sel_i[2]  | ~\new_[18125]_ );
  assign \new_[11932]_  = ~\new_[16566]_  | ~\new_[27642]_  | ~\new_[21447]_ ;
  assign \new_[11933]_  = (~\m4_sel_i[0]  | ~\new_[16306]_ ) & (~\m3_sel_i[0]  | ~\new_[18846]_ );
  assign \new_[11934]_  = (~\m5_data_i[27]  | ~\new_[18014]_ ) & (~\m6_data_i[27]  | ~\new_[17229]_ );
  assign \new_[11935]_  = ~\new_[28124]_  & (~\new_[16572]_  | ~\new_[24278]_ );
  assign \new_[11936]_  = (~\m2_data_i[29]  | ~\new_[17222]_ ) & (~\m1_data_i[29]  | ~\new_[17273]_ );
  assign \new_[11937]_  = ~\new_[29805]_  & (~\new_[16576]_  | ~\new_[23095]_ );
  assign \new_[11938]_  = (~\m2_data_i[26]  | ~\new_[17222]_ ) & (~\m1_data_i[26]  | ~\new_[18906]_ );
  assign \new_[11939]_  = ~\new_[28037]_  & (~\new_[16579]_  | ~\new_[23180]_ );
  assign \new_[11940]_  = ~\new_[29364]_  & (~\new_[16581]_  | ~\new_[22671]_ );
  assign \new_[11941]_  = ~\new_[16354]_  | ~\new_[15099]_ ;
  assign \new_[11942]_  = ~\new_[30143]_  & (~\new_[16584]_  | ~\new_[22975]_ );
  assign \new_[11943]_  = ~\new_[16585]_  | ~\new_[27951]_  | ~\new_[22767]_ ;
  assign \new_[11944]_  = ~\new_[16586]_  | ~\new_[26424]_  | ~\new_[22728]_ ;
  assign \new_[11945]_  = ~\new_[16360]_  | ~\new_[15103]_ ;
  assign \new_[11946]_  = ~\new_[28106]_  | (~\new_[16587]_  & ~\new_[25031]_ );
  assign \new_[11947]_  = (~\m7_data_i[1]  | ~\new_[18108]_ ) & (~\m0_data_i[1]  | ~\new_[18026]_ );
  assign \new_[11948]_  = (~\m2_data_i[16]  | ~\new_[17222]_ ) & (~\m1_data_i[16]  | ~\new_[18906]_ );
  assign \new_[11949]_  = ~\new_[16589]_  | ~\new_[29460]_  | ~\new_[24052]_ ;
  assign \new_[11950]_  = ~\new_[16352]_  | ~\new_[15109]_ ;
  assign \new_[11951]_  = ~\new_[30358]_  & (~\new_[16592]_  | ~\new_[20464]_ );
  assign \new_[11952]_  = ~\new_[16593]_  | ~\new_[29413]_  | ~\new_[24229]_ ;
  assign \new_[11953]_  = (~\m7_data_i[12]  | ~\new_[19584]_ ) & (~\m0_data_i[12]  | ~\new_[18026]_ );
  assign \new_[11954]_  = ~\new_[30090]_  & (~\new_[16594]_  | ~\new_[20413]_ );
  assign \new_[11955]_  = ~\new_[27379]_  | (~\new_[16596]_  & ~\new_[23692]_ );
  assign \new_[11956]_  = ~\new_[29236]_  & (~\new_[16597]_  | ~\new_[22866]_ );
  assign \new_[11957]_  = ~\new_[16598]_  | ~\new_[28523]_  | ~\new_[21450]_ ;
  assign \new_[11958]_  = (~\m2_data_i[30]  | ~\new_[18078]_ ) & (~\m1_data_i[30]  | ~\new_[19632]_ );
  assign \new_[11959]_  = ~\new_[16358]_  | ~\new_[15117]_ ;
  assign \new_[11960]_  = ~\new_[28148]_  | (~\new_[16565]_  & ~\new_[25058]_ );
  assign \new_[11961]_  = ~\new_[16601]_  | ~\new_[27694]_  | ~\new_[22768]_ ;
  assign \new_[11962]_  = ~\new_[16602]_  | ~\new_[29284]_  | ~\new_[24079]_ ;
  assign \new_[11963]_  = ~\new_[16604]_  | ~\new_[27578]_  | ~\new_[22845]_ ;
  assign \new_[11964]_  = ~\new_[16605]_  | ~\new_[27741]_  | ~\new_[22737]_ ;
  assign \new_[11965]_  = \new_[6185]_  ? \new_[27997]_  : \new_[16324]_ ;
  assign \new_[11966]_  = (~\m2_data_i[8]  | ~\new_[18068]_ ) & (~\m1_data_i[8]  | ~\new_[20573]_ );
  assign \new_[11967]_  = ~\new_[28044]_  & (~\new_[16610]_  | ~\new_[21568]_ );
  assign \new_[11968]_  = ~\new_[16611]_  | ~\new_[29464]_  | ~\new_[26183]_ ;
  assign \new_[11969]_  = ~\new_[28066]_  & (~\new_[16612]_  | ~\new_[22818]_ );
  assign \new_[11970]_  = (~\new_[18035]_  | ~\m6_addr_i[28] ) & (~\new_[16276]_  | ~\new_[31276]_ );
  assign \new_[11971]_  = \new_[15170]_  | \new_[27372]_ ;
  assign \new_[11972]_  = ~\new_[23103]_  & (~\new_[15949]_  | ~\new_[28522]_ );
  assign \new_[11973]_  = (~\m3_data_i[31]  | ~\new_[32350]_ ) & (~\m2_data_i[31]  | ~\new_[17223]_ );
  assign \new_[11974]_  = ~\new_[26499]_  & (~\new_[15950]_  | ~\new_[28772]_ );
  assign \new_[11975]_  = ~\new_[27363]_  & (~\new_[15951]_  | ~\new_[26362]_ );
  assign \new_[11976]_  = (~\m7_data_i[31]  | ~\new_[17240]_ ) & (~\m6_data_i[31]  | ~\new_[19581]_ );
  assign \new_[11977]_  = (~\m5_data_i[31]  | ~\new_[17202]_ ) & (~\m4_data_i[31]  | ~\new_[16309]_ );
  assign \new_[11978]_  = ~\new_[24682]_  | ~\new_[15053]_ ;
  assign \new_[11979]_  = ~\new_[25193]_  | ~\new_[15059]_ ;
  assign \new_[11980]_  = ~\new_[25173]_  | ~\new_[15065]_ ;
  assign \new_[11981]_  = ~\new_[19386]_  | ~\new_[15072]_ ;
  assign \new_[11982]_  = ~\new_[20373]_  | ~\new_[15081]_ ;
  assign \new_[11983]_  = ~\new_[20375]_  | ~\new_[15088]_ ;
  assign \new_[11984]_  = ~\new_[19396]_  | ~\new_[15094]_ ;
  assign \new_[11985]_  = ~\new_[19399]_  | ~\new_[15100]_ ;
  assign \new_[11986]_  = (~\m3_data_i[30]  | ~\new_[32350]_ ) & (~\m2_data_i[30]  | ~\new_[17223]_ );
  assign \new_[11987]_  = ~\new_[25192]_  | ~\new_[15107]_ ;
  assign \new_[11988]_  = ~\new_[19388]_  | ~\new_[15111]_ ;
  assign \new_[11989]_  = ~\new_[25171]_  | ~\new_[15119]_ ;
  assign \new_[11990]_  = ~\new_[20382]_  | ~\new_[15123]_ ;
  assign \new_[11991]_  = ~\new_[20388]_  | ~\new_[15127]_ ;
  assign \new_[11992]_  = (~\m5_data_i[30]  | ~\new_[18745]_ ) & (~\m4_data_i[30]  | ~\new_[17270]_ );
  assign \new_[11993]_  = ~\new_[29555]_  & (~\new_[16310]_  | ~\new_[21532]_ );
  assign \new_[11994]_  = (~\m2_addr_i[22]  | ~\new_[17222]_ ) & (~\m1_addr_i[22]  | ~\new_[17273]_ );
  assign \new_[11995]_  = ~\new_[23072]_  & (~\new_[16533]_  | ~\new_[20496]_ );
  assign \new_[11996]_  = ~\new_[28647]_  & (~\new_[16521]_  | ~\new_[21523]_ );
  assign \new_[11997]_  = (~\m7_data_i[10]  | ~\new_[18098]_ ) & (~\m0_data_i[10]  | ~\new_[18026]_ );
  assign \new_[11998]_  = (~\m3_data_i[29]  | ~\new_[18936]_ ) & (~\m2_data_i[29]  | ~\new_[18808]_ );
  assign \new_[11999]_  = ~\new_[28673]_  & (~\new_[16335]_  | ~\new_[19448]_ );
  assign \new_[12000]_  = ~\new_[28738]_  & (~\new_[16329]_  | ~\new_[21484]_ );
  assign \new_[12001]_  = (~\m2_addr_i[20]  | ~\new_[17222]_ ) & (~\m1_addr_i[20]  | ~\new_[17273]_ );
  assign \new_[12002]_  = ~\new_[30406]_  & (~\new_[15940]_  | ~\new_[28740]_ );
  assign \new_[12003]_  = (~\m5_data_i[29]  | ~\new_[17203]_ ) & (~\m4_data_i[29]  | ~\new_[16309]_ );
  assign \new_[12004]_  = ~\new_[15052]_  & (~\new_[28992]_  | ~\new_[5895]_ );
  assign \new_[12005]_  = \new_[15140]_  & \new_[27876]_ ;
  assign \new_[12006]_  = (~\m3_data_i[28]  | ~\new_[32350]_ ) & (~\m2_data_i[28]  | ~\new_[17223]_ );
  assign \new_[12007]_  = ~\new_[15057]_  & (~\new_[29541]_  | ~\new_[5896]_ );
  assign \new_[12008]_  = \new_[15148]_  & \new_[27933]_ ;
  assign \new_[12009]_  = ~\new_[28780]_  & (~\new_[15944]_  | ~\new_[28492]_ );
  assign \new_[12010]_  = ~\new_[15064]_  & (~\new_[29217]_  | ~\new_[5897]_ );
  assign \new_[12011]_  = (~\m5_data_i[28]  | ~\new_[17202]_ ) & (~\m4_data_i[28]  | ~\new_[17270]_ );
  assign \new_[12012]_  = \new_[15156]_  & \new_[26748]_ ;
  assign \new_[12013]_  = (~\m2_addr_i[17]  | ~\new_[17222]_ ) & (~\m1_addr_i[17]  | ~\new_[18906]_ );
  assign \new_[12014]_  = (~\m7_data_i[28]  | ~\new_[17240]_ ) & (~\m6_data_i[28]  | ~\new_[18089]_ );
  assign \new_[12015]_  = \new_[15164]_  & \new_[29066]_ ;
  assign \new_[12016]_  = (~\m2_addr_i[16]  | ~\new_[17222]_ ) & (~\m1_addr_i[16]  | ~\new_[18906]_ );
  assign \new_[12017]_  = \new_[15169]_  & \new_[28879]_ ;
  assign \new_[12018]_  = ~\new_[15079]_  & (~\new_[29700]_  | ~\new_[5900]_ );
  assign \new_[12019]_  = (~\m3_data_i[27]  | ~\new_[32350]_ ) & (~\m2_data_i[27]  | ~\new_[17223]_ );
  assign \new_[12020]_  = ~\new_[29584]_  & (~\new_[15952]_  | ~\new_[28048]_ );
  assign \new_[12021]_  = (~\m2_addr_i[15]  | ~\new_[17222]_ ) & (~\m1_addr_i[15]  | ~\new_[17273]_ );
  assign \new_[12022]_  = \new_[15185]_  & \new_[28758]_ ;
  assign \new_[12023]_  = ~\new_[15087]_  & (~\new_[29157]_  | ~\new_[5901]_ );
  assign \new_[12024]_  = (~\m7_data_i[27]  | ~\new_[17240]_ ) & (~\m6_data_i[27]  | ~\new_[19581]_ );
  assign \new_[12025]_  = ~\new_[29446]_  & (~\new_[15954]_  | ~\new_[28559]_ );
  assign \new_[12026]_  = \new_[15191]_  & \new_[29586]_ ;
  assign \new_[12027]_  = (~\m5_data_i[27]  | ~\new_[17202]_ ) & (~\m4_data_i[27]  | ~\new_[16309]_ );
  assign \new_[12028]_  = \new_[15194]_  & \new_[29196]_ ;
  assign \new_[12029]_  = (~\m2_addr_i[13]  | ~\new_[17222]_ ) & (~\m1_addr_i[13]  | ~\new_[17273]_ );
  assign \new_[12030]_  = (~\m3_data_i[26]  | ~\new_[32350]_ ) & (~\m2_data_i[26]  | ~\new_[17223]_ );
  assign \new_[12031]_  = \new_[15203]_  & \new_[26589]_ ;
  assign \new_[12032]_  = ~\new_[15104]_  & (~\new_[29101]_  | ~\new_[5904]_ );
  assign \new_[12033]_  = \new_[15212]_  & \new_[26823]_ ;
  assign \new_[12034]_  = ~\new_[29250]_  & (~\new_[15957]_  | ~\new_[28708]_ );
  assign \new_[12035]_  = \new_[15219]_  & \new_[28030]_ ;
  assign \new_[12036]_  = \new_[15221]_  & \new_[27767]_ ;
  assign \new_[12037]_  = (~\m5_data_i[26]  | ~\new_[17203]_ ) & (~\m4_data_i[26]  | ~\new_[16309]_ );
  assign \new_[12038]_  = ~\new_[15115]_  & (~\new_[29671]_  | ~\new_[5933]_ );
  assign \new_[12039]_  = (~\m2_addr_i[10]  | ~\new_[17222]_ ) & (~\m1_addr_i[10]  | ~\new_[17273]_ );
  assign \new_[12040]_  = ~\new_[29612]_  & (~\new_[15963]_  | ~\new_[28305]_ );
  assign \new_[12041]_  = (~\m5_data_i[25]  | ~\new_[17203]_ ) & (~\m4_data_i[25]  | ~\new_[17270]_ );
  assign \new_[12042]_  = (~\m5_data_i[25]  | ~\new_[18738]_ ) & (~\m6_data_i[25]  | ~\new_[18031]_ );
  assign \new_[12043]_  = ~\new_[15118]_  & (~\new_[29167]_  | ~\new_[5906]_ );
  assign \new_[12044]_  = (~\m3_data_i[25]  | ~\new_[18936]_ ) & (~\m2_data_i[25]  | ~\new_[18808]_ );
  assign \new_[12045]_  = \new_[15238]_  & \new_[27819]_ ;
  assign \new_[12046]_  = ~\new_[26640]_  & (~\new_[15961]_  | ~\new_[28154]_ );
  assign \new_[12047]_  = \new_[15243]_  & \new_[28854]_ ;
  assign \new_[12048]_  = ~\new_[15121]_  & (~\new_[29047]_  | ~\new_[5907]_ );
  assign \new_[12049]_  = ~\new_[29138]_  & (~\new_[15943]_  | ~\new_[28501]_ );
  assign \new_[12050]_  = (~\m2_addr_i[8]  | ~\new_[17222]_ ) & (~\m1_addr_i[8]  | ~\new_[18906]_ );
  assign \new_[12051]_  = ~\new_[15126]_  & (~\new_[29354]_  | ~\new_[5908]_ );
  assign \new_[12052]_  = ~\new_[30073]_  & (~\new_[15964]_  | ~\new_[28475]_ );
  assign \new_[12053]_  = (~\m2_addr_i[7]  | ~\new_[17222]_ ) & (~\m1_addr_i[7]  | ~\new_[17273]_ );
  assign \new_[12054]_  = (~\m7_data_i[25]  | ~\new_[17240]_ ) & (~\m6_data_i[25]  | ~\new_[18089]_ );
  assign \new_[12055]_  = (~\m3_data_i[24]  | ~\new_[32350]_ ) & (~\m2_data_i[24]  | ~\new_[17223]_ );
  assign \new_[12056]_  = ~\new_[15131]_  & (~\new_[29172]_  | ~\new_[5894]_ );
  assign \new_[12057]_  = (~\m2_addr_i[6]  | ~\new_[17222]_ ) & (~\m1_addr_i[6]  | ~\new_[18906]_ );
  assign \new_[12058]_  = ~\new_[26699]_  & (~\new_[15966]_  | ~\new_[22554]_ );
  assign \new_[12059]_  = ~\new_[17527]_  | ~\new_[17528]_  | ~\new_[17526]_  | ~\new_[18465]_ ;
  assign \new_[12060]_  = (~\m5_data_i[24]  | ~\new_[17202]_ ) & (~\m4_data_i[24]  | ~\new_[16309]_ );
  assign \new_[12061]_  = ~\new_[27851]_  & (~\new_[15967]_  | ~\new_[24126]_ );
  assign \new_[12062]_  = ~\new_[26603]_  & (~\new_[15968]_  | ~\new_[26186]_ );
  assign \new_[12063]_  = (~\m3_data_i[23]  | ~\new_[32350]_ ) & (~\m2_data_i[23]  | ~\new_[17223]_ );
  assign \new_[12064]_  = ~\new_[18468]_  | ~\new_[18469]_  | ~\new_[18467]_  | ~\new_[16645]_ ;
  assign \new_[12065]_  = ~\new_[27877]_  & (~\new_[15969]_  | ~\new_[24253]_ );
  assign \new_[12066]_  = (~\m7_data_i[23]  | ~\new_[17240]_ ) & (~\m6_data_i[23]  | ~\new_[18090]_ );
  assign \new_[12067]_  = ~\new_[28024]_  & (~\new_[15984]_  | ~\new_[24370]_ );
  assign \new_[12068]_  = ~\new_[26540]_  & (~\new_[15970]_  | ~\new_[22733]_ );
  assign \new_[12069]_  = (~\m5_data_i[23]  | ~\new_[17202]_ ) & (~\m4_data_i[23]  | ~\new_[16309]_ );
  assign \new_[12070]_  = ~\new_[28661]_  & (~\new_[15971]_  | ~\new_[22748]_ );
  assign \new_[12071]_  = ~\new_[28268]_  & (~\new_[15972]_  | ~\new_[24234]_ );
  assign \new_[12072]_  = (~\m3_data_i[22]  | ~\new_[32350]_ ) & (~\m2_data_i[22]  | ~\new_[17223]_ );
  assign \new_[12073]_  = ~\new_[26781]_  & (~\new_[15973]_  | ~\new_[21421]_ );
  assign \new_[12074]_  = (~\m2_sel_i[3]  | ~\new_[17222]_ ) & (~\m1_sel_i[3]  | ~\new_[18906]_ );
  assign \new_[12075]_  = (~\m5_data_i[22]  | ~\new_[17202]_ ) & (~\m4_data_i[22]  | ~\new_[16309]_ );
  assign \new_[12076]_  = (~\new_[15974]_  | ~\new_[28742]_ ) & (~\new_[24321]_  | ~\new_[28742]_ );
  assign \new_[12077]_  = (~\m7_data_i[22]  | ~\new_[17240]_ ) & (~\m6_data_i[22]  | ~\new_[18090]_ );
  assign \new_[12078]_  = (~\m2_sel_i[1]  | ~\new_[17222]_ ) & (~\m1_sel_i[1]  | ~\new_[17273]_ );
  assign \new_[12079]_  = ~\new_[28737]_  & (~\new_[15975]_  | ~\new_[24209]_ );
  assign \new_[12080]_  = (~\m7_data_i[21]  | ~\new_[17240]_ ) & (~\m6_data_i[21]  | ~\new_[19581]_ );
  assign \new_[12081]_  = (~\m2_sel_i[0]  | ~\new_[17222]_ ) & (~\m1_sel_i[0]  | ~\new_[18906]_ );
  assign \new_[12082]_  = ~\new_[28430]_  & (~\new_[15985]_  | ~\new_[24454]_ );
  assign \new_[12083]_  = ~\new_[26871]_  & (~\new_[15976]_  | ~\new_[22608]_ );
  assign \new_[12084]_  = (~\m5_data_i[20]  | ~\new_[17203]_ ) & (~\m4_data_i[20]  | ~\new_[16309]_ );
  assign \new_[12085]_  = ~\new_[28765]_  & (~\new_[15977]_  | ~\new_[22639]_ );
  assign \new_[12086]_  = (~\m7_data_i[20]  | ~\new_[17240]_ ) & (~\m6_data_i[20]  | ~\new_[19581]_ );
  assign \new_[12087]_  = ~\new_[27702]_  & (~\new_[15979]_  | ~\new_[22615]_ );
  assign \new_[12088]_  = (~\m7_data_i[31]  | ~\new_[19606]_ ) & (~\m0_data_i[31]  | ~\new_[18781]_ );
  assign \new_[12089]_  = ~\new_[18474]_  | ~\new_[17550]_  | ~\new_[17548]_  | ~\new_[17549]_ ;
  assign \new_[12090]_  = (~\m4_data_i[31]  | ~\new_[18156]_ ) & (~\m3_data_i[31]  | ~\new_[18130]_ );
  assign \new_[12091]_  = ~\new_[17551]_  | ~\new_[17552]_  | ~\new_[18470]_  | ~\new_[18475]_ ;
  assign \new_[12092]_  = (~\m7_data_i[30]  | ~\new_[19606]_ ) & (~\m0_data_i[30]  | ~\new_[18781]_ );
  assign \new_[12093]_  = ~\new_[28637]_  & (~\new_[15980]_  | ~\new_[22718]_ );
  assign \new_[12094]_  = ~\new_[28696]_  & (~\new_[15982]_  | ~\new_[24251]_ );
  assign \new_[12095]_  = (~\m4_data_i[29]  | ~\new_[18155]_ ) & (~\m3_data_i[29]  | ~\new_[18130]_ );
  assign \new_[12096]_  = (~\m3_data_i[18]  | ~\new_[32350]_ ) & (~\m2_data_i[18]  | ~\new_[17223]_ );
  assign \new_[12097]_  = (~\m7_data_i[28]  | ~\new_[19606]_ ) & (~\m0_data_i[28]  | ~\new_[18781]_ );
  assign \new_[12098]_  = ~\new_[15443]_  & ~\new_[16532]_ ;
  assign \new_[12099]_  = (~\m5_data_i[18]  | ~\new_[17202]_ ) & (~\m4_data_i[18]  | ~\new_[17270]_ );
  assign \new_[12100]_  = (~\m4_data_i[27]  | ~\new_[18156]_ ) & (~\m3_data_i[27]  | ~\new_[18130]_ );
  assign \new_[12101]_  = ~\new_[27831]_  & (~\new_[15978]_  | ~\new_[22765]_ );
  assign \new_[12102]_  = (~\m5_data_i[17]  | ~\new_[17202]_ ) & (~\m4_data_i[17]  | ~\new_[17270]_ );
  assign \new_[12103]_  = ~\new_[27834]_  & (~\new_[15981]_  | ~\new_[22721]_ );
  assign \new_[12104]_  = (~\m4_data_i[26]  | ~\new_[18157]_ ) & (~\m3_data_i[26]  | ~\new_[18130]_ );
  assign \new_[12105]_  = (~\m7_data_i[26]  | ~\new_[19606]_ ) & (~\m0_data_i[26]  | ~\new_[19557]_ );
  assign \new_[12106]_  = (~\m4_data_i[25]  | ~\new_[18157]_ ) & (~\m3_data_i[25]  | ~\new_[18130]_ );
  assign \new_[12107]_  = ~\new_[16692]_  | ~\new_[16693]_  | ~\new_[16690]_  | ~\new_[16691]_ ;
  assign \new_[12108]_  = (~\m7_data_i[25]  | ~\new_[19606]_ ) & (~\m0_data_i[25]  | ~\new_[19557]_ );
  assign \new_[12109]_  = (~\m7_data_i[24]  | ~\new_[19606]_ ) & (~\m0_data_i[24]  | ~\new_[18781]_ );
  assign \new_[12110]_  = ~\new_[16694]_  | ~\new_[16695]_  | ~\new_[14507]_  | ~\new_[15899]_ ;
  assign \new_[12111]_  = ~\new_[17559]_  | ~\new_[17560]_  | ~\new_[16696]_  | ~\new_[15900]_ ;
  assign \new_[12112]_  = (~\m2_data_i[7]  | ~\new_[18077]_ ) & (~\m1_data_i[7]  | ~\new_[18186]_ );
  assign \new_[12113]_  = (~\m4_data_i[23]  | ~\new_[18155]_ ) & (~\m3_data_i[23]  | ~\new_[18130]_ );
  assign \new_[12114]_  = (~\m7_data_i[22]  | ~\new_[19606]_ ) & (~\m0_data_i[22]  | ~\new_[18781]_ );
  assign \new_[12115]_  = (~\m4_data_i[22]  | ~\new_[18156]_ ) & (~\m3_data_i[22]  | ~\new_[18130]_ );
  assign \new_[12116]_  = (~\m3_data_i[16]  | ~\new_[32350]_ ) & (~\m2_data_i[16]  | ~\new_[17223]_ );
  assign \new_[12117]_  = (~\m4_data_i[21]  | ~\new_[18155]_ ) & (~\m3_data_i[21]  | ~\new_[18130]_ );
  assign \new_[12118]_  = (~\m5_data_i[16]  | ~\new_[17203]_ ) & (~\m4_data_i[16]  | ~\new_[17270]_ );
  assign \new_[12119]_  = (~\m4_data_i[20]  | ~\new_[18155]_ ) & (~\m3_data_i[20]  | ~\new_[18130]_ );
  assign \new_[12120]_  = (~\m7_data_i[15]  | ~\new_[17240]_ ) & (~\m6_data_i[15]  | ~\new_[18090]_ );
  assign \new_[12121]_  = (~\m7_data_i[19]  | ~\new_[19606]_ ) & (~\m0_data_i[19]  | ~\new_[18781]_ );
  assign \new_[12122]_  = (~\m4_data_i[19]  | ~\new_[18155]_ ) & (~\m3_data_i[19]  | ~\new_[18130]_ );
  assign \new_[12123]_  = (~\m3_data_i[15]  | ~\new_[18936]_ ) & (~\m2_data_i[15]  | ~\new_[17224]_ );
  assign \new_[12124]_  = (~\m7_data_i[17]  | ~\new_[19606]_ ) & (~\m0_data_i[17]  | ~\new_[18781]_ );
  assign \new_[12125]_  = (~\m4_data_i[17]  | ~\new_[18155]_ ) & (~\m3_data_i[17]  | ~\new_[18130]_ );
  assign \new_[12126]_  = (~\m7_data_i[16]  | ~\new_[19606]_ ) & (~\m0_data_i[16]  | ~\new_[18781]_ );
  assign \new_[12127]_  = (~\m7_data_i[15]  | ~\new_[19606]_ ) & (~\m0_data_i[15]  | ~\new_[18781]_ );
  assign \new_[12128]_  = (~\m4_data_i[15]  | ~\new_[18156]_ ) & (~\m3_data_i[15]  | ~\new_[18130]_ );
  assign \new_[12129]_  = ~\new_[16699]_  | ~\new_[17561]_  | ~\new_[15906]_  | ~\new_[15907]_ ;
  assign \new_[12130]_  = (~\m3_data_i[9]  | ~\new_[32350]_ ) & (~\m2_data_i[9]  | ~\new_[18808]_ );
  assign \new_[12131]_  = (~\m4_data_i[14]  | ~\new_[18157]_ ) & (~\m3_data_i[14]  | ~\new_[18130]_ );
  assign \new_[12132]_  = (~\m4_data_i[13]  | ~\new_[18155]_ ) & (~\m3_data_i[13]  | ~\new_[18130]_ );
  assign \new_[12133]_  = ~\new_[16702]_  | ~\new_[16704]_  | ~\new_[16703]_  | ~\new_[16701]_ ;
  assign \new_[12134]_  = (~\m5_data_i[9]  | ~\new_[18756]_ ) & (~\m6_data_i[9]  | ~\new_[17213]_ );
  assign \new_[12135]_  = ~\new_[27932]_  & (~\new_[15983]_  | ~\new_[24245]_ );
  assign \new_[12136]_  = (~\m4_data_i[12]  | ~\new_[18156]_ ) & (~\m3_data_i[12]  | ~\new_[18130]_ );
  assign \new_[12137]_  = ~\new_[15265]_  & (~\new_[30145]_  | ~\new_[6174]_ );
  assign \new_[12138]_  = ~\new_[15267]_  & (~\new_[29992]_  | ~\new_[6035]_ );
  assign \new_[12139]_  = (~\m5_data_i[2]  | ~\new_[18752]_ ) & (~\m6_data_i[2]  | ~\new_[17213]_ );
  assign \new_[12140]_  = (~\m4_data_i[11]  | ~\new_[18157]_ ) & (~\m3_data_i[11]  | ~\new_[18130]_ );
  assign \new_[12141]_  = ~\new_[15271]_  & (~\new_[29907]_  | ~\new_[6037]_ );
  assign \new_[12142]_  = (~\m7_data_i[12]  | ~\new_[17240]_ ) & (~\m6_data_i[12]  | ~\new_[19581]_ );
  assign \new_[12143]_  = ~\new_[28263]_  & (~\new_[15936]_  | ~\new_[19431]_ );
  assign \new_[12144]_  = (~\m4_data_i[10]  | ~\new_[18157]_ ) & (~\m3_data_i[10]  | ~\new_[18130]_ );
  assign \new_[12145]_  = ~\new_[15273]_  & (~\new_[29826]_  | ~\new_[6039]_ );
  assign \new_[12146]_  = (~\m3_data_i[12]  | ~\new_[32350]_ ) & (~\m2_data_i[12]  | ~\new_[18808]_ );
  assign \new_[12147]_  = (~\m4_data_i[9]  | ~\new_[18155]_ ) & (~\m3_data_i[9]  | ~\new_[18130]_ );
  assign \new_[12148]_  = ~\new_[15277]_  & (~\new_[29810]_  | ~\new_[6043]_ );
  assign \new_[12149]_  = ~\new_[15281]_  & (~\new_[29848]_  | ~\new_[6044]_ );
  assign \new_[12150]_  = (~\m5_data_i[12]  | ~\new_[17202]_ ) & (~\m4_data_i[12]  | ~\new_[16309]_ );
  assign \new_[12151]_  = (~\m4_data_i[8]  | ~\new_[18157]_ ) & (~\m3_data_i[8]  | ~\new_[18130]_ );
  assign \new_[12152]_  = ~\new_[28913]_  & (~\new_[15937]_  | ~\new_[19443]_ );
  assign \new_[12153]_  = ~\new_[15287]_  & (~\new_[30236]_  | ~\new_[6047]_ );
  assign \new_[12154]_  = (~\m4_data_i[7]  | ~\new_[18155]_ ) & (~\m3_data_i[7]  | ~\new_[18130]_ );
  assign \new_[12155]_  = (~\m7_data_i[6]  | ~\new_[19606]_ ) & (~\m0_data_i[6]  | ~\new_[18781]_ );
  assign \new_[12156]_  = ~\new_[15290]_  & (~\new_[29889]_  | ~\new_[6049]_ );
  assign \new_[12157]_  = (~\m4_data_i[6]  | ~\new_[18156]_ ) & (~\m3_data_i[6]  | ~\new_[18130]_ );
  assign \new_[12158]_  = ~\new_[15297]_  & (~\new_[30733]_  | ~\new_[6053]_ );
  assign \new_[12159]_  = (~\m4_data_i[5]  | ~\new_[18155]_ ) & (~\m3_data_i[5]  | ~\new_[18130]_ );
  assign \new_[12160]_  = (~\m7_data_i[5]  | ~\new_[19606]_ ) & (~\m0_data_i[5]  | ~\new_[18781]_ );
  assign \new_[12161]_  = ~\new_[15304]_  & (~\new_[30033]_  | ~\new_[6197]_ );
  assign \new_[12162]_  = (~\m4_data_i[4]  | ~\new_[18155]_ ) & (~\m3_data_i[4]  | ~\new_[18130]_ );
  assign \new_[12163]_  = ~\new_[15306]_  & (~\new_[30328]_  | ~\new_[6058]_ );
  assign \new_[12164]_  = ~\new_[15310]_  & (~\new_[30718]_  | ~\new_[6195]_ );
  assign \new_[12165]_  = (~\m4_data_i[3]  | ~\new_[18155]_ ) & (~\m3_data_i[3]  | ~\new_[18130]_ );
  assign \new_[12166]_  = ~\new_[29646]_  & (~\new_[16419]_  | ~\new_[24366]_ );
  assign \new_[12167]_  = ~\new_[15315]_  & (~\new_[30251]_  | ~\new_[6063]_ );
  assign \new_[12168]_  = (~\m4_data_i[2]  | ~\new_[18157]_ ) & (~\m3_data_i[2]  | ~\new_[18130]_ );
  assign \new_[12169]_  = (~\m7_data_i[1]  | ~\new_[19606]_ ) & (~\m0_data_i[1]  | ~\new_[18781]_ );
  assign \new_[12170]_  = ~\new_[15318]_  & (~\new_[30326]_  | ~\new_[6194]_ );
  assign \new_[12171]_  = ~\new_[26634]_  & (~\new_[16337]_  | ~\new_[20492]_ );
  assign \new_[12172]_  = (~\m4_data_i[1]  | ~\new_[18156]_ ) & (~\m3_data_i[1]  | ~\new_[18130]_ );
  assign \new_[12173]_  = ~\new_[15322]_  & (~\new_[30308]_  | ~\new_[6068]_ );
  assign \new_[12174]_  = (~\m7_data_i[0]  | ~\new_[19606]_ ) & (~\m0_data_i[0]  | ~\new_[18781]_ );
  assign \new_[12175]_  = (~\m4_data_i[0]  | ~\new_[18156]_ ) & (~\m3_data_i[0]  | ~\new_[18130]_ );
  assign \new_[12176]_  = ~\new_[15326]_  & (~\new_[30375]_  | ~\new_[31400]_ );
  assign \new_[12177]_  = ~\new_[28936]_  & (~\new_[16332]_  | ~\new_[21548]_ );
  assign \new_[12178]_  = (~\new_[18155]_  | ~\m4_addr_i[31] ) & (~\new_[18130]_  | ~\m3_addr_i[31] );
  assign \new_[12179]_  = (~\m5_data_i[9]  | ~\new_[17202]_ ) & (~\m4_data_i[9]  | ~\new_[16309]_ );
  assign \new_[12180]_  = (~\m3_data_i[8]  | ~\new_[32350]_ ) & (~\m2_data_i[8]  | ~\new_[18808]_ );
  assign \new_[12181]_  = ~\new_[15334]_  & (~\new_[30275]_  | ~\new_[6073]_ );
  assign \new_[12182]_  = (~\new_[19606]_  | ~\new_[31885]_ ) & (~\new_[18781]_  | ~\new_[31292]_ );
  assign \new_[12183]_  = ~\new_[15336]_  & (~\new_[29290]_  | ~\new_[6189]_ );
  assign \new_[12184]_  = (~\new_[18157]_  | ~\m4_addr_i[30] ) & (~\new_[18130]_  | ~\m3_addr_i[30] );
  assign \new_[12185]_  = ~\new_[15339]_  & (~\new_[30788]_  | ~\new_[5992]_ );
  assign \new_[12186]_  = ~\new_[15343]_  & (~\new_[29792]_  | ~\new_[6076]_ );
  assign \new_[12187]_  = (~\new_[18155]_  | ~\m4_addr_i[29] ) & (~\new_[18130]_  | ~\m3_addr_i[29] );
  assign \new_[12188]_  = ~\new_[29313]_  & (~\new_[15896]_  | ~\new_[20463]_ );
  assign \new_[12189]_  = (~\m5_data_i[8]  | ~\new_[17202]_ ) & (~\m4_data_i[8]  | ~\new_[16309]_ );
  assign \new_[12190]_  = ~\new_[15348]_  & (~\new_[30121]_  | ~\new_[6077]_ );
  assign \new_[12191]_  = (~\new_[18157]_  | ~\m4_addr_i[28] ) & (~\new_[18130]_  | ~\m3_addr_i[28] );
  assign \new_[12192]_  = (~\m3_data_i[7]  | ~\new_[32350]_ ) & (~\m2_data_i[7]  | ~\new_[18808]_ );
  assign \new_[12193]_  = ~\new_[15358]_  & (~\new_[30151]_  | ~\new_[6079]_ );
  assign \new_[12194]_  = (~\new_[18156]_  | ~\m4_addr_i[27] ) & (~\new_[18130]_  | ~\m3_addr_i[27] );
  assign \new_[12195]_  = ~\new_[15362]_  & (~\new_[29968]_  | ~\new_[6081]_ );
  assign \new_[12196]_  = (~\new_[19606]_  | ~\m7_addr_i[27] ) & (~\new_[20547]_  | ~\m0_addr_i[27] );
  assign \new_[12197]_  = ~\new_[15365]_  & (~\new_[30737]_  | ~\new_[6082]_ );
  assign \new_[12198]_  = (~\new_[18155]_  | ~\m4_addr_i[26] ) & (~\new_[18130]_  | ~\m3_addr_i[26] );
  assign \new_[12199]_  = ~\new_[15369]_  & (~\new_[29997]_  | ~\new_[6186]_ );
  assign \new_[12200]_  = ~\new_[26649]_  & (~\new_[16318]_  | ~\new_[19430]_ );
  assign \new_[12201]_  = ~\new_[15371]_  & (~\new_[28999]_  | ~\new_[6185]_ );
  assign \new_[12202]_  = (~\m7_data_i[27]  | ~\new_[18112]_ ) & (~\m0_data_i[27]  | ~\new_[18019]_ );
  assign \new_[12203]_  = (~\m5_data_i[7]  | ~\new_[17202]_ ) & (~\m4_data_i[7]  | ~\new_[18884]_ );
  assign \new_[12204]_  = ~\new_[15375]_  & (~\new_[30652]_  | ~\new_[6086]_ );
  assign \new_[12205]_  = (~\new_[19606]_  | ~\m7_addr_i[25] ) & (~\new_[20547]_  | ~\m0_addr_i[25] );
  assign \new_[12206]_  = ~\new_[15382]_  & (~\new_[30201]_  | ~\new_[31499]_ );
  assign \new_[12207]_  = (~\new_[19606]_  | ~\m7_addr_i[24] ) & (~\new_[18781]_  | ~\m0_addr_i[24] );
  assign \new_[12208]_  = (~\new_[18157]_  | ~\m4_addr_i[24] ) & (~\new_[18130]_  | ~\m3_addr_i[24] );
  assign \new_[12209]_  = ~\new_[15386]_  & (~\new_[30502]_  | ~\new_[6183]_ );
  assign \new_[12210]_  = ~\new_[15392]_  & (~\new_[30325]_  | ~\new_[6093]_ );
  assign \new_[12211]_  = ~\new_[27874]_  & (~\new_[16328]_  | ~\new_[20456]_ );
  assign \new_[12212]_  = (~\m7_addr_i[23]  | ~\new_[19606]_ ) & (~\m0_addr_i[23]  | ~\new_[19557]_ );
  assign \new_[12213]_  = (~\m4_addr_i[22]  | ~\new_[18155]_ ) & (~\m3_addr_i[22]  | ~\new_[18130]_ );
  assign \new_[12214]_  = ~\new_[15396]_  & (~\new_[30706]_  | ~\new_[6095]_ );
  assign \new_[12215]_  = (~\m3_data_i[6]  | ~\new_[18936]_ ) & (~\m2_data_i[6]  | ~\new_[17224]_ );
  assign \new_[12216]_  = ~\new_[23345]_  & (~\new_[16136]_  | ~\new_[30164]_ );
  assign \new_[12217]_  = (~\m7_addr_i[21]  | ~\new_[19606]_ ) & (~\m0_addr_i[21]  | ~\new_[18781]_ );
  assign \new_[12218]_  = ~\new_[22573]_  & (~\new_[16145]_  | ~\new_[29219]_ );
  assign \new_[12219]_  = (~\m3_data_i[5]  | ~\new_[18936]_ ) & (~\m2_data_i[5]  | ~\new_[18808]_ );
  assign \new_[12220]_  = ~\new_[21222]_  & (~\new_[16147]_  | ~\new_[30426]_ );
  assign \new_[12221]_  = ~\new_[22146]_  & (~\new_[16148]_  | ~\new_[28989]_ );
  assign \new_[12222]_  = (~\m4_addr_i[20]  | ~\new_[18155]_ ) & (~\m3_addr_i[20]  | ~\new_[18130]_ );
  assign \new_[12223]_  = ~\new_[22309]_  & (~\new_[16153]_  | ~\new_[29032]_ );
  assign \new_[12224]_  = (~\m5_data_i[5]  | ~\new_[17202]_ ) & (~\m4_data_i[5]  | ~\new_[18884]_ );
  assign \new_[12225]_  = ~\new_[21194]_  & (~\new_[16154]_  | ~\new_[29401]_ );
  assign \new_[12226]_  = (~\m4_addr_i[19]  | ~\new_[18155]_ ) & (~\m3_addr_i[19]  | ~\new_[18130]_ );
  assign \new_[12227]_  = (~\m7_data_i[4]  | ~\new_[17240]_ ) & (~\m6_data_i[4]  | ~\new_[19581]_ );
  assign \new_[12228]_  = ~\new_[23545]_  & (~\new_[16202]_  | ~\new_[29221]_ );
  assign \new_[12229]_  = ~\new_[22139]_  & (~\new_[16163]_  | ~\new_[29171]_ );
  assign \new_[12230]_  = ~\new_[22358]_  & (~\new_[16174]_  | ~\new_[29082]_ );
  assign \new_[12231]_  = (~\m4_addr_i[17]  | ~\new_[18155]_ ) & (~\m3_addr_i[17]  | ~\new_[18130]_ );
  assign \new_[12232]_  = (~\m7_addr_i[13]  | ~\new_[18100]_ ) & (~\m0_addr_i[13]  | ~\new_[18026]_ );
  assign \new_[12233]_  = (~\m2_data_i[24]  | ~\new_[18078]_ ) & (~\m1_data_i[24]  | ~\new_[19632]_ );
  assign \new_[12234]_  = ~\new_[22361]_  & (~\new_[16181]_  | ~\new_[30034]_ );
  assign \new_[12235]_  = (~\m5_data_i[4]  | ~\new_[17202]_ ) & (~\m4_data_i[4]  | ~\new_[16309]_ );
  assign \new_[12236]_  = (~\m4_addr_i[16]  | ~\new_[18155]_ ) & (~\m3_addr_i[16]  | ~\new_[18130]_ );
  assign \new_[12237]_  = ~\new_[22443]_  & (~\new_[16155]_  | ~\new_[29061]_ );
  assign \new_[12238]_  = ~\new_[23754]_  & (~\new_[16186]_  | ~\new_[29038]_ );
  assign \new_[12239]_  = (~\m4_addr_i[15]  | ~\new_[18155]_ ) & (~\m3_addr_i[15]  | ~\new_[18130]_ );
  assign \new_[12240]_  = ~\new_[22354]_  & (~\new_[16198]_  | ~\new_[28007]_ );
  assign \new_[12241]_  = (~\m7_addr_i[14]  | ~\new_[19606]_ ) & (~\m0_addr_i[14]  | ~\new_[18781]_ );
  assign \new_[12242]_  = (~\m4_addr_i[14]  | ~\new_[18157]_ ) & (~\m3_addr_i[14]  | ~\new_[18130]_ );
  assign \new_[12243]_  = (~\m3_data_i[3]  | ~\new_[32350]_ ) & (~\m2_data_i[3]  | ~\new_[18808]_ );
  assign \new_[12244]_  = ~\new_[23867]_  & (~\new_[16226]_  | ~\new_[28850]_ );
  assign \new_[12245]_  = (~\m5_data_i[3]  | ~\new_[17202]_ ) & (~\m4_data_i[3]  | ~\new_[16309]_ );
  assign \new_[12246]_  = (~\m7_addr_i[12]  | ~\new_[19606]_ ) & (~\m0_addr_i[12]  | ~\new_[18781]_ );
  assign \new_[12247]_  = (~\m4_addr_i[12]  | ~\new_[18156]_ ) & (~\m3_addr_i[12]  | ~\new_[18130]_ );
  assign \new_[12248]_  = ~\new_[28183]_  | ~\new_[15859]_  | ~\new_[30111]_ ;
  assign \new_[12249]_  = (~\m7_addr_i[11]  | ~\new_[19606]_ ) & (~\m0_addr_i[11]  | ~\new_[18781]_ );
  assign \new_[12250]_  = (~\m7_addr_i[10]  | ~\new_[19606]_ ) & (~\m0_addr_i[10]  | ~\new_[18781]_ );
  assign \new_[12251]_  = (~\m4_addr_i[10]  | ~\new_[18155]_ ) & (~\m3_addr_i[10]  | ~\new_[18130]_ );
  assign \new_[12252]_  = ~\new_[29746]_  | ~\new_[15860]_  | ~\new_[30318]_ ;
  assign \new_[12253]_  = (~\m4_addr_i[9]  | ~\new_[18155]_ ) & (~\m3_addr_i[9]  | ~\new_[18130]_ );
  assign \new_[12254]_  = (~\m7_addr_i[9]  | ~\new_[19606]_ ) & (~\m0_addr_i[9]  | ~\new_[18781]_ );
  assign \new_[12255]_  = (~\m3_data_i[1]  | ~\new_[32350]_ ) & (~\m2_data_i[1]  | ~\new_[18808]_ );
  assign \new_[12256]_  = (~\m4_addr_i[8]  | ~\new_[18155]_ ) & (~\m3_addr_i[8]  | ~\new_[18130]_ );
  assign \new_[12257]_  = ~\new_[29251]_  | ~\new_[15861]_  | ~\new_[29780]_ ;
  assign \new_[12258]_  = (~\m4_addr_i[7]  | ~\new_[18155]_ ) & (~\m3_addr_i[7]  | ~\new_[18130]_ );
  assign \new_[12259]_  = (~\m5_data_i[1]  | ~\new_[18745]_ ) & (~\m4_data_i[1]  | ~\new_[17270]_ );
  assign \new_[12260]_  = (~\m7_data_i[0]  | ~\new_[17240]_ ) & (~\m6_data_i[0]  | ~\new_[19581]_ );
  assign \new_[12261]_  = ~\new_[15810]_  & ~\new_[16056]_ ;
  assign \new_[12262]_  = (~\m4_addr_i[6]  | ~\new_[18156]_ ) & (~\m3_addr_i[6]  | ~\new_[18130]_ );
  assign \new_[12263]_  = (~\m4_addr_i[5]  | ~\new_[18156]_ ) & (~\m3_addr_i[5]  | ~\new_[18130]_ );
  assign \new_[12264]_  = ~\new_[30697]_  | ~\new_[15866]_  | ~\new_[30146]_ ;
  assign \new_[12265]_  = (~\m3_data_i[0]  | ~\new_[32350]_ ) & (~\m2_data_i[0]  | ~\new_[18808]_ );
  assign \new_[12266]_  = (~\m5_data_i[0]  | ~\new_[17202]_ ) & (~\m4_data_i[0]  | ~\new_[18884]_ );
  assign \new_[12267]_  = ~\new_[29904]_  | ~\new_[15867]_  | ~\new_[30005]_ ;
  assign \new_[12268]_  = (~\m4_addr_i[4]  | ~\new_[18156]_ ) & (~\m3_addr_i[4]  | ~\new_[18130]_ );
  assign \new_[12269]_  = (~\m4_addr_i[3]  | ~\new_[18155]_ ) & (~\m3_addr_i[3]  | ~\new_[18130]_ );
  assign \new_[12270]_  = ~\new_[15812]_  & ~\new_[16078]_ ;
  assign \new_[12271]_  = ~\new_[29404]_  | ~\new_[15871]_  | ~\new_[30086]_ ;
  assign \new_[12272]_  = (~\new_[17270]_  | ~\m4_addr_i[31] ) & (~\new_[18936]_  | ~\m3_addr_i[31] );
  assign \new_[12273]_  = (~\new_[17223]_  | ~\m2_addr_i[31] ) & (~\new_[17277]_  | ~\new_[31447]_ );
  assign \new_[12274]_  = (~\new_[18067]_  | ~\m2_addr_i[27] ) & (~\new_[20573]_  | ~\m1_addr_i[27] );
  assign \new_[12275]_  = ~\new_[15813]_  & ~\new_[16083]_ ;
  assign \new_[12276]_  = (~\m4_addr_i[1]  | ~\new_[18155]_ ) & (~\m3_addr_i[1]  | ~\new_[18130]_ );
  assign \new_[12277]_  = (~\new_[17223]_  | ~\new_[31486]_ ) & (~\new_[17277]_  | ~\new_[31308]_ );
  assign \new_[12278]_  = (~\m4_addr_i[0]  | ~\new_[18155]_ ) & (~\m3_addr_i[0]  | ~\new_[18130]_ );
  assign \new_[12279]_  = ~\new_[30572]_  | ~\new_[15877]_  | ~\new_[30071]_ ;
  assign \new_[12280]_  = ~\new_[15814]_  & ~\new_[16845]_ ;
  assign \new_[12281]_  = (~\m4_sel_i[2]  | ~\new_[18155]_ ) & (~\m3_sel_i[2]  | ~\new_[18130]_ );
  assign \new_[12282]_  = (~\new_[17270]_  | ~\m4_addr_i[29] ) & (~\new_[32350]_  | ~\m3_addr_i[29] );
  assign \new_[12283]_  = (~\new_[17223]_  | ~\new_[31000]_ ) & (~\new_[18192]_  | ~\new_[31538]_ );
  assign \new_[12284]_  = ~\new_[29299]_  | ~\new_[15884]_  | ~\new_[30180]_ ;
  assign \new_[12285]_  = (~\m4_sel_i[1]  | ~\new_[18155]_ ) & (~\m3_sel_i[1]  | ~\new_[18130]_ );
  assign \new_[12286]_  = (~\new_[17270]_  | ~\m4_addr_i[28] ) & (~\new_[18936]_  | ~\m3_addr_i[28] );
  assign \new_[12287]_  = (~\m7_data_i[3]  | ~\new_[18107]_ ) & (~\m0_data_i[3]  | ~\new_[18026]_ );
  assign \new_[12288]_  = (~\new_[17223]_  | ~\new_[31547]_ ) & (~\new_[17277]_  | ~\new_[31458]_ );
  assign \new_[12289]_  = (~\m4_sel_i[0]  | ~\new_[18156]_ ) & (~\m3_sel_i[0]  | ~\new_[18130]_ );
  assign \new_[12290]_  = (~m7_we_i | ~\new_[19606]_ ) & (~m0_we_i | ~\new_[18781]_ );
  assign \new_[12291]_  = ~\new_[30786]_  | ~\new_[15887]_  | ~\new_[30278]_ ;
  assign \new_[12292]_  = (~\new_[17270]_  | ~\m4_addr_i[27] ) & (~\new_[18936]_  | ~\m3_addr_i[27] );
  assign \new_[12293]_  = (~m4_we_i | ~\new_[18157]_ ) & (~m3_we_i | ~\new_[18130]_ );
  assign \new_[12294]_  = (~\new_[17223]_  | ~\m2_addr_i[27] ) & (~\new_[17277]_  | ~\m1_addr_i[27] );
  assign \new_[12295]_  = ~\new_[15817]_  & ~\new_[16930]_ ;
  assign \new_[12296]_  = (~\new_[17270]_  | ~\m4_addr_i[26] ) & (~\new_[18936]_  | ~\m3_addr_i[26] );
  assign \new_[12297]_  = (~\new_[17223]_  | ~\m2_addr_i[26] ) & (~\new_[17277]_  | ~\m1_addr_i[26] );
  assign \new_[12298]_  = (~\new_[17270]_  | ~\m4_addr_i[25] ) & (~\new_[18936]_  | ~\m3_addr_i[25] );
  assign \new_[12299]_  = ~\new_[30016]_  | ~\new_[15892]_  | ~\new_[30280]_ ;
  assign \new_[12300]_  = (~\m5_data_i[30]  | ~\new_[18014]_ ) & (~\m6_data_i[30]  | ~\new_[17229]_ );
  assign \new_[12301]_  = (~\m4_data_i[30]  | ~\new_[18149]_ ) & (~\m3_data_i[30]  | ~\new_[18929]_ );
  assign \new_[12302]_  = ~\new_[30444]_  | ~\new_[15893]_  | ~\new_[30218]_ ;
  assign \new_[12303]_  = (~\new_[17223]_  | ~\m2_addr_i[25] ) & (~\new_[18192]_  | ~\m1_addr_i[25] );
  assign \new_[12304]_  = ~\new_[15821]_  & ~\new_[16837]_ ;
  assign \new_[12305]_  = (~\m7_data_i[30]  | ~\new_[17232]_ ) & (~\m0_data_i[30]  | ~\new_[20580]_ );
  assign \new_[12306]_  = (~\m5_data_i[29]  | ~\new_[18014]_ ) & (~\m6_data_i[29]  | ~\new_[17229]_ );
  assign \new_[12307]_  = (~\m4_data_i[29]  | ~\new_[18149]_ ) & (~\m3_data_i[29]  | ~\new_[18929]_ );
  assign \new_[12308]_  = (~\new_[17270]_  | ~\m4_addr_i[24] ) & (~\new_[32350]_  | ~\m3_addr_i[24] );
  assign \new_[12309]_  = (~\m7_data_i[29]  | ~\new_[17232]_ ) & (~\m0_data_i[29]  | ~\new_[20580]_ );
  assign \new_[12310]_  = (~\m5_data_i[28]  | ~\new_[18014]_ ) & (~\m6_data_i[28]  | ~\new_[17229]_ );
  assign \new_[12311]_  = ~\new_[29557]_  | ~\new_[14517]_  | ~\new_[30123]_ ;
  assign \new_[12312]_  = (~\new_[17223]_  | ~\m2_addr_i[24] ) & (~\new_[18192]_  | ~\m1_addr_i[24] );
  assign \new_[12313]_  = (~\m4_data_i[28]  | ~\new_[18149]_ ) & (~\m3_data_i[28]  | ~\new_[18929]_ );
  assign \new_[12314]_  = (~\m3_addr_i[23]  | ~\new_[32350]_ ) & (~\m2_addr_i[23]  | ~\new_[17223]_ );
  assign \new_[12315]_  = (~\m7_data_i[28]  | ~\new_[17232]_ ) & (~\m0_data_i[28]  | ~\new_[18941]_ );
  assign \new_[12316]_  = (~\m4_data_i[27]  | ~\new_[18149]_ ) & (~\m3_data_i[27]  | ~\new_[18928]_ );
  assign \new_[12317]_  = ~\new_[15822]_  & ~\new_[16980]_ ;
  assign \new_[12318]_  = ~\new_[29900]_  | ~\new_[14521]_  | ~\new_[30104]_ ;
  assign \new_[12319]_  = (~\m5_data_i[26]  | ~\new_[18014]_ ) & (~\m6_data_i[26]  | ~\new_[17229]_ );
  assign \new_[12320]_  = (~\m4_data_i[26]  | ~\new_[18149]_ ) & (~\m3_data_i[26]  | ~\new_[18928]_ );
  assign \new_[12321]_  = (~\m7_data_i[26]  | ~\new_[17232]_ ) & (~\m0_data_i[26]  | ~\new_[19648]_ );
  assign \new_[12322]_  = ~\new_[13853]_ ;
  assign \new_[12323]_  = (~\m5_data_i[25]  | ~\new_[18015]_ ) & (~\m6_data_i[25]  | ~\new_[17229]_ );
  assign \new_[12324]_  = ~\new_[21121]_  & (~\new_[16015]_  | ~\new_[28845]_ );
  assign \new_[12325]_  = (~\m4_data_i[25]  | ~\new_[18149]_ ) & (~\m3_data_i[25]  | ~\new_[18928]_ );
  assign \new_[12326]_  = (~\m5_addr_i[22]  | ~\new_[17202]_ ) & (~\m4_addr_i[22]  | ~\new_[17270]_ );
  assign \new_[12327]_  = (~\m7_data_i[24]  | ~\new_[17232]_ ) & (~\m0_data_i[24]  | ~\new_[20580]_ );
  assign \new_[12328]_  = (~\m4_data_i[24]  | ~\new_[18149]_ ) & (~\m3_data_i[24]  | ~\new_[18928]_ );
  assign \new_[12329]_  = (~\m5_data_i[24]  | ~\new_[18016]_ ) & (~\m6_data_i[24]  | ~\new_[17229]_ );
  assign \new_[12330]_  = (~\m5_data_i[23]  | ~\new_[18014]_ ) & (~\m6_data_i[23]  | ~\new_[17229]_ );
  assign \new_[12331]_  = (~\m7_addr_i[22]  | ~\new_[17240]_ ) & (~\m6_addr_i[22]  | ~\new_[17227]_ );
  assign \new_[12332]_  = (~\m4_data_i[23]  | ~\new_[18149]_ ) & (~\m3_data_i[23]  | ~\new_[18929]_ );
  assign \new_[12333]_  = (~\m5_data_i[22]  | ~\new_[18014]_ ) & (~\m6_data_i[22]  | ~\new_[17229]_ );
  assign \new_[12334]_  = ~\new_[13861]_ ;
  assign \new_[12335]_  = (~\m4_data_i[22]  | ~\new_[18149]_ ) & (~\m3_data_i[22]  | ~\new_[18929]_ );
  assign \new_[12336]_  = ~\new_[13862]_ ;
  assign \new_[12337]_  = (~\m5_addr_i[21]  | ~\new_[17203]_ ) & (~\m4_addr_i[21]  | ~\new_[17270]_ );
  assign \new_[12338]_  = (~\m4_data_i[21]  | ~\new_[18149]_ ) & (~\m3_data_i[21]  | ~\new_[18928]_ );
  assign \new_[12339]_  = (~\m3_addr_i[21]  | ~\new_[18936]_ ) & (~\m2_addr_i[21]  | ~\new_[18808]_ );
  assign \new_[12340]_  = (~\m5_data_i[20]  | ~\new_[18014]_ ) & (~\m6_data_i[20]  | ~\new_[17229]_ );
  assign \new_[12341]_  = (~\m4_data_i[20]  | ~\new_[18149]_ ) & (~\m3_data_i[20]  | ~\new_[18928]_ );
  assign \new_[12342]_  = ~\new_[13866]_ ;
  assign \new_[12343]_  = (~\m4_data_i[19]  | ~\new_[18149]_ ) & (~\m3_data_i[19]  | ~\new_[18929]_ );
  assign \new_[12344]_  = (~\m3_addr_i[20]  | ~\new_[32350]_ ) & (~\m2_addr_i[20]  | ~\new_[17223]_ );
  assign \new_[12345]_  = (~\m5_data_i[18]  | ~\new_[18014]_ ) & (~\m6_data_i[18]  | ~\new_[17229]_ );
  assign \new_[12346]_  = (~\m7_data_i[18]  | ~\new_[17232]_ ) & (~\m0_data_i[18]  | ~\new_[19648]_ );
  assign \new_[12347]_  = ~\new_[15730]_  & ~\new_[23693]_ ;
  assign \new_[12348]_  = (~\m7_addr_i[20]  | ~\new_[17240]_ ) & (~\m6_addr_i[20]  | ~\new_[18090]_ );
  assign \new_[12349]_  = ~\new_[13875]_ ;
  assign \new_[12350]_  = (~\m5_addr_i[20]  | ~\new_[17203]_ ) & (~\m4_addr_i[20]  | ~\new_[17270]_ );
  assign \new_[12351]_  = (~\m7_data_i[30]  | ~\new_[19584]_ ) & (~\m0_data_i[30]  | ~\new_[18026]_ );
  assign \new_[12352]_  = ~\new_[21164]_  & (~\new_[16044]_  | ~\new_[28880]_ );
  assign \new_[12353]_  = (~\m5_data_i[16]  | ~\new_[18014]_ ) & (~\m6_data_i[16]  | ~\new_[17229]_ );
  assign \new_[12354]_  = (~\m4_data_i[16]  | ~\new_[18149]_ ) & (~\m3_data_i[16]  | ~\new_[18928]_ );
  assign \new_[12355]_  = ~\new_[13884]_ ;
  assign \new_[12356]_  = ~\new_[13885]_ ;
  assign \new_[12357]_  = (~\m5_addr_i[19]  | ~\new_[17202]_ ) & (~\m4_addr_i[19]  | ~\new_[16309]_ );
  assign \new_[12358]_  = (~\m5_data_i[12]  | ~\new_[18016]_ ) & (~\m6_data_i[12]  | ~\new_[17229]_ );
  assign \new_[12359]_  = (~\m4_data_i[12]  | ~\new_[18149]_ ) & (~\m3_data_i[12]  | ~\new_[18928]_ );
  assign \new_[12360]_  = (~\m5_addr_i[18]  | ~\new_[17203]_ ) & (~\m4_addr_i[18]  | ~\new_[16309]_ );
  assign \new_[12361]_  = ~\new_[15742]_  & ~\new_[26955]_ ;
  assign \new_[12362]_  = ~\new_[13895]_ ;
  assign \new_[12363]_  = (~\m4_data_i[10]  | ~\new_[18149]_ ) & (~\m3_data_i[10]  | ~\new_[18928]_ );
  assign \new_[12364]_  = ~\new_[13897]_ ;
  assign \new_[12365]_  = (~\m7_data_i[10]  | ~\new_[17232]_ ) & (~\m0_data_i[10]  | ~\new_[18941]_ );
  assign \new_[12366]_  = (~\m3_addr_i[17]  | ~\new_[32350]_ ) & (~\m2_addr_i[17]  | ~\new_[17223]_ );
  assign \new_[12367]_  = (~\m5_data_i[8]  | ~\new_[18016]_ ) & (~\m6_data_i[8]  | ~\new_[17229]_ );
  assign \new_[12368]_  = (~\m5_addr_i[17]  | ~\new_[17202]_ ) & (~\m4_addr_i[17]  | ~\new_[17270]_ );
  assign \new_[12369]_  = (~\m7_data_i[8]  | ~\new_[17232]_ ) & (~\m0_data_i[8]  | ~\new_[18941]_ );
  assign \new_[12370]_  = (~\m5_data_i[7]  | ~\new_[18016]_ ) & (~\m6_data_i[7]  | ~\new_[17229]_ );
  assign \new_[12371]_  = (~\m7_data_i[6]  | ~\new_[17232]_ ) & (~\m0_data_i[6]  | ~\new_[20580]_ );
  assign \new_[12372]_  = ~\new_[13911]_ ;
  assign \new_[12373]_  = (~\m4_data_i[5]  | ~\new_[18149]_ ) & (~\m3_data_i[5]  | ~\new_[18929]_ );
  assign \new_[12374]_  = ~\new_[21183]_  & (~\new_[16080]_  | ~\new_[30279]_ );
  assign \new_[12375]_  = (~\m3_addr_i[16]  | ~\new_[32350]_ ) & (~\m2_addr_i[16]  | ~\new_[17223]_ );
  assign \new_[12376]_  = (~\m7_data_i[5]  | ~\new_[17232]_ ) & (~\m0_data_i[5]  | ~\new_[18941]_ );
  assign \new_[12377]_  = (~\m5_addr_i[16]  | ~\new_[17202]_ ) & (~\m4_addr_i[16]  | ~\new_[16309]_ );
  assign \new_[12378]_  = (~\m4_data_i[4]  | ~\new_[18149]_ ) & (~\m3_data_i[4]  | ~\new_[18928]_ );
  assign \new_[12379]_  = (~\m5_addr_i[15]  | ~\new_[17202]_ ) & (~\m4_addr_i[15]  | ~\new_[17270]_ );
  assign \new_[12380]_  = (~\m4_data_i[3]  | ~\new_[18149]_ ) & (~\m3_data_i[3]  | ~\new_[18929]_ );
  assign \new_[12381]_  = ~\new_[13919]_ ;
  assign \new_[12382]_  = (~\m4_data_i[2]  | ~\new_[18149]_ ) & (~\m3_data_i[2]  | ~\new_[18929]_ );
  assign \new_[12383]_  = ~\new_[13923]_ ;
  assign \new_[12384]_  = (~\m7_data_i[2]  | ~\new_[17232]_ ) & (~\m0_data_i[2]  | ~\new_[18941]_ );
  assign \new_[12385]_  = ~\new_[13927]_ ;
  assign \new_[12386]_  = (~\m7_data_i[3]  | ~\new_[17240]_ ) & (~\m6_data_i[3]  | ~\new_[19581]_ );
  assign \new_[12387]_  = \new_[14570]_  | \new_[24550]_ ;
  assign \new_[12388]_  = (~\m5_addr_i[14]  | ~\new_[18745]_ ) & (~\m4_addr_i[14]  | ~\new_[18884]_ );
  assign \new_[12389]_  = (~\new_[17232]_  | ~\m7_addr_i[31] ) & (~\new_[19648]_  | ~\m0_addr_i[31] );
  assign \new_[12390]_  = (~\m3_addr_i[13]  | ~\new_[32350]_ ) & (~\m2_addr_i[13]  | ~\new_[17223]_ );
  assign \new_[12391]_  = ~\new_[15770]_  & ~\new_[23729]_ ;
  assign \new_[12392]_  = (~\new_[17232]_  | ~\new_[31531]_ ) & (~\new_[20580]_  | ~\new_[31481]_ );
  assign \new_[12393]_  = (~\new_[18149]_  | ~\m4_addr_i[29] ) & (~\new_[18930]_  | ~\m3_addr_i[29] );
  assign \new_[12394]_  = (~\new_[17232]_  | ~\new_[30577]_ ) & (~\new_[20580]_  | ~\new_[30957]_ );
  assign \new_[12395]_  = ~\new_[22307]_  & (~\new_[16042]_  | ~\new_[29225]_ );
  assign \new_[12396]_  = \new_[14572]_  | \new_[23997]_ ;
  assign \new_[12397]_  = ~\new_[13935]_ ;
  assign \new_[12398]_  = (~\m7_addr_i[13]  | ~\new_[17240]_ ) & (~\m6_addr_i[13]  | ~\new_[19581]_ );
  assign \new_[12399]_  = (~\new_[17232]_  | ~\m7_addr_i[27] ) & (~\new_[20580]_  | ~\m0_addr_i[27] );
  assign \new_[12400]_  = (~\m5_addr_i[13]  | ~\new_[17202]_ ) & (~\m4_addr_i[13]  | ~\new_[16309]_ );
  assign \new_[12401]_  = (~\new_[17232]_  | ~\m7_addr_i[26] ) & (~\new_[20580]_  | ~\m0_addr_i[26] );
  assign \new_[12402]_  = ~\new_[23786]_  & (~\new_[16091]_  | ~\new_[30158]_ );
  assign \new_[12403]_  = (~\m3_addr_i[12]  | ~\new_[32350]_ ) & (~\m2_addr_i[12]  | ~\new_[17223]_ );
  assign \new_[12404]_  = (~\m7_data_i[24]  | ~\new_[18106]_ ) & (~\m0_data_i[24]  | ~\new_[18026]_ );
  assign \new_[12405]_  = ~\new_[13947]_ ;
  assign \new_[12406]_  = (~\new_[17232]_  | ~\m7_addr_i[25] ) & (~\new_[19648]_  | ~\m0_addr_i[25] );
  assign \new_[12407]_  = (~\m7_addr_i[12]  | ~\new_[17240]_ ) & (~\m6_addr_i[12]  | ~\new_[17227]_ );
  assign \new_[12408]_  = (~\new_[18149]_  | ~\m4_addr_i[24] ) & (~\new_[18928]_  | ~\m3_addr_i[24] );
  assign \new_[12409]_  = (~\m5_addr_i[12]  | ~\new_[17202]_ ) & (~\m4_addr_i[12]  | ~\new_[17270]_ );
  assign \new_[12410]_  = (~\new_[17232]_  | ~\m7_addr_i[24] ) & (~\new_[18941]_  | ~\m0_addr_i[24] );
  assign \new_[12411]_  = (~\m5_addr_i[23]  | ~\new_[18016]_ ) & (~\m6_addr_i[23]  | ~\new_[17229]_ );
  assign \new_[12412]_  = (~\m7_data_i[7]  | ~\new_[19584]_ ) & (~\m0_data_i[7]  | ~\new_[18026]_ );
  assign \new_[12413]_  = (~\m7_addr_i[21]  | ~\new_[17232]_ ) & (~\m0_addr_i[21]  | ~\new_[20580]_ );
  assign \new_[12414]_  = ~\new_[15787]_  & ~\new_[22379]_ ;
  assign \new_[12415]_  = (~\m5_addr_i[21]  | ~\new_[18016]_ ) & (~\m6_addr_i[21]  | ~\new_[17229]_ );
  assign \new_[12416]_  = (~\m2_data_i[26]  | ~\new_[18077]_ ) & (~\m1_data_i[26]  | ~\new_[19632]_ );
  assign \new_[12417]_  = (~\m5_addr_i[20]  | ~\new_[18015]_ ) & (~\m6_addr_i[20]  | ~\new_[17229]_ );
  assign \new_[12418]_  = ~\new_[13959]_ ;
  assign \new_[12419]_  = (~\m7_addr_i[11]  | ~\new_[17240]_ ) & (~\m6_addr_i[11]  | ~\new_[18089]_ );
  assign \new_[12420]_  = (~\m7_addr_i[20]  | ~\new_[17232]_ ) & (~\m0_addr_i[20]  | ~\new_[19648]_ );
  assign \new_[12421]_  = \new_[14575]_  | \new_[26416]_ ;
  assign \new_[12422]_  = ~\new_[13961]_ ;
  assign \new_[12423]_  = (~\m7_addr_i[10]  | ~\new_[17240]_ ) & (~\m6_addr_i[10]  | ~\new_[18819]_ );
  assign \new_[12424]_  = ~\new_[22854]_  & (~\new_[16075]_  | ~\new_[26535]_ );
  assign \new_[12425]_  = ~\new_[22227]_  & (~\new_[16027]_  | ~\new_[29386]_ );
  assign \new_[12426]_  = (~\m4_addr_i[19]  | ~\new_[18149]_ ) & (~\m3_addr_i[19]  | ~\new_[18928]_ );
  assign \new_[12427]_  = (~\m5_addr_i[19]  | ~\new_[18015]_ ) & (~\m6_addr_i[19]  | ~\new_[17229]_ );
  assign \new_[12428]_  = (~\m4_addr_i[18]  | ~\new_[18149]_ ) & (~\m3_addr_i[18]  | ~\new_[18928]_ );
  assign \new_[12429]_  = (~\m5_addr_i[18]  | ~\new_[18016]_ ) & (~\m6_addr_i[18]  | ~\new_[17229]_ );
  assign \new_[12430]_  = ~\new_[22456]_  & (~\new_[16082]_  | ~\new_[29563]_ );
  assign \new_[12431]_  = (~\m7_data_i[14]  | ~\new_[18108]_ ) & (~\m0_data_i[14]  | ~\new_[18026]_ );
  assign \new_[12432]_  = (~\m7_addr_i[9]  | ~\new_[17240]_ ) & (~\m6_addr_i[9]  | ~\new_[18819]_ );
  assign \new_[12433]_  = (~\m5_addr_i[17]  | ~\new_[18016]_ ) & (~\m6_addr_i[17]  | ~\new_[17229]_ );
  assign \new_[12434]_  = (~\m4_addr_i[16]  | ~\new_[18149]_ ) & (~\m3_addr_i[16]  | ~\new_[18929]_ );
  assign \new_[12435]_  = (~\m7_addr_i[15]  | ~\new_[17232]_ ) & (~\m0_addr_i[15]  | ~\new_[20580]_ );
  assign \new_[12436]_  = (~\m5_data_i[11]  | ~\new_[18015]_ ) & (~\m6_data_i[11]  | ~\new_[17229]_ );
  assign \new_[12437]_  = (~\m5_addr_i[15]  | ~\new_[18016]_ ) & (~\m6_addr_i[15]  | ~\new_[17229]_ );
  assign \new_[12438]_  = (~\m5_addr_i[14]  | ~\new_[18014]_ ) & (~\m6_addr_i[14]  | ~\new_[17229]_ );
  assign \new_[12439]_  = (~\m3_addr_i[8]  | ~\new_[32350]_ ) & (~\m2_addr_i[8]  | ~\new_[18808]_ );
  assign \new_[12440]_  = (~\m7_addr_i[14]  | ~\new_[17232]_ ) & (~\m0_addr_i[14]  | ~\new_[20580]_ );
  assign \new_[12441]_  = (~\m5_addr_i[13]  | ~\new_[18014]_ ) & (~\m6_addr_i[13]  | ~\new_[17229]_ );
  assign \new_[12442]_  = (~\m7_addr_i[13]  | ~\new_[17232]_ ) & (~\m0_addr_i[13]  | ~\new_[19648]_ );
  assign \new_[12443]_  = ~\new_[15823]_  | ~\new_[21544]_ ;
  assign \new_[12444]_  = (~\m4_addr_i[12]  | ~\new_[18149]_ ) & (~\m3_addr_i[12]  | ~\new_[18929]_ );
  assign \new_[12445]_  = (~\m7_addr_i[11]  | ~\new_[17232]_ ) & (~\m0_addr_i[11]  | ~\new_[20580]_ );
  assign \new_[12446]_  = (~\m5_addr_i[11]  | ~\new_[18016]_ ) & (~\m6_addr_i[11]  | ~\new_[17229]_ );
  assign \new_[12447]_  = (~\m5_addr_i[7]  | ~\new_[17202]_ ) & (~\m4_addr_i[7]  | ~\new_[17270]_ );
  assign \new_[12448]_  = ~\new_[26626]_  & (~\new_[16016]_  | ~\new_[22709]_ );
  assign \new_[12449]_  = (~\m7_addr_i[10]  | ~\new_[17232]_ ) & (~\m0_addr_i[10]  | ~\new_[20580]_ );
  assign \new_[12450]_  = (~\m4_addr_i[10]  | ~\new_[18149]_ ) & (~\m3_addr_i[10]  | ~\new_[18929]_ );
  assign \new_[12451]_  = (~\m7_addr_i[9]  | ~\new_[17232]_ ) & (~\m0_addr_i[9]  | ~\new_[20580]_ );
  assign \new_[12452]_  = (~\m5_addr_i[9]  | ~\new_[18016]_ ) & (~\m6_addr_i[9]  | ~\new_[17229]_ );
  assign \new_[12453]_  = ~\new_[15824]_  | ~\new_[22860]_ ;
  assign \new_[12454]_  = ~\new_[15825]_  | ~\new_[21535]_ ;
  assign \new_[12455]_  = (~\m4_addr_i[8]  | ~\new_[18149]_ ) & (~\m3_addr_i[8]  | ~\new_[18928]_ );
  assign \new_[12456]_  = (~\m5_addr_i[6]  | ~\new_[17202]_ ) & (~\m4_addr_i[6]  | ~\new_[17270]_ );
  assign \new_[12457]_  = (~\m7_addr_i[7]  | ~\new_[17232]_ ) & (~\m0_addr_i[7]  | ~\new_[20580]_ );
  assign \new_[12458]_  = ~\new_[26652]_  & (~\new_[16025]_  | ~\new_[21413]_ );
  assign \new_[12459]_  = (~\m7_data_i[5]  | ~\new_[19584]_ ) & (~\m0_data_i[5]  | ~\new_[18026]_ );
  assign \new_[12460]_  = (~\m5_addr_i[6]  | ~\new_[18014]_ ) & (~\m6_addr_i[6]  | ~\new_[17229]_ );
  assign \new_[12461]_  = (~\m7_addr_i[6]  | ~\new_[17232]_ ) & (~\m0_addr_i[6]  | ~\new_[19648]_ );
  assign \new_[12462]_  = ~\new_[26774]_  & (~\new_[16028]_  | ~\new_[19406]_ );
  assign \new_[12463]_  = ~\new_[15827]_  | ~\new_[21504]_ ;
  assign \new_[12464]_  = ~\new_[15828]_  | ~\new_[21540]_ ;
  assign \new_[12465]_  = ~\new_[15830]_  | ~\new_[22969]_ ;
  assign \new_[12466]_  = (~\m7_addr_i[5]  | ~\new_[17232]_ ) & (~\m0_addr_i[5]  | ~\new_[18941]_ );
  assign \new_[12467]_  = (~\m4_addr_i[4]  | ~\new_[18149]_ ) & (~\m3_addr_i[4]  | ~\new_[18929]_ );
  assign \new_[12468]_  = (~\m7_addr_i[4]  | ~\new_[17232]_ ) & (~\m0_addr_i[4]  | ~\new_[18941]_ );
  assign \new_[12469]_  = (~\m3_addr_i[5]  | ~\new_[18936]_ ) & (~\new_[31095]_  | ~\new_[17224]_ );
  assign \new_[12470]_  = ~\new_[28304]_  & (~\new_[16036]_  | ~\new_[21350]_ );
  assign \new_[12471]_  = (~\m7_data_i[14]  | ~\new_[19606]_ ) & (~\m0_data_i[14]  | ~\new_[18781]_ );
  assign \new_[12472]_  = (~\m4_addr_i[3]  | ~\new_[18149]_ ) & (~\m3_addr_i[3]  | ~\new_[18928]_ );
  assign \new_[12473]_  = (~\m2_addr_i[15]  | ~\new_[18078]_ ) & (~\m1_addr_i[15]  | ~\new_[18184]_ );
  assign \new_[12474]_  = ~\new_[15831]_  | ~\new_[22886]_ ;
  assign \new_[12475]_  = ~\new_[15832]_  | ~\new_[21475]_ ;
  assign \new_[12476]_  = ~\new_[15833]_  | ~\new_[21782]_ ;
  assign \new_[12477]_  = (~\m4_addr_i[1]  | ~\new_[18149]_ ) & (~\m3_addr_i[1]  | ~\new_[18928]_ );
  assign \new_[12478]_  = (~\m5_addr_i[1]  | ~\new_[18015]_ ) & (~\m6_addr_i[1]  | ~\new_[17229]_ );
  assign \new_[12479]_  = (~\m7_addr_i[4]  | ~\new_[17240]_ ) & (~\m6_addr_i[4]  | ~\new_[18090]_ );
  assign \new_[12480]_  = (~\m4_addr_i[0]  | ~\new_[18149]_ ) & (~\m3_addr_i[0]  | ~\new_[18929]_ );
  assign \new_[12481]_  = (~\m3_addr_i[4]  | ~\new_[18936]_ ) & (~\m2_addr_i[4]  | ~\new_[17224]_ );
  assign \new_[12482]_  = ~\new_[27395]_  & (~\new_[16045]_  | ~\new_[22676]_ );
  assign \new_[12483]_  = (~\m5_sel_i[3]  | ~\new_[18016]_ ) & (~\m6_sel_i[3]  | ~\new_[17229]_ );
  assign \new_[12484]_  = (~\m5_sel_i[2]  | ~\new_[18014]_ ) & (~\m6_sel_i[2]  | ~\new_[17229]_ );
  assign \new_[12485]_  = (~\m7_addr_i[3]  | ~\new_[17240]_ ) & (~\m6_addr_i[3]  | ~\new_[18090]_ );
  assign \new_[12486]_  = ~\new_[15834]_  | ~\new_[20454]_ ;
  assign \new_[12487]_  = (~\m3_addr_i[3]  | ~\new_[18936]_ ) & (~\m2_addr_i[3]  | ~\new_[17224]_ );
  assign \new_[12488]_  = (~\m4_sel_i[1]  | ~\new_[18149]_ ) & (~\m3_sel_i[1]  | ~\new_[18928]_ );
  assign \new_[12489]_  = (~\m4_sel_i[0]  | ~\new_[18149]_ ) & (~\m3_sel_i[0]  | ~\new_[18928]_ );
  assign \new_[12490]_  = (~\m2_addr_i[8]  | ~\new_[18069]_ ) & (~\m1_addr_i[8]  | ~\new_[18897]_ );
  assign \new_[12491]_  = (~\m5_sel_i[0]  | ~\new_[18015]_ ) & (~\m6_sel_i[0]  | ~\new_[17229]_ );
  assign \new_[12492]_  = ~\new_[28691]_  & (~\new_[16052]_  | ~\new_[19408]_ );
  assign \new_[12493]_  = (~\m7_data_i[13]  | ~\new_[19584]_ ) & (~\m0_data_i[13]  | ~\new_[18026]_ );
  assign \new_[12494]_  = (~\m2_data_i[28]  | ~\new_[18069]_ ) & (~\m1_data_i[28]  | ~\new_[18897]_ );
  assign \new_[12495]_  = (~\m7_addr_i[2]  | ~\new_[17240]_ ) & (~\m6_addr_i[2]  | ~\new_[19581]_ );
  assign \new_[12496]_  = (~m7_we_i | ~\new_[17232]_ ) & (~m0_we_i | ~\new_[18941]_ );
  assign \new_[12497]_  = (~m5_we_i | ~\new_[18015]_ ) & (~m6_we_i | ~\new_[17229]_ );
  assign \new_[12498]_  = ~\new_[15837]_  | ~\new_[22863]_ ;
  assign \new_[12499]_  = ~\new_[15811]_  & (~\new_[29959]_  | ~\new_[31422]_ );
  assign \new_[12500]_  = (~\m5_addr_i[1]  | ~\new_[17202]_ ) & (~\m4_addr_i[1]  | ~\new_[17270]_ );
  assign \new_[12501]_  = (~\m2_data_i[30]  | ~\new_[18067]_ ) & (~\m1_data_i[30]  | ~\new_[20573]_ );
  assign \new_[12502]_  = (~\m2_data_i[29]  | ~\new_[18069]_ ) & (~\m1_data_i[29]  | ~\new_[18901]_ );
  assign \new_[12503]_  = ~\new_[15838]_  | ~\new_[20504]_ ;
  assign \new_[12504]_  = ~\new_[26754]_  & (~\new_[16076]_  | ~\new_[22804]_ );
  assign \new_[12505]_  = (~\m2_data_i[27]  | ~\new_[18068]_ ) & (~\m1_data_i[27]  | ~\new_[20573]_ );
  assign \new_[12506]_  = (~\m2_data_i[26]  | ~\new_[18068]_ ) & (~\m1_data_i[26]  | ~\new_[19625]_ );
  assign \new_[12507]_  = ~\new_[15840]_  | ~\new_[20461]_ ;
  assign \new_[12508]_  = ~\new_[28848]_  & (~\new_[16050]_  | ~\new_[22776]_ );
  assign \new_[12509]_  = (~\m2_data_i[23]  | ~\new_[18069]_ ) & (~\m1_data_i[23]  | ~\new_[20573]_ );
  assign \new_[12510]_  = ~\new_[15841]_  | ~\new_[20457]_ ;
  assign \new_[12511]_  = ~\new_[15842]_  | ~\new_[23055]_ ;
  assign \new_[12512]_  = (~\m7_sel_i[3]  | ~\new_[18116]_ ) & (~\m0_sel_i[3]  | ~\new_[18932]_ );
  assign \new_[12513]_  = (~\m3_sel_i[1]  | ~\new_[32350]_ ) & (~\m2_sel_i[1]  | ~\new_[17223]_ );
  assign \new_[12514]_  = (~\m2_data_i[20]  | ~\new_[18067]_ ) & (~\m1_data_i[20]  | ~\new_[20573]_ );
  assign \new_[12515]_  = ~\new_[26644]_  & (~\new_[16089]_  | ~\new_[22773]_ );
  assign \new_[12516]_  = ~\new_[15843]_  | ~\new_[20507]_ ;
  assign \new_[12517]_  = ~\new_[15844]_  | ~\new_[20525]_ ;
  assign \new_[12518]_  = (~\m2_data_i[16]  | ~\new_[18067]_ ) & (~\m1_data_i[16]  | ~\new_[20573]_ );
  assign \new_[12519]_  = (~\m2_data_i[14]  | ~\new_[18069]_ ) & (~\m1_data_i[14]  | ~\new_[18899]_ );
  assign \new_[12520]_  = ~\new_[15845]_  | ~\new_[21546]_ ;
  assign \new_[12521]_  = ~\new_[15846]_  | ~\new_[21533]_ ;
  assign \new_[12522]_  = ~\new_[15847]_  | ~\new_[22911]_ ;
  assign \new_[12523]_  = ~\new_[15848]_  | ~\new_[24298]_ ;
  assign \new_[12524]_  = ~\new_[15815]_  & (~\new_[30188]_  | ~\new_[5989]_ );
  assign \new_[12525]_  = (~\m7_data_i[13]  | ~\new_[18095]_ ) & (~\m0_data_i[13]  | ~\new_[18767]_ );
  assign \new_[12526]_  = (~\m2_data_i[11]  | ~\new_[18068]_ ) & (~\m1_data_i[11]  | ~\new_[18901]_ );
  assign \new_[12527]_  = (~\m7_data_i[11]  | ~\new_[18095]_ ) & (~\m0_data_i[11]  | ~\new_[20545]_ );
  assign \new_[12528]_  = ~\new_[15849]_  | ~\new_[21472]_ ;
  assign \new_[12529]_  = ~\new_[15850]_  | ~\new_[21502]_ ;
  assign \new_[12530]_  = (~\m2_data_i[9]  | ~\new_[18068]_ ) & (~\m1_data_i[9]  | ~\new_[20573]_ );
  assign \new_[12531]_  = (~\m7_data_i[9]  | ~\new_[18095]_ ) & (~\m0_data_i[9]  | ~\new_[20545]_ );
  assign \new_[12532]_  = (~\m7_data_i[8]  | ~\new_[18095]_ ) & (~\m0_data_i[8]  | ~\new_[18767]_ );
  assign \new_[12533]_  = ~\new_[28053]_  & (~\new_[16014]_  | ~\new_[22786]_ );
  assign \new_[12534]_  = (~\m7_data_i[7]  | ~\new_[18095]_ ) & (~\m0_data_i[7]  | ~\new_[20545]_ );
  assign \new_[12535]_  = (~\m2_data_i[6]  | ~\new_[18067]_ ) & (~\m1_data_i[6]  | ~\new_[20573]_ );
  assign \new_[12536]_  = ~\new_[29054]_  & (~\new_[16105]_  | ~\new_[19418]_ );
  assign \new_[12537]_  = (~\m7_data_i[5]  | ~\new_[18095]_ ) & (~\m0_data_i[5]  | ~\new_[18767]_ );
  assign \new_[12538]_  = ~\new_[15851]_  | ~\new_[21527]_ ;
  assign \new_[12539]_  = ~\new_[27240]_  & (~\new_[16061]_  | ~\new_[22766]_ );
  assign \new_[12540]_  = ~\new_[15852]_  | ~\new_[21541]_ ;
  assign \new_[12541]_  = ~\new_[15853]_  | ~\new_[21518]_ ;
  assign \new_[12542]_  = ~\new_[15839]_  | ~\new_[22950]_ ;
  assign \new_[12543]_  = (~\m7_data_i[0]  | ~\new_[18095]_ ) & (~\m0_data_i[0]  | ~\new_[20545]_ );
  assign \new_[12544]_  = (~\m2_data_i[31]  | ~\new_[18078]_ ) & (~\m1_data_i[31]  | ~\new_[19632]_ );
  assign \new_[12545]_  = ~\new_[15820]_  & (~\new_[30265]_  | ~\new_[5928]_ );
  assign \new_[12546]_  = ~\new_[15854]_  | ~\new_[20474]_ ;
  assign \new_[12547]_  = ~\new_[28426]_  & (~\new_[16128]_  | ~\new_[21453]_ );
  assign \new_[12548]_  = ~\new_[29156]_  & (~\new_[16108]_  | ~\new_[29808]_ );
  assign \new_[12549]_  = (~\new_[18067]_  | ~\m2_addr_i[25] ) & (~\new_[20573]_  | ~\m1_addr_i[25] );
  assign \new_[12550]_  = ~\new_[15855]_  | ~\new_[20453]_ ;
  assign \new_[12551]_  = (~\m2_addr_i[23]  | ~\new_[18067]_ ) & (~\m1_addr_i[23]  | ~\new_[20573]_ );
  assign \new_[12552]_  = ~\new_[27533]_  & (~\new_[16124]_  | ~\new_[29151]_ );
  assign \new_[12553]_  = ~\new_[26713]_  & (~\new_[16127]_  | ~\new_[22744]_ );
  assign \new_[12554]_  = ~\new_[29533]_  & (~\new_[16135]_  | ~\new_[19435]_ );
  assign \new_[12555]_  = ~\new_[23109]_  & (~\new_[16157]_  | ~\new_[20485]_ );
  assign \new_[12556]_  = ~\new_[28613]_  & (~\new_[16207]_  | ~\new_[18427]_ );
  assign \new_[12557]_  = (~\m5_data_i[24]  | ~\new_[18738]_ ) & (~\m6_data_i[24]  | ~\new_[18031]_ );
  assign \new_[12558]_  = ~\new_[28599]_  & (~\new_[16225]_  | ~\new_[18426]_ );
  assign \new_[12559]_  = ~\new_[15718]_  | ~\new_[22860]_ ;
  assign \new_[12560]_  = (~\m7_addr_i[5]  | ~\new_[18115]_ ) & (~\new_[31848]_  | ~\new_[18932]_ );
  assign \new_[12561]_  = ~\new_[15720]_  & ~\new_[26351]_ ;
  assign \new_[12562]_  = ~\new_[15722]_  | ~\new_[21504]_ ;
  assign \new_[12563]_  = ~\new_[15724]_  & ~\new_[29561]_ ;
  assign \new_[12564]_  = (~\m5_data_i[31]  | ~\new_[18016]_ ) & (~\m6_data_i[31]  | ~\new_[17229]_ );
  assign \new_[12565]_  = ~\new_[15727]_  | ~\new_[22886]_ ;
  assign \new_[12566]_  = (~\m5_data_i[22]  | ~\new_[18738]_ ) & (~\m6_data_i[22]  | ~\new_[18031]_ );
  assign \new_[12567]_  = ~\new_[15731]_  & ~\new_[28576]_ ;
  assign \new_[12568]_  = ~\new_[15737]_  | ~\new_[20454]_ ;
  assign \new_[12569]_  = (~\m5_data_i[21]  | ~\new_[18014]_ ) & (~\m6_data_i[21]  | ~\new_[17229]_ );
  assign \new_[12570]_  = ~\new_[24770]_  & (~\new_[16235]_  | ~\new_[29904]_ );
  assign \new_[12571]_  = ~\new_[26313]_  & (~\new_[16237]_  | ~\new_[29404]_ );
  assign \new_[12572]_  = (~\new_[19606]_  | ~\new_[30577]_ ) & (~\new_[18781]_  | ~\new_[30957]_ );
  assign \new_[12573]_  = ~\new_[15759]_  | ~\new_[20457]_ ;
  assign \new_[12574]_  = (~\m2_addr_i[9]  | ~\new_[18067]_ ) & (~\m1_addr_i[9]  | ~\new_[20573]_ );
  assign \new_[12575]_  = (~\m2_addr_i[16]  | ~\new_[18077]_ ) & (~\m1_addr_i[16]  | ~\new_[18182]_ );
  assign \new_[12576]_  = ~\new_[15760]_  & ~\new_[28221]_ ;
  assign \new_[12577]_  = ~\new_[15764]_  | ~\new_[20507]_ ;
  assign \new_[12578]_  = (~\m5_data_i[19]  | ~\new_[18016]_ ) & (~\m6_data_i[19]  | ~\new_[17229]_ );
  assign \new_[12579]_  = ~\new_[15768]_  | ~\new_[21546]_ ;
  assign \new_[12580]_  = (~\m2_addr_i[7]  | ~\new_[18068]_ ) & (~\m1_addr_i[7]  | ~\new_[19625]_ );
  assign \new_[12581]_  = ~\new_[15771]_  & ~\new_[27663]_ ;
  assign \new_[12582]_  = (~\m2_addr_i[6]  | ~\new_[18069]_ ) & (~\m1_addr_i[6]  | ~\new_[18897]_ );
  assign \new_[12583]_  = ~\new_[15775]_  | ~\new_[21472]_ ;
  assign \new_[12584]_  = ~\new_[22884]_  | (~\new_[16095]_  & ~\new_[29989]_ );
  assign \new_[12585]_  = ~\new_[15776]_  & ~\new_[28784]_ ;
  assign \new_[12586]_  = (~\new_[31095]_  | ~\new_[18069]_ ) & (~\m1_addr_i[5]  | ~\new_[19626]_ );
  assign \new_[12587]_  = ~\new_[15784]_  | ~\new_[21541]_ ;
  assign \new_[12588]_  = (~\new_[31399]_  | ~\new_[18069]_ ) & (~\m1_addr_i[3]  | ~\new_[18900]_ );
  assign \new_[12589]_  = ~\new_[15788]_  & ~\new_[27634]_ ;
  assign \new_[12590]_  = ~\new_[24542]_  & (~\new_[16240]_  | ~\new_[30016]_ );
  assign \new_[12591]_  = (~\m2_addr_i[2]  | ~\new_[18069]_ ) & (~\new_[31477]_  | ~\new_[18899]_ );
  assign \new_[12592]_  = ~\new_[24692]_  & (~\new_[16241]_  | ~\new_[29557]_ );
  assign \new_[12593]_  = (~\m2_sel_i[3]  | ~\new_[18069]_ ) & (~\m1_sel_i[3]  | ~\new_[18897]_ );
  assign \new_[12594]_  = ~\new_[29027]_  & (~\new_[16021]_  | ~\new_[30030]_ );
  assign \new_[12595]_  = (~\m5_data_i[14]  | ~\new_[18738]_ ) & (~\m6_data_i[14]  | ~\new_[18031]_ );
  assign \new_[12596]_  = ~\new_[28994]_  & (~\new_[16030]_  | ~\new_[28872]_ );
  assign \new_[12597]_  = ~\new_[29137]_  & (~\new_[16039]_  | ~\new_[30057]_ );
  assign \new_[12598]_  = ~\new_[30447]_  & (~\new_[16047]_  | ~\new_[28883]_ );
  assign \new_[12599]_  = (~\m2_sel_i[1]  | ~\new_[18069]_ ) & (~\m1_sel_i[1]  | ~\new_[18900]_ );
  assign \new_[12600]_  = (~\m5_data_i[13]  | ~\new_[18738]_ ) & (~\m6_data_i[13]  | ~\new_[18030]_ );
  assign \new_[12601]_  = (~\m2_sel_i[0]  | ~\new_[18069]_ ) & (~\m1_sel_i[0]  | ~\new_[18900]_ );
  assign \new_[12602]_  = ~\new_[30742]_  & (~\new_[16092]_  | ~\new_[28939]_ );
  assign \new_[12603]_  = ~\new_[29049]_  & (~\new_[16090]_  | ~\new_[28887]_ );
  assign \new_[12604]_  = ~\new_[29325]_  & (~\new_[16100]_  | ~\new_[29248]_ );
  assign \new_[12605]_  = (~\m5_data_i[12]  | ~\new_[18738]_ ) & (~\m6_data_i[12]  | ~\new_[18031]_ );
  assign \new_[12606]_  = ~\new_[29282]_  & (~\new_[16094]_  | ~\new_[28924]_ );
  assign \new_[12607]_  = (~\m5_data_i[21]  | ~\new_[18738]_ ) & (~\m6_data_i[21]  | ~\new_[18031]_ );
  assign \new_[12608]_  = ~\new_[29486]_  & (~\new_[16102]_  | ~\new_[29268]_ );
  assign \new_[12609]_  = (~\m2_addr_i[1]  | ~\new_[18069]_ ) & (~\m1_addr_i[1]  | ~\new_[19626]_ );
  assign \new_[12610]_  = (~\m5_data_i[10]  | ~\new_[18738]_ ) & (~\m6_data_i[10]  | ~\new_[18031]_ );
  assign \new_[12611]_  = ~\new_[14524]_  & (~\new_[30230]_  | ~\new_[6033]_ );
  assign \new_[12612]_  = (~\new_[15999]_  | ~\new_[29527]_ ) & (~\new_[30285]_  | ~\new_[5909]_ );
  assign \new_[12613]_  = ~\new_[14525]_  & (~\new_[29909]_  | ~\new_[6040]_ );
  assign \new_[12614]_  = (~\m7_data_i[28]  | ~\new_[18112]_ ) & (~\m0_data_i[28]  | ~\new_[18019]_ );
  assign \new_[12615]_  = (~\m2_data_i[28]  | ~\new_[16291]_ ) & (~\m1_data_i[28]  | ~\new_[18905]_ );
  assign \new_[12616]_  = (~\new_[16000]_  | ~\new_[29320]_ ) & (~\new_[30334]_  | ~\new_[5911]_ );
  assign \new_[12617]_  = ~\new_[14526]_  & (~\new_[29815]_  | ~\new_[6032]_ );
  assign \new_[12618]_  = (~\m5_data_i[8]  | ~\new_[18738]_ ) & (~\m6_data_i[8]  | ~\new_[18031]_ );
  assign \new_[12619]_  = (~\new_[16001]_  | ~\new_[29228]_ ) & (~\new_[30192]_  | ~\new_[5912]_ );
  assign \new_[12620]_  = (~\m7_data_i[26]  | ~\new_[18112]_ ) & (~\m0_data_i[26]  | ~\new_[18019]_ );
  assign \new_[12621]_  = (~\m5_data_i[7]  | ~\new_[18738]_ ) & (~\m6_data_i[7]  | ~\new_[18031]_ );
  assign \new_[12622]_  = (~\new_[16003]_  | ~\new_[29103]_ ) & (~\new_[30249]_  | ~\new_[5914]_ );
  assign \new_[12623]_  = (~\m7_data_i[25]  | ~\new_[18112]_ ) & (~\m0_data_i[25]  | ~\new_[18019]_ );
  assign \new_[12624]_  = (~\m2_data_i[25]  | ~\new_[16291]_ ) & (~\m1_data_i[25]  | ~\new_[18905]_ );
  assign \new_[12625]_  = ~\new_[14528]_  & (~\new_[29700]_  | ~\new_[5978]_ );
  assign \new_[12626]_  = (~\m7_data_i[24]  | ~\new_[18113]_ ) & (~\m0_data_i[24]  | ~\new_[18019]_ );
  assign \new_[12627]_  = (~\new_[16004]_  | ~\new_[29441]_ ) & (~\new_[30219]_  | ~\new_[5978]_ );
  assign \new_[12628]_  = ~\new_[15251]_  & (~\new_[30199]_  | ~\new_[6196]_ );
  assign \new_[12629]_  = (~\m5_data_i[6]  | ~\new_[18738]_ ) & (~\m6_data_i[6]  | ~\new_[18030]_ );
  assign \new_[12630]_  = ~\new_[14530]_  & (~\new_[29157]_  | ~\new_[5983]_ );
  assign \new_[12631]_  = (~\new_[16005]_  | ~\new_[28828]_ ) & (~\new_[30087]_  | ~\new_[5983]_ );
  assign \new_[12632]_  = (~\m5_data_i[23]  | ~\new_[17194]_ ) & (~\m6_data_i[23]  | ~\new_[18792]_ );
  assign \new_[12633]_  = (~\m2_data_i[23]  | ~\new_[17219]_ ) & (~\m1_data_i[23]  | ~\new_[18905]_ );
  assign \new_[12634]_  = (~\new_[16006]_  | ~\new_[28963]_ ) & (~\new_[30319]_  | ~\new_[5917]_ );
  assign \new_[12635]_  = ~\new_[15028]_  & (~\new_[30010]_  | ~\new_[31157]_ );
  assign \new_[12636]_  = (~\m5_data_i[22]  | ~\new_[17194]_ ) & (~\m6_data_i[22]  | ~\new_[18042]_ );
  assign \new_[12637]_  = (~\m5_data_i[5]  | ~\new_[18738]_ ) & (~\m6_data_i[5]  | ~\new_[18031]_ );
  assign \new_[12638]_  = (~\new_[16002]_  | ~\new_[29721]_ ) & (~\new_[30069]_  | ~\new_[5918]_ );
  assign \new_[12639]_  = (~\m2_data_i[22]  | ~\new_[17219]_ ) & (~\m1_data_i[22]  | ~\new_[18905]_ );
  assign \new_[12640]_  = ~\new_[14993]_  & (~\new_[30066]_  | ~\new_[6069]_ );
  assign \new_[12641]_  = (~\m5_data_i[21]  | ~\new_[17194]_ ) & (~\m6_data_i[21]  | ~\new_[18792]_ );
  assign \new_[12642]_  = (~\new_[16007]_  | ~\new_[29006]_ ) & (~\new_[29934]_  | ~\new_[5921]_ );
  assign \new_[12643]_  = (~\m2_data_i[21]  | ~\new_[17219]_ ) & (~\m1_data_i[21]  | ~\new_[18905]_ );
  assign \new_[12644]_  = ~\new_[14531]_  & (~\new_[30188]_  | ~\new_[6072]_ );
  assign \new_[12645]_  = (~\m5_data_i[4]  | ~\new_[18738]_ ) & (~\m6_data_i[4]  | ~\new_[18030]_ );
  assign \new_[12646]_  = (~\new_[16009]_  | ~\new_[29695]_ ) & (~\new_[30008]_  | ~\new_[5923]_ );
  assign \new_[12647]_  = (~\m5_data_i[20]  | ~\new_[17194]_ ) & (~\m6_data_i[20]  | ~\new_[18792]_ );
  assign \new_[12648]_  = ~\new_[14532]_  & (~\new_[30075]_  | ~\new_[5924]_ );
  assign \new_[12649]_  = (~\m2_data_i[20]  | ~\new_[17219]_ ) & (~\m1_data_i[20]  | ~\new_[18905]_ );
  assign \new_[12650]_  = (~\m7_data_i[19]  | ~\new_[18112]_ ) & (~\m0_data_i[19]  | ~\new_[18019]_ );
  assign \new_[12651]_  = (~\new_[16008]_  | ~\new_[30009]_ ) & (~\new_[29652]_  | ~\new_[5926]_ );
  assign \new_[12652]_  = ~\new_[14916]_  & (~\new_[30115]_  | ~\new_[6078]_ );
  assign \new_[12653]_  = (~\new_[16011]_  | ~\new_[29456]_ ) & (~\new_[30272]_  | ~\new_[5927]_ );
  assign \new_[12654]_  = ~\new_[14536]_  & (~\new_[30265]_  | ~\new_[6084]_ );
  assign \new_[12655]_  = (~\m5_data_i[3]  | ~\new_[18738]_ ) & (~\m6_data_i[3]  | ~\new_[18030]_ );
  assign \new_[12656]_  = (~\m7_data_i[18]  | ~\new_[18112]_ ) & (~\m0_data_i[18]  | ~\new_[18019]_ );
  assign \new_[12657]_  = (~\m2_data_i[18]  | ~\new_[16291]_ ) & (~\m1_data_i[18]  | ~\new_[18905]_ );
  assign \new_[12658]_  = ~\new_[15808]_  & (~\new_[29047]_  | ~\new_[31648]_ );
  assign \new_[12659]_  = (~\new_[16010]_  | ~\new_[28898]_ ) & (~\new_[30339]_  | ~\new_[31648]_ );
  assign \new_[12660]_  = ~\new_[14539]_  & (~\new_[29354]_  | ~\new_[31763]_ );
  assign \new_[12661]_  = (~\m7_data_i[17]  | ~\new_[18112]_ ) & (~\m0_data_i[17]  | ~\new_[18019]_ );
  assign \new_[12662]_  = (~\new_[16012]_  | ~\new_[29226]_ ) & (~\new_[30305]_  | ~\new_[31763]_ );
  assign \new_[12663]_  = (~\m2_data_i[17]  | ~\new_[16291]_ ) & (~\m1_data_i[17]  | ~\new_[18905]_ );
  assign \new_[12664]_  = (~\m7_data_i[16]  | ~\new_[18112]_ ) & (~\m0_data_i[16]  | ~\new_[18019]_ );
  assign \new_[12665]_  = (~\new_[16013]_  | ~\new_[30150]_ ) & (~\new_[28933]_  | ~\new_[6094]_ );
  assign \new_[12666]_  = (~\m2_data_i[16]  | ~\new_[16291]_ ) & (~\m1_data_i[16]  | ~\new_[18905]_ );
  assign \new_[12667]_  = (~\m5_data_i[2]  | ~\new_[18738]_ ) & (~\m6_data_i[2]  | ~\new_[18031]_ );
  assign \new_[12668]_  = (~\m7_data_i[15]  | ~\new_[18112]_ ) & (~\m0_data_i[15]  | ~\new_[18020]_ );
  assign \new_[12669]_  = \new_[5909]_  ? \new_[28908]_  : \new_[16022]_ ;
  assign \new_[12670]_  = (~\m7_data_i[14]  | ~\new_[18112]_ ) & (~\m0_data_i[14]  | ~\new_[18020]_ );
  assign \new_[12671]_  = (~\m5_data_i[1]  | ~\new_[18738]_ ) & (~\m6_data_i[1]  | ~\new_[18030]_ );
  assign \new_[12672]_  = \new_[5911]_  ? \new_[29112]_  : \new_[16031]_ ;
  assign \new_[12673]_  = (~\new_[16032]_  | ~\new_[30318]_ ) & (~\new_[30575]_  | ~\new_[31148]_ );
  assign \new_[12674]_  = (~\m5_data_i[13]  | ~\new_[17194]_ ) & (~\m6_data_i[13]  | ~\new_[18792]_ );
  assign \new_[12675]_  = (~\m2_data_i[13]  | ~\new_[16291]_ ) & (~\m1_data_i[13]  | ~\new_[18905]_ );
  assign \new_[12676]_  = \new_[5912]_  ? \new_[28968]_  : \new_[16040]_ ;
  assign \new_[12677]_  = (~\new_[16041]_  | ~\new_[29780]_ ) & (~\new_[30769]_  | ~\new_[6096]_ );
  assign \new_[12678]_  = (~\m5_data_i[12]  | ~\new_[17194]_ ) & (~\m6_data_i[12]  | ~\new_[18042]_ );
  assign \new_[12679]_  = \new_[5914]_  ? \new_[28835]_  : \new_[16048]_ ;
  assign \new_[12680]_  = (~\m5_data_i[11]  | ~\new_[17194]_ ) & (~\m6_data_i[11]  | ~\new_[18792]_ );
  assign \new_[12681]_  = (~\m2_data_i[11]  | ~\new_[17219]_ ) & (~\m1_data_i[11]  | ~\new_[18905]_ );
  assign \new_[12682]_  = (~\new_[18030]_  | ~\m6_addr_i[31] ) & (~\new_[18738]_  | ~\new_[31001]_ );
  assign \new_[12683]_  = (~\m4_data_i[9]  | ~\new_[17265]_ ) & (~\m3_data_i[9]  | ~\new_[17248]_ );
  assign \new_[12684]_  = (~\new_[18030]_  | ~\m6_addr_i[30] ) & (~\new_[18738]_  | ~\new_[31147]_ );
  assign \new_[12685]_  = (~\m5_data_i[8]  | ~\new_[17194]_ ) & (~\m6_data_i[8]  | ~\new_[18792]_ );
  assign \new_[12686]_  = (~\new_[16086]_  | ~\new_[30178]_ ) & (~\new_[30696]_  | ~\new_[6066]_ );
  assign \new_[12687]_  = \new_[5917]_  ? \new_[28911]_  : \new_[16084]_ ;
  assign \new_[12688]_  = (~\m2_data_i[8]  | ~\new_[17219]_ ) & (~\m1_data_i[8]  | ~\new_[18905]_ );
  assign \new_[12689]_  = (~\m3_addr_i[1]  | ~\new_[32350]_ ) & (~\m2_addr_i[1]  | ~\new_[17223]_ );
  assign \new_[12690]_  = \new_[5918]_  ? \new_[29633]_  : \new_[16018]_ ;
  assign \new_[12691]_  = (~\m7_data_i[7]  | ~\new_[18113]_ ) & (~\m0_data_i[7]  | ~\new_[18020]_ );
  assign \new_[12692]_  = \new_[5921]_  ? \new_[28864]_  : \new_[16060]_ ;
  assign \new_[12693]_  = (~\new_[16043]_  | ~\new_[30180]_ ) & (~\new_[30661]_  | ~\new_[6072]_ );
  assign \new_[12694]_  = (~\m5_data_i[6]  | ~\new_[17194]_ ) & (~\m6_data_i[6]  | ~\new_[18042]_ );
  assign \new_[12695]_  = \new_[5923]_  ? \new_[28844]_  : \new_[16065]_ ;
  assign \new_[12696]_  = (~\new_[18030]_  | ~\m6_addr_i[29] ) & (~\new_[18738]_  | ~\new_[31407]_ );
  assign \new_[12697]_  = (~\new_[16023]_  | ~\new_[30343]_ ) & (~\new_[30837]_  | ~\new_[5924]_ );
  assign \new_[12698]_  = (~\m5_data_i[5]  | ~\new_[17194]_ ) & (~\m6_data_i[5]  | ~\new_[18792]_ );
  assign \new_[12699]_  = (~\new_[18030]_  | ~\m6_addr_i[28] ) & (~\new_[18738]_  | ~\new_[31276]_ );
  assign \new_[12700]_  = (~\new_[16125]_  | ~\new_[29979]_ ) & (~\new_[30637]_  | ~\new_[5924]_ );
  assign \new_[12701]_  = (~\m2_data_i[5]  | ~\new_[17219]_ ) & (~\m1_data_i[5]  | ~\new_[18905]_ );
  assign \new_[12702]_  = (~\new_[16099]_  | ~\new_[30105]_ ) & (~\new_[29606]_  | ~\new_[5926]_ );
  assign \new_[12703]_  = (~\m4_data_i[5]  | ~\new_[17265]_ ) & (~\m3_data_i[5]  | ~\new_[17248]_ );
  assign \new_[12704]_  = (~\m7_data_i[4]  | ~\new_[18113]_ ) & (~\m0_data_i[4]  | ~\new_[18020]_ );
  assign \new_[12705]_  = \new_[5927]_  ? \new_[29189]_  : \new_[16104]_ ;
  assign \new_[12706]_  = (~\m2_addr_i[18]  | ~\new_[18077]_ ) & (~\m1_addr_i[18]  | ~\new_[18183]_ );
  assign \new_[12707]_  = (~\m2_data_i[4]  | ~\new_[17219]_ ) & (~\m1_data_i[4]  | ~\new_[18905]_ );
  assign \new_[12708]_  = (~\m2_data_i[3]  | ~\new_[17219]_ ) & (~\m1_data_i[3]  | ~\new_[18905]_ );
  assign \new_[12709]_  = (~\m4_data_i[3]  | ~\new_[17265]_ ) & (~\m3_data_i[3]  | ~\new_[18128]_ );
  assign \new_[12710]_  = (~\new_[18030]_  | ~\m6_addr_i[27] ) & (~\new_[18738]_  | ~\m5_addr_i[27] );
  assign \new_[12711]_  = (~\m5_data_i[2]  | ~\new_[17194]_ ) & (~\m6_data_i[2]  | ~\new_[18042]_ );
  assign \new_[12712]_  = (~\m2_data_i[2]  | ~\new_[17219]_ ) & (~\m1_data_i[2]  | ~\new_[18905]_ );
  assign \new_[12713]_  = (~\m5_data_i[1]  | ~\new_[17194]_ ) & (~\m6_data_i[1]  | ~\new_[18042]_ );
  assign \new_[12714]_  = (~\new_[18030]_  | ~\m6_addr_i[26] ) & (~\new_[18738]_  | ~\m5_addr_i[26] );
  assign \new_[12715]_  = (~\m2_data_i[1]  | ~\new_[17219]_ ) & (~\m1_data_i[1]  | ~\new_[18905]_ );
  assign \new_[12716]_  = ~\new_[24674]_  & (~\new_[16257]_  | ~\new_[29550]_ );
  assign \new_[12717]_  = (~\m7_data_i[0]  | ~\new_[18112]_ ) & (~\m0_data_i[0]  | ~\new_[18020]_ );
  assign \new_[12718]_  = (~\new_[17219]_  | ~\m2_addr_i[31] ) & (~\new_[18905]_  | ~\new_[31447]_ );
  assign \new_[12719]_  = (~\new_[18113]_  | ~\m7_addr_i[31] ) & (~\new_[18020]_  | ~\m0_addr_i[31] );
  assign \new_[12720]_  = (~\new_[18030]_  | ~\m6_addr_i[25] ) & (~\new_[18738]_  | ~\m5_addr_i[25] );
  assign \new_[12721]_  = ~\new_[26543]_  & (~\new_[16258]_  | ~\new_[29159]_ );
  assign \new_[12722]_  = (~\new_[17219]_  | ~\new_[31486]_ ) & (~\new_[18905]_  | ~\new_[31308]_ );
  assign \new_[12723]_  = ~\new_[27896]_  & (~\new_[16259]_  | ~\new_[30000]_ );
  assign \new_[12724]_  = ~\new_[24570]_  & (~\new_[16266]_  | ~\new_[29168]_ );
  assign \new_[12725]_  = (~\new_[16291]_  | ~\m2_addr_i[29] ) & (~\new_[18905]_  | ~\new_[31538]_ );
  assign \new_[12726]_  = ~\new_[28489]_  & (~\new_[16260]_  | ~\new_[30446]_ );
  assign \new_[12727]_  = (~\new_[18113]_  | ~\new_[30577]_ ) & (~\new_[18020]_  | ~\new_[30957]_ );
  assign \new_[12728]_  = (~\new_[18030]_  | ~\m6_addr_i[24] ) & (~\new_[18738]_  | ~\m5_addr_i[24] );
  assign \new_[12729]_  = (~\new_[18792]_  | ~\m6_addr_i[28] ) & (~\new_[17194]_  | ~\new_[31276]_ );
  assign \new_[12730]_  = (~\new_[18113]_  | ~\m7_addr_i[27] ) & (~\new_[18020]_  | ~\m0_addr_i[27] );
  assign \new_[12731]_  = (~\new_[17219]_  | ~\m2_addr_i[27] ) & (~\new_[18905]_  | ~\m1_addr_i[27] );
  assign \new_[12732]_  = (~\new_[17265]_  | ~\m4_addr_i[27] ) & (~\new_[18849]_  | ~\m3_addr_i[27] );
  assign \new_[12733]_  = (~\new_[18792]_  | ~\m6_addr_i[27] ) & (~\new_[17194]_  | ~\m5_addr_i[27] );
  assign \new_[12734]_  = (~\new_[18113]_  | ~\m7_addr_i[26] ) & (~\new_[18020]_  | ~\m0_addr_i[26] );
  assign \new_[12735]_  = (~\new_[17219]_  | ~\m2_addr_i[26] ) & (~\new_[18905]_  | ~\m1_addr_i[26] );
  assign \new_[12736]_  = (~\new_[18792]_  | ~\m6_addr_i[26] ) & (~\new_[17194]_  | ~\m5_addr_i[26] );
  assign \new_[12737]_  = (~\new_[18113]_  | ~\m7_addr_i[25] ) & (~\new_[18020]_  | ~\m0_addr_i[25] );
  assign \new_[12738]_  = (~\new_[17219]_  | ~\m2_addr_i[25] ) & (~\new_[18905]_  | ~\m1_addr_i[25] );
  assign \new_[12739]_  = ~\new_[26548]_  & (~\new_[16263]_  | ~\new_[28877]_ );
  assign \new_[12740]_  = (~\new_[18792]_  | ~\m6_addr_i[25] ) & (~\new_[17194]_  | ~\m5_addr_i[25] );
  assign \new_[12741]_  = (~\new_[18113]_  | ~\m7_addr_i[24] ) & (~\new_[18020]_  | ~\m0_addr_i[24] );
  assign \new_[12742]_  = (~\new_[17219]_  | ~\m2_addr_i[24] ) & (~\new_[18905]_  | ~\m1_addr_i[24] );
  assign \new_[12743]_  = ~\new_[28794]_  & (~\new_[16264]_  | ~\new_[30554]_ );
  assign \new_[12744]_  = (~\new_[18792]_  | ~\m6_addr_i[24] ) & (~\new_[17194]_  | ~\m5_addr_i[24] );
  assign \new_[12745]_  = (~\m7_addr_i[23]  | ~\new_[18112]_ ) & (~\m0_addr_i[23]  | ~\new_[18019]_ );
  assign \new_[12746]_  = (~\m7_addr_i[22]  | ~\new_[18112]_ ) & (~\m0_addr_i[22]  | ~\new_[18019]_ );
  assign \new_[12747]_  = ~\new_[27923]_  & (~\new_[16269]_  | ~\new_[29787]_ );
  assign \new_[12748]_  = ~\new_[26961]_  & (~\new_[16261]_  | ~\new_[28337]_ );
  assign \new_[12749]_  = (~\m7_addr_i[21]  | ~\new_[18112]_ ) & (~\m0_addr_i[21]  | ~\new_[18019]_ );
  assign \new_[12750]_  = ~\new_[28216]_  & (~\new_[16265]_  | ~\new_[28985]_ );
  assign \new_[12751]_  = ~\new_[28583]_  & (~\new_[16267]_  | ~\new_[30751]_ );
  assign \new_[12752]_  = (~\m7_addr_i[20]  | ~\new_[18112]_ ) & (~\m0_addr_i[20]  | ~\new_[18019]_ );
  assign \new_[12753]_  = (~\m2_addr_i[20]  | ~\new_[16291]_ ) & (~\m1_addr_i[20]  | ~\new_[18905]_ );
  assign \new_[12754]_  = (~\m7_addr_i[19]  | ~\new_[18112]_ ) & (~\m0_addr_i[19]  | ~\new_[18019]_ );
  assign \new_[12755]_  = (~\m2_addr_i[19]  | ~\new_[16291]_ ) & (~\m1_addr_i[19]  | ~\new_[18905]_ );
  assign \new_[12756]_  = (~\m2_data_i[11]  | ~\new_[18078]_ ) & (~\m1_data_i[11]  | ~\new_[18185]_ );
  assign \new_[12757]_  = (~\m5_data_i[6]  | ~\new_[18755]_ ) & (~\m6_data_i[6]  | ~\new_[17213]_ );
  assign \new_[12758]_  = (~\m7_addr_i[18]  | ~\new_[18112]_ ) & (~\m0_addr_i[18]  | ~\new_[18019]_ );
  assign \new_[12759]_  = (~\m2_addr_i[18]  | ~\new_[16291]_ ) & (~\m1_addr_i[18]  | ~\new_[18905]_ );
  assign \new_[12760]_  = ~\new_[27378]_  & (~\new_[16262]_  | ~\new_[30411]_ );
  assign \new_[12761]_  = (~\m5_addr_i[19]  | ~\new_[18738]_ ) & (~\m6_addr_i[19]  | ~\new_[18031]_ );
  assign \new_[12762]_  = ~\new_[28240]_  & (~\new_[16270]_  | ~\new_[30727]_ );
  assign \new_[12763]_  = (~\m7_addr_i[17]  | ~\new_[18112]_ ) & (~\m0_addr_i[17]  | ~\new_[18019]_ );
  assign \new_[12764]_  = (~\m2_addr_i[17]  | ~\new_[16291]_ ) & (~\m1_addr_i[17]  | ~\new_[18905]_ );
  assign \new_[12765]_  = ~\new_[28286]_  & (~\new_[16268]_  | ~\new_[29455]_ );
  assign \new_[12766]_  = (~\m7_addr_i[16]  | ~\new_[18113]_ ) & (~\m0_addr_i[16]  | ~\new_[18019]_ );
  assign \new_[12767]_  = (~\m5_addr_i[18]  | ~\new_[18738]_ ) & (~\m6_addr_i[18]  | ~\new_[16285]_ );
  assign \new_[12768]_  = (~\m7_addr_i[15]  | ~\new_[18113]_ ) & (~\m0_addr_i[15]  | ~\new_[18019]_ );
  assign \new_[12769]_  = (~\m7_addr_i[14]  | ~\new_[18112]_ ) & (~\m0_addr_i[14]  | ~\new_[18019]_ );
  assign \new_[12770]_  = ~\new_[27925]_  & (~\new_[16243]_  | ~\new_[17407]_ );
  assign \new_[12771]_  = (~\m5_addr_i[17]  | ~\new_[18738]_ ) & (~\m6_addr_i[17]  | ~\new_[18031]_ );
  assign \new_[12772]_  = (~\m7_addr_i[13]  | ~\new_[18112]_ ) & (~\m0_addr_i[13]  | ~\new_[18019]_ );
  assign \new_[12773]_  = (~\m7_addr_i[12]  | ~\new_[18112]_ ) & (~\m0_addr_i[12]  | ~\new_[18019]_ );
  assign \new_[12774]_  = ~\new_[27940]_  & (~\new_[16244]_  | ~\new_[19439]_ );
  assign \new_[12775]_  = (~\m7_addr_i[11]  | ~\new_[18112]_ ) & (~\m0_addr_i[11]  | ~\new_[18019]_ );
  assign \new_[12776]_  = (~\m5_addr_i[16]  | ~\new_[18738]_ ) & (~\m6_addr_i[16]  | ~\new_[18031]_ );
  assign \new_[12777]_  = (~\m7_data_i[9]  | ~\new_[18107]_ ) & (~\m0_data_i[9]  | ~\new_[18026]_ );
  assign \new_[12778]_  = (~\m7_addr_i[10]  | ~\new_[18112]_ ) & (~\m0_addr_i[10]  | ~\new_[18019]_ );
  assign \new_[12779]_  = ~\new_[26925]_  & (~\new_[16246]_  | ~\new_[17489]_ );
  assign \new_[12780]_  = (~\m7_addr_i[9]  | ~\new_[18112]_ ) & (~\m0_addr_i[9]  | ~\new_[18019]_ );
  assign \new_[12781]_  = (~\m5_addr_i[15]  | ~\new_[18738]_ ) & (~\m6_addr_i[15]  | ~\new_[18031]_ );
  assign \new_[12782]_  = (~\m2_addr_i[8]  | ~\new_[17219]_ ) & (~\m1_addr_i[8]  | ~\new_[18905]_ );
  assign \new_[12783]_  = ~\new_[22685]_  & (~\new_[16049]_  | ~\new_[28835]_ );
  assign \new_[12784]_  = ~\new_[29689]_  & (~\new_[16248]_  | ~\new_[19304]_ );
  assign \new_[12785]_  = (~\m7_data_i[2]  | ~\new_[18095]_ ) & (~\m0_data_i[2]  | ~\new_[20545]_ );
  assign \new_[12786]_  = (~\m7_addr_i[7]  | ~\new_[18112]_ ) & (~\m0_addr_i[7]  | ~\new_[18019]_ );
  assign \new_[12787]_  = (~\m5_addr_i[14]  | ~\new_[18738]_ ) & (~\m6_addr_i[14]  | ~\new_[18031]_ );
  assign \new_[12788]_  = (~\m2_addr_i[7]  | ~\new_[16291]_ ) & (~\m1_addr_i[7]  | ~\new_[18905]_ );
  assign \new_[12789]_  = ~\new_[17125]_  | ~\new_[29925]_  | ~\new_[29922]_  | ~\new_[30022]_ ;
  assign \new_[12790]_  = (~\m7_addr_i[6]  | ~\new_[18112]_ ) & (~\m0_addr_i[6]  | ~\new_[18019]_ );
  assign \new_[12791]_  = ~\new_[15712]_  | (~\new_[30409]_  & ~\new_[31429]_ );
  assign \new_[12792]_  = (~\m2_addr_i[6]  | ~\new_[17219]_ ) & (~\m1_addr_i[6]  | ~\new_[18905]_ );
  assign \new_[12793]_  = (~\m5_addr_i[13]  | ~\new_[18738]_ ) & (~\m6_addr_i[13]  | ~\new_[16285]_ );
  assign \new_[12794]_  = (~\m7_addr_i[5]  | ~\new_[18112]_ ) & (~\new_[31848]_  | ~\new_[18019]_ );
  assign \new_[12795]_  = (~\new_[16158]_  | ~\new_[29212]_ ) & (~\new_[30270]_  | ~\new_[31394]_ );
  assign \new_[12796]_  = ~\new_[17119]_  | ~\new_[28730]_  | ~\new_[29682]_  | ~\new_[29593]_ ;
  assign \new_[12797]_  = ~\new_[15744]_  | (~\new_[29682]_  & ~\new_[31033]_ );
  assign \new_[12798]_  = (~\m7_addr_i[4]  | ~\new_[18113]_ ) & (~\m0_addr_i[4]  | ~\new_[18020]_ );
  assign \new_[12799]_  = (~\m2_addr_i[4]  | ~\new_[16291]_ ) & (~\m1_addr_i[4]  | ~\new_[18905]_ );
  assign \new_[12800]_  = (~\new_[31726]_  | ~\new_[18113]_ ) & (~\m0_addr_i[3]  | ~\new_[18020]_ );
  assign \new_[12801]_  = ~\new_[27857]_  & (~\new_[16249]_  | ~\new_[21463]_ );
  assign \new_[12802]_  = (~\m4_addr_i[6]  | ~\new_[17260]_ ) & (~\m3_addr_i[6]  | ~\new_[18175]_ );
  assign \new_[12803]_  = (~\m7_addr_i[2]  | ~\new_[18113]_ ) & (~\m0_addr_i[2]  | ~\new_[18020]_ );
  assign \new_[12804]_  = (~\m2_addr_i[2]  | ~\new_[16291]_ ) & (~\m1_addr_i[2]  | ~\new_[18905]_ );
  assign \new_[12805]_  = (~\m4_addr_i[2]  | ~\new_[17265]_ ) & (~\m3_addr_i[2]  | ~\new_[18128]_ );
  assign \new_[12806]_  = (~\m5_addr_i[11]  | ~\new_[18738]_ ) & (~\m6_addr_i[11]  | ~\new_[18031]_ );
  assign \new_[12807]_  = (~\m7_addr_i[1]  | ~\new_[18113]_ ) & (~\m0_addr_i[1]  | ~\new_[18019]_ );
  assign \new_[12808]_  = (~\m2_addr_i[1]  | ~\new_[16291]_ ) & (~\m1_addr_i[1]  | ~\new_[18905]_ );
  assign \new_[12809]_  = ~\new_[28975]_  & (~\new_[16252]_  | ~\new_[22977]_ );
  assign \new_[12810]_  = (~\m2_addr_i[0]  | ~\new_[17219]_ ) & (~\m1_addr_i[0]  | ~\new_[18905]_ );
  assign \new_[12811]_  = ~\new_[17120]_  | ~\new_[30045]_  | ~\new_[30083]_  | ~\new_[28039]_ ;
  assign \new_[12812]_  = (~\m2_sel_i[3]  | ~\new_[17219]_ ) & (~\m1_sel_i[3]  | ~\new_[18905]_ );
  assign \new_[12813]_  = (~\m5_addr_i[10]  | ~\new_[18738]_ ) & (~\m6_addr_i[10]  | ~\new_[16285]_ );
  assign \new_[12814]_  = ~\new_[22815]_  & (~\new_[16085]_  | ~\new_[28911]_ );
  assign \new_[12815]_  = ~\new_[29060]_  & (~\new_[16250]_  | ~\new_[19422]_ );
  assign \new_[12816]_  = (~\m2_sel_i[2]  | ~\new_[17219]_ ) & (~\m1_sel_i[2]  | ~\new_[18905]_ );
  assign \new_[12817]_  = (~\m5_addr_i[9]  | ~\new_[18738]_ ) & (~\m6_addr_i[9]  | ~\new_[18031]_ );
  assign \new_[12818]_  = (~\m7_sel_i[1]  | ~\new_[18112]_ ) & (~\m0_sel_i[1]  | ~\new_[18019]_ );
  assign \new_[12819]_  = (~\m7_sel_i[0]  | ~\new_[18112]_ ) & (~\m0_sel_i[0]  | ~\new_[18020]_ );
  assign \new_[12820]_  = ~\new_[26582]_  & (~\new_[16245]_  | ~\new_[19440]_ );
  assign \new_[12821]_  = (~m7_we_i | ~\new_[18113]_ ) & (~m0_we_i | ~\new_[18020]_ );
  assign \new_[12822]_  = (~\m5_addr_i[8]  | ~\new_[18738]_ ) & (~\m6_addr_i[8]  | ~\new_[16285]_ );
  assign \new_[12823]_  = (~m4_we_i | ~\new_[17265]_ ) & (~m3_we_i | ~\new_[17248]_ );
  assign \new_[12824]_  = ~\new_[26670]_  & (~\new_[16251]_  | ~\new_[17404]_ );
  assign \new_[12825]_  = (~\m5_addr_i[7]  | ~\new_[18738]_ ) & (~\m6_addr_i[7]  | ~\new_[18031]_ );
  assign \new_[12826]_  = (~\m7_data_i[29]  | ~\new_[18112]_ ) & (~\m0_data_i[29]  | ~\new_[18019]_ );
  assign \new_[12827]_  = (~\m5_addr_i[6]  | ~\new_[18738]_ ) & (~\m6_addr_i[6]  | ~\new_[18031]_ );
  assign \new_[12828]_  = ~\new_[27701]_  & (~\new_[16247]_  | ~\new_[17410]_ );
  assign \new_[12829]_  = (~\m5_addr_i[5]  | ~\new_[18738]_ ) & (~\m6_addr_i[5]  | ~\new_[16285]_ );
  assign \new_[12830]_  = (~\m5_data_i[31]  | ~\new_[18737]_ ) & (~\m6_data_i[31]  | ~\new_[16286]_ );
  assign \new_[12831]_  = (~\m5_data_i[30]  | ~\new_[17190]_ ) & (~\m6_data_i[30]  | ~\new_[16286]_ );
  assign \new_[12832]_  = ~\new_[17136]_  | ~\new_[30220]_  | ~\new_[30138]_  | ~\new_[28935]_ ;
  assign \new_[12833]_  = (~\m5_data_i[29]  | ~\new_[17190]_ ) & (~\m6_data_i[29]  | ~\new_[16286]_ );
  assign \new_[12834]_  = ~\new_[27861]_  & (~\new_[16253]_  | ~\new_[22932]_ );
  assign \new_[12835]_  = (~\m5_addr_i[4]  | ~\new_[18738]_ ) & (~\m6_addr_i[4]  | ~\new_[18031]_ );
  assign \new_[12836]_  = (~\m5_data_i[28]  | ~\new_[17191]_ ) & (~\m6_data_i[28]  | ~\new_[16286]_ );
  assign \new_[12837]_  = ~\new_[26765]_  & (~\new_[16254]_  | ~\new_[17416]_ );
  assign \new_[12838]_  = (~\m5_data_i[27]  | ~\new_[17191]_ ) & (~\m6_data_i[27]  | ~\new_[16286]_ );
  assign \new_[12839]_  = (~\m5_addr_i[3]  | ~\new_[18738]_ ) & (~\m6_addr_i[3]  | ~\new_[16285]_ );
  assign \new_[12840]_  = ~\new_[17131]_  | ~\new_[28282]_  | ~\new_[28889]_  | ~\new_[28280]_ ;
  assign \new_[12841]_  = (~\m5_data_i[26]  | ~\new_[17191]_ ) & (~\m6_data_i[26]  | ~\new_[16286]_ );
  assign \new_[12842]_  = (~\m5_data_i[25]  | ~\new_[17190]_ ) & (~\m6_data_i[25]  | ~\new_[16286]_ );
  assign \new_[12843]_  = ~\new_[28006]_  & (~\new_[16256]_  | ~\new_[21511]_ );
  assign \new_[12844]_  = (~\m5_addr_i[2]  | ~\new_[18738]_ ) & (~\m6_addr_i[2]  | ~\new_[18031]_ );
  assign \new_[12845]_  = (~\m5_data_i[24]  | ~\new_[17191]_ ) & (~\m6_data_i[24]  | ~\new_[16286]_ );
  assign \new_[12846]_  = (~\m5_addr_i[1]  | ~\new_[18738]_ ) & (~\m6_addr_i[1]  | ~\new_[18031]_ );
  assign \new_[12847]_  = (~\m5_data_i[23]  | ~\new_[17191]_ ) & (~\m6_data_i[23]  | ~\new_[16286]_ );
  assign \new_[12848]_  = ~\new_[29752]_  & (~\new_[16255]_  | ~\new_[21578]_ );
  assign \new_[12849]_  = (~\m5_data_i[22]  | ~\new_[17191]_ ) & (~\m6_data_i[22]  | ~\new_[16286]_ );
  assign \new_[12850]_  = (~\m5_data_i[21]  | ~\new_[17191]_ ) & (~\m6_data_i[21]  | ~\new_[16286]_ );
  assign \new_[12851]_  = (~\m5_addr_i[0]  | ~\new_[18738]_ ) & (~\m6_addr_i[0]  | ~\new_[18031]_ );
  assign \new_[12852]_  = (~\m5_data_i[20]  | ~\new_[17191]_ ) & (~\m6_data_i[20]  | ~\new_[16286]_ );
  assign \new_[12853]_  = (~\m2_data_i[25]  | ~\new_[18077]_ ) & (~\m1_data_i[25]  | ~\new_[18182]_ );
  assign \new_[12854]_  = (~\m5_data_i[19]  | ~\new_[18737]_ ) & (~\m6_data_i[19]  | ~\new_[18032]_ );
  assign \new_[12855]_  = (~\m5_sel_i[3]  | ~\new_[18738]_ ) & (~\m6_sel_i[3]  | ~\new_[18031]_ );
  assign \new_[12856]_  = ~\new_[17030]_  | ~\new_[17031]_  | ~\new_[14616]_  | ~\new_[16149]_ ;
  assign \new_[12857]_  = (~\m5_data_i[18]  | ~\new_[17191]_ ) & (~\m6_data_i[18]  | ~\new_[16286]_ );
  assign \new_[12858]_  = (~\m5_data_i[17]  | ~\new_[17191]_ ) & (~\m6_data_i[17]  | ~\new_[16286]_ );
  assign \new_[12859]_  = (~\m5_data_i[16]  | ~\new_[17191]_ ) & (~\m6_data_i[16]  | ~\new_[18032]_ );
  assign \new_[12860]_  = (~\m5_sel_i[1]  | ~\new_[18738]_ ) & (~\m6_sel_i[1]  | ~\new_[16285]_ );
  assign \new_[12861]_  = (~\m5_data_i[15]  | ~\new_[18737]_ ) & (~\m6_data_i[15]  | ~\new_[16286]_ );
  assign \new_[12862]_  = ~\new_[16863]_  | ~\new_[17732]_  | ~\new_[14653]_  | ~\new_[17728]_ ;
  assign \new_[12863]_  = ~\new_[16875]_  | ~\new_[17736]_  | ~\new_[14661]_  | ~\new_[17735]_ ;
  assign \new_[12864]_  = (~\m5_data_i[14]  | ~\new_[18737]_ ) & (~\m6_data_i[14]  | ~\new_[16286]_ );
  assign \new_[12865]_  = ~\new_[16880]_  | ~\new_[17739]_  | ~\new_[16879]_  | ~\new_[18569]_ ;
  assign \new_[12866]_  = (~\m5_data_i[13]  | ~\new_[18737]_ ) & (~\m6_data_i[13]  | ~\new_[16286]_ );
  assign \new_[12867]_  = (~\m5_sel_i[0]  | ~\new_[18738]_ ) & (~\m6_sel_i[0]  | ~\new_[18031]_ );
  assign \new_[12868]_  = (~\new_[16077]_  | ~s2_err_i) & (~\new_[18578]_  | ~s1_err_i);
  assign \new_[12869]_  = (~\m5_data_i[12]  | ~\new_[18737]_ ) & (~\m6_data_i[12]  | ~\new_[16286]_ );
  assign \new_[12870]_  = (~\new_[17759]_  | ~s4_err_i) & (~\new_[16079]_  | ~s0_err_i);
  assign \new_[12871]_  = (~\m5_data_i[11]  | ~\new_[18737]_ ) & (~\m6_data_i[11]  | ~\new_[16286]_ );
  assign \new_[12872]_  = (~\new_[18660]_  | ~s10_err_i) & (~\new_[16179]_  | ~s9_err_i);
  assign \new_[12873]_  = (~m5_we_i | ~\new_[18738]_ ) & (~m6_we_i | ~\new_[16285]_ );
  assign \new_[12874]_  = (~\m4_data_i[10]  | ~\new_[17272]_ ) & (~\m3_data_i[10]  | ~\new_[17280]_ );
  assign \new_[12875]_  = (~\m5_data_i[10]  | ~\new_[18737]_ ) & (~\m6_data_i[10]  | ~\new_[16286]_ );
  assign \new_[12876]_  = (~\new_[16077]_  | ~s2_rty_i) & (~\new_[18578]_  | ~s1_rty_i);
  assign \new_[12877]_  = (~\m4_data_i[9]  | ~\new_[17272]_ ) & (~\m3_data_i[9]  | ~\new_[17280]_ );
  assign \new_[12878]_  = (~\m5_data_i[9]  | ~\new_[18737]_ ) & (~\m6_data_i[9]  | ~\new_[16286]_ );
  assign \new_[12879]_  = (~\new_[18660]_  | ~s10_rty_i) & (~\new_[16179]_  | ~s9_rty_i);
  assign \new_[12880]_  = (~\m7_data_i[31]  | ~\new_[19584]_ ) & (~\m0_data_i[31]  | ~\new_[18026]_ );
  assign \new_[12881]_  = (~\m5_data_i[8]  | ~\new_[17190]_ ) & (~\m6_data_i[8]  | ~\new_[16286]_ );
  assign \new_[12882]_  = (~\m5_data_i[7]  | ~\new_[17190]_ ) & (~\m6_data_i[7]  | ~\new_[18032]_ );
  assign \new_[12883]_  = (~\new_[17759]_  | ~s4_rty_i) & (~\new_[16079]_  | ~s0_rty_i);
  assign \new_[12884]_  = (~\m5_data_i[6]  | ~\new_[18737]_ ) & (~\m6_data_i[6]  | ~\new_[16286]_ );
  assign \new_[12885]_  = (~\m5_data_i[5]  | ~\new_[18737]_ ) & (~\m6_data_i[5]  | ~\new_[16286]_ );
  assign \new_[12886]_  = ~\new_[17051]_  | ~\new_[17052]_  | ~\new_[16172]_  | ~\new_[17873]_ ;
  assign \new_[12887]_  = (~\m5_data_i[4]  | ~\new_[17190]_ ) & (~\m6_data_i[4]  | ~\new_[18032]_ );
  assign \new_[12888]_  = (~\m7_addr_i[6]  | ~\new_[18115]_ ) & (~\m0_addr_i[6]  | ~\new_[19637]_ );
  assign \new_[12889]_  = (~\m4_data_i[3]  | ~\new_[17272]_ ) & (~\m3_data_i[3]  | ~\new_[17280]_ );
  assign \new_[12890]_  = (~\m5_data_i[3]  | ~\new_[18737]_ ) & (~\m6_data_i[3]  | ~\new_[16286]_ );
  assign \new_[12891]_  = (~\m5_data_i[2]  | ~\new_[18737]_ ) & (~\m6_data_i[2]  | ~\new_[16286]_ );
  assign \new_[12892]_  = (~\m4_data_i[1]  | ~\new_[17272]_ ) & (~\m3_data_i[1]  | ~\new_[17280]_ );
  assign \new_[12893]_  = (~\m5_data_i[1]  | ~\new_[18737]_ ) & (~\m6_data_i[1]  | ~\new_[16286]_ );
  assign \new_[12894]_  = ~\new_[17101]_  | ~\new_[18662]_  | ~\new_[16188]_  | ~\new_[17890]_ ;
  assign \new_[12895]_  = (~\m7_data_i[31]  | ~\new_[18825]_ ) & (~\m0_data_i[31]  | ~\new_[18010]_ );
  assign \new_[12896]_  = ~\new_[17063]_  | ~\new_[18663]_  | ~\new_[16146]_  | ~\new_[17879]_ ;
  assign \new_[12897]_  = (~\m5_data_i[0]  | ~\new_[18737]_ ) & (~\m6_data_i[0]  | ~\new_[16286]_ );
  assign \new_[12898]_  = (~\new_[16286]_  | ~\m6_addr_i[31] ) & (~\new_[17192]_  | ~\new_[31001]_ );
  assign \new_[12899]_  = (~\new_[16286]_  | ~\m6_addr_i[30] ) & (~\new_[17192]_  | ~\new_[31147]_ );
  assign \new_[12900]_  = (~\m4_data_i[30]  | ~\new_[16305]_ ) & (~\m3_data_i[30]  | ~\new_[18200]_ );
  assign \new_[12901]_  = (~\new_[16286]_  | ~\m6_addr_i[29] ) & (~\new_[17192]_  | ~\new_[31407]_ );
  assign \new_[12902]_  = (~\m7_data_i[11]  | ~\new_[18108]_ ) & (~\m0_data_i[11]  | ~\new_[18026]_ );
  assign \new_[12903]_  = (~\m4_data_i[29]  | ~\new_[16305]_ ) & (~\m3_data_i[29]  | ~\new_[18200]_ );
  assign \new_[12904]_  = (~\new_[16286]_  | ~\m6_addr_i[28] ) & (~\new_[17192]_  | ~\new_[31276]_ );
  assign \new_[12905]_  = (~\new_[16286]_  | ~\m6_addr_i[27] ) & (~\new_[17192]_  | ~\m5_addr_i[27] );
  assign \new_[12906]_  = (~\m7_addr_i[15]  | ~\new_[18099]_ ) & (~\m0_addr_i[15]  | ~\new_[18026]_ );
  assign \new_[12907]_  = ~\new_[17072]_  | ~\new_[17073]_  | ~\new_[17070]_  | ~\new_[17071]_ ;
  assign \new_[12908]_  = (~\new_[16286]_  | ~\m6_addr_i[26] ) & (~\new_[17192]_  | ~\m5_addr_i[26] );
  assign \new_[12909]_  = (~\new_[16286]_  | ~\m6_addr_i[25] ) & (~\new_[17192]_  | ~\m5_addr_i[25] );
  assign \new_[12910]_  = ~\new_[17095]_  | ~\new_[17096]_  | ~\new_[17887]_  | ~\new_[16218]_ ;
  assign \new_[12911]_  = (~\m2_data_i[27]  | ~\new_[17216]_ ) & (~\m1_data_i[27]  | ~\new_[18888]_ );
  assign \new_[12912]_  = ~\new_[17103]_  | ~\new_[18667]_  | ~\new_[17099]_  | ~\new_[17100]_ ;
  assign \new_[12913]_  = (~\new_[16286]_  | ~\m6_addr_i[24] ) & (~\new_[17192]_  | ~\m5_addr_i[24] );
  assign \new_[12914]_  = (~\m5_addr_i[23]  | ~\new_[17191]_ ) & (~\m6_addr_i[23]  | ~\new_[16286]_ );
  assign \new_[12915]_  = (~\m5_addr_i[22]  | ~\new_[17191]_ ) & (~\m6_addr_i[22]  | ~\new_[16286]_ );
  assign \new_[12916]_  = (~\m7_data_i[25]  | ~\new_[18825]_ ) & (~\m0_data_i[25]  | ~\new_[18010]_ );
  assign \new_[12917]_  = (~\m5_addr_i[21]  | ~\new_[17191]_ ) & (~\m6_addr_i[21]  | ~\new_[16286]_ );
  assign \new_[12918]_  = (~\m5_addr_i[20]  | ~\new_[17191]_ ) & (~\m6_addr_i[20]  | ~\new_[16286]_ );
  assign \new_[12919]_  = (~\m4_data_i[25]  | ~\new_[18877]_ ) & (~\m3_data_i[25]  | ~\new_[18200]_ );
  assign \new_[12920]_  = (~\m5_addr_i[19]  | ~\new_[17191]_ ) & (~\m6_addr_i[19]  | ~\new_[16286]_ );
  assign \new_[12921]_  = (~\m7_data_i[24]  | ~\new_[18824]_ ) & (~\m0_data_i[24]  | ~\new_[18010]_ );
  assign \new_[12922]_  = (~\m5_addr_i[18]  | ~\new_[18737]_ ) & (~\m6_addr_i[18]  | ~\new_[16286]_ );
  assign \new_[12923]_  = (~\m4_data_i[24]  | ~\new_[18877]_ ) & (~\m3_data_i[24]  | ~\new_[18200]_ );
  assign \new_[12924]_  = (~\m5_addr_i[17]  | ~\new_[17191]_ ) & (~\m6_addr_i[17]  | ~\new_[16286]_ );
  assign \new_[12925]_  = (~\m7_data_i[23]  | ~\new_[18825]_ ) & (~\m0_data_i[23]  | ~\new_[18010]_ );
  assign \new_[12926]_  = (~\m4_data_i[23]  | ~\new_[18877]_ ) & (~\m3_data_i[23]  | ~\new_[18200]_ );
  assign \new_[12927]_  = (~\m5_addr_i[16]  | ~\new_[17191]_ ) & (~\m6_addr_i[16]  | ~\new_[16286]_ );
  assign \new_[12928]_  = (~\m5_addr_i[15]  | ~\new_[18737]_ ) & (~\m6_addr_i[15]  | ~\new_[18032]_ );
  assign \new_[12929]_  = (~\m7_data_i[22]  | ~\new_[18825]_ ) & (~\m0_data_i[22]  | ~\new_[18010]_ );
  assign \new_[12930]_  = (~\m4_data_i[22]  | ~\new_[16305]_ ) & (~\m3_data_i[22]  | ~\new_[19638]_ );
  assign \new_[12931]_  = (~\m5_addr_i[14]  | ~\new_[17191]_ ) & (~\m6_addr_i[14]  | ~\new_[16286]_ );
  assign \new_[12932]_  = (~\m5_addr_i[13]  | ~\new_[17191]_ ) & (~\m6_addr_i[13]  | ~\new_[16286]_ );
  assign \new_[12933]_  = (~\m7_data_i[21]  | ~\new_[18825]_ ) & (~\m0_data_i[21]  | ~\new_[18010]_ );
  assign \new_[12934]_  = (~\m4_data_i[21]  | ~\new_[16305]_ ) & (~\m3_data_i[21]  | ~\new_[18200]_ );
  assign \new_[12935]_  = (~\m5_addr_i[12]  | ~\new_[17191]_ ) & (~\m6_addr_i[12]  | ~\new_[16286]_ );
  assign \new_[12936]_  = (~\m5_addr_i[11]  | ~\new_[17191]_ ) & (~\m6_addr_i[11]  | ~\new_[16286]_ );
  assign \new_[12937]_  = (~\m5_addr_i[10]  | ~\new_[17191]_ ) & (~\m6_addr_i[10]  | ~\new_[16286]_ );
  assign \new_[12938]_  = (~\m4_data_i[20]  | ~\new_[16305]_ ) & (~\m3_data_i[20]  | ~\new_[18200]_ );
  assign \new_[12939]_  = (~\m5_addr_i[13]  | ~\new_[18748]_ ) & (~\m6_addr_i[13]  | ~\new_[17213]_ );
  assign \new_[12940]_  = (~\m5_addr_i[9]  | ~\new_[17191]_ ) & (~\m6_addr_i[9]  | ~\new_[16286]_ );
  assign \new_[12941]_  = (~\m5_data_i[19]  | ~\new_[18738]_ ) & (~\m6_data_i[19]  | ~\new_[18031]_ );
  assign \new_[12942]_  = (~\m7_addr_i[14]  | ~\new_[18099]_ ) & (~\m0_addr_i[14]  | ~\new_[18026]_ );
  assign \new_[12943]_  = (~\m5_addr_i[8]  | ~\new_[17191]_ ) & (~\m6_addr_i[8]  | ~\new_[16286]_ );
  assign \new_[12944]_  = (~\m7_data_i[18]  | ~\new_[18824]_ ) & (~\m0_data_i[18]  | ~\new_[18010]_ );
  assign \new_[12945]_  = (~\m5_addr_i[7]  | ~\new_[17191]_ ) & (~\m6_addr_i[7]  | ~\new_[16286]_ );
  assign \new_[12946]_  = (~\m5_addr_i[6]  | ~\new_[17191]_ ) & (~\m6_addr_i[6]  | ~\new_[16286]_ );
  assign \new_[12947]_  = (~\m4_addr_i[5]  | ~\new_[17272]_ ) & (~\m3_addr_i[5]  | ~\new_[17280]_ );
  assign \new_[12948]_  = (~\m5_addr_i[5]  | ~\new_[18737]_ ) & (~\m6_addr_i[5]  | ~\new_[18032]_ );
  assign \new_[12949]_  = (~\m7_data_i[17]  | ~\new_[18825]_ ) & (~\m0_data_i[17]  | ~\new_[18010]_ );
  assign \new_[12950]_  = (~\m5_addr_i[4]  | ~\new_[17190]_ ) & (~\m6_addr_i[4]  | ~\new_[18032]_ );
  assign \new_[12951]_  = (~\m4_data_i[17]  | ~\new_[16305]_ ) & (~\m3_data_i[17]  | ~\new_[19638]_ );
  assign \new_[12952]_  = (~\m5_addr_i[3]  | ~\new_[18737]_ ) & (~\m6_addr_i[3]  | ~\new_[16286]_ );
  assign \new_[12953]_  = (~\m7_data_i[16]  | ~\new_[18825]_ ) & (~\m0_data_i[16]  | ~\new_[18010]_ );
  assign \new_[12954]_  = \new_[14745]_  & \new_[17014]_ ;
  assign \new_[12955]_  = (~\m5_addr_i[2]  | ~\new_[17190]_ ) & (~\m6_addr_i[2]  | ~\new_[18032]_ );
  assign \new_[12956]_  = (~\m4_data_i[16]  | ~\new_[16305]_ ) & (~\m3_data_i[16]  | ~\new_[18200]_ );
  assign \new_[12957]_  = (~\m7_data_i[25]  | ~\new_[18103]_ ) & (~\m0_data_i[25]  | ~\new_[18026]_ );
  assign \new_[12958]_  = (~\m5_addr_i[1]  | ~\new_[17191]_ ) & (~\m6_addr_i[1]  | ~\new_[18032]_ );
  assign \new_[12959]_  = (~\m7_data_i[15]  | ~\new_[18824]_ ) & (~\m0_data_i[15]  | ~\new_[18011]_ );
  assign \new_[12960]_  = (~\m4_data_i[15]  | ~\new_[18877]_ ) & (~\m3_data_i[15]  | ~\new_[18200]_ );
  assign \new_[12961]_  = (~\m5_addr_i[0]  | ~\new_[17191]_ ) & (~\m6_addr_i[0]  | ~\new_[16286]_ );
  assign \new_[12962]_  = (~\m2_addr_i[0]  | ~\new_[18069]_ ) & (~\m1_addr_i[0]  | ~\new_[18900]_ );
  assign \new_[12963]_  = (~\m7_data_i[14]  | ~\new_[18824]_ ) & (~\m0_data_i[14]  | ~\new_[18011]_ );
  assign \new_[12964]_  = (~\m5_sel_i[3]  | ~\new_[17191]_ ) & (~\m6_sel_i[3]  | ~\new_[18032]_ );
  assign \new_[12965]_  = (~\m5_sel_i[2]  | ~\new_[18737]_ ) & (~\m6_sel_i[2]  | ~\new_[18032]_ );
  assign \new_[12966]_  = (~\m4_data_i[14]  | ~\new_[18877]_ ) & (~\m3_data_i[14]  | ~\new_[18200]_ );
  assign \new_[12967]_  = (~\m5_sel_i[1]  | ~\new_[17191]_ ) & (~\m6_sel_i[1]  | ~\new_[16286]_ );
  assign \new_[12968]_  = (~\m7_data_i[13]  | ~\new_[18824]_ ) & (~\m0_data_i[13]  | ~\new_[18011]_ );
  assign \new_[12969]_  = (~\m4_data_i[13]  | ~\new_[18877]_ ) & (~\m3_data_i[13]  | ~\new_[18200]_ );
  assign \new_[12970]_  = (~\m5_sel_i[0]  | ~\new_[17191]_ ) & (~\m6_sel_i[0]  | ~\new_[16286]_ );
  assign \new_[12971]_  = (~\m7_data_i[12]  | ~\new_[18824]_ ) & (~\m0_data_i[12]  | ~\new_[18011]_ );
  assign \new_[12972]_  = (~m5_we_i | ~\new_[18737]_ ) & (~m6_we_i | ~\new_[16286]_ );
  assign \new_[12973]_  = (~\m2_data_i[12]  | ~\new_[17216]_ ) & (~\m1_data_i[12]  | ~\new_[18888]_ );
  assign \new_[12974]_  = (~\m4_data_i[12]  | ~\new_[18877]_ ) & (~\m3_data_i[12]  | ~\new_[18200]_ );
  assign \new_[12975]_  = (~\m7_data_i[11]  | ~\new_[18824]_ ) & (~\m0_data_i[11]  | ~\new_[18011]_ );
  assign \new_[12976]_  = (~\m4_data_i[11]  | ~\new_[18877]_ ) & (~\m3_data_i[11]  | ~\new_[18200]_ );
  assign \new_[12977]_  = (~\m7_data_i[10]  | ~\new_[18824]_ ) & (~\m0_data_i[10]  | ~\new_[18011]_ );
  assign \new_[12978]_  = (~\m4_data_i[10]  | ~\new_[18877]_ ) & (~\m3_data_i[10]  | ~\new_[18200]_ );
  assign \new_[12979]_  = (~\m5_data_i[9]  | ~\new_[18738]_ ) & (~\m6_data_i[9]  | ~\new_[18031]_ );
  assign \new_[12980]_  = (~\m7_data_i[9]  | ~\new_[18824]_ ) & (~\m0_data_i[9]  | ~\new_[18011]_ );
  assign \new_[12981]_  = (~\m2_data_i[9]  | ~\new_[17216]_ ) & (~\m1_data_i[9]  | ~\new_[19618]_ );
  assign \new_[12982]_  = (~\m4_data_i[9]  | ~\new_[18877]_ ) & (~\m3_data_i[9]  | ~\new_[18200]_ );
  assign \new_[12983]_  = (~\m7_data_i[8]  | ~\new_[18824]_ ) & (~\m0_data_i[8]  | ~\new_[18011]_ );
  assign \new_[12984]_  = \new_[16859]_  & \new_[14652]_ ;
  assign \new_[12985]_  = (~\m2_data_i[8]  | ~\new_[17216]_ ) & (~\m1_data_i[8]  | ~\new_[19618]_ );
  assign \new_[12986]_  = (~\m4_data_i[8]  | ~\new_[18877]_ ) & (~\m3_data_i[8]  | ~\new_[18200]_ );
  assign \new_[12987]_  = (~\m7_data_i[7]  | ~\new_[18824]_ ) & (~\m0_data_i[7]  | ~\new_[18011]_ );
  assign \new_[12988]_  = (~\m2_data_i[7]  | ~\new_[17216]_ ) & (~\m1_data_i[7]  | ~\new_[19618]_ );
  assign \new_[12989]_  = (~\m4_data_i[7]  | ~\new_[18877]_ ) & (~\m3_data_i[7]  | ~\new_[18200]_ );
  assign \new_[12990]_  = (~\m7_data_i[6]  | ~\new_[18824]_ ) & (~\m0_data_i[6]  | ~\new_[18011]_ );
  assign \new_[12991]_  = (~\m2_data_i[6]  | ~\new_[17216]_ ) & (~\m1_data_i[6]  | ~\new_[19619]_ );
  assign \new_[12992]_  = (~\m4_data_i[6]  | ~\new_[18877]_ ) & (~\m3_data_i[6]  | ~\new_[18200]_ );
  assign \new_[12993]_  = (~\m7_data_i[5]  | ~\new_[18824]_ ) & (~\m0_data_i[5]  | ~\new_[18011]_ );
  assign \new_[12994]_  = (~\m2_data_i[5]  | ~\new_[17216]_ ) & (~\m1_data_i[5]  | ~\new_[19619]_ );
  assign \new_[12995]_  = (~\m4_data_i[5]  | ~\new_[18877]_ ) & (~\m3_data_i[5]  | ~\new_[18200]_ );
  assign \new_[12996]_  = (~\m7_data_i[4]  | ~\new_[18824]_ ) & (~\m0_data_i[4]  | ~\new_[18011]_ );
  assign \new_[12997]_  = (~\m2_data_i[4]  | ~\new_[17216]_ ) & (~\m1_data_i[4]  | ~\new_[19619]_ );
  assign \new_[12998]_  = (~\m4_data_i[4]  | ~\new_[18877]_ ) & (~\m3_data_i[4]  | ~\new_[18200]_ );
  assign \new_[12999]_  = (~\m7_data_i[3]  | ~\new_[18824]_ ) & (~\m0_data_i[3]  | ~\new_[18011]_ );
  assign \new_[13000]_  = (~\m4_data_i[3]  | ~\new_[18877]_ ) & (~\m3_data_i[3]  | ~\new_[18200]_ );
  assign \new_[13001]_  = (~\m7_data_i[2]  | ~\new_[18824]_ ) & (~\m0_data_i[2]  | ~\new_[18011]_ );
  assign \new_[13002]_  = (~\m2_data_i[2]  | ~\new_[17216]_ ) & (~\m1_data_i[2]  | ~\new_[19618]_ );
  assign \new_[13003]_  = (~\m4_data_i[2]  | ~\new_[18877]_ ) & (~\m3_data_i[2]  | ~\new_[18200]_ );
  assign \new_[13004]_  = (~\m7_data_i[1]  | ~\new_[18824]_ ) & (~\m0_data_i[1]  | ~\new_[18011]_ );
  assign \new_[13005]_  = (~\m4_data_i[1]  | ~\new_[18877]_ ) & (~\m3_data_i[1]  | ~\new_[18200]_ );
  assign \new_[13006]_  = ~\new_[27697]_  & (~\new_[16271]_  | ~\new_[29355]_ );
  assign \new_[13007]_  = (~\m7_data_i[0]  | ~\new_[18824]_ ) & (~\m0_data_i[0]  | ~\new_[18011]_ );
  assign \new_[13008]_  = (~\m4_data_i[0]  | ~\new_[18877]_ ) & (~\m3_data_i[0]  | ~\new_[18200]_ );
  assign \new_[13009]_  = (~\new_[18824]_  | ~\new_[31496]_ ) & (~\new_[18010]_  | ~\m0_addr_i[31] );
  assign \new_[13010]_  = (~\new_[16305]_  | ~\m4_addr_i[31] ) & (~\new_[19638]_  | ~\m3_addr_i[31] );
  assign \new_[13011]_  = ~\new_[24583]_  & (~\new_[16272]_  | ~\new_[30210]_ );
  assign \new_[13012]_  = (~\new_[18824]_  | ~\new_[31885]_ ) & (~\new_[18010]_  | ~\new_[31292]_ );
  assign \new_[13013]_  = (~\new_[16305]_  | ~\m4_addr_i[30] ) & (~\new_[18200]_  | ~\m3_addr_i[30] );
  assign \new_[13014]_  = (~\new_[18824]_  | ~\new_[31531]_ ) & (~\new_[18010]_  | ~\new_[31481]_ );
  assign \new_[13015]_  = (~\new_[16305]_  | ~\m4_addr_i[29] ) & (~\new_[19638]_  | ~\m3_addr_i[29] );
  assign \new_[13016]_  = (~\m3_addr_i[9]  | ~\new_[32350]_ ) & (~\m2_addr_i[9]  | ~\new_[17223]_ );
  assign \new_[13017]_  = (~\new_[18824]_  | ~\new_[30577]_ ) & (~\new_[18010]_  | ~\new_[30957]_ );
  assign \new_[13018]_  = (~\new_[18824]_  | ~\m7_addr_i[27] ) & (~\new_[18010]_  | ~\m0_addr_i[27] );
  assign \new_[13019]_  = (~\new_[18824]_  | ~\m7_addr_i[26] ) & (~\new_[18010]_  | ~\m0_addr_i[26] );
  assign \new_[13020]_  = (~\m7_addr_i[16]  | ~\new_[18103]_ ) & (~\m0_addr_i[16]  | ~\new_[18026]_ );
  assign \new_[13021]_  = ~m1_stb_i | ~\new_[26173]_  | ~\new_[18192]_ ;
  assign \new_[13022]_  = (~\new_[18824]_  | ~\m7_addr_i[25] ) & (~\new_[18010]_  | ~\m0_addr_i[25] );
  assign \new_[13023]_  = (~\m7_addr_i[18]  | ~\new_[18105]_ ) & (~\m0_addr_i[18]  | ~\new_[18026]_ );
  assign \new_[13024]_  = (~\new_[18824]_  | ~\m7_addr_i[24] ) & (~\new_[18010]_  | ~\m0_addr_i[24] );
  assign \new_[13025]_  = (~\m7_addr_i[17]  | ~\new_[18102]_ ) & (~\m0_addr_i[17]  | ~\new_[18026]_ );
  assign \new_[13026]_  = \new_[14706]_  & \new_[16113]_ ;
  assign \new_[13027]_  = (~\new_[16305]_  | ~\m4_addr_i[24] ) & (~\new_[19638]_  | ~\m3_addr_i[24] );
  assign \new_[13028]_  = (~\m7_addr_i[23]  | ~\new_[18825]_ ) & (~\m0_addr_i[23]  | ~\new_[18010]_ );
  assign \new_[13029]_  = \new_[14811]_  & \new_[17086]_ ;
  assign \new_[13030]_  = (~\m4_addr_i[23]  | ~\new_[16305]_ ) & (~\m3_addr_i[23]  | ~\new_[18200]_ );
  assign \new_[13031]_  = (~\m7_addr_i[22]  | ~\new_[18825]_ ) & (~\m0_addr_i[22]  | ~\new_[18010]_ );
  assign \new_[13032]_  = (~\m4_addr_i[22]  | ~\new_[16305]_ ) & (~\m3_addr_i[22]  | ~\new_[19638]_ );
  assign \new_[13033]_  = ~\new_[27555]_  & (~\new_[16273]_  | ~\new_[28850]_ );
  assign \new_[13034]_  = (~\m7_addr_i[21]  | ~\new_[18825]_ ) & (~\m0_addr_i[21]  | ~\new_[18010]_ );
  assign \new_[13035]_  = (~\m4_addr_i[21]  | ~\new_[16305]_ ) & (~\m3_addr_i[21]  | ~\new_[18200]_ );
  assign \new_[13036]_  = ~\new_[14624]_  & ~\new_[17323]_ ;
  assign \new_[13037]_  = (~\m7_addr_i[20]  | ~\new_[18825]_ ) & (~\m0_addr_i[20]  | ~\new_[18010]_ );
  assign \new_[13038]_  = ~\new_[14627]_  & ~\new_[17329]_ ;
  assign \new_[13039]_  = (~\m7_addr_i[19]  | ~\new_[18825]_ ) & (~\m0_addr_i[19]  | ~\new_[18010]_ );
  assign \new_[13040]_  = (~\m7_addr_i[18]  | ~\new_[18825]_ ) & (~\m0_addr_i[18]  | ~\new_[18010]_ );
  assign \new_[13041]_  = (~\m7_addr_i[17]  | ~\new_[18825]_ ) & (~\m0_addr_i[17]  | ~\new_[18010]_ );
  assign \new_[13042]_  = (~\m4_addr_i[17]  | ~\new_[16305]_ ) & (~\m3_addr_i[17]  | ~\new_[18200]_ );
  assign \new_[13043]_  = (~\m4_addr_i[0]  | ~\new_[17260]_ ) & (~\m3_addr_i[0]  | ~\new_[18175]_ );
  assign \new_[13044]_  = (~\m4_addr_i[16]  | ~\new_[16305]_ ) & (~\m3_addr_i[16]  | ~\new_[19638]_ );
  assign \new_[13045]_  = (~\m4_addr_i[15]  | ~\new_[16305]_ ) & (~\m3_addr_i[15]  | ~\new_[19638]_ );
  assign \new_[13046]_  = (~\m4_addr_i[14]  | ~\new_[16305]_ ) & (~\m3_addr_i[14]  | ~\new_[18200]_ );
  assign \new_[13047]_  = (~\m7_addr_i[13]  | ~\new_[18825]_ ) & (~\m0_addr_i[13]  | ~\new_[18010]_ );
  assign \new_[13048]_  = ~\new_[14611]_  & (~\new_[17295]_  | ~\new_[31564]_ );
  assign \new_[13049]_  = (~\m5_data_i[14]  | ~\new_[18759]_ ) & (~\m6_data_i[14]  | ~\new_[18787]_ );
  assign \new_[13050]_  = (~\m4_addr_i[13]  | ~\new_[16305]_ ) & (~\m3_addr_i[13]  | ~\new_[18200]_ );
  assign \new_[13051]_  = (~\m7_addr_i[12]  | ~\new_[18825]_ ) & (~\m0_addr_i[12]  | ~\new_[18010]_ );
  assign \new_[13052]_  = (~\m4_addr_i[12]  | ~\new_[16305]_ ) & (~\m3_addr_i[12]  | ~\new_[19638]_ );
  assign \new_[13053]_  = ~\new_[14618]_  & (~\new_[17301]_  | ~\new_[31846]_ );
  assign \new_[13054]_  = ~\new_[14625]_  & (~\new_[17323]_  | ~\new_[31810]_ );
  assign \new_[13055]_  = (~\m7_addr_i[10]  | ~\new_[18825]_ ) & (~\m0_addr_i[10]  | ~\new_[18010]_ );
  assign \new_[13056]_  = (~\m5_addr_i[3]  | ~\new_[18016]_ ) & (~\m6_addr_i[3]  | ~\new_[17229]_ );
  assign \new_[13057]_  = (~\m4_addr_i[9]  | ~\new_[16305]_ ) & (~\m3_addr_i[9]  | ~\new_[18200]_ );
  assign \new_[13058]_  = (~\m7_addr_i[8]  | ~\new_[18825]_ ) & (~\m0_addr_i[8]  | ~\new_[18011]_ );
  assign \new_[13059]_  = (~\m4_addr_i[8]  | ~\new_[16305]_ ) & (~\m3_addr_i[8]  | ~\new_[18200]_ );
  assign \new_[13060]_  = (~\m7_addr_i[7]  | ~\new_[18825]_ ) & (~\m0_addr_i[7]  | ~\new_[18011]_ );
  assign \new_[13061]_  = (~\m4_addr_i[6]  | ~\new_[18877]_ ) & (~\m3_addr_i[6]  | ~\new_[18200]_ );
  assign \new_[13062]_  = (~\m7_addr_i[5]  | ~\new_[18824]_ ) & (~\new_[31848]_  | ~\new_[18011]_ );
  assign \new_[13063]_  = (~\new_[31095]_  | ~\new_[17216]_ ) & (~\m1_addr_i[5]  | ~\new_[18888]_ );
  assign \new_[13064]_  = (~\m4_addr_i[5]  | ~\new_[18877]_ ) & (~\m3_addr_i[5]  | ~\new_[18200]_ );
  assign \new_[13065]_  = (~\m7_addr_i[4]  | ~\new_[18824]_ ) & (~\m0_addr_i[4]  | ~\new_[18011]_ );
  assign \new_[13066]_  = (~\m2_addr_i[4]  | ~\new_[17216]_ ) & (~\m1_addr_i[4]  | ~\new_[19618]_ );
  assign \new_[13067]_  = (~\m4_addr_i[4]  | ~\new_[18877]_ ) & (~\m3_addr_i[4]  | ~\new_[18200]_ );
  assign \new_[13068]_  = (~\new_[31726]_  | ~\new_[18824]_ ) & (~\m0_addr_i[3]  | ~\new_[18011]_ );
  assign \new_[13069]_  = (~\m4_addr_i[3]  | ~\new_[18877]_ ) & (~\m3_addr_i[3]  | ~\new_[18200]_ );
  assign \new_[13070]_  = (~\m7_addr_i[2]  | ~\new_[18824]_ ) & (~\m0_addr_i[2]  | ~\new_[18011]_ );
  assign \new_[13071]_  = (~\m2_addr_i[2]  | ~\new_[17216]_ ) & (~\new_[31477]_  | ~\new_[19618]_ );
  assign \new_[13072]_  = (~\m4_addr_i[2]  | ~\new_[18877]_ ) & (~\m3_addr_i[2]  | ~\new_[18200]_ );
  assign \new_[13073]_  = (~\m7_addr_i[1]  | ~\new_[18824]_ ) & (~\m0_addr_i[1]  | ~\new_[18010]_ );
  assign \new_[13074]_  = (~\m4_addr_i[1]  | ~\new_[16305]_ ) & (~\m3_addr_i[1]  | ~\new_[18200]_ );
  assign \new_[13075]_  = ~\new_[14677]_  & (~\new_[17329]_  | ~\new_[31718]_ );
  assign \new_[13076]_  = (~\m7_addr_i[0]  | ~\new_[18825]_ ) & (~\m0_addr_i[0]  | ~\new_[18010]_ );
  assign \new_[13077]_  = (~\m4_addr_i[0]  | ~\new_[16305]_ ) & (~\m3_addr_i[0]  | ~\new_[18200]_ );
  assign \new_[13078]_  = (~\m7_sel_i[3]  | ~\new_[18825]_ ) & (~\m0_sel_i[3]  | ~\new_[18010]_ );
  assign \new_[13079]_  = (~\m4_sel_i[3]  | ~\new_[16305]_ ) & (~\m3_sel_i[3]  | ~\new_[18200]_ );
  assign \new_[13080]_  = (~\m7_sel_i[2]  | ~\new_[18825]_ ) & (~\m0_sel_i[2]  | ~\new_[18010]_ );
  assign \new_[13081]_  = (~\new_[17193]_  | ~\m2_addr_i[25] ) & (~\new_[18193]_  | ~\m1_addr_i[25] );
  assign \new_[13082]_  = (~\m4_sel_i[2]  | ~\new_[16305]_ ) & (~\m3_sel_i[2]  | ~\new_[18200]_ );
  assign \new_[13083]_  = (~\m7_sel_i[1]  | ~\new_[18825]_ ) & (~\m0_sel_i[1]  | ~\new_[18010]_ );
  assign \new_[13084]_  = (~\m4_sel_i[1]  | ~\new_[16305]_ ) & (~\m3_sel_i[1]  | ~\new_[18200]_ );
  assign \new_[13085]_  = (~\m7_sel_i[0]  | ~\new_[18825]_ ) & (~\m0_sel_i[0]  | ~\new_[18011]_ );
  assign \new_[13086]_  = (~\m4_sel_i[0]  | ~\new_[16305]_ ) & (~\m3_sel_i[0]  | ~\new_[18200]_ );
  assign \new_[13087]_  = ~\new_[14685]_  & (~\new_[17347]_  | ~\new_[31597]_ );
  assign \new_[13088]_  = (~m7_we_i | ~\new_[18824]_ ) & (~m0_we_i | ~\new_[18011]_ );
  assign \new_[13089]_  = (~m2_we_i | ~\new_[17216]_ ) & (~m1_we_i | ~\new_[18888]_ );
  assign \new_[13090]_  = (~m4_we_i | ~\new_[18877]_ ) & (~m3_we_i | ~\new_[18200]_ );
  assign \new_[13091]_  = ~\new_[29125]_  & (~\new_[23676]_  | ~\new_[16330]_ );
  assign \new_[13092]_  = (~\m7_data_i[31]  | ~\new_[18115]_ ) & (~\m0_data_i[31]  | ~\new_[18932]_ );
  assign \new_[13093]_  = (~\m7_data_i[30]  | ~\new_[18115]_ ) & (~\m0_data_i[30]  | ~\new_[18932]_ );
  assign \new_[13094]_  = (~\m7_data_i[29]  | ~\new_[18115]_ ) & (~\m0_data_i[29]  | ~\new_[18932]_ );
  assign \new_[13095]_  = ~\new_[14691]_  & (~\new_[17335]_  | ~\new_[31575]_ );
  assign \new_[13096]_  = (~\m7_data_i[28]  | ~\new_[18115]_ ) & (~\m0_data_i[28]  | ~\new_[18932]_ );
  assign \new_[13097]_  = (~\m7_data_i[27]  | ~\new_[18116]_ ) & (~\m0_data_i[27]  | ~\new_[19637]_ );
  assign \new_[13098]_  = (~\m4_data_i[27]  | ~\new_[17260]_ ) & (~\m3_data_i[27]  | ~\new_[18175]_ );
  assign \new_[13099]_  = (~\m7_data_i[26]  | ~\new_[18115]_ ) & (~\m0_data_i[26]  | ~\new_[18932]_ );
  assign \new_[13100]_  = (~\m7_data_i[24]  | ~\new_[18115]_ ) & (~\m0_data_i[24]  | ~\new_[18932]_ );
  assign \new_[13101]_  = (~\m5_sel_i[1]  | ~\new_[18014]_ ) & (~\m6_sel_i[1]  | ~\new_[17229]_ );
  assign \new_[13102]_  = (~\m7_data_i[23]  | ~\new_[18115]_ ) & (~\m0_data_i[23]  | ~\new_[18932]_ );
  assign \new_[13103]_  = (~\m7_data_i[22]  | ~\new_[18115]_ ) & (~\m0_data_i[22]  | ~\new_[18932]_ );
  assign \new_[13104]_  = (~\m5_data_i[22]  | ~\new_[17187]_ ) & (~\m6_data_i[22]  | ~\new_[19563]_ );
  assign \new_[13105]_  = (~\m4_data_i[21]  | ~\new_[17260]_ ) & (~\m3_data_i[21]  | ~\new_[18175]_ );
  assign \new_[13106]_  = (~\m5_data_i[21]  | ~\new_[17187]_ ) & (~\m6_data_i[21]  | ~\new_[18049]_ );
  assign \new_[13107]_  = (~\m5_data_i[20]  | ~\new_[17187]_ ) & (~\m6_data_i[20]  | ~\new_[18051]_ );
  assign \new_[13108]_  = (~\m4_data_i[19]  | ~\new_[17260]_ ) & (~\m3_data_i[19]  | ~\new_[18175]_ );
  assign \new_[13109]_  = (~\m7_data_i[18]  | ~\new_[18116]_ ) & (~\m0_data_i[18]  | ~\new_[18932]_ );
  assign \new_[13110]_  = (~\m4_data_i[18]  | ~\new_[17260]_ ) & (~\m3_data_i[18]  | ~\new_[18175]_ );
  assign \new_[13111]_  = (~\m5_data_i[18]  | ~\new_[17188]_ ) & (~\m6_data_i[18]  | ~\new_[18050]_ );
  assign \new_[13112]_  = (~\m4_sel_i[3]  | ~\new_[18149]_ ) & (~\m3_sel_i[3]  | ~\new_[18928]_ );
  assign \new_[13113]_  = ~m5_stb_i | ~\new_[26243]_  | ~\new_[18738]_ ;
  assign \new_[13114]_  = ~m2_stb_i | ~\new_[27055]_  | ~\new_[18799]_ ;
  assign \new_[13115]_  = (~\m5_data_i[17]  | ~\new_[17188]_ ) & (~\m6_data_i[17]  | ~\new_[18048]_ );
  assign \new_[13116]_  = (~\m4_data_i[16]  | ~\new_[17260]_ ) & (~\m3_data_i[16]  | ~\new_[18175]_ );
  assign \new_[13117]_  = (~\m5_data_i[16]  | ~\new_[17188]_ ) & (~\m6_data_i[16]  | ~\new_[18048]_ );
  assign \new_[13118]_  = ~m6_stb_i | ~\new_[26689]_  | ~\new_[18031]_ ;
  assign \new_[13119]_  = (~\m5_data_i[15]  | ~\new_[17189]_ ) & (~\m6_data_i[15]  | ~\new_[18051]_ );
  assign \new_[13120]_  = (~\m7_data_i[14]  | ~\new_[18116]_ ) & (~\m0_data_i[14]  | ~\new_[18932]_ );
  assign \new_[13121]_  = (~\m5_data_i[14]  | ~\new_[17189]_ ) & (~\m6_data_i[14]  | ~\new_[18051]_ );
  assign \new_[13122]_  = (~\m7_data_i[13]  | ~\new_[18116]_ ) & (~\m0_data_i[13]  | ~\new_[18932]_ );
  assign \new_[13123]_  = (~\m5_data_i[13]  | ~\new_[17189]_ ) & (~\m6_data_i[13]  | ~\new_[18051]_ );
  assign \new_[13124]_  = (~\m7_data_i[12]  | ~\new_[18116]_ ) & (~\m0_data_i[12]  | ~\new_[18932]_ );
  assign \new_[13125]_  = (~\m5_data_i[12]  | ~\new_[17189]_ ) & (~\m6_data_i[12]  | ~\new_[18051]_ );
  assign \new_[13126]_  = (~\m4_data_i[11]  | ~\new_[17260]_ ) & (~\m3_data_i[11]  | ~\new_[18175]_ );
  assign \new_[13127]_  = (~\m5_data_i[11]  | ~\new_[17189]_ ) & (~\m6_data_i[11]  | ~\new_[18051]_ );
  assign \new_[13128]_  = (~\m7_data_i[10]  | ~\new_[18116]_ ) & (~\m0_data_i[10]  | ~\new_[18932]_ );
  assign \new_[13129]_  = (~\m4_addr_i[13]  | ~\new_[18149]_ ) & (~\m3_addr_i[13]  | ~\new_[18928]_ );
  assign \new_[13130]_  = (~\m5_data_i[10]  | ~\new_[18735]_ ) & (~\m6_data_i[10]  | ~\new_[18051]_ );
  assign \new_[13131]_  = (~\m7_data_i[9]  | ~\new_[18116]_ ) & (~\m0_data_i[9]  | ~\new_[18932]_ );
  assign \new_[13132]_  = (~\m5_data_i[9]  | ~\new_[17189]_ ) & (~\m6_data_i[9]  | ~\new_[18051]_ );
  assign \new_[13133]_  = (~\m4_addr_i[7]  | ~\new_[17260]_ ) & (~\m3_addr_i[7]  | ~\new_[18175]_ );
  assign \new_[13134]_  = (~\m5_data_i[8]  | ~\new_[18735]_ ) & (~\m6_data_i[8]  | ~\new_[18051]_ );
  assign \new_[13135]_  = (~\m5_data_i[7]  | ~\new_[17189]_ ) & (~\m6_data_i[7]  | ~\new_[18051]_ );
  assign \new_[13136]_  = ~\new_[16980]_  & (~\new_[17348]_  | ~\new_[31804]_ );
  assign \new_[13137]_  = (~\m5_data_i[6]  | ~\new_[18735]_ ) & (~\m6_data_i[6]  | ~\new_[18051]_ );
  assign \new_[13138]_  = (~\m5_data_i[5]  | ~\new_[17189]_ ) & (~\m6_data_i[5]  | ~\new_[18051]_ );
  assign \new_[13139]_  = (~\m7_data_i[4]  | ~\new_[18116]_ ) & (~\m0_data_i[4]  | ~\new_[18932]_ );
  assign \new_[13140]_  = (~\m5_data_i[4]  | ~\new_[17189]_ ) & (~\m6_data_i[4]  | ~\new_[18050]_ );
  assign \new_[13141]_  = (~\m5_data_i[3]  | ~\new_[17189]_ ) & (~\m6_data_i[3]  | ~\new_[18051]_ );
  assign \new_[13142]_  = (~\new_[17227]_  | ~\m6_addr_i[30] ) & (~\new_[17202]_  | ~\new_[31147]_ );
  assign \new_[13143]_  = (~\m7_data_i[2]  | ~\new_[18116]_ ) & (~\m0_data_i[2]  | ~\new_[18932]_ );
  assign \new_[13144]_  = (~\m5_data_i[2]  | ~\new_[18735]_ ) & (~\m6_data_i[2]  | ~\new_[18050]_ );
  assign \new_[13145]_  = (~\m7_data_i[1]  | ~\new_[18116]_ ) & (~\m0_data_i[1]  | ~\new_[18932]_ );
  assign \new_[13146]_  = (~\m5_data_i[1]  | ~\new_[17189]_ ) & (~\m6_data_i[1]  | ~\new_[18050]_ );
  assign \new_[13147]_  = (~\m5_data_i[0]  | ~\new_[17189]_ ) & (~\m6_data_i[0]  | ~\new_[18051]_ );
  assign \new_[13148]_  = (~\new_[18116]_  | ~\m7_addr_i[31] ) & (~\new_[18932]_  | ~\m0_addr_i[31] );
  assign \new_[13149]_  = (~\m5_addr_i[1]  | ~\new_[17188]_ ) & (~\m6_addr_i[1]  | ~\new_[18051]_ );
  assign \new_[13150]_  = (~\new_[19563]_  | ~\m6_addr_i[31] ) & (~\new_[18735]_  | ~\new_[31001]_ );
  assign \new_[13151]_  = (~\new_[18116]_  | ~\new_[31885]_ ) & (~\new_[18932]_  | ~\new_[31292]_ );
  assign \new_[13152]_  = (~\new_[19563]_  | ~\m6_addr_i[30] ) & (~\new_[18735]_  | ~\new_[31147]_ );
  assign \new_[13153]_  = (~\new_[18116]_  | ~\new_[31531]_ ) & (~\new_[18932]_  | ~\new_[31481]_ );
  assign \new_[13154]_  = ~\new_[28992]_  & (~\new_[20745]_  | ~\new_[17290]_ );
  assign \new_[13155]_  = (~\new_[19563]_  | ~\m6_addr_i[29] ) & (~\new_[18735]_  | ~\new_[31407]_ );
  assign \new_[13156]_  = (~\new_[18116]_  | ~\new_[30577]_ ) & (~\new_[18932]_  | ~\new_[30957]_ );
  assign \new_[13157]_  = ~\new_[29541]_  & (~\new_[20763]_  | ~\new_[17297]_ );
  assign \new_[13158]_  = (~\new_[19563]_  | ~\m6_addr_i[28] ) & (~\new_[18735]_  | ~\new_[31276]_ );
  assign \new_[13159]_  = (~\new_[18116]_  | ~\m7_addr_i[25] ) & (~\new_[18932]_  | ~\m0_addr_i[25] );
  assign \new_[13160]_  = (~\new_[18116]_  | ~\m7_addr_i[27] ) & (~\new_[18932]_  | ~\m0_addr_i[27] );
  assign \new_[13161]_  = ~\new_[29217]_  & (~\new_[20780]_  | ~\new_[17303]_ );
  assign \new_[13162]_  = (~\new_[19563]_  | ~\m6_addr_i[27] ) & (~\new_[18735]_  | ~\m5_addr_i[27] );
  assign \new_[13163]_  = (~\new_[18149]_  | ~\m4_addr_i[28] ) & (~\new_[18929]_  | ~\m3_addr_i[28] );
  assign \new_[13164]_  = (~\new_[18116]_  | ~\m7_addr_i[26] ) & (~\new_[18932]_  | ~\m0_addr_i[26] );
  assign \new_[13165]_  = ~\new_[29058]_  & (~\new_[20837]_  | ~\new_[17307]_ );
  assign \new_[13166]_  = (~\new_[19563]_  | ~\m6_addr_i[25] ) & (~\new_[18735]_  | ~\m5_addr_i[25] );
  assign \new_[13167]_  = (~\new_[18116]_  | ~\m7_addr_i[24] ) & (~\new_[18932]_  | ~\m0_addr_i[24] );
  assign \new_[13168]_  = (~\m4_addr_i[23]  | ~\new_[17260]_ ) & (~\m3_addr_i[23]  | ~\new_[18175]_ );
  assign \new_[13169]_  = (~\m5_addr_i[23]  | ~\new_[17188]_ ) & (~\m6_addr_i[23]  | ~\new_[18049]_ );
  assign \new_[13170]_  = ~\new_[29254]_  & (~\new_[20739]_  | ~\new_[17325]_ );
  assign \new_[13171]_  = (~\m5_addr_i[22]  | ~\new_[17188]_ ) & (~\m6_addr_i[22]  | ~\new_[19563]_ );
  assign \new_[13172]_  = (~\m4_addr_i[21]  | ~\new_[17260]_ ) & (~\m3_addr_i[21]  | ~\new_[18175]_ );
  assign \new_[13173]_  = ~\new_[20306]_  & (~\new_[17208]_  | ~\new_[30057]_ );
  assign \new_[13174]_  = ~\new_[29115]_  & (~\new_[20798]_  | ~\new_[17330]_ );
  assign \new_[13175]_  = ~\new_[29101]_  & (~\new_[20869]_  | ~\new_[17332]_ );
  assign \new_[13176]_  = (~\m4_addr_i[19]  | ~\new_[17260]_ ) & (~\m3_addr_i[19]  | ~\new_[18175]_ );
  assign \new_[13177]_  = (~\m5_addr_i[19]  | ~\new_[17187]_ ) & (~\m6_addr_i[19]  | ~\new_[18050]_ );
  assign \new_[13178]_  = ~\new_[29229]_  & (~\new_[20929]_  | ~\new_[17338]_ );
  assign \new_[13179]_  = (~\m4_addr_i[18]  | ~\new_[17260]_ ) & (~\m3_addr_i[18]  | ~\new_[18175]_ );
  assign \new_[13180]_  = (~\m5_addr_i[18]  | ~\new_[17188]_ ) & (~\m6_addr_i[18]  | ~\new_[18050]_ );
  assign \new_[13181]_  = (~\m4_addr_i[17]  | ~\new_[17260]_ ) & (~\m3_addr_i[17]  | ~\new_[18175]_ );
  assign \new_[13182]_  = (~\m5_addr_i[17]  | ~\new_[17188]_ ) & (~\m6_addr_i[17]  | ~\new_[18050]_ );
  assign \new_[13183]_  = (~\m4_addr_i[16]  | ~\new_[17260]_ ) & (~\m3_addr_i[16]  | ~\new_[18175]_ );
  assign \new_[13184]_  = ~\new_[29167]_  & (~\new_[20980]_  | ~\new_[17337]_ );
  assign \new_[13185]_  = (~\m2_addr_i[18]  | ~\new_[18069]_ ) & (~\m1_addr_i[18]  | ~\new_[19625]_ );
  assign \new_[13186]_  = (~\m5_addr_i[14]  | ~\new_[17187]_ ) & (~\m6_addr_i[14]  | ~\new_[18049]_ );
  assign \new_[13187]_  = (~\m4_addr_i[13]  | ~\new_[17260]_ ) & (~\m3_addr_i[13]  | ~\new_[18175]_ );
  assign \new_[13188]_  = (~\m5_addr_i[13]  | ~\new_[17187]_ ) & (~\m6_addr_i[13]  | ~\new_[18050]_ );
  assign \new_[13189]_  = ~\new_[20296]_  & (~\new_[17242]_  | ~\new_[28872]_ );
  assign \new_[13190]_  = \new_[6035]_  ? \new_[29029]_  : \new_[17289]_ ;
  assign \new_[13191]_  = (~\m4_addr_i[12]  | ~\new_[17260]_ ) & (~\m3_addr_i[12]  | ~\new_[18175]_ );
  assign \new_[13192]_  = (~\m5_addr_i[12]  | ~\new_[17187]_ ) & (~\m6_addr_i[12]  | ~\new_[18050]_ );
  assign \new_[13193]_  = \new_[6039]_  ? \new_[29291]_  : \new_[17292]_ ;
  assign \new_[13194]_  = (~\m4_addr_i[11]  | ~\new_[17260]_ ) & (~\m3_addr_i[11]  | ~\new_[18175]_ );
  assign \new_[13195]_  = \new_[6044]_  ? \new_[28934]_  : \new_[17299]_ ;
  assign \new_[13196]_  = (~\m4_addr_i[10]  | ~\new_[17260]_ ) & (~\m3_addr_i[10]  | ~\new_[18175]_ );
  assign \new_[13197]_  = \new_[17291]_  ? \new_[30785]_  : \new_[6199]_ ;
  assign \new_[13198]_  = \new_[6047]_  ? \new_[29381]_  : \new_[17305]_ ;
  assign \new_[13199]_  = (~\m4_addr_i[9]  | ~\new_[17260]_ ) & (~\m3_addr_i[9]  | ~\new_[18175]_ );
  assign \new_[13200]_  = (~\m5_addr_i[9]  | ~\new_[17188]_ ) & (~\m6_addr_i[9]  | ~\new_[18049]_ );
  assign \new_[13201]_  = \new_[5973]_  ? \new_[28993]_  : \new_[17314]_ ;
  assign \new_[13202]_  = (~\m5_addr_i[8]  | ~\new_[17188]_ ) & (~\m6_addr_i[8]  | ~\new_[18049]_ );
  assign \new_[13203]_  = \new_[6058]_  ? \new_[28110]_  : \new_[17318]_ ;
  assign \new_[13204]_  = (~\m4_addr_i[1]  | ~\new_[17260]_ ) & (~\m3_addr_i[1]  | ~\new_[18175]_ );
  assign \new_[13205]_  = ~\new_[16293]_  & ~\new_[31619]_ ;
  assign \new_[13206]_  = ~\new_[31990]_  & ~\new_[31667]_ ;
  assign \new_[13207]_  = ~\new_[31688]_  & ~\new_[16321]_ ;
  assign \new_[13208]_  = ~\new_[16304]_  & ~\new_[31739]_ ;
  assign \new_[13209]_  = ~\new_[16304]_  & ~\new_[31790]_ ;
  assign \new_[13210]_  = ~\new_[31907]_  & ~\new_[16303]_ ;
  assign \new_[13211]_  = (~\m4_addr_i[21]  | ~\new_[18156]_ ) & (~\m3_addr_i[21]  | ~\new_[18130]_ );
  assign \new_[13212]_  = ~\new_[31750]_  & ~\new_[16321]_ ;
  assign \new_[13213]_  = ~\new_[16304]_  & ~\new_[31913]_ ;
  assign \new_[13214]_  = ~\new_[16326]_  & ~\new_[31745]_ ;
  assign \new_[13215]_  = ~\new_[16326]_  & ~\new_[31644]_ ;
  assign \new_[13216]_  = ~\new_[31609]_  & ~\new_[16321]_ ;
  assign \new_[13217]_  = ~\new_[16326]_  & ~\new_[31612]_ ;
  assign \new_[13218]_  = (~\m2_data_i[4]  | ~\new_[18068]_ ) & (~\m1_data_i[4]  | ~\new_[20573]_ );
  assign \new_[13219]_  = (~\m4_data_i[31]  | ~\new_[19608]_ ) & (~\m3_data_i[31]  | ~\new_[18002]_ );
  assign \new_[13220]_  = (~\m4_data_i[30]  | ~\new_[17261]_ ) & (~\m3_data_i[30]  | ~\new_[18002]_ );
  assign \new_[13221]_  = (~\m5_data_i[30]  | ~\new_[18871]_ ) & (~\m6_data_i[30]  | ~\new_[20552]_ );
  assign \new_[13222]_  = (~\m4_data_i[29]  | ~\new_[17261]_ ) & (~\m3_data_i[29]  | ~\new_[18002]_ );
  assign \new_[13223]_  = (~\m4_data_i[28]  | ~\new_[17261]_ ) & (~\m3_data_i[28]  | ~\new_[18002]_ );
  assign \new_[13224]_  = (~\m4_data_i[27]  | ~\new_[17261]_ ) & (~\m3_data_i[27]  | ~\new_[18002]_ );
  assign \new_[13225]_  = (~\m4_data_i[26]  | ~\new_[17261]_ ) & (~\m3_data_i[26]  | ~\new_[18002]_ );
  assign \new_[13226]_  = ~m6_stb_i | ~\new_[17213]_  | ~\new_[29149]_ ;
  assign \new_[13227]_  = ~m2_stb_i | ~\new_[18078]_  | ~\new_[29963]_ ;
  assign \new_[13228]_  = (~\m4_data_i[25]  | ~\new_[17261]_ ) & (~\m3_data_i[25]  | ~\new_[18002]_ );
  assign \new_[13229]_  = (~\m4_data_i[24]  | ~\new_[17261]_ ) & (~\m3_data_i[24]  | ~\new_[18002]_ );
  assign \new_[13230]_  = (~\m4_data_i[23]  | ~\new_[19608]_ ) & (~\m3_data_i[23]  | ~\new_[19539]_ );
  assign \new_[13231]_  = (~\m5_data_i[23]  | ~\new_[18871]_ ) & (~\m6_data_i[23]  | ~\new_[18794]_ );
  assign \new_[13232]_  = (~\m7_data_i[23]  | ~\new_[18835]_ ) & (~\m0_data_i[23]  | ~\new_[19642]_ );
  assign \new_[13233]_  = (~\m4_data_i[22]  | ~\new_[17261]_ ) & (~\m3_data_i[22]  | ~\new_[18002]_ );
  assign \new_[13234]_  = (~\m4_data_i[21]  | ~\new_[17261]_ ) & (~\m3_data_i[21]  | ~\new_[18002]_ );
  assign \new_[13235]_  = (~\m5_data_i[21]  | ~\new_[18871]_ ) & (~\m6_data_i[21]  | ~\new_[18794]_ );
  assign \new_[13236]_  = ~\new_[27983]_  & ~\new_[16293]_ ;
  assign \new_[13237]_  = (~\m4_data_i[20]  | ~\new_[17261]_ ) & (~\m3_data_i[20]  | ~\new_[19539]_ );
  assign \new_[13238]_  = (~\m5_data_i[20]  | ~\new_[18871]_ ) & (~\m6_data_i[20]  | ~\new_[18052]_ );
  assign \new_[13239]_  = (~\m4_data_i[19]  | ~\new_[17261]_ ) & (~\m3_data_i[19]  | ~\new_[18002]_ );
  assign \new_[13240]_  = (~\m4_data_i[18]  | ~\new_[17261]_ ) & (~\m3_data_i[18]  | ~\new_[18002]_ );
  assign \new_[13241]_  = (~\m5_data_i[18]  | ~\new_[18871]_ ) & (~\m6_data_i[18]  | ~\new_[20552]_ );
  assign \new_[13242]_  = (~\m2_addr_i[21]  | ~\new_[18067]_ ) & (~\m1_addr_i[21]  | ~\new_[19625]_ );
  assign \new_[13243]_  = (~\m4_data_i[17]  | ~\new_[17261]_ ) & (~\m3_data_i[17]  | ~\new_[18002]_ );
  assign \new_[13244]_  = (~\m4_data_i[16]  | ~\new_[17261]_ ) & (~\m3_data_i[16]  | ~\new_[18002]_ );
  assign \new_[13245]_  = ~\new_[28927]_  & ~\new_[16293]_ ;
  assign \new_[13246]_  = (~\m4_data_i[15]  | ~\new_[17261]_ ) & (~\m3_data_i[15]  | ~\new_[18002]_ );
  assign \new_[13247]_  = ~s1_ack_i | ~\new_[18030]_  | ~\new_[30108]_ ;
  assign \new_[13248]_  = (~\m4_data_i[14]  | ~\new_[17261]_ ) & (~\m3_data_i[14]  | ~\new_[18002]_ );
  assign \new_[13249]_  = ~s14_ack_i | ~\new_[18032]_  | ~\new_[29631]_ ;
  assign \new_[13250]_  = ~s8_ack_i | ~\new_[16287]_  | ~\new_[29420]_ ;
  assign \new_[13251]_  = (~\m4_data_i[13]  | ~\new_[17261]_ ) & (~\m3_data_i[13]  | ~\new_[18002]_ );
  assign \new_[13252]_  = ~s14_err_i | ~\new_[16286]_  | ~\new_[29631]_ ;
  assign \new_[13253]_  = (~\m4_data_i[12]  | ~\new_[17261]_ ) & (~\m3_data_i[12]  | ~\new_[18002]_ );
  assign \new_[13254]_  = ~s1_err_i | ~\new_[18030]_  | ~\new_[30108]_ ;
  assign \new_[13255]_  = (~\m4_data_i[11]  | ~\new_[19608]_ ) & (~\m3_data_i[11]  | ~\new_[18002]_ );
  assign \new_[13256]_  = ~s14_rty_i | ~\new_[18032]_  | ~\new_[29631]_ ;
  assign \new_[13257]_  = ~s8_rty_i | ~\new_[16287]_  | ~\new_[29420]_ ;
  assign \new_[13258]_  = ~s11_rty_i | ~\new_[17229]_  | ~\new_[30284]_ ;
  assign \new_[13259]_  = (~\m4_data_i[10]  | ~\new_[17261]_ ) & (~\m3_data_i[10]  | ~\new_[18002]_ );
  assign \new_[13260]_  = ~s1_rty_i | ~\new_[18030]_  | ~\new_[30108]_ ;
  assign \new_[13261]_  = ~s14_ack_i | ~\new_[16290]_  | ~\new_[29807]_ ;
  assign \new_[13262]_  = (~\m4_data_i[9]  | ~\new_[17261]_ ) & (~\m3_data_i[9]  | ~\new_[18002]_ );
  assign \new_[13263]_  = (~\m4_data_i[8]  | ~\new_[17261]_ ) & (~\m3_data_i[8]  | ~\new_[18002]_ );
  assign \new_[13264]_  = (~\m4_data_i[7]  | ~\new_[17261]_ ) & (~\m3_data_i[7]  | ~\new_[18002]_ );
  assign \new_[13265]_  = ~s14_err_i | ~\new_[16290]_  | ~\new_[29807]_ ;
  assign \new_[13266]_  = (~\m4_data_i[6]  | ~\new_[19608]_ ) & (~\m3_data_i[6]  | ~\new_[18002]_ );
  assign \new_[13267]_  = ~s2_rty_i | ~\new_[17216]_  | ~\new_[29788]_ ;
  assign \new_[13268]_  = (~\m4_data_i[5]  | ~\new_[17261]_ ) & (~\m3_data_i[5]  | ~\new_[18002]_ );
  assign \new_[13269]_  = (~\m7_data_i[4]  | ~\new_[18835]_ ) & (~\m0_data_i[4]  | ~\new_[18937]_ );
  assign \new_[13270]_  = (~\m4_data_i[4]  | ~\new_[19608]_ ) & (~\m3_data_i[4]  | ~\new_[19539]_ );
  assign \new_[13271]_  = ~s14_rty_i | ~\new_[16290]_  | ~\new_[29807]_ ;
  assign \new_[13272]_  = ~m6_stb_i | ~\new_[16289]_  | ~\new_[29823]_ ;
  assign \new_[13273]_  = (~\m7_data_i[3]  | ~\new_[18835]_ ) & (~\m0_data_i[3]  | ~\new_[18937]_ );
  assign \new_[13274]_  = (~\m4_data_i[3]  | ~\new_[17261]_ ) & (~\m3_data_i[3]  | ~\new_[18002]_ );
  assign \new_[13275]_  = ~\new_[27213]_  & ~\new_[31990]_ ;
  assign \new_[13276]_  = (~\m4_data_i[2]  | ~\new_[17261]_ ) & (~\m3_data_i[2]  | ~\new_[19539]_ );
  assign \new_[13277]_  = (~\m7_data_i[2]  | ~\new_[18835]_ ) & (~\m0_data_i[2]  | ~\new_[19642]_ );
  assign \new_[13278]_  = (~\m4_data_i[1]  | ~\new_[17261]_ ) & (~\m3_data_i[1]  | ~\new_[18734]_ );
  assign \new_[13279]_  = (~\m7_data_i[1]  | ~\new_[18835]_ ) & (~\m0_data_i[1]  | ~\new_[18937]_ );
  assign \new_[13280]_  = (~\m4_data_i[0]  | ~\new_[17261]_ ) & (~\m3_data_i[0]  | ~\new_[19539]_ );
  assign \new_[13281]_  = (~\m7_data_i[0]  | ~\new_[18835]_ ) & (~\m0_data_i[0]  | ~\new_[19642]_ );
  assign \new_[13282]_  = ~m4_stb_i | ~\new_[18878]_  | ~\new_[29627]_ ;
  assign \new_[13283]_  = \new_[16325]_  & \new_[31935]_ ;
  assign \new_[13284]_  = (~\new_[18795]_  | ~\m6_addr_i[31] ) & (~\new_[18871]_  | ~\new_[31001]_ );
  assign \new_[13285]_  = (~\new_[17261]_  | ~\m4_addr_i[31] ) & (~\new_[18002]_  | ~\m3_addr_i[31] );
  assign \new_[13286]_  = (~\new_[17261]_  | ~\m4_addr_i[30] ) & (~\new_[18734]_  | ~\m3_addr_i[30] );
  assign \new_[13287]_  = (~\new_[18795]_  | ~\m6_addr_i[30] ) & (~\new_[18871]_  | ~\new_[31147]_ );
  assign \new_[13288]_  = (~\new_[17261]_  | ~\m4_addr_i[29] ) & (~\new_[19539]_  | ~\m3_addr_i[29] );
  assign \new_[13289]_  = (~\new_[18835]_  | ~\new_[31531]_ ) & (~\new_[18937]_  | ~\new_[31481]_ );
  assign \new_[13290]_  = (~\new_[18795]_  | ~\m6_addr_i[29] ) & (~\new_[18871]_  | ~\new_[31407]_ );
  assign \new_[13291]_  = (~\new_[18795]_  | ~\m6_addr_i[28] ) & (~\new_[18871]_  | ~\new_[31276]_ );
  assign \new_[13292]_  = (~\new_[19608]_  | ~\m4_addr_i[28] ) & (~\new_[18002]_  | ~\m3_addr_i[28] );
  assign \new_[13293]_  = ~\new_[30683]_  & ~\new_[16274]_ ;
  assign \new_[13294]_  = (~\new_[18795]_  | ~\m6_addr_i[27] ) & (~\new_[18871]_  | ~\m5_addr_i[27] );
  assign \new_[13295]_  = (~\new_[19608]_  | ~\m4_addr_i[27] ) & (~\new_[18002]_  | ~\m3_addr_i[27] );
  assign \new_[13296]_  = (~\new_[17261]_  | ~\m4_addr_i[26] ) & (~\new_[18734]_  | ~\m3_addr_i[26] );
  assign \new_[13297]_  = (~\new_[18795]_  | ~\m6_addr_i[26] ) & (~\new_[18871]_  | ~\m5_addr_i[26] );
  assign \new_[13298]_  = (~\m2_data_i[30]  | ~\new_[18799]_ ) & (~\m1_data_i[30]  | ~\new_[18887]_ );
  assign \new_[13299]_  = (~\new_[17261]_  | ~\m4_addr_i[25] ) & (~\new_[18734]_  | ~\m3_addr_i[25] );
  assign \new_[13300]_  = (~\new_[18794]_  | ~\m6_addr_i[25] ) & (~\new_[18871]_  | ~\m5_addr_i[25] );
  assign \new_[13301]_  = (~\new_[18795]_  | ~\m6_addr_i[24] ) & (~\new_[18871]_  | ~\m5_addr_i[24] );
  assign \new_[13302]_  = (~\new_[19608]_  | ~\m4_addr_i[24] ) & (~\new_[18002]_  | ~\m3_addr_i[24] );
  assign \new_[13303]_  = (~\m4_addr_i[23]  | ~\new_[17261]_ ) & (~\m3_addr_i[23]  | ~\new_[18002]_ );
  assign \new_[13304]_  = (~\m4_addr_i[22]  | ~\new_[17261]_ ) & (~\m3_addr_i[22]  | ~\new_[18734]_ );
  assign \new_[13305]_  = (~\m4_addr_i[21]  | ~\new_[17261]_ ) & (~\m3_addr_i[21]  | ~\new_[18002]_ );
  assign \new_[13306]_  = ~m2_stb_i | ~\new_[17219]_  | ~\new_[32056]_ ;
  assign \new_[13307]_  = ~m6_stb_i | ~\new_[18032]_  | ~\new_[29631]_ ;
  assign \new_[13308]_  = ~m2_stb_i | ~\new_[18068]_  | ~\new_[30626]_ ;
  assign \new_[13309]_  = (~\m4_addr_i[20]  | ~\new_[17261]_ ) & (~\m3_addr_i[20]  | ~\new_[18002]_ );
  assign \new_[13310]_  = (~\m5_addr_i[20]  | ~\new_[18871]_ ) & (~\m6_addr_i[20]  | ~\new_[18794]_ );
  assign \new_[13311]_  = ~s2_ack_i | ~\new_[18877]_  | ~\new_[30088]_ ;
  assign \new_[13312]_  = (~\m4_addr_i[19]  | ~\new_[17261]_ ) & (~\m3_addr_i[19]  | ~\new_[18002]_ );
  assign \new_[13313]_  = ~s9_ack_i | ~\new_[16308]_  | ~\new_[29185]_ ;
  assign \new_[13314]_  = (~\m5_addr_i[19]  | ~\new_[18871]_ ) & (~\m6_addr_i[19]  | ~\new_[18794]_ );
  assign \new_[13315]_  = ~s14_ack_i | ~\new_[17272]_  | ~\new_[29641]_ ;
  assign \new_[13316]_  = ~s2_err_i | ~\new_[18877]_  | ~\new_[30088]_ ;
  assign \new_[13317]_  = ~s8_err_i | ~\new_[18878]_  | ~\new_[29627]_ ;
  assign \new_[13318]_  = (~\m4_addr_i[18]  | ~\new_[17261]_ ) & (~\m3_addr_i[18]  | ~\new_[18002]_ );
  assign \new_[13319]_  = (~\m4_addr_i[17]  | ~\new_[19608]_ ) & (~\m3_addr_i[17]  | ~\new_[19539]_ );
  assign \new_[13320]_  = ~s2_rty_i | ~\new_[18877]_  | ~\new_[30088]_ ;
  assign \new_[13321]_  = ~m2_stb_i | ~\new_[17216]_  | ~\new_[29788]_ ;
  assign \new_[13322]_  = (~\m5_addr_i[17]  | ~\new_[18871]_ ) & (~\m6_addr_i[17]  | ~\new_[18794]_ );
  assign \new_[13323]_  = ~m4_stb_i | ~\new_[18877]_  | ~\new_[30088]_ ;
  assign \new_[13324]_  = ~s9_rty_i | ~\new_[16308]_  | ~\new_[29185]_ ;
  assign \new_[13325]_  = (~\m4_addr_i[16]  | ~\new_[17261]_ ) & (~\m3_addr_i[16]  | ~\new_[18002]_ );
  assign \new_[13326]_  = (~\m5_addr_i[16]  | ~\new_[18871]_ ) & (~\m6_addr_i[16]  | ~\new_[18794]_ );
  assign \new_[13327]_  = (~\m5_addr_i[15]  | ~\new_[18871]_ ) & (~\m6_addr_i[15]  | ~\new_[18795]_ );
  assign \new_[13328]_  = (~\m4_addr_i[15]  | ~\new_[17261]_ ) & (~\m3_addr_i[15]  | ~\new_[18002]_ );
  assign \new_[13329]_  = (~\m4_addr_i[14]  | ~\new_[17261]_ ) & (~\m3_addr_i[14]  | ~\new_[19539]_ );
  assign \new_[13330]_  = (~\m5_addr_i[14]  | ~\new_[18871]_ ) & (~\m6_addr_i[14]  | ~\new_[18052]_ );
  assign \new_[13331]_  = (~\m4_addr_i[13]  | ~\new_[19608]_ ) & (~\m3_addr_i[13]  | ~\new_[19539]_ );
  assign \new_[13332]_  = (~\m7_addr_i[13]  | ~\new_[18835]_ ) & (~\m0_addr_i[13]  | ~\new_[19642]_ );
  assign \new_[13333]_  = (~\m5_addr_i[13]  | ~\new_[18871]_ ) & (~\m6_addr_i[13]  | ~\new_[18795]_ );
  assign \new_[13334]_  = (~\m4_addr_i[12]  | ~\new_[19608]_ ) & (~\m3_addr_i[12]  | ~\new_[19539]_ );
  assign \new_[13335]_  = (~\m5_addr_i[12]  | ~\new_[18871]_ ) & (~\m6_addr_i[12]  | ~\new_[18794]_ );
  assign \new_[13336]_  = (~\m4_addr_i[11]  | ~\new_[17261]_ ) & (~\m3_addr_i[11]  | ~\new_[18002]_ );
  assign \new_[13337]_  = ~m4_stb_i | ~\new_[18157]_  | ~\new_[29012]_ ;
  assign \new_[13338]_  = (~\m4_addr_i[10]  | ~\new_[19608]_ ) & (~\m3_addr_i[10]  | ~\new_[18002]_ );
  assign \new_[13339]_  = (~\m4_addr_i[9]  | ~\new_[19608]_ ) & (~\m3_addr_i[9]  | ~\new_[19539]_ );
  assign \new_[13340]_  = (~\m5_addr_i[9]  | ~\new_[18871]_ ) & (~\m6_addr_i[9]  | ~\new_[18794]_ );
  assign \new_[13341]_  = (~\m7_addr_i[9]  | ~\new_[18835]_ ) & (~\m0_addr_i[9]  | ~\new_[18937]_ );
  assign \new_[13342]_  = (~\m4_addr_i[8]  | ~\new_[17261]_ ) & (~\m3_addr_i[8]  | ~\new_[18002]_ );
  assign \new_[13343]_  = (~\m4_addr_i[7]  | ~\new_[17261]_ ) & (~\m3_addr_i[7]  | ~\new_[18002]_ );
  assign \new_[13344]_  = (~\m4_addr_i[6]  | ~\new_[19608]_ ) & (~\m3_addr_i[6]  | ~\new_[19539]_ );
  assign \new_[13345]_  = ~s12_ack_i | ~\new_[18004]_  | ~\new_[29640]_ ;
  assign \new_[13346]_  = (~\m5_addr_i[6]  | ~\new_[18871]_ ) & (~\m6_addr_i[6]  | ~\new_[18795]_ );
  assign \new_[13347]_  = (~\m2_addr_i[14]  | ~\new_[18068]_ ) & (~\m1_addr_i[14]  | ~\new_[18901]_ );
  assign \new_[13348]_  = (~\m7_addr_i[6]  | ~\new_[18835]_ ) & (~\m0_addr_i[6]  | ~\new_[18937]_ );
  assign \new_[13349]_  = ~s9_ack_i | ~\new_[16277]_  | ~\new_[29951]_ ;
  assign \new_[13350]_  = ~\new_[30335]_  | ~\new_[18026]_  | ~m0_stb_i;
  assign \new_[13351]_  = (~\m4_addr_i[5]  | ~\new_[19608]_ ) & (~\m3_addr_i[5]  | ~\new_[18002]_ );
  assign \new_[13352]_  = (~\m5_addr_i[5]  | ~\new_[18871]_ ) & (~\m6_addr_i[5]  | ~\new_[18795]_ );
  assign \new_[13353]_  = ~s11_ack_i | ~\new_[18015]_  | ~\new_[30311]_ ;
  assign \new_[13354]_  = (~\m4_addr_i[4]  | ~\new_[19608]_ ) & (~\m3_addr_i[4]  | ~\new_[18002]_ );
  assign \new_[13355]_  = ~s12_err_i | ~\new_[18004]_  | ~\new_[29640]_ ;
  assign \new_[13356]_  = (~\m5_addr_i[4]  | ~\new_[18871]_ ) & (~\m6_addr_i[4]  | ~\new_[18795]_ );
  assign \new_[13357]_  = ~s9_err_i | ~\new_[18008]_  | ~\new_[29951]_ ;
  assign \new_[13358]_  = (~\m7_addr_i[4]  | ~\new_[18835]_ ) & (~\m0_addr_i[4]  | ~\new_[19642]_ );
  assign \new_[13359]_  = \new_[16300]_  | \new_[23747]_ ;
  assign \new_[13360]_  = ~s1_rty_i | ~\new_[18738]_  | ~\new_[29769]_ ;
  assign \new_[13361]_  = (~\m4_addr_i[3]  | ~\new_[19608]_ ) & (~\m3_addr_i[3]  | ~\new_[18002]_ );
  assign \new_[13362]_  = (~\m7_addr_i[3]  | ~\new_[18835]_ ) & (~\new_[31884]_  | ~\new_[18937]_ );
  assign \new_[13363]_  = \new_[16294]_  | \new_[23366]_ ;
  assign \new_[13364]_  = ~s9_rty_i | ~\new_[16277]_  | ~\new_[29951]_ ;
  assign \new_[13365]_  = (~\m4_addr_i[2]  | ~\new_[17261]_ ) & (~\m3_addr_i[2]  | ~\new_[18734]_ );
  assign \new_[13366]_  = ~s12_rty_i | ~\new_[18004]_  | ~\new_[29640]_ ;
  assign \new_[13367]_  = ~\new_[30589]_  & ~\new_[16316]_ ;
  assign \new_[13368]_  = ~\new_[29603]_  | ~\new_[16279]_  | ~s0_ack_i;
  assign \new_[13369]_  = \new_[16281]_  | \new_[23398]_ ;
  assign \new_[13370]_  = (~\m4_addr_i[1]  | ~\new_[17261]_ ) & (~\m3_addr_i[1]  | ~\new_[18002]_ );
  assign \new_[13371]_  = \new_[16282]_  | \new_[23434]_ ;
  assign \new_[13372]_  = ~\new_[29034]_  | ~\new_[18027]_  | ~s9_ack_i;
  assign \new_[13373]_  = (~\m4_addr_i[0]  | ~\new_[19608]_ ) & (~\m3_addr_i[0]  | ~\new_[18002]_ );
  assign \new_[13374]_  = \new_[16283]_  | \new_[22189]_ ;
  assign \new_[13375]_  = ~\new_[29708]_  | ~\new_[16284]_  | ~m0_stb_i;
  assign \new_[13376]_  = (~\m4_sel_i[3]  | ~\new_[17261]_ ) & (~\m3_sel_i[3]  | ~\new_[18734]_ );
  assign \new_[13377]_  = ~m3_stb_i | ~\new_[18206]_  | ~\new_[29939]_ ;
  assign \new_[13378]_  = (~\m7_sel_i[3]  | ~\new_[18835]_ ) & (~\m0_sel_i[3]  | ~\new_[18937]_ );
  assign \new_[13379]_  = \new_[16298]_  | \new_[22232]_ ;
  assign \new_[13380]_  = (~\m4_sel_i[2]  | ~\new_[19608]_ ) & (~\m3_sel_i[2]  | ~\new_[19539]_ );
  assign \new_[13381]_  = (~\m7_sel_i[2]  | ~\new_[18835]_ ) & (~\m0_sel_i[2]  | ~\new_[19642]_ );
  assign \new_[13382]_  = (~\m4_sel_i[1]  | ~\new_[17261]_ ) & (~\m3_sel_i[1]  | ~\new_[18002]_ );
  assign \new_[13383]_  = (~\m4_sel_i[0]  | ~\new_[19608]_ ) & (~\m3_sel_i[0]  | ~\new_[19539]_ );
  assign \new_[13384]_  = \new_[16311]_  | \new_[22207]_ ;
  assign \new_[13385]_  = (~\m7_sel_i[0]  | ~\new_[18835]_ ) & (~\m0_sel_i[0]  | ~\new_[19642]_ );
  assign \new_[13386]_  = ~s12_ack_i | ~\new_[16296]_  | ~\new_[27347]_ ;
  assign \new_[13387]_  = (~m4_we_i | ~\new_[19608]_ ) & (~m3_we_i | ~\new_[19539]_ );
  assign \new_[13388]_  = ~s12_err_i | ~\new_[16296]_  | ~\new_[27347]_ ;
  assign \new_[13389]_  = (~m7_we_i | ~\new_[18835]_ ) & (~m0_we_i | ~\new_[19642]_ );
  assign \new_[13390]_  = ~s14_err_i | ~\new_[16297]_  | ~\new_[30106]_ ;
  assign \new_[13391]_  = (~\m5_data_i[31]  | ~\new_[18007]_ ) & (~\m6_data_i[31]  | ~\new_[19577]_ );
  assign \new_[13392]_  = (~\m4_data_i[31]  | ~\new_[17267]_ ) & (~\m3_data_i[31]  | ~\new_[18206]_ );
  assign \new_[13393]_  = ~m7_stb_i | ~\new_[18111]_  | ~\new_[29905]_ ;
  assign \new_[13394]_  = \new_[16299]_  | \new_[23608]_ ;
  assign \new_[13395]_  = (~\m5_data_i[30]  | ~\new_[18007]_ ) & (~\m6_data_i[30]  | ~\new_[18086]_ );
  assign \new_[13396]_  = ~s3_ack_i | ~\new_[18175]_  | ~\new_[29947]_ ;
  assign \new_[13397]_  = (~\m5_data_i[28]  | ~\new_[18007]_ ) & (~\m6_data_i[28]  | ~\new_[18086]_ );
  assign \new_[13398]_  = (~\m4_data_i[28]  | ~\new_[17267]_ ) & (~\m3_data_i[28]  | ~\new_[18206]_ );
  assign \new_[13399]_  = ~s14_rty_i | ~\new_[16297]_  | ~\new_[30106]_ ;
  assign \new_[13400]_  = ~s3_rty_i | ~\new_[18175]_  | ~\new_[29947]_ ;
  assign \new_[13401]_  = ~s12_rty_i | ~\new_[16296]_  | ~\new_[27347]_ ;
  assign \new_[13402]_  = (~\m5_data_i[27]  | ~\new_[18007]_ ) & (~\m6_data_i[27]  | ~\new_[18087]_ );
  assign \new_[13403]_  = (~\m4_data_i[26]  | ~\new_[17267]_ ) & (~\m3_data_i[26]  | ~\new_[18206]_ );
  assign \new_[13404]_  = ~\new_[27760]_  & ~\new_[16316]_ ;
  assign \new_[13405]_  = (~\m5_data_i[26]  | ~\new_[18007]_ ) & (~\m6_data_i[26]  | ~\new_[18086]_ );
  assign \new_[13406]_  = ~m3_stb_i | ~\new_[18130]_  | ~\new_[29710]_ ;
  assign \new_[13407]_  = ~\new_[29476]_  & ~\new_[16303]_ ;
  assign \new_[13408]_  = ~m5_stb_i | ~\new_[17194]_  | ~\new_[32267]_ ;
  assign \new_[13409]_  = ~\new_[27565]_  & ~\new_[32345]_ ;
  assign \new_[13410]_  = ~s14_ack_i | ~\new_[16297]_  | ~\new_[30106]_ ;
  assign \new_[13411]_  = ~\new_[28874]_  & ~\new_[16304]_ ;
  assign \new_[13412]_  = (~\m5_data_i[23]  | ~\new_[18007]_ ) & (~\m6_data_i[23]  | ~\new_[19577]_ );
  assign \new_[13413]_  = ~s3_err_i | ~\new_[18175]_  | ~\new_[29947]_ ;
  assign \new_[13414]_  = (~\m2_data_i[15]  | ~\new_[18799]_ ) & (~\m1_data_i[15]  | ~\new_[20571]_ );
  assign \new_[13415]_  = (~\m5_data_i[21]  | ~\new_[18007]_ ) & (~\m6_data_i[21]  | ~\new_[18087]_ );
  assign \new_[13416]_  = (~\m5_data_i[20]  | ~\new_[18007]_ ) & (~\m6_data_i[20]  | ~\new_[18086]_ );
  assign \new_[13417]_  = \new_[16313]_  | \new_[22320]_ ;
  assign \new_[13418]_  = ~m3_stb_i | ~\new_[18175]_  | ~\new_[29947]_ ;
  assign \new_[13419]_  = (~\m4_data_i[17]  | ~\new_[17267]_ ) & (~\m3_data_i[17]  | ~\new_[18206]_ );
  assign \new_[13420]_  = (~\m5_data_i[17]  | ~\new_[18007]_ ) & (~\m6_data_i[17]  | ~\new_[18086]_ );
  assign \new_[13421]_  = (~\m4_data_i[16]  | ~\new_[18881]_ ) & (~\m3_data_i[16]  | ~\new_[18206]_ );
  assign \new_[13422]_  = (~\m2_data_i[13]  | ~\new_[17221]_ ) & (~\m1_data_i[13]  | ~\new_[17275]_ );
  assign \new_[13423]_  = (~\m5_data_i[12]  | ~\new_[18007]_ ) & (~\m6_data_i[12]  | ~\new_[19577]_ );
  assign \new_[13424]_  = ~\new_[23388]_  & (~\new_[17370]_  | ~\new_[28134]_ );
  assign \new_[13425]_  = (~\m5_data_i[11]  | ~\new_[18007]_ ) & (~\m6_data_i[11]  | ~\new_[19577]_ );
  assign \new_[13426]_  = (~\m4_data_i[10]  | ~\new_[17267]_ ) & (~\m3_data_i[10]  | ~\new_[18206]_ );
  assign \new_[13427]_  = (~\m2_data_i[10]  | ~\new_[17221]_ ) & (~\m1_data_i[10]  | ~\new_[17275]_ );
  assign \new_[13428]_  = ~\new_[22246]_  & (~\new_[17371]_  | ~\new_[24356]_ );
  assign \new_[13429]_  = (~\m5_data_i[10]  | ~\new_[18007]_ ) & (~\m6_data_i[10]  | ~\new_[19577]_ );
  assign \new_[13430]_  = (~\m5_data_i[9]  | ~\new_[18007]_ ) & (~\m6_data_i[9]  | ~\new_[18086]_ );
  assign \new_[13431]_  = (~\m4_data_i[9]  | ~\new_[17267]_ ) & (~\m3_data_i[9]  | ~\new_[18206]_ );
  assign \new_[13432]_  = (~\m5_data_i[8]  | ~\new_[18007]_ ) & (~\m6_data_i[8]  | ~\new_[18086]_ );
  assign \new_[13433]_  = (~\m4_data_i[8]  | ~\new_[17267]_ ) & (~\m3_data_i[8]  | ~\new_[18206]_ );
  assign \new_[13434]_  = ~\new_[25123]_  & (~\new_[17372]_  | ~\new_[23096]_ );
  assign \new_[13435]_  = (~\m4_data_i[6]  | ~\new_[17267]_ ) & (~\m3_data_i[6]  | ~\new_[18206]_ );
  assign \new_[13436]_  = (~\m2_data_i[6]  | ~\new_[17221]_ ) & (~\m1_data_i[6]  | ~\new_[17275]_ );
  assign \new_[13437]_  = (~\m4_addr_i[21]  | ~\new_[18149]_ ) & (~\m3_addr_i[21]  | ~\new_[18930]_ );
  assign \new_[13438]_  = (~\m5_data_i[5]  | ~\new_[18007]_ ) & (~\m6_data_i[5]  | ~\new_[18086]_ );
  assign \new_[13439]_  = (~\m4_data_i[5]  | ~\new_[17267]_ ) & (~\m3_data_i[5]  | ~\new_[18206]_ );
  assign \new_[13440]_  = (~\m4_data_i[4]  | ~\new_[17267]_ ) & (~\m3_data_i[4]  | ~\new_[18206]_ );
  assign \new_[13441]_  = (~\new_[19563]_  | ~\m6_addr_i[26] ) & (~\new_[18735]_  | ~\m5_addr_i[26] );
  assign \new_[13442]_  = (~\m4_data_i[3]  | ~\new_[17267]_ ) & (~\m3_data_i[3]  | ~\new_[18206]_ );
  assign \new_[13443]_  = (~\m5_data_i[3]  | ~\new_[18007]_ ) & (~\m6_data_i[3]  | ~\new_[18086]_ );
  assign \new_[13444]_  = (~\m5_addr_i[16]  | ~\new_[17188]_ ) & (~\m6_addr_i[16]  | ~\new_[18050]_ );
  assign \new_[13445]_  = (~\m5_data_i[2]  | ~\new_[18007]_ ) & (~\m6_data_i[2]  | ~\new_[18086]_ );
  assign \new_[13446]_  = (~\m4_data_i[2]  | ~\new_[17267]_ ) & (~\m3_data_i[2]  | ~\new_[18206]_ );
  assign \new_[13447]_  = (~\m5_data_i[1]  | ~\new_[18007]_ ) & (~\m6_data_i[1]  | ~\new_[18086]_ );
  assign \new_[13448]_  = (~\m4_data_i[1]  | ~\new_[17267]_ ) & (~\m3_data_i[1]  | ~\new_[18206]_ );
  assign \new_[13449]_  = (~\new_[19577]_  | ~\m6_addr_i[31] ) & (~\new_[18007]_  | ~\new_[31001]_ );
  assign \new_[13450]_  = (~\new_[17221]_  | ~\m2_addr_i[31] ) & (~\new_[17274]_  | ~\new_[31447]_ );
  assign \new_[13451]_  = (~\new_[17267]_  | ~\m4_addr_i[31] ) & (~\new_[18206]_  | ~\m3_addr_i[31] );
  assign \new_[13452]_  = (~\new_[17267]_  | ~\m4_addr_i[30] ) & (~\new_[18206]_  | ~\m3_addr_i[30] );
  assign \new_[13453]_  = (~\new_[17221]_  | ~\m2_addr_i[29] ) & (~\new_[17274]_  | ~\new_[31538]_ );
  assign \new_[13454]_  = (~\new_[19577]_  | ~\m6_addr_i[28] ) & (~\new_[18007]_  | ~\new_[31276]_ );
  assign \new_[13455]_  = (~\new_[19577]_  | ~\m6_addr_i[27] ) & (~\new_[18007]_  | ~\m5_addr_i[27] );
  assign \new_[13456]_  = (~\new_[19577]_  | ~\m6_addr_i[26] ) & (~\new_[18007]_  | ~\m5_addr_i[26] );
  assign \new_[13457]_  = (~\new_[17267]_  | ~\m4_addr_i[26] ) & (~\new_[18206]_  | ~\m3_addr_i[26] );
  assign \new_[13458]_  = (~\new_[17221]_  | ~\m2_addr_i[26] ) & (~\new_[18180]_  | ~\m1_addr_i[26] );
  assign \new_[13459]_  = (~\m3_sel_i[3]  | ~\new_[32350]_ ) & (~\m2_sel_i[3]  | ~\new_[18808]_ );
  assign \new_[13460]_  = (~\new_[17221]_  | ~\m2_addr_i[25] ) & (~\new_[17274]_  | ~\m1_addr_i[25] );
  assign \new_[13461]_  = (~\new_[17221]_  | ~\m2_addr_i[24] ) & (~\new_[18180]_  | ~\m1_addr_i[24] );
  assign \new_[13462]_  = (~\m5_addr_i[23]  | ~\new_[18007]_ ) & (~\m6_addr_i[23]  | ~\new_[18087]_ );
  assign \new_[13463]_  = (~\m5_addr_i[22]  | ~\new_[18007]_ ) & (~\m6_addr_i[22]  | ~\new_[18087]_ );
  assign \new_[13464]_  = ~\new_[28938]_  | (~\new_[17421]_  & ~\new_[24780]_ );
  assign \new_[13465]_  = ~\new_[30303]_  & (~\new_[17397]_  | ~\new_[23051]_ );
  assign \new_[13466]_  = (~\m5_addr_i[19]  | ~\new_[18007]_ ) & (~\m6_addr_i[19]  | ~\new_[18086]_ );
  assign \new_[13467]_  = (~\m5_addr_i[16]  | ~\new_[18007]_ ) & (~\m6_addr_i[16]  | ~\new_[18086]_ );
  assign \new_[13468]_  = (~\m5_addr_i[15]  | ~\new_[18007]_ ) & (~\m6_addr_i[15]  | ~\new_[18086]_ );
  assign \new_[13469]_  = (~\m5_addr_i[14]  | ~\new_[18007]_ ) & (~\m6_addr_i[14]  | ~\new_[18086]_ );
  assign \new_[13470]_  = (~\m5_addr_i[12]  | ~\new_[18007]_ ) & (~\m6_addr_i[12]  | ~\new_[18086]_ );
  assign \new_[13471]_  = (~\m5_addr_i[9]  | ~\new_[18007]_ ) & (~\m6_addr_i[9]  | ~\new_[18087]_ );
  assign \new_[13472]_  = (~\m5_addr_i[5]  | ~\new_[18007]_ ) & (~\m6_addr_i[5]  | ~\new_[18087]_ );
  assign \new_[13473]_  = (~\m4_addr_i[4]  | ~\new_[17267]_ ) & (~\m3_addr_i[4]  | ~\new_[18206]_ );
  assign \new_[13474]_  = (~\m2_addr_i[2]  | ~\new_[17221]_ ) & (~\new_[31477]_  | ~\new_[17275]_ );
  assign \new_[13475]_  = ~\new_[29986]_  & (~\new_[17398]_  | ~\new_[20743]_ );
  assign \new_[13476]_  = (~\m5_addr_i[1]  | ~\new_[18007]_ ) & (~\m6_addr_i[1]  | ~\new_[18087]_ );
  assign \new_[13477]_  = (~\m5_addr_i[0]  | ~\new_[18007]_ ) & (~\m6_addr_i[0]  | ~\new_[18086]_ );
  assign \new_[13478]_  = (~\m5_sel_i[3]  | ~\new_[18007]_ ) & (~\m6_sel_i[3]  | ~\new_[19577]_ );
  assign \new_[13479]_  = (~\m5_sel_i[2]  | ~\new_[18007]_ ) & (~\m6_sel_i[2]  | ~\new_[19577]_ );
  assign \new_[13480]_  = (~\m4_sel_i[2]  | ~\new_[17267]_ ) & (~\m3_sel_i[2]  | ~\new_[18206]_ );
  assign \new_[13481]_  = (~\m5_sel_i[1]  | ~\new_[18007]_ ) & (~\m6_sel_i[1]  | ~\new_[19577]_ );
  assign \new_[13482]_  = (~\m4_sel_i[1]  | ~\new_[17267]_ ) & (~\m3_sel_i[1]  | ~\new_[18206]_ );
  assign \new_[13483]_  = (~\m2_data_i[31]  | ~\new_[18805]_ ) & (~\m1_data_i[31]  | ~\new_[18913]_ );
  assign \new_[13484]_  = (~\m7_data_i[25]  | ~\new_[18832]_ ) & (~\m0_data_i[25]  | ~\new_[18066]_ );
  assign \new_[13485]_  = ~\new_[28443]_  & (~\new_[17399]_  | ~\new_[20502]_ );
  assign \new_[13486]_  = (~\m7_data_i[24]  | ~\new_[18832]_ ) & (~\m0_data_i[24]  | ~\new_[18066]_ );
  assign \new_[13487]_  = ~\new_[14852]_ ;
  assign \new_[13488]_  = (~\m2_data_i[22]  | ~\new_[20555]_ ) & (~\m1_data_i[22]  | ~\new_[18913]_ );
  assign \new_[13489]_  = (~\m7_data_i[20]  | ~\new_[18832]_ ) & (~\m0_data_i[20]  | ~\new_[18066]_ );
  assign \new_[13490]_  = (~\m7_addr_i[1]  | ~\new_[18116]_ ) & (~\m0_addr_i[1]  | ~\new_[18932]_ );
  assign \new_[13491]_  = ~\new_[20288]_  & (~\new_[17206]_  | ~\new_[30030]_ );
  assign \new_[13492]_  = ~\new_[30122]_  & (~\new_[17400]_  | ~\new_[24315]_ );
  assign \new_[13493]_  = ~\new_[17269]_ ;
  assign \new_[13494]_  = (~\m2_data_i[18]  | ~\new_[20555]_ ) & (~\m1_data_i[18]  | ~\new_[18913]_ );
  assign \new_[13495]_  = ~\new_[28697]_  & (~\new_[17408]_  | ~\new_[22730]_ );
  assign \new_[13496]_  = (~\m7_data_i[16]  | ~\new_[18832]_ ) & (~\m0_data_i[16]  | ~\new_[18066]_ );
  assign \new_[13497]_  = (~\m2_data_i[16]  | ~\new_[18799]_ ) & (~\m1_data_i[16]  | ~\new_[18887]_ );
  assign \new_[13498]_  = (~\m2_data_i[15]  | ~\new_[18804]_ ) & (~\m1_data_i[15]  | ~\new_[17276]_ );
  assign \new_[13499]_  = (~\m7_data_i[15]  | ~\new_[18832]_ ) & (~\m0_data_i[15]  | ~\new_[18066]_ );
  assign \new_[13500]_  = (~\m2_data_i[14]  | ~\new_[20555]_ ) & (~\m1_data_i[14]  | ~\new_[17276]_ );
  assign \new_[13501]_  = (~\m7_data_i[14]  | ~\new_[18832]_ ) & (~\m0_data_i[14]  | ~\new_[18066]_ );
  assign \new_[13502]_  = (~\m2_data_i[13]  | ~\new_[20555]_ ) & (~\m1_data_i[13]  | ~\new_[17276]_ );
  assign \new_[13503]_  = (~\m7_data_i[13]  | ~\new_[18832]_ ) & (~\m0_data_i[13]  | ~\new_[18066]_ );
  assign \new_[13504]_  = (~\new_[17388]_  | ~\new_[29694]_ ) & (~\new_[26152]_  | ~\new_[29694]_ );
  assign \new_[13505]_  = (~\m7_data_i[12]  | ~\new_[18832]_ ) & (~\m0_data_i[12]  | ~\new_[18066]_ );
  assign \new_[13506]_  = (~\m5_addr_i[2]  | ~\new_[17189]_ ) & (~\m6_addr_i[2]  | ~\new_[18051]_ );
  assign \new_[13507]_  = (~\m2_data_i[11]  | ~\new_[20555]_ ) & (~\m1_data_i[11]  | ~\new_[18913]_ );
  assign \new_[13508]_  = (~\new_[17389]_  | ~\new_[29194]_ ) & (~\new_[22785]_  | ~\new_[29194]_ );
  assign \new_[13509]_  = (~\m2_data_i[9]  | ~\new_[18805]_ ) & (~\m1_data_i[9]  | ~\new_[18913]_ );
  assign \new_[13510]_  = (~\m7_data_i[7]  | ~\new_[18832]_ ) & (~\m0_data_i[7]  | ~\new_[18066]_ );
  assign \new_[13511]_  = (~\m7_data_i[6]  | ~\new_[18832]_ ) & (~\m0_data_i[6]  | ~\new_[18066]_ );
  assign \new_[13512]_  = (~\m2_data_i[6]  | ~\new_[20555]_ ) & (~\m1_data_i[6]  | ~\new_[18913]_ );
  assign \new_[13513]_  = (~\m2_data_i[5]  | ~\new_[18804]_ ) & (~\m1_data_i[5]  | ~\new_[17276]_ );
  assign \new_[13514]_  = (~\m7_data_i[5]  | ~\new_[18832]_ ) & (~\m0_data_i[5]  | ~\new_[18066]_ );
  assign \new_[13515]_  = (~\m2_data_i[4]  | ~\new_[18804]_ ) & (~\m1_data_i[4]  | ~\new_[17276]_ );
  assign \new_[13516]_  = (~\m2_data_i[3]  | ~\new_[20555]_ ) & (~\m1_data_i[3]  | ~\new_[18913]_ );
  assign \new_[13517]_  = (~\m2_data_i[2]  | ~\new_[18804]_ ) & (~\m1_data_i[2]  | ~\new_[17276]_ );
  assign \new_[13518]_  = (~\m7_data_i[2]  | ~\new_[18832]_ ) & (~\m0_data_i[2]  | ~\new_[18066]_ );
  assign \new_[13519]_  = (~\m2_data_i[0]  | ~\new_[20555]_ ) & (~\m1_data_i[0]  | ~\new_[18913]_ );
  assign \new_[13520]_  = (~\new_[20555]_  | ~\m2_addr_i[31] ) & (~\new_[18913]_  | ~\new_[31447]_ );
  assign \new_[13521]_  = (~\new_[18832]_  | ~\new_[31531]_ ) & (~\new_[18066]_  | ~\new_[31481]_ );
  assign \new_[13522]_  = (~\new_[20555]_  | ~\m2_addr_i[29] ) & (~\new_[18913]_  | ~\new_[31538]_ );
  assign \new_[13523]_  = (~\new_[17394]_  | ~\new_[29494]_ ) & (~\new_[21423]_  | ~\new_[29494]_ );
  assign \new_[13524]_  = (~\new_[18804]_  | ~\m2_addr_i[25] ) & (~\new_[18913]_  | ~\m1_addr_i[25] );
  assign \new_[13525]_  = \new_[14880]_ ;
  assign \new_[13526]_  = \new_[14880]_ ;
  assign \new_[13527]_  = ~\new_[16336]_  & ~\new_[19372]_ ;
  assign \new_[13528]_  = (~\m4_sel_i[0]  | ~\new_[17260]_ ) & (~\m3_sel_i[0]  | ~\new_[18175]_ );
  assign \new_[13529]_  = (~\m2_addr_i[16]  | ~\new_[18804]_ ) & (~\m1_addr_i[16]  | ~\new_[18913]_ );
  assign \new_[13530]_  = ~\new_[14888]_ ;
  assign \new_[13531]_  = \new_[6006]_  ? \new_[29130]_  : \new_[17345]_ ;
  assign \new_[13532]_  = (~\m2_addr_i[15]  | ~\new_[18804]_ ) & (~\m1_addr_i[15]  | ~\new_[18913]_ );
  assign \new_[13533]_  = (~\m2_addr_i[14]  | ~\new_[18804]_ ) & (~\m1_addr_i[14]  | ~\new_[18913]_ );
  assign \new_[13534]_  = (~\m2_addr_i[13]  | ~\new_[18805]_ ) & (~\m1_addr_i[13]  | ~\new_[18913]_ );
  assign \new_[13535]_  = (~\new_[17380]_  | ~\new_[29662]_ ) & (~\new_[22714]_  | ~\new_[29662]_ );
  assign \new_[13536]_  = (~\new_[17381]_  | ~\new_[29000]_ ) & (~\new_[22784]_  | ~\new_[29000]_ );
  assign \new_[13537]_  = (~\m2_addr_i[8]  | ~\new_[20555]_ ) & (~\m1_addr_i[8]  | ~\new_[18913]_ );
  assign \new_[13538]_  = (~\m2_addr_i[7]  | ~\new_[18804]_ ) & (~\m1_addr_i[7]  | ~\new_[17276]_ );
  assign \new_[13539]_  = ~\new_[14895]_ ;
  assign \new_[13540]_  = (~\m2_addr_i[6]  | ~\new_[20555]_ ) & (~\m1_addr_i[6]  | ~\new_[17276]_ );
  assign \new_[13541]_  = (~\new_[31095]_  | ~\new_[20555]_ ) & (~\m1_addr_i[5]  | ~\new_[18913]_ );
  assign \new_[13542]_  = (~\m2_addr_i[4]  | ~\new_[18805]_ ) & (~\m1_addr_i[4]  | ~\new_[18913]_ );
  assign \new_[13543]_  = (~\new_[31399]_  | ~\new_[18805]_ ) & (~\m1_addr_i[3]  | ~\new_[18913]_ );
  assign \new_[13544]_  = (~\m2_addr_i[2]  | ~\new_[20555]_ ) & (~\new_[31477]_  | ~\new_[18913]_ );
  assign \new_[13545]_  = (~\m5_addr_i[3]  | ~\new_[17189]_ ) & (~\m6_addr_i[3]  | ~\new_[18051]_ );
  assign \new_[13546]_  = (~\m5_sel_i[1]  | ~\new_[17188]_ ) & (~\m6_sel_i[1]  | ~\new_[19563]_ );
  assign \new_[13547]_  = (~\m2_addr_i[1]  | ~\new_[18804]_ ) & (~\m1_addr_i[1]  | ~\new_[18913]_ );
  assign \new_[13548]_  = (~\m2_sel_i[0]  | ~\new_[20555]_ ) & (~\m1_sel_i[0]  | ~\new_[18913]_ );
  assign \new_[13549]_  = (~m7_we_i | ~\new_[18832]_ ) & (~m0_we_i | ~\new_[18066]_ );
  assign \new_[13550]_  = (~m2_we_i | ~\new_[20555]_ ) & (~m1_we_i | ~\new_[17276]_ );
  assign \new_[13551]_  = (~\m2_data_i[24]  | ~\new_[18799]_ ) & (~\m1_data_i[24]  | ~\new_[18887]_ );
  assign \new_[13552]_  = (~\new_[17385]_  | ~\new_[30027]_ ) & (~\new_[21388]_  | ~\new_[30027]_ );
  assign \new_[13553]_  = (~\new_[17386]_  | ~\new_[28901]_ ) & (~\new_[21433]_  | ~\new_[28901]_ );
  assign \new_[13554]_  = ~\new_[16426]_  | ~\new_[28247]_ ;
  assign \new_[13555]_  = ~\new_[16428]_  | ~\new_[28670]_ ;
  assign \new_[13556]_  = ~\new_[16430]_  | ~\new_[28279]_ ;
  assign \new_[13557]_  = ~\new_[16437]_  | ~\new_[30194]_ ;
  assign \new_[13558]_  = ~\new_[16379]_  | ~\new_[24653]_ ;
  assign \new_[13559]_  = ~\new_[16443]_  | ~\new_[28071]_ ;
  assign \new_[13560]_  = ~\new_[16451]_  | ~\new_[30300]_ ;
  assign \new_[13561]_  = ~\new_[16453]_  | ~\new_[28671]_ ;
  assign \new_[13562]_  = ~\new_[16455]_  | ~\new_[30156]_ ;
  assign \new_[13563]_  = ~\new_[16460]_  | ~\new_[29078]_ ;
  assign \new_[13564]_  = ~\new_[16461]_  | ~\new_[28299]_ ;
  assign \new_[13565]_  = ~\new_[21516]_  | ~\new_[26570]_  | ~\new_[17457]_ ;
  assign \new_[13566]_  = ~\new_[16478]_  & ~\new_[28301]_ ;
  assign \new_[13567]_  = ~\new_[16493]_  | ~\new_[28585]_ ;
  assign \new_[13568]_  = ~\new_[16705]_  | ~\new_[28527]_  | ~\new_[22703]_ ;
  assign \new_[13569]_  = \new_[16510]_  | \new_[24008]_ ;
  assign \new_[13570]_  = \new_[16512]_  | \new_[24998]_ ;
  assign \new_[13571]_  = ~\new_[20295]_  & (~\new_[17259]_  | ~\new_[29268]_ );
  assign \new_[13572]_  = ~\new_[16479]_  & ~\new_[28228]_ ;
  assign \new_[13573]_  = ~\new_[16706]_  | ~\new_[28586]_  | ~\new_[24231]_ ;
  assign \new_[13574]_  = ~\new_[16707]_  | ~\new_[29026]_  | ~\new_[26216]_ ;
  assign \new_[13575]_  = \new_[6003]_  ? \new_[29569]_  : \new_[17340]_ ;
  assign \new_[13576]_  = ~\new_[16480]_  & ~\new_[28803]_ ;
  assign \new_[13577]_  = (~\m2_data_i[31]  | ~\new_[18069]_ ) & (~\m1_data_i[31]  | ~\new_[20573]_ );
  assign \new_[13578]_  = ~\new_[16708]_  | ~\new_[26901]_  | ~\new_[24203]_ ;
  assign \new_[13579]_  = ~\new_[16481]_  & ~\new_[28531]_ ;
  assign \new_[13580]_  = ~\new_[16709]_  | ~\new_[27552]_  | ~\new_[22692]_ ;
  assign \new_[13581]_  = ~\new_[16482]_  & ~\new_[26453]_ ;
  assign \new_[13582]_  = ~\new_[16710]_  | ~\new_[29311]_  | ~\new_[24117]_ ;
  assign \new_[13583]_  = ~\new_[16439]_  | ~\new_[26789]_ ;
  assign \new_[13584]_  = ~\new_[16440]_  | ~\new_[27792]_ ;
  assign \new_[13585]_  = ~\new_[16484]_  & ~\new_[27707]_ ;
  assign \new_[13586]_  = ~\new_[16711]_  | ~\new_[28116]_  | ~\new_[21391]_ ;
  assign \new_[13587]_  = ~\new_[16712]_  | ~\new_[29249]_  | ~\new_[24238]_ ;
  assign \new_[13588]_  = ~\new_[16485]_  & ~\new_[27801]_ ;
  assign \new_[13589]_  = ~\new_[16497]_  | ~\new_[28550]_ ;
  assign \new_[13590]_  = ~\new_[16445]_  | ~\new_[28416]_ ;
  assign \new_[13591]_  = ~\new_[16713]_  | ~\new_[27646]_  | ~\new_[24198]_ ;
  assign \new_[13592]_  = (~\m5_sel_i[2]  | ~\new_[17187]_ ) & (~\m6_sel_i[2]  | ~\new_[19563]_ );
  assign \new_[13593]_  = ~\new_[16486]_  & ~\new_[25466]_ ;
  assign \new_[13594]_  = ~\new_[16714]_  | ~\new_[28480]_  | ~\new_[22580]_ ;
  assign \new_[13595]_  = (~\m5_addr_i[4]  | ~\new_[17189]_ ) & (~\m6_addr_i[4]  | ~\new_[18051]_ );
  assign \new_[13596]_  = ~\new_[16487]_  & ~\new_[25006]_ ;
  assign \new_[13597]_  = \new_[16523]_  | \new_[26426]_ ;
  assign \new_[13598]_  = ~\new_[16488]_  & ~\new_[28340]_ ;
  assign \new_[13599]_  = ~\new_[16489]_  & ~\new_[26254]_ ;
  assign \new_[13600]_  = \new_[6068]_  ? \new_[29145]_  : \new_[17333]_ ;
  assign \new_[13601]_  = (~\m4_sel_i[2]  | ~\new_[17260]_ ) & (~\m3_sel_i[2]  | ~\new_[18175]_ );
  assign \new_[13602]_  = ~\new_[16715]_  | ~\new_[28632]_  | ~\new_[22839]_ ;
  assign \new_[13603]_  = ~\new_[16716]_  | ~\new_[28523]_  | ~\new_[21440]_ ;
  assign \new_[13604]_  = \new_[16526]_  | \new_[27677]_ ;
  assign \new_[13605]_  = ~\new_[16490]_  & ~\new_[28584]_ ;
  assign \new_[13606]_  = \new_[6086]_  ? \new_[30149]_  : \new_[17322]_ ;
  assign \new_[13607]_  = ~\new_[16717]_  | ~\new_[27694]_  | ~\new_[22667]_ ;
  assign \new_[13608]_  = ~\new_[22133]_  & (~\new_[17243]_  | ~\new_[28924]_ );
  assign \new_[13609]_  = ~\new_[16491]_  & ~\new_[27690]_ ;
  assign \new_[13610]_  = ~\new_[16718]_  | ~\new_[27578]_  | ~\new_[22570]_ ;
  assign \new_[13611]_  = ~\new_[16719]_  | ~\new_[29449]_  | ~\new_[25590]_ ;
  assign \new_[13612]_  = ~\new_[16492]_  & ~\new_[27622]_ ;
  assign \new_[13613]_  = \new_[17343]_  ? \new_[30618]_  : \new_[6194]_ ;
  assign \new_[13614]_  = ~\new_[16720]_  | ~\new_[28569]_  | ~\new_[24244]_ ;
  assign \new_[13615]_  = (~\m7_addr_i[4]  | ~\new_[18116]_ ) & (~\m0_addr_i[4]  | ~\new_[18932]_ );
  assign \new_[13616]_  = \new_[16531]_  | \new_[24780]_ ;
  assign \new_[13617]_  = ~\new_[17436]_  | ~\new_[26303]_  | ~\new_[21359]_ ;
  assign \new_[13618]_  = ~\new_[28680]_  & (~\new_[17437]_  | ~\new_[22813]_ );
  assign \new_[13619]_  = ~\new_[17440]_  | ~\new_[28586]_  | ~\new_[24215]_ ;
  assign \new_[13620]_  = ~\new_[17441]_  | ~\new_[29026]_  | ~\new_[26155]_ ;
  assign \new_[13621]_  = ~\new_[17444]_  | ~\new_[26901]_  | ~\new_[23128]_ ;
  assign \new_[13622]_  = ~\new_[17445]_  | ~\new_[26580]_  | ~\new_[22758]_ ;
  assign \new_[13623]_  = (~\m2_data_i[10]  | ~\new_[18799]_ ) & (~\m1_data_i[10]  | ~\new_[20571]_ );
  assign \new_[13624]_  = ~\new_[17449]_  | ~\new_[27552]_  | ~\new_[22731]_ ;
  assign \new_[13625]_  = ~\new_[28028]_  & (~\new_[17450]_  | ~\new_[22342]_ );
  assign \new_[13626]_  = ~\new_[17455]_  | ~\new_[29311]_  | ~\new_[24239]_ ;
  assign \new_[13627]_  = ~\new_[17456]_  | ~\new_[26865]_  | ~\new_[21384]_ ;
  assign \new_[13628]_  = ~\new_[17461]_  | ~\new_[28144]_  | ~\new_[22760]_ ;
  assign \new_[13629]_  = ~\new_[17465]_  | ~\new_[28116]_  | ~\new_[21426]_ ;
  assign \new_[13630]_  = ~\new_[17466]_  | ~\new_[24684]_  | ~\new_[22742]_ ;
  assign \new_[13631]_  = ~\new_[17467]_  | ~\new_[29249]_  | ~\new_[24224]_ ;
  assign \new_[13632]_  = ~\new_[17468]_  | ~\new_[27627]_  | ~\new_[21399]_ ;
  assign \new_[13633]_  = ~\new_[17473]_  | ~\new_[27646]_  | ~\new_[24232]_ ;
  assign \new_[13634]_  = ~\new_[17474]_  | ~\new_[24441]_  | ~\new_[20411]_ ;
  assign \new_[13635]_  = ~\new_[17477]_  | ~\new_[28480]_  | ~\new_[22759]_ ;
  assign \new_[13636]_  = ~\new_[17478]_  | ~\new_[26312]_  | ~\new_[22565]_ ;
  assign \new_[13637]_  = ~\new_[17482]_  | ~\new_[28540]_  | ~\new_[24250]_ ;
  assign \new_[13638]_  = ~\new_[17485]_  | ~\new_[27648]_  | ~\new_[22212]_ ;
  assign \new_[13639]_  = ~\new_[17486]_  | ~\new_[26338]_  | ~\new_[21406]_ ;
  assign \new_[13640]_  = ~\new_[17487]_  | ~\new_[24364]_  | ~\new_[22770]_ ;
  assign \new_[13641]_  = ~\new_[17491]_  | ~\new_[28632]_  | ~\new_[22747]_ ;
  assign \new_[13642]_  = ~\new_[17492]_  | ~\new_[26520]_  | ~\new_[22740]_ ;
  assign \new_[13643]_  = (~\m2_data_i[11]  | ~\new_[18806]_ ) & (~\m1_data_i[11]  | ~\new_[17273]_ );
  assign \new_[13644]_  = ~\new_[17494]_  | ~\new_[26435]_  | ~\new_[22376]_ ;
  assign \new_[13645]_  = ~\new_[17497]_  | ~\new_[26346]_  | ~\new_[21235]_ ;
  assign \new_[13646]_  = (~\m2_data_i[4]  | ~\new_[18806]_ ) & (~\m1_data_i[4]  | ~\new_[17273]_ );
  assign \new_[13647]_  = ~\new_[17498]_  | ~\new_[23135]_  | ~\new_[21366]_ ;
  assign \new_[13648]_  = ~\new_[29838]_  & (~\new_[17501]_  | ~\new_[23039]_ );
  assign \new_[13649]_  = ~\new_[17502]_  | ~\new_[26594]_  | ~\new_[24220]_ ;
  assign \new_[13650]_  = (~\m5_addr_i[5]  | ~\new_[17189]_ ) & (~\m6_addr_i[5]  | ~\new_[18051]_ );
  assign \new_[13651]_  = ~\new_[17508]_  | ~\new_[26205]_  | ~\new_[22701]_ ;
  assign \new_[13652]_  = ~\new_[21220]_  | ~\new_[16378]_ ;
  assign \new_[13653]_  = ~\new_[26642]_  & (~\new_[16748]_  | ~\new_[27662]_ );
  assign \new_[13654]_  = ~\new_[26989]_  | ~\new_[16372]_ ;
  assign \new_[13655]_  = ~\new_[20343]_  & (~\new_[17244]_  | ~\new_[29248]_ );
  assign \new_[13656]_  = ~\new_[25264]_  | ~\new_[16389]_ ;
  assign \new_[13657]_  = (~\new_[18806]_  | ~\m2_addr_i[24] ) & (~\new_[17273]_  | ~\m1_addr_i[24] );
  assign \new_[13658]_  = (~\m5_addr_i[22]  | ~\new_[17199]_ ) & (~\m6_addr_i[22]  | ~\new_[20551]_ );
  assign \new_[13659]_  = ~\new_[29942]_  & (~\new_[17402]_  | ~\new_[21499]_ );
  assign \new_[13660]_  = (~\m2_data_i[22]  | ~\new_[18068]_ ) & (~\m1_data_i[22]  | ~\new_[20573]_ );
  assign \new_[13661]_  = ~\new_[29076]_  & (~\new_[17349]_  | ~\new_[21525]_ );
  assign \new_[13662]_  = ~\new_[28875]_  & (~\new_[16740]_  | ~\new_[28585]_ );
  assign \new_[13663]_  = \new_[16397]_  & \new_[28693]_ ;
  assign \new_[13664]_  = \new_[16398]_  & \new_[28701]_ ;
  assign \new_[13665]_  = (~\m2_addr_i[18]  | ~\new_[18806]_ ) & (~\m1_addr_i[18]  | ~\new_[17273]_ );
  assign \new_[13666]_  = \new_[16399]_  & \new_[30077]_ ;
  assign \new_[13667]_  = \new_[16401]_  & \new_[29658]_ ;
  assign \new_[13668]_  = ~\new_[23097]_  & (~\new_[16746]_  | ~\new_[28167]_ );
  assign \new_[13669]_  = ~\new_[26665]_  & (~\new_[16749]_  | ~\new_[28164]_ );
  assign \new_[13670]_  = ~\new_[28991]_  & (~\new_[16751]_  | ~\new_[28550]_ );
  assign \new_[13671]_  = \new_[16409]_  & \new_[29301]_ ;
  assign \new_[13672]_  = ~\new_[29716]_  & (~\new_[16742]_  | ~\new_[28122]_ );
  assign \new_[13673]_  = \new_[16413]_  & \new_[29193]_ ;
  assign \new_[13674]_  = ~\new_[28763]_  & (~\new_[16758]_  | ~\new_[28297]_ );
  assign \new_[13675]_  = \new_[16418]_  & \new_[29630]_ ;
  assign \new_[13676]_  = ~\new_[28026]_  & (~\new_[16761]_  | ~\new_[28306]_ );
  assign \new_[13677]_  = \new_[16406]_  & \new_[28200]_ ;
  assign \new_[13678]_  = ~\new_[27871]_  & (~\new_[16762]_  | ~\new_[28241]_ );
  assign \new_[13679]_  = \new_[16425]_  & \new_[28938]_ ;
  assign \new_[13680]_  = ~\new_[26682]_  & (~\new_[16763]_  | ~\new_[24194]_ );
  assign \new_[13681]_  = ~\new_[29620]_  & (~\new_[16775]_  | ~\new_[24382]_ );
  assign \new_[13682]_  = (~\m4_sel_i[3]  | ~\new_[17260]_ ) & (~\m3_sel_i[3]  | ~\new_[18175]_ );
  assign \new_[13683]_  = (~\new_[31399]_  | ~\new_[18806]_ ) & (~\m1_addr_i[3]  | ~\new_[18906]_ );
  assign \new_[13684]_  = ~\new_[26669]_  & (~\new_[16776]_  | ~\new_[24381]_ );
  assign \new_[13685]_  = ~\new_[28258]_  & (~\new_[16764]_  | ~\new_[24212]_ );
  assign \new_[13686]_  = ~\new_[27921]_  & (~\new_[16765]_  | ~\new_[25313]_ );
  assign \new_[13687]_  = \new_[6063]_  ? \new_[28865]_  : \new_[17321]_ ;
  assign \new_[13688]_  = ~\new_[26621]_  & (~\new_[16766]_  | ~\new_[21380]_ );
  assign \new_[13689]_  = ~\new_[26542]_  & (~\new_[16767]_  | ~\new_[24005]_ );
  assign \new_[13690]_  = (~\m4_addr_i[17]  | ~\new_[18149]_ ) & (~\m3_addr_i[17]  | ~\new_[18930]_ );
  assign \new_[13691]_  = ~\new_[28146]_  & (~\new_[16768]_  | ~\new_[26249]_ );
  assign \new_[13692]_  = (~\m3_data_i[21]  | ~\new_[32350]_ ) & (~\m2_data_i[21]  | ~\new_[18808]_ );
  assign \new_[13693]_  = (~\m3_data_i[20]  | ~\new_[32350]_ ) & (~\m2_data_i[20]  | ~\new_[18808]_ );
  assign \new_[13694]_  = ~\new_[28315]_  & (~\new_[16769]_  | ~\new_[24020]_ );
  assign \new_[13695]_  = ~\new_[28104]_  & (~\new_[16778]_  | ~\new_[24297]_ );
  assign \new_[13696]_  = (~\m3_data_i[19]  | ~\new_[32350]_ ) & (~\m2_data_i[19]  | ~\new_[17224]_ );
  assign \new_[13697]_  = ~\new_[26816]_  & (~\new_[16770]_  | ~\new_[24091]_ );
  assign \new_[13698]_  = (~\m5_data_i[31]  | ~\new_[17199]_ ) & (~\m6_data_i[31]  | ~\new_[18789]_ );
  assign \new_[13699]_  = ~\new_[30330]_  & (~\new_[16777]_  | ~\new_[24271]_ );
  assign \new_[13700]_  = (~\m4_data_i[30]  | ~\new_[18156]_ ) & (~\m3_data_i[30]  | ~\new_[18130]_ );
  assign \new_[13701]_  = (~\m5_data_i[29]  | ~\new_[17199]_ ) & (~\m6_data_i[29]  | ~\new_[20551]_ );
  assign \new_[13702]_  = ~\new_[27764]_  & (~\new_[16771]_  | ~\new_[21351]_ );
  assign \new_[13703]_  = ~\new_[27886]_  & (~\new_[16772]_  | ~\new_[24248]_ );
  assign \new_[13704]_  = ~\new_[18476]_  | ~\new_[18477]_  | ~\new_[16677]_  | ~\new_[17553]_ ;
  assign \new_[13705]_  = ~\new_[24660]_  & (~\new_[16779]_  | ~\new_[24375]_ );
  assign \new_[13706]_  = (~\m4_data_i[28]  | ~\new_[18156]_ ) & (~\m3_data_i[28]  | ~\new_[18130]_ );
  assign \new_[13707]_  = (~\m5_data_i[27]  | ~\new_[17199]_ ) & (~\m6_data_i[27]  | ~\new_[18789]_ );
  assign \new_[13708]_  = (~\m5_data_i[26]  | ~\new_[17199]_ ) & (~\m6_data_i[26]  | ~\new_[20551]_ );
  assign \new_[13709]_  = (~\m5_data_i[25]  | ~\new_[17199]_ ) & (~\m6_data_i[25]  | ~\new_[19561]_ );
  assign \new_[13710]_  = ~\new_[27856]_  & (~\new_[16773]_  | ~\new_[26165]_ );
  assign \new_[13711]_  = (~\m3_data_i[17]  | ~\new_[32350]_ ) & (~\m2_data_i[17]  | ~\new_[18808]_ );
  assign \new_[13712]_  = (~\m5_data_i[24]  | ~\new_[17199]_ ) & (~\m6_data_i[24]  | ~\new_[20551]_ );
  assign \new_[13713]_  = (~\m4_data_i[24]  | ~\new_[18156]_ ) & (~\m3_data_i[24]  | ~\new_[18130]_ );
  assign \new_[13714]_  = (~\m5_data_i[23]  | ~\new_[17199]_ ) & (~\m6_data_i[23]  | ~\new_[19561]_ );
  assign \new_[13715]_  = (~\m5_data_i[22]  | ~\new_[17201]_ ) & (~\m6_data_i[22]  | ~\new_[20551]_ );
  assign \new_[13716]_  = (~\m5_data_i[21]  | ~\new_[17199]_ ) & (~\m6_data_i[21]  | ~\new_[18789]_ );
  assign \new_[13717]_  = (~\m5_data_i[20]  | ~\new_[17199]_ ) & (~\m6_data_i[20]  | ~\new_[18789]_ );
  assign \new_[13718]_  = (~\m5_addr_i[20]  | ~\new_[17187]_ ) & (~\m6_addr_i[20]  | ~\new_[18050]_ );
  assign \new_[13719]_  = (~\m5_data_i[18]  | ~\new_[17199]_ ) & (~\m6_data_i[18]  | ~\new_[18789]_ );
  assign \new_[13720]_  = (~\m4_data_i[18]  | ~\new_[18156]_ ) & (~\m3_data_i[18]  | ~\new_[18130]_ );
  assign \new_[13721]_  = (~\m5_data_i[17]  | ~\new_[17201]_ ) & (~\m6_data_i[17]  | ~\new_[20551]_ );
  assign \new_[13722]_  = (~\m5_data_i[16]  | ~\new_[17199]_ ) & (~\m6_data_i[16]  | ~\new_[18789]_ );
  assign \new_[13723]_  = (~\m4_data_i[16]  | ~\new_[18156]_ ) & (~\m3_data_i[16]  | ~\new_[18130]_ );
  assign \new_[13724]_  = (~\m4_addr_i[20]  | ~\new_[17260]_ ) & (~\m3_addr_i[20]  | ~\new_[18175]_ );
  assign \new_[13725]_  = (~\m3_data_i[14]  | ~\new_[32350]_ ) & (~\m2_data_i[14]  | ~\new_[17224]_ );
  assign \new_[13726]_  = (~\m5_data_i[15]  | ~\new_[19544]_ ) & (~\m6_data_i[15]  | ~\new_[18789]_ );
  assign \new_[13727]_  = (~\m5_data_i[14]  | ~\new_[19544]_ ) & (~\m6_data_i[14]  | ~\new_[20551]_ );
  assign \new_[13728]_  = (~\m5_data_i[13]  | ~\new_[17201]_ ) & (~\m6_data_i[13]  | ~\new_[20551]_ );
  assign \new_[13729]_  = (~\m5_data_i[12]  | ~\new_[17199]_ ) & (~\m6_data_i[12]  | ~\new_[19561]_ );
  assign \new_[13730]_  = ~\new_[27899]_  & (~\new_[16774]_  | ~\new_[26185]_ );
  assign \new_[13731]_  = (~\m3_data_i[13]  | ~\new_[18936]_ ) & (~\m2_data_i[13]  | ~\new_[17224]_ );
  assign \new_[13732]_  = ~\new_[29659]_  & (~\new_[17379]_  | ~\new_[22947]_ );
  assign \new_[13733]_  = (~\m5_data_i[11]  | ~\new_[17199]_ ) & (~\m6_data_i[11]  | ~\new_[19561]_ );
  assign \new_[13734]_  = ~\new_[16427]_  & (~\new_[30541]_  | ~\new_[6203]_ );
  assign \new_[13735]_  = (~\m5_data_i[10]  | ~\new_[17199]_ ) & (~\m6_data_i[10]  | ~\new_[19561]_ );
  assign \new_[13736]_  = ~\new_[16431]_  & (~\new_[30420]_  | ~\new_[6041]_ );
  assign \new_[13737]_  = (~\m5_data_i[9]  | ~\new_[19544]_ ) & (~\m6_data_i[9]  | ~\new_[18789]_ );
  assign \new_[13738]_  = ~\new_[28356]_  & (~\new_[16739]_  | ~\new_[21455]_ );
  assign \new_[13739]_  = ~\new_[16433]_  & (~\new_[30648]_  | ~\new_[31143]_ );
  assign \new_[13740]_  = (~\m5_data_i[8]  | ~\new_[17199]_ ) & (~\m6_data_i[8]  | ~\new_[19561]_ );
  assign \new_[13741]_  = ~\new_[16434]_  & (~\new_[30336]_  | ~\new_[6199]_ );
  assign \new_[13742]_  = ~\new_[16436]_  & (~\new_[29926]_  | ~\new_[6200]_ );
  assign \new_[13743]_  = (~\m5_data_i[6]  | ~\new_[19544]_ ) & (~\m6_data_i[6]  | ~\new_[18789]_ );
  assign \new_[13744]_  = ~\new_[26598]_  & (~\new_[17293]_  | ~\new_[20478]_ );
  assign \new_[13745]_  = (~\m3_data_i[11]  | ~\new_[32350]_ ) & (~\m2_data_i[11]  | ~\new_[17224]_ );
  assign \new_[13746]_  = ~\new_[16438]_  & (~\new_[30038]_  | ~\new_[6208]_ );
  assign \new_[13747]_  = (~\m5_data_i[5]  | ~\new_[19544]_ ) & (~\m6_data_i[5]  | ~\new_[20551]_ );
  assign \new_[13748]_  = ~\new_[16441]_  & (~\new_[29828]_  | ~\new_[31406]_ );
  assign \new_[13749]_  = ~\new_[26645]_  & (~\new_[17417]_  | ~\new_[20499]_ );
  assign \new_[13750]_  = (~\m3_data_i[10]  | ~\new_[18936]_ ) & (~\m2_data_i[10]  | ~\new_[18808]_ );
  assign \new_[13751]_  = (~\m5_data_i[4]  | ~\new_[19544]_ ) & (~\m6_data_i[4]  | ~\new_[18789]_ );
  assign \new_[13752]_  = (~\m5_data_i[3]  | ~\new_[17200]_ ) & (~\m6_data_i[3]  | ~\new_[18789]_ );
  assign \new_[13753]_  = ~\new_[16446]_  & (~\new_[30029]_  | ~\new_[6211]_ );
  assign \new_[13754]_  = (~\m5_data_i[2]  | ~\new_[17200]_ ) & (~\m6_data_i[2]  | ~\new_[18789]_ );
  assign \new_[13755]_  = ~\new_[16448]_  & (~\new_[30002]_  | ~\new_[6273]_ );
  assign \new_[13756]_  = (~\m5_data_i[1]  | ~\new_[19544]_ ) & (~\m6_data_i[1]  | ~\new_[18789]_ );
  assign \new_[13757]_  = ~\new_[16450]_  & (~\new_[30553]_  | ~\new_[6213]_ );
  assign \new_[13758]_  = (~\m5_data_i[0]  | ~\new_[19544]_ ) & (~\m6_data_i[0]  | ~\new_[18789]_ );
  assign \new_[13759]_  = (~\m5_sel_i[3]  | ~\new_[17187]_ ) & (~\m6_sel_i[3]  | ~\new_[18050]_ );
  assign \new_[13760]_  = (~\m5_addr_i[21]  | ~\new_[17187]_ ) & (~\m6_addr_i[21]  | ~\new_[18049]_ );
  assign \new_[13761]_  = ~\new_[16452]_  & (~\new_[29790]_  | ~\new_[6214]_ );
  assign \new_[13762]_  = ~\new_[29407]_  & (~\new_[17309]_  | ~\new_[20470]_ );
  assign \new_[13763]_  = (~\new_[20551]_  | ~\m6_addr_i[30] ) & (~\new_[17201]_  | ~\new_[31147]_ );
  assign \new_[13764]_  = (~\new_[19561]_  | ~\m6_addr_i[29] ) & (~\new_[17200]_  | ~\new_[31407]_ );
  assign \new_[13765]_  = ~\new_[16456]_  & (~\new_[30466]_  | ~\new_[6268]_ );
  assign \new_[13766]_  = (~\new_[19561]_  | ~\m6_addr_i[27] ) & (~\new_[17200]_  | ~\m5_addr_i[27] );
  assign \new_[13767]_  = ~\new_[28257]_  & (~\new_[17412]_  | ~\new_[22693]_ );
  assign \new_[13768]_  = (~\new_[19561]_  | ~\m6_addr_i[25] ) & (~\new_[17200]_  | ~\m5_addr_i[25] );
  assign \new_[13769]_  = ~\new_[29297]_  & (~\new_[17365]_  | ~\new_[22948]_ );
  assign \new_[13770]_  = (~\new_[20551]_  | ~\m6_addr_i[24] ) & (~\new_[17201]_  | ~\m5_addr_i[24] );
  assign \new_[13771]_  = (~\m5_addr_i[23]  | ~\new_[17199]_ ) & (~\m6_addr_i[23]  | ~\new_[19561]_ );
  assign \new_[13772]_  = (~\m4_addr_i[23]  | ~\new_[18156]_ ) & (~\m3_addr_i[23]  | ~\new_[18130]_ );
  assign \new_[13773]_  = (~\m5_addr_i[21]  | ~\new_[17199]_ ) & (~\m6_addr_i[21]  | ~\new_[20551]_ );
  assign \new_[13774]_  = (~\m5_addr_i[20]  | ~\new_[17199]_ ) & (~\m6_addr_i[20]  | ~\new_[20551]_ );
  assign \new_[13775]_  = ~\new_[22151]_  & (~\new_[17033]_  | ~\new_[30550]_ );
  assign \new_[13776]_  = ~\new_[21565]_  & (~\new_[17036]_  | ~\new_[30410]_ );
  assign \new_[13777]_  = (~\m5_addr_i[19]  | ~\new_[17201]_ ) & (~\m6_addr_i[19]  | ~\new_[20551]_ );
  assign \new_[13778]_  = ~\new_[22131]_  & (~\new_[17042]_  | ~\new_[29212]_ );
  assign \new_[13779]_  = (~\m5_addr_i[18]  | ~\new_[17199]_ ) & (~\m6_addr_i[18]  | ~\new_[18789]_ );
  assign \new_[13780]_  = (~\m4_addr_i[18]  | ~\new_[18156]_ ) & (~\m3_addr_i[18]  | ~\new_[18130]_ );
  assign \new_[13781]_  = ~\new_[24301]_  & (~\new_[17049]_  | ~\new_[28967]_ );
  assign \new_[13782]_  = (~\m5_addr_i[17]  | ~\new_[17199]_ ) & (~\m6_addr_i[17]  | ~\new_[18789]_ );
  assign \new_[13783]_  = (~\m3_data_i[4]  | ~\new_[18936]_ ) & (~\m2_data_i[4]  | ~\new_[17224]_ );
  assign \new_[13784]_  = ~\new_[23633]_  & (~\new_[17029]_  | ~\new_[30107]_ );
  assign \new_[13785]_  = (~\m5_addr_i[16]  | ~\new_[17201]_ ) & (~\m6_addr_i[16]  | ~\new_[20551]_ );
  assign \new_[13786]_  = (~\m5_addr_i[15]  | ~\new_[17199]_ ) & (~\m6_addr_i[15]  | ~\new_[18789]_ );
  assign \new_[13787]_  = ~\new_[23817]_  & (~\new_[17077]_  | ~\new_[29972]_ );
  assign \new_[13788]_  = ~\new_[22269]_  & (~\new_[17067]_  | ~\new_[29040]_ );
  assign \new_[13789]_  = (~\m5_addr_i[14]  | ~\new_[17200]_ ) & (~\m6_addr_i[14]  | ~\new_[20551]_ );
  assign \new_[13790]_  = ~\new_[23573]_  & (~\new_[17048]_  | ~\new_[30723]_ );
  assign \new_[13791]_  = (~\m4_addr_i[13]  | ~\new_[18156]_ ) & (~\m3_addr_i[13]  | ~\new_[18130]_ );
  assign \new_[13792]_  = (~\m5_addr_i[13]  | ~\new_[17200]_ ) & (~\m6_addr_i[13]  | ~\new_[18789]_ );
  assign \new_[13793]_  = ~\new_[30152]_  | ~\new_[16639]_  | ~\new_[29794]_ ;
  assign \new_[13794]_  = (~\m5_addr_i[12]  | ~\new_[17199]_ ) & (~\m6_addr_i[12]  | ~\new_[18789]_ );
  assign \new_[13795]_  = ~\new_[16614]_  & ~\new_[16020]_ ;
  assign \new_[13796]_  = (~\m4_addr_i[22]  | ~\new_[17260]_ ) & (~\m3_addr_i[22]  | ~\new_[18175]_ );
  assign \new_[13797]_  = ~\new_[16642]_  & ~\new_[21267]_ ;
  assign \new_[13798]_  = (~\m5_addr_i[11]  | ~\new_[17199]_ ) & (~\m6_addr_i[11]  | ~\new_[18789]_ );
  assign \new_[13799]_  = (~\m4_addr_i[11]  | ~\new_[18156]_ ) & (~\m3_addr_i[11]  | ~\new_[18130]_ );
  assign \new_[13800]_  = (~\m3_data_i[2]  | ~\new_[32350]_ ) & (~\m2_data_i[2]  | ~\new_[18808]_ );
  assign \new_[13801]_  = ~\new_[16643]_  & ~\new_[21301]_ ;
  assign \new_[13802]_  = ~\new_[16646]_  & ~\new_[21270]_ ;
  assign \new_[13803]_  = (~\m5_addr_i[7]  | ~\new_[17200]_ ) & (~\m6_addr_i[7]  | ~\new_[20551]_ );
  assign \new_[13804]_  = ~\new_[29762]_  | ~\new_[16647]_  | ~\new_[28835]_ ;
  assign \new_[13805]_  = ~\new_[16160]_  & ~\new_[29058]_ ;
  assign \new_[13806]_  = ~\new_[16648]_  & ~\new_[21324]_ ;
  assign \new_[13807]_  = (~\m5_addr_i[6]  | ~\new_[17199]_ ) & (~\m6_addr_i[6]  | ~\new_[19561]_ );
  assign \new_[13808]_  = ~\new_[30011]_  | ~\new_[16649]_  | ~\new_[30160]_ ;
  assign \new_[13809]_  = ~\new_[29984]_  | ~\new_[16656]_  | ~\new_[30409]_ ;
  assign \new_[13810]_  = ~\new_[16599]_  & ~\new_[30130]_ ;
  assign \new_[13811]_  = (~\m5_addr_i[5]  | ~\new_[17199]_ ) & (~\m6_addr_i[5]  | ~\new_[19561]_ );
  assign \new_[13812]_  = ~\new_[21592]_  & (~\new_[16868]_  | ~\new_[29831]_ );
  assign \new_[13813]_  = (~\m5_addr_i[4]  | ~\new_[17199]_ ) & (~\m6_addr_i[4]  | ~\new_[18789]_ );
  assign \new_[13814]_  = ~\new_[16660]_  & ~\new_[23947]_ ;
  assign \new_[13815]_  = ~\new_[30717]_  | ~\new_[16661]_  | ~\new_[30349]_ ;
  assign \new_[13816]_  = (~\m5_addr_i[3]  | ~\new_[19544]_ ) & (~\m6_addr_i[3]  | ~\new_[20551]_ );
  assign \new_[13817]_  = (~\new_[17227]_  | ~\m6_addr_i[31] ) & (~\new_[18745]_  | ~\new_[31001]_ );
  assign \new_[13818]_  = ~\new_[16662]_  & ~\new_[23914]_ ;
  assign \new_[13819]_  = ~\new_[30213]_  | ~\new_[16663]_  | ~\new_[29877]_ ;
  assign \new_[13820]_  = ~\new_[30092]_  | ~\new_[16667]_  | ~\new_[28911]_ ;
  assign \new_[13821]_  = ~\new_[16371]_  & ~\new_[29254]_ ;
  assign \new_[13822]_  = ~\new_[16668]_  & ~\new_[21294]_ ;
  assign \new_[13823]_  = ~\new_[28888]_  | ~\new_[16669]_  | ~\new_[30178]_ ;
  assign \new_[13824]_  = (~\m5_addr_i[0]  | ~\new_[17199]_ ) & (~\m6_addr_i[0]  | ~\new_[19561]_ );
  assign \new_[13825]_  = ~\new_[16357]_  & ~\new_[29115]_ ;
  assign \new_[13826]_  = (~\m4_sel_i[3]  | ~\new_[18156]_ ) & (~\m3_sel_i[3]  | ~\new_[18130]_ );
  assign \new_[13827]_  = ~\new_[16670]_  & ~\new_[21276]_ ;
  assign \new_[13828]_  = (~\new_[17227]_  | ~\m6_addr_i[29] ) & (~\new_[18745]_  | ~\new_[31407]_ );
  assign \new_[13829]_  = (~\m5_sel_i[2]  | ~\new_[17199]_ ) & (~\m6_sel_i[2]  | ~\new_[18789]_ );
  assign \new_[13830]_  = ~\new_[16674]_  & ~\new_[20561]_ ;
  assign \new_[13831]_  = (~\m5_sel_i[1]  | ~\new_[17199]_ ) & (~\m6_sel_i[1]  | ~\new_[18789]_ );
  assign \new_[13832]_  = ~\new_[15925]_  & ~\new_[29229]_ ;
  assign \new_[13833]_  = (~\m5_sel_i[0]  | ~\new_[17199]_ ) & (~\m6_sel_i[0]  | ~\new_[18789]_ );
  assign \new_[13834]_  = ~\new_[16675]_  & ~\new_[21315]_ ;
  assign \new_[13835]_  = ~\new_[21480]_  & (~\new_[16924]_  | ~\new_[30751]_ );
  assign \new_[13836]_  = (~\new_[19581]_  | ~\m6_addr_i[28] ) & (~\new_[18745]_  | ~\new_[31276]_ );
  assign \new_[13837]_  = ~\new_[16676]_  & ~\new_[23920]_ ;
  assign \new_[13838]_  = (~m5_we_i | ~\new_[19544]_ ) & (~m6_we_i | ~\new_[20551]_ );
  assign \new_[13839]_  = (~\new_[17227]_  | ~\m6_addr_i[27] ) & (~\new_[17202]_  | ~\m5_addr_i[27] );
  assign \new_[13840]_  = (~\new_[17227]_  | ~\m6_addr_i[26] ) & (~\new_[18745]_  | ~\m5_addr_i[26] );
  assign \new_[13841]_  = ~\new_[16681]_  & ~\new_[21314]_ ;
  assign \new_[13842]_  = ~\new_[28001]_  | ~\new_[16682]_  | ~\new_[30089]_ ;
  assign \new_[13843]_  = (~\new_[17227]_  | ~\m6_addr_i[25] ) & (~\new_[18745]_  | ~\m5_addr_i[25] );
  assign \new_[13844]_  = ~\new_[23050]_  & (~\new_[16932]_  | ~\new_[29571]_ );
  assign \new_[13845]_  = (~\m4_data_i[31]  | ~\new_[18149]_ ) & (~\m3_data_i[31]  | ~\new_[18930]_ );
  assign \new_[13846]_  = ~\new_[22367]_  & (~\new_[17251]_  | ~\new_[28887]_ );
  assign \new_[13847]_  = ~\new_[16686]_  & ~\new_[23905]_ ;
  assign \new_[13848]_  = (~\new_[17227]_  | ~\m6_addr_i[24] ) & (~\new_[18745]_  | ~\m5_addr_i[24] );
  assign \new_[13849]_  = (~\m5_data_i[7]  | ~\new_[17200]_ ) & (~\m6_data_i[7]  | ~\new_[18789]_ );
  assign \new_[13850]_  = ~\new_[15913]_  & ~\new_[23951]_ ;
  assign \new_[13851]_  = ~\new_[29798]_  | ~\new_[15914]_  | ~\new_[29897]_ ;
  assign \new_[13852]_  = ~\new_[24794]_  & (~\new_[16789]_  | ~\new_[30150]_ );
  assign \new_[13853]_  = ~\new_[22409]_  & (~\new_[16795]_  | ~\new_[23064]_ );
  assign \new_[13854]_  = \new_[15941]_  | \new_[24008]_ ;
  assign \new_[13855]_  = ~\new_[23355]_  & (~\new_[16798]_  | ~\new_[30020]_ );
  assign \new_[13856]_  = ~\new_[22124]_  & (~\new_[16807]_  | ~\new_[30337]_ );
  assign \new_[13857]_  = ~\new_[15143]_ ;
  assign \new_[13858]_  = ~\new_[15144]_ ;
  assign \new_[13859]_  = (~\m3_addr_i[22]  | ~\new_[32350]_ ) & (~\m2_addr_i[22]  | ~\new_[18808]_ );
  assign \new_[13860]_  = \new_[15942]_  | \new_[25439]_ ;
  assign \new_[13861]_  = ~\new_[27692]_  & (~\new_[16810]_  | ~\new_[23088]_ );
  assign \new_[13862]_  = ~\new_[24387]_  & (~\new_[16811]_  | ~\new_[24467]_ );
  assign \new_[13863]_  = ~\new_[21136]_  & (~\new_[16812]_  | ~\new_[30232]_ );
  assign \new_[13864]_  = ~\new_[16555]_  & ~\new_[23404]_ ;
  assign \new_[13865]_  = ~\new_[26893]_  & (~\new_[16824]_  | ~\new_[29975]_ );
  assign \new_[13866]_  = ~\new_[22694]_  & (~\new_[16826]_  | ~\new_[26274]_ );
  assign \new_[13867]_  = ~\new_[15150]_ ;
  assign \new_[13868]_  = \new_[15945]_  | \new_[24761]_ ;
  assign \new_[13869]_  = ~\new_[15153]_ ;
  assign \new_[13870]_  = ~\new_[15154]_ ;
  assign \new_[13871]_  = ~\new_[22149]_  & (~\new_[16831]_  | ~\new_[30665]_ );
  assign \new_[13872]_  = (~\m4_data_i[18]  | ~\new_[18149]_ ) & (~\m3_data_i[18]  | ~\new_[18930]_ );
  assign \new_[13873]_  = (~\m4_data_i[17]  | ~\new_[18149]_ ) & (~\m3_data_i[17]  | ~\new_[18930]_ );
  assign \new_[13874]_  = ~\new_[24869]_  & (~\new_[16839]_  | ~\new_[30505]_ );
  assign \new_[13875]_  = ~\new_[23062]_  & (~\new_[16841]_  | ~\new_[22899]_ );
  assign \new_[13876]_  = ~\new_[15158]_ ;
  assign \new_[13877]_  = \new_[15947]_  | \new_[23162]_ ;
  assign \new_[13878]_  = ~\new_[15161]_ ;
  assign \new_[13879]_  = ~\new_[23458]_  & (~\new_[16842]_  | ~\new_[30255]_ );
  assign \new_[13880]_  = (~\m4_data_i[15]  | ~\new_[18149]_ ) & (~\m3_data_i[15]  | ~\new_[18928]_ );
  assign \new_[13881]_  = ~\new_[16559]_  & ~\new_[24892]_ ;
  assign \new_[13882]_  = (~\m4_data_i[14]  | ~\new_[18149]_ ) & (~\m3_data_i[14]  | ~\new_[18930]_ );
  assign \new_[13883]_  = (~\m3_addr_i[19]  | ~\new_[32350]_ ) & (~\m2_addr_i[19]  | ~\new_[18808]_ );
  assign \new_[13884]_  = ~\new_[21921]_  & (~\new_[16848]_  | ~\new_[23084]_ );
  assign \new_[13885]_  = ~\new_[19445]_  & (~\new_[16849]_  | ~\new_[26726]_ );
  assign \new_[13886]_  = ~\new_[22264]_  & (~\new_[16850]_  | ~\new_[29150]_ );
  assign \new_[13887]_  = (~\m4_data_i[13]  | ~\new_[18149]_ ) & (~\m3_data_i[13]  | ~\new_[18930]_ );
  assign \new_[13888]_  = \new_[15948]_  | \new_[26405]_ ;
  assign \new_[13889]_  = ~\new_[15167]_ ;
  assign \new_[13890]_  = ~\new_[15168]_ ;
  assign \new_[13891]_  = ~\new_[23485]_  & (~\new_[16853]_  | ~\new_[29782]_ );
  assign \new_[13892]_  = (~\m3_addr_i[18]  | ~\new_[32350]_ ) & (~\m2_addr_i[18]  | ~\new_[18808]_ );
  assign \new_[13893]_  = ~\new_[15173]_ ;
  assign \new_[13894]_  = (~\m4_data_i[11]  | ~\new_[18149]_ ) & (~\m3_data_i[11]  | ~\new_[18928]_ );
  assign \new_[13895]_  = ~\new_[21592]_  & (~\new_[16869]_  | ~\new_[25129]_ );
  assign \new_[13896]_  = ~\new_[22226]_  & (~\new_[16870]_  | ~\new_[30217]_ );
  assign \new_[13897]_  = ~\new_[23183]_  & (~\new_[16876]_  | ~\new_[27706]_ );
  assign \new_[13898]_  = ~\new_[23527]_  & (~\new_[16884]_  | ~\new_[29441]_ );
  assign \new_[13899]_  = (~\m4_data_i[9]  | ~\new_[18149]_ ) & (~\m3_data_i[9]  | ~\new_[18930]_ );
  assign \new_[13900]_  = ~\new_[16571]_  & ~\new_[26969]_ ;
  assign \new_[13901]_  = ~\new_[15178]_ ;
  assign \new_[13902]_  = ~\new_[15179]_ ;
  assign \new_[13903]_  = ~\new_[23544]_  & (~\new_[16944]_  | ~\new_[28870]_ );
  assign \new_[13904]_  = (~\m4_data_i[8]  | ~\new_[18149]_ ) & (~\m3_data_i[8]  | ~\new_[18930]_ );
  assign \new_[13905]_  = \new_[15953]_  | \new_[25127]_ ;
  assign \new_[13906]_  = ~\new_[15181]_ ;
  assign \new_[13907]_  = ~\new_[15182]_ ;
  assign \new_[13908]_  = (~\m4_data_i[7]  | ~\new_[18149]_ ) & (~\m3_data_i[7]  | ~\new_[18930]_ );
  assign \new_[13909]_  = ~\new_[23567]_  & (~\new_[16895]_  | ~\new_[28828]_ );
  assign \new_[13910]_  = (~\m4_data_i[6]  | ~\new_[18149]_ ) & (~\m3_data_i[6]  | ~\new_[18928]_ );
  assign \new_[13911]_  = ~\new_[22210]_  & (~\new_[16873]_  | ~\new_[22137]_ );
  assign \new_[13912]_  = ~\new_[15187]_ ;
  assign \new_[13913]_  = \new_[15955]_  | \new_[24511]_ ;
  assign \new_[13914]_  = ~\new_[15188]_ ;
  assign \new_[13915]_  = ~\new_[15190]_ ;
  assign \new_[13916]_  = ~\new_[22263]_  & (~\new_[16898]_  | ~\new_[30636]_ );
  assign \new_[13917]_  = ~\new_[16578]_  & ~\new_[23778]_ ;
  assign \new_[13918]_  = ~\new_[25102]_  & (~\new_[16904]_  | ~\new_[29867]_ );
  assign \new_[13919]_  = ~\new_[22942]_  & (~\new_[16905]_  | ~\new_[25660]_ );
  assign \new_[13920]_  = ~\new_[15196]_ ;
  assign \new_[13921]_  = \new_[15956]_  | \new_[26561]_ ;
  assign \new_[13922]_  = (~\m3_addr_i[15]  | ~\new_[32350]_ ) & (~\m2_addr_i[15]  | ~\new_[18808]_ );
  assign \new_[13923]_  = ~\new_[23182]_  & (~\new_[16900]_  | ~\new_[27953]_ );
  assign \new_[13924]_  = ~\new_[23615]_  & (~\new_[16908]_  | ~\new_[30595]_ );
  assign \new_[13925]_  = (~\m4_data_i[1]  | ~\new_[18149]_ ) & (~\m3_data_i[1]  | ~\new_[18928]_ );
  assign \new_[13926]_  = ~\new_[16583]_  & ~\new_[26853]_ ;
  assign \new_[13927]_  = ~\new_[21556]_  & (~\new_[16913]_  | ~\new_[26169]_ );
  assign \new_[13928]_  = ~\new_[15205]_ ;
  assign \new_[13929]_  = (~\new_[18149]_  | ~\m4_addr_i[31] ) & (~\new_[18930]_  | ~\m3_addr_i[31] );
  assign \new_[13930]_  = (~\new_[18149]_  | ~\m4_addr_i[30] ) & (~\new_[18930]_  | ~\m3_addr_i[30] );
  assign \new_[13931]_  = ~\new_[23631]_  & (~\new_[16797]_  | ~\new_[30600]_ );
  assign \new_[13932]_  = ~\new_[23647]_  & (~\new_[16823]_  | ~\new_[30321]_ );
  assign \new_[13933]_  = ~\new_[15214]_ ;
  assign \new_[13934]_  = ~\new_[15215]_ ;
  assign \new_[13935]_  = ~\new_[24746]_  & (~\new_[16911]_  | ~\new_[24348]_ );
  assign \new_[13936]_  = ~\new_[15218]_ ;
  assign \new_[13937]_  = ~\new_[22314]_  & (~\new_[16917]_  | ~\new_[29912]_ );
  assign \new_[13938]_  = (~\new_[18149]_  | ~\m4_addr_i[27] ) & (~\new_[18929]_  | ~\m3_addr_i[27] );
  assign \new_[13939]_  = (~\new_[19563]_  | ~\m6_addr_i[24] ) & (~\new_[18735]_  | ~\m5_addr_i[24] );
  assign \new_[13940]_  = ~\new_[16591]_  & ~\new_[22363]_ ;
  assign \new_[13941]_  = ~\new_[25025]_  & (~\new_[16923]_  | ~\new_[29979]_ );
  assign \new_[13942]_  = ~\new_[15222]_ ;
  assign \new_[13943]_  = ~\new_[15224]_ ;
  assign \new_[13944]_  = (~\new_[18149]_  | ~\m4_addr_i[26] ) & (~\new_[18929]_  | ~\m3_addr_i[26] );
  assign \new_[13945]_  = \new_[15958]_  | \new_[23924]_ ;
  assign \new_[13946]_  = (~\new_[18149]_  | ~\m4_addr_i[25] ) & (~\new_[18930]_  | ~\m3_addr_i[25] );
  assign \new_[13947]_  = ~\new_[21480]_  & (~\new_[16886]_  | ~\new_[26744]_ );
  assign \new_[13948]_  = ~\new_[23837]_  & (~\new_[16967]_  | ~\new_[30702]_ );
  assign \new_[13949]_  = \new_[15959]_  | \new_[25065]_ ;
  assign \new_[13950]_  = ~\new_[26488]_  & (~\new_[16968]_  | ~\new_[30009]_ );
  assign \new_[13951]_  = ~\new_[15229]_ ;
  assign \new_[13952]_  = ~\new_[15230]_ ;
  assign \new_[13953]_  = (~\m4_addr_i[23]  | ~\new_[18149]_ ) & (~\m3_addr_i[23]  | ~\new_[18928]_ );
  assign \new_[13954]_  = \new_[15960]_  | \new_[26829]_ ;
  assign \new_[13955]_  = (~\m4_addr_i[22]  | ~\new_[18149]_ ) & (~\m3_addr_i[22]  | ~\new_[18930]_ );
  assign \new_[13956]_  = (~\m3_addr_i[11]  | ~\new_[32350]_ ) & (~\m2_addr_i[11]  | ~\new_[17224]_ );
  assign \new_[13957]_  = ~\new_[23384]_  & (~\new_[16966]_  | ~\new_[30142]_ );
  assign \new_[13958]_  = ~\new_[15240]_ ;
  assign \new_[13959]_  = ~\new_[23050]_  & (~\new_[16959]_  | ~\new_[27909]_ );
  assign \new_[13960]_  = ~\new_[23726]_  & (~\new_[16938]_  | ~\new_[29685]_ );
  assign \new_[13961]_  = ~\new_[24345]_  & (~\new_[16935]_  | ~\new_[23059]_ );
  assign \new_[13962]_  = (~\m4_addr_i[20]  | ~\new_[18149]_ ) & (~\m3_addr_i[20]  | ~\new_[18930]_ );
  assign \new_[13963]_  = (~\m3_addr_i[10]  | ~\new_[32350]_ ) & (~\m2_addr_i[10]  | ~\new_[17224]_ );
  assign \new_[13964]_  = ~\new_[23761]_  & (~\new_[16936]_  | ~\new_[28898]_ );
  assign \new_[13965]_  = ~\new_[15246]_ ;
  assign \new_[13966]_  = ~\new_[15247]_ ;
  assign \new_[13967]_  = \new_[15962]_  | \new_[24337]_ ;
  assign \new_[13968]_  = ~\new_[15249]_ ;
  assign \new_[13969]_  = ~\new_[23748]_  & (~\new_[16814]_  | ~\new_[29927]_ );
  assign \new_[13970]_  = ~\new_[23843]_  & (~\new_[16974]_  | ~\new_[29226]_ );
  assign \new_[13971]_  = ~\new_[16609]_  & ~\new_[25138]_ ;
  assign \new_[13972]_  = ~\new_[15253]_ ;
  assign \new_[13973]_  = ~\new_[15255]_ ;
  assign \new_[13974]_  = (~\m4_addr_i[15]  | ~\new_[18149]_ ) & (~\m3_addr_i[15]  | ~\new_[18930]_ );
  assign \new_[13975]_  = \new_[15965]_  | \new_[26752]_ ;
  assign \new_[13976]_  = ~\new_[23164]_  & (~\new_[16979]_  | ~\new_[29118]_ );
  assign \new_[13977]_  = ~\new_[16622]_  | ~\new_[22873]_ ;
  assign \new_[13978]_  = ~\new_[27750]_  & (~\new_[16794]_  | ~\new_[29028]_ );
  assign \new_[13979]_  = (~\m4_addr_i[11]  | ~\new_[18149]_ ) & (~\m3_addr_i[11]  | ~\new_[18930]_ );
  assign \new_[13980]_  = (~\m3_addr_i[7]  | ~\new_[32350]_ ) & (~\m2_addr_i[7]  | ~\new_[18808]_ );
  assign \new_[13981]_  = (~\m4_addr_i[9]  | ~\new_[18149]_ ) & (~\m3_addr_i[9]  | ~\new_[18930]_ );
  assign \new_[13982]_  = ~\new_[28189]_  & (~\new_[16808]_  | ~\new_[20500]_ );
  assign \new_[13983]_  = (~\m4_addr_i[7]  | ~\new_[18149]_ ) & (~\m3_addr_i[7]  | ~\new_[18930]_ );
  assign \new_[13984]_  = (~\m3_addr_i[6]  | ~\new_[32350]_ ) & (~\m2_addr_i[6]  | ~\new_[18808]_ );
  assign \new_[13985]_  = (~\m4_addr_i[6]  | ~\new_[18149]_ ) & (~\m3_addr_i[6]  | ~\new_[18930]_ );
  assign \new_[13986]_  = (~\m4_addr_i[5]  | ~\new_[18149]_ ) & (~\m3_addr_i[5]  | ~\new_[18930]_ );
  assign \new_[13987]_  = ~\new_[29218]_  & (~\new_[16825]_  | ~\new_[21466]_ );
  assign \new_[13988]_  = (~\m4_addr_i[2]  | ~\new_[18149]_ ) & (~\m3_addr_i[2]  | ~\new_[18930]_ );
  assign \new_[13989]_  = ~\new_[16623]_  | ~\new_[22927]_ ;
  assign \new_[13990]_  = ~\new_[16615]_  & (~\new_[29930]_  | ~\new_[5970]_ );
  assign \new_[13991]_  = ~\new_[23062]_  & (~\new_[16840]_  | ~\new_[28050]_ );
  assign \new_[13992]_  = (~\m4_sel_i[2]  | ~\new_[18149]_ ) & (~\m3_sel_i[2]  | ~\new_[18928]_ );
  assign \new_[13993]_  = ~\new_[16624]_  | ~\new_[22995]_ ;
  assign \new_[13994]_  = ~\new_[16625]_  | ~\new_[24317]_ ;
  assign \new_[13995]_  = ~\new_[16616]_  & (~\new_[30093]_  | ~\new_[6050]_ );
  assign \new_[13996]_  = ~\new_[23121]_  | ~\new_[24356]_  | ~\new_[16781]_ ;
  assign \new_[13997]_  = ~\new_[28995]_  & (~\new_[16855]_  | ~\new_[21396]_ );
  assign \new_[13998]_  = (~m4_we_i | ~\new_[18149]_ ) & (~m3_we_i | ~\new_[18930]_ );
  assign \new_[13999]_  = (~\m3_addr_i[2]  | ~\new_[18936]_ ) & (~\m2_addr_i[2]  | ~\new_[17224]_ );
  assign \new_[14000]_  = ~\new_[28754]_  & (~\new_[16865]_  | ~\new_[20469]_ );
  assign \new_[14001]_  = ~\new_[26382]_  & (~\new_[16866]_  | ~\new_[29593]_ );
  assign \new_[14002]_  = ~\new_[23173]_  & (~\new_[16867]_  | ~\new_[29868]_ );
  assign \new_[14003]_  = ~\new_[26275]_  | ~\new_[26359]_  | ~\new_[16783]_ ;
  assign \new_[14004]_  = ~\new_[26643]_  & (~\new_[16874]_  | ~\new_[21424]_ );
  assign \new_[14005]_  = ~\new_[26447]_  & (~\new_[16792]_  | ~\new_[21358]_ );
  assign \new_[14006]_  = ~\new_[16628]_  | ~\new_[20449]_ ;
  assign \new_[14007]_  = (~\m3_addr_i[0]  | ~\new_[32350]_ ) & (~\m2_addr_i[0]  | ~\new_[17224]_ );
  assign \new_[14008]_  = ~\new_[16629]_  | ~\new_[24268]_ ;
  assign \new_[14009]_  = ~\new_[16617]_  & (~\new_[30199]_  | ~\new_[6057]_ );
  assign \new_[14010]_  = ~\new_[28303]_  & (~\new_[16887]_  | ~\new_[20445]_ );
  assign \new_[14011]_  = ~\new_[26583]_  & (~\new_[16889]_  | ~\new_[22536]_ );
  assign \new_[14012]_  = ~\new_[16630]_  | ~\new_[20446]_ ;
  assign \new_[14013]_  = (~\m2_data_i[25]  | ~\new_[18068]_ ) & (~\m1_data_i[25]  | ~\new_[18901]_ );
  assign \new_[14014]_  = ~\new_[16632]_  | ~\new_[21560]_ ;
  assign \new_[14015]_  = ~\new_[29986]_  & (~\new_[16896]_  | ~\new_[21494]_ );
  assign \new_[14016]_  = (~\m2_data_i[24]  | ~\new_[18067]_ ) & (~\m1_data_i[24]  | ~\new_[19626]_ );
  assign \new_[14017]_  = (~\m3_sel_i[2]  | ~\new_[32350]_ ) & (~\m2_sel_i[2]  | ~\new_[18808]_ );
  assign \new_[14018]_  = ~\new_[29154]_  & (~\new_[16804]_  | ~\new_[22274]_ );
  assign \new_[14019]_  = ~\new_[16633]_  | ~\new_[24451]_ ;
  assign \new_[14020]_  = ~\new_[16618]_  & (~\new_[30010]_  | ~\new_[5984]_ );
  assign \new_[14021]_  = (~\m2_data_i[21]  | ~\new_[18067]_ ) & (~\m1_data_i[21]  | ~\new_[19625]_ );
  assign \new_[14022]_  = (~m5_we_i | ~\new_[18735]_ ) & (~m6_we_i | ~\new_[18051]_ );
  assign \new_[14023]_  = (~\m2_data_i[19]  | ~\new_[18068]_ ) & (~\m1_data_i[19]  | ~\new_[20573]_ );
  assign \new_[14024]_  = (~\m2_data_i[18]  | ~\new_[18069]_ ) & (~\m1_data_i[18]  | ~\new_[20573]_ );
  assign \new_[14025]_  = ~\new_[27984]_  & (~\new_[16877]_  | ~\new_[20424]_ );
  assign \new_[14026]_  = ~\new_[16634]_  | ~\new_[22966]_ ;
  assign \new_[14027]_  = (~\m2_data_i[17]  | ~\new_[18069]_ ) & (~\m1_data_i[17]  | ~\new_[19625]_ );
  assign \new_[14028]_  = ~\new_[16619]_  & (~\new_[30066]_  | ~\new_[6070]_ );
  assign \new_[14029]_  = (~\m3_sel_i[0]  | ~\new_[32350]_ ) & (~\m2_sel_i[0]  | ~\new_[17224]_ );
  assign \new_[14030]_  = ~\new_[30238]_  & (~\new_[16828]_  | ~\new_[20455]_ );
  assign \new_[14031]_  = ~\new_[21556]_  & (~\new_[16912]_  | ~\new_[28073]_ );
  assign \new_[14032]_  = ~\new_[22982]_  | ~\new_[21584]_  | ~\new_[16784]_ ;
  assign \new_[14033]_  = ~\new_[22439]_  & (~\new_[17230]_  | ~\new_[28939]_ );
  assign \new_[14034]_  = (~m3_we_i | ~\new_[32350]_ ) & (~m2_we_i | ~\new_[17224]_ );
  assign \new_[14035]_  = ~\new_[29932]_  & (~\new_[16977]_  | ~\new_[20700]_ );
  assign \new_[14036]_  = (~\m2_data_i[13]  | ~\new_[18068]_ ) & (~\m1_data_i[13]  | ~\new_[20573]_ );
  assign \new_[14037]_  = (~\m2_data_i[12]  | ~\new_[18069]_ ) & (~\m1_data_i[12]  | ~\new_[19625]_ );
  assign \new_[14038]_  = (~\m2_data_i[10]  | ~\new_[18069]_ ) & (~\m1_data_i[10]  | ~\new_[19625]_ );
  assign \new_[14039]_  = ~\new_[16635]_  | ~\new_[20506]_ ;
  assign \new_[14040]_  = ~\new_[16620]_  & (~\new_[30075]_  | ~\new_[5925]_ );
  assign \new_[14041]_  = (~\m2_data_i[7]  | ~\new_[19567]_ ) & (~\m1_data_i[7]  | ~\new_[18899]_ );
  assign \new_[14042]_  = ~\new_[29414]_  & (~\new_[16817]_  | ~\new_[29851]_ );
  assign \new_[14043]_  = (~\m2_data_i[5]  | ~\new_[19567]_ ) & (~\m1_data_i[5]  | ~\new_[19626]_ );
  assign \new_[14044]_  = ~\new_[28443]_  & (~\new_[16927]_  | ~\new_[20510]_ );
  assign \new_[14045]_  = (~\m2_data_i[3]  | ~\new_[18069]_ ) & (~\m1_data_i[3]  | ~\new_[19625]_ );
  assign \new_[14046]_  = ~\new_[26779]_  & (~\new_[16928]_  | ~\new_[29583]_ );
  assign \new_[14047]_  = (~\m2_data_i[2]  | ~\new_[18068]_ ) & (~\m1_data_i[2]  | ~\new_[18901]_ );
  assign \new_[14048]_  = (~\m7_data_i[31]  | ~\new_[18823]_ ) & (~\m0_data_i[31]  | ~\new_[20539]_ );
  assign \new_[14049]_  = (~\m2_data_i[1]  | ~\new_[18069]_ ) & (~\m1_data_i[1]  | ~\new_[19625]_ );
  assign \new_[14050]_  = (~\m2_data_i[31]  | ~\new_[18799]_ ) & (~\m1_data_i[31]  | ~\new_[18887]_ );
  assign \new_[14051]_  = ~\new_[28804]_  & (~\new_[16965]_  | ~\new_[20481]_ );
  assign \new_[14052]_  = ~\new_[26721]_  & (~\new_[16960]_  | ~\new_[28675]_ );
  assign \new_[14053]_  = (~\new_[19567]_  | ~\new_[31537]_ ) & (~\new_[19626]_  | ~\m1_addr_i[31] );
  assign \new_[14054]_  = (~\new_[19567]_  | ~\new_[31486]_ ) & (~\new_[19626]_  | ~\new_[31308]_ );
  assign \new_[14055]_  = (~\m2_data_i[29]  | ~\new_[18799]_ ) & (~\m1_data_i[29]  | ~\new_[18887]_ );
  assign \new_[14056]_  = ~\new_[16631]_  | ~\new_[19444]_ ;
  assign \new_[14057]_  = ~\new_[30122]_  & (~\new_[16800]_  | ~\new_[24457]_ );
  assign \new_[14058]_  = ~\new_[23056]_  & (~\new_[16939]_  | ~\new_[30117]_ );
  assign \new_[14059]_  = (~\m2_data_i[28]  | ~\new_[18799]_ ) & (~\m1_data_i[28]  | ~\new_[20571]_ );
  assign \new_[14060]_  = ~\new_[26817]_  & (~\new_[16888]_  | ~\new_[29421]_ );
  assign \new_[14061]_  = ~\new_[23118]_  | ~\new_[23122]_  | ~\new_[16780]_ ;
  assign \new_[14062]_  = (~\m7_data_i[28]  | ~\new_[17236]_ ) & (~\m0_data_i[28]  | ~\new_[20539]_ );
  assign \new_[14063]_  = (~\new_[19567]_  | ~\m2_addr_i[26] ) & (~\new_[19626]_  | ~\m1_addr_i[26] );
  assign \new_[14064]_  = ~\new_[28697]_  & (~\new_[16941]_  | ~\new_[22812]_ );
  assign \new_[14065]_  = ~\new_[16636]_  | ~\new_[19447]_ ;
  assign \new_[14066]_  = ~\new_[16637]_  | ~\new_[22104]_ ;
  assign \new_[14067]_  = ~\new_[16638]_  | ~\new_[23124]_ ;
  assign \new_[14068]_  = ~\new_[16621]_  & (~\new_[30047]_  | ~\new_[6092]_ );
  assign \new_[14069]_  = (~\m7_data_i[26]  | ~\new_[17235]_ ) & (~\m0_data_i[26]  | ~\new_[19535]_ );
  assign \new_[14070]_  = (~\new_[19567]_  | ~\m2_addr_i[24] ) & (~\new_[19626]_  | ~\m1_addr_i[24] );
  assign \new_[14071]_  = ~\new_[23569]_  | ~\new_[23120]_  | ~\new_[16788]_ ;
  assign \new_[14072]_  = (~\m2_data_i[26]  | ~\new_[18799]_ ) & (~\m1_data_i[26]  | ~\new_[18887]_ );
  assign \new_[14073]_  = ~\new_[29009]_  & (~\new_[16978]_  | ~\new_[30233]_ );
  assign \new_[14074]_  = (~\m2_addr_i[22]  | ~\new_[18068]_ ) & (~\m1_addr_i[22]  | ~\new_[18898]_ );
  assign \new_[14075]_  = (~\m7_data_i[25]  | ~\new_[17236]_ ) & (~\m0_data_i[25]  | ~\new_[20539]_ );
  assign \new_[14076]_  = (~\m2_addr_i[20]  | ~\new_[18067]_ ) & (~\m1_addr_i[20]  | ~\new_[19626]_ );
  assign \new_[14077]_  = (~\m7_data_i[24]  | ~\new_[17235]_ ) & (~\m0_data_i[24]  | ~\new_[19535]_ );
  assign \new_[14078]_  = ~\new_[28607]_  & (~\new_[17047]_  | ~\new_[18428]_ );
  assign \new_[14079]_  = ~\new_[28087]_  & (~\new_[17058]_  | ~\new_[19428]_ );
  assign \new_[14080]_  = ~\new_[30165]_  & (~\new_[17111]_  | ~\new_[18420]_ );
  assign \new_[14081]_  = (~\m2_addr_i[17]  | ~\new_[18068]_ ) & (~\m1_addr_i[17]  | ~\new_[18898]_ );
  assign \new_[14082]_  = (~\new_[19567]_  | ~\new_[31547]_ ) & (~\new_[19626]_  | ~\new_[31458]_ );
  assign \new_[14083]_  = (~\m7_data_i[23]  | ~\new_[18823]_ ) & (~\m0_data_i[23]  | ~\new_[18731]_ );
  assign \new_[14084]_  = (~\m2_data_i[23]  | ~\new_[18799]_ ) & (~\m1_data_i[23]  | ~\new_[20571]_ );
  assign \new_[14085]_  = (~\m2_addr_i[16]  | ~\new_[18068]_ ) & (~\m1_addr_i[16]  | ~\new_[20573]_ );
  assign \new_[14086]_  = ~\new_[24276]_  & (~\new_[17140]_  | ~\new_[28183]_ );
  assign \new_[14087]_  = (~\m7_data_i[22]  | ~\new_[17235]_ ) & (~\m0_data_i[22]  | ~\new_[19535]_ );
  assign \new_[14088]_  = (~\m2_addr_i[15]  | ~\new_[18068]_ ) & (~\m1_addr_i[15]  | ~\new_[20573]_ );
  assign \new_[14089]_  = ~\new_[22969]_  | (~\new_[16821]_  & ~\new_[30633]_ );
  assign \new_[14090]_  = ~\new_[21782]_  | (~\new_[16836]_  & ~\new_[30253]_ );
  assign \new_[14091]_  = ~\new_[26636]_  & (~\new_[17144]_  | ~\new_[29762]_ );
  assign \new_[14092]_  = (~\m7_data_i[21]  | ~\new_[17236]_ ) & (~\m0_data_i[21]  | ~\new_[19537]_ );
  assign \new_[14093]_  = (~\m2_addr_i[12]  | ~\new_[18068]_ ) & (~\m1_addr_i[12]  | ~\new_[18898]_ );
  assign \new_[14094]_  = ~\new_[16568]_  | ~\new_[20449]_ ;
  assign \new_[14095]_  = (~\m2_addr_i[11]  | ~\new_[18068]_ ) & (~\m1_addr_i[11]  | ~\new_[19625]_ );
  assign \new_[14096]_  = ~\new_[16574]_  | ~\new_[20446]_ ;
  assign \new_[14097]_  = (~\m2_data_i[20]  | ~\new_[18799]_ ) & (~\m1_data_i[20]  | ~\new_[20571]_ );
  assign \new_[14098]_  = ~\new_[27752]_  & (~\new_[17149]_  | ~\new_[30092]_ );
  assign \new_[14099]_  = ~\new_[23055]_  | (~\new_[16949]_  & ~\new_[30350]_ );
  assign \new_[14100]_  = ~\new_[26913]_  & (~\new_[17151]_  | ~\new_[29888]_ );
  assign \new_[14101]_  = ~\new_[24298]_  | (~\new_[16940]_  & ~\new_[29238]_ );
  assign \new_[14102]_  = (~\m7_data_i[18]  | ~\new_[17236]_ ) & (~\m0_data_i[18]  | ~\new_[19537]_ );
  assign \new_[14103]_  = ~\new_[27664]_  & (~\new_[17152]_  | ~\new_[30061]_ );
  assign \new_[14104]_  = (~\m2_addr_i[4]  | ~\new_[19567]_ ) & (~\m1_addr_i[4]  | ~\new_[18899]_ );
  assign \new_[14105]_  = ~\new_[16580]_  | ~\new_[19444]_ ;
  assign \new_[14106]_  = (~\m7_data_i[16]  | ~\new_[17236]_ ) & (~\m0_data_i[16]  | ~\new_[18731]_ );
  assign \new_[14107]_  = ~\new_[16607]_  | ~\new_[19447]_ ;
  assign \new_[14108]_  = (~\m7_data_i[15]  | ~\new_[17236]_ ) & (~\m0_data_i[15]  | ~\new_[18731]_ );
  assign \new_[14109]_  = ~\new_[16613]_  | ~\new_[20458]_ ;
  assign \new_[14110]_  = (~\m7_data_i[14]  | ~\new_[17233]_ ) & (~\m0_data_i[14]  | ~\new_[20539]_ );
  assign \new_[14111]_  = (~\m2_data_i[14]  | ~\new_[18799]_ ) & (~\m1_data_i[14]  | ~\new_[20571]_ );
  assign \new_[14112]_  = ~\new_[28996]_  & (~\new_[16882]_  | ~\new_[28962]_ );
  assign \new_[14113]_  = (~\m7_data_i[13]  | ~\new_[17236]_ ) & (~\m0_data_i[13]  | ~\new_[20539]_ );
  assign \new_[14114]_  = ~\new_[16532]_  & (~\new_[17317]_  | ~\new_[6274]_ );
  assign \new_[14115]_  = ~\new_[28858]_  & (~\new_[16892]_  | ~\new_[29202]_ );
  assign \new_[14116]_  = (~\m5_sel_i[3]  | ~\new_[17199]_ ) & (~\m6_sel_i[3]  | ~\new_[18789]_ );
  assign \new_[14117]_  = (~m2_we_i | ~\new_[19567]_ ) & (~m1_we_i | ~\new_[19626]_ );
  assign \new_[14118]_  = (~\m7_data_i[12]  | ~\new_[18823]_ ) & (~\m0_data_i[12]  | ~\new_[20539]_ );
  assign \new_[14119]_  = (~\m7_data_i[11]  | ~\new_[17236]_ ) & (~\m0_data_i[11]  | ~\new_[20539]_ );
  assign \new_[14120]_  = (~\m2_data_i[11]  | ~\new_[18799]_ ) & (~\m1_data_i[11]  | ~\new_[18887]_ );
  assign \new_[14121]_  = ~\new_[29030]_  & (~\new_[16969]_  | ~\new_[29744]_ );
  assign \new_[14122]_  = ~\new_[30100]_  & (~\new_[16971]_  | ~\new_[29350]_ );
  assign \new_[14123]_  = (~\m7_data_i[9]  | ~\new_[17233]_ ) & (~\m0_data_i[9]  | ~\new_[18732]_ );
  assign \new_[14124]_  = ~\new_[15920]_  & (~\new_[30598]_  | ~\new_[6033]_ );
  assign \new_[14125]_  = (~\m2_data_i[9]  | ~\new_[18799]_ ) & (~\m1_data_i[9]  | ~\new_[20571]_ );
  assign \new_[14126]_  = ~\new_[15921]_  & (~\new_[30287]_  | ~\new_[6040]_ );
  assign \new_[14127]_  = (~\m7_data_i[8]  | ~\new_[18823]_ ) & (~\m0_data_i[8]  | ~\new_[18732]_ );
  assign \new_[14128]_  = ~\new_[15922]_  & (~\new_[30109]_  | ~\new_[6032]_ );
  assign \new_[14129]_  = (~\m7_data_i[7]  | ~\new_[17233]_ ) & (~\m0_data_i[7]  | ~\new_[20539]_ );
  assign \new_[14130]_  = (~\m2_data_i[7]  | ~\new_[18799]_ ) & (~\m1_data_i[7]  | ~\new_[18887]_ );
  assign \new_[14131]_  = ~\new_[16232]_  & (~\new_[30093]_  | ~\new_[31712]_ );
  assign \new_[14132]_  = ~\new_[16687]_  & (~\new_[30130]_  | ~\new_[31232]_ );
  assign \new_[14133]_  = ~\new_[16641]_  & (~\new_[29181]_  | ~\new_[31232]_ );
  assign \new_[14134]_  = ~\new_[16573]_  & (~\new_[29959]_  | ~\new_[31440]_ );
  assign \new_[14135]_  = (~\m7_data_i[6]  | ~\new_[17233]_ ) & (~\m0_data_i[6]  | ~\new_[20539]_ );
  assign \new_[14136]_  = ~\new_[15924]_  & (~\new_[30515]_  | ~\new_[6196]_ );
  assign \new_[14137]_  = (~\m5_addr_i[6]  | ~\new_[17187]_ ) & (~\m6_addr_i[6]  | ~\new_[18048]_ );
  assign \new_[14138]_  = ~\new_[16382]_  & (~\new_[30254]_  | ~\new_[30897]_ );
  assign \new_[14139]_  = (~\m7_data_i[23]  | ~\new_[18113]_ ) & (~\m0_data_i[23]  | ~\new_[19552]_ );
  assign \new_[14140]_  = ~\new_[16364]_  & (~\new_[30423]_  | ~\new_[31157]_ );
  assign \new_[14141]_  = ~\new_[15930]_  & (~\new_[30157]_  | ~\new_[6184]_ );
  assign \new_[14142]_  = (~\m7_data_i[22]  | ~\new_[18113]_ ) & (~\m0_data_i[22]  | ~\new_[19552]_ );
  assign \new_[14143]_  = (~\m7_data_i[5]  | ~\new_[17236]_ ) & (~\m0_data_i[5]  | ~\new_[20539]_ );
  assign \new_[14144]_  = ~\new_[16347]_  & (~\new_[30063]_  | ~\new_[6069]_ );
  assign \new_[14145]_  = (~\m7_data_i[4]  | ~\new_[17233]_ ) & (~\m0_data_i[4]  | ~\new_[20539]_ );
  assign \new_[14146]_  = (~\m7_data_i[21]  | ~\new_[18113]_ ) & (~\m0_data_i[21]  | ~\new_[18018]_ );
  assign \new_[14147]_  = ~\new_[15926]_  & (~\new_[28204]_  | ~\new_[5924]_ );
  assign \new_[14148]_  = (~\m7_data_i[20]  | ~\new_[18113]_ ) & (~\m0_data_i[20]  | ~\new_[18018]_ );
  assign \new_[14149]_  = ~\new_[15927]_  & (~\new_[29671]_  | ~\new_[5926]_ );
  assign \new_[14150]_  = (~\m2_data_i[4]  | ~\new_[18799]_ ) & (~\m1_data_i[4]  | ~\new_[20571]_ );
  assign \new_[14151]_  = ~\new_[15928]_  & (~\new_[30309]_  | ~\new_[6078]_ );
  assign \new_[14152]_  = ~\new_[15929]_  & (~\new_[30445]_  | ~\new_[6084]_ );
  assign \new_[14153]_  = (~\m7_data_i[3]  | ~\new_[17236]_ ) & (~\m0_data_i[3]  | ~\new_[20539]_ );
  assign \new_[14154]_  = ~\new_[15931]_  & (~\new_[30047]_  | ~\new_[6216]_ );
  assign \new_[14155]_  = (~\m7_data_i[2]  | ~\new_[18823]_ ) & (~\m0_data_i[2]  | ~\new_[18732]_ );
  assign \new_[14156]_  = ~\new_[15933]_  & (~\new_[29172]_  | ~\new_[6094]_ );
  assign \new_[14157]_  = (~\m5_addr_i[0]  | ~\new_[17188]_ ) & (~\m6_addr_i[0]  | ~\new_[18050]_ );
  assign \new_[14158]_  = (~\new_[16806]_  | ~\new_[30111]_ ) & (~\new_[30694]_  | ~\new_[6040]_ );
  assign \new_[14159]_  = (~\m7_data_i[1]  | ~\new_[17233]_ ) & (~\m0_data_i[1]  | ~\new_[19537]_ );
  assign \new_[14160]_  = (~\new_[16953]_  | ~\new_[30280]_ ) & (~\new_[29582]_  | ~\new_[31648]_ );
  assign \new_[14161]_  = (~\new_[16822]_  | ~\new_[29975]_ ) & (~\new_[30747]_  | ~\new_[31148]_ );
  assign \new_[14162]_  = (~\m2_data_i[1]  | ~\new_[18799]_ ) & (~\m1_data_i[1]  | ~\new_[20571]_ );
  assign \new_[14163]_  = (~\m7_data_i[13]  | ~\new_[18113]_ ) & (~\m0_data_i[13]  | ~\new_[18018]_ );
  assign \new_[14164]_  = (~\new_[16838]_  | ~\new_[30505]_ ) & (~\new_[28317]_  | ~\new_[6096]_ );
  assign \new_[14165]_  = (~\m7_data_i[12]  | ~\new_[18113]_ ) & (~\m0_data_i[12]  | ~\new_[18018]_ );
  assign \new_[14166]_  = ~\new_[16564]_  & (~\new_[30044]_  | ~\new_[31232]_ );
  assign \new_[14167]_  = (~\new_[16858]_  | ~\new_[30409]_ ) & (~\new_[29576]_  | ~\new_[31232]_ );
  assign \new_[14168]_  = (~\new_[17235]_  | ~\m7_addr_i[31] ) & (~\new_[18732]_  | ~\m0_addr_i[31] );
  assign \new_[14169]_  = (~\m7_data_i[11]  | ~\new_[18114]_ ) & (~\m0_data_i[11]  | ~\new_[18018]_ );
  assign \new_[14170]_  = ~\new_[16569]_  & (~\new_[28982]_  | ~\new_[5978]_ );
  assign \new_[14171]_  = (~\new_[16976]_  | ~\new_[30005]_ ) & (~\new_[29089]_  | ~\new_[5978]_ );
  assign \new_[14172]_  = (~\m7_data_i[10]  | ~\new_[18114]_ ) & (~\m0_data_i[10]  | ~\new_[18018]_ );
  assign \new_[14173]_  = (~\new_[18799]_  | ~\new_[31537]_ ) & (~\new_[18887]_  | ~\m1_addr_i[31] );
  assign \new_[14174]_  = ~\new_[16575]_  & (~\new_[29331]_  | ~\new_[5983]_ );
  assign \new_[14175]_  = (~\m7_data_i[9]  | ~\new_[18113]_ ) & (~\m0_data_i[9]  | ~\new_[18020]_ );
  assign \new_[14176]_  = (~\new_[16894]_  | ~\new_[30086]_ ) & (~\new_[29639]_  | ~\new_[5983]_ );
  assign \new_[14177]_  = (~\m7_data_i[8]  | ~\new_[18114]_ ) & (~\m0_data_i[8]  | ~\new_[18018]_ );
  assign \new_[14178]_  = (~\new_[16947]_  | ~\new_[29867]_ ) & (~\new_[30632]_  | ~\new_[6066]_ );
  assign \new_[14179]_  = (~\new_[18823]_  | ~\new_[31885]_ ) & (~\new_[19537]_  | ~\new_[31292]_ );
  assign \new_[14180]_  = (~\new_[16925]_  | ~\new_[30321]_ ) & (~\new_[30656]_  | ~\new_[6072]_ );
  assign \new_[14181]_  = (~\m7_data_i[6]  | ~\new_[18113]_ ) & (~\m0_data_i[6]  | ~\new_[18018]_ );
  assign \new_[14182]_  = (~\m7_data_i[5]  | ~\new_[18113]_ ) & (~\m0_data_i[5]  | ~\new_[18020]_ );
  assign \new_[14183]_  = ~\new_[16595]_  & (~\new_[28950]_  | ~\new_[5926]_ );
  assign \new_[14184]_  = (~\new_[18799]_  | ~\new_[31547]_ ) & (~\new_[20571]_  | ~\new_[31458]_ );
  assign \new_[14185]_  = (~\new_[16929]_  | ~\new_[30089]_ ) & (~\new_[30543]_  | ~\new_[6084]_ );
  assign \new_[14186]_  = (~\new_[17235]_  | ~\new_[30577]_ ) & (~\new_[19537]_  | ~\new_[30957]_ );
  assign \new_[14187]_  = (~\m7_data_i[3]  | ~\new_[18113]_ ) & (~\m0_data_i[3]  | ~\new_[18020]_ );
  assign \new_[14188]_  = ~\new_[16603]_  & (~\new_[29096]_  | ~\new_[31648]_ );
  assign \new_[14189]_  = ~\new_[16608]_  & (~\new_[29166]_  | ~\new_[31763]_ );
  assign \new_[14190]_  = (~\new_[16973]_  | ~\new_[30123]_ ) & (~\new_[29333]_  | ~\new_[31763]_ );
  assign \new_[14191]_  = (~\new_[18799]_  | ~\m2_addr_i[27] ) & (~\new_[20571]_  | ~\m1_addr_i[27] );
  assign \new_[14192]_  = (~\m7_data_i[2]  | ~\new_[18114]_ ) & (~\m0_data_i[2]  | ~\new_[18018]_ );
  assign \new_[14193]_  = (~\new_[17235]_  | ~\m7_addr_i[27] ) & (~\new_[19537]_  | ~\m0_addr_i[27] );
  assign \new_[14194]_  = (~\new_[16982]_  | ~\new_[30104]_ ) & (~\new_[29676]_  | ~\new_[6094]_ );
  assign \new_[14195]_  = \new_[16790]_  ? \new_[30042]_  : \new_[6202]_ ;
  assign \new_[14196]_  = (~\m7_data_i[1]  | ~\new_[18113]_ ) & (~\m0_data_i[1]  | ~\new_[18018]_ );
  assign \new_[14197]_  = (~\m7_data_i[19]  | ~\new_[17236]_ ) & (~\m0_data_i[19]  | ~\new_[19535]_ );
  assign \new_[14198]_  = (~\new_[17233]_  | ~\m7_addr_i[26] ) & (~\new_[19537]_  | ~\m0_addr_i[26] );
  assign \new_[14199]_  = ~\new_[28385]_  & (~\new_[17159]_  | ~\new_[30582]_ );
  assign \new_[14200]_  = (~\new_[18799]_  | ~\m2_addr_i[26] ) & (~\new_[18887]_  | ~\m1_addr_i[26] );
  assign \new_[14201]_  = ~\new_[28473]_  & (~\new_[17160]_  | ~\new_[29003]_ );
  assign \new_[14202]_  = ~\new_[26387]_  & (~\new_[17161]_  | ~\new_[29192]_ );
  assign \new_[14203]_  = (~\new_[17235]_  | ~\m7_addr_i[25] ) & (~\new_[19537]_  | ~\m0_addr_i[25] );
  assign \new_[14204]_  = (~\new_[18113]_  | ~\new_[31885]_ ) & (~\new_[18020]_  | ~\new_[31292]_ );
  assign \new_[14205]_  = (~\new_[18799]_  | ~\m2_addr_i[25] ) & (~\new_[20571]_  | ~\m1_addr_i[25] );
  assign \new_[14206]_  = (~\new_[18114]_  | ~\new_[31531]_ ) & (~\new_[18018]_  | ~\new_[31481]_ );
  assign \new_[14207]_  = (~\new_[17233]_  | ~\m7_addr_i[24] ) & (~\new_[19537]_  | ~\m0_addr_i[24] );
  assign \new_[14208]_  = \new_[6081]_  ? \new_[29042]_  : \new_[17308]_ ;
  assign \new_[14209]_  = ~\new_[28799]_  & (~\new_[17162]_  | ~\new_[30497]_ );
  assign \new_[14210]_  = \new_[16860]_  ? \new_[29777]_  : \new_[31423]_ ;
  assign \new_[14211]_  = (~\new_[18799]_  | ~\m2_addr_i[24] ) & (~\new_[20571]_  | ~\m1_addr_i[24] );
  assign \new_[14212]_  = ~\new_[26846]_  & (~\new_[17163]_  | ~\new_[29831]_ );
  assign \new_[14213]_  = \new_[16885]_  ? \new_[29865]_  : \new_[6056]_ ;
  assign \new_[14214]_  = (~\m2_addr_i[23]  | ~\new_[18799]_ ) & (~\m1_addr_i[23]  | ~\new_[18887]_ );
  assign \new_[14215]_  = ~\new_[28381]_  & (~\new_[17164]_  | ~\new_[29271]_ );
  assign \new_[14216]_  = \new_[16916]_  ? \new_[29994]_  : \new_[6062]_ ;
  assign \new_[14217]_  = ~\new_[27971]_  & (~\new_[17165]_  | ~\new_[30329]_ );
  assign \new_[14218]_  = (~\m7_addr_i[22]  | ~\new_[17234]_ ) & (~\m0_addr_i[22]  | ~\new_[19537]_ );
  assign \new_[14219]_  = ~\new_[24754]_  & (~\new_[17166]_  | ~\new_[28930]_ );
  assign \new_[14220]_  = (~\m2_addr_i[22]  | ~\new_[18799]_ ) & (~\m1_addr_i[22]  | ~\new_[20571]_ );
  assign \new_[14221]_  = ~\new_[27698]_  & (~\new_[17171]_  | ~\new_[28073]_ );
  assign \new_[14222]_  = ~\new_[26767]_  & (~\new_[17167]_  | ~\new_[28285]_ );
  assign \new_[14223]_  = ~\new_[28703]_  & (~\new_[17158]_  | ~\new_[30842]_ );
  assign \new_[14224]_  = ~\new_[26943]_  & (~\new_[17168]_  | ~\new_[27802]_ );
  assign \new_[14225]_  = (~\m2_addr_i[21]  | ~\new_[18799]_ ) & (~\m1_addr_i[21]  | ~\new_[20571]_ );
  assign \new_[14226]_  = ~\new_[24704]_  & (~\new_[17173]_  | ~\new_[28935]_ );
  assign \new_[14227]_  = (~\m7_addr_i[20]  | ~\new_[17234]_ ) & (~\m0_addr_i[20]  | ~\new_[19537]_ );
  assign \new_[14228]_  = \new_[16963]_  ? \new_[30277]_  : \new_[6080]_ ;
  assign \new_[14229]_  = ~\new_[28383]_  & (~\new_[17169]_  | ~\new_[29608]_ );
  assign \new_[14230]_  = (~\m2_addr_i[20]  | ~\new_[18799]_ ) & (~\m1_addr_i[20]  | ~\new_[20571]_ );
  assign \new_[14231]_  = ~\new_[27534]_  & (~\new_[17172]_  | ~\new_[28280]_ );
  assign \new_[14232]_  = (~\m7_addr_i[19]  | ~\new_[17234]_ ) & (~\m0_addr_i[19]  | ~\new_[19535]_ );
  assign \new_[14233]_  = ~\new_[28731]_  & (~\new_[17170]_  | ~\new_[29571]_ );
  assign \new_[14234]_  = \new_[16809]_  ? \new_[29772]_  : \new_[6087]_ ;
  assign \new_[14235]_  = \new_[16975]_  ? \new_[30208]_  : \new_[6091]_ ;
  assign \new_[14236]_  = (~\m7_addr_i[18]  | ~\new_[17235]_ ) & (~\m0_addr_i[18]  | ~\new_[19535]_ );
  assign \new_[14237]_  = ~\new_[28227]_  & (~\new_[17174]_  | ~\new_[30764]_ );
  assign \new_[14238]_  = ~\new_[16548]_  | ~\new_[22229]_ ;
  assign \new_[14239]_  = ~\new_[26794]_  | (~\new_[16791]_  & ~\new_[30145]_ );
  assign \new_[14240]_  = ~\new_[21535]_  | (~\new_[16802]_  & ~\new_[29841]_ );
  assign \new_[14241]_  = ~\new_[22811]_  & (~\new_[16803]_  | ~\new_[28908]_ );
  assign \new_[14242]_  = ~\new_[16552]_  | ~\new_[22892]_ ;
  assign \new_[14243]_  = ~\new_[22961]_  | (~\new_[16805]_  & ~\new_[29907]_ );
  assign \new_[14244]_  = (~\m7_addr_i[17]  | ~\new_[17236]_ ) & (~\m0_addr_i[17]  | ~\new_[20539]_ );
  assign \new_[14245]_  = (~\m7_addr_i[16]  | ~\new_[17234]_ ) & (~\m0_addr_i[16]  | ~\new_[18732]_ );
  assign \new_[14246]_  = ~\new_[21540]_  | (~\new_[16816]_  & ~\new_[30415]_ );
  assign \new_[14247]_  = (~\m2_addr_i[16]  | ~\new_[18799]_ ) & (~\m1_addr_i[16]  | ~\new_[18887]_ );
  assign \new_[14248]_  = ~\new_[22769]_  & (~\new_[16818]_  | ~\new_[29112]_ );
  assign \new_[14249]_  = ~\new_[16554]_  | ~\new_[22973]_ ;
  assign \new_[14250]_  = ~\new_[24721]_  | (~\new_[16820]_  & ~\new_[29810]_ );
  assign \new_[14251]_  = (~\m7_addr_i[15]  | ~\new_[17235]_ ) & (~\m0_addr_i[15]  | ~\new_[18732]_ );
  assign \new_[14252]_  = ~\new_[21475]_  | (~\new_[16834]_  & ~\new_[30202]_ );
  assign \new_[14253]_  = ~\new_[22752]_  & (~\new_[16835]_  | ~\new_[28968]_ );
  assign \new_[14254]_  = (~\m7_addr_i[14]  | ~\new_[17235]_ ) & (~\m0_addr_i[14]  | ~\new_[18732]_ );
  assign \new_[14255]_  = ~\new_[17896]_  | ~\new_[28753]_  | ~\new_[28969]_  | ~\new_[28050]_ ;
  assign \new_[14256]_  = (~\m7_data_i[17]  | ~\new_[17236]_ ) & (~\m0_data_i[17]  | ~\new_[20539]_ );
  assign \new_[14257]_  = ~\new_[17905]_  | ~\new_[28202]_  | ~\new_[29783]_  | ~\new_[26655]_ ;
  assign \new_[14258]_  = ~\new_[21507]_  | (~\new_[16844]_  & ~\new_[29931]_ );
  assign \new_[14259]_  = (~\m7_addr_i[8]  | ~\new_[18113]_ ) & (~\m0_addr_i[8]  | ~\new_[18018]_ );
  assign \new_[14260]_  = ~\new_[17909]_  | ~\new_[29756]_  | ~\new_[28840]_  | ~\new_[29186]_ ;
  assign \new_[14261]_  = (~\m7_addr_i[13]  | ~\new_[17234]_ ) & (~\m0_addr_i[13]  | ~\new_[18732]_ );
  assign \new_[14262]_  = ~\new_[28775]_  & (~\new_[17157]_  | ~\new_[21456]_ );
  assign \new_[14263]_  = (~\m2_addr_i[12]  | ~\new_[18799]_ ) & (~\m1_addr_i[12]  | ~\new_[20571]_ );
  assign \new_[14264]_  = (~\m7_addr_i[12]  | ~\new_[17236]_ ) & (~\m0_addr_i[12]  | ~\new_[18731]_ );
  assign \new_[14265]_  = ~\new_[20504]_  | (~\new_[16883]_  & ~\new_[29445]_ );
  assign \new_[14266]_  = ~\new_[22723]_  & (~\new_[16933]_  | ~\new_[29189]_ );
  assign \new_[14267]_  = ~\new_[16570]_  | ~\new_[24268]_ ;
  assign \new_[14268]_  = ~\new_[26324]_  | (~\new_[16946]_  & ~\new_[30033]_ );
  assign \new_[14269]_  = ~\new_[17912]_  | ~\new_[28161]_  | ~\new_[30344]_  | ~\new_[28684]_ ;
  assign \new_[14270]_  = (~\m7_addr_i[11]  | ~\new_[18823]_ ) & (~\m0_addr_i[11]  | ~\new_[20539]_ );
  assign \new_[14271]_  = ~\new_[17914]_  | ~\new_[27981]_  | ~\new_[30294]_  | ~\new_[30628]_ ;
  assign \new_[14272]_  = ~\new_[20461]_  | (~\new_[16893]_  & ~\new_[29174]_ );
  assign \new_[14273]_  = (~\m7_addr_i[10]  | ~\new_[17234]_ ) & (~\m0_addr_i[10]  | ~\new_[18732]_ );
  assign \new_[14274]_  = ~\new_[17916]_  | ~\new_[29786]_  | ~\new_[29162]_  | ~\new_[28121]_ ;
  assign \new_[14275]_  = (~\m7_addr_i[0]  | ~\new_[18113]_ ) & (~\m0_addr_i[0]  | ~\new_[18018]_ );
  assign \new_[14276]_  = ~\new_[21508]_  | (~\new_[16907]_  & ~\new_[30053]_ );
  assign \new_[14277]_  = (~\m7_addr_i[9]  | ~\new_[17234]_ ) & (~\m0_addr_i[9]  | ~\new_[19535]_ );
  assign \new_[14278]_  = (~\m7_sel_i[3]  | ~\new_[18113]_ ) & (~\m0_sel_i[3]  | ~\new_[19552]_ );
  assign \new_[14279]_  = ~\new_[16577]_  | ~\new_[24451]_ ;
  assign \new_[14280]_  = (~\m2_addr_i[9]  | ~\new_[18799]_ ) & (~\m1_addr_i[9]  | ~\new_[18887]_ );
  assign \new_[14281]_  = ~\new_[24748]_  | (~\new_[16903]_  & ~\new_[30326]_ );
  assign \new_[14282]_  = ~\new_[17931]_  | ~\new_[28040]_  | ~\new_[29086]_  | ~\new_[28245]_ ;
  assign \new_[14283]_  = (~\m7_sel_i[2]  | ~\new_[18113]_ ) & (~\m0_sel_i[2]  | ~\new_[19552]_ );
  assign \new_[14284]_  = ~\new_[20525]_  | (~\new_[16819]_  & ~\new_[30212]_ );
  assign \new_[14285]_  = (~\m2_addr_i[8]  | ~\new_[18799]_ ) & (~\m1_addr_i[8]  | ~\new_[18887]_ );
  assign \new_[14286]_  = ~\new_[22828]_  & (~\new_[16909]_  | ~\new_[29633]_ );
  assign \new_[14287]_  = ~\new_[16582]_  | ~\new_[22966]_ ;
  assign \new_[14288]_  = ~\new_[24673]_  | (~\new_[16937]_  & ~\new_[30375]_ );
  assign \new_[14289]_  = ~\new_[17919]_  | ~\new_[28951]_  | ~\new_[29175]_  | ~\new_[28073]_ ;
  assign \new_[14290]_  = (~\m7_addr_i[8]  | ~\new_[17235]_ ) & (~\m0_addr_i[8]  | ~\new_[19535]_ );
  assign \new_[14291]_  = (~\m7_addr_i[7]  | ~\new_[17235]_ ) & (~\m0_addr_i[7]  | ~\new_[20539]_ );
  assign \new_[14292]_  = ~\new_[21533]_  | (~\new_[16906]_  & ~\new_[30058]_ );
  assign \new_[14293]_  = ~\new_[22656]_  & (~\new_[16934]_  | ~\new_[28864]_ );
  assign \new_[14294]_  = ~\new_[16588]_  | ~\new_[22911]_ ;
  assign \new_[14295]_  = (~\m7_addr_i[6]  | ~\new_[17235]_ ) & (~\m0_addr_i[6]  | ~\new_[20539]_ );
  assign \new_[14296]_  = (~\m2_addr_i[6]  | ~\new_[18799]_ ) & (~\m1_addr_i[6]  | ~\new_[18887]_ );
  assign \new_[14297]_  = (~\m7_addr_i[5]  | ~\new_[17233]_ ) & (~\new_[31848]_  | ~\new_[20539]_ );
  assign \new_[14298]_  = (~\m2_addr_i[5]  | ~\new_[18799]_ ) & (~\m1_addr_i[5]  | ~\new_[20571]_ );
  assign \new_[14299]_  = ~\new_[21502]_  | (~\new_[16919]_  & ~\new_[30114]_ );
  assign \new_[14300]_  = ~\new_[22817]_  & (~\new_[16793]_  | ~\new_[28844]_ );
  assign \new_[14301]_  = ~\new_[16590]_  | ~\new_[20506]_ ;
  assign \new_[14302]_  = ~\new_[26245]_  | (~\new_[16796]_  & ~\new_[29792]_ );
  assign \new_[14303]_  = ~\new_[17907]_  | ~\new_[28932]_  | ~\new_[28878]_  | ~\new_[28732]_ ;
  assign \new_[14304]_  = (~\m7_addr_i[4]  | ~\new_[17233]_ ) & (~\m0_addr_i[4]  | ~\new_[19537]_ );
  assign \new_[14305]_  = (~\m2_addr_i[4]  | ~\new_[18799]_ ) & (~\m1_addr_i[4]  | ~\new_[20571]_ );
  assign \new_[14306]_  = ~\new_[22937]_  & (~\new_[16787]_  | ~\new_[30138]_ );
  assign \new_[14307]_  = ~\new_[21527]_  | (~\new_[16970]_  & ~\new_[29944]_ );
  assign \new_[14308]_  = ~\new_[16606]_  | ~\new_[22587]_ ;
  assign \new_[14309]_  = ~\new_[26653]_  | (~\new_[16926]_  & ~\new_[30151]_ );
  assign \new_[14310]_  = ~\new_[17936]_  | ~\new_[28345]_  | ~\new_[30126]_  | ~\new_[28640]_ ;
  assign \new_[14311]_  = (~\new_[31726]_  | ~\new_[17233]_ ) & (~\m0_addr_i[3]  | ~\new_[20539]_ );
  assign \new_[14312]_  = (~\m2_addr_i[3]  | ~\new_[18799]_ ) & (~\m1_addr_i[3]  | ~\new_[18887]_ );
  assign \new_[14313]_  = ~\new_[16545]_  | (~\new_[30343]_  & ~\new_[5925]_ );
  assign \new_[14314]_  = ~\new_[21518]_  | (~\new_[16931]_  & ~\new_[30140]_ );
  assign \new_[14315]_  = ~\new_[16600]_  | ~\new_[22950]_ ;
  assign \new_[14316]_  = ~\new_[23145]_  | (~\new_[16943]_  & ~\new_[29997]_ );
  assign \new_[14317]_  = (~\m7_addr_i[2]  | ~\new_[17236]_ ) & (~\m0_addr_i[2]  | ~\new_[19537]_ );
  assign \new_[14318]_  = ~\new_[21474]_  & (~\new_[16785]_  | ~\new_[28889]_ );
  assign \new_[14319]_  = (~\m2_addr_i[2]  | ~\new_[18799]_ ) & (~\m1_addr_i[2]  | ~\new_[18887]_ );
  assign \new_[14320]_  = ~\new_[17925]_  | ~\new_[28288]_  | ~\new_[29886]_  | ~\new_[28535]_ ;
  assign \new_[14321]_  = ~\new_[22897]_  & (~\new_[16786]_  | ~\new_[29886]_ );
  assign \new_[14322]_  = ~\new_[20474]_  | (~\new_[16952]_  & ~\new_[29629]_ );
  assign \new_[14323]_  = (~\m7_addr_i[1]  | ~\new_[17236]_ ) & (~\m0_addr_i[1]  | ~\new_[20539]_ );
  assign \new_[14324]_  = ~\new_[17924]_  | ~\new_[29433]_  | ~\new_[30333]_  | ~\new_[30117]_ ;
  assign \new_[14325]_  = ~\new_[20453]_  | (~\new_[16972]_  & ~\new_[29564]_ );
  assign \new_[14326]_  = (~\m7_addr_i[0]  | ~\new_[17236]_ ) & (~\m0_addr_i[0]  | ~\new_[19535]_ );
  assign \new_[14327]_  = ~\new_[21544]_  | (~\new_[16981]_  & ~\new_[29861]_ );
  assign \new_[14328]_  = (~\m7_sel_i[3]  | ~\new_[17235]_ ) & (~\m0_sel_i[3]  | ~\new_[19535]_ );
  assign \new_[14329]_  = (~\m2_sel_i[2]  | ~\new_[18799]_ ) & (~\m1_sel_i[2]  | ~\new_[18887]_ );
  assign \new_[14330]_  = (~\m7_sel_i[2]  | ~\new_[17233]_ ) & (~\m0_sel_i[2]  | ~\new_[19537]_ );
  assign \new_[14331]_  = (~\m7_sel_i[0]  | ~\new_[17235]_ ) & (~\m0_sel_i[0]  | ~\new_[19535]_ );
  assign \new_[14332]_  = (~m7_we_i | ~\new_[17233]_ ) & (~m0_we_i | ~\new_[20539]_ );
  assign \new_[14333]_  = ~\new_[15662]_ ;
  assign \new_[14334]_  = (~m2_we_i | ~\new_[18799]_ ) & (~m1_we_i | ~\new_[18887]_ );
  assign \new_[14335]_  = (~\new_[17758]_  | ~s7_err_i) & (~\new_[17046]_  | ~s6_err_i);
  assign \new_[14336]_  = ~\new_[15666]_ ;
  assign \new_[14337]_  = (~\new_[17758]_  | ~s7_rty_i) & (~\new_[17046]_  | ~s6_rty_i);
  assign \new_[14338]_  = (~\m5_data_i[31]  | ~\new_[18740]_ ) & (~\m6_data_i[31]  | ~\new_[20550]_ );
  assign \new_[14339]_  = (~\m7_data_i[30]  | ~\new_[18824]_ ) & (~\m0_data_i[30]  | ~\new_[18011]_ );
  assign \new_[14340]_  = (~\m7_data_i[29]  | ~\new_[18824]_ ) & (~\m0_data_i[29]  | ~\new_[18011]_ );
  assign \new_[14341]_  = (~\m5_data_i[29]  | ~\new_[18740]_ ) & (~\m6_data_i[29]  | ~\new_[18786]_ );
  assign \new_[14342]_  = (~\m7_data_i[28]  | ~\new_[18824]_ ) & (~\m0_data_i[28]  | ~\new_[18011]_ );
  assign \new_[14343]_  = (~\m7_data_i[27]  | ~\new_[18824]_ ) & (~\m0_data_i[27]  | ~\new_[18011]_ );
  assign \new_[14344]_  = (~\m5_data_i[27]  | ~\new_[18740]_ ) & (~\m6_data_i[27]  | ~\new_[18786]_ );
  assign \new_[14345]_  = \new_[5964]_  ? \new_[28845]_  : \new_[17115]_ ;
  assign \new_[14346]_  = \new_[30511]_  ? \new_[30139]_  : \new_[17117]_ ;
  assign \new_[14347]_  = \new_[5913]_  ? \new_[28880]_  : \new_[17122]_ ;
  assign \new_[14348]_  = \new_[6206]_  ? \new_[29783]_  : \new_[17123]_ ;
  assign \new_[14349]_  = \new_[6031]_  ? \new_[29922]_  : \new_[17124]_ ;
  assign \new_[14350]_  = (~\new_[17137]_  | ~\new_[29682]_ ) & (~\new_[30068]_  | ~\new_[31394]_ );
  assign \new_[14351]_  = \new_[5981]_  ? \new_[29162]_  : \new_[17127]_ ;
  assign \new_[14352]_  = \new_[5981]_  ? \new_[30279]_  : \new_[17126]_ ;
  assign \new_[14353]_  = \new_[6064]_  ? \new_[30083]_  : \new_[17118]_ ;
  assign \new_[14354]_  = (~\m5_data_i[23]  | ~\new_[18740]_ ) & (~\m6_data_i[23]  | ~\new_[18786]_ );
  assign \new_[14355]_  = (~\m5_data_i[22]  | ~\new_[18740]_ ) & (~\m6_data_i[22]  | ~\new_[20550]_ );
  assign \new_[14356]_  = \new_[6190]_  ? \new_[29225]_  : \new_[17116]_ ;
  assign \new_[14357]_  = \new_[5991]_  ? \new_[29785]_  : \new_[17128]_ ;
  assign \new_[14358]_  = \new_[5994]_  ? \new_[30158]_  : \new_[17129]_ ;
  assign \new_[14359]_  = \new_[5996]_  ? \new_[30138]_  : \new_[17135]_ ;
  assign \new_[14360]_  = \new_[5996]_  ? \new_[30702]_  : \new_[17130]_ ;
  assign \new_[14361]_  = (~\m5_data_i[21]  | ~\new_[18740]_ ) & (~\m6_data_i[21]  | ~\new_[20550]_ );
  assign \new_[14362]_  = (~\m7_data_i[20]  | ~\new_[18825]_ ) & (~\m0_data_i[20]  | ~\new_[18011]_ );
  assign \new_[14363]_  = \new_[5999]_  ? \new_[28889]_  : \new_[17134]_ ;
  assign \new_[14364]_  = \new_[5999]_  ? \new_[29685]_  : \new_[17132]_ ;
  assign \new_[14365]_  = \new_[6001]_  ? \new_[29886]_  : \new_[17133]_ ;
  assign \new_[14366]_  = \new_[5931]_  ? \new_[29563]_  : \new_[17121]_ ;
  assign \new_[14367]_  = (~\m7_data_i[19]  | ~\new_[18825]_ ) & (~\m0_data_i[19]  | ~\new_[18011]_ );
  assign \new_[14368]_  = (~\m5_data_i[19]  | ~\new_[18740]_ ) & (~\m6_data_i[19]  | ~\new_[18786]_ );
  assign \new_[14369]_  = \new_[17012]_  & \new_[16137]_ ;
  assign \new_[14370]_  = \new_[27750]_  | \new_[16017]_ ;
  assign \new_[14371]_  = ~\new_[26679]_  & (~\new_[17175]_  | ~\new_[30164]_ );
  assign \new_[14372]_  = (~\m5_data_i[16]  | ~\new_[18740]_ ) & (~\m6_data_i[16]  | ~\new_[18786]_ );
  assign \new_[14373]_  = \new_[17023]_  & \new_[16142]_ ;
  assign \new_[14374]_  = ~\new_[30287]_  & (~\new_[17254]_  | ~\new_[26320]_ );
  assign \new_[14375]_  = ~\new_[16143]_  & ~\new_[23113]_ ;
  assign \new_[14376]_  = ~\new_[28727]_  & (~\new_[17176]_  | ~\new_[29219]_ );
  assign \new_[14377]_  = \new_[27824]_  | \new_[16026]_ ;
  assign \new_[14378]_  = (~\m5_data_i[15]  | ~\new_[18740]_ ) & (~\m6_data_i[15]  | ~\new_[18786]_ );
  assign \new_[14379]_  = ~\new_[27562]_  & (~\new_[17177]_  | ~\new_[30426]_ );
  assign \new_[14380]_  = (~\m7_data_i[10]  | ~\new_[17236]_ ) & (~\m0_data_i[10]  | ~\new_[20539]_ );
  assign \new_[14381]_  = (~\m5_data_i[14]  | ~\new_[18740]_ ) & (~\m6_data_i[14]  | ~\new_[18786]_ );
  assign \new_[14382]_  = ~\new_[27978]_  & (~\new_[17184]_  | ~\new_[28989]_ );
  assign \new_[14383]_  = \new_[26592]_  | \new_[16037]_ ;
  assign \new_[14384]_  = \new_[26614]_  | \new_[16046]_ ;
  assign \new_[14385]_  = ~\new_[28899]_  & (~\new_[17281]_  | ~\new_[28181]_ );
  assign \new_[14386]_  = ~\new_[16214]_  & ~\new_[24771]_ ;
  assign \new_[14387]_  = ~\new_[29977]_  | (~\new_[20887]_  & ~\new_[17310]_ );
  assign \new_[14388]_  = \new_[27574]_  | \new_[16074]_ ;
  assign \new_[14389]_  = ~\new_[27638]_  & (~\new_[17180]_  | ~\new_[29401]_ );
  assign \new_[14390]_  = \new_[16054]_  & \new_[16851]_ ;
  assign \new_[14391]_  = ~m2_stb_i | ~\new_[26175]_  | ~\new_[17224]_ ;
  assign \new_[14392]_  = (~\m5_data_i[9]  | ~\new_[18740]_ ) & (~\m6_data_i[9]  | ~\new_[18786]_ );
  assign \new_[14393]_  = (~\m5_data_i[8]  | ~\new_[18740]_ ) & (~\m6_data_i[8]  | ~\new_[18786]_ );
  assign \new_[14394]_  = \new_[23173]_  | \new_[16066]_ ;
  assign \new_[14395]_  = (~\m5_data_i[7]  | ~\new_[18740]_ ) & (~\m6_data_i[7]  | ~\new_[18786]_ );
  assign \new_[14396]_  = ~\new_[27610]_  & (~\new_[17182]_  | ~\new_[29221]_ );
  assign \new_[14397]_  = (~\m5_data_i[5]  | ~\new_[18740]_ ) & (~\m6_data_i[5]  | ~\new_[18786]_ );
  assign \new_[14398]_  = ~\new_[26575]_  & (~\new_[17178]_  | ~\new_[29171]_ );
  assign \new_[14399]_  = \new_[26751]_  | \new_[16081]_ ;
  assign \new_[14400]_  = ~\new_[29573]_  & (~\new_[17228]_  | ~\new_[28631]_ );
  assign \new_[14401]_  = ~\new_[16167]_  & ~\new_[24661]_ ;
  assign \new_[14402]_  = (~\m4_data_i[0]  | ~\new_[18149]_ ) & (~\m3_data_i[0]  | ~\new_[18930]_ );
  assign \new_[14403]_  = (~\m5_data_i[3]  | ~\new_[18740]_ ) & (~\m6_data_i[3]  | ~\new_[18786]_ );
  assign \new_[14404]_  = \new_[27410]_  | \new_[16097]_ ;
  assign \new_[14405]_  = (~\m7_addr_i[0]  | ~\new_[18116]_ ) & (~\m0_addr_i[0]  | ~\new_[18932]_ );
  assign \new_[14406]_  = (~\m5_data_i[2]  | ~\new_[18740]_ ) & (~\m6_data_i[2]  | ~\new_[18786]_ );
  assign \new_[14407]_  = ~\new_[29767]_  & (~\new_[17250]_  | ~\new_[28575]_ );
  assign \new_[14408]_  = ~\new_[16180]_  & ~\new_[25602]_ ;
  assign \new_[14409]_  = \new_[26438]_  | \new_[16087]_ ;
  assign \new_[14410]_  = (~\m5_data_i[0]  | ~\new_[18740]_ ) & (~\m6_data_i[0]  | ~\new_[18786]_ );
  assign \new_[14411]_  = \new_[28563]_  | \new_[16093]_ ;
  assign \new_[14412]_  = (~\new_[18786]_  | ~\m6_addr_i[31] ) & (~\new_[18740]_  | ~\new_[31001]_ );
  assign \new_[14413]_  = ~\new_[29565]_  & (~\new_[17209]_  | ~\new_[28373]_ );
  assign \new_[14414]_  = ~\new_[16197]_  & ~\new_[26345]_ ;
  assign \new_[14415]_  = (~\new_[18786]_  | ~\m6_addr_i[30] ) & (~\new_[18740]_  | ~\new_[31147]_ );
  assign \new_[14416]_  = \new_[26661]_  | \new_[16107]_ ;
  assign \new_[14417]_  = ~\new_[27679]_  & (~\new_[17179]_  | ~\new_[29061]_ );
  assign \new_[14418]_  = ~\new_[28305]_  | ~\new_[28964]_  | ~\new_[17351]_ ;
  assign \new_[14419]_  = (~\new_[18786]_  | ~\m6_addr_i[29] ) & (~\new_[18740]_  | ~\new_[31407]_ );
  assign \new_[14420]_  = ~\new_[16221]_  & ~\new_[23381]_ ;
  assign \new_[14421]_  = ~\new_[27356]_  & (~\new_[17186]_  | ~\new_[29038]_ );
  assign \new_[14422]_  = (~\new_[18786]_  | ~\m6_addr_i[28] ) & (~\new_[18740]_  | ~\new_[31276]_ );
  assign \new_[14423]_  = \new_[16191]_  & \new_[16192]_ ;
  assign \new_[14424]_  = \new_[16193]_  & \new_[16194]_ ;
  assign \new_[14425]_  = (~\new_[18786]_  | ~\m6_addr_i[27] ) & (~\new_[18740]_  | ~\m5_addr_i[27] );
  assign \new_[14426]_  = \new_[26721]_  | \new_[16106]_ ;
  assign \new_[14427]_  = ~m5_stb_i | ~\new_[24201]_  | ~\new_[17202]_ ;
  assign \new_[14428]_  = ~\new_[27689]_  & (~\new_[17181]_  | ~\new_[28007]_ );
  assign \new_[14429]_  = ~m3_stb_i | ~\new_[27519]_  | ~\new_[32350]_ ;
  assign \new_[14430]_  = (~\new_[18786]_  | ~\m6_addr_i[26] ) & (~\new_[18740]_  | ~\m5_addr_i[26] );
  assign \new_[14431]_  = (~\new_[18786]_  | ~\m6_addr_i[25] ) & (~\new_[18740]_  | ~\m5_addr_i[25] );
  assign \new_[14432]_  = \new_[26817]_  | \new_[16111]_ ;
  assign \new_[14433]_  = (~\new_[18786]_  | ~\m6_addr_i[24] ) & (~\new_[18740]_  | ~\m5_addr_i[24] );
  assign \new_[14434]_  = \new_[17075]_  & \new_[16199]_ ;
  assign \new_[14435]_  = \new_[16219]_  & \new_[17097]_ ;
  assign \new_[14436]_  = \new_[27533]_  | \new_[16126]_ ;
  assign \new_[14437]_  = ~\new_[16024]_  & ~\new_[29909]_ ;
  assign \new_[14438]_  = ~\new_[16029]_  & ~\new_[17295]_ ;
  assign \new_[14439]_  = ~\new_[16038]_  & ~\new_[17301]_ ;
  assign \new_[14440]_  = (~\m5_addr_i[21]  | ~\new_[18740]_ ) & (~\m6_addr_i[21]  | ~\new_[18786]_ );
  assign \new_[14441]_  = ~\new_[16098]_  & ~\new_[17335]_ ;
  assign \new_[14442]_  = ~\new_[16034]_  & ~\new_[17347]_ ;
  assign \new_[14443]_  = ~\new_[16088]_  & ~\new_[16323]_ ;
  assign \new_[14444]_  = ~\new_[16129]_  | ~\new_[26320]_ ;
  assign \new_[14445]_  = \new_[16130]_  | \new_[26351]_ ;
  assign \new_[14446]_  = \new_[16131]_  | \new_[26453]_ ;
  assign \new_[14447]_  = (~\m5_addr_i[18]  | ~\new_[18740]_ ) & (~\m6_addr_i[18]  | ~\new_[20550]_ );
  assign \new_[14448]_  = (~\m5_addr_i[7]  | ~\new_[17188]_ ) & (~\m6_addr_i[7]  | ~\new_[18049]_ );
  assign \new_[14449]_  = \new_[16132]_  | \new_[25466]_ ;
  assign \new_[14450]_  = (~\m5_addr_i[17]  | ~\new_[18740]_ ) & (~\m6_addr_i[17]  | ~\new_[20550]_ );
  assign \new_[14451]_  = (~\m7_addr_i[16]  | ~\new_[18825]_ ) & (~\m0_addr_i[16]  | ~\new_[18011]_ );
  assign \new_[14452]_  = \new_[16133]_  | \new_[28784]_ ;
  assign \new_[14453]_  = \new_[16134]_  | \new_[27634]_ ;
  assign \new_[14454]_  = (~\m7_addr_i[15]  | ~\new_[18825]_ ) & (~\m0_addr_i[15]  | ~\new_[18011]_ );
  assign \new_[14455]_  = ~\new_[16837]_  & (~\new_[17294]_  | ~\new_[31678]_ );
  assign \new_[14456]_  = ~\new_[15997]_  & (~\new_[17255]_  | ~\m1_addr_i[4] );
  assign \new_[14457]_  = ~\new_[15994]_  & (~\new_[17226]_  | ~\m3_addr_i[4] );
  assign \new_[14458]_  = (~\m7_addr_i[14]  | ~\new_[18825]_ ) & (~\m0_addr_i[14]  | ~\new_[18011]_ );
  assign \new_[14459]_  = ~\new_[15990]_  & (~\new_[17342]_  | ~\m6_addr_i[4] );
  assign \new_[14460]_  = ~\new_[15991]_  & (~\new_[17311]_  | ~\m4_addr_i[4] );
  assign \new_[14461]_  = ~\new_[15995]_  & (~\new_[31996]_  | ~\m7_addr_i[3] );
  assign \new_[14462]_  = ~\new_[16020]_  & (~\new_[18227]_  | ~\new_[31853]_ );
  assign \new_[14463]_  = (~\m5_addr_i[13]  | ~\new_[18740]_ ) & (~\m6_addr_i[13]  | ~\new_[18786]_ );
  assign \new_[14464]_  = ~\new_[22381]_  & (~\new_[17258]_  | ~\new_[28883]_ );
  assign \new_[14465]_  = (~\m5_addr_i[12]  | ~\new_[18740]_ ) & (~\m6_addr_i[12]  | ~\new_[20550]_ );
  assign \new_[14466]_  = (~\m7_addr_i[11]  | ~\new_[18825]_ ) & (~\m0_addr_i[11]  | ~\new_[18011]_ );
  assign \new_[14467]_  = (~\m5_addr_i[11]  | ~\new_[18740]_ ) & (~\m6_addr_i[11]  | ~\new_[18786]_ );
  assign \new_[14468]_  = \new_[6077]_  ? \new_[29589]_  : \new_[17334]_ ;
  assign \new_[14469]_  = ~\new_[16056]_  & (~\new_[17316]_  | ~\new_[31888]_ );
  assign \new_[14470]_  = (~\m5_addr_i[10]  | ~\new_[18740]_ ) & (~\m6_addr_i[10]  | ~\new_[18786]_ );
  assign \new_[14471]_  = (~\m7_addr_i[9]  | ~\new_[18825]_ ) & (~\m0_addr_i[9]  | ~\new_[18011]_ );
  assign \new_[14472]_  = (~\m5_addr_i[8]  | ~\new_[18740]_ ) & (~\m6_addr_i[8]  | ~\new_[20550]_ );
  assign \new_[14473]_  = (~\m7_addr_i[6]  | ~\new_[18825]_ ) & (~\m0_addr_i[6]  | ~\new_[18011]_ );
  assign \new_[14474]_  = (~\m5_addr_i[6]  | ~\new_[18740]_ ) & (~\m6_addr_i[6]  | ~\new_[20550]_ );
  assign \new_[14475]_  = ~\new_[16078]_  & (~\new_[17319]_  | ~\new_[31576]_ );
  assign \new_[14476]_  = (~\m5_addr_i[4]  | ~\new_[18740]_ ) & (~\m6_addr_i[4]  | ~\new_[18786]_ );
  assign \new_[14477]_  = ~\new_[17231]_  | ~\new_[31368]_  | ~n8694;
  assign \new_[14478]_  = ~\new_[16083]_  & (~\new_[18272]_  | ~\new_[31759]_ );
  assign \new_[14479]_  = (~\m5_addr_i[2]  | ~\new_[18740]_ ) & (~\m6_addr_i[2]  | ~\new_[18786]_ );
  assign \new_[14480]_  = (~\m5_addr_i[0]  | ~\new_[18740]_ ) & (~\m6_addr_i[0]  | ~\new_[18786]_ );
  assign \new_[14481]_  = ~\new_[16845]_  & (~\new_[17304]_  | ~\new_[31830]_ );
  assign \new_[14482]_  = (~\m5_sel_i[1]  | ~\new_[18740]_ ) & (~\m6_sel_i[1]  | ~\new_[20550]_ );
  assign \new_[14483]_  = (~\m5_addr_i[15]  | ~\new_[17187]_ ) & (~\m6_addr_i[15]  | ~\new_[18051]_ );
  assign \new_[14484]_  = (~\m5_sel_i[0]  | ~\new_[18740]_ ) & (~\m6_sel_i[0]  | ~\new_[20550]_ );
  assign \new_[14485]_  = (~m5_we_i | ~\new_[18740]_ ) & (~m6_we_i | ~\new_[20550]_ );
  assign \new_[14486]_  = (~\m7_data_i[20]  | ~\new_[17234]_ ) & (~\m0_data_i[20]  | ~\new_[19535]_ );
  assign \new_[14487]_  = (~\m4_data_i[31]  | ~\new_[17260]_ ) & (~\m3_data_i[31]  | ~\new_[18175]_ );
  assign \new_[14488]_  = (~\m5_data_i[30]  | ~\new_[17188]_ ) & (~\m6_data_i[30]  | ~\new_[19563]_ );
  assign \new_[14489]_  = ~\new_[27861]_  & (~\new_[24763]_  | ~\new_[17352]_ );
  assign \new_[14490]_  = (~\m2_addr_i[10]  | ~\new_[19567]_ ) & (~\m1_addr_i[10]  | ~\new_[19626]_ );
  assign \new_[14491]_  = ~\new_[16930]_  & (~\new_[17336]_  | ~\new_[31698]_ );
  assign \new_[14492]_  = (~\m4_data_i[28]  | ~\new_[17260]_ ) & (~\m3_data_i[28]  | ~\new_[18175]_ );
  assign \new_[14493]_  = (~\m5_data_i[28]  | ~\new_[17187]_ ) & (~\m6_data_i[28]  | ~\new_[18048]_ );
  assign \new_[14494]_  = (~\m5_data_i[27]  | ~\new_[17187]_ ) & (~\m6_data_i[27]  | ~\new_[19563]_ );
  assign \new_[14495]_  = (~\m4_data_i[26]  | ~\new_[17260]_ ) & (~\m3_data_i[26]  | ~\new_[18175]_ );
  assign \new_[14496]_  = (~\m7_data_i[25]  | ~\new_[18116]_ ) & (~\m0_data_i[25]  | ~\new_[18932]_ );
  assign \new_[14497]_  = (~\m4_data_i[25]  | ~\new_[17260]_ ) & (~\m3_data_i[25]  | ~\new_[18175]_ );
  assign \new_[14498]_  = (~\m5_data_i[25]  | ~\new_[17188]_ ) & (~\m6_data_i[25]  | ~\new_[18048]_ );
  assign \new_[14499]_  = (~\m4_data_i[24]  | ~\new_[17260]_ ) & (~\m3_data_i[24]  | ~\new_[18175]_ );
  assign \new_[14500]_  = (~\m4_data_i[23]  | ~\new_[17260]_ ) & (~\m3_data_i[23]  | ~\new_[18175]_ );
  assign \new_[14501]_  = (~\m5_data_i[23]  | ~\new_[17187]_ ) & (~\m6_data_i[23]  | ~\new_[18048]_ );
  assign \new_[14502]_  = (~\m4_data_i[22]  | ~\new_[17260]_ ) & (~\m3_data_i[22]  | ~\new_[18175]_ );
  assign \new_[14503]_  = (~\m2_addr_i[11]  | ~\new_[18119]_ ) & (~\m1_addr_i[11]  | ~\new_[18892]_ );
  assign \new_[14504]_  = ~\new_[18004]_  | ~\new_[30549]_  | ~n8344;
  assign \new_[14505]_  = (~\m2_sel_i[2]  | ~\new_[18119]_ ) & (~\m1_sel_i[2]  | ~\new_[18894]_ );
  assign \new_[14506]_  = ~\new_[17195]_  | ~\new_[30488]_  | ~n8324;
  assign \new_[14507]_  = ~\new_[16285]_  | ~\new_[31450]_  | ~n8799;
  assign \new_[14508]_  = (~\m5_data_i[19]  | ~\new_[18735]_ ) & (~\m6_data_i[19]  | ~\new_[18051]_ );
  assign \new_[14509]_  = ~m4_stb_i | ~\new_[27586]_  | ~\new_[18143]_ ;
  assign \new_[14510]_  = ~m3_stb_i | ~\new_[28766]_  | ~\new_[18201]_ ;
  assign \new_[14511]_  = ~m7_stb_i | ~\new_[26856]_  | ~\new_[18823]_ ;
  assign \new_[14512]_  = ~\new_[18070]_  | ~\new_[31463]_  | ~n8824;
  assign \new_[14513]_  = (~\m2_addr_i[14]  | ~\new_[18119]_ ) & (~\m1_addr_i[14]  | ~\new_[18891]_ );
  assign \new_[14514]_  = ~\new_[18032]_  | ~\new_[31291]_  | ~n8549;
  assign \new_[14515]_  = ~\new_[18096]_  | ~\new_[31524]_  | ~n8894;
  assign \new_[14516]_  = \new_[31235]_  ? \new_[29197]_  : \new_[18260]_ ;
  assign \new_[14517]_  = ~\new_[29752]_  & (~\new_[23840]_  | ~\new_[18354]_ );
  assign \new_[14518]_  = ~\new_[17260]_  | ~\new_[31385]_  | ~n8764;
  assign \new_[14519]_  = ~\new_[18175]_  | ~\new_[31365]_  | ~n8679;
  assign \new_[14520]_  = (~\m4_addr_i[23]  | ~\new_[19613]_ ) & (~\m3_addr_i[23]  | ~\new_[18866]_ );
  assign \new_[14521]_  = ~\new_[29278]_  & (~\new_[25150]_  | ~\new_[18357]_ );
  assign \new_[14522]_  = (~\new_[31399]_  | ~\new_[18119]_ ) & (~\m1_addr_i[3]  | ~\new_[20572]_ );
  assign \new_[14523]_  = ~\new_[29181]_  & (~\new_[18358]_  | ~\new_[27576]_ );
  assign \new_[14524]_  = ~\new_[30230]_  & (~\new_[21634]_  | ~\new_[18222]_ );
  assign \new_[14525]_  = ~\new_[29909]_  & (~\new_[20747]_  | ~\new_[18232]_ );
  assign \new_[14526]_  = ~\new_[29815]_  & (~\new_[20017]_  | ~\new_[18240]_ );
  assign \new_[14527]_  = (~\m4_data_i[1]  | ~\new_[19612]_ ) & (~\m3_data_i[1]  | ~\new_[18861]_ );
  assign \new_[14528]_  = ~\new_[29700]_  & (~\new_[20836]_  | ~\new_[18263]_ );
  assign \new_[14529]_  = (~\m4_addr_i[22]  | ~\new_[19614]_ ) & (~\m3_addr_i[22]  | ~\new_[20568]_ );
  assign \new_[14530]_  = ~\new_[29157]_  & (~\new_[20908]_  | ~\new_[18268]_ );
  assign \new_[14531]_  = ~\new_[30188]_  & (~\new_[20116]_  | ~\new_[18289]_ );
  assign \new_[14532]_  = ~\new_[30075]_  & (~\new_[20093]_  | ~\new_[18291]_ );
  assign \new_[14533]_  = (~\new_[19614]_  | ~\m4_addr_i[31] ) & (~\new_[20568]_  | ~\m3_addr_i[31] );
  assign \new_[14534]_  = (~\new_[19614]_  | ~\m4_addr_i[25] ) & (~\new_[20568]_  | ~\m3_addr_i[25] );
  assign \new_[14535]_  = (~\new_[19612]_  | ~\m4_addr_i[30] ) & (~\new_[20568]_  | ~\m3_addr_i[30] );
  assign \new_[14536]_  = ~\new_[30265]_  & (~\new_[20940]_  | ~\new_[18304]_ );
  assign \new_[14537]_  = (~\m4_data_i[19]  | ~\new_[19613]_ ) & (~\m3_data_i[19]  | ~\new_[18856]_ );
  assign \new_[14538]_  = (~\m4_addr_i[21]  | ~\new_[19614]_ ) & (~\m3_addr_i[21]  | ~\new_[18855]_ );
  assign \new_[14539]_  = ~\new_[29354]_  & (~\new_[20986]_  | ~\new_[18320]_ );
  assign \new_[14540]_  = (~\m4_data_i[26]  | ~\new_[19609]_ ) & (~\m3_data_i[26]  | ~\new_[18201]_ );
  assign \new_[14541]_  = (~\m4_addr_i[11]  | ~\new_[19613]_ ) & (~\m3_addr_i[11]  | ~\new_[20568]_ );
  assign \new_[14542]_  = \new_[18234]_  ? \new_[30660]_  : \new_[6037]_ ;
  assign \new_[14543]_  = \new_[6041]_  ? \new_[29223]_  : \new_[18235]_ ;
  assign \new_[14544]_  = (~\m5_addr_i[11]  | ~\new_[18735]_ ) & (~\m6_addr_i[11]  | ~\new_[18050]_ );
  assign \new_[14545]_  = (~\m4_data_i[20]  | ~\new_[19613]_ ) & (~\m3_data_i[20]  | ~\new_[18855]_ );
  assign \new_[14546]_  = \new_[18280]_  ? \new_[30629]_  : \new_[6043]_ ;
  assign \new_[14547]_  = \new_[31143]_  ? \new_[30604]_  : \new_[18244]_ ;
  assign \new_[14548]_  = (~\new_[18079]_  | ~\new_[31486]_ ) & (~\new_[19632]_  | ~\new_[31308]_ );
  assign \new_[14549]_  = \new_[6200]_  ? \new_[29763]_  : \new_[18252]_ ;
  assign \new_[14550]_  = \new_[18292]_  ? \new_[30662]_  : \new_[6076]_ ;
  assign \new_[14551]_  = (~\m4_data_i[27]  | ~\new_[19613]_ ) & (~\m3_data_i[27]  | ~\new_[20568]_ );
  assign \new_[14552]_  = (~\m2_data_i[6]  | ~\new_[19572]_ ) & (~\m1_data_i[6]  | ~\new_[18187]_ );
  assign \new_[14553]_  = (~\new_[18079]_  | ~\new_[31000]_ ) & (~\new_[19632]_  | ~\new_[31538]_ );
  assign \new_[14554]_  = (~\new_[19614]_  | ~\m4_addr_i[29] ) & (~\new_[18865]_  | ~\m3_addr_i[29] );
  assign \new_[14555]_  = (~\new_[18079]_  | ~\new_[31547]_ ) & (~\new_[19632]_  | ~\new_[31458]_ );
  assign \new_[14556]_  = (~\new_[19612]_  | ~\m4_addr_i[28] ) & (~\new_[18865]_  | ~\m3_addr_i[28] );
  assign \new_[14557]_  = (~\new_[18079]_  | ~\m2_addr_i[27] ) & (~\new_[19632]_  | ~\m1_addr_i[27] );
  assign \new_[14558]_  = (~\new_[19612]_  | ~\m4_addr_i[27] ) & (~\new_[18865]_  | ~\m3_addr_i[27] );
  assign \new_[14559]_  = (~\m4_addr_i[9]  | ~\new_[19613]_ ) & (~\m3_addr_i[9]  | ~\new_[20568]_ );
  assign \new_[14560]_  = (~\new_[18079]_  | ~\m2_addr_i[26] ) & (~\new_[19632]_  | ~\m1_addr_i[26] );
  assign \new_[14561]_  = (~\new_[19612]_  | ~\m4_addr_i[26] ) & (~\new_[18865]_  | ~\m3_addr_i[26] );
  assign \new_[14562]_  = (~\m4_addr_i[8]  | ~\new_[19614]_ ) & (~\m3_addr_i[8]  | ~\new_[20568]_ );
  assign \new_[14563]_  = (~\new_[18233]_  | ~\new_[30111]_ ) & (~\new_[30694]_  | ~\new_[6037]_ );
  assign \new_[14564]_  = (~\m4_addr_i[7]  | ~\new_[19613]_ ) & (~\m3_addr_i[7]  | ~\new_[20568]_ );
  assign \new_[14565]_  = (~\new_[18231]_  | ~\new_[29780]_ ) & (~\new_[30769]_  | ~\new_[6199]_ );
  assign \new_[14566]_  = (~\new_[31095]_  | ~\new_[18119]_ ) & (~\m1_addr_i[5]  | ~\new_[20572]_ );
  assign \new_[14567]_  = (~\m2_addr_i[8]  | ~\new_[18119]_ ) & (~\m1_addr_i[8]  | ~\new_[18893]_ );
  assign \new_[14568]_  = (~\m4_addr_i[6]  | ~\new_[19613]_ ) & (~\m3_addr_i[6]  | ~\new_[18856]_ );
  assign \new_[14569]_  = (~\new_[18310]_  | ~\new_[30178]_ ) & (~\new_[30696]_  | ~\new_[6194]_ );
  assign \new_[14570]_  = \new_[5988]_  ? \new_[29175]_  : \new_[18286]_ ;
  assign \new_[14571]_  = (~\m4_addr_i[5]  | ~\new_[19613]_ ) & (~\m3_addr_i[5]  | ~\new_[18859]_ );
  assign \new_[14572]_  = \new_[6189]_  ? \new_[29656]_  : \new_[18306]_ ;
  assign \new_[14573]_  = (~\new_[18270]_  | ~\new_[30343]_ ) & (~\new_[30837]_  | ~\new_[6076]_ );
  assign \new_[14574]_  = (~\m4_addr_i[4]  | ~\new_[19612]_ ) & (~\m3_addr_i[4]  | ~\new_[18862]_ );
  assign \new_[14575]_  = \new_[6185]_  ? \new_[28889]_  : \new_[18302]_ ;
  assign \new_[14576]_  = (~\m2_addr_i[3]  | ~\new_[19572]_ ) & (~\m1_addr_i[3]  | ~\new_[18191]_ );
  assign \new_[14577]_  = (~\m4_addr_i[3]  | ~\new_[19613]_ ) & (~\m3_addr_i[3]  | ~\new_[18860]_ );
  assign \new_[14578]_  = (~\m4_addr_i[2]  | ~\new_[19614]_ ) & (~\m3_addr_i[2]  | ~\new_[18864]_ );
  assign \new_[14579]_  = (~\new_[18266]_  | ~\new_[30765]_ ) & (~\new_[28568]_  | ~\new_[30765]_ );
  assign \new_[14580]_  = (~\m4_addr_i[1]  | ~\new_[19612]_ ) & (~\m3_addr_i[1]  | ~\new_[18857]_ );
  assign \new_[14581]_  = (~\new_[18315]_  | ~\new_[30707]_ ) & (~\new_[27954]_  | ~\new_[30707]_ );
  assign \new_[14582]_  = (~\m4_addr_i[0]  | ~\new_[19614]_ ) & (~\m3_addr_i[0]  | ~\new_[18857]_ );
  assign \new_[14583]_  = (~\m4_sel_i[3]  | ~\new_[19614]_ ) & (~\m3_sel_i[3]  | ~\new_[18857]_ );
  assign \new_[14584]_  = ~\new_[17253]_  & ~\new_[31563]_ ;
  assign \new_[14585]_  = ~\new_[17253]_  & ~\new_[31626]_ ;
  assign \new_[14586]_  = ~\new_[21049]_  | ~\new_[19377]_  | ~\m3_addr_i[3]  | ~\new_[21241]_ ;
  assign \new_[14587]_  = ~\new_[17252]_  | ~\m5_addr_i[3] ;
  assign \new_[14588]_  = ~\new_[17253]_  & ~\new_[31794]_ ;
  assign \new_[14589]_  = ~\new_[31793]_  & ~\new_[17253]_ ;
  assign \new_[14590]_  = (~\m4_sel_i[0]  | ~\new_[19612]_ ) & (~\m3_sel_i[0]  | ~\new_[18860]_ );
  assign \new_[14591]_  = ~\new_[17342]_  | ~\m6_addr_i[5] ;
  assign \new_[14592]_  = ~\new_[17313]_  | ~\m4_addr_i[5] ;
  assign \new_[14593]_  = ~\new_[17256]_  | ~\m1_addr_i[3] ;
  assign \new_[14594]_  = ~\new_[17326]_  | ~\m2_addr_i[3] ;
  assign \new_[14595]_  = ~\new_[17311]_  | ~\m4_addr_i[3] ;
  assign \new_[14596]_  = ~\new_[32349]_  | ~\m0_addr_i[3] ;
  assign \new_[14597]_  = (~m2_we_i | ~\new_[19572]_ ) & (~m1_we_i | ~\new_[18187]_ );
  assign \new_[14598]_  = (~m4_we_i | ~\new_[19613]_ ) & (~m3_we_i | ~\new_[18860]_ );
  assign \new_[14599]_  = (~\m2_data_i[31]  | ~\new_[18061]_ ) & (~\m1_data_i[31]  | ~\new_[18921]_ );
  assign \new_[14600]_  = (~\m2_data_i[30]  | ~\new_[18058]_ ) & (~\m1_data_i[30]  | ~\new_[18921]_ );
  assign \new_[14601]_  = (~\m2_data_i[29]  | ~\new_[18062]_ ) & (~\m1_data_i[29]  | ~\new_[18921]_ );
  assign \new_[14602]_  = (~\m2_data_i[28]  | ~\new_[18063]_ ) & (~\m1_data_i[28]  | ~\new_[20576]_ );
  assign \new_[14603]_  = (~\m2_data_i[27]  | ~\new_[18064]_ ) & (~\m1_data_i[27]  | ~\new_[18920]_ );
  assign \new_[14604]_  = \new_[22532]_  & \new_[17283]_ ;
  assign \new_[14605]_  = (~\m2_data_i[26]  | ~\new_[18058]_ ) & (~\m1_data_i[26]  | ~\new_[18922]_ );
  assign \new_[14606]_  = (~\m2_data_i[25]  | ~\new_[18058]_ ) & (~\m1_data_i[25]  | ~\new_[18921]_ );
  assign \new_[14607]_  = (~\m2_data_i[24]  | ~\new_[18062]_ ) & (~\m1_data_i[24]  | ~\new_[18920]_ );
  assign \new_[14608]_  = ~\new_[17355]_  & ~\new_[23366]_ ;
  assign \new_[14609]_  = (~\m2_data_i[23]  | ~\new_[18057]_ ) & (~\m1_data_i[23]  | ~\new_[18923]_ );
  assign \new_[14610]_  = (~\m2_data_i[22]  | ~\new_[18063]_ ) & (~\m1_data_i[22]  | ~\new_[20576]_ );
  assign \new_[14611]_  = \new_[17296]_  & \new_[31564]_ ;
  assign \new_[14612]_  = ~\new_[17357]_  & ~\new_[23398]_ ;
  assign \new_[14613]_  = (~\m2_data_i[21]  | ~\new_[18064]_ ) & (~\m1_data_i[21]  | ~\new_[20576]_ );
  assign \new_[14614]_  = (~\m2_data_i[20]  | ~\new_[18064]_ ) & (~\m1_data_i[20]  | ~\new_[20576]_ );
  assign \new_[14615]_  = ~\new_[17356]_  & ~\new_[22320]_ ;
  assign \new_[14616]_  = ~m6_stb_i | ~\new_[18794]_  | ~\new_[29036]_ ;
  assign \new_[14617]_  = (~\m2_data_i[19]  | ~\new_[18058]_ ) & (~\m1_data_i[19]  | ~\new_[18921]_ );
  assign \new_[14618]_  = \new_[17302]_  & \new_[31846]_ ;
  assign \new_[14619]_  = (~\m2_data_i[18]  | ~\new_[18054]_ ) & (~\m1_data_i[18]  | ~\new_[18922]_ );
  assign \new_[14620]_  = ~\new_[17358]_  & ~\new_[23434]_ ;
  assign \new_[14621]_  = (~\m2_data_i[17]  | ~\new_[18060]_ ) & (~\m1_data_i[17]  | ~\new_[18919]_ );
  assign \new_[14622]_  = \new_[22515]_  & \new_[17282]_ ;
  assign \new_[14623]_  = (~\m2_data_i[16]  | ~\new_[18060]_ ) & (~\m1_data_i[16]  | ~\new_[18921]_ );
  assign \new_[14624]_  = ~\new_[17306]_  | ~\new_[31810]_ ;
  assign \new_[14625]_  = \new_[17320]_  & \new_[31810]_ ;
  assign \new_[14626]_  = (~\m2_data_i[15]  | ~\new_[18065]_ ) & (~\m1_data_i[15]  | ~\new_[20576]_ );
  assign \new_[14627]_  = ~\new_[17328]_  | ~\new_[31718]_ ;
  assign \new_[14628]_  = ~m2_stb_i | ~\new_[18803]_  | ~\new_[29298]_ ;
  assign \new_[14629]_  = ~m4_stb_i | ~\new_[18881]_  | ~\new_[28767]_ ;
  assign \new_[14630]_  = (~\m2_data_i[14]  | ~\new_[18065]_ ) & (~\m1_data_i[14]  | ~\new_[20576]_ );
  assign \new_[14631]_  = ~s12_ack_i | ~\new_[17241]_  | ~\new_[29621]_ ;
  assign \new_[14632]_  = ~\new_[27638]_  & (~\new_[18367]_  | ~\new_[29401]_ );
  assign \new_[14633]_  = ~s11_ack_i | ~\new_[17229]_  | ~\new_[30284]_ ;
  assign \new_[14634]_  = ~s4_ack_i | ~\new_[17213]_  | ~\new_[29149]_ ;
  assign \new_[14635]_  = (~\m2_data_i[13]  | ~\new_[18053]_ ) & (~\m1_data_i[13]  | ~\new_[20576]_ );
  assign \new_[14636]_  = ~s7_ack_i | ~\new_[16289]_  | ~\new_[29823]_ ;
  assign \new_[14637]_  = ~s5_ack_i | ~\new_[18794]_  | ~\new_[29036]_ ;
  assign \new_[14638]_  = ~s12_err_i | ~\new_[18836]_  | ~\new_[29621]_ ;
  assign \new_[14639]_  = (~\m7_data_i[12]  | ~\new_[18835]_ ) & (~\m0_data_i[12]  | ~\new_[18937]_ );
  assign \new_[14640]_  = (~\m2_data_i[12]  | ~\new_[18053]_ ) & (~\m1_data_i[12]  | ~\new_[20576]_ );
  assign \new_[14641]_  = ~s4_err_i | ~\new_[17213]_  | ~\new_[29149]_ ;
  assign \new_[14642]_  = (~\m7_data_i[11]  | ~\new_[18835]_ ) & (~\m0_data_i[11]  | ~\new_[18937]_ );
  assign \new_[14643]_  = ~s7_err_i | ~\new_[16289]_  | ~\new_[29823]_ ;
  assign \new_[14644]_  = (~\m2_data_i[11]  | ~\new_[18065]_ ) & (~\m1_data_i[11]  | ~\new_[20576]_ );
  assign \new_[14645]_  = ~s5_rty_i | ~\new_[18794]_  | ~\new_[29036]_ ;
  assign \new_[14646]_  = ~s12_rty_i | ~\new_[17241]_  | ~\new_[29621]_ ;
  assign \new_[14647]_  = (~\m7_data_i[10]  | ~\new_[18835]_ ) & (~\m0_data_i[10]  | ~\new_[18937]_ );
  assign \new_[14648]_  = (~\m2_data_i[10]  | ~\new_[18065]_ ) & (~\m1_data_i[10]  | ~\new_[20576]_ );
  assign \new_[14649]_  = ~s4_rty_i | ~\new_[17213]_  | ~\new_[29149]_ ;
  assign \new_[14650]_  = ~s7_rty_i | ~\new_[16289]_  | ~\new_[29823]_ ;
  assign \new_[14651]_  = (~\m2_data_i[9]  | ~\new_[18053]_ ) & (~\m1_data_i[9]  | ~\new_[18918]_ );
  assign \new_[14652]_  = ~s2_ack_i | ~\new_[17215]_  | ~\new_[29788]_ ;
  assign \new_[14653]_  = ~s9_ack_i | ~\new_[17222]_  | ~\new_[29709]_ ;
  assign \new_[14654]_  = (~\m2_data_i[8]  | ~\new_[19565]_ ) & (~\m1_data_i[8]  | ~\new_[20576]_ );
  assign \new_[14655]_  = (~\m4_data_i[14]  | ~\new_[19613]_ ) & (~\m3_data_i[14]  | ~\new_[20568]_ );
  assign \new_[14656]_  = (~\m7_data_i[7]  | ~\new_[18835]_ ) & (~\m0_data_i[7]  | ~\new_[18937]_ );
  assign \new_[14657]_  = ~s1_err_i | ~\new_[18799]_  | ~\new_[30357]_ ;
  assign \new_[14658]_  = (~\m2_data_i[7]  | ~\new_[19565]_ ) & (~\m1_data_i[7]  | ~\new_[20576]_ );
  assign \new_[14659]_  = ~s13_err_i | ~\new_[18801]_  | ~\new_[32056]_ ;
  assign \new_[14660]_  = (~\m2_data_i[6]  | ~\new_[19565]_ ) & (~\m1_data_i[6]  | ~\new_[18918]_ );
  assign \new_[14661]_  = ~s9_err_i | ~\new_[17222]_  | ~\new_[29709]_ ;
  assign \new_[14662]_  = (~\m2_data_i[5]  | ~\new_[18053]_ ) & (~\m1_data_i[5]  | ~\new_[20576]_ );
  assign \new_[14663]_  = (~\m2_data_i[4]  | ~\new_[19565]_ ) & (~\m1_data_i[4]  | ~\new_[20576]_ );
  assign \new_[14664]_  = (~\m2_data_i[3]  | ~\new_[19565]_ ) & (~\m1_data_i[3]  | ~\new_[20576]_ );
  assign \new_[14665]_  = (~\m2_data_i[2]  | ~\new_[18055]_ ) & (~\m1_data_i[2]  | ~\new_[18925]_ );
  assign \new_[14666]_  = ~\new_[17362]_  & ~\new_[23608]_ ;
  assign \new_[14667]_  = (~\m2_data_i[1]  | ~\new_[19565]_ ) & (~\m1_data_i[1]  | ~\new_[18924]_ );
  assign \new_[14668]_  = (~\m2_data_i[0]  | ~\new_[18055]_ ) & (~\m1_data_i[0]  | ~\new_[18925]_ );
  assign \new_[14669]_  = (~\new_[18835]_  | ~\new_[31496]_ ) & (~\new_[20578]_  | ~\m0_addr_i[31] );
  assign \new_[14670]_  = (~\new_[18054]_  | ~\m2_addr_i[31] ) & (~\new_[20576]_  | ~\new_[31447]_ );
  assign \new_[14671]_  = ~\new_[17360]_  & ~\new_[22207]_ ;
  assign \new_[14672]_  = (~\new_[18056]_  | ~\new_[31486]_ ) & (~\new_[18923]_  | ~\new_[31308]_ );
  assign \new_[14673]_  = \new_[22498]_  & \new_[17288]_ ;
  assign \new_[14674]_  = (~\m4_addr_i[14]  | ~\new_[19612]_ ) & (~\m3_addr_i[14]  | ~\new_[18858]_ );
  assign \new_[14675]_  = (~\new_[18835]_  | ~\new_[31885]_ ) & (~\new_[18937]_  | ~\new_[31292]_ );
  assign \new_[14676]_  = (~\new_[18056]_  | ~\m2_addr_i[29] ) & (~\new_[18923]_  | ~\new_[31538]_ );
  assign \new_[14677]_  = \new_[17315]_  & \new_[31718]_ ;
  assign \new_[14678]_  = ~\new_[17361]_  & ~\new_[22232]_ ;
  assign \new_[14679]_  = \new_[23916]_  & \new_[17285]_ ;
  assign \new_[14680]_  = (~\new_[18835]_  | ~\new_[30577]_ ) & (~\new_[18937]_  | ~\new_[30957]_ );
  assign \new_[14681]_  = (~\new_[19565]_  | ~\new_[31547]_ ) & (~\new_[18918]_  | ~\new_[31458]_ );
  assign \new_[14682]_  = (~\new_[18056]_  | ~\m2_addr_i[27] ) & (~\new_[18923]_  | ~\m1_addr_i[27] );
  assign \new_[14683]_  = ~m6_stb_i | ~\new_[18836]_  | ~\new_[29621]_ ;
  assign \new_[14684]_  = (~\new_[18835]_  | ~\m7_addr_i[27] ) & (~\new_[18937]_  | ~\m0_addr_i[27] );
  assign \new_[14685]_  = \new_[17344]_  & \new_[31597]_ ;
  assign \new_[14686]_  = (~\new_[18835]_  | ~\m7_addr_i[26] ) & (~\new_[20578]_  | ~\m0_addr_i[26] );
  assign \new_[14687]_  = ~\new_[29491]_  & ~\new_[17253]_ ;
  assign \new_[14688]_  = \new_[22509]_  & \new_[17284]_ ;
  assign \new_[14689]_  = (~\m4_addr_i[2]  | ~\new_[18165]_ ) & (~\m3_addr_i[2]  | ~\new_[19636]_ );
  assign \new_[14690]_  = (~\new_[19565]_  | ~\m2_addr_i[26] ) & (~\new_[18926]_  | ~\m1_addr_i[26] );
  assign \new_[14691]_  = \new_[17298]_  & \new_[31575]_ ;
  assign \new_[14692]_  = (~\new_[18056]_  | ~\m2_addr_i[25] ) & (~\new_[18923]_  | ~\m1_addr_i[25] );
  assign \new_[14693]_  = \new_[21309]_  & \new_[17287]_ ;
  assign \new_[14694]_  = (~\new_[18835]_  | ~\m7_addr_i[25] ) & (~\new_[18937]_  | ~\m0_addr_i[25] );
  assign \new_[14695]_  = (~\new_[18835]_  | ~\m7_addr_i[24] ) & (~\new_[20578]_  | ~\m0_addr_i[24] );
  assign \new_[14696]_  = (~\new_[18054]_  | ~\m2_addr_i[24] ) & (~\new_[20576]_  | ~\m1_addr_i[24] );
  assign \new_[14697]_  = ~\new_[17354]_  & ~\new_[23747]_ ;
  assign \new_[14698]_  = (~\m2_addr_i[23]  | ~\new_[18063]_ ) & (~\m1_addr_i[23]  | ~\new_[20576]_ );
  assign \new_[14699]_  = (~\m2_addr_i[22]  | ~\new_[18063]_ ) & (~\m1_addr_i[22]  | ~\new_[18922]_ );
  assign \new_[14700]_  = (~\m7_addr_i[22]  | ~\new_[18835]_ ) & (~\m0_addr_i[22]  | ~\new_[18937]_ );
  assign \new_[14701]_  = \new_[21284]_  & \new_[17286]_ ;
  assign \new_[14702]_  = (~\m2_addr_i[21]  | ~\new_[18061]_ ) & (~\m1_addr_i[21]  | ~\new_[18920]_ );
  assign \new_[14703]_  = (~\m2_addr_i[20]  | ~\new_[18061]_ ) & (~\m1_addr_i[20]  | ~\new_[18922]_ );
  assign \new_[14704]_  = ~s3_ack_i | ~\new_[17260]_  | ~\new_[30457]_ ;
  assign \new_[14705]_  = ~s5_ack_i | ~\new_[19608]_  | ~\new_[28768]_ ;
  assign \new_[14706]_  = ~s8_ack_i | ~\new_[17263]_  | ~\new_[29627]_ ;
  assign \new_[14707]_  = ~s13_ack_i | ~\new_[17266]_  | ~\new_[28851]_ ;
  assign \new_[14708]_  = (~\m2_addr_i[19]  | ~\new_[18059]_ ) & (~\m1_addr_i[19]  | ~\new_[20576]_ );
  assign \new_[14709]_  = ~s7_ack_i | ~\new_[18882]_  | ~\new_[28223]_ ;
  assign \new_[14710]_  = (~\m4_data_i[15]  | ~\new_[19613]_ ) & (~\m3_data_i[15]  | ~\new_[18859]_ );
  assign \new_[14711]_  = ~s0_ack_i | ~\new_[16309]_  | ~\new_[29349]_ ;
  assign \new_[14712]_  = (~\m2_addr_i[18]  | ~\new_[18059]_ ) & (~\m1_addr_i[18]  | ~\new_[20576]_ );
  assign \new_[14713]_  = ~s3_err_i | ~\new_[17260]_  | ~\new_[30457]_ ;
  assign \new_[14714]_  = ~s13_err_i | ~\new_[17266]_  | ~\new_[28851]_ ;
  assign \new_[14715]_  = ~s0_err_i | ~\new_[17271]_  | ~\new_[29349]_ ;
  assign \new_[14716]_  = (~\m7_addr_i[17]  | ~\new_[18835]_ ) & (~\m0_addr_i[17]  | ~\new_[20578]_ );
  assign \new_[14717]_  = ~s7_err_i | ~\new_[18882]_  | ~\new_[28223]_ ;
  assign \new_[14718]_  = ~s3_rty_i | ~\new_[17260]_  | ~\new_[30457]_ ;
  assign \new_[14719]_  = ~s8_rty_i | ~\new_[17263]_  | ~\new_[29627]_ ;
  assign \new_[14720]_  = (~\m2_addr_i[17]  | ~\new_[19565]_ ) & (~\m1_addr_i[17]  | ~\new_[18926]_ );
  assign \new_[14721]_  = ~s13_rty_i | ~\new_[17266]_  | ~\new_[28851]_ ;
  assign \new_[14722]_  = ~s0_rty_i | ~\new_[17270]_  | ~\new_[29349]_ ;
  assign \new_[14723]_  = (~\m7_addr_i[16]  | ~\new_[18835]_ ) & (~\m0_addr_i[16]  | ~\new_[20578]_ );
  assign \new_[14724]_  = (~\m2_addr_i[16]  | ~\new_[18064]_ ) & (~\m1_addr_i[16]  | ~\new_[20576]_ );
  assign \new_[14725]_  = ~s7_rty_i | ~\new_[18882]_  | ~\new_[28223]_ ;
  assign \new_[14726]_  = (~\m7_addr_i[15]  | ~\new_[18835]_ ) & (~\m0_addr_i[15]  | ~\new_[20578]_ );
  assign \new_[14727]_  = (~\m2_addr_i[15]  | ~\new_[18062]_ ) & (~\m1_addr_i[15]  | ~\new_[18922]_ );
  assign \new_[14728]_  = (~\m7_addr_i[14]  | ~\new_[18835]_ ) & (~\m0_addr_i[14]  | ~\new_[19642]_ );
  assign \new_[14729]_  = (~\m2_addr_i[14]  | ~\new_[18062]_ ) & (~\m1_addr_i[14]  | ~\new_[20576]_ );
  assign \new_[14730]_  = (~\m2_addr_i[13]  | ~\new_[18057]_ ) & (~\m1_addr_i[13]  | ~\new_[18923]_ );
  assign \new_[14731]_  = ~m4_stb_i | ~\new_[17260]_  | ~\new_[30457]_ ;
  assign \new_[14732]_  = ~\new_[17359]_  & ~\new_[22189]_ ;
  assign \new_[14733]_  = (~\m4_data_i[21]  | ~\new_[18163]_ ) & (~\m3_data_i[21]  | ~\new_[18198]_ );
  assign \new_[14734]_  = (~\m2_addr_i[12]  | ~\new_[19565]_ ) & (~\m1_addr_i[12]  | ~\new_[18926]_ );
  assign \new_[14735]_  = (~\m2_addr_i[11]  | ~\new_[18060]_ ) & (~\m1_addr_i[11]  | ~\new_[18920]_ );
  assign \new_[14736]_  = (~\m2_addr_i[10]  | ~\new_[18059]_ ) & (~\m1_addr_i[10]  | ~\new_[18920]_ );
  assign \new_[14737]_  = (~\m2_addr_i[9]  | ~\new_[18057]_ ) & (~\m1_addr_i[9]  | ~\new_[18923]_ );
  assign \new_[14738]_  = (~\m2_addr_i[8]  | ~\new_[18055]_ ) & (~\m1_addr_i[8]  | ~\new_[18925]_ );
  assign \new_[14739]_  = (~\m7_addr_i[8]  | ~\new_[18835]_ ) & (~\m0_addr_i[8]  | ~\new_[18937]_ );
  assign \new_[14740]_  = (~\m2_addr_i[7]  | ~\new_[19565]_ ) & (~\m1_addr_i[7]  | ~\new_[18926]_ );
  assign \new_[14741]_  = (~\m2_addr_i[6]  | ~\new_[18055]_ ) & (~\m1_addr_i[6]  | ~\new_[18925]_ );
  assign \new_[14742]_  = ~s3_ack_i | ~\new_[18735]_  | ~\new_[29928]_ ;
  assign \new_[14743]_  = ~s5_ack_i | ~\new_[18871]_  | ~\new_[28136]_ ;
  assign \new_[14744]_  = ~s14_ack_i | ~\new_[17192]_  | ~\new_[30181]_ ;
  assign \new_[14745]_  = ~s1_ack_i | ~\new_[18738]_  | ~\new_[29769]_ ;
  assign \new_[14746]_  = ~s13_ack_i | ~\new_[17194]_  | ~\new_[32267]_ ;
  assign \new_[14747]_  = (~\m7_addr_i[5]  | ~\new_[18835]_ ) & (~\new_[31848]_  | ~\new_[18937]_ );
  assign \new_[14748]_  = (~\new_[31095]_  | ~\new_[19565]_ ) & (~\m1_addr_i[5]  | ~\new_[20576]_ );
  assign \new_[14749]_  = ~s8_ack_i | ~\new_[17204]_  | ~\new_[29636]_ ;
  assign \new_[14750]_  = ~s1_err_i | ~\new_[18738]_  | ~\new_[29769]_ ;
  assign \new_[14751]_  = ~s2_err_i | ~\new_[18740]_  | ~\new_[30013]_ ;
  assign \new_[14752]_  = ~s14_err_i | ~\new_[17192]_  | ~\new_[30181]_ ;
  assign \new_[14753]_  = (~\m2_addr_i[4]  | ~\new_[18055]_ ) & (~\m1_addr_i[4]  | ~\new_[18925]_ );
  assign \new_[14754]_  = ~s13_err_i | ~\new_[17194]_  | ~\new_[32267]_ ;
  assign \new_[14755]_  = ~s2_rty_i | ~\new_[18740]_  | ~\new_[30013]_ ;
  assign \new_[14756]_  = ~s8_rty_i | ~\new_[17204]_  | ~\new_[29636]_ ;
  assign \new_[14757]_  = (~\new_[31399]_  | ~\new_[19565]_ ) & (~\m1_addr_i[3]  | ~\new_[18924]_ );
  assign \new_[14758]_  = ~s14_rty_i | ~\new_[17192]_  | ~\new_[30181]_ ;
  assign \new_[14759]_  = ~\new_[20334]_  & (~\new_[18368]_  | ~\new_[26322]_ );
  assign \new_[14760]_  = (~\m7_addr_i[2]  | ~\new_[18835]_ ) & (~\m0_addr_i[2]  | ~\new_[20578]_ );
  assign \new_[14761]_  = (~\m2_addr_i[2]  | ~\new_[19565]_ ) & (~\m1_addr_i[2]  | ~\new_[20576]_ );
  assign \new_[14762]_  = ~\new_[21562]_  & (~\new_[18374]_  | ~\new_[26328]_ );
  assign \new_[14763]_  = (~\m2_addr_i[1]  | ~\new_[18059]_ ) & (~\m1_addr_i[1]  | ~\new_[18922]_ );
  assign \new_[14764]_  = ~m5_stb_i | ~\new_[18871]_  | ~\new_[28136]_ ;
  assign \new_[14765]_  = (~\m2_addr_i[0]  | ~\new_[18057]_ ) & (~\m1_addr_i[0]  | ~\new_[18923]_ );
  assign \new_[14766]_  = (~\m7_addr_i[0]  | ~\new_[18835]_ ) & (~\m0_addr_i[0]  | ~\new_[18937]_ );
  assign \new_[14767]_  = ~\new_[22416]_  & (~\new_[18372]_  | ~\new_[23046]_ );
  assign \new_[14768]_  = ~\new_[23391]_  & (~\new_[18376]_  | ~\new_[24792]_ );
  assign \new_[14769]_  = ~\new_[22186]_  & (~\new_[18369]_  | ~\new_[24745]_ );
  assign \new_[14770]_  = ~m1_stb_i | ~\new_[17274]_  | ~\new_[29052]_ ;
  assign \new_[14771]_  = (~\m2_sel_i[3]  | ~\new_[18060]_ ) & (~\m1_sel_i[3]  | ~\new_[18920]_ );
  assign \new_[14772]_  = ~m5_stb_i | ~\new_[18007]_  | ~\new_[29704]_ ;
  assign \new_[14773]_  = ~\new_[21181]_  & (~\new_[18370]_  | ~\new_[24632]_ );
  assign \new_[14774]_  = ~\new_[17346]_  | ~\new_[27706]_ ;
  assign \new_[14775]_  = ~s6_rty_i | ~\new_[18207]_  | ~\new_[29939]_ ;
  assign \new_[14776]_  = (~\m2_sel_i[2]  | ~\new_[19565]_ ) & (~\m1_sel_i[2]  | ~\new_[18924]_ );
  assign \new_[14777]_  = ~\new_[27985]_  | ~\new_[18066]_  | ~m0_stb_i;
  assign \new_[14778]_  = ~m7_stb_i | ~\new_[18832]_  | ~\new_[28313]_ ;
  assign \new_[14779]_  = ~\new_[22245]_  & (~\new_[18371]_  | ~\new_[27525]_ );
  assign \new_[14780]_  = (~\m2_sel_i[1]  | ~\new_[18061]_ ) & (~\m1_sel_i[1]  | ~\new_[18919]_ );
  assign \new_[14781]_  = (~\m7_sel_i[1]  | ~\new_[18835]_ ) & (~\m0_sel_i[1]  | ~\new_[18937]_ );
  assign \new_[14782]_  = (~\m2_sel_i[0]  | ~\new_[19565]_ ) & (~\m1_sel_i[0]  | ~\new_[18924]_ );
  assign \new_[14783]_  = ~m5_stb_i | ~\new_[17204]_  | ~\new_[29636]_ ;
  assign \new_[14784]_  = ~s2_ack_i | ~\new_[18824]_  | ~\new_[30113]_ ;
  assign \new_[14785]_  = ~s0_ack_i | ~\new_[18826]_  | ~\new_[27879]_ ;
  assign \new_[14786]_  = ~s3_ack_i | ~\new_[18116]_  | ~\new_[29579]_ ;
  assign \new_[14787]_  = (~\m4_addr_i[19]  | ~\new_[19613]_ ) & (~\m3_addr_i[19]  | ~\new_[20568]_ );
  assign \new_[14788]_  = ~s3_err_i | ~\new_[18116]_  | ~\new_[29579]_ ;
  assign \new_[14789]_  = (~m2_we_i | ~\new_[19565]_ ) & (~m1_we_i | ~\new_[18924]_ );
  assign \new_[14790]_  = ~s2_err_i | ~\new_[18824]_  | ~\new_[30113]_ ;
  assign \new_[14791]_  = ~m1_stb_i | ~\new_[18906]_  | ~\new_[30354]_ ;
  assign \new_[14792]_  = ~m3_stb_i | ~\new_[17249]_  | ~\new_[29024]_ ;
  assign \new_[14793]_  = ~\new_[21206]_  & (~\new_[18375]_  | ~\new_[26226]_ );
  assign \new_[14794]_  = ~\new_[17324]_  | ~\new_[24348]_ ;
  assign \new_[14795]_  = ~m5_stb_i | ~\new_[17201]_  | ~\new_[29045]_ ;
  assign \new_[14796]_  = ~s0_rty_i | ~\new_[18826]_  | ~\new_[27879]_ ;
  assign \new_[14797]_  = ~s11_err_i | ~\new_[18930]_  | ~\new_[30200]_ ;
  assign \new_[14798]_  = (~\m2_data_i[28]  | ~\new_[18803]_ ) & (~\m1_data_i[28]  | ~\new_[18910]_ );
  assign \new_[14799]_  = ~\new_[17331]_  | ~\new_[26169]_ ;
  assign \new_[14800]_  = ~s14_rty_i | ~\new_[18927]_  | ~\new_[30166]_ ;
  assign \new_[14801]_  = ~m3_stb_i | ~\new_[18928]_  | ~\new_[30200]_ ;
  assign \new_[14802]_  = ~s3_rty_i | ~\new_[18116]_  | ~\new_[29579]_ ;
  assign \new_[14803]_  = ~\new_[17339]_  | ~\new_[23059]_ ;
  assign \new_[14804]_  = ~m7_stb_i | ~\new_[18114]_  | ~\new_[32338]_ ;
  assign \new_[14805]_  = ~\new_[28726]_  | ~\new_[18020]_  | ~m0_stb_i;
  assign \new_[14806]_  = ~m1_stb_i | ~\new_[18905]_  | ~\new_[32327]_ ;
  assign \new_[14807]_  = ~m5_stb_i | ~\new_[18737]_  | ~\new_[30181]_ ;
  assign \new_[14808]_  = ~m3_stb_i | ~\new_[17280]_  | ~\new_[30166]_ ;
  assign \new_[14809]_  = ~m5_stb_i | ~\new_[18740]_  | ~\new_[30013]_ ;
  assign \new_[14810]_  = ~s14_ack_i | ~\new_[17280]_  | ~\new_[30166]_ ;
  assign \new_[14811]_  = ~s8_ack_i | ~\new_[18846]_  | ~\new_[29428]_ ;
  assign \new_[14812]_  = ~s11_rty_i | ~\new_[18930]_  | ~\new_[30200]_ ;
  assign \new_[14813]_  = ~\new_[21248]_  & (~\new_[18373]_  | ~\new_[27705]_ );
  assign \new_[14814]_  = ~m5_stb_i | ~\new_[18735]_  | ~\new_[29928]_ ;
  assign \new_[14815]_  = ~m7_stb_i | ~\new_[18116]_  | ~\new_[29579]_ ;
  assign \new_[14816]_  = ~s14_err_i | ~\new_[17280]_  | ~\new_[30166]_ ;
  assign \new_[14817]_  = (~\m2_data_i[9]  | ~\new_[18803]_ ) & (~\m1_data_i[9]  | ~\new_[18180]_ );
  assign \new_[14818]_  = ~\new_[24940]_  & (~\new_[18380]_  | ~\new_[27846]_ );
  assign \new_[14819]_  = ~\new_[25014]_  & (~\new_[18381]_  | ~\new_[22891]_ );
  assign \new_[14820]_  = (~\m2_data_i[8]  | ~\new_[18803]_ ) & (~\m1_data_i[8]  | ~\new_[18910]_ );
  assign \new_[14821]_  = (~\m2_data_i[17]  | ~\new_[18074]_ ) & (~\m1_data_i[17]  | ~\new_[18908]_ );
  assign \new_[14822]_  = ~\new_[30297]_  | ~\new_[17185]_  | ~\new_[21343]_ ;
  assign \new_[14823]_  = ~\new_[29020]_  | ~\new_[17183]_  | ~\new_[22258]_ ;
  assign \new_[14824]_  = (~\m2_data_i[3]  | ~\new_[18803]_ ) & (~\m1_data_i[3]  | ~\new_[18910]_ );
  assign \new_[14825]_  = (~\m2_data_i[22]  | ~\new_[18119]_ ) & (~\m1_data_i[22]  | ~\new_[20572]_ );
  assign \new_[14826]_  = (~\m2_data_i[1]  | ~\new_[18803]_ ) & (~\m1_data_i[1]  | ~\new_[18180]_ );
  assign \new_[14827]_  = (~\m4_data_i[16]  | ~\new_[19612]_ ) & (~\m3_data_i[16]  | ~\new_[18858]_ );
  assign \new_[14828]_  = (~\new_[18086]_  | ~\m6_addr_i[29] ) & (~\new_[18007]_  | ~\new_[31407]_ );
  assign \new_[14829]_  = (~\m2_addr_i[22]  | ~\new_[18803]_ ) & (~\m1_addr_i[22]  | ~\new_[18180]_ );
  assign \new_[14830]_  = ~\new_[31990]_ ;
  assign \new_[14831]_  = (~\m2_data_i[25]  | ~\new_[18119]_ ) & (~\m1_data_i[25]  | ~\new_[18891]_ );
  assign \new_[14832]_  = (~\m2_addr_i[15]  | ~\new_[18803]_ ) & (~\m1_addr_i[15]  | ~\new_[18910]_ );
  assign \new_[14833]_  = ~\new_[19372]_  & ~\new_[17363]_ ;
  assign \new_[14834]_  = ~\new_[17207]_ ;
  assign \new_[14835]_  = (~\m4_data_i[17]  | ~\new_[19613]_ ) & (~\m3_data_i[17]  | ~\new_[20568]_ );
  assign \new_[14836]_  = ~\new_[17212]_ ;
  assign \new_[14837]_  = ~\new_[19569]_ ;
  assign \new_[14838]_  = ~\new_[19372]_  & ~\new_[17366]_ ;
  assign \new_[14839]_  = ~\new_[16293]_ ;
  assign \new_[14840]_  = (~\m2_sel_i[2]  | ~\new_[18803]_ ) & (~\m1_sel_i[2]  | ~\new_[18180]_ );
  assign \new_[14841]_  = (~\m2_data_i[30]  | ~\new_[18805]_ ) & (~\m1_data_i[30]  | ~\new_[18912]_ );
  assign \new_[14842]_  = (~\m2_data_i[29]  | ~\new_[18804]_ ) & (~\m1_data_i[29]  | ~\new_[18912]_ );
  assign \new_[14843]_  = (~\m2_data_i[28]  | ~\new_[18805]_ ) & (~\m1_data_i[28]  | ~\new_[18912]_ );
  assign \new_[14844]_  = ~\new_[20353]_  & ~\new_[17366]_ ;
  assign \new_[14845]_  = (~\m2_data_i[27]  | ~\new_[18804]_ ) & (~\m1_data_i[27]  | ~\new_[18913]_ );
  assign \new_[14846]_  = (~\m2_data_i[26]  | ~\new_[18804]_ ) & (~\m1_data_i[26]  | ~\new_[18913]_ );
  assign \new_[14847]_  = (~\m2_data_i[25]  | ~\new_[20555]_ ) & (~\m1_data_i[25]  | ~\new_[18913]_ );
  assign \new_[14848]_  = ~\new_[16302]_ ;
  assign \new_[14849]_  = ~\new_[16302]_ ;
  assign \new_[14850]_  = ~\new_[16302]_ ;
  assign \new_[14851]_  = (~\m2_data_i[24]  | ~\new_[20555]_ ) & (~\m1_data_i[24]  | ~\new_[18912]_ );
  assign \new_[14852]_  = \new_[16303]_ ;
  assign \new_[14853]_  = (~\m2_data_i[23]  | ~\new_[20555]_ ) & (~\m1_data_i[23]  | ~\new_[18912]_ );
  assign \new_[14854]_  = (~\m2_data_i[21]  | ~\new_[20555]_ ) & (~\m1_data_i[21]  | ~\new_[18912]_ );
  assign \new_[14855]_  = (~\m2_data_i[20]  | ~\new_[18804]_ ) & (~\m1_data_i[20]  | ~\new_[18912]_ );
  assign \new_[14856]_  = \new_[20353]_  & \new_[17367]_ ;
  assign \new_[14857]_  = (~\m2_data_i[19]  | ~\new_[18804]_ ) & (~\m1_data_i[19]  | ~\new_[18913]_ );
  assign \new_[14858]_  = (~\m2_data_i[17]  | ~\new_[18804]_ ) & (~\m1_data_i[17]  | ~\new_[18912]_ );
  assign \new_[14859]_  = (~\m2_data_i[16]  | ~\new_[18805]_ ) & (~\m1_data_i[16]  | ~\new_[18912]_ );
  assign \new_[14860]_  = \new_[5992]_  ? \new_[29893]_  : \new_[18226]_ ;
  assign \new_[14861]_  = ~\new_[20353]_  & ~\new_[17363]_ ;
  assign \new_[14862]_  = (~\m2_data_i[12]  | ~\new_[20555]_ ) & (~\m1_data_i[12]  | ~\new_[18912]_ );
  assign \new_[14863]_  = (~\m2_data_i[10]  | ~\new_[20555]_ ) & (~\m1_data_i[10]  | ~\new_[18912]_ );
  assign \new_[14864]_  = (~\m2_data_i[8]  | ~\new_[18804]_ ) & (~\m1_data_i[8]  | ~\new_[18912]_ );
  assign \new_[14865]_  = (~\m2_data_i[7]  | ~\new_[18804]_ ) & (~\m1_data_i[7]  | ~\new_[18912]_ );
  assign \new_[14866]_  = (~\m2_sel_i[1]  | ~\new_[18074]_ ) & (~\m1_sel_i[1]  | ~\new_[18909]_ );
  assign \new_[14867]_  = (~\m2_data_i[1]  | ~\new_[18805]_ ) & (~\m1_data_i[1]  | ~\new_[18912]_ );
  assign \new_[14868]_  = (~\m4_data_i[18]  | ~\new_[19615]_ ) & (~\m3_data_i[18]  | ~\new_[18198]_ );
  assign \new_[14869]_  = (~\m5_sel_i[0]  | ~\new_[18735]_ ) & (~\m6_sel_i[0]  | ~\new_[19563]_ );
  assign \new_[14870]_  = (~\new_[18805]_  | ~\new_[31486]_ ) & (~\new_[18912]_  | ~\new_[31308]_ );
  assign \new_[14871]_  = (~\m4_data_i[18]  | ~\new_[19613]_ ) & (~\m3_data_i[18]  | ~\new_[18856]_ );
  assign \new_[14872]_  = (~\new_[18079]_  | ~\m2_addr_i[25] ) & (~\new_[19632]_  | ~\m1_addr_i[25] );
  assign \new_[14873]_  = (~\new_[18805]_  | ~\new_[31547]_ ) & (~\new_[18913]_  | ~\new_[31458]_ );
  assign \new_[14874]_  = (~\new_[18805]_  | ~\m2_addr_i[27] ) & (~\new_[18912]_  | ~\m1_addr_i[27] );
  assign \new_[14875]_  = (~\new_[20555]_  | ~\m2_addr_i[26] ) & (~\new_[18913]_  | ~\m1_addr_i[26] );
  assign \new_[14876]_  = \new_[18295]_  ? \new_[30710]_  : \new_[6073]_ ;
  assign \new_[14877]_  = (~\new_[20555]_  | ~\m2_addr_i[24] ) & (~\new_[18913]_  | ~\m1_addr_i[24] );
  assign \new_[14878]_  = ~\new_[16316]_ ;
  assign \new_[14879]_  = (~\m2_addr_i[23]  | ~\new_[18804]_ ) & (~\m1_addr_i[23]  | ~\new_[18912]_ );
  assign \new_[14880]_  = ~\new_[16316]_ ;
  assign \new_[14881]_  = (~\m2_addr_i[22]  | ~\new_[18804]_ ) & (~\m1_addr_i[22]  | ~\new_[18912]_ );
  assign \new_[14882]_  = (~\m2_addr_i[21]  | ~\new_[18805]_ ) & (~\m1_addr_i[21]  | ~\new_[18912]_ );
  assign \new_[14883]_  = (~\m2_addr_i[20]  | ~\new_[18804]_ ) & (~\m1_addr_i[20]  | ~\new_[18913]_ );
  assign \new_[14884]_  = (~\m2_addr_i[19]  | ~\new_[18805]_ ) & (~\m1_addr_i[19]  | ~\new_[18912]_ );
  assign \new_[14885]_  = (~\m4_addr_i[12]  | ~\new_[19615]_ ) & (~\m3_addr_i[12]  | ~\new_[18198]_ );
  assign \new_[14886]_  = (~\m2_addr_i[18]  | ~\new_[18804]_ ) & (~\m1_addr_i[18]  | ~\new_[18913]_ );
  assign \new_[14887]_  = (~\m2_addr_i[17]  | ~\new_[18804]_ ) & (~\m1_addr_i[17]  | ~\new_[18912]_ );
  assign \new_[14888]_  = ~\new_[16322]_ ;
  assign \new_[14889]_  = (~\m4_data_i[3]  | ~\new_[19613]_ ) & (~\m3_data_i[3]  | ~\new_[18861]_ );
  assign \new_[14890]_  = (~\m2_addr_i[12]  | ~\new_[18804]_ ) & (~\m1_addr_i[12]  | ~\new_[18913]_ );
  assign \new_[14891]_  = (~\m2_addr_i[11]  | ~\new_[20555]_ ) & (~\m1_addr_i[11]  | ~\new_[18912]_ );
  assign \new_[14892]_  = (~\m2_addr_i[10]  | ~\new_[18805]_ ) & (~\m1_addr_i[10]  | ~\new_[18912]_ );
  assign \new_[14893]_  = (~\m2_addr_i[9]  | ~\new_[18804]_ ) & (~\m1_addr_i[9]  | ~\new_[18913]_ );
  assign \new_[14894]_  = (~\m4_data_i[21]  | ~\new_[19613]_ ) & (~\m3_data_i[21]  | ~\new_[20568]_ );
  assign \new_[14895]_  = ~\new_[16326]_ ;
  assign \new_[14896]_  = (~\m2_addr_i[0]  | ~\new_[18805]_ ) & (~\m1_addr_i[0]  | ~\new_[18912]_ );
  assign \new_[14897]_  = (~\m4_addr_i[15]  | ~\new_[19612]_ ) & (~\m3_addr_i[15]  | ~\new_[18855]_ );
  assign \new_[14898]_  = (~\m2_sel_i[3]  | ~\new_[18804]_ ) & (~\m1_sel_i[3]  | ~\new_[18913]_ );
  assign \new_[14899]_  = (~\m2_sel_i[2]  | ~\new_[18804]_ ) & (~\m1_sel_i[2]  | ~\new_[18913]_ );
  assign \new_[14900]_  = (~\m2_sel_i[1]  | ~\new_[18804]_ ) & (~\m1_sel_i[1]  | ~\new_[18913]_ );
  assign \new_[14901]_  = (~\new_[18079]_  | ~\m2_addr_i[31] ) & (~\new_[19632]_  | ~\new_[31447]_ );
  assign \new_[14902]_  = (~\m4_data_i[29]  | ~\new_[19613]_ ) & (~\m3_data_i[29]  | ~\new_[20568]_ );
  assign \new_[14903]_  = (~\m4_data_i[7]  | ~\new_[19613]_ ) & (~\m3_data_i[7]  | ~\new_[18862]_ );
  assign \new_[14904]_  = (~\m4_data_i[12]  | ~\new_[19612]_ ) & (~\m3_data_i[12]  | ~\new_[18864]_ );
  assign \new_[14905]_  = ~\new_[17387]_  | ~\new_[28002]_ ;
  assign \new_[14906]_  = ~\new_[17390]_  | ~\new_[29091]_ ;
  assign \new_[14907]_  = ~\new_[17391]_  | ~\new_[28741]_ ;
  assign \new_[14908]_  = ~\new_[17392]_  | ~\new_[30369]_ ;
  assign \new_[14909]_  = ~\new_[17393]_  | ~\new_[29121]_ ;
  assign \new_[14910]_  = ~\new_[17395]_  | ~\new_[28679]_ ;
  assign \new_[14911]_  = ~\new_[17396]_  | ~\new_[28717]_ ;
  assign \new_[14912]_  = (~\m4_addr_i[20]  | ~\new_[19614]_ ) & (~\m3_addr_i[20]  | ~\new_[18858]_ );
  assign \new_[14913]_  = ~\new_[17565]_  | ~\new_[29448]_  | ~\new_[24192]_ ;
  assign \new_[14914]_  = (~\m4_data_i[5]  | ~\new_[19613]_ ) & (~\m3_data_i[5]  | ~\new_[18864]_ );
  assign \new_[14915]_  = ~\new_[17566]_  | ~\new_[29454]_  | ~\new_[24226]_ ;
  assign \new_[14916]_  = ~\new_[30115]_  & (~\new_[21937]_  | ~\new_[18317]_ );
  assign \new_[14917]_  = ~\new_[17567]_  | ~\new_[28218]_  | ~\new_[25248]_ ;
  assign \new_[14918]_  = (~\m5_addr_i[10]  | ~\new_[18735]_ ) & (~\m6_addr_i[10]  | ~\new_[18049]_ );
  assign \new_[14919]_  = ~\new_[17568]_  | ~\new_[27642]_  | ~\new_[21451]_ ;
  assign \new_[14920]_  = \new_[6213]_  ? \new_[30243]_  : \new_[18258]_ ;
  assign \new_[14921]_  = ~\new_[17569]_  | ~\new_[28634]_  | ~\new_[25658]_ ;
  assign \new_[14922]_  = ~\new_[17570]_  | ~\new_[29499]_  | ~\new_[24099]_ ;
  assign \new_[14923]_  = (~\m2_data_i[3]  | ~\new_[19572]_ ) & (~\m1_data_i[3]  | ~\new_[18191]_ );
  assign \new_[14924]_  = ~\new_[17571]_  | ~\new_[28540]_  | ~\new_[24233]_ ;
  assign \new_[14925]_  = ~\new_[17572]_  | ~\new_[27648]_  | ~\new_[22739]_ ;
  assign \new_[14926]_  = (~\m2_addr_i[12]  | ~\new_[18075]_ ) & (~\m1_addr_i[12]  | ~\new_[20575]_ );
  assign \new_[14927]_  = ~\new_[17573]_  | ~\new_[29413]_  | ~\new_[24252]_ ;
  assign \new_[14928]_  = ~\new_[17401]_  & ~\new_[28558]_ ;
  assign \new_[14929]_  = ~\new_[17574]_  | ~\new_[28838]_  | ~\new_[24006]_ ;
  assign \new_[14930]_  = \new_[17415]_  | \new_[24854]_ ;
  assign \new_[14931]_  = ~\new_[17575]_  | ~\new_[29464]_  | ~\new_[26184]_ ;
  assign \new_[14932]_  = ~\new_[18450]_  | ~\new_[27730]_  | ~\new_[21398]_ ;
  assign \new_[14933]_  = ~\new_[18442]_  | ~\new_[29448]_  | ~\new_[24242]_ ;
  assign \new_[14934]_  = ~\new_[18443]_  | ~\new_[25013]_  | ~\new_[22702]_ ;
  assign \new_[14935]_  = ~\new_[18444]_  | ~\new_[27676]_  | ~\new_[22575]_ ;
  assign \new_[14936]_  = ~\new_[18445]_  | ~\new_[26120]_  | ~\new_[24237]_ ;
  assign \new_[14937]_  = (~\m4_addr_i[3]  | ~\new_[18164]_ ) & (~\m3_addr_i[3]  | ~\new_[19636]_ );
  assign \new_[14938]_  = ~\new_[18446]_  | ~\new_[29454]_  | ~\new_[24207]_ ;
  assign \new_[14939]_  = ~\new_[18447]_  | ~\new_[24094]_  | ~\new_[24204]_ ;
  assign \new_[14940]_  = ~\new_[18448]_  | ~\new_[28218]_  | ~\new_[26160]_ ;
  assign \new_[14941]_  = ~\new_[18449]_  | ~\new_[24438]_  | ~\new_[22844]_ ;
  assign \new_[14942]_  = (~\m2_data_i[18]  | ~\new_[18799]_ ) & (~\m1_data_i[18]  | ~\new_[18887]_ );
  assign \new_[14943]_  = ~\new_[18453]_  | ~\new_[28634]_  | ~\new_[26161]_ ;
  assign \new_[14944]_  = ~\new_[18454]_  | ~\new_[26423]_  | ~\new_[21361]_ ;
  assign \new_[14945]_  = ~\new_[18455]_  | ~\new_[29499]_  | ~\new_[24228]_ ;
  assign \new_[14946]_  = ~\new_[18456]_  | ~\new_[24722]_  | ~\new_[22646]_ ;
  assign \new_[14947]_  = (~\m4_data_i[8]  | ~\new_[19613]_ ) & (~\m3_data_i[8]  | ~\new_[18859]_ );
  assign \new_[14948]_  = (~\m2_data_i[21]  | ~\new_[18806]_ ) & (~\m1_data_i[21]  | ~\new_[18177]_ );
  assign \new_[14949]_  = ~\new_[18457]_  | ~\new_[28324]_  | ~\new_[22749]_ ;
  assign \new_[14950]_  = ~\new_[18458]_  | ~\new_[26210]_  | ~\new_[20436]_ ;
  assign \new_[14951]_  = (~\m2_data_i[10]  | ~\new_[18806]_ ) & (~\m1_data_i[10]  | ~\new_[18177]_ );
  assign \new_[14952]_  = ~\new_[18460]_  | ~\new_[28838]_  | ~\new_[23984]_ ;
  assign \new_[14953]_  = ~\new_[18461]_  | ~\new_[27669]_  | ~\new_[22710]_ ;
  assign \new_[14954]_  = (~\m2_data_i[7]  | ~\new_[18806]_ ) & (~\m1_data_i[7]  | ~\new_[18177]_ );
  assign \new_[14955]_  = (~\m2_data_i[2]  | ~\new_[18806]_ ) & (~\m1_data_i[2]  | ~\new_[18177]_ );
  assign \new_[14956]_  = (~\m4_data_i[0]  | ~\new_[18160]_ ) & (~\m3_data_i[0]  | ~\new_[18199]_ );
  assign \new_[14957]_  = ~\new_[18462]_  | ~\new_[28142]_  | ~\new_[22843]_ ;
  assign \new_[14958]_  = (~\new_[18451]_  | ~\new_[27792]_ ) & (~\new_[21375]_  | ~\new_[27792]_ );
  assign \new_[14959]_  = (~\m4_data_i[0]  | ~\new_[19613]_ ) & (~\m3_data_i[0]  | ~\new_[18862]_ );
  assign \new_[14960]_  = (~\m2_addr_i[12]  | ~\new_[18806]_ ) & (~\m1_addr_i[12]  | ~\new_[18177]_ );
  assign \new_[14961]_  = ~\new_[28055]_  & (~\new_[17592]_  | ~\new_[24472]_ );
  assign \new_[14962]_  = (~\m4_addr_i[16]  | ~\new_[19613]_ ) & (~\m3_addr_i[16]  | ~\new_[18855]_ );
  assign \new_[14963]_  = (~\m2_data_i[5]  | ~\new_[19572]_ ) & (~\m1_data_i[5]  | ~\new_[18187]_ );
  assign \new_[14964]_  = ~\new_[24667]_  & (~\new_[17594]_  | ~\new_[24497]_ );
  assign \new_[14965]_  = ~\new_[24573]_  & (~\new_[17595]_  | ~\new_[23204]_ );
  assign \new_[14966]_  = ~\new_[28095]_  & (~\new_[17582]_  | ~\new_[20479]_ );
  assign \new_[14967]_  = ~\new_[24568]_  & (~\new_[17596]_  | ~\new_[24349]_ );
  assign \new_[14968]_  = ~\new_[27988]_  & (~\new_[17597]_  | ~\new_[24409]_ );
  assign \new_[14969]_  = ~\new_[30187]_  & (~\new_[17593]_  | ~\new_[24309]_ );
  assign \new_[14970]_  = (~\m2_data_i[31]  | ~\new_[18075]_ ) & (~\m1_data_i[31]  | ~\new_[19630]_ );
  assign \new_[14971]_  = (~\m5_data_i[30]  | ~\new_[19544]_ ) & (~\m6_data_i[30]  | ~\new_[19561]_ );
  assign \new_[14972]_  = ~\new_[29552]_  & (~\new_[17598]_  | ~\new_[23171]_ );
  assign \new_[14973]_  = (~\m2_data_i[29]  | ~\new_[18075]_ ) & (~\m1_data_i[29]  | ~\new_[19630]_ );
  assign \new_[14974]_  = (~\m4_data_i[24]  | ~\new_[19613]_ ) & (~\m3_data_i[24]  | ~\new_[20568]_ );
  assign \new_[14975]_  = (~\m7_data_i[29]  | ~\new_[19606]_ ) & (~\m0_data_i[29]  | ~\new_[18781]_ );
  assign \new_[14976]_  = (~\m5_data_i[28]  | ~\new_[19544]_ ) & (~\m6_data_i[28]  | ~\new_[19561]_ );
  assign \new_[14977]_  = (~\m7_data_i[27]  | ~\new_[19606]_ ) & (~\m0_data_i[27]  | ~\new_[18781]_ );
  assign \new_[14978]_  = (~\m4_sel_i[3]  | ~\new_[18163]_ ) & (~\m3_sel_i[3]  | ~\new_[18198]_ );
  assign \new_[14979]_  = ~\new_[28769]_  & (~\new_[17599]_  | ~\new_[24323]_ );
  assign \new_[14980]_  = (~\m2_data_i[25]  | ~\new_[18074]_ ) & (~\m1_data_i[25]  | ~\new_[20575]_ );
  assign \new_[14981]_  = (~\m2_data_i[24]  | ~\new_[18074]_ ) & (~\m1_data_i[24]  | ~\new_[18908]_ );
  assign \new_[14982]_  = (~\m2_data_i[23]  | ~\new_[18075]_ ) & (~\m1_data_i[23]  | ~\new_[20575]_ );
  assign \new_[14983]_  = (~\m7_data_i[23]  | ~\new_[19606]_ ) & (~\m0_data_i[23]  | ~\new_[18781]_ );
  assign \new_[14984]_  = (~\m2_data_i[22]  | ~\new_[18074]_ ) & (~\m1_data_i[22]  | ~\new_[19629]_ );
  assign \new_[14985]_  = (~\m7_data_i[21]  | ~\new_[19606]_ ) & (~\m0_data_i[21]  | ~\new_[18781]_ );
  assign \new_[14986]_  = (~\m7_data_i[20]  | ~\new_[19606]_ ) & (~\m0_data_i[20]  | ~\new_[20547]_ );
  assign \new_[14987]_  = (~\m2_data_i[20]  | ~\new_[18074]_ ) & (~\m1_data_i[20]  | ~\new_[18909]_ );
  assign \new_[14988]_  = (~\m2_data_i[19]  | ~\new_[18075]_ ) & (~\m1_data_i[19]  | ~\new_[19630]_ );
  assign \new_[14989]_  = (~\m5_data_i[19]  | ~\new_[19544]_ ) & (~\m6_data_i[19]  | ~\new_[19561]_ );
  assign \new_[14990]_  = (~\m7_data_i[18]  | ~\new_[19606]_ ) & (~\m0_data_i[18]  | ~\new_[20547]_ );
  assign \new_[14991]_  = (~\m2_data_i[18]  | ~\new_[18074]_ ) & (~\m1_data_i[18]  | ~\new_[20575]_ );
  assign \new_[14992]_  = (~\new_[18806]_  | ~\m2_addr_i[26] ) & (~\new_[18177]_  | ~\m1_addr_i[26] );
  assign \new_[14993]_  = ~\new_[30066]_  & (~\new_[21827]_  | ~\new_[18284]_ );
  assign \new_[14994]_  = (~\m2_data_i[16]  | ~\new_[18074]_ ) & (~\m1_data_i[16]  | ~\new_[19630]_ );
  assign \new_[14995]_  = (~\m7_data_i[13]  | ~\new_[19606]_ ) & (~\m0_data_i[13]  | ~\new_[20547]_ );
  assign \new_[14996]_  = (~\m2_data_i[13]  | ~\new_[18074]_ ) & (~\m1_data_i[13]  | ~\new_[18909]_ );
  assign \new_[14997]_  = ~\new_[26529]_  & (~\new_[17600]_  | ~\new_[23594]_ );
  assign \new_[14998]_  = (~\m7_data_i[12]  | ~\new_[19606]_ ) & (~\m0_data_i[12]  | ~\new_[18781]_ );
  assign \new_[14999]_  = \new_[18319]_  ? \new_[30591]_  : \new_[6186]_ ;
  assign \new_[15000]_  = (~\m2_data_i[11]  | ~\new_[18075]_ ) & (~\m1_data_i[11]  | ~\new_[20575]_ );
  assign \new_[15001]_  = (~\m7_data_i[11]  | ~\new_[19606]_ ) & (~\m0_data_i[11]  | ~\new_[18781]_ );
  assign \new_[15002]_  = (~\m7_data_i[10]  | ~\new_[19606]_ ) & (~\m0_data_i[10]  | ~\new_[20547]_ );
  assign \new_[15003]_  = (~\m2_data_i[10]  | ~\new_[18074]_ ) & (~\m1_data_i[10]  | ~\new_[18908]_ );
  assign \new_[15004]_  = (~\m7_data_i[9]  | ~\new_[19606]_ ) & (~\m0_data_i[9]  | ~\new_[20547]_ );
  assign \new_[15005]_  = (~\m2_data_i[9]  | ~\new_[18074]_ ) & (~\m1_data_i[9]  | ~\new_[18908]_ );
  assign \new_[15006]_  = (~\m2_data_i[8]  | ~\new_[18075]_ ) & (~\m1_data_i[8]  | ~\new_[20575]_ );
  assign \new_[15007]_  = (~\m7_data_i[8]  | ~\new_[19606]_ ) & (~\m0_data_i[8]  | ~\new_[18781]_ );
  assign \new_[15008]_  = (~\m2_data_i[7]  | ~\new_[18075]_ ) & (~\m1_data_i[7]  | ~\new_[20575]_ );
  assign \new_[15009]_  = (~\m7_data_i[7]  | ~\new_[19606]_ ) & (~\m0_data_i[7]  | ~\new_[18781]_ );
  assign \new_[15010]_  = (~\m4_data_i[28]  | ~\new_[18162]_ ) & (~\m3_data_i[28]  | ~\new_[19636]_ );
  assign \new_[15011]_  = (~\m2_data_i[6]  | ~\new_[18074]_ ) & (~\m1_data_i[6]  | ~\new_[18908]_ );
  assign \new_[15012]_  = (~\m2_data_i[5]  | ~\new_[18074]_ ) & (~\m1_data_i[5]  | ~\new_[18908]_ );
  assign \new_[15013]_  = (~\m7_data_i[4]  | ~\new_[19606]_ ) & (~\m0_data_i[4]  | ~\new_[18781]_ );
  assign \new_[15014]_  = (~\m7_data_i[3]  | ~\new_[19606]_ ) & (~\m0_data_i[3]  | ~\new_[20547]_ );
  assign \new_[15015]_  = (~\m7_data_i[2]  | ~\new_[19606]_ ) & (~\m0_data_i[2]  | ~\new_[18781]_ );
  assign \new_[15016]_  = (~\m2_data_i[1]  | ~\new_[18074]_ ) & (~\m1_data_i[1]  | ~\new_[19630]_ );
  assign \new_[15017]_  = (~\m4_addr_i[17]  | ~\new_[19613]_ ) & (~\m3_addr_i[17]  | ~\new_[20568]_ );
  assign \new_[15018]_  = (~\new_[18789]_  | ~\m6_addr_i[31] ) & (~\new_[19544]_  | ~\new_[31001]_ );
  assign \new_[15019]_  = (~\new_[19606]_  | ~\m7_addr_i[31] ) & (~\new_[20547]_  | ~\m0_addr_i[31] );
  assign \new_[15020]_  = (~\m4_data_i[23]  | ~\new_[19613]_ ) & (~\m3_data_i[23]  | ~\new_[18856]_ );
  assign \new_[15021]_  = (~\new_[19606]_  | ~\new_[31531]_ ) & (~\new_[20547]_  | ~\new_[31481]_ );
  assign \new_[15022]_  = (~\new_[18074]_  | ~\m2_addr_i[29] ) & (~\new_[20575]_  | ~\new_[31538]_ );
  assign \new_[15023]_  = (~\new_[20551]_  | ~\m6_addr_i[28] ) & (~\new_[19544]_  | ~\new_[31276]_ );
  assign \new_[15024]_  = (~\new_[18074]_  | ~\m2_addr_i[27] ) & (~\new_[18909]_  | ~\m1_addr_i[27] );
  assign \new_[15025]_  = (~\new_[20551]_  | ~\m6_addr_i[26] ) & (~\new_[19544]_  | ~\m5_addr_i[26] );
  assign \new_[15026]_  = (~\new_[18074]_  | ~\m2_addr_i[25] ) & (~\new_[20575]_  | ~\m1_addr_i[25] );
  assign \new_[15027]_  = (~\m2_addr_i[22]  | ~\new_[18075]_ ) & (~\m1_addr_i[22]  | ~\new_[19630]_ );
  assign \new_[15028]_  = ~\new_[30010]_  & (~\new_[20138]_  | ~\new_[18278]_ );
  assign \new_[15029]_  = (~\m7_addr_i[22]  | ~\new_[19606]_ ) & (~\m0_addr_i[22]  | ~\new_[19557]_ );
  assign \new_[15030]_  = ~\new_[23356]_  & (~\new_[17860]_  | ~\new_[30296]_ );
  assign \new_[15031]_  = (~\m2_addr_i[21]  | ~\new_[18074]_ ) & (~\m1_addr_i[21]  | ~\new_[19630]_ );
  assign \new_[15032]_  = (~\m2_addr_i[20]  | ~\new_[18075]_ ) & (~\m1_addr_i[20]  | ~\new_[19630]_ );
  assign \new_[15033]_  = (~\m7_addr_i[20]  | ~\new_[19606]_ ) & (~\m0_addr_i[20]  | ~\new_[19557]_ );
  assign \new_[15034]_  = ~\new_[22172]_  & (~\new_[17864]_  | ~\new_[28837]_ );
  assign \new_[15035]_  = (~\m7_addr_i[19]  | ~\new_[19606]_ ) & (~\m0_addr_i[19]  | ~\new_[19557]_ );
  assign \new_[15036]_  = ~\new_[23556]_  & (~\new_[17881]_  | ~\new_[29015]_ );
  assign \new_[15037]_  = (~\m2_addr_i[18]  | ~\new_[18074]_ ) & (~\m1_addr_i[18]  | ~\new_[18909]_ );
  assign \new_[15038]_  = (~\m7_addr_i[17]  | ~\new_[19606]_ ) & (~\m0_addr_i[17]  | ~\new_[20547]_ );
  assign \new_[15039]_  = ~\new_[21217]_  & (~\new_[17875]_  | ~\new_[29978]_ );
  assign \new_[15040]_  = (~\m2_addr_i[17]  | ~\new_[18074]_ ) & (~\m1_addr_i[17]  | ~\new_[18908]_ );
  assign \new_[15041]_  = (~\m2_addr_i[16]  | ~\new_[18074]_ ) & (~\m1_addr_i[16]  | ~\new_[19629]_ );
  assign \new_[15042]_  = (~\m7_addr_i[16]  | ~\new_[19606]_ ) & (~\m0_addr_i[16]  | ~\new_[19557]_ );
  assign \new_[15043]_  = ~\new_[21188]_  & (~\new_[17891]_  | ~\new_[28188]_ );
  assign \new_[15044]_  = (~\m2_addr_i[15]  | ~\new_[18075]_ ) & (~\m1_addr_i[15]  | ~\new_[19630]_ );
  assign \new_[15045]_  = (~\m7_addr_i[15]  | ~\new_[19606]_ ) & (~\m0_addr_i[15]  | ~\new_[18781]_ );
  assign \new_[15046]_  = (~\m2_addr_i[14]  | ~\new_[18074]_ ) & (~\m1_addr_i[14]  | ~\new_[18909]_ );
  assign \new_[15047]_  = ~\new_[23793]_  & (~\new_[17894]_  | ~\new_[29996]_ );
  assign \new_[15048]_  = (~\m2_addr_i[13]  | ~\new_[18074]_ ) & (~\m1_addr_i[13]  | ~\new_[19629]_ );
  assign \new_[15049]_  = ~\new_[17525]_  & ~\new_[23887]_ ;
  assign \new_[15050]_  = (~\m7_addr_i[13]  | ~\new_[19606]_ ) & (~\m0_addr_i[13]  | ~\new_[18781]_ );
  assign \new_[15051]_  = ~\new_[30097]_  | ~\new_[17531]_  | ~\new_[28908]_ ;
  assign \new_[15052]_  = ~\new_[16722]_  & ~\new_[28992]_ ;
  assign \new_[15053]_  = ~\new_[17439]_  | ~\new_[27898]_ ;
  assign \new_[15054]_  = (~\m2_addr_i[11]  | ~\new_[18074]_ ) & (~\m1_addr_i[11]  | ~\new_[20575]_ );
  assign \new_[15055]_  = ~\new_[30320]_  | ~\new_[17532]_  | ~\new_[29112]_ ;
  assign \new_[15056]_  = (~\m4_addr_i[18]  | ~\new_[19613]_ ) & (~\m3_addr_i[18]  | ~\new_[18866]_ );
  assign \new_[15057]_  = ~\new_[16723]_  & ~\new_[29541]_ ;
  assign \new_[15058]_  = (~\m2_addr_i[10]  | ~\new_[18075]_ ) & (~\m1_addr_i[10]  | ~\new_[19630]_ );
  assign \new_[15059]_  = ~\new_[17443]_  | ~\new_[27231]_ ;
  assign \new_[15060]_  = (~\m5_addr_i[10]  | ~\new_[19544]_ ) & (~\m6_addr_i[10]  | ~\new_[19561]_ );
  assign \new_[15061]_  = (~\m2_addr_i[9]  | ~\new_[18075]_ ) & (~\m1_addr_i[9]  | ~\new_[19630]_ );
  assign \new_[15062]_  = ~\new_[30172]_  | ~\new_[17536]_  | ~\new_[28968]_ ;
  assign \new_[15063]_  = (~\m5_addr_i[9]  | ~\new_[19544]_ ) & (~\m6_addr_i[9]  | ~\new_[19561]_ );
  assign \new_[15064]_  = ~\new_[16724]_  & ~\new_[29217]_ ;
  assign \new_[15065]_  = ~\new_[17447]_  | ~\new_[26803]_ ;
  assign \new_[15066]_  = (~\m2_addr_i[8]  | ~\new_[18074]_ ) & (~\m1_addr_i[8]  | ~\new_[18907]_ );
  assign \new_[15067]_  = (~\m7_addr_i[8]  | ~\new_[19606]_ ) & (~\m0_addr_i[8]  | ~\new_[20547]_ );
  assign \new_[15068]_  = ~\new_[22904]_  & (~\new_[17694]_  | ~\new_[29168]_ );
  assign \new_[15069]_  = (~\m5_addr_i[8]  | ~\new_[19544]_ ) & (~\m6_addr_i[8]  | ~\new_[19561]_ );
  assign \new_[15070]_  = (~\m7_addr_i[7]  | ~\new_[19606]_ ) & (~\m0_addr_i[7]  | ~\new_[20547]_ );
  assign \new_[15071]_  = (~\m2_addr_i[7]  | ~\new_[18074]_ ) & (~\m1_addr_i[7]  | ~\new_[18908]_ );
  assign \new_[15072]_  = ~\new_[17452]_  | ~\new_[26192]_ ;
  assign \new_[15073]_  = (~\m2_addr_i[6]  | ~\new_[18074]_ ) & (~\m1_addr_i[6]  | ~\new_[18907]_ );
  assign \new_[15074]_  = ~\new_[19445]_  & (~\new_[17705]_  | ~\new_[29397]_ );
  assign \new_[15075]_  = ~\new_[22930]_  & (~\new_[17712]_  | ~\new_[30497]_ );
  assign \new_[15076]_  = (~\m7_addr_i[6]  | ~\new_[19606]_ ) & (~\m0_addr_i[6]  | ~\new_[20547]_ );
  assign \new_[15077]_  = ~\new_[17538]_  & ~\new_[23901]_ ;
  assign \new_[15078]_  = (~\new_[31095]_  | ~\new_[18075]_ ) & (~\m1_addr_i[5]  | ~\new_[20575]_ );
  assign \new_[15079]_  = ~\new_[17382]_  & ~\new_[29700]_ ;
  assign \new_[15080]_  = (~\m7_addr_i[4]  | ~\new_[19606]_ ) & (~\m0_addr_i[4]  | ~\new_[18781]_ );
  assign \new_[15081]_  = ~\new_[17463]_  | ~\new_[24256]_ ;
  assign \new_[15082]_  = (~\m2_addr_i[3]  | ~\new_[18074]_ ) & (~\m1_addr_i[3]  | ~\new_[18909]_ );
  assign \new_[15083]_  = ~\new_[22913]_  & (~\new_[17747]_  | ~\new_[29271]_ );
  assign \new_[15084]_  = ~\new_[22596]_  & (~\new_[17753]_  | ~\new_[30627]_ );
  assign \new_[15085]_  = (~\m7_addr_i[3]  | ~\new_[19606]_ ) & (~\new_[31884]_  | ~\new_[18781]_ );
  assign \new_[15086]_  = (~\m2_addr_i[2]  | ~\new_[18074]_ ) & (~\new_[31477]_  | ~\new_[18909]_ );
  assign \new_[15087]_  = ~\new_[17384]_  & ~\new_[29157]_ ;
  assign \new_[15088]_  = ~\new_[17469]_  | ~\new_[24295]_ ;
  assign \new_[15089]_  = (~\m7_addr_i[2]  | ~\new_[19606]_ ) & (~\m0_addr_i[2]  | ~\new_[20547]_ );
  assign \new_[15090]_  = ~\new_[21486]_  & (~\new_[17762]_  | ~\new_[28877]_ );
  assign \new_[15091]_  = (~\m5_addr_i[2]  | ~\new_[19544]_ ) & (~\m6_addr_i[2]  | ~\new_[20551]_ );
  assign \new_[15092]_  = ~\new_[23011]_  & (~\new_[17763]_  | ~\new_[30329]_ );
  assign \new_[15093]_  = (~\m7_addr_i[1]  | ~\new_[19606]_ ) & (~\m0_addr_i[1]  | ~\new_[20547]_ );
  assign \new_[15094]_  = ~\new_[17476]_  | ~\new_[26247]_ ;
  assign \new_[15095]_  = (~\m5_addr_i[1]  | ~\new_[19544]_ ) & (~\m6_addr_i[1]  | ~\new_[19561]_ );
  assign \new_[15096]_  = ~\new_[22972]_  & (~\new_[17807]_  | ~\new_[28930]_ );
  assign \new_[15097]_  = (~\m2_addr_i[0]  | ~\new_[18075]_ ) & (~\m1_addr_i[0]  | ~\new_[20575]_ );
  assign \new_[15098]_  = (~\m7_addr_i[0]  | ~\new_[19606]_ ) & (~\m0_addr_i[0]  | ~\new_[18781]_ );
  assign \new_[15099]_  = ~\new_[29888]_  | ~\new_[17544]_  | ~\new_[29633]_ ;
  assign \new_[15100]_  = ~\new_[17480]_  | ~\new_[26437]_ ;
  assign \new_[15101]_  = (~\m7_sel_i[3]  | ~\new_[19606]_ ) & (~\m0_sel_i[3]  | ~\new_[19557]_ );
  assign \new_[15102]_  = ~\new_[21478]_  & (~\new_[17776]_  | ~\new_[28285]_ );
  assign \new_[15103]_  = ~\new_[29863]_  | ~\new_[17546]_  | ~\new_[28864]_ ;
  assign \new_[15104]_  = ~\new_[16731]_  & ~\new_[29101]_ ;
  assign \new_[15105]_  = (~\m2_sel_i[2]  | ~\new_[18075]_ ) & (~\m1_sel_i[2]  | ~\new_[19630]_ );
  assign \new_[15106]_  = (~\m7_sel_i[2]  | ~\new_[19606]_ ) & (~\m0_sel_i[2]  | ~\new_[20547]_ );
  assign \new_[15107]_  = ~\new_[17484]_  | ~\new_[27609]_ ;
  assign \new_[15108]_  = (~\m7_sel_i[1]  | ~\new_[19606]_ ) & (~\m0_sel_i[1]  | ~\new_[20547]_ );
  assign \new_[15109]_  = ~\new_[30061]_  | ~\new_[17547]_  | ~\new_[28844]_ ;
  assign \new_[15110]_  = (~\m7_addr_i[5]  | ~\new_[19606]_ ) & (~\m0_addr_i[5]  | ~\new_[20547]_ );
  assign \new_[15111]_  = ~\new_[17490]_  | ~\new_[26211]_ ;
  assign \new_[15112]_  = ~\new_[22971]_  & (~\new_[17787]_  | ~\new_[28985]_ );
  assign \new_[15113]_  = (~\m7_sel_i[0]  | ~\new_[19606]_ ) & (~\m0_sel_i[0]  | ~\new_[20547]_ );
  assign \new_[15114]_  = (~m2_we_i | ~\new_[18074]_ ) & (~m1_we_i | ~\new_[19629]_ );
  assign \new_[15115]_  = ~\new_[17364]_  & ~\new_[29671]_ ;
  assign \new_[15116]_  = ~\new_[23117]_  & (~\new_[17823]_  | ~\new_[29608]_ );
  assign \new_[15117]_  = ~\new_[30159]_  | ~\new_[17554]_  | ~\new_[29189]_ ;
  assign \new_[15118]_  = ~\new_[16733]_  & ~\new_[29167]_ ;
  assign \new_[15119]_  = ~\new_[17496]_  | ~\new_[27703]_ ;
  assign \new_[15120]_  = ~\new_[22854]_  & (~\new_[17826]_  | ~\new_[29817]_ );
  assign \new_[15121]_  = ~\new_[16734]_  & ~\new_[29047]_ ;
  assign \new_[15122]_  = (~\m2_data_i[31]  | ~\new_[18119]_ ) & (~\m1_data_i[31]  | ~\new_[18891]_ );
  assign \new_[15123]_  = ~\new_[17499]_  | ~\new_[24440]_ ;
  assign \new_[15124]_  = ~\new_[23031]_  & (~\new_[17710]_  | ~\new_[30411]_ );
  assign \new_[15125]_  = (~\m2_data_i[29]  | ~\new_[18119]_ ) & (~\m1_data_i[29]  | ~\new_[18891]_ );
  assign \new_[15126]_  = ~\new_[16736]_  & ~\new_[29354]_ ;
  assign \new_[15127]_  = ~\new_[17505]_  | ~\new_[24316]_ ;
  assign \new_[15128]_  = (~\m2_data_i[28]  | ~\new_[18119]_ ) & (~\m1_data_i[28]  | ~\new_[18891]_ );
  assign \new_[15129]_  = (~\m4_data_i[22]  | ~\new_[19613]_ ) & (~\m3_data_i[22]  | ~\new_[20568]_ );
  assign \new_[15130]_  = (~\m2_data_i[27]  | ~\new_[19590]_ ) & (~\m1_data_i[27]  | ~\new_[18892]_ );
  assign \new_[15131]_  = ~\new_[16738]_  & ~\new_[29172]_ ;
  assign \new_[15132]_  = ~\new_[17434]_  & ~\new_[24601]_ ;
  assign \new_[15133]_  = (~\m4_data_i[26]  | ~\new_[19614]_ ) & (~\m3_data_i[26]  | ~\new_[20568]_ );
  assign \new_[15134]_  = (~\m2_data_i[26]  | ~\new_[18119]_ ) & (~\m1_data_i[26]  | ~\new_[18896]_ );
  assign \new_[15135]_  = ~\new_[16394]_ ;
  assign \new_[15136]_  = ~\new_[16395]_ ;
  assign \new_[15137]_  = ~\new_[16396]_ ;
  assign \new_[15138]_  = (~\m2_data_i[24]  | ~\new_[18119]_ ) & (~\m1_data_i[24]  | ~\new_[18896]_ );
  assign \new_[15139]_  = ~\new_[25088]_  & (~\new_[17664]_  | ~\new_[29527]_ );
  assign \new_[15140]_  = \new_[16741]_  | \new_[26250]_ ;
  assign \new_[15141]_  = (~\m2_data_i[14]  | ~\new_[18074]_ ) & (~\m1_data_i[14]  | ~\new_[20575]_ );
  assign \new_[15142]_  = (~\m2_data_i[23]  | ~\new_[18119]_ ) & (~\m1_data_i[23]  | ~\new_[18891]_ );
  assign \new_[15143]_  = ~\new_[23015]_  & (~\new_[17670]_  | ~\new_[25315]_ );
  assign \new_[15144]_  = ~\new_[24305]_  & (~\new_[17671]_  | ~\new_[26924]_ );
  assign \new_[15145]_  = ~\new_[23375]_  & (~\new_[17672]_  | ~\new_[29220]_ );
  assign \new_[15146]_  = (~\m2_data_i[21]  | ~\new_[18119]_ ) & (~\m1_data_i[21]  | ~\new_[18891]_ );
  assign \new_[15147]_  = ~\new_[24840]_  & (~\new_[17675]_  | ~\new_[29320]_ );
  assign \new_[15148]_  = \new_[16743]_  | \new_[25351]_ ;
  assign \new_[15149]_  = (~\m2_data_i[20]  | ~\new_[18119]_ ) & (~\m1_data_i[20]  | ~\new_[18891]_ );
  assign \new_[15150]_  = ~\new_[24260]_  & (~\new_[17682]_  | ~\new_[24043]_ );
  assign \new_[15151]_  = ~\new_[21148]_  & (~\new_[17683]_  | ~\new_[30386]_ );
  assign \new_[15152]_  = (~\m2_data_i[19]  | ~\new_[18119]_ ) & (~\m1_data_i[19]  | ~\new_[18891]_ );
  assign \new_[15153]_  = ~\new_[27958]_  & (~\new_[17684]_  | ~\new_[23127]_ );
  assign \new_[15154]_  = ~\new_[21611]_  & (~\new_[17686]_  | ~\new_[26372]_ );
  assign \new_[15155]_  = ~\new_[24864]_  & (~\new_[17688]_  | ~\new_[29228]_ );
  assign \new_[15156]_  = \new_[16744]_  | \new_[26206]_ ;
  assign \new_[15157]_  = (~\m2_data_i[17]  | ~\new_[18119]_ ) & (~\m1_data_i[17]  | ~\new_[18894]_ );
  assign \new_[15158]_  = ~\new_[22904]_  & (~\new_[17695]_  | ~\new_[24367]_ );
  assign \new_[15159]_  = ~\new_[16400]_ ;
  assign \new_[15160]_  = (~\m2_data_i[16]  | ~\new_[18119]_ ) & (~\m1_data_i[16]  | ~\new_[18891]_ );
  assign \new_[15161]_  = ~\new_[22919]_  & (~\new_[17696]_  | ~\new_[27508]_ );
  assign \new_[15162]_  = ~\new_[22187]_  & (~\new_[17698]_  | ~\new_[29103]_ );
  assign \new_[15163]_  = (~\m2_data_i[15]  | ~\new_[18119]_ ) & (~\m1_data_i[15]  | ~\new_[20572]_ );
  assign \new_[15164]_  = \new_[16745]_  | \new_[24812]_ ;
  assign \new_[15165]_  = (~\m2_data_i[14]  | ~\new_[19590]_ ) & (~\m1_data_i[14]  | ~\new_[20572]_ );
  assign \new_[15166]_  = (~\m2_data_i[13]  | ~\new_[19590]_ ) & (~\m1_data_i[13]  | ~\new_[20572]_ );
  assign \new_[15167]_  = ~\new_[24351]_  & (~\new_[17715]_  | ~\new_[24314]_ );
  assign \new_[15168]_  = ~\new_[22930]_  & (~\new_[17719]_  | ~\new_[27952]_ );
  assign \new_[15169]_  = \new_[16747]_  | \new_[24744]_ ;
  assign \new_[15170]_  = ~\new_[17458]_  & ~\new_[23491]_ ;
  assign \new_[15171]_  = (~\m2_data_i[12]  | ~\new_[18119]_ ) & (~\m1_data_i[12]  | ~\new_[20572]_ );
  assign \new_[15172]_  = ~\new_[23873]_  & (~\new_[17733]_  | ~\new_[30728]_ );
  assign \new_[15173]_  = ~\new_[26382]_  & (~\new_[17734]_  | ~\new_[24340]_ );
  assign \new_[15174]_  = (~\m2_data_i[11]  | ~\new_[18119]_ ) & (~\m1_data_i[11]  | ~\new_[18895]_ );
  assign \new_[15175]_  = (~\m2_data_i[10]  | ~\new_[18119]_ ) & (~\m1_data_i[10]  | ~\new_[20572]_ );
  assign \new_[15176]_  = ~\new_[16403]_ ;
  assign \new_[15177]_  = ~\new_[22112]_  & (~\new_[17737]_  | ~\new_[30617]_ );
  assign \new_[15178]_  = ~\new_[22618]_  & (~\new_[17748]_  | ~\new_[24354]_ );
  assign \new_[15179]_  = ~\new_[22913]_  & (~\new_[17749]_  | ~\new_[27782]_ );
  assign \new_[15180]_  = (~\m2_data_i[8]  | ~\new_[18119]_ ) & (~\m1_data_i[8]  | ~\new_[20572]_ );
  assign \new_[15181]_  = ~\new_[24427]_  & (~\new_[17754]_  | ~\new_[26198]_ );
  assign \new_[15182]_  = ~\new_[22596]_  & (~\new_[17755]_  | ~\new_[26863]_ );
  assign \new_[15183]_  = (~\m2_data_i[7]  | ~\new_[19590]_ ) & (~\m1_data_i[7]  | ~\new_[18892]_ );
  assign \new_[15184]_  = ~\new_[23555]_  & (~\new_[17798]_  | ~\new_[29967]_ );
  assign \new_[15185]_  = \new_[16750]_  | \new_[27581]_ ;
  assign \new_[15186]_  = (~\m2_data_i[6]  | ~\new_[18119]_ ) & (~\m1_data_i[6]  | ~\new_[20572]_ );
  assign \new_[15187]_  = ~\new_[21486]_  & (~\new_[17727]_  | ~\new_[24386]_ );
  assign \new_[15188]_  = ~\new_[24372]_  & (~\new_[17764]_  | ~\new_[24376]_ );
  assign \new_[15189]_  = (~\m2_data_i[5]  | ~\new_[19590]_ ) & (~\m1_data_i[5]  | ~\new_[20572]_ );
  assign \new_[15190]_  = ~\new_[23011]_  & (~\new_[17765]_  | ~\new_[26323]_ );
  assign \new_[15191]_  = \new_[16752]_  | \new_[26393]_ ;
  assign \new_[15192]_  = ~\new_[22270]_  & (~\new_[17766]_  | ~\new_[28963]_ );
  assign \new_[15193]_  = (~\m2_data_i[4]  | ~\new_[19590]_ ) & (~\m1_data_i[4]  | ~\new_[20572]_ );
  assign \new_[15194]_  = \new_[16753]_  | \new_[26204]_ ;
  assign \new_[15195]_  = (~\m2_data_i[30]  | ~\new_[18119]_ ) & (~\m1_data_i[30]  | ~\new_[20572]_ );
  assign \new_[15196]_  = ~\new_[22972]_  & (~\new_[17800]_  | ~\new_[24510]_ );
  assign \new_[15197]_  = ~\new_[21229]_  & (~\new_[17772]_  | ~\new_[29506]_ );
  assign \new_[15198]_  = (~\m2_data_i[3]  | ~\new_[18119]_ ) & (~\m1_data_i[3]  | ~\new_[20572]_ );
  assign \new_[15199]_  = ~\new_[16408]_ ;
  assign \new_[15200]_  = (~\m2_data_i[2]  | ~\new_[18119]_ ) & (~\m1_data_i[2]  | ~\new_[20572]_ );
  assign \new_[15201]_  = (~\m2_data_i[1]  | ~\new_[18119]_ ) & (~\m1_data_i[1]  | ~\new_[18895]_ );
  assign \new_[15202]_  = ~\new_[22289]_  & (~\new_[17661]_  | ~\new_[29721]_ );
  assign \new_[15203]_  = \new_[16754]_  | \new_[26200]_ ;
  assign \new_[15204]_  = (~\m2_data_i[0]  | ~\new_[18119]_ ) & (~\m1_data_i[0]  | ~\new_[18895]_ );
  assign \new_[15205]_  = ~\new_[21478]_  & (~\new_[17791]_  | ~\new_[26266]_ );
  assign \new_[15206]_  = ~\new_[22295]_  & (~\new_[17777]_  | ~\new_[29974]_ );
  assign \new_[15207]_  = (~\new_[19590]_  | ~\m2_addr_i[31] ) & (~\new_[18892]_  | ~\new_[31447]_ );
  assign \new_[15208]_  = ~\new_[16411]_ ;
  assign \new_[15209]_  = ~\new_[16412]_ ;
  assign \new_[15210]_  = (~\new_[18119]_  | ~\new_[31486]_ ) & (~\new_[18892]_  | ~\new_[31308]_ );
  assign \new_[15211]_  = ~\new_[25000]_  & (~\new_[17781]_  | ~\new_[29006]_ );
  assign \new_[15212]_  = \new_[16755]_  | \new_[24768]_ ;
  assign \new_[15213]_  = (~\new_[18119]_  | ~\m2_addr_i[29] ) & (~\new_[18892]_  | ~\new_[31538]_ );
  assign \new_[15214]_  = ~\new_[21468]_  & (~\new_[17804]_  | ~\new_[22980]_ );
  assign \new_[15215]_  = ~\new_[22896]_  & (~\new_[17783]_  | ~\new_[26334]_ );
  assign \new_[15216]_  = (~\new_[18119]_  | ~\new_[31547]_ ) & (~\new_[18892]_  | ~\new_[31458]_ );
  assign \new_[15217]_  = (~\new_[18119]_  | ~\m2_addr_i[27] ) & (~\new_[18893]_  | ~\m1_addr_i[27] );
  assign \new_[15218]_  = ~\new_[23037]_  & (~\new_[17785]_  | ~\new_[26404]_ );
  assign \new_[15219]_  = \new_[16756]_  | \new_[26450]_ ;
  assign \new_[15220]_  = ~\new_[22140]_  & (~\new_[17689]_  | ~\new_[29695]_ );
  assign \new_[15221]_  = \new_[16757]_  | \new_[26233]_ ;
  assign \new_[15222]_  = ~\new_[23001]_  & (~\new_[17788]_  | ~\new_[22934]_ );
  assign \new_[15223]_  = (~\new_[18119]_  | ~\m2_addr_i[26] ) & (~\new_[18892]_  | ~\m1_addr_i[26] );
  assign \new_[15224]_  = ~\new_[22971]_  & (~\new_[17751]_  | ~\new_[27407]_ );
  assign \new_[15225]_  = ~\new_[16414]_ ;
  assign \new_[15226]_  = (~\new_[19590]_  | ~\m2_addr_i[25] ) & (~\new_[18895]_  | ~\m1_addr_i[25] );
  assign \new_[15227]_  = ~\new_[17503]_  & ~\new_[26976]_ ;
  assign \new_[15228]_  = (~\new_[18119]_  | ~\m2_addr_i[24] ) & (~\new_[18892]_  | ~\m1_addr_i[24] );
  assign \new_[15229]_  = ~\new_[22850]_  & (~\new_[17816]_  | ~\new_[26085]_ );
  assign \new_[15230]_  = ~\new_[23117]_  & (~\new_[17817]_  | ~\new_[27241]_ );
  assign \new_[15231]_  = ~\new_[23680]_  & (~\new_[17793]_  | ~\new_[28926]_ );
  assign \new_[15232]_  = (~\m2_addr_i[23]  | ~\new_[18119]_ ) & (~\m1_addr_i[23]  | ~\new_[18896]_ );
  assign \new_[15233]_  = ~\new_[16416]_ ;
  assign \new_[15234]_  = (~\m2_addr_i[22]  | ~\new_[18119]_ ) & (~\m1_addr_i[22]  | ~\new_[18894]_ );
  assign \new_[15235]_  = ~\new_[16417]_ ;
  assign \new_[15236]_  = ~\new_[25115]_  & (~\new_[17794]_  | ~\new_[29210]_ );
  assign \new_[15237]_  = ~\new_[24981]_  & (~\new_[17767]_  | ~\new_[29456]_ );
  assign \new_[15238]_  = \new_[16759]_  | \new_[26279]_ ;
  assign \new_[15239]_  = (~\m2_addr_i[21]  | ~\new_[18119]_ ) & (~\m1_addr_i[21]  | ~\new_[18891]_ );
  assign \new_[15240]_  = ~\new_[21531]_  & (~\new_[17801]_  | ~\new_[23538]_ );
  assign \new_[15241]_  = (~\m2_addr_i[20]  | ~\new_[18119]_ ) & (~\m1_addr_i[20]  | ~\new_[18891]_ );
  assign \new_[15242]_  = (~\m2_addr_i[19]  | ~\new_[18119]_ ) & (~\m1_addr_i[19]  | ~\new_[18893]_ );
  assign \new_[15243]_  = \new_[16760]_  | \new_[25386]_ ;
  assign \new_[15244]_  = ~\new_[17504]_  & ~\new_[26934]_ ;
  assign \new_[15245]_  = (~\m2_addr_i[18]  | ~\new_[18119]_ ) & (~\m1_addr_i[18]  | ~\new_[18893]_ );
  assign \new_[15246]_  = ~\new_[23056]_  & (~\new_[17827]_  | ~\new_[22175]_ );
  assign \new_[15247]_  = ~\new_[23031]_  & (~\new_[17805]_  | ~\new_[25996]_ );
  assign \new_[15248]_  = (~\m2_addr_i[17]  | ~\new_[18119]_ ) & (~\m1_addr_i[17]  | ~\new_[18892]_ );
  assign \new_[15249]_  = ~\new_[27653]_  & (~\new_[17779]_  | ~\new_[24437]_ );
  assign \new_[15250]_  = ~\new_[16421]_ ;
  assign \new_[15251]_  = ~\new_[30199]_  & (~\new_[21914]_  | ~\new_[18265]_ );
  assign \new_[15252]_  = (~\m2_addr_i[16]  | ~\new_[18119]_ ) & (~\m1_addr_i[16]  | ~\new_[18896]_ );
  assign \new_[15253]_  = ~\new_[22851]_  & (~\new_[17834]_  | ~\new_[26400]_ );
  assign \new_[15254]_  = (~\m2_addr_i[15]  | ~\new_[18119]_ ) & (~\m1_addr_i[15]  | ~\new_[18892]_ );
  assign \new_[15255]_  = ~\new_[22848]_  & (~\new_[17835]_  | ~\new_[27550]_ );
  assign \new_[15256]_  = ~\new_[23866]_  & (~\new_[17837]_  | ~\new_[28371]_ );
  assign \new_[15257]_  = ~\new_[16423]_ ;
  assign \new_[15258]_  = ~\new_[16424]_ ;
  assign \new_[15259]_  = (~\m4_data_i[9]  | ~\new_[19612]_ ) & (~\m3_data_i[9]  | ~\new_[18860]_ );
  assign \new_[15260]_  = (~\m2_addr_i[13]  | ~\new_[18119]_ ) & (~\m1_addr_i[13]  | ~\new_[18896]_ );
  assign \new_[15261]_  = ~\new_[17514]_  | ~\new_[20458]_ ;
  assign \new_[15262]_  = (~\m2_addr_i[12]  | ~\new_[18119]_ ) & (~\m1_addr_i[12]  | ~\new_[18896]_ );
  assign \new_[15263]_  = ~\new_[17515]_  | ~\new_[22229]_ ;
  assign \new_[15264]_  = ~\new_[17510]_  & (~\new_[30230]_  | ~\new_[6034]_ );
  assign \new_[15265]_  = ~\new_[24465]_  | ~\new_[27463]_  | ~\new_[17657]_ ;
  assign \new_[15266]_  = ~\new_[30303]_  & (~\new_[17658]_  | ~\new_[23063]_ );
  assign \new_[15267]_  = ~\new_[23417]_  | ~\new_[24162]_  | ~\new_[17601]_ ;
  assign \new_[15268]_  = (~\m2_addr_i[10]  | ~\new_[18119]_ ) & (~\m1_addr_i[10]  | ~\new_[18891]_ );
  assign \new_[15269]_  = ~\new_[26650]_  & (~\new_[17660]_  | ~\new_[22729]_ );
  assign \new_[15270]_  = (~\m2_addr_i[9]  | ~\new_[18119]_ ) & (~\m1_addr_i[9]  | ~\new_[18891]_ );
  assign \new_[15271]_  = ~\new_[22967]_  | ~\new_[26322]_  | ~\new_[17668]_ ;
  assign \new_[15272]_  = (~\m2_addr_i[7]  | ~\new_[18119]_ ) & (~\m1_addr_i[7]  | ~\new_[18892]_ );
  assign \new_[15273]_  = ~\new_[24097]_  | ~\new_[24471]_  | ~\new_[17604]_ ;
  assign \new_[15274]_  = (~\m2_addr_i[6]  | ~\new_[18119]_ ) & (~\m1_addr_i[6]  | ~\new_[18892]_ );
  assign \new_[15275]_  = ~\new_[17516]_  | ~\new_[22973]_ ;
  assign \new_[15276]_  = ~\new_[17511]_  & (~\new_[29815]_  | ~\new_[5967]_ );
  assign \new_[15277]_  = ~\new_[23048]_  | ~\new_[26328]_  | ~\new_[17678]_ ;
  assign \new_[15278]_  = ~\new_[22694]_  & (~\new_[17680]_  | ~\new_[29983]_ );
  assign \new_[15279]_  = (~\m2_addr_i[4]  | ~\new_[18119]_ ) & (~\m1_addr_i[4]  | ~\new_[20572]_ );
  assign \new_[15280]_  = ~\new_[26592]_  & (~\new_[17681]_  | ~\new_[28918]_ );
  assign \new_[15281]_  = ~\new_[23090]_  | ~\new_[23413]_  | ~\new_[17609]_ ;
  assign \new_[15282]_  = (~\m2_addr_i[2]  | ~\new_[18119]_ ) & (~\new_[31477]_  | ~\new_[20572]_ );
  assign \new_[15283]_  = ~\new_[28408]_  & (~\new_[17687]_  | ~\new_[21383]_ );
  assign \new_[15284]_  = (~\m2_addr_i[1]  | ~\new_[18119]_ ) & (~\m1_addr_i[1]  | ~\new_[18896]_ );
  assign \new_[15285]_  = ~\new_[26614]_  & (~\new_[17693]_  | ~\new_[28836]_ );
  assign \new_[15286]_  = (~\m2_addr_i[0]  | ~\new_[18119]_ ) & (~\m1_addr_i[0]  | ~\new_[18891]_ );
  assign \new_[15287]_  = ~\new_[24491]_  | ~\new_[24450]_  | ~\new_[17614]_ ;
  assign \new_[15288]_  = (~\m2_sel_i[3]  | ~\new_[19590]_ ) & (~\m1_sel_i[3]  | ~\new_[18892]_ );
  assign \new_[15289]_  = ~\new_[26615]_  & (~\new_[17697]_  | ~\new_[21400]_ );
  assign \new_[15290]_  = ~\new_[23267]_  | ~\new_[27640]_  | ~\new_[17702]_ ;
  assign \new_[15291]_  = (~\m2_sel_i[1]  | ~\new_[18119]_ ) & (~\m1_sel_i[1]  | ~\new_[18892]_ );
  assign \new_[15292]_  = ~\new_[28651]_  & (~\new_[17703]_  | ~\new_[22983]_ );
  assign \new_[15293]_  = ~\new_[21921]_  & (~\new_[17704]_  | ~\new_[29186]_ );
  assign \new_[15294]_  = (~\m2_sel_i[0]  | ~\new_[18119]_ ) & (~\m1_sel_i[0]  | ~\new_[18896]_ );
  assign \new_[15295]_  = (~m2_we_i | ~\new_[18119]_ ) & (~m1_we_i | ~\new_[20572]_ );
  assign \new_[15296]_  = ~\new_[29206]_  & (~\new_[17711]_  | ~\new_[30242]_ );
  assign \new_[15297]_  = ~\new_[26693]_  | ~\new_[26271]_  | ~\new_[17619]_ ;
  assign \new_[15298]_  = ~\new_[17517]_  | ~\new_[24425]_ ;
  assign \new_[15299]_  = (~\m4_data_i[31]  | ~\new_[18159]_ ) & (~\m3_data_i[31]  | ~\new_[18197]_ );
  assign \new_[15300]_  = (~\m4_data_i[30]  | ~\new_[19615]_ ) & (~\m3_data_i[30]  | ~\new_[18198]_ );
  assign \new_[15301]_  = (~\m4_data_i[29]  | ~\new_[19615]_ ) & (~\m3_data_i[29]  | ~\new_[18198]_ );
  assign \new_[15302]_  = ~\new_[17519]_  | ~\new_[22865]_ ;
  assign \new_[15303]_  = (~\m4_data_i[11]  | ~\new_[19612]_ ) & (~\m3_data_i[11]  | ~\new_[20568]_ );
  assign \new_[15304]_  = ~\new_[24410]_  | ~\new_[27525]_  | ~\new_[17745]_ ;
  assign \new_[15305]_  = ~\new_[22618]_  & (~\new_[17746]_  | ~\new_[28684]_ );
  assign \new_[15306]_  = ~\new_[24378]_  | ~\new_[23155]_  | ~\new_[17624]_ ;
  assign \new_[15307]_  = (~\m4_data_i[27]  | ~\new_[18159]_ ) & (~\m3_data_i[27]  | ~\new_[18196]_ );
  assign \new_[15308]_  = (~\m4_data_i[26]  | ~\new_[18160]_ ) & (~\m3_data_i[26]  | ~\new_[18199]_ );
  assign \new_[15309]_  = ~\new_[28942]_  & (~\new_[17752]_  | ~\new_[30198]_ );
  assign \new_[15310]_  = ~\new_[28353]_  | ~\new_[26220]_  | ~\new_[17626]_ ;
  assign \new_[15311]_  = (~\m4_data_i[25]  | ~\new_[18162]_ ) & (~\m3_data_i[25]  | ~\new_[19636]_ );
  assign \new_[15312]_  = (~\m4_data_i[24]  | ~\new_[19615]_ ) & (~\m3_data_i[24]  | ~\new_[18198]_ );
  assign \new_[15313]_  = ~\new_[22210]_  & (~\new_[17743]_  | ~\new_[28121]_ );
  assign \new_[15314]_  = ~\new_[26751]_  & (~\new_[17740]_  | ~\new_[29276]_ );
  assign \new_[15315]_  = ~\new_[23621]_  | ~\new_[23078]_  | ~\new_[17629]_ ;
  assign \new_[15316]_  = (~\m4_data_i[23]  | ~\new_[19615]_ ) & (~\m3_data_i[23]  | ~\new_[18198]_ );
  assign \new_[15317]_  = (~\m4_data_i[22]  | ~\new_[18159]_ ) & (~\m3_data_i[22]  | ~\new_[19636]_ );
  assign \new_[15318]_  = ~\new_[21465]_  | ~\new_[27418]_  | ~\new_[17810]_ ;
  assign \new_[15319]_  = (~\m4_data_i[20]  | ~\new_[18159]_ ) & (~\m3_data_i[20]  | ~\new_[18197]_ );
  assign \new_[15320]_  = ~\new_[22942]_  & (~\new_[17808]_  | ~\new_[28245]_ );
  assign \new_[15321]_  = ~\new_[27410]_  & (~\new_[17770]_  | ~\new_[29410]_ );
  assign \new_[15322]_  = ~\new_[24065]_  | ~\new_[24081]_  | ~\new_[17633]_ ;
  assign \new_[15323]_  = (~\m4_data_i[19]  | ~\new_[18159]_ ) & (~\m3_data_i[19]  | ~\new_[18198]_ );
  assign \new_[15324]_  = (~\m4_data_i[17]  | ~\new_[19615]_ ) & (~\m3_data_i[17]  | ~\new_[18198]_ );
  assign \new_[15325]_  = ~\new_[17520]_  | ~\new_[22990]_ ;
  assign \new_[15326]_  = ~\new_[23134]_  | ~\new_[24745]_  | ~\new_[17774]_ ;
  assign \new_[15327]_  = ~\new_[26438]_  & (~\new_[17775]_  | ~\new_[28595]_ );
  assign \new_[15328]_  = (~\m4_data_i[16]  | ~\new_[18159]_ ) & (~\m3_data_i[16]  | ~\new_[19636]_ );
  assign \new_[15329]_  = (~\m4_data_i[15]  | ~\new_[19615]_ ) & (~\m3_data_i[15]  | ~\new_[18198]_ );
  assign \new_[15330]_  = ~\new_[29319]_  & (~\new_[17723]_  | ~\new_[30693]_ );
  assign \new_[15331]_  = ~\new_[28895]_  & (~\new_[17778]_  | ~\new_[22699]_ );
  assign \new_[15332]_  = (~\m4_data_i[14]  | ~\new_[18164]_ ) & (~\m3_data_i[14]  | ~\new_[18198]_ );
  assign \new_[15333]_  = (~\m4_data_i[13]  | ~\new_[19615]_ ) & (~\m3_data_i[13]  | ~\new_[18199]_ );
  assign \new_[15334]_  = ~\new_[21798]_  | ~\new_[26226]_  | ~\new_[17780]_ ;
  assign \new_[15335]_  = (~\m4_data_i[12]  | ~\new_[19615]_ ) & (~\m3_data_i[12]  | ~\new_[18198]_ );
  assign \new_[15336]_  = ~\new_[22887]_  | ~\new_[22891]_  | ~\new_[17638]_ ;
  assign \new_[15337]_  = (~\m4_data_i[11]  | ~\new_[18160]_ ) & (~\m3_data_i[11]  | ~\new_[18199]_ );
  assign \new_[15338]_  = ~\new_[24746]_  & (~\new_[17784]_  | ~\new_[27802]_ );
  assign \new_[15339]_  = ~\new_[26285]_  | ~\new_[26701]_  | ~\new_[17610]_ ;
  assign \new_[15340]_  = ~\new_[27870]_  & (~\new_[17663]_  | ~\new_[21364]_ );
  assign \new_[15341]_  = (~\m4_data_i[10]  | ~\new_[19615]_ ) & (~\m3_data_i[10]  | ~\new_[18199]_ );
  assign \new_[15342]_  = (~\m4_data_i[9]  | ~\new_[19615]_ ) & (~\m3_data_i[9]  | ~\new_[18198]_ );
  assign \new_[15343]_  = ~\new_[22880]_  | ~\new_[23046]_  | ~\new_[17790]_ ;
  assign \new_[15344]_  = (~\m2_data_i[0]  | ~\new_[19572]_ ) & (~\m1_data_i[0]  | ~\new_[18187]_ );
  assign \new_[15345]_  = ~\new_[23001]_  & (~\new_[17674]_  | ~\new_[28732]_ );
  assign \new_[15346]_  = (~\m4_data_i[8]  | ~\new_[19615]_ ) & (~\m3_data_i[8]  | ~\new_[18198]_ );
  assign \new_[15347]_  = ~\new_[26661]_  & (~\new_[17677]_  | ~\new_[29623]_ );
  assign \new_[15348]_  = ~\new_[23152]_  | ~\new_[24213]_  | ~\new_[17644]_ ;
  assign \new_[15349]_  = (~\m4_data_i[7]  | ~\new_[18164]_ ) & (~\m3_data_i[7]  | ~\new_[18198]_ );
  assign \new_[15350]_  = (~\m4_data_i[6]  | ~\new_[18164]_ ) & (~\m3_data_i[6]  | ~\new_[18198]_ );
  assign \new_[15351]_  = (~\m4_data_i[5]  | ~\new_[18165]_ ) & (~\m3_data_i[5]  | ~\new_[18198]_ );
  assign \new_[15352]_  = ~\new_[17521]_  | ~\new_[19446]_ ;
  assign \new_[15353]_  = ~\new_[17522]_  | ~\new_[22587]_ ;
  assign \new_[15354]_  = (~\m4_data_i[4]  | ~\new_[19615]_ ) & (~\m3_data_i[4]  | ~\new_[18199]_ );
  assign \new_[15355]_  = ~\new_[17523]_  | ~\new_[22846]_ ;
  assign \new_[15356]_  = ~\new_[17512]_  & (~\new_[30115]_  | ~\new_[6270]_ );
  assign \new_[15357]_  = (~\m4_data_i[3]  | ~\new_[18161]_ ) & (~\m3_data_i[3]  | ~\new_[18199]_ );
  assign \new_[15358]_  = ~\new_[24462]_  | ~\new_[24792]_  | ~\new_[17771]_ ;
  assign \new_[15359]_  = (~\m2_data_i[2]  | ~\new_[18074]_ ) & (~\m1_data_i[2]  | ~\new_[19629]_ );
  assign \new_[15360]_  = ~\new_[22850]_  & (~\new_[17792]_  | ~\new_[28640]_ );
  assign \new_[15361]_  = (~\m4_data_i[2]  | ~\new_[18160]_ ) & (~\m3_data_i[2]  | ~\new_[18199]_ );
  assign \new_[15362]_  = ~\new_[24445]_  | ~\new_[24290]_  | ~\new_[17622]_ ;
  assign \new_[15363]_  = (~\m4_data_i[31]  | ~\new_[19609]_ ) & (~\m3_data_i[31]  | ~\new_[18201]_ );
  assign \new_[15364]_  = (~\m4_data_i[1]  | ~\new_[18164]_ ) & (~\m3_data_i[1]  | ~\new_[18198]_ );
  assign \new_[15365]_  = ~\new_[28065]_  | ~\new_[27907]_  | ~\new_[17648]_ ;
  assign \new_[15366]_  = ~\new_[27015]_  & (~\new_[17815]_  | ~\new_[24247]_ );
  assign \new_[15367]_  = (~\m4_data_i[30]  | ~\new_[19609]_ ) & (~\m3_data_i[30]  | ~\new_[18201]_ );
  assign \new_[15368]_  = (~\new_[19615]_  | ~\m4_addr_i[31] ) & (~\new_[18198]_  | ~\m3_addr_i[31] );
  assign \new_[15369]_  = ~\new_[21585]_  | ~\new_[27705]_  | ~\new_[17799]_ ;
  assign \new_[15370]_  = (~\m7_data_i[30]  | ~\new_[18823]_ ) & (~\m0_data_i[30]  | ~\new_[18731]_ );
  assign \new_[15371]_  = ~\new_[21884]_  | ~\new_[22926]_  | ~\new_[17642]_ ;
  assign \new_[15372]_  = (~\new_[18159]_  | ~\m4_addr_i[30] ) & (~\new_[18197]_  | ~\m3_addr_i[30] );
  assign \new_[15373]_  = ~\new_[24345]_  & (~\new_[17659]_  | ~\new_[28535]_ );
  assign \new_[15374]_  = (~\m4_data_i[29]  | ~\new_[19609]_ ) & (~\m3_data_i[29]  | ~\new_[18201]_ );
  assign \new_[15375]_  = ~\new_[24444]_  | ~\new_[26572]_  | ~\new_[17643]_ ;
  assign \new_[15376]_  = (~\m7_data_i[29]  | ~\new_[18823]_ ) & (~\m0_data_i[29]  | ~\new_[19537]_ );
  assign \new_[15377]_  = ~\new_[17524]_  | ~\new_[21994]_ ;
  assign \new_[15378]_  = (~\new_[18161]_  | ~\m4_addr_i[28] ) & (~\new_[18196]_  | ~\m3_addr_i[28] );
  assign \new_[15379]_  = ~\new_[17518]_  | ~\new_[24446]_ ;
  assign \new_[15380]_  = ~\new_[17513]_  & (~\new_[30157]_  | ~\new_[6215]_ );
  assign \new_[15381]_  = (~\m4_data_i[28]  | ~\new_[19609]_ ) & (~\m3_data_i[28]  | ~\new_[18201]_ );
  assign \new_[15382]_  = ~\new_[24399]_  | ~\new_[26355]_  | ~\new_[17789]_ ;
  assign \new_[15383]_  = (~\m2_data_i[18]  | ~\new_[18119]_ ) & (~\m1_data_i[18]  | ~\new_[18891]_ );
  assign \new_[15384]_  = (~\new_[18159]_  | ~\m4_addr_i[27] ) & (~\new_[18196]_  | ~\m3_addr_i[27] );
  assign \new_[15385]_  = (~\new_[18161]_  | ~\m4_addr_i[26] ) & (~\new_[18196]_  | ~\m3_addr_i[26] );
  assign \new_[15386]_  = ~\new_[28419]_  | ~\new_[28133]_  | ~\new_[17645]_ ;
  assign \new_[15387]_  = (~\m2_data_i[27]  | ~\new_[18799]_ ) & (~\m1_data_i[27]  | ~\new_[18887]_ );
  assign \new_[15388]_  = ~\new_[21531]_  & (~\new_[17824]_  | ~\new_[28280]_ );
  assign \new_[15389]_  = (~\m7_data_i[27]  | ~\new_[18823]_ ) & (~\m0_data_i[27]  | ~\new_[18731]_ );
  assign \new_[15390]_  = (~\new_[18161]_  | ~\m4_addr_i[25] ) & (~\new_[18196]_  | ~\m3_addr_i[25] );
  assign \new_[15391]_  = (~\m4_data_i[27]  | ~\new_[19609]_ ) & (~\m3_data_i[27]  | ~\new_[19639]_ );
  assign \new_[15392]_  = ~\new_[24275]_  | ~\new_[26632]_  | ~\new_[17831]_ ;
  assign \new_[15393]_  = ~\new_[28677]_  & (~\new_[17832]_  | ~\new_[23065]_ );
  assign \new_[15394]_  = (~\new_[18159]_  | ~\m4_addr_i[24] ) & (~\new_[19636]_  | ~\m3_addr_i[24] );
  assign \new_[15395]_  = (~\m4_addr_i[23]  | ~\new_[18159]_ ) & (~\m3_addr_i[23]  | ~\new_[19636]_ );
  assign \new_[15396]_  = ~\new_[28289]_  | ~\new_[27606]_  | ~\new_[17653]_ ;
  assign \new_[15397]_  = (~\m4_addr_i[22]  | ~\new_[18159]_ ) & (~\m3_addr_i[22]  | ~\new_[18196]_ );
  assign \new_[15398]_  = ~\new_[26763]_  & (~\new_[17838]_  | ~\new_[21435]_ );
  assign \new_[15399]_  = (~\m4_addr_i[21]  | ~\new_[18159]_ ) & (~\m3_addr_i[21]  | ~\new_[18197]_ );
  assign \new_[15400]_  = (~\m2_data_i[25]  | ~\new_[18799]_ ) & (~\m1_data_i[25]  | ~\new_[18887]_ );
  assign \new_[15401]_  = (~\m4_data_i[25]  | ~\new_[18143]_ ) & (~\m3_data_i[25]  | ~\new_[18201]_ );
  assign \new_[15402]_  = (~\m4_addr_i[20]  | ~\new_[18159]_ ) & (~\m3_addr_i[20]  | ~\new_[18199]_ );
  assign \new_[15403]_  = (~\m4_data_i[24]  | ~\new_[18143]_ ) & (~\m3_data_i[24]  | ~\new_[18201]_ );
  assign \new_[15404]_  = (~\m4_addr_i[19]  | ~\new_[18159]_ ) & (~\m3_addr_i[19]  | ~\new_[18199]_ );
  assign \new_[15405]_  = (~\m4_addr_i[18]  | ~\new_[19615]_ ) & (~\m3_addr_i[18]  | ~\new_[18198]_ );
  assign \new_[15406]_  = (~\m4_data_i[23]  | ~\new_[19609]_ ) & (~\m3_data_i[23]  | ~\new_[18201]_ );
  assign \new_[15407]_  = ~\new_[26379]_  & (~\new_[17939]_  | ~\new_[29900]_ );
  assign \new_[15408]_  = (~\m4_addr_i[17]  | ~\new_[18163]_ ) & (~\m3_addr_i[17]  | ~\new_[19636]_ );
  assign \new_[15409]_  = ~\new_[17435]_  & ~\new_[28687]_ ;
  assign \new_[15410]_  = ~\new_[26668]_  & (~\new_[17940]_  | ~\new_[30097]_ );
  assign \new_[15411]_  = ~\new_[23022]_  | (~\new_[17666]_  & ~\new_[28397]_ );
  assign \new_[15412]_  = (~\m4_addr_i[16]  | ~\new_[19615]_ ) & (~\m3_addr_i[16]  | ~\new_[18198]_ );
  assign \new_[15413]_  = (~\m2_data_i[22]  | ~\new_[18799]_ ) & (~\m1_data_i[22]  | ~\new_[18887]_ );
  assign \new_[15414]_  = (~\m4_data_i[22]  | ~\new_[18145]_ ) & (~\m3_data_i[22]  | ~\new_[18201]_ );
  assign \new_[15415]_  = (~\m4_addr_i[15]  | ~\new_[18165]_ ) & (~\m3_addr_i[15]  | ~\new_[19636]_ );
  assign \new_[15416]_  = ~\new_[27626]_  & (~\new_[17943]_  | ~\new_[30172]_ );
  assign \new_[15417]_  = (~\m4_addr_i[14]  | ~\new_[19615]_ ) & (~\m3_addr_i[14]  | ~\new_[19636]_ );
  assign \new_[15418]_  = ~\new_[26352]_  & (~\new_[17944]_  | ~\new_[29251]_ );
  assign \new_[15419]_  = (~\m2_data_i[21]  | ~\new_[18799]_ ) & (~\m1_data_i[21]  | ~\new_[18887]_ );
  assign \new_[15420]_  = (~\m4_data_i[21]  | ~\new_[18143]_ ) & (~\m3_data_i[21]  | ~\new_[18201]_ );
  assign \new_[15421]_  = (~\m4_addr_i[13]  | ~\new_[18162]_ ) & (~\m3_addr_i[13]  | ~\new_[19636]_ );
  assign \new_[15422]_  = ~\new_[17454]_  & ~\new_[28566]_ ;
  assign \new_[15423]_  = ~\new_[25892]_  & (~\new_[17945]_  | ~\new_[29984]_ );
  assign \new_[15424]_  = ~\new_[24425]_  | (~\new_[17730]_  & ~\new_[28944]_ );
  assign \new_[15425]_  = (~\m4_data_i[31]  | ~\new_[19613]_ ) & (~\m3_data_i[31]  | ~\new_[20568]_ );
  assign \new_[15426]_  = ~\new_[27979]_  & (~\new_[17947]_  | ~\new_[30697]_ );
  assign \new_[15427]_  = ~\new_[17460]_  & ~\new_[26999]_ ;
  assign \new_[15428]_  = (~\m4_data_i[20]  | ~\new_[18146]_ ) & (~\m3_data_i[20]  | ~\new_[18201]_ );
  assign \new_[15429]_  = ~\new_[17464]_  & ~\new_[28341]_ ;
  assign \new_[15430]_  = ~\new_[17472]_  & ~\new_[28978]_ ;
  assign \new_[15431]_  = (~\m4_addr_i[10]  | ~\new_[18162]_ ) & (~\m3_addr_i[10]  | ~\new_[19636]_ );
  assign \new_[15432]_  = (~\m2_data_i[19]  | ~\new_[18799]_ ) & (~\m1_data_i[19]  | ~\new_[18887]_ );
  assign \new_[15433]_  = (~\m4_addr_i[11]  | ~\new_[18160]_ ) & (~\m3_addr_i[11]  | ~\new_[18199]_ );
  assign \new_[15434]_  = (~\m4_addr_i[9]  | ~\new_[18159]_ ) & (~\m3_addr_i[9]  | ~\new_[18198]_ );
  assign \new_[15435]_  = (~\m4_data_i[19]  | ~\new_[18147]_ ) & (~\m3_data_i[19]  | ~\new_[18201]_ );
  assign \new_[15436]_  = (~\m4_addr_i[8]  | ~\new_[18160]_ ) & (~\m3_addr_i[8]  | ~\new_[18199]_ );
  assign \new_[15437]_  = ~\new_[22990]_  | (~\new_[17802]_  & ~\new_[30348]_ );
  assign \new_[15438]_  = ~\new_[17481]_  & ~\new_[27994]_ ;
  assign \new_[15439]_  = (~\m4_addr_i[7]  | ~\new_[19615]_ ) & (~\m3_addr_i[7]  | ~\new_[18198]_ );
  assign \new_[15440]_  = (~\m4_data_i[18]  | ~\new_[18143]_ ) & (~\m3_data_i[18]  | ~\new_[19639]_ );
  assign \new_[15441]_  = ~\new_[26276]_  & (~\new_[17946]_  | ~\new_[29299]_ );
  assign \new_[15442]_  = (~\m4_addr_i[6]  | ~\new_[18163]_ ) & (~\m3_addr_i[6]  | ~\new_[18198]_ );
  assign \new_[15443]_  = ~\new_[17419]_  & ~\new_[17317]_ ;
  assign \new_[15444]_  = (~\m2_data_i[17]  | ~\new_[18799]_ ) & (~\m1_data_i[17]  | ~\new_[18887]_ );
  assign \new_[15445]_  = ~\new_[22846]_  | (~\new_[17819]_  & ~\new_[30620]_ );
  assign \new_[15446]_  = (~\m4_addr_i[5]  | ~\new_[18164]_ ) & (~\m3_addr_i[5]  | ~\new_[18198]_ );
  assign \new_[15447]_  = (~\m4_data_i[17]  | ~\new_[18142]_ ) & (~\m3_data_i[17]  | ~\new_[19639]_ );
  assign \new_[15448]_  = ~\new_[17493]_  & ~\new_[29632]_ ;
  assign \new_[15449]_  = (~\m4_addr_i[4]  | ~\new_[18165]_ ) & (~\m3_addr_i[4]  | ~\new_[18198]_ );
  assign \new_[15450]_  = ~\new_[27667]_  & (~\new_[17941]_  | ~\new_[30159]_ );
  assign \new_[15451]_  = ~\new_[22642]_  | (~\new_[17655]_  & ~\new_[29508]_ );
  assign \new_[15452]_  = ~\new_[24414]_  & (~\new_[17942]_  | ~\new_[28001]_ );
  assign \new_[15453]_  = (~\m4_data_i[16]  | ~\new_[19609]_ ) & (~\m3_data_i[16]  | ~\new_[18201]_ );
  assign \new_[15454]_  = ~\new_[24446]_  | (~\new_[17685]_  & ~\new_[30755]_ );
  assign \new_[15455]_  = ~\new_[17500]_  & ~\new_[29468]_ ;
  assign \new_[15456]_  = (~\m4_addr_i[1]  | ~\new_[18162]_ ) & (~\m3_addr_i[1]  | ~\new_[18198]_ );
  assign \new_[15457]_  = (~\m4_data_i[15]  | ~\new_[18144]_ ) & (~\m3_data_i[15]  | ~\new_[18201]_ );
  assign \new_[15458]_  = ~\new_[17507]_  & ~\new_[28454]_ ;
  assign \new_[15459]_  = (~\m4_data_i[14]  | ~\new_[18143]_ ) & (~\m3_data_i[14]  | ~\new_[18201]_ );
  assign \new_[15460]_  = (~\m4_sel_i[2]  | ~\new_[18163]_ ) & (~\m3_sel_i[2]  | ~\new_[19636]_ );
  assign \new_[15461]_  = (~\m2_data_i[13]  | ~\new_[18799]_ ) & (~\m1_data_i[13]  | ~\new_[18887]_ );
  assign \new_[15462]_  = (~\m4_data_i[13]  | ~\new_[19609]_ ) & (~\m3_data_i[13]  | ~\new_[18201]_ );
  assign \new_[15463]_  = (~\m4_sel_i[0]  | ~\new_[18165]_ ) & (~\m3_sel_i[0]  | ~\new_[18198]_ );
  assign \new_[15464]_  = (~\m2_data_i[12]  | ~\new_[18799]_ ) & (~\m1_data_i[12]  | ~\new_[18887]_ );
  assign \new_[15465]_  = (~\m4_data_i[12]  | ~\new_[18143]_ ) & (~\m3_data_i[12]  | ~\new_[18201]_ );
  assign \new_[15466]_  = (~m4_we_i | ~\new_[18165]_ ) & (~m3_we_i | ~\new_[18198]_ );
  assign \new_[15467]_  = ~\new_[29453]_  & (~\new_[17821]_  | ~\new_[30363]_ );
  assign \new_[15468]_  = (~\m4_data_i[11]  | ~\new_[18144]_ ) & (~\m3_data_i[11]  | ~\new_[19639]_ );
  assign \new_[15469]_  = (~\m4_data_i[10]  | ~\new_[18143]_ ) & (~\m3_data_i[10]  | ~\new_[18201]_ );
  assign \new_[15470]_  = (~\m4_data_i[9]  | ~\new_[19609]_ ) & (~\m3_data_i[9]  | ~\new_[18201]_ );
  assign \new_[15471]_  = ~\new_[30259]_  & (~\new_[17840]_  | ~\new_[29357]_ );
  assign \new_[15472]_  = (~\m2_data_i[8]  | ~\new_[18799]_ ) & (~\m1_data_i[8]  | ~\new_[18887]_ );
  assign \new_[15473]_  = (~\m4_data_i[8]  | ~\new_[18144]_ ) & (~\m3_data_i[8]  | ~\new_[19639]_ );
  assign \new_[15474]_  = ~\new_[16725]_  & (~\new_[29930]_  | ~\new_[6096]_ );
  assign \new_[15475]_  = ~\new_[16726]_  & (~\new_[30174]_  | ~\new_[6096]_ );
  assign \new_[15476]_  = ~\new_[16721]_  & (~\new_[30564]_  | ~\new_[31712]_ );
  assign \new_[15477]_  = (~\m4_data_i[7]  | ~\new_[18144]_ ) & (~\m3_data_i[7]  | ~\new_[19639]_ );
  assign \new_[15478]_  = ~\new_[17420]_  & (~\new_[30185]_  | ~\new_[31440]_ );
  assign \new_[15479]_  = (~\m2_data_i[6]  | ~\new_[18799]_ ) & (~\m1_data_i[6]  | ~\new_[18887]_ );
  assign \new_[15480]_  = (~\m4_data_i[6]  | ~\new_[18144]_ ) & (~\m3_data_i[6]  | ~\new_[19639]_ );
  assign \new_[15481]_  = ~\new_[17383]_  & (~\new_[30651]_  | ~\new_[30897]_ );
  assign \new_[15482]_  = (~\m2_data_i[5]  | ~\new_[18799]_ ) & (~\m1_data_i[5]  | ~\new_[18887]_ );
  assign \new_[15483]_  = (~\m4_data_i[5]  | ~\new_[18143]_ ) & (~\m3_data_i[5]  | ~\new_[18201]_ );
  assign \new_[15484]_  = ~\new_[16732]_  & (~\new_[29916]_  | ~\new_[6072]_ );
  assign \new_[15485]_  = (~\m4_data_i[4]  | ~\new_[19609]_ ) & (~\m3_data_i[4]  | ~\new_[18201]_ );
  assign \new_[15486]_  = (~\m4_data_i[3]  | ~\new_[19609]_ ) & (~\m3_data_i[3]  | ~\new_[18201]_ );
  assign \new_[15487]_  = (~\m2_data_i[3]  | ~\new_[18799]_ ) & (~\m1_data_i[3]  | ~\new_[18887]_ );
  assign \new_[15488]_  = ~\new_[16735]_  & (~\new_[30225]_  | ~\new_[6184]_ );
  assign \new_[15489]_  = (~\m2_data_i[2]  | ~\new_[18799]_ ) & (~\m1_data_i[2]  | ~\new_[18887]_ );
  assign \new_[15490]_  = ~\new_[16737]_  & (~\new_[30708]_  | ~\new_[6216]_ );
  assign \new_[15491]_  = (~\m4_data_i[2]  | ~\new_[18144]_ ) & (~\m3_data_i[2]  | ~\new_[19639]_ );
  assign \new_[15492]_  = ~\new_[17438]_  & (~\new_[29855]_  | ~\new_[5909]_ );
  assign \new_[15493]_  = (~\new_[17667]_  | ~\new_[30337]_ ) & (~\new_[30663]_  | ~\new_[6040]_ );
  assign \new_[15494]_  = ~\new_[17442]_  & (~\new_[29100]_  | ~\new_[5911]_ );
  assign \new_[15495]_  = (~\m4_data_i[1]  | ~\new_[18144]_ ) & (~\m3_data_i[1]  | ~\new_[18201]_ );
  assign \new_[15496]_  = ~\new_[17446]_  & (~\new_[30389]_  | ~\new_[5912]_ );
  assign \new_[15497]_  = (~\m4_data_i[0]  | ~\new_[18143]_ ) & (~\m3_data_i[0]  | ~\new_[18201]_ );
  assign \new_[15498]_  = ~\new_[17451]_  & (~\new_[28899]_  | ~\new_[5914]_ );
  assign \new_[15499]_  = (~\m2_data_i[0]  | ~\new_[18799]_ ) & (~\m1_data_i[0]  | ~\new_[18887]_ );
  assign \new_[15500]_  = (~\new_[17700]_  | ~\new_[30160]_ ) & (~\new_[30711]_  | ~\new_[31712]_ );
  assign \new_[15501]_  = (~\m7_data_i[0]  | ~\new_[18823]_ ) & (~\m0_data_i[0]  | ~\new_[18731]_ );
  assign \new_[15502]_  = (~\new_[17679]_  | ~\new_[30146]_ ) & (~\new_[30443]_  | ~\new_[31440]_ );
  assign \new_[15503]_  = (~\new_[17731]_  | ~\new_[30728]_ ) & (~\new_[28846]_  | ~\new_[31440]_ );
  assign \new_[15504]_  = (~\new_[19609]_  | ~\m4_addr_i[31] ) & (~\new_[18201]_  | ~\m3_addr_i[31] );
  assign \new_[15505]_  = (~\new_[17742]_  | ~\new_[30349]_ ) & (~\new_[30675]_  | ~\new_[30884]_ );
  assign \new_[15506]_  = (~\new_[18799]_  | ~\new_[31486]_ ) & (~\new_[18887]_  | ~\new_[31308]_ );
  assign \new_[15507]_  = ~\new_[17475]_  & (~\new_[29573]_  | ~\new_[5917]_ );
  assign \new_[15508]_  = (~\new_[18143]_  | ~\m4_addr_i[30] ) & (~\new_[19639]_  | ~\m3_addr_i[30] );
  assign \new_[15509]_  = ~\new_[17479]_  & (~\new_[29767]_  | ~\new_[5918]_ );
  assign \new_[15510]_  = (~\new_[17725]_  | ~\new_[30071]_ ) & (~\new_[30780]_  | ~\new_[6069]_ );
  assign \new_[15511]_  = (~\new_[17773]_  | ~\new_[29802]_ ) & (~\new_[30684]_  | ~\new_[6069]_ );
  assign \new_[15512]_  = (~\new_[18799]_  | ~\m2_addr_i[29] ) & (~\new_[18887]_  | ~\new_[31538]_ );
  assign \new_[15513]_  = ~\new_[17483]_  & (~\new_[29648]_  | ~\new_[5921]_ );
  assign \new_[15514]_  = (~\new_[19609]_  | ~\m4_addr_i[29] ) & (~\new_[18201]_  | ~\m3_addr_i[29] );
  assign \new_[15515]_  = (~\new_[18823]_  | ~\new_[31531]_ ) & (~\new_[20539]_  | ~\new_[31481]_ );
  assign \new_[15516]_  = ~\new_[17488]_  & (~\new_[29565]_  | ~\new_[5923]_ );
  assign \new_[15517]_  = (~\m2_data_i[9]  | ~\new_[19572]_ ) & (~\m1_data_i[9]  | ~\new_[18191]_ );
  assign \new_[15518]_  = (~\new_[19609]_  | ~\m4_addr_i[28] ) & (~\new_[18201]_  | ~\m3_addr_i[28] );
  assign \new_[15519]_  = (~\new_[17818]_  | ~\new_[29813]_ ) & (~\new_[30682]_  | ~\new_[6078]_ );
  assign \new_[15520]_  = ~\new_[17495]_  & (~\new_[29898]_  | ~\new_[5927]_ );
  assign \new_[15521]_  = (~\new_[17796]_  | ~\new_[30142]_ ) & (~\new_[30840]_  | ~\new_[6084]_ );
  assign \new_[15522]_  = (~\new_[17803]_  | ~\new_[30218]_ ) & (~\new_[30713]_  | ~\new_[30998]_ );
  assign \new_[15523]_  = (~\new_[19609]_  | ~\m4_addr_i[27] ) & (~\new_[18201]_  | ~\m3_addr_i[27] );
  assign \new_[15524]_  = (~\new_[17714]_  | ~\new_[30352]_ ) & (~\new_[30557]_  | ~\new_[30998]_ );
  assign \new_[15525]_  = (~\new_[17820]_  | ~\new_[30278]_ ) & (~\new_[30501]_  | ~\new_[6078]_ );
  assign \new_[15526]_  = (~\new_[17829]_  | ~\new_[29897]_ ) & (~\new_[30545]_  | ~\new_[31045]_ );
  assign \new_[15527]_  = ~\new_[17509]_  & (~\new_[29119]_  | ~\new_[6094]_ );
  assign \new_[15528]_  = (~\new_[18143]_  | ~\m4_addr_i[26] ) & (~\new_[19639]_  | ~\m3_addr_i[26] );
  assign \new_[15529]_  = ~\new_[27518]_  & (~\new_[17952]_  | ~\new_[29969]_ );
  assign \new_[15530]_  = ~\new_[24566]_  & (~\new_[17953]_  | ~\new_[29435]_ );
  assign \new_[15531]_  = ~\new_[27773]_  & (~\new_[17954]_  | ~\new_[29983]_ );
  assign \new_[15532]_  = (~\new_[19609]_  | ~\m4_addr_i[25] ) & (~\new_[18201]_  | ~\m3_addr_i[25] );
  assign \new_[15533]_  = ~\new_[27571]_  & (~\new_[17955]_  | ~\new_[28050]_ );
  assign \new_[15534]_  = ~\new_[24752]_  & (~\new_[17956]_  | ~\new_[29186]_ );
  assign \new_[15535]_  = (~\new_[19609]_  | ~\m4_addr_i[24] ) & (~\new_[18201]_  | ~\m3_addr_i[24] );
  assign \new_[15536]_  = ~\new_[26815]_  & (~\new_[17951]_  | ~\new_[30022]_ );
  assign \new_[15537]_  = ~\new_[27325]_  & (~\new_[17958]_  | ~\new_[29593]_ );
  assign \new_[15538]_  = (~\m4_addr_i[23]  | ~\new_[19609]_ ) & (~\m3_addr_i[23]  | ~\new_[19639]_ );
  assign \new_[15539]_  = ~\new_[28369]_  & (~\new_[17966]_  | ~\new_[30552]_ );
  assign \new_[15540]_  = ~\new_[26686]_  & (~\new_[17959]_  | ~\new_[28806]_ );
  assign \new_[15541]_  = ~\new_[28274]_  & (~\new_[17960]_  | ~\new_[28684]_ );
  assign \new_[15542]_  = (~\m4_data_i[25]  | ~\new_[19614]_ ) & (~\m3_data_i[25]  | ~\new_[20568]_ );
  assign \new_[15543]_  = ~\new_[28217]_  & (~\new_[17961]_  | ~\new_[30628]_ );
  assign \new_[15544]_  = ~\new_[28287]_  & (~\new_[17962]_  | ~\new_[30627]_ );
  assign \new_[15545]_  = ~\new_[26604]_  & (~\new_[17957]_  | ~\new_[28121]_ );
  assign \new_[15546]_  = (~\m7_addr_i[23]  | ~\new_[18823]_ ) & (~\m0_addr_i[23]  | ~\new_[19537]_ );
  assign \new_[15547]_  = ~\new_[28548]_  & (~\new_[17963]_  | ~\new_[28039]_ );
  assign \new_[15548]_  = ~\new_[27624]_  & (~\new_[17967]_  | ~\new_[28245]_ );
  assign \new_[15549]_  = (~\m4_addr_i[22]  | ~\new_[19609]_ ) & (~\m3_addr_i[22]  | ~\new_[18201]_ );
  assign \new_[15550]_  = (~\m4_addr_i[21]  | ~\new_[19609]_ ) & (~\m3_addr_i[21]  | ~\new_[19639]_ );
  assign \new_[15551]_  = (~\m7_addr_i[21]  | ~\new_[18823]_ ) & (~\m0_addr_i[21]  | ~\new_[18731]_ );
  assign \new_[15552]_  = ~\new_[27700]_  & (~\new_[17950]_  | ~\new_[28732]_ );
  assign \new_[15553]_  = ~\new_[28081]_  & (~\new_[17969]_  | ~\new_[28640]_ );
  assign \new_[15554]_  = ~\new_[29470]_  & (~\new_[17965]_  | ~\new_[30205]_ );
  assign \new_[15555]_  = (~\m4_addr_i[20]  | ~\new_[19609]_ ) & (~\m3_addr_i[20]  | ~\new_[19639]_ );
  assign \new_[15556]_  = ~\new_[24363]_  & (~\new_[17964]_  | ~\new_[28535]_ );
  assign \new_[15557]_  = (~\m2_addr_i[19]  | ~\new_[18799]_ ) & (~\m1_addr_i[19]  | ~\new_[18887]_ );
  assign \new_[15558]_  = (~\m4_addr_i[19]  | ~\new_[18146]_ ) & (~\m3_addr_i[19]  | ~\new_[18201]_ );
  assign \new_[15559]_  = ~\new_[27629]_  & (~\new_[17968]_  | ~\new_[30117]_ );
  assign \new_[15560]_  = (~\m4_data_i[2]  | ~\new_[19612]_ ) & (~\m3_data_i[2]  | ~\new_[18862]_ );
  assign \new_[15561]_  = (~\m4_data_i[13]  | ~\new_[19613]_ ) & (~\m3_data_i[13]  | ~\new_[18859]_ );
  assign \new_[15562]_  = ~\new_[28118]_  & (~\new_[17970]_  | ~\new_[28355]_ );
  assign \new_[15563]_  = (~\m2_addr_i[18]  | ~\new_[18799]_ ) & (~\m1_addr_i[18]  | ~\new_[18887]_ );
  assign \new_[15564]_  = ~\new_[17422]_  | (~\new_[30104]_  & ~\new_[5894]_ );
  assign \new_[15565]_  = ~\new_[29278]_  & (~\new_[17949]_  | ~\new_[21555]_ );
  assign \new_[15566]_  = (~\m4_addr_i[18]  | ~\new_[18145]_ ) & (~\m3_addr_i[18]  | ~\new_[19639]_ );
  assign \new_[15567]_  = ~\new_[18669]_  | ~\new_[28010]_  | ~\new_[30221]_  | ~\new_[28114]_ ;
  assign \new_[15568]_  = (~\m2_addr_i[17]  | ~\new_[18799]_ ) & (~\m1_addr_i[17]  | ~\new_[18887]_ );
  assign \new_[15569]_  = (~\m4_addr_i[17]  | ~\new_[18143]_ ) & (~\m3_addr_i[17]  | ~\new_[18201]_ );
  assign \new_[15570]_  = ~\new_[17423]_  | (~\new_[30111]_  & ~\new_[5910]_ );
  assign \new_[15571]_  = ~\new_[18670]_  | ~\new_[28046]_  | ~\new_[29079]_  | ~\new_[29969]_ ;
  assign \new_[15572]_  = ~\new_[21587]_  & (~\new_[17603]_  | ~\new_[29079]_ );
  assign \new_[15573]_  = ~\new_[24332]_  & (~\new_[17605]_  | ~\new_[30135]_ );
  assign \new_[15574]_  = (~\m4_addr_i[16]  | ~\new_[19609]_ ) & (~\m3_addr_i[16]  | ~\new_[19639]_ );
  assign \new_[15575]_  = ~\new_[17424]_  | (~\new_[30318]_  & ~\new_[5967]_ );
  assign \new_[15576]_  = ~\new_[18674]_  | ~\new_[29488]_  | ~\new_[28866]_  | ~\new_[29983]_ ;
  assign \new_[15577]_  = ~\new_[22964]_  & (~\new_[17608]_  | ~\new_[28866]_ );
  assign \new_[15578]_  = ~\new_[24449]_  & (~\new_[17611]_  | ~\new_[30139]_ );
  assign \new_[15579]_  = (~\m2_addr_i[15]  | ~\new_[18799]_ ) & (~\m1_addr_i[15]  | ~\new_[18887]_ );
  assign \new_[15580]_  = (~\m4_addr_i[15]  | ~\new_[18147]_ ) & (~\m3_addr_i[15]  | ~\new_[18201]_ );
  assign \new_[15581]_  = ~\new_[17448]_  | ~\new_[22927]_ ;
  assign \new_[15582]_  = ~\new_[17425]_  | (~\new_[29780]_  & ~\new_[5970]_ );
  assign \new_[15583]_  = ~\new_[21503]_  & (~\new_[17613]_  | ~\new_[28969]_ );
  assign \new_[15584]_  = (~\m2_addr_i[14]  | ~\new_[18799]_ ) & (~\m1_addr_i[14]  | ~\new_[18887]_ );
  assign \new_[15585]_  = ~\new_[22902]_  & (~\new_[17615]_  | ~\new_[29783]_ );
  assign \new_[15586]_  = (~\m4_addr_i[14]  | ~\new_[18145]_ ) & (~\m3_addr_i[14]  | ~\new_[19639]_ );
  assign \new_[15587]_  = ~\new_[17453]_  | ~\new_[22995]_ ;
  assign \new_[15588]_  = ~\new_[26399]_  | (~\new_[17699]_  & ~\new_[29889]_ );
  assign \new_[15589]_  = (~\m2_addr_i[13]  | ~\new_[18799]_ ) & (~\m1_addr_i[13]  | ~\new_[18887]_ );
  assign \new_[15590]_  = ~\new_[21344]_  & (~\new_[17617]_  | ~\new_[28840]_ );
  assign \new_[15591]_  = ~\new_[21575]_  & (~\new_[17618]_  | ~\new_[29922]_ );
  assign \new_[15592]_  = (~\m4_addr_i[13]  | ~\new_[18147]_ ) & (~\m3_addr_i[13]  | ~\new_[18201]_ );
  assign \new_[15593]_  = ~\new_[17459]_  | ~\new_[22863]_ ;
  assign \new_[15594]_  = ~\new_[24347]_  | (~\new_[17729]_  & ~\new_[30038]_ );
  assign \new_[15595]_  = (~\m4_addr_i[12]  | ~\new_[19609]_ ) & (~\m3_addr_i[12]  | ~\new_[18201]_ );
  assign \new_[15596]_  = (~\new_[17865]_  | ~\new_[30432]_ ) & (~\new_[28849]_  | ~\new_[31491]_ );
  assign \new_[15597]_  = ~\new_[18678]_  | ~\new_[27928]_  | ~\new_[30207]_  | ~\new_[30552]_ ;
  assign \new_[15598]_  = ~\new_[17462]_  | (~\new_[30207]_  & ~\new_[31121]_ );
  assign \new_[15599]_  = ~\new_[17426]_  | (~\new_[30005]_  & ~\new_[5900]_ );
  assign \new_[15600]_  = (~\m4_addr_i[11]  | ~\new_[19609]_ ) & (~\m3_addr_i[11]  | ~\new_[19639]_ );
  assign \new_[15601]_  = (~\m2_addr_i[11]  | ~\new_[18799]_ ) & (~\m1_addr_i[11]  | ~\new_[18887]_ );
  assign \new_[15602]_  = ~\new_[22945]_  & (~\new_[17623]_  | ~\new_[30344]_ );
  assign \new_[15603]_  = ~\new_[23035]_  & (~\new_[17625]_  | ~\new_[30294]_ );
  assign \new_[15604]_  = ~\new_[17427]_  | (~\new_[30086]_  & ~\new_[5901]_ );
  assign \new_[15605]_  = ~\new_[17470]_  | ~\new_[22888]_ ;
  assign \new_[15606]_  = (~\m2_addr_i[10]  | ~\new_[18799]_ ) & (~\m1_addr_i[10]  | ~\new_[18887]_ );
  assign \new_[15607]_  = ~\new_[28817]_  | (~\new_[17760]_  & ~\new_[30029]_ );
  assign \new_[15608]_  = (~\m4_addr_i[10]  | ~\new_[18143]_ ) & (~\m3_addr_i[10]  | ~\new_[19639]_ );
  assign \new_[15609]_  = ~\new_[21595]_  & (~\new_[17628]_  | ~\new_[29162]_ );
  assign \new_[15610]_  = ~\new_[23000]_  & (~\new_[17630]_  | ~\new_[30083]_ );
  assign \new_[15611]_  = ~\new_[17428]_  | (~\new_[30178]_  & ~\new_[5984]_ );
  assign \new_[15612]_  = ~\new_[21517]_  & (~\new_[17632]_  | ~\new_[29086]_ );
  assign \new_[15613]_  = ~\new_[18683]_  | ~\new_[28832]_  | ~\new_[29891]_  | ~\new_[29064]_ ;
  assign \new_[15614]_  = (~\m4_addr_i[9]  | ~\new_[18142]_ ) & (~\m3_addr_i[9]  | ~\new_[18201]_ );
  assign \new_[15615]_  = ~\new_[21566]_  & (~\new_[17634]_  | ~\new_[29891]_ );
  assign \new_[15616]_  = (~\m4_addr_i[8]  | ~\new_[18146]_ ) & (~\m3_addr_i[8]  | ~\new_[18201]_ );
  assign \new_[15617]_  = ~\new_[21510]_  & (~\new_[17636]_  | ~\new_[29175]_ );
  assign \new_[15618]_  = ~\new_[18682]_  | ~\new_[30110]_  | ~\new_[29892]_  | ~\new_[30491]_ ;
  assign \new_[15619]_  = (~\m2_addr_i[7]  | ~\new_[18799]_ ) & (~\m1_addr_i[7]  | ~\new_[18887]_ );
  assign \new_[15620]_  = (~\m4_addr_i[7]  | ~\new_[18147]_ ) & (~\m3_addr_i[7]  | ~\new_[18201]_ );
  assign \new_[15621]_  = ~\new_[24412]_  | (~\new_[17839]_  & ~\new_[30275]_ );
  assign \new_[15622]_  = ~\new_[17429]_  | (~\new_[30180]_  & ~\new_[5989]_ );
  assign \new_[15623]_  = (~\m4_addr_i[6]  | ~\new_[18146]_ ) & (~\m3_addr_i[6]  | ~\new_[18201]_ );
  assign \new_[15624]_  = ~\new_[18677]_  | ~\new_[28751]_  | ~\new_[29656]_  | ~\new_[28023]_ ;
  assign \new_[15625]_  = ~\new_[22992]_  & (~\new_[17606]_  | ~\new_[29656]_ );
  assign \new_[15626]_  = (~\m4_addr_i[0]  | ~\new_[18162]_ ) & (~\m3_addr_i[0]  | ~\new_[18198]_ );
  assign \new_[15627]_  = ~\new_[18684]_  | ~\new_[28702]_  | ~\new_[29785]_  | ~\new_[27802]_ ;
  assign \new_[15628]_  = ~\new_[24355]_  & (~\new_[17620]_  | ~\new_[29785]_ );
  assign \new_[15629]_  = (~\m4_addr_i[5]  | ~\new_[18144]_ ) & (~\m3_addr_i[5]  | ~\new_[18201]_ );
  assign \new_[15630]_  = ~\new_[21473]_  & (~\new_[17640]_  | ~\new_[28878]_ );
  assign \new_[15631]_  = (~\m4_addr_i[4]  | ~\new_[19609]_ ) & (~\m3_addr_i[4]  | ~\new_[18201]_ );
  assign \new_[15632]_  = ~\new_[17430]_  | (~\new_[30105]_  & ~\new_[5933]_ );
  assign \new_[15633]_  = ~\new_[23023]_  & (~\new_[17647]_  | ~\new_[30126]_ );
  assign \new_[15634]_  = ~\new_[18688]_  | ~\new_[28502]_  | ~\new_[29913]_  | ~\new_[29537]_ ;
  assign \new_[15635]_  = (~\m4_addr_i[3]  | ~\new_[18144]_ ) & (~\m3_addr_i[3]  | ~\new_[18201]_ );
  assign \new_[15636]_  = ~\new_[17431]_  | (~\new_[30089]_  & ~\new_[5928]_ );
  assign \new_[15637]_  = (~\m4_addr_i[2]  | ~\new_[19609]_ ) & (~\m3_addr_i[2]  | ~\new_[18201]_ );
  assign \new_[15638]_  = ~\new_[17432]_  | (~\new_[30280]_  & ~\new_[5907]_ );
  assign \new_[15639]_  = ~\new_[17471]_  | ~\new_[21994]_ ;
  assign \new_[15640]_  = ~\new_[27548]_  | (~\new_[17806]_  & ~\new_[30201]_ );
  assign \new_[15641]_  = (~\m2_data_i[9]  | ~\new_[19590]_ ) & (~\m1_data_i[9]  | ~\new_[20572]_ );
  assign \new_[15642]_  = ~\new_[22959]_  & (~\new_[17637]_  | ~\new_[30333]_ );
  assign \new_[15643]_  = (~\m2_addr_i[1]  | ~\new_[18799]_ ) & (~\m1_addr_i[1]  | ~\new_[18887]_ );
  assign \new_[15644]_  = ~\new_[18679]_  | ~\new_[29622]_  | ~\new_[30437]_  | ~\new_[30544]_ ;
  assign \new_[15645]_  = (~\m4_addr_i[1]  | ~\new_[18142]_ ) & (~\m3_addr_i[1]  | ~\new_[18201]_ );
  assign \new_[15646]_  = ~\new_[17433]_  | (~\new_[30123]_  & ~\new_[5908]_ );
  assign \new_[15647]_  = ~\new_[17506]_  | ~\new_[22104]_ ;
  assign \new_[15648]_  = ~\new_[26284]_  | (~\new_[17828]_  & ~\new_[30325]_ );
  assign \new_[15649]_  = (~\m2_addr_i[0]  | ~\new_[18799]_ ) & (~\m1_addr_i[0]  | ~\new_[18887]_ );
  assign \new_[15650]_  = ~\new_[18689]_  | ~\new_[28262]_  | ~\new_[30025]_  | ~\new_[28355]_ ;
  assign \new_[15651]_  = ~\new_[24515]_  & (~\new_[17651]_  | ~\new_[30025]_ );
  assign \new_[15652]_  = (~\m4_addr_i[0]  | ~\new_[18143]_ ) & (~\m3_addr_i[0]  | ~\new_[19639]_ );
  assign \new_[15653]_  = (~\m2_sel_i[3]  | ~\new_[18799]_ ) & (~\m1_sel_i[3]  | ~\new_[18887]_ );
  assign \new_[15654]_  = (~\m4_sel_i[3]  | ~\new_[18143]_ ) & (~\m3_sel_i[3]  | ~\new_[19639]_ );
  assign \new_[15655]_  = (~\m4_sel_i[2]  | ~\new_[19609]_ ) & (~\m3_sel_i[2]  | ~\new_[18201]_ );
  assign \new_[15656]_  = (~\m4_sel_i[1]  | ~\new_[19609]_ ) & (~\m3_sel_i[1]  | ~\new_[18201]_ );
  assign \new_[15657]_  = (~\m2_sel_i[1]  | ~\new_[18799]_ ) & (~\m1_sel_i[1]  | ~\new_[18887]_ );
  assign \new_[15658]_  = (~\m7_sel_i[1]  | ~\new_[18823]_ ) & (~\m0_sel_i[1]  | ~\new_[18731]_ );
  assign \new_[15659]_  = (~\m2_sel_i[0]  | ~\new_[18799]_ ) & (~\m1_sel_i[0]  | ~\new_[18887]_ );
  assign \new_[15660]_  = (~\m4_sel_i[0]  | ~\new_[18145]_ ) & (~\m3_sel_i[0]  | ~\new_[18201]_ );
  assign \new_[15661]_  = (~\new_[18577]_  | ~s11_err_i) & (~\new_[17750]_  | ~s8_err_i);
  assign \new_[15662]_  = (~\new_[17756]_  | ~s14_err_i) & (~\new_[18659]_  | ~s12_err_i);
  assign \new_[15663]_  = (~m4_we_i | ~\new_[18144]_ ) & (~m3_we_i | ~\new_[18201]_ );
  assign \new_[15664]_  = (~\new_[18661]_  | ~s5_err_i) & (~\new_[17870]_  | ~s3_err_i);
  assign \new_[15665]_  = (~\new_[17756]_  | ~s14_rty_i) & (~\new_[18659]_  | ~s12_rty_i);
  assign \new_[15666]_  = (~\new_[18577]_  | ~s11_rty_i) & (~\new_[17750]_  | ~s8_rty_i);
  assign \new_[15667]_  = (~\new_[18661]_  | ~s5_rty_i) & (~\new_[17870]_  | ~s3_rty_i);
  assign \new_[15668]_  = (~\m4_data_i[31]  | ~\new_[18877]_ ) & (~\m3_data_i[31]  | ~\new_[18200]_ );
  assign \new_[15669]_  = (~\m5_data_i[30]  | ~\new_[18740]_ ) & (~\m6_data_i[30]  | ~\new_[18786]_ );
  assign \new_[15670]_  = (~\m5_data_i[28]  | ~\new_[18740]_ ) & (~\m6_data_i[28]  | ~\new_[18786]_ );
  assign \new_[15671]_  = (~\m4_data_i[28]  | ~\new_[18877]_ ) & (~\m3_data_i[28]  | ~\new_[19638]_ );
  assign \new_[15672]_  = (~\m4_data_i[27]  | ~\new_[18877]_ ) & (~\m3_data_i[27]  | ~\new_[19638]_ );
  assign \new_[15673]_  = \new_[5964]_  ? \new_[30221]_  : \new_[17895]_ ;
  assign \new_[15674]_  = (~\m5_data_i[26]  | ~\new_[18740]_ ) & (~\m6_data_i[26]  | ~\new_[18786]_ );
  assign \new_[15675]_  = \new_[6246]_  ? \new_[30730]_  : \new_[17897]_ ;
  assign \new_[15676]_  = (~\m4_data_i[26]  | ~\new_[18877]_ ) & (~\m3_data_i[26]  | ~\new_[18200]_ );
  assign \new_[15677]_  = \new_[6246]_  ? \new_[30020]_  : \new_[17898]_ ;
  assign \new_[15678]_  = (~\m7_data_i[26]  | ~\new_[18824]_ ) & (~\m0_data_i[26]  | ~\new_[18010]_ );
  assign \new_[15679]_  = \new_[6038]_  ? \new_[29220]_  : \new_[17900]_ ;
  assign \new_[15680]_  = \new_[6176]_  ? \new_[30135]_  : \new_[17901]_ ;
  assign \new_[15681]_  = \new_[5968]_  ? \new_[30386]_  : \new_[17903]_ ;
  assign \new_[15682]_  = \new_[5913]_  ? \new_[28969]_  : \new_[17904]_ ;
  assign \new_[15683]_  = \new_[6206]_  ? \new_[30255]_  : \new_[17906]_ ;
  assign \new_[15684]_  = (~\m5_data_i[25]  | ~\new_[18740]_ ) & (~\m6_data_i[25]  | ~\new_[18786]_ );
  assign \new_[15685]_  = \new_[5830]_  ? \new_[28840]_  : \new_[17910]_ ;
  assign \new_[15686]_  = \new_[5830]_  ? \new_[29150]_  : \new_[17911]_ ;
  assign \new_[15687]_  = \new_[6031]_  ? \new_[29782]_  : \new_[17908]_ ;
  assign \new_[15688]_  = (~\m5_data_i[24]  | ~\new_[18740]_ ) & (~\m6_data_i[24]  | ~\new_[18786]_ );
  assign \new_[15689]_  = \new_[5979]_  ? \new_[30344]_  : \new_[17913]_ ;
  assign \new_[15690]_  = \new_[5979]_  ? \new_[28870]_  : \new_[17932]_ ;
  assign \new_[15691]_  = \new_[6059]_  ? \new_[30294]_  : \new_[17915]_ ;
  assign \new_[15692]_  = \new_[6059]_  ? \new_[29967]_  : \new_[17927]_ ;
  assign \new_[15693]_  = \new_[6064]_  ? \new_[30636]_  : \new_[17917]_ ;
  assign \new_[15694]_  = \new_[5985]_  ? \new_[29086]_  : \new_[17930]_ ;
  assign \new_[15695]_  = \new_[5985]_  ? \new_[29506]_  : \new_[17928]_ ;
  assign \new_[15696]_  = \new_[6212]_  ? \new_[29891]_  : \new_[17918]_ ;
  assign \new_[15697]_  = \new_[5919]_  ? \new_[29175]_  : \new_[17920]_ ;
  assign \new_[15698]_  = \new_[5919]_  ? \new_[29974]_  : \new_[17921]_ ;
  assign \new_[15699]_  = \new_[6071]_  ? \new_[30600]_  : \new_[17922]_ ;
  assign \new_[15700]_  = \new_[6190]_  ? \new_[29656]_  : \new_[17923]_ ;
  assign \new_[15701]_  = \new_[5991]_  ? \new_[29912]_  : \new_[17902]_ ;
  assign \new_[15702]_  = \new_[5994]_  ? \new_[28878]_  : \new_[17899]_ ;
  assign \new_[15703]_  = \new_[5997]_  ? \new_[28926]_  : \new_[17934]_ ;
  assign \new_[15704]_  = \new_[6001]_  ? \new_[29386]_  : \new_[17926]_ ;
  assign \new_[15705]_  = \new_[5931]_  ? \new_[30333]_  : \new_[17929]_ ;
  assign \new_[15706]_  = (~\m5_data_i[20]  | ~\new_[18740]_ ) & (~\m6_data_i[20]  | ~\new_[18786]_ );
  assign \new_[15707]_  = \new_[5930]_  ? \new_[29927]_  : \new_[17933]_ ;
  assign \new_[15708]_  = \new_[5997]_  ? \new_[30126]_  : \new_[17935]_ ;
  assign \new_[15709]_  = \new_[5932]_  ? \new_[30025]_  : \new_[17937]_ ;
  assign \new_[15710]_  = (~\m4_data_i[19]  | ~\new_[18877]_ ) & (~\m3_data_i[19]  | ~\new_[19638]_ );
  assign \new_[15711]_  = \new_[6007]_  ? \new_[29118]_  : \new_[17938]_ ;
  assign \new_[15712]_  = ~\new_[16902]_  | ~\new_[30409]_ ;
  assign \new_[15713]_  = (~\m4_data_i[18]  | ~\new_[18877]_ ) & (~\m3_data_i[18]  | ~\new_[18200]_ );
  assign \new_[15714]_  = (~\m5_data_i[18]  | ~\new_[18740]_ ) & (~\m6_data_i[18]  | ~\new_[18786]_ );
  assign \new_[15715]_  = (~\new_[18159]_  | ~\m4_addr_i[29] ) & (~\new_[19636]_  | ~\m3_addr_i[29] );
  assign \new_[15716]_  = (~\m5_data_i[17]  | ~\new_[18740]_ ) & (~\m6_data_i[17]  | ~\new_[18786]_ );
  assign \new_[15717]_  = \new_[29479]_  | \new_[16799]_ ;
  assign \new_[15718]_  = ~\new_[16801]_  | ~\new_[30097]_ ;
  assign \new_[15719]_  = ~\new_[17024]_  & ~\new_[24710]_ ;
  assign \new_[15720]_  = ~\new_[28397]_  & (~\new_[20009]_  | ~\new_[18017]_ );
  assign \new_[15721]_  = \new_[27686]_  | \new_[16813]_ ;
  assign \new_[15722]_  = ~\new_[16815]_  | ~\new_[30320]_ ;
  assign \new_[15723]_  = ~\new_[17028]_  & ~\new_[24783]_ ;
  assign \new_[15724]_  = ~\new_[30633]_  & (~\new_[20770]_  | ~\new_[18024]_ );
  assign \new_[15725]_  = ~\new_[26381]_  & (~\new_[17975]_  | ~\new_[30550]_ );
  assign \new_[15726]_  = \new_[28130]_  | \new_[16832]_ ;
  assign \new_[15727]_  = ~\new_[16833]_  | ~\new_[30172]_ ;
  assign \new_[15728]_  = ~\new_[17034]_  & ~\new_[25925]_ ;
  assign \new_[15729]_  = (~\m5_data_i[13]  | ~\new_[18740]_ ) & (~\m6_data_i[13]  | ~\new_[18786]_ );
  assign \new_[15730]_  = ~\new_[30174]_  & (~\new_[18028]_  | ~\new_[26281]_ );
  assign \new_[15731]_  = ~\new_[30253]_  & (~\new_[20755]_  | ~\new_[18029]_ );
  assign \new_[15732]_  = ~\new_[17035]_  & ~\new_[22987]_ ;
  assign \new_[15733]_  = (~\m5_data_i[12]  | ~\new_[18740]_ ) & (~\m6_data_i[12]  | ~\new_[18786]_ );
  assign \new_[15734]_  = ~\new_[26951]_  & (~\new_[17977]_  | ~\new_[29032]_ );
  assign \new_[15735]_  = (~\m5_data_i[11]  | ~\new_[18740]_ ) & (~\m6_data_i[11]  | ~\new_[18786]_ );
  assign \new_[15736]_  = \new_[29430]_  | \new_[16918]_ ;
  assign \new_[15737]_  = ~\new_[16843]_  | ~\new_[29762]_ ;
  assign \new_[15738]_  = (~\m5_data_i[10]  | ~\new_[18740]_ ) & (~\m6_data_i[10]  | ~\new_[18786]_ );
  assign \new_[15739]_  = ~\new_[28479]_  & (~\new_[17972]_  | ~\new_[28837]_ );
  assign \new_[15740]_  = \new_[29206]_  | \new_[16856]_ ;
  assign \new_[15741]_  = ~\new_[17039]_  & ~\new_[28578]_ ;
  assign \new_[15742]_  = ~\new_[30185]_  & (~\new_[18001]_  | ~\new_[28579]_ );
  assign \new_[15743]_  = ~\new_[17040]_  & ~\new_[26314]_ ;
  assign \new_[15744]_  = ~\new_[16782]_  | ~\new_[29682]_ ;
  assign \new_[15745]_  = ~\new_[26419]_  & (~\new_[17979]_  | ~\new_[29212]_ );
  assign \new_[15746]_  = ~\new_[26979]_  & (~\new_[17980]_  | ~\new_[30432]_ );
  assign \new_[15747]_  = ~\new_[28982]_  & (~\new_[18195]_  | ~\new_[28538]_ );
  assign \new_[15748]_  = ~\new_[17074]_  & ~\new_[24469]_ ;
  assign \new_[15749]_  = \new_[6268]_  ? \new_[29825]_  : \new_[18246]_ ;
  assign \new_[15750]_  = (~\m5_data_i[6]  | ~\new_[18740]_ ) & (~\m6_data_i[6]  | ~\new_[18786]_ );
  assign \new_[15751]_  = \new_[26685]_  | \new_[16942]_ ;
  assign \new_[15752]_  = ~\new_[28707]_  & (~\new_[17981]_  | ~\new_[29015]_ );
  assign \new_[15753]_  = \new_[28942]_  | \new_[16890]_ ;
  assign \new_[15754]_  = ~\new_[29331]_  & (~\new_[18122]_  | ~\new_[26768]_ );
  assign \new_[15755]_  = ~\new_[17055]_  & ~\new_[23174]_ ;
  assign \new_[15756]_  = (~\m5_data_i[4]  | ~\new_[18740]_ ) & (~\m6_data_i[4]  | ~\new_[18786]_ );
  assign \new_[15757]_  = \new_[28485]_  | \new_[16899]_ ;
  assign \new_[15758]_  = ~\new_[27388]_  & (~\new_[17984]_  | ~\new_[28967]_ );
  assign \new_[15759]_  = ~\new_[16922]_  | ~\new_[30092]_ ;
  assign \new_[15760]_  = ~\new_[30350]_  & (~\new_[20948]_  | ~\new_[18136]_ );
  assign \new_[15761]_  = ~\new_[26629]_  & (~\new_[17985]_  | ~\new_[29082]_ );
  assign \new_[15762]_  = \new_[31406]_  ? \new_[30293]_  : \new_[18257]_ ;
  assign \new_[15763]_  = \new_[29558]_  | \new_[16871]_ ;
  assign \new_[15764]_  = ~\new_[16830]_  | ~\new_[29888]_ ;
  assign \new_[15765]_  = (~\m5_data_i[1]  | ~\new_[18740]_ ) & (~\m6_data_i[1]  | ~\new_[18786]_ );
  assign \new_[15766]_  = \new_[29319]_  | \new_[16914]_ ;
  assign \new_[15767]_  = ~\new_[29338]_  & (~\new_[17991]_  | ~\new_[30107]_ );
  assign \new_[15768]_  = ~\new_[16915]_  | ~\new_[29863]_ ;
  assign \new_[15769]_  = ~\new_[17027]_  & ~\new_[26257]_ ;
  assign \new_[15770]_  = ~\new_[29916]_  & (~\new_[18120]_  | ~\new_[26538]_ );
  assign \new_[15771]_  = ~\new_[29238]_  & (~\new_[20744]_  | ~\new_[18121]_ );
  assign \new_[15772]_  = ~\new_[17037]_  & ~\new_[23053]_ ;
  assign \new_[15773]_  = ~\new_[27860]_  & (~\new_[17988]_  | ~\new_[30034]_ );
  assign \new_[15774]_  = \new_[26388]_  | \new_[16948]_ ;
  assign \new_[15775]_  = ~\new_[16910]_  | ~\new_[30061]_ ;
  assign \new_[15776]_  = ~\new_[29989]_  & (~\new_[20095]_  | ~\new_[18123]_ );
  assign \new_[15777]_  = \new_[29414]_  | \new_[16962]_ ;
  assign \new_[15778]_  = (~\m2_data_i[2]  | ~\new_[19572]_ ) & (~\m1_data_i[2]  | ~\new_[18191]_ );
  assign \new_[15779]_  = (~\m4_data_i[4]  | ~\new_[19612]_ ) & (~\m3_data_i[4]  | ~\new_[18861]_ );
  assign \new_[15780]_  = \new_[26779]_  | \new_[16862]_ ;
  assign \new_[15781]_  = (~\new_[18877]_  | ~\m4_addr_i[28] ) & (~\new_[18200]_  | ~\m3_addr_i[28] );
  assign \new_[15782]_  = ~\new_[28800]_  & (~\new_[17995]_  | ~\new_[29972]_ );
  assign \new_[15783]_  = \new_[28484]_  | \new_[16958]_ ;
  assign \new_[15784]_  = ~\new_[16964]_  | ~\new_[30159]_ ;
  assign \new_[15785]_  = ~\new_[17064]_  & ~\new_[26439]_ ;
  assign \new_[15786]_  = (~\new_[18877]_  | ~\m4_addr_i[27] ) & (~\new_[18200]_  | ~\m3_addr_i[27] );
  assign \new_[15787]_  = ~\new_[30445]_  & (~\new_[18021]_  | ~\new_[26410]_ );
  assign \new_[15788]_  = ~\new_[29508]_  & (~\new_[20065]_  | ~\new_[18132]_ );
  assign \new_[15789]_  = ~\new_[17066]_  & ~\new_[24341]_ ;
  assign \new_[15790]_  = (~\new_[18877]_  | ~\m4_addr_i[26] ) & (~\new_[18200]_  | ~\m3_addr_i[26] );
  assign \new_[15791]_  = ~m6_stb_i | ~\new_[25239]_  | ~\new_[18089]_ ;
  assign \new_[15792]_  = ~\new_[24662]_  & (~\new_[17996]_  | ~\new_[29701]_ );
  assign \new_[15793]_  = \new_[26311]_  | \new_[16961]_ ;
  assign \new_[15794]_  = ~\new_[29096]_  & (~\new_[18081]_  | ~\new_[28490]_ );
  assign \new_[15795]_  = (~\new_[18877]_  | ~\m4_addr_i[25] ) & (~\new_[18200]_  | ~\m3_addr_i[25] );
  assign \new_[15796]_  = ~\new_[17105]_  & ~\new_[23082]_ ;
  assign \new_[15797]_  = ~\new_[28251]_  & (~\new_[17992]_  | ~\new_[29040]_ );
  assign \new_[15798]_  = ~\new_[30507]_  | (~\new_[20932]_  & ~\new_[18307]_ );
  assign \new_[15799]_  = ~\new_[27993]_  & (~\new_[17994]_  | ~\new_[30723]_ );
  assign \new_[15800]_  = \new_[29156]_  | \new_[16897]_ ;
  assign \new_[15801]_  = (~\m4_data_i[6]  | ~\new_[19613]_ ) & (~\m3_data_i[6]  | ~\new_[18861]_ );
  assign \new_[15802]_  = \new_[17092]_  & \new_[17093]_ ;
  assign \new_[15803]_  = ~\new_[29166]_  & (~\new_[18202]_  | ~\new_[26790]_ );
  assign \new_[15804]_  = ~\new_[17109]_  & ~\new_[23239]_ ;
  assign \new_[15805]_  = (~\m5_addr_i[23]  | ~\new_[18740]_ ) & (~\m6_addr_i[23]  | ~\new_[18786]_ );
  assign \new_[15806]_  = ~\new_[30021]_  | (~\new_[21977]_  & ~\new_[18322]_ );
  assign \new_[15807]_  = (~\m5_addr_i[22]  | ~\new_[18740]_ ) & (~\m6_addr_i[22]  | ~\new_[18786]_ );
  assign \new_[15808]_  = ~\new_[29047]_  & (~\new_[20926]_  | ~\new_[18241]_ );
  assign \new_[15809]_  = \new_[29009]_  | \new_[16945]_ ;
  assign \new_[15810]_  = ~\new_[18558]_  & ~\new_[17316]_ ;
  assign \new_[15811]_  = ~\new_[16864]_  & ~\new_[29959]_ ;
  assign \new_[15812]_  = ~\new_[16891]_  & ~\new_[17319]_ ;
  assign \new_[15813]_  = ~\new_[16901]_  & ~\new_[18272]_ ;
  assign \new_[15814]_  = ~\new_[16881]_  & ~\new_[17304]_ ;
  assign \new_[15815]_  = ~\new_[16847]_  & ~\new_[30188]_ ;
  assign \new_[15816]_  = (~\m4_addr_i[20]  | ~\new_[18877]_ ) & (~\m3_addr_i[20]  | ~\new_[18200]_ );
  assign \new_[15817]_  = ~\new_[16829]_  & ~\new_[17336]_ ;
  assign \new_[15818]_  = (~\m4_data_i[10]  | ~\new_[19614]_ ) & (~\m3_data_i[10]  | ~\new_[18864]_ );
  assign \new_[15819]_  = (~\m5_addr_i[20]  | ~\new_[18740]_ ) & (~\m6_addr_i[20]  | ~\new_[18786]_ );
  assign \new_[15820]_  = ~\new_[16852]_  & ~\new_[30265]_ ;
  assign \new_[15821]_  = ~\new_[17692]_  & ~\new_[17294]_ ;
  assign \new_[15822]_  = ~\new_[18640]_  & ~\new_[17348]_ ;
  assign \new_[15823]_  = \new_[16983]_  | \new_[28301]_ ;
  assign \new_[15824]_  = ~\new_[16984]_  | ~\new_[28412]_ ;
  assign \new_[15825]_  = \new_[16985]_  | \new_[28228]_ ;
  assign \new_[15826]_  = (~\m4_addr_i[19]  | ~\new_[18877]_ ) & (~\m3_addr_i[19]  | ~\new_[18200]_ );
  assign \new_[15827]_  = ~\new_[16986]_  | ~\new_[28222]_ ;
  assign \new_[15828]_  = \new_[16987]_  | \new_[28803]_ ;
  assign \new_[15829]_  = (~\m5_addr_i[19]  | ~\new_[18740]_ ) & (~\m6_addr_i[19]  | ~\new_[18786]_ );
  assign \new_[15830]_  = \new_[16989]_  | \new_[29561]_ ;
  assign \new_[15831]_  = ~\new_[16990]_  | ~\new_[28500]_ ;
  assign \new_[15832]_  = \new_[16991]_  | \new_[28531]_ ;
  assign \new_[15833]_  = \new_[16992]_  | \new_[28576]_ ;
  assign \new_[15834]_  = ~\new_[16993]_  | ~\new_[28181]_ ;
  assign \new_[15835]_  = (~\m4_addr_i[18]  | ~\new_[18877]_ ) & (~\m3_addr_i[18]  | ~\new_[19638]_ );
  assign \new_[15836]_  = (~\new_[18079]_  | ~\m2_addr_i[24] ) & (~\new_[19632]_  | ~\m1_addr_i[24] );
  assign \new_[15837]_  = ~\new_[16994]_  | ~\new_[28579]_ ;
  assign \new_[15838]_  = \new_[17009]_  | \new_[27707]_ ;
  assign \new_[15839]_  = ~\new_[17005]_  | ~\new_[26410]_ ;
  assign \new_[15840]_  = \new_[16997]_  | \new_[27801]_ ;
  assign \new_[15841]_  = ~\new_[16998]_  | ~\new_[28631]_ ;
  assign \new_[15842]_  = \new_[17007]_  | \new_[28221]_ ;
  assign \new_[15843]_  = ~\new_[17006]_  | ~\new_[28575]_ ;
  assign \new_[15844]_  = \new_[17003]_  | \new_[25006]_ ;
  assign \new_[15845]_  = ~\new_[16999]_  | ~\new_[28474]_ ;
  assign \new_[15846]_  = \new_[17002]_  | \new_[28340]_ ;
  assign \new_[15847]_  = ~\new_[17000]_  | ~\new_[26538]_ ;
  assign \new_[15848]_  = \new_[16995]_  | \new_[27663]_ ;
  assign \new_[15849]_  = ~\new_[17008]_  | ~\new_[28373]_ ;
  assign \new_[15850]_  = \new_[17001]_  | \new_[26254]_ ;
  assign \new_[15851]_  = \new_[17010]_  | \new_[28558]_ ;
  assign \new_[15852]_  = ~\new_[16988]_  | ~\new_[28108]_ ;
  assign \new_[15853]_  = \new_[17004]_  | \new_[28584]_ ;
  assign \new_[15854]_  = \new_[16996]_  | \new_[27690]_ ;
  assign \new_[15855]_  = \new_[17011]_  | \new_[27622]_ ;
  assign \new_[15856]_  = (~\m5_addr_i[16]  | ~\new_[18740]_ ) & (~\m6_addr_i[16]  | ~\new_[20550]_ );
  assign \new_[15857]_  = (~\m5_addr_i[15]  | ~\new_[18740]_ ) & (~\m6_addr_i[15]  | ~\new_[18786]_ );
  assign \new_[15858]_  = (~\m5_addr_i[14]  | ~\new_[18740]_ ) & (~\m6_addr_i[14]  | ~\new_[18786]_ );
  assign \new_[15859]_  = ~\new_[28189]_  & (~\new_[21129]_  | ~\new_[18325]_ );
  assign \new_[15860]_  = ~\new_[29218]_  & (~\new_[23399]_  | ~\new_[18327]_ );
  assign \new_[15861]_  = ~\new_[30144]_  & (~\new_[23436]_  | ~\new_[18330]_ );
  assign \new_[15862]_  = (~\m4_sel_i[1]  | ~\new_[18163]_ ) & (~\m3_sel_i[1]  | ~\new_[19636]_ );
  assign \new_[15863]_  = (~\m4_addr_i[11]  | ~\new_[18877]_ ) & (~\m3_addr_i[11]  | ~\new_[18200]_ );
  assign \new_[15864]_  = ~\new_[18207]_  | ~\new_[31357]_  | ~n8649;
  assign \new_[15865]_  = (~\m4_addr_i[10]  | ~\new_[18877]_ ) & (~\m3_addr_i[10]  | ~\new_[18200]_ );
  assign \new_[15866]_  = ~\new_[28754]_  & (~\new_[22230]_  | ~\new_[18333]_ );
  assign \new_[15867]_  = ~\new_[27857]_  & (~\new_[23479]_  | ~\new_[18335]_ );
  assign \new_[15868]_  = (~\m5_addr_i[9]  | ~\new_[18740]_ ) & (~\m6_addr_i[9]  | ~\new_[18786]_ );
  assign \new_[15869]_  = (~\m4_addr_i[7]  | ~\new_[18877]_ ) & (~\m3_addr_i[7]  | ~\new_[18200]_ );
  assign \new_[15870]_  = (~\m5_addr_i[7]  | ~\new_[18740]_ ) & (~\m6_addr_i[7]  | ~\new_[18786]_ );
  assign \new_[15871]_  = ~\new_[28975]_  & (~\new_[23563]_  | ~\new_[18338]_ );
  assign \new_[15872]_  = (~\m5_addr_i[5]  | ~\new_[18740]_ ) & (~\m6_addr_i[5]  | ~\new_[18786]_ );
  assign \new_[15873]_  = ~\new_[18080]_  | ~\new_[30486]_  | ~n8314;
  assign \new_[15874]_  = ~\new_[18033]_  | ~\new_[31360]_  | ~n8659;
  assign \new_[15875]_  = (~\m5_addr_i[3]  | ~\new_[18740]_ ) & (~\m6_addr_i[3]  | ~\new_[18786]_ );
  assign \new_[15876]_  = (~\m5_addr_i[1]  | ~\new_[18740]_ ) & (~\m6_addr_i[1]  | ~\new_[20550]_ );
  assign \new_[15877]_  = ~\new_[30238]_  & (~\new_[23716]_  | ~\new_[18355]_ );
  assign \new_[15878]_  = ~\new_[18027]_  | ~\new_[31283]_  | ~n8514;
  assign \new_[15879]_  = (~\m5_sel_i[3]  | ~\new_[18740]_ ) & (~\m6_sel_i[3]  | ~\new_[18786]_ );
  assign \new_[15880]_  = ~\new_[18111]_  | ~\new_[31241]_  | ~n8444;
  assign \new_[15881]_  = ~\new_[18154]_  | ~\new_[31249]_  | ~n8479;
  assign \new_[15882]_  = (~\m5_sel_i[2]  | ~\new_[18740]_ ) & (~\m6_sel_i[2]  | ~\new_[18786]_ );
  assign \new_[15883]_  = ~\new_[18008]_  | ~\new_[31532]_  | ~n8924;
  assign \new_[15884]_  = ~\new_[29932]_  & (~\new_[20301]_  | ~\new_[18341]_ );
  assign \new_[15885]_  = (~\m5_data_i[31]  | ~\new_[18735]_ ) & (~\m6_data_i[31]  | ~\new_[18048]_ );
  assign \new_[15886]_  = (~\m5_data_i[29]  | ~\new_[18735]_ ) & (~\m6_data_i[29]  | ~\new_[19563]_ );
  assign \new_[15887]_  = ~\new_[28443]_  & (~\new_[23811]_  | ~\new_[18352]_ );
  assign \new_[15888]_  = (~\m5_data_i[26]  | ~\new_[18735]_ ) & (~\m6_data_i[26]  | ~\new_[18051]_ );
  assign \new_[15889]_  = ~\new_[18023]_  | ~\new_[31234]_  | ~n8414;
  assign \new_[15890]_  = (~\m5_data_i[24]  | ~\new_[18735]_ ) & (~\m6_data_i[24]  | ~\new_[18048]_ );
  assign \new_[15891]_  = ~\new_[18192]_  | ~\new_[31316]_  | ~n8589;
  assign \new_[15892]_  = ~\new_[28006]_  & (~\new_[24135]_  | ~\new_[18337]_ );
  assign \new_[15893]_  = ~\new_[30122]_  & (~\new_[21126]_  | ~\new_[18324]_ );
  assign \new_[15894]_  = ~\new_[18095]_  | ~\new_[31527]_  | ~n8909;
  assign \new_[15895]_  = ~\new_[18801]_  | ~\new_[31247]_  | ~n8469;
  assign \new_[15896]_  = ~\new_[26245]_  | ~\new_[17786]_ ;
  assign \new_[15897]_  = ~\new_[18849]_  | ~\new_[31288]_  | ~n8534;
  assign \new_[15898]_  = ~\new_[18880]_  | ~\new_[31243]_  | ~n8454;
  assign \new_[15899]_  = ~\new_[18823]_  | ~\new_[31367]_  | ~n8689;
  assign \new_[15900]_  = ~\new_[18738]_  | ~\new_[31343]_  | ~n8619;
  assign \new_[15901]_  = ~m0_stb_i | ~\new_[26918]_  | ~\new_[18732]_ ;
  assign \new_[15902]_  = ~m1_stb_i | ~\new_[27538]_  | ~\new_[18887]_ ;
  assign \new_[15903]_  = ~\new_[18927]_  | ~\new_[31344]_  | ~n8624;
  assign \new_[15904]_  = ~\new_[18886]_  | ~\new_[31381]_  | ~n8749;
  assign \new_[15905]_  = ~\new_[18737]_  | ~\new_[31239]_  | ~n8434;
  assign \new_[15906]_  = ~\new_[16305]_  | ~\new_[31379]_  | ~n8739;
  assign \new_[15907]_  = ~\new_[18740]_  | ~\new_[31377]_  | ~n8734;
  assign \new_[15908]_  = ~\new_[14837]_  | ~\new_[31386]_  | ~n8769;
  assign \new_[15909]_  = ~\new_[18808]_  | ~\new_[31248]_  | ~n8474;
  assign \new_[15910]_  = ~\new_[18826]_  | ~\new_[31395]_  | ~n8789;
  assign \new_[15911]_  = ~\new_[18735]_  | ~\new_[30490]_  | ~n8329;
  assign \new_[15912]_  = ~\new_[18739]_  | ~\new_[31372]_  | ~n8714;
  assign \new_[15913]_  = \new_[17650]_  & \new_[29350]_ ;
  assign \new_[15914]_  = ~\new_[28677]_  & (~\new_[21145]_  | ~\new_[19190]_ );
  assign \new_[15915]_  = ~\new_[29977]_  | (~\new_[19113]_  & ~\new_[21194]_ );
  assign \new_[15916]_  = ~\new_[30434]_  | (~\new_[19116]_  & ~\new_[23859]_ );
  assign \new_[15917]_  = ~\new_[28905]_  | (~\new_[19114]_  & ~\new_[22340]_ );
  assign \new_[15918]_  = ~\new_[30784]_  | (~\new_[19111]_  & ~\new_[22254]_ );
  assign \new_[15919]_  = ~\new_[30707]_  | (~\new_[19118]_  & ~\new_[20348]_ );
  assign \new_[15920]_  = ~\new_[30598]_  & (~\new_[21635]_  | ~\new_[18962]_ );
  assign \new_[15921]_  = ~\new_[30287]_  & (~\new_[20004]_  | ~\new_[18974]_ );
  assign \new_[15922]_  = ~\new_[30109]_  & (~\new_[21683]_  | ~\new_[18983]_ );
  assign \new_[15923]_  = (~\m4_addr_i[12]  | ~\new_[19614]_ ) & (~\m3_addr_i[12]  | ~\new_[18863]_ );
  assign \new_[15924]_  = ~\new_[30515]_  & (~\new_[21909]_  | ~\new_[19014]_ );
  assign \new_[15925]_  = ~\new_[26518]_  & (~\new_[19142]_  | ~\new_[30061]_ );
  assign \new_[15926]_  = ~\new_[28204]_  & (~\new_[21984]_  | ~\new_[19102]_ );
  assign \new_[15927]_  = ~\new_[29671]_  & (~\new_[20985]_  | ~\new_[19095]_ );
  assign \new_[15928]_  = ~\new_[30309]_  & (~\new_[21936]_  | ~\new_[19055]_ );
  assign \new_[15929]_  = ~\new_[30445]_  & (~\new_[20987]_  | ~\new_[19096]_ );
  assign \new_[15930]_  = ~\new_[30157]_  & (~\new_[21968]_  | ~\new_[19076]_ );
  assign \new_[15931]_  = ~\new_[30047]_  & (~\new_[21972]_  | ~\new_[19100]_ );
  assign \new_[15932]_  = \new_[19005]_  ? \new_[30597]_  : \new_[31438]_ ;
  assign \new_[15933]_  = ~\new_[29172]_  & (~\new_[21003]_  | ~\new_[19107]_ );
  assign \new_[15934]_  = \new_[18964]_  ? \new_[30540]_  : \new_[6174]_ ;
  assign \new_[15935]_  = \new_[6203]_  ? \new_[29911]_  : \new_[18971]_ ;
  assign \new_[15936]_  = ~\new_[22961]_  | ~\new_[17669]_ ;
  assign \new_[15937]_  = ~\new_[24328]_  | ~\new_[17691]_ ;
  assign \new_[15938]_  = \new_[6053]_  ? \new_[29771]_  : \new_[19000]_ ;
  assign \new_[15939]_  = (~\m4_addr_i[10]  | ~\new_[19614]_ ) & (~\m3_addr_i[10]  | ~\new_[18863]_ );
  assign \new_[15940]_  = (~\new_[19206]_  | ~\new_[30104]_ ) & (~\new_[29676]_  | ~\new_[6202]_ );
  assign \new_[15941]_  = \new_[6035]_  ? \new_[30221]_  : \new_[18968]_ ;
  assign \new_[15942]_  = \new_[6039]_  ? \new_[29079]_  : \new_[18978]_ ;
  assign \new_[15943]_  = (~\new_[19216]_  | ~\new_[30280]_ ) & (~\new_[29582]_  | ~\new_[6087]_ );
  assign \new_[15944]_  = (~\new_[18986]_  | ~\new_[30318]_ ) & (~\new_[30575]_  | ~\new_[6043]_ );
  assign \new_[15945]_  = \new_[6044]_  ? \new_[28866]_  : \new_[18988]_ ;
  assign \new_[15946]_  = (~\m2_data_i[21]  | ~\new_[19571]_ ) & (~\m1_data_i[21]  | ~\new_[19630]_ );
  assign \new_[15947]_  = \new_[6047]_  ? \new_[28969]_  : \new_[18981]_ ;
  assign \new_[15948]_  = \new_[5973]_  ? \new_[28840]_  : \new_[19006]_ ;
  assign \new_[15949]_  = (~\new_[19209]_  | ~\new_[30409]_ ) & (~\new_[29576]_  | ~\new_[31423]_ );
  assign \new_[15950]_  = (~\new_[19004]_  | ~\new_[30146]_ ) & (~\new_[30443]_  | ~\new_[6208]_ );
  assign \new_[15951]_  = (~\new_[19042]_  | ~\new_[29682]_ ) & (~\new_[30068]_  | ~\new_[31235]_ );
  assign \new_[15952]_  = (~\new_[19212]_  | ~\new_[30005]_ ) & (~\new_[29089]_  | ~\new_[6056]_ );
  assign \new_[15953]_  = \new_[6058]_  ? \new_[30344]_  : \new_[19071]_ ;
  assign \new_[15954]_  = (~\new_[19213]_  | ~\new_[30086]_ ) & (~\new_[29639]_  | ~\new_[6062]_ );
  assign \new_[15955]_  = \new_[6063]_  ? \new_[29162]_  : \new_[19024]_ ;
  assign \new_[15956]_  = \new_[6068]_  ? \new_[29086]_  : \new_[19049]_ ;
  assign \new_[15957]_  = (~\new_[19066]_  | ~\new_[30180]_ ) & (~\new_[30661]_  | ~\new_[6073]_ );
  assign \new_[15958]_  = \new_[6077]_  ? \new_[28878]_  : \new_[19101]_ ;
  assign \new_[15959]_  = \new_[6268]_  ? \new_[30138]_  : \new_[19059]_ ;
  assign \new_[15960]_  = \new_[6081]_  ? \new_[30126]_  : \new_[19081]_ ;
  assign \new_[15961]_  = (~\new_[19064]_  | ~\new_[30089]_ ) & (~\new_[30543]_  | ~\new_[6186]_ );
  assign \new_[15962]_  = \new_[6003]_  ? \new_[30333]_  : \new_[19074]_ ;
  assign \new_[15963]_  = (~\new_[19215]_  | ~\new_[30105]_ ) & (~\new_[29606]_  | ~\new_[6080]_ );
  assign \new_[15964]_  = (~\new_[19220]_  | ~\new_[30123]_ ) & (~\new_[29333]_  | ~\new_[6091]_ );
  assign \new_[15965]_  = \new_[6006]_  ? \new_[30025]_  : \new_[19104]_ ;
  assign \new_[15966]_  = (~\new_[18967]_  | ~\new_[29874]_ ) & (~\new_[26038]_  | ~\new_[29874]_ );
  assign \new_[15967]_  = (~\new_[18977]_  | ~\new_[30215]_ ) & (~\new_[26440]_  | ~\new_[30215]_ );
  assign \new_[15968]_  = (~\new_[19052]_  | ~\new_[30508]_ ) & (~\new_[29450]_  | ~\new_[30508]_ );
  assign \new_[15969]_  = (~\new_[18987]_  | ~\new_[29260]_ ) & (~\new_[24852]_  | ~\new_[29260]_ );
  assign \new_[15970]_  = (~\new_[19021]_  | ~\new_[29692]_ ) & (~\new_[24760]_  | ~\new_[29692]_ );
  assign \new_[15971]_  = (~\new_[19012]_  | ~\new_[29977]_ ) & (~\new_[24596]_  | ~\new_[29977]_ );
  assign \new_[15972]_  = (~\new_[18979]_  | ~\new_[30774]_ ) & (~\new_[27570]_  | ~\new_[30774]_ );
  assign \new_[15973]_  = (~\new_[19056]_  | ~\new_[29233]_ ) & (~\new_[27680]_  | ~\new_[29233]_ );
  assign \new_[15974]_  = ~\new_[30167]_  & (~\new_[19027]_  | ~\new_[27914]_ );
  assign \new_[15975]_  = (~\new_[19023]_  | ~\new_[29139]_ ) & (~\new_[26321]_  | ~\new_[29139]_ );
  assign \new_[15976]_  = (~\new_[19054]_  | ~\new_[29887]_ ) & (~\new_[26383]_  | ~\new_[29887]_ );
  assign \new_[15977]_  = (~\new_[19041]_  | ~\new_[28905]_ ) & (~\new_[23136]_  | ~\new_[28905]_ );
  assign \new_[15978]_  = (~\new_[19067]_  | ~\new_[30147]_ ) & (~\new_[23110]_  | ~\new_[30147]_ );
  assign \new_[15979]_  = (~\new_[19002]_  | ~\new_[30125]_ ) & (~\new_[23163]_  | ~\new_[30125]_ );
  assign \new_[15980]_  = (~\new_[18993]_  | ~\new_[30316]_ ) & (~\new_[26163]_  | ~\new_[30316]_ );
  assign \new_[15981]_  = (~\new_[19015]_  | ~\new_[29560]_ ) & (~\new_[26289]_  | ~\new_[29560]_ );
  assign \new_[15982]_  = (~\new_[19093]_  | ~\new_[30610]_ ) & (~\new_[26310]_  | ~\new_[30610]_ );
  assign \new_[15983]_  = (~\new_[19103]_  | ~\new_[30021]_ ) & (~\new_[26293]_  | ~\new_[30021]_ );
  assign \new_[15984]_  = ~\new_[22167]_  & (~\new_[18769]_  | ~\new_[30573]_ );
  assign \new_[15985]_  = ~\new_[23768]_  & (~\new_[18870]_  | ~\new_[30814]_ );
  assign \new_[15986]_  = (~\m4_sel_i[2]  | ~\new_[19614]_ ) & (~\m3_sel_i[2]  | ~\new_[18857]_ );
  assign \new_[15987]_  = (~\m4_sel_i[1]  | ~\new_[19614]_ ) & (~\m3_sel_i[1]  | ~\new_[18863]_ );
  assign \new_[15988]_  = ~\new_[21049]_  | ~\new_[20357]_  | ~\m7_addr_i[5]  | ~\new_[21241]_ ;
  assign \new_[15989]_  = ~\m5_addr_i[5]  | ~\new_[20357]_  | ~\new_[20355]_  | ~\new_[21241]_ ;
  assign \new_[15990]_  = ~\new_[31991]_  & ~\new_[31782]_ ;
  assign \new_[15991]_  = ~\new_[18135]_  & ~\new_[31671]_ ;
  assign \new_[15992]_  = ~\new_[31991]_  & ~\new_[31585]_ ;
  assign \new_[15993]_  = ~\new_[31747]_  & ~\new_[18135]_ ;
  assign \new_[15994]_  = ~\new_[18279]_  & ~\new_[31703]_ ;
  assign \new_[15995]_  = ~\new_[18308]_  & ~\new_[31874]_ ;
  assign \new_[15996]_  = ~\new_[18279]_  & ~\new_[31592]_ ;
  assign \new_[15997]_  = ~\new_[32308]_  & ~\new_[31647]_ ;
  assign \new_[15998]_  = ~\new_[32308]_  & ~\new_[31812]_ ;
  assign \new_[15999]_  = ~\new_[26839]_  | ~\new_[18229]_  | ~\new_[22387]_ ;
  assign \new_[16000]_  = ~\new_[28541]_  | ~\new_[18238]_  | ~\new_[22321]_ ;
  assign \new_[16001]_  = ~\new_[27602]_  | ~\new_[18248]_  | ~\new_[22195]_ ;
  assign \new_[16002]_  = ~\new_[28186]_  | ~\new_[18283]_  | ~\new_[22171]_ ;
  assign \new_[16003]_  = ~\new_[28510]_  | ~\new_[18250]_  | ~\new_[22202]_ ;
  assign \new_[16004]_  = ~\new_[28420]_  | ~\new_[18264]_  | ~\new_[21260]_ ;
  assign \new_[16005]_  = ~\new_[28574]_  | ~\new_[18269]_  | ~\new_[21216]_ ;
  assign \new_[16006]_  = ~\new_[28554]_  | ~\new_[18275]_  | ~\new_[22268]_ ;
  assign \new_[16007]_  = ~\new_[28384]_  | ~\new_[18298]_  | ~\new_[22366]_ ;
  assign \new_[16008]_  = ~\new_[27130]_  | ~\new_[18293]_  | ~\new_[20358]_ ;
  assign \new_[16009]_  = ~\new_[28291]_  | ~\new_[18288]_  | ~\new_[22330]_ ;
  assign \new_[16010]_  = ~\new_[28606]_  | ~\new_[18318]_  | ~\new_[21205]_ ;
  assign \new_[16011]_  = ~\new_[28294]_  | ~\new_[18297]_  | ~\new_[22430]_ ;
  assign \new_[16012]_  = ~\new_[28346]_  | ~\new_[18321]_  | ~\new_[21252]_ ;
  assign \new_[16013]_  = ~\new_[28193]_  | ~\new_[18323]_  | ~\new_[21173]_ ;
  assign \new_[16014]_  = \new_[21285]_  & \new_[18217]_ ;
  assign \new_[16015]_  = \new_[18365]_  | \new_[26513]_ ;
  assign \new_[16016]_  = \new_[21316]_  & \new_[18209]_ ;
  assign \new_[16017]_  = \new_[18140]_  & \new_[24162]_ ;
  assign \new_[16018]_  = ~\new_[27613]_  | ~\new_[18340]_  | ~\new_[22288]_ ;
  assign \new_[16019]_  = ~m4_stb_i | ~\new_[19614]_  | ~\new_[28392]_ ;
  assign \new_[16020]_  = \new_[18312]_  & \new_[31853]_ ;
  assign \new_[16021]_  = ~\new_[18230]_  & ~\new_[24710]_ ;
  assign \new_[16022]_  = ~\new_[26822]_  | ~\new_[18349]_  | ~\new_[22383]_ ;
  assign \new_[16023]_  = ~\new_[28139]_  | ~\new_[18343]_  | ~\new_[25059]_ ;
  assign \new_[16024]_  = ~\new_[22276]_  & (~\new_[19248]_  | ~\new_[23020]_ );
  assign \new_[16025]_  = \new_[23890]_  & \new_[18210]_ ;
  assign \new_[16026]_  = \new_[18022]_  & \new_[24471]_ ;
  assign \new_[16027]_  = \new_[18364]_  | \new_[24431]_ ;
  assign \new_[16028]_  = \new_[22471]_  & \new_[18211]_ ;
  assign \new_[16029]_  = ~\new_[18236]_  | ~\new_[31564]_ ;
  assign \new_[16030]_  = ~\new_[18239]_  & ~\new_[24783]_ ;
  assign \new_[16031]_  = ~\new_[27758]_  | ~\new_[18326]_  | ~\new_[22135]_ ;
  assign \new_[16032]_  = ~\new_[28525]_  | ~\new_[18328]_  | ~\new_[24843]_ ;
  assign \new_[16033]_  = (~\m4_addr_i[13]  | ~\new_[19614]_ ) & (~\m3_addr_i[13]  | ~\new_[18858]_ );
  assign \new_[16034]_  = ~\new_[18299]_  | ~\new_[31597]_ ;
  assign \new_[16035]_  = ~m2_stb_i | ~\new_[19565]_  | ~\new_[28714]_ ;
  assign \new_[16036]_  = \new_[23908]_  & \new_[18212]_ ;
  assign \new_[16037]_  = \new_[18025]_  & \new_[23413]_ ;
  assign \new_[16038]_  = ~\new_[18245]_  | ~\new_[31846]_ ;
  assign \new_[16039]_  = ~\new_[18249]_  & ~\new_[25925]_ ;
  assign \new_[16040]_  = ~\new_[26735]_  | ~\new_[18329]_  | ~\new_[22181]_ ;
  assign \new_[16041]_  = ~\new_[28551]_  | ~\new_[18331]_  | ~\new_[24867]_ ;
  assign \new_[16042]_  = \new_[18362]_  | \new_[26341]_ ;
  assign \new_[16043]_  = ~\new_[24461]_  | ~\new_[18342]_  | ~\new_[24836]_ ;
  assign \new_[16044]_  = \new_[18361]_  | \new_[25975]_ ;
  assign \new_[16045]_  = \new_[21273]_  & \new_[18208]_ ;
  assign \new_[16046]_  = \new_[18000]_  & \new_[24450]_ ;
  assign \new_[16047]_  = ~\new_[18254]_  & ~\new_[24771]_ ;
  assign \new_[16048]_  = ~\new_[27608]_  | ~\new_[18332]_  | ~\new_[22184]_ ;
  assign \new_[16049]_  = ~\new_[22187]_  & (~\new_[19257]_  | ~\new_[23068]_ );
  assign \new_[16050]_  = \new_[21278]_  & \new_[18215]_ ;
  assign \new_[16051]_  = ~m6_stb_i | ~\new_[18087]_  | ~\new_[29954]_ ;
  assign \new_[16052]_  = \new_[22481]_  & \new_[18214]_ ;
  assign \new_[16053]_  = ~s3_ack_i | ~\new_[18051]_  | ~\new_[30429]_ ;
  assign \new_[16054]_  = ~s3_err_i | ~\new_[19563]_  | ~\new_[30429]_ ;
  assign \new_[16055]_  = ~s3_rty_i | ~\new_[18051]_  | ~\new_[30429]_ ;
  assign \new_[16056]_  = \new_[18225]_  & \new_[31888]_ ;
  assign \new_[16057]_  = ~s5_ack_i | ~\new_[19565]_  | ~\new_[28714]_ ;
  assign \new_[16058]_  = ~s12_ack_i | ~\new_[18067]_  | ~\new_[30626]_ ;
  assign \new_[16059]_  = ~s13_ack_i | ~\new_[18801]_  | ~\new_[32056]_ ;
  assign \new_[16060]_  = ~\new_[27641]_  | ~\new_[18350]_  | ~\new_[22255]_ ;
  assign \new_[16061]_  = \new_[23921]_  & \new_[18221]_ ;
  assign \new_[16062]_  = ~s11_ack_i | ~\new_[18119]_  | ~\new_[29876]_ ;
  assign \new_[16063]_  = ~s5_err_i | ~\new_[19565]_  | ~\new_[28714]_ ;
  assign \new_[16064]_  = ~s12_err_i | ~\new_[18067]_  | ~\new_[30626]_ ;
  assign \new_[16065]_  = ~\new_[27632]_  | ~\new_[18334]_  | ~\new_[22319]_ ;
  assign \new_[16066]_  = \new_[18082]_  & \new_[26359]_ ;
  assign \new_[16067]_  = ~s11_err_i | ~\new_[18119]_  | ~\new_[29876]_ ;
  assign \new_[16068]_  = ~s5_rty_i | ~\new_[19565]_  | ~\new_[28714]_ ;
  assign \new_[16069]_  = ~s1_rty_i | ~\new_[18799]_  | ~\new_[30357]_ ;
  assign \new_[16070]_  = ~s11_rty_i | ~\new_[18119]_  | ~\new_[29876]_ ;
  assign \new_[16071]_  = ~s13_rty_i | ~\new_[18801]_  | ~\new_[32056]_ ;
  assign \new_[16072]_  = ~s12_rty_i | ~\new_[18067]_  | ~\new_[30626]_ ;
  assign \new_[16073]_  = ~m2_stb_i | ~\new_[20555]_  | ~\new_[30193]_ ;
  assign \new_[16074]_  = \new_[18084]_  & \new_[24356]_ ;
  assign \new_[16075]_  = ~\new_[24431]_  & (~\new_[19263]_  | ~\new_[29817]_ );
  assign \new_[16076]_  = \new_[21590]_  & \new_[18219]_ ;
  assign \new_[16077]_  = \new_[18010]_  & \new_[29625]_ ;
  assign \new_[16078]_  = \new_[18267]_  & \new_[31576]_ ;
  assign \new_[16079]_  = \new_[18023]_  & \new_[29603]_ ;
  assign \new_[16080]_  = \new_[18363]_  | \new_[24668]_ ;
  assign \new_[16081]_  = \new_[18088]_  & \new_[23078]_ ;
  assign \new_[16082]_  = \new_[18360]_  | \new_[26617]_ ;
  assign \new_[16083]_  = \new_[18273]_  & \new_[31759]_ ;
  assign \new_[16084]_  = ~\new_[27621]_  | ~\new_[18336]_  | ~\new_[22259]_ ;
  assign \new_[16085]_  = ~\new_[22270]_  & (~\new_[19274]_  | ~\new_[23014]_ );
  assign \new_[16086]_  = ~\new_[28743]_  | ~\new_[18351]_  | ~\new_[25106]_ ;
  assign \new_[16087]_  = \new_[18137]_  & \new_[21584]_ ;
  assign \new_[16088]_  = ~\new_[18281]_  | ~\new_[31935]_ ;
  assign \new_[16089]_  = \new_[23911]_  & \new_[18216]_ ;
  assign \new_[16090]_  = ~\new_[18242]_  & ~\new_[25602]_ ;
  assign \new_[16091]_  = \new_[18359]_  | \new_[25674]_ ;
  assign \new_[16092]_  = ~\new_[18276]_  & ~\new_[24661]_ ;
  assign \new_[16093]_  = \new_[18131]_  & \new_[22891]_ ;
  assign \new_[16094]_  = ~\new_[18277]_  & ~\new_[26345]_ ;
  assign \new_[16095]_  = ~\new_[28564]_  | (~\new_[19273]_  & ~\new_[30075]_ );
  assign \new_[16096]_  = ~m4_stb_i | ~\new_[18149]_  | ~\new_[29953]_ ;
  assign \new_[16097]_  = \new_[18126]_  & \new_[24081]_ ;
  assign \new_[16098]_  = ~\new_[18261]_  | ~\new_[31575]_ ;
  assign \new_[16099]_  = ~\new_[28429]_  | ~\new_[18353]_  | ~\new_[22218]_ ;
  assign \new_[16100]_  = ~\new_[18285]_  & ~\new_[26257]_ ;
  assign \new_[16101]_  = ~m6_stb_i | ~\new_[18035]_  | ~\new_[29706]_ ;
  assign \new_[16102]_  = ~\new_[18311]_  & ~\new_[26439]_ ;
  assign \new_[16103]_  = ~m2_stb_i | ~\new_[19590]_  | ~\new_[29876]_ ;
  assign \new_[16104]_  = ~\new_[27644]_  | ~\new_[18345]_  | ~\new_[22349]_ ;
  assign \new_[16105]_  = \new_[22537]_  & \new_[18218]_ ;
  assign \new_[16106]_  = \new_[18118]_  & \new_[22926]_ ;
  assign \new_[16107]_  = \new_[18134]_  & \new_[24213]_ ;
  assign \new_[16108]_  = ~\new_[27993]_  & (~\new_[19277]_  | ~\new_[30723]_ );
  assign \new_[16109]_  = ~m4_stb_i | ~\new_[19615]_  | ~\new_[29317]_ ;
  assign \new_[16110]_  = ~m6_stb_i | ~\new_[18043]_  | ~\new_[32134]_ ;
  assign \new_[16111]_  = \new_[18139]_  & \new_[23122]_ ;
  assign \new_[16112]_  = ~s1_ack_i | ~\new_[18143]_  | ~\new_[29779]_ ;
  assign \new_[16113]_  = ~s11_ack_i | ~\new_[18149]_  | ~\new_[29953]_ ;
  assign \new_[16114]_  = ~s10_ack_i | ~\new_[18157]_  | ~\new_[29012]_ ;
  assign \new_[16115]_  = ~s12_ack_i | ~\new_[19615]_  | ~\new_[29317]_ ;
  assign \new_[16116]_  = ~s1_err_i | ~\new_[18142]_  | ~\new_[29779]_ ;
  assign \new_[16117]_  = ~s11_err_i | ~\new_[18149]_  | ~\new_[29953]_ ;
  assign \new_[16118]_  = ~s9_err_i | ~\new_[18154]_  | ~\new_[29185]_ ;
  assign \new_[16119]_  = ~s10_err_i | ~\new_[19611]_  | ~\new_[29012]_ ;
  assign \new_[16120]_  = ~s1_rty_i | ~\new_[18143]_  | ~\new_[29779]_ ;
  assign \new_[16121]_  = ~s11_rty_i | ~\new_[18149]_  | ~\new_[29953]_ ;
  assign \new_[16122]_  = ~s10_rty_i | ~\new_[18157]_  | ~\new_[29012]_ ;
  assign \new_[16123]_  = ~m6_stb_i | ~\new_[18051]_  | ~\new_[30429]_ ;
  assign \new_[16124]_  = ~\new_[27555]_  & (~\new_[19284]_  | ~\new_[28850]_ );
  assign \new_[16125]_  = ~\new_[28564]_  | ~\new_[18344]_  | ~\new_[21172]_ ;
  assign \new_[16126]_  = \new_[18205]_  & \new_[23120]_ ;
  assign \new_[16127]_  = \new_[23079]_  & \new_[18220]_ ;
  assign \new_[16128]_  = \new_[21286]_  & \new_[18213]_ ;
  assign \new_[16129]_  = ~\new_[24276]_  & (~\new_[19275]_  | ~\new_[28183]_ );
  assign \new_[16130]_  = \new_[18348]_  | \new_[22978]_ ;
  assign \new_[16131]_  = \new_[18356]_  | \new_[26187]_ ;
  assign \new_[16132]_  = \new_[18339]_  | \new_[26568]_ ;
  assign \new_[16133]_  = \new_[18346]_  | \new_[26504]_ ;
  assign \new_[16134]_  = \new_[18347]_  | \new_[24002]_ ;
  assign \new_[16135]_  = \new_[17999]_  | \new_[23334]_ ;
  assign \new_[16136]_  = ~\new_[18224]_  | ~\new_[23064]_ ;
  assign \new_[16137]_  = ~\new_[29625]_  | ~\new_[18010]_  | ~s2_ack_i;
  assign \new_[16138]_  = ~m7_stb_i | ~\new_[19584]_  | ~\new_[27855]_ ;
  assign \new_[16139]_  = ~m1_stb_i | ~\new_[19632]_  | ~\new_[28842]_ ;
  assign \new_[16140]_  = ~s5_err_i | ~\new_[18871]_  | ~\new_[28136]_ ;
  assign \new_[16141]_  = ~s11_rty_i | ~\new_[19547]_  | ~\new_[30311]_ ;
  assign \new_[16142]_  = ~s5_rty_i | ~\new_[18871]_  | ~\new_[28136]_ ;
  assign \new_[16143]_  = ~\new_[30287]_  & (~\new_[19333]_  | ~\new_[29483]_ );
  assign \new_[16144]_  = ~\new_[28726]_  | ~\new_[18020]_  | ~s13_ack_i;
  assign \new_[16145]_  = ~\new_[18305]_  | ~\new_[25315]_ ;
  assign \new_[16146]_  = ~s6_err_i | ~\new_[18206]_  | ~\new_[29939]_ ;
  assign \new_[16147]_  = ~\new_[18294]_  | ~\new_[23088]_ ;
  assign \new_[16148]_  = ~\new_[18243]_  | ~\new_[26274]_ ;
  assign \new_[16149]_  = ~m7_stb_i | ~\new_[18835]_  | ~\new_[29534]_ ;
  assign \new_[16150]_  = ~\new_[30335]_  | ~\new_[19554]_  | ~s4_ack_i;
  assign \new_[16151]_  = ~s12_rty_i | ~\new_[18198]_  | ~\new_[30298]_ ;
  assign \new_[16152]_  = ~s13_ack_i | ~\new_[19587]_  | ~\new_[32338]_ ;
  assign \new_[16153]_  = ~\new_[18251]_  | ~\new_[22899]_ ;
  assign \new_[16154]_  = ~\new_[18255]_  | ~\new_[23084]_ ;
  assign \new_[16155]_  = ~\new_[18223]_  | ~\new_[22934]_ ;
  assign \new_[16156]_  = ~\new_[27985]_  | ~\new_[18066]_  | ~s7_ack_i;
  assign \new_[16157]_  = \new_[18071]_  | \new_[22214]_ ;
  assign \new_[16158]_  = ~\new_[26362]_  | ~\new_[18259]_  | ~\new_[23589]_ ;
  assign \new_[16159]_  = ~\new_[30026]_  | ~\new_[18083]_  | ~s14_ack_i;
  assign \new_[16160]_  = ~\new_[24885]_  & (~\new_[19139]_  | ~\new_[29762]_ );
  assign \new_[16161]_  = ~m1_stb_i | ~\new_[18913]_  | ~\new_[30031]_ ;
  assign \new_[16162]_  = ~\new_[22260]_  & (~\new_[19295]_  | ~\new_[27901]_ );
  assign \new_[16163]_  = ~\new_[18271]_  | ~\new_[22137]_ ;
  assign \new_[16164]_  = ~m3_stb_i | ~\new_[18846]_  | ~\new_[29428]_ ;
  assign \new_[16165]_  = ~\new_[29241]_  | ~\new_[19643]_  | ~m0_stb_i;
  assign \new_[16166]_  = ~m1_stb_i | ~\new_[18167]_  | ~\new_[29670]_ ;
  assign \new_[16167]_  = ~\new_[29573]_  & (~\new_[19286]_  | ~\new_[26392]_ );
  assign \new_[16168]_  = ~s9_ack_i | ~\new_[18111]_  | ~\new_[29905]_ ;
  assign \new_[16169]_  = ~s5_ack_i | ~\new_[18835]_  | ~\new_[29534]_ ;
  assign \new_[16170]_  = ~s5_err_i | ~\new_[18835]_  | ~\new_[29534]_ ;
  assign \new_[16171]_  = ~s1_err_i | ~\new_[18823]_  | ~\new_[30124]_ ;
  assign \new_[16172]_  = ~s9_err_i | ~\new_[18111]_  | ~\new_[29905]_ ;
  assign \new_[16173]_  = ~s5_rty_i | ~\new_[18835]_  | ~\new_[29534]_ ;
  assign \new_[16174]_  = ~\new_[18303]_  | ~\new_[25660]_ ;
  assign \new_[16175]_  = ~s13_rty_i | ~\new_[18114]_  | ~\new_[32338]_ ;
  assign \new_[16176]_  = ~s9_rty_i | ~\new_[18111]_  | ~\new_[29905]_ ;
  assign \new_[16177]_  = ~s2_rty_i | ~\new_[18824]_  | ~\new_[30113]_ ;
  assign \new_[16178]_  = ~s1_rty_i | ~\new_[18823]_  | ~\new_[30124]_ ;
  assign \new_[16179]_  = \new_[18027]_  & \new_[29034]_ ;
  assign \new_[16180]_  = ~\new_[29767]_  & (~\new_[19301]_  | ~\new_[26261]_ );
  assign \new_[16181]_  = ~\new_[18290]_  | ~\new_[22980]_ ;
  assign \new_[16182]_  = ~s0_err_i | ~\new_[18192]_  | ~\new_[29434]_ ;
  assign \new_[16183]_  = ~\new_[29708]_  | ~\new_[18784]_  | ~s6_ack_i;
  assign \new_[16184]_  = ~m7_stb_i | ~\new_[19606]_  | ~\new_[29949]_ ;
  assign \new_[16185]_  = ~s2_ack_i | ~\new_[19638]_  | ~\new_[29846]_ ;
  assign \new_[16186]_  = ~\new_[18316]_  | ~\new_[26085]_ ;
  assign \new_[16187]_  = ~s10_ack_i | ~\new_[19595]_  | ~\new_[29710]_ ;
  assign \new_[16188]_  = ~s6_ack_i | ~\new_[18206]_  | ~\new_[29939]_ ;
  assign \new_[16189]_  = ~s12_err_i | ~\new_[18197]_  | ~\new_[30298]_ ;
  assign \new_[16190]_  = ~m5_stb_i | ~\new_[19547]_  | ~\new_[30311]_ ;
  assign \new_[16191]_  = ~s1_err_i | ~\new_[19639]_  | ~\new_[30001]_ ;
  assign \new_[16192]_  = ~s2_err_i | ~\new_[19638]_  | ~\new_[29846]_ ;
  assign \new_[16193]_  = ~s1_rty_i | ~\new_[19639]_  | ~\new_[30001]_ ;
  assign \new_[16194]_  = ~s2_rty_i | ~\new_[19638]_  | ~\new_[29846]_ ;
  assign \new_[16195]_  = ~s10_rty_i | ~\new_[19595]_  | ~\new_[29710]_ ;
  assign \new_[16196]_  = ~s10_err_i | ~\new_[19595]_  | ~\new_[29710]_ ;
  assign \new_[16197]_  = ~\new_[29565]_  & (~\new_[19307]_  | ~\new_[24785]_ );
  assign \new_[16198]_  = ~\new_[18300]_  | ~\new_[23538]_ ;
  assign \new_[16199]_  = ~s14_ack_i | ~\new_[18174]_  | ~\new_[29976]_ ;
  assign \new_[16200]_  = ~s8_err_i | ~\new_[18125]_  | ~\new_[29428]_ ;
  assign \new_[16201]_  = ~s0_rty_i | ~\new_[18936]_  | ~\new_[29819]_ ;
  assign \new_[16202]_  = ~\new_[18309]_  | ~\new_[24354]_ ;
  assign \new_[16203]_  = ~m3_stb_i | ~\new_[18849]_  | ~\new_[32168]_ ;
  assign \new_[16204]_  = ~m3_stb_i | ~\new_[18197]_  | ~\new_[30298]_ ;
  assign \new_[16205]_  = ~\new_[30026]_  | ~\new_[18083]_  | ~m0_stb_i;
  assign \new_[16206]_  = ~m1_stb_i | ~\new_[19627]_  | ~\new_[29976]_ ;
  assign \new_[16207]_  = \new_[18152]_  | \new_[21242]_ ;
  assign \new_[16208]_  = ~m7_stb_i | ~\new_[18824]_  | ~\new_[30113]_ ;
  assign \new_[16209]_  = ~\new_[29625]_  | ~\new_[18010]_  | ~m0_stb_i;
  assign \new_[16210]_  = ~m3_stb_i | ~\new_[19638]_  | ~\new_[29846]_ ;
  assign \new_[16211]_  = ~s0_ack_i | ~\new_[18192]_  | ~\new_[29434]_ ;
  assign \new_[16212]_  = ~s3_err_i | ~\new_[19633]_  | ~\new_[30469]_ ;
  assign \new_[16213]_  = ~s14_err_i | ~\new_[19627]_  | ~\new_[29976]_ ;
  assign \new_[16214]_  = ~\new_[28899]_  & (~\new_[19291]_  | ~\new_[26337]_ );
  assign \new_[16215]_  = ~s1_ack_i | ~\new_[18823]_  | ~\new_[30124]_ ;
  assign \new_[16216]_  = ~s9_err_i | ~\new_[18177]_  | ~\new_[30354]_ ;
  assign \new_[16217]_  = ~s12_ack_i | ~\new_[19636]_  | ~\new_[30298]_ ;
  assign \new_[16218]_  = ~s14_rty_i | ~\new_[19627]_  | ~\new_[29976]_ ;
  assign \new_[16219]_  = ~s8_rty_i | ~\new_[18167]_  | ~\new_[29670]_ ;
  assign \new_[16220]_  = ~s0_rty_i | ~\new_[18192]_  | ~\new_[29434]_ ;
  assign \new_[16221]_  = ~\new_[28950]_  & (~\new_[19310]_  | ~\new_[26852]_ );
  assign \new_[16222]_  = ~s1_ack_i | ~\new_[18201]_  | ~\new_[30001]_ ;
  assign \new_[16223]_  = ~s8_rty_i | ~\new_[18846]_  | ~\new_[29428]_ ;
  assign \new_[16224]_  = ~\new_[29241]_  | ~\new_[18204]_  | ~s8_ack_i;
  assign \new_[16225]_  = \new_[18133]_  | \new_[21234]_ ;
  assign \new_[16226]_  = ~\new_[18313]_  | ~\new_[26400]_ ;
  assign \new_[16227]_  = ~\new_[23378]_  & (~\new_[19312]_  | ~\new_[24471]_ );
  assign \new_[16228]_  = ~\new_[23382]_  & (~\new_[19313]_  | ~\new_[26271]_ );
  assign \new_[16229]_  = ~\new_[23744]_  & (~\new_[19314]_  | ~\new_[23122]_ );
  assign \new_[16230]_  = ~\new_[23418]_  & (~\new_[19320]_  | ~\new_[23413]_ );
  assign \new_[16231]_  = ~\new_[24863]_  & (~\new_[19317]_  | ~\new_[27973]_ );
  assign \new_[16232]_  = ~\new_[30093]_  & (~\new_[21727]_  | ~\new_[18994]_ );
  assign \new_[16233]_  = ~\new_[21202]_  & (~\new_[19318]_  | ~\new_[26359]_ );
  assign \new_[16234]_  = ~\new_[26907]_  & (~\new_[19324]_  | ~\new_[26776]_ );
  assign \new_[16235]_  = ~\new_[20979]_  | (~\new_[19326]_  & ~\new_[30219]_ );
  assign \new_[16236]_  = ~\new_[23549]_  & (~\new_[19319]_  | ~\new_[23155]_ );
  assign \new_[16237]_  = ~\new_[20853]_  | (~\new_[19323]_  & ~\new_[30087]_ );
  assign \new_[16238]_  = ~\new_[22275]_  & (~\new_[19322]_  | ~\new_[21584]_ );
  assign \new_[16239]_  = ~\new_[22316]_  & (~\new_[19321]_  | ~\new_[26701]_ );
  assign \new_[16240]_  = ~\new_[20879]_  | (~\new_[19325]_  & ~\new_[30339]_ );
  assign \new_[16241]_  = ~\new_[20989]_  | (~\new_[19327]_  & ~\new_[30305]_ );
  assign \new_[16242]_  = ~\new_[25147]_  & (~\new_[19328]_  | ~\new_[27606]_ );
  assign \new_[16243]_  = ~\new_[24716]_  & (~\new_[19276]_  | ~\new_[23365]_ );
  assign \new_[16244]_  = ~\new_[25195]_  & (~\new_[19267]_  | ~\new_[22424]_ );
  assign \new_[16245]_  = ~\new_[25159]_  & (~\new_[19252]_  | ~\new_[22324]_ );
  assign \new_[16246]_  = ~\new_[25168]_  & (~\new_[19254]_  | ~\new_[24528]_ );
  assign \new_[16247]_  = ~\new_[25179]_  & (~\new_[19283]_  | ~\new_[22241]_ );
  assign \new_[16248]_  = ~\new_[25265]_  & (~\new_[19259]_  | ~\new_[22157]_ );
  assign \new_[16249]_  = ~\new_[21317]_  & (~\new_[19279]_  | ~\new_[21186]_ );
  assign \new_[16250]_  = ~\new_[25190]_  & (~\new_[19250]_  | ~\new_[22273]_ );
  assign \new_[16251]_  = ~\new_[25206]_  & (~\new_[19247]_  | ~\new_[22251]_ );
  assign \new_[16252]_  = ~\new_[20531]_  & (~\new_[19266]_  | ~\new_[21207]_ );
  assign \new_[16253]_  = ~\new_[21321]_  & (~\new_[19280]_  | ~\new_[21221]_ );
  assign \new_[16254]_  = ~\new_[25187]_  & (~\new_[19264]_  | ~\new_[22423]_ );
  assign \new_[16255]_  = ~\new_[21271]_  & (~\new_[19253]_  | ~\new_[21254]_ );
  assign \new_[16256]_  = ~\new_[21295]_  & (~\new_[19281]_  | ~\new_[21138]_ );
  assign \new_[16257]_  = ~\new_[29028]_  | ~\new_[17971]_  | ~\new_[24807]_ ;
  assign \new_[16258]_  = ~\new_[30229]_  | ~\new_[17973]_  | ~\new_[22341]_ ;
  assign \new_[16259]_  = ~\new_[30222]_  | ~\new_[17974]_  | ~\new_[23424]_ ;
  assign \new_[16260]_  = ~\new_[30525]_  | ~\new_[17978]_  | ~\new_[23080]_ ;
  assign \new_[16261]_  = ~\new_[29987]_  | ~\new_[17989]_  | ~\new_[23572]_ ;
  assign \new_[16262]_  = ~\new_[29421]_  | ~\new_[17986]_  | ~\new_[23787]_ ;
  assign \new_[16263]_  = ~\new_[29276]_  | ~\new_[17983]_  | ~\new_[23401]_ ;
  assign \new_[16264]_  = ~\new_[29869]_  | ~\new_[17982]_  | ~\new_[22333]_ ;
  assign \new_[16265]_  = ~\new_[29623]_  | ~\new_[17990]_  | ~\new_[23860]_ ;
  assign \new_[16266]_  = ~\new_[28836]_  | ~\new_[17976]_  | ~\new_[23657]_ ;
  assign \new_[16267]_  = ~\new_[29851]_  | ~\new_[17997]_  | ~\new_[22239]_ ;
  assign \new_[16268]_  = ~\new_[29151]_  | ~\new_[17998]_  | ~\new_[24737]_ ;
  assign \new_[16269]_  = ~\new_[28278]_  | ~\new_[17987]_  | ~\new_[23736]_ ;
  assign \new_[16270]_  = ~\new_[29808]_  | ~\new_[17993]_  | ~\new_[24955]_ ;
  assign \new_[16271]_  = ~\new_[18383]_  | ~\new_[26239]_ ;
  assign \new_[16272]_  = ~\new_[18382]_  | ~\new_[27561]_ ;
  assign \new_[16273]_  = ~\new_[18384]_  | ~\new_[27594]_ ;
  assign \new_[16274]_  = ~\new_[31996]_ ;
  assign \new_[16275]_  = ~\new_[17197]_ ;
  assign \new_[16276]_  = ~\new_[17198]_ ;
  assign \new_[16277]_  = ~\new_[17198]_ ;
  assign \new_[16278]_  = ~\new_[17198]_ ;
  assign \new_[16279]_  = ~\new_[17207]_ ;
  assign \new_[16280]_  = ~\new_[17207]_ ;
  assign \new_[16281]_  = ~\new_[28422]_  & (~\new_[19346]_  | ~\new_[28872]_ );
  assign \new_[16282]_  = ~\new_[28815]_  & (~\new_[19348]_  | ~\new_[30057]_ );
  assign \new_[16283]_  = ~\new_[26857]_  & (~\new_[19349]_  | ~\new_[28883]_ );
  assign \new_[16284]_  = ~\new_[17210]_ ;
  assign \new_[16285]_  = ~\new_[18785]_ ;
  assign \new_[16286]_  = ~\new_[17211]_ ;
  assign \new_[16287]_  = ~\new_[17212]_ ;
  assign \new_[16288]_  = ~\new_[17212]_ ;
  assign \new_[16289]_  = ~\new_[18041]_ ;
  assign \new_[16290]_  = ~\new_[17214]_ ;
  assign \new_[16291]_  = ~\new_[17217]_ ;
  assign \new_[16292]_  = ~\new_[17225]_ ;
  assign \new_[16293]_  = ~\new_[17226]_ ;
  assign \new_[16294]_  = ~\new_[28113]_  & (~\new_[19371]_  | ~\new_[30030]_ );
  assign \new_[16295]_  = \new_[17231]_ ;
  assign \new_[16296]_  = ~\new_[17237]_ ;
  assign \new_[16297]_  = ~\new_[17238]_ ;
  assign \new_[16298]_  = ~\new_[27959]_  & (~\new_[19370]_  | ~\new_[28887]_ );
  assign \new_[16299]_  = ~\new_[28797]_  & (~\new_[19367]_  | ~\new_[29248]_ );
  assign \new_[16300]_  = ~\new_[26824]_  & (~\new_[19369]_  | ~\new_[29268]_ );
  assign \new_[16301]_  = ~\new_[17253]_ ;
  assign \new_[16302]_  = \new_[17253]_ ;
  assign \new_[16303]_  = ~\new_[17255]_ ;
  assign \new_[16304]_  = ~\new_[17255]_ ;
  assign \new_[16305]_  = ~\new_[19610]_ ;
  assign \new_[16306]_  = ~\new_[18148]_ ;
  assign \new_[16307]_  = ~\new_[17269]_ ;
  assign \new_[16308]_  = ~\new_[17269]_ ;
  assign \new_[16309]_  = ~\new_[18158]_ ;
  assign \new_[16310]_  = ~\new_[20359]_  & (~\new_[18730]_  | ~\new_[29357]_ );
  assign \new_[16311]_  = ~\new_[26788]_  & (~\new_[19342]_  | ~\new_[28939]_ );
  assign \new_[16312]_  = ~\new_[18942]_ ;
  assign \new_[16313]_  = ~\new_[28361]_  & (~\new_[19368]_  | ~\new_[28924]_ );
  assign \new_[16314]_  = \new_[18998]_  ? \new_[30649]_  : \new_[6049]_ ;
  assign \new_[16315]_  = ~\new_[25014]_  & (~\new_[19400]_  | ~\new_[21300]_ );
  assign \new_[16316]_  = ~\new_[17311]_ ;
  assign \new_[16317]_  = \new_[6214]_  ? \new_[29781]_  : \new_[19020]_ ;
  assign \new_[16318]_  = ~\new_[23145]_  | ~\new_[17825]_ ;
  assign \new_[16319]_  = (~\m4_data_i[28]  | ~\new_[19614]_ ) & (~\m3_data_i[28]  | ~\new_[18866]_ );
  assign \new_[16320]_  = ~\new_[22275]_  & (~\new_[19401]_  | ~\new_[21297]_ );
  assign \new_[16321]_  = ~\new_[17327]_ ;
  assign \new_[16322]_  = \new_[17327]_ ;
  assign \new_[16323]_  = ~\new_[20328]_  | ~\new_[23016]_  | ~\new_[26395]_  | ~\new_[28675]_ ;
  assign \new_[16324]_  = ~\new_[23720]_  & (~\new_[19402]_  | ~\new_[21311]_ );
  assign \new_[16325]_  = ~\new_[20325]_  | ~\new_[24255]_  | ~\new_[27691]_  | ~\new_[30297]_ ;
  assign \new_[16326]_  = ~\new_[17342]_ ;
  assign \new_[16327]_  = \new_[18970]_  ? \new_[30521]_  : \new_[6093]_ ;
  assign \new_[16328]_  = ~\new_[26284]_  | ~\new_[17833]_ ;
  assign \new_[16329]_  = ~\new_[20363]_  & (~\new_[18845]_  | ~\new_[29744]_ );
  assign \new_[16330]_  = ~\new_[18366]_  | ~\new_[29979]_ ;
  assign \new_[16331]_  = \new_[18960]_  ? \new_[30581]_  : \new_[31400]_ ;
  assign \new_[16332]_  = ~\new_[24673]_  | ~\new_[17673]_ ;
  assign \new_[16333]_  = (~\m4_data_i[30]  | ~\new_[19614]_ ) & (~\m3_data_i[30]  | ~\new_[18866]_ );
  assign \new_[16334]_  = \new_[19072]_  ? \new_[30642]_  : \new_[31499]_ ;
  assign \new_[16335]_  = ~\new_[18400]_  & (~\new_[18848]_  | ~\new_[30363]_ );
  assign \new_[16336]_  = ~\new_[19373]_  | ~\new_[18402]_ ;
  assign \new_[16337]_  = ~\new_[24748]_  | ~\new_[17809]_ ;
  assign \new_[16338]_  = ~\new_[17368]_ ;
  assign \new_[16339]_  = ~\new_[17369]_ ;
  assign \new_[16340]_  = ~\new_[18397]_  | ~\new_[30297]_ ;
  assign \new_[16341]_  = \new_[6273]_  ? \new_[30048]_  : \new_[19029]_ ;
  assign n8804 = m5_s0_cyc_o_reg;
  assign \new_[16343]_  = (~\m2_data_i[30]  | ~\new_[19571]_ ) & (~\m1_data_i[30]  | ~\new_[19629]_ );
  assign \new_[16344]_  = (~\m2_data_i[28]  | ~\new_[19571]_ ) & (~\m1_data_i[28]  | ~\new_[19629]_ );
  assign \new_[16345]_  = (~\m2_data_i[27]  | ~\new_[19571]_ ) & (~\m1_data_i[27]  | ~\new_[19630]_ );
  assign \new_[16346]_  = (~\m2_data_i[26]  | ~\new_[19571]_ ) & (~\m1_data_i[26]  | ~\new_[19629]_ );
  assign \new_[16347]_  = ~\new_[30063]_  & (~\new_[21721]_  | ~\new_[19037]_ );
  assign \new_[16348]_  = (~\m2_data_i[15]  | ~\new_[19571]_ ) & (~\m1_data_i[15]  | ~\new_[19630]_ );
  assign \new_[16349]_  = ~\new_[5917]_  | ~\new_[28248]_  | ~\new_[29227]_ ;
  assign \new_[16350]_  = ~\new_[5909]_  | ~\new_[26534]_  | ~\new_[29195]_ ;
  assign \new_[16351]_  = (~\m2_data_i[12]  | ~\new_[19571]_ ) & (~\m1_data_i[12]  | ~\new_[20575]_ );
  assign \new_[16352]_  = ~\new_[5923]_  | ~\new_[26530]_  | ~\new_[29068]_ ;
  assign \new_[16353]_  = ~\new_[5911]_  | ~\new_[26554]_  | ~\new_[29394]_ ;
  assign \new_[16354]_  = ~\new_[5918]_  | ~\new_[26496]_  | ~\new_[29578]_ ;
  assign \new_[16355]_  = ~\new_[5914]_  | ~\new_[28244]_  | ~\new_[29465]_ ;
  assign \new_[16356]_  = ~\new_[5912]_  | ~\new_[26446]_  | ~\new_[28833]_ ;
  assign \new_[16357]_  = ~\new_[24989]_  & (~\new_[19162]_  | ~\new_[29888]_ );
  assign \new_[16358]_  = ~\new_[5927]_  | ~\new_[24693]_  | ~\new_[29056]_ ;
  assign \new_[16359]_  = (~\m2_data_i[4]  | ~\new_[19571]_ ) & (~\m1_data_i[4]  | ~\new_[20575]_ );
  assign \new_[16360]_  = ~\new_[5921]_  | ~\new_[24585]_  | ~\new_[29663]_ ;
  assign \new_[16361]_  = (~\m2_data_i[3]  | ~\new_[19571]_ ) & (~\m1_data_i[3]  | ~\new_[19630]_ );
  assign \new_[16362]_  = (~\m2_data_i[0]  | ~\new_[19571]_ ) & (~\m1_data_i[0]  | ~\new_[19630]_ );
  assign \new_[16363]_  = (~\new_[19571]_  | ~\m2_addr_i[31] ) & (~\new_[19629]_  | ~\new_[31447]_ );
  assign \new_[16364]_  = ~\new_[30423]_  & (~\new_[21933]_  | ~\new_[19032]_ );
  assign \new_[16365]_  = (~\new_[19571]_  | ~\new_[31486]_ ) & (~\new_[19630]_  | ~\new_[31308]_ );
  assign \new_[16366]_  = (~\new_[19571]_  | ~\new_[31547]_ ) & (~\new_[19629]_  | ~\new_[31458]_ );
  assign \new_[16367]_  = (~\new_[19571]_  | ~\m2_addr_i[26] ) & (~\new_[18907]_  | ~\m1_addr_i[26] );
  assign \new_[16368]_  = (~\new_[19571]_  | ~\m2_addr_i[24] ) & (~\new_[19629]_  | ~\m1_addr_i[24] );
  assign \new_[16369]_  = (~\m2_addr_i[23]  | ~\new_[19571]_ ) & (~\m1_addr_i[23]  | ~\new_[19630]_ );
  assign \new_[16370]_  = (~\m2_addr_i[19]  | ~\new_[19571]_ ) & (~\m1_addr_i[19]  | ~\new_[19629]_ );
  assign \new_[16371]_  = ~\new_[24964]_  & (~\new_[19140]_  | ~\new_[30092]_ );
  assign \new_[16372]_  = ~\new_[18441]_  | ~\new_[27544]_ ;
  assign \new_[16373]_  = ~\new_[22857]_  & (~\new_[18509]_  | ~\new_[29550]_ );
  assign \new_[16374]_  = ~\new_[24305]_  & (~\new_[18522]_  | ~\new_[29003]_ );
  assign \new_[16375]_  = ~\new_[24260]_  & (~\new_[18533]_  | ~\new_[29192]_ );
  assign \new_[16376]_  = ~\new_[21611]_  & (~\new_[18535]_  | ~\new_[30000]_ );
  assign \new_[16377]_  = ~\new_[22919]_  & (~\new_[18544]_  | ~\new_[30446]_ );
  assign \new_[16378]_  = ~\new_[28266]_  | ~\new_[26375]_  | ~\new_[18559]_ ;
  assign \new_[16379]_  = ~\new_[24868]_  & (~\new_[18567]_  | ~\new_[28806]_ );
  assign \new_[16380]_  = (~\m2_addr_i[4]  | ~\new_[19571]_ ) & (~\m1_addr_i[4]  | ~\new_[20575]_ );
  assign \new_[16381]_  = (~\m2_addr_i[1]  | ~\new_[19571]_ ) & (~\m1_addr_i[1]  | ~\new_[20575]_ );
  assign \new_[16382]_  = ~\new_[30254]_  & (~\new_[21779]_  | ~\new_[19019]_ );
  assign \new_[16383]_  = ~\new_[23182]_  & (~\new_[18593]_  | ~\new_[30554]_ );
  assign \new_[16384]_  = (~\m2_sel_i[3]  | ~\new_[19571]_ ) & (~\m1_sel_i[3]  | ~\new_[20575]_ );
  assign \new_[16385]_  = ~\new_[22882]_  & (~\new_[18556]_  | ~\new_[30842]_ );
  assign \new_[16386]_  = ~\new_[22896]_  & (~\new_[18611]_  | ~\new_[29787]_ );
  assign \new_[16387]_  = ~\new_[23037]_  & (~\new_[18600]_  | ~\new_[28337]_ );
  assign \new_[16388]_  = (~\m2_sel_i[0]  | ~\new_[19571]_ ) & (~\m1_sel_i[0]  | ~\new_[18907]_ );
  assign \new_[16389]_  = ~\new_[18459]_  | ~\new_[24330]_ ;
  assign \new_[16390]_  = ~\new_[22981]_  & (~\new_[18624]_  | ~\new_[30205]_ );
  assign \new_[16391]_  = ~\new_[22848]_  & (~\new_[18636]_  | ~\new_[29455]_ );
  assign \new_[16392]_  = \new_[19022]_  ? \new_[30703]_  : \new_[6211]_ ;
  assign \new_[16393]_  = ~\new_[25116]_  & (~\new_[18507]_  | ~\new_[30283]_ );
  assign \new_[16394]_  = ~\new_[22857]_  & (~\new_[18510]_  | ~\new_[23146]_ );
  assign \new_[16395]_  = ~\new_[26224]_  & (~\new_[18512]_  | ~\new_[24283]_ );
  assign \new_[16396]_  = ~\new_[23058]_  & (~\new_[18513]_  | ~\new_[27264]_ );
  assign \new_[16397]_  = \new_[17583]_  | \new_[24998]_ ;
  assign \new_[16398]_  = \new_[17584]_  | \new_[27572]_ ;
  assign \new_[16399]_  = \new_[17585]_  | \new_[27615]_ ;
  assign \new_[16400]_  = ~\new_[24324]_  & (~\new_[18547]_  | ~\new_[23937]_ );
  assign \new_[16401]_  = \new_[17586]_  | \new_[26409]_ ;
  assign \new_[16402]_  = ~\new_[24862]_  & (~\new_[18551]_  | ~\new_[30037]_ );
  assign \new_[16403]_  = ~\new_[24868]_  & (~\new_[18568]_  | ~\new_[26252]_ );
  assign \new_[16404]_  = ~\new_[24937]_  & (~\new_[18536]_  | ~\new_[29870]_ );
  assign \new_[16405]_  = ~\new_[18452]_  & ~\new_[24976]_ ;
  assign \new_[16406]_  = \new_[17590]_  | \new_[24854]_ ;
  assign \new_[16407]_  = ~\new_[26930]_  & (~\new_[18586]_  | ~\new_[30645]_ );
  assign \new_[16408]_  = ~\new_[24563]_  & (~\new_[18589]_  | ~\new_[24443]_ );
  assign \new_[16409]_  = \new_[17588]_  | \new_[27965]_ ;
  assign \new_[16410]_  = ~\new_[25026]_  & (~\new_[18584]_  | ~\new_[29802]_ );
  assign \new_[16411]_  = ~\new_[23273]_  & (~\new_[18594]_  | ~\new_[24475]_ );
  assign \new_[16412]_  = ~\new_[22882]_  & (~\new_[18527]_  | ~\new_[27360]_ );
  assign \new_[16413]_  = \new_[17587]_  | \new_[26426]_ ;
  assign \new_[16414]_  = ~\new_[23066]_  & (~\new_[18602]_  | ~\new_[24417]_ );
  assign \new_[16415]_  = ~\new_[26998]_  & (~\new_[18605]_  | ~\new_[29813]_ );
  assign \new_[16416]_  = ~\new_[26380]_  & (~\new_[18623]_  | ~\new_[26390]_ );
  assign \new_[16417]_  = ~\new_[22981]_  & (~\new_[18622]_  | ~\new_[28253]_ );
  assign \new_[16418]_  = \new_[17589]_  | \new_[27677]_ ;
  assign \new_[16419]_  = ~\new_[28817]_  | ~\new_[17761]_ ;
  assign \new_[16420]_  = ~\new_[26960]_  & (~\new_[18618]_  | ~\new_[30352]_ );
  assign \new_[16421]_  = ~\new_[20489]_  & (~\new_[18616]_  | ~\new_[27584]_ );
  assign \new_[16422]_  = ~\new_[25137]_  & (~\new_[18633]_  | ~\new_[30262]_ );
  assign \new_[16423]_  = ~\new_[24929]_  & (~\new_[18638]_  | ~\new_[24458]_ );
  assign \new_[16424]_  = ~\new_[21545]_  & (~\new_[18639]_  | ~\new_[26807]_ );
  assign \new_[16425]_  = \new_[17591]_  | \new_[24780]_ ;
  assign \new_[16426]_  = ~\new_[22409]_  & (~\new_[18621]_  | ~\new_[28114]_ );
  assign \new_[16427]_  = ~\new_[26905]_  | ~\new_[26811]_  | ~\new_[18486]_ ;
  assign \new_[16428]_  = ~\new_[23015]_  & (~\new_[18520]_  | ~\new_[29969]_ );
  assign \new_[16429]_  = ~\new_[27824]_  & (~\new_[18521]_  | ~\new_[28894]_ );
  assign \new_[16430]_  = ~\new_[27692]_  & (~\new_[18525]_  | ~\new_[29435]_ );
  assign \new_[16431]_  = ~\new_[26251]_  | ~\new_[28134]_  | ~\new_[18487]_ ;
  assign \new_[16432]_  = ~\new_[28130]_  & (~\new_[18534]_  | ~\new_[30222]_ );
  assign \new_[16433]_  = ~\new_[26246]_  | ~\new_[27973]_  | ~\new_[18488]_ ;
  assign \new_[16434]_  = ~\new_[21509]_  | ~\new_[26213]_  | ~\new_[18519]_ ;
  assign \new_[16435]_  = ~\new_[29430]_  & (~\new_[18543]_  | ~\new_[30525]_ );
  assign \new_[16436]_  = ~\new_[26223]_  | ~\new_[26776]_  | ~\new_[18489]_ ;
  assign \new_[16437]_  = ~\new_[24351]_  & (~\new_[18554]_  | ~\new_[30022]_ );
  assign \new_[16438]_  = ~\new_[23187]_  | ~\new_[24632]_  | ~\new_[18562]_ ;
  assign \new_[16439]_  = ~\new_[23183]_  & (~\new_[18565]_  | ~\new_[30552]_ );
  assign \new_[16440]_  = ~\new_[26270]_  & (~\new_[18566]_  | ~\new_[30467]_ );
  assign \new_[16441]_  = ~\new_[26260]_  | ~\new_[27914]_  | ~\new_[18492]_ ;
  assign \new_[16442]_  = ~\new_[26685]_  & (~\new_[18574]_  | ~\new_[28818]_ );
  assign \new_[16443]_  = ~\new_[24427]_  & (~\new_[18576]_  | ~\new_[30628]_ );
  assign \new_[16444]_  = ~\new_[18464]_  | ~\new_[22888]_ ;
  assign \new_[16445]_  = ~\new_[18463]_  & (~\new_[30254]_  | ~\new_[6061]_ );
  assign \new_[16446]_  = ~\new_[24365]_  | ~\new_[27901]_  | ~\new_[18585]_ ;
  assign \new_[16447]_  = ~\new_[28485]_  & (~\new_[18537]_  | ~\new_[30599]_ );
  assign \new_[16448]_  = ~\new_[26835]_  | ~\new_[26283]_  | ~\new_[18493]_ ;
  assign \new_[16449]_  = ~\new_[29558]_  & (~\new_[18590]_  | ~\new_[29869]_ );
  assign \new_[16450]_  = ~\new_[24613]_  | ~\new_[27846]_  | ~\new_[18494]_ ;
  assign \new_[16451]_  = ~\new_[23273]_  & (~\new_[18563]_  | ~\new_[30491]_ );
  assign \new_[16452]_  = ~\new_[27772]_  | ~\new_[27425]_  | ~\new_[18496]_ ;
  assign \new_[16453]_  = ~\new_[21468]_  & (~\new_[18596]_  | ~\new_[28023]_ );
  assign \new_[16454]_  = ~\new_[28563]_  & (~\new_[18597]_  | ~\new_[28278]_ );
  assign \new_[16455]_  = ~\new_[23066]_  & (~\new_[18603]_  | ~\new_[28935]_ );
  assign \new_[16456]_  = ~\new_[25505]_  | ~\new_[23096]_  | ~\new_[18498]_ ;
  assign \new_[16457]_  = \new_[6082]_  ? \new_[30579]_  : \new_[19105]_ ;
  assign \new_[16458]_  = ~\new_[28484]_  & (~\new_[18607]_  | ~\new_[30248]_ );
  assign \new_[16459]_  = ~\new_[26311]_  & (~\new_[18634]_  | ~\new_[30297]_ );
  assign \new_[16460]_  = ~\new_[27653]_  & (~\new_[18615]_  | ~\new_[30544]_ );
  assign \new_[16461]_  = ~\new_[22851]_  & (~\new_[18635]_  | ~\new_[28355]_ );
  assign \new_[16462]_  = ~\new_[22873]_  | (~\new_[18502]_  & ~\new_[29853]_ );
  assign \new_[16463]_  = ~\new_[27733]_  & (~\new_[18691]_  | ~\new_[30320]_ );
  assign \new_[16464]_  = ~\new_[26541]_  & (~\new_[18692]_  | ~\new_[29746]_ );
  assign \new_[16465]_  = ~\new_[24317]_  | (~\new_[18549]_  & ~\new_[29935]_ );
  assign \new_[16466]_  = ~\new_[27625]_  & (~\new_[18693]_  | ~\new_[30011]_ );
  assign \new_[16467]_  = ~\new_[22865]_  | (~\new_[18572]_  & ~\new_[30070]_ );
  assign \new_[16468]_  = ~\new_[28612]_  & (~\new_[18694]_  | ~\new_[30717]_ );
  assign \new_[16469]_  = ~\new_[21560]_  | (~\new_[18581]_  & ~\new_[30526]_ );
  assign \new_[16470]_  = ~\new_[24861]_  & (~\new_[18695]_  | ~\new_[28888]_ );
  assign \new_[16471]_  = ~\new_[28417]_  & (~\new_[18696]_  | ~\new_[30572]_ );
  assign \new_[16472]_  = ~\new_[27665]_  & (~\new_[18697]_  | ~\new_[29863]_ );
  assign \new_[16473]_  = ~\new_[24322]_  & (~\new_[18698]_  | ~\new_[28762]_ );
  assign \new_[16474]_  = ~\new_[25213]_  & (~\new_[18699]_  | ~\new_[28964]_ );
  assign \new_[16475]_  = \new_[6195]_  ? \new_[29332]_  : \new_[19016]_ ;
  assign \new_[16476]_  = ~\new_[23124]_  | (~\new_[18631]_  & ~\new_[30003]_ );
  assign \new_[16477]_  = ~\new_[27543]_  & (~\new_[18700]_  | ~\new_[29798]_ );
  assign \new_[16478]_  = ~\new_[29861]_  & (~\new_[18500]_  | ~\new_[29357]_ );
  assign \new_[16479]_  = ~\new_[29841]_  & (~\new_[18515]_  | ~\new_[30030]_ );
  assign \new_[16480]_  = ~\new_[30415]_  & (~\new_[18528]_  | ~\new_[28872]_ );
  assign \new_[16481]_  = ~\new_[30202]_  & (~\new_[18538]_  | ~\new_[30057]_ );
  assign \new_[16482]_  = ~\new_[29931]_  & (~\new_[18546]_  | ~\new_[28883]_ );
  assign \new_[16483]_  = ~\new_[29902]_  & (~\new_[18504]_  | ~\new_[29104]_ );
  assign \new_[16484]_  = ~\new_[29445]_  & (~\new_[18625]_  | ~\new_[28962]_ );
  assign \new_[16485]_  = ~\new_[29174]_  & (~\new_[18579]_  | ~\new_[29202]_ );
  assign \new_[16486]_  = ~\new_[30053]_  & (~\new_[18587]_  | ~\new_[28939]_ );
  assign \new_[16487]_  = ~\new_[30212]_  & (~\new_[18511]_  | ~\new_[28887]_ );
  assign \new_[16488]_  = ~\new_[30058]_  & (~\new_[18517]_  | ~\new_[29248]_ );
  assign \new_[16489]_  = ~\new_[30114]_  & (~\new_[18523]_  | ~\new_[28924]_ );
  assign \new_[16490]_  = ~\new_[30140]_  & (~\new_[18575]_  | ~\new_[29268]_ );
  assign \new_[16491]_  = ~\new_[29629]_  & (~\new_[18614]_  | ~\new_[29744]_ );
  assign \new_[16492]_  = ~\new_[29564]_  & (~\new_[18627]_  | ~\new_[29350]_ );
  assign \new_[16493]_  = (~\new_[18503]_  | ~\new_[29794]_ ) & (~\new_[30612]_  | ~\new_[6033]_ );
  assign \new_[16494]_  = (~\new_[18505]_  | ~\new_[30283]_ ) & (~\new_[30566]_  | ~\new_[6033]_ );
  assign \new_[16495]_  = (~\new_[18550]_  | ~\new_[30037]_ ) & (~\new_[30616]_  | ~\new_[31712]_ );
  assign \new_[16496]_  = (~\new_[18620]_  | ~\new_[29870]_ ) & (~\new_[30688]_  | ~\new_[30884]_ );
  assign \new_[16497]_  = (~\new_[18582]_  | ~\new_[29877]_ ) & (~\new_[30478]_  | ~\new_[30897]_ );
  assign \new_[16498]_  = (~\new_[18583]_  | ~\new_[30645]_ ) & (~\new_[30028]_  | ~\new_[30897]_ );
  assign \new_[16499]_  = (~\new_[18632]_  | ~\new_[30262]_ ) & (~\new_[30607]_  | ~\new_[31045]_ );
  assign \new_[16500]_  = ~\new_[28162]_  & (~\new_[18701]_  | ~\new_[28114]_ );
  assign \new_[16501]_  = ~\new_[28495]_  & (~\new_[18702]_  | ~\new_[28069]_ );
  assign \new_[16502]_  = ~\new_[26597]_  & (~\new_[18704]_  | ~\new_[27787]_ );
  assign \new_[16503]_  = ~\new_[27601]_  & (~\new_[18705]_  | ~\new_[26655]_ );
  assign \new_[16504]_  = ~\new_[26394]_  & (~\new_[18706]_  | ~\new_[29064]_ );
  assign \new_[16505]_  = ~\new_[27991]_  & (~\new_[18703]_  | ~\new_[30491]_ );
  assign \new_[16506]_  = ~\new_[27628]_  & (~\new_[18707]_  | ~\new_[28023]_ );
  assign \new_[16507]_  = ~\new_[28233]_  & (~\new_[18708]_  | ~\new_[29537]_ );
  assign \new_[16508]_  = ~\new_[28229]_  & (~\new_[18709]_  | ~\new_[30735]_ );
  assign \new_[16509]_  = ~\new_[18432]_  | (~\new_[29794]_  & ~\new_[6034]_ );
  assign \new_[16510]_  = ~\new_[24266]_  & (~\new_[18484]_  | ~\new_[30221]_ );
  assign \new_[16511]_  = ~\new_[19500]_  | ~\new_[28042]_  | ~\new_[30730]_  | ~\new_[28069]_ ;
  assign \new_[16512]_  = ~\new_[26365]_  & (~\new_[18485]_  | ~\new_[30730]_ );
  assign \new_[16513]_  = ~\new_[19501]_  | ~\new_[28192]_  | ~\new_[30135]_  | ~\new_[29435]_ ;
  assign \new_[16514]_  = ~\new_[19502]_  | ~\new_[29642]_  | ~\new_[30139]_  | ~\new_[27787]_ ;
  assign \new_[16515]_  = ~\new_[24328]_  | (~\new_[18541]_  & ~\new_[30336]_ );
  assign \new_[16516]_  = ~\new_[18433]_  | (~\new_[30160]_  & ~\new_[6050]_ );
  assign \new_[16517]_  = ~\new_[18434]_  | (~\new_[30146]_  & ~\new_[31422]_ );
  assign \new_[16518]_  = (~\new_[19614]_  | ~\m4_addr_i[24] ) & (~\new_[18863]_  | ~\m3_addr_i[24] );
  assign \new_[16519]_  = ~\new_[18435]_  | (~\new_[30349]_  & ~\new_[6057]_ );
  assign \new_[16520]_  = ~\new_[18436]_  | (~\new_[29877]_  & ~\new_[6061]_ );
  assign \new_[16521]_  = ~\new_[20356]_  & (~\new_[18812]_  | ~\new_[28962]_ );
  assign \new_[16522]_  = ~\new_[18437]_  | (~\new_[30071]_  & ~\new_[6070]_ );
  assign \new_[16523]_  = ~\new_[23028]_  & (~\new_[18495]_  | ~\new_[29892]_ );
  assign \new_[16524]_  = \new_[19092]_  ? \new_[30677]_  : \new_[6079]_ ;
  assign \new_[16525]_  = ~\new_[18438]_  | (~\new_[30278]_  & ~\new_[6270]_ );
  assign \new_[16526]_  = ~\new_[23012]_  & (~\new_[18497]_  | ~\new_[29913]_ );
  assign \new_[16527]_  = ~\new_[18439]_  | (~\new_[30218]_  & ~\new_[6215]_ );
  assign \new_[16528]_  = \new_[19075]_  ? \new_[30568]_  : \new_[6197]_ ;
  assign \new_[16529]_  = ~\new_[18440]_  | (~\new_[29897]_  & ~\new_[6092]_ );
  assign \new_[16530]_  = ~\new_[19503]_  | ~\new_[28760]_  | ~\new_[30724]_  | ~\new_[30735]_ ;
  assign \new_[16531]_  = ~\new_[26268]_  & (~\new_[18499]_  | ~\new_[30724]_ );
  assign \new_[16532]_  = \new_[18262]_  & \new_[6274]_ ;
  assign \new_[16533]_  = ~\new_[19361]_  & (~\new_[18802]_  | ~\new_[29104]_ );
  assign \new_[16534]_  = \new_[6038]_  ? \new_[29079]_  : \new_[18671]_ ;
  assign \new_[16535]_  = \new_[6176]_  ? \new_[30232]_  : \new_[18672]_ ;
  assign \new_[16536]_  = \new_[5968]_  ? \new_[28866]_  : \new_[18675]_ ;
  assign \new_[16537]_  = \new_[30511]_  ? \new_[30665]_  : \new_[18676]_ ;
  assign \new_[16538]_  = (~\new_[18673]_  | ~\new_[30207]_ ) & (~\new_[30701]_  | ~\new_[31491]_ );
  assign \new_[16539]_  = \new_[6212]_  ? \new_[30595]_  : \new_[18681]_ ;
  assign \new_[16540]_  = \new_[6071]_  ? \new_[29892]_  : \new_[18680]_ ;
  assign \new_[16541]_  = \new_[6269]_  ? \new_[29913]_  : \new_[18687]_ ;
  assign \new_[16542]_  = \new_[6269]_  ? \new_[29210]_  : \new_[18686]_ ;
  assign \new_[16543]_  = \new_[5930]_  ? \new_[30437]_  : \new_[18685]_ ;
  assign \new_[16544]_  = \new_[5932]_  ? \new_[28371]_  : \new_[18690]_ ;
  assign \new_[16545]_  = ~\new_[17795]_  | ~\new_[30343]_ ;
  assign \new_[16546]_  = ~\new_[29119]_  & (~\new_[18729]_  | ~\new_[28049]_ );
  assign \new_[16547]_  = ~\new_[17858]_  & ~\new_[23160]_ ;
  assign \new_[16548]_  = ~\new_[17656]_  | ~\new_[30152]_ ;
  assign \new_[16549]_  = ~\new_[17859]_  & ~\new_[27540]_ ;
  assign \new_[16550]_  = ~\new_[29874]_  | (~\new_[20121]_  & ~\new_[18965]_ );
  assign \new_[16551]_  = ~\new_[29855]_  & (~\new_[18869]_  | ~\new_[28412]_ );
  assign \new_[16552]_  = ~\new_[17665]_  | ~\new_[28183]_ ;
  assign \new_[16553]_  = ~\new_[29100]_  & (~\new_[18773]_  | ~\new_[28222]_ );
  assign \new_[16554]_  = ~\new_[17676]_  | ~\new_[29746]_ ;
  assign \new_[16555]_  = ~\new_[30109]_  & (~\new_[18774]_  | ~\new_[26305]_ );
  assign \new_[16556]_  = ~\new_[17862]_  & ~\new_[22939]_ ;
  assign \new_[16557]_  = ~\new_[30389]_  & (~\new_[18779]_  | ~\new_[28500]_ );
  assign \new_[16558]_  = ~\new_[29032]_  | (~\new_[20000]_  & ~\new_[18969]_ );
  assign \new_[16559]_  = ~\new_[30564]_  & (~\new_[18783]_  | ~\new_[28275]_ );
  assign \new_[16560]_  = ~\new_[17863]_  & ~\new_[25488]_ ;
  assign \new_[16561]_  = ~\new_[29401]_  | (~\new_[20079]_  & ~\new_[18999]_ );
  assign \new_[16562]_  = ~\new_[28522]_  | ~\new_[29984]_  | ~\new_[19145]_ ;
  assign \new_[16563]_  = ~\new_[17724]_  | ~\new_[29104]_ ;
  assign \new_[16564]_  = ~\new_[30044]_  & (~\new_[21795]_  | ~\new_[19161]_ );
  assign \new_[16565]_  = ~\new_[29898]_  & (~\new_[18778]_  | ~\new_[28108]_ );
  assign \new_[16566]_  = ~\new_[29233]_  | (~\new_[20881]_  & ~\new_[19034]_ );
  assign \new_[16567]_  = ~\new_[30217]_  | (~\new_[19272]_  & ~\new_[19852]_ );
  assign \new_[16568]_  = ~\new_[28048]_  | ~\new_[29904]_  | ~\new_[19148]_ ;
  assign \new_[16569]_  = ~\new_[28982]_  & (~\new_[20990]_  | ~\new_[19149]_ );
  assign \new_[16570]_  = ~\new_[17741]_  | ~\new_[30717]_ ;
  assign \new_[16571]_  = ~\new_[30515]_  & (~\new_[18872]_  | ~\new_[27990]_ );
  assign \new_[16572]_  = ~\new_[17868]_  & ~\new_[24558]_ ;
  assign \new_[16573]_  = ~\new_[29959]_  & (~\new_[21750]_  | ~\new_[19003]_ );
  assign \new_[16574]_  = ~\new_[28559]_  | ~\new_[29404]_  | ~\new_[19154]_ ;
  assign \new_[16575]_  = ~\new_[29331]_  & (~\new_[20901]_  | ~\new_[19155]_ );
  assign \new_[16576]_  = ~\new_[17871]_  & ~\new_[26825]_ ;
  assign \new_[16577]_  = ~\new_[17812]_  | ~\new_[28888]_ ;
  assign \new_[16578]_  = ~\new_[30423]_  & (~\new_[18873]_  | ~\new_[24612]_ );
  assign \new_[16579]_  = ~\new_[17866]_  & ~\new_[23045]_ ;
  assign \new_[16580]_  = ~\new_[28501]_  | ~\new_[30016]_  | ~\new_[19127]_ ;
  assign \new_[16581]_  = ~\new_[26804]_  & (~\new_[18725]_  | ~\new_[29978]_ );
  assign \new_[16582]_  = ~\new_[17836]_  | ~\new_[30572]_ ;
  assign \new_[16583]_  = ~\new_[30063]_  & (~\new_[18839]_  | ~\new_[28178]_ );
  assign \new_[16584]_  = ~\new_[17876]_  & ~\new_[26431]_ ;
  assign \new_[16585]_  = ~\new_[28905]_  | (~\new_[20966]_  & ~\new_[19039]_ );
  assign \new_[16586]_  = ~\new_[29355]_  | (~\new_[20067]_  & ~\new_[19040]_ );
  assign \new_[16587]_  = ~\new_[29648]_  & (~\new_[18842]_  | ~\new_[28474]_ );
  assign \new_[16588]_  = ~\new_[17782]_  | ~\new_[29299]_ ;
  assign \new_[16589]_  = ~\new_[30784]_  | (~\new_[20894]_  & ~\new_[19046]_ );
  assign \new_[16590]_  = ~\new_[17726]_  | ~\new_[28762]_ ;
  assign \new_[16591]_  = ~\new_[28204]_  & (~\new_[18843]_  | ~\new_[26420]_ );
  assign \new_[16592]_  = ~\new_[17869]_  & ~\new_[24346]_ ;
  assign \new_[16593]_  = ~\new_[30610]_  | (~\new_[20087]_  & ~\new_[19051]_ );
  assign \new_[16594]_  = ~\new_[27559]_  & (~\new_[18726]_  | ~\new_[28188]_ );
  assign \new_[16595]_  = ~\new_[28950]_  & (~\new_[21962]_  | ~\new_[19185]_ );
  assign \new_[16596]_  = ~\new_[28950]_  & (~\new_[18938]_  | ~\new_[26812]_ );
  assign \new_[16597]_  = ~\new_[17889]_  & ~\new_[24644]_ ;
  assign \new_[16598]_  = ~\new_[30084]_  | (~\new_[21946]_  & ~\new_[19057]_ );
  assign \new_[16599]_  = ~\new_[23491]_  & (~\new_[19131]_  | ~\new_[29984]_ );
  assign \new_[16600]_  = ~\new_[17797]_  | ~\new_[28001]_ ;
  assign \new_[16601]_  = ~\new_[30147]_  | (~\new_[20974]_  & ~\new_[19065]_ );
  assign \new_[16602]_  = ~\new_[30707]_  | (~\new_[20797]_  & ~\new_[19068]_ );
  assign \new_[16603]_  = ~\new_[29096]_  & (~\new_[20746]_  | ~\new_[19143]_ );
  assign \new_[16604]_  = ~\new_[29560]_  | (~\new_[20115]_  & ~\new_[19070]_ );
  assign \new_[16605]_  = ~\new_[29040]_  | (~\new_[20122]_  & ~\new_[19073]_ );
  assign \new_[16606]_  = ~\new_[17822]_  | ~\new_[30786]_ ;
  assign \new_[16607]_  = ~\new_[28475]_  | ~\new_[29557]_  | ~\new_[19186]_ ;
  assign \new_[16608]_  = ~\new_[29166]_  & (~\new_[21557]_  | ~\new_[19187]_ );
  assign \new_[16609]_  = ~\new_[30708]_  & (~\new_[18771]_  | ~\new_[28128]_ );
  assign \new_[16610]_  = ~\new_[17892]_  & ~\new_[25573]_ ;
  assign \new_[16611]_  = ~\new_[30820]_  | (~\new_[21001]_  & ~\new_[19106]_ );
  assign \new_[16612]_  = ~\new_[29372]_  & (~\new_[18728]_  | ~\new_[29996]_ );
  assign \new_[16613]_  = ~\new_[28740]_  | ~\new_[29900]_  | ~\new_[19191]_ ;
  assign \new_[16614]_  = ~\new_[18514]_  & ~\new_[18227]_ ;
  assign \new_[16615]_  = ~\new_[17690]_  & ~\new_[29930]_ ;
  assign \new_[16616]_  = ~\new_[17701]_  & ~\new_[30093]_ ;
  assign \new_[16617]_  = ~\new_[17744]_  & ~\new_[30199]_ ;
  assign \new_[16618]_  = ~\new_[17768]_  & ~\new_[30010]_ ;
  assign \new_[16619]_  = ~\new_[17769]_  & ~\new_[30066]_ ;
  assign \new_[16620]_  = ~\new_[17654]_  & ~\new_[30075]_ ;
  assign \new_[16621]_  = ~\new_[17830]_  & ~\new_[30047]_ ;
  assign \new_[16622]_  = \new_[17841]_  | \new_[28687]_ ;
  assign \new_[16623]_  = ~\new_[17842]_  | ~\new_[26281]_ ;
  assign \new_[16624]_  = ~\new_[17843]_  | ~\new_[28275]_ ;
  assign \new_[16625]_  = \new_[17844]_  | \new_[28566]_ ;
  assign \new_[16626]_  = ~\new_[17845]_  | ~\new_[28508]_ ;
  assign \new_[16627]_  = \new_[17846]_  | \new_[26366]_ ;
  assign \new_[16628]_  = ~\new_[17847]_  | ~\new_[28538]_ ;
  assign \new_[16629]_  = ~\new_[17848]_  | ~\new_[27990]_ ;
  assign \new_[16630]_  = ~\new_[17851]_  | ~\new_[26768]_ ;
  assign \new_[16631]_  = ~\new_[17853]_  | ~\new_[28490]_ ;
  assign \new_[16632]_  = \new_[17849]_  | \new_[28978]_ ;
  assign \new_[16633]_  = ~\new_[17854]_  | ~\new_[24612]_ ;
  assign \new_[16634]_  = ~\new_[17850]_  | ~\new_[28178]_ ;
  assign \new_[16635]_  = ~\new_[17852]_  | ~\new_[26420]_ ;
  assign \new_[16636]_  = ~\new_[17855]_  | ~\new_[26790]_ ;
  assign \new_[16637]_  = ~\new_[17856]_  | ~\new_[28128]_ ;
  assign \new_[16638]_  = \new_[17857]_  | \new_[28454]_ ;
  assign \new_[16639]_  = ~\new_[30303]_  & (~\new_[23335]_  | ~\new_[19124]_ );
  assign \new_[16640]_  = ~\new_[18787]_  | ~\new_[31314]_  | ~n8584;
  assign \new_[16641]_  = ~\new_[29181]_  & (~\new_[20736]_  | ~\new_[19001]_ );
  assign \new_[16642]_  = \new_[17602]_  & \new_[30030]_ ;
  assign \new_[16643]_  = \new_[17607]_  & \new_[28872]_ ;
  assign \new_[16644]_  = ~\new_[18871]_  | ~\new_[30487]_  | ~n8319;
  assign \new_[16645]_  = ~\new_[18835]_  | ~\new_[31236]_  | ~n8419;
  assign \new_[16646]_  = \new_[17612]_  & \new_[30057]_ ;
  assign \new_[16647]_  = ~\new_[29689]_  & (~\new_[23622]_  | ~\new_[19138]_ );
  assign \new_[16648]_  = \new_[17616]_  & \new_[28883]_ ;
  assign \new_[16649]_  = ~\new_[28651]_  & (~\new_[21223]_  | ~\new_[19141]_ );
  assign \new_[16650]_  = ~\new_[18784]_  | ~\new_[31363]_  | ~n8669;
  assign \new_[16651]_  = ~\new_[18910]_  | ~\new_[31520]_  | ~n8879;
  assign \new_[16652]_  = ~\new_[18803]_  | ~\new_[31472]_  | ~n8834;
  assign \new_[16653]_  = ~\new_[18831]_  | ~\new_[31286]_  | ~n8524;
  assign \new_[16654]_  = ~\new_[18881]_  | ~\new_[30484]_  | ~n8304;
  assign \new_[16655]_  = ~\new_[18742]_  | ~\new_[30792]_  | ~n8364;
  assign \new_[16656]_  = ~\new_[28775]_  & (~\new_[24951]_  | ~\new_[19156]_ );
  assign \new_[16657]_  = ~\new_[18790]_  | ~\new_[31307]_  | ~n8574;
  assign \new_[16658]_  = ~\new_[17276]_  | ~\new_[31223]_  | ~n8394;
  assign \new_[16659]_  = ~\new_[18882]_  | ~\new_[31528]_  | ~n8914;
  assign \new_[16660]_  = \new_[17621]_  & \new_[28962]_ ;
  assign \new_[16661]_  = ~\new_[28303]_  & (~\new_[23785]_  | ~\new_[19181]_ );
  assign \new_[16662]_  = \new_[17627]_  & \new_[29202]_ ;
  assign \new_[16663]_  = ~\new_[29986]_  & (~\new_[22292]_  | ~\new_[19157]_ );
  assign \new_[16664]_  = ~\new_[18846]_  | ~\new_[31530]_  | ~n8919;
  assign \new_[16665]_  = ~\new_[18878]_  | ~\new_[31515]_  | ~n8859;
  assign \new_[16666]_  = ~\new_[18760]_  | ~\new_[30793]_  | ~n8369;
  assign \new_[16667]_  = ~\new_[29060]_  & (~\new_[23707]_  | ~\new_[19160]_ );
  assign \new_[16668]_  = \new_[17631]_  & \new_[28939]_ ;
  assign \new_[16669]_  = ~\new_[28043]_  & (~\new_[23764]_  | ~\new_[19182]_ );
  assign \new_[16670]_  = \new_[17635]_  & \new_[28887]_ ;
  assign \new_[16671]_  = ~\new_[18806]_  | ~\new_[31336]_  | ~n8614;
  assign \new_[16672]_  = ~\new_[18850]_  | ~\new_[31313]_  | ~n8579;
  assign \new_[16673]_  = ~\new_[18906]_  | ~\new_[31349]_  | ~n8634;
  assign \new_[16674]_  = \new_[17652]_  & \new_[29248]_ ;
  assign \new_[16675]_  = \new_[17639]_  & \new_[28924]_ ;
  assign \new_[16676]_  = \new_[17649]_  & \new_[30363]_ ;
  assign \new_[16677]_  = ~\new_[18879]_  | ~\new_[31238]_  | ~n8429;
  assign \new_[16678]_  = ~\new_[18821]_  | ~\new_[31330]_  | ~n8604;
  assign \new_[16679]_  = ~\new_[18822]_  | ~\new_[31534]_  | ~n8934;
  assign \new_[16680]_  = ~\new_[18929]_  | ~\new_[31296]_  | ~n8564;
  assign \new_[16681]_  = \new_[17641]_  & \new_[29268]_ ;
  assign \new_[16682]_  = ~\new_[28804]_  & (~\new_[22427]_  | ~\new_[19184]_ );
  assign \new_[16683]_  = ~\new_[18745]_  | ~\new_[31453]_  | ~n8804;
  assign \new_[16684]_  = ~\new_[18884]_  | ~\new_[31242]_  | ~n8449;
  assign \new_[16685]_  = ~\new_[18936]_  | ~\new_[31516]_  | ~n8864;
  assign \new_[16686]_  = \new_[17646]_  & \new_[29744]_ ;
  assign \new_[16687]_  = ~\new_[30130]_  & (~\new_[20741]_  | ~\new_[18963]_ );
  assign \new_[16688]_  = ~\new_[18836]_  | ~\new_[31542]_  | ~n8939;
  assign \new_[16689]_  = ~\new_[19615]_  | ~\new_[31525]_  | ~n8899;
  assign \new_[16690]_  = ~\new_[19562]_  | ~\new_[31373]_  | ~n8719;
  assign \new_[16691]_  = ~\new_[19587]_  | ~\new_[31255]_  | ~n8489;
  assign \new_[16692]_  = ~\new_[19552]_  | ~\new_[31448]_  | ~n8794;
  assign \new_[16693]_  = ~\new_[19628]_  | ~\new_[31508]_  | ~n8844;
  assign \new_[16694]_  = ~\new_[19568]_  | ~\new_[31318]_  | ~n8594;
  assign \new_[16695]_  = ~\new_[19639]_  | ~\new_[31370]_  | ~n8704;
  assign \new_[16696]_  = ~\new_[19609]_  | ~\new_[31361]_  | ~n8664;
  assign \new_[16697]_  = ~\new_[19575]_  | ~\new_[31382]_  | ~n8754;
  assign \new_[16698]_  = ~\new_[19627]_  | ~\new_[31523]_  | ~n8889;
  assign \new_[16699]_  = ~\new_[19545]_  | ~\new_[31369]_  | ~n8699;
  assign \new_[16700]_  = ~\new_[19638]_  | ~\new_[31244]_  | ~n8459;
  assign \new_[16701]_  = ~\new_[19588]_  | ~\new_[31459]_  | ~n8814;
  assign \new_[16702]_  = ~\new_[19637]_  | ~\new_[31376]_  | ~n8729;
  assign \new_[16703]_  = ~\new_[19563]_  | ~\new_[31352]_  | ~n8639;
  assign \new_[16704]_  = ~\new_[19633]_  | ~\new_[31282]_  | ~n8509;
  assign \new_[16705]_  = ~\new_[29874]_  | (~\new_[19762]_  & ~\new_[23345]_ );
  assign \new_[16706]_  = ~\new_[30215]_  | (~\new_[19764]_  & ~\new_[22573]_ );
  assign \new_[16707]_  = ~\new_[30508]_  | (~\new_[19768]_  & ~\new_[21222]_ );
  assign \new_[16708]_  = ~\new_[29260]_  | (~\new_[19773]_  & ~\new_[22146]_ );
  assign \new_[16709]_  = ~\new_[29692]_  | (~\new_[19778]_  & ~\new_[22309]_ );
  assign \new_[16710]_  = ~\new_[30774]_  | (~\new_[19777]_  & ~\new_[22172]_ );
  assign \new_[16711]_  = ~\new_[30246]_  | (~\new_[19788]_  & ~\new_[23545]_ );
  assign \new_[16712]_  = ~\new_[30615]_  | (~\new_[19791]_  & ~\new_[23556]_ );
  assign \new_[16713]_  = ~\new_[29139]_  | (~\new_[19796]_  & ~\new_[22139]_ );
  assign \new_[16714]_  = ~\new_[29887]_  | (~\new_[19808]_  & ~\new_[22358]_ );
  assign \new_[16715]_  = ~\new_[30316]_  | (~\new_[19797]_  & ~\new_[22443]_ );
  assign \new_[16716]_  = ~\new_[30084]_  | (~\new_[19812]_  & ~\new_[23754]_ );
  assign \new_[16717]_  = ~\new_[30147]_  | (~\new_[19809]_  & ~\new_[22354]_ );
  assign \new_[16718]_  = ~\new_[29560]_  | (~\new_[19795]_  & ~\new_[22269]_ );
  assign \new_[16719]_  = ~\new_[30507]_  | (~\new_[19782]_  & ~\new_[23573]_ );
  assign \new_[16720]_  = ~\new_[30021]_  | (~\new_[19815]_  & ~\new_[23867]_ );
  assign \new_[16721]_  = ~\new_[30564]_  & (~\new_[20799]_  | ~\new_[19685]_ );
  assign \new_[16722]_  = ~\new_[24820]_  & (~\new_[19825]_  | ~\new_[30097]_ );
  assign \new_[16723]_  = ~\new_[24839]_  & (~\new_[19831]_  | ~\new_[30320]_ );
  assign \new_[16724]_  = ~\new_[24881]_  & (~\new_[19837]_  | ~\new_[30172]_ );
  assign \new_[16725]_  = ~\new_[29930]_  & (~\new_[20023]_  | ~\new_[19678]_ );
  assign \new_[16726]_  = ~\new_[30174]_  & (~\new_[21693]_  | ~\new_[19675]_ );
  assign n8474 = m2_s0_cyc_o_reg;
  assign n8449 = m4_s0_cyc_o_reg;
  assign n8619 = m5_s1_cyc_o_reg;
  assign n8789 = m7_s0_cyc_o_reg;
  assign \new_[16731]_  = ~\new_[25031]_  & (~\new_[19849]_  | ~\new_[29863]_ );
  assign \new_[16732]_  = ~\new_[29916]_  & (~\new_[20031]_  | ~\new_[19686]_ );
  assign \new_[16733]_  = ~\new_[25058]_  & (~\new_[19887]_  | ~\new_[30159]_ );
  assign \new_[16734]_  = ~\new_[23827]_  & (~\new_[19902]_  | ~\new_[30016]_ );
  assign \new_[16735]_  = ~\new_[30225]_  & (~\new_[20777]_  | ~\new_[19670]_ );
  assign \new_[16736]_  = ~\new_[23842]_  & (~\new_[19903]_  | ~\new_[29557]_ );
  assign \new_[16737]_  = ~\new_[30708]_  & (~\new_[20772]_  | ~\new_[19751]_ );
  assign \new_[16738]_  = ~\new_[23170]_  & (~\new_[19910]_  | ~\new_[29900]_ );
  assign \new_[16739]_  = ~\new_[24721]_  | ~\new_[18532]_ ;
  assign \new_[16740]_  = (~\new_[19662]_  | ~\new_[29794]_ ) & (~\new_[30612]_  | ~\new_[6174]_ );
  assign \new_[16741]_  = \new_[6036]_  ? \new_[28908]_  : \new_[19923]_ ;
  assign \new_[16742]_  = (~\new_[19718]_  | ~\new_[30071]_ ) & (~\new_[30780]_  | ~\new_[31400]_ );
  assign \new_[16743]_  = \new_[6042]_  ? \new_[29112]_  : \new_[19927]_ ;
  assign \new_[16744]_  = \new_[6045]_  ? \new_[28968]_  : \new_[19932]_ ;
  assign \new_[16745]_  = \new_[6051]_  ? \new_[28835]_  : \new_[19936]_ ;
  assign \new_[16746]_  = (~\new_[19715]_  | ~\new_[30160]_ ) & (~\new_[30711]_  | ~\new_[6049]_ );
  assign \new_[16747]_  = \new_[6053]_  ? \new_[29922]_  : \new_[19666]_ ;
  assign \new_[16748]_  = (~\new_[19680]_  | ~\new_[30207]_ ) & (~\new_[30701]_  | ~\new_[31406]_ );
  assign \new_[16749]_  = (~\new_[19739]_  | ~\new_[30349]_ ) & (~\new_[30675]_  | ~\new_[6197]_ );
  assign \new_[16750]_  = \new_[6195]_  ? \new_[30294]_  : \new_[19727]_ ;
  assign \new_[16751]_  = (~\new_[19705]_  | ~\new_[29877]_ ) & (~\new_[30478]_  | ~\new_[6211]_ );
  assign \new_[16752]_  = \new_[6273]_  ? \new_[30083]_  : \new_[19659]_ ;
  assign \new_[16753]_  = \new_[6067]_  ? \new_[28911]_  : \new_[19941]_ ;
  assign \new_[16754]_  = \new_[6193]_  ? \new_[29633]_  : \new_[19925]_ ;
  assign \new_[16755]_  = \new_[6074]_  ? \new_[28864]_  : \new_[19950]_ ;
  assign \new_[16756]_  = \new_[5992]_  ? \new_[29785]_  : \new_[19729]_ ;
  assign \new_[16757]_  = \new_[6075]_  ? \new_[28844]_  : \new_[19934]_ ;
  assign \new_[16758]_  = (~\new_[19717]_  | ~\new_[30278]_ ) & (~\new_[30501]_  | ~\new_[6079]_ );
  assign \new_[16759]_  = \new_[6083]_  ? \new_[29189]_  : \new_[19956]_ ;
  assign \new_[16760]_  = \new_[6086]_  ? \new_[29886]_  : \new_[19733]_ ;
  assign \new_[16761]_  = (~\new_[19676]_  | ~\new_[30218]_ ) & (~\new_[30713]_  | ~\new_[31499]_ );
  assign \new_[16762]_  = (~\new_[19754]_  | ~\new_[29897]_ ) & (~\new_[30545]_  | ~\new_[6093]_ );
  assign \new_[16763]_  = (~\new_[19665]_  | ~\new_[30726]_ ) & (~\new_[28672]_  | ~\new_[30726]_ );
  assign \new_[16764]_  = (~\new_[19677]_  | ~\new_[30750]_ ) & (~\new_[29123]_  | ~\new_[30750]_ );
  assign \new_[16765]_  = (~\new_[19725]_  | ~\new_[30721]_ ) & (~\new_[28515]_  | ~\new_[30721]_ );
  assign \new_[16766]_  = (~\new_[19736]_  | ~\new_[30246]_ ) & (~\new_[26263]_  | ~\new_[30246]_ );
  assign \new_[16767]_  = (~\new_[19730]_  | ~\new_[30615]_ ) & (~\new_[27835]_  | ~\new_[30615]_ );
  assign \new_[16768]_  = (~\new_[19708]_  | ~\new_[30574]_ ) & (~\new_[26725]_  | ~\new_[30574]_ );
  assign \new_[16769]_  = (~\new_[19721]_  | ~\new_[30538]_ ) & (~\new_[28655]_  | ~\new_[30538]_ );
  assign \new_[16770]_  = (~\new_[19671]_  | ~\new_[30784]_ ) & (~\new_[28103]_  | ~\new_[30784]_ );
  assign \new_[16771]_  = (~\new_[19697]_  | ~\new_[30084]_ ) & (~\new_[26222]_  | ~\new_[30084]_ );
  assign \new_[16772]_  = (~\new_[19737]_  | ~\new_[30789]_ ) & (~\new_[28238]_  | ~\new_[30789]_ );
  assign \new_[16773]_  = (~\new_[19738]_  | ~\new_[30507]_ ) & (~\new_[29051]_  | ~\new_[30507]_ );
  assign \new_[16774]_  = (~\new_[19758]_  | ~\new_[30820]_ ) & (~\new_[28407]_  | ~\new_[30820]_ );
  assign \new_[16775]_  = ~\new_[22372]_  & (~\new_[19550]_  | ~\new_[30754]_ );
  assign \new_[16776]_  = ~\new_[22143]_  & (~\new_[19553]_  | ~\new_[30676]_ );
  assign \new_[16777]_  = ~\new_[20311]_  & (~\new_[19592]_  | ~\new_[30563]_ );
  assign \new_[16778]_  = ~\new_[22243]_  & (~\new_[19574]_  | ~\new_[30775]_ );
  assign \new_[16779]_  = ~\new_[23833]_  & (~\new_[19602]_  | ~\new_[30725]_ );
  assign \new_[16780]_  = \new_[19119]_  | \new_[30078]_ ;
  assign \new_[16781]_  = \new_[19112]_  | \new_[30206]_ ;
  assign \new_[16782]_  = ~\new_[19110]_  & ~\new_[22226]_ ;
  assign \new_[16783]_  = \new_[19117]_  | \new_[29169]_ ;
  assign \new_[16784]_  = \new_[19115]_  | \new_[29300]_ ;
  assign \new_[16785]_  = ~\new_[19120]_  & ~\new_[23726]_ ;
  assign \new_[16786]_  = ~\new_[19109]_  & ~\new_[22227]_ ;
  assign \new_[16787]_  = ~\new_[19121]_  & ~\new_[23837]_ ;
  assign \new_[16788]_  = \new_[19122]_  | \new_[30072]_ ;
  assign \new_[16789]_  = \new_[19193]_  | \new_[27639]_ ;
  assign \new_[16790]_  = ~\new_[19221]_  & ~\new_[23334]_ ;
  assign \new_[16791]_  = \new_[19094]_  | \new_[27540]_ ;
  assign \new_[16792]_  = \new_[25178]_  & \new_[18947]_ ;
  assign \new_[16793]_  = ~\new_[22140]_  & (~\new_[20001]_  | ~\new_[22868]_ );
  assign \new_[16794]_  = ~\new_[26679]_  & (~\new_[20129]_  | ~\new_[30164]_ );
  assign \new_[16795]_  = ~\new_[28162]_  & (~\new_[19997]_  | ~\new_[28114]_ );
  assign \new_[16796]_  = \new_[19048]_  | \new_[24346]_ ;
  assign \new_[16797]_  = \new_[19231]_  | \new_[26673]_ ;
  assign \new_[16798]_  = \new_[19222]_  | \new_[28398]_ ;
  assign \new_[16799]_  = \new_[18746]_  & \new_[26811]_ ;
  assign \new_[16800]_  = \new_[25211]_  & \new_[18948]_ ;
  assign \new_[16801]_  = ~\new_[26250]_  & (~\new_[20002]_  | ~\new_[28908]_ );
  assign \new_[16802]_  = ~\new_[26839]_  | (~\new_[20041]_  & ~\new_[28992]_ );
  assign \new_[16803]_  = ~\new_[25088]_  & (~\new_[20119]_  | ~\new_[24319]_ );
  assign \new_[16804]_  = \new_[22470]_  & \new_[18951]_ ;
  assign \new_[16805]_  = \new_[18975]_  | \new_[23113]_ ;
  assign \new_[16806]_  = ~\new_[24675]_  | ~\new_[19129]_  | ~\new_[24824]_ ;
  assign \new_[16807]_  = \new_[19194]_  | \new_[22978]_ ;
  assign \new_[16808]_  = \new_[22466]_  & \new_[18944]_ ;
  assign \new_[16809]_  = ~\new_[19236]_  & ~\new_[21234]_ ;
  assign \new_[16810]_  = ~\new_[24566]_  & (~\new_[20100]_  | ~\new_[29435]_ );
  assign \new_[16811]_  = ~\new_[26225]_  & (~\new_[20012]_  | ~\new_[29159]_ );
  assign \new_[16812]_  = \new_[19234]_  | \new_[26225]_ ;
  assign \new_[16813]_  = \new_[18847]_  & \new_[28134]_ ;
  assign \new_[16814]_  = \new_[19223]_  | \new_[28654]_ ;
  assign \new_[16815]_  = ~\new_[25351]_  & (~\new_[20092]_  | ~\new_[29112]_ );
  assign \new_[16816]_  = ~\new_[28541]_  | (~\new_[20013]_  & ~\new_[29541]_ );
  assign \new_[16817]_  = ~\new_[27559]_  & (~\new_[20047]_  | ~\new_[28188]_ );
  assign \new_[16818]_  = ~\new_[24840]_  & (~\new_[20015]_  | ~\new_[24313]_ );
  assign \new_[16819]_  = ~\new_[28186]_  | (~\new_[20077]_  & ~\new_[29115]_ );
  assign \new_[16820]_  = \new_[18985]_  | \new_[22939]_ ;
  assign \new_[16821]_  = ~\new_[28722]_  | (~\new_[20019]_  & ~\new_[29815]_ );
  assign \new_[16822]_  = ~\new_[28722]_  | ~\new_[19833]_  | ~\new_[20286]_ ;
  assign \new_[16823]_  = \new_[19195]_  | \new_[24352]_ ;
  assign \new_[16824]_  = \new_[19196]_  | \new_[27591]_ ;
  assign \new_[16825]_  = \new_[22501]_  & \new_[18946]_ ;
  assign \new_[16826]_  = ~\new_[27773]_  & (~\new_[20021]_  | ~\new_[29983]_ );
  assign \new_[16827]_  = ~m4_stb_i | ~\new_[19608]_  | ~\new_[28768]_ ;
  assign \new_[16828]_  = \new_[25198]_  & \new_[18953]_ ;
  assign \new_[16829]_  = ~\new_[19060]_  | ~\new_[31698]_ ;
  assign \new_[16830]_  = ~\new_[26200]_  & (~\new_[20022]_  | ~\new_[29633]_ );
  assign \new_[16831]_  = \new_[19225]_  | \new_[27821]_ ;
  assign \new_[16832]_  = \new_[18777]_  & \new_[27973]_ ;
  assign \new_[16833]_  = ~\new_[26206]_  & (~\new_[20025]_  | ~\new_[28968]_ );
  assign \new_[16834]_  = ~\new_[27602]_  | (~\new_[20033]_  & ~\new_[29217]_ );
  assign \new_[16835]_  = ~\new_[24864]_  & (~\new_[20026]_  | ~\new_[24272]_ );
  assign \new_[16836]_  = ~\new_[28210]_  | (~\new_[20016]_  & ~\new_[29930]_ );
  assign \new_[16837]_  = \new_[18991]_  & \new_[31678]_ ;
  assign \new_[16838]_  = ~\new_[28210]_  | ~\new_[19839]_  | ~\new_[20309]_ ;
  assign \new_[16839]_  = \new_[19197]_  | \new_[26552]_ ;
  assign \new_[16840]_  = ~\new_[23162]_  & (~\new_[20126]_  | ~\new_[28969]_ );
  assign \new_[16841]_  = ~\new_[27571]_  & (~\new_[19991]_  | ~\new_[28050]_ );
  assign \new_[16842]_  = \new_[19226]_  | \new_[27597]_ ;
  assign \new_[16843]_  = ~\new_[24812]_  & (~\new_[19994]_  | ~\new_[28835]_ );
  assign \new_[16844]_  = ~\new_[28510]_  | (~\new_[20099]_  & ~\new_[29058]_ );
  assign \new_[16845]_  = \new_[18995]_  & \new_[31830]_ ;
  assign \new_[16846]_  = ~s2_ack_i | ~\new_[18786]_  | ~\new_[30085]_ ;
  assign \new_[16847]_  = ~\new_[23729]_  & (~\new_[20088]_  | ~\new_[22962]_ );
  assign \new_[16848]_  = ~\new_[24752]_  & (~\new_[20039]_  | ~\new_[29186]_ );
  assign \new_[16849]_  = ~\new_[24677]_  & (~\new_[20068]_  | ~\new_[29397]_ );
  assign \new_[16850]_  = \new_[19227]_  | \new_[24677]_ ;
  assign \new_[16851]_  = ~s5_err_i | ~\new_[18795]_  | ~\new_[29036]_ ;
  assign \new_[16852]_  = ~\new_[22379]_  & (~\new_[19995]_  | ~\new_[23002]_ );
  assign \new_[16853]_  = \new_[19224]_  | \new_[28406]_ ;
  assign \new_[16854]_  = ~s2_err_i | ~\new_[18786]_  | ~\new_[30085]_ ;
  assign \new_[16855]_  = \new_[22492]_  & \new_[18945]_ ;
  assign \new_[16856]_  = \new_[18768]_  & \new_[26271]_ ;
  assign \new_[16857]_  = ~s2_rty_i | ~\new_[18786]_  | ~\new_[30085]_ ;
  assign \new_[16858]_  = ~\new_[28570]_  | ~\new_[19146]_  | ~\new_[22261]_ ;
  assign \new_[16859]_  = ~s1_ack_i | ~\new_[18799]_  | ~\new_[30357]_ ;
  assign \new_[16860]_  = ~\new_[19237]_  & ~\new_[22214]_ ;
  assign \new_[16861]_  = ~s6_ack_i | ~\new_[18803]_  | ~\new_[29298]_ ;
  assign \new_[16862]_  = \new_[18800]_  & \new_[24290]_ ;
  assign \new_[16863]_  = ~s0_ack_i | ~\new_[18808]_  | ~\new_[30481]_ ;
  assign \new_[16864]_  = ~\new_[26955]_  & (~\new_[19998]_  | ~\new_[23184]_ );
  assign \new_[16865]_  = \new_[24537]_  & \new_[18943]_ ;
  assign \new_[16866]_  = ~\new_[26729]_  & (~\new_[20106]_  | ~\new_[29682]_ );
  assign \new_[16867]_  = ~\new_[26419]_  & (~\new_[20080]_  | ~\new_[29212]_ );
  assign \new_[16868]_  = \new_[19211]_  & \new_[27642]_ ;
  assign \new_[16869]_  = ~\new_[26732]_  & (~\new_[20049]_  | ~\new_[29831]_ );
  assign \new_[16870]_  = \new_[19243]_  | \new_[26732]_ ;
  assign \new_[16871]_  = \new_[18838]_  & \new_[27846]_ ;
  assign \new_[16872]_  = ~s6_err_i | ~\new_[18803]_  | ~\new_[29298]_ ;
  assign \new_[16873]_  = ~\new_[26604]_  & (~\new_[20069]_  | ~\new_[28121]_ );
  assign \new_[16874]_  = \new_[22489]_  & \new_[18949]_ ;
  assign \new_[16875]_  = ~s0_err_i | ~\new_[18808]_  | ~\new_[30481]_ ;
  assign \new_[16876]_  = ~\new_[28369]_  & (~\new_[19999]_  | ~\new_[30552]_ );
  assign \new_[16877]_  = \new_[22500]_  & \new_[18952]_ ;
  assign \new_[16878]_  = ~s9_rty_i | ~\new_[18806]_  | ~\new_[29709]_ ;
  assign \new_[16879]_  = ~s6_rty_i | ~\new_[18803]_  | ~\new_[29298]_ ;
  assign \new_[16880]_  = ~s0_rty_i | ~\new_[18808]_  | ~\new_[30481]_ ;
  assign \new_[16881]_  = ~\new_[19011]_  | ~\new_[31830]_ ;
  assign \new_[16882]_  = ~\new_[19010]_  & ~\new_[24469]_ ;
  assign \new_[16883]_  = ~\new_[28420]_  | (~\new_[20144]_  & ~\new_[29700]_ );
  assign \new_[16884]_  = \new_[19203]_  | \new_[24343]_ ;
  assign \new_[16885]_  = ~\new_[19228]_  & ~\new_[21242]_ ;
  assign \new_[16886]_  = ~\new_[28135]_  & (~\new_[20139]_  | ~\new_[30751]_ );
  assign \new_[16887]_  = \new_[25166]_  & \new_[18955]_ ;
  assign \new_[16888]_  = ~\new_[28251]_  & (~\new_[20072]_  | ~\new_[29040]_ );
  assign \new_[16889]_  = \new_[23148]_  & \new_[18954]_ ;
  assign \new_[16890]_  = \new_[18815]_  & \new_[26220]_ ;
  assign \new_[16891]_  = ~\new_[19058]_  | ~\new_[31576]_ ;
  assign \new_[16892]_  = ~\new_[19050]_  & ~\new_[23174]_ ;
  assign \new_[16893]_  = ~\new_[28574]_  | (~\new_[20096]_  & ~\new_[29157]_ );
  assign \new_[16894]_  = ~\new_[26741]_  | ~\new_[19167]_  | ~\new_[21213]_ ;
  assign \new_[16895]_  = \new_[19198]_  | \new_[24359]_ ;
  assign \new_[16896]_  = \new_[24670]_  & \new_[18950]_ ;
  assign \new_[16897]_  = \new_[18816]_  & \new_[28133]_ ;
  assign \new_[16898]_  = \new_[19230]_  | \new_[27580]_ ;
  assign \new_[16899]_  = \new_[18770]_  & \new_[26283]_ ;
  assign \new_[16900]_  = ~\new_[28546]_  & (~\new_[20074]_  | ~\new_[30554]_ );
  assign \new_[16901]_  = ~\new_[18966]_  | ~\new_[31759]_ ;
  assign \new_[16902]_  = ~\new_[23798]_  & (~\new_[20082]_  | ~\new_[26297]_ );
  assign \new_[16903]_  = \new_[19033]_  | \new_[23045]_ ;
  assign \new_[16904]_  = \new_[19201]_  | \new_[26547]_ ;
  assign \new_[16905]_  = ~\new_[27624]_  & (~\new_[20110]_  | ~\new_[28245]_ );
  assign \new_[16906]_  = ~\new_[28384]_  | (~\new_[20133]_  & ~\new_[29101]_ );
  assign \new_[16907]_  = ~\new_[28554]_  | (~\new_[20075]_  & ~\new_[29254]_ );
  assign \new_[16908]_  = \new_[19229]_  | \new_[28546]_ ;
  assign \new_[16909]_  = ~\new_[22289]_  & (~\new_[20078]_  | ~\new_[22915]_ );
  assign \new_[16910]_  = ~\new_[26233]_  & (~\new_[20148]_  | ~\new_[28844]_ );
  assign \new_[16911]_  = ~\new_[26943]_  & (~\new_[20081]_  | ~\new_[27802]_ );
  assign \new_[16912]_  = ~\new_[24550]_  & (~\new_[20150]_  | ~\new_[29175]_ );
  assign \new_[16913]_  = ~\new_[27698]_  & (~\new_[20083]_  | ~\new_[28073]_ );
  assign \new_[16914]_  = \new_[18844]_  & \new_[27425]_ ;
  assign \new_[16915]_  = ~\new_[24768]_  & (~\new_[20090]_  | ~\new_[28864]_ );
  assign \new_[16916]_  = ~\new_[19233]_  & ~\new_[21240]_ ;
  assign \new_[16917]_  = \new_[19232]_  | \new_[24374]_ ;
  assign \new_[16918]_  = \new_[18782]_  & \new_[26776]_ ;
  assign \new_[16919]_  = ~\new_[28291]_  | (~\new_[20064]_  & ~\new_[29229]_ );
  assign \new_[16920]_  = ~m6_stb_i | ~\new_[18789]_  | ~\new_[30227]_ ;
  assign \new_[16921]_  = ~m2_stb_i | ~\new_[19571]_  | ~\new_[29021]_ ;
  assign \new_[16922]_  = ~\new_[26204]_  & (~\new_[20070]_  | ~\new_[28911]_ );
  assign \new_[16923]_  = \new_[19199]_  | \new_[26504]_ ;
  assign \new_[16924]_  = \new_[19219]_  & \new_[29413]_ ;
  assign \new_[16925]_  = ~\new_[28176]_  | ~\new_[19873]_  | ~\new_[20339]_ ;
  assign \new_[16926]_  = \new_[19088]_  | \new_[24644]_ ;
  assign \new_[16927]_  = \new_[25200]_  & \new_[18957]_ ;
  assign \new_[16928]_  = ~\new_[27356]_  & (~\new_[20135]_  | ~\new_[29038]_ );
  assign \new_[16929]_  = ~\new_[26757]_  | ~\new_[19177]_  | ~\new_[25060]_ ;
  assign \new_[16930]_  = \new_[18976]_  & \new_[31698]_ ;
  assign \new_[16931]_  = ~\new_[28294]_  | (~\new_[20101]_  & ~\new_[29167]_ );
  assign \new_[16932]_  = \new_[19217]_  & \new_[27694]_ ;
  assign \new_[16933]_  = ~\new_[24981]_  & (~\new_[20066]_  | ~\new_[24287]_ );
  assign \new_[16934]_  = ~\new_[25000]_  & (~\new_[20105]_  | ~\new_[24344]_ );
  assign \new_[16935]_  = ~\new_[24363]_  & (~\new_[19993]_  | ~\new_[28535]_ );
  assign \new_[16936]_  = \new_[19202]_  | \new_[24362]_ ;
  assign \new_[16937]_  = \new_[19038]_  | \new_[26431]_ ;
  assign \new_[16938]_  = \new_[19235]_  | \new_[26414]_ ;
  assign \new_[16939]_  = ~\new_[24337]_  & (~\new_[20111]_  | ~\new_[30333]_ );
  assign \new_[16940]_  = ~\new_[28176]_  | (~\new_[20091]_  & ~\new_[30188]_ );
  assign \new_[16941]_  = \new_[22462]_  & \new_[18956]_ ;
  assign \new_[16942]_  = \new_[18840]_  & \new_[23155]_ ;
  assign \new_[16943]_  = \new_[19063]_  | \new_[24341]_ ;
  assign \new_[16944]_  = \new_[19238]_  | \new_[26560]_ ;
  assign \new_[16945]_  = \new_[18874]_  & \new_[27606]_ ;
  assign \new_[16946]_  = \new_[19080]_  | \new_[24558]_ ;
  assign \new_[16947]_  = ~\new_[28674]_  | ~\new_[20687]_  | ~\new_[20352]_ ;
  assign \new_[16948]_  = \new_[18939]_  & \new_[26701]_ ;
  assign \new_[16949]_  = ~\new_[28674]_  | (~\new_[20127]_  & ~\new_[30010]_ );
  assign \new_[16950]_  = ~s6_ack_i | ~\new_[18881]_  | ~\new_[28767]_ ;
  assign \new_[16951]_  = ~s5_err_i | ~\new_[19608]_  | ~\new_[28768]_ ;
  assign \new_[16952]_  = ~\new_[28606]_  | (~\new_[20137]_  & ~\new_[29047]_ );
  assign \new_[16953]_  = ~\new_[26874]_  | ~\new_[19176]_  | ~\new_[21185]_ ;
  assign \new_[16954]_  = ~s6_err_i | ~\new_[18881]_  | ~\new_[28767]_ ;
  assign \new_[16955]_  = ~m6_stb_i | ~\new_[18786]_  | ~\new_[30085]_ ;
  assign \new_[16956]_  = ~s5_rty_i | ~\new_[19608]_  | ~\new_[28768]_ ;
  assign \new_[16957]_  = ~s6_rty_i | ~\new_[18881]_  | ~\new_[28767]_ ;
  assign \new_[16958]_  = \new_[18867]_  & \new_[27907]_ ;
  assign \new_[16959]_  = ~\new_[26414]_  & (~\new_[20132]_  | ~\new_[29571]_ );
  assign \new_[16960]_  = ~\new_[27689]_  & (~\new_[20103]_  | ~\new_[28007]_ );
  assign \new_[16961]_  = \new_[18868]_  & \new_[26572]_ ;
  assign \new_[16962]_  = \new_[18911]_  & \new_[23096]_ ;
  assign \new_[16963]_  = ~\new_[19240]_  & ~\new_[21247]_ ;
  assign \new_[16964]_  = ~\new_[26279]_  & (~\new_[20136]_  | ~\new_[29189]_ );
  assign \new_[16965]_  = \new_[22490]_  & \new_[18958]_ ;
  assign \new_[16966]_  = \new_[19200]_  | \new_[24002]_ ;
  assign \new_[16967]_  = \new_[19241]_  | \new_[28135]_ ;
  assign \new_[16968]_  = \new_[19204]_  | \new_[27765]_ ;
  assign \new_[16969]_  = ~\new_[19028]_  & ~\new_[23082]_ ;
  assign \new_[16970]_  = ~\new_[27130]_  | (~\new_[20140]_  & ~\new_[29671]_ );
  assign \new_[16971]_  = ~\new_[18996]_  & ~\new_[23239]_ ;
  assign \new_[16972]_  = ~\new_[28346]_  | (~\new_[20035]_  & ~\new_[29354]_ );
  assign \new_[16973]_  = ~\new_[26704]_  | ~\new_[19188]_  | ~\new_[21169]_ ;
  assign \new_[16974]_  = \new_[19205]_  | \new_[23512]_ ;
  assign \new_[16975]_  = ~\new_[19242]_  & ~\new_[21159]_ ;
  assign \new_[16976]_  = ~\new_[27950]_  | ~\new_[19150]_  | ~\new_[21158]_ ;
  assign \new_[16977]_  = \new_[22467]_  & \new_[18959]_ ;
  assign \new_[16978]_  = ~\new_[29372]_  & (~\new_[20124]_  | ~\new_[29996]_ );
  assign \new_[16979]_  = \new_[19239]_  | \new_[28092]_ ;
  assign \new_[16980]_  = \new_[19079]_  & \new_[31804]_ ;
  assign \new_[16981]_  = ~\new_[28193]_  | (~\new_[20152]_  & ~\new_[29172]_ );
  assign \new_[16982]_  = ~\new_[28074]_  | ~\new_[19192]_  | ~\new_[22459]_ ;
  assign \new_[16983]_  = \new_[19123]_  | \new_[27639]_ ;
  assign \new_[16984]_  = ~\new_[26668]_  & (~\new_[21653]_  | ~\new_[30097]_ );
  assign \new_[16985]_  = \new_[19128]_  | \new_[28380]_ ;
  assign \new_[16986]_  = ~\new_[27733]_  & (~\new_[21817]_  | ~\new_[30320]_ );
  assign \new_[16987]_  = \new_[19165]_  | \new_[27962]_ ;
  assign \new_[16988]_  = ~\new_[27667]_  & (~\new_[21692]_  | ~\new_[30159]_ );
  assign \new_[16989]_  = \new_[19133]_  | \new_[27591]_ ;
  assign \new_[16990]_  = ~\new_[27626]_  & (~\new_[21715]_  | ~\new_[30172]_ );
  assign \new_[16991]_  = \new_[19135]_  | \new_[28098]_ ;
  assign \new_[16992]_  = \new_[19132]_  | \new_[26552]_ ;
  assign \new_[16993]_  = ~\new_[26636]_  & (~\new_[20147]_  | ~\new_[29762]_ );
  assign \new_[16994]_  = ~\new_[27979]_  & (~\new_[20142]_  | ~\new_[30697]_ );
  assign \new_[16995]_  = \new_[19125]_  | \new_[24352]_ ;
  assign \new_[16996]_  = \new_[19153]_  | \new_[24362]_ ;
  assign \new_[16997]_  = \new_[19163]_  | \new_[24359]_ ;
  assign \new_[16998]_  = ~\new_[27752]_  & (~\new_[20089]_  | ~\new_[30092]_ );
  assign \new_[16999]_  = ~\new_[27665]_  & (~\new_[21852]_  | ~\new_[29863]_ );
  assign \new_[17000]_  = ~\new_[26276]_  & (~\new_[20007]_  | ~\new_[29299]_ );
  assign \new_[17001]_  = \new_[19174]_  | \new_[26195]_ ;
  assign \new_[17002]_  = \new_[19172]_  | \new_[27582]_ ;
  assign \new_[17003]_  = \new_[19173]_  | \new_[26208]_ ;
  assign \new_[17004]_  = \new_[19130]_  | \new_[27743]_ ;
  assign \new_[17005]_  = ~\new_[24414]_  & (~\new_[20052]_  | ~\new_[28001]_ );
  assign \new_[17006]_  = ~\new_[26913]_  & (~\new_[20109]_  | ~\new_[29888]_ );
  assign \new_[17007]_  = \new_[19180]_  | \new_[26547]_ ;
  assign \new_[17008]_  = ~\new_[27664]_  & (~\new_[20104]_  | ~\new_[30061]_ );
  assign \new_[17009]_  = \new_[19152]_  | \new_[24343]_ ;
  assign \new_[17010]_  = \new_[19171]_  | \new_[27765]_ ;
  assign \new_[17011]_  = \new_[19189]_  | \new_[23512]_ ;
  assign \new_[17012]_  = ~\new_[29215]_  | ~\new_[20539]_  | ~s1_ack_i;
  assign \new_[17013]_  = ~\new_[23339]_  & (~\new_[20153]_  | ~\new_[27463]_ );
  assign \new_[17014]_  = ~s2_ack_i | ~\new_[18740]_  | ~\new_[30013]_ ;
  assign \new_[17015]_  = ~s6_ack_i | ~\new_[18742]_  | ~\new_[29704]_ ;
  assign \new_[17016]_  = ~s0_ack_i | ~\new_[18745]_  | ~\new_[29258]_ ;
  assign \new_[17017]_  = ~m5_stb_i | ~\new_[20544]_  | ~\new_[29628]_ ;
  assign \new_[17018]_  = ~s10_ack_i | ~\new_[19544]_  | ~\new_[29045]_ ;
  assign \new_[17019]_  = ~s3_err_i | ~\new_[18735]_  | ~\new_[29928]_ ;
  assign \new_[17020]_  = ~s0_err_i | ~\new_[18745]_  | ~\new_[29258]_ ;
  assign \new_[17021]_  = ~s10_err_i | ~\new_[19544]_  | ~\new_[29045]_ ;
  assign \new_[17022]_  = ~s6_err_i | ~\new_[18742]_  | ~\new_[29704]_ ;
  assign \new_[17023]_  = ~s3_rty_i | ~\new_[18735]_  | ~\new_[29928]_ ;
  assign \new_[17024]_  = ~\new_[29855]_  & (~\new_[20185]_  | ~\new_[26262]_ );
  assign \new_[17025]_  = ~s10_rty_i | ~\new_[19544]_  | ~\new_[29045]_ ;
  assign \new_[17026]_  = ~s0_rty_i | ~\new_[18745]_  | ~\new_[29258]_ ;
  assign \new_[17027]_  = ~\new_[29648]_  & (~\new_[20158]_  | ~\new_[26430]_ );
  assign \new_[17028]_  = ~\new_[29100]_  & (~\new_[20174]_  | ~\new_[26515]_ );
  assign \new_[17029]_  = ~\new_[19043]_  | ~\new_[24475]_ ;
  assign \new_[17030]_  = ~\new_[29649]_  | ~\new_[18937]_  | ~m0_stb_i;
  assign \new_[17031]_  = ~m1_stb_i | ~\new_[18919]_  | ~\new_[29025]_ ;
  assign \new_[17032]_  = ~m3_stb_i | ~\new_[18734]_  | ~\new_[29948]_ ;
  assign \new_[17033]_  = ~\new_[18989]_  | ~\new_[23127]_ ;
  assign \new_[17034]_  = ~\new_[30389]_  & (~\new_[20159]_  | ~\new_[26342]_ );
  assign \new_[17035]_  = ~\new_[30174]_  & (~\new_[20269]_  | ~\new_[29305]_ );
  assign \new_[17036]_  = ~\new_[19099]_  | ~\new_[23937]_ ;
  assign \new_[17037]_  = ~\new_[29916]_  & (~\new_[20271]_  | ~\new_[29601]_ );
  assign \new_[17038]_  = ~m7_stb_i | ~\new_[18830]_  | ~\new_[29707]_ ;
  assign \new_[17039]_  = ~\new_[30044]_  & (~\new_[20180]_  | ~\new_[27353]_ );
  assign \new_[17040]_  = ~\new_[30185]_  & (~\new_[20279]_  | ~\new_[29351]_ );
  assign \new_[17041]_  = ~\new_[29711]_  | ~\new_[18766]_  | ~s12_ack_i;
  assign \new_[17042]_  = ~\new_[18997]_  | ~\new_[24340]_ ;
  assign \new_[17043]_  = ~s13_ack_i | ~\new_[18849]_  | ~\new_[32168]_ ;
  assign \new_[17044]_  = ~m3_stb_i | ~\new_[20567]_  | ~\new_[30131]_ ;
  assign \new_[17045]_  = ~s9_rty_i | ~\new_[18850]_  | ~\new_[29024]_ ;
  assign \new_[17046]_  = \new_[18784]_  & \new_[29708]_ ;
  assign \new_[17047]_  = \new_[18841]_  | \new_[21240]_ ;
  assign \new_[17048]_  = ~\new_[19025]_  | ~\new_[24437]_ ;
  assign \new_[17049]_  = ~\new_[19026]_  | ~\new_[24376]_ ;
  assign \new_[17050]_  = ~s7_ack_i | ~\new_[18832]_  | ~\new_[28313]_ ;
  assign \new_[17051]_  = ~s6_err_i | ~\new_[18831]_  | ~\new_[29707]_ ;
  assign \new_[17052]_  = ~s7_err_i | ~\new_[18832]_  | ~\new_[28313]_ ;
  assign \new_[17053]_  = ~s6_rty_i | ~\new_[18831]_  | ~\new_[29707]_ ;
  assign \new_[17054]_  = ~s7_rty_i | ~\new_[18832]_  | ~\new_[28313]_ ;
  assign \new_[17055]_  = ~\new_[29331]_  & (~\new_[20168]_  | ~\new_[27725]_ );
  assign \new_[17056]_  = ~\new_[22194]_  & (~\new_[20176]_  | ~\new_[27640]_ );
  assign \new_[17057]_  = ~m1_stb_i | ~\new_[18907]_  | ~\new_[29705]_ ;
  assign \new_[17058]_  = \new_[18934]_  | \new_[21247]_ ;
  assign \new_[17059]_  = ~s9_ack_i | ~\new_[18850]_  | ~\new_[29024]_ ;
  assign \new_[17060]_  = ~s5_err_i | ~\new_[19539]_  | ~\new_[29948]_ ;
  assign \new_[17061]_  = ~s13_err_i | ~\new_[18849]_  | ~\new_[32168]_ ;
  assign \new_[17062]_  = ~m1_stb_i | ~\new_[20572]_  | ~\new_[30260]_ ;
  assign \new_[17063]_  = ~s0_err_i | ~\new_[18936]_  | ~\new_[29819]_ ;
  assign \new_[17064]_  = ~\new_[29898]_  & (~\new_[20172]_  | ~\new_[26358]_ );
  assign \new_[17065]_  = ~s13_rty_i | ~\new_[18849]_  | ~\new_[32168]_ ;
  assign \new_[17066]_  = ~\new_[30445]_  & (~\new_[20282]_  | ~\new_[29536]_ );
  assign \new_[17067]_  = ~\new_[19077]_  | ~\new_[22175]_ ;
  assign \new_[17068]_  = ~s6_ack_i | ~\new_[18829]_  | ~\new_[29707]_ ;
  assign \new_[17069]_  = ~m1_stb_i | ~\new_[18888]_  | ~\new_[30189]_ ;
  assign \new_[17070]_  = ~s1_ack_i | ~\new_[18887]_  | ~\new_[30195]_ ;
  assign \new_[17071]_  = ~s2_ack_i | ~\new_[20541]_  | ~\new_[30189]_ ;
  assign \new_[17072]_  = ~s8_ack_i | ~\new_[19621]_  | ~\new_[29670]_ ;
  assign \new_[17073]_  = ~s11_ack_i | ~\new_[18894]_  | ~\new_[30260]_ ;
  assign \new_[17074]_  = ~\new_[28982]_  & (~\new_[20199]_  | ~\new_[27721]_ );
  assign \new_[17075]_  = ~s12_ack_i | ~\new_[20573]_  | ~\new_[28957]_ ;
  assign \new_[17076]_  = ~s5_ack_i | ~\new_[18734]_  | ~\new_[29948]_ ;
  assign \new_[17077]_  = ~\new_[19089]_  | ~\new_[26390]_ ;
  assign \new_[17078]_  = ~s13_ack_i | ~\new_[18905]_  | ~\new_[32327]_ ;
  assign \new_[17079]_  = ~s9_ack_i | ~\new_[18906]_  | ~\new_[30354]_ ;
  assign \new_[17080]_  = ~s6_ack_i | ~\new_[18910]_  | ~\new_[29052]_ ;
  assign \new_[17081]_  = ~s7_ack_i | ~\new_[18912]_  | ~\new_[30031]_ ;
  assign \new_[17082]_  = ~s3_ack_i | ~\new_[19633]_  | ~\new_[30469]_ ;
  assign \new_[17083]_  = ~s5_ack_i | ~\new_[18925]_  | ~\new_[29025]_ ;
  assign \new_[17084]_  = ~s8_err_i | ~\new_[18890]_  | ~\new_[29670]_ ;
  assign \new_[17085]_  = ~s11_err_i | ~\new_[20572]_  | ~\new_[30260]_ ;
  assign \new_[17086]_  = ~s11_ack_i | ~\new_[18929]_  | ~\new_[30200]_ ;
  assign \new_[17087]_  = ~s5_err_i | ~\new_[18919]_  | ~\new_[29025]_ ;
  assign \new_[17088]_  = ~\new_[29035]_  | ~\new_[18932]_  | ~s3_ack_i;
  assign \new_[17089]_  = ~s13_err_i | ~\new_[18905]_  | ~\new_[32327]_ ;
  assign \new_[17090]_  = ~s6_err_i | ~\new_[18910]_  | ~\new_[29052]_ ;
  assign \new_[17091]_  = ~s7_err_i | ~\new_[18912]_  | ~\new_[30031]_ ;
  assign \new_[17092]_  = ~s1_err_i | ~\new_[18887]_  | ~\new_[30195]_ ;
  assign \new_[17093]_  = ~s2_err_i | ~\new_[20541]_  | ~\new_[30189]_ ;
  assign \new_[17094]_  = ~s5_rty_i | ~\new_[19539]_  | ~\new_[29948]_ ;
  assign \new_[17095]_  = ~s1_rty_i | ~\new_[18887]_  | ~\new_[30195]_ ;
  assign \new_[17096]_  = ~s2_rty_i | ~\new_[18888]_  | ~\new_[30189]_ ;
  assign \new_[17097]_  = ~s11_rty_i | ~\new_[20572]_  | ~\new_[30260]_ ;
  assign \new_[17098]_  = ~s13_rty_i | ~\new_[18905]_  | ~\new_[32327]_ ;
  assign \new_[17099]_  = ~s6_rty_i | ~\new_[18910]_  | ~\new_[29052]_ ;
  assign \new_[17100]_  = ~s7_rty_i | ~\new_[18912]_  | ~\new_[30031]_ ;
  assign \new_[17101]_  = ~s0_ack_i | ~\new_[18936]_  | ~\new_[29819]_ ;
  assign \new_[17102]_  = ~s3_rty_i | ~\new_[19633]_  | ~\new_[30469]_ ;
  assign \new_[17103]_  = ~s9_rty_i | ~\new_[18906]_  | ~\new_[30354]_ ;
  assign \new_[17104]_  = ~s5_rty_i | ~\new_[20576]_  | ~\new_[29025]_ ;
  assign \new_[17105]_  = ~\new_[29096]_  & (~\new_[20200]_  | ~\new_[27553]_ );
  assign \new_[17106]_  = ~\new_[29649]_  | ~\new_[18937]_  | ~s5_ack_i;
  assign \new_[17107]_  = ~s9_err_i | ~\new_[18850]_  | ~\new_[29024]_ ;
  assign \new_[17108]_  = ~\new_[29035]_  | ~\new_[18932]_  | ~m0_stb_i;
  assign \new_[17109]_  = ~\new_[29166]_  & (~\new_[20202]_  | ~\new_[26813]_ );
  assign \new_[17110]_  = ~m1_stb_i | ~\new_[19633]_  | ~\new_[30469]_ ;
  assign \new_[17111]_  = \new_[18775]_  | \new_[21159]_ ;
  assign \new_[17112]_  = ~\new_[22444]_  & (~\new_[20203]_  | ~\new_[26632]_ );
  assign \new_[17113]_  = ~\new_[29749]_  | ~\new_[20547]_  | ~m0_stb_i;
  assign \new_[17114]_  = ~\new_[23739]_  & (~\new_[20171]_  | ~\new_[26355]_ );
  assign \new_[17115]_  = ~\new_[28527]_  | ~\new_[19126]_  | ~\new_[23792]_ ;
  assign \new_[17116]_  = ~\new_[27648]_  | ~\new_[19164]_  | ~\new_[23654]_ ;
  assign \new_[17117]_  = \new_[21764]_  | \new_[19134]_ ;
  assign \new_[17118]_  = \new_[21703]_  | \new_[19159]_ ;
  assign \new_[17119]_  = ~\new_[29197]_  | ~\new_[19210]_  | ~\new_[27620]_ ;
  assign \new_[17120]_  = \new_[22165]_  | \new_[19207]_ ;
  assign \new_[17121]_  = ~\new_[27578]_  | ~\new_[19178]_  | ~\new_[23663]_ ;
  assign \new_[17122]_  = ~\new_[27552]_  | ~\new_[19136]_  | ~\new_[23447]_ ;
  assign \new_[17123]_  = \new_[21725]_  | \new_[19137]_ ;
  assign \new_[17124]_  = \new_[20802]_  | \new_[19144]_ ;
  assign \new_[17125]_  = \new_[22205]_  | \new_[19208]_ ;
  assign \new_[17126]_  = ~\new_[27646]_  | ~\new_[19158]_  | ~\new_[22279]_ ;
  assign \new_[17127]_  = \new_[20835]_  | \new_[19151]_ ;
  assign \new_[17128]_  = \new_[20896]_  | \new_[19166]_ ;
  assign \new_[17129]_  = ~\new_[28632]_  | ~\new_[19168]_  | ~\new_[23343]_ ;
  assign \new_[17130]_  = ~\new_[29413]_  | ~\new_[19170]_  | ~\new_[23839]_ ;
  assign \new_[17131]_  = \new_[22420]_  | \new_[19218]_ ;
  assign \new_[17132]_  = ~\new_[27694]_  | ~\new_[19175]_  | ~\new_[23735]_ ;
  assign \new_[17133]_  = \new_[20888]_  | \new_[19179]_ ;
  assign \new_[17134]_  = \new_[20927]_  | \new_[19183]_ ;
  assign \new_[17135]_  = \new_[21964]_  | \new_[19169]_ ;
  assign \new_[17136]_  = \new_[22433]_  | \new_[19214]_ ;
  assign \new_[17137]_  = ~\new_[27620]_  | ~\new_[19147]_  | ~\new_[23507]_ ;
  assign \new_[17138]_  = ~\new_[23350]_  & (~\new_[20208]_  | ~\new_[24162]_ );
  assign \new_[17139]_  = ~\new_[26880]_  & (~\new_[20256]_  | ~\new_[26811]_ );
  assign \new_[17140]_  = ~\new_[20118]_  | (~\new_[20253]_  & ~\new_[30663]_ );
  assign \new_[17141]_  = ~\new_[23406]_  & (~\new_[20247]_  | ~\new_[24290]_ );
  assign \new_[17142]_  = ~\new_[23746]_  & (~\new_[20222]_  | ~\new_[24213]_ );
  assign \new_[17143]_  = ~\new_[23452]_  & (~\new_[20218]_  | ~\new_[24450]_ );
  assign \new_[17144]_  = ~\new_[20145]_  | (~\new_[20219]_  & ~\new_[30249]_ );
  assign \new_[17145]_  = ~\new_[23582]_  & (~\new_[20220]_  | ~\new_[23078]_ );
  assign \new_[17146]_  = ~\new_[22280]_  & (~\new_[20223]_  | ~\new_[27914]_ );
  assign \new_[17147]_  = ~\new_[23559]_  & (~\new_[20248]_  | ~\new_[26220]_ );
  assign \new_[17148]_  = ~\new_[24827]_  & (~\new_[20210]_  | ~\new_[26283]_ );
  assign \new_[17149]_  = ~\new_[20073]_  | (~\new_[20226]_  & ~\new_[30319]_ );
  assign \new_[17150]_  = ~\new_[23683]_  & (~\new_[20230]_  | ~\new_[24081]_ );
  assign \new_[17151]_  = ~\new_[20084]_  | (~\new_[20236]_  & ~\new_[30069]_ );
  assign \new_[17152]_  = ~\new_[20085]_  | (~\new_[20239]_  & ~\new_[30008]_ );
  assign \new_[17153]_  = ~\new_[25062]_  & (~\new_[20244]_  | ~\new_[27425]_ );
  assign \new_[17154]_  = ~\new_[23720]_  & (~\new_[20262]_  | ~\new_[22926]_ );
  assign \new_[17155]_  = ~\new_[23751]_  & (~\new_[20254]_  | ~\new_[28133]_ );
  assign \new_[17156]_  = ~\new_[23869]_  & (~\new_[20212]_  | ~\new_[23120]_ );
  assign \new_[17157]_  = ~\new_[21308]_  & (~\new_[20107]_  | ~\new_[21180]_ );
  assign \new_[17158]_  = ~\new_[30693]_  | ~\new_[18719]_  | ~\new_[26022]_ ;
  assign \new_[17159]_  = ~\new_[30015]_  | ~\new_[18710]_  | ~\new_[24814]_ ;
  assign \new_[17160]_  = ~\new_[28894]_  | ~\new_[18711]_  | ~\new_[23737]_ ;
  assign \new_[17161]_  = ~\new_[28918]_  | ~\new_[18713]_  | ~\new_[23414]_ ;
  assign \new_[17162]_  = ~\new_[30242]_  | ~\new_[18712]_  | ~\new_[23448]_ ;
  assign \new_[17163]_  = ~\new_[20117]_  | (~\new_[20235]_  & ~\new_[30270]_ );
  assign \new_[17164]_  = ~\new_[28818]_  | ~\new_[18714]_  | ~\new_[24942]_ ;
  assign \new_[17165]_  = ~\new_[30599]_  | ~\new_[18715]_  | ~\new_[24961]_ ;
  assign \new_[17166]_  = ~\new_[29410]_  | ~\new_[18722]_  | ~\new_[23732]_ ;
  assign \new_[17167]_  = ~\new_[28595]_  | ~\new_[18718]_  | ~\new_[23698]_ ;
  assign \new_[17168]_  = ~\new_[29893]_  | ~\new_[18720]_  | ~\new_[23662]_ ;
  assign \new_[17169]_  = ~\new_[29583]_  | ~\new_[18716]_  | ~\new_[25253]_ ;
  assign \new_[17170]_  = ~\new_[28675]_  | ~\new_[18723]_  | ~\new_[23727]_ ;
  assign \new_[17171]_  = ~\new_[29681]_  | ~\new_[18717]_  | ~\new_[23628]_ ;
  assign \new_[17172]_  = ~\new_[27997]_  | ~\new_[18724]_  | ~\new_[25469]_ ;
  assign \new_[17173]_  = ~\new_[29825]_  | ~\new_[18721]_  | ~\new_[25131]_ ;
  assign \new_[17174]_  = ~\new_[30233]_  | ~\new_[18727]_  | ~\new_[26522]_ ;
  assign \new_[17175]_  = ~\new_[19338]_  | ~\new_[26374]_ ;
  assign \new_[17176]_  = ~\new_[19337]_  | ~\new_[26292]_ ;
  assign \new_[17177]_  = ~\new_[19336]_  | ~\new_[27926]_ ;
  assign \new_[17178]_  = ~\new_[19331]_  | ~\new_[26347]_ ;
  assign \new_[17179]_  = ~\new_[19339]_  | ~\new_[26443]_ ;
  assign \new_[17180]_  = ~\new_[19329]_  | ~\new_[26309]_ ;
  assign \new_[17181]_  = ~\new_[19334]_  | ~\new_[26395]_ ;
  assign \new_[17182]_  = ~\new_[19332]_  | ~\new_[27635]_ ;
  assign \new_[17183]_  = ~\new_[19316]_  | ~\new_[29401]_ ;
  assign \new_[17184]_  = ~\new_[19330]_  | ~\new_[26083]_ ;
  assign \new_[17185]_  = ~\new_[19315]_  | ~\new_[29701]_ ;
  assign \new_[17186]_  = ~\new_[19335]_  | ~\new_[27596]_ ;
  assign \new_[17187]_  = ~\new_[18003]_ ;
  assign \new_[17188]_  = ~\new_[18003]_ ;
  assign \new_[17189]_  = ~\new_[18003]_ ;
  assign \new_[17190]_  = ~\new_[18005]_ ;
  assign \new_[17191]_  = ~\new_[18005]_ ;
  assign \new_[17192]_  = ~\new_[18005]_ ;
  assign \new_[17193]_  = ~\new_[18006]_ ;
  assign \new_[17194]_  = ~\new_[18741]_ ;
  assign \new_[17195]_  = ~\new_[18741]_ ;
  assign \new_[17196]_  = ~\new_[18741]_ ;
  assign \new_[17197]_  = ~\new_[18742]_ ;
  assign \new_[17198]_  = ~\new_[18008]_ ;
  assign \new_[17199]_  = ~\new_[18009]_ ;
  assign \new_[17200]_  = ~\new_[18009]_ ;
  assign \new_[17201]_  = ~\new_[18009]_ ;
  assign \new_[17202]_  = ~\new_[18012]_ ;
  assign \new_[17203]_  = ~\new_[18012]_ ;
  assign \new_[17204]_  = ~\new_[18013]_ ;
  assign \new_[17205]_  = ~\new_[18013]_ ;
  assign \new_[17206]_  = ~\new_[28992]_  & (~\new_[20289]_  | ~\new_[23367]_ );
  assign \new_[17207]_  = ~\new_[18023]_ ;
  assign \new_[17208]_  = ~\new_[29217]_  & (~\new_[20317]_  | ~\new_[23435]_ );
  assign \new_[17209]_  = ~\new_[29695]_  | ~\new_[19306]_  | ~\new_[30061]_ ;
  assign \new_[17210]_  = ~\new_[18784]_ ;
  assign \new_[17211]_  = ~\new_[18032]_ ;
  assign \new_[17212]_  = ~\new_[18033]_ ;
  assign \new_[17213]_  = ~\new_[18034]_ ;
  assign \new_[17214]_  = ~\new_[18070]_ ;
  assign \new_[17215]_  = ~\new_[19569]_ ;
  assign \new_[17216]_  = ~\new_[19569]_ ;
  assign \new_[17217]_  = ~\new_[18801]_ ;
  assign \new_[17218]_  = ~\new_[17217]_ ;
  assign \new_[17219]_  = ~\new_[17217]_ ;
  assign \new_[17220]_  = ~\new_[18072]_ ;
  assign \new_[17221]_  = ~\new_[18072]_ ;
  assign \new_[17222]_  = ~\new_[18073]_ ;
  assign \new_[17223]_  = ~\new_[18076]_ ;
  assign \new_[17224]_  = ~\new_[18076]_ ;
  assign \new_[17225]_  = ~\new_[18080]_ ;
  assign \new_[17226]_  = ~\new_[18085]_ ;
  assign \new_[17227]_  = ~\new_[18818]_ ;
  assign \new_[17228]_  = ~\new_[28963]_  | ~\new_[19297]_  | ~\new_[30092]_ ;
  assign \new_[17229]_  = ~\new_[18091]_ ;
  assign \new_[17230]_  = ~\new_[29254]_  & (~\new_[20329]_  | ~\new_[23794]_ );
  assign \new_[17231]_  = ~\new_[24610]_  & ~\new_[19260]_ ;
  assign \new_[17232]_  = ~\new_[18092]_ ;
  assign \new_[17233]_  = ~\new_[18093]_ ;
  assign \new_[17234]_  = ~\new_[18093]_ ;
  assign \new_[17235]_  = ~\new_[18093]_ ;
  assign \new_[17236]_  = ~\new_[18094]_ ;
  assign \new_[17237]_  = ~\new_[18095]_ ;
  assign \new_[17238]_  = ~\new_[18096]_ ;
  assign \new_[17239]_  = ~\new_[18097]_ ;
  assign \new_[17240]_  = ~\new_[18097]_ ;
  assign \new_[17241]_  = ~\new_[18117]_ ;
  assign \new_[17242]_  = ~\new_[29541]_  & (~\new_[20337]_  | ~\new_[23644]_ );
  assign \new_[17243]_  = ~\new_[29229]_  & (~\new_[20347]_  | ~\new_[23709]_ );
  assign \new_[17244]_  = ~\new_[29101]_  & (~\new_[20344]_  | ~\new_[23724]_ );
  assign \new_[17245]_  = ~\new_[18124]_ ;
  assign \new_[17246]_  = ~\new_[18124]_ ;
  assign \new_[17247]_  = ~\new_[18124]_ ;
  assign \new_[17248]_  = ~\new_[18127]_ ;
  assign \new_[17249]_  = ~\new_[18129]_ ;
  assign \new_[17250]_  = ~\new_[29721]_  | ~\new_[19311]_  | ~\new_[29888]_ ;
  assign \new_[17251]_  = ~\new_[29115]_  & (~\new_[20349]_  | ~\new_[23795]_ );
  assign \new_[17252]_  = ~\new_[18135]_ ;
  assign \new_[17253]_  = \new_[18135]_ ;
  assign \new_[17254]_  = ~\new_[28183]_  | ~\new_[19287]_  | ~\new_[30337]_ ;
  assign \new_[17255]_  = ~\new_[18138]_ ;
  assign \new_[17256]_  = ~\new_[18138]_ ;
  assign \new_[17257]_  = ~\new_[18138]_ ;
  assign \new_[17258]_  = ~\new_[29058]_  & (~\new_[20351]_  | ~\new_[23466]_ );
  assign \new_[17259]_  = ~\new_[29167]_  & (~\new_[20297]_  | ~\new_[23635]_ );
  assign \new_[17260]_  = ~\new_[18875]_ ;
  assign \new_[17261]_  = ~\new_[18141]_ ;
  assign \new_[17262]_  = ~\new_[18148]_ ;
  assign \new_[17263]_  = ~\new_[18148]_ ;
  assign \new_[17264]_  = ~\new_[18150]_ ;
  assign \new_[17265]_  = ~\new_[18150]_ ;
  assign \new_[17266]_  = ~\new_[18150]_ ;
  assign \new_[17267]_  = ~\new_[18151]_ ;
  assign \new_[17268]_  = ~\new_[18153]_ ;
  assign \new_[17269]_  = ~\new_[18154]_ ;
  assign \new_[17270]_  = ~\new_[18158]_ ;
  assign \new_[17271]_  = ~\new_[18158]_ ;
  assign \new_[17272]_  = ~\new_[18166]_ ;
  assign \new_[17273]_  = ~\new_[18176]_ ;
  assign \new_[17274]_  = ~\new_[18178]_ ;
  assign \new_[17275]_  = ~\new_[18179]_ ;
  assign \new_[17276]_  = ~\new_[19631]_ ;
  assign \new_[17277]_  = \new_[18192]_ ;
  assign \new_[17278]_  = ~\new_[18194]_ ;
  assign \new_[17279]_  = ~\new_[18194]_ ;
  assign \new_[17280]_  = ~\new_[18194]_ ;
  assign \new_[17281]_  = ~\new_[29103]_  | ~\new_[19290]_  | ~\new_[29762]_ ;
  assign \new_[17282]_  = ~\new_[30573]_  | ~\new_[29251]_  | ~\new_[20942]_  | ~\new_[30767]_ ;
  assign \new_[17283]_  = ~\new_[30147]_  | ~\new_[28280]_  | ~\new_[19244]_  | ~\new_[29571]_ ;
  assign \new_[17284]_  = ~\new_[30563]_  | ~\new_[28762]_  | ~\new_[19269]_  | ~\new_[30578]_ ;
  assign \new_[17285]_  = ~\new_[28905]_  | ~\new_[28073]_  | ~\new_[19246]_  | ~\new_[28285]_ ;
  assign \new_[17286]_  = ~\new_[30707]_  | ~\new_[28535]_  | ~\new_[20731]_  | ~\new_[29817]_ ;
  assign \new_[17287]_  = ~\new_[30125]_  | ~\new_[28023]_  | ~\new_[19245]_  | ~\new_[29787]_ ;
  assign \new_[17288]_  = ~\new_[30814]_  | ~\new_[28888]_  | ~\new_[21794]_  | ~\new_[30613]_ ;
  assign \new_[17289]_  = ~\new_[23350]_  & (~\new_[20395]_  | ~\new_[22463]_ );
  assign \new_[17290]_  = ~\new_[18228]_ ;
  assign \new_[17291]_  = ~\new_[21163]_  & (~\new_[20407]_  | ~\new_[23898]_ );
  assign \new_[17292]_  = ~\new_[23378]_  & (~\new_[20403]_  | ~\new_[22513]_ );
  assign \new_[17293]_  = ~\new_[26399]_  | ~\new_[18552]_ ;
  assign \new_[17294]_  = ~\new_[21155]_  | ~\new_[24442]_  | ~\new_[26267]_  | ~\new_[29421]_ ;
  assign \new_[17295]_  = ~\new_[21214]_  | ~\new_[22870]_  | ~\new_[26292]_  | ~\new_[28894]_ ;
  assign \new_[17296]_  = ~\new_[21140]_  | ~\new_[23004]_  | ~\new_[27926]_  | ~\new_[30229]_ ;
  assign \new_[17297]_  = ~\new_[18237]_ ;
  assign \new_[17298]_  = ~\new_[21157]_  | ~\new_[24617]_  | ~\new_[27848]_  | ~\new_[29851]_ ;
  assign \new_[17299]_  = ~\new_[23418]_  & (~\new_[20397]_  | ~\new_[22473]_ );
  assign \new_[17300]_  = \new_[6095]_  ? \new_[29768]_  : \new_[19759]_ ;
  assign \new_[17301]_  = ~\new_[21154]_  | ~\new_[22999]_  | ~\new_[26083]_  | ~\new_[28918]_ ;
  assign \new_[17302]_  = ~\new_[21176]_  | ~\new_[23140]_  | ~\new_[27736]_  | ~\new_[30222]_ ;
  assign \new_[17303]_  = ~\new_[18247]_ ;
  assign \new_[17304]_  = ~\new_[21174]_  | ~\new_[21506]_  | ~\new_[26239]_  | ~\new_[28595]_ ;
  assign \new_[17305]_  = ~\new_[23452]_  & (~\new_[20396]_  | ~\new_[22474]_ );
  assign \new_[17306]_  = ~\new_[30573]_  | ~\new_[21520]_  | ~\new_[23592]_  | ~\new_[24401]_ ;
  assign \new_[17307]_  = ~\new_[18253]_ ;
  assign \new_[17308]_  = ~\new_[23406]_  & (~\new_[20394]_  | ~\new_[22468]_ );
  assign \new_[17309]_  = ~\new_[24412]_  | ~\new_[18595]_ ;
  assign \new_[17310]_  = ~\new_[30204]_  & (~\new_[20335]_  | ~\new_[22196]_ );
  assign \new_[17311]_  = ~\new_[18256]_ ;
  assign \new_[17312]_  = ~\new_[18256]_ ;
  assign \new_[17313]_  = ~\new_[18256]_ ;
  assign \new_[17314]_  = ~\new_[22246]_  & (~\new_[20398]_  | ~\new_[22482]_ );
  assign \new_[17315]_  = ~\new_[21199]_  | ~\new_[26402]_  | ~\new_[27593]_  | ~\new_[29869]_ ;
  assign \new_[17316]_  = ~\new_[21178]_  | ~\new_[23060]_  | ~\new_[26309]_  | ~\new_[29020]_ ;
  assign \new_[17317]_  = ~\new_[21149]_  | ~\new_[24455]_  | ~\new_[24782]_  | ~\new_[29868]_ ;
  assign \new_[17318]_  = ~\new_[23549]_  & (~\new_[20404]_  | ~\new_[22516]_ );
  assign \new_[17319]_  = ~\new_[21233]_  | ~\new_[21823]_  | ~\new_[27635]_  | ~\new_[28818]_ ;
  assign \new_[17320]_  = ~\new_[21191]_  | ~\new_[27605]_  | ~\new_[26940]_  | ~\new_[30525]_ ;
  assign \new_[17321]_  = ~\new_[23582]_  & (~\new_[20400]_  | ~\new_[22495]_ );
  assign \new_[17322]_  = ~\new_[22440]_  & (~\new_[20402]_  | ~\new_[23919]_ );
  assign \new_[17323]_  = ~\new_[21196]_  | ~\new_[24310]_  | ~\new_[26300]_  | ~\new_[28836]_ ;
  assign \new_[17324]_  = ~\new_[27802]_  | ~\new_[19305]_  | ~\new_[29912]_ ;
  assign \new_[17325]_  = ~\new_[18274]_ ;
  assign \new_[17326]_  = ~\new_[18279]_ ;
  assign \new_[17327]_  = ~\new_[18279]_ ;
  assign \new_[17328]_  = ~\new_[30814]_  | ~\new_[21547]_  | ~\new_[24819]_  | ~\new_[26244]_ ;
  assign \new_[17329]_  = ~\new_[21177]_  | ~\new_[24257]_  | ~\new_[26360]_  | ~\new_[29410]_ ;
  assign \new_[17330]_  = ~\new_[18282]_ ;
  assign \new_[17331]_  = ~\new_[28073]_  | ~\new_[19302]_  | ~\new_[29974]_ ;
  assign \new_[17332]_  = ~\new_[18287]_ ;
  assign \new_[17333]_  = ~\new_[23683]_  & (~\new_[20401]_  | ~\new_[22506]_ );
  assign \new_[17334]_  = ~\new_[23746]_  & (~\new_[20399]_  | ~\new_[22514]_ );
  assign \new_[17335]_  = ~\new_[21119]_  | ~\new_[22861]_  | ~\new_[26443]_  | ~\new_[29623]_ ;
  assign \new_[17336]_  = ~\new_[21226]_  | ~\new_[22998]_  | ~\new_[27596]_  | ~\new_[29583]_ ;
  assign \new_[17337]_  = ~\new_[18296]_ ;
  assign \new_[17338]_  = ~\new_[18301]_ ;
  assign \new_[17339]_  = ~\new_[28535]_  | ~\new_[19300]_  | ~\new_[29386]_ ;
  assign \new_[17340]_  = ~\new_[23744]_  & (~\new_[20406]_  | ~\new_[22521]_ );
  assign \new_[17341]_  = ~\new_[18308]_ ;
  assign \new_[17342]_  = ~\new_[18308]_ ;
  assign \new_[17343]_  = ~\new_[22204]_  & (~\new_[20405]_  | ~\new_[24685]_ );
  assign \new_[17344]_  = ~\new_[21253]_  | ~\new_[21538]_  | ~\new_[27561]_  | ~\new_[29987]_ ;
  assign \new_[17345]_  = ~\new_[23869]_  & (~\new_[20408]_  | ~\new_[22522]_ );
  assign \new_[17346]_  = ~\new_[30552]_  | ~\new_[19293]_  | ~\new_[30617]_ ;
  assign \new_[17347]_  = ~\new_[22455]_  | ~\new_[26215]_  | ~\new_[26333]_  | ~\new_[28278]_ ;
  assign \new_[17348]_  = ~\new_[21236]_  | ~\new_[20523]_  | ~\new_[27594]_  | ~\new_[29151]_ ;
  assign \new_[17349]_  = ~\new_[20302]_  & (~\new_[19644]_  | ~\new_[29350]_ );
  assign \new_[17350]_  = \new_[6183]_  ? \new_[30269]_  : \new_[19688]_ ;
  assign \new_[17351]_  = ~\new_[19271]_  | ~\new_[30105]_ ;
  assign \new_[17352]_  = ~\new_[19270]_  | ~\new_[30009]_ ;
  assign \new_[17353]_  = ~\new_[29227]_  | ~\new_[5902]_ ;
  assign \new_[17354]_  = ~\new_[19265]_  & (~\new_[29268]_  | ~\new_[30080]_ );
  assign \new_[17355]_  = ~\new_[19262]_  & (~\new_[30030]_  | ~\new_[29839]_ );
  assign \new_[17356]_  = ~\new_[19268]_  & (~\new_[28924]_  | ~\new_[30043]_ );
  assign \new_[17357]_  = ~\new_[19251]_  & (~\new_[28872]_  | ~\new_[30040]_ );
  assign \new_[17358]_  = ~\new_[19255]_  & (~\new_[30057]_  | ~\new_[29899]_ );
  assign \new_[17359]_  = ~\new_[19258]_  & (~\new_[28883]_  | ~\new_[30203]_ );
  assign \new_[17360]_  = ~\new_[19256]_  & (~\new_[28939]_  | ~\new_[29833]_ );
  assign \new_[17361]_  = ~\new_[19261]_  & (~\new_[28887]_  | ~\new_[30292]_ );
  assign \new_[17362]_  = ~\new_[19278]_  & (~\new_[29248]_  | ~\new_[30307]_ );
  assign \new_[17363]_  = ~\new_[20355]_  | ~\new_[19378]_ ;
  assign \new_[17364]_  = ~\new_[23692]_  & (~\new_[19853]_  | ~\new_[28964]_ );
  assign \new_[17365]_  = ~\new_[27548]_  | ~\new_[18545]_ ;
  assign \new_[17366]_  = ~\new_[19373]_  | ~\new_[19378]_ ;
  assign \new_[17367]_  = ~\new_[19373]_  & ~\new_[19378]_ ;
  assign \new_[17368]_  = ~\new_[30336]_  & (~\new_[20473]_  | ~\new_[29305]_ );
  assign \new_[17369]_  = ~\new_[30326]_  & (~\new_[20490]_  | ~\new_[29461]_ );
  assign \new_[17370]_  = ~\new_[19366]_  | ~\new_[30229]_ ;
  assign \new_[17371]_  = ~\new_[19355]_  | ~\new_[29020]_ ;
  assign \new_[17372]_  = ~\new_[19375]_  | ~\new_[29851]_ ;
  assign \new_[17373]_  = ~\new_[5973]_  | ~\new_[30237]_  | ~\new_[28718]_ ;
  assign n8849 = m6_s0_cyc_o_reg;
  assign n8414 = m0_s0_cyc_o_reg;
  assign n8589 = m1_s0_cyc_o_reg;
  assign \new_[17377]_  = ~\new_[6001]_  | ~\new_[28288]_  | ~\new_[27778]_ ;
  assign \new_[17378]_  = ~\new_[5919]_  | ~\new_[28910]_  | ~\new_[29300]_ ;
  assign \new_[17379]_  = ~\new_[26794]_  | ~\new_[18508]_ ;
  assign \new_[17380]_  = ~\new_[23058]_  & (~\new_[19473]_  | ~\new_[30582]_ );
  assign \new_[17381]_  = ~\new_[24387]_  & (~\new_[19475]_  | ~\new_[29159]_ );
  assign \new_[17382]_  = ~\new_[23526]_  & (~\new_[19855]_  | ~\new_[29904]_ );
  assign \new_[17383]_  = ~\new_[30651]_  & (~\new_[21807]_  | ~\new_[19719]_ );
  assign \new_[17384]_  = ~\new_[23566]_  & (~\new_[19878]_  | ~\new_[29404]_ );
  assign \new_[17385]_  = ~\new_[20489]_  & (~\new_[19488]_  | ~\new_[30727]_ );
  assign \new_[17386]_  = ~\new_[21545]_  & (~\new_[19497]_  | ~\new_[30764]_ );
  assign \new_[17387]_  = ~\new_[26224]_  & (~\new_[19490]_  | ~\new_[28069]_ );
  assign \new_[17388]_  = ~\new_[29479]_  & (~\new_[19472]_  | ~\new_[30015]_ );
  assign \new_[17389]_  = ~\new_[27686]_  & (~\new_[19474]_  | ~\new_[30229]_ );
  assign \new_[17390]_  = ~\new_[27958]_  & (~\new_[19476]_  | ~\new_[27787]_ );
  assign \new_[17391]_  = ~\new_[24324]_  & (~\new_[19478]_  | ~\new_[26655]_ );
  assign \new_[17392]_  = ~\new_[24372]_  & (~\new_[19477]_  | ~\new_[28039]_ );
  assign \new_[17393]_  = ~\new_[24563]_  & (~\new_[19485]_  | ~\new_[29064]_ );
  assign \new_[17394]_  = ~\new_[26388]_  & (~\new_[19486]_  | ~\new_[29987]_ );
  assign \new_[17395]_  = ~\new_[26380]_  & (~\new_[19487]_  | ~\new_[29537]_ );
  assign \new_[17396]_  = ~\new_[24929]_  & (~\new_[19496]_  | ~\new_[30735]_ );
  assign \new_[17397]_  = ~\new_[27650]_  & (~\new_[19505]_  | ~\new_[30152]_ );
  assign \new_[17398]_  = ~\new_[26826]_  & (~\new_[19508]_  | ~\new_[30213]_ );
  assign \new_[17399]_  = ~\new_[28486]_  & (~\new_[19509]_  | ~\new_[30786]_ );
  assign \new_[17400]_  = ~\new_[28296]_  & (~\new_[19507]_  | ~\new_[30444]_ );
  assign \new_[17401]_  = ~\new_[29944]_  & (~\new_[19494]_  | ~\new_[30363]_ );
  assign \new_[17402]_  = ~\new_[20336]_  & (~\new_[19593]_  | ~\new_[29202]_ );
  assign \new_[17403]_  = ~\new_[29195]_  | ~\new_[5895]_ ;
  assign \new_[17404]_  = ~\new_[29663]_  | ~\new_[6074]_ ;
  assign \new_[17405]_  = ~\new_[28833]_  | ~\new_[5897]_ ;
  assign \new_[17406]_  = ~\new_[29578]_  | ~\new_[5903]_ ;
  assign \new_[17407]_  = ~\new_[29195]_  | ~\new_[6036]_ ;
  assign \new_[17408]_  = ~\new_[28668]_  & (~\new_[19510]_  | ~\new_[30544]_ );
  assign \new_[17409]_  = ~\new_[29465]_  | ~\new_[5898]_ ;
  assign \new_[17410]_  = ~\new_[29068]_  | ~\new_[6075]_ ;
  assign \new_[17411]_  = ~\new_[29056]_  | ~\new_[5906]_ ;
  assign \new_[17412]_  = ~\new_[26653]_  | ~\new_[18606]_ ;
  assign \new_[17413]_  = ~\new_[29394]_  | ~\new_[5896]_ ;
  assign \new_[17414]_  = ~\new_[29068]_  | ~\new_[5905]_ ;
  assign \new_[17415]_  = ~\new_[26331]_  & (~\new_[19469]_  | ~\new_[30437]_ );
  assign \new_[17416]_  = ~\new_[29056]_  | ~\new_[6083]_ ;
  assign \new_[17417]_  = ~\new_[26324]_  | ~\new_[18573]_ ;
  assign \new_[17418]_  = ~\new_[29663]_  | ~\new_[5904]_ ;
  assign \new_[17419]_  = ~\new_[19007]_  | ~\new_[6274]_ ;
  assign \new_[17420]_  = ~\new_[30185]_  & (~\new_[20907]_  | ~\new_[19692]_ );
  assign \new_[17421]_  = \new_[6007]_  ? \new_[30724]_  : \new_[19504]_ ;
  assign \new_[17422]_  = ~\new_[18501]_  | ~\new_[30104]_ ;
  assign \new_[17423]_  = ~\new_[18518]_  | ~\new_[30111]_ ;
  assign \new_[17424]_  = ~\new_[18531]_  | ~\new_[30318]_ ;
  assign \new_[17425]_  = ~\new_[18524]_  | ~\new_[29780]_ ;
  assign \new_[17426]_  = ~\new_[18570]_  | ~\new_[30005]_ ;
  assign \new_[17427]_  = ~\new_[18598]_  | ~\new_[30086]_ ;
  assign \new_[17428]_  = ~\new_[18588]_  | ~\new_[30178]_ ;
  assign \new_[17429]_  = ~\new_[18526]_  | ~\new_[30180]_ ;
  assign \new_[17430]_  = ~\new_[18626]_  | ~\new_[30105]_ ;
  assign \new_[17431]_  = ~\new_[18609]_  | ~\new_[30089]_ ;
  assign \new_[17432]_  = ~\new_[18608]_  | ~\new_[30280]_ ;
  assign \new_[17433]_  = ~\new_[18628]_  | ~\new_[30123]_ ;
  assign \new_[17434]_  = ~\new_[30598]_  & (~\new_[19534]_  | ~\new_[28127]_ );
  assign \new_[17435]_  = ~\new_[29853]_  & (~\new_[21932]_  | ~\new_[19538]_ );
  assign \new_[17436]_  = ~\new_[30164]_  | (~\new_[19996]_  & ~\new_[20584]_ );
  assign \new_[17437]_  = ~\new_[26948]_  & (~\new_[19512]_  | ~\new_[30296]_ );
  assign \new_[17438]_  = ~\new_[29855]_  & (~\new_[20820]_  | ~\new_[19824]_ );
  assign \new_[17439]_  = ~\new_[18516]_  & ~\new_[29027]_ ;
  assign \new_[17440]_  = ~\new_[30215]_  | (~\new_[20752]_  & ~\new_[19668]_ );
  assign \new_[17441]_  = ~\new_[30508]_  | (~\new_[21670]_  & ~\new_[19669]_ );
  assign \new_[17442]_  = ~\new_[29100]_  & (~\new_[20897]_  | ~\new_[19830]_ );
  assign \new_[17443]_  = ~\new_[18529]_  & ~\new_[28994]_ ;
  assign \new_[17444]_  = ~\new_[29260]_  | (~\new_[20771]_  & ~\new_[19673]_ );
  assign \new_[17445]_  = ~\new_[28989]_  | (~\new_[20871]_  & ~\new_[19674]_ );
  assign \new_[17446]_  = ~\new_[30389]_  & (~\new_[20781]_  | ~\new_[19836]_ );
  assign \new_[17447]_  = ~\new_[18539]_  & ~\new_[29137]_ ;
  assign \new_[17448]_  = ~\new_[18540]_  | ~\new_[29251]_ ;
  assign \new_[17449]_  = ~\new_[29692]_  | (~\new_[20028]_  & ~\new_[19679]_ );
  assign \new_[17450]_  = ~\new_[25460]_  & (~\new_[19528]_  | ~\new_[30410]_ );
  assign \new_[17451]_  = ~\new_[28899]_  & (~\new_[20851]_  | ~\new_[19843]_ );
  assign \new_[17452]_  = ~\new_[18548]_  & ~\new_[30447]_ ;
  assign \new_[17453]_  = ~\new_[18610]_  | ~\new_[30011]_ ;
  assign \new_[17454]_  = ~\new_[29935]_  & (~\new_[21830]_  | ~\new_[19594]_ );
  assign \new_[17455]_  = ~\new_[30774]_  | (~\new_[20831]_  & ~\new_[19693]_ );
  assign \new_[17456]_  = ~\new_[28837]_  | (~\new_[20814]_  & ~\new_[19689]_ );
  assign \new_[17457]_  = \new_[18601]_  | \new_[29902]_ ;
  assign \new_[17458]_  = ~\new_[30044]_  & (~\new_[19582]_  | ~\new_[28508]_ );
  assign \new_[17459]_  = ~\new_[18561]_  | ~\new_[30697]_ ;
  assign \new_[17460]_  = ~\new_[28944]_  & (~\new_[23192]_  | ~\new_[19573]_ );
  assign \new_[17461]_  = ~\new_[30434]_  | (~\new_[22931]_  & ~\new_[19695]_ );
  assign \new_[17462]_  = ~\new_[18491]_  | ~\new_[30207]_ ;
  assign \new_[17463]_  = ~\new_[18571]_  & ~\new_[28996]_ ;
  assign \new_[17464]_  = ~\new_[30070]_  & (~\new_[23246]_  | ~\new_[19576]_ );
  assign \new_[17465]_  = ~\new_[30246]_  | (~\new_[20844]_  & ~\new_[19700]_ );
  assign \new_[17466]_  = ~\new_[29221]_  | (~\new_[20946]_  & ~\new_[19701]_ );
  assign \new_[17467]_  = ~\new_[30615]_  | (~\new_[20847]_  & ~\new_[19702]_ );
  assign \new_[17468]_  = ~\new_[29015]_  | (~\new_[20930]_  & ~\new_[19703]_ );
  assign \new_[17469]_  = ~\new_[18580]_  & ~\new_[28858]_ ;
  assign \new_[17470]_  = ~\new_[18591]_  | ~\new_[30213]_ ;
  assign \new_[17471]_  = ~\new_[18613]_  | ~\new_[30444]_ ;
  assign \new_[17472]_  = ~\new_[30526]_  & (~\new_[21789]_  | ~\new_[19579]_ );
  assign \new_[17473]_  = ~\new_[29139]_  | (~\new_[20062]_  & ~\new_[19704]_ );
  assign \new_[17474]_  = ~\new_[29171]_  | (~\new_[20061]_  & ~\new_[19707]_ );
  assign \new_[17475]_  = ~\new_[29573]_  & (~\new_[20859]_  | ~\new_[19862]_ );
  assign \new_[17476]_  = ~\new_[18637]_  & ~\new_[30742]_ ;
  assign \new_[17477]_  = ~\new_[29887]_  | (~\new_[20855]_  & ~\new_[19711]_ );
  assign \new_[17478]_  = ~\new_[29082]_  | (~\new_[20872]_  & ~\new_[19712]_ );
  assign \new_[17479]_  = ~\new_[29767]_  & (~\new_[20761]_  | ~\new_[19867]_ );
  assign \new_[17480]_  = ~\new_[18542]_  & ~\new_[29049]_ ;
  assign \new_[17481]_  = ~\new_[30348]_  & (~\new_[21882]_  | ~\new_[19591]_ );
  assign \new_[17482]_  = ~\new_[30538]_  | (~\new_[20857]_  & ~\new_[19720]_ );
  assign \new_[17483]_  = ~\new_[29648]_  & (~\new_[20784]_  | ~\new_[19870]_ );
  assign \new_[17484]_  = ~\new_[18612]_  & ~\new_[29325]_ ;
  assign \new_[17485]_  = ~\new_[30125]_  | (~\new_[20086]_  & ~\new_[20621]_ );
  assign \new_[17486]_  = ~\new_[30034]_  | (~\new_[20053]_  & ~\new_[19698]_ );
  assign \new_[17487]_  = ~\new_[30210]_  | (~\new_[20112]_  & ~\new_[21603]_ );
  assign \new_[17488]_  = ~\new_[29565]_  & (~\new_[20816]_  | ~\new_[19877]_ );
  assign \new_[17489]_  = ~\new_[28833]_  | ~\new_[6045]_ ;
  assign \new_[17490]_  = ~\new_[18599]_  & ~\new_[29282]_ ;
  assign \new_[17491]_  = ~\new_[30316]_  | (~\new_[20054]_  & ~\new_[19694]_ );
  assign \new_[17492]_  = ~\new_[29061]_  | (~\new_[20040]_  & ~\new_[19687]_ );
  assign \new_[17493]_  = ~\new_[30620]_  & (~\new_[24021]_  | ~\new_[19601]_ );
  assign \new_[17494]_  = ~\new_[29038]_  | (~\new_[20976]_  & ~\new_[19726]_ );
  assign \new_[17495]_  = ~\new_[29898]_  & (~\new_[20918]_  | ~\new_[19886]_ );
  assign \new_[17496]_  = ~\new_[18592]_  & ~\new_[29486]_ ;
  assign \new_[17497]_  = ~\new_[28007]_  | (~\new_[20973]_  & ~\new_[19731]_ );
  assign \new_[17498]_  = ~\new_[29701]_  | (~\new_[20010]_  & ~\new_[20625]_ );
  assign \new_[17499]_  = ~\new_[18617]_  & ~\new_[29030]_ ;
  assign \new_[17500]_  = ~\new_[30755]_  & (~\new_[23244]_  | ~\new_[19604]_ );
  assign \new_[17501]_  = ~\new_[18658]_  & ~\new_[25966]_ ;
  assign \new_[17502]_  = ~\new_[30723]_  | (~\new_[20734]_  & ~\new_[19735]_ );
  assign \new_[17503]_  = ~\new_[30309]_  & (~\new_[19620]_  | ~\new_[28411]_ );
  assign \new_[17504]_  = ~\new_[30225]_  & (~\new_[19616]_  | ~\new_[28276]_ );
  assign \new_[17505]_  = ~\new_[18629]_  & ~\new_[30100]_ ;
  assign \new_[17506]_  = ~\new_[18630]_  | ~\new_[29798]_ ;
  assign \new_[17507]_  = ~\new_[30003]_  & (~\new_[21659]_  | ~\new_[19645]_ );
  assign \new_[17508]_  = ~\new_[28850]_  | (~\new_[20998]_  & ~\new_[19755]_ );
  assign \new_[17509]_  = ~\new_[29119]_  & (~\new_[21987]_  | ~\new_[19909]_ );
  assign \new_[17510]_  = ~\new_[18506]_  & ~\new_[30230]_ ;
  assign \new_[17511]_  = ~\new_[18530]_  & ~\new_[29815]_ ;
  assign \new_[17512]_  = ~\new_[18604]_  & ~\new_[30115]_ ;
  assign \new_[17513]_  = ~\new_[18619]_  & ~\new_[30157]_ ;
  assign \new_[17514]_  = ~\new_[18651]_  | ~\new_[28049]_ ;
  assign \new_[17515]_  = ~\new_[18642]_  | ~\new_[28127]_ ;
  assign \new_[17516]_  = ~\new_[18643]_  | ~\new_[26305]_ ;
  assign \new_[17517]_  = \new_[18644]_  | \new_[26999]_ ;
  assign \new_[17518]_  = \new_[18648]_  | \new_[29468]_ ;
  assign \new_[17519]_  = \new_[18645]_  | \new_[28341]_ ;
  assign \new_[17520]_  = \new_[18641]_  | \new_[27994]_ ;
  assign \new_[17521]_  = ~\new_[18650]_  | ~\new_[26812]_ ;
  assign \new_[17522]_  = ~\new_[18649]_  | ~\new_[28411]_ ;
  assign \new_[17523]_  = \new_[18647]_  | \new_[29632]_ ;
  assign \new_[17524]_  = ~\new_[18646]_  | ~\new_[28276]_ ;
  assign \new_[17525]_  = \new_[18483]_  & \new_[29357]_ ;
  assign \new_[17526]_  = ~\new_[19612]_  | ~\new_[31334]_  | ~n8609;
  assign \new_[17527]_  = ~\new_[19554]_  | ~\new_[31222]_  | ~n8389;
  assign \new_[17528]_  = ~\new_[19632]_  | ~\new_[31522]_  | ~n8884;
  assign \new_[17529]_  = ~\new_[19572]_  | ~\new_[31298]_  | ~n8569;
  assign \new_[17530]_  = ~\new_[19584]_  | ~\new_[31251]_  | ~n8484;
  assign \new_[17531]_  = ~\new_[27925]_  & (~\new_[23477]_  | ~\new_[19823]_ );
  assign \new_[17532]_  = ~\new_[27940]_  & (~\new_[23393]_  | ~\new_[19829]_ );
  assign \new_[17533]_  = ~\new_[19565]_  | ~\new_[30795]_  | ~n8379;
  assign \new_[17534]_  = ~\new_[19539]_  | ~\new_[31387]_  | ~n8774;
  assign \new_[17535]_  = ~\new_[19608]_  | ~\new_[31224]_  | ~n8399;
  assign \new_[17536]_  = ~\new_[26925]_  & (~\new_[23429]_  | ~\new_[19835]_ );
  assign \new_[17537]_  = ~\new_[19577]_  | ~\new_[31359]_  | ~n8654;
  assign \new_[17538]_  = \new_[18490]_  & \new_[29104]_ ;
  assign \new_[17539]_  = ~\new_[19586]_  | ~\new_[31237]_  | ~n8424;
  assign \new_[17540]_  = ~\new_[19566]_  | ~\new_[31526]_  | ~n8904;
  assign \new_[17541]_  = ~\new_[19567]_  | ~\new_[31348]_  | ~n8629;
  assign \new_[17542]_  = ~\new_[19643]_  | ~\new_[31258]_  | ~n8494;
  assign \new_[17543]_  = ~\new_[19621]_  | ~\new_[30926]_  | ~n8384;
  assign \new_[17544]_  = ~\new_[26582]_  & (~\new_[23431]_  | ~\new_[19866]_ );
  assign \new_[17545]_  = ~\new_[19559]_  | ~\new_[31462]_  | ~n8819;
  assign \new_[17546]_  = ~\new_[26670]_  & (~\new_[23700]_  | ~\new_[19869]_ );
  assign \new_[17547]_  = ~\new_[27701]_  & (~\new_[23595]_  | ~\new_[19876]_ );
  assign \new_[17548]_  = ~\new_[19571]_  | ~\new_[31289]_  | ~n8539;
  assign \new_[17549]_  = ~\new_[19595]_  | ~\new_[31233]_  | ~n8409;
  assign \new_[17550]_  = ~\new_[19606]_  | ~\new_[31325]_  | ~n8599;
  assign \new_[17551]_  = ~\new_[19611]_  | ~\new_[30777]_  | ~n8359;
  assign \new_[17552]_  = ~\new_[19544]_  | ~\new_[30794]_  | ~n8374;
  assign \new_[17553]_  = ~\new_[19547]_  | ~\new_[30548]_  | ~n8339;
  assign \new_[17554]_  = ~\new_[26765]_  & (~\new_[23836]_  | ~\new_[19901]_ );
  assign \new_[17555]_  = ~\new_[19590]_  | ~\new_[31287]_  | ~n8529;
  assign \new_[17556]_  = ~\new_[19581]_  | ~\new_[31511]_  | ~n8849;
  assign \new_[17557]_  = ~\new_[19636]_  | ~\new_[31290]_  | ~n8544;
  assign \new_[17558]_  = ~\new_[20573]_  | ~\new_[31389]_  | ~n8779;
  assign \new_[17559]_  = ~\new_[20539]_  | ~\new_[31371]_  | ~n8709;
  assign \new_[17560]_  = ~\new_[20571]_  | ~\new_[30546]_  | ~n8334;
  assign \new_[17561]_  = ~\new_[20541]_  | ~\new_[31374]_  | ~n8724;
  assign \new_[17562]_  = ~\new_[20550]_  | ~\new_[31354]_  | ~n8644;
  assign \new_[17563]_  = ~\new_[20560]_  | ~\new_[31364]_  | ~n8674;
  assign \new_[17564]_  = ~\new_[20545]_  | ~\new_[31366]_  | ~n8684;
  assign \new_[17565]_  = ~\new_[30726]_  | (~\new_[20638]_  & ~\new_[23356]_ );
  assign \new_[17566]_  = ~\new_[30750]_  | (~\new_[20643]_  & ~\new_[22151]_ );
  assign \new_[17567]_  = ~\new_[30721]_  | (~\new_[20645]_  & ~\new_[21565]_ );
  assign \new_[17568]_  = ~\new_[29233]_  | (~\new_[20648]_  & ~\new_[22131]_ );
  assign \new_[17569]_  = ~\new_[30574]_  | (~\new_[20649]_  & ~\new_[24301]_ );
  assign \new_[17570]_  = ~\new_[30765]_  | (~\new_[20650]_  & ~\new_[21217]_ );
  assign \new_[17571]_  = ~\new_[30538]_  | (~\new_[20653]_  & ~\new_[23633]_ );
  assign \new_[17572]_  = ~\new_[30125]_  | (~\new_[20646]_  & ~\new_[22361]_ );
  assign \new_[17573]_  = ~\new_[30610]_  | (~\new_[20660]_  & ~\new_[21188]_ );
  assign \new_[17574]_  = ~\new_[30789]_  | (~\new_[20658]_  & ~\new_[23817]_ );
  assign \new_[17575]_  = ~\new_[30820]_  | (~\new_[20661]_  & ~\new_[23793]_ );
  assign n8594 = m2_s1_cyc_o_reg;
  assign n8689 = m7_s1_cyc_o_reg;
  assign n8404 = m2_s15_cyc_o_reg;
  assign n8759 = m4_s15_cyc_o_reg;
  assign n8909 = m7_s12_cyc_o_reg;
  assign n8694 = m7_s8_cyc_o_reg;
  assign \new_[17582]_  = ~\new_[24347]_  | ~\new_[19481]_ ;
  assign \new_[17583]_  = \new_[6203]_  ? \new_[30730]_  : \new_[20604]_ ;
  assign \new_[17584]_  = \new_[6041]_  ? \new_[30135]_  : \new_[20591]_ ;
  assign \new_[17585]_  = \new_[31143]_  ? \new_[30139]_  : \new_[20598]_ ;
  assign \new_[17586]_  = \new_[6200]_  ? \new_[29783]_  : \new_[20618]_ ;
  assign \new_[17587]_  = \new_[6214]_  ? \new_[29892]_  : \new_[20620]_ ;
  assign \new_[17588]_  = \new_[6213]_  ? \new_[29891]_  : \new_[20624]_ ;
  assign \new_[17589]_  = \new_[6082]_  ? \new_[29913]_  : \new_[20605]_ ;
  assign \new_[17590]_  = \new_[6183]_  ? \new_[30437]_  : \new_[20583]_ ;
  assign \new_[17591]_  = \new_[6095]_  ? \new_[30724]_  : \new_[20636]_ ;
  assign \new_[17592]_  = ~\new_[23108]_  & (~\new_[20540]_  | ~\new_[30416]_ );
  assign \new_[17593]_  = ~\new_[22115]_  & (~\new_[20563]_  | ~\new_[30647]_ );
  assign \new_[17594]_  = ~\new_[23648]_  & (~\new_[20564]_  | ~\new_[30695]_ );
  assign \new_[17595]_  = ~\new_[22200]_  & (~\new_[20556]_  | ~\new_[30555]_ );
  assign \new_[17596]_  = ~\new_[23775]_  & (~\new_[20569]_  | ~\new_[30752]_ );
  assign \new_[17597]_  = ~\new_[23576]_  & (~\new_[20559]_  | ~\new_[30782]_ );
  assign \new_[17598]_  = ~\new_[22446]_  & (~\new_[20581]_  | ~\new_[30630]_ );
  assign \new_[17599]_  = ~\new_[22343]_  & (~\new_[20553]_  | ~\new_[30719]_ );
  assign \new_[17600]_  = ~\new_[23861]_  & (~\new_[20579]_  | ~\new_[30799]_ );
  assign \new_[17601]_  = \new_[19763]_  | \new_[29992]_ ;
  assign \new_[17602]_  = \new_[19826]_  | \new_[30245]_ ;
  assign \new_[17603]_  = ~\new_[19765]_  & ~\new_[23375]_ ;
  assign \new_[17604]_  = \new_[19766]_  | \new_[29826]_ ;
  assign \new_[17605]_  = ~\new_[19769]_  & ~\new_[21136]_ ;
  assign \new_[17606]_  = ~\new_[19803]_  & ~\new_[22307]_ ;
  assign \new_[17607]_  = \new_[19832]_  | \new_[29908]_ ;
  assign \new_[17608]_  = ~\new_[19774]_  & ~\new_[21148]_ ;
  assign \new_[17609]_  = \new_[19775]_  | \new_[29848]_ ;
  assign \new_[17610]_  = \new_[19806]_  | \new_[30788]_ ;
  assign \new_[17611]_  = ~\new_[19776]_  & ~\new_[22149]_ ;
  assign \new_[17612]_  = \new_[19838]_  | \new_[29765]_ ;
  assign \new_[17613]_  = ~\new_[19779]_  & ~\new_[21164]_ ;
  assign \new_[17614]_  = \new_[19780]_  | \new_[30236]_ ;
  assign \new_[17615]_  = ~\new_[19781]_  & ~\new_[23458]_ ;
  assign \new_[17616]_  = \new_[19899]_  | \new_[30268]_ ;
  assign \new_[17617]_  = ~\new_[19794]_  & ~\new_[22264]_ ;
  assign \new_[17618]_  = ~\new_[19783]_  & ~\new_[23485]_ ;
  assign \new_[17619]_  = \new_[19771]_  | \new_[30733]_ ;
  assign \new_[17620]_  = ~\new_[19805]_  & ~\new_[22314]_ ;
  assign \new_[17621]_  = \new_[19856]_  | \new_[29865]_ ;
  assign \new_[17622]_  = \new_[19785]_  | \new_[29968]_ ;
  assign \new_[17623]_  = ~\new_[19789]_  & ~\new_[23544]_ ;
  assign \new_[17624]_  = \new_[19790]_  | \new_[30328]_ ;
  assign \new_[17625]_  = ~\new_[19792]_  & ~\new_[23555]_ ;
  assign \new_[17626]_  = \new_[19793]_  | \new_[30718]_ ;
  assign \new_[17627]_  = \new_[19871]_  | \new_[29994]_ ;
  assign \new_[17628]_  = ~\new_[19784]_  & ~\new_[21183]_ ;
  assign \new_[17629]_  = \new_[19787]_  | \new_[30251]_ ;
  assign \new_[17630]_  = ~\new_[19770]_  & ~\new_[22263]_ ;
  assign \new_[17631]_  = \new_[19863]_  | \new_[29914]_ ;
  assign \new_[17632]_  = ~\new_[19798]_  & ~\new_[21229]_ ;
  assign \new_[17633]_  = \new_[19807]_  | \new_[30308]_ ;
  assign \new_[17634]_  = ~\new_[19799]_  & ~\new_[23615]_ ;
  assign \new_[17635]_  = \new_[19860]_  | \new_[30304]_ ;
  assign \new_[17636]_  = ~\new_[19801]_  & ~\new_[22295]_ ;
  assign \new_[17637]_  = ~\new_[19800]_  & ~\new_[22456]_ ;
  assign \new_[17638]_  = \new_[19804]_  | \new_[29290]_ ;
  assign \new_[17639]_  = \new_[19828]_  | \new_[30267]_ ;
  assign \new_[17640]_  = ~\new_[19772]_  & ~\new_[23786]_ ;
  assign \new_[17641]_  = \new_[19897]_  | \new_[30024]_ ;
  assign \new_[17642]_  = \new_[19802]_  | \new_[28999]_ ;
  assign \new_[17643]_  = \new_[19814]_  | \new_[30652]_ ;
  assign \new_[17644]_  = \new_[19767]_  | \new_[30121]_ ;
  assign \new_[17645]_  = \new_[19810]_  | \new_[30502]_ ;
  assign \new_[17646]_  = \new_[19891]_  | \new_[29772]_ ;
  assign \new_[17647]_  = ~\new_[19811]_  & ~\new_[23680]_ ;
  assign \new_[17648]_  = \new_[19813]_  | \new_[30737]_ ;
  assign \new_[17649]_  = \new_[19900]_  | \new_[30277]_ ;
  assign \new_[17650]_  = \new_[19904]_  | \new_[30208]_ ;
  assign \new_[17651]_  = ~\new_[19816]_  & ~\new_[23866]_ ;
  assign \new_[17652]_  = \new_[19872]_  | \new_[30062]_ ;
  assign \new_[17653]_  = \new_[19817]_  | \new_[30706]_ ;
  assign \new_[17654]_  = ~\new_[22363]_  & (~\new_[20875]_  | ~\new_[22952]_ );
  assign \new_[17655]_  = ~\new_[28643]_  | (~\new_[20919]_  & ~\new_[30265]_ );
  assign \new_[17656]_  = ~\new_[26841]_  & (~\new_[20983]_  | ~\new_[29794]_ );
  assign \new_[17657]_  = \new_[19921]_  | \new_[30145]_ ;
  assign \new_[17658]_  = \new_[25152]_  & \new_[19649]_ ;
  assign \new_[17659]_  = ~\new_[25386]_  & (~\new_[20824]_  | ~\new_[29886]_ );
  assign \new_[17660]_  = \new_[22520]_  & \new_[19656]_ ;
  assign \new_[17661]_  = \new_[19911]_  | \new_[26208]_ ;
  assign \new_[17662]_  = ~s9_rty_i | ~\new_[19559]_  | ~\new_[29706]_ ;
  assign \new_[17663]_  = \new_[22485]_  & \new_[19650]_ ;
  assign \new_[17664]_  = \new_[19920]_  | \new_[28380]_ ;
  assign \new_[17665]_  = ~\new_[27549]_  & (~\new_[20748]_  | ~\new_[30111]_ );
  assign \new_[17666]_  = ~\new_[28532]_  | (~\new_[20937]_  & ~\new_[29909]_ );
  assign \new_[17667]_  = ~\new_[28532]_  | ~\new_[19895]_  | ~\new_[21232]_ ;
  assign \new_[17668]_  = \new_[19924]_  | \new_[29907]_ ;
  assign \new_[17669]_  = ~\new_[19551]_  | ~\new_[26322]_ ;
  assign \new_[17670]_  = ~\new_[27518]_  & (~\new_[20902]_  | ~\new_[29969]_ );
  assign \new_[17671]_  = ~\new_[26391]_  & (~\new_[20757]_  | ~\new_[29003]_ );
  assign \new_[17672]_  = \new_[19974]_  | \new_[26391]_ ;
  assign \new_[17673]_  = ~\new_[19549]_  | ~\new_[24745]_ ;
  assign \new_[17674]_  = ~\new_[23924]_  & (~\new_[20782]_  | ~\new_[28878]_ );
  assign \new_[17675]_  = \new_[19912]_  | \new_[27962]_ ;
  assign \new_[17676]_  = ~\new_[27918]_  & (~\new_[20889]_  | ~\new_[30318]_ );
  assign \new_[17677]_  = ~\new_[27679]_  & (~\new_[20768]_  | ~\new_[29061]_ );
  assign \new_[17678]_  = \new_[19928]_  | \new_[29810]_ ;
  assign \new_[17679]_  = ~\new_[26607]_  | ~\new_[19850]_  | ~\new_[24912]_ ;
  assign \new_[17680]_  = ~\new_[24761]_  & (~\new_[20863]_  | ~\new_[28866]_ );
  assign \new_[17681]_  = ~\new_[27978]_  & (~\new_[20773]_  | ~\new_[28989]_ );
  assign \new_[17682]_  = ~\new_[26531]_  & (~\new_[20858]_  | ~\new_[29192]_ );
  assign \new_[17683]_  = \new_[19969]_  | \new_[26531]_ ;
  assign \new_[17684]_  = ~\new_[26597]_  & (~\new_[20778]_  | ~\new_[27787]_ );
  assign \new_[17685]_  = ~\new_[28587]_  | (~\new_[20865]_  & ~\new_[30157]_ );
  assign \new_[17686]_  = ~\new_[27821]_  & (~\new_[20833]_  | ~\new_[30000]_ );
  assign \new_[17687]_  = \new_[22487]_  & \new_[19653]_ ;
  assign \new_[17688]_  = \new_[19915]_  | \new_[28098]_ ;
  assign \new_[17689]_  = \new_[19919]_  | \new_[26195]_ ;
  assign \new_[17690]_  = ~\new_[23693]_  & (~\new_[20786]_  | ~\new_[21520]_ );
  assign \new_[17691]_  = ~\new_[19555]_  | ~\new_[26213]_ ;
  assign \new_[17692]_  = ~\new_[19682]_  | ~\new_[31678]_ ;
  assign \new_[17693]_  = ~\new_[26951]_  & (~\new_[20790]_  | ~\new_[29032]_ );
  assign \new_[17694]_  = \new_[19922]_  & \new_[27552]_ ;
  assign \new_[17695]_  = ~\new_[25975]_  & (~\new_[20846]_  | ~\new_[29168]_ );
  assign \new_[17696]_  = ~\new_[27597]_  & (~\new_[20965]_  | ~\new_[30446]_ );
  assign \new_[17697]_  = \new_[22477]_  & \new_[19651]_ ;
  assign \new_[17698]_  = \new_[19917]_  | \new_[26187]_ ;
  assign \new_[17699]_  = \new_[19732]_  | \new_[25488]_ ;
  assign \new_[17700]_  = ~\new_[24705]_  | ~\new_[19845]_  | ~\new_[24889]_ ;
  assign \new_[17701]_  = ~\new_[24892]_  & (~\new_[20905]_  | ~\new_[27946]_ );
  assign \new_[17702]_  = \new_[19953]_  | \new_[29889]_ ;
  assign \new_[17703]_  = \new_[24649]_  & \new_[19652]_ ;
  assign \new_[17704]_  = ~\new_[26405]_  & (~\new_[20877]_  | ~\new_[28840]_ );
  assign \new_[17705]_  = \new_[19938]_  & \new_[28091]_ ;
  assign \new_[17706]_  = ~s0_ack_i | ~\new_[19581]_  | ~\new_[29651]_ ;
  assign \new_[17707]_  = ~s9_ack_i | ~\new_[19559]_  | ~\new_[29706]_ ;
  assign \new_[17708]_  = ~s6_ack_i | ~\new_[19577]_  | ~\new_[29954]_ ;
  assign \new_[17709]_  = ~s13_ack_i | ~\new_[19562]_  | ~\new_[32134]_ ;
  assign \new_[17710]_  = \new_[19940]_  & \new_[27578]_ ;
  assign \new_[17711]_  = ~\new_[28479]_  & (~\new_[20809]_  | ~\new_[28837]_ );
  assign \new_[17712]_  = \new_[19939]_  & \new_[29311]_ ;
  assign \new_[17713]_  = ~s13_err_i | ~\new_[19562]_  | ~\new_[32134]_ ;
  assign \new_[17714]_  = ~\new_[28587]_  | ~\new_[19889]_  | ~\new_[22362]_ ;
  assign \new_[17715]_  = ~\new_[26815]_  & (~\new_[20815]_  | ~\new_[30022]_ );
  assign \new_[17716]_  = ~s0_err_i | ~\new_[19581]_  | ~\new_[29651]_ ;
  assign \new_[17717]_  = ~s9_err_i | ~\new_[19559]_  | ~\new_[29706]_ ;
  assign \new_[17718]_  = ~s6_err_i | ~\new_[19577]_  | ~\new_[29954]_ ;
  assign \new_[17719]_  = ~\new_[28406]_  & (~\new_[20783]_  | ~\new_[30497]_ );
  assign \new_[17720]_  = ~s13_rty_i | ~\new_[19562]_  | ~\new_[32134]_ ;
  assign \new_[17721]_  = ~s0_rty_i | ~\new_[19581]_  | ~\new_[29651]_ ;
  assign \new_[17722]_  = ~s6_rty_i | ~\new_[19577]_  | ~\new_[29954]_ ;
  assign \new_[17723]_  = ~\new_[29338]_  & (~\new_[20916]_  | ~\new_[30107]_ );
  assign \new_[17724]_  = ~\new_[19734]_  & ~\new_[28578]_ ;
  assign \new_[17725]_  = ~\new_[28604]_  | ~\new_[19874]_  | ~\new_[26097]_ ;
  assign \new_[17726]_  = ~\new_[27232]_  & (~\new_[20822]_  | ~\new_[30343]_ );
  assign \new_[17727]_  = ~\new_[24668]_  & (~\new_[20826]_  | ~\new_[28877]_ );
  assign \new_[17728]_  = ~s10_ack_i | ~\new_[19571]_  | ~\new_[29021]_ ;
  assign \new_[17729]_  = \new_[19681]_  | \new_[26314]_ ;
  assign \new_[17730]_  = ~\new_[28496]_  | (~\new_[20774]_  & ~\new_[29959]_ );
  assign \new_[17731]_  = ~\new_[28496]_  | ~\new_[19851]_  | ~\new_[22215]_ ;
  assign \new_[17732]_  = ~s4_ack_i | ~\new_[19572]_  | ~\new_[29963]_ ;
  assign \new_[17733]_  = \new_[19918]_  | \new_[24063]_ ;
  assign \new_[17734]_  = ~\new_[27325]_  & (~\new_[20880]_  | ~\new_[29593]_ );
  assign \new_[17735]_  = ~s10_err_i | ~\new_[19571]_  | ~\new_[29021]_ ;
  assign \new_[17736]_  = ~s4_err_i | ~\new_[19572]_  | ~\new_[29963]_ ;
  assign \new_[17737]_  = \new_[19971]_  | \new_[24273]_ ;
  assign \new_[17738]_  = ~s10_rty_i | ~\new_[19571]_  | ~\new_[29021]_ ;
  assign \new_[17739]_  = ~s4_rty_i | ~\new_[19572]_  | ~\new_[29963]_ ;
  assign \new_[17740]_  = ~\new_[26575]_  & (~\new_[20959]_  | ~\new_[29171]_ );
  assign \new_[17741]_  = ~\new_[27617]_  & (~\new_[20842]_  | ~\new_[30349]_ );
  assign \new_[17742]_  = ~\new_[28802]_  | ~\new_[19898]_  | ~\new_[26408]_ ;
  assign \new_[17743]_  = ~\new_[24511]_  & (~\new_[20843]_  | ~\new_[29162]_ );
  assign \new_[17744]_  = ~\new_[26969]_  & (~\new_[20951]_  | ~\new_[24432]_ );
  assign \new_[17745]_  = \new_[19942]_  | \new_[30033]_ ;
  assign \new_[17746]_  = ~\new_[25127]_  & (~\new_[20944]_  | ~\new_[30344]_ );
  assign \new_[17747]_  = \new_[19944]_  & \new_[28116]_ ;
  assign \new_[17748]_  = ~\new_[28274]_  & (~\new_[20939]_  | ~\new_[28684]_ );
  assign \new_[17749]_  = ~\new_[26560]_  & (~\new_[20845]_  | ~\new_[29271]_ );
  assign \new_[17750]_  = \new_[19643]_  & \new_[29241]_ ;
  assign \new_[17751]_  = ~\new_[25674]_  & (~\new_[20886]_  | ~\new_[28985]_ );
  assign \new_[17752]_  = ~\new_[28707]_  & (~\new_[20848]_  | ~\new_[29015]_ );
  assign \new_[17753]_  = \new_[19946]_  & \new_[29249]_ ;
  assign \new_[17754]_  = ~\new_[28217]_  & (~\new_[20925]_  | ~\new_[30628]_ );
  assign \new_[17755]_  = ~\new_[28572]_  & (~\new_[20850]_  | ~\new_[30627]_ );
  assign \new_[17756]_  = \new_[19575]_  & \new_[30026]_ ;
  assign \new_[17757]_  = \new_[19552]_  & \new_[28726]_ ;
  assign \new_[17758]_  = \new_[19566]_  & \new_[27985]_ ;
  assign \new_[17759]_  = \new_[19554]_  & \new_[30335]_ ;
  assign \new_[17760]_  = \new_[19714]_  | \new_[26825]_ ;
  assign \new_[17761]_  = ~\new_[19578]_  | ~\new_[27901]_ ;
  assign \new_[17762]_  = \new_[19960]_  & \new_[27646]_ ;
  assign \new_[17763]_  = \new_[19931]_  & \new_[28634]_ ;
  assign \new_[17764]_  = ~\new_[28548]_  & (~\new_[20860]_  | ~\new_[28039]_ );
  assign \new_[17765]_  = ~\new_[27580]_  & (~\new_[20765]_  | ~\new_[30329]_ );
  assign \new_[17766]_  = \new_[19913]_  | \new_[26568]_ ;
  assign \new_[17767]_  = \new_[19916]_  | \new_[27743]_ ;
  assign \new_[17768]_  = ~\new_[23778]_  & (~\new_[20950]_  | ~\new_[21547]_ );
  assign \new_[17769]_  = ~\new_[26853]_  & (~\new_[20941]_  | ~\new_[24423]_ );
  assign \new_[17770]_  = ~\new_[26629]_  & (~\new_[20934]_  | ~\new_[29082]_ );
  assign \new_[17771]_  = \new_[19952]_  | \new_[30151]_ ;
  assign \new_[17772]_  = \new_[19972]_  | \new_[26209]_ ;
  assign \new_[17773]_  = ~\new_[28097]_  | ~\new_[19885]_  | ~\new_[22338]_ ;
  assign \new_[17774]_  = \new_[19929]_  | \new_[30375]_ ;
  assign \new_[17775]_  = ~\new_[27697]_  & (~\new_[20994]_  | ~\new_[29355]_ );
  assign \new_[17776]_  = \new_[19963]_  & \new_[27951]_ ;
  assign \new_[17777]_  = \new_[19970]_  | \new_[24430]_ ;
  assign \new_[17778]_  = \new_[22464]_  & \new_[19654]_ ;
  assign \new_[17779]_  = ~\new_[28668]_  & (~\new_[20913]_  | ~\new_[30544]_ );
  assign \new_[17780]_  = \new_[19951]_  | \new_[30275]_ ;
  assign \new_[17781]_  = \new_[19914]_  | \new_[27582]_ ;
  assign \new_[17782]_  = ~\new_[26832]_  & (~\new_[20754]_  | ~\new_[30180]_ );
  assign \new_[17783]_  = ~\new_[26341]_  & (~\new_[20839]_  | ~\new_[29787]_ );
  assign \new_[17784]_  = ~\new_[26450]_  & (~\new_[20915]_  | ~\new_[29785]_ );
  assign \new_[17785]_  = ~\new_[24374]_  & (~\new_[20911]_  | ~\new_[28337]_ );
  assign \new_[17786]_  = ~\new_[19580]_  | ~\new_[23046]_ ;
  assign \new_[17787]_  = \new_[19926]_  & \new_[28632]_ ;
  assign \new_[17788]_  = ~\new_[27700]_  & (~\new_[20904]_  | ~\new_[28732]_ );
  assign \new_[17789]_  = \new_[19957]_  | \new_[30201]_ ;
  assign \new_[17790]_  = \new_[19964]_  | \new_[29792]_ ;
  assign \new_[17791]_  = ~\new_[24430]_  & (~\new_[20910]_  | ~\new_[28285]_ );
  assign \new_[17792]_  = ~\new_[26829]_  & (~\new_[20912]_  | ~\new_[30126]_ );
  assign \new_[17793]_  = \new_[19977]_  | \new_[26308]_ ;
  assign \new_[17794]_  = \new_[19976]_  | \new_[26730]_ ;
  assign \new_[17795]_  = ~\new_[25025]_  & (~\new_[20900]_  | ~\new_[26302]_ );
  assign \new_[17796]_  = ~\new_[28643]_  | ~\new_[20683]_  | ~\new_[21209]_ ;
  assign \new_[17797]_  = ~\new_[27734]_  & (~\new_[20953]_  | ~\new_[30089]_ );
  assign \new_[17798]_  = \new_[19973]_  | \new_[28572]_ ;
  assign \new_[17799]_  = \new_[19968]_  | \new_[29997]_ ;
  assign \new_[17800]_  = ~\new_[26209]_  & (~\new_[20874]_  | ~\new_[28930]_ );
  assign \new_[17801]_  = ~\new_[27534]_  & (~\new_[20922]_  | ~\new_[28280]_ );
  assign \new_[17802]_  = ~\new_[28097]_  | (~\new_[20883]_  & ~\new_[30066]_ );
  assign \new_[17803]_  = ~\new_[24615]_  | ~\new_[19819]_  | ~\new_[25121]_ ;
  assign \new_[17804]_  = ~\new_[27628]_  & (~\new_[20924]_  | ~\new_[28023]_ );
  assign \new_[17805]_  = ~\new_[26617]_  & (~\new_[20938]_  | ~\new_[30411]_ );
  assign \new_[17806]_  = \new_[19663]_  | \new_[25966]_ ;
  assign \new_[17807]_  = \new_[19949]_  & \new_[28480]_ ;
  assign \new_[17808]_  = ~\new_[26561]_  & (~\new_[20873]_  | ~\new_[29086]_ );
  assign \new_[17809]_  = ~\new_[19603]_  | ~\new_[27418]_ ;
  assign \new_[17810]_  = \new_[19948]_  | \new_[30326]_ ;
  assign \new_[17811]_  = ~s4_ack_i | ~\new_[19612]_  | ~\new_[28392]_ ;
  assign \new_[17812]_  = ~\new_[27751]_  & (~\new_[20868]_  | ~\new_[30178]_ );
  assign \new_[17813]_  = ~s4_err_i | ~\new_[19614]_  | ~\new_[28392]_ ;
  assign \new_[17814]_  = ~s4_rty_i | ~\new_[19612]_  | ~\new_[28392]_ ;
  assign \new_[17815]_  = \new_[23922]_  & \new_[19655]_ ;
  assign \new_[17816]_  = ~\new_[28081]_  & (~\new_[20968]_  | ~\new_[28640]_ );
  assign \new_[17817]_  = ~\new_[26308]_  & (~\new_[20936]_  | ~\new_[29608]_ );
  assign \new_[17818]_  = ~\new_[28477]_  | ~\new_[19882]_  | ~\new_[22412]_ ;
  assign \new_[17819]_  = ~\new_[28477]_  | (~\new_[20967]_  & ~\new_[30115]_ );
  assign \new_[17820]_  = ~\new_[28230]_  | ~\new_[19881]_  | ~\new_[25042]_ ;
  assign \new_[17821]_  = ~\new_[19723]_  & ~\new_[23381]_ ;
  assign \new_[17822]_  = ~\new_[26879]_  & (~\new_[20909]_  | ~\new_[30278]_ );
  assign \new_[17823]_  = \new_[19955]_  & \new_[28523]_ ;
  assign \new_[17824]_  = ~\new_[26416]_  & (~\new_[20970]_  | ~\new_[28889]_ );
  assign \new_[17825]_  = ~\new_[19640]_  | ~\new_[27705]_ ;
  assign \new_[17826]_  = \new_[19962]_  & \new_[29284]_ ;
  assign \new_[17827]_  = ~\new_[27629]_  & (~\new_[21002]_  | ~\new_[30117]_ );
  assign \new_[17828]_  = \new_[19752]_  | \new_[25573]_ ;
  assign \new_[17829]_  = ~\new_[25564]_  | ~\new_[19905]_  | ~\new_[24849]_ ;
  assign \new_[17830]_  = ~\new_[25138]_  & (~\new_[20996]_  | ~\new_[27563]_ );
  assign \new_[17831]_  = \new_[19966]_  | \new_[30325]_ ;
  assign \new_[17832]_  = \new_[25269]_  & \new_[19657]_ ;
  assign \new_[17833]_  = ~\new_[19646]_  | ~\new_[26632]_ ;
  assign \new_[17834]_  = ~\new_[28118]_  & (~\new_[20958]_  | ~\new_[28355]_ );
  assign \new_[17835]_  = ~\new_[24586]_  & (~\new_[21000]_  | ~\new_[29455]_ );
  assign \new_[17836]_  = ~\new_[26731]_  & (~\new_[20997]_  | ~\new_[30071]_ );
  assign \new_[17837]_  = \new_[19975]_  | \new_[24586]_ ;
  assign \new_[17838]_  = \new_[22543]_  & \new_[19658]_ ;
  assign \new_[17839]_  = \new_[19756]_  | \new_[23053]_ ;
  assign \new_[17840]_  = ~\new_[19761]_  & ~\new_[23160]_ ;
  assign \new_[17841]_  = \new_[19818]_  | \new_[28503]_ ;
  assign \new_[17842]_  = ~\new_[26352]_  & (~\new_[20764]_  | ~\new_[29251]_ );
  assign \new_[17843]_  = ~\new_[27625]_  & (~\new_[20801]_  | ~\new_[30011]_ );
  assign \new_[17844]_  = \new_[19846]_  | \new_[26385]_ ;
  assign \new_[17845]_  = ~\new_[25892]_  & (~\new_[20828]_  | ~\new_[29984]_ );
  assign \new_[17846]_  = ~\new_[27576]_  | (~\new_[20817]_  & ~\new_[29902]_ );
  assign \new_[17847]_  = ~\new_[24770]_  & (~\new_[20975]_  | ~\new_[29904]_ );
  assign \new_[17848]_  = ~\new_[28612]_  & (~\new_[20952]_  | ~\new_[30717]_ );
  assign \new_[17849]_  = \new_[19859]_  | \new_[29624]_ ;
  assign \new_[17850]_  = ~\new_[28417]_  & (~\new_[20891]_  | ~\new_[30572]_ );
  assign \new_[17851]_  = ~\new_[26313]_  & (~\new_[20893]_  | ~\new_[29404]_ );
  assign \new_[17852]_  = ~\new_[24322]_  & (~\new_[20899]_  | ~\new_[28762]_ );
  assign \new_[17853]_  = ~\new_[24542]_  & (~\new_[20750]_  | ~\new_[30016]_ );
  assign \new_[17854]_  = ~\new_[24861]_  & (~\new_[20957]_  | ~\new_[28888]_ );
  assign \new_[17855]_  = ~\new_[24692]_  & (~\new_[20991]_  | ~\new_[29557]_ );
  assign \new_[17856]_  = ~\new_[27543]_  & (~\new_[20995]_  | ~\new_[29798]_ );
  assign \new_[17857]_  = \new_[19906]_  | \new_[26231]_ ;
  assign \new_[17858]_  = ~\new_[29119]_  & (~\new_[21004]_  | ~\new_[27585]_ );
  assign \new_[17859]_  = ~\new_[30598]_  & (~\new_[21102]_  | ~\new_[29500]_ );
  assign \new_[17860]_  = ~\new_[19664]_  | ~\new_[24283]_ ;
  assign \new_[17861]_  = ~m3_stb_i | ~\new_[20568]_  | ~\new_[29961]_ ;
  assign \new_[17862]_  = ~\new_[30109]_  & (~\new_[21104]_  | ~\new_[29294]_ );
  assign \new_[17863]_  = ~\new_[30564]_  & (~\new_[21105]_  | ~\new_[29344]_ );
  assign \new_[17864]_  = ~\new_[19683]_  | ~\new_[24314]_ ;
  assign \new_[17865]_  = ~\new_[27662]_  | ~\new_[19696]_  | ~\new_[23568]_ ;
  assign \new_[17866]_  = ~\new_[30423]_  & (~\new_[21109]_  | ~\new_[29461]_ );
  assign \new_[17867]_  = ~m5_stb_i | ~\new_[20542]_  | ~\new_[30060]_ ;
  assign \new_[17868]_  = ~\new_[30515]_  & (~\new_[21107]_  | ~\new_[29489]_ );
  assign \new_[17869]_  = ~\new_[28204]_  & (~\new_[21110]_  | ~\new_[29474]_ );
  assign \new_[17870]_  = \new_[19637]_  & \new_[29035]_ ;
  assign \new_[17871]_  = ~\new_[30651]_  & (~\new_[21108]_  | ~\new_[29528]_ );
  assign \new_[17872]_  = ~s10_ack_i | ~\new_[19606]_  | ~\new_[29949]_ ;
  assign \new_[17873]_  = ~s10_err_i | ~\new_[19606]_  | ~\new_[29949]_ ;
  assign \new_[17874]_  = ~s10_rty_i | ~\new_[19606]_  | ~\new_[29949]_ ;
  assign \new_[17875]_  = ~\new_[19713]_  | ~\new_[24443]_ ;
  assign \new_[17876]_  = ~\new_[30063]_  & (~\new_[21103]_  | ~\new_[29480]_ );
  assign \new_[17877]_  = ~s4_rty_i | ~\new_[19584]_  | ~\new_[27855]_ ;
  assign \new_[17878]_  = ~s12_err_i | ~\new_[19626]_  | ~\new_[28957]_ ;
  assign \new_[17879]_  = ~s7_err_i | ~\new_[20567]_  | ~\new_[30131]_ ;
  assign \new_[17880]_  = ~\new_[29205]_  | ~\new_[19648]_  | ~m0_stb_i;
  assign \new_[17881]_  = ~\new_[19728]_  | ~\new_[26198]_ ;
  assign \new_[17882]_  = ~m1_stb_i | ~\new_[19626]_  | ~\new_[28957]_ ;
  assign \new_[17883]_  = ~\new_[29711]_  | ~\new_[20545]_  | ~m0_stb_i;
  assign \new_[17884]_  = ~s4_ack_i | ~\new_[19584]_  | ~\new_[27855]_ ;
  assign \new_[17885]_  = ~s4_ack_i | ~\new_[19632]_  | ~\new_[28842]_ ;
  assign \new_[17886]_  = ~s4_err_i | ~\new_[19632]_  | ~\new_[28842]_ ;
  assign \new_[17887]_  = ~s12_rty_i | ~\new_[20573]_  | ~\new_[28957]_ ;
  assign \new_[17888]_  = ~s4_rty_i | ~\new_[19632]_  | ~\new_[28842]_ ;
  assign \new_[17889]_  = ~\new_[30309]_  & (~\new_[21114]_  | ~\new_[29390]_ );
  assign \new_[17890]_  = ~s7_ack_i | ~\new_[20567]_  | ~\new_[30131]_ ;
  assign \new_[17891]_  = ~\new_[19722]_  | ~\new_[24417]_ ;
  assign \new_[17892]_  = ~\new_[30708]_  & (~\new_[21115]_  | ~\new_[28871]_ );
  assign \new_[17893]_  = ~\new_[29205]_  | ~\new_[19648]_  | ~s11_ack_i;
  assign \new_[17894]_  = ~\new_[19757]_  | ~\new_[24458]_ ;
  assign \new_[17895]_  = \new_[21913]_  | \new_[19820]_ ;
  assign \new_[17896]_  = \new_[22170]_  | \new_[19933]_ ;
  assign \new_[17897]_  = \new_[23248]_  | \new_[19821]_ ;
  assign \new_[17898]_  = ~\new_[29448]_  | ~\new_[19822]_  | ~\new_[23780]_ ;
  assign \new_[17899]_  = \new_[21652]_  | \new_[19879]_ ;
  assign \new_[17900]_  = ~\new_[28586]_  | ~\new_[19888]_  | ~\new_[24831]_ ;
  assign \new_[17901]_  = \new_[21674]_  | \new_[19827]_ ;
  assign \new_[17902]_  = ~\new_[29460]_  | ~\new_[19875]_  | ~\new_[22313]_ ;
  assign \new_[17903]_  = ~\new_[26901]_  | ~\new_[19834]_  | ~\new_[24822]_ ;
  assign \new_[17904]_  = \new_[20738]_  | \new_[19840]_ ;
  assign \new_[17905]_  = \new_[22177]_  | \new_[19935]_ ;
  assign \new_[17906]_  = ~\new_[28218]_  | ~\new_[19841]_  | ~\new_[22178]_ ;
  assign \new_[17907]_  = \new_[22327]_  | \new_[19954]_ ;
  assign \new_[17908]_  = ~\new_[29311]_  | ~\new_[19844]_  | ~\new_[25073]_ ;
  assign \new_[17909]_  = \new_[21259]_  | \new_[19937]_ ;
  assign \new_[17910]_  = \new_[20071]_  | \new_[19847]_ ;
  assign \new_[17911]_  = ~\new_[28091]_  | ~\new_[19848]_  | ~\new_[23598]_ ;
  assign \new_[17912]_  = \new_[22219]_  | \new_[19943]_ ;
  assign \new_[17913]_  = \new_[21879]_  | \new_[19896]_ ;
  assign \new_[17914]_  = \new_[22364]_  | \new_[19945]_ ;
  assign \new_[17915]_  = \new_[20906]_  | \new_[19499]_ ;
  assign \new_[17916]_  = \new_[22384]_  | \new_[19947]_ ;
  assign \new_[17917]_  = ~\new_[28634]_  | ~\new_[19861]_  | ~\new_[23423]_ ;
  assign \new_[17918]_  = \new_[21806]_  | \new_[19865]_ ;
  assign \new_[17919]_  = \new_[21192]_  | \new_[19930]_ ;
  assign \new_[17920]_  = \new_[20933]_  | \new_[19894]_ ;
  assign \new_[17921]_  = ~\new_[27951]_  | ~\new_[19868]_  | ~\new_[23750]_ ;
  assign \new_[17922]_  = ~\new_[28540]_  | ~\new_[19854]_  | ~\new_[26911]_ ;
  assign \new_[17923]_  = \new_[20737]_  | \new_[19880]_ ;
  assign \new_[17924]_  = \new_[21184]_  | \new_[19958]_ ;
  assign \new_[17925]_  = \new_[21200]_  | \new_[19967]_ ;
  assign \new_[17926]_  = ~\new_[29284]_  | ~\new_[19893]_  | ~\new_[22395]_ ;
  assign \new_[17927]_  = ~\new_[29249]_  | ~\new_[19858]_  | ~\new_[24947]_ ;
  assign \new_[17928]_  = ~\new_[28480]_  | ~\new_[19890]_  | ~\new_[23741]_ ;
  assign \new_[17929]_  = \new_[20794]_  | \new_[19842]_ ;
  assign \new_[17930]_  = \new_[21820]_  | \new_[19864]_ ;
  assign \new_[17931]_  = \new_[22374]_  | \new_[19959]_ ;
  assign \new_[17932]_  = ~\new_[28116]_  | ~\new_[19857]_  | ~\new_[23543]_ ;
  assign \new_[17933]_  = ~\new_[29449]_  | ~\new_[19892]_  | ~\new_[25079]_ ;
  assign \new_[17934]_  = ~\new_[28523]_  | ~\new_[19884]_  | ~\new_[23810]_ ;
  assign \new_[17935]_  = \new_[21934]_  | \new_[19883]_ ;
  assign \new_[17936]_  = \new_[22418]_  | \new_[19961]_ ;
  assign \new_[17937]_  = \new_[20999]_  | \new_[19907]_ ;
  assign \new_[17938]_  = ~\new_[29464]_  | ~\new_[19908]_  | ~\new_[26986]_ ;
  assign \new_[17939]_  = ~\new_[21633]_  | (~\new_[21099]_  & ~\new_[28933]_ );
  assign \new_[17940]_  = ~\new_[21654]_  | (~\new_[21069]_  & ~\new_[30285]_ );
  assign \new_[17941]_  = ~\new_[21656]_  | (~\new_[21057]_  & ~\new_[30272]_ );
  assign \new_[17942]_  = ~\new_[20762]_  | (~\new_[21088]_  & ~\new_[30840]_ );
  assign \new_[17943]_  = ~\new_[21717]_  | (~\new_[21063]_  & ~\new_[30192]_ );
  assign \new_[17944]_  = ~\new_[21719]_  | (~\new_[21060]_  & ~\new_[28317]_ );
  assign \new_[17945]_  = ~\new_[20931]_  | (~\new_[21059]_  & ~\new_[29181]_ );
  assign \new_[17946]_  = ~\new_[20856]_  | (~\new_[21075]_  & ~\new_[30656]_ );
  assign \new_[17947]_  = ~\new_[20898]_  | (~\new_[21080]_  & ~\new_[28846]_ );
  assign \new_[17948]_  = ~\new_[25084]_  & (~\new_[21086]_  | ~\new_[27907]_ );
  assign \new_[17949]_  = ~\new_[21326]_  & (~\new_[20735]_  | ~\new_[21257]_ );
  assign \new_[17950]_  = ~\new_[29589]_  | ~\new_[19529]_  | ~\new_[24973]_ ;
  assign \new_[17951]_  = ~\new_[29771]_  | ~\new_[19519]_  | ~\new_[24902]_ ;
  assign \new_[17952]_  = ~\new_[29291]_  | ~\new_[19513]_  | ~\new_[24832]_ ;
  assign \new_[17953]_  = ~\new_[29223]_  | ~\new_[19514]_  | ~\new_[22129]_ ;
  assign \new_[17954]_  = ~\new_[28934]_  | ~\new_[19515]_  | ~\new_[21561]_ ;
  assign \new_[17955]_  = ~\new_[29381]_  | ~\new_[19516]_  | ~\new_[22173]_ ;
  assign \new_[17956]_  = ~\new_[28993]_  | ~\new_[19518]_  | ~\new_[23590]_ ;
  assign \new_[17957]_  = ~\new_[28865]_  | ~\new_[19522]_  | ~\new_[22228]_ ;
  assign \new_[17958]_  = ~\new_[29197]_  | ~\new_[19520]_  | ~\new_[23510]_ ;
  assign \new_[17959]_  = ~\new_[20895]_  | (~\new_[21078]_  & ~\new_[28849]_ );
  assign \new_[17960]_  = ~\new_[28110]_  | ~\new_[19524]_  | ~\new_[24941]_ ;
  assign \new_[17961]_  = ~\new_[29332]_  | ~\new_[19531]_  | ~\new_[24948]_ ;
  assign \new_[17962]_  = ~\new_[30198]_  | ~\new_[19525]_  | ~\new_[24949]_ ;
  assign \new_[17963]_  = ~\new_[30048]_  | ~\new_[19526]_  | ~\new_[23586]_ ;
  assign \new_[17964]_  = ~\new_[30149]_  | ~\new_[19521]_  | ~\new_[24484]_ ;
  assign \new_[17965]_  = ~\new_[30248]_  | ~\new_[19532]_  | ~\new_[25112]_ ;
  assign \new_[17966]_  = ~\new_[30293]_  | ~\new_[19523]_  | ~\new_[23348]_ ;
  assign \new_[17967]_  = ~\new_[29145]_  | ~\new_[19527]_  | ~\new_[22360]_ ;
  assign \new_[17968]_  = ~\new_[29569]_  | ~\new_[19517]_  | ~\new_[23879]_ ;
  assign \new_[17969]_  = ~\new_[29042]_  | ~\new_[19530]_  | ~\new_[25029]_ ;
  assign \new_[17970]_  = ~\new_[29130]_  | ~\new_[19533]_  | ~\new_[24738]_ ;
  assign \new_[17971]_  = ~\new_[20207]_  | ~\new_[30164]_ ;
  assign \new_[17972]_  = ~\new_[20272]_  | ~\new_[27577]_ ;
  assign \new_[17973]_  = ~\new_[20245]_  | ~\new_[30426]_ ;
  assign \new_[17974]_  = ~\new_[20215]_  | ~\new_[30550]_ ;
  assign \new_[17975]_  = ~\new_[20267]_  | ~\new_[27736]_ ;
  assign \new_[17976]_  = ~\new_[20217]_  | ~\new_[29032]_ ;
  assign \new_[17977]_  = ~\new_[20270]_  | ~\new_[26300]_ ;
  assign \new_[17978]_  = ~\new_[20252]_  | ~\new_[30410]_ ;
  assign \new_[17979]_  = ~\new_[20275]_  | ~\new_[24782]_ ;
  assign \new_[17980]_  = ~\new_[20273]_  | ~\new_[27673]_ ;
  assign \new_[17981]_  = ~\new_[20277]_  | ~\new_[27568]_ ;
  assign \new_[17982]_  = ~\new_[20224]_  | ~\new_[29978]_ ;
  assign \new_[17983]_  = ~\new_[20227]_  | ~\new_[29171]_ ;
  assign \new_[17984]_  = ~\new_[20265]_  | ~\new_[27845]_ ;
  assign \new_[17985]_  = ~\new_[20276]_  | ~\new_[26360]_ ;
  assign \new_[17986]_  = ~\new_[20246]_  | ~\new_[29040]_ ;
  assign \new_[17987]_  = ~\new_[20251]_  | ~\new_[30034]_ ;
  assign \new_[17988]_  = ~\new_[20266]_  | ~\new_[26333]_ ;
  assign \new_[17989]_  = ~\new_[20216]_  | ~\new_[30210]_ ;
  assign \new_[17990]_  = ~\new_[20240]_  | ~\new_[29061]_ ;
  assign \new_[17991]_  = ~\new_[20268]_  | ~\new_[27769]_ ;
  assign \new_[17992]_  = ~\new_[20278]_  | ~\new_[26267]_ ;
  assign \new_[17993]_  = ~\new_[20263]_  | ~\new_[30723]_ ;
  assign \new_[17994]_  = ~\new_[20274]_  | ~\new_[26745]_ ;
  assign \new_[17995]_  = ~\new_[20280]_  | ~\new_[27474]_ ;
  assign \new_[17996]_  = ~\new_[20281]_  | ~\new_[27691]_ ;
  assign \new_[17997]_  = ~\new_[20242]_  | ~\new_[28188]_ ;
  assign \new_[17998]_  = ~\new_[20260]_  | ~\new_[28850]_ ;
  assign \new_[17999]_  = ~\new_[24756]_  & (~\new_[21118]_  | ~\new_[29357]_ );
  assign \new_[18000]_  = \new_[20205]_  & \new_[24491]_ ;
  assign \new_[18001]_  = ~\new_[30697]_  | ~\new_[20173]_  | ~\new_[30728]_ ;
  assign \new_[18002]_  = ~\new_[18733]_ ;
  assign \new_[18003]_  = ~\new_[18735]_ ;
  assign \new_[18004]_  = ~\new_[18736]_ ;
  assign \new_[18005]_  = ~\new_[18737]_ ;
  assign \new_[18006]_  = ~\new_[18739]_ ;
  assign \new_[18007]_  = \new_[18742]_ ;
  assign \new_[18008]_  = \new_[23441]_  & \new_[20131]_ ;
  assign \new_[18009]_  = ~\new_[19544]_ ;
  assign \new_[18010]_  = ~\new_[20543]_ ;
  assign \new_[18011]_  = ~\new_[20543]_ ;
  assign \new_[18012]_  = ~\new_[18745]_ ;
  assign \new_[18013]_  = ~\new_[18760]_ ;
  assign \new_[18014]_  = ~\new_[18761]_ ;
  assign \new_[18015]_  = ~\new_[18761]_ ;
  assign \new_[18016]_  = ~\new_[18761]_ ;
  assign \new_[18017]_  = \new_[20231]_  | \new_[30287]_ ;
  assign \new_[18018]_  = ~\new_[18772]_ ;
  assign \new_[18019]_  = ~\new_[18772]_ ;
  assign \new_[18020]_  = ~\new_[18772]_ ;
  assign \new_[18021]_  = ~\new_[28001]_  | ~\new_[20181]_  | ~\new_[30142]_ ;
  assign \new_[18022]_  = \new_[20249]_  & \new_[24097]_ ;
  assign \new_[18023]_  = \new_[23639]_  & \new_[20020]_ ;
  assign \new_[18024]_  = \new_[20213]_  | \new_[30109]_ ;
  assign \new_[18025]_  = \new_[20214]_  & \new_[23090]_ ;
  assign \new_[18026]_  = ~\new_[18776]_ ;
  assign \new_[18027]_  = ~\new_[18780]_ ;
  assign \new_[18028]_  = ~\new_[29251]_  | ~\new_[20160]_  | ~\new_[30505]_ ;
  assign \new_[18029]_  = \new_[20211]_  | \new_[30174]_ ;
  assign \new_[18030]_  = ~\new_[18785]_ ;
  assign \new_[18031]_  = ~\new_[18785]_ ;
  assign \new_[18032]_  = ~\new_[26413]_  & ~\new_[20037]_ ;
  assign \new_[18033]_  = \new_[24610]_  & \new_[20038]_ ;
  assign \new_[18034]_  = ~\new_[18787]_ ;
  assign \new_[18035]_  = ~\new_[18788]_ ;
  assign \new_[18036]_  = ~\new_[18788]_ ;
  assign \new_[18037]_  = ~\new_[18788]_ ;
  assign \new_[18038]_  = ~\new_[18788]_ ;
  assign \new_[18039]_  = ~\new_[18788]_ ;
  assign \new_[18040]_  = ~\new_[18788]_ ;
  assign \new_[18041]_  = ~\new_[18790]_ ;
  assign \new_[18042]_  = ~\new_[18791]_ ;
  assign \new_[18043]_  = ~\new_[18791]_ ;
  assign \new_[18044]_  = ~\new_[18791]_ ;
  assign \new_[18045]_  = ~\new_[18791]_ ;
  assign \new_[18046]_  = ~\new_[18791]_ ;
  assign \new_[18047]_  = ~\new_[18791]_ ;
  assign \new_[18048]_  = ~\new_[18793]_ ;
  assign \new_[18049]_  = ~\new_[18793]_ ;
  assign \new_[18050]_  = ~\new_[18793]_ ;
  assign \new_[18051]_  = ~\new_[18793]_ ;
  assign \new_[18052]_  = ~\new_[19564]_ ;
  assign \new_[18053]_  = ~\new_[18796]_ ;
  assign \new_[18054]_  = ~\new_[18796]_ ;
  assign \new_[18055]_  = ~\new_[18796]_ ;
  assign \new_[18056]_  = ~\new_[18796]_ ;
  assign \new_[18057]_  = ~\new_[18796]_ ;
  assign \new_[18058]_  = ~\new_[18796]_ ;
  assign \new_[18059]_  = ~\new_[18796]_ ;
  assign \new_[18060]_  = ~\new_[18796]_ ;
  assign \new_[18061]_  = ~\new_[18796]_ ;
  assign \new_[18062]_  = ~\new_[18796]_ ;
  assign \new_[18063]_  = ~\new_[18796]_ ;
  assign \new_[18064]_  = ~\new_[18796]_ ;
  assign \new_[18065]_  = ~\new_[18796]_ ;
  assign \new_[18066]_  = ~\new_[18797]_ ;
  assign \new_[18067]_  = ~\new_[18798]_ ;
  assign \new_[18068]_  = ~\new_[18798]_ ;
  assign \new_[18069]_  = ~\new_[18798]_ ;
  assign \new_[18070]_  = ~\new_[26413]_  & ~\new_[20796]_ ;
  assign \new_[18071]_  = ~\new_[26269]_  & (~\new_[21210]_  | ~\new_[29104]_ );
  assign \new_[18072]_  = ~\new_[18803]_ ;
  assign \new_[18073]_  = ~\new_[18806]_ ;
  assign \new_[18074]_  = ~\new_[18807]_ ;
  assign \new_[18075]_  = ~\new_[18807]_ ;
  assign \new_[18076]_  = ~\new_[18808]_ ;
  assign \new_[18077]_  = ~\new_[18809]_ ;
  assign \new_[18078]_  = ~\new_[18809]_ ;
  assign \new_[18079]_  = ~\new_[18809]_ ;
  assign \new_[18080]_  = \new_[24610]_  & \new_[20045]_ ;
  assign \new_[18081]_  = ~\new_[28898]_  | ~\new_[20163]_  | ~\new_[30016]_ ;
  assign \new_[18082]_  = \new_[20237]_  & \new_[26275]_ ;
  assign \new_[18083]_  = ~\new_[18810]_ ;
  assign \new_[18084]_  = \new_[20221]_  & \new_[23121]_ ;
  assign \new_[18085]_  = ~\new_[21250]_  | ~\new_[22102]_  | ~\new_[22413]_ ;
  assign \new_[18086]_  = ~\new_[18813]_ ;
  assign \new_[18087]_  = ~\new_[18814]_ ;
  assign \new_[18088]_  = \new_[20228]_  & \new_[23621]_ ;
  assign \new_[18089]_  = ~\new_[18817]_ ;
  assign \new_[18090]_  = ~\new_[18820]_ ;
  assign \new_[18091]_  = ~\new_[18821]_ ;
  assign \new_[18092]_  = ~\new_[18822]_ ;
  assign \new_[18093]_  = ~\new_[18823]_ ;
  assign \new_[18094]_  = ~\new_[18823]_ ;
  assign \new_[18095]_  = \new_[26956]_  & \new_[20036]_ ;
  assign \new_[18096]_  = ~\new_[23529]_  & ~\new_[20037]_ ;
  assign \new_[18097]_  = ~\new_[18826]_ ;
  assign \new_[18098]_  = ~\new_[18827]_ ;
  assign \new_[18099]_  = ~\new_[18827]_ ;
  assign \new_[18100]_  = ~\new_[18827]_ ;
  assign \new_[18101]_  = ~\new_[18827]_ ;
  assign \new_[18102]_  = ~\new_[18827]_ ;
  assign \new_[18103]_  = ~\new_[18827]_ ;
  assign \new_[18104]_  = ~\new_[18827]_ ;
  assign \new_[18105]_  = ~\new_[18827]_ ;
  assign \new_[18106]_  = ~\new_[18827]_ ;
  assign \new_[18107]_  = ~\new_[18827]_ ;
  assign \new_[18108]_  = ~\new_[18827]_ ;
  assign \new_[18109]_  = ~\new_[18827]_ ;
  assign \new_[18110]_  = ~\new_[18827]_ ;
  assign \new_[18111]_  = ~\new_[18828]_ ;
  assign \new_[18112]_  = ~\new_[18833]_ ;
  assign \new_[18113]_  = ~\new_[18833]_ ;
  assign \new_[18114]_  = ~\new_[18833]_ ;
  assign \new_[18115]_  = ~\new_[18834]_ ;
  assign \new_[18116]_  = ~\new_[18834]_ ;
  assign \new_[18117]_  = ~\new_[18836]_ ;
  assign \new_[18118]_  = \new_[20229]_  & \new_[21884]_ ;
  assign \new_[18119]_  = ~\new_[18837]_ ;
  assign \new_[18120]_  = ~\new_[29299]_  | ~\new_[20166]_  | ~\new_[30321]_ ;
  assign \new_[18121]_  = \new_[20250]_  | \new_[29916]_ ;
  assign \new_[18122]_  = ~\new_[28828]_  | ~\new_[20167]_  | ~\new_[29404]_ ;
  assign \new_[18123]_  = \new_[20258]_  | \new_[28204]_ ;
  assign \new_[18124]_  = ~\new_[18846]_ ;
  assign \new_[18125]_  = \new_[18846]_ ;
  assign \new_[18126]_  = \new_[20243]_  & \new_[24065]_ ;
  assign \new_[18127]_  = ~\new_[18849]_ ;
  assign \new_[18128]_  = \new_[18849]_ ;
  assign \new_[18129]_  = ~\new_[18850]_ ;
  assign \new_[18130]_  = ~\new_[18851]_ ;
  assign \new_[18131]_  = \new_[20238]_  & \new_[22887]_ ;
  assign \new_[18132]_  = \new_[20232]_  | \new_[30445]_ ;
  assign \new_[18133]_  = ~\new_[26349]_  & (~\new_[21230]_  | ~\new_[29744]_ );
  assign \new_[18134]_  = \new_[20241]_  & \new_[23152]_ ;
  assign \new_[18135]_  = ~\new_[20813]_  | ~\new_[21243]_  | ~\new_[22102]_ ;
  assign \new_[18136]_  = \new_[20255]_  | \new_[30423]_ ;
  assign \new_[18137]_  = \new_[20234]_  & \new_[22982]_ ;
  assign \new_[18138]_  = ~\new_[21250]_  | ~\new_[21245]_  | ~\new_[22102]_ ;
  assign \new_[18139]_  = \new_[20257]_  & \new_[23118]_ ;
  assign \new_[18140]_  = \new_[20209]_  & \new_[23417]_ ;
  assign \new_[18141]_  = ~\new_[19608]_ ;
  assign \new_[18142]_  = ~\new_[18876]_ ;
  assign \new_[18143]_  = ~\new_[18876]_ ;
  assign \new_[18144]_  = ~\new_[18876]_ ;
  assign \new_[18145]_  = ~\new_[18876]_ ;
  assign \new_[18146]_  = ~\new_[18876]_ ;
  assign \new_[18147]_  = ~\new_[18876]_ ;
  assign \new_[18148]_  = ~\new_[18878]_ ;
  assign \new_[18149]_  = \new_[18879]_ ;
  assign \new_[18150]_  = ~\new_[18880]_ ;
  assign \new_[18151]_  = ~\new_[18881]_ ;
  assign \new_[18152]_  = ~\new_[24965]_  & (~\new_[21187]_  | ~\new_[28962]_ );
  assign \new_[18153]_  = ~\new_[18882]_ ;
  assign \new_[18154]_  = \new_[24870]_  & \new_[20131]_ ;
  assign \new_[18155]_  = ~\new_[18883]_ ;
  assign \new_[18156]_  = ~\new_[18883]_ ;
  assign \new_[18157]_  = ~\new_[18883]_ ;
  assign \new_[18158]_  = ~\new_[18884]_ ;
  assign \new_[18159]_  = ~\new_[18885]_ ;
  assign \new_[18160]_  = ~\new_[18885]_ ;
  assign \new_[18161]_  = ~\new_[18885]_ ;
  assign \new_[18162]_  = ~\new_[18885]_ ;
  assign \new_[18163]_  = ~\new_[18885]_ ;
  assign \new_[18164]_  = ~\new_[18885]_ ;
  assign \new_[18165]_  = ~\new_[18885]_ ;
  assign \new_[18166]_  = ~\new_[18886]_ ;
  assign \new_[18167]_  = ~\new_[18889]_ ;
  assign \new_[18168]_  = ~\new_[18902]_ ;
  assign \new_[18169]_  = ~\new_[18902]_ ;
  assign \new_[18170]_  = ~\new_[18902]_ ;
  assign \new_[18171]_  = ~\new_[18902]_ ;
  assign \new_[18172]_  = ~\new_[18902]_ ;
  assign \new_[18173]_  = ~\new_[18902]_ ;
  assign \new_[18174]_  = ~\new_[18903]_ ;
  assign \new_[18175]_  = ~\new_[18904]_ ;
  assign \new_[18176]_  = ~\new_[18906]_ ;
  assign \new_[18177]_  = \new_[18906]_ ;
  assign \new_[18178]_  = ~\new_[18910]_ ;
  assign \new_[18179]_  = ~\new_[18910]_ ;
  assign \new_[18180]_  = \new_[18910]_ ;
  assign \new_[18181]_  = ~\new_[18914]_ ;
  assign \new_[18182]_  = ~\new_[18914]_ ;
  assign \new_[18183]_  = ~\new_[18914]_ ;
  assign \new_[18184]_  = ~\new_[18914]_ ;
  assign \new_[18185]_  = ~\new_[18914]_ ;
  assign \new_[18186]_  = ~\new_[18914]_ ;
  assign \new_[18187]_  = ~\new_[18914]_ ;
  assign \new_[18188]_  = ~\new_[18914]_ ;
  assign \new_[18189]_  = ~\new_[18914]_ ;
  assign \new_[18190]_  = ~\new_[18914]_ ;
  assign \new_[18191]_  = ~\new_[18914]_ ;
  assign \new_[18192]_  = \new_[25999]_  & \new_[20020]_ ;
  assign \new_[18193]_  = ~\new_[18915]_ ;
  assign \new_[18194]_  = ~\new_[18927]_ ;
  assign \new_[18195]_  = ~\new_[29441]_  | ~\new_[20164]_  | ~\new_[29904]_ ;
  assign \new_[18196]_  = ~\new_[18931]_ ;
  assign \new_[18197]_  = ~\new_[18931]_ ;
  assign \new_[18198]_  = ~\new_[18931]_ ;
  assign \new_[18199]_  = ~\new_[18931]_ ;
  assign \new_[18200]_  = ~\new_[18933]_ ;
  assign \new_[18201]_  = ~\new_[18935]_ ;
  assign \new_[18202]_  = ~\new_[29226]_  | ~\new_[20201]_  | ~\new_[29557]_ ;
  assign \new_[18203]_  = ~\new_[18940]_ ;
  assign \new_[18204]_  = ~\new_[18940]_ ;
  assign \new_[18205]_  = \new_[20259]_  & \new_[23569]_ ;
  assign \new_[18206]_  = ~\new_[18942]_ ;
  assign \new_[18207]_  = ~\new_[18942]_ ;
  assign \new_[18208]_  = ~\new_[29692]_  | ~\new_[28050]_  | ~\new_[19979]_  | ~\new_[29168]_ ;
  assign \new_[18209]_  = ~\new_[29874]_  | ~\new_[28114]_  | ~\new_[19987]_  | ~\new_[29550]_ ;
  assign \new_[18210]_  = ~\new_[30215]_  | ~\new_[29969]_  | ~\new_[19985]_  | ~\new_[29003]_ ;
  assign \new_[18211]_  = ~\new_[30508]_  | ~\new_[29435]_  | ~\new_[23189]_  | ~\new_[29159]_ ;
  assign \new_[18212]_  = ~\new_[29260]_  | ~\new_[29983]_  | ~\new_[19978]_  | ~\new_[29192]_ ;
  assign \new_[18213]_  = ~\new_[29560]_  | ~\new_[30117]_  | ~\new_[19990]_  | ~\new_[30411]_ ;
  assign \new_[18214]_  = ~\new_[29977]_  | ~\new_[29186]_  | ~\new_[19981]_  | ~\new_[29397]_ ;
  assign \new_[18215]_  = ~\new_[29139]_  | ~\new_[28121]_  | ~\new_[19980]_  | ~\new_[28877]_ ;
  assign \new_[18216]_  = ~\new_[29887]_  | ~\new_[28245]_  | ~\new_[19984]_  | ~\new_[28930]_ ;
  assign \new_[18217]_  = ~\new_[30316]_  | ~\new_[28732]_  | ~\new_[19982]_  | ~\new_[28985]_ ;
  assign \new_[18218]_  = ~\new_[30610]_  | ~\new_[28935]_  | ~\new_[19986]_  | ~\new_[30751]_ ;
  assign \new_[18219]_  = ~\new_[30246]_  | ~\new_[28684]_  | ~\new_[19983]_  | ~\new_[29271]_ ;
  assign \new_[18220]_  = ~\new_[30021]_  | ~\new_[28355]_  | ~\new_[19988]_  | ~\new_[29455]_ ;
  assign \new_[18221]_  = ~\new_[30084]_  | ~\new_[28640]_  | ~\new_[19989]_  | ~\new_[29608]_ ;
  assign \new_[18222]_  = ~\new_[18961]_ ;
  assign \new_[18223]_  = ~\new_[28732]_  | ~\new_[20178]_  | ~\new_[30158]_ ;
  assign \new_[18224]_  = ~\new_[28114]_  | ~\new_[20154]_  | ~\new_[28845]_ ;
  assign \new_[18225]_  = ~\new_[22392]_  | ~\new_[24184]_  | ~\new_[27577]_  | ~\new_[30242]_ ;
  assign \new_[18226]_  = ~\new_[22316]_  & (~\new_[21340]_  | ~\new_[25197]_ );
  assign \new_[18227]_  = ~\new_[22388]_  | ~\new_[22877]_  | ~\new_[26374]_  | ~\new_[29028]_ ;
  assign \new_[18228]_  = ~\new_[29855]_  & (~\new_[21266]_  | ~\new_[23360]_ );
  assign \new_[18229]_  = ~\new_[18972]_ ;
  assign \new_[18230]_  = ~\new_[29855]_  & (~\new_[21266]_  | ~\new_[26664]_ );
  assign \new_[18231]_  = ~\new_[21163]_  & (~\new_[21509]_  | ~\new_[23898]_ );
  assign \new_[18232]_  = ~\new_[18973]_ ;
  assign \new_[18233]_  = ~\new_[20334]_  & (~\new_[22967]_  | ~\new_[23928]_ );
  assign \new_[18234]_  = ~\new_[20334]_  & (~\new_[21329]_  | ~\new_[23928]_ );
  assign \new_[18235]_  = ~\new_[23388]_  & (~\new_[21337]_  | ~\new_[27001]_ );
  assign \new_[18236]_  = ~\new_[30754]_  | ~\new_[23020]_  | ~\new_[23684]_  | ~\new_[22974]_ ;
  assign \new_[18237]_  = ~\new_[29100]_  & (~\new_[21302]_  | ~\new_[23392]_ );
  assign \new_[18238]_  = ~\new_[18980]_ ;
  assign \new_[18239]_  = ~\new_[29100]_  & (~\new_[21302]_  | ~\new_[27093]_ );
  assign \new_[18240]_  = ~\new_[18982]_ ;
  assign \new_[18241]_  = ~\new_[18984]_ ;
  assign \new_[18242]_  = ~\new_[29767]_  & (~\new_[21274]_  | ~\new_[26710]_ );
  assign \new_[18243]_  = ~\new_[29983]_  | ~\new_[20157]_  | ~\new_[30386]_ ;
  assign \new_[18244]_  = ~\new_[24863]_  & (~\new_[21331]_  | ~\new_[27003]_ );
  assign \new_[18245]_  = ~\new_[30676]_  | ~\new_[22957]_  | ~\new_[24903]_  | ~\new_[26556]_ ;
  assign \new_[18246]_  = ~\new_[25123]_  & (~\new_[21338]_  | ~\new_[22507]_ );
  assign \new_[18247]_  = ~\new_[30389]_  & (~\new_[21269]_  | ~\new_[24531]_ );
  assign \new_[18248]_  = ~\new_[18990]_ ;
  assign \new_[18249]_  = ~\new_[30389]_  & (~\new_[21269]_  | ~\new_[27556]_ );
  assign \new_[18250]_  = ~\new_[18992]_ ;
  assign \new_[18251]_  = ~\new_[28050]_  | ~\new_[20161]_  | ~\new_[28880]_ ;
  assign \new_[18252]_  = ~\new_[26907]_  & (~\new_[21335]_  | ~\new_[24652]_ );
  assign \new_[18253]_  = ~\new_[28899]_  & (~\new_[21275]_  | ~\new_[23459]_ );
  assign \new_[18254]_  = ~\new_[28899]_  & (~\new_[21275]_  | ~\new_[26675]_ );
  assign \new_[18255]_  = ~\new_[29186]_  | ~\new_[20169]_  | ~\new_[29150]_ ;
  assign \new_[18256]_  = ~\new_[20813]_  | ~\new_[21055]_  | ~\new_[22411]_ ;
  assign \new_[18257]_  = ~\new_[22280]_  & (~\new_[21332]_  | ~\new_[24600]_ );
  assign \new_[18258]_  = ~\new_[24940]_  & (~\new_[21333]_  | ~\new_[25266]_ );
  assign \new_[18259]_  = ~\new_[20046]_  | ~\new_[29682]_ ;
  assign \new_[18260]_  = ~\new_[21202]_  & (~\new_[21336]_  | ~\new_[23917]_ );
  assign \new_[18261]_  = ~\new_[30563]_  | ~\new_[22952]_  | ~\new_[23486]_  | ~\new_[26302]_ ;
  assign \new_[18262]_  = ~\new_[22147]_  | ~\new_[24406]_  | ~\new_[27673]_  | ~\new_[30467]_ ;
  assign \new_[18263]_  = ~\new_[19008]_ ;
  assign \new_[18264]_  = ~\new_[19009]_ ;
  assign \new_[18265]_  = ~\new_[19013]_ ;
  assign \new_[18266]_  = ~\new_[30553]_  & (~\new_[21190]_  | ~\new_[24982]_ );
  assign \new_[18267]_  = ~\new_[22337]_  | ~\new_[24398]_  | ~\new_[27568]_  | ~\new_[30198]_ ;
  assign \new_[18268]_  = ~\new_[19017]_ ;
  assign \new_[18269]_  = ~\new_[19018]_ ;
  assign \new_[18270]_  = ~\new_[22416]_  & (~\new_[22880]_  | ~\new_[21291]_ );
  assign \new_[18271]_  = ~\new_[28121]_  | ~\new_[20162]_  | ~\new_[30279]_ ;
  assign \new_[18272]_  = ~\new_[22398]_  | ~\new_[22960]_  | ~\new_[26347]_  | ~\new_[29276]_ ;
  assign \new_[18273]_  = ~\new_[22404]_  | ~\new_[24153]_  | ~\new_[27845]_  | ~\new_[30599]_ ;
  assign \new_[18274]_  = ~\new_[29573]_  & (~\new_[21292]_  | ~\new_[23593]_ );
  assign \new_[18275]_  = ~\new_[19030]_ ;
  assign \new_[18276]_  = ~\new_[29573]_  & (~\new_[21292]_  | ~\new_[26755]_ );
  assign \new_[18277]_  = ~\new_[29565]_  & (~\new_[21310]_  | ~\new_[26727]_ );
  assign \new_[18278]_  = ~\new_[19031]_ ;
  assign \new_[18279]_  = ~\new_[22411]_  | ~\new_[22413]_  | ~\new_[21250]_ ;
  assign \new_[18280]_  = ~\new_[21562]_  & (~\new_[21330]_  | ~\new_[23894]_ );
  assign \new_[18281]_  = ~\new_[30725]_  | ~\new_[23002]_  | ~\new_[23421]_  | ~\new_[24498]_ ;
  assign \new_[18282]_  = ~\new_[29767]_  & (~\new_[21274]_  | ~\new_[23617]_ );
  assign \new_[18283]_  = ~\new_[19035]_ ;
  assign \new_[18284]_  = ~\new_[19036]_ ;
  assign \new_[18285]_  = ~\new_[29648]_  & (~\new_[21290]_  | ~\new_[26847]_ );
  assign \new_[18286]_  = ~\new_[22275]_  & (~\new_[22982]_  | ~\new_[21297]_ );
  assign \new_[18287]_  = ~\new_[29648]_  & (~\new_[21290]_  | ~\new_[23791]_ );
  assign \new_[18288]_  = ~\new_[19044]_ ;
  assign \new_[18289]_  = ~\new_[19045]_ ;
  assign \new_[18290]_  = ~\new_[28023]_  | ~\new_[20175]_  | ~\new_[29225]_ ;
  assign \new_[18291]_  = ~\new_[19047]_ ;
  assign \new_[18292]_  = ~\new_[22416]_  & (~\new_[21334]_  | ~\new_[21291]_ );
  assign \new_[18293]_  = ~\new_[19053]_ ;
  assign \new_[18294]_  = ~\new_[29435]_  | ~\new_[20156]_  | ~\new_[30232]_ ;
  assign \new_[18295]_  = ~\new_[21206]_  & (~\new_[21341]_  | ~\new_[23952]_ );
  assign \new_[18296]_  = ~\new_[29898]_  & (~\new_[21323]_  | ~\new_[23499]_ );
  assign \new_[18297]_  = ~\new_[19061]_ ;
  assign \new_[18298]_  = ~\new_[19062]_ ;
  assign \new_[18299]_  = ~\new_[30775]_  | ~\new_[22962]_  | ~\new_[23858]_  | ~\new_[24416]_ ;
  assign \new_[18300]_  = ~\new_[28280]_  | ~\new_[20183]_  | ~\new_[29685]_ ;
  assign \new_[18301]_  = ~\new_[29565]_  & (~\new_[21310]_  | ~\new_[23665]_ );
  assign \new_[18302]_  = ~\new_[23720]_  & (~\new_[21884]_  | ~\new_[21311]_ );
  assign \new_[18303]_  = ~\new_[28245]_  | ~\new_[20182]_  | ~\new_[29506]_ ;
  assign \new_[18304]_  = ~\new_[19069]_ ;
  assign \new_[18305]_  = ~\new_[29969]_  | ~\new_[20155]_  | ~\new_[29220]_ ;
  assign \new_[18306]_  = ~\new_[25014]_  & (~\new_[22887]_  | ~\new_[21300]_ );
  assign \new_[18307]_  = ~\new_[28867]_  & (~\new_[21201]_  | ~\new_[23652]_ );
  assign \new_[18308]_  = ~\new_[22413]_  | ~\new_[20813]_  | ~\new_[22411]_ ;
  assign \new_[18309]_  = ~\new_[28684]_  | ~\new_[20165]_  | ~\new_[28870]_ ;
  assign \new_[18310]_  = ~\new_[22204]_  & (~\new_[21465]_  | ~\new_[24685]_ );
  assign \new_[18311]_  = ~\new_[29898]_  & (~\new_[21323]_  | ~\new_[26738]_ );
  assign \new_[18312]_  = ~\new_[22183]_  | ~\new_[27587]_  | ~\new_[27904]_  | ~\new_[30015]_ ;
  assign \new_[18313]_  = ~\new_[28355]_  | ~\new_[20204]_  | ~\new_[28371]_ ;
  assign n7664 = ~\new_[28916]_  | ~\new_[20191]_ ;
  assign \new_[18315]_  = ~\new_[30652]_  & (~\new_[21203]_  | ~\new_[23604]_ );
  assign \new_[18316]_  = ~\new_[28640]_  | ~\new_[20179]_  | ~\new_[28926]_ ;
  assign \new_[18317]_  = ~\new_[19090]_ ;
  assign \new_[18318]_  = ~\new_[19091]_ ;
  assign \new_[18319]_  = ~\new_[21248]_  & (~\new_[21339]_  | ~\new_[25188]_ );
  assign \new_[18320]_  = ~\new_[19097]_ ;
  assign \new_[18321]_  = ~\new_[19098]_ ;
  assign \new_[18322]_  = ~\new_[29906]_  & (~\new_[21256]_  | ~\new_[23862]_ );
  assign \new_[18323]_  = ~\new_[19108]_ ;
  assign \new_[18324]_  = ~\new_[20003]_  | ~\new_[30352]_ ;
  assign \new_[18325]_  = ~\new_[20006]_  | ~\new_[30337]_ ;
  assign \new_[18326]_  = ~\new_[20014]_  | ~\new_[29320]_ ;
  assign \new_[18327]_  = ~\new_[20018]_  | ~\new_[29975]_ ;
  assign \new_[18328]_  = ~\new_[29975]_  | (~\new_[21128]_  & ~\new_[23400]_ );
  assign \new_[18329]_  = ~\new_[20030]_  | ~\new_[29228]_ ;
  assign \new_[18330]_  = ~\new_[20027]_  | ~\new_[30505]_ ;
  assign \new_[18331]_  = ~\new_[30505]_  | (~\new_[21559]_  & ~\new_[23408]_ );
  assign \new_[18332]_  = ~\new_[20032]_  | ~\new_[29103]_ ;
  assign \new_[18333]_  = ~\new_[20048]_  | ~\new_[30728]_ ;
  assign \new_[18334]_  = ~\new_[20060]_  | ~\new_[29695]_ ;
  assign \new_[18335]_  = ~\new_[20149]_  | ~\new_[29441]_ ;
  assign \new_[18336]_  = ~\new_[20029]_  | ~\new_[28963]_ ;
  assign \new_[18337]_  = ~\new_[20125]_  | ~\new_[28898]_ ;
  assign \new_[18338]_  = ~\new_[20097]_  | ~\new_[28828]_ ;
  assign \new_[18339]_  = ~\new_[20076]_  & ~\new_[30053]_ ;
  assign \new_[18340]_  = ~\new_[20011]_  | ~\new_[29721]_ ;
  assign \new_[18341]_  = ~\new_[20024]_  | ~\new_[30321]_ ;
  assign \new_[18342]_  = ~\new_[30321]_  | (~\new_[21204]_  & ~\new_[23536]_ );
  assign \new_[18343]_  = ~\new_[29979]_  | (~\new_[22190]_  & ~\new_[21198]_ );
  assign \new_[18344]_  = ~\new_[30563]_  | (~\new_[22296]_  & ~\new_[21219]_ );
  assign \new_[18345]_  = ~\new_[20102]_  | ~\new_[29456]_ ;
  assign \new_[18346]_  = ~\new_[20108]_  & ~\new_[29989]_ ;
  assign \new_[18347]_  = ~\new_[20098]_  & ~\new_[29508]_ ;
  assign \new_[18348]_  = ~\new_[20008]_  & ~\new_[28397]_ ;
  assign \new_[18349]_  = ~\new_[20120]_  | ~\new_[29527]_ ;
  assign \new_[18350]_  = ~\new_[20057]_  | ~\new_[29006]_ ;
  assign \new_[18351]_  = ~\new_[29867]_  | (~\new_[21238]_  & ~\new_[25108]_ );
  assign \new_[18352]_  = ~\new_[20134]_  | ~\new_[29813]_ ;
  assign \new_[18353]_  = ~\new_[30009]_  | (~\new_[21251]_  & ~\new_[22256]_ );
  assign \new_[18354]_  = ~\new_[20141]_  | ~\new_[29226]_ ;
  assign \new_[18355]_  = ~\new_[20143]_  | ~\new_[29802]_ ;
  assign \new_[18356]_  = ~\new_[20146]_  & ~\new_[29931]_ ;
  assign \new_[18357]_  = ~\new_[20151]_  | ~\new_[30150]_ ;
  assign \new_[18358]_  = ~\new_[24360]_  | ~\new_[20042]_ ;
  assign \new_[18359]_  = ~\new_[24080]_  & (~\new_[21285]_  | ~\new_[26315]_ );
  assign \new_[18360]_  = ~\new_[24293]_  & (~\new_[21286]_  | ~\new_[24564]_ );
  assign \new_[18361]_  = ~\new_[24418]_  & (~\new_[21273]_  | ~\new_[26121]_ );
  assign \new_[18362]_  = ~\new_[24507]_  & (~\new_[21309]_  | ~\new_[26287]_ );
  assign \new_[18363]_  = ~\new_[23007]_  & (~\new_[21278]_  | ~\new_[26330]_ );
  assign \new_[18364]_  = ~\new_[24284]_  & (~\new_[21284]_  | ~\new_[22956]_ );
  assign \new_[18365]_  = ~\new_[24261]_  & (~\new_[21316]_  | ~\new_[25767]_ );
  assign \new_[18366]_  = ~\new_[20330]_  | ~\new_[28564]_ ;
  assign \new_[18367]_  = ~\new_[20335]_  | ~\new_[26995]_ ;
  assign \new_[18368]_  = ~\new_[19288]_ ;
  assign \new_[18369]_  = ~\new_[19289]_ ;
  assign \new_[18370]_  = ~\new_[19292]_ ;
  assign \new_[18371]_  = ~\new_[19294]_ ;
  assign \new_[18372]_  = ~\new_[19296]_ ;
  assign \new_[18373]_  = ~\new_[19298]_ ;
  assign \new_[18374]_  = ~\new_[19299]_ ;
  assign \new_[18375]_  = ~\new_[19303]_ ;
  assign \new_[18376]_  = ~\new_[19308]_ ;
  assign n8484 = m7_s4_cyc_o_reg;
  assign n8554 = m7_s15_cyc_o_reg;
  assign n8309 = m6_s15_cyc_o_reg;
  assign \new_[18380]_  = ~\new_[20323]_  | ~\new_[29869]_ ;
  assign \new_[18381]_  = ~\new_[22355]_  | ~\new_[28278]_ ;
  assign \new_[18382]_  = ~\new_[30784]_  | ~\new_[5992]_  | ~\new_[29987]_  | ~\new_[21538]_ ;
  assign \new_[18383]_  = ~\new_[28905]_  | ~\new_[5988]_  | ~\new_[28595]_  | ~\new_[21506]_ ;
  assign \new_[18384]_  = ~\new_[30021]_  | ~\new_[6006]_  | ~\new_[29151]_  | ~\new_[20523]_ ;
  assign \new_[18385]_  = ~\new_[5894]_  | ~\new_[28271]_  | ~\new_[29119]_ ;
  assign \new_[18386]_  = ~\new_[5898]_  | ~\new_[30412]_  | ~\new_[28899]_ ;
  assign \new_[18387]_  = ~\new_[31491]_  | ~\new_[27792]_  | ~\new_[29750]_ ;
  assign n8799 = m6_s1_cyc_o_reg;
  assign \new_[18389]_  = ~\new_[5900]_  | ~\new_[26904]_  | ~\new_[28982]_ ;
  assign \new_[18390]_  = ~\new_[5901]_  | ~\new_[29330]_  | ~\new_[29331]_ ;
  assign n8664 = m4_s1_cyc_o_reg;
  assign \new_[18392]_  = ~\new_[5902]_  | ~\new_[30345]_  | ~\new_[29573]_ ;
  assign n8334 = m1_s1_cyc_o_reg;
  assign n8864 = m3_s0_cyc_o_reg;
  assign n8709 = m0_s1_cyc_o_reg;
  assign \new_[18396]_  = ~\new_[5907]_  | ~\new_[28242]_  | ~\new_[29096]_ ;
  assign \new_[18397]_  = ~\new_[31789]_  | ~\new_[27691]_  | ~\new_[28535]_ ;
  assign \new_[18398]_  = ~\new_[31235]_  | ~\new_[28332]_  | ~\new_[28402]_ ;
  assign \new_[18399]_  = ~\new_[6183]_  | ~\new_[29542]_  | ~\new_[29367]_ ;
  assign \new_[18400]_  = \new_[29840]_  & \new_[26571]_ ;
  assign \new_[18401]_  = ~\new_[5933]_  | ~\new_[27379]_  | ~\new_[28950]_ ;
  assign \new_[18402]_  = ~\new_[19378]_ ;
  assign \new_[18403]_  = ~\new_[5908]_  | ~\new_[27974]_  | ~\new_[29166]_ ;
  assign \new_[18404]_  = ~\new_[5913]_  | ~\new_[28093]_  | ~\new_[30236]_ ;
  assign \new_[18405]_  = ~\new_[6176]_  | ~\new_[28192]_  | ~\new_[28816]_ ;
  assign \new_[18406]_  = ~\new_[6190]_  | ~\new_[28671]_  | ~\new_[29290]_ ;
  assign \new_[18407]_  = \new_[20471]_  | \new_[30144]_ ;
  assign \new_[18408]_  = ~\new_[5830]_  | ~\new_[29756]_  | ~\new_[28232]_ ;
  assign \new_[18409]_  = ~\new_[5830]_  | ~\new_[29616]_  | ~\new_[30206]_ ;
  assign \new_[18410]_  = \new_[20497]_  | \new_[28804]_ ;
  assign \new_[18411]_  = ~\new_[5981]_  | ~\new_[29858]_  | ~\new_[30251]_ ;
  assign \new_[18412]_  = ~\new_[5968]_  | ~\new_[28961]_  | ~\new_[29848]_ ;
  assign \new_[18413]_  = ~\new_[5985]_  | ~\new_[28082]_  | ~\new_[30308]_ ;
  assign \new_[18414]_  = \new_[20468]_  | \new_[29125]_ ;
  assign \new_[18415]_  = ~\new_[5996]_  | ~\new_[30220]_  | ~\new_[28052]_ ;
  assign \new_[18416]_  = ~\new_[5999]_  | ~\new_[28224]_  | ~\new_[28999]_ ;
  assign \new_[18417]_  = \new_[19965]_  | \new_[28043]_ ;
  assign \new_[18418]_  = \new_[20467]_  | \new_[28189]_ ;
  assign \new_[18419]_  = ~\new_[5931]_  | ~\new_[29686]_  | ~\new_[30078]_ ;
  assign \new_[18420]_  = ~\new_[30305]_  | ~\new_[6091]_ ;
  assign \new_[18421]_  = ~\new_[27778]_  | ~\new_[6086]_ ;
  assign \new_[18422]_  = ~\new_[29300]_  | ~\new_[5920]_ ;
  assign \new_[18423]_  = ~\new_[27778]_  | ~\new_[5929]_ ;
  assign \new_[18424]_  = ~\new_[28718]_  | ~\new_[5972]_ ;
  assign \new_[18425]_  = ~\new_[26842]_  | ~\new_[5970]_ ;
  assign \new_[18426]_  = ~\new_[30339]_  | ~\new_[6087]_ ;
  assign \new_[18427]_  = ~\new_[30219]_  | ~\new_[6056]_ ;
  assign \new_[18428]_  = ~\new_[30087]_  | ~\new_[6062]_ ;
  assign \new_[18429]_  = ~\new_[26638]_  | ~\new_[6194]_ ;
  assign \new_[18430]_  = ~\new_[26638]_  | ~\new_[5984]_ ;
  assign \new_[18431]_  = ~\new_[26842]_  | ~\new_[6199]_ ;
  assign \new_[18432]_  = ~\new_[19471]_  | ~\new_[29794]_ ;
  assign \new_[18433]_  = ~\new_[19479]_  | ~\new_[30160]_ ;
  assign \new_[18434]_  = ~\new_[19480]_  | ~\new_[30146]_ ;
  assign \new_[18435]_  = ~\new_[19489]_  | ~\new_[30349]_ ;
  assign \new_[18436]_  = ~\new_[19482]_  | ~\new_[29877]_ ;
  assign \new_[18437]_  = ~\new_[19484]_  | ~\new_[30071]_ ;
  assign \new_[18438]_  = ~\new_[19493]_  | ~\new_[30278]_ ;
  assign \new_[18439]_  = ~\new_[19491]_  | ~\new_[30218]_ ;
  assign \new_[18440]_  = ~\new_[19495]_  | ~\new_[29897]_ ;
  assign \new_[18441]_  = ~\new_[19470]_  & ~\new_[30259]_ ;
  assign \new_[18442]_  = ~\new_[30726]_  | (~\new_[20956]_  & ~\new_[21597]_ );
  assign \new_[18443]_  = ~\new_[30296]_  | (~\new_[20742]_  & ~\new_[21598]_ );
  assign \new_[18444]_  = ~\new_[29219]_  | (~\new_[20753]_  & ~\new_[20587]_ );
  assign \new_[18445]_  = ~\new_[30426]_  | (~\new_[20759]_  & ~\new_[21599]_ );
  assign \new_[18446]_  = ~\new_[30750]_  | (~\new_[21698]_  & ~\new_[20596]_ );
  assign \new_[18447]_  = ~\new_[30550]_  | (~\new_[21699]_  & ~\new_[20597]_ );
  assign \new_[18448]_  = ~\new_[30721]_  | (~\new_[20792]_  & ~\new_[20602]_ );
  assign \new_[18449]_  = ~\new_[30410]_  | (~\new_[20849]_  & ~\new_[20603]_ );
  assign \new_[18450]_  = ~\new_[30617]_  | (~\new_[20812]_  & ~\new_[20674]_ );
  assign \new_[18451]_  = ~\new_[26270]_  & (~\new_[20558]_  | ~\new_[27914]_ );
  assign \new_[18452]_  = ~\new_[30651]_  & (~\new_[20562]_  | ~\new_[28524]_ );
  assign \new_[18453]_  = ~\new_[30574]_  | (~\new_[20793]_  & ~\new_[20613]_ );
  assign \new_[18454]_  = ~\new_[28967]_  | (~\new_[20789]_  & ~\new_[20601]_ );
  assign \new_[18455]_  = ~\new_[30765]_  | (~\new_[21825]_  & ~\new_[20615]_ );
  assign \new_[18456]_  = ~\new_[29978]_  | (~\new_[21815]_  & ~\new_[20616]_ );
  assign \new_[18457]_  = ~\new_[30107]_  | (~\new_[20840]_  & ~\new_[20619]_ );
  assign \new_[18458]_  = ~\new_[28188]_  | (~\new_[20740]_  & ~\new_[20628]_ );
  assign \new_[18459]_  = ~\new_[19492]_  & ~\new_[29453]_ ;
  assign \new_[18460]_  = ~\new_[30789]_  | (~\new_[21846]_  & ~\new_[20627]_ );
  assign \new_[18461]_  = ~\new_[29972]_  | (~\new_[21953]_  & ~\new_[20626]_ );
  assign \new_[18462]_  = ~\new_[29996]_  | (~\new_[20955]_  & ~\new_[20635]_ );
  assign \new_[18463]_  = ~\new_[19483]_  & ~\new_[30254]_ ;
  assign \new_[18464]_  = ~\new_[19498]_  | ~\new_[28524]_ ;
  assign \new_[18465]_  = ~\new_[20544]_  | ~\new_[31517]_  | ~n8869;
  assign \new_[18466]_  = ~\new_[20568]_  | ~\new_[31466]_  | ~n8829;
  assign \new_[18467]_  = ~\new_[20552]_  | ~\new_[31380]_  | ~n8744;
  assign \new_[18468]_  = ~\new_[20578]_  | ~\new_[31392]_  | ~n8784;
  assign \new_[18469]_  = ~\new_[20576]_  | ~\new_[31519]_  | ~n8874;
  assign \new_[18470]_  = ~\new_[20547]_  | ~\new_[31295]_  | ~n8559;
  assign \new_[18471]_  = ~\new_[20555]_  | ~\new_[31261]_  | ~n8499;
  assign \new_[18472]_  = ~\new_[20567]_  | ~\new_[31279]_  | ~n8504;
  assign \new_[18473]_  = ~\new_[20542]_  | ~\new_[31503]_  | ~n8839;
  assign \new_[18474]_  = ~\new_[20551]_  | ~\new_[31513]_  | ~n8854;
  assign \new_[18475]_  = ~\new_[20575]_  | ~\new_[31285]_  | ~n8519;
  assign \new_[18476]_  = ~\new_[20580]_  | ~\new_[31533]_  | ~n8929;
  assign \new_[18477]_  = ~\new_[20572]_  | ~\new_[31246]_  | ~n8464;
  assign n8794 = m0_s13_cyc_o_reg;
  assign n8439 = m0_s15_cyc_o_reg;
  assign n8904 = m0_s7_cyc_o_reg;
  assign n8304 = m4_s6_cyc_o_reg;
  assign n8319 = m5_s5_cyc_o_reg;
  assign \new_[18483]_  = \new_[20663]_  | \new_[30042]_ ;
  assign \new_[18484]_  = ~\new_[20592]_  & ~\new_[21121]_ ;
  assign \new_[18485]_  = ~\new_[20639]_  & ~\new_[23355]_ ;
  assign \new_[18486]_  = \new_[20640]_  | \new_[30541]_ ;
  assign \new_[18487]_  = \new_[20642]_  | \new_[30420]_ ;
  assign \new_[18488]_  = \new_[20644]_  | \new_[30648]_ ;
  assign \new_[18489]_  = \new_[20647]_  | \new_[29926]_ ;
  assign \new_[18490]_  = \new_[20681]_  | \new_[29777]_ ;
  assign \new_[18491]_  = ~\new_[20654]_  & ~\new_[22112]_ ;
  assign \new_[18492]_  = \new_[20652]_  | \new_[29828]_ ;
  assign \new_[18493]_  = \new_[20641]_  | \new_[30002]_ ;
  assign \new_[18494]_  = \new_[20651]_  | \new_[30553]_ ;
  assign \new_[18495]_  = ~\new_[20656]_  & ~\new_[23631]_ ;
  assign \new_[18496]_  = \new_[20655]_  | \new_[29790]_ ;
  assign \new_[18497]_  = ~\new_[20657]_  & ~\new_[25115]_ ;
  assign \new_[18498]_  = \new_[20659]_  | \new_[30466]_ ;
  assign \new_[18499]_  = ~\new_[20662]_  & ~\new_[23164]_ ;
  assign \new_[18500]_  = ~\new_[20582]_  & ~\new_[23170]_ ;
  assign \new_[18501]_  = ~\new_[24794]_  & (~\new_[21632]_  | ~\new_[26674]_ );
  assign \new_[18502]_  = ~\new_[28555]_  | (~\new_[21787]_  & ~\new_[30230]_ );
  assign \new_[18503]_  = ~\new_[28644]_  | ~\new_[20664]_  | ~\new_[24797]_ ;
  assign \new_[18504]_  = ~\new_[20610]_  & ~\new_[23491]_ ;
  assign \new_[18505]_  = ~\new_[28555]_  | ~\new_[20665]_  | ~\new_[23830]_ ;
  assign \new_[18506]_  = ~\new_[24601]_  & (~\new_[21638]_  | ~\new_[27573]_ );
  assign \new_[18507]_  = \new_[20697]_  | \new_[28503]_ ;
  assign \new_[18508]_  = ~\new_[20574]_  | ~\new_[27463]_ ;
  assign \new_[18509]_  = \new_[20722]_  & \new_[28527]_ ;
  assign \new_[18510]_  = ~\new_[26513]_  & (~\new_[21643]_  | ~\new_[29550]_ );
  assign \new_[18511]_  = ~\new_[20520]_  & ~\new_[24989]_ ;
  assign \new_[18512]_  = ~\new_[28495]_  & (~\new_[21648]_  | ~\new_[28069]_ );
  assign \new_[18513]_  = ~\new_[28398]_  & (~\new_[21649]_  | ~\new_[30582]_ );
  assign \new_[18514]_  = ~\new_[20585]_  | ~\new_[31853]_ ;
  assign \new_[18515]_  = ~\new_[20586]_  & ~\new_[24820]_ ;
  assign \new_[18516]_  = ~\new_[21267]_  & (~\new_[21992]_  | ~\new_[30030]_ );
  assign \new_[18517]_  = ~\new_[20588]_  & ~\new_[25031]_ ;
  assign \new_[18518]_  = ~\new_[22124]_  & (~\new_[21792]_  | ~\new_[22974]_ );
  assign \new_[18519]_  = \new_[20705]_  | \new_[30336]_ ;
  assign \new_[18520]_  = ~\new_[25439]_  & (~\new_[21662]_  | ~\new_[29079]_ );
  assign \new_[18521]_  = ~\new_[28727]_  & (~\new_[21821]_  | ~\new_[29219]_ );
  assign \new_[18522]_  = \new_[20702]_  & \new_[28586]_ ;
  assign \new_[18523]_  = ~\new_[20589]_  & ~\new_[26518]_ ;
  assign \new_[18524]_  = ~\new_[24869]_  & (~\new_[21667]_  | ~\new_[24401]_ );
  assign \new_[18525]_  = ~\new_[27572]_  & (~\new_[21672]_  | ~\new_[30135]_ );
  assign \new_[18526]_  = ~\new_[23647]_  & (~\new_[21708]_  | ~\new_[24416]_ );
  assign \new_[18527]_  = ~\new_[26673]_  & (~\new_[21677]_  | ~\new_[30842]_ );
  assign \new_[18528]_  = ~\new_[20593]_  & ~\new_[24839]_ ;
  assign \new_[18529]_  = ~\new_[21301]_  & (~\new_[21996]_  | ~\new_[28872]_ );
  assign \new_[18530]_  = ~\new_[23404]_  & (~\new_[21801]_  | ~\new_[22957]_ );
  assign \new_[18531]_  = ~\new_[26893]_  & (~\new_[21689]_  | ~\new_[26556]_ );
  assign \new_[18532]_  = ~\new_[20546]_  | ~\new_[26328]_ ;
  assign \new_[18533]_  = \new_[20704]_  & \new_[26901]_ ;
  assign \new_[18534]_  = ~\new_[26381]_  & (~\new_[21701]_  | ~\new_[30550]_ );
  assign \new_[18535]_  = \new_[20710]_  & \new_[29454]_ ;
  assign \new_[18536]_  = \new_[20695]_  | \new_[26228]_ ;
  assign \new_[18537]_  = ~\new_[27388]_  & (~\new_[21712]_  | ~\new_[28967]_ );
  assign \new_[18538]_  = ~\new_[20599]_  & ~\new_[24881]_ ;
  assign \new_[18539]_  = ~\new_[21270]_  & (~\new_[21999]_  | ~\new_[30057]_ );
  assign \new_[18540]_  = ~\new_[27481]_  & (~\new_[21686]_  | ~\new_[29780]_ );
  assign \new_[18541]_  = \new_[20594]_  | \new_[22987]_ ;
  assign \new_[18542]_  = ~\new_[21276]_  & (~\new_[22009]_  | ~\new_[28887]_ );
  assign \new_[18543]_  = ~\new_[25460]_  & (~\new_[21724]_  | ~\new_[30410]_ );
  assign \new_[18544]_  = \new_[20706]_  & \new_[28218]_ ;
  assign \new_[18545]_  = ~\new_[20548]_  | ~\new_[26355]_ ;
  assign \new_[18546]_  = ~\new_[20606]_  & ~\new_[24885]_ ;
  assign \new_[18547]_  = ~\new_[27601]_  & (~\new_[21745]_  | ~\new_[26655]_ );
  assign \new_[18548]_  = ~\new_[21324]_  & (~\new_[22001]_  | ~\new_[28883]_ );
  assign \new_[18549]_  = ~\new_[28231]_  | (~\new_[21729]_  & ~\new_[30093]_ );
  assign \new_[18550]_  = ~\new_[28231]_  | ~\new_[20670]_  | ~\new_[22350]_ ;
  assign \new_[18551]_  = \new_[20691]_  | \new_[26385]_ ;
  assign \new_[18552]_  = ~\new_[20565]_  | ~\new_[27640]_ ;
  assign \new_[18553]_  = ~s10_ack_i | ~\new_[20551]_  | ~\new_[30227]_ ;
  assign \new_[18554]_  = ~\new_[24744]_  & (~\new_[23032]_  | ~\new_[29922]_ );
  assign \new_[18555]_  = ~s10_err_i | ~\new_[20551]_  | ~\new_[30227]_ ;
  assign \new_[18556]_  = \new_[20707]_  & \new_[28540]_ ;
  assign \new_[18557]_  = ~s10_rty_i | ~\new_[20551]_  | ~\new_[30227]_ ;
  assign \new_[18558]_  = ~\new_[20629]_  | ~\new_[31888]_ ;
  assign \new_[18559]_  = \new_[20554]_  | \new_[23901]_ ;
  assign \new_[18560]_  = ~s7_ack_i | ~\new_[20555]_  | ~\new_[30193]_ ;
  assign \new_[18561]_  = ~\new_[27937]_  & (~\new_[21752]_  | ~\new_[30146]_ );
  assign \new_[18562]_  = \new_[20714]_  | \new_[30038]_ ;
  assign \new_[18563]_  = ~\new_[26426]_  & (~\new_[21753]_  | ~\new_[29892]_ );
  assign \new_[18564]_  = ~s7_err_i | ~\new_[20555]_  | ~\new_[30193]_ ;
  assign \new_[18565]_  = ~\new_[27976]_  & (~\new_[21743]_  | ~\new_[30207]_ );
  assign \new_[18566]_  = ~\new_[26979]_  & (~\new_[21757]_  | ~\new_[30432]_ );
  assign \new_[18567]_  = \new_[20709]_  & \new_[28144]_ ;
  assign \new_[18568]_  = ~\new_[24273]_  & (~\new_[21761]_  | ~\new_[28806]_ );
  assign \new_[18569]_  = ~s7_rty_i | ~\new_[20555]_  | ~\new_[30193]_ ;
  assign \new_[18570]_  = ~\new_[23527]_  & (~\new_[21952]_  | ~\new_[24421]_ );
  assign \new_[18571]_  = ~\new_[23947]_  & (~\new_[22047]_  | ~\new_[28962]_ );
  assign \new_[18572]_  = ~\new_[28494]_  | (~\new_[21904]_  & ~\new_[30199]_ );
  assign \new_[18573]_  = ~\new_[20557]_  | ~\new_[27525]_ ;
  assign \new_[18574]_  = ~\new_[27610]_  & (~\new_[21760]_  | ~\new_[29221]_ );
  assign \new_[18575]_  = ~\new_[20609]_  & ~\new_[25058]_ ;
  assign \new_[18576]_  = ~\new_[27581]_  & (~\new_[21858]_  | ~\new_[30294]_ );
  assign \new_[18577]_  = \new_[20580]_  & \new_[29205]_ ;
  assign \new_[18578]_  = \new_[20539]_  & \new_[29215]_ ;
  assign \new_[18579]_  = ~\new_[20622]_  & ~\new_[23566]_ ;
  assign \new_[18580]_  = ~\new_[23914]_  & (~\new_[21596]_  | ~\new_[29202]_ );
  assign \new_[18581]_  = ~\new_[28416]_  | (~\new_[21781]_  & ~\new_[30254]_ );
  assign \new_[18582]_  = ~\new_[27633]_  | ~\new_[20677]_  | ~\new_[24954]_ ;
  assign \new_[18583]_  = ~\new_[28416]_  | ~\new_[20678]_  | ~\new_[23616]_ ;
  assign \new_[18584]_  = \new_[20694]_  | \new_[26421]_ ;
  assign \new_[18585]_  = \new_[20711]_  | \new_[30029]_ ;
  assign \new_[18586]_  = \new_[20693]_  | \new_[29624]_ ;
  assign \new_[18587]_  = ~\new_[20614]_  & ~\new_[24964]_ ;
  assign \new_[18588]_  = ~\new_[25102]_  & (~\new_[21894]_  | ~\new_[26244]_ );
  assign \new_[18589]_  = ~\new_[26394]_  & (~\new_[22677]_  | ~\new_[29064]_ );
  assign \new_[18590]_  = ~\new_[26804]_  & (~\new_[21802]_  | ~\new_[29978]_ );
  assign \new_[18591]_  = ~\new_[27905]_  & (~\new_[21804]_  | ~\new_[29877]_ );
  assign \new_[18592]_  = ~\new_[21314]_  & (~\new_[22016]_  | ~\new_[29268]_ );
  assign \new_[18593]_  = \new_[20713]_  & \new_[29499]_ ;
  assign \new_[18594]_  = ~\new_[27991]_  & (~\new_[21706]_  | ~\new_[30491]_ );
  assign \new_[18595]_  = ~\new_[20566]_  | ~\new_[26226]_ ;
  assign \new_[18596]_  = ~\new_[23997]_  & (~\new_[21642]_  | ~\new_[29656]_ );
  assign \new_[18597]_  = ~\new_[27860]_  & (~\new_[21864]_  | ~\new_[30034]_ );
  assign \new_[18598]_  = ~\new_[23567]_  & (~\new_[21777]_  | ~\new_[23254]_ );
  assign \new_[18599]_  = ~\new_[21315]_  & (~\new_[22011]_  | ~\new_[28924]_ );
  assign \new_[18600]_  = \new_[20717]_  & \new_[29460]_ ;
  assign \new_[18601]_  = ~\new_[26769]_  | (~\new_[21828]_  & ~\new_[30130]_ );
  assign \new_[18602]_  = ~\new_[24704]_  & (~\new_[21834]_  | ~\new_[28935]_ );
  assign \new_[18603]_  = ~\new_[25065]_  & (~\new_[21705]_  | ~\new_[30138]_ );
  assign \new_[18604]_  = ~\new_[26976]_  & (~\new_[21844]_  | ~\new_[24499]_ );
  assign \new_[18605]_  = \new_[20692]_  | \new_[27616]_ ;
  assign \new_[18606]_  = ~\new_[20577]_  | ~\new_[24792]_ ;
  assign \new_[18607]_  = ~\new_[28800]_  & (~\new_[21950]_  | ~\new_[29972]_ );
  assign \new_[18608]_  = ~\new_[23761]_  & (~\new_[21912]_  | ~\new_[24520]_ );
  assign \new_[18609]_  = ~\new_[23384]_  & (~\new_[21945]_  | ~\new_[24498]_ );
  assign \new_[18610]_  = ~\new_[27614]_  & (~\new_[21850]_  | ~\new_[30160]_ );
  assign \new_[18611]_  = \new_[20720]_  & \new_[27648]_ ;
  assign \new_[18612]_  = ~\new_[20561]_  & (~\new_[22018]_  | ~\new_[29248]_ );
  assign \new_[18613]_  = ~\new_[26734]_  & (~\new_[21771]_  | ~\new_[30218]_ );
  assign \new_[18614]_  = ~\new_[20623]_  & ~\new_[23827]_ ;
  assign \new_[18615]_  = ~\new_[24854]_  & (~\new_[21714]_  | ~\new_[30437]_ );
  assign \new_[18616]_  = ~\new_[28654]_  & (~\new_[21735]_  | ~\new_[30727]_ );
  assign \new_[18617]_  = ~\new_[23905]_  & (~\new_[22010]_  | ~\new_[29744]_ );
  assign \new_[18618]_  = \new_[20696]_  | \new_[27643]_ ;
  assign \new_[18619]_  = ~\new_[26934]_  & (~\new_[21979]_  | ~\new_[26318]_ );
  assign \new_[18620]_  = ~\new_[28494]_  | ~\new_[20676]_  | ~\new_[22242]_ ;
  assign \new_[18621]_  = ~\new_[24008]_  & (~\new_[21641]_  | ~\new_[30221]_ );
  assign \new_[18622]_  = ~\new_[26730]_  & (~\new_[21840]_  | ~\new_[30205]_ );
  assign \new_[18623]_  = ~\new_[28233]_  & (~\new_[22199]_  | ~\new_[29537]_ );
  assign \new_[18624]_  = \new_[20721]_  & \new_[28838]_ ;
  assign \new_[18625]_  = ~\new_[20632]_  & ~\new_[23526]_ ;
  assign \new_[18626]_  = ~\new_[26488]_  & (~\new_[21959]_  | ~\new_[27727]_ );
  assign \new_[18627]_  = ~\new_[20633]_  & ~\new_[23842]_ ;
  assign \new_[18628]_  = ~\new_[23843]_  & (~\new_[21970]_  | ~\new_[24312]_ );
  assign \new_[18629]_  = ~\new_[23951]_  & (~\new_[21998]_  | ~\new_[29350]_ );
  assign \new_[18630]_  = ~\new_[27583]_  & (~\new_[21973]_  | ~\new_[29897]_ );
  assign \new_[18631]_  = ~\new_[28368]_  | (~\new_[21974]_  & ~\new_[30047]_ );
  assign \new_[18632]_  = ~\new_[28368]_  | ~\new_[20689]_  | ~\new_[22441]_ ;
  assign \new_[18633]_  = \new_[20698]_  | \new_[26231]_ ;
  assign \new_[18634]_  = ~\new_[24662]_  & (~\new_[21967]_  | ~\new_[29701]_ );
  assign \new_[18635]_  = ~\new_[26752]_  & (~\new_[21978]_  | ~\new_[30025]_ );
  assign \new_[18636]_  = \new_[20724]_  & \new_[28569]_ ;
  assign \new_[18637]_  = ~\new_[21294]_  & (~\new_[22076]_  | ~\new_[28939]_ );
  assign \new_[18638]_  = ~\new_[28229]_  & (~\new_[21982]_  | ~\new_[30735]_ );
  assign \new_[18639]_  = ~\new_[28092]_  & (~\new_[21915]_  | ~\new_[30764]_ );
  assign \new_[18640]_  = ~\new_[20637]_  | ~\new_[31804]_ ;
  assign \new_[18641]_  = \new_[20679]_  | \new_[26421]_ ;
  assign \new_[18642]_  = ~\new_[27650]_  & (~\new_[21636]_  | ~\new_[30152]_ );
  assign \new_[18643]_  = ~\new_[26541]_  & (~\new_[21687]_  | ~\new_[29746]_ );
  assign \new_[18644]_  = \new_[20672]_  | \new_[24063]_ ;
  assign \new_[18645]_  = \new_[20686]_  | \new_[26228]_ ;
  assign \new_[18646]_  = ~\new_[28296]_  & (~\new_[21841]_  | ~\new_[30444]_ );
  assign \new_[18647]_  = \new_[20685]_  | \new_[27616]_ ;
  assign \new_[18648]_  = \new_[20675]_  | \new_[27643]_ ;
  assign \new_[18649]_  = ~\new_[28486]_  & (~\new_[21928]_  | ~\new_[30786]_ );
  assign \new_[18650]_  = ~\new_[25213]_  & (~\new_[21956]_  | ~\new_[28964]_ );
  assign \new_[18651]_  = ~\new_[26379]_  & (~\new_[21980]_  | ~\new_[29900]_ );
  assign \new_[18652]_  = ~s7_ack_i | ~\new_[20542]_  | ~\new_[30060]_ ;
  assign \new_[18653]_  = ~s4_ack_i | ~\new_[20544]_  | ~\new_[29628]_ ;
  assign \new_[18654]_  = ~s4_err_i | ~\new_[20544]_  | ~\new_[29628]_ ;
  assign \new_[18655]_  = ~s7_err_i | ~\new_[20542]_  | ~\new_[30060]_ ;
  assign \new_[18656]_  = ~s4_rty_i | ~\new_[20544]_  | ~\new_[29628]_ ;
  assign \new_[18657]_  = ~\new_[29749]_  | ~\new_[20547]_  | ~s10_ack_i;
  assign \new_[18658]_  = ~\new_[30225]_  & (~\new_[22103]_  | ~\new_[29577]_ );
  assign \new_[18659]_  = \new_[20545]_  & \new_[29711]_ ;
  assign \new_[18660]_  = \new_[20547]_  & \new_[29749]_ ;
  assign \new_[18661]_  = \new_[20578]_  & \new_[29649]_ ;
  assign \new_[18662]_  = ~s4_ack_i | ~\new_[20568]_  | ~\new_[29961]_ ;
  assign \new_[18663]_  = ~s4_err_i | ~\new_[20568]_  | ~\new_[29961]_ ;
  assign \new_[18664]_  = ~s4_rty_i | ~\new_[20568]_  | ~\new_[29961]_ ;
  assign \new_[18665]_  = ~s10_ack_i | ~\new_[20575]_  | ~\new_[29705]_ ;
  assign \new_[18666]_  = ~s10_err_i | ~\new_[20575]_  | ~\new_[29705]_ ;
  assign \new_[18667]_  = ~s10_rty_i | ~\new_[20575]_  | ~\new_[29705]_ ;
  assign \new_[18668]_  = ~s7_rty_i | ~\new_[20567]_  | ~\new_[30131]_ ;
  assign \new_[18669]_  = \new_[22110]_  | \new_[20699]_ ;
  assign \new_[18670]_  = \new_[22126]_  | \new_[20701]_ ;
  assign \new_[18671]_  = \new_[21663]_  | \new_[20666]_ ;
  assign \new_[18672]_  = ~\new_[29026]_  | ~\new_[20667]_  | ~\new_[23705]_ ;
  assign \new_[18673]_  = ~\new_[27730]_  | ~\new_[20673]_  | ~\new_[24922]_ ;
  assign \new_[18674]_  = \new_[22145]_  | \new_[20703]_ ;
  assign \new_[18675]_  = \new_[20861]_  | \new_[20668]_ ;
  assign \new_[18676]_  = ~\new_[29454]_  | ~\new_[20669]_  | ~\new_[22238]_ ;
  assign \new_[18677]_  = \new_[22161]_  | \new_[20716]_ ;
  assign \new_[18678]_  = ~\new_[30293]_  | ~\new_[20708]_  | ~\new_[27730]_ ;
  assign \new_[18679]_  = \new_[22179]_  | \new_[20719]_ ;
  assign \new_[18680]_  = \new_[21731]_  | \new_[20671]_ ;
  assign \new_[18681]_  = ~\new_[29499]_  | ~\new_[20680]_  | ~\new_[23623]_ ;
  assign \new_[18682]_  = \new_[22142]_  | \new_[20725]_ ;
  assign \new_[18683]_  = \new_[23649]_  | \new_[20715]_ ;
  assign \new_[18684]_  = \new_[21227]_  | \new_[21621]_ ;
  assign \new_[18685]_  = \new_[20954]_  | \new_[20684]_ ;
  assign \new_[18686]_  = ~\new_[28838]_  | ~\new_[20688]_  | ~\new_[25011]_ ;
  assign \new_[18687]_  = \new_[21944]_  | \new_[20682]_ ;
  assign \new_[18688]_  = \new_[23831]_  | \new_[20712]_ ;
  assign \new_[18689]_  = \new_[22448]_  | \new_[20723]_ ;
  assign \new_[18690]_  = ~\new_[28569]_  | ~\new_[20690]_  | ~\new_[23864]_ ;
  assign \new_[18691]_  = ~\new_[21816]_  | (~\new_[22080]_  & ~\new_[30334]_ );
  assign \new_[18692]_  = ~\new_[23206]_  | (~\new_[22081]_  & ~\new_[30747]_ );
  assign \new_[18693]_  = ~\new_[21838]_  | (~\new_[22082]_  & ~\new_[30616]_ );
  assign \new_[18694]_  = ~\new_[21897]_  | (~\new_[22096]_  & ~\new_[30688]_ );
  assign \new_[18695]_  = ~\new_[21898]_  | (~\new_[22097]_  & ~\new_[30632]_ );
  assign \new_[18696]_  = ~\new_[21808]_  | (~\new_[22085]_  & ~\new_[30684]_ );
  assign \new_[18697]_  = ~\new_[21824]_  | (~\new_[22086]_  & ~\new_[29934]_ );
  assign \new_[18698]_  = ~\new_[21929]_  | (~\new_[22087]_  & ~\new_[30637]_ );
  assign \new_[18699]_  = ~\new_[21958]_  | (~\new_[22088]_  & ~\new_[29652]_ );
  assign \new_[18700]_  = ~\new_[21675]_  | (~\new_[22099]_  & ~\new_[30607]_ );
  assign \new_[18701]_  = ~\new_[29029]_  | ~\new_[20529]_  | ~\new_[22111]_ ;
  assign \new_[18702]_  = ~\new_[29911]_  | ~\new_[20530]_  | ~\new_[24813]_ ;
  assign \new_[18703]_  = ~\new_[29781]_  | ~\new_[20532]_  | ~\new_[24997]_ ;
  assign \new_[18704]_  = ~\new_[30604]_  | ~\new_[20533]_  | ~\new_[23422]_ ;
  assign \new_[18705]_  = ~\new_[29763]_  | ~\new_[20534]_  | ~\new_[24880]_ ;
  assign \new_[18706]_  = ~\new_[30243]_  | ~\new_[20535]_  | ~\new_[24983]_ ;
  assign \new_[18707]_  = ~\new_[29505]_  | ~\new_[20536]_  | ~\new_[23655]_ ;
  assign \new_[18708]_  = ~\new_[30579]_  | ~\new_[20537]_  | ~\new_[26978]_ ;
  assign \new_[18709]_  = ~\new_[29768]_  | ~\new_[20538]_  | ~\new_[24620]_ ;
  assign \new_[18710]_  = ~\new_[21056]_  | ~\new_[30296]_ ;
  assign \new_[18711]_  = ~\new_[21090]_  | ~\new_[29219]_ ;
  assign \new_[18712]_  = ~\new_[21067]_  | ~\new_[28837]_ ;
  assign \new_[18713]_  = ~\new_[21061]_  | ~\new_[28989]_ ;
  assign \new_[18714]_  = ~\new_[21093]_  | ~\new_[29221]_ ;
  assign \new_[18715]_  = ~\new_[21072]_  | ~\new_[28967]_ ;
  assign \new_[18716]_  = ~\new_[21076]_  | ~\new_[29038]_ ;
  assign \new_[18717]_  = ~\new_[29974]_  | (~\new_[22371]_  & ~\new_[24430]_ );
  assign \new_[18718]_  = ~\new_[21081]_  | ~\new_[29355]_ ;
  assign \new_[18719]_  = ~\new_[21077]_  | ~\new_[30107]_ ;
  assign \new_[18720]_  = ~\new_[29912]_  | (~\new_[22262]_  & ~\new_[24374]_ );
  assign \new_[18721]_  = ~\new_[30702]_  | (~\new_[22431]_  & ~\new_[28135]_ );
  assign \new_[18722]_  = ~\new_[21084]_  | ~\new_[29082]_ ;
  assign \new_[18723]_  = ~\new_[21064]_  | ~\new_[28007]_ ;
  assign \new_[18724]_  = ~\new_[29685]_  | (~\new_[22410]_  & ~\new_[26414]_ );
  assign \new_[18725]_  = ~\new_[21106]_  | ~\new_[27593]_ ;
  assign \new_[18726]_  = ~\new_[21111]_  | ~\new_[27848]_ ;
  assign \new_[18727]_  = ~\new_[21100]_  | ~\new_[29996]_ ;
  assign \new_[18728]_  = ~\new_[21112]_  | ~\new_[27546]_ ;
  assign \new_[18729]_  = ~\new_[30150]_  | ~\new_[21988]_  | ~\new_[29900]_ ;
  assign \new_[18730]_  = ~\new_[29172]_  & (~\new_[22438]_  | ~\new_[25139]_ );
  assign \new_[18731]_  = ~\new_[19536]_ ;
  assign \new_[18732]_  = ~\new_[19536]_ ;
  assign \new_[18733]_  = ~\new_[19539]_ ;
  assign \new_[18734]_  = \new_[19539]_ ;
  assign \new_[18735]_  = ~\new_[25113]_  & ~\new_[20982]_ ;
  assign \new_[18736]_  = ~\new_[26956]_  | ~\new_[20963]_ ;
  assign \new_[18737]_  = \new_[26413]_  & \new_[20964]_ ;
  assign \new_[18738]_  = ~\new_[19540]_ ;
  assign \new_[18739]_  = \new_[25113]_  & \new_[20819]_ ;
  assign \new_[18740]_  = ~\new_[19541]_ ;
  assign \new_[18741]_  = ~\new_[23089]_  | ~\new_[20969]_ ;
  assign \new_[18742]_  = \new_[26517]_  & \new_[20961]_ ;
  assign \new_[18743]_  = ~\new_[19543]_ ;
  assign \new_[18744]_  = ~\new_[19543]_ ;
  assign \new_[18745]_  = ~\new_[23639]_  & ~\new_[20962]_ ;
  assign \new_[18746]_  = \new_[21095]_  & \new_[26905]_ ;
  assign \new_[18747]_  = ~\new_[19546]_ ;
  assign \new_[18748]_  = ~\new_[19546]_ ;
  assign \new_[18749]_  = ~\new_[19546]_ ;
  assign \new_[18750]_  = ~\new_[19546]_ ;
  assign \new_[18751]_  = ~\new_[19546]_ ;
  assign \new_[18752]_  = ~\new_[19546]_ ;
  assign \new_[18753]_  = ~\new_[19546]_ ;
  assign \new_[18754]_  = ~\new_[19546]_ ;
  assign \new_[18755]_  = ~\new_[19546]_ ;
  assign \new_[18756]_  = ~\new_[19546]_ ;
  assign \new_[18757]_  = ~\new_[19546]_ ;
  assign \new_[18758]_  = ~\new_[19546]_ ;
  assign \new_[18759]_  = ~\new_[19546]_ ;
  assign \new_[18760]_  = ~\new_[24610]_  & ~\new_[20960]_ ;
  assign \new_[18761]_  = ~\new_[19547]_ ;
  assign \new_[18762]_  = ~\new_[19548]_ ;
  assign \new_[18763]_  = ~\new_[19548]_ ;
  assign \new_[18764]_  = ~\new_[19548]_ ;
  assign \new_[18765]_  = ~\new_[19548]_ ;
  assign \new_[18766]_  = ~\new_[19548]_ ;
  assign \new_[18767]_  = ~\new_[19548]_ ;
  assign \new_[18768]_  = \new_[21068]_  & \new_[26693]_ ;
  assign \new_[18769]_  = ~\new_[30336]_  & (~\new_[22122]_  | ~\new_[26902]_ );
  assign \new_[18770]_  = \new_[21073]_  & \new_[26835]_ ;
  assign \new_[18771]_  = ~\new_[29798]_  | ~\new_[21053]_  | ~\new_[30262]_ ;
  assign \new_[18772]_  = ~\new_[19552]_ ;
  assign \new_[18773]_  = ~\new_[29320]_  | ~\new_[21995]_  | ~\new_[30320]_ ;
  assign \new_[18774]_  = ~\new_[29746]_  | ~\new_[21006]_  | ~\new_[29975]_ ;
  assign \new_[18775]_  = ~\new_[26203]_  & (~\new_[22150]_  | ~\new_[29350]_ );
  assign \new_[18776]_  = ~\new_[19554]_ ;
  assign \new_[18777]_  = \new_[21062]_  & \new_[26246]_ ;
  assign \new_[18778]_  = ~\new_[29456]_  | ~\new_[22002]_  | ~\new_[30159]_ ;
  assign \new_[18779]_  = ~\new_[29228]_  | ~\new_[22000]_  | ~\new_[30172]_ ;
  assign \new_[18780]_  = \new_[23441]_  | \new_[20791]_ ;
  assign \new_[18781]_  = ~\new_[19556]_ ;
  assign \new_[18782]_  = \new_[20527]_  & \new_[26223]_ ;
  assign \new_[18783]_  = ~\new_[30011]_  | ~\new_[21009]_  | ~\new_[30037]_ ;
  assign \new_[18784]_  = ~\new_[26517]_  & ~\new_[20830]_ ;
  assign \new_[18785]_  = \new_[25114]_  | \new_[20804]_ ;
  assign \new_[18786]_  = ~\new_[19558]_ ;
  assign \new_[18787]_  = \new_[24860]_  & \new_[20807]_ ;
  assign \new_[18788]_  = ~\new_[19559]_ ;
  assign \new_[18789]_  = ~\new_[19560]_ ;
  assign \new_[18790]_  = \new_[24907]_  & \new_[20811]_ ;
  assign \new_[18791]_  = ~\new_[19562]_ ;
  assign \new_[18792]_  = \new_[19562]_ ;
  assign \new_[18793]_  = ~\new_[19563]_ ;
  assign \new_[18794]_  = ~\new_[19564]_ ;
  assign \new_[18795]_  = ~\new_[19564]_ ;
  assign \new_[18796]_  = ~\new_[19565]_ ;
  assign \new_[18797]_  = ~\new_[19566]_ ;
  assign \new_[18798]_  = ~\new_[19567]_ ;
  assign \new_[18799]_  = \new_[19568]_ ;
  assign \new_[18800]_  = \new_[21091]_  & \new_[24445]_ ;
  assign \new_[18801]_  = ~\new_[23089]_  & ~\new_[20921]_ ;
  assign \new_[18802]_  = ~\new_[30130]_  & (~\new_[22301]_  | ~\new_[24909]_ );
  assign \new_[18803]_  = ~\new_[26517]_  & ~\new_[20825]_ ;
  assign \new_[18804]_  = ~\new_[19570]_ ;
  assign \new_[18805]_  = ~\new_[19570]_ ;
  assign \new_[18806]_  = ~\new_[23441]_  & ~\new_[20769]_ ;
  assign \new_[18807]_  = ~\new_[19571]_ ;
  assign \new_[18808]_  = \new_[23639]_  & \new_[20827]_ ;
  assign \new_[18809]_  = ~\new_[19572]_ ;
  assign \new_[18810]_  = ~\new_[19575]_ ;
  assign \new_[18811]_  = \new_[19575]_ ;
  assign \new_[18812]_  = ~\new_[29700]_  & (~\new_[22240]_  | ~\new_[23796]_ );
  assign \new_[18813]_  = ~\new_[19577]_ ;
  assign \new_[18814]_  = ~\new_[19577]_ ;
  assign \new_[18815]_  = \new_[21085]_  & \new_[28353]_ ;
  assign \new_[18816]_  = \new_[21071]_  & \new_[28419]_ ;
  assign \new_[18817]_  = ~\new_[19581]_ ;
  assign \new_[18818]_  = ~\new_[19581]_ ;
  assign \new_[18819]_  = \new_[19581]_ ;
  assign \new_[18820]_  = ~\new_[19581]_ ;
  assign \new_[18821]_  = ~\new_[23874]_  & ~\new_[20806]_ ;
  assign \new_[18822]_  = ~\new_[24732]_  & ~\new_[20806]_ ;
  assign \new_[18823]_  = ~\new_[26849]_  & ~\new_[20804]_ ;
  assign \new_[18824]_  = ~\new_[19583]_ ;
  assign \new_[18825]_  = ~\new_[19583]_ ;
  assign \new_[18826]_  = ~\new_[23639]_  & ~\new_[21734]_ ;
  assign \new_[18827]_  = ~\new_[19584]_ ;
  assign \new_[18828]_  = ~\new_[23441]_  | ~\new_[20808]_ ;
  assign \new_[18829]_  = ~\new_[19585]_ ;
  assign \new_[18830]_  = ~\new_[19585]_ ;
  assign \new_[18831]_  = ~\new_[19585]_ ;
  assign \new_[18832]_  = \new_[19586]_ ;
  assign \new_[18833]_  = ~\new_[19587]_ ;
  assign \new_[18834]_  = ~\new_[19588]_ ;
  assign \new_[18835]_  = ~\new_[19589]_ ;
  assign \new_[18836]_  = ~\new_[26956]_  & ~\new_[20805]_ ;
  assign \new_[18837]_  = ~\new_[19590]_ ;
  assign \new_[18838]_  = \new_[21092]_  & \new_[24613]_ ;
  assign \new_[18839]_  = ~\new_[30572]_  | ~\new_[21018]_  | ~\new_[29802]_ ;
  assign \new_[18840]_  = \new_[21070]_  & \new_[24378]_ ;
  assign \new_[18841]_  = ~\new_[25800]_  & (~\new_[22253]_  | ~\new_[29202]_ );
  assign \new_[18842]_  = ~\new_[29006]_  | ~\new_[22015]_  | ~\new_[29863]_ ;
  assign \new_[18843]_  = ~\new_[28762]_  | ~\new_[21022]_  | ~\new_[29979]_ ;
  assign \new_[18844]_  = \new_[21082]_  & \new_[27772]_ ;
  assign \new_[18845]_  = ~\new_[29047]_  & (~\new_[22168]_  | ~\new_[23763]_ );
  assign \new_[18846]_  = ~\new_[24610]_  & ~\new_[20829]_ ;
  assign \new_[18847]_  = \new_[21083]_  & \new_[26251]_ ;
  assign \new_[18848]_  = ~\new_[29671]_  & (~\new_[23823]_  | ~\new_[25039]_ );
  assign \new_[18849]_  = ~\new_[24830]_  & ~\new_[20921]_ ;
  assign \new_[18850]_  = ~\new_[24870]_  & ~\new_[20769]_ ;
  assign \new_[18851]_  = ~\new_[19595]_ ;
  assign \new_[18852]_  = ~\new_[19596]_ ;
  assign \new_[18853]_  = ~\new_[19596]_ ;
  assign \new_[18854]_  = ~\new_[19596]_ ;
  assign \new_[18855]_  = ~\new_[19598]_ ;
  assign \new_[18856]_  = ~\new_[19598]_ ;
  assign \new_[18857]_  = ~\new_[19598]_ ;
  assign \new_[18858]_  = ~\new_[19598]_ ;
  assign \new_[18859]_  = ~\new_[19599]_ ;
  assign \new_[18860]_  = ~\new_[19599]_ ;
  assign \new_[18861]_  = ~\new_[19599]_ ;
  assign \new_[18862]_  = ~\new_[19599]_ ;
  assign \new_[18863]_  = ~\new_[19600]_ ;
  assign \new_[18864]_  = ~\new_[19600]_ ;
  assign \new_[18865]_  = ~\new_[19600]_ ;
  assign \new_[18866]_  = ~\new_[19600]_ ;
  assign \new_[18867]_  = \new_[21097]_  & \new_[28065]_ ;
  assign \new_[18868]_  = \new_[21094]_  & \new_[24444]_ ;
  assign \new_[18869]_  = ~\new_[29527]_  | ~\new_[21991]_  | ~\new_[30097]_ ;
  assign \new_[18870]_  = ~\new_[30326]_  & (~\new_[22208]_  | ~\new_[24971]_ );
  assign \new_[18871]_  = ~\new_[19607]_ ;
  assign \new_[18872]_  = ~\new_[30717]_  | ~\new_[21013]_  | ~\new_[29870]_ ;
  assign \new_[18873]_  = ~\new_[28888]_  | ~\new_[21028]_  | ~\new_[29867]_ ;
  assign \new_[18874]_  = \new_[21101]_  & \new_[28289]_ ;
  assign \new_[18875]_  = \new_[23818]_  | \new_[20982]_ ;
  assign \new_[18876]_  = ~\new_[19609]_ ;
  assign \new_[18877]_  = ~\new_[19610]_ ;
  assign \new_[18878]_  = ~\new_[23848]_  & ~\new_[20960]_ ;
  assign \new_[18879]_  = \new_[24732]_  & \new_[21920]_ ;
  assign \new_[18880]_  = \new_[22128]_  & \new_[20969]_ ;
  assign \new_[18881]_  = \new_[23472]_  & \new_[20961]_ ;
  assign \new_[18882]_  = ~\new_[23488]_  & ~\new_[23252]_ ;
  assign \new_[18883]_  = ~\new_[19611]_ ;
  assign \new_[18884]_  = ~\new_[25999]_  & ~\new_[20962]_ ;
  assign \new_[18885]_  = ~\new_[19615]_ ;
  assign \new_[18886]_  = \new_[23529]_  & \new_[20964]_ ;
  assign \new_[18887]_  = ~\new_[19542]_ ;
  assign \new_[18888]_  = ~\new_[19617]_ ;
  assign \new_[18889]_  = ~\new_[19621]_ ;
  assign \new_[18890]_  = \new_[19621]_ ;
  assign \new_[18891]_  = ~\new_[19622]_ ;
  assign \new_[18892]_  = ~\new_[19622]_ ;
  assign \new_[18893]_  = ~\new_[19622]_ ;
  assign \new_[18894]_  = ~\new_[19622]_ ;
  assign \new_[18895]_  = ~\new_[19622]_ ;
  assign \new_[18896]_  = ~\new_[19622]_ ;
  assign \new_[18897]_  = ~\new_[19623]_ ;
  assign \new_[18898]_  = ~\new_[19623]_ ;
  assign \new_[18899]_  = ~\new_[19623]_ ;
  assign \new_[18900]_  = ~\new_[19623]_ ;
  assign \new_[18901]_  = ~\new_[19624]_ ;
  assign \new_[18902]_  = ~\new_[19627]_ ;
  assign \new_[18903]_  = ~\new_[19627]_ ;
  assign \new_[18904]_  = ~\new_[23818]_  | ~\new_[20819]_ ;
  assign \new_[18905]_  = \new_[19628]_ ;
  assign \new_[18906]_  = ~\new_[24870]_  & ~\new_[20791]_ ;
  assign \new_[18907]_  = ~\new_[19506]_ ;
  assign \new_[18908]_  = ~\new_[19506]_ ;
  assign \new_[18909]_  = ~\new_[19506]_ ;
  assign \new_[18910]_  = ~\new_[23472]_  & ~\new_[20830]_ ;
  assign \new_[18911]_  = \new_[21098]_  & \new_[25505]_ ;
  assign \new_[18912]_  = ~\new_[19631]_ ;
  assign \new_[18913]_  = ~\new_[19631]_ ;
  assign \new_[18914]_  = ~\new_[19632]_ ;
  assign \new_[18915]_  = ~\new_[19633]_ ;
  assign \new_[18916]_  = \new_[19633]_ ;
  assign \new_[18917]_  = \new_[19633]_ ;
  assign \new_[18918]_  = ~\new_[19634]_ ;
  assign \new_[18919]_  = ~\new_[19634]_ ;
  assign \new_[18920]_  = ~\new_[19634]_ ;
  assign \new_[18921]_  = ~\new_[19634]_ ;
  assign \new_[18922]_  = ~\new_[19634]_ ;
  assign \new_[18923]_  = ~\new_[19634]_ ;
  assign \new_[18924]_  = ~\new_[19634]_ ;
  assign \new_[18925]_  = ~\new_[19634]_ ;
  assign \new_[18926]_  = ~\new_[19634]_ ;
  assign \new_[18927]_  = ~\new_[23529]_  & ~\new_[20796]_ ;
  assign \new_[18928]_  = ~\new_[19635]_ ;
  assign \new_[18929]_  = ~\new_[19635]_ ;
  assign \new_[18930]_  = ~\new_[19635]_ ;
  assign \new_[18931]_  = ~\new_[19636]_ ;
  assign \new_[18932]_  = \new_[19637]_ ;
  assign \new_[18933]_  = ~\new_[19638]_ ;
  assign \new_[18934]_  = ~\new_[26571]_  & (~\new_[22318]_  | ~\new_[30363]_ );
  assign \new_[18935]_  = ~\new_[19639]_ ;
  assign \new_[18936]_  = \new_[25999]_  & \new_[20827]_ ;
  assign \new_[18937]_  = ~\new_[19641]_ ;
  assign \new_[18938]_  = ~\new_[30009]_  | ~\new_[22008]_  | ~\new_[28964]_ ;
  assign \new_[18939]_  = \new_[21087]_  & \new_[26285]_ ;
  assign \new_[18940]_  = ~\new_[19643]_ ;
  assign \new_[18941]_  = ~\new_[19647]_ ;
  assign \new_[18942]_  = \new_[23472]_  | \new_[20825]_ ;
  assign \new_[18943]_  = ~\new_[30555]_  | ~\new_[30697]_  | ~\new_[20758]_  | ~\new_[28057]_ ;
  assign \new_[18944]_  = ~\new_[30754]_  | ~\new_[28183]_  | ~\new_[20751]_  | ~\new_[27883]_ ;
  assign \new_[18945]_  = ~\new_[30774]_  | ~\new_[30022]_  | ~\new_[20727]_  | ~\new_[30497]_ ;
  assign \new_[18946]_  = ~\new_[30676]_  | ~\new_[29746]_  | ~\new_[20876]_  | ~\new_[30132]_ ;
  assign \new_[18947]_  = ~\new_[30434]_  | ~\new_[30552]_  | ~\new_[21629]_  | ~\new_[28806]_ ;
  assign \new_[18948]_  = ~\new_[30719]_  | ~\new_[30444]_  | ~\new_[20928]_  | ~\new_[30367]_ ;
  assign \new_[18949]_  = ~\new_[29233]_  | ~\new_[29593]_  | ~\new_[20728]_  | ~\new_[29831]_ ;
  assign \new_[18950]_  = ~\new_[30782]_  | ~\new_[30213]_  | ~\new_[20878]_  | ~\new_[29553]_ ;
  assign \new_[18951]_  = ~\new_[30574]_  | ~\new_[28039]_  | ~\new_[20726]_  | ~\new_[30329]_ ;
  assign \new_[18952]_  = ~\new_[30765]_  | ~\new_[29064]_  | ~\new_[21628]_  | ~\new_[30554]_ ;
  assign \new_[18953]_  = ~\new_[30647]_  | ~\new_[30572]_  | ~\new_[20779]_  | ~\new_[29050]_ ;
  assign \new_[18954]_  = ~\new_[30615]_  | ~\new_[30628]_  | ~\new_[20729]_  | ~\new_[30627]_ ;
  assign \new_[18955]_  = ~\new_[30752]_  | ~\new_[30717]_  | ~\new_[21889]_  | ~\new_[30519]_ ;
  assign \new_[18956]_  = ~\new_[30507]_  | ~\new_[30544]_  | ~\new_[20730]_  | ~\new_[30727]_ ;
  assign \new_[18957]_  = ~\new_[30630]_  | ~\new_[30786]_  | ~\new_[20971]_  | ~\new_[30290]_ ;
  assign \new_[18958]_  = ~\new_[30725]_  | ~\new_[28001]_  | ~\new_[21845]_  | ~\new_[30099]_ ;
  assign \new_[18959]_  = ~\new_[30775]_  | ~\new_[29299]_  | ~\new_[21349]_  | ~\new_[28215]_ ;
  assign \new_[18960]_  = ~\new_[22186]_  & (~\new_[22556]_  | ~\new_[23912]_ );
  assign \new_[18961]_  = ~\new_[30598]_  & (~\new_[22460]_  | ~\new_[24796]_ );
  assign \new_[18962]_  = ~\new_[19660]_ ;
  assign \new_[18963]_  = ~\new_[19661]_ ;
  assign \new_[18964]_  = ~\new_[23339]_  & (~\new_[22547]_  | ~\new_[25153]_ );
  assign \new_[18965]_  = ~\new_[28270]_  & (~\new_[22109]_  | ~\new_[23342]_ );
  assign \new_[18966]_  = ~\new_[30782]_  | ~\new_[24357]_  | ~\new_[23106]_  | ~\new_[26367]_ ;
  assign \new_[18967]_  = ~\new_[29992]_  & (~\new_[22394]_  | ~\new_[23349]_ );
  assign \new_[18968]_  = ~\new_[23350]_  & (~\new_[23417]_  | ~\new_[22463]_ );
  assign \new_[18969]_  = ~\new_[28678]_  & (~\new_[22169]_  | ~\new_[24524]_ );
  assign \new_[18970]_  = ~\new_[22444]_  & (~\new_[22548]_  | ~\new_[25270]_ );
  assign \new_[18971]_  = ~\new_[26880]_  & (~\new_[22551]_  | ~\new_[25170]_ );
  assign \new_[18972]_  = ~\new_[28992]_  & (~\new_[22519]_  | ~\new_[23773]_ );
  assign \new_[18973]_  = ~\new_[30287]_  & (~\new_[22465]_  | ~\new_[22121]_ );
  assign \new_[18974]_  = ~\new_[19667]_ ;
  assign \new_[18975]_  = ~\new_[30287]_  & (~\new_[22465]_  | ~\new_[28115]_ );
  assign \new_[18976]_  = ~\new_[23347]_  | ~\new_[24478]_  | ~\new_[27474]_  | ~\new_[30248]_ ;
  assign \new_[18977]_  = ~\new_[29826]_  & (~\new_[22356]_  | ~\new_[23377]_ );
  assign \new_[18978]_  = ~\new_[23378]_  & (~\new_[24097]_  | ~\new_[22513]_ );
  assign \new_[18979]_  = ~\new_[30733]_  & (~\new_[22206]_  | ~\new_[23642]_ );
  assign \new_[18980]_  = ~\new_[29541]_  & (~\new_[22472]_  | ~\new_[23679]_ );
  assign \new_[18981]_  = ~\new_[23452]_  & (~\new_[24491]_  | ~\new_[22474]_ );
  assign \new_[18982]_  = ~\new_[30109]_  & (~\new_[21593]_  | ~\new_[24842]_ );
  assign \new_[18983]_  = ~\new_[19672]_ ;
  assign \new_[18984]_  = ~\new_[29096]_  & (~\new_[22497]_  | ~\new_[23390]_ );
  assign \new_[18985]_  = ~\new_[30109]_  & (~\new_[21593]_  | ~\new_[28492]_ );
  assign \new_[18986]_  = ~\new_[21562]_  & (~\new_[23048]_  | ~\new_[23894]_ );
  assign \new_[18987]_  = ~\new_[29848]_  & (~\new_[22252]_  | ~\new_[23570]_ );
  assign \new_[18988]_  = ~\new_[23418]_  & (~\new_[23090]_  | ~\new_[22473]_ );
  assign \new_[18989]_  = ~\new_[27787]_  | ~\new_[21007]_  | ~\new_[30665]_ ;
  assign \new_[18990]_  = ~\new_[29217]_  & (~\new_[22480]_  | ~\new_[23480]_ );
  assign \new_[18991]_  = ~\new_[23495]_  | ~\new_[23186]_  | ~\new_[26745]_  | ~\new_[29808]_ ;
  assign \new_[18992]_  = ~\new_[29058]_  & (~\new_[22478]_  | ~\new_[23524]_ );
  assign \new_[18993]_  = ~\new_[30121]_  & (~\new_[22382]_  | ~\new_[23668]_ );
  assign \new_[18994]_  = ~\new_[19684]_ ;
  assign \new_[18995]_  = ~\new_[23461]_  | ~\new_[24402]_  | ~\new_[27769]_  | ~\new_[30693]_ ;
  assign \new_[18996]_  = ~\new_[29166]_  & (~\new_[22483]_  | ~\new_[28475]_ );
  assign \new_[18997]_  = ~\new_[29593]_  | ~\new_[21011]_  | ~\new_[30217]_ ;
  assign \new_[18998]_  = ~\new_[22194]_  & (~\new_[22552]_  | ~\new_[24691]_ );
  assign \new_[18999]_  = ~\new_[28021]_  & (~\new_[23473]_  | ~\new_[22197]_ );
  assign \new_[19000]_  = ~\new_[23382]_  & (~\new_[22550]_  | ~\new_[23167]_ );
  assign \new_[19001]_  = ~\new_[19690]_ ;
  assign \new_[19002]_  = ~\new_[29290]_  & (~\new_[22193]_  | ~\new_[23674]_ );
  assign \new_[19003]_  = ~\new_[19691]_ ;
  assign \new_[19004]_  = ~\new_[21181]_  & (~\new_[23187]_  | ~\new_[23895]_ );
  assign \new_[19005]_  = ~\new_[21181]_  & (~\new_[22558]_  | ~\new_[23895]_ );
  assign \new_[19006]_  = ~\new_[22246]_  & (~\new_[23121]_  | ~\new_[22482]_ );
  assign \new_[19007]_  = ~\new_[30555]_  | ~\new_[23184]_  | ~\new_[23442]_  | ~\new_[24487]_ ;
  assign \new_[19008]_  = ~\new_[28982]_  & (~\new_[21576]_  | ~\new_[23522]_ );
  assign \new_[19009]_  = ~\new_[29700]_  & (~\new_[22544]_  | ~\new_[23725]_ );
  assign \new_[19010]_  = ~\new_[28982]_  & (~\new_[21576]_  | ~\new_[28048]_ );
  assign \new_[19011]_  = ~\new_[30647]_  | ~\new_[24423]_  | ~\new_[23489]_  | ~\new_[26396]_ ;
  assign \new_[19012]_  = ~\new_[30206]_  & (~\new_[22201]_  | ~\new_[22247]_ );
  assign \new_[19013]_  = ~\new_[30515]_  & (~\new_[22523]_  | ~\new_[24933]_ );
  assign \new_[19014]_  = ~\new_[19699]_ ;
  assign \new_[19015]_  = ~\new_[30078]_  & (~\new_[22370]_  | ~\new_[22345]_ );
  assign \new_[19016]_  = ~\new_[23559]_  & (~\new_[22559]_  | ~\new_[23906]_ );
  assign \new_[19017]_  = ~\new_[29331]_  & (~\new_[22510]_  | ~\new_[23562]_ );
  assign \new_[19018]_  = ~\new_[29157]_  & (~\new_[22493]_  | ~\new_[23560]_ );
  assign \new_[19019]_  = ~\new_[19706]_ ;
  assign \new_[19020]_  = ~\new_[25062]_  & (~\new_[22557]_  | ~\new_[25194]_ );
  assign \new_[19021]_  = ~\new_[30236]_  & (~\new_[22265]_  | ~\new_[24521]_ );
  assign \new_[19022]_  = ~\new_[22260]_  & (~\new_[22555]_  | ~\new_[25185]_ );
  assign \new_[19023]_  = ~\new_[30251]_  & (~\new_[22153]_  | ~\new_[23478]_ );
  assign \new_[19024]_  = ~\new_[23582]_  & (~\new_[23621]_  | ~\new_[22495]_ );
  assign \new_[19025]_  = ~\new_[30544]_  | ~\new_[22013]_  | ~\new_[29927]_ ;
  assign \new_[19026]_  = ~\new_[28039]_  | ~\new_[21017]_  | ~\new_[30636]_ ;
  assign \new_[19027]_  = ~\new_[21014]_  | ~\new_[30467]_ ;
  assign \new_[19028]_  = ~\new_[29096]_  & (~\new_[22497]_  | ~\new_[28501]_ );
  assign \new_[19029]_  = ~\new_[24827]_  & (~\new_[22561]_  | ~\new_[23889]_ );
  assign \new_[19030]_  = ~\new_[29254]_  & (~\new_[22511]_  | ~\new_[23337]_ );
  assign \new_[19031]_  = ~\new_[30423]_  & (~\new_[22533]_  | ~\new_[24968]_ );
  assign \new_[19032]_  = ~\new_[19710]_ ;
  assign \new_[19033]_  = ~\new_[30423]_  & (~\new_[22533]_  | ~\new_[28556]_ );
  assign \new_[19034]_  = ~\new_[30270]_  & (~\new_[22223]_  | ~\new_[23589]_ );
  assign \new_[19035]_  = ~\new_[29115]_  & (~\new_[22469]_  | ~\new_[23444]_ );
  assign \new_[19036]_  = ~\new_[30063]_  & (~\new_[22502]_  | ~\new_[24990]_ );
  assign \new_[19037]_  = ~\new_[19716]_ ;
  assign \new_[19038]_  = ~\new_[30063]_  & (~\new_[22502]_  | ~\new_[28122]_ );
  assign \new_[19039]_  = ~\new_[29773]_  & (~\new_[23685]_  | ~\new_[22310]_ );
  assign \new_[19040]_  = ~\new_[28357]_  & (~\new_[22294]_  | ~\new_[23626]_ );
  assign \new_[19041]_  = ~\new_[29300]_  & (~\new_[22234]_  | ~\new_[22302]_ );
  assign \new_[19042]_  = ~\new_[21202]_  & (~\new_[26275]_  | ~\new_[23917]_ );
  assign \new_[19043]_  = ~\new_[30491]_  | ~\new_[21012]_  | ~\new_[30600]_ ;
  assign \new_[19044]_  = ~\new_[29229]_  & (~\new_[22503]_  | ~\new_[23962]_ );
  assign \new_[19045]_  = ~\new_[29916]_  & (~\new_[23927]_  | ~\new_[22267]_ );
  assign \new_[19046]_  = ~\new_[30741]_  & (~\new_[26984]_  | ~\new_[22312]_ );
  assign \new_[19047]_  = ~\new_[28204]_  & (~\new_[22504]_  | ~\new_[25003]_ );
  assign \new_[19048]_  = ~\new_[28204]_  & (~\new_[22504]_  | ~\new_[28573]_ );
  assign \new_[19049]_  = ~\new_[23683]_  & (~\new_[24065]_  | ~\new_[22506]_ );
  assign \new_[19050]_  = ~\new_[29331]_  & (~\new_[22510]_  | ~\new_[28559]_ );
  assign \new_[19051]_  = ~\new_[29113]_  & (~\new_[22164]_  | ~\new_[25034]_ );
  assign \new_[19052]_  = ~\new_[30420]_  & (~\new_[22332]_  | ~\new_[24549]_ );
  assign \new_[19053]_  = ~\new_[29671]_  & (~\new_[22538]_  | ~\new_[23838]_ );
  assign \new_[19054]_  = ~\new_[30308]_  & (~\new_[22334]_  | ~\new_[23611]_ );
  assign \new_[19055]_  = ~\new_[19724]_ ;
  assign \new_[19056]_  = ~\new_[29169]_  & (~\new_[22329]_  | ~\new_[24483]_ );
  assign \new_[19057]_  = ~\new_[29955]_  & (~\new_[22339]_  | ~\new_[23826]_ );
  assign \new_[19058]_  = ~\new_[30752]_  | ~\new_[24432]_  | ~\new_[25043]_  | ~\new_[26212]_ ;
  assign \new_[19059]_  = ~\new_[25123]_  & (~\new_[25505]_  | ~\new_[22507]_ );
  assign \new_[19060]_  = ~\new_[30630]_  | ~\new_[24499]_  | ~\new_[23659]_  | ~\new_[25357]_ ;
  assign \new_[19061]_  = ~\new_[29167]_  & (~\new_[22539]_  | ~\new_[23851]_ );
  assign \new_[19062]_  = ~\new_[29101]_  & (~\new_[22512]_  | ~\new_[23371]_ );
  assign \new_[19063]_  = ~\new_[30445]_  & (~\new_[21580]_  | ~\new_[28154]_ );
  assign \new_[19064]_  = ~\new_[21248]_  & (~\new_[21585]_  | ~\new_[25188]_ );
  assign \new_[19065]_  = ~\new_[29277]_  & (~\new_[22317]_  | ~\new_[23666]_ );
  assign \new_[19066]_  = ~\new_[21206]_  & (~\new_[21798]_  | ~\new_[23952]_ );
  assign \new_[19067]_  = ~\new_[28999]_  & (~\new_[22291]_  | ~\new_[23682]_ );
  assign \new_[19068]_  = ~\new_[29970]_  & (~\new_[24884]_  | ~\new_[22155]_ );
  assign \new_[19069]_  = ~\new_[30445]_  & (~\new_[21580]_  | ~\new_[23718]_ );
  assign \new_[19070]_  = ~\new_[29985]_  & (~\new_[22399]_  | ~\new_[22365]_ );
  assign \new_[19071]_  = ~\new_[23549]_  & (~\new_[24378]_  | ~\new_[22516]_ );
  assign \new_[19072]_  = ~\new_[23739]_  & (~\new_[22549]_  | ~\new_[23930]_ );
  assign \new_[19073]_  = ~\new_[28998]_  & (~\new_[22248]_  | ~\new_[23770]_ );
  assign \new_[19074]_  = ~\new_[23744]_  & (~\new_[23118]_  | ~\new_[22521]_ );
  assign \new_[19075]_  = ~\new_[22245]_  & (~\new_[22553]_  | ~\new_[25207]_ );
  assign \new_[19076]_  = ~\new_[19740]_ ;
  assign \new_[19077]_  = ~\new_[30117]_  | ~\new_[21023]_  | ~\new_[29563]_ ;
  assign n7679 = ~\new_[29376]_  | ~\new_[21044]_ ;
  assign \new_[19079]_  = ~\new_[23880]_  | ~\new_[25209]_  | ~\new_[27546]_  | ~\new_[30233]_ ;
  assign \new_[19080]_  = ~\new_[30515]_  & (~\new_[22523]_  | ~\new_[28164]_ );
  assign \new_[19081]_  = ~\new_[23406]_  & (~\new_[24445]_  | ~\new_[22468]_ );
  assign n7694 = ~\new_[29163]_  | ~\new_[21031]_ ;
  assign n7699 = ~\new_[29409]_  | ~\new_[21035]_ ;
  assign n7669 = ~\new_[29280]_  | ~\new_[21038]_ ;
  assign n7674 = ~\new_[29323]_  | ~\new_[21030]_ ;
  assign n7689 = ~\new_[29037]_  | ~\new_[21046]_ ;
  assign n7684 = ~\new_[28921]_  | ~\new_[21048]_ ;
  assign \new_[19088]_  = ~\new_[30309]_  & (~\new_[22534]_  | ~\new_[28297]_ );
  assign \new_[19089]_  = ~\new_[29537]_  | ~\new_[21021]_  | ~\new_[29210]_ ;
  assign \new_[19090]_  = ~\new_[30309]_  & (~\new_[22534]_  | ~\new_[25041]_ );
  assign \new_[19091]_  = ~\new_[29047]_  & (~\new_[22535]_  | ~\new_[23514]_ );
  assign \new_[19092]_  = ~\new_[23391]_  & (~\new_[22562]_  | ~\new_[23950]_ );
  assign \new_[19093]_  = ~\new_[30466]_  & (~\new_[22425]_  | ~\new_[25126]_ );
  assign \new_[19094]_  = ~\new_[30598]_  & (~\new_[22460]_  | ~\new_[28585]_ );
  assign \new_[19095]_  = ~\new_[19748]_ ;
  assign \new_[19096]_  = ~\new_[19749]_ ;
  assign \new_[19097]_  = ~\new_[29166]_  & (~\new_[22483]_  | ~\new_[23351]_ );
  assign \new_[19098]_  = ~\new_[29354]_  & (~\new_[22541]_  | ~\new_[23483]_ );
  assign \new_[19099]_  = ~\new_[26655]_  | ~\new_[21008]_  | ~\new_[30255]_ ;
  assign \new_[19100]_  = ~\new_[19750]_ ;
  assign \new_[19101]_  = ~\new_[23746]_  & (~\new_[23152]_  | ~\new_[22514]_ );
  assign \new_[19102]_  = ~\new_[19753]_ ;
  assign \new_[19103]_  = ~\new_[30072]_  & (~\new_[23789]_  | ~\new_[22396]_ );
  assign \new_[19104]_  = ~\new_[23869]_  & (~\new_[23569]_  | ~\new_[22522]_ );
  assign \new_[19105]_  = ~\new_[25084]_  & (~\new_[22560]_  | ~\new_[24578]_ );
  assign \new_[19106]_  = ~\new_[30584]_  & (~\new_[22451]_  | ~\new_[25143]_ );
  assign \new_[19107]_  = ~\new_[19760]_ ;
  assign \new_[19108]_  = ~\new_[29172]_  & (~\new_[22545]_  | ~\new_[23882]_ );
  assign \new_[19109]_  = ~\new_[26188]_  & (~\new_[22405]_  | ~\new_[30297]_ );
  assign \new_[19110]_  = ~\new_[24788]_  & (~\new_[22315]_  | ~\new_[29868]_ );
  assign \new_[19111]_  = ~\new_[24525]_  & (~\new_[22290]_  | ~\new_[29893]_ );
  assign \new_[19112]_  = \new_[20810]_  & \new_[26309]_ ;
  assign \new_[19113]_  = ~\new_[24157]_  & (~\new_[22266]_  | ~\new_[28993]_ );
  assign \new_[19114]_  = ~\new_[24311]_  & (~\new_[22352]_  | ~\new_[29681]_ );
  assign \new_[19115]_  = \new_[20890]_  & \new_[26239]_ ;
  assign \new_[19116]_  = ~\new_[26378]_  & (~\new_[22231]_  | ~\new_[30293]_ );
  assign \new_[19117]_  = \new_[20923]_  & \new_[24782]_ ;
  assign \new_[19118]_  = ~\new_[22909]_  & (~\new_[22432]_  | ~\new_[30149]_ );
  assign \new_[19119]_  = \new_[20795]_  & \new_[26267]_ ;
  assign \new_[19120]_  = ~\new_[24428]_  & (~\new_[22380]_  | ~\new_[28675]_ );
  assign \new_[19121]_  = ~\new_[26707]_  & (~\new_[22429]_  | ~\new_[29851]_ );
  assign \new_[19122]_  = \new_[20949]_  & \new_[27594]_ ;
  assign \new_[19123]_  = ~\new_[20732]_  & ~\new_[29861]_ ;
  assign \new_[19124]_  = ~\new_[20984]_  | ~\new_[30283]_ ;
  assign \new_[19125]_  = ~\new_[20832]_  & ~\new_[29238]_ ;
  assign \new_[19126]_  = ~\new_[29874]_  | (~\new_[22108]_  & ~\new_[25104]_ );
  assign \new_[19127]_  = ~\new_[20885]_  | ~\new_[30280]_ ;
  assign \new_[19128]_  = ~\new_[20834]_  & ~\new_[29841]_ ;
  assign \new_[19129]_  = ~\new_[30337]_  | (~\new_[22375]_  & ~\new_[23759]_ );
  assign \new_[19130]_  = ~\new_[20756]_  & ~\new_[30140]_ ;
  assign \new_[19131]_  = ~\new_[20823]_  & ~\new_[30044]_ ;
  assign \new_[19132]_  = ~\new_[20760]_  & ~\new_[30253]_ ;
  assign \new_[19133]_  = ~\new_[20882]_  & ~\new_[30633]_ ;
  assign \new_[19134]_  = ~\new_[30289]_  & (~\new_[22238]_  | ~\new_[26896]_ );
  assign \new_[19135]_  = ~\new_[20788]_  & ~\new_[30202]_ ;
  assign \new_[19136]_  = ~\new_[29692]_  | (~\new_[22119]_  & ~\new_[23446]_ );
  assign \new_[19137]_  = ~\new_[30757]_  & (~\new_[22178]_  | ~\new_[23521]_ );
  assign \new_[19138]_  = ~\new_[20767]_  | ~\new_[29103]_ ;
  assign \new_[19139]_  = ~\new_[20977]_  & ~\new_[28899]_ ;
  assign \new_[19140]_  = ~\new_[20803]_  & ~\new_[29573]_ ;
  assign \new_[19141]_  = ~\new_[20800]_  | ~\new_[30037]_ ;
  assign \new_[19142]_  = ~\new_[20787]_  & ~\new_[29565]_ ;
  assign \new_[19143]_  = ~\new_[30280]_  | (~\new_[22233]_  & ~\new_[24914]_ );
  assign \new_[19144]_  = ~\new_[29544]_  & (~\new_[25073]_  | ~\new_[22203]_ );
  assign \new_[19145]_  = ~\new_[20914]_  | ~\new_[30409]_ ;
  assign \new_[19146]_  = \new_[20818]_  | \new_[29181]_ ;
  assign \new_[19147]_  = ~\new_[30217]_  | (~\new_[22225]_  & ~\new_[22224]_ );
  assign \new_[19148]_  = ~\new_[20838]_  | ~\new_[30005]_ ;
  assign \new_[19149]_  = ~\new_[30005]_  | (~\new_[22162]_  & ~\new_[25141]_ );
  assign \new_[19150]_  = ~\new_[29441]_  | (~\new_[22457]_  & ~\new_[23872]_ );
  assign \new_[19151]_  = ~\new_[29222]_  & (~\new_[22279]_  | ~\new_[23468]_ );
  assign \new_[19152]_  = ~\new_[20972]_  & ~\new_[29445]_ ;
  assign \new_[19153]_  = ~\new_[20947]_  & ~\new_[29629]_ ;
  assign \new_[19154]_  = ~\new_[20852]_  | ~\new_[30086]_ ;
  assign \new_[19155]_  = ~\new_[30086]_  | (~\new_[22323]_  & ~\new_[24950]_ );
  assign \new_[19156]_  = \new_[20821]_  | \new_[29181]_ ;
  assign \new_[19157]_  = ~\new_[20884]_  | ~\new_[30645]_ ;
  assign \new_[19158]_  = ~\new_[29139]_  | (~\new_[22257]_  & ~\new_[23523]_ );
  assign \new_[19159]_  = ~\new_[30342]_  & (~\new_[23423]_  | ~\new_[22293]_ );
  assign \new_[19160]_  = ~\new_[20862]_  | ~\new_[28963]_ ;
  assign \new_[19161]_  = ~\new_[30409]_  | (~\new_[23584]_  & ~\new_[22132]_ );
  assign \new_[19162]_  = ~\new_[20749]_  & ~\new_[29767]_ ;
  assign \new_[19163]_  = ~\new_[20892]_  & ~\new_[29174]_ ;
  assign \new_[19164]_  = ~\new_[30125]_  | (~\new_[22249]_  & ~\new_[25010]_ );
  assign \new_[19165]_  = ~\new_[20766]_  & ~\new_[30415]_ ;
  assign \new_[19166]_  = ~\new_[30438]_  & (~\new_[22313]_  | ~\new_[27547]_ );
  assign \new_[19167]_  = ~\new_[28828]_  | (~\new_[22331]_  & ~\new_[23687]_ );
  assign \new_[19168]_  = ~\new_[30316]_  | (~\new_[22325]_  & ~\new_[23379]_ );
  assign \new_[19169]_  = ~\new_[30162]_  & (~\new_[23839]_  | ~\new_[22369]_ );
  assign \new_[19170]_  = ~\new_[30610]_  | (~\new_[22328]_  & ~\new_[22209]_ );
  assign \new_[19171]_  = ~\new_[20864]_  & ~\new_[29944]_ ;
  assign \new_[19172]_  = ~\new_[20917]_  & ~\new_[30058]_ ;
  assign \new_[19173]_  = ~\new_[20903]_  & ~\new_[30212]_ ;
  assign \new_[19174]_  = ~\new_[20775]_  & ~\new_[30114]_ ;
  assign \new_[19175]_  = ~\new_[30147]_  | (~\new_[23824]_  & ~\new_[22414]_ );
  assign \new_[19176]_  = ~\new_[28898]_  | (~\new_[22304]_  & ~\new_[23834]_ );
  assign \new_[19177]_  = ~\new_[30142]_  | (~\new_[22308]_  & ~\new_[25061]_ );
  assign \new_[19178]_  = ~\new_[29560]_  | (~\new_[22406]_  & ~\new_[23470]_ );
  assign \new_[19179]_  = ~\new_[30036]_  & (~\new_[22395]_  | ~\new_[23712]_ );
  assign \new_[19180]_  = ~\new_[20870]_  & ~\new_[30350]_ ;
  assign \new_[19181]_  = ~\new_[20841]_  | ~\new_[29870]_ ;
  assign \new_[19182]_  = ~\new_[20867]_  | ~\new_[29867]_ ;
  assign \new_[19183]_  = ~\new_[30055]_  & (~\new_[23735]_  | ~\new_[22353]_ );
  assign \new_[19184]_  = ~\new_[20981]_  | ~\new_[30142]_ ;
  assign \new_[19185]_  = ~\new_[30105]_  | (~\new_[23503]_  & ~\new_[22408]_ );
  assign \new_[19186]_  = ~\new_[20988]_  | ~\new_[30123]_ ;
  assign \new_[19187]_  = ~\new_[30123]_  | (~\new_[22180]_  & ~\new_[24895]_ );
  assign \new_[19188]_  = ~\new_[29226]_  | (~\new_[22434]_  & ~\new_[23475]_ );
  assign \new_[19189]_  = ~\new_[20992]_  & ~\new_[29564]_ ;
  assign \new_[19190]_  = ~\new_[20993]_  | ~\new_[30262]_ ;
  assign \new_[19191]_  = ~\new_[20776]_  | ~\new_[30104]_ ;
  assign \new_[19192]_  = ~\new_[30150]_  | (~\new_[22191]_  & ~\new_[23883]_ );
  assign \new_[19193]_  = ~\new_[24282]_  & (~\new_[22546]_  | ~\new_[28049]_ );
  assign \new_[19194]_  = ~\new_[21470]_  & (~\new_[22466]_  | ~\new_[25811]_ );
  assign \new_[19195]_  = ~\new_[22988]_  & (~\new_[22467]_  | ~\new_[25413]_ );
  assign \new_[19196]_  = ~\new_[24415]_  & (~\new_[22501]_  | ~\new_[26170]_ );
  assign \new_[19197]_  = ~\new_[22869]_  & (~\new_[22515]_  | ~\new_[26237]_ );
  assign \new_[19198]_  = ~\new_[23018]_  & (~\new_[22527]_  | ~\new_[26768]_ );
  assign \new_[19199]_  = ~\new_[21512]_  & (~\new_[22509]_  | ~\new_[25483]_ );
  assign \new_[19200]_  = ~\new_[23009]_  & (~\new_[22490]_  | ~\new_[26168]_ );
  assign \new_[19201]_  = ~\new_[23085]_  & (~\new_[22498]_  | ~\new_[26159]_ );
  assign \new_[19202]_  = ~\new_[21775]_  & (~\new_[22508]_  | ~\new_[28490]_ );
  assign \new_[19203]_  = ~\new_[22917]_  & (~\new_[22491]_  | ~\new_[28538]_ );
  assign \new_[19204]_  = ~\new_[24342]_  & (~\new_[22540]_  | ~\new_[26812]_ );
  assign \new_[19205]_  = ~\new_[22855]_  & (~\new_[22542]_  | ~\new_[26790]_ );
  assign \new_[19206]_  = ~\new_[23334]_  & (~\new_[22450]_  | ~\new_[27636]_ );
  assign \new_[19207]_  = ~\new_[30342]_  & (~\new_[22293]_  | ~\new_[28634]_ );
  assign \new_[19208]_  = ~\new_[29544]_  & (~\new_[22203]_  | ~\new_[29311]_ );
  assign \new_[19209]_  = ~\new_[22214]_  & (~\new_[22213]_  | ~\new_[27745]_ );
  assign \new_[19210]_  = ~\new_[21010]_  | ~\new_[30217]_ ;
  assign \new_[19211]_  = ~\new_[21020]_  | ~\new_[29233]_ ;
  assign \new_[19212]_  = ~\new_[21242]_  & (~\new_[22237]_  | ~\new_[27762]_ );
  assign \new_[19213]_  = ~\new_[21240]_  & (~\new_[22305]_  | ~\new_[27746]_ );
  assign \new_[19214]_  = ~\new_[30162]_  & (~\new_[22369]_  | ~\new_[29413]_ );
  assign \new_[19215]_  = ~\new_[21247]_  & (~\new_[22335]_  | ~\new_[28507]_ );
  assign \new_[19216]_  = ~\new_[21234]_  & (~\new_[22130]_  | ~\new_[27619]_ );
  assign \new_[19217]_  = ~\new_[30147]_  | (~\new_[22414]_  & ~\new_[27689]_ );
  assign \new_[19218]_  = ~\new_[30055]_  & (~\new_[22353]_  | ~\new_[27694]_ );
  assign \new_[19219]_  = ~\new_[30610]_  | (~\new_[22209]_  & ~\new_[27559]_ );
  assign \new_[19220]_  = ~\new_[21159]_  & (~\new_[22437]_  | ~\new_[27589]_ );
  assign \new_[19221]_  = ~\new_[20733]_  & (~\new_[29357]_  | ~\new_[29676]_ );
  assign \new_[19222]_  = ~\new_[26573]_  & (~\new_[22520]_  | ~\new_[26218]_ );
  assign \new_[19223]_  = ~\new_[27254]_  & (~\new_[22462]_  | ~\new_[27611]_ );
  assign \new_[19224]_  = ~\new_[24320]_  & (~\new_[22492]_  | ~\new_[25046]_ );
  assign \new_[19225]_  = ~\new_[25598]_  & (~\new_[22487]_  | ~\new_[24513]_ );
  assign \new_[19226]_  = ~\new_[26369]_  & (~\new_[22477]_  | ~\new_[24389]_ );
  assign \new_[19227]_  = ~\new_[24302]_  & (~\new_[22481]_  | ~\new_[24391]_ );
  assign \new_[19228]_  = ~\new_[20935]_  & (~\new_[28962]_  | ~\new_[29089]_ );
  assign \new_[19229]_  = ~\new_[26288]_  & (~\new_[22500]_  | ~\new_[23142]_ );
  assign \new_[19230]_  = ~\new_[24259]_  & (~\new_[22470]_  | ~\new_[26238]_ );
  assign \new_[19231]_  = ~\new_[26370]_  & (~\new_[22464]_  | ~\new_[26667]_ );
  assign \new_[19232]_  = ~\new_[22221]_  & (~\new_[22485]_  | ~\new_[24383]_ );
  assign \new_[19233]_  = ~\new_[20854]_  & (~\new_[29202]_  | ~\new_[29639]_ );
  assign \new_[19234]_  = ~\new_[24263]_  & (~\new_[22471]_  | ~\new_[24039]_ );
  assign \new_[19235]_  = ~\new_[22878]_  & (~\new_[22532]_  | ~\new_[24591]_ );
  assign \new_[19236]_  = ~\new_[20943]_  & (~\new_[29744]_  | ~\new_[29582]_ );
  assign \new_[19237]_  = ~\new_[20920]_  & (~\new_[29104]_  | ~\new_[29576]_ );
  assign \new_[19238]_  = ~\new_[24308]_  & (~\new_[21590]_  | ~\new_[26255]_ );
  assign \new_[19239]_  = ~\new_[26265]_  & (~\new_[22543]_  | ~\new_[27531]_ );
  assign \new_[19240]_  = ~\new_[20978]_  & (~\new_[30363]_  | ~\new_[29606]_ );
  assign \new_[19241]_  = ~\new_[23006]_  & (~\new_[22537]_  | ~\new_[24407]_ );
  assign \new_[19242]_  = ~\new_[20785]_  & (~\new_[29350]_  | ~\new_[29333]_ );
  assign \new_[19243]_  = ~\new_[22874]_  & (~\new_[22489]_  | ~\new_[27854]_ );
  assign \new_[19244]_  = ~\new_[21311]_  & ~\new_[30055]_ ;
  assign \new_[19245]_  = ~\new_[21300]_  & ~\new_[30240]_ ;
  assign \new_[19246]_  = ~\new_[21297]_  & ~\new_[28857]_ ;
  assign \new_[19247]_  = ~\new_[23608]_  & ~\new_[29663]_ ;
  assign \new_[19248]_  = \new_[21130]_  | \new_[30660]_ ;
  assign n8609 = m4_s4_cyc_o_reg;
  assign \new_[19250]_  = ~\new_[22207]_  & ~\new_[29227]_ ;
  assign \new_[19251]_  = \new_[21301]_  | \new_[27529]_ ;
  assign \new_[19252]_  = ~\new_[22232]_  & ~\new_[29578]_ ;
  assign \new_[19253]_  = ~\new_[21159]_  & ~\new_[29774]_ ;
  assign \new_[19254]_  = ~\new_[23434]_  & ~\new_[28833]_ ;
  assign \new_[19255]_  = \new_[21270]_  | \new_[28470]_ ;
  assign \new_[19256]_  = \new_[21294]_  | \new_[27500]_ ;
  assign \new_[19257]_  = ~\new_[21170]_  | ~\new_[28883]_ ;
  assign \new_[19258]_  = \new_[21324]_  | \new_[27511]_ ;
  assign \new_[19259]_  = ~\new_[22189]_  & ~\new_[29465]_ ;
  assign \new_[19260]_  = ~\new_[20038]_ ;
  assign \new_[19261]_  = \new_[21276]_  | \new_[27509]_ ;
  assign \new_[19262]_  = \new_[21267]_  | \new_[28352]_ ;
  assign \new_[19263]_  = ~\new_[22405]_  | ~\new_[21343]_ ;
  assign \new_[19264]_  = ~\new_[23747]_  & ~\new_[29056]_ ;
  assign \new_[19265]_  = \new_[21314]_  | \new_[27441]_ ;
  assign \new_[19266]_  = ~\new_[21240]_  & ~\new_[30176]_ ;
  assign \new_[19267]_  = ~\new_[23398]_  & ~\new_[29394]_ ;
  assign \new_[19268]_  = \new_[21315]_  | \new_[27517]_ ;
  assign \new_[19269]_  = ~\new_[21291]_  & ~\new_[30637]_ ;
  assign \new_[19270]_  = ~\new_[21193]_  | ~\new_[27130]_ ;
  assign \new_[19271]_  = ~\new_[21239]_  | ~\new_[28429]_ ;
  assign \new_[19272]_  = ~\new_[21182]_  | ~\new_[27642]_ ;
  assign \new_[19273]_  = ~\new_[21219]_  & ~\new_[24346]_ ;
  assign \new_[19274]_  = ~\new_[21197]_  | ~\new_[28939]_ ;
  assign \new_[19275]_  = \new_[21130]_  | \new_[22124]_ ;
  assign \new_[19276]_  = ~\new_[23366]_  & ~\new_[29195]_ ;
  assign \new_[19277]_  = ~\new_[21201]_  | ~\new_[26581]_ ;
  assign \new_[19278]_  = \new_[20561]_  | \new_[27311]_ ;
  assign \new_[19279]_  = ~\new_[21242]_  & ~\new_[28979]_ ;
  assign \new_[19280]_  = ~\new_[21247]_  & ~\new_[30032]_ ;
  assign \new_[19281]_  = ~\new_[21234]_  & ~\new_[29745]_ ;
  assign n8399 = m4_s5_cyc_o_reg;
  assign \new_[19283]_  = ~\new_[22320]_  & ~\new_[29068]_ ;
  assign \new_[19284]_  = ~\new_[21256]_  | ~\new_[28483]_ ;
  assign n8424 = m7_s7_cyc_o_reg;
  assign \new_[19286]_  = ~\new_[30258]_  | ~\new_[27500]_  | ~\new_[23014]_ ;
  assign \new_[19287]_  = \new_[21131]_  | \new_[26351]_ ;
  assign \new_[19288]_  = ~\new_[29907]_  & (~\new_[22963]_  | ~\new_[29483]_ );
  assign \new_[19289]_  = ~\new_[30375]_  & (~\new_[22852]_  | ~\new_[29480]_ );
  assign \new_[19290]_  = \new_[21171]_  | \new_[26187]_ ;
  assign \new_[19291]_  = ~\new_[30094]_  | ~\new_[27511]_  | ~\new_[23068]_ ;
  assign \new_[19292]_  = ~\new_[30038]_  & (~\new_[22114]_  | ~\new_[29351]_ );
  assign \new_[19293]_  = ~\new_[22867]_  | ~\new_[26252]_  | ~\new_[26189]_ ;
  assign \new_[19294]_  = ~\new_[30033]_  & (~\new_[22928]_  | ~\new_[29489]_ );
  assign \new_[19295]_  = ~\new_[20170]_ ;
  assign \new_[19296]_  = ~\new_[29792]_  & (~\new_[23038]_  | ~\new_[29474]_ );
  assign \new_[19297]_  = \new_[21224]_  | \new_[26568]_ ;
  assign \new_[19298]_  = ~\new_[29997]_  & (~\new_[22935]_  | ~\new_[29536]_ );
  assign \new_[19299]_  = ~\new_[29810]_  & (~\new_[22106]_  | ~\new_[29294]_ );
  assign \new_[19300]_  = ~\new_[23024]_  | ~\new_[26535]_  | ~\new_[24636]_ ;
  assign \new_[19301]_  = ~\new_[30381]_  | ~\new_[27509]_  | ~\new_[22915]_ ;
  assign \new_[19302]_  = ~\new_[23017]_  | ~\new_[26266]_  | ~\new_[26296]_ ;
  assign \new_[19303]_  = ~\new_[30275]_  & (~\new_[21571]_  | ~\new_[29601]_ );
  assign \new_[19304]_  = ~\new_[29465]_  | ~\new_[6051]_ ;
  assign \new_[19305]_  = ~\new_[21563]_  | ~\new_[26404]_  | ~\new_[26339]_ ;
  assign \new_[19306]_  = \new_[21215]_  | \new_[26195]_ ;
  assign \new_[19307]_  = ~\new_[30211]_  | ~\new_[27517]_  | ~\new_[22868]_ ;
  assign \new_[19308]_  = ~\new_[30151]_  & (~\new_[22883]_  | ~\new_[29390]_ );
  assign n8914 = m4_s7_cyc_o_reg;
  assign \new_[19310]_  = ~\new_[29840]_  | ~\new_[27341]_  | ~\new_[27727]_ ;
  assign \new_[19311]_  = \new_[21255]_  | \new_[26208]_ ;
  assign \new_[19312]_  = ~\new_[21228]_  | ~\new_[28894]_ ;
  assign \new_[19313]_  = ~\new_[21142]_  | ~\new_[30242]_ ;
  assign \new_[19314]_  = ~\new_[21160]_  | ~\new_[29421]_ ;
  assign \new_[19315]_  = ~\new_[23059]_  | (~\new_[22956]_  & ~\new_[30036]_ );
  assign \new_[19316]_  = ~\new_[23084]_  | (~\new_[24391]_  & ~\new_[28718]_ );
  assign \new_[19317]_  = ~\new_[21153]_  | ~\new_[30222]_ ;
  assign \new_[19318]_  = ~\new_[21218]_  | ~\new_[29868]_ ;
  assign \new_[19319]_  = ~\new_[22282]_  | ~\new_[28818]_ ;
  assign \new_[19320]_  = ~\new_[21150]_  | ~\new_[28918]_ ;
  assign \new_[19321]_  = ~\new_[21152]_  | ~\new_[29987]_ ;
  assign \new_[19322]_  = ~\new_[22297]_  | ~\new_[28595]_ ;
  assign \new_[19323]_  = ~\new_[21211]_  & ~\new_[24359]_ ;
  assign \new_[19324]_  = ~\new_[21225]_  | ~\new_[30525]_ ;
  assign \new_[19325]_  = ~\new_[21208]_  & ~\new_[24362]_ ;
  assign \new_[19326]_  = ~\new_[21246]_  & ~\new_[24343]_ ;
  assign \new_[19327]_  = ~\new_[21166]_  & ~\new_[23512]_ ;
  assign \new_[19328]_  = ~\new_[21237]_  | ~\new_[30233]_ ;
  assign \new_[19329]_  = ~\new_[29977]_  | ~\new_[5973]_  | ~\new_[29020]_  | ~\new_[23060]_ ;
  assign \new_[19330]_  = ~\new_[29260]_  | ~\new_[6044]_  | ~\new_[28918]_  | ~\new_[22999]_ ;
  assign \new_[19331]_  = ~\new_[29139]_  | ~\new_[6063]_  | ~\new_[29276]_  | ~\new_[22960]_ ;
  assign \new_[19332]_  = ~\new_[30246]_  | ~\new_[6058]_  | ~\new_[28818]_  | ~\new_[21823]_ ;
  assign \new_[19333]_  = ~\new_[30754]_  | ~\new_[6037]_  | ~\new_[30513]_  | ~\new_[22974]_ ;
  assign \new_[19334]_  = ~\new_[30147]_  | ~\new_[6185]_  | ~\new_[28675]_  | ~\new_[23016]_ ;
  assign \new_[19335]_  = ~\new_[30084]_  | ~\new_[6081]_  | ~\new_[29583]_  | ~\new_[22998]_ ;
  assign \new_[19336]_  = ~\new_[30508]_  | ~\new_[6041]_  | ~\new_[30229]_  | ~\new_[23004]_ ;
  assign \new_[19337]_  = ~\new_[30215]_  | ~\new_[6039]_  | ~\new_[28894]_  | ~\new_[22870]_ ;
  assign \new_[19338]_  = ~\new_[29874]_  | ~\new_[6035]_  | ~\new_[29028]_  | ~\new_[22877]_ ;
  assign \new_[19339]_  = ~\new_[30316]_  | ~\new_[6077]_  | ~\new_[29623]_  | ~\new_[22861]_ ;
  assign \new_[19340]_  = ~\new_[5903]_  | ~\new_[28656]_  | ~\new_[29767]_ ;
  assign \new_[19341]_  = ~\new_[6174]_  | ~\new_[29090]_  | ~\new_[30566]_ ;
  assign \new_[19342]_  = ~\new_[21461]_  | ~\new_[26392]_ ;
  assign n8379 = m2_s5_cyc_o_reg;
  assign n8354 = m3_s15_cyc_o_reg;
  assign \new_[19345]_  = ~\new_[6037]_  | ~\new_[26786]_  | ~\new_[30663]_ ;
  assign \new_[19346]_  = ~\new_[21513]_  | ~\new_[26515]_ ;
  assign \new_[19347]_  = ~\new_[6043]_  | ~\new_[27085]_  | ~\new_[30747]_ ;
  assign \new_[19348]_  = ~\new_[21482]_  | ~\new_[26342]_ ;
  assign \new_[19349]_  = ~\new_[21537]_  | ~\new_[26337]_ ;
  assign \new_[19350]_  = ~\new_[6063]_  | ~\new_[28156]_  | ~\new_[29222]_ ;
  assign \new_[19351]_  = ~\new_[31429]_  | ~\new_[26465]_  | ~\new_[29181]_ ;
  assign \new_[19352]_  = ~\new_[31394]_  | ~\new_[28158]_  | ~\new_[28909]_ ;
  assign \new_[19353]_  = ~\new_[31400]_  | ~\new_[29283]_  | ~\new_[30684]_ ;
  assign \new_[19354]_  = ~\new_[31491]_  | ~\new_[26789]_  | ~\new_[29828]_ ;
  assign \new_[19355]_  = ~\new_[31431]_  | ~\new_[26309]_  | ~\new_[29186]_ ;
  assign \new_[19356]_  = ~\new_[6197]_  | ~\new_[27814]_  | ~\new_[30688]_ ;
  assign \new_[19357]_  = ~\new_[6195]_  | ~\new_[28662]_  | ~\new_[29375]_ ;
  assign \new_[19358]_  = ~\new_[6186]_  | ~\new_[26711]_  | ~\new_[30840]_ ;
  assign n8704 = m3_s1_cyc_o_reg;
  assign \new_[19360]_  = ~\new_[6194]_  | ~\new_[26455]_  | ~\new_[30632]_ ;
  assign \new_[19361]_  = \new_[29590]_  & \new_[26269]_ ;
  assign \new_[19362]_  = ~\new_[5988]_  | ~\new_[30281]_  | ~\new_[28857]_ ;
  assign \new_[19363]_  = ~\new_[6076]_  | ~\new_[28117]_  | ~\new_[30637]_ ;
  assign \new_[19364]_  = ~\new_[6079]_  | ~\new_[27939]_  | ~\new_[30682]_ ;
  assign \new_[19365]_  = ~\new_[6003]_  | ~\new_[28986]_  | ~\new_[28236]_ ;
  assign \new_[19366]_  = ~\new_[31617]_  | ~\new_[27926]_  | ~\new_[29435]_ ;
  assign \new_[19367]_  = ~\new_[21550]_  | ~\new_[26430]_ ;
  assign \new_[19368]_  = ~\new_[21501]_  | ~\new_[24785]_ ;
  assign \new_[19369]_  = ~\new_[21487]_  | ~\new_[26358]_ ;
  assign \new_[19370]_  = ~\new_[21554]_  | ~\new_[26261]_ ;
  assign \new_[19371]_  = ~\new_[21189]_  | ~\new_[26262]_ ;
  assign \new_[19372]_  = ~\new_[20353]_ ;
  assign \new_[19373]_  = ~\new_[20355]_ ;
  assign \new_[19374]_  = ~\new_[6053]_  | ~\new_[28827]_  | ~\new_[29544]_ ;
  assign \new_[19375]_  = ~\new_[31890]_  | ~\new_[27848]_  | ~\new_[28935]_ ;
  assign \new_[19376]_  = ~\new_[6268]_  | ~\new_[29143]_  | ~\new_[30162]_ ;
  assign \new_[19377]_  = ~\new_[20357]_ ;
  assign \new_[19378]_  = ~\new_[20357]_ ;
  assign \new_[19379]_  = ~\new_[6095]_  | ~\new_[29155]_  | ~\new_[30276]_ ;
  assign \new_[19380]_  = ~\new_[5964]_  | ~\new_[28247]_  | ~\new_[29992]_ ;
  assign \new_[19381]_  = \new_[20522]_  | \new_[29218]_ ;
  assign \new_[19382]_  = ~\new_[28899]_  | ~\new_[6051]_ ;
  assign \new_[19383]_  = ~\new_[6064]_  | ~\new_[30369]_  | ~\new_[30002]_ ;
  assign \new_[19384]_  = \new_[21462]_  | \new_[29932]_ ;
  assign \new_[19385]_  = ~\new_[5914]_  | ~\new_[30091]_  | ~\new_[29931]_ ;
  assign \new_[19386]_  = ~\new_[6051]_  | ~\new_[30091]_  | ~\new_[29931]_ ;
  assign \new_[19387]_  = ~\new_[6206]_  | ~\new_[28741]_  | ~\new_[29926]_ ;
  assign \new_[19388]_  = ~\new_[6075]_  | ~\new_[28646]_  | ~\new_[30114]_ ;
  assign \new_[19389]_  = ~\new_[5979]_  | ~\new_[28246]_  | ~\new_[30328]_ ;
  assign \new_[19390]_  = ~\new_[6071]_  | ~\new_[30300]_  | ~\new_[29790]_ ;
  assign \new_[19391]_  = ~\new_[5917]_  | ~\new_[29801]_  | ~\new_[30053]_ ;
  assign \new_[19392]_  = ~\new_[5918]_  | ~\new_[28163]_  | ~\new_[30212]_ ;
  assign \new_[19393]_  = ~\new_[5923]_  | ~\new_[28646]_  | ~\new_[30114]_ ;
  assign \new_[19394]_  = ~\new_[30839]_  | ~\new_[29001]_  | ~\new_[30121]_ ;
  assign \new_[19395]_  = ~\new_[5997]_  | ~\new_[28728]_  | ~\new_[29968]_ ;
  assign \new_[19396]_  = ~\new_[6067]_  | ~\new_[29801]_  | ~\new_[30053]_ ;
  assign \new_[19397]_  = ~\new_[6212]_  | ~\new_[28832]_  | ~\new_[28609]_ ;
  assign \new_[19398]_  = ~\new_[5932]_  | ~\new_[28299]_  | ~\new_[30072]_ ;
  assign \new_[19399]_  = ~\new_[6193]_  | ~\new_[28163]_  | ~\new_[30212]_ ;
  assign \new_[19400]_  = ~\new_[21469]_  & (~\new_[27897]_  | ~\new_[28278]_ );
  assign \new_[19401]_  = ~\new_[21558]_  & (~\new_[28357]_  | ~\new_[28595]_ );
  assign \new_[19402]_  = ~\new_[20945]_  & (~\new_[28029]_  | ~\new_[28675]_ );
  assign \new_[19403]_  = ~\new_[28402]_  | ~\new_[31394]_ ;
  assign \new_[19404]_  = ~\new_[29508]_  | ~\new_[6084]_ ;
  assign \new_[19405]_  = ~\new_[30236]_  | ~\new_[5971]_ ;
  assign \new_[19406]_  = ~\new_[28816]_  | ~\new_[6041]_ ;
  assign \new_[19407]_  = ~\new_[29367]_  | ~\new_[6090]_ ;
  assign \new_[19408]_  = ~\new_[28232]_  | ~\new_[5973]_ ;
  assign \new_[19409]_  = ~\new_[29750]_  | ~\new_[31121]_ ;
  assign \new_[19410]_  = ~\new_[29848]_  | ~\new_[5969]_ ;
  assign \new_[19411]_  = ~\new_[28232]_  | ~\new_[5972]_ ;
  assign \new_[19412]_  = ~\new_[30206]_  | ~\new_[5972]_ ;
  assign \new_[19413]_  = ~\new_[28999]_  | ~\new_[6000]_ ;
  assign \new_[19414]_  = ~\new_[30251]_  | ~\new_[5982]_ ;
  assign \new_[19415]_  = ~\new_[30308]_  | ~\new_[5986]_ ;
  assign \new_[19416]_  = ~\new_[29290]_  | ~\new_[5990]_ ;
  assign \new_[19417]_  = ~\new_[28816]_  | ~\new_[5966]_ ;
  assign \new_[19418]_  = ~\new_[28052]_  | ~\new_[6268]_ ;
  assign \new_[19419]_  = ~\new_[30078]_  | ~\new_[6088]_ ;
  assign \new_[19420]_  = ~\new_[28052]_  | ~\new_[5995]_ ;
  assign \new_[19421]_  = ~\new_[28402]_  | ~\new_[31033]_ ;
  assign \new_[19422]_  = ~\new_[29227]_  | ~\new_[6067]_ ;
  assign \new_[19423]_  = ~\new_[28397]_  | ~\new_[5910]_ ;
  assign \new_[19424]_  = ~\new_[28982]_  | ~\new_[6056]_ ;
  assign \new_[19425]_  = ~\new_[29814]_  | ~\new_[5898]_ ;
  assign \new_[19426]_  = ~\new_[30253]_  | ~\new_[5970]_ ;
  assign \new_[19427]_  = ~\new_[29573]_  | ~\new_[6067]_ ;
  assign \new_[19428]_  = ~\new_[29652]_  | ~\new_[6080]_ ;
  assign \new_[19429]_  = ~\new_[30253]_  | ~\new_[6096]_ ;
  assign \new_[19430]_  = ~\new_[29508]_  | ~\new_[6186]_ ;
  assign \new_[19431]_  = ~\new_[28397]_  | ~\new_[6037]_ ;
  assign \new_[19432]_  = ~\new_[28950]_  | ~\new_[6080]_ ;
  assign \new_[19433]_  = ~\new_[29508]_  | ~\new_[5928]_ ;
  assign \new_[19434]_  = ~\new_[28397]_  | ~\new_[6040]_ ;
  assign \new_[19435]_  = ~\new_[28933]_  | ~\new_[6202]_ ;
  assign \new_[19436]_  = ~\new_[29119]_  | ~\new_[6202]_ ;
  assign \new_[19437]_  = ~\new_[29166]_  | ~\new_[6091]_ ;
  assign \new_[19438]_  = ~\new_[30141]_  | ~\new_[5903]_ ;
  assign \new_[19439]_  = ~\new_[29394]_  | ~\new_[6042]_ ;
  assign \new_[19440]_  = ~\new_[29578]_  | ~\new_[6193]_ ;
  assign \new_[19441]_  = ~\new_[29096]_  | ~\new_[6087]_ ;
  assign \new_[19442]_  = ~\new_[30052]_  | ~\new_[5902]_ ;
  assign \new_[19443]_  = ~\new_[30253]_  | ~\new_[6199]_ ;
  assign \new_[19444]_  = ~\new_[29096]_  & ~\new_[30399]_ ;
  assign \new_[19445]_  = ~\new_[28993]_  | ~\new_[29150]_ ;
  assign \new_[19446]_  = ~\new_[28950]_  & ~\new_[28031]_ ;
  assign \new_[19447]_  = ~\new_[29166]_  & ~\new_[30148]_ ;
  assign \new_[19448]_  = ~\new_[29671]_  | ~\new_[6080]_ ;
  assign \new_[19449]_  = ~\new_[29882]_  | ~\new_[5906]_ ;
  assign \new_[19450]_  = ~\new_[29331]_  | ~\new_[6062]_ ;
  assign n8699 = m0_s2_cyc_o_reg;
  assign n8669 = m0_s6_cyc_o_reg;
  assign n8349 = m1_s15_cyc_o_reg;
  assign n8884 = m1_s4_cyc_o_reg;
  assign n8384 = m1_s8_cyc_o_reg;
  assign n8539 = m2_s10_cyc_o_reg;
  assign n8359 = m4_s10_cyc_o_reg;
  assign n8899 = m4_s12_cyc_o_reg;
  assign n8859 = m4_s8_cyc_o_reg;
  assign n8374 = m5_s10_cyc_o_reg;
  assign n8344 = m5_s12_cyc_o_reg;
  assign n8809 = m5_s15_cyc_o_reg;
  assign n8369 = m5_s8_cyc_o_reg;
  assign n8939 = m6_s12_cyc_o_reg;
  assign n8584 = m6_s4_cyc_o_reg;
  assign n8934 = m7_s11_cyc_o_reg;
  assign n8419 = m7_s5_cyc_o_reg;
  assign \new_[19468]_  = ~\new_[29055]_  | ~\new_[5910]_ ;
  assign \new_[19469]_  = ~\new_[21605]_  & ~\new_[23748]_ ;
  assign \new_[19470]_  = ~\new_[23887]_  & (~\new_[23266]_  | ~\new_[29357]_ );
  assign \new_[19471]_  = ~\new_[25116]_  & (~\new_[23194]_  | ~\new_[26550]_ );
  assign \new_[19472]_  = ~\new_[26948]_  & (~\new_[23249]_  | ~\new_[30296]_ );
  assign \new_[19473]_  = \new_[21612]_  & \new_[29448]_ ;
  assign \new_[19474]_  = ~\new_[27562]_  & (~\new_[23235]_  | ~\new_[30426]_ );
  assign \new_[19475]_  = \new_[21614]_  & \new_[29026]_ ;
  assign \new_[19476]_  = ~\new_[27615]_  & (~\new_[23215]_  | ~\new_[30139]_ );
  assign \new_[19477]_  = ~\new_[26393]_  & (~\new_[24496]_  | ~\new_[30083]_ );
  assign \new_[19478]_  = ~\new_[26409]_  & (~\new_[24485]_  | ~\new_[29783]_ );
  assign \new_[19479]_  = ~\new_[24862]_  & (~\new_[23212]_  | ~\new_[25475]_ );
  assign \new_[19480]_  = ~\new_[23873]_  & (~\new_[23202]_  | ~\new_[24487]_ );
  assign \new_[19481]_  = ~\new_[21591]_  | ~\new_[24632]_ ;
  assign \new_[19482]_  = ~\new_[26930]_  & (~\new_[23222]_  | ~\new_[26367]_ );
  assign \new_[19483]_  = ~\new_[24976]_  & (~\new_[23225]_  | ~\new_[24357]_ );
  assign \new_[19484]_  = ~\new_[25026]_  & (~\new_[23200]_  | ~\new_[26396]_ );
  assign \new_[19485]_  = ~\new_[27965]_  & (~\new_[23226]_  | ~\new_[29891]_ );
  assign \new_[19486]_  = ~\new_[24583]_  & (~\new_[23230]_  | ~\new_[30210]_ );
  assign \new_[19487]_  = ~\new_[27677]_  & (~\new_[23236]_  | ~\new_[29913]_ );
  assign \new_[19488]_  = \new_[21622]_  & \new_[29449]_ ;
  assign \new_[19489]_  = ~\new_[24937]_  & (~\new_[23207]_  | ~\new_[26212]_ );
  assign \new_[19490]_  = ~\new_[24998]_  & (~\new_[23250]_  | ~\new_[30730]_ );
  assign \new_[19491]_  = ~\new_[26960]_  & (~\new_[23243]_  | ~\new_[27506]_ );
  assign \new_[19492]_  = ~\new_[23920]_  & (~\new_[23278]_  | ~\new_[30363]_ );
  assign \new_[19493]_  = ~\new_[26998]_  & (~\new_[23219]_  | ~\new_[25357]_ );
  assign \new_[19494]_  = ~\new_[21601]_  & ~\new_[23692]_ ;
  assign \new_[19495]_  = ~\new_[25137]_  & (~\new_[24517]_  | ~\new_[24764]_ );
  assign \new_[19496]_  = ~\new_[24780]_  & (~\new_[23262]_  | ~\new_[30724]_ );
  assign \new_[19497]_  = \new_[21623]_  & \new_[29464]_ ;
  assign \new_[19498]_  = ~\new_[26826]_  & (~\new_[23221]_  | ~\new_[30213]_ );
  assign \new_[19499]_  = ~\new_[29375]_  & (~\new_[24947]_  | ~\new_[23740]_ );
  assign \new_[19500]_  = \new_[22117]_  | \new_[21610]_ ;
  assign \new_[19501]_  = \new_[22348]_  | \new_[21613]_ ;
  assign \new_[19502]_  = \new_[23420]_  | \new_[21617]_ ;
  assign \new_[19503]_  = \new_[22453]_  | \new_[21624]_ ;
  assign \new_[19504]_  = \new_[21981]_  | \new_[21608]_ ;
  assign \new_[19505]_  = ~\new_[21637]_  | (~\new_[23326]_  & ~\new_[30566]_ );
  assign \new_[19506]_  = ~\new_[20575]_ ;
  assign \new_[19507]_  = ~\new_[23210]_  | (~\new_[23327]_  & ~\new_[30557]_ );
  assign \new_[19508]_  = ~\new_[24166]_  | (~\new_[24646]_  & ~\new_[30028]_ );
  assign \new_[19509]_  = ~\new_[23253]_  | (~\new_[23329]_  & ~\new_[30682]_ );
  assign \new_[19510]_  = ~\new_[30269]_  | ~\new_[21588]_  | ~\new_[25080]_ ;
  assign \new_[19511]_  = ~\new_[28944]_  | ~\new_[31422]_ ;
  assign \new_[19512]_  = ~\new_[22101]_  | ~\new_[27904]_ ;
  assign \new_[19513]_  = ~\new_[29220]_  | (~\new_[23376]_  & ~\new_[26391]_ );
  assign \new_[19514]_  = ~\new_[30232]_  | (~\new_[23385]_  & ~\new_[26225]_ );
  assign \new_[19515]_  = ~\new_[30386]_  | (~\new_[23415]_  & ~\new_[26531]_ );
  assign \new_[19516]_  = ~\new_[28880]_  | (~\new_[23853]_  & ~\new_[25975]_ );
  assign \new_[19517]_  = ~\new_[29563]_  | (~\new_[23743]_  & ~\new_[26617]_ );
  assign \new_[19518]_  = ~\new_[29150]_  | (~\new_[23585]_  & ~\new_[24677]_ );
  assign \new_[19519]_  = ~\new_[29782]_  | (~\new_[23443]_  & ~\new_[28406]_ );
  assign \new_[19520]_  = ~\new_[30217]_  | (~\new_[23531]_  & ~\new_[26732]_ );
  assign \new_[19521]_  = ~\new_[29386]_  | (~\new_[23565]_  & ~\new_[24431]_ );
  assign \new_[19522]_  = ~\new_[30279]_  | (~\new_[23502]_  & ~\new_[24668]_ );
  assign \new_[19523]_  = ~\new_[30617]_  | (~\new_[23653]_  & ~\new_[24273]_ );
  assign \new_[19524]_  = ~\new_[28870]_  | (~\new_[23546]_  & ~\new_[26560]_ );
  assign \new_[19525]_  = ~\new_[22089]_  | ~\new_[29015]_ ;
  assign \new_[19526]_  = ~\new_[30636]_  | (~\new_[23587]_  & ~\new_[27580]_ );
  assign \new_[19527]_  = ~\new_[29506]_  | (~\new_[23730]_  & ~\new_[26209]_ );
  assign \new_[19528]_  = ~\new_[22105]_  | ~\new_[26940]_ ;
  assign \new_[19529]_  = ~\new_[30158]_  | (~\new_[23695]_  & ~\new_[25674]_ );
  assign \new_[19530]_  = ~\new_[28926]_  | (~\new_[23805]_  & ~\new_[26308]_ );
  assign \new_[19531]_  = ~\new_[29967]_  | (~\new_[23557]_  & ~\new_[28572]_ );
  assign \new_[19532]_  = ~\new_[22098]_  | ~\new_[29972]_ ;
  assign \new_[19533]_  = ~\new_[28371]_  | (~\new_[23868]_  & ~\new_[24586]_ );
  assign \new_[19534]_  = ~\new_[30152]_  | ~\new_[21989]_  | ~\new_[30283]_ ;
  assign \new_[19535]_  = \new_[20539]_ ;
  assign \new_[19536]_  = ~\new_[20539]_ ;
  assign \new_[19537]_  = \new_[20539]_ ;
  assign \new_[19538]_  = \new_[22078]_  | \new_[30598]_ ;
  assign \new_[19539]_  = ~\new_[26931]_  & ~\new_[21867]_ ;
  assign \new_[19540]_  = ~\new_[25114]_  | ~\new_[21918]_ ;
  assign \new_[19541]_  = ~\new_[24817]_  | ~\new_[21919]_ ;
  assign \new_[19542]_  = ~\new_[20571]_ ;
  assign \new_[19543]_  = ~\new_[20542]_ ;
  assign \new_[19544]_  = \new_[26947]_  & \new_[21924]_ ;
  assign \new_[19545]_  = ~\new_[20543]_ ;
  assign \new_[19546]_  = ~\new_[20544]_ ;
  assign \new_[19547]_  = \new_[23874]_  & \new_[21920]_ ;
  assign \new_[19548]_  = ~\new_[20545]_ ;
  assign \new_[19549]_  = ~\new_[22012]_  & ~\new_[25182]_ ;
  assign \new_[19550]_  = ~\new_[29907]_  & (~\new_[23939]_  | ~\new_[24826]_ );
  assign \new_[19551]_  = ~\new_[21993]_  & ~\new_[24388]_ ;
  assign \new_[19552]_  = ~\new_[23089]_  & ~\new_[21671]_ ;
  assign \new_[19553]_  = ~\new_[29810]_  & (~\new_[23407]_  | ~\new_[24985]_ );
  assign \new_[19554]_  = \new_[24860]_  & \new_[21709]_ ;
  assign \new_[19555]_  = ~\new_[22019]_  & ~\new_[23074]_ ;
  assign \new_[19556]_  = ~\new_[20547]_ ;
  assign \new_[19557]_  = \new_[20547]_ ;
  assign \new_[19558]_  = ~\new_[20550]_ ;
  assign \new_[19559]_  = ~\new_[23441]_  & ~\new_[21738]_ ;
  assign \new_[19560]_  = ~\new_[20551]_ ;
  assign \new_[19561]_  = \new_[20551]_ ;
  assign \new_[19562]_  = ~\new_[23089]_  & ~\new_[21740]_ ;
  assign \new_[19563]_  = ~\new_[23818]_  & ~\new_[21742]_ ;
  assign \new_[19564]_  = ~\new_[20552]_ ;
  assign \new_[19565]_  = ~\new_[24956]_  & ~\new_[21867]_ ;
  assign \new_[19566]_  = \new_[24907]_  & \new_[21751]_ ;
  assign \new_[19567]_  = ~\new_[26956]_  & ~\new_[21695]_ ;
  assign \new_[19568]_  = ~\new_[25114]_  & ~\new_[21748]_ ;
  assign \new_[19569]_  = \new_[24817]_  | \new_[21749]_ ;
  assign \new_[19570]_  = ~\new_[20555]_ ;
  assign \new_[19571]_  = ~\new_[26947]_  & ~\new_[21847]_ ;
  assign \new_[19572]_  = \new_[24860]_  & \new_[21746]_ ;
  assign \new_[19573]_  = \new_[22090]_  | \new_[30185]_ ;
  assign \new_[19574]_  = ~\new_[30275]_  & (~\new_[23450]_  | ~\new_[25051]_ );
  assign \new_[19575]_  = ~\new_[26413]_  & ~\new_[21769]_ ;
  assign \new_[19576]_  = \new_[22094]_  | \new_[30515]_ ;
  assign \new_[19577]_  = ~\new_[26517]_  & ~\new_[21881]_ ;
  assign \new_[19578]_  = ~\new_[22007]_  & ~\new_[26307]_ ;
  assign \new_[19579]_  = \new_[22084]_  | \new_[30651]_ ;
  assign \new_[19580]_  = ~\new_[22005]_  & ~\new_[23181]_ ;
  assign \new_[19581]_  = ~\new_[25999]_  & ~\new_[21734]_ ;
  assign \new_[19582]_  = ~\new_[24269]_  | ~\new_[22004]_ ;
  assign \new_[19583]_  = ~\new_[20560]_ ;
  assign \new_[19584]_  = ~\new_[24860]_  & ~\new_[21737]_ ;
  assign \new_[19585]_  = \new_[23472]_  | \new_[21881]_ ;
  assign \new_[19586]_  = ~\new_[24907]_  & ~\new_[21739]_ ;
  assign \new_[19587]_  = ~\new_[22128]_  & ~\new_[21740]_ ;
  assign \new_[19588]_  = ~\new_[25113]_  & ~\new_[21742]_ ;
  assign \new_[19589]_  = ~\new_[24956]_  | ~\new_[24371]_ ;
  assign \new_[19590]_  = ~\new_[23874]_  & ~\new_[22955]_ ;
  assign \new_[19591]_  = \new_[22095]_  | \new_[30063]_ ;
  assign \new_[19592]_  = ~\new_[29792]_  & (~\new_[23875]_  | ~\new_[25004]_ );
  assign \new_[19593]_  = ~\new_[29157]_  & (~\new_[23637]_  | ~\new_[23641]_ );
  assign \new_[19594]_  = \new_[22083]_  | \new_[30564]_ ;
  assign \new_[19595]_  = ~\new_[25024]_  & ~\new_[21847]_ ;
  assign \new_[19596]_  = ~\new_[20567]_ ;
  assign \new_[19597]_  = \new_[20567]_ ;
  assign \new_[19598]_  = ~\new_[20568]_ ;
  assign \new_[19599]_  = ~\new_[20568]_ ;
  assign \new_[19600]_  = ~\new_[20568]_ ;
  assign \new_[19601]_  = \new_[22092]_  | \new_[30309]_ ;
  assign \new_[19602]_  = ~\new_[29997]_  & (~\new_[23832]_  | ~\new_[24700]_ );
  assign \new_[19603]_  = ~\new_[23281]_  & ~\new_[22875]_ ;
  assign \new_[19604]_  = \new_[22093]_  | \new_[30225]_ ;
  assign \new_[19605]_  = ~\new_[6038]_  | ~\new_[28046]_  | ~\new_[29597]_ ;
  assign \new_[19606]_  = ~\new_[20570]_ ;
  assign \new_[19607]_  = ~\new_[24956]_  | ~\new_[21917]_ ;
  assign \new_[19608]_  = \new_[23577]_  & \new_[21917]_ ;
  assign \new_[19609]_  = \new_[26849]_  & \new_[21918]_ ;
  assign \new_[19610]_  = ~\new_[26881]_  | ~\new_[21919]_ ;
  assign \new_[19611]_  = \new_[25024]_  & \new_[21924]_ ;
  assign \new_[19612]_  = ~\new_[20549]_ ;
  assign \new_[19613]_  = ~\new_[20549]_ ;
  assign \new_[19614]_  = ~\new_[20549]_ ;
  assign \new_[19615]_  = ~\new_[26956]_  & ~\new_[21925]_ ;
  assign \new_[19616]_  = ~\new_[30444]_  | ~\new_[22025]_  | ~\new_[30352]_ ;
  assign \new_[19617]_  = ~\new_[20541]_ ;
  assign \new_[19618]_  = \new_[20541]_ ;
  assign \new_[19619]_  = \new_[20541]_ ;
  assign \new_[19620]_  = ~\new_[30786]_  | ~\new_[22071]_  | ~\new_[29813]_ ;
  assign \new_[19621]_  = ~\new_[24610]_  & ~\new_[21976]_ ;
  assign \new_[19622]_  = ~\new_[20572]_ ;
  assign \new_[19623]_  = ~\new_[20573]_ ;
  assign \new_[19624]_  = ~\new_[20573]_ ;
  assign \new_[19625]_  = \new_[20573]_ ;
  assign \new_[19626]_  = \new_[20573]_ ;
  assign \new_[19627]_  = ~\new_[23529]_  & ~\new_[21769]_ ;
  assign \new_[19628]_  = ~\new_[22128]_  & ~\new_[21671]_ ;
  assign \new_[19629]_  = \new_[20575]_ ;
  assign \new_[19630]_  = \new_[20575]_ ;
  assign \new_[19631]_  = ~\new_[23488]_  | ~\new_[21751]_ ;
  assign \new_[19632]_  = \new_[26897]_  & \new_[21709]_ ;
  assign \new_[19633]_  = ~\new_[25113]_  & ~\new_[22116]_ ;
  assign \new_[19634]_  = ~\new_[20576]_ ;
  assign \new_[19635]_  = \new_[24732]_  | \new_[22955]_ ;
  assign \new_[19636]_  = ~\new_[25063]_  & ~\new_[21695]_ ;
  assign \new_[19637]_  = ~\new_[23818]_  & ~\new_[22116]_ ;
  assign \new_[19638]_  = ~\new_[26881]_  & ~\new_[21749]_ ;
  assign \new_[19639]_  = ~\new_[26849]_  & ~\new_[21748]_ ;
  assign \new_[19640]_  = ~\new_[22017]_  & ~\new_[23144]_ ;
  assign \new_[19641]_  = ~\new_[20578]_ ;
  assign \new_[19642]_  = \new_[20578]_ ;
  assign \new_[19643]_  = ~\new_[23848]_  & ~\new_[21976]_ ;
  assign \new_[19644]_  = ~\new_[29354]_  & (~\new_[23847]_  | ~\new_[23846]_ );
  assign \new_[19645]_  = \new_[22100]_  | \new_[30708]_ ;
  assign \new_[19646]_  = ~\new_[21990]_  & ~\new_[24960]_ ;
  assign \new_[19647]_  = ~\new_[20580]_ ;
  assign \new_[19648]_  = \new_[20580]_ ;
  assign \new_[19649]_  = ~\new_[30416]_  | ~\new_[30152]_  | ~\new_[21640]_  | ~\new_[28045]_ ;
  assign \new_[19650]_  = ~\new_[30784]_  | ~\new_[27802]_  | ~\new_[21627]_  | ~\new_[28337]_ ;
  assign \new_[19651]_  = ~\new_[30721]_  | ~\new_[26655]_  | ~\new_[21626]_  | ~\new_[30446]_ ;
  assign \new_[19652]_  = ~\new_[30695]_  | ~\new_[30011]_  | ~\new_[21813]_  | ~\new_[30731]_ ;
  assign \new_[19653]_  = ~\new_[30750]_  | ~\new_[27787]_  | ~\new_[23190]_  | ~\new_[30000]_ ;
  assign \new_[19654]_  = ~\new_[30538]_  | ~\new_[30491]_  | ~\new_[21630]_  | ~\new_[30842]_ ;
  assign \new_[19655]_  = ~\new_[30789]_  | ~\new_[29537]_  | ~\new_[21631]_  | ~\new_[30205]_ ;
  assign \new_[19656]_  = ~\new_[30726]_  | ~\new_[28069]_  | ~\new_[21625]_  | ~\new_[30582]_ ;
  assign \new_[19657]_  = ~\new_[30799]_  | ~\new_[29798]_  | ~\new_[21650]_  | ~\new_[30586]_ ;
  assign \new_[19658]_  = ~\new_[30820]_  | ~\new_[30735]_  | ~\new_[23075]_  | ~\new_[30764]_ ;
  assign \new_[19659]_  = ~\new_[24827]_  & (~\new_[26835]_  | ~\new_[23889]_ );
  assign \new_[19660]_  = ~\new_[30612]_  & (~\new_[23886]_  | ~\new_[24797]_ );
  assign \new_[19661]_  = ~\new_[30044]_  & (~\new_[23900]_  | ~\new_[24905]_ );
  assign \new_[19662]_  = ~\new_[23339]_  & (~\new_[24465]_  | ~\new_[25153]_ );
  assign \new_[19663]_  = ~\new_[30225]_  & (~\new_[23904]_  | ~\new_[28306]_ );
  assign \new_[19664]_  = ~\new_[28069]_  | ~\new_[21606]_  | ~\new_[30020]_ ;
  assign \new_[19665]_  = ~\new_[30541]_  & (~\new_[23358]_  | ~\new_[24816]_ );
  assign \new_[19666]_  = ~\new_[23382]_  & (~\new_[26693]_  | ~\new_[23167]_ );
  assign \new_[19667]_  = ~\new_[30694]_  & (~\new_[23929]_  | ~\new_[24824]_ );
  assign \new_[19668]_  = ~\new_[30095]_  & (~\new_[24828]_  | ~\new_[23373]_ );
  assign \new_[19669]_  = ~\new_[29743]_  & (~\new_[26889]_  | ~\new_[23380]_ );
  assign \new_[19670]_  = ~\new_[20590]_ ;
  assign \new_[19671]_  = ~\new_[30788]_  & (~\new_[23395]_  | ~\new_[23437]_ );
  assign \new_[19672]_  = ~\new_[30575]_  & (~\new_[23893]_  | ~\new_[24843]_ );
  assign \new_[19673]_  = ~\new_[30168]_  & (~\new_[23605]_  | ~\new_[23410]_ );
  assign \new_[19674]_  = ~\new_[26627]_  & (~\new_[23411]_  | ~\new_[23412]_ );
  assign \new_[19675]_  = ~\new_[20595]_ ;
  assign \new_[19676]_  = ~\new_[23739]_  & (~\new_[24399]_  | ~\new_[23930]_ );
  assign \new_[19677]_  = ~\new_[30648]_  & (~\new_[23426]_  | ~\new_[24886]_ );
  assign \new_[19678]_  = ~\new_[20600]_ ;
  assign \new_[19679]_  = ~\new_[29952]_  & (~\new_[23357]_  | ~\new_[23445]_ );
  assign \new_[19680]_  = ~\new_[22280]_  & (~\new_[26260]_  | ~\new_[24600]_ );
  assign \new_[19681]_  = ~\new_[30185]_  & (~\new_[23909]_  | ~\new_[28772]_ );
  assign \new_[19682]_  = ~\new_[30719]_  | ~\new_[26318]_  | ~\new_[23451]_  | ~\new_[27506]_ ;
  assign \new_[19683]_  = ~\new_[30022]_  | ~\new_[22003]_  | ~\new_[29782]_ ;
  assign \new_[19684]_  = ~\new_[30564]_  & (~\new_[23926]_  | ~\new_[23745]_ );
  assign \new_[19685]_  = ~\new_[20607]_ ;
  assign \new_[19686]_  = ~\new_[20608]_ ;
  assign \new_[19687]_  = ~\new_[28027]_  & (~\new_[23678]_  | ~\new_[24897]_ );
  assign \new_[19688]_  = ~\new_[23751]_  & (~\new_[23955]_  | ~\new_[26994]_ );
  assign \new_[19689]_  = ~\new_[29013]_  & (~\new_[24901]_  | ~\new_[23487]_ );
  assign \new_[19690]_  = ~\new_[30130]_  & (~\new_[25199]_  | ~\new_[23352]_ );
  assign \new_[19691]_  = ~\new_[30185]_  & (~\new_[23909]_  | ~\new_[23496]_ );
  assign \new_[19692]_  = ~\new_[20611]_ ;
  assign \new_[19693]_  = ~\new_[29776]_  & (~\new_[23500]_  | ~\new_[23482]_ );
  assign \new_[19694]_  = ~\new_[30118]_  & (~\new_[23706]_  | ~\new_[23677]_ );
  assign \new_[19695]_  = ~\new_[28849]_  & (~\new_[24921]_  | ~\new_[23568]_ );
  assign \new_[19696]_  = ~\new_[21768]_  | ~\new_[30207]_ ;
  assign \new_[19697]_  = ~\new_[29968]_  & (~\new_[23661]_  | ~\new_[23476]_ );
  assign \new_[19698]_  = ~\new_[27897]_  & (~\new_[24918]_  | ~\new_[23511]_ );
  assign \new_[19699]_  = ~\new_[30675]_  & (~\new_[23933]_  | ~\new_[26408]_ );
  assign \new_[19700]_  = ~\new_[30301]_  & (~\new_[24939]_  | ~\new_[23541]_ );
  assign \new_[19701]_  = ~\new_[29371]_  & (~\new_[23769]_  | ~\new_[24911]_ );
  assign \new_[19702]_  = ~\new_[30247]_  & (~\new_[23550]_  | ~\new_[23454]_ );
  assign \new_[19703]_  = ~\new_[28829]_  & (~\new_[25077]_  | ~\new_[23742]_ );
  assign \new_[19704]_  = ~\new_[26660]_  & (~\new_[23558]_  | ~\new_[23579]_ );
  assign \new_[19705]_  = ~\new_[22260]_  & (~\new_[24365]_  | ~\new_[25185]_ );
  assign \new_[19706]_  = ~\new_[30651]_  & (~\new_[23907]_  | ~\new_[26059]_ );
  assign \new_[19707]_  = ~\new_[26651]_  & (~\new_[23580]_  | ~\new_[23515]_ );
  assign \new_[19708]_  = ~\new_[30002]_  & (~\new_[23591]_  | ~\new_[25076]_ );
  assign \new_[19709]_  = ~\new_[30127]_  | ~\new_[5904]_ ;
  assign \new_[19710]_  = ~\new_[30696]_  & (~\new_[23949]_  | ~\new_[25106]_ );
  assign \new_[19711]_  = ~\new_[30302]_  & (~\new_[23606]_  | ~\new_[23607]_ );
  assign \new_[19712]_  = ~\new_[28166]_  & (~\new_[23599]_  | ~\new_[25086]_ );
  assign \new_[19713]_  = ~\new_[29064]_  | ~\new_[22014]_  | ~\new_[30595]_ ;
  assign \new_[19714]_  = ~\new_[30651]_  & (~\new_[23907]_  | ~\new_[28550]_ );
  assign \new_[19715]_  = ~\new_[22194]_  & (~\new_[23267]_  | ~\new_[24691]_ );
  assign \new_[19716]_  = ~\new_[30780]_  & (~\new_[23892]_  | ~\new_[26097]_ );
  assign \new_[19717]_  = ~\new_[23391]_  & (~\new_[24462]_  | ~\new_[23950]_ );
  assign \new_[19718]_  = ~\new_[22186]_  & (~\new_[23134]_  | ~\new_[23912]_ );
  assign \new_[19719]_  = ~\new_[20617]_ ;
  assign \new_[19720]_  = ~\new_[30746]_  & (~\new_[23561]_  | ~\new_[25071]_ );
  assign \new_[19721]_  = ~\new_[29790]_  & (~\new_[23681]_  | ~\new_[25380]_ );
  assign \new_[19722]_  = ~\new_[28935]_  | ~\new_[22075]_  | ~\new_[30702]_ ;
  assign \new_[19723]_  = ~\new_[28950]_  & (~\new_[23918]_  | ~\new_[28305]_ );
  assign \new_[19724]_  = ~\new_[30501]_  & (~\new_[23948]_  | ~\new_[25042]_ );
  assign \new_[19725]_  = ~\new_[29926]_  & (~\new_[23691]_  | ~\new_[24883]_ );
  assign \new_[19726]_  = ~\new_[29384]_  & (~\new_[23825]_  | ~\new_[25047]_ );
  assign \new_[19727]_  = ~\new_[23559]_  & (~\new_[28353]_  | ~\new_[23906]_ );
  assign \new_[19728]_  = ~\new_[30628]_  | ~\new_[22006]_  | ~\new_[29967]_ ;
  assign \new_[19729]_  = ~\new_[22316]_  & (~\new_[26285]_  | ~\new_[25197]_ );
  assign \new_[19730]_  = ~\new_[30718]_  & (~\new_[23710]_  | ~\new_[23749]_ );
  assign \new_[19731]_  = ~\new_[28029]_  & (~\new_[23821]_  | ~\new_[23723]_ );
  assign \new_[19732]_  = ~\new_[30564]_  & (~\new_[23926]_  | ~\new_[28167]_ );
  assign \new_[19733]_  = ~\new_[22440]_  & (~\new_[24444]_  | ~\new_[23919]_ );
  assign \new_[19734]_  = ~\new_[30044]_  & (~\new_[23900]_  | ~\new_[28522]_ );
  assign \new_[19735]_  = ~\new_[28859]_  & (~\new_[24935]_  | ~\new_[23650]_ );
  assign \new_[19736]_  = ~\new_[30328]_  & (~\new_[23755]_  | ~\new_[23548]_ );
  assign \new_[19737]_  = ~\new_[30737]_  & (~\new_[23804]_  | ~\new_[23708]_ );
  assign \new_[19738]_  = ~\new_[30502]_  & (~\new_[23346]_  | ~\new_[23782]_ );
  assign \new_[19739]_  = ~\new_[22245]_  & (~\new_[24410]_  | ~\new_[25207]_ );
  assign \new_[19740]_  = ~\new_[30225]_  & (~\new_[23904]_  | ~\new_[23850]_ );
  assign n7769 = ~\new_[29240]_  | ~\new_[22029]_ ;
  assign n7704 = ~\new_[29285]_  | ~\new_[22043]_ ;
  assign n7764 = ~\new_[29683]_  | ~\new_[22069]_ ;
  assign n7754 = ~\new_[29307]_  | ~\new_[22053]_ ;
  assign n7749 = ~\new_[29418]_  | ~\new_[22062]_ ;
  assign n7709 = ~\new_[29267]_  | ~\new_[22067]_ ;
  assign n7759 = ~\new_[29245]_  | ~\new_[22037]_ ;
  assign \new_[19748]_  = ~\new_[28950]_  & (~\new_[23918]_  | ~\new_[25036]_ );
  assign \new_[19749]_  = ~\new_[30543]_  & (~\new_[23903]_  | ~\new_[25060]_ );
  assign \new_[19750]_  = ~\new_[30708]_  & (~\new_[23896]_  | ~\new_[23849]_ );
  assign \new_[19751]_  = ~\new_[20634]_ ;
  assign \new_[19752]_  = ~\new_[30708]_  & (~\new_[23896]_  | ~\new_[28241]_ );
  assign \new_[19753]_  = ~\new_[30837]_  & (~\new_[23915]_  | ~\new_[25059]_ );
  assign \new_[19754]_  = ~\new_[22444]_  & (~\new_[24275]_  | ~\new_[25270]_ );
  assign \new_[19755]_  = ~\new_[28191]_  & (~\new_[24799]_  | ~\new_[23341]_ );
  assign \new_[19756]_  = ~\new_[29916]_  & (~\new_[23927]_  | ~\new_[28708]_ );
  assign \new_[19757]_  = ~\new_[30735]_  | ~\new_[22077]_  | ~\new_[29118]_ ;
  assign \new_[19758]_  = ~\new_[30706]_  & (~\new_[23783]_  | ~\new_[23876]_ );
  assign \new_[19759]_  = ~\new_[25147]_  & (~\new_[23956]_  | ~\new_[25214]_ );
  assign \new_[19760]_  = ~\new_[29119]_  & (~\new_[23954]_  | ~\new_[24726]_ );
  assign \new_[19761]_  = ~\new_[29119]_  & (~\new_[23954]_  | ~\new_[28740]_ );
  assign \new_[19762]_  = ~\new_[24774]_  & (~\new_[23344]_  | ~\new_[29029]_ );
  assign \new_[19763]_  = \new_[21644]_  & \new_[26374]_ ;
  assign \new_[19764]_  = ~\new_[24264]_  & (~\new_[23374]_  | ~\new_[29291]_ );
  assign \new_[19765]_  = ~\new_[24286]_  & (~\new_[23689]_  | ~\new_[28894]_ );
  assign \new_[19766]_  = \new_[21666]_  & \new_[26292]_ ;
  assign \new_[19767]_  = \new_[21833]_  & \new_[26443]_ ;
  assign \new_[19768]_  = ~\new_[24433]_  & (~\new_[23383]_  | ~\new_[29223]_ );
  assign \new_[19769]_  = ~\new_[24508]_  & (~\new_[23696]_  | ~\new_[30229]_ );
  assign \new_[19770]_  = ~\new_[26077]_  & (~\new_[23083]_  | ~\new_[30599]_ );
  assign \new_[19771]_  = \new_[21744]_  & \new_[27577]_ ;
  assign \new_[19772]_  = ~\new_[23126]_  & (~\new_[23490]_  | ~\new_[29623]_ );
  assign \new_[19773]_  = ~\new_[24419]_  & (~\new_[23501]_  | ~\new_[28934]_ );
  assign \new_[19774]_  = ~\new_[24408]_  & (~\new_[23416]_  | ~\new_[28918]_ );
  assign \new_[19775]_  = \new_[21696]_  & \new_[26083]_ ;
  assign \new_[19776]_  = ~\new_[26273]_  & (~\new_[23425]_  | ~\new_[30222]_ );
  assign \new_[19777]_  = ~\new_[26234]_  & (~\new_[23614]_  | ~\new_[29771]_ );
  assign \new_[19778]_  = ~\new_[24292]_  & (~\new_[23852]_  | ~\new_[29381]_ );
  assign \new_[19779]_  = ~\new_[26253]_  & (~\new_[23575]_  | ~\new_[28836]_ );
  assign \new_[19780]_  = \new_[21723]_  & \new_[26300]_ ;
  assign \new_[19781]_  = ~\new_[28514]_  & (~\new_[23797]_  | ~\new_[30525]_ );
  assign \new_[19782]_  = ~\new_[27722]_  & (~\new_[23643]_  | ~\new_[30269]_ );
  assign \new_[19783]_  = ~\new_[26132]_  & (~\new_[23430]_  | ~\new_[30242]_ );
  assign \new_[19784]_  = ~\new_[24529]_  & (~\new_[23494]_  | ~\new_[29276]_ );
  assign \new_[19785]_  = \new_[22938]_  & \new_[27596]_ ;
  assign \new_[19786]_  = ~\new_[30840]_  | ~\new_[5928]_ ;
  assign \new_[19787]_  = \new_[21785]_  & \new_[26347]_ ;
  assign \new_[19788]_  = ~\new_[23081]_  & (~\new_[23762]_  | ~\new_[28110]_ );
  assign \new_[19789]_  = ~\new_[24280]_  & (~\new_[23757]_  | ~\new_[28818]_ );
  assign \new_[19790]_  = \new_[21797]_  & \new_[27635]_ ;
  assign \new_[19791]_  = ~\new_[26397]_  & (~\new_[23554]_  | ~\new_[29332]_ );
  assign \new_[19792]_  = ~\new_[26470]_  & (~\new_[23728]_  | ~\new_[30198]_ );
  assign \new_[19793]_  = \new_[21843]_  & \new_[27568]_ ;
  assign \new_[19794]_  = ~\new_[24468]_  & (~\new_[23578]_  | ~\new_[29020]_ );
  assign \new_[19795]_  = ~\new_[24403]_  & (~\new_[23784]_  | ~\new_[29569]_ );
  assign \new_[19796]_  = ~\new_[25829]_  & (~\new_[23513]_  | ~\new_[28865]_ );
  assign \new_[19797]_  = ~\new_[23258]_  & (~\new_[23774]_  | ~\new_[29589]_ );
  assign \new_[19798]_  = ~\new_[24946]_  & (~\new_[23722]_  | ~\new_[29410]_ );
  assign \new_[19799]_  = ~\new_[27728]_  & (~\new_[23597]_  | ~\new_[29869]_ );
  assign \new_[19800]_  = ~\new_[26398]_  & (~\new_[23553]_  | ~\new_[29421]_ );
  assign \new_[19801]_  = ~\new_[23077]_  & (~\new_[23629]_  | ~\new_[28595]_ );
  assign \new_[19802]_  = \new_[21660]_  & \new_[26395]_ ;
  assign \new_[19803]_  = ~\new_[27566]_  & (~\new_[24893]_  | ~\new_[28278]_ );
  assign \new_[19804]_  = \new_[21829]_  & \new_[26333]_ ;
  assign \new_[19805]_  = ~\new_[22496]_  & (~\new_[23363]_  | ~\new_[29987]_ );
  assign \new_[19806]_  = \new_[21716]_  & \new_[27561]_ ;
  assign \new_[19807]_  = \new_[21837]_  & \new_[26360]_ ;
  assign \new_[19808]_  = ~\new_[24390]_  & (~\new_[23610]_  | ~\new_[29145]_ );
  assign \new_[19809]_  = ~\new_[22905]_  & (~\new_[23808]_  | ~\new_[27997]_ );
  assign \new_[19810]_  = \new_[21906]_  & \new_[26745]_ ;
  assign \new_[19811]_  = ~\new_[24405]_  & (~\new_[23758]_  | ~\new_[29583]_ );
  assign \new_[19812]_  = ~\new_[24452]_  & (~\new_[24028]_  | ~\new_[29042]_ );
  assign \new_[19813]_  = \new_[21871]_  & \new_[27474]_ ;
  assign \new_[19814]_  = \new_[21645]_  & \new_[27691]_ ;
  assign \new_[19815]_  = ~\new_[24470]_  & (~\new_[23865]_  | ~\new_[29130]_ );
  assign \new_[19816]_  = ~\new_[22918]_  & (~\new_[23855]_  | ~\new_[29151]_ );
  assign \new_[19817]_  = \new_[21985]_  & \new_[27546]_ ;
  assign \new_[19818]_  = ~\new_[21941]_  & ~\new_[29853]_ ;
  assign \new_[19819]_  = ~\new_[30352]_  | (~\new_[23738]_  & ~\new_[23819]_ );
  assign \new_[19820]_  = ~\new_[29784]_  & (~\new_[23792]_  | ~\new_[24806]_ );
  assign \new_[19821]_  = ~\new_[30736]_  & (~\new_[23780]_  | ~\new_[26680]_ );
  assign \new_[19822]_  = ~\new_[30726]_  | (~\new_[23354]_  & ~\new_[26600]_ );
  assign \new_[19823]_  = ~\new_[21886]_  | ~\new_[29527]_ ;
  assign \new_[19824]_  = ~\new_[28908]_  | (~\new_[23771]_  & ~\new_[23772]_ );
  assign \new_[19825]_  = ~\new_[21651]_  & ~\new_[29855]_ ;
  assign \new_[19826]_  = ~\new_[28908]_  | (~\new_[23367]_  & ~\new_[28992]_ );
  assign \new_[19827]_  = ~\new_[30425]_  & (~\new_[23705]_  | ~\new_[26618]_ );
  assign \new_[19828]_  = ~\new_[28844]_  | (~\new_[23709]_  & ~\new_[29229]_ );
  assign \new_[19829]_  = ~\new_[21679]_  | ~\new_[29320]_ ;
  assign \new_[19830]_  = ~\new_[29112]_  | (~\new_[23396]_  & ~\new_[23394]_ );
  assign \new_[19831]_  = ~\new_[21822]_  & ~\new_[29100]_ ;
  assign \new_[19832]_  = ~\new_[29112]_  | (~\new_[23644]_  & ~\new_[29541]_ );
  assign \new_[19833]_  = ~\new_[30676]_  | (~\new_[25993]_  & ~\new_[23402]_ );
  assign \new_[19834]_  = ~\new_[29260]_  | (~\new_[23609]_  & ~\new_[24855]_ );
  assign \new_[19835]_  = ~\new_[21728]_  | ~\new_[29228]_ ;
  assign \new_[19836]_  = ~\new_[28968]_  | (~\new_[23460]_  & ~\new_[23467]_ );
  assign \new_[19837]_  = ~\new_[21713]_  & ~\new_[30389]_ ;
  assign \new_[19838]_  = ~\new_[28968]_  | (~\new_[23435]_  & ~\new_[29217]_ );
  assign \new_[19839]_  = ~\new_[30573]_  | (~\new_[24920]_  & ~\new_[23438]_ );
  assign \new_[19840]_  = ~\new_[29827]_  & (~\new_[23447]_  | ~\new_[23790]_ );
  assign \new_[19841]_  = ~\new_[30721]_  | (~\new_[23753]_  & ~\new_[24879]_ );
  assign \new_[19842]_  = ~\new_[28236]_  & (~\new_[23663]_  | ~\new_[23588]_ );
  assign \new_[19843]_  = ~\new_[28835]_  | (~\new_[23464]_  & ~\new_[23463]_ );
  assign \new_[19844]_  = ~\new_[30774]_  | (~\new_[23508]_  & ~\new_[23474]_ );
  assign \new_[19845]_  = ~\new_[30037]_  | (~\new_[23717]_  & ~\new_[25068]_ );
  assign \new_[19846]_  = ~\new_[21730]_  & ~\new_[29935]_ ;
  assign \new_[19847]_  = ~\new_[28718]_  & (~\new_[23598]_  | ~\new_[23613]_ );
  assign \new_[19848]_  = ~\new_[29977]_  | (~\new_[24506]_  & ~\new_[23603]_ );
  assign \new_[19849]_  = ~\new_[21811]_  & ~\new_[29648]_ ;
  assign \new_[19850]_  = ~\new_[30728]_  | (~\new_[23498]_  & ~\new_[24490]_ );
  assign \new_[19851]_  = ~\new_[30555]_  | (~\new_[24910]_  & ~\new_[23520]_ );
  assign \new_[19852]_  = ~\new_[30323]_  & (~\new_[23361]_  | ~\new_[23419]_ );
  assign \new_[19853]_  = ~\new_[21961]_  & ~\new_[28950]_ ;
  assign \new_[19854]_  = ~\new_[30538]_  | (~\new_[23601]_  & ~\new_[26511]_ );
  assign \new_[19855]_  = ~\new_[21762]_  & ~\new_[28982]_ ;
  assign \new_[19856]_  = ~\new_[30005]_  | (~\new_[23796]_  & ~\new_[29700]_ );
  assign \new_[19857]_  = ~\new_[30246]_  | (~\new_[23539]_  & ~\new_[23542]_ );
  assign \new_[19858]_  = ~\new_[30615]_  | (~\new_[23645]_  & ~\new_[23552]_ );
  assign \new_[19859]_  = ~\new_[21793]_  & ~\new_[30526]_ ;
  assign \new_[19860]_  = ~\new_[29633]_  | (~\new_[23795]_  & ~\new_[29115]_ );
  assign \new_[19861]_  = ~\new_[30574]_  | (~\new_[23583]_  & ~\new_[23534]_ );
  assign \new_[19862]_  = ~\new_[28911]_  | (~\new_[23581]_  & ~\new_[23632]_ );
  assign \new_[19863]_  = ~\new_[28911]_  | (~\new_[23794]_  & ~\new_[29254]_ );
  assign \new_[19864]_  = ~\new_[30173]_  & (~\new_[23741]_  | ~\new_[23756]_ );
  assign \new_[19865]_  = ~\new_[30014]_  & (~\new_[23623]_  | ~\new_[25005]_ );
  assign \new_[19866]_  = ~\new_[21707]_  | ~\new_[29721]_ ;
  assign \new_[19867]_  = ~\new_[29633]_  | (~\new_[23620]_  & ~\new_[23619]_ );
  assign \new_[19868]_  = ~\new_[28905]_  | (~\new_[23701]_  & ~\new_[23841]_ );
  assign \new_[19869]_  = ~\new_[21810]_  | ~\new_[29006]_ ;
  assign \new_[19870]_  = ~\new_[28864]_  | (~\new_[23574]_  & ~\new_[23799]_ );
  assign \new_[19871]_  = ~\new_[30086]_  | (~\new_[23641]_  & ~\new_[29157]_ );
  assign \new_[19872]_  = ~\new_[28864]_  | (~\new_[23724]_  & ~\new_[29101]_ );
  assign \new_[19873]_  = ~\new_[30775]_  | (~\new_[24919]_  & ~\new_[23646]_ );
  assign \new_[19874]_  = ~\new_[29802]_  | (~\new_[23697]_  & ~\new_[23863]_ );
  assign \new_[19875]_  = ~\new_[30784]_  | (~\new_[23881]_  & ~\new_[26945]_ );
  assign \new_[19876]_  = ~\new_[21812]_  | ~\new_[29695]_ ;
  assign \new_[19877]_  = ~\new_[28844]_  | (~\new_[23667]_  & ~\new_[23618]_ );
  assign \new_[19878]_  = ~\new_[21826]_  & ~\new_[29331]_ ;
  assign \new_[19879]_  = ~\new_[29272]_  & (~\new_[23343]_  | ~\new_[23455]_ );
  assign \new_[19880]_  = ~\new_[30240]_  & (~\new_[23654]_  | ~\new_[24844]_ );
  assign \new_[19881]_  = ~\new_[29813]_  | (~\new_[23806]_  & ~\new_[23814]_ );
  assign \new_[19882]_  = ~\new_[30630]_  | (~\new_[25040]_  & ~\new_[23809]_ );
  assign \new_[19883]_  = ~\new_[30400]_  & (~\new_[23810]_  | ~\new_[23820]_ );
  assign \new_[19884]_  = ~\new_[30084]_  | (~\new_[25120]_  & ~\new_[23815]_ );
  assign \new_[19885]_  = ~\new_[30647]_  | (~\new_[24999]_  & ~\new_[23985]_ );
  assign \new_[19886]_  = ~\new_[29189]_  | (~\new_[23713]_  & ~\new_[24016]_ );
  assign \new_[19887]_  = ~\new_[21986]_  & ~\new_[29898]_ ;
  assign \new_[19888]_  = ~\new_[30215]_  | (~\new_[23752]_  & ~\new_[25075]_ );
  assign \new_[19889]_  = ~\new_[30719]_  | (~\new_[24594]_  & ~\new_[23359]_ );
  assign \new_[19890]_  = ~\new_[29887]_  | (~\new_[23571]_  & ~\new_[23715]_ );
  assign \new_[19891]_  = ~\new_[30280]_  | (~\new_[23763]_  & ~\new_[29047]_ );
  assign \new_[19892]_  = ~\new_[30507]_  | (~\new_[23331]_  & ~\new_[26927]_ );
  assign \new_[19893]_  = ~\new_[30707]_  | (~\new_[23734]_  & ~\new_[23803]_ );
  assign \new_[19894]_  = ~\new_[28857]_  & (~\new_[23750]_  | ~\new_[23627]_ );
  assign \new_[19895]_  = ~\new_[30754]_  | (~\new_[24823]_  & ~\new_[23370]_ );
  assign \new_[19896]_  = ~\new_[30407]_  & (~\new_[23543]_  | ~\new_[23767]_ );
  assign \new_[19897]_  = ~\new_[29189]_  | (~\new_[23635]_  & ~\new_[29167]_ );
  assign \new_[19898]_  = ~\new_[29870]_  | (~\new_[23532]_  & ~\new_[24803]_ );
  assign \new_[19899]_  = ~\new_[28835]_  | (~\new_[23466]_  & ~\new_[29058]_ );
  assign \new_[19900]_  = ~\new_[30105]_  | (~\new_[25039]_  & ~\new_[29671]_ );
  assign \new_[19901]_  = ~\new_[21784]_  | ~\new_[29456]_ ;
  assign \new_[19902]_  = ~\new_[21855]_  & ~\new_[29096]_ ;
  assign \new_[19903]_  = ~\new_[21969]_  & ~\new_[29166]_ ;
  assign \new_[19904]_  = ~\new_[30123]_  | (~\new_[23846]_  & ~\new_[29354]_ );
  assign \new_[19905]_  = ~\new_[30262]_  | (~\new_[23854]_  & ~\new_[24846]_ );
  assign \new_[19906]_  = ~\new_[21975]_  & ~\new_[30003]_ ;
  assign \new_[19907]_  = ~\new_[29383]_  & (~\new_[23864]_  | ~\new_[24802]_ );
  assign \new_[19908]_  = ~\new_[30820]_  | (~\new_[23871]_  & ~\new_[27426]_ );
  assign \new_[19909]_  = ~\new_[30104]_  | (~\new_[23885]_  & ~\new_[25151]_ );
  assign \new_[19910]_  = ~\new_[21655]_  & ~\new_[29119]_ ;
  assign \new_[19911]_  = ~\new_[27660]_  & (~\new_[23899]_  | ~\new_[28575]_ );
  assign \new_[19912]_  = ~\new_[27739]_  & (~\new_[23891]_  | ~\new_[28222]_ );
  assign \new_[19913]_  = ~\new_[26304]_  & (~\new_[23923]_  | ~\new_[28631]_ );
  assign \new_[19914]_  = ~\new_[27631]_  & (~\new_[23913]_  | ~\new_[28474]_ );
  assign \new_[19915]_  = ~\new_[28659]_  & (~\new_[23897]_  | ~\new_[28500]_ );
  assign \new_[19916]_  = ~\new_[28577]_  & (~\new_[23910]_  | ~\new_[28108]_ );
  assign \new_[19917]_  = ~\new_[26286]_  & (~\new_[23925]_  | ~\new_[28181]_ );
  assign \new_[19918]_  = ~\new_[22912]_  & (~\new_[24537]_  | ~\new_[28498]_ );
  assign \new_[19919]_  = ~\new_[27805]_  & (~\new_[23902]_  | ~\new_[28373]_ );
  assign \new_[19920]_  = ~\new_[28401]_  & (~\new_[23888]_  | ~\new_[28412]_ );
  assign \new_[19921]_  = \new_[21639]_  & \new_[29500]_ ;
  assign \new_[19922]_  = ~\new_[29692]_  | (~\new_[23446]_  & ~\new_[26951]_ );
  assign \new_[19923]_  = ~\new_[23366]_  & (~\new_[24821]_  | ~\new_[24368]_ );
  assign \new_[19924]_  = \new_[21872]_  & \new_[29483]_ ;
  assign \new_[19925]_  = ~\new_[22232]_  & (~\new_[24074]_  | ~\new_[24333]_ );
  assign \new_[19926]_  = ~\new_[30316]_  | (~\new_[23379]_  & ~\new_[27679]_ );
  assign \new_[19927]_  = ~\new_[23398]_  & (~\new_[23227]_  | ~\new_[24459]_ );
  assign \new_[19928]_  = \new_[21690]_  & \new_[29294]_ ;
  assign \new_[19929]_  = \new_[21736]_  & \new_[29480]_ ;
  assign \new_[19930]_  = ~\new_[28857]_  & (~\new_[23627]_  | ~\new_[27951]_ );
  assign \new_[19931]_  = ~\new_[30574]_  | (~\new_[23534]_  & ~\new_[27388]_ );
  assign \new_[19932]_  = ~\new_[23434]_  & (~\new_[26557]_  | ~\new_[24514]_ );
  assign \new_[19933]_  = ~\new_[29827]_  & (~\new_[23790]_  | ~\new_[27552]_ );
  assign \new_[19934]_  = ~\new_[22320]_  & (~\new_[23530]_  | ~\new_[24289]_ );
  assign \new_[19935]_  = ~\new_[30757]_  & (~\new_[23521]_  | ~\new_[28218]_ );
  assign \new_[19936]_  = ~\new_[22189]_  & (~\new_[23428]_  | ~\new_[24523]_ );
  assign \new_[19937]_  = ~\new_[28718]_  & (~\new_[23613]_  | ~\new_[28091]_ );
  assign \new_[19938]_  = ~\new_[29977]_  | (~\new_[23603]_  & ~\new_[27638]_ );
  assign \new_[19939]_  = ~\new_[30774]_  | (~\new_[23474]_  & ~\new_[28479]_ );
  assign \new_[19940]_  = ~\new_[29560]_  | (~\new_[23470]_  & ~\new_[28251]_ );
  assign \new_[19941]_  = ~\new_[22207]_  & (~\new_[23596]_  | ~\new_[23131]_ );
  assign \new_[19942]_  = \new_[21720]_  & \new_[29489]_ ;
  assign \new_[19943]_  = ~\new_[30407]_  & (~\new_[23767]_  | ~\new_[28116]_ );
  assign \new_[19944]_  = ~\new_[30246]_  | (~\new_[23542]_  & ~\new_[27610]_ );
  assign \new_[19945]_  = ~\new_[29375]_  & (~\new_[23740]_  | ~\new_[29249]_ );
  assign \new_[19946]_  = ~\new_[30615]_  | (~\new_[23552]_  & ~\new_[28707]_ );
  assign \new_[19947]_  = ~\new_[29222]_  & (~\new_[23468]_  | ~\new_[27646]_ );
  assign \new_[19948]_  = \new_[21733]_  & \new_[29461]_ ;
  assign \new_[19949]_  = ~\new_[29887]_  | (~\new_[23715]_  & ~\new_[26629]_ );
  assign \new_[19950]_  = ~\new_[23608]_  & (~\new_[23551]_  | ~\new_[23630]_ );
  assign \new_[19951]_  = \new_[21836]_  & \new_[29601]_ ;
  assign \new_[19952]_  = \new_[21774]_  & \new_[29390]_ ;
  assign \new_[19953]_  = \new_[21732]_  & \new_[29344]_ ;
  assign \new_[19954]_  = ~\new_[29272]_  & (~\new_[23455]_  | ~\new_[28632]_ );
  assign \new_[19955]_  = ~\new_[30084]_  | (~\new_[23815]_  & ~\new_[27356]_ );
  assign \new_[19956]_  = ~\new_[23747]_  & (~\new_[23835]_  | ~\new_[24466]_ );
  assign \new_[19957]_  = \new_[21963]_  & \new_[29577]_ ;
  assign \new_[19958]_  = ~\new_[28236]_  & (~\new_[23588]_  | ~\new_[27578]_ );
  assign \new_[19959]_  = ~\new_[30173]_  & (~\new_[23756]_  | ~\new_[28480]_ );
  assign \new_[19960]_  = ~\new_[29139]_  | (~\new_[23523]_  & ~\new_[26575]_ );
  assign \new_[19961]_  = ~\new_[30400]_  & (~\new_[23820]_  | ~\new_[28523]_ );
  assign \new_[19962]_  = ~\new_[30707]_  | (~\new_[23803]_  & ~\new_[24662]_ );
  assign \new_[19963]_  = ~\new_[28905]_  | (~\new_[23841]_  & ~\new_[27697]_ );
  assign \new_[19964]_  = \new_[21831]_  & \new_[29474]_ ;
  assign \new_[19965]_  = ~\new_[26638]_  | ~\new_[6066]_ ;
  assign \new_[19966]_  = \new_[21657]_  & \new_[28871]_ ;
  assign \new_[19967]_  = ~\new_[30036]_  & (~\new_[23712]_  | ~\new_[29284]_ );
  assign \new_[19968]_  = \new_[21983]_  & \new_[29536]_ ;
  assign \new_[19969]_  = ~\new_[23104]_  & (~\new_[23908]_  | ~\new_[26361]_ );
  assign \new_[19970]_  = ~\new_[22996]_  & (~\new_[23916]_  | ~\new_[24640]_ );
  assign \new_[19971]_  = ~\new_[22951]_  & (~\new_[25178]_  | ~\new_[27807]_ );
  assign \new_[19972]_  = ~\new_[24400]_  & (~\new_[23911]_  | ~\new_[26377]_ );
  assign \new_[19973]_  = ~\new_[24424]_  & (~\new_[23148]_  | ~\new_[27272]_ );
  assign \new_[19974]_  = ~\new_[24044]_  & (~\new_[23890]_  | ~\new_[26406]_ );
  assign \new_[19975]_  = ~\new_[24396]_  & (~\new_[23079]_  | ~\new_[26432]_ );
  assign \new_[19976]_  = ~\new_[26471]_  & (~\new_[23922]_  | ~\new_[27002]_ );
  assign \new_[19977]_  = ~\new_[24447]_  & (~\new_[23921]_  | ~\new_[26368]_ );
  assign \new_[19978]_  = ~\new_[22473]_  & ~\new_[29736]_ ;
  assign \new_[19979]_  = ~\new_[22474]_  & ~\new_[29827]_ ;
  assign \new_[19980]_  = ~\new_[22495]_  & ~\new_[29222]_ ;
  assign \new_[19981]_  = ~\new_[22482]_  & ~\new_[28718]_ ;
  assign \new_[19982]_  = ~\new_[22514]_  & ~\new_[29272]_ ;
  assign \new_[19983]_  = ~\new_[22516]_  & ~\new_[30407]_ ;
  assign \new_[19984]_  = ~\new_[22506]_  & ~\new_[30173]_ ;
  assign \new_[19985]_  = ~\new_[22513]_  & ~\new_[29966]_ ;
  assign \new_[19986]_  = ~\new_[22507]_  & ~\new_[30162]_ ;
  assign \new_[19987]_  = ~\new_[22463]_  & ~\new_[29784]_ ;
  assign \new_[19988]_  = ~\new_[22522]_  & ~\new_[29383]_ ;
  assign \new_[19989]_  = ~\new_[22468]_  & ~\new_[30400]_ ;
  assign \new_[19990]_  = ~\new_[22521]_  & ~\new_[28236]_ ;
  assign \new_[19991]_  = ~\new_[23852]_  | ~\new_[22173]_ ;
  assign \new_[19992]_  = \new_[22605]_  & \new_[22595]_ ;
  assign \new_[19993]_  = ~\new_[22432]_  | ~\new_[24484]_ ;
  assign \new_[19994]_  = ~\new_[22182]_  | ~\new_[27608]_ ;
  assign \new_[19995]_  = \new_[22235]_  | \new_[30591]_ ;
  assign \new_[19996]_  = ~\new_[23342]_  | ~\new_[26389]_ ;
  assign \new_[19997]_  = ~\new_[23344]_  | ~\new_[22111]_ ;
  assign \new_[19998]_  = \new_[22216]_  | \new_[30597]_ ;
  assign \new_[19999]_  = ~\new_[22231]_  | ~\new_[23348]_ ;
  assign \new_[20000]_  = ~\new_[23445]_  | ~\new_[26256]_ ;
  assign \new_[20001]_  = ~\new_[22402]_  | ~\new_[28924]_ ;
  assign \new_[20002]_  = ~\new_[22385]_  | ~\new_[26822]_ ;
  assign \new_[20003]_  = ~\new_[22419]_  | ~\new_[28587]_ ;
  assign \new_[20004]_  = \new_[22121]_  & \new_[28115]_ ;
  assign \new_[20005]_  = ~\new_[30747]_  | ~\new_[5967]_ ;
  assign \new_[20006]_  = ~\new_[22378]_  | ~\new_[28532]_ ;
  assign \new_[20007]_  = \new_[22426]_  | \new_[23647]_ ;
  assign \new_[20008]_  = ~\new_[25085]_  & ~\new_[22276]_ ;
  assign \new_[20009]_  = ~\new_[22276]_  & ~\new_[29907]_ ;
  assign \new_[20010]_  = ~\new_[22155]_  | ~\new_[27564]_ ;
  assign \new_[20011]_  = ~\new_[22171]_  | ~\new_[24987]_ ;
  assign \new_[20012]_  = ~\new_[23696]_  | ~\new_[22341]_ ;
  assign \new_[20013]_  = \new_[22472]_  & \new_[24456]_ ;
  assign \new_[20014]_  = ~\new_[22321]_  | ~\new_[25023]_ ;
  assign \new_[20015]_  = ~\new_[22311]_  | ~\new_[28872]_ ;
  assign \new_[20016]_  = ~\new_[23438]_  & ~\new_[22987]_ ;
  assign \new_[20017]_  = ~\new_[25993]_  & ~\new_[22939]_ ;
  assign \new_[20018]_  = ~\new_[22138]_  | ~\new_[28722]_ ;
  assign \new_[20019]_  = ~\new_[23402]_  & ~\new_[22939]_ ;
  assign \new_[20020]_  = ~\new_[24851]_  & ~\new_[24957]_ ;
  assign \new_[20021]_  = ~\new_[23501]_  | ~\new_[21561]_ ;
  assign \new_[20022]_  = ~\new_[22287]_  | ~\new_[27613]_ ;
  assign \new_[20023]_  = ~\new_[24920]_  & ~\new_[22987]_ ;
  assign \new_[20024]_  = ~\new_[22244]_  | ~\new_[28176]_ ;
  assign \new_[20025]_  = ~\new_[22192]_  | ~\new_[26735]_ ;
  assign \new_[20026]_  = ~\new_[22159]_  | ~\new_[30057]_ ;
  assign \new_[20027]_  = ~\new_[22144]_  | ~\new_[28210]_ ;
  assign \new_[20028]_  = \new_[22119]_  | \new_[26951]_ ;
  assign \new_[20029]_  = ~\new_[22268]_  | ~\new_[23703]_ ;
  assign \new_[20030]_  = ~\new_[22195]_  | ~\new_[24891]_ ;
  assign \new_[20031]_  = \new_[22267]_  & \new_[28708]_ ;
  assign \new_[20032]_  = ~\new_[22202]_  | ~\new_[23462]_ ;
  assign \new_[20033]_  = \new_[22480]_  & \new_[24281]_ ;
  assign \new_[20034]_  = ~\new_[29699]_  | ~\new_[6076]_ ;
  assign \new_[20035]_  = \new_[22541]_  & \new_[26428]_ ;
  assign \new_[20036]_  = ~\new_[20805]_ ;
  assign \new_[20037]_  = ~\new_[26384]_  | ~\new_[24924]_ ;
  assign \new_[20038]_  = \new_[24811]_  & \new_[25100]_ ;
  assign \new_[20039]_  = ~\new_[22266]_  | ~\new_[23590]_ ;
  assign \new_[20040]_  = ~\new_[23677]_  | ~\new_[26403]_ ;
  assign \new_[20041]_  = \new_[22519]_  & \new_[23165]_ ;
  assign \new_[20042]_  = ~\new_[22484]_  | ~\new_[28508]_ ;
  assign \new_[20043]_  = \new_[22590]_  & \new_[22591]_ ;
  assign \new_[20044]_  = \new_[21615]_  & \new_[22611]_ ;
  assign \new_[20045]_  = ~\new_[20829]_ ;
  assign \new_[20046]_  = ~\new_[22123]_  | ~\new_[23507]_ ;
  assign \new_[20047]_  = ~\new_[22164]_  | ~\new_[26973]_ ;
  assign \new_[20048]_  = ~\new_[22222]_  | ~\new_[28496]_ ;
  assign \new_[20049]_  = ~\new_[22315]_  | ~\new_[23386]_ ;
  assign \new_[20050]_  = \new_[22602]_  & \new_[22643]_ ;
  assign \new_[20051]_  = \new_[22597]_  & \new_[22648]_ ;
  assign \new_[20052]_  = \new_[22235]_  | \new_[23384]_ ;
  assign \new_[20053]_  = ~\new_[25007]_  | ~\new_[26219]_ ;
  assign \new_[20054]_  = \new_[22325]_  | \new_[27679]_ ;
  assign \new_[20055]_  = \new_[22689]_  & \new_[22681]_ ;
  assign \new_[20056]_  = \new_[22663]_  & \new_[22627]_ ;
  assign \new_[20057]_  = ~\new_[22366]_  | ~\new_[25037]_ ;
  assign \new_[20058]_  = \new_[22607]_  & \new_[22659]_ ;
  assign \new_[20059]_  = \new_[22593]_  & \new_[22653]_ ;
  assign \new_[20060]_  = ~\new_[22330]_  | ~\new_[25019]_ ;
  assign \new_[20061]_  = ~\new_[23579]_  | ~\new_[26336]_ ;
  assign \new_[20062]_  = \new_[22257]_  | \new_[26575]_ ;
  assign \new_[20063]_  = \new_[22600]_  & \new_[22185]_ ;
  assign \new_[20064]_  = \new_[22503]_  & \new_[24307]_ ;
  assign \new_[20065]_  = ~\new_[22379]_  & ~\new_[29997]_ ;
  assign \new_[20066]_  = ~\new_[22174]_  | ~\new_[29268]_ ;
  assign \new_[20067]_  = ~\new_[22310]_  | ~\new_[26590]_ ;
  assign \new_[20068]_  = ~\new_[23578]_  | ~\new_[22258]_ ;
  assign \new_[20069]_  = ~\new_[23513]_  | ~\new_[22228]_ ;
  assign \new_[20070]_  = ~\new_[22299]_  | ~\new_[27621]_ ;
  assign \new_[20071]_  = ~\new_[22197]_  | ~\new_[24274]_ ;
  assign \new_[20072]_  = ~\new_[22399]_  | ~\new_[24656]_ ;
  assign \new_[20073]_  = ~\new_[22270]_  & ~\new_[29914]_ ;
  assign \new_[20074]_  = ~\new_[23597]_  | ~\new_[22333]_ ;
  assign \new_[20075]_  = \new_[22511]_  & \new_[23137]_ ;
  assign \new_[20076]_  = ~\new_[22271]_  & ~\new_[24964]_ ;
  assign \new_[20077]_  = \new_[22469]_  & \new_[23968]_ ;
  assign \new_[20078]_  = ~\new_[22107]_  | ~\new_[28887]_ ;
  assign \new_[20079]_  = ~\new_[22196]_  | ~\new_[26995]_ ;
  assign \new_[20080]_  = ~\new_[22223]_  | ~\new_[26362]_ ;
  assign \new_[20081]_  = ~\new_[22290]_  | ~\new_[23662]_ ;
  assign \new_[20082]_  = ~\new_[22211]_  | ~\new_[29104]_ ;
  assign \new_[20083]_  = ~\new_[22352]_  | ~\new_[23628]_ ;
  assign \new_[20084]_  = ~\new_[22289]_  & ~\new_[30304]_ ;
  assign \new_[20085]_  = ~\new_[22140]_  & ~\new_[30267]_ ;
  assign \new_[20086]_  = \new_[22249]_  | \new_[27860]_ ;
  assign \new_[20087]_  = \new_[22328]_  | \new_[27559]_ ;
  assign \new_[20088]_  = \new_[22426]_  | \new_[30710]_ ;
  assign \new_[20089]_  = \new_[22270]_  | \new_[23440]_ ;
  assign \new_[20090]_  = ~\new_[22407]_  | ~\new_[27641]_ ;
  assign \new_[20091]_  = ~\new_[23646]_  & ~\new_[23053]_ ;
  assign \new_[20092]_  = ~\new_[22134]_  | ~\new_[27758]_ ;
  assign \new_[20093]_  = ~\new_[22296]_  & ~\new_[24346]_ ;
  assign \new_[20094]_  = \new_[22686]_  & \new_[22635]_ ;
  assign \new_[20095]_  = ~\new_[22363]_  & ~\new_[29792]_ ;
  assign \new_[20096]_  = \new_[22493]_  & \new_[26248]_ ;
  assign \new_[20097]_  = ~\new_[22628]_  | ~\new_[28574]_ ;
  assign \new_[20098]_  = ~\new_[25977]_  & ~\new_[22379]_ ;
  assign \new_[20099]_  = \new_[22478]_  & \new_[23268]_ ;
  assign \new_[20100]_  = ~\new_[23383]_  | ~\new_[22129]_ ;
  assign \new_[20101]_  = \new_[22539]_  & \new_[23087]_ ;
  assign \new_[20102]_  = ~\new_[22430]_  | ~\new_[25056]_ ;
  assign \new_[20103]_  = ~\new_[22317]_  | ~\new_[26866]_ ;
  assign \new_[20104]_  = \new_[22140]_  | \new_[23457]_ ;
  assign \new_[20105]_  = ~\new_[22393]_  | ~\new_[29248]_ ;
  assign \new_[20106]_  = ~\new_[22123]_  | ~\new_[27620]_ ;
  assign \new_[20107]_  = ~\new_[22214]_  & ~\new_[29062]_ ;
  assign \new_[20108]_  = ~\new_[23733]_  & ~\new_[22363]_ ;
  assign \new_[20109]_  = \new_[22289]_  | \new_[23372]_ ;
  assign \new_[20110]_  = ~\new_[23610]_  | ~\new_[22360]_ ;
  assign \new_[20111]_  = ~\new_[22248]_  | ~\new_[24464]_ ;
  assign \new_[20112]_  = ~\new_[22312]_  | ~\new_[27696]_ ;
  assign \new_[20113]_  = \new_[22631]_  & \new_[22598]_ ;
  assign \new_[20114]_  = \new_[22634]_  & \new_[22601]_ ;
  assign \new_[20115]_  = \new_[22406]_  | \new_[28251]_ ;
  assign \new_[20116]_  = ~\new_[24919]_  & ~\new_[23053]_ ;
  assign \new_[20117]_  = ~\new_[22131]_  & ~\new_[29169]_ ;
  assign \new_[20118]_  = ~\new_[22124]_  & ~\new_[30660]_ ;
  assign \new_[20119]_  = ~\new_[22120]_  | ~\new_[30030]_ ;
  assign \new_[20120]_  = ~\new_[22387]_  | ~\new_[25091]_ ;
  assign \new_[20121]_  = \new_[22108]_  | \new_[26679]_ ;
  assign \new_[20122]_  = ~\new_[22365]_  | ~\new_[24656]_ ;
  assign \new_[20123]_  = \new_[22670]_  & \new_[22669]_ ;
  assign \new_[20124]_  = ~\new_[22451]_  | ~\new_[27557]_ ;
  assign \new_[20125]_  = ~\new_[22422]_  | ~\new_[28606]_ ;
  assign \new_[20126]_  = ~\new_[22169]_  | ~\new_[26201]_ ;
  assign \new_[20127]_  = ~\new_[25105]_  & ~\new_[23045]_ ;
  assign \new_[20128]_  = \new_[22678]_  & \new_[22606]_ ;
  assign \new_[20129]_  = ~\new_[22109]_  | ~\new_[26389]_ ;
  assign \new_[20130]_  = \new_[22687]_  & \new_[22688]_ ;
  assign \new_[20131]_  = ~\new_[25149]_  & ~\new_[23453]_ ;
  assign \new_[20132]_  = ~\new_[22380]_  | ~\new_[23727]_ ;
  assign \new_[20133]_  = \new_[22512]_  & \new_[23166]_ ;
  assign \new_[20134]_  = ~\new_[22415]_  | ~\new_[28477]_ ;
  assign \new_[20135]_  = ~\new_[22339]_  | ~\new_[28086]_ ;
  assign \new_[20136]_  = ~\new_[22347]_  | ~\new_[27644]_ ;
  assign \new_[20137]_  = \new_[22535]_  & \new_[24541]_ ;
  assign \new_[20138]_  = ~\new_[24966]_  & ~\new_[23045]_ ;
  assign \new_[20139]_  = ~\new_[22429]_  | ~\new_[22239]_ ;
  assign \new_[20140]_  = \new_[22538]_  & \new_[24544]_ ;
  assign \new_[20141]_  = ~\new_[22198]_  | ~\new_[28346]_ ;
  assign \new_[20142]_  = \new_[22216]_  | \new_[23873]_ ;
  assign \new_[20143]_  = ~\new_[22447]_  | ~\new_[28097]_ ;
  assign \new_[20144]_  = \new_[22544]_  & \new_[24751]_ ;
  assign \new_[20145]_  = ~\new_[22187]_  & ~\new_[30268]_ ;
  assign \new_[20146]_  = ~\new_[22188]_  & ~\new_[24885]_ ;
  assign \new_[20147]_  = \new_[22187]_  | \new_[23465]_ ;
  assign \new_[20148]_  = ~\new_[22284]_  | ~\new_[27632]_ ;
  assign \new_[20149]_  = ~\new_[22452]_  | ~\new_[28420]_ ;
  assign \new_[20150]_  = ~\new_[22294]_  | ~\new_[23086]_ ;
  assign \new_[20151]_  = ~\new_[22458]_  | ~\new_[28193]_ ;
  assign \new_[20152]_  = \new_[22545]_  & \new_[24709]_ ;
  assign \new_[20153]_  = ~\new_[21005]_ ;
  assign \new_[20154]_  = ~\new_[23208]_  | ~\new_[23146]_  | ~\new_[27761]_ ;
  assign \new_[20155]_  = ~\new_[23992]_  | ~\new_[26924]_  | ~\new_[27808]_ ;
  assign \new_[20156]_  = ~\new_[24294]_  | ~\new_[24467]_  | ~\new_[27678]_ ;
  assign \new_[20157]_  = ~\new_[24262]_  | ~\new_[24043]_  | ~\new_[27651]_ ;
  assign \new_[20158]_  = ~\new_[29881]_  | ~\new_[27311]_  | ~\new_[24344]_ ;
  assign \new_[20159]_  = ~\new_[30282]_  | ~\new_[28470]_  | ~\new_[24272]_ ;
  assign \new_[20160]_  = \new_[22166]_  | \new_[28576]_ ;
  assign \new_[20161]_  = ~\new_[24429]_  | ~\new_[24367]_  | ~\new_[26709]_ ;
  assign \new_[20162]_  = ~\new_[23141]_  | ~\new_[24386]_  | ~\new_[27656]_ ;
  assign \new_[20163]_  = \new_[22442]_  | \new_[24362]_ ;
  assign \new_[20164]_  = \new_[22417]_  | \new_[24343]_ ;
  assign \new_[20165]_  = ~\new_[24422]_  | ~\new_[27782]_  | ~\new_[27757]_ ;
  assign \new_[20166]_  = \new_[22428]_  | \new_[27663]_ ;
  assign \new_[20167]_  = \new_[22306]_  | \new_[24359]_ ;
  assign \new_[20168]_  = ~\new_[29941]_  | ~\new_[27281]_  | ~\new_[23254]_ ;
  assign \new_[20169]_  = ~\new_[23139]_  | ~\new_[26726]_  | ~\new_[27004]_ ;
  assign \new_[20170]_  = ~\new_[30029]_  & (~\new_[24358]_  | ~\new_[29528]_ );
  assign \new_[20171]_  = ~\new_[21015]_ ;
  assign \new_[20172]_  = ~\new_[30317]_  | ~\new_[27441]_  | ~\new_[24287]_ ;
  assign \new_[20173]_  = \new_[22217]_  | \new_[26999]_ ;
  assign \new_[20174]_  = ~\new_[30102]_  | ~\new_[27529]_  | ~\new_[24313]_ ;
  assign \new_[20175]_  = ~\new_[24395]_  | ~\new_[26334]_  | ~\new_[28528]_ ;
  assign \new_[20176]_  = ~\new_[21019]_ ;
  assign n8549 = m6_s14_cyc_o_reg;
  assign \new_[20178]_  = ~\new_[24054]_  | ~\new_[27407]_  | ~\new_[26838]_ ;
  assign \new_[20179]_  = ~\new_[23099]_  | ~\new_[27241]_  | ~\new_[27560]_ ;
  assign \new_[20180]_  = ~\new_[29590]_  | ~\new_[26178]_  | ~\new_[26297]_ ;
  assign \new_[20181]_  = \new_[22386]_  | \new_[27634]_ ;
  assign \new_[20182]_  = ~\new_[24420]_  | ~\new_[24510]_  | ~\new_[27699]_ ;
  assign \new_[20183]_  = ~\new_[23439]_  | ~\new_[27909]_  | ~\new_[27655]_ ;
  assign n8524 = m7_s6_cyc_o_reg;
  assign \new_[20185]_  = ~\new_[29924]_  | ~\new_[28352]_  | ~\new_[24319]_ ;
  assign n7724 = ~\new_[29328]_  | ~\new_[22518]_ ;
  assign n7714 = ~\new_[28923]_  | ~\new_[22525]_ ;
  assign n8659 = m6_s8_cyc_o_reg;
  assign n8819 = m6_s9_cyc_o_reg;
  assign n7719 = ~\new_[29644]_  | ~\new_[22528]_ ;
  assign \new_[20191]_  = ~\new_[24201]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign n8744 = m6_s5_cyc_o_reg;
  assign n7744 = ~\new_[29275]_  | ~\new_[22529]_ ;
  assign n8869 = m5_s4_cyc_o_reg;
  assign n7739 = ~\new_[29698]_  | ~\new_[22530]_ ;
  assign n7734 = ~\new_[29109]_  | ~\new_[22531]_ ;
  assign n8719 = m6_s13_cyc_o_reg;
  assign n7729 = ~\new_[29687]_  | ~\new_[22517]_ ;
  assign \new_[20199]_  = ~\new_[30183]_  | ~\new_[27521]_  | ~\new_[24421]_ ;
  assign \new_[20200]_  = ~\new_[30054]_  | ~\new_[27494]_  | ~\new_[24520]_ ;
  assign \new_[20201]_  = \new_[22436]_  | \new_[23512]_ ;
  assign \new_[20202]_  = ~\new_[30299]_  | ~\new_[27496]_  | ~\new_[24312]_ ;
  assign \new_[20203]_  = ~\new_[21054]_ ;
  assign \new_[20204]_  = ~\new_[24361]_  | ~\new_[27550]_  | ~\new_[27652]_ ;
  assign \new_[20205]_  = ~\new_[22176]_  | ~\new_[28836]_ ;
  assign n8364 = m5_s6_cyc_o_reg;
  assign \new_[20207]_  = ~\new_[23064]_  | (~\new_[25767]_  & ~\new_[29784]_ );
  assign \new_[20208]_  = ~\new_[22113]_  | ~\new_[29028]_ ;
  assign \new_[20209]_  = ~\new_[22397]_  | ~\new_[29028]_ ;
  assign \new_[20210]_  = ~\new_[22125]_  | ~\new_[30599]_ ;
  assign \new_[20211]_  = \new_[22127]_  & \new_[26281]_ ;
  assign \new_[20212]_  = ~\new_[22403]_  | ~\new_[29151]_ ;
  assign \new_[20213]_  = \new_[22283]_  & \new_[26305]_ ;
  assign \new_[20214]_  = ~\new_[22148]_  | ~\new_[28918]_ ;
  assign \new_[20215]_  = ~\new_[23127]_  | (~\new_[24513]_  & ~\new_[30289]_ );
  assign \new_[20216]_  = ~\new_[24348]_  | (~\new_[24383]_  & ~\new_[30438]_ );
  assign \new_[20217]_  = ~\new_[22899]_  | (~\new_[26121]_  & ~\new_[29827]_ );
  assign \new_[20218]_  = ~\new_[22285]_  | ~\new_[28836]_ ;
  assign \new_[20219]_  = ~\new_[22445]_  & ~\new_[26187]_ ;
  assign \new_[20220]_  = ~\new_[22278]_  | ~\new_[29276]_ ;
  assign \new_[20221]_  = ~\new_[22236]_  | ~\new_[29020]_ ;
  assign \new_[20222]_  = ~\new_[22326]_  | ~\new_[29623]_ ;
  assign \new_[20223]_  = ~\new_[30467]_  | (~\new_[24218]_  & ~\new_[28745]_ );
  assign \new_[20224]_  = ~\new_[24443]_  | (~\new_[23142]_  & ~\new_[30014]_ );
  assign n8479 = m4_s9_cyc_o_reg;
  assign \new_[20226]_  = ~\new_[22272]_  & ~\new_[26568]_ ;
  assign \new_[20227]_  = ~\new_[22137]_  | (~\new_[26330]_  & ~\new_[29222]_ );
  assign \new_[20228]_  = ~\new_[22118]_  | ~\new_[29276]_ ;
  assign \new_[20229]_  = ~\new_[22377]_  | ~\new_[28675]_ ;
  assign \new_[20230]_  = ~\new_[22336]_  | ~\new_[29410]_ ;
  assign \new_[20231]_  = \new_[22373]_  & \new_[26320]_ ;
  assign \new_[20232]_  = \new_[22277]_  & \new_[26410]_ ;
  assign \new_[20233]_  = ~\new_[30566]_  | ~\new_[6034]_ ;
  assign \new_[20234]_  = ~\new_[22298]_  | ~\new_[28595]_ ;
  assign \new_[20235]_  = \new_[22359]_  & \new_[24340]_ ;
  assign \new_[20236]_  = ~\new_[22250]_  & ~\new_[26208]_ ;
  assign \new_[20237]_  = ~\new_[22303]_  | ~\new_[29868]_ ;
  assign \new_[20238]_  = ~\new_[22368]_  | ~\new_[28278]_ ;
  assign \new_[20239]_  = ~\new_[22158]_  & ~\new_[26195]_ ;
  assign \new_[20240]_  = ~\new_[22934]_  | (~\new_[26315]_  & ~\new_[29272]_ );
  assign \new_[20241]_  = ~\new_[22136]_  | ~\new_[29623]_ ;
  assign \new_[20242]_  = ~\new_[24417]_  | (~\new_[24407]_  & ~\new_[30162]_ );
  assign \new_[20243]_  = ~\new_[22281]_  | ~\new_[29410]_ ;
  assign \new_[20244]_  = ~\new_[22300]_  | ~\new_[30693]_ ;
  assign \new_[20245]_  = ~\new_[23088]_  | (~\new_[24039]_  & ~\new_[30425]_ );
  assign \new_[20246]_  = ~\new_[22175]_  | (~\new_[24564]_  & ~\new_[28236]_ );
  assign \new_[20247]_  = ~\new_[22163]_  | ~\new_[29583]_ ;
  assign \new_[20248]_  = ~\new_[22346]_  | ~\new_[30198]_ ;
  assign \new_[20249]_  = ~\new_[22351]_  | ~\new_[28894]_ ;
  assign \new_[20250]_  = \new_[22435]_  & \new_[26538]_ ;
  assign \new_[20251]_  = ~\new_[22980]_  | (~\new_[26287]_  & ~\new_[30240]_ );
  assign \new_[20252]_  = ~\new_[23937]_  | (~\new_[24389]_  & ~\new_[30757]_ );
  assign \new_[20253]_  = ~\new_[22978]_  & (~\new_[29442]_  | ~\new_[27883]_ );
  assign \new_[20254]_  = ~\new_[22389]_  | ~\new_[29808]_ ;
  assign \new_[20255]_  = \new_[22390]_  & \new_[24612]_ ;
  assign \new_[20256]_  = ~\new_[22391]_  | ~\new_[30015]_ ;
  assign \new_[20257]_  = ~\new_[22152]_  | ~\new_[29421]_ ;
  assign \new_[20258]_  = \new_[22322]_  & \new_[26420]_ ;
  assign \new_[20259]_  = ~\new_[22401]_  | ~\new_[29151]_ ;
  assign \new_[20260]_  = ~\new_[26400]_  | (~\new_[26432]_  & ~\new_[29383]_ );
  assign n8454 = m4_s13_cyc_o_reg;
  assign \new_[20262]_  = ~\new_[22357]_  | ~\new_[28675]_ ;
  assign \new_[20263]_  = ~\new_[24437]_  | (~\new_[27611]_  & ~\new_[29367]_ );
  assign n8749 = m4_s14_cyc_o_reg;
  assign \new_[20265]_  = ~\new_[30574]_  | ~\new_[6273]_  | ~\new_[30599]_  | ~\new_[24153]_ ;
  assign \new_[20266]_  = ~\new_[30125]_  | ~\new_[6189]_  | ~\new_[28278]_  | ~\new_[26215]_ ;
  assign \new_[20267]_  = ~\new_[30750]_  | ~\new_[31143]_  | ~\new_[30222]_  | ~\new_[23140]_ ;
  assign \new_[20268]_  = ~\new_[30538]_  | ~\new_[6214]_  | ~\new_[30693]_  | ~\new_[24402]_ ;
  assign \new_[20269]_  = ~\new_[30573]_  | ~\new_[6199]_  | ~\new_[30640]_  | ~\new_[24401]_ ;
  assign \new_[20270]_  = ~\new_[29692]_  | ~\new_[6047]_  | ~\new_[28836]_  | ~\new_[24310]_ ;
  assign \new_[20271]_  = ~\new_[30775]_  | ~\new_[6073]_  | ~\new_[30494]_  | ~\new_[24416]_ ;
  assign \new_[20272]_  = ~\new_[30774]_  | ~\new_[6053]_  | ~\new_[30242]_  | ~\new_[24184]_ ;
  assign \new_[20273]_  = ~\new_[30434]_  | ~\new_[31406]_  | ~\new_[30467]_  | ~\new_[24406]_ ;
  assign \new_[20274]_  = ~\new_[30507]_  | ~\new_[6183]_  | ~\new_[29808]_  | ~\new_[23186]_ ;
  assign \new_[20275]_  = ~\new_[29233]_  | ~\new_[31235]_  | ~\new_[29868]_  | ~\new_[24455]_ ;
  assign \new_[20276]_  = ~\new_[29887]_  | ~\new_[6068]_  | ~\new_[29410]_  | ~\new_[24257]_ ;
  assign \new_[20277]_  = ~\new_[30615]_  | ~\new_[6195]_  | ~\new_[30198]_  | ~\new_[24398]_ ;
  assign \new_[20278]_  = ~\new_[29560]_  | ~\new_[6003]_  | ~\new_[29421]_  | ~\new_[24442]_ ;
  assign \new_[20279]_  = ~\new_[30555]_  | ~\new_[6208]_  | ~\new_[30686]_  | ~\new_[24487]_ ;
  assign \new_[20280]_  = ~\new_[30789]_  | ~\new_[6082]_  | ~\new_[30248]_  | ~\new_[24478]_ ;
  assign \new_[20281]_  = ~\new_[30707]_  | ~\new_[6086]_  | ~\new_[30297]_  | ~\new_[24255]_ ;
  assign \new_[20282]_  = ~\new_[30725]_  | ~\new_[6186]_  | ~\new_[30571]_  | ~\new_[24498]_ ;
  assign n8579 = m3_s9_cyc_o_reg;
  assign n8919 = m3_s8_cyc_o_reg;
  assign \new_[20285]_  = ~\new_[31394]_  | ~\new_[28014]_  | ~\new_[29169]_ ;
  assign \new_[20286]_  = ~\new_[21128]_ ;
  assign \new_[20287]_  = ~\new_[5895]_  | ~\new_[28265]_  | ~\new_[29855]_ ;
  assign \new_[20288]_  = \new_[29924]_  & \new_[28113]_ ;
  assign \new_[20289]_  = \new_[26262]_  & \new_[30097]_ ;
  assign n8409 = m3_s10_cyc_o_reg;
  assign n8834 = m2_s6_cyc_o_reg;
  assign n8614 = m2_s9_cyc_o_reg;
  assign n8879 = m1_s6_cyc_o_reg;
  assign \new_[20294]_  = ~\new_[5896]_  | ~\new_[28209]_  | ~\new_[29100]_ ;
  assign \new_[20295]_  = \new_[30317]_  & \new_[26824]_ ;
  assign \new_[20296]_  = \new_[30102]_  & \new_[28422]_ ;
  assign \new_[20297]_  = \new_[26358]_  & \new_[30159]_ ;
  assign \new_[20298]_  = ~\new_[6044]_  | ~\new_[28971]_  | ~\new_[29736]_ ;
  assign n8494 = m0_s8_cyc_o_reg;
  assign n8874 = m1_s5_cyc_o_reg;
  assign \new_[20301]_  = ~\new_[26427]_  & ~\new_[30710]_ ;
  assign \new_[20302]_  = \new_[30299]_  & \new_[26203]_ ;
  assign \new_[20303]_  = ~\new_[31143]_  | ~\new_[30182]_  | ~\new_[30289]_ ;
  assign \new_[20304]_  = ~\new_[5897]_  | ~\new_[28688]_  | ~\new_[30389]_ ;
  assign n8514 = m0_s9_cyc_o_reg;
  assign \new_[20306]_  = \new_[30282]_  & \new_[28815]_ ;
  assign n8779 = m1_s12_cyc_o_reg;
  assign n8519 = m1_s10_cyc_o_reg;
  assign \new_[20309]_  = ~\new_[21559]_ ;
  assign \new_[20310]_  = ~\new_[6047]_  | ~\new_[28629]_  | ~\new_[29827]_ ;
  assign \new_[20311]_  = ~\new_[23046]_  & ~\new_[30075]_ ;
  assign \new_[20312]_  = ~\new_[6049]_  | ~\new_[27852]_  | ~\new_[30616]_ ;
  assign n8729 = m0_s3_cyc_o_reg;
  assign \new_[20314]_  = ~\new_[5905]_  | ~\new_[27992]_  | ~\new_[29565]_ ;
  assign n8784 = m0_s5_cyc_o_reg;
  assign \new_[20316]_  = ~\new_[31232]_  | ~\new_[26549]_  | ~\new_[30355]_ ;
  assign \new_[20317]_  = \new_[26342]_  & \new_[30172]_ ;
  assign n8684 = m0_s12_cyc_o_reg;
  assign \new_[20319]_  = ~\new_[5906]_  | ~\new_[28148]_  | ~\new_[29898]_ ;
  assign n8929 = m0_s11_cyc_o_reg;
  assign n8559 = m0_s10_cyc_o_reg;
  assign n8814 = m7_s3_cyc_o_reg;
  assign \new_[20323]_  = ~\new_[31410]_  | ~\new_[27593]_  | ~\new_[29064]_ ;
  assign \new_[20324]_  = ~\new_[6058]_  | ~\new_[29362]_  | ~\new_[30407]_ ;
  assign \new_[20325]_  = ~\new_[30186]_  & ~\new_[22909]_ ;
  assign \new_[20326]_  = ~\new_[31429]_  | ~\new_[26549]_  | ~\new_[30355]_ ;
  assign \new_[20327]_  = ~\new_[6211]_  | ~\new_[28100]_  | ~\new_[30028]_ ;
  assign \new_[20328]_  = ~\new_[28893]_  & ~\new_[22905]_ ;
  assign \new_[20329]_  = \new_[26392]_  & \new_[30092]_ ;
  assign \new_[20330]_  = ~\new_[21198]_ ;
  assign \new_[20331]_  = ~\new_[6068]_  | ~\new_[29348]_  | ~\new_[30173]_ ;
  assign \new_[20332]_  = ~\new_[6213]_  | ~\new_[29160]_  | ~\new_[30014]_ ;
  assign \new_[20333]_  = ~\new_[6086]_  | ~\new_[28970]_  | ~\new_[30036]_ ;
  assign \new_[20334]_  = ~\new_[22961]_  | ~\new_[30337]_ ;
  assign \new_[20335]_  = ~\new_[5830]_  | ~\new_[28840]_  | ~\new_[29150]_ ;
  assign \new_[20336]_  = \new_[29941]_  & \new_[25800]_ ;
  assign \new_[20337]_  = \new_[26515]_  & \new_[30320]_ ;
  assign \new_[20338]_  = ~\new_[31406]_  | ~\new_[26484]_  | ~\new_[30224]_ ;
  assign \new_[20339]_  = ~\new_[21204]_ ;
  assign \new_[20340]_  = ~\new_[6073]_  | ~\new_[29073]_  | ~\new_[30656]_ ;
  assign \new_[20341]_  = ~\new_[6189]_  | ~\new_[27999]_  | ~\new_[30240]_ ;
  assign \new_[20342]_  = ~\new_[31438]_  | ~\new_[27894]_  | ~\new_[28846]_ ;
  assign \new_[20343]_  = \new_[29881]_  & \new_[28797]_ ;
  assign \new_[20344]_  = \new_[26430]_  & \new_[29863]_ ;
  assign \new_[20345]_  = ~\new_[5904]_  | ~\new_[28106]_  | ~\new_[29648]_ ;
  assign \new_[20346]_  = ~\new_[6273]_  | ~\new_[29110]_  | ~\new_[30342]_ ;
  assign \new_[20347]_  = \new_[24785]_  & \new_[30061]_ ;
  assign \new_[20348]_  = ~\new_[21343]_ ;
  assign \new_[20349]_  = \new_[26261]_  & \new_[29888]_ ;
  assign \new_[20350]_  = ~\new_[31499]_  | ~\new_[28058]_  | ~\new_[30557]_ ;
  assign \new_[20351]_  = \new_[26337]_  & \new_[29762]_ ;
  assign \new_[20352]_  = ~\new_[21238]_ ;
  assign \new_[20353]_  = ~\new_[21241]_ ;
  assign \new_[20354]_  = ~\new_[6082]_  | ~\new_[29353]_  | ~\new_[30244]_ ;
  assign \new_[20355]_  = ~\new_[21049]_ ;
  assign \new_[20356]_  = \new_[30183]_  & \new_[24965]_ ;
  assign \new_[20357]_  = ~\new_[21250]_ ;
  assign \new_[20358]_  = ~\new_[21251]_ ;
  assign \new_[20359]_  = \new_[29873]_  & \new_[24756]_ ;
  assign \new_[20360]_  = ~\new_[6093]_  | ~\new_[26259]_  | ~\new_[30607]_ ;
  assign \new_[20361]_  = ~\new_[6006]_  | ~\new_[26759]_  | ~\new_[29383]_ ;
  assign \new_[20362]_  = ~\new_[6214]_  | ~\new_[29538]_  | ~\new_[30273]_ ;
  assign \new_[20363]_  = \new_[30054]_  & \new_[26349]_ ;
  assign \new_[20364]_  = ~\new_[5931]_  | ~\new_[29433]_  | ~\new_[29672]_ ;
  assign \new_[20365]_  = ~\new_[6206]_  | ~\new_[28202]_  | ~\new_[29360]_ ;
  assign \new_[20366]_  = ~\new_[6038]_  | ~\new_[28670]_  | ~\new_[29826]_ ;
  assign \new_[20367]_  = ~\new_[30511]_  | ~\new_[29642]_  | ~\new_[29019]_ ;
  assign \new_[20368]_  = ~\new_[6031]_  | ~\new_[29925]_  | ~\new_[29122]_ ;
  assign \new_[20369]_  = ~\new_[31429]_  | ~\new_[26493]_  | ~\new_[30044]_ ;
  assign \new_[20370]_  = \new_[22916]_  | \new_[28754]_ ;
  assign \new_[20371]_  = ~\new_[31648]_  | ~\new_[28721]_  | ~\new_[29629]_ ;
  assign \new_[20372]_  = ~\new_[5978]_  | ~\new_[26524]_  | ~\new_[28979]_ ;
  assign \new_[20373]_  = ~\new_[6056]_  | ~\new_[28281]_  | ~\new_[29445]_ ;
  assign \new_[20374]_  = \new_[22879]_  | \new_[28303]_ ;
  assign \new_[20375]_  = ~\new_[6062]_  | ~\new_[28739]_  | ~\new_[29174]_ ;
  assign \new_[20376]_  = ~\new_[5968]_  | ~\new_[29488]_  | ~\new_[29501]_ ;
  assign \new_[20377]_  = ~\new_[31232]_  | ~\new_[27920]_  | ~\new_[29062]_ ;
  assign \new_[20378]_  = \new_[22958]_  | \new_[30238]_ ;
  assign \new_[20379]_  = ~\new_[5983]_  | ~\new_[28739]_  | ~\new_[29174]_ ;
  assign \new_[20380]_  = ~\new_[31648]_  | ~\new_[26620]_  | ~\new_[29745]_ ;
  assign \new_[20381]_  = ~\new_[5991]_  | ~\new_[28702]_  | ~\new_[28873]_ ;
  assign \new_[20382]_  = ~\new_[6087]_  | ~\new_[28721]_  | ~\new_[29629]_ ;
  assign \new_[20383]_  = ~\new_[29790]_  | ~\new_[6192]_ ;
  assign \new_[20384]_  = ~\new_[28609]_  | ~\new_[5987]_ ;
  assign \new_[20385]_  = \new_[22968]_  | \new_[28443]_ ;
  assign \new_[20386]_  = ~\new_[31394]_  | ~\new_[28730]_  | ~\new_[30331]_ ;
  assign \new_[20387]_  = ~\new_[31763]_  | ~\new_[28912]_  | ~\new_[29564]_ ;
  assign \new_[20388]_  = ~\new_[6091]_  | ~\new_[28912]_  | ~\new_[29564]_ ;
  assign \new_[20389]_  = \new_[22954]_  | \new_[28677]_ ;
  assign \new_[20390]_  = ~\new_[31491]_  | ~\new_[27928]_  | ~\new_[30340]_ ;
  assign \new_[20391]_  = ~\new_[5978]_  | ~\new_[28281]_  | ~\new_[29445]_ ;
  assign \new_[20392]_  = ~\new_[6007]_  | ~\new_[28760]_  | ~\new_[29956]_ ;
  assign \new_[20393]_  = ~\new_[6094]_  | ~\new_[28379]_  | ~\new_[29748]_ ;
  assign \new_[20394]_  = ~\new_[22400]_  & (~\new_[29384]_  | ~\new_[29583]_ );
  assign \new_[20395]_  = ~\new_[22856]_  & (~\new_[28658]_  | ~\new_[29028]_ );
  assign \new_[20396]_  = ~\new_[22220]_  & (~\new_[28678]_  | ~\new_[28836]_ );
  assign \new_[20397]_  = ~\new_[21569]_  & (~\new_[26627]_  | ~\new_[28918]_ );
  assign \new_[20398]_  = ~\new_[22920]_  & (~\new_[28021]_  | ~\new_[29020]_ );
  assign \new_[20399]_  = ~\new_[22900]_  & (~\new_[28027]_  | ~\new_[29623]_ );
  assign \new_[20400]_  = ~\new_[22286]_  & (~\new_[26651]_  | ~\new_[29276]_ );
  assign \new_[20401]_  = ~\new_[22633]_  & (~\new_[28166]_  | ~\new_[29410]_ );
  assign \new_[20402]_  = ~\new_[23040]_  & (~\new_[29359]_  | ~\new_[30297]_ );
  assign \new_[20403]_  = ~\new_[22652]_  & (~\new_[27427]_  | ~\new_[28894]_ );
  assign \new_[20404]_  = ~\new_[23076]_  & (~\new_[29371]_  | ~\new_[28818]_ );
  assign \new_[20405]_  = ~\new_[22875]_  & (~\new_[30696]_  | ~\new_[30653]_ );
  assign \new_[20406]_  = ~\new_[22921]_  & (~\new_[28998]_  | ~\new_[29421]_ );
  assign \new_[20407]_  = ~\new_[23074]_  & (~\new_[30769]_  | ~\new_[30640]_ );
  assign \new_[20408]_  = ~\new_[22847]_  & (~\new_[28191]_  | ~\new_[29151]_ );
  assign \new_[20409]_  = ~\new_[29375]_  | ~\new_[6060]_ ;
  assign \new_[20410]_  = ~\new_[30328]_  | ~\new_[5980]_ ;
  assign \new_[20411]_  = ~\new_[26660]_  | ~\new_[5981]_ ;
  assign \new_[20412]_  = ~\new_[30121]_  | ~\new_[5993]_ ;
  assign \new_[20413]_  = ~\new_[29113]_  | ~\new_[6268]_ ;
  assign \new_[20414]_  = ~\new_[30059]_  | ~\new_[5993]_ ;
  assign \new_[20415]_  = ~\new_[28819]_  | ~\new_[5922]_ ;
  assign \new_[20416]_  = ~\new_[28909]_  | ~\new_[31033]_ ;
  assign \new_[20417]_  = ~\new_[29595]_  | ~\new_[5988]_ ;
  assign \new_[20418]_  = ~\new_[30002]_  | ~\new_[6065]_ ;
  assign \new_[20419]_  = ~\new_[29544]_  | ~\new_[6052]_ ;
  assign \new_[20420]_  = ~\new_[28020]_  | ~\new_[6063]_ ;
  assign \new_[20421]_  = ~\new_[29222]_  | ~\new_[5982]_ ;
  assign \new_[20422]_  = ~\new_[28020]_  | ~\new_[5982]_ ;
  assign \new_[20423]_  = ~\new_[29926]_  | ~\new_[6048]_ ;
  assign \new_[20424]_  = ~\new_[28609]_  | ~\new_[6213]_ ;
  assign \new_[20425]_  = ~\new_[26660]_  | ~\new_[5982]_ ;
  assign \new_[20426]_  = ~\new_[28362]_  | ~\new_[6044]_ ;
  assign \new_[20427]_  = ~\new_[28362]_  | ~\new_[5969]_ ;
  assign \new_[20428]_  = ~\new_[28884]_  | ~\new_[5929]_ ;
  assign \new_[20429]_  = ~\new_[29828]_  | ~\new_[31121]_ ;
  assign \new_[20430]_  = ~\new_[28909]_  | ~\new_[31235]_ ;
  assign \new_[20431]_  = ~\new_[29595]_  | ~\new_[5920]_ ;
  assign \new_[20432]_  = ~\new_[28857]_  | ~\new_[5920]_ ;
  assign \new_[20433]_  = ~\new_[28331]_  | ~\new_[5966]_ ;
  assign \new_[20434]_  = ~\new_[28884]_  | ~\new_[6086]_ ;
  assign \new_[20435]_  = ~\new_[30059]_  | ~\new_[6077]_ ;
  assign \new_[20436]_  = ~\new_[29113]_  | ~\new_[5996]_ ;
  assign \new_[20437]_  = ~\new_[30072]_  | ~\new_[6005]_ ;
  assign \new_[20438]_  = ~\new_[26660]_  | ~\new_[6063]_ ;
  assign \new_[20439]_  = ~\new_[28236]_  | ~\new_[6088]_ ;
  assign \new_[20440]_  = ~\new_[29992]_  | ~\new_[5963]_ ;
  assign \new_[20441]_  = ~\new_[29968]_  | ~\new_[5998]_ ;
  assign \new_[20442]_  = ~\new_[30162]_  | ~\new_[5995]_ ;
  assign \new_[20443]_  = ~\new_[29113]_  | ~\new_[5995]_ ;
  assign \new_[20444]_  = ~\new_[30276]_  | ~\new_[6217]_ ;
  assign \new_[20445]_  = ~\new_[29452]_  | ~\new_[6197]_ ;
  assign \new_[20446]_  = \new_[30163]_  & \new_[29202]_ ;
  assign \new_[20447]_  = ~\new_[30076]_  | ~\new_[5905]_ ;
  assign \new_[20448]_  = ~\new_[30070]_  | ~\new_[6196]_ ;
  assign \new_[20449]_  = \new_[29943]_  & \new_[28962]_ ;
  assign \new_[20450]_  = ~\new_[29935]_  | ~\new_[31712]_ ;
  assign \new_[20451]_  = ~\new_[29598]_  | ~\new_[31422]_ ;
  assign \new_[20452]_  = ~\new_[30003]_  | ~\new_[6092]_ ;
  assign \new_[20453]_  = ~\new_[30208]_  & ~\new_[30305]_ ;
  assign \new_[20454]_  = \new_[30312]_  & \new_[28883]_ ;
  assign \new_[20455]_  = ~\new_[29077]_  | ~\new_[31400]_ ;
  assign \new_[20456]_  = ~\new_[30003]_  | ~\new_[6093]_ ;
  assign \new_[20457]_  = \new_[30006]_  & \new_[28939]_ ;
  assign \new_[20458]_  = \new_[30019]_  & \new_[29357]_ ;
  assign \new_[20459]_  = ~\new_[29767]_  | ~\new_[6193]_ ;
  assign \new_[20460]_  = ~\new_[29935]_  | ~\new_[6050]_ ;
  assign \new_[20461]_  = ~\new_[29994]_  & ~\new_[30087]_ ;
  assign \new_[20462]_  = ~\new_[30219]_  | ~\new_[5900]_ ;
  assign \new_[20463]_  = ~\new_[29989]_  | ~\new_[6076]_ ;
  assign \new_[20464]_  = ~\new_[28204]_  | ~\new_[6076]_ ;
  assign \new_[20465]_  = ~\new_[30003]_  | ~\new_[6216]_ ;
  assign \new_[20466]_  = ~\new_[29699]_  | ~\new_[5925]_ ;
  assign \new_[20467]_  = ~\new_[29055]_  | ~\new_[6040]_ ;
  assign \new_[20468]_  = ~\new_[29699]_  | ~\new_[5924]_ ;
  assign \new_[20469]_  = ~\new_[29598]_  | ~\new_[31438]_ ;
  assign \new_[20470]_  = ~\new_[29238]_  | ~\new_[6073]_ ;
  assign \new_[20471]_  = ~\new_[26842]_  | ~\new_[6096]_ ;
  assign \new_[20472]_  = ~\new_[30350]_  | ~\new_[5984]_ ;
  assign \new_[20473]_  = ~\new_[26842]_  & ~\new_[6199]_ ;
  assign \new_[20474]_  = ~\new_[29772]_  & ~\new_[30339]_ ;
  assign \new_[20475]_  = ~\new_[30305]_  | ~\new_[5908]_ ;
  assign \new_[20476]_  = ~\new_[30663]_  | ~\new_[5910]_ ;
  assign \new_[20477]_  = ~\new_[29238]_  | ~\new_[5989]_ ;
  assign \new_[20478]_  = ~\new_[29935]_  | ~\new_[6049]_ ;
  assign \new_[20479]_  = ~\new_[28944]_  | ~\new_[31438]_ ;
  assign \new_[20480]_  = ~\new_[28204]_  | ~\new_[5925]_ ;
  assign \new_[20481]_  = ~\new_[29611]_  | ~\new_[6186]_ ;
  assign \new_[20482]_  = ~\new_[28944]_  | ~\new_[31440]_ ;
  assign \new_[20483]_  = ~\new_[30087]_  | ~\new_[5901]_ ;
  assign \new_[20484]_  = ~\new_[30070]_  | ~\new_[6057]_ ;
  assign \new_[20485]_  = ~\new_[29181]_  | ~\new_[31423]_ ;
  assign \new_[20486]_  = ~\new_[30339]_  | ~\new_[5907]_ ;
  assign \new_[20487]_  = ~\new_[30684]_  | ~\new_[6070]_ ;
  assign \new_[20488]_  = ~\new_[29611]_  | ~\new_[5928]_ ;
  assign \new_[20489]_  = ~\new_[30269]_  | ~\new_[29927]_ ;
  assign \new_[20490]_  = ~\new_[26638]_  & ~\new_[6194]_ ;
  assign \new_[20491]_  = ~\new_[30637]_  | ~\new_[5925]_ ;
  assign \new_[20492]_  = ~\new_[30350]_  | ~\new_[6194]_ ;
  assign \new_[20493]_  = ~\new_[30350]_  | ~\new_[31157]_ ;
  assign \new_[20494]_  = ~\new_[29989]_  | ~\new_[5924]_ ;
  assign \new_[20495]_  = ~\new_[30688]_  | ~\new_[6057]_ ;
  assign \new_[20496]_  = ~\new_[30130]_  | ~\new_[31423]_ ;
  assign \new_[20497]_  = ~\new_[29611]_  | ~\new_[6084]_ ;
  assign \new_[20498]_  = ~\new_[29238]_  | ~\new_[6072]_ ;
  assign \new_[20499]_  = ~\new_[30070]_  | ~\new_[6197]_ ;
  assign \new_[20500]_  = ~\new_[29055]_  | ~\new_[6037]_ ;
  assign \new_[20501]_  = ~\new_[29452]_  | ~\new_[6057]_ ;
  assign \new_[20502]_  = ~\new_[29647]_  | ~\new_[6270]_ ;
  assign \new_[20503]_  = ~\new_[29989]_  | ~\new_[5925]_ ;
  assign \new_[20504]_  = ~\new_[29865]_  & ~\new_[30219]_ ;
  assign \new_[20505]_  = ~\new_[30682]_  | ~\new_[6270]_ ;
  assign \new_[20506]_  = ~\new_[29792]_  & ~\new_[28204]_ ;
  assign \new_[20507]_  = ~\new_[29767]_  & ~\new_[30141]_ ;
  assign \new_[20508]_  = ~\new_[29077]_  | ~\new_[6070]_ ;
  assign \new_[20509]_  = ~\new_[30632]_  | ~\new_[5984]_ ;
  assign \new_[20510]_  = ~\new_[29647]_  | ~\new_[6079]_ ;
  assign \new_[20511]_  = ~\new_[28846]_  | ~\new_[31422]_ ;
  assign \new_[20512]_  = ~\new_[29882]_  | ~\new_[6083]_ ;
  assign n8844 = m1_s13_cyc_o_reg;
  assign n8529 = m2_s11_cyc_o_reg;
  assign n8564 = m3_s11_cyc_o_reg;
  assign n8534 = m3_s13_cyc_o_reg;
  assign n8829 = m3_s4_cyc_o_reg;
  assign n8734 = m5_s2_cyc_o_reg;
  assign n8644 = m6_s2_cyc_o_reg;
  assign \new_[20520]_  = ~\new_[29767]_  & (~\new_[25154]_  | ~\new_[28575]_ );
  assign \new_[20521]_  = ~\new_[30633]_  | ~\new_[6032]_ ;
  assign \new_[20522]_  = ~\new_[26563]_  | ~\new_[31148]_ ;
  assign \new_[20523]_  = ~\new_[22918]_ ;
  assign \new_[20524]_  = ~\new_[28979]_  | ~\new_[5900]_ ;
  assign \new_[20525]_  = ~\new_[30304]_  & ~\new_[30069]_ ;
  assign \new_[20526]_  = ~\new_[29564]_  | ~\new_[5908]_ ;
  assign \new_[20527]_  = ~\new_[23675]_  | ~\new_[30525]_ ;
  assign \new_[20528]_  = ~\new_[30249]_  | ~\new_[6051]_ ;
  assign \new_[20529]_  = ~\new_[28845]_  | (~\new_[24945]_  & ~\new_[26513]_ );
  assign \new_[20530]_  = ~\new_[30020]_  | (~\new_[25097]_  & ~\new_[28398]_ );
  assign \new_[20531]_  = ~\new_[26623]_  | ~\new_[26768]_ ;
  assign \new_[20532]_  = ~\new_[30600]_  | (~\new_[24845]_  & ~\new_[26673]_ );
  assign \new_[20533]_  = ~\new_[30665]_  | (~\new_[24926]_  & ~\new_[27821]_ );
  assign \new_[20534]_  = ~\new_[30255]_  | (~\new_[24882]_  & ~\new_[27597]_ );
  assign \new_[20535]_  = ~\new_[30595]_  | (~\new_[24749]_  & ~\new_[28546]_ );
  assign \new_[20536]_  = ~\new_[29225]_  | (~\new_[25012]_  & ~\new_[26341]_ );
  assign \new_[20537]_  = ~\new_[29210]_  | (~\new_[25053]_  & ~\new_[26730]_ );
  assign \new_[20538]_  = ~\new_[29118]_  | (~\new_[25145]_  & ~\new_[28092]_ );
  assign \new_[20539]_  = ~\new_[25114]_  & ~\new_[23195]_ ;
  assign \new_[20540]_  = ~\new_[30145]_  & (~\new_[26869]_  | ~\new_[24790]_ );
  assign \new_[20541]_  = ~\new_[26881]_  & ~\new_[23198]_ ;
  assign \new_[20542]_  = ~\new_[24907]_  & ~\new_[23252]_ ;
  assign \new_[20543]_  = \new_[24817]_  | \new_[23198]_ ;
  assign \new_[20544]_  = ~\new_[24860]_  & ~\new_[23251]_ ;
  assign \new_[20545]_  = ~\new_[26956]_  & ~\new_[24186]_ ;
  assign \new_[20546]_  = ~\new_[23276]_  & ~\new_[24453]_ ;
  assign \new_[20547]_  = ~\new_[26947]_  & ~\new_[23211]_ ;
  assign \new_[20548]_  = ~\new_[23280]_  & ~\new_[26467]_ ;
  assign \new_[20549]_  = \new_[26897]_  | \new_[23251]_ ;
  assign \new_[20550]_  = ~\new_[24817]_  & ~\new_[23213]_ ;
  assign \new_[20551]_  = ~\new_[26947]_  & ~\new_[23218]_ ;
  assign \new_[20552]_  = \new_[23577]_  & \new_[24371]_ ;
  assign \new_[20553]_  = ~\new_[30201]_  & (~\new_[26928]_  | ~\new_[25015]_ );
  assign \new_[20554]_  = \new_[23149]_  & \new_[29104]_ ;
  assign \new_[20555]_  = \new_[24907]_  & \new_[24394]_ ;
  assign \new_[20556]_  = ~\new_[30038]_  & (~\new_[24906]_  | ~\new_[26923]_ );
  assign \new_[20557]_  = ~\new_[23270]_  & ~\new_[26356]_ ;
  assign \new_[20558]_  = \new_[23328]_  & \new_[26260]_ ;
  assign \new_[20559]_  = ~\new_[30029]_  & (~\new_[26290]_  | ~\new_[27599]_ );
  assign \new_[20560]_  = ~\new_[26881]_  & ~\new_[23213]_ ;
  assign \new_[20561]_  = ~\new_[23630]_  | ~\new_[27670]_ ;
  assign \new_[20562]_  = ~\new_[30213]_  | ~\new_[23274]_  | ~\new_[30645]_ ;
  assign \new_[20563]_  = ~\new_[30375]_  & (~\new_[24850]_  | ~\new_[24900]_ );
  assign \new_[20564]_  = ~\new_[29889]_  & (~\new_[27377]_  | ~\new_[24896]_ );
  assign \new_[20565]_  = ~\new_[23271]_  & ~\new_[24555]_ ;
  assign \new_[20566]_  = ~\new_[23169]_  & ~\new_[24149]_ ;
  assign \new_[20567]_  = \new_[23488]_  & \new_[24394]_ ;
  assign \new_[20568]_  = ~\new_[24860]_  & ~\new_[24411]_ ;
  assign \new_[20569]_  = ~\new_[30033]_  & (~\new_[25092]_  | ~\new_[25094]_ );
  assign \new_[20570]_  = \new_[25024]_  | \new_[23218]_ ;
  assign \new_[20571]_  = ~\new_[26849]_  & ~\new_[23195]_ ;
  assign \new_[20572]_  = ~\new_[24732]_  & ~\new_[23265]_ ;
  assign \new_[20573]_  = ~\new_[25063]_  & ~\new_[24186]_ ;
  assign \new_[20574]_  = ~\new_[23321]_  & ~\new_[24758]_ ;
  assign \new_[20575]_  = ~\new_[25024]_  & ~\new_[23211]_ ;
  assign \new_[20576]_  = \new_[24956]_  & \new_[23256]_ ;
  assign \new_[20577]_  = ~\new_[23279]_  & ~\new_[25775]_ ;
  assign \new_[20578]_  = \new_[26931]_  & \new_[23256]_ ;
  assign \new_[20579]_  = ~\new_[30325]_  & (~\new_[26883]_  | ~\new_[24689]_ );
  assign \new_[20580]_  = ~\new_[26987]_  & ~\new_[23265]_ ;
  assign \new_[20581]_  = ~\new_[30151]_  & (~\new_[25463]_  | ~\new_[25045]_ );
  assign \new_[20582]_  = ~\new_[29119]_  & (~\new_[25271]_  | ~\new_[28049]_ );
  assign \new_[20583]_  = ~\new_[23751]_  & (~\new_[28419]_  | ~\new_[26994]_ );
  assign \new_[20584]_  = ~\new_[28658]_  & (~\new_[24804]_  | ~\new_[24805]_ );
  assign \new_[20585]_  = ~\new_[30416]_  | ~\new_[27573]_  | ~\new_[25093]_  | ~\new_[26550]_ ;
  assign \new_[20586]_  = ~\new_[29855]_  & (~\new_[25157]_  | ~\new_[28412]_ );
  assign \new_[20587]_  = ~\new_[27427]_  & (~\new_[25081]_  | ~\new_[24565]_ );
  assign \new_[20588]_  = ~\new_[29648]_  & (~\new_[25191]_  | ~\new_[28474]_ );
  assign \new_[20589]_  = ~\new_[29565]_  & (~\new_[24635]_  | ~\new_[28373]_ );
  assign \new_[20590]_  = ~\new_[30713]_  & (~\new_[25162]_  | ~\new_[25121]_ );
  assign \new_[20591]_  = ~\new_[23388]_  & (~\new_[26251]_  | ~\new_[27001]_ );
  assign \new_[20592]_  = ~\new_[24300]_  & (~\new_[24808]_  | ~\new_[29028]_ );
  assign \new_[20593]_  = ~\new_[29100]_  & (~\new_[24657]_  | ~\new_[28222]_ );
  assign \new_[20594]_  = ~\new_[30174]_  & (~\new_[25202]_  | ~\new_[28481]_ );
  assign \new_[20595]_  = ~\new_[30769]_  & (~\new_[25169]_  | ~\new_[24867]_ );
  assign \new_[20596]_  = ~\new_[29199]_  & (~\new_[24943]_  | ~\new_[24858]_ );
  assign \new_[20597]_  = ~\new_[28685]_  & (~\new_[26895]_  | ~\new_[24859]_ );
  assign \new_[20598]_  = ~\new_[24863]_  & (~\new_[26246]_  | ~\new_[27003]_ );
  assign \new_[20599]_  = ~\new_[30389]_  & (~\new_[25167]_  | ~\new_[28500]_ );
  assign \new_[20600]_  = ~\new_[30174]_  & (~\new_[25202]_  | ~\new_[24866]_ );
  assign \new_[20601]_  = ~\new_[29132]_  & (~\new_[26965]_  | ~\new_[24872]_ );
  assign \new_[20602]_  = ~\new_[30762]_  & (~\new_[24875]_  | ~\new_[24876]_ );
  assign \new_[20603]_  = ~\new_[29315]_  & (~\new_[27458]_  | ~\new_[24877]_ );
  assign \new_[20604]_  = ~\new_[26880]_  & (~\new_[26905]_  | ~\new_[25170]_ );
  assign \new_[20605]_  = ~\new_[25084]_  & (~\new_[28065]_  | ~\new_[24578]_ );
  assign \new_[20606]_  = ~\new_[28899]_  & (~\new_[25161]_  | ~\new_[28181]_ );
  assign \new_[20607]_  = ~\new_[30711]_  & (~\new_[25175]_  | ~\new_[24889]_ );
  assign \new_[20608]_  = ~\new_[30661]_  & (~\new_[24687]_  | ~\new_[24836]_ );
  assign \new_[20609]_  = ~\new_[29898]_  & (~\new_[25183]_  | ~\new_[28108]_ );
  assign \new_[20610]_  = ~\new_[30044]_  & (~\new_[25177]_  | ~\new_[28508]_ );
  assign \new_[20611]_  = ~\new_[30443]_  & (~\new_[25180]_  | ~\new_[24912]_ );
  assign \new_[20612]_  = ~\new_[30044]_  & ~\new_[30355]_ ;
  assign \new_[20613]_  = ~\new_[30209]_  & (~\new_[24873]_  | ~\new_[24958]_ );
  assign \new_[20614]_  = ~\new_[29573]_  & (~\new_[25156]_  | ~\new_[28631]_ );
  assign \new_[20615]_  = ~\new_[30569]_  & (~\new_[24978]_  | ~\new_[25016]_ );
  assign \new_[20616]_  = ~\new_[28960]_  & (~\new_[26942]_  | ~\new_[24979]_ );
  assign \new_[20617]_  = ~\new_[30478]_  & (~\new_[25208]_  | ~\new_[24954]_ );
  assign \new_[20618]_  = ~\new_[26907]_  & (~\new_[26223]_  | ~\new_[24652]_ );
  assign \new_[20619]_  = ~\new_[29370]_  & (~\new_[25072]_  | ~\new_[24934]_ );
  assign \new_[20620]_  = ~\new_[25062]_  & (~\new_[27772]_  | ~\new_[25194]_ );
  assign \new_[20621]_  = ~\new_[28211]_  & (~\new_[24975]_  | ~\new_[25007]_ );
  assign \new_[20622]_  = ~\new_[29331]_  & (~\new_[24654]_  | ~\new_[26768]_ );
  assign \new_[20623]_  = ~\new_[29096]_  & (~\new_[25267]_  | ~\new_[28490]_ );
  assign \new_[20624]_  = ~\new_[24940]_  & (~\new_[24613]_  | ~\new_[25266]_ );
  assign \new_[20625]_  = ~\new_[29359]_  & (~\new_[25083]_  | ~\new_[25069]_ );
  assign \new_[20626]_  = ~\new_[28984]_  & (~\new_[26981]_  | ~\new_[25050]_ );
  assign \new_[20627]_  = ~\new_[30771]_  & (~\new_[25049]_  | ~\new_[25133]_ );
  assign \new_[20628]_  = ~\new_[29165]_  & (~\new_[25035]_  | ~\new_[24904]_ );
  assign \new_[20629]_  = ~\new_[30695]_  | ~\new_[27946]_  | ~\new_[24818]_  | ~\new_[25475]_ ;
  assign n7829 = ~\new_[28937]_  | ~\new_[23302]_ ;
  assign \new_[20631]_  = ~\new_[28992]_  | ~\new_[6036]_ ;
  assign \new_[20632]_  = ~\new_[28982]_  & (~\new_[25181]_  | ~\new_[28538]_ );
  assign \new_[20633]_  = ~\new_[29166]_  & (~\new_[25268]_  | ~\new_[26790]_ );
  assign \new_[20634]_  = ~\new_[30545]_  & (~\new_[25163]_  | ~\new_[24849]_ );
  assign \new_[20635]_  = ~\new_[28988]_  & (~\new_[26972]_  | ~\new_[25947]_ );
  assign \new_[20636]_  = ~\new_[25147]_  & (~\new_[28289]_  | ~\new_[25214]_ );
  assign \new_[20637]_  = ~\new_[30799]_  | ~\new_[27563]_  | ~\new_[23690]_  | ~\new_[24764]_ ;
  assign \new_[20638]_  = ~\new_[26494]_  & (~\new_[26968]_  | ~\new_[29911]_ );
  assign \new_[20639]_  = ~\new_[28499]_  & (~\new_[24815]_  | ~\new_[30015]_ );
  assign \new_[20640]_  = \new_[24526]_  & \new_[27904]_ ;
  assign \new_[20641]_  = \new_[23224]_  & \new_[27845]_ ;
  assign \new_[20642]_  = \new_[23203]_  & \new_[27926]_ ;
  assign \new_[20643]_  = ~\new_[24331]_  & (~\new_[24927]_  | ~\new_[30604]_ );
  assign \new_[20644]_  = \new_[23209]_  & \new_[27736]_ ;
  assign \new_[20645]_  = ~\new_[24303]_  & (~\new_[26909]_  | ~\new_[29763]_ );
  assign \new_[20646]_  = ~\new_[26242]_  & (~\new_[25099]_  | ~\new_[29505]_ );
  assign \new_[20647]_  = \new_[23238]_  & \new_[26940]_ ;
  assign \new_[20648]_  = ~\new_[24436]_  & (~\new_[24917]_  | ~\new_[29197]_ );
  assign \new_[20649]_  = ~\new_[26294]_  & (~\new_[24535]_  | ~\new_[30048]_ );
  assign \new_[20650]_  = ~\new_[24460]_  & (~\new_[24980]_  | ~\new_[30243]_ );
  assign \new_[20651]_  = \new_[23217]_  & \new_[27593]_ ;
  assign \new_[20652]_  = ~\new_[28745]_  & (~\new_[26444]_  | ~\new_[30434]_ );
  assign \new_[20653]_  = ~\new_[26717]_  & (~\new_[26565]_  | ~\new_[29781]_ );
  assign \new_[20654]_  = ~\new_[26354]_  & (~\new_[25070]_  | ~\new_[30467]_ );
  assign \new_[20655]_  = \new_[23237]_  & \new_[27769]_ ;
  assign \new_[20656]_  = ~\new_[26350]_  & (~\new_[25048]_  | ~\new_[30693]_ );
  assign \new_[20657]_  = ~\new_[26459]_  & (~\new_[25111]_  | ~\new_[30248]_ );
  assign \new_[20658]_  = ~\new_[26814]_  & (~\new_[25052]_  | ~\new_[30579]_ );
  assign \new_[20659]_  = \new_[23255]_  & \new_[27848]_ ;
  assign \new_[20660]_  = ~\new_[23114]_  & (~\new_[25132]_  | ~\new_[29825]_ );
  assign \new_[20661]_  = ~\new_[27783]_  & (~\new_[25144]_  | ~\new_[29768]_ );
  assign \new_[20662]_  = ~\new_[26728]_  & (~\new_[25103]_  | ~\new_[30233]_ );
  assign \new_[20663]_  = ~\new_[30104]_  | (~\new_[25139]_  & ~\new_[29172]_ );
  assign \new_[20664]_  = ~\new_[30283]_  | (~\new_[25122]_  & ~\new_[24798]_ );
  assign \new_[20665]_  = ~\new_[30416]_  | (~\new_[24888]_  & ~\new_[24963]_ );
  assign \new_[20666]_  = ~\new_[29966]_  & (~\new_[24831]_  | ~\new_[24829]_ );
  assign \new_[20667]_  = ~\new_[30508]_  | (~\new_[24835]_  & ~\new_[26891]_ );
  assign \new_[20668]_  = ~\new_[29736]_  & (~\new_[24822]_  | ~\new_[24853]_ );
  assign \new_[20669]_  = ~\new_[30750]_  | (~\new_[24857]_  & ~\new_[26898]_ );
  assign \new_[20670]_  = ~\new_[30695]_  | (~\new_[25078]_  & ~\new_[25064]_ );
  assign \new_[20671]_  = ~\new_[30273]_  & (~\new_[26911]_  | ~\new_[24995]_ );
  assign \new_[20672]_  = ~\new_[23214]_  & ~\new_[28944]_ ;
  assign \new_[20673]_  = ~\new_[30617]_  | (~\new_[24925]_  & ~\new_[24923]_ );
  assign \new_[20674]_  = ~\new_[30167]_  & (~\new_[24972]_  | ~\new_[27774]_ );
  assign \new_[20675]_  = ~\new_[24476]_  & ~\new_[30755]_ ;
  assign \new_[20676]_  = ~\new_[30752]_  | (~\new_[24932]_  & ~\new_[24936]_ );
  assign \new_[20677]_  = ~\new_[30645]_  | (~\new_[24986]_  & ~\new_[24991]_ );
  assign \new_[20678]_  = ~\new_[30782]_  | (~\new_[24996]_  & ~\new_[24988]_ );
  assign \new_[20679]_  = ~\new_[24170]_  & ~\new_[30348]_ ;
  assign \new_[20680]_  = ~\new_[30765]_  | (~\new_[25021]_  & ~\new_[26051]_ );
  assign \new_[20681]_  = ~\new_[30409]_  | (~\new_[24909]_  & ~\new_[30130]_ );
  assign \new_[20682]_  = ~\new_[30244]_  & (~\new_[25011]_  | ~\new_[25109]_ );
  assign \new_[20683]_  = ~\new_[30725]_  | (~\new_[24604]_  & ~\new_[25110]_ );
  assign \new_[20684]_  = ~\new_[29367]_  & (~\new_[25079]_  | ~\new_[26903]_ );
  assign \new_[20685]_  = ~\new_[23234]_  & ~\new_[30620]_ ;
  assign \new_[20686]_  = ~\new_[23247]_  & ~\new_[30070]_ ;
  assign \new_[20687]_  = ~\new_[30814]_  | (~\new_[24966]_  & ~\new_[25105]_ );
  assign \new_[20688]_  = ~\new_[30789]_  | (~\new_[26553]_  & ~\new_[25117]_ );
  assign \new_[20689]_  = ~\new_[30799]_  | (~\new_[24605]_  & ~\new_[25136]_ );
  assign \new_[20690]_  = ~\new_[30021]_  | (~\new_[24809]_  & ~\new_[24739]_ );
  assign \new_[20691]_  = ~\new_[24377]_  & (~\new_[24649]_  | ~\new_[28445]_ );
  assign \new_[20692]_  = ~\new_[23946]_  & (~\new_[25200]_  | ~\new_[28807]_ );
  assign \new_[20693]_  = ~\new_[26532]_  & (~\new_[24670]_  | ~\new_[28185]_ );
  assign \new_[20694]_  = ~\new_[24339]_  & (~\new_[25198]_  | ~\new_[28359]_ );
  assign \new_[20695]_  = ~\new_[24306]_  & (~\new_[25166]_  | ~\new_[28434]_ );
  assign \new_[20696]_  = ~\new_[24335]_  & (~\new_[25211]_  | ~\new_[28452]_ );
  assign \new_[20697]_  = ~\new_[26386]_  & (~\new_[25152]_  | ~\new_[28463]_ );
  assign \new_[20698]_  = ~\new_[24279]_  & (~\new_[25269]_  | ~\new_[28427]_ );
  assign \new_[20699]_  = ~\new_[29784]_  & (~\new_[24806]_  | ~\new_[28527]_ );
  assign \new_[20700]_  = ~\new_[24759]_  | ~\new_[6073]_ ;
  assign \new_[20701]_  = ~\new_[29966]_  & (~\new_[24829]_  | ~\new_[28586]_ );
  assign \new_[20702]_  = ~\new_[30215]_  | (~\new_[25075]_  & ~\new_[28727]_ );
  assign \new_[20703]_  = ~\new_[29736]_  & (~\new_[24853]_  | ~\new_[26901]_ );
  assign \new_[20704]_  = ~\new_[29260]_  | (~\new_[24855]_  & ~\new_[27978]_ );
  assign \new_[20705]_  = \new_[23241]_  & \new_[29305]_ ;
  assign \new_[20706]_  = ~\new_[30721]_  | (~\new_[24879]_  & ~\new_[25460]_ );
  assign \new_[20707]_  = ~\new_[30538]_  | (~\new_[26511]_  & ~\new_[29338]_ );
  assign \new_[20708]_  = ~\new_[23269]_  | ~\new_[30617]_ ;
  assign \new_[20709]_  = ~\new_[23272]_  | ~\new_[30434]_ ;
  assign \new_[20710]_  = ~\new_[30750]_  | (~\new_[26898]_  & ~\new_[26381]_ );
  assign \new_[20711]_  = \new_[23223]_  & \new_[29528]_ ;
  assign \new_[20712]_  = ~\new_[30244]_  & (~\new_[25109]_  | ~\new_[28838]_ );
  assign \new_[20713]_  = ~\new_[30765]_  | (~\new_[26051]_  & ~\new_[26804]_ );
  assign \new_[20714]_  = \new_[23229]_  & \new_[29351]_ ;
  assign \new_[20715]_  = ~\new_[30014]_  & (~\new_[25005]_  | ~\new_[29499]_ );
  assign \new_[20716]_  = ~\new_[30240]_  & (~\new_[24844]_  | ~\new_[27648]_ );
  assign \new_[20717]_  = ~\new_[30784]_  | (~\new_[26945]_  & ~\new_[24583]_ );
  assign \new_[20718]_  = ~\new_[29062]_  | ~\new_[31429]_ ;
  assign \new_[20719]_  = ~\new_[29367]_  & (~\new_[26903]_  | ~\new_[29449]_ );
  assign \new_[20720]_  = ~\new_[30125]_  | (~\new_[25010]_  & ~\new_[27860]_ );
  assign \new_[20721]_  = ~\new_[30789]_  | (~\new_[25117]_  & ~\new_[28800]_ );
  assign \new_[20722]_  = ~\new_[29874]_  | (~\new_[25104]_  & ~\new_[26679]_ );
  assign \new_[20723]_  = ~\new_[29383]_  & (~\new_[24802]_  | ~\new_[28569]_ );
  assign \new_[20724]_  = ~\new_[30021]_  | (~\new_[24739]_  & ~\new_[27555]_ );
  assign \new_[20725]_  = ~\new_[30273]_  & (~\new_[24995]_  | ~\new_[28540]_ );
  assign \new_[20726]_  = ~\new_[23889]_  & ~\new_[30342]_ ;
  assign \new_[20727]_  = ~\new_[23167]_  & ~\new_[29544]_ ;
  assign \new_[20728]_  = ~\new_[23917]_  & ~\new_[28402]_ ;
  assign \new_[20729]_  = ~\new_[23906]_  & ~\new_[29375]_ ;
  assign \new_[20730]_  = ~\new_[26994]_  & ~\new_[29367]_ ;
  assign \new_[20731]_  = ~\new_[23919]_  & ~\new_[30036]_ ;
  assign \new_[20732]_  = ~\new_[23332]_  & ~\new_[23170]_ ;
  assign \new_[20733]_  = \new_[23887]_  | \new_[26840]_ ;
  assign \new_[20734]_  = ~\new_[23652]_  | ~\new_[26581]_ ;
  assign \new_[20735]_  = ~\new_[23334]_  & ~\new_[29748]_ ;
  assign \new_[20736]_  = \new_[23634]_  & \new_[26769]_ ;
  assign \new_[20737]_  = ~\new_[23511]_  | ~\new_[27359]_ ;
  assign \new_[20738]_  = ~\new_[24524]_  | ~\new_[26201]_ ;
  assign \new_[20739]_  = \new_[23337]_  & \new_[23137]_ ;
  assign \new_[20740]_  = ~\new_[25034]_  | ~\new_[26973]_ ;
  assign \new_[20741]_  = \new_[23352]_  & \new_[26806]_ ;
  assign \new_[20742]_  = ~\new_[26875]_  | ~\new_[27431]_ ;
  assign \new_[20743]_  = ~\new_[30835]_  | ~\new_[6061]_ ;
  assign \new_[20744]_  = ~\new_[23729]_  & ~\new_[30275]_ ;
  assign \new_[20745]_  = \new_[23773]_  & \new_[23165]_ ;
  assign \new_[20746]_  = \new_[23390]_  & \new_[28501]_ ;
  assign \new_[20747]_  = ~\new_[24823]_  & ~\new_[23113]_ ;
  assign \new_[20748]_  = ~\new_[23929]_  | ~\new_[24675]_ ;
  assign \new_[20749]_  = ~\new_[23372]_  & ~\new_[30304]_ ;
  assign \new_[20750]_  = \new_[23761]_  | \new_[25107]_ ;
  assign \new_[20751]_  = ~\new_[23928]_  & ~\new_[30663]_ ;
  assign \new_[20752]_  = \new_[23752]_  | \new_[28727]_ ;
  assign \new_[20753]_  = ~\new_[23373]_  | ~\new_[27724]_ ;
  assign \new_[20754]_  = ~\new_[24687]_  | ~\new_[24461]_ ;
  assign \new_[20755]_  = ~\new_[23693]_  & ~\new_[30336]_ ;
  assign \new_[20756]_  = ~\new_[23449]_  & ~\new_[25058]_ ;
  assign \new_[20757]_  = ~\new_[23689]_  | ~\new_[23737]_ ;
  assign \new_[20758]_  = ~\new_[23895]_  & ~\new_[28846]_ ;
  assign \new_[20759]_  = ~\new_[23380]_  | ~\new_[28259]_ ;
  assign \new_[20760]_  = ~\new_[25054]_  & ~\new_[23693]_ ;
  assign \new_[20761]_  = \new_[23617]_  & \new_[26710]_ ;
  assign \new_[20762]_  = ~\new_[23384]_  & ~\new_[30591]_ ;
  assign \new_[20763]_  = \new_[23679]_  & \new_[24456]_ ;
  assign \new_[20764]_  = \new_[23671]_  | \new_[24869]_ ;
  assign \new_[20765]_  = ~\new_[23083]_  | ~\new_[24961]_ ;
  assign \new_[20766]_  = ~\new_[23660]_  & ~\new_[24839]_ ;
  assign \new_[20767]_  = ~\new_[23462]_  | ~\new_[28510]_ ;
  assign \new_[20768]_  = ~\new_[23706]_  | ~\new_[26403]_ ;
  assign \new_[20769]_  = ~\new_[25149]_  | ~\new_[23453]_ ;
  assign \new_[20770]_  = ~\new_[23404]_  & ~\new_[29810]_ ;
  assign \new_[20771]_  = \new_[23609]_  | \new_[27978]_ ;
  assign \new_[20772]_  = \new_[23849]_  & \new_[28241]_ ;
  assign \new_[20773]_  = ~\new_[23605]_  | ~\new_[27753]_ ;
  assign \new_[20774]_  = ~\new_[23520]_  & ~\new_[26314]_ ;
  assign \new_[20775]_  = ~\new_[23788]_  & ~\new_[26518]_ ;
  assign \new_[20776]_  = ~\new_[23884]_  | ~\new_[28074]_ ;
  assign \new_[20777]_  = \new_[23850]_  & \new_[28306]_ ;
  assign \new_[20778]_  = ~\new_[24927]_  | ~\new_[23422]_ ;
  assign \new_[20779]_  = ~\new_[23912]_  & ~\new_[30684]_ ;
  assign \new_[20780]_  = \new_[23480]_  & \new_[24281]_ ;
  assign \new_[20781]_  = \new_[24531]_  & \new_[27556]_ ;
  assign \new_[20782]_  = ~\new_[23678]_  | ~\new_[24665]_ ;
  assign \new_[20783]_  = ~\new_[23430]_  | ~\new_[23448]_ ;
  assign \new_[20784]_  = \new_[23791]_  & \new_[26847]_ ;
  assign \new_[20785]_  = \new_[23951]_  | \new_[27496]_ ;
  assign \new_[20786]_  = \new_[23671]_  | \new_[30785]_ ;
  assign \new_[20787]_  = ~\new_[23457]_  & ~\new_[30267]_ ;
  assign \new_[20788]_  = ~\new_[23432]_  & ~\new_[24881]_ ;
  assign \new_[20789]_  = ~\new_[24958]_  | ~\new_[27098]_ ;
  assign \new_[20790]_  = ~\new_[23357]_  | ~\new_[26256]_ ;
  assign \new_[20791]_  = ~\new_[23877]_  | ~\new_[23453]_ ;
  assign \new_[20792]_  = \new_[23753]_  | \new_[25460]_ ;
  assign \new_[20793]_  = \new_[23583]_  | \new_[27388]_ ;
  assign \new_[20794]_  = ~\new_[23770]_  | ~\new_[24464]_ ;
  assign \new_[20795]_  = ~\new_[23711]_  | ~\new_[29560]_ ;
  assign \new_[20796]_  = ~\new_[23537]_  | ~\new_[24924]_ ;
  assign \new_[20797]_  = \new_[23734]_  | \new_[24662]_ ;
  assign \new_[20798]_  = \new_[23444]_  & \new_[23968]_ ;
  assign \new_[20799]_  = \new_[23745]_  & \new_[28167]_ ;
  assign \new_[20800]_  = ~\new_[23731]_  | ~\new_[28231]_ ;
  assign \new_[20801]_  = \new_[23469]_  | \new_[24862]_ ;
  assign \new_[20802]_  = ~\new_[23487]_  | ~\new_[26418]_ ;
  assign \new_[20803]_  = ~\new_[23440]_  & ~\new_[29914]_ ;
  assign \new_[20804]_  = ~\new_[26873]_  | ~\new_[26878]_ ;
  assign \new_[20805]_  = ~\new_[26908]_  | ~\new_[26894]_ ;
  assign \new_[20806]_  = ~\new_[26736]_  | ~\new_[26867]_ ;
  assign \new_[20807]_  = ~\new_[21737]_ ;
  assign \new_[20808]_  = ~\new_[21738]_ ;
  assign \new_[20809]_  = ~\new_[23500]_  | ~\new_[26750]_ ;
  assign \new_[20810]_  = ~\new_[23540]_  | ~\new_[29977]_ ;
  assign \new_[20811]_  = ~\new_[21739]_ ;
  assign \new_[20812]_  = ~\new_[23516]_  | ~\new_[28144]_ ;
  assign \new_[20813]_  = \new_[32314]_ ;
  assign \new_[20814]_  = ~\new_[23482]_  | ~\new_[26750]_ ;
  assign \new_[20815]_  = ~\new_[23614]_  | ~\new_[24902]_ ;
  assign \new_[20816]_  = \new_[23665]_  & \new_[26727]_ ;
  assign \new_[20817]_  = ~\new_[23492]_  & ~\new_[23491]_ ;
  assign \new_[20818]_  = \new_[23634]_  & \new_[23766]_ ;
  assign \new_[20819]_  = ~\new_[23828]_  & ~\new_[25124]_ ;
  assign \new_[20820]_  = \new_[23360]_  & \new_[26664]_ ;
  assign \new_[20821]_  = \new_[23766]_  & \new_[26769]_ ;
  assign \new_[20822]_  = ~\new_[23915]_  | ~\new_[28139]_ ;
  assign \new_[20823]_  = ~\new_[23777]_  & ~\new_[29777]_ ;
  assign \new_[20824]_  = ~\new_[25083]_  | ~\new_[24329]_ ;
  assign \new_[20825]_  = ~\new_[26506]_  | ~\new_[23484]_ ;
  assign \new_[20826]_  = ~\new_[23494]_  | ~\new_[23401]_ ;
  assign \new_[20827]_  = ~\new_[23409]_  & ~\new_[24957]_ ;
  assign \new_[20828]_  = \new_[23798]_  | \new_[23777]_ ;
  assign \new_[20829]_  = ~\new_[24811]_  | ~\new_[23669]_ ;
  assign \new_[20830]_  = ~\new_[23481]_  | ~\new_[23484]_ ;
  assign \new_[20831]_  = \new_[23508]_  | \new_[28479]_ ;
  assign \new_[20832]_  = ~\new_[24913]_  & ~\new_[23729]_ ;
  assign \new_[20833]_  = ~\new_[23425]_  | ~\new_[23424]_ ;
  assign \new_[20834]_  = ~\new_[23362]_  & ~\new_[24820]_ ;
  assign \new_[20835]_  = ~\new_[23515]_  | ~\new_[24778]_ ;
  assign \new_[20836]_  = \new_[23725]_  & \new_[24751]_ ;
  assign \new_[20837]_  = \new_[23524]_  & \new_[23268]_ ;
  assign \new_[20838]_  = ~\new_[23870]_  | ~\new_[27950]_ ;
  assign \new_[20839]_  = ~\new_[24893]_  | ~\new_[23736]_ ;
  assign \new_[20840]_  = ~\new_[25071]_  | ~\new_[26941]_ ;
  assign \new_[20841]_  = ~\new_[23340]_  | ~\new_[28494]_ ;
  assign \new_[20842]_  = ~\new_[23933]_  | ~\new_[28802]_ ;
  assign \new_[20843]_  = ~\new_[23580]_  | ~\new_[24778]_ ;
  assign \new_[20844]_  = \new_[23539]_  | \new_[27610]_ ;
  assign \new_[20845]_  = ~\new_[23757]_  | ~\new_[24942]_ ;
  assign \new_[20846]_  = ~\new_[23575]_  | ~\new_[23657]_ ;
  assign \new_[20847]_  = \new_[23645]_  | \new_[28707]_ ;
  assign \new_[20848]_  = ~\new_[23550]_  | ~\new_[28565]_ ;
  assign \new_[20849]_  = ~\new_[24876]_  | ~\new_[26933]_ ;
  assign \new_[20850]_  = ~\new_[23728]_  | ~\new_[24949]_ ;
  assign \new_[20851]_  = \new_[23459]_  & \new_[26675]_ ;
  assign \new_[20852]_  = ~\new_[23564]_  | ~\new_[26741]_ ;
  assign \new_[20853]_  = ~\new_[23567]_  & ~\new_[29994]_ ;
  assign \new_[20854]_  = \new_[23914]_  | \new_[27281]_ ;
  assign \new_[20855]_  = \new_[23571]_  | \new_[26629]_ ;
  assign \new_[20856]_  = ~\new_[23647]_  & ~\new_[30710]_ ;
  assign \new_[20857]_  = \new_[23601]_  | \new_[29338]_ ;
  assign \new_[20858]_  = ~\new_[23416]_  | ~\new_[23414]_ ;
  assign \new_[20859]_  = \new_[23593]_  & \new_[26755]_ ;
  assign \new_[20860]_  = ~\new_[24535]_  | ~\new_[23586]_ ;
  assign \new_[20861]_  = ~\new_[23412]_  | ~\new_[24967]_ ;
  assign \new_[20862]_  = ~\new_[23703]_  | ~\new_[28554]_ ;
  assign \new_[20863]_  = ~\new_[23411]_  | ~\new_[24967]_ ;
  assign \new_[20864]_  = ~\new_[23694]_  & ~\new_[23692]_ ;
  assign \new_[20865]_  = ~\new_[23359]_  & ~\new_[25966]_ ;
  assign \new_[20866]_  = ~\new_[29629]_  | ~\new_[5907]_ ;
  assign \new_[20867]_  = ~\new_[23801]_  | ~\new_[28674]_ ;
  assign \new_[20868]_  = ~\new_[23949]_  | ~\new_[28743]_ ;
  assign \new_[20869]_  = \new_[23371]_  & \new_[23166]_ ;
  assign \new_[20870]_  = ~\new_[25098]_  & ~\new_[23778]_ ;
  assign \new_[20871]_  = ~\new_[23410]_  | ~\new_[27753]_ ;
  assign \new_[20872]_  = ~\new_[23607]_  | ~\new_[26809]_ ;
  assign \new_[20873]_  = ~\new_[23599]_  | ~\new_[26319]_ ;
  assign \new_[20874]_  = ~\new_[23722]_  | ~\new_[23732]_ ;
  assign \new_[20875]_  = \new_[23504]_  | \new_[30662]_ ;
  assign \new_[20876]_  = ~\new_[23894]_  & ~\new_[30747]_ ;
  assign \new_[20877]_  = ~\new_[23473]_  | ~\new_[24274]_ ;
  assign \new_[20878]_  = ~\new_[25185]_  & ~\new_[30028]_ ;
  assign \new_[20879]_  = ~\new_[23761]_  & ~\new_[29772]_ ;
  assign \new_[20880]_  = ~\new_[24917]_  | ~\new_[23510]_ ;
  assign \new_[20881]_  = ~\new_[23361]_  | ~\new_[26795]_ ;
  assign \new_[20882]_  = ~\new_[24848]_  & ~\new_[23404]_ ;
  assign \new_[20883]_  = ~\new_[23985]_  & ~\new_[26431]_ ;
  assign \new_[20884]_  = ~\new_[23625]_  | ~\new_[28416]_ ;
  assign \new_[20885]_  = ~\new_[23497]_  | ~\new_[26874]_ ;
  assign \new_[20886]_  = ~\new_[23490]_  | ~\new_[23860]_ ;
  assign \new_[20887]_  = \new_[24506]_  | \new_[27638]_ ;
  assign \new_[20888]_  = ~\new_[25069]_  | ~\new_[24329]_ ;
  assign \new_[20889]_  = ~\new_[23893]_  | ~\new_[28525]_ ;
  assign \new_[20890]_  = ~\new_[23640]_  | ~\new_[28905]_ ;
  assign \new_[20891]_  = \new_[23658]_  | \new_[25026]_ ;
  assign \new_[20892]_  = ~\new_[23664]_  & ~\new_[23566]_ ;
  assign \new_[20893]_  = \new_[23567]_  | \new_[24952]_ ;
  assign \new_[20894]_  = \new_[23881]_  | \new_[24583]_ ;
  assign \new_[20895]_  = ~\new_[23859]_  & ~\new_[29828]_ ;
  assign \new_[20896]_  = ~\new_[26959]_  | ~\new_[24500]_ ;
  assign \new_[20897]_  = \new_[23392]_  & \new_[27093]_ ;
  assign \new_[20898]_  = ~\new_[23873]_  & ~\new_[30597]_ ;
  assign \new_[20899]_  = \new_[23504]_  | \new_[25025]_ ;
  assign \new_[20900]_  = \new_[23733]_  | \new_[29792]_ ;
  assign \new_[20901]_  = \new_[23562]_  & \new_[28559]_ ;
  assign \new_[20902]_  = ~\new_[23374]_  | ~\new_[24832]_ ;
  assign \new_[20903]_  = ~\new_[23338]_  & ~\new_[24989]_ ;
  assign \new_[20904]_  = ~\new_[23774]_  | ~\new_[24973]_ ;
  assign \new_[20905]_  = \new_[23469]_  | \new_[30649]_ ;
  assign \new_[20906]_  = ~\new_[23742]_  | ~\new_[26373]_ ;
  assign \new_[20907]_  = \new_[23496]_  & \new_[28772]_ ;
  assign \new_[20908]_  = \new_[23560]_  & \new_[26248]_ ;
  assign \new_[20909]_  = ~\new_[23948]_  | ~\new_[28230]_ ;
  assign \new_[20910]_  = ~\new_[23629]_  | ~\new_[23698]_ ;
  assign \new_[20911]_  = ~\new_[23363]_  | ~\new_[23572]_ ;
  assign \new_[20912]_  = ~\new_[23825]_  | ~\new_[25708]_ ;
  assign \new_[20913]_  = ~\new_[23643]_  | ~\new_[25080]_ ;
  assign \new_[20914]_  = ~\new_[23389]_  | ~\new_[28570]_ ;
  assign \new_[20915]_  = ~\new_[26949]_  | ~\new_[24500]_ ;
  assign \new_[20916]_  = ~\new_[23561]_  | ~\new_[26941]_ ;
  assign \new_[20917]_  = ~\new_[23779]_  & ~\new_[25031]_ ;
  assign \new_[20918]_  = \new_[23499]_  & \new_[26738]_ ;
  assign \new_[20919]_  = ~\new_[25110]_  & ~\new_[24341]_ ;
  assign \new_[20920]_  = \new_[23901]_  | \new_[26178]_ ;
  assign \new_[20921]_  = ~\new_[24837]_  | ~\new_[23387]_ ;
  assign \new_[20922]_  = ~\new_[23808]_  | ~\new_[25469]_ ;
  assign \new_[20923]_  = \new_[24483]_  | \new_[30323]_ ;
  assign \new_[20924]_  = ~\new_[25099]_  | ~\new_[23655]_ ;
  assign \new_[20925]_  = ~\new_[23554]_  | ~\new_[24948]_ ;
  assign \new_[20926]_  = \new_[23514]_  & \new_[24541]_ ;
  assign \new_[20927]_  = ~\new_[23723]_  | ~\new_[24993]_ ;
  assign \new_[20928]_  = ~\new_[23930]_  & ~\new_[30557]_ ;
  assign \new_[20929]_  = \new_[23962]_  & \new_[24307]_ ;
  assign \new_[20930]_  = ~\new_[23454]_  | ~\new_[28565]_ ;
  assign \new_[20931]_  = ~\new_[23798]_  & ~\new_[29777]_ ;
  assign \new_[20932]_  = \new_[23331]_  | \new_[27993]_ ;
  assign \new_[20933]_  = ~\new_[23626]_  | ~\new_[23086]_ ;
  assign \new_[20934]_  = ~\new_[23606]_  | ~\new_[26809]_ ;
  assign \new_[20935]_  = \new_[23947]_  | \new_[27521]_ ;
  assign \new_[20936]_  = ~\new_[23758]_  | ~\new_[25253]_ ;
  assign \new_[20937]_  = ~\new_[23370]_  & ~\new_[23113]_ ;
  assign \new_[20938]_  = ~\new_[23553]_  | ~\new_[23787]_ ;
  assign \new_[20939]_  = ~\new_[23762]_  | ~\new_[24941]_ ;
  assign \new_[20940]_  = ~\new_[24604]_  & ~\new_[24341]_ ;
  assign \new_[20941]_  = \new_[23658]_  | \new_[30581]_ ;
  assign \new_[20942]_  = ~\new_[23898]_  & ~\new_[28317]_ ;
  assign \new_[20943]_  = \new_[23905]_  | \new_[27494]_ ;
  assign \new_[20944]_  = ~\new_[23769]_  | ~\new_[26197]_ ;
  assign \new_[20945]_  = ~\new_[21884]_ ;
  assign \new_[20946]_  = ~\new_[23541]_  | ~\new_[26980]_ ;
  assign \new_[20947]_  = ~\new_[23670]_  & ~\new_[23827]_ ;
  assign \new_[20948]_  = ~\new_[23778]_  & ~\new_[30326]_ ;
  assign \new_[20949]_  = ~\new_[23781]_  | ~\new_[30021]_ ;
  assign \new_[20950]_  = \new_[23600]_  | \new_[30618]_ ;
  assign \new_[20951]_  = \new_[23533]_  | \new_[30568]_ ;
  assign \new_[20952]_  = \new_[23533]_  | \new_[24937]_ ;
  assign \new_[20953]_  = ~\new_[23903]_  | ~\new_[26757]_ ;
  assign \new_[20954]_  = ~\new_[23650]_  | ~\new_[24577]_ ;
  assign \new_[20955]_  = ~\new_[25143]_  | ~\new_[27557]_ ;
  assign \new_[20956]_  = \new_[23354]_  | \new_[26948]_ ;
  assign \new_[20957]_  = \new_[23600]_  | \new_[25102]_ ;
  assign \new_[20958]_  = ~\new_[23865]_  | ~\new_[24738]_ ;
  assign \new_[20959]_  = ~\new_[23558]_  | ~\new_[26336]_ ;
  assign \new_[20960]_  = \new_[24811]_  | \new_[23669]_ ;
  assign \new_[20961]_  = ~\new_[26506]_  & ~\new_[23484]_ ;
  assign \new_[20962]_  = ~\new_[23409]_  | ~\new_[24957]_ ;
  assign \new_[20963]_  = ~\new_[21925]_ ;
  assign \new_[20964]_  = ~\new_[23537]_  & ~\new_[24924]_ ;
  assign \new_[20965]_  = ~\new_[23797]_  | ~\new_[23080]_ ;
  assign \new_[20966]_  = \new_[23701]_  | \new_[27697]_ ;
  assign \new_[20967]_  = ~\new_[23809]_  & ~\new_[24644]_ ;
  assign \new_[20968]_  = ~\new_[24028]_  | ~\new_[25029]_ ;
  assign \new_[20969]_  = ~\new_[24837]_  & ~\new_[23387]_ ;
  assign \new_[20970]_  = ~\new_[23821]_  | ~\new_[24993]_ ;
  assign \new_[20971]_  = ~\new_[23950]_  & ~\new_[30682]_ ;
  assign \new_[20972]_  = ~\new_[23528]_  & ~\new_[23526]_ ;
  assign \new_[20973]_  = ~\new_[23666]_  | ~\new_[26866]_ ;
  assign \new_[20974]_  = \new_[23824]_  | \new_[27689]_ ;
  assign \new_[20975]_  = \new_[23527]_  | \new_[24928]_ ;
  assign \new_[20976]_  = ~\new_[23826]_  | ~\new_[28086]_ ;
  assign \new_[20977]_  = ~\new_[23465]_  & ~\new_[30268]_ ;
  assign \new_[20978]_  = \new_[23920]_  | \new_[27341]_ ;
  assign \new_[20979]_  = ~\new_[23527]_  & ~\new_[29865]_ ;
  assign \new_[20980]_  = \new_[23851]_  & \new_[23087]_ ;
  assign \new_[20981]_  = ~\new_[23719]_  | ~\new_[28643]_ ;
  assign \new_[20982]_  = ~\new_[23828]_  | ~\new_[25124]_ ;
  assign \new_[20983]_  = ~\new_[23886]_  | ~\new_[28644]_ ;
  assign \new_[20984]_  = ~\new_[23336]_  | ~\new_[28555]_ ;
  assign \new_[20985]_  = \new_[23838]_  & \new_[24544]_ ;
  assign \new_[20986]_  = \new_[23483]_  & \new_[26428]_ ;
  assign \new_[20987]_  = \new_[23718]_  & \new_[28154]_ ;
  assign \new_[20988]_  = ~\new_[23471]_  | ~\new_[26704]_ ;
  assign \new_[20989]_  = ~\new_[23843]_  & ~\new_[30208]_ ;
  assign \new_[20990]_  = \new_[23522]_  & \new_[28048]_ ;
  assign \new_[20991]_  = \new_[23843]_  | \new_[25134]_ ;
  assign \new_[20992]_  = ~\new_[23844]_  & ~\new_[23842]_ ;
  assign \new_[20993]_  = ~\new_[23405]_  | ~\new_[28368]_ ;
  assign \new_[20994]_  = ~\new_[23685]_  | ~\new_[26590]_ ;
  assign \new_[20995]_  = \new_[23856]_  | \new_[25137]_ ;
  assign \new_[20996]_  = \new_[23856]_  | \new_[30521]_ ;
  assign \new_[20997]_  = ~\new_[23892]_  | ~\new_[28604]_ ;
  assign \new_[20998]_  = ~\new_[23862]_  | ~\new_[28483]_ ;
  assign \new_[20999]_  = ~\new_[23341]_  | ~\new_[26194]_ ;
  assign \new_[21000]_  = ~\new_[23855]_  | ~\new_[24737]_ ;
  assign \new_[21001]_  = \new_[23871]_  | \new_[29372]_ ;
  assign \new_[21002]_  = ~\new_[23784]_  | ~\new_[23879]_ ;
  assign \new_[21003]_  = \new_[23882]_  & \new_[24709]_ ;
  assign \new_[21004]_  = ~\new_[29873]_  | ~\new_[26840]_  | ~\new_[26674]_ ;
  assign \new_[21005]_  = ~\new_[30145]_  & (~\new_[25944]_  | ~\new_[29500]_ );
  assign \new_[21006]_  = \new_[23624]_  | \new_[29561]_ ;
  assign \new_[21007]_  = ~\new_[26489]_  | ~\new_[26372]_  | ~\new_[28378]_ ;
  assign \new_[21008]_  = ~\new_[24720]_  | ~\new_[27508]_  | ~\new_[29117]_ ;
  assign \new_[21009]_  = \new_[23702]_  | \new_[28566]_ ;
  assign \new_[21010]_  = ~\new_[23509]_  | ~\new_[27642]_ ;
  assign \new_[21011]_  = ~\new_[26282]_  | ~\new_[25129]_  | ~\new_[28511]_ ;
  assign \new_[21012]_  = ~\new_[24683]_  | ~\new_[27360]_  | ~\new_[29128]_ ;
  assign \new_[21013]_  = \new_[23535]_  | \new_[28341]_ ;
  assign \new_[21014]_  = ~\new_[30552]_  | ~\new_[23518]_  | ~\new_[27673]_ ;
  assign \new_[21015]_  = ~\new_[30201]_  & (~\new_[26325]_  | ~\new_[29577]_ );
  assign n8444 = m7_s9_cyc_o_reg;
  assign \new_[21017]_  = ~\new_[26235]_  | ~\new_[26323]_  | ~\new_[28187]_ ;
  assign \new_[21018]_  = \new_[23822]_  | \new_[27994]_ ;
  assign \new_[21019]_  = ~\new_[29889]_  & (~\new_[26415]_  | ~\new_[29344]_ );
  assign \new_[21020]_  = ~\new_[23419]_  | ~\new_[26795]_ ;
  assign \new_[21021]_  = ~\new_[26202]_  | ~\new_[28253]_  | ~\new_[28567]_ ;
  assign \new_[21022]_  = \new_[23673]_  | \new_[28784]_ ;
  assign \new_[21023]_  = ~\new_[24557]_  | ~\new_[25996]_  | ~\new_[28413]_ ;
  assign n7809 = ~\new_[29093]_  | ~\new_[23945]_ ;
  assign n8489 = m7_s13_cyc_o_reg;
  assign n8674 = m7_s2_cyc_o_reg;
  assign n7789 = ~\new_[29497]_  | ~\new_[23943]_ ;
  assign \new_[21028]_  = \new_[23602]_  | \new_[28221]_ ;
  assign n7799 = ~\new_[28892]_  | ~\new_[23931]_ ;
  assign \new_[21030]_  = ~\new_[26164]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[21031]_  = ~\new_[26156]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign n8894 = m7_s14_cyc_o_reg;
  assign n7779 = ~\new_[29734]_  | ~\new_[23935]_ ;
  assign n7784 = ~\new_[28902]_  | ~\new_[23936]_ ;
  assign \new_[21035]_  = ~\new_[26173]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign n8599 = m7_s10_cyc_o_reg;
  assign n8574 = m6_s7_cyc_o_reg;
  assign \new_[21038]_  = ~\new_[26175]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign n7819 = ~\new_[29618]_  | ~\new_[23938]_ ;
  assign n7824 = ~\new_[29312]_  | ~\new_[23112]_ ;
  assign n8654 = m6_s6_cyc_o_reg;
  assign n7804 = ~\new_[29075]_  | ~\new_[23942]_ ;
  assign n7814 = ~\new_[29288]_  | ~\new_[23932]_ ;
  assign \new_[21044]_  = ~\new_[26243]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign n7794 = ~\new_[29654]_  | ~\new_[23944]_ ;
  assign \new_[21046]_  = ~\new_[25239]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign n8604 = m6_s11_cyc_o_reg;
  assign \new_[21048]_  = ~\new_[25155]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[21049]_  = \new_[22413]_ ;
  assign n8924 = m5_s9_cyc_o_reg;
  assign n7774 = ~\new_[29198]_  | ~\new_[23934]_ ;
  assign n8854 = m6_s10_cyc_o_reg;
  assign \new_[21053]_  = \new_[23857]_  | \new_[28454]_ ;
  assign \new_[21054]_  = ~\new_[30325]_  & (~\new_[26442]_  | ~\new_[28871]_ );
  assign \new_[21055]_  = ~\new_[22413]_ ;
  assign \new_[21056]_  = ~\new_[24283]_  | (~\new_[26218]_  & ~\new_[30736]_ );
  assign \new_[21057]_  = ~\new_[23353]_  & ~\new_[27743]_ ;
  assign n8839 = m5_s7_cyc_o_reg;
  assign \new_[21059]_  = \new_[23493]_  & \new_[27576]_ ;
  assign \new_[21060]_  = ~\new_[26552]_  & (~\new_[29572]_  | ~\new_[30767]_ );
  assign \new_[21061]_  = ~\new_[26274]_  | (~\new_[26361]_  & ~\new_[29736]_ );
  assign \new_[21062]_  = ~\new_[23427]_  | ~\new_[30222]_ ;
  assign \new_[21063]_  = ~\new_[23433]_  & ~\new_[28098]_ ;
  assign \new_[21064]_  = ~\new_[23538]_  | (~\new_[24591]_  & ~\new_[30055]_ );
  assign n8434 = m5_s14_cyc_o_reg;
  assign n8329 = m5_s3_cyc_o_reg;
  assign \new_[21067]_  = ~\new_[24314]_  | (~\new_[25046]_  & ~\new_[29544]_ );
  assign \new_[21068]_  = ~\new_[23368]_  | ~\new_[30242]_ ;
  assign \new_[21069]_  = ~\new_[23765]_  & ~\new_[28380]_ ;
  assign \new_[21070]_  = ~\new_[23638]_  | ~\new_[28818]_ ;
  assign \new_[21071]_  = ~\new_[23699]_  | ~\new_[29808]_ ;
  assign \new_[21072]_  = ~\new_[24376]_  | (~\new_[26238]_  & ~\new_[30342]_ );
  assign \new_[21073]_  = ~\new_[23364]_  | ~\new_[30599]_ ;
  assign n8324 = m5_s13_cyc_o_reg;
  assign \new_[21075]_  = ~\new_[24352]_  & (~\new_[29531]_  | ~\new_[28215]_ );
  assign \new_[21076]_  = ~\new_[26085]_  | (~\new_[26368]_  & ~\new_[30400]_ );
  assign \new_[21077]_  = ~\new_[24475]_  | (~\new_[26667]_  & ~\new_[30273]_ );
  assign \new_[21078]_  = \new_[23656]_  & \new_[27706]_ ;
  assign n8339 = m5_s11_cyc_o_reg;
  assign \new_[21080]_  = ~\new_[24063]_  & (~\new_[29439]_  | ~\new_[28057]_ );
  assign \new_[21081]_  = ~\new_[26169]_  | (~\new_[24640]_  & ~\new_[28857]_ );
  assign \new_[21082]_  = ~\new_[23672]_  | ~\new_[30693]_ ;
  assign \new_[21083]_  = ~\new_[23688]_  | ~\new_[30229]_ ;
  assign \new_[21084]_  = ~\new_[25660]_  | (~\new_[26377]_  & ~\new_[30173]_ );
  assign \new_[21085]_  = ~\new_[23704]_  | ~\new_[30198]_ ;
  assign \new_[21086]_  = ~\new_[23807]_  | ~\new_[30248]_ ;
  assign \new_[21087]_  = ~\new_[23636]_  | ~\new_[29987]_ ;
  assign \new_[21088]_  = ~\new_[24002]_  & (~\new_[29566]_  | ~\new_[30099]_ );
  assign n8429 = m4_s11_cyc_o_reg;
  assign \new_[21090]_  = ~\new_[25315]_  | (~\new_[26406]_  & ~\new_[29966]_ );
  assign \new_[21091]_  = ~\new_[23829]_  | ~\new_[29583]_ ;
  assign \new_[21092]_  = ~\new_[23505]_  | ~\new_[29869]_ ;
  assign \new_[21093]_  = ~\new_[24354]_  | (~\new_[26255]_  & ~\new_[30407]_ );
  assign \new_[21094]_  = ~\new_[23760]_  | ~\new_[30297]_ ;
  assign \new_[21095]_  = ~\new_[23776]_  | ~\new_[30015]_ ;
  assign n8739 = m4_s2_cyc_o_reg;
  assign \new_[21097]_  = ~\new_[23800]_  | ~\new_[30248]_ ;
  assign \new_[21098]_  = ~\new_[23816]_  | ~\new_[29851]_ ;
  assign \new_[21099]_  = ~\new_[23333]_  & ~\new_[27639]_ ;
  assign \new_[21100]_  = ~\new_[24458]_  | (~\new_[27531]_  & ~\new_[30276]_ );
  assign \new_[21101]_  = ~\new_[23878]_  | ~\new_[30233]_ ;
  assign \new_[21102]_  = ~\new_[30416]_  | ~\new_[6174]_  | ~\new_[30828]_  | ~\new_[26550]_ ;
  assign \new_[21103]_  = ~\new_[30647]_  | ~\new_[31400]_  | ~\new_[30667]_  | ~\new_[26396]_ ;
  assign \new_[21104]_  = ~\new_[30676]_  | ~\new_[6043]_  | ~\new_[30678]_  | ~\new_[26556]_ ;
  assign \new_[21105]_  = ~\new_[30695]_  | ~\new_[6049]_  | ~\new_[30499]_  | ~\new_[25475]_ ;
  assign \new_[21106]_  = ~\new_[30765]_  | ~\new_[6213]_  | ~\new_[29869]_  | ~\new_[26402]_ ;
  assign \new_[21107]_  = ~\new_[30752]_  | ~\new_[6197]_  | ~\new_[30691]_  | ~\new_[26212]_ ;
  assign \new_[21108]_  = ~\new_[30782]_  | ~\new_[6211]_  | ~\new_[30638]_  | ~\new_[26367]_ ;
  assign \new_[21109]_  = ~\new_[30814]_  | ~\new_[6194]_  | ~\new_[30653]_  | ~\new_[26244]_ ;
  assign \new_[21110]_  = ~\new_[30563]_  | ~\new_[6076]_  | ~\new_[30846]_  | ~\new_[26302]_ ;
  assign \new_[21111]_  = ~\new_[30610]_  | ~\new_[6268]_  | ~\new_[29851]_  | ~\new_[24617]_ ;
  assign \new_[21112]_  = ~\new_[30820]_  | ~\new_[6095]_  | ~\new_[30233]_  | ~\new_[25209]_ ;
  assign \new_[21113]_  = \new_[30057]_  | \new_[31569]_ ;
  assign \new_[21114]_  = ~\new_[30630]_  | ~\new_[6079]_  | ~\new_[30635]_  | ~\new_[25357]_ ;
  assign \new_[21115]_  = ~\new_[30799]_  | ~\new_[6093]_  | ~\new_[30641]_  | ~\new_[24764]_ ;
  assign n8569 = m2_s4_cyc_o_reg;
  assign n8774 = m3_s5_cyc_o_reg;
  assign \new_[21118]_  = ~\new_[24379]_  | ~\new_[27585]_ ;
  assign \new_[21119]_  = ~\new_[29293]_  & ~\new_[23258]_ ;
  assign n8649 = m3_s6_cyc_o_reg;
  assign \new_[21121]_  = ~\new_[22111]_ ;
  assign \new_[21122]_  = ~\new_[6035]_  | ~\new_[28064]_  | ~\new_[29784]_ ;
  assign n8504 = m3_s7_cyc_o_reg;
  assign \new_[21124]_  = ~\new_[6203]_  | ~\new_[29547]_  | ~\new_[30736]_ ;
  assign n8679 = m3_s3_cyc_o_reg;
  assign \new_[21126]_  = ~\new_[27637]_  & ~\new_[30642]_ ;
  assign n8624 = m3_s14_cyc_o_reg;
  assign \new_[21128]_  = ~\new_[23093]_  & ~\new_[29815]_ ;
  assign \new_[21129]_  = ~\new_[24325]_  & ~\new_[30660]_ ;
  assign \new_[21130]_  = ~\new_[24240]_  & ~\new_[30663]_ ;
  assign \new_[21131]_  = ~\new_[24240]_  | ~\new_[24512]_ ;
  assign n8544 = m3_s12_cyc_o_reg;
  assign n8314 = m2_s8_cyc_o_reg;
  assign \new_[21134]_  = ~\new_[6039]_  | ~\new_[26672]_  | ~\new_[29966]_ ;
  assign n8499 = m2_s7_cyc_o_reg;
  assign \new_[21136]_  = ~\new_[22129]_ ;
  assign \new_[21137]_  = ~\new_[29565]_  | ~\new_[6075]_ ;
  assign \new_[21138]_  = ~\new_[22130]_ ;
  assign \new_[21139]_  = ~\new_[6041]_  | ~\new_[28034]_  | ~\new_[30425]_ ;
  assign \new_[21140]_  = ~\new_[28078]_  & ~\new_[24433]_ ;
  assign n8469 = m2_s13_cyc_o_reg;
  assign \new_[21142]_  = ~\new_[31733]_  | ~\new_[27577]_  | ~\new_[30022]_ ;
  assign n8824 = m2_s14_cyc_o_reg;
  assign n8769 = m2_s2_cyc_o_reg;
  assign \new_[21145]_  = ~\new_[27196]_  & ~\new_[30521]_ ;
  assign n8394 = m1_s7_cyc_o_reg;
  assign n8634 = m1_s9_cyc_o_reg;
  assign \new_[21148]_  = ~\new_[21561]_ ;
  assign \new_[21149]_  = ~\new_[30323]_  & ~\new_[24436]_ ;
  assign \new_[21150]_  = ~\new_[31751]_  | ~\new_[26083]_  | ~\new_[29983]_ ;
  assign n8724 = m1_s2_cyc_o_reg;
  assign \new_[21152]_  = ~\new_[31819]_  | ~\new_[27561]_  | ~\new_[27802]_ ;
  assign \new_[21153]_  = ~\new_[31551]_  | ~\new_[27736]_  | ~\new_[27787]_ ;
  assign \new_[21154]_  = ~\new_[30404]_  & ~\new_[24419]_ ;
  assign \new_[21155]_  = ~\new_[30261]_  & ~\new_[24403]_ ;
  assign n8889 = m1_s14_cyc_o_reg;
  assign \new_[21157]_  = ~\new_[29999]_  & ~\new_[23114]_ ;
  assign \new_[21158]_  = ~\new_[22162]_ ;
  assign \new_[21159]_  = ~\new_[24316]_  | ~\new_[29226]_ ;
  assign \new_[21160]_  = ~\new_[31521]_  | ~\new_[26267]_  | ~\new_[30117]_ ;
  assign n8464 = m1_s11_cyc_o_reg;
  assign \new_[21162]_  = ~\new_[6199]_  | ~\new_[28367]_  | ~\new_[28317]_ ;
  assign \new_[21163]_  = ~\new_[24328]_  | ~\new_[30505]_ ;
  assign \new_[21164]_  = ~\new_[22173]_ ;
  assign n8459 = m3_s2_cyc_o_reg;
  assign \new_[21166]_  = ~\new_[28404]_  & ~\new_[29564]_ ;
  assign n8754 = m0_s14_cyc_o_reg;
  assign \new_[21168]_  = ~\new_[6200]_  | ~\new_[29760]_  | ~\new_[30757]_ ;
  assign \new_[21169]_  = ~\new_[22180]_ ;
  assign \new_[21170]_  = ~\new_[22188]_ ;
  assign \new_[21171]_  = ~\new_[24392]_  | ~\new_[26715]_ ;
  assign \new_[21172]_  = ~\new_[22190]_ ;
  assign \new_[21173]_  = ~\new_[22191]_ ;
  assign \new_[21174]_  = ~\new_[29830]_  & ~\new_[24311]_ ;
  assign n8389 = m0_s4_cyc_o_reg;
  assign \new_[21176]_  = ~\new_[28981]_  & ~\new_[24331]_ ;
  assign \new_[21177]_  = ~\new_[29568]_  & ~\new_[24390]_ ;
  assign \new_[21178]_  = ~\new_[29069]_  & ~\new_[24157]_ ;
  assign \new_[21179]_  = ~\new_[31429]_  | ~\new_[28266]_  | ~\new_[29902]_ ;
  assign \new_[21180]_  = ~\new_[22213]_ ;
  assign \new_[21181]_  = ~\new_[24347]_  | ~\new_[30728]_ ;
  assign \new_[21182]_  = ~\new_[22225]_ ;
  assign \new_[21183]_  = ~\new_[22228]_ ;
  assign \new_[21184]_  = ~\new_[24464]_  | ~\new_[29569]_ ;
  assign \new_[21185]_  = ~\new_[22233]_ ;
  assign \new_[21186]_  = ~\new_[22237]_ ;
  assign \new_[21187]_  = ~\new_[24434]_  | ~\new_[27721]_ ;
  assign \new_[21188]_  = ~\new_[22239]_ ;
  assign \new_[21189]_  = ~\new_[29195]_  & ~\new_[6036]_ ;
  assign \new_[21190]_  = \new_[27593]_  & \new_[29064]_ ;
  assign \new_[21191]_  = ~\new_[28801]_  & ~\new_[24303]_ ;
  assign \new_[21192]_  = ~\new_[23086]_  | ~\new_[29681]_ ;
  assign \new_[21193]_  = ~\new_[22256]_ ;
  assign \new_[21194]_  = ~\new_[22258]_ ;
  assign \new_[21195]_  = ~\new_[6081]_  | ~\new_[26977]_  | ~\new_[30400]_ ;
  assign \new_[21196]_  = ~\new_[30064]_  & ~\new_[24292]_ ;
  assign \new_[21197]_  = ~\new_[22271]_ ;
  assign \new_[21198]_  = ~\new_[24193]_  & ~\new_[30075]_ ;
  assign \new_[21199]_  = ~\new_[29540]_  & ~\new_[24460]_ ;
  assign \new_[21200]_  = ~\new_[24329]_  | ~\new_[30149]_ ;
  assign \new_[21201]_  = ~\new_[5930]_  | ~\new_[30437]_  | ~\new_[29927]_ ;
  assign \new_[21202]_  = \new_[23173]_  | \new_[28402]_ ;
  assign \new_[21203]_  = \new_[27691]_  & \new_[28535]_ ;
  assign \new_[21204]_  = ~\new_[23245]_  & ~\new_[30188]_ ;
  assign \new_[21205]_  = ~\new_[22304]_ ;
  assign \new_[21206]_  = ~\new_[24412]_  | ~\new_[30321]_ ;
  assign \new_[21207]_  = ~\new_[22305]_ ;
  assign \new_[21208]_  = ~\new_[28447]_  & ~\new_[29629]_ ;
  assign \new_[21209]_  = ~\new_[22308]_ ;
  assign \new_[21210]_  = ~\new_[24265]_  | ~\new_[27353]_ ;
  assign \new_[21211]_  = ~\new_[28444]_  & ~\new_[29174]_ ;
  assign \new_[21212]_  = ~\new_[5992]_  | ~\new_[29085]_  | ~\new_[30438]_ ;
  assign \new_[21213]_  = ~\new_[22323]_ ;
  assign \new_[21214]_  = ~\new_[28393]_  & ~\new_[24264]_ ;
  assign \new_[21215]_  = ~\new_[23168]_  | ~\new_[27489]_ ;
  assign \new_[21216]_  = ~\new_[22331]_ ;
  assign \new_[21217]_  = ~\new_[22333]_ ;
  assign \new_[21218]_  = ~\new_[31870]_  | ~\new_[24782]_  | ~\new_[29593]_ ;
  assign \new_[21219]_  = ~\new_[24193]_  & ~\new_[30837]_ ;
  assign \new_[21220]_  = ~\new_[31423]_  | ~\new_[28266]_  | ~\new_[29902]_ ;
  assign \new_[21221]_  = ~\new_[22335]_ ;
  assign \new_[21222]_  = ~\new_[22341]_ ;
  assign \new_[21223]_  = ~\new_[27604]_  & ~\new_[30649]_ ;
  assign \new_[21224]_  = ~\new_[23999]_  | ~\new_[26953]_ ;
  assign \new_[21225]_  = ~\new_[31928]_  | ~\new_[26940]_  | ~\new_[26655]_ ;
  assign \new_[21226]_  = ~\new_[29398]_  & ~\new_[24452]_ ;
  assign \new_[21227]_  = ~\new_[24500]_  | ~\new_[29893]_ ;
  assign \new_[21228]_  = ~\new_[31616]_  | ~\new_[26292]_  | ~\new_[29969]_ ;
  assign \new_[21229]_  = ~\new_[22360]_ ;
  assign \new_[21230]_  = ~\new_[24380]_  | ~\new_[27553]_ ;
  assign \new_[21231]_  = ~\new_[6077]_  | ~\new_[29265]_  | ~\new_[29272]_ ;
  assign \new_[21232]_  = ~\new_[22375]_ ;
  assign \new_[21233]_  = ~\new_[28966]_  & ~\new_[23081]_ ;
  assign \new_[21234]_  = ~\new_[24440]_  | ~\new_[28898]_ ;
  assign \new_[21235]_  = ~\new_[29277]_  | ~\new_[5999]_ ;
  assign \new_[21236]_  = ~\new_[28067]_  & ~\new_[24470]_ ;
  assign \new_[21237]_  = ~\new_[31799]_  | ~\new_[27546]_  | ~\new_[30735]_ ;
  assign \new_[21238]_  = ~\new_[23547]_  & ~\new_[30010]_ ;
  assign \new_[21239]_  = ~\new_[22408]_ ;
  assign \new_[21240]_  = ~\new_[24295]_  | ~\new_[28828]_ ;
  assign \new_[21241]_  = ~\new_[22411]_ ;
  assign \new_[21242]_  = ~\new_[24256]_  | ~\new_[29441]_ ;
  assign \new_[21243]_  = ~\new_[22413]_ ;
  assign \new_[21244]_  = ~\new_[22413]_ ;
  assign \new_[21245]_  = ~\new_[22413]_ ;
  assign \new_[21246]_  = ~\new_[27505]_  & ~\new_[29445]_ ;
  assign \new_[21247]_  = ~\new_[24330]_  | ~\new_[30009]_ ;
  assign \new_[21248]_  = ~\new_[23145]_  | ~\new_[30142]_ ;
  assign \new_[21249]_  = ~\new_[6185]_  | ~\new_[29373]_  | ~\new_[30055]_ ;
  assign \new_[21250]_  = ~\new_[32313]_ ;
  assign \new_[21251]_  = ~\new_[24544]_  & ~\new_[29671]_ ;
  assign \new_[21252]_  = ~\new_[22434]_ ;
  assign \new_[21253]_  = ~\new_[29660]_  & ~\new_[24525]_ ;
  assign \new_[21254]_  = ~\new_[22437]_ ;
  assign \new_[21255]_  = ~\new_[24448]_  | ~\new_[27526]_ ;
  assign \new_[21256]_  = ~\new_[5932]_  | ~\new_[30025]_  | ~\new_[28371]_ ;
  assign \new_[21257]_  = ~\new_[22450]_ ;
  assign \new_[21258]_  = ~\new_[31232]_  | ~\new_[28266]_  | ~\new_[29902]_ ;
  assign \new_[21259]_  = ~\new_[24274]_  | ~\new_[28993]_ ;
  assign \new_[21260]_  = ~\new_[22457]_ ;
  assign \new_[21261]_  = \new_[28366]_  & \new_[5913]_ ;
  assign \new_[21262]_  = ~\new_[5964]_  | ~\new_[28010]_  | ~\new_[30332]_ ;
  assign \new_[21263]_  = ~\new_[5913]_  | ~\new_[28753]_  | ~\new_[30327]_ ;
  assign \new_[21264]_  = ~\new_[6246]_  | ~\new_[28042]_  | ~\new_[29880]_ ;
  assign \new_[21265]_  = ~\new_[6246]_  | ~\new_[28002]_  | ~\new_[30541]_ ;
  assign \new_[21266]_  = ~\new_[5909]_  | ~\new_[28908]_  | ~\new_[29527]_ ;
  assign \new_[21267]_  = ~\new_[24368]_  | ~\new_[27595]_ ;
  assign \new_[21268]_  = ~\new_[6176]_  | ~\new_[28279]_  | ~\new_[30420]_ ;
  assign \new_[21269]_  = ~\new_[5912]_  | ~\new_[28968]_  | ~\new_[29228]_ ;
  assign \new_[21270]_  = ~\new_[24514]_  | ~\new_[27592]_ ;
  assign \new_[21271]_  = ~\new_[26782]_  | ~\new_[26790]_ ;
  assign \new_[21272]_  = ~\new_[6190]_  | ~\new_[28751]_  | ~\new_[30129]_ ;
  assign \new_[21273]_  = ~\new_[27571]_  & ~\new_[23154]_ ;
  assign \new_[21274]_  = ~\new_[5918]_  | ~\new_[29633]_  | ~\new_[29721]_ ;
  assign \new_[21275]_  = ~\new_[5914]_  | ~\new_[28835]_  | ~\new_[29103]_ ;
  assign \new_[21276]_  = ~\new_[24333]_  | ~\new_[26329]_ ;
  assign \new_[21277]_  = ~\new_[6031]_  | ~\new_[30194]_  | ~\new_[30733]_ ;
  assign \new_[21278]_  = ~\new_[26604]_  & ~\new_[23403]_ ;
  assign \new_[21279]_  = ~\new_[6071]_  | ~\new_[30110]_  | ~\new_[30291]_ ;
  assign \new_[21280]_  = ~\new_[5996]_  | ~\new_[30156]_  | ~\new_[30466]_ ;
  assign \new_[21281]_  = ~\new_[6204]_  | ~\new_[29091]_  | ~\new_[30648]_ ;
  assign \new_[21282]_  = ~\new_[5979]_  | ~\new_[28161]_  | ~\new_[29854]_ ;
  assign \new_[21283]_  = ~\new_[31176]_  | ~\new_[28071]_  | ~\new_[30718]_ ;
  assign \new_[21284]_  = ~\new_[24363]_  & ~\new_[23185]_ ;
  assign \new_[21285]_  = ~\new_[27700]_  & ~\new_[23102]_ ;
  assign \new_[21286]_  = ~\new_[27629]_  & ~\new_[23456]_ ;
  assign \new_[21287]_  = \new_[24196]_  | \new_[29986]_ ;
  assign \new_[21288]_  = ~\new_[5981]_  | ~\new_[29786]_  | ~\new_[29965]_ ;
  assign \new_[21289]_  = ~\new_[6064]_  | ~\new_[30045]_  | ~\new_[30235]_ ;
  assign \new_[21290]_  = ~\new_[5921]_  | ~\new_[28864]_  | ~\new_[29006]_ ;
  assign \new_[21291]_  = ~\new_[23517]_  & (~\new_[30846]_  | ~\new_[6076]_ );
  assign \new_[21292]_  = ~\new_[5917]_  | ~\new_[28911]_  | ~\new_[28963]_ ;
  assign \new_[21293]_  = ~\new_[5919]_  | ~\new_[28951]_  | ~\new_[30101]_ ;
  assign \new_[21294]_  = ~\new_[23131]_  | ~\new_[24699]_ ;
  assign \new_[21295]_  = ~\new_[26591]_  | ~\new_[28490]_ ;
  assign \new_[21296]_  = ~\new_[5985]_  | ~\new_[28040]_  | ~\new_[30413]_ ;
  assign \new_[21297]_  = ~\new_[23136]_  & (~\new_[28595]_  | ~\new_[5988]_ );
  assign \new_[21298]_  = \new_[24426]_  | \new_[30122]_ ;
  assign \new_[21299]_  = ~\new_[30848]_  | ~\new_[29121]_  | ~\new_[30553]_ ;
  assign \new_[21300]_  = ~\new_[23163]_  & (~\new_[28278]_  | ~\new_[6189]_ );
  assign \new_[21301]_  = ~\new_[24459]_  | ~\new_[27465]_ ;
  assign \new_[21302]_  = ~\new_[5911]_  | ~\new_[29112]_  | ~\new_[29320]_ ;
  assign \new_[21303]_  = ~\new_[5994]_  | ~\new_[28932]_  | ~\new_[29809]_ ;
  assign \new_[21304]_  = ~\new_[5930]_  | ~\new_[29622]_  | ~\new_[29915]_ ;
  assign \new_[21305]_  = ~\new_[5983]_  | ~\new_[28633]_  | ~\new_[30176]_ ;
  assign \new_[21306]_  = ~\new_[5991]_  | ~\new_[28243]_  | ~\new_[30788]_ ;
  assign \new_[21307]_  = ~\new_[6269]_  | ~\new_[28679]_  | ~\new_[30737]_ ;
  assign \new_[21308]_  = ~\new_[27718]_  | ~\new_[28508]_ ;
  assign \new_[21309]_  = ~\new_[27628]_  & ~\new_[24505]_ ;
  assign \new_[21310]_  = ~\new_[5923]_  | ~\new_[28844]_  | ~\new_[29695]_ ;
  assign \new_[21311]_  = ~\new_[23110]_  & (~\new_[28675]_  | ~\new_[6185]_ );
  assign \new_[21312]_  = ~\new_[6059]_  | ~\new_[27981]_  | ~\new_[30250]_ ;
  assign \new_[21313]_  = ~\new_[31132]_  | ~\new_[29078]_  | ~\new_[30502]_ ;
  assign \new_[21314]_  = ~\new_[24466]_  | ~\new_[26236]_ ;
  assign \new_[21315]_  = ~\new_[24289]_  | ~\new_[27791]_ ;
  assign \new_[21316]_  = ~\new_[28162]_  & ~\new_[24474]_ ;
  assign \new_[21317]_  = ~\new_[27748]_  | ~\new_[28538]_ ;
  assign \new_[21318]_  = ~\new_[6001]_  | ~\new_[27996]_  | ~\new_[30652]_ ;
  assign \new_[21319]_  = ~\new_[5999]_  | ~\new_[28282]_  | ~\new_[29918]_ ;
  assign \new_[21320]_  = ~\new_[5997]_  | ~\new_[28345]_  | ~\new_[30315]_ ;
  assign \new_[21321]_  = ~\new_[27731]_  | ~\new_[26812]_ ;
  assign \new_[21322]_  = ~\new_[5926]_  | ~\new_[24547]_  | ~\new_[30032]_ ;
  assign \new_[21323]_  = ~\new_[5927]_  | ~\new_[29189]_  | ~\new_[29456]_ ;
  assign \new_[21324]_  = ~\new_[24523]_  | ~\new_[26241]_ ;
  assign \new_[21325]_  = ~\new_[31763]_  | ~\new_[28652]_  | ~\new_[29774]_ ;
  assign \new_[21326]_  = ~\new_[27375]_  | ~\new_[28049]_ ;
  assign \new_[21327]_  = ~\new_[5932]_  | ~\new_[28262]_  | ~\new_[29789]_ ;
  assign \new_[21328]_  = ~\new_[6007]_  | ~\new_[28717]_  | ~\new_[30706]_ ;
  assign \new_[21329]_  = ~\new_[24388]_  & (~\new_[30694]_  | ~\new_[30513]_ );
  assign \new_[21330]_  = ~\new_[24453]_  & (~\new_[30575]_  | ~\new_[30678]_ );
  assign \new_[21331]_  = ~\new_[24106]_  & (~\new_[28685]_  | ~\new_[30222]_ );
  assign \new_[21332]_  = ~\new_[24318]_  & (~\new_[30701]_  | ~\new_[30467]_ );
  assign \new_[21333]_  = ~\new_[23115]_  & (~\new_[28960]_  | ~\new_[29869]_ );
  assign \new_[21334]_  = ~\new_[23181]_  & (~\new_[30837]_  | ~\new_[30846]_ );
  assign \new_[21335]_  = ~\new_[24291]_  & (~\new_[29315]_  | ~\new_[30525]_ );
  assign \new_[21336]_  = ~\new_[24334]_  & (~\new_[30068]_  | ~\new_[29868]_ );
  assign \new_[21337]_  = ~\new_[23105]_  & (~\new_[28686]_  | ~\new_[30229]_ );
  assign \new_[21338]_  = ~\new_[24435]_  & (~\new_[29165]_  | ~\new_[29851]_ );
  assign \new_[21339]_  = ~\new_[23144]_  & (~\new_[30543]_  | ~\new_[30571]_ );
  assign \new_[21340]_  = ~\new_[23123]_  & (~\new_[28076]_  | ~\new_[29987]_ );
  assign \new_[21341]_  = ~\new_[24149]_  & (~\new_[30661]_  | ~\new_[30494]_ );
  assign \new_[21342]_  = ~\new_[30240]_  | ~\new_[5990]_ ;
  assign \new_[21343]_  = ~\new_[24363]_  | ~\new_[29701]_ ;
  assign \new_[21344]_  = ~\new_[28840]_  & ~\new_[5972]_ ;
  assign \new_[21345]_  = ~\new_[30247]_  | ~\new_[6195]_ ;
  assign \new_[21346]_  = ~\new_[29776]_  | ~\new_[6052]_ ;
  assign \new_[21347]_  = \new_[29159]_  | \new_[31617]_ ;
  assign \new_[21348]_  = ~\new_[29545]_  | ~\new_[6192]_ ;
  assign \new_[21349]_  = ~\new_[23952]_  & ~\new_[30656]_ ;
  assign \new_[21350]_  = ~\new_[29501]_  | ~\new_[6044]_ ;
  assign \new_[21351]_  = ~\new_[29398]_  | ~\new_[6081]_ ;
  assign \new_[21352]_  = ~\new_[29885]_  | ~\new_[6005]_ ;
  assign \new_[21353]_  = ~\new_[29306]_  | ~\new_[6046]_ ;
  assign \new_[21354]_  = ~\new_[30289]_  | ~\new_[6046]_ ;
  assign \new_[21355]_  = ~\new_[29306]_  | ~\new_[31143]_ ;
  assign \new_[21356]_  = ~\new_[30141]_  | ~\new_[5918]_ ;
  assign \new_[21357]_  = \new_[28337]_  | \new_[31819]_ ;
  assign \new_[21358]_  = ~\new_[30340]_  | ~\new_[31406]_ ;
  assign \new_[21359]_  = ~\new_[28270]_  | ~\new_[5964]_ ;
  assign \new_[21360]_  = ~\new_[28270]_  | ~\new_[5963]_ ;
  assign \new_[21361]_  = ~\new_[30209]_  | ~\new_[6064]_ ;
  assign \new_[21362]_  = ~\new_[28285]_  & ~\new_[30874]_ ;
  assign \new_[21363]_  = ~\new_[30209]_  | ~\new_[6273]_ ;
  assign \new_[21364]_  = ~\new_[28873]_  | ~\new_[5992]_ ;
  assign \new_[21365]_  = ~\new_[28293]_  | ~\new_[6088]_ ;
  assign \new_[21366]_  = ~\new_[29970]_  | ~\new_[6001]_ ;
  assign \new_[21367]_  = ~\new_[29776]_  | ~\new_[6053]_ ;
  assign \new_[21368]_  = ~\new_[29597]_  | ~\new_[5965]_ ;
  assign \new_[21369]_  = ~\new_[29672]_  | ~\new_[6088]_ ;
  assign \new_[21370]_  = ~\new_[29360]_  | ~\new_[6048]_ ;
  assign \new_[21371]_  = ~\new_[30209]_  | ~\new_[6065]_ ;
  assign \new_[21372]_  = ~\new_[28012]_  | ~\new_[5982]_ ;
  assign \new_[21373]_  = ~\new_[26657]_  | ~\new_[5971]_ ;
  assign \new_[21374]_  = ~\new_[28610]_  | ~\new_[5990]_ ;
  assign \new_[21375]_  = \new_[29750]_  & \new_[31406]_ ;
  assign \new_[21376]_  = ~\new_[29122]_  | ~\new_[6052]_ ;
  assign \new_[21377]_  = ~\new_[28366]_  | ~\new_[5971]_ ;
  assign \new_[21378]_  = ~\new_[26657]_  | ~\new_[6047]_ ;
  assign \new_[21379]_  = ~\new_[29019]_  | ~\new_[6046]_ ;
  assign \new_[21380]_  = ~\new_[28966]_  | ~\new_[6058]_ ;
  assign \new_[21381]_  = ~\new_[29956]_  | ~\new_[6217]_ ;
  assign \new_[21382]_  = ~\new_[28830]_  | ~\new_[6217]_ ;
  assign \new_[21383]_  = ~\new_[29019]_  | ~\new_[31143]_ ;
  assign \new_[21384]_  = ~\new_[29776]_  | ~\new_[6031]_ ;
  assign \new_[21385]_  = ~\new_[29184]_  | ~\new_[6090]_ ;
  assign \new_[21386]_  = ~\new_[30331]_  | ~\new_[31033]_ ;
  assign \new_[21387]_  = ~\new_[30266]_  | ~\new_[5973]_ ;
  assign \new_[21388]_  = \new_[29184]_  & \new_[31132]_ ;
  assign \new_[21389]_  = \new_[28012]_  & \new_[5981]_ ;
  assign \new_[21390]_  = ~\new_[29256]_  | ~\new_[5980]_ ;
  assign \new_[21391]_  = ~\new_[28966]_  | ~\new_[5980]_ ;
  assign \new_[21392]_  = ~\new_[29277]_  | ~\new_[6185]_ ;
  assign \new_[21393]_  = ~\new_[28682]_  | ~\new_[5986]_ ;
  assign \new_[21394]_  = ~\new_[28834]_  | ~\new_[6052]_ ;
  assign \new_[21395]_  = \new_[28293]_  & \new_[5931]_ ;
  assign \new_[21396]_  = ~\new_[29122]_  | ~\new_[6053]_ ;
  assign \new_[21397]_  = ~\new_[29071]_  | ~\new_[6065]_ ;
  assign \new_[21398]_  = ~\new_[30224]_  | ~\new_[31491]_ ;
  assign \new_[21399]_  = ~\new_[30247]_  | ~\new_[6059]_ ;
  assign \new_[21400]_  = ~\new_[29360]_  | ~\new_[6200]_ ;
  assign \new_[21401]_  = ~\new_[29169]_  | ~\new_[31033]_ ;
  assign \new_[21402]_  = ~\new_[30014]_  | ~\new_[5987]_ ;
  assign \new_[21403]_  = ~\new_[28211]_  | ~\new_[5990]_ ;
  assign \new_[21404]_  = ~\new_[29736]_  | ~\new_[5969]_ ;
  assign \new_[21405]_  = ~\new_[30004]_  | ~\new_[5965]_ ;
  assign \new_[21406]_  = ~\new_[28211]_  | ~\new_[6190]_ ;
  assign \new_[21407]_  = ~\new_[30173]_  | ~\new_[5986]_ ;
  assign \new_[21408]_  = ~\new_[30340]_  | ~\new_[31121]_ ;
  assign \new_[21409]_  = ~\new_[29995]_  | ~\new_[6000]_ ;
  assign \new_[21410]_  = ~\new_[30244]_  | ~\new_[6085]_ ;
  assign \new_[21411]_  = ~\new_[29799]_  | ~\new_[5998]_ ;
  assign \new_[21412]_  = ~\new_[30004]_  | ~\new_[6039]_ ;
  assign \new_[21413]_  = ~\new_[29597]_  | ~\new_[6039]_ ;
  assign \new_[21414]_  = ~\new_[30247]_  | ~\new_[6060]_ ;
  assign \new_[21415]_  = ~\new_[28234]_  | ~\new_[5993]_ ;
  assign \new_[21416]_  = ~\new_[29758]_  | ~\new_[6088]_ ;
  assign \new_[21417]_  = \new_[28234]_  & \new_[5994]_ ;
  assign \new_[21418]_  = ~\new_[29791]_  | ~\new_[5980]_ ;
  assign \new_[21419]_  = ~\new_[28873]_  | ~\new_[5922]_ ;
  assign \new_[21420]_  = ~\new_[30407]_  | ~\new_[5980]_ ;
  assign \new_[21421]_  = ~\new_[30323]_  | ~\new_[31235]_ ;
  assign \new_[21422]_  = ~\new_[29970]_  | ~\new_[5929]_ ;
  assign \new_[21423]_  = ~\new_[28337]_  & ~\new_[31787]_ ;
  assign \new_[21424]_  = ~\new_[30331]_  | ~\new_[31235]_ ;
  assign \new_[21425]_  = ~\new_[30342]_  | ~\new_[6065]_ ;
  assign \new_[21426]_  = ~\new_[28966]_  | ~\new_[5979]_ ;
  assign \new_[21427]_  = ~\new_[30224]_  | ~\new_[31121]_ ;
  assign \new_[21428]_  = ~\new_[29826]_  | ~\new_[5965]_ ;
  assign \new_[21429]_  = ~\new_[29501]_  | ~\new_[5969]_ ;
  assign \new_[21430]_  = ~\new_[29722]_  | ~\new_[6245]_ ;
  assign \new_[21431]_  = ~\new_[29266]_  | ~\new_[5929]_ ;
  assign \new_[21432]_  = ~\new_[28211]_  | ~\new_[6189]_ ;
  assign \new_[21433]_  = \new_[28830]_  & \new_[6007]_ ;
  assign \new_[21434]_  = ~\new_[29758]_  | ~\new_[6003]_ ;
  assign \new_[21435]_  = ~\new_[29956]_  | ~\new_[6095]_ ;
  assign \new_[21436]_  = ~\new_[28409]_  | ~\new_[5963]_ ;
  assign \new_[21437]_  = ~\new_[28250]_  | ~\new_[5963]_ ;
  assign \new_[21438]_  = \new_[28250]_  & \new_[5964]_ ;
  assign \new_[21439]_  = ~\new_[30036]_  | ~\new_[5929]_ ;
  assign \new_[21440]_  = ~\new_[29398]_  | ~\new_[5998]_ ;
  assign \new_[21441]_  = ~\new_[29613]_  | ~\new_[6000]_ ;
  assign \new_[21442]_  = ~\new_[29347]_  | ~\new_[6048]_ ;
  assign \new_[21443]_  = ~\new_[29277]_  | ~\new_[6000]_ ;
  assign \new_[21444]_  = ~\new_[29970]_  | ~\new_[6086]_ ;
  assign \new_[21445]_  = ~\new_[28977]_  | ~\new_[5922]_ ;
  assign \new_[21446]_  = \new_[28610]_  & \new_[6190]_ ;
  assign \new_[21447]_  = ~\new_[30323]_  | ~\new_[31394]_ ;
  assign \new_[21448]_  = ~\new_[28891]_  | ~\new_[5995]_ ;
  assign \new_[21449]_  = ~\new_[30266]_  | ~\new_[5972]_ ;
  assign \new_[21450]_  = ~\new_[29398]_  | ~\new_[5997]_ ;
  assign \new_[21451]_  = ~\new_[30323]_  | ~\new_[31033]_ ;
  assign \new_[21452]_  = ~\new_[29827]_  | ~\new_[5971]_ ;
  assign \new_[21453]_  = ~\new_[29672]_  | ~\new_[6003]_ ;
  assign \new_[21454]_  = ~\new_[29383]_  | ~\new_[6005]_ ;
  assign \new_[21455]_  = ~\new_[30633]_  | ~\new_[6043]_ ;
  assign \new_[21456]_  = ~\new_[29062]_  | ~\new_[31423]_ ;
  assign \new_[21457]_  = ~\new_[30607]_  | ~\new_[6092]_ ;
  assign \new_[21458]_  = ~\new_[24759]_  | ~\new_[5989]_ ;
  assign \new_[21459]_  = ~\new_[30319]_  | ~\new_[6067]_ ;
  assign \new_[21460]_  = ~\new_[29648]_  | ~\new_[6074]_ ;
  assign \new_[21461]_  = ~\new_[29227]_  & ~\new_[6067]_ ;
  assign \new_[21462]_  = ~\new_[24759]_  | ~\new_[6072]_ ;
  assign \new_[21463]_  = ~\new_[28979]_  | ~\new_[6056]_ ;
  assign \new_[21464]_  = ~\new_[30616]_  | ~\new_[6050]_ ;
  assign \new_[21465]_  = ~\new_[22875]_ ;
  assign \new_[21466]_  = ~\new_[26563]_  | ~\new_[6043]_ ;
  assign \new_[21467]_  = ~\new_[29174]_  | ~\new_[5901]_ ;
  assign \new_[21468]_  = ~\new_[28278]_  | ~\new_[30034]_ ;
  assign \new_[21469]_  = ~\new_[22887]_ ;
  assign \new_[21470]_  = ~\new_[27883]_  | ~\new_[30763]_ ;
  assign \new_[21471]_  = ~\new_[30389]_  | ~\new_[6045]_ ;
  assign \new_[21472]_  = ~\new_[29565]_  & ~\new_[30076]_ ;
  assign \new_[21473]_  = ~\new_[28878]_  & ~\new_[5993]_ ;
  assign \new_[21474]_  = ~\new_[28889]_  & ~\new_[6000]_ ;
  assign \new_[21475]_  = ~\new_[29765]_  & ~\new_[30192]_ ;
  assign \new_[21476]_  = ~\new_[30192]_  | ~\new_[6045]_ ;
  assign \new_[21477]_  = ~\new_[26563]_  | ~\new_[5967]_ ;
  assign \new_[21478]_  = ~\new_[29681]_  | ~\new_[29974]_ ;
  assign \new_[21479]_  = ~\new_[29217]_  | ~\new_[6045]_ ;
  assign \new_[21480]_  = ~\new_[29825]_  | ~\new_[30702]_ ;
  assign \new_[21481]_  = ~\new_[28933]_  | ~\new_[5894]_ ;
  assign \new_[21482]_  = ~\new_[28833]_  & ~\new_[6045]_ ;
  assign \new_[21483]_  = ~\new_[28270]_  | ~\new_[6035]_ ;
  assign \new_[21484]_  = ~\new_[29047]_  | ~\new_[6087]_ ;
  assign \new_[21485]_  = ~\new_[30052]_  | ~\new_[6067]_ ;
  assign \new_[21486]_  = ~\new_[28865]_  | ~\new_[30279]_ ;
  assign \new_[21487]_  = ~\new_[29056]_  & ~\new_[6083]_ ;
  assign \new_[21488]_  = ~\new_[30273]_  | ~\new_[6192]_ ;
  assign \new_[21489]_  = ~\new_[29541]_  | ~\new_[6042]_ ;
  assign \new_[21490]_  = ~\new_[30334]_  | ~\new_[6042]_ ;
  assign \new_[21491]_  = \new_[30030]_  | \new_[31800]_ ;
  assign \new_[21492]_  = ~\new_[30557]_  | ~\new_[6215]_ ;
  assign \new_[21493]_  = ~\new_[30028]_  | ~\new_[6061]_ ;
  assign \new_[21494]_  = ~\new_[30835]_  | ~\new_[6211]_ ;
  assign \new_[21495]_  = ~\new_[29445]_  | ~\new_[5900]_ ;
  assign \new_[21496]_  = ~\new_[30008]_  | ~\new_[6075]_ ;
  assign \new_[21497]_  = ~\new_[30285]_  | ~\new_[6036]_ ;
  assign \new_[21498]_  = ~\new_[30656]_  | ~\new_[5989]_ ;
  assign \new_[21499]_  = ~\new_[29157]_  | ~\new_[6062]_ ;
  assign \new_[21500]_  = ~\new_[29100]_  | ~\new_[6042]_ ;
  assign \new_[21501]_  = ~\new_[29068]_  & ~\new_[6075]_ ;
  assign \new_[21502]_  = ~\new_[30267]_  & ~\new_[30008]_ ;
  assign \new_[21503]_  = ~\new_[28969]_  & ~\new_[5971]_ ;
  assign \new_[21504]_  = ~\new_[29100]_  & ~\new_[30314]_ ;
  assign \new_[21505]_  = ~\new_[30633]_  | ~\new_[5967]_ ;
  assign \new_[21506]_  = ~\new_[23077]_ ;
  assign \new_[21507]_  = ~\new_[30268]_  & ~\new_[30249]_ ;
  assign \new_[21508]_  = ~\new_[29914]_  & ~\new_[30319]_ ;
  assign \new_[21509]_  = ~\new_[23074]_ ;
  assign \new_[21510]_  = ~\new_[29175]_  & ~\new_[5920]_ ;
  assign \new_[21511]_  = ~\new_[29745]_  | ~\new_[6087]_ ;
  assign \new_[21512]_  = ~\new_[30578]_  | ~\new_[29324]_ ;
  assign \new_[21513]_  = ~\new_[29394]_  & ~\new_[6042]_ ;
  assign \new_[21514]_  = ~\new_[29748]_  | ~\new_[5894]_ ;
  assign \new_[21515]_  = ~\new_[30272]_  | ~\new_[6083]_ ;
  assign \new_[21516]_  = ~\new_[29777]_  & ~\new_[29181]_ ;
  assign \new_[21517]_  = ~\new_[29086]_  & ~\new_[5986]_ ;
  assign \new_[21518]_  = ~\new_[30024]_  & ~\new_[30272]_ ;
  assign \new_[21519]_  = ~\new_[29934]_  | ~\new_[6074]_ ;
  assign \new_[21520]_  = ~\new_[30174]_  & ~\new_[26842]_ ;
  assign \new_[21521]_  = ~\new_[29745]_  | ~\new_[5907]_ ;
  assign \new_[21522]_  = ~\new_[30141]_  | ~\new_[6193]_ ;
  assign \new_[21523]_  = ~\new_[29700]_  | ~\new_[6056]_ ;
  assign \new_[21524]_  = ~\new_[29652]_  | ~\new_[5933]_ ;
  assign \new_[21525]_  = ~\new_[29354]_  | ~\new_[6091]_ ;
  assign \new_[21526]_  = ~\new_[30348]_  | ~\new_[6069]_ ;
  assign \new_[21527]_  = ~\new_[30277]_  & ~\new_[29652]_ ;
  assign \new_[21528]_  = ~\new_[29855]_  | ~\new_[6036]_ ;
  assign \new_[21529]_  = ~\new_[29167]_  | ~\new_[6083]_ ;
  assign \new_[21530]_  = ~\new_[30355]_  | ~\new_[31423]_ ;
  assign \new_[21531]_  = ~\new_[28675]_  | ~\new_[28007]_ ;
  assign \new_[21532]_  = ~\new_[29172]_  | ~\new_[6202]_ ;
  assign \new_[21533]_  = ~\new_[30062]_  & ~\new_[29934]_ ;
  assign \new_[21534]_  = ~\new_[29882]_  | ~\new_[5927]_ ;
  assign \new_[21535]_  = ~\new_[30245]_  & ~\new_[30285]_ ;
  assign \new_[21536]_  = ~\new_[30044]_  | ~\new_[31423]_ ;
  assign \new_[21537]_  = ~\new_[29465]_  & ~\new_[6051]_ ;
  assign \new_[21538]_  = ~\new_[22496]_ ;
  assign \new_[21539]_  = ~\new_[29814]_  | ~\new_[5914]_ ;
  assign \new_[21540]_  = ~\new_[29908]_  & ~\new_[30334]_ ;
  assign \new_[21541]_  = ~\new_[29898]_  & ~\new_[29882]_ ;
  assign \new_[21542]_  = ~\new_[30348]_  | ~\new_[6070]_ ;
  assign \new_[21543]_  = ~\new_[29814]_  | ~\new_[6051]_ ;
  assign \new_[21544]_  = ~\new_[30042]_  & ~\new_[28933]_ ;
  assign \new_[21545]_  = ~\new_[29768]_  | ~\new_[29118]_ ;
  assign \new_[21546]_  = ~\new_[29648]_  & ~\new_[30127]_ ;
  assign \new_[21547]_  = ~\new_[30423]_  & ~\new_[26638]_ ;
  assign \new_[21548]_  = ~\new_[30348]_  | ~\new_[31400]_ ;
  assign \new_[21549]_  = ~\new_[29101]_  | ~\new_[6074]_ ;
  assign \new_[21550]_  = ~\new_[29663]_  & ~\new_[6074]_ ;
  assign \new_[21551]_  = ~\new_[30069]_  | ~\new_[6193]_ ;
  assign \new_[21552]_  = ~\new_[30052]_  | ~\new_[5917]_ ;
  assign \new_[21553]_  = ~\new_[29898]_  | ~\new_[6083]_ ;
  assign \new_[21554]_  = ~\new_[29578]_  & ~\new_[6193]_ ;
  assign \new_[21555]_  = ~\new_[29748]_  | ~\new_[6202]_ ;
  assign \new_[21556]_  = ~\new_[28595]_  | ~\new_[29355]_ ;
  assign \new_[21557]_  = \new_[23351]_  & \new_[28475]_ ;
  assign \new_[21558]_  = ~\new_[22982]_ ;
  assign \new_[21559]_  = ~\new_[24413]_  & ~\new_[29930]_ ;
  assign \new_[21560]_  = ~\new_[30703]_  & ~\new_[30028]_ ;
  assign \new_[21561]_  = ~\new_[26387]_  | ~\new_[30386]_ ;
  assign \new_[21562]_  = ~\new_[24721]_  | ~\new_[29975]_ ;
  assign \new_[21563]_  = ~\new_[24374]_ ;
  assign \new_[21564]_  = ~\new_[30598]_  | ~\new_[6034]_ ;
  assign \new_[21565]_  = ~\new_[23080]_ ;
  assign \new_[21566]_  = ~\new_[29891]_  & ~\new_[5987]_ ;
  assign \new_[21567]_  = ~\new_[28004]_  | ~\new_[6036]_ ;
  assign \new_[21568]_  = ~\new_[30708]_  | ~\new_[6093]_ ;
  assign \new_[21569]_  = ~\new_[23090]_ ;
  assign \new_[21570]_  = ~\new_[30755]_  | ~\new_[6184]_ ;
  assign \new_[21571]_  = ~\new_[24759]_  & ~\new_[6073]_ ;
  assign \new_[21572]_  = ~\new_[30326]_  | ~\new_[5984]_ ;
  assign \new_[21573]_  = ~\new_[30032]_  | ~\new_[5933]_ ;
  assign \new_[21574]_  = ~\new_[30234]_  | ~\new_[5900]_ ;
  assign \new_[21575]_  = ~\new_[29922]_  & ~\new_[6052]_ ;
  assign \new_[21576]_  = ~\new_[5978]_  | ~\new_[30005]_  | ~\new_[29441]_ ;
  assign \new_[21577]_  = (~\new_[27855]_  | ~\s4_data_i[8] ) & (~\new_[27879]_  | ~\s0_data_i[8] );
  assign \new_[21578]_  = ~\new_[29774]_  | ~\new_[6091]_ ;
  assign \new_[21579]_  = (~\new_[30106]_  | ~\s14_data_i[0] ) & (~\new_[27347]_  | ~\s12_data_i[0] );
  assign \new_[21580]_  = ~\new_[6084]_  | ~\new_[30089]_  | ~\new_[30142]_ ;
  assign \new_[21581]_  = (~\new_[27855]_  | ~\s4_data_i[20] ) & (~\new_[27879]_  | ~\s0_data_i[20] );
  assign \new_[21582]_  = ~\new_[30029]_  | ~\new_[30897]_ ;
  assign \new_[21583]_  = (~\new_[29604]_  | ~\s11_data_i[8] ) & (~\new_[27337]_  | ~\s8_data_i[8] );
  assign \new_[21584]_  = ~\new_[23136]_ ;
  assign \new_[21585]_  = ~\new_[23144]_ ;
  assign \new_[21586]_  = (~\new_[30106]_  | ~\s14_data_i[7] ) & (~\new_[27347]_  | ~\s12_data_i[7] );
  assign \new_[21587]_  = ~\new_[29079]_  & ~\new_[5965]_ ;
  assign \new_[21588]_  = ~\new_[29927]_  | (~\new_[26962]_  & ~\new_[28654]_ );
  assign \new_[21589]_  = ~\new_[30231]_  | ~\new_[6094]_ ;
  assign \new_[21590]_  = ~\new_[28274]_  & ~\new_[24599]_ ;
  assign \new_[21591]_  = ~\new_[24777]_  & ~\new_[25770]_ ;
  assign \new_[21592]_  = ~\new_[29197]_  | ~\new_[30217]_ ;
  assign \new_[21593]_  = ~\new_[6032]_  | ~\new_[30318]_  | ~\new_[29975]_ ;
  assign \new_[21594]_  = \new_[28872]_  | \new_[31903]_ ;
  assign \new_[21595]_  = ~\new_[29162]_  & ~\new_[5982]_ ;
  assign \new_[21596]_  = ~\new_[30086]_  | ~\new_[28641]_  | ~\new_[27513]_ ;
  assign \new_[21597]_  = ~\new_[30845]_  & (~\new_[26681]_  | ~\new_[26875]_ );
  assign \new_[21598]_  = ~\new_[29016]_  & (~\new_[26876]_  | ~\new_[26971]_ );
  assign \new_[21599]_  = ~\new_[28686]_  & (~\new_[27170]_  | ~\new_[26890]_ );
  assign \new_[21600]_  = ~\new_[30076]_  | ~\new_[6075]_ ;
  assign \new_[21601]_  = ~\new_[28950]_  & (~\new_[26996]_  | ~\new_[26812]_ );
  assign \new_[21602]_  = ~\new_[30708]_  | ~\new_[6092]_ ;
  assign \new_[21603]_  = ~\new_[28076]_  & (~\new_[26949]_  | ~\new_[26959]_ );
  assign \new_[21604]_  = ~\new_[30375]_  | ~\new_[6070]_ ;
  assign \new_[21605]_  = ~\new_[26227]_  & (~\new_[26919]_  | ~\new_[29808]_ );
  assign \new_[21606]_  = ~\new_[27600]_  | ~\new_[27264]_  | ~\new_[29600]_ ;
  assign \new_[21607]_  = ~\new_[30275]_  | ~\new_[6072]_ ;
  assign \new_[21608]_  = ~\new_[30276]_  & (~\new_[26986]_  | ~\new_[26970]_ );
  assign \new_[21609]_  = ~\new_[30325]_  | ~\new_[6092]_ ;
  assign \new_[21610]_  = ~\new_[30736]_  & (~\new_[26680]_  | ~\new_[29448]_ );
  assign \new_[21611]_  = ~\new_[30604]_  | ~\new_[30665]_ ;
  assign \new_[21612]_  = ~\new_[30726]_  | (~\new_[26600]_  & ~\new_[26948]_ );
  assign \new_[21613]_  = ~\new_[30425]_  & (~\new_[26618]_  | ~\new_[29026]_ );
  assign \new_[21614]_  = ~\new_[30508]_  | (~\new_[26891]_  & ~\new_[27562]_ );
  assign \new_[21615]_  = (~\new_[29604]_  | ~\s11_data_i[29] ) & (~\new_[27337]_  | ~\s8_data_i[29] );
  assign \new_[21616]_  = ~\new_[30245]_  | ~\new_[5895]_ ;
  assign \new_[21617]_  = ~\new_[30289]_  & (~\new_[26896]_  | ~\new_[29454]_ );
  assign \new_[21618]_  = ~\new_[30336]_  | ~\new_[5970]_ ;
  assign n8764 = m4_s3_cyc_o_reg;
  assign \new_[21620]_  = ~\new_[29997]_  | ~\new_[6084]_ ;
  assign \new_[21621]_  = ~\new_[30438]_  & (~\new_[27547]_  | ~\new_[29460]_ );
  assign \new_[21622]_  = ~\new_[30507]_  | (~\new_[26927]_  & ~\new_[27993]_ );
  assign \new_[21623]_  = ~\new_[30820]_  | (~\new_[27426]_  & ~\new_[29372]_ );
  assign \new_[21624]_  = ~\new_[30276]_  & (~\new_[26970]_  | ~\new_[29464]_ );
  assign \new_[21625]_  = ~\new_[25170]_  & ~\new_[30736]_ ;
  assign \new_[21626]_  = ~\new_[24652]_  & ~\new_[30757]_ ;
  assign \new_[21627]_  = ~\new_[25197]_  & ~\new_[30438]_ ;
  assign \new_[21628]_  = ~\new_[25266]_  & ~\new_[30014]_ ;
  assign \new_[21629]_  = ~\new_[24600]_  & ~\new_[30224]_ ;
  assign \new_[21630]_  = ~\new_[25194]_  & ~\new_[30273]_ ;
  assign \new_[21631]_  = ~\new_[24578]_  & ~\new_[30244]_ ;
  assign \new_[21632]_  = ~\new_[24795]_  | ~\new_[29357]_ ;
  assign \new_[21633]_  = ~\new_[24794]_  & ~\new_[30042]_ ;
  assign \new_[21634]_  = ~\new_[24888]_  & ~\new_[27540]_ ;
  assign \new_[21635]_  = \new_[24796]_  & \new_[28585]_ ;
  assign \new_[21636]_  = \new_[24994]_  | \new_[25116]_ ;
  assign \new_[21637]_  = ~\new_[25116]_  & ~\new_[30540]_ ;
  assign \new_[21638]_  = \new_[24994]_  | \new_[30540]_ ;
  assign \new_[21639]_  = \new_[24790]_  | \new_[30230]_ ;
  assign \new_[21640]_  = ~\new_[25153]_  & ~\new_[30566]_ ;
  assign \new_[21641]_  = ~\new_[24804]_  | ~\new_[24974]_ ;
  assign \new_[21642]_  = ~\new_[24918]_  | ~\new_[27359]_ ;
  assign \new_[21643]_  = ~\new_[24808]_  | ~\new_[24807]_ ;
  assign \new_[21644]_  = ~\new_[24593]_  | ~\new_[29874]_ ;
  assign \new_[21645]_  = ~\new_[24970]_  | ~\new_[30707]_ ;
  assign \new_[21646]_  = \new_[24639]_  & \new_[25310]_ ;
  assign \new_[21647]_  = \new_[25303]_  & \new_[25480]_ ;
  assign \new_[21648]_  = ~\new_[26968]_  | ~\new_[24813]_ ;
  assign \new_[21649]_  = ~\new_[24815]_  | ~\new_[24814]_ ;
  assign \new_[21650]_  = ~\new_[25270]_  & ~\new_[30607]_ ;
  assign \new_[21651]_  = ~\new_[25089]_  & ~\new_[30245]_ ;
  assign \new_[21652]_  = ~\new_[24897]_  | ~\new_[24665]_ ;
  assign \new_[21653]_  = \new_[25088]_  | \new_[25089]_ ;
  assign \new_[21654]_  = ~\new_[25088]_  & ~\new_[30245]_ ;
  assign \new_[21655]_  = ~\new_[24724]_  & ~\new_[30042]_ ;
  assign \new_[21656]_  = ~\new_[24981]_  & ~\new_[30024]_ ;
  assign \new_[21657]_  = \new_[24689]_  | \new_[30047]_ ;
  assign \new_[21658]_  = \new_[25839]_  & \new_[25328]_ ;
  assign \new_[21659]_  = ~\new_[25138]_  & ~\new_[30325]_ ;
  assign \new_[21660]_  = ~\new_[25030]_  | ~\new_[30147]_ ;
  assign \new_[21661]_  = \new_[25334]_  & \new_[26567]_ ;
  assign \new_[21662]_  = ~\new_[25081]_  | ~\new_[26363]_ ;
  assign \new_[21663]_  = ~\new_[24565]_  | ~\new_[26363]_ ;
  assign \new_[21664]_  = \new_[25959]_  & \new_[26327]_ ;
  assign \new_[21665]_  = \new_[25912]_  & \new_[24590]_ ;
  assign \new_[21666]_  = ~\new_[24833]_  | ~\new_[30215]_ ;
  assign \new_[21667]_  = \new_[25054]_  | \new_[30336]_ ;
  assign \new_[21668]_  = \new_[25346]_  & \new_[25924]_ ;
  assign \new_[21669]_  = \new_[25329]_  & \new_[25990]_ ;
  assign \new_[21670]_  = \new_[24835]_  | \new_[27562]_ ;
  assign \new_[21671]_  = \new_[24837]_  | \new_[24838]_ ;
  assign \new_[21672]_  = ~\new_[27170]_  | ~\new_[26344]_ ;
  assign \new_[21673]_  = \new_[26264]_  & \new_[25761]_ ;
  assign \new_[21674]_  = ~\new_[26890]_  | ~\new_[26344]_ ;
  assign \new_[21675]_  = ~\new_[25137]_  & ~\new_[30521]_ ;
  assign \new_[21676]_  = \new_[25354]_  & \new_[25355]_ ;
  assign \new_[21677]_  = ~\new_[25048]_  | ~\new_[26022]_ ;
  assign \new_[21678]_  = \new_[26196]_  & \new_[25363]_ ;
  assign \new_[21679]_  = ~\new_[25023]_  | ~\new_[28541]_ ;
  assign \new_[21680]_  = \new_[25720]_  & \new_[25370]_ ;
  assign \new_[21681]_  = \new_[25372]_  & \new_[25378]_ ;
  assign \new_[21682]_  = \new_[25375]_  & \new_[25697]_ ;
  assign \new_[21683]_  = \new_[24842]_  & \new_[28492]_ ;
  assign \new_[21684]_  = \new_[25710]_  & \new_[26118]_ ;
  assign \new_[21685]_  = \new_[25679]_  & \new_[25381]_ ;
  assign \new_[21686]_  = ~\new_[25169]_  | ~\new_[28551]_ ;
  assign \new_[21687]_  = \new_[24992]_  | \new_[26893]_ ;
  assign \new_[21688]_  = \new_[25664]_  & \new_[25665]_ ;
  assign \new_[21689]_  = \new_[24848]_  | \new_[29810]_ ;
  assign \new_[21690]_  = \new_[24985]_  | \new_[29815]_ ;
  assign \new_[21691]_  = \new_[25396]_  & \new_[25397]_ ;
  assign \new_[21692]_  = \new_[24981]_  | \new_[25057]_ ;
  assign \new_[21693]_  = \new_[24866]_  & \new_[28481]_ ;
  assign \new_[21694]_  = \new_[25400]_  & \new_[25401]_ ;
  assign \new_[21695]_  = ~\new_[26908]_  | ~\new_[26576]_ ;
  assign \new_[21696]_  = ~\new_[24953]_  | ~\new_[29260]_ ;
  assign \new_[21697]_  = \new_[26411]_  & \new_[25408]_ ;
  assign \new_[21698]_  = \new_[24857]_  | \new_[26381]_ ;
  assign \new_[21699]_  = ~\new_[24858]_  | ~\new_[28519]_ ;
  assign \new_[21700]_  = \new_[25795]_  & \new_[25416]_ ;
  assign \new_[21701]_  = ~\new_[24943]_  | ~\new_[28519]_ ;
  assign \new_[21702]_  = \new_[24669]_  & \new_[26371]_ ;
  assign \new_[21703]_  = ~\new_[24872]_  | ~\new_[27737]_ ;
  assign \new_[21704]_  = \new_[25553]_  & \new_[25543]_ ;
  assign \new_[21705]_  = ~\new_[25035]_  | ~\new_[27709]_ ;
  assign \new_[21706]_  = ~\new_[26565]_  | ~\new_[24997]_ ;
  assign \new_[21707]_  = ~\new_[24987]_  | ~\new_[28186]_ ;
  assign \new_[21708]_  = \new_[24913]_  | \new_[30275]_ ;
  assign \new_[21709]_  = ~\new_[26915]_  & ~\new_[26564]_ ;
  assign \new_[21710]_  = \new_[24707]_  & \new_[25320]_ ;
  assign \new_[21711]_  = \new_[25309]_  & \new_[25429]_ ;
  assign \new_[21712]_  = ~\new_[24873]_  | ~\new_[27098]_ ;
  assign \new_[21713]_  = ~\new_[24878]_  & ~\new_[29765]_ ;
  assign \new_[21714]_  = ~\new_[24935]_  | ~\new_[24577]_ ;
  assign \new_[21715]_  = \new_[24864]_  | \new_[24878]_ ;
  assign \new_[21716]_  = ~\new_[26562]_  | ~\new_[30784]_ ;
  assign \new_[21717]_  = ~\new_[24864]_  & ~\new_[29765]_ ;
  assign \new_[21718]_  = \new_[25424]_  & \new_[25342]_ ;
  assign \new_[21719]_  = ~\new_[24869]_  & ~\new_[30785]_ ;
  assign \new_[21720]_  = \new_[25094]_  | \new_[30199]_ ;
  assign \new_[21721]_  = \new_[24990]_  & \new_[28122]_ ;
  assign \new_[21722]_  = \new_[24801]_  & \new_[25911]_ ;
  assign \new_[21723]_  = ~\new_[26551]_  | ~\new_[29692]_ ;
  assign \new_[21724]_  = ~\new_[24875]_  | ~\new_[26933]_ ;
  assign \new_[21725]_  = ~\new_[24877]_  | ~\new_[28542]_ ;
  assign \new_[21726]_  = \new_[24552]_  & \new_[26013]_ ;
  assign \new_[21727]_  = ~\new_[25078]_  & ~\new_[25488]_ ;
  assign \new_[21728]_  = ~\new_[24891]_  | ~\new_[27602]_ ;
  assign \new_[21729]_  = ~\new_[25064]_  & ~\new_[25488]_ ;
  assign \new_[21730]_  = ~\new_[26914]_  & ~\new_[24892]_ ;
  assign \new_[21731]_  = ~\new_[24934]_  | ~\new_[27401]_ ;
  assign \new_[21732]_  = \new_[24896]_  | \new_[30093]_ ;
  assign \new_[21733]_  = \new_[24971]_  | \new_[30010]_ ;
  assign \new_[21734]_  = ~\new_[24851]_  | ~\new_[24957]_ ;
  assign \new_[21735]_  = ~\new_[26919]_  | ~\new_[24955]_ ;
  assign \new_[21736]_  = \new_[24900]_  | \new_[30066]_ ;
  assign \new_[21737]_  = ~\new_[26915]_  | ~\new_[26564]_ ;
  assign \new_[21738]_  = ~\new_[25149]_  | ~\new_[24874]_ ;
  assign \new_[21739]_  = ~\new_[26487]_  | ~\new_[26922]_ ;
  assign \new_[21740]_  = ~\new_[24837]_  | ~\new_[24838]_ ;
  assign \new_[21741]_  = \new_[24757]_  & \new_[25790]_ ;
  assign \new_[21742]_  = ~\new_[25119]_  | ~\new_[25124]_ ;
  assign \new_[21743]_  = ~\new_[24938]_  | ~\new_[27730]_ ;
  assign \new_[21744]_  = ~\new_[25001]_  | ~\new_[30774]_ ;
  assign \new_[21745]_  = ~\new_[26909]_  | ~\new_[24880]_ ;
  assign \new_[21746]_  = ~\new_[24411]_ ;
  assign \new_[21747]_  = \new_[25536]_  & \new_[25533]_ ;
  assign \new_[21748]_  = ~\new_[26873]_  | ~\new_[24810]_ ;
  assign \new_[21749]_  = ~\new_[26884]_  | ~\new_[24825]_ ;
  assign \new_[21750]_  = ~\new_[24910]_  & ~\new_[26314]_ ;
  assign \new_[21751]_  = ~\new_[26487]_  & ~\new_[26922]_ ;
  assign \new_[21752]_  = ~\new_[25180]_  | ~\new_[26607]_ ;
  assign \new_[21753]_  = ~\new_[25072]_  | ~\new_[27401]_ ;
  assign \new_[21754]_  = \new_[25301]_  & \new_[26111]_ ;
  assign \new_[21755]_  = \new_[25394]_  & \new_[25706]_ ;
  assign \new_[21756]_  = \new_[25425]_  & \new_[26797]_ ;
  assign \new_[21757]_  = ~\new_[24921]_  | ~\new_[27662]_ ;
  assign \new_[21758]_  = \new_[25555]_  & \new_[26569]_ ;
  assign \new_[21759]_  = ~\new_[30127]_  | ~\new_[5921]_ ;
  assign \new_[21760]_  = ~\new_[24939]_  | ~\new_[26980]_ ;
  assign \new_[21761]_  = ~\new_[25070]_  | ~\new_[24743]_ ;
  assign \new_[21762]_  = ~\new_[24928]_  & ~\new_[29865]_ ;
  assign \new_[21763]_  = \new_[25701]_  & \new_[24622]_ ;
  assign \new_[21764]_  = ~\new_[24859]_  | ~\new_[26609]_ ;
  assign \new_[21765]_  = \new_[25578]_  & \new_[27199]_ ;
  assign \new_[21766]_  = ~\new_[28004]_  | ~\new_[5909]_ ;
  assign \new_[21767]_  = \new_[25868]_  & \new_[25871]_ ;
  assign \new_[21768]_  = ~\new_[24938]_  | ~\new_[24922]_ ;
  assign \new_[21769]_  = \new_[26384]_  | \new_[24924]_ ;
  assign \new_[21770]_  = \new_[25541]_  & \new_[26696]_ ;
  assign \new_[21771]_  = ~\new_[25162]_  | ~\new_[24615]_ ;
  assign \new_[21772]_  = \new_[26010]_  & \new_[25331]_ ;
  assign \new_[21773]_  = \new_[25592]_  & \new_[27139]_ ;
  assign \new_[21774]_  = \new_[25045]_  | \new_[30115]_ ;
  assign \new_[21775]_  = ~\new_[30103]_  | ~\new_[30046]_ ;
  assign \new_[21776]_  = \new_[24695]_  & \new_[26783]_ ;
  assign \new_[21777]_  = ~\new_[25018]_  | ~\new_[29202]_ ;
  assign \new_[21778]_  = \new_[25645]_  & \new_[25343]_ ;
  assign \new_[21779]_  = ~\new_[24996]_  & ~\new_[26825]_ ;
  assign \new_[21780]_  = \new_[25605]_  & \new_[25620]_ ;
  assign \new_[21781]_  = ~\new_[24988]_  & ~\new_[26825]_ ;
  assign \new_[21782]_  = ~\new_[30785]_  & ~\new_[28317]_ ;
  assign \new_[21783]_  = \new_[25612]_  & \new_[27216]_ ;
  assign \new_[21784]_  = ~\new_[25056]_  | ~\new_[28294]_ ;
  assign \new_[21785]_  = ~\new_[24899]_  | ~\new_[29139]_ ;
  assign \new_[21786]_  = \new_[25499]_  & \new_[27156]_ ;
  assign \new_[21787]_  = ~\new_[24963]_  & ~\new_[27540]_ ;
  assign \new_[21788]_  = \new_[25625]_  & \new_[27073]_ ;
  assign \new_[21789]_  = ~\new_[24976]_  & ~\new_[30029]_ ;
  assign \new_[21790]_  = \new_[25316]_  & \new_[27249]_ ;
  assign \new_[21791]_  = \new_[24641]_  & \new_[25848]_ ;
  assign \new_[21792]_  = \new_[25085]_  | \new_[29907]_ ;
  assign \new_[21793]_  = ~\new_[27527]_  & ~\new_[24976]_ ;
  assign \new_[21794]_  = ~\new_[24685]_  & ~\new_[30632]_ ;
  assign \new_[21795]_  = \new_[24905]_  & \new_[28522]_ ;
  assign \new_[21796]_  = \new_[25902]_  & \new_[27716]_ ;
  assign \new_[21797]_  = ~\new_[24944]_  | ~\new_[30246]_ ;
  assign \new_[21798]_  = ~\new_[24149]_ ;
  assign \new_[21799]_  = \new_[25427]_  & \new_[25831]_ ;
  assign \new_[21800]_  = \new_[25606]_  & \new_[27233]_ ;
  assign \new_[21801]_  = \new_[24992]_  | \new_[30629]_ ;
  assign \new_[21802]_  = ~\new_[24978]_  | ~\new_[28798]_ ;
  assign \new_[21803]_  = \new_[25433]_  & \new_[27071]_ ;
  assign \new_[21804]_  = ~\new_[25208]_  | ~\new_[27633]_ ;
  assign \new_[21805]_  = \new_[25804]_  & \new_[25353]_ ;
  assign \new_[21806]_  = ~\new_[24979]_  | ~\new_[27510]_ ;
  assign \new_[21807]_  = \new_[26059]_  & \new_[28550]_ ;
  assign \new_[21808]_  = ~\new_[25026]_  & ~\new_[30581]_ ;
  assign \new_[21809]_  = \new_[25364]_  & \new_[27082]_ ;
  assign \new_[21810]_  = ~\new_[25037]_  | ~\new_[28384]_ ;
  assign \new_[21811]_  = ~\new_[25201]_  & ~\new_[30062]_ ;
  assign \new_[21812]_  = ~\new_[25019]_  | ~\new_[28291]_ ;
  assign \new_[21813]_  = ~\new_[24691]_  & ~\new_[30616]_ ;
  assign \new_[21814]_  = \new_[24597]_  & \new_[25067]_ ;
  assign \new_[21815]_  = ~\new_[25016]_  | ~\new_[28798]_ ;
  assign \new_[21816]_  = ~\new_[24840]_  & ~\new_[29908]_ ;
  assign \new_[21817]_  = \new_[24840]_  | \new_[25017]_ ;
  assign \new_[21818]_  = \new_[25722]_  & \new_[25724]_ ;
  assign \new_[21819]_  = \new_[24534]_  & \new_[27969]_ ;
  assign \new_[21820]_  = ~\new_[25086]_  | ~\new_[26319]_ ;
  assign \new_[21821]_  = ~\new_[24828]_  | ~\new_[27724]_ ;
  assign \new_[21822]_  = ~\new_[25017]_  & ~\new_[29908]_ ;
  assign \new_[21823]_  = ~\new_[24280]_ ;
  assign \new_[21824]_  = ~\new_[25000]_  & ~\new_[30062]_ ;
  assign \new_[21825]_  = \new_[25021]_  | \new_[26804]_ ;
  assign \new_[21826]_  = ~\new_[24952]_  & ~\new_[29994]_ ;
  assign \new_[21827]_  = ~\new_[24999]_  & ~\new_[26431]_ ;
  assign \new_[21828]_  = \new_[25199]_  & \new_[26806]_ ;
  assign \new_[21829]_  = ~\new_[25027]_  | ~\new_[30125]_ ;
  assign \new_[21830]_  = ~\new_[24892]_  & ~\new_[29889]_ ;
  assign \new_[21831]_  = \new_[25004]_  | \new_[30075]_ ;
  assign \new_[21832]_  = \new_[25518]_  & \new_[25312]_ ;
  assign \new_[21833]_  = ~\new_[25020]_  | ~\new_[30316]_ ;
  assign \new_[21834]_  = ~\new_[25132]_  | ~\new_[25131]_ ;
  assign \new_[21835]_  = ~\new_[29914]_  | ~\new_[5917]_ ;
  assign \new_[21836]_  = \new_[25051]_  | \new_[30188]_ ;
  assign \new_[21837]_  = ~\new_[24977]_  | ~\new_[29887]_ ;
  assign \new_[21838]_  = ~\new_[24862]_  & ~\new_[30649]_ ;
  assign \new_[21839]_  = \new_[25700]_  & \new_[25801]_ ;
  assign \new_[21840]_  = ~\new_[25111]_  | ~\new_[25112]_ ;
  assign \new_[21841]_  = \new_[25028]_  | \new_[26960]_ ;
  assign \new_[21842]_  = \new_[25755]_  & \new_[25420]_ ;
  assign \new_[21843]_  = ~\new_[25082]_  | ~\new_[30615]_ ;
  assign \new_[21844]_  = \new_[25044]_  | \new_[30677]_ ;
  assign \new_[21845]_  = ~\new_[25188]_  & ~\new_[30840]_ ;
  assign \new_[21846]_  = \new_[26553]_  | \new_[28800]_ ;
  assign \new_[21847]_  = ~\new_[26985]_  | ~\new_[24890]_ ;
  assign \new_[21848]_  = \new_[25714]_  & \new_[25308]_ ;
  assign \new_[21849]_  = \new_[25781]_  & \new_[25957]_ ;
  assign \new_[21850]_  = ~\new_[25175]_  | ~\new_[24705]_ ;
  assign \new_[21851]_  = \new_[25889]_  & \new_[25854]_ ;
  assign \new_[21852]_  = \new_[25000]_  | \new_[25201]_ ;
  assign \new_[21853]_  = \new_[25793]_  & \new_[26514]_ ;
  assign \new_[21854]_  = ~\new_[30231]_  | ~\new_[5894]_ ;
  assign \new_[21855]_  = ~\new_[25107]_  & ~\new_[29772]_ ;
  assign \new_[21856]_  = \new_[25662]_  & \new_[25616]_ ;
  assign \new_[21857]_  = \new_[24625]_  & \new_[26042]_ ;
  assign \new_[21858]_  = ~\new_[25077]_  | ~\new_[26373]_ ;
  assign \new_[21859]_  = \new_[24701]_  & \new_[25913]_ ;
  assign \new_[21860]_  = \new_[26091]_  & \new_[25719]_ ;
  assign \new_[21861]_  = \new_[25798]_  & \new_[25464]_ ;
  assign \new_[21862]_  = \new_[26574]_  & \new_[25387]_ ;
  assign \new_[21863]_  = \new_[25791]_  & \new_[26100]_ ;
  assign \new_[21864]_  = ~\new_[24975]_  | ~\new_[26219]_ ;
  assign \new_[21865]_  = \new_[25402]_  & \new_[25326]_ ;
  assign \new_[21866]_  = \new_[25821]_  & \new_[27554]_ ;
  assign \new_[21867]_  = ~\new_[26983]_  | ~\new_[24887]_ ;
  assign \new_[21868]_  = \new_[25760]_  & \new_[25826]_ ;
  assign \new_[21869]_  = \new_[25734]_  & \new_[25749]_ ;
  assign \new_[21870]_  = \new_[25827]_  & \new_[25738]_ ;
  assign \new_[21871]_  = ~\new_[25055]_  | ~\new_[30789]_ ;
  assign \new_[21872]_  = \new_[24826]_  | \new_[29909]_ ;
  assign \new_[21873]_  = \new_[24611]_  & \new_[25841]_ ;
  assign \new_[21874]_  = \new_[25610]_  & \new_[25842]_ ;
  assign \new_[21875]_  = \new_[26024]_  & \new_[25851]_ ;
  assign \new_[21876]_  = \new_[25859]_  & \new_[26046]_ ;
  assign \new_[21877]_  = \new_[25860]_  & \new_[27151]_ ;
  assign \new_[21878]_  = \new_[25872]_  & \new_[25873]_ ;
  assign \new_[21879]_  = ~\new_[24911]_  | ~\new_[26197]_ ;
  assign \new_[21880]_  = \new_[25212]_  & \new_[25879]_ ;
  assign \new_[21881]_  = ~\new_[26506]_  | ~\new_[26502]_ ;
  assign \new_[21882]_  = ~\new_[26853]_  & ~\new_[30375]_ ;
  assign \new_[21883]_  = \new_[25174]_  & \new_[25882]_ ;
  assign \new_[21884]_  = ~\new_[28675]_  | ~\new_[29918]_ ;
  assign \new_[21885]_  = \new_[25528]_  & \new_[25894]_ ;
  assign \new_[21886]_  = ~\new_[25091]_  | ~\new_[26839]_ ;
  assign \new_[21887]_  = \new_[25903]_  & \new_[25904]_ ;
  assign \new_[21888]_  = \new_[25909]_  & \new_[25434]_ ;
  assign \new_[21889]_  = ~\new_[25207]_  & ~\new_[30688]_ ;
  assign \new_[21890]_  = \new_[25908]_  & \new_[24856]_ ;
  assign \new_[21891]_  = \new_[25498]_  & \new_[25493]_ ;
  assign \new_[21892]_  = \new_[24834]_  & \new_[25914]_ ;
  assign \new_[21893]_  = \new_[25919]_  & \new_[25431]_ ;
  assign \new_[21894]_  = \new_[25098]_  | \new_[30326]_ ;
  assign \new_[21895]_  = \new_[24767]_  & \new_[25926]_ ;
  assign \new_[21896]_  = \new_[25933]_  & \new_[25935]_ ;
  assign \new_[21897]_  = ~\new_[24937]_  & ~\new_[30568]_ ;
  assign \new_[21898]_  = ~\new_[25102]_  & ~\new_[30618]_ ;
  assign \new_[21899]_  = ~\new_[29916]_  | ~\new_[6073]_ ;
  assign \new_[21900]_  = \new_[26232]_  & \new_[27409]_ ;
  assign \new_[21901]_  = \new_[25148]_  & \new_[25953]_ ;
  assign \new_[21902]_  = \new_[25956]_  & \new_[24676]_ ;
  assign \new_[21903]_  = \new_[25530]_  & \new_[25613]_ ;
  assign \new_[21904]_  = ~\new_[24936]_  & ~\new_[24558]_ ;
  assign \new_[21905]_  = \new_[24727]_  & \new_[25970]_ ;
  assign \new_[21906]_  = ~\new_[25101]_  | ~\new_[30507]_ ;
  assign \new_[21907]_  = \new_[25978]_  & \new_[25980]_ ;
  assign \new_[21908]_  = \new_[24696]_  & \new_[25984]_ ;
  assign \new_[21909]_  = \new_[24933]_  & \new_[28164]_ ;
  assign \new_[21910]_  = \new_[26131]_  & \new_[26138]_ ;
  assign \new_[21911]_  = \new_[25991]_  & \new_[24679]_ ;
  assign \new_[21912]_  = ~\new_[25022]_  | ~\new_[29744]_ ;
  assign \new_[21913]_  = ~\new_[24805]_  | ~\new_[24974]_ ;
  assign \new_[21914]_  = ~\new_[24932]_  & ~\new_[24558]_ ;
  assign \new_[21915]_  = ~\new_[25103]_  | ~\new_[26522]_ ;
  assign \new_[21916]_  = \new_[26005]_  & \new_[26007]_ ;
  assign \new_[21917]_  = ~\new_[26983]_  & ~\new_[24887]_ ;
  assign \new_[21918]_  = ~\new_[26873]_  & ~\new_[24810]_ ;
  assign \new_[21919]_  = ~\new_[26884]_  & ~\new_[24825]_ ;
  assign \new_[21920]_  = ~\new_[26736]_  & ~\new_[24607]_ ;
  assign \new_[21921]_  = ~\new_[29020]_  | ~\new_[29401]_ ;
  assign \new_[21922]_  = \new_[26021]_  & \new_[24678]_ ;
  assign \new_[21923]_  = \new_[24655]_  & \new_[26015]_ ;
  assign \new_[21924]_  = ~\new_[26985]_  & ~\new_[24890]_ ;
  assign \new_[21925]_  = \new_[26908]_  | \new_[26576]_ ;
  assign \new_[21926]_  = \new_[25838]_  & \new_[26036]_ ;
  assign \new_[21927]_  = \new_[25950]_  & \new_[25506]_ ;
  assign \new_[21928]_  = \new_[25044]_  | \new_[26998]_ ;
  assign \new_[21929]_  = ~\new_[25025]_  & ~\new_[30662]_ ;
  assign \new_[21930]_  = \new_[25696]_  & \new_[26039]_ ;
  assign \new_[21931]_  = \new_[25823]_  & \new_[25282]_ ;
  assign \new_[21932]_  = ~\new_[24601]_  & ~\new_[30145]_ ;
  assign \new_[21933]_  = \new_[24968]_  & \new_[28556]_ ;
  assign \new_[21934]_  = ~\new_[25047]_  | ~\new_[25708]_ ;
  assign \new_[21935]_  = \new_[24616]_  & \new_[24614]_ ;
  assign \new_[21936]_  = \new_[25041]_  & \new_[28297]_ ;
  assign \new_[21937]_  = ~\new_[25040]_  & ~\new_[24644]_ ;
  assign \new_[21938]_  = \new_[26054]_  & \new_[24608]_ ;
  assign \new_[21939]_  = ~\new_[30109]_  | ~\new_[5967]_ ;
  assign \new_[21940]_  = \new_[25733]_  & \new_[24592]_ ;
  assign \new_[21941]_  = ~\new_[26868]_  & ~\new_[24601]_ ;
  assign \new_[21942]_  = \new_[25751]_  & \new_[25642]_ ;
  assign \new_[21943]_  = \new_[24574]_  & \new_[26061]_ ;
  assign \new_[21944]_  = ~\new_[25050]_  | ~\new_[26760]_ ;
  assign \new_[21945]_  = \new_[25977]_  | \new_[29997]_ ;
  assign \new_[21946]_  = \new_[25120]_  | \new_[27356]_ ;
  assign \new_[21947]_  = \new_[25802]_  & \new_[26033]_ ;
  assign \new_[21948]_  = \new_[25681]_  & \new_[26068]_ ;
  assign \new_[21949]_  = \new_[24650]_  & \new_[26073]_ ;
  assign \new_[21950]_  = ~\new_[25049]_  | ~\new_[28700]_ ;
  assign \new_[21951]_  = \new_[25657]_  & \new_[25654]_ ;
  assign \new_[21952]_  = ~\new_[24930]_  | ~\new_[28962]_ ;
  assign \new_[21953]_  = ~\new_[25133]_  | ~\new_[28700]_ ;
  assign \new_[21954]_  = \new_[26076]_  & \new_[24581]_ ;
  assign \new_[21955]_  = \new_[26081]_  & \new_[26082]_ ;
  assign \new_[21956]_  = \new_[26488]_  | \new_[25130]_ ;
  assign \new_[21957]_  = \new_[25683]_  & \new_[26089]_ ;
  assign \new_[21958]_  = ~\new_[26488]_  & ~\new_[30277]_ ;
  assign \new_[21959]_  = ~\new_[25038]_  | ~\new_[30363]_ ;
  assign \new_[21960]_  = \new_[26096]_  & \new_[25582]_ ;
  assign \new_[21961]_  = ~\new_[25130]_  & ~\new_[30277]_ ;
  assign \new_[21962]_  = \new_[25036]_  & \new_[28305]_ ;
  assign \new_[21963]_  = \new_[25015]_  | \new_[30157]_ ;
  assign \new_[21964]_  = ~\new_[24904]_  | ~\new_[27709]_ ;
  assign \new_[21965]_  = \new_[26546]_  & \new_[26105]_ ;
  assign \new_[21966]_  = \new_[25502]_  & \new_[26537]_ ;
  assign \new_[21967]_  = ~\new_[24884]_  | ~\new_[27564]_ ;
  assign \new_[21968]_  = ~\new_[24594]_  & ~\new_[25966]_ ;
  assign \new_[21969]_  = ~\new_[25134]_  & ~\new_[30208]_ ;
  assign \new_[21970]_  = ~\new_[25135]_  | ~\new_[29350]_ ;
  assign \new_[21971]_  = \new_[24562]_  & \new_[26114]_ ;
  assign \new_[21972]_  = ~\new_[24605]_  & ~\new_[25573]_ ;
  assign \new_[21973]_  = ~\new_[25163]_  | ~\new_[25564]_ ;
  assign \new_[21974]_  = ~\new_[25136]_  & ~\new_[25573]_ ;
  assign \new_[21975]_  = ~\new_[26888]_  & ~\new_[25138]_ ;
  assign \new_[21976]_  = \new_[24811]_  | \new_[25100]_ ;
  assign \new_[21977]_  = \new_[24809]_  | \new_[27555]_ ;
  assign \new_[21978]_  = ~\new_[24799]_  | ~\new_[26194]_ ;
  assign \new_[21979]_  = \new_[25028]_  | \new_[30642]_ ;
  assign \new_[21980]_  = \new_[24794]_  | \new_[24724]_ ;
  assign \new_[21981]_  = ~\new_[25947]_  | ~\new_[27726]_ ;
  assign \new_[21982]_  = ~\new_[25144]_  | ~\new_[24620]_ ;
  assign \new_[21983]_  = \new_[24700]_  | \new_[30265]_ ;
  assign \new_[21984]_  = \new_[25003]_  & \new_[28573]_ ;
  assign \new_[21985]_  = ~\new_[25146]_  | ~\new_[30820]_ ;
  assign \new_[21986]_  = ~\new_[25057]_  & ~\new_[30024]_ ;
  assign \new_[21987]_  = \new_[24726]_  & \new_[28740]_ ;
  assign \new_[21988]_  = \new_[25142]_  | \new_[27639]_ ;
  assign \new_[21989]_  = \new_[24800]_  | \new_[28687]_ ;
  assign \new_[21990]_  = ~\new_[30325]_  & (~\new_[28509]_  | ~\new_[28871]_ );
  assign \new_[21991]_  = \new_[25087]_  | \new_[28380]_ ;
  assign \new_[21992]_  = ~\new_[28908]_  | ~\new_[27384]_  | ~\new_[27944]_ ;
  assign \new_[21993]_  = ~\new_[29907]_  & (~\new_[28394]_  | ~\new_[29483]_ );
  assign \new_[21994]_  = ~\new_[30201]_  & ~\new_[30225]_ ;
  assign \new_[21995]_  = \new_[24841]_  | \new_[27962]_ ;
  assign \new_[21996]_  = ~\new_[29112]_  | ~\new_[27942]_  | ~\new_[27495]_ ;
  assign n7889 = ~\new_[29326]_  | ~\new_[25245]_ ;
  assign \new_[21998]_  = ~\new_[30123]_  | ~\new_[28307]_  | ~\new_[27497]_ ;
  assign \new_[21999]_  = ~\new_[28968]_  | ~\new_[26845]_  | ~\new_[27394]_ ;
  assign \new_[22000]_  = \new_[24871]_  | \new_[28098]_ ;
  assign \new_[22001]_  = ~\new_[28835]_  | ~\new_[27826]_  | ~\new_[27498]_ ;
  assign \new_[22002]_  = \new_[24984]_  | \new_[27743]_ ;
  assign \new_[22003]_  = ~\new_[27740]_  | ~\new_[27952]_  | ~\new_[29415]_ ;
  assign \new_[22004]_  = ~\new_[27158]_  | ~\new_[27576]_  | ~\new_[26706]_ ;
  assign \new_[22005]_  = ~\new_[29792]_  & (~\new_[28512]_  | ~\new_[29474]_ );
  assign \new_[22006]_  = ~\new_[27365]_  | ~\new_[26863]_  | ~\new_[29665]_ ;
  assign \new_[22007]_  = ~\new_[30029]_  & (~\new_[29422]_  | ~\new_[29528]_ );
  assign \new_[22008]_  = \new_[24969]_  | \new_[27765]_ ;
  assign \new_[22009]_  = ~\new_[29633]_  | ~\new_[27191]_  | ~\new_[27492]_ ;
  assign \new_[22010]_  = ~\new_[30280]_  | ~\new_[28194]_  | ~\new_[27966]_ ;
  assign \new_[22011]_  = ~\new_[28844]_  | ~\new_[27285]_  | ~\new_[27464]_ ;
  assign \new_[22012]_  = ~\new_[30375]_  & (~\new_[28442]_  | ~\new_[29480]_ );
  assign \new_[22013]_  = ~\new_[27683]_  | ~\new_[27584]_  | ~\new_[28855]_ ;
  assign \new_[22014]_  = ~\new_[27693]_  | ~\new_[27953]_  | ~\new_[29469]_ ;
  assign \new_[22015]_  = \new_[25066]_  | \new_[27582]_ ;
  assign \new_[22016]_  = ~\new_[29189]_  | ~\new_[26596]_  | ~\new_[27524]_ ;
  assign \new_[22017]_  = ~\new_[29997]_  & (~\new_[28405]_  | ~\new_[29536]_ );
  assign \new_[22018]_  = ~\new_[28864]_  | ~\new_[26821]_  | ~\new_[26793]_ ;
  assign \new_[22019]_  = ~\new_[30336]_  & (~\new_[29478]_  | ~\new_[29305]_ );
  assign n7914 = ~\new_[29295]_  | ~\new_[25259]_ ;
  assign n7929 = ~\new_[29592]_  | ~\new_[25255]_ ;
  assign n7884 = ~\new_[29213]_  | ~\new_[25210]_ ;
  assign n7959 = ~\new_[29308]_  | ~\new_[25243]_ ;
  assign n7874 = ~\new_[29615]_  | ~\new_[25242]_ ;
  assign \new_[22025]_  = \new_[25074]_  | \new_[29468]_ ;
  assign n7964 = ~\new_[29391]_  | ~\new_[25240]_ ;
  assign n8049 = ~\new_[29080]_  | ~\new_[25216]_ ;
  assign n8044 = ~\new_[29081]_  | ~\new_[25218]_ ;
  assign \new_[22029]_  = ~\new_[26918]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign n7834 = ~\new_[29263]_  | ~\new_[25220]_ ;
  assign n8029 = ~\new_[29607]_  | ~\new_[25221]_ ;
  assign n8034 = ~\new_[29747]_  | ~\new_[25222]_ ;
  assign n7839 = ~\new_[29732]_  | ~\new_[25223]_ ;
  assign n8004 = ~\new_[29207]_  | ~\new_[25224]_ ;
  assign n8024 = ~\new_[29562]_  | ~\new_[25263]_ ;
  assign n7844 = ~\new_[29309]_  | ~\new_[25227]_ ;
  assign \new_[22037]_  = ~\new_[27538]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign n7849 = ~\new_[29270]_  | ~\new_[25262]_ ;
  assign n8009 = ~\new_[29690]_  | ~\new_[25228]_ ;
  assign n7999 = ~\new_[29259]_  | ~\new_[25229]_ ;
  assign n7854 = ~\new_[29018]_  | ~\new_[25230]_ ;
  assign n7859 = ~\new_[29023]_  | ~\new_[25231]_ ;
  assign \new_[22043]_  = ~\new_[27055]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign n7989 = ~\new_[29072]_  | ~\new_[25261]_ ;
  assign n7994 = ~\new_[28954]_  | ~\new_[25232]_ ;
  assign n7984 = ~\new_[29340]_  | ~\new_[25234]_ ;
  assign \new_[22047]_  = ~\new_[30005]_  | ~\new_[28054]_  | ~\new_[27028]_ ;
  assign n7979 = ~\new_[29610]_  | ~\new_[25235]_ ;
  assign n7974 = ~\new_[29377]_  | ~\new_[25236]_ ;
  assign n7864 = ~\new_[29141]_  | ~\new_[25237]_ ;
  assign n7869 = ~\new_[29559]_  | ~\new_[25238]_ ;
  assign n7969 = ~\new_[29239]_  | ~\new_[25241]_ ;
  assign \new_[22053]_  = ~\new_[27586]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign n8639 = m6_s3_cyc_o_reg;
  assign n7879 = ~\new_[29164]_  | ~\new_[25244]_ ;
  assign n7944 = ~\new_[29048]_  | ~\new_[25246]_ ;
  assign n7954 = ~\new_[29429]_  | ~\new_[24631]_ ;
  assign n7894 = ~\new_[29341]_  | ~\new_[25247]_ ;
  assign n7899 = ~\new_[28906]_  | ~\new_[25249]_ ;
  assign n7949 = ~\new_[28928]_  | ~\new_[25172]_ ;
  assign n7919 = ~\new_[29684]_  | ~\new_[24589]_ ;
  assign \new_[22062]_  = ~\new_[26689]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign n7904 = ~\new_[29591]_  | ~\new_[25250]_ ;
  assign n7939 = ~\new_[29653]_  | ~\new_[25252]_ ;
  assign n7934 = ~\new_[29231]_  | ~\new_[25256]_ ;
  assign n7909 = ~\new_[29253]_  | ~\new_[25257]_ ;
  assign \new_[22067]_  = ~\new_[26856]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign n8054 = ~\new_[29626]_  | ~\new_[25258]_ ;
  assign \new_[22069]_  = ~\new_[27519]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign n7924 = ~\new_[29216]_  | ~\new_[25260]_ ;
  assign \new_[22071]_  = \new_[25164]_  | \new_[29632]_ ;
  assign n8019 = ~\new_[29417]_  | ~\new_[25226]_ ;
  assign n8014 = ~\new_[29680]_  | ~\new_[25225]_ ;
  assign n8039 = ~\new_[29111]_  | ~\new_[25219]_ ;
  assign \new_[22075]_  = ~\new_[26742]_  | ~\new_[26744]_  | ~\new_[29467]_ ;
  assign \new_[22076]_  = ~\new_[28911]_  | ~\new_[27915]_  | ~\new_[27528]_ ;
  assign \new_[22077]_  = ~\new_[26828]_  | ~\new_[26807]_  | ~\new_[28847]_ ;
  assign \new_[22078]_  = \new_[25509]_  & \new_[28127]_ ;
  assign \new_[22079]_  = ~\new_[29955]_  | ~\new_[5998]_ ;
  assign \new_[22080]_  = ~\new_[25009]_  & ~\new_[27962]_ ;
  assign \new_[22081]_  = ~\new_[27591]_  & (~\new_[29444]_  | ~\new_[30132]_ );
  assign \new_[22082]_  = ~\new_[26385]_  & (~\new_[29440]_  | ~\new_[30731]_ );
  assign \new_[22083]_  = \new_[24894]_  & \new_[28275]_ ;
  assign \new_[22084]_  = \new_[24962]_  & \new_[28524]_ ;
  assign \new_[22085]_  = ~\new_[26421]_  & (~\new_[29437]_  | ~\new_[29050]_ );
  assign \new_[22086]_  = ~\new_[25008]_  & ~\new_[27582]_ ;
  assign \new_[22087]_  = ~\new_[26504]_  & (~\new_[27512]_  | ~\new_[30578]_ );
  assign \new_[22088]_  = ~\new_[26278]_  & ~\new_[27765]_ ;
  assign \new_[22089]_  = ~\new_[26198]_  | (~\new_[27272]_  & ~\new_[29375]_ );
  assign \new_[22090]_  = \new_[24916]_  & \new_[28579]_ ;
  assign n8714 = m2_s3_cyc_o_reg;
  assign \new_[22092]_  = \new_[25824]_  & \new_[28411]_ ;
  assign \new_[22093]_  = \new_[25090]_  & \new_[28276]_ ;
  assign \new_[22094]_  = \new_[25096]_  & \new_[27990]_ ;
  assign \new_[22095]_  = \new_[24931]_  & \new_[28178]_ ;
  assign \new_[22096]_  = ~\new_[26228]_  & (~\new_[29443]_  | ~\new_[30519]_ );
  assign \new_[22097]_  = ~\new_[26547]_  & (~\new_[29451]_  | ~\new_[30613]_ );
  assign \new_[22098]_  = ~\new_[26390]_  | (~\new_[27002]_  & ~\new_[30244]_ );
  assign \new_[22099]_  = ~\new_[26231]_  & (~\new_[29457]_  | ~\new_[30586]_ );
  assign \new_[22100]_  = \new_[25140]_  & \new_[28128]_ ;
  assign \new_[22101]_  = ~\new_[30726]_  | ~\new_[6203]_  | ~\new_[30015]_  | ~\new_[27587]_ ;
  assign \new_[22102]_  = \new_[23802]_ ;
  assign \new_[22103]_  = ~\new_[30719]_  | ~\new_[31499]_  | ~\new_[30603]_  | ~\new_[27506]_ ;
  assign \new_[22104]_  = ~\new_[30325]_  & ~\new_[30708]_ ;
  assign \new_[22105]_  = ~\new_[30721]_  | ~\new_[6200]_  | ~\new_[30525]_  | ~\new_[27605]_ ;
  assign \new_[22106]_  = ~\new_[26563]_  & ~\new_[6043]_ ;
  assign \new_[22107]_  = ~\new_[23338]_ ;
  assign \new_[22108]_  = ~\new_[26389]_  & ~\new_[28270]_ ;
  assign \new_[22109]_  = ~\new_[5964]_  | ~\new_[30221]_  | ~\new_[28845]_ ;
  assign \new_[22110]_  = ~\new_[24974]_  | ~\new_[29029]_ ;
  assign \new_[22111]_  = ~\new_[24674]_  | ~\new_[28845]_ ;
  assign \new_[22112]_  = ~\new_[23348]_ ;
  assign \new_[22113]_  = ~\new_[31669]_  | ~\new_[26374]_  | ~\new_[28114]_ ;
  assign \new_[22114]_  = ~\new_[29598]_  & ~\new_[31438]_ ;
  assign \new_[22115]_  = ~\new_[24745]_  & ~\new_[30066]_ ;
  assign \new_[22116]_  = \new_[25119]_  | \new_[25124]_ ;
  assign \new_[22117]_  = ~\new_[28395]_  | ~\new_[29911]_ ;
  assign \new_[22118]_  = ~\new_[28560]_  | ~\new_[26347]_ ;
  assign \new_[22119]_  = ~\new_[26256]_  & ~\new_[29952]_ ;
  assign \new_[22120]_  = ~\new_[23362]_ ;
  assign \new_[22121]_  = \new_[24675]_  | \new_[30694]_ ;
  assign \new_[22122]_  = \new_[29305]_  & \new_[29251]_ ;
  assign \new_[22123]_  = ~\new_[31394]_  | ~\new_[30217]_  | ~\new_[29233]_ ;
  assign \new_[22124]_  = \new_[26351]_  & \new_[30337]_ ;
  assign \new_[22125]_  = ~\new_[31719]_  | ~\new_[27845]_  | ~\new_[28039]_ ;
  assign \new_[22126]_  = ~\new_[26363]_  | ~\new_[29291]_ ;
  assign \new_[22127]_  = \new_[26237]_  | \new_[28317]_ ;
  assign \new_[22128]_  = ~\new_[23089]_ ;
  assign \new_[22129]_  = ~\new_[26543]_  | ~\new_[30232]_ ;
  assign \new_[22130]_  = ~\new_[27494]_  & ~\new_[26349]_ ;
  assign \new_[22131]_  = ~\new_[23386]_ ;
  assign \new_[22132]_  = ~\new_[23389]_ ;
  assign \new_[22133]_  = \new_[30211]_  & \new_[28361]_ ;
  assign \new_[22134]_  = ~\new_[23394]_ ;
  assign \new_[22135]_  = ~\new_[23396]_ ;
  assign \new_[22136]_  = ~\new_[28749]_  | ~\new_[26443]_ ;
  assign \new_[22137]_  = ~\new_[23403]_ ;
  assign \new_[22138]_  = ~\new_[23400]_ ;
  assign \new_[22139]_  = ~\new_[23401]_ ;
  assign \new_[22140]_  = \new_[26254]_  & \new_[29695]_ ;
  assign n8629 = m2_s12_cyc_o_reg;
  assign \new_[22142]_  = ~\new_[27401]_  | ~\new_[29781]_ ;
  assign \new_[22143]_  = ~\new_[26328]_  & ~\new_[29815]_ ;
  assign \new_[22144]_  = ~\new_[23408]_ ;
  assign \new_[22145]_  = ~\new_[24967]_  | ~\new_[28934]_ ;
  assign \new_[22146]_  = ~\new_[23414]_ ;
  assign \new_[22147]_  = ~\new_[30167]_  & ~\new_[26378]_ ;
  assign \new_[22148]_  = ~\new_[28090]_  | ~\new_[26083]_ ;
  assign \new_[22149]_  = ~\new_[23422]_ ;
  assign \new_[22150]_  = ~\new_[26117]_  | ~\new_[26813]_ ;
  assign \new_[22151]_  = ~\new_[23424]_ ;
  assign \new_[22152]_  = ~\new_[27567]_  | ~\new_[26267]_ ;
  assign \new_[22153]_  = \new_[26347]_  & \new_[28121]_ ;
  assign n8509 = m1_s3_cyc_o_reg;
  assign \new_[22155]_  = ~\new_[26272]_  | ~\new_[29886]_ ;
  assign \new_[22156]_  = ~\new_[30063]_  | ~\new_[6070]_ ;
  assign \new_[22157]_  = ~\new_[23428]_ ;
  assign \new_[22158]_  = ~\new_[28536]_  & ~\new_[30114]_ ;
  assign \new_[22159]_  = ~\new_[23432]_ ;
  assign \new_[22160]_  = ~\new_[30325]_  | ~\new_[6216]_ ;
  assign \new_[22161]_  = ~\new_[27359]_  | ~\new_[29505]_ ;
  assign \new_[22162]_  = ~\new_[28420]_  & ~\new_[30219]_ ;
  assign \new_[22163]_  = ~\new_[31553]_  | ~\new_[27596]_  | ~\new_[28640]_ ;
  assign \new_[22164]_  = ~\new_[5996]_  | ~\new_[30138]_  | ~\new_[30702]_ ;
  assign \new_[22165]_  = ~\new_[27737]_  | ~\new_[30048]_ ;
  assign \new_[22166]_  = \new_[27515]_  | \new_[26552]_ ;
  assign \new_[22167]_  = ~\new_[26213]_  & ~\new_[29930]_ ;
  assign \new_[22168]_  = \new_[27553]_  & \new_[30016]_ ;
  assign \new_[22169]_  = ~\new_[5913]_  | ~\new_[28880]_  | ~\new_[29692]_ ;
  assign \new_[22170]_  = ~\new_[26201]_  | ~\new_[29381]_ ;
  assign \new_[22171]_  = ~\new_[25602]_  | ~\new_[30381]_ ;
  assign \new_[22172]_  = ~\new_[23448]_ ;
  assign \new_[22173]_  = ~\new_[24570]_  | ~\new_[28880]_ ;
  assign \new_[22174]_  = ~\new_[23449]_ ;
  assign \new_[22175]_  = ~\new_[23456]_ ;
  assign \new_[22176]_  = ~\new_[27539]_  | ~\new_[26300]_ ;
  assign \new_[22177]_  = ~\new_[28542]_  | ~\new_[29763]_ ;
  assign \new_[22178]_  = ~\new_[25460]_  | ~\new_[30721]_ ;
  assign \new_[22179]_  = ~\new_[24577]_  | ~\new_[30269]_ ;
  assign \new_[22180]_  = ~\new_[28346]_  & ~\new_[30305]_ ;
  assign \new_[22181]_  = ~\new_[23460]_ ;
  assign \new_[22182]_  = ~\new_[23463]_ ;
  assign \new_[22183]_  = ~\new_[28953]_  & ~\new_[26494]_ ;
  assign \new_[22184]_  = ~\new_[23464]_ ;
  assign \new_[22185]_  = (~\new_[30106]_  | ~\s14_data_i[31] ) & (~\new_[27347]_  | ~\s12_data_i[31] );
  assign \new_[22186]_  = ~\new_[24673]_  | ~\new_[29802]_ ;
  assign \new_[22187]_  = \new_[26453]_  & \new_[29103]_ ;
  assign \new_[22188]_  = ~\new_[26162]_  & ~\new_[29465]_ ;
  assign \new_[22189]_  = ~\new_[26192]_  | ~\new_[29103]_ ;
  assign \new_[22190]_  = ~\new_[24621]_  & ~\new_[30075]_ ;
  assign \new_[22191]_  = ~\new_[24709]_  & ~\new_[29172]_ ;
  assign \new_[22192]_  = ~\new_[23467]_ ;
  assign \new_[22193]_  = \new_[26333]_  & \new_[28023]_ ;
  assign \new_[22194]_  = ~\new_[26399]_  | ~\new_[30037]_ ;
  assign \new_[22195]_  = ~\new_[25925]_  | ~\new_[30282]_ ;
  assign \new_[22196]_  = ~\new_[24787]_  | ~\new_[28840]_ ;
  assign \new_[22197]_  = \new_[28091]_  | \new_[28718]_ ;
  assign \new_[22198]_  = ~\new_[23475]_ ;
  assign \new_[22199]_  = ~\new_[25052]_  | ~\new_[26978]_ ;
  assign \new_[22200]_  = ~\new_[24632]_  & ~\new_[29959]_ ;
  assign \new_[22201]_  = \new_[26309]_  & \new_[29186]_ ;
  assign \new_[22202]_  = ~\new_[24771]_  | ~\new_[30094]_ ;
  assign \new_[22203]_  = ~\new_[26193]_  | ~\new_[30774]_ ;
  assign \new_[22204]_  = ~\new_[24748]_  | ~\new_[29867]_ ;
  assign \new_[22205]_  = ~\new_[26418]_  | ~\new_[29771]_ ;
  assign \new_[22206]_  = \new_[27577]_  & \new_[30022]_ ;
  assign \new_[22207]_  = ~\new_[26247]_  | ~\new_[28963]_ ;
  assign \new_[22208]_  = \new_[29461]_  & \new_[28888]_ ;
  assign \new_[22209]_  = ~\new_[26291]_  & ~\new_[29165]_ ;
  assign \new_[22210]_  = ~\new_[29276]_  | ~\new_[29171]_ ;
  assign \new_[22211]_  = ~\new_[23492]_ ;
  assign \new_[22212]_  = ~\new_[28089]_  | ~\new_[6190]_ ;
  assign \new_[22213]_  = ~\new_[26178]_  & ~\new_[26269]_ ;
  assign \new_[22214]_  = ~\new_[26375]_  | ~\new_[29929]_ ;
  assign \new_[22215]_  = ~\new_[23498]_ ;
  assign \new_[22216]_  = ~\new_[26258]_  & ~\new_[28846]_ ;
  assign \new_[22217]_  = ~\new_[26258]_  | ~\new_[25715]_ ;
  assign \new_[22218]_  = ~\new_[23503]_ ;
  assign \new_[22219]_  = ~\new_[26197]_  | ~\new_[28110]_ ;
  assign \new_[22220]_  = ~\new_[24491]_ ;
  assign \new_[22221]_  = ~\new_[28337]_  | ~\new_[30210]_ ;
  assign \new_[22222]_  = ~\new_[24490]_ ;
  assign \new_[22223]_  = ~\new_[31394]_  | ~\new_[29682]_  | ~\new_[30217]_ ;
  assign \new_[22224]_  = ~\new_[23509]_ ;
  assign \new_[22225]_  = ~\new_[26795]_  & ~\new_[30323]_ ;
  assign \new_[22226]_  = ~\new_[23510]_ ;
  assign \new_[22227]_  = ~\new_[24484]_ ;
  assign \new_[22228]_  = ~\new_[26548]_  | ~\new_[30279]_ ;
  assign \new_[22229]_  = ~\new_[30145]_  & ~\new_[30598]_ ;
  assign \new_[22230]_  = ~\new_[26317]_  & ~\new_[30597]_ ;
  assign \new_[22231]_  = \new_[26189]_  | \new_[30224]_ ;
  assign \new_[22232]_  = ~\new_[26437]_  | ~\new_[29721]_ ;
  assign \new_[22233]_  = ~\new_[28606]_  & ~\new_[30339]_ ;
  assign \new_[22234]_  = \new_[26239]_  & \new_[28073]_ ;
  assign \new_[22235]_  = ~\new_[26158]_  & ~\new_[30840]_ ;
  assign \new_[22236]_  = ~\new_[26613]_  | ~\new_[26309]_ ;
  assign \new_[22237]_  = ~\new_[27521]_  & ~\new_[24965]_ ;
  assign \new_[22238]_  = ~\new_[26381]_  | ~\new_[30750]_ ;
  assign \new_[22239]_  = ~\new_[24704]_  | ~\new_[28188]_ ;
  assign \new_[22240]_  = \new_[27721]_  & \new_[29904]_ ;
  assign \new_[22241]_  = ~\new_[23530]_ ;
  assign \new_[22242]_  = ~\new_[23532]_ ;
  assign \new_[22243]_  = ~\new_[26226]_  & ~\new_[30188]_ ;
  assign \new_[22244]_  = ~\new_[23536]_ ;
  assign \new_[22245]_  = ~\new_[26324]_  | ~\new_[29870]_ ;
  assign \new_[22246]_  = \new_[27574]_  | \new_[28718]_ ;
  assign \new_[22247]_  = ~\new_[23540]_ ;
  assign \new_[22248]_  = ~\new_[5931]_  | ~\new_[29563]_  | ~\new_[29560]_ ;
  assign \new_[22249]_  = ~\new_[26219]_  & ~\new_[28211]_ ;
  assign \new_[22250]_  = ~\new_[27329]_  & ~\new_[30212]_ ;
  assign \new_[22251]_  = ~\new_[23551]_ ;
  assign \new_[22252]_  = \new_[26083]_  & \new_[29983]_ ;
  assign \new_[22253]_  = ~\new_[24624]_  | ~\new_[27725]_ ;
  assign \new_[22254]_  = ~\new_[23572]_ ;
  assign \new_[22255]_  = ~\new_[23574]_ ;
  assign \new_[22256]_  = ~\new_[25861]_  & ~\new_[28950]_ ;
  assign \new_[22257]_  = ~\new_[26336]_  & ~\new_[26660]_ ;
  assign \new_[22258]_  = ~\new_[24752]_  | ~\new_[29401]_ ;
  assign \new_[22259]_  = ~\new_[23581]_ ;
  assign \new_[22260]_  = ~\new_[28817]_  | ~\new_[30645]_ ;
  assign \new_[22261]_  = ~\new_[23584]_ ;
  assign \new_[22262]_  = \new_[28513]_  & \new_[28337]_ ;
  assign \new_[22263]_  = ~\new_[23586]_ ;
  assign \new_[22264]_  = ~\new_[23590]_ ;
  assign \new_[22265]_  = \new_[26300]_  & \new_[28050]_ ;
  assign \new_[22266]_  = \new_[27004]_  | \new_[28718]_ ;
  assign \new_[22267]_  = ~\new_[26427]_  | ~\new_[30180]_ ;
  assign \new_[22268]_  = ~\new_[24661]_  | ~\new_[30258]_ ;
  assign \new_[22269]_  = ~\new_[23787]_ ;
  assign \new_[22270]_  = \new_[25466]_  & \new_[28963]_ ;
  assign \new_[22271]_  = ~\new_[25711]_  & ~\new_[29227]_ ;
  assign \new_[22272]_  = ~\new_[25711]_  & ~\new_[30053]_ ;
  assign \new_[22273]_  = ~\new_[23596]_ ;
  assign \new_[22274]_  = ~\new_[30235]_  | ~\new_[6273]_ ;
  assign \new_[22275]_  = \new_[26438]_  | \new_[28857]_ ;
  assign \new_[22276]_  = ~\new_[26214]_  & ~\new_[30287]_ ;
  assign \new_[22277]_  = \new_[26168]_  | \new_[30840]_ ;
  assign \new_[22278]_  = ~\new_[31695]_  | ~\new_[26347]_  | ~\new_[28121]_ ;
  assign \new_[22279]_  = ~\new_[26575]_  | ~\new_[29139]_ ;
  assign \new_[22280]_  = \new_[26270]_  | \new_[30224]_ ;
  assign \new_[22281]_  = ~\new_[27911]_  | ~\new_[26360]_ ;
  assign \new_[22282]_  = ~\new_[31608]_  | ~\new_[27635]_  | ~\new_[28684]_ ;
  assign \new_[22283]_  = \new_[26170]_  | \new_[30747]_ ;
  assign \new_[22284]_  = ~\new_[23618]_ ;
  assign \new_[22285]_  = ~\new_[31660]_  | ~\new_[26300]_  | ~\new_[28050]_ ;
  assign \new_[22286]_  = ~\new_[23621]_ ;
  assign \new_[22287]_  = ~\new_[23619]_ ;
  assign \new_[22288]_  = ~\new_[23620]_ ;
  assign \new_[22289]_  = \new_[25006]_  & \new_[29721]_ ;
  assign \new_[22290]_  = \new_[26339]_  | \new_[30438]_ ;
  assign \new_[22291]_  = \new_[26395]_  & \new_[28280]_ ;
  assign \new_[22292]_  = ~\new_[28111]_  & ~\new_[30703]_ ;
  assign \new_[22293]_  = ~\new_[26521]_  | ~\new_[30574]_ ;
  assign \new_[22294]_  = ~\new_[5919]_  | ~\new_[29974]_  | ~\new_[28905]_ ;
  assign \new_[22295]_  = ~\new_[23628]_ ;
  assign \new_[22296]_  = ~\new_[28573]_  & ~\new_[28204]_ ;
  assign \new_[22297]_  = ~\new_[31408]_  | ~\new_[26239]_  | ~\new_[28073]_ ;
  assign \new_[22298]_  = ~\new_[28153]_  | ~\new_[26239]_ ;
  assign \new_[22299]_  = ~\new_[23632]_ ;
  assign \new_[22300]_  = ~\new_[31624]_  | ~\new_[27769]_  | ~\new_[30491]_ ;
  assign \new_[22301]_  = \new_[27353]_  & \new_[29984]_ ;
  assign \new_[22302]_  = ~\new_[23640]_ ;
  assign \new_[22303]_  = ~\new_[26412]_  | ~\new_[24782]_ ;
  assign \new_[22304]_  = ~\new_[24541]_  & ~\new_[29047]_ ;
  assign \new_[22305]_  = ~\new_[27281]_  & ~\new_[25800]_ ;
  assign \new_[22306]_  = ~\new_[26348]_  | ~\new_[28382]_ ;
  assign \new_[22307]_  = ~\new_[23655]_ ;
  assign \new_[22308]_  = ~\new_[24633]_  & ~\new_[30265]_ ;
  assign \new_[22309]_  = ~\new_[23657]_ ;
  assign \new_[22310]_  = ~\new_[24554]_  | ~\new_[29175]_ ;
  assign \new_[22311]_  = ~\new_[23660]_ ;
  assign \new_[22312]_  = ~\new_[26509]_  | ~\new_[29785]_ ;
  assign \new_[22313]_  = ~\new_[24583]_  | ~\new_[30784]_ ;
  assign \new_[22314]_  = ~\new_[23662]_ ;
  assign \new_[22315]_  = ~\new_[26295]_  | ~\new_[29593]_ ;
  assign \new_[22316]_  = \new_[26388]_  | \new_[30438]_ ;
  assign \new_[22317]_  = ~\new_[5999]_  | ~\new_[28889]_  | ~\new_[29685]_ ;
  assign \new_[22318]_  = ~\new_[26476]_  | ~\new_[26852]_ ;
  assign \new_[22319]_  = ~\new_[23667]_ ;
  assign \new_[22320]_  = ~\new_[26211]_  | ~\new_[29695]_ ;
  assign \new_[22321]_  = ~\new_[24783]_  | ~\new_[30102]_ ;
  assign \new_[22322]_  = \new_[25483]_  | \new_[30637]_ ;
  assign \new_[22323]_  = ~\new_[28574]_  & ~\new_[30087]_ ;
  assign \new_[22324]_  = ~\new_[24074]_ ;
  assign \new_[22325]_  = ~\new_[26403]_  & ~\new_[30118]_ ;
  assign \new_[22326]_  = ~\new_[31229]_  | ~\new_[26443]_  | ~\new_[28732]_ ;
  assign \new_[22327]_  = ~\new_[24665]_  | ~\new_[29589]_ ;
  assign \new_[22328]_  = ~\new_[26973]_  & ~\new_[29113]_ ;
  assign \new_[22329]_  = \new_[24782]_  & \new_[29593]_ ;
  assign \new_[22330]_  = ~\new_[26345]_  | ~\new_[30211]_ ;
  assign \new_[22331]_  = ~\new_[26248]_  & ~\new_[29157]_ ;
  assign \new_[22332]_  = \new_[27926]_  & \new_[29435]_ ;
  assign \new_[22333]_  = ~\new_[26394]_  | ~\new_[29978]_ ;
  assign \new_[22334]_  = \new_[26360]_  & \new_[28245]_ ;
  assign \new_[22335]_  = ~\new_[27341]_  & ~\new_[26571]_ ;
  assign \new_[22336]_  = ~\new_[31643]_  | ~\new_[26360]_  | ~\new_[28245]_ ;
  assign \new_[22337]_  = ~\new_[29754]_  & ~\new_[26397]_ ;
  assign \new_[22338]_  = ~\new_[23697]_ ;
  assign \new_[22339]_  = ~\new_[5997]_  | ~\new_[30126]_  | ~\new_[28926]_ ;
  assign \new_[22340]_  = ~\new_[23698]_ ;
  assign \new_[22341]_  = ~\new_[24566]_  | ~\new_[30426]_ ;
  assign \new_[22342]_  = ~\new_[30762]_  | ~\new_[6200]_ ;
  assign \new_[22343]_  = ~\new_[26355]_  & ~\new_[30157]_ ;
  assign \new_[22344]_  = \new_[26030]_  & \new_[26031]_ ;
  assign \new_[22345]_  = ~\new_[23711]_ ;
  assign \new_[22346]_  = ~\new_[31725]_  | ~\new_[27568]_  | ~\new_[30628]_ ;
  assign \new_[22347]_  = ~\new_[24016]_ ;
  assign \new_[22348]_  = ~\new_[26344]_  | ~\new_[29223]_ ;
  assign \new_[22349]_  = ~\new_[23713]_ ;
  assign \new_[22350]_  = ~\new_[23717]_ ;
  assign \new_[22351]_  = ~\new_[27284]_  | ~\new_[26292]_ ;
  assign \new_[22352]_  = \new_[26296]_  | \new_[28857]_ ;
  assign \new_[22353]_  = \new_[26422]_  | \new_[28893]_ ;
  assign \new_[22354]_  = ~\new_[23727]_ ;
  assign \new_[22355]_  = ~\new_[31837]_  | ~\new_[26333]_  | ~\new_[28023]_ ;
  assign \new_[22356]_  = \new_[26292]_  & \new_[29969]_ ;
  assign \new_[22357]_  = ~\new_[31862]_  | ~\new_[26395]_  | ~\new_[28280]_ ;
  assign \new_[22358]_  = ~\new_[23732]_ ;
  assign \new_[22359]_  = \new_[27854]_  | \new_[28402]_ ;
  assign \new_[22360]_  = ~\new_[24754]_  | ~\new_[29506]_ ;
  assign \new_[22361]_  = ~\new_[23736]_ ;
  assign \new_[22362]_  = ~\new_[23738]_ ;
  assign \new_[22363]_  = ~\new_[24688]_  & ~\new_[28204]_ ;
  assign \new_[22364]_  = ~\new_[26373]_  | ~\new_[29332]_ ;
  assign \new_[22365]_  = ~\new_[26433]_  | ~\new_[30333]_ ;
  assign \new_[22366]_  = ~\new_[26257]_  | ~\new_[29881]_ ;
  assign \new_[22367]_  = \new_[30381]_  & \new_[27959]_ ;
  assign \new_[22368]_  = ~\new_[26831]_  | ~\new_[26333]_ ;
  assign \new_[22369]_  = \new_[26291]_  | \new_[29999]_ ;
  assign \new_[22370]_  = \new_[26267]_  & \new_[30117]_ ;
  assign \new_[22371]_  = \new_[26843]_  & \new_[28285]_ ;
  assign \new_[22372]_  = ~\new_[26322]_  & ~\new_[29909]_ ;
  assign \new_[22373]_  = \new_[25811]_  | \new_[30663]_ ;
  assign \new_[22374]_  = ~\new_[26319]_  | ~\new_[29145]_ ;
  assign \new_[22375]_  = ~\new_[26299]_  & ~\new_[29909]_ ;
  assign \new_[22376]_  = ~\new_[29955]_  | ~\new_[5997]_ ;
  assign \new_[22377]_  = ~\new_[27729]_  | ~\new_[26395]_ ;
  assign \new_[22378]_  = ~\new_[23759]_ ;
  assign \new_[22379]_  = ~\new_[25330]_  & ~\new_[30445]_ ;
  assign \new_[22380]_  = ~\new_[26468]_  | ~\new_[28280]_ ;
  assign \new_[22381]_  = \new_[30094]_  & \new_[26857]_ ;
  assign \new_[22382]_  = \new_[26443]_  & \new_[28732]_ ;
  assign \new_[22383]_  = ~\new_[23771]_ ;
  assign \new_[22384]_  = ~\new_[24778]_  | ~\new_[28865]_ ;
  assign \new_[22385]_  = ~\new_[23772]_ ;
  assign \new_[22386]_  = ~\new_[26158]_  | ~\new_[25550]_ ;
  assign \new_[22387]_  = ~\new_[24710]_  | ~\new_[29924]_ ;
  assign \new_[22388]_  = ~\new_[28748]_  & ~\new_[24774]_ ;
  assign \new_[22389]_  = ~\new_[31362]_  | ~\new_[26745]_  | ~\new_[30544]_ ;
  assign \new_[22390]_  = \new_[26159]_  | \new_[30632]_ ;
  assign \new_[22391]_  = ~\new_[31915]_  | ~\new_[27904]_  | ~\new_[28069]_ ;
  assign \new_[22392]_  = ~\new_[28824]_  & ~\new_[26234]_ ;
  assign \new_[22393]_  = ~\new_[23779]_ ;
  assign \new_[22394]_  = \new_[26374]_  & \new_[28114]_ ;
  assign \new_[22395]_  = ~\new_[24662]_  | ~\new_[30707]_ ;
  assign \new_[22396]_  = ~\new_[23781]_ ;
  assign \new_[22397]_  = ~\new_[27551]_  | ~\new_[26374]_ ;
  assign \new_[22398]_  = ~\new_[30074]_  & ~\new_[25829]_ ;
  assign \new_[22399]_  = ~\new_[5931]_  | ~\new_[30333]_  | ~\new_[29563]_ ;
  assign \new_[22400]_  = ~\new_[24445]_ ;
  assign \new_[22401]_  = ~\new_[26199]_  | ~\new_[27594]_ ;
  assign \new_[22402]_  = ~\new_[23788]_ ;
  assign \new_[22403]_  = ~\new_[31683]_  | ~\new_[27594]_  | ~\new_[28355]_ ;
  assign \new_[22404]_  = ~\new_[28358]_  & ~\new_[26294]_ ;
  assign \new_[22405]_  = ~\new_[26724]_  | ~\new_[28535]_ ;
  assign \new_[22406]_  = ~\new_[24656]_  & ~\new_[29985]_ ;
  assign \new_[22407]_  = ~\new_[23799]_ ;
  assign \new_[22408]_  = ~\new_[25861]_  & ~\new_[29652]_ ;
  assign \new_[22409]_  = ~\new_[29028]_  | ~\new_[30164]_ ;
  assign \new_[22410]_  = \new_[26468]_  & \new_[29571]_ ;
  assign \new_[22411]_  = ~\new_[23802]_ ;
  assign \new_[22412]_  = ~\new_[23806]_ ;
  assign \new_[22413]_  = \new_[23812]_ ;
  assign \new_[22414]_  = ~\new_[26422]_  & ~\new_[28029]_ ;
  assign \new_[22415]_  = ~\new_[23814]_ ;
  assign \new_[22416]_  = ~\new_[26245]_  | ~\new_[29979]_ ;
  assign \new_[22417]_  = ~\new_[26364]_  | ~\new_[28437]_ ;
  assign \new_[22418]_  = ~\new_[25708]_  | ~\new_[29042]_ ;
  assign \new_[22419]_  = ~\new_[23819]_ ;
  assign \new_[22420]_  = ~\new_[24993]_  | ~\new_[27997]_ ;
  assign \new_[22421]_  = ~\new_[30315]_  | ~\new_[5998]_ ;
  assign \new_[22422]_  = ~\new_[23834]_ ;
  assign \new_[22423]_  = ~\new_[23835]_ ;
  assign \new_[22424]_  = ~\new_[23227]_ ;
  assign \new_[22425]_  = \new_[27848]_  & \new_[28935]_ ;
  assign \new_[22426]_  = ~\new_[26172]_  & ~\new_[30656]_ ;
  assign \new_[22427]_  = ~\new_[24740]_  & ~\new_[30591]_ ;
  assign \new_[22428]_  = ~\new_[26172]_  | ~\new_[24609]_ ;
  assign \new_[22429]_  = ~\new_[26357]_  | ~\new_[28935]_ ;
  assign \new_[22430]_  = ~\new_[26439]_  | ~\new_[30317]_ ;
  assign \new_[22431]_  = \new_[26357]_  & \new_[30751]_ ;
  assign \new_[22432]_  = \new_[24636]_  | \new_[30036]_ ;
  assign \new_[22433]_  = ~\new_[27709]_  | ~\new_[29825]_ ;
  assign \new_[22434]_  = ~\new_[26428]_  & ~\new_[29354]_ ;
  assign \new_[22435]_  = \new_[25413]_  | \new_[30656]_ ;
  assign \new_[22436]_  = ~\new_[24766]_  | ~\new_[28423]_ ;
  assign \new_[22437]_  = ~\new_[27496]_  & ~\new_[26203]_ ;
  assign \new_[22438]_  = \new_[27585]_  & \new_[29900]_ ;
  assign \new_[22439]_  = \new_[30258]_  & \new_[26788]_ ;
  assign \new_[22440]_  = \new_[26311]_  | \new_[30036]_ ;
  assign \new_[22441]_  = ~\new_[23854]_ ;
  assign \new_[22442]_  = ~\new_[26479]_  | ~\new_[28360]_ ;
  assign \new_[22443]_  = ~\new_[23860]_ ;
  assign \new_[22444]_  = ~\new_[26284]_  | ~\new_[30262]_ ;
  assign \new_[22445]_  = ~\new_[26162]_  & ~\new_[29931]_ ;
  assign \new_[22446]_  = ~\new_[24792]_  & ~\new_[30115]_ ;
  assign \new_[22447]_  = ~\new_[23863]_ ;
  assign \new_[22448]_  = ~\new_[26194]_  | ~\new_[29130]_ ;
  assign \new_[22449]_  = \new_[28020]_  & \new_[5981]_ ;
  assign \new_[22450]_  = ~\new_[26840]_  & ~\new_[24756]_ ;
  assign \new_[22451]_  = ~\new_[6007]_  | ~\new_[30724]_  | ~\new_[29118]_ ;
  assign \new_[22452]_  = ~\new_[23872]_ ;
  assign \new_[22453]_  = ~\new_[27726]_  | ~\new_[29768]_ ;
  assign \new_[22454]_  = ~\new_[30336]_  | ~\new_[6096]_ ;
  assign \new_[22455]_  = ~\new_[28089]_  & ~\new_[26242]_ ;
  assign \new_[22456]_  = ~\new_[23879]_ ;
  assign \new_[22457]_  = ~\new_[24751]_  & ~\new_[29700]_ ;
  assign \new_[22458]_  = ~\new_[23883]_ ;
  assign \new_[22459]_  = ~\new_[23885]_ ;
  assign \new_[22460]_  = ~\new_[6033]_  | ~\new_[29794]_  | ~\new_[30283]_ ;
  assign \new_[22461]_  = \new_[25846]_  | \new_[30303]_ ;
  assign \new_[22462]_  = ~\new_[28668]_  & ~\new_[25508]_ ;
  assign \new_[22463]_  = ~\new_[26038]_  & (~\new_[29028]_  | ~\new_[6035]_ );
  assign \new_[22464]_  = ~\new_[27991]_  & ~\new_[26353]_ ;
  assign \new_[22465]_  = ~\new_[6040]_  | ~\new_[30111]_  | ~\new_[30337]_ ;
  assign \new_[22466]_  = \new_[26214]_  & \new_[26320]_ ;
  assign \new_[22467]_  = \new_[26746]_  & \new_[26538]_ ;
  assign \new_[22468]_  = ~\new_[26222]_  & (~\new_[29583]_  | ~\new_[6081]_ );
  assign \new_[22469]_  = ~\new_[5918]_  | ~\new_[29619]_  | ~\new_[29633]_ ;
  assign \new_[22470]_  = ~\new_[28548]_  & ~\new_[26326]_ ;
  assign \new_[22471]_  = ~\new_[24566]_  & ~\new_[24561]_ ;
  assign \new_[22472]_  = ~\new_[5911]_  | ~\new_[30079]_  | ~\new_[29112]_ ;
  assign \new_[22473]_  = ~\new_[24852]_  & (~\new_[28918]_  | ~\new_[6044]_ );
  assign \new_[22474]_  = ~\new_[24760]_  & (~\new_[28836]_  | ~\new_[6047]_ );
  assign \new_[22475]_  = ~\new_[29880]_  | ~\new_[6245]_ ;
  assign \new_[22476]_  = ~\new_[31491]_  | ~\new_[24653]_  | ~\new_[28344]_ ;
  assign \new_[22477]_  = ~\new_[27601]_  & ~\new_[26401]_ ;
  assign \new_[22478]_  = ~\new_[5914]_  | ~\new_[30312]_  | ~\new_[28835]_ ;
  assign \new_[22479]_  = \new_[25621]_  | \new_[28651]_ ;
  assign \new_[22480]_  = ~\new_[5912]_  | ~\new_[28070]_  | ~\new_[28968]_ ;
  assign \new_[22481]_  = ~\new_[24752]_  & ~\new_[26316]_ ;
  assign \new_[22482]_  = ~\new_[24596]_  & (~\new_[29020]_  | ~\new_[5973]_ );
  assign \new_[22483]_  = ~\new_[31763]_  | ~\new_[30123]_  | ~\new_[29226]_ ;
  assign \new_[22484]_  = ~\new_[25892]_  & (~\new_[29984]_  | ~\new_[31429]_ );
  assign \new_[22485]_  = ~\new_[26943]_  & ~\new_[24619]_ ;
  assign \new_[22486]_  = ~\new_[31429]_  | ~\new_[26570]_  | ~\new_[29777]_ ;
  assign \new_[22487]_  = ~\new_[26597]_  & ~\new_[26277]_ ;
  assign \new_[22488]_  = ~\new_[31394]_  | ~\new_[27989]_  | ~\new_[27892]_ ;
  assign \new_[22489]_  = ~\new_[27325]_  & ~\new_[24642]_ ;
  assign \new_[22490]_  = \new_[25330]_  & \new_[26410]_ ;
  assign \new_[22491]_  = ~\new_[24770]_  & (~\new_[29904]_  | ~\new_[5900]_ );
  assign \new_[22492]_  = ~\new_[26815]_  & ~\new_[24712]_ ;
  assign \new_[22493]_  = ~\new_[5983]_  | ~\new_[30163]_  | ~\new_[30086]_ ;
  assign \new_[22494]_  = ~\new_[30151]_  | ~\new_[6078]_ ;
  assign \new_[22495]_  = ~\new_[26321]_  & (~\new_[29276]_  | ~\new_[6063]_ );
  assign \new_[22496]_  = ~\new_[29912]_  | ~\new_[28337]_ ;
  assign \new_[22497]_  = ~\new_[31648]_  | ~\new_[30280]_  | ~\new_[28898]_ ;
  assign \new_[22498]_  = \new_[27537]_  & \new_[24612]_ ;
  assign \new_[22499]_  = ~\new_[6269]_  | ~\new_[28502]_  | ~\new_[30732]_ ;
  assign \new_[22500]_  = ~\new_[26394]_  & ~\new_[25254]_ ;
  assign \new_[22501]_  = \new_[27674]_  & \new_[26305]_ ;
  assign \new_[22502]_  = ~\new_[6069]_  | ~\new_[30071]_  | ~\new_[29802]_ ;
  assign \new_[22503]_  = ~\new_[5923]_  | ~\new_[30257]_  | ~\new_[28844]_ ;
  assign \new_[22504]_  = ~\new_[5924]_  | ~\new_[30343]_  | ~\new_[29979]_ ;
  assign \new_[22505]_  = ~\new_[31232]_  | ~\new_[26570]_  | ~\new_[29777]_ ;
  assign \new_[22506]_  = ~\new_[26383]_  & (~\new_[29410]_  | ~\new_[6068]_ );
  assign \new_[22507]_  = ~\new_[26310]_  & (~\new_[29851]_  | ~\new_[6268]_ );
  assign \new_[22508]_  = ~\new_[24542]_  & (~\new_[30016]_  | ~\new_[5907]_ );
  assign \new_[22509]_  = \new_[24688]_  & \new_[26420]_ ;
  assign \new_[22510]_  = ~\new_[5983]_  | ~\new_[30086]_  | ~\new_[28828]_ ;
  assign \new_[22511]_  = ~\new_[5917]_  | ~\new_[30006]_  | ~\new_[28911]_ ;
  assign \new_[22512]_  = ~\new_[5921]_  | ~\new_[29910]_  | ~\new_[28864]_ ;
  assign \new_[22513]_  = ~\new_[26440]_  & (~\new_[28894]_  | ~\new_[6039]_ );
  assign \new_[22514]_  = ~\new_[26163]_  & (~\new_[29623]_  | ~\new_[6077]_ );
  assign \new_[22515]_  = \new_[27695]_  & \new_[26281]_ ;
  assign \new_[22516]_  = ~\new_[26263]_  & (~\new_[28818]_  | ~\new_[6058]_ );
  assign \new_[22517]_  = ~\new_[27337]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[22518]_  = ~\new_[27347]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[22519]_  = ~\new_[5909]_  | ~\new_[28249]_  | ~\new_[28908]_ ;
  assign \new_[22520]_  = ~\new_[28495]_  & ~\new_[26217]_ ;
  assign \new_[22521]_  = ~\new_[26289]_  & (~\new_[29421]_  | ~\new_[6003]_ );
  assign \new_[22522]_  = ~\new_[26293]_  & (~\new_[29151]_  | ~\new_[6006]_ );
  assign \new_[22523]_  = ~\new_[6196]_  | ~\new_[30349]_  | ~\new_[29870]_ ;
  assign \new_[22524]_  = ~\new_[29272]_  | ~\new_[5993]_ ;
  assign \new_[22525]_  = ~\new_[32049]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[22526]_  = ~\new_[30541]_  | ~\new_[6245]_ ;
  assign \new_[22527]_  = ~\new_[26313]_  & (~\new_[29404]_  | ~\new_[5901]_ );
  assign \new_[22528]_  = ~\new_[27781]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[22529]_  = ~\new_[32127]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[22530]_  = ~\new_[32343]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[22531]_  = ~\new_[27855]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[22532]_  = ~\new_[27534]_  & ~\new_[26153]_ ;
  assign \new_[22533]_  = ~\new_[6066]_  | ~\new_[30178]_  | ~\new_[29867]_ ;
  assign \new_[22534]_  = ~\new_[6078]_  | ~\new_[30278]_  | ~\new_[29813]_ ;
  assign \new_[22535]_  = ~\new_[31648]_  | ~\new_[30046]_  | ~\new_[30280]_ ;
  assign \new_[22536]_  = ~\new_[30250]_  | ~\new_[6195]_ ;
  assign \new_[22537]_  = ~\new_[24704]_  & ~\new_[24627]_ ;
  assign \new_[22538]_  = ~\new_[5926]_  | ~\new_[30196]_  | ~\new_[30105]_ ;
  assign \new_[22539]_  = ~\new_[5927]_  | ~\new_[28724]_  | ~\new_[29189]_ ;
  assign \new_[22540]_  = ~\new_[25213]_  & (~\new_[28964]_  | ~\new_[5933]_ );
  assign \new_[22541]_  = ~\new_[31763]_  | ~\new_[30161]_  | ~\new_[30123]_ ;
  assign \new_[22542]_  = ~\new_[24692]_  & (~\new_[29557]_  | ~\new_[5908]_ );
  assign \new_[22543]_  = ~\new_[28229]_  & ~\new_[24776]_ ;
  assign \new_[22544]_  = ~\new_[5978]_  | ~\new_[29943]_  | ~\new_[30005]_ ;
  assign \new_[22545]_  = ~\new_[6094]_  | ~\new_[30019]_  | ~\new_[30104]_ ;
  assign \new_[22546]_  = ~\new_[26379]_  & (~\new_[29900]_  | ~\new_[5894]_ );
  assign \new_[22547]_  = ~\new_[24758]_  & (~\new_[30612]_  | ~\new_[30828]_ );
  assign \new_[22548]_  = ~\new_[24960]_  & (~\new_[30545]_  | ~\new_[30641]_ );
  assign \new_[22549]_  = ~\new_[26467]_  & (~\new_[30713]_  | ~\new_[30603]_ );
  assign \new_[22550]_  = ~\new_[26229]_  & (~\new_[29013]_  | ~\new_[30242]_ );
  assign \new_[22551]_  = ~\new_[26191]_  & (~\new_[29016]_  | ~\new_[30015]_ );
  assign \new_[22552]_  = ~\new_[24555]_  & (~\new_[30711]_  | ~\new_[30499]_ );
  assign \new_[22553]_  = ~\new_[26356]_  & (~\new_[30675]_  | ~\new_[30691]_ );
  assign \new_[22554]_  = ~\new_[28748]_  | ~\new_[6035]_ ;
  assign \new_[22555]_  = ~\new_[26307]_  & (~\new_[30478]_  | ~\new_[30638]_ );
  assign \new_[22556]_  = ~\new_[25182]_  & (~\new_[30780]_  | ~\new_[30667]_ );
  assign \new_[22557]_  = ~\new_[26449]_  & (~\new_[29370]_  | ~\new_[30693]_ );
  assign \new_[22558]_  = ~\new_[25770]_  & (~\new_[30443]_  | ~\new_[30686]_ );
  assign \new_[22559]_  = ~\new_[27658]_  & (~\new_[28829]_  | ~\new_[30198]_ );
  assign \new_[22560]_  = ~\new_[27647]_  & (~\new_[28984]_  | ~\new_[30248]_ );
  assign \new_[22561]_  = ~\new_[26230]_  & (~\new_[29132]_  | ~\new_[30599]_ );
  assign \new_[22562]_  = ~\new_[25775]_  & (~\new_[30501]_  | ~\new_[30635]_ );
  assign \new_[22563]_  = ~\new_[30301]_  | ~\new_[5980]_ ;
  assign \new_[22564]_  = (~\new_[27855]_  | ~\s4_data_i[24] ) & (~\new_[27879]_  | ~\s0_data_i[24] );
  assign \new_[22565]_  = ~\new_[30302]_  | ~\new_[5985]_ ;
  assign \new_[22566]_  = (~\new_[30106]_  | ~\s14_data_i[1] ) & (~\new_[27347]_  | ~\s12_data_i[1] );
  assign \new_[22567]_  = (~\new_[30106]_  | ~\s14_data_i[3] ) & (~\new_[27347]_  | ~\s12_data_i[3] );
  assign \new_[22568]_  = (~\new_[27855]_  | ~\s4_data_i[26] ) & (~\new_[27879]_  | ~\s0_data_i[26] );
  assign \new_[22569]_  = (~\new_[29604]_  | ~\s11_data_i[3] ) & (~\new_[27337]_  | ~\s8_data_i[3] );
  assign \new_[22570]_  = ~\new_[30261]_  | ~\new_[6088]_ ;
  assign \new_[22571]_  = ~\new_[30553]_  | ~\new_[5987]_ ;
  assign \new_[22572]_  = ~\new_[29946]_  | ~\new_[5998]_ ;
  assign \new_[22573]_  = ~\new_[23737]_ ;
  assign \new_[22574]_  = (~\new_[29604]_  | ~\s11_data_i[14] ) & (~\new_[27337]_  | ~\s8_data_i[14] );
  assign \new_[22575]_  = ~\new_[30095]_  | ~\new_[6038]_ ;
  assign \new_[22576]_  = (~\new_[27855]_  | ~\s4_data_i[16] ) & (~\new_[27879]_  | ~\s0_data_i[16] );
  assign \new_[22577]_  = ~\new_[29763]_  & ~\new_[31165]_ ;
  assign \new_[22578]_  = (~\new_[30106]_  | ~\s14_data_i[4] ) & (~\new_[27347]_  | ~\s12_data_i[4] );
  assign \new_[22579]_  = (~\new_[29604]_  | ~\s11_data_i[4] ) & (~\new_[27337]_  | ~\s8_data_i[4] );
  assign \new_[22580]_  = ~\new_[29568]_  | ~\new_[5986]_ ;
  assign \new_[22581]_  = ~\new_[30718]_  | ~\new_[6060]_ ;
  assign \new_[22582]_  = \new_[25617]_  & \new_[25853]_ ;
  assign \new_[22583]_  = ~\new_[30149]_  & ~\new_[31416]_ ;
  assign \new_[22584]_  = (~\new_[27855]_  | ~\s4_data_i[29] ) & (~\new_[27879]_  | ~\s0_data_i[29] );
  assign \new_[22585]_  = (~\new_[27855]_  | ~\s4_data_i[4] ) & (~\new_[27879]_  | ~\s0_data_i[4] );
  assign \new_[22586]_  = ~\new_[30239]_  | ~\new_[5986]_ ;
  assign \new_[22587]_  = ~\new_[30151]_  & ~\new_[30309]_ ;
  assign \new_[22588]_  = (~\new_[27855]_  | ~\s4_data_i[5] ) & (~\new_[27879]_  | ~\s0_data_i[5] );
  assign \new_[22589]_  = (~\new_[30106]_  | ~\s14_data_i[6] ) & (~\new_[27347]_  | ~\s12_data_i[6] );
  assign \new_[22590]_  = (~\new_[29604]_  | ~\s11_data_i[30] ) & (~\new_[27337]_  | ~\s8_data_i[30] );
  assign \new_[22591]_  = (~\new_[30106]_  | ~\s14_data_i[30] ) & (~\new_[27347]_  | ~\s12_data_i[30] );
  assign \new_[22592]_  = ~\new_[30286]_  | ~\new_[6195]_ ;
  assign \new_[22593]_  = (~\new_[29604]_  | ~\s11_data_i[16] ) & (~\new_[27337]_  | ~\s8_data_i[16] );
  assign \new_[22594]_  = ~\new_[30390]_  | ~\new_[5920]_ ;
  assign \new_[22595]_  = (~\new_[30106]_  | ~\s14_data_i[25] ) & (~\new_[27347]_  | ~\s12_data_i[25] );
  assign \new_[22596]_  = ~\new_[29332]_  | ~\new_[29967]_ ;
  assign \new_[22597]_  = (~\new_[29604]_  | ~\s11_data_i[27] ) & (~\new_[27337]_  | ~\s8_data_i[27] );
  assign \new_[22598]_  = (~\new_[30106]_  | ~\s14_data_i[26] ) & (~\new_[27347]_  | ~\s12_data_i[26] );
  assign \new_[22599]_  = (~\new_[27855]_  | ~\s4_data_i[25] ) & (~\new_[27879]_  | ~\s0_data_i[25] );
  assign \new_[22600]_  = (~\new_[29604]_  | ~\s11_data_i[31] ) & (~\new_[27337]_  | ~\s8_data_i[31] );
  assign \new_[22601]_  = (~\new_[30106]_  | ~\s14_data_i[24] ) & (~\new_[27347]_  | ~\s12_data_i[24] );
  assign \new_[22602]_  = (~\new_[29604]_  | ~\s11_data_i[23] ) & (~\new_[27337]_  | ~\s8_data_i[23] );
  assign \new_[22603]_  = (~\new_[27855]_  | ~\s4_data_i[22] ) & (~\new_[27879]_  | ~\s0_data_i[22] );
  assign \new_[22604]_  = (~\new_[27855]_  | ~\s4_data_i[27] ) & (~\new_[27879]_  | ~\s0_data_i[27] );
  assign \new_[22605]_  = (~\new_[29604]_  | ~\s11_data_i[25] ) & (~\new_[27337]_  | ~\s8_data_i[25] );
  assign \new_[22606]_  = (~\new_[30106]_  | ~\s14_data_i[20] ) & (~\new_[27347]_  | ~\s12_data_i[20] );
  assign \new_[22607]_  = (~\new_[29604]_  | ~\s11_data_i[17] ) & (~\new_[27337]_  | ~\s8_data_i[17] );
  assign \new_[22608]_  = ~\new_[29568]_  | ~\new_[6068]_ ;
  assign \new_[22609]_  = (~\new_[27855]_  | ~\s4_data_i[0] ) & (~\new_[27879]_  | ~\s0_data_i[0] );
  assign \new_[22610]_  = (~\new_[30106]_  | ~\s14_data_i[15] ) & (~\new_[27347]_  | ~\s12_data_i[15] );
  assign \new_[22611]_  = (~\new_[30106]_  | ~\s14_data_i[29] ) & (~\new_[27347]_  | ~\s12_data_i[29] );
  assign \new_[22612]_  = (~\new_[29604]_  | ~\s11_data_i[13] ) & (~\new_[27337]_  | ~\s8_data_i[13] );
  assign \new_[22613]_  = ~\new_[30129]_  | ~\new_[6189]_ ;
  assign \new_[22614]_  = (~\new_[27855]_  | ~\s4_data_i[7] ) & (~\new_[27879]_  | ~\s0_data_i[7] );
  assign \new_[22615]_  = ~\new_[28089]_  | ~\new_[6189]_ ;
  assign \new_[22616]_  = (~\new_[29604]_  | ~\s11_data_i[10] ) & (~\new_[27337]_  | ~\s8_data_i[10] );
  assign \new_[22617]_  = (~\new_[30106]_  | ~\s14_data_i[9] ) & (~\new_[27347]_  | ~\s12_data_i[9] );
  assign \new_[22618]_  = ~\new_[28818]_  | ~\new_[29221]_ ;
  assign \new_[22619]_  = (~\new_[30106]_  | ~\s14_data_i[8] ) & (~\new_[27347]_  | ~\s12_data_i[8] );
  assign \new_[22620]_  = (~\new_[29604]_  | ~\s11_data_i[2] ) & (~\new_[27337]_  | ~\s8_data_i[2] );
  assign \new_[22621]_  = (~\new_[27855]_  | ~\s4_data_i[1] ) & (~\new_[27879]_  | ~\s0_data_i[1] );
  assign \new_[22622]_  = (~\new_[30106]_  | ~\s14_data_i[10] ) & (~\new_[27347]_  | ~\s12_data_i[10] );
  assign \new_[22623]_  = (~\new_[29604]_  | ~\s11_data_i[9] ) & (~\new_[27337]_  | ~\s8_data_i[9] );
  assign \new_[22624]_  = (~\new_[27855]_  | ~\s4_data_i[15] ) & (~\new_[27879]_  | ~\s0_data_i[15] );
  assign \new_[22625]_  = (~\new_[27855]_  | ~\s4_data_i[9] ) & (~\new_[27879]_  | ~\s0_data_i[9] );
  assign \new_[22626]_  = (~\new_[27855]_  | ~\s4_data_i[23] ) & (~\new_[27879]_  | ~\s0_data_i[23] );
  assign \new_[22627]_  = (~\new_[30106]_  | ~\s14_data_i[18] ) & (~\new_[27347]_  | ~\s12_data_i[18] );
  assign \new_[22628]_  = ~\new_[23687]_ ;
  assign \new_[22629]_  = (~\new_[29604]_  | ~\s11_data_i[15] ) & (~\new_[27337]_  | ~\s8_data_i[15] );
  assign \new_[22630]_  = (~\new_[27855]_  | ~\s4_data_i[10] ) & (~\new_[27879]_  | ~\s0_data_i[10] );
  assign \new_[22631]_  = (~\new_[29604]_  | ~\s11_data_i[26] ) & (~\new_[27337]_  | ~\s8_data_i[26] );
  assign \new_[22632]_  = \new_[29571]_  | \new_[31862]_ ;
  assign \new_[22633]_  = ~\new_[24065]_ ;
  assign \new_[22634]_  = (~\new_[29604]_  | ~\s11_data_i[24] ) & (~\new_[27337]_  | ~\s8_data_i[24] );
  assign \new_[22635]_  = (~\new_[30106]_  | ~\s14_data_i[28] ) & (~\new_[27347]_  | ~\s12_data_i[28] );
  assign \new_[22636]_  = (~\new_[29604]_  | ~\s11_data_i[6] ) & (~\new_[27337]_  | ~\s8_data_i[6] );
  assign \new_[22637]_  = (~\new_[27855]_  | ~\s4_data_i[30] ) & (~\new_[27879]_  | ~\s0_data_i[30] );
  assign \new_[22638]_  = (~\new_[27855]_  | ~\s4_data_i[12] ) & (~\new_[27879]_  | ~\s0_data_i[12] );
  assign \new_[22639]_  = ~\new_[29830]_  | ~\new_[5988]_ ;
  assign \new_[22640]_  = (~\new_[29604]_  | ~\s11_data_i[1] ) & (~\new_[27337]_  | ~\s8_data_i[1] );
  assign \new_[22641]_  = (~\new_[27855]_  | ~\s4_data_i[13] ) & (~\new_[27879]_  | ~\s0_data_i[13] );
  assign \new_[22642]_  = ~\new_[30591]_  & ~\new_[30840]_ ;
  assign \new_[22643]_  = (~\new_[30106]_  | ~\s14_data_i[23] ) & (~\new_[27347]_  | ~\s12_data_i[23] );
  assign \new_[22644]_  = (~\new_[27855]_  | ~\s4_data_i[28] ) & (~\new_[27879]_  | ~\s0_data_i[28] );
  assign \new_[22645]_  = ~\new_[30204]_  | ~\new_[5830]_ ;
  assign \new_[22646]_  = ~\new_[30569]_  | ~\new_[6212]_ ;
  assign \new_[22647]_  = (~\new_[30106]_  | ~\s14_data_i[2] ) & (~\new_[27347]_  | ~\s12_data_i[2] );
  assign \new_[22648]_  = (~\new_[30106]_  | ~\s14_data_i[27] ) & (~\new_[27347]_  | ~\s12_data_i[27] );
  assign \new_[22649]_  = ~\new_[29962]_  | ~\new_[5987]_ ;
  assign \new_[22650]_  = (~\new_[30106]_  | ~\s14_data_i[14] ) & (~\new_[27347]_  | ~\s12_data_i[14] );
  assign \new_[22651]_  = ~\new_[30235]_  | ~\new_[6065]_ ;
  assign \new_[22652]_  = ~\new_[24097]_ ;
  assign \new_[22653]_  = (~\new_[30106]_  | ~\s14_data_i[16] ) & (~\new_[27347]_  | ~\s12_data_i[16] );
  assign \new_[22654]_  = ~\new_[29962]_  | ~\new_[6213]_ ;
  assign \new_[22655]_  = ~\new_[30204]_  | ~\new_[5972]_ ;
  assign \new_[22656]_  = ~\new_[28864]_  & ~\new_[5904]_ ;
  assign \new_[22657]_  = ~\new_[29069]_  | ~\new_[5972]_ ;
  assign \new_[22658]_  = \new_[29608]_  | \new_[31553]_ ;
  assign \new_[22659]_  = (~\new_[30106]_  | ~\s14_data_i[17] ) & (~\new_[27347]_  | ~\s12_data_i[17] );
  assign \new_[22660]_  = (~\new_[27855]_  | ~\s4_data_i[17] ) & (~\new_[27879]_  | ~\s0_data_i[17] );
  assign \new_[22661]_  = \new_[26065]_  & \new_[24560]_ ;
  assign \new_[22662]_  = (~\new_[30106]_  | ~\s14_data_i[12] ) & (~\new_[27347]_  | ~\s12_data_i[12] );
  assign \new_[22663]_  = (~\new_[29604]_  | ~\s11_data_i[18] ) & (~\new_[27337]_  | ~\s8_data_i[18] );
  assign \new_[22664]_  = (~\new_[29604]_  | ~\s11_data_i[7] ) & (~\new_[27337]_  | ~\s8_data_i[7] );
  assign \new_[22665]_  = (~\new_[27855]_  | ~\s4_data_i[31] ) & (~\new_[27879]_  | ~\s0_data_i[31] );
  assign \new_[22666]_  = (~\new_[27855]_  | ~\s4_data_i[14] ) & (~\new_[27879]_  | ~\s0_data_i[14] );
  assign \new_[22667]_  = ~\new_[28893]_  | ~\new_[6000]_ ;
  assign \new_[22668]_  = (~\new_[27855]_  | ~\s4_data_i[18] ) & (~\new_[27879]_  | ~\s0_data_i[18] );
  assign \new_[22669]_  = (~\new_[30106]_  | ~\s14_data_i[19] ) & (~\new_[27347]_  | ~\s12_data_i[19] );
  assign \new_[22670]_  = (~\new_[29604]_  | ~\s11_data_i[19] ) & (~\new_[27337]_  | ~\s8_data_i[19] );
  assign \new_[22671]_  = ~\new_[30569]_  | ~\new_[6213]_ ;
  assign \new_[22672]_  = (~\new_[27855]_  | ~\s4_data_i[11] ) & (~\new_[27879]_  | ~\s0_data_i[11] );
  assign \new_[22673]_  = (~\new_[27855]_  | ~\s4_data_i[2] ) & (~\new_[27879]_  | ~\s0_data_i[2] );
  assign \new_[22674]_  = (~\new_[27855]_  | ~\s4_data_i[19] ) & (~\new_[27879]_  | ~\s0_data_i[19] );
  assign \new_[22675]_  = \new_[25669]_  & \new_[25656]_ ;
  assign \new_[22676]_  = ~\new_[30327]_  | ~\new_[6047]_ ;
  assign \new_[22677]_  = ~\new_[24980]_  | ~\new_[24983]_ ;
  assign \new_[22678]_  = (~\new_[29604]_  | ~\s11_data_i[20] ) & (~\new_[27337]_  | ~\s8_data_i[20] );
  assign \new_[22679]_  = ~\new_[30620]_  | ~\new_[6270]_ ;
  assign \new_[22680]_  = ~\new_[29773]_  | ~\new_[5988]_ ;
  assign \new_[22681]_  = (~\new_[30106]_  | ~\s14_data_i[21] ) & (~\new_[27347]_  | ~\s12_data_i[21] );
  assign \new_[22682]_  = ~\new_[30757]_  | ~\new_[6048]_ ;
  assign \new_[22683]_  = (~\new_[27855]_  | ~\s4_data_i[6] ) & (~\new_[27879]_  | ~\s0_data_i[6] );
  assign \new_[22684]_  = (~\new_[27855]_  | ~\s4_data_i[21] ) & (~\new_[27879]_  | ~\s0_data_i[21] );
  assign \new_[22685]_  = ~\new_[28835]_  & ~\new_[5898]_ ;
  assign \new_[22686]_  = (~\new_[29604]_  | ~\s11_data_i[28] ) & (~\new_[27337]_  | ~\s8_data_i[28] );
  assign \new_[22687]_  = (~\new_[29604]_  | ~\s11_data_i[22] ) & (~\new_[27337]_  | ~\s8_data_i[22] );
  assign \new_[22688]_  = (~\new_[30106]_  | ~\s14_data_i[22] ) & (~\new_[27347]_  | ~\s12_data_i[22] );
  assign \new_[22689]_  = (~\new_[29604]_  | ~\s11_data_i[21] ) & (~\new_[27337]_  | ~\s8_data_i[21] );
  assign \new_[22690]_  = (~\new_[29604]_  | ~\s11_data_i[12] ) & (~\new_[27337]_  | ~\s8_data_i[12] );
  assign \new_[22691]_  = (~\new_[29604]_  | ~\s11_data_i[0] ) & (~\new_[27337]_  | ~\s8_data_i[0] );
  assign \new_[22692]_  = ~\new_[30064]_  | ~\new_[5971]_ ;
  assign \new_[22693]_  = ~\new_[30620]_  | ~\new_[6079]_ ;
  assign \new_[22694]_  = ~\new_[28918]_  | ~\new_[28989]_ ;
  assign \new_[22695]_  = ~\new_[30327]_  | ~\new_[5971]_ ;
  assign \new_[22696]_  = ~\new_[29455]_  & ~\new_[31724]_ ;
  assign \new_[22697]_  = \new_[29455]_  | \new_[31683]_ ;
  assign \new_[22698]_  = ~\new_[29784]_  | ~\new_[5963]_ ;
  assign \new_[22699]_  = ~\new_[30291]_  | ~\new_[6214]_ ;
  assign \new_[22700]_  = ~\new_[30118]_  | ~\new_[5993]_ ;
  assign \new_[22701]_  = ~\new_[29906]_  | ~\new_[5932]_ ;
  assign \new_[22702]_  = ~\new_[30845]_  | ~\new_[6246]_ ;
  assign \new_[22703]_  = ~\new_[28748]_  | ~\new_[5963]_ ;
  assign \new_[22704]_  = ~\new_[30302]_  | ~\new_[6068]_ ;
  assign \new_[22705]_  = ~\new_[30845]_  | ~\new_[6245]_ ;
  assign \new_[22706]_  = \new_[28930]_  | \new_[31643]_ ;
  assign \new_[22707]_  = ~\new_[30741]_  | ~\new_[5922]_ ;
  assign \new_[22708]_  = ~\new_[28110]_  & ~\new_[31014]_ ;
  assign \new_[22709]_  = ~\new_[30332]_  | ~\new_[6035]_ ;
  assign \new_[22710]_  = ~\new_[30771]_  | ~\new_[6269]_ ;
  assign \new_[22711]_  = ~\new_[30095]_  | ~\new_[5965]_ ;
  assign \new_[22712]_  = ~\new_[30095]_  | ~\new_[6039]_ ;
  assign \new_[22713]_  = ~\new_[29397]_  & ~\new_[30925]_ ;
  assign \new_[22714]_  = ~\new_[29911]_  & ~\new_[31645]_ ;
  assign \new_[22715]_  = ~\new_[29781]_  & ~\new_[31180]_ ;
  assign \new_[22716]_  = ~\new_[30741]_  | ~\new_[5992]_ ;
  assign \new_[22717]_  = ~\new_[30291]_  | ~\new_[6192]_ ;
  assign \new_[22718]_  = ~\new_[29293]_  | ~\new_[6077]_ ;
  assign \new_[22719]_  = \new_[28362]_  & \new_[5968]_ ;
  assign \new_[22720]_  = ~\new_[30067]_  | ~\new_[5969]_ ;
  assign \new_[22721]_  = ~\new_[30261]_  | ~\new_[6003]_ ;
  assign \new_[22722]_  = ~\new_[30118]_  | ~\new_[6077]_ ;
  assign \new_[22723]_  = ~\new_[29189]_  & ~\new_[5906]_ ;
  assign \new_[22724]_  = ~\new_[29650]_  | ~\new_[6065]_ ;
  assign \new_[22725]_  = ~\new_[30048]_  & ~\new_[31042]_ ;
  assign \new_[22726]_  = ~\new_[30746]_  | ~\new_[6214]_ ;
  assign \new_[22727]_  = ~\new_[30746]_  | ~\new_[6192]_ ;
  assign \new_[22728]_  = ~\new_[29773]_  | ~\new_[5919]_ ;
  assign \new_[22729]_  = ~\new_[29880]_  | ~\new_[6203]_ ;
  assign \new_[22730]_  = ~\new_[29915]_  | ~\new_[6090]_ ;
  assign \new_[22731]_  = ~\new_[30064]_  | ~\new_[5913]_ ;
  assign \new_[22732]_  = ~\new_[29960]_  | ~\new_[6005]_ ;
  assign \new_[22733]_  = ~\new_[30064]_  | ~\new_[6047]_ ;
  assign \new_[22734]_  = ~\new_[29952]_  | ~\new_[6047]_ ;
  assign \new_[22735]_  = ~\new_[30167]_  | ~\new_[31121]_ ;
  assign \new_[22736]_  = ~\new_[30762]_  | ~\new_[6048]_ ;
  assign \new_[22737]_  = ~\new_[29985]_  | ~\new_[5931]_ ;
  assign \new_[22738]_  = ~\new_[29771]_  & ~\new_[31039]_ ;
  assign \new_[22739]_  = ~\new_[28089]_  | ~\new_[5990]_ ;
  assign \new_[22740]_  = ~\new_[30118]_  | ~\new_[5994]_ ;
  assign \new_[22741]_  = ~\new_[29825]_  & ~\new_[31108]_ ;
  assign \new_[22742]_  = ~\new_[30301]_  | ~\new_[5979]_ ;
  assign \new_[22743]_  = ~\new_[29950]_  | ~\new_[6046]_ ;
  assign \new_[22744]_  = ~\new_[29789]_  | ~\new_[6006]_ ;
  assign \new_[22745]_  = ~\new_[30648]_  | ~\new_[6046]_ ;
  assign \new_[22746]_  = ~\new_[30204]_  | ~\new_[5973]_ ;
  assign \new_[22747]_  = ~\new_[29293]_  | ~\new_[30839]_ ;
  assign \new_[22748]_  = ~\new_[29069]_  | ~\new_[5973]_ ;
  assign \new_[22749]_  = ~\new_[30746]_  | ~\new_[6071]_ ;
  assign \new_[22750]_  = ~\new_[29918]_  | ~\new_[6185]_ ;
  assign \new_[22751]_  = ~\new_[30502]_  | ~\new_[6090]_ ;
  assign \new_[22752]_  = ~\new_[28968]_  & ~\new_[5897]_ ;
  assign \new_[22753]_  = ~\new_[30168]_  | ~\new_[6044]_ ;
  assign \new_[22754]_  = ~\new_[30733]_  | ~\new_[6052]_ ;
  assign \new_[22755]_  = ~\new_[29854]_  | ~\new_[5980]_ ;
  assign \new_[22756]_  = ~\new_[29965]_  | ~\new_[5982]_ ;
  assign \new_[22757]_  = ~\new_[29919]_  | ~\new_[5972]_ ;
  assign \new_[22758]_  = ~\new_[30168]_  | ~\new_[5968]_ ;
  assign \new_[22759]_  = ~\new_[29568]_  | ~\new_[5985]_ ;
  assign \new_[22760]_  = ~\new_[30167]_  | ~\new_[31491]_ ;
  assign \new_[22761]_  = ~\new_[29883]_  | ~\new_[6183]_ ;
  assign \new_[22762]_  = ~\new_[30301]_  | ~\new_[6058]_ ;
  assign \new_[22763]_  = ~\new_[30771]_  | ~\new_[6082]_ ;
  assign \new_[22764]_  = ~\new_[30438]_  | ~\new_[5922]_ ;
  assign \new_[22765]_  = ~\new_[28893]_  | ~\new_[6185]_ ;
  assign \new_[22766]_  = ~\new_[30315]_  | ~\new_[6081]_ ;
  assign \new_[22767]_  = ~\new_[29830]_  | ~\new_[5919]_ ;
  assign \new_[22768]_  = ~\new_[28893]_  | ~\new_[5999]_ ;
  assign \new_[22769]_  = ~\new_[29112]_  & ~\new_[5896]_ ;
  assign \new_[22770]_  = ~\new_[30741]_  | ~\new_[5991]_ ;
  assign \new_[22771]_  = ~\new_[30055]_  | ~\new_[6000]_ ;
  assign \new_[22772]_  = ~\new_[29893]_  & ~\new_[31787]_ ;
  assign \new_[22773]_  = ~\new_[30413]_  | ~\new_[6068]_ ;
  assign \new_[22774]_  = ~\new_[30569]_  | ~\new_[5987]_ ;
  assign \new_[22775]_  = ~\new_[29830]_  | ~\new_[5920]_ ;
  assign \new_[22776]_  = ~\new_[29965]_  | ~\new_[6063]_ ;
  assign \new_[22777]_  = ~\new_[30425]_  | ~\new_[5966]_ ;
  assign \new_[22778]_  = ~\new_[29966]_  | ~\new_[5965]_ ;
  assign \new_[22779]_  = ~\new_[29981]_  | ~\new_[5966]_ ;
  assign \new_[22780]_  = \new_[30059]_  & \new_[5994]_ ;
  assign \new_[22781]_  = ~\new_[30170]_  | ~\new_[6085]_ ;
  assign \new_[22782]_  = ~\new_[30420]_  | ~\new_[5966]_ ;
  assign \new_[22783]_  = ~\new_[30413]_  | ~\new_[5986]_ ;
  assign \new_[22784]_  = \new_[29981]_  & \new_[6176]_ ;
  assign \new_[22785]_  = \new_[28331]_  & \new_[6176]_ ;
  assign \new_[22786]_  = ~\new_[29809]_  | ~\new_[6077]_ ;
  assign \new_[22787]_  = ~\new_[29955]_  | ~\new_[6081]_ ;
  assign \new_[22788]_  = ~\new_[30788]_  | ~\new_[5922]_ ;
  assign \new_[22789]_  = ~\new_[30216]_  | ~\new_[6060]_ ;
  assign \new_[22790]_  = ~\new_[30286]_  | ~\new_[6060]_ ;
  assign \new_[22791]_  = ~\new_[27997]_  & ~\new_[31140]_ ;
  assign \new_[22792]_  = ~\new_[30101]_  | ~\new_[5920]_ ;
  assign \new_[22793]_  = ~\new_[28856]_  | ~\new_[5990]_ ;
  assign \new_[22794]_  = ~\new_[29571]_  & ~\new_[31140]_ ;
  assign \new_[22795]_  = \new_[28884]_  & \new_[6001]_ ;
  assign \new_[22796]_  = ~\new_[30168]_  | ~\new_[5969]_ ;
  assign \new_[22797]_  = ~\new_[29952]_  | ~\new_[5971]_ ;
  assign \new_[22798]_  = ~\new_[30400]_  | ~\new_[5998]_ ;
  assign \new_[22799]_  = ~\new_[30214]_  | ~\new_[5965]_ ;
  assign \new_[22800]_  = ~\new_[30652]_  | ~\new_[5929]_ ;
  assign \new_[22801]_  = \new_[30216]_  & \new_[6059]_ ;
  assign \new_[22802]_  = ~\new_[29809]_  | ~\new_[5993]_ ;
  assign \new_[22803]_  = \new_[29950]_  & \new_[6204]_ ;
  assign \new_[22804]_  = ~\new_[29854]_  | ~\new_[6058]_ ;
  assign \new_[22805]_  = ~\new_[30250]_  | ~\new_[6060]_ ;
  assign \new_[22806]_  = \new_[29271]_  | \new_[31608]_ ;
  assign \new_[22807]_  = ~\new_[29773]_  | ~\new_[5920]_ ;
  assign \new_[22808]_  = ~\new_[30051]_  | ~\new_[6053]_ ;
  assign \new_[22809]_  = ~\new_[30302]_  | ~\new_[5986]_ ;
  assign \new_[22810]_  = ~\new_[29271]_  & ~\new_[31014]_ ;
  assign \new_[22811]_  = ~\new_[28908]_  & ~\new_[5895]_ ;
  assign \new_[22812]_  = ~\new_[29915]_  | ~\new_[6183]_ ;
  assign \new_[22813]_  = ~\new_[30845]_  | ~\new_[6203]_ ;
  assign \new_[22814]_  = ~\new_[30051]_  | ~\new_[6052]_ ;
  assign \new_[22815]_  = ~\new_[28911]_  & ~\new_[5902]_ ;
  assign \new_[22816]_  = ~\new_[30706]_  | ~\new_[6217]_ ;
  assign \new_[22817]_  = ~\new_[28844]_  & ~\new_[5905]_ ;
  assign \new_[22818]_  = ~\new_[30584]_  | ~\new_[6095]_ ;
  assign \new_[22819]_  = \new_[29550]_  | \new_[31669]_ ;
  assign \new_[22820]_  = ~\new_[30332]_  | ~\new_[5963]_ ;
  assign \new_[22821]_  = ~\new_[29883]_  | ~\new_[6090]_ ;
  assign \new_[22822]_  = ~\new_[29985]_  | ~\new_[6088]_ ;
  assign \new_[22823]_  = ~\new_[30584]_  | ~\new_[6217]_ ;
  assign \new_[22824]_  = ~\new_[28748]_  | ~\new_[5964]_ ;
  assign \new_[22825]_  = ~\new_[29650]_  | ~\new_[6273]_ ;
  assign \new_[22826]_  = ~\new_[29952]_  | ~\new_[5913]_ ;
  assign \new_[22827]_  = ~\new_[29918]_  | ~\new_[6000]_ ;
  assign \new_[22828]_  = ~\new_[29633]_  & ~\new_[5903]_ ;
  assign \new_[22829]_  = ~\new_[30715]_  | ~\new_[6085]_ ;
  assign \new_[22830]_  = ~\new_[29003]_  & ~\new_[31665]_ ;
  assign \new_[22831]_  = ~\new_[30101]_  | ~\new_[5988]_ ;
  assign \new_[22832]_  = ~\new_[30771]_  | ~\new_[6085]_ ;
  assign \new_[22833]_  = ~\new_[29608]_  & ~\new_[31421]_ ;
  assign \new_[22834]_  = ~\new_[30737]_  | ~\new_[6085]_ ;
  assign \new_[22835]_  = ~\new_[30736]_  | ~\new_[6245]_ ;
  assign \new_[22836]_  = ~\new_[29985]_  | ~\new_[6003]_ ;
  assign \new_[22837]_  = ~\new_[30466]_  | ~\new_[5995]_ ;
  assign \new_[22838]_  = ~\new_[29069]_  | ~\new_[5830]_ ;
  assign \new_[22839]_  = ~\new_[29293]_  | ~\new_[5993]_ ;
  assign \new_[22840]_  = ~\new_[29906]_  | ~\new_[6005]_ ;
  assign \new_[22841]_  = ~\new_[29789]_  | ~\new_[6005]_ ;
  assign \new_[22842]_  = ~\new_[29906]_  | ~\new_[6006]_ ;
  assign \new_[22843]_  = ~\new_[30584]_  | ~\new_[6007]_ ;
  assign \new_[22844]_  = ~\new_[30762]_  | ~\new_[6206]_ ;
  assign \new_[22845]_  = ~\new_[30261]_  | ~\new_[5931]_ ;
  assign \new_[22846]_  = ~\new_[30677]_  & ~\new_[30682]_ ;
  assign \new_[22847]_  = ~\new_[23569]_ ;
  assign \new_[22848]_  = ~\new_[29130]_  | ~\new_[28371]_ ;
  assign \new_[22849]_  = ~\new_[30114]_  | ~\new_[5905]_ ;
  assign \new_[22850]_  = ~\new_[29583]_  | ~\new_[29038]_ ;
  assign \new_[22851]_  = ~\new_[29151]_  | ~\new_[28850]_ ;
  assign \new_[22852]_  = ~\new_[29077]_  & ~\new_[31400]_ ;
  assign \new_[22853]_  = ~\new_[29907]_  | ~\new_[5910]_ ;
  assign \new_[22854]_  = ~\new_[30149]_  | ~\new_[29386]_ ;
  assign \new_[22855]_  = ~\new_[30128]_  | ~\new_[30161]_ ;
  assign \new_[22856]_  = ~\new_[23417]_ ;
  assign \new_[22857]_  = ~\new_[29029]_  | ~\new_[28845]_ ;
  assign \new_[22858]_  = ~\new_[30185]_  | ~\new_[31438]_ ;
  assign \new_[22859]_  = ~\new_[30033]_  | ~\new_[6196]_ ;
  assign \new_[22860]_  = \new_[28249]_  & \new_[30030]_ ;
  assign \new_[22861]_  = ~\new_[23126]_ ;
  assign \new_[22862]_  = ~\new_[30174]_  | ~\new_[5970]_ ;
  assign \new_[22863]_  = ~\new_[30038]_  & ~\new_[30185]_ ;
  assign \new_[22864]_  = ~\new_[30399]_  | ~\new_[6087]_ ;
  assign \new_[22865]_  = ~\new_[30568]_  & ~\new_[30688]_ ;
  assign \new_[22866]_  = ~\new_[30309]_  | ~\new_[6079]_ ;
  assign \new_[22867]_  = ~\new_[24273]_ ;
  assign \new_[22868]_  = ~\new_[30114]_  & ~\new_[30008]_ ;
  assign \new_[22869]_  = ~\new_[30767]_  | ~\new_[30623]_ ;
  assign \new_[22870]_  = ~\new_[24286]_ ;
  assign \new_[22871]_  = ~\new_[30062]_  | ~\new_[5921]_ ;
  assign \new_[22872]_  = ~\new_[30029]_  | ~\new_[6061]_ ;
  assign \new_[22873]_  = ~\new_[30540]_  & ~\new_[30566]_ ;
  assign \new_[22874]_  = ~\new_[29831]_  | ~\new_[29212]_ ;
  assign \new_[22875]_  = ~\new_[30326]_  & ~\new_[28888]_ ;
  assign \new_[22876]_  = ~\new_[30201]_  | ~\new_[6184]_ ;
  assign \new_[22877]_  = ~\new_[24300]_ ;
  assign \new_[22878]_  = ~\new_[29571]_  | ~\new_[28007]_ ;
  assign \new_[22879]_  = ~\new_[29452]_  | ~\new_[30884]_ ;
  assign \new_[22880]_  = ~\new_[23181]_ ;
  assign \new_[22881]_  = ~\new_[29792]_  | ~\new_[5924]_ ;
  assign \new_[22882]_  = ~\new_[29781]_  | ~\new_[30600]_ ;
  assign \new_[22883]_  = ~\new_[29647]_  & ~\new_[6079]_ ;
  assign \new_[22884]_  = ~\new_[30662]_  & ~\new_[30637]_ ;
  assign \new_[22885]_  = ~\new_[29908]_  | ~\new_[5911]_ ;
  assign \new_[22886]_  = \new_[28070]_  & \new_[30057]_ ;
  assign \new_[22887]_  = ~\new_[28278]_  | ~\new_[30129]_ ;
  assign \new_[22888]_  = ~\new_[30029]_  & ~\new_[30651]_ ;
  assign \new_[22889]_  = ~\new_[30304]_  | ~\new_[5903]_ ;
  assign \new_[22890]_  = ~\new_[29765]_  | ~\new_[5912]_ ;
  assign \new_[22891]_  = ~\new_[23163]_ ;
  assign \new_[22892]_  = ~\new_[29907]_  & ~\new_[30287]_ ;
  assign \new_[22893]_  = ~\new_[28284]_  | ~\new_[5912]_ ;
  assign \new_[22894]_  = ~\new_[30225]_  | ~\new_[6215]_ ;
  assign \new_[22895]_  = ~\new_[30148]_  | ~\new_[31763]_ ;
  assign \new_[22896]_  = ~\new_[29505]_  | ~\new_[29225]_ ;
  assign \new_[22897]_  = ~\new_[29886]_  & ~\new_[5929]_ ;
  assign \new_[22898]_  = ~\new_[30127]_  | ~\new_[6074]_ ;
  assign \new_[22899]_  = ~\new_[23154]_ ;
  assign \new_[22900]_  = ~\new_[23152]_ ;
  assign \new_[22901]_  = ~\new_[30245]_  | ~\new_[5909]_ ;
  assign \new_[22902]_  = ~\new_[29783]_  & ~\new_[6048]_ ;
  assign \new_[22903]_  = ~\new_[30267]_  | ~\new_[5923]_ ;
  assign \new_[22904]_  = ~\new_[29381]_  | ~\new_[28880]_ ;
  assign \new_[22905]_  = ~\new_[28007]_  | ~\new_[28280]_ ;
  assign \new_[22906]_  = ~\new_[30129]_  | ~\new_[5990]_ ;
  assign \new_[22907]_  = ~\new_[30304]_  | ~\new_[5918]_ ;
  assign \new_[22908]_  = ~\new_[30268]_  | ~\new_[5914]_ ;
  assign \new_[22909]_  = ~\new_[29701]_  | ~\new_[28535]_ ;
  assign \new_[22910]_  = ~\new_[30024]_  | ~\new_[5906]_ ;
  assign \new_[22911]_  = ~\new_[30275]_  & ~\new_[29916]_ ;
  assign \new_[22912]_  = ~\new_[28057]_  | ~\new_[30608]_ ;
  assign \new_[22913]_  = ~\new_[28110]_  | ~\new_[28870]_ ;
  assign \new_[22914]_  = ~\new_[30076]_  | ~\new_[5923]_ ;
  assign \new_[22915]_  = ~\new_[30212]_  & ~\new_[30069]_ ;
  assign \new_[22916]_  = ~\new_[29598]_  | ~\new_[31440]_ ;
  assign \new_[22917]_  = ~\new_[30223]_  | ~\new_[29943]_ ;
  assign \new_[22918]_  = ~\new_[28371]_  | ~\new_[29455]_ ;
  assign \new_[22919]_  = ~\new_[29763]_  | ~\new_[30255]_ ;
  assign \new_[22920]_  = ~\new_[23121]_ ;
  assign \new_[22921]_  = ~\new_[23118]_ ;
  assign \new_[22922]_  = ~\new_[29774]_  | ~\new_[5908]_ ;
  assign \new_[22923]_  = ~\new_[30275]_  | ~\new_[5989]_ ;
  assign \new_[22924]_  = ~\new_[30176]_  | ~\new_[5901]_ ;
  assign \new_[22925]_  = ~\new_[29914]_  | ~\new_[5902]_ ;
  assign \new_[22926]_  = ~\new_[23110]_ ;
  assign \new_[22927]_  = ~\new_[30336]_  & ~\new_[30174]_ ;
  assign \new_[22928]_  = ~\new_[29452]_  & ~\new_[6197]_ ;
  assign \new_[22929]_  = ~\new_[30148]_  | ~\new_[5908]_ ;
  assign \new_[22930]_  = ~\new_[29771]_  | ~\new_[29782]_ ;
  assign \new_[22931]_  = ~\new_[24972]_  | ~\new_[28370]_ ;
  assign \new_[22932]_  = ~\new_[30032]_  | ~\new_[6080]_ ;
  assign \new_[22933]_  = ~\new_[30234]_  | ~\new_[6056]_ ;
  assign \new_[22934]_  = ~\new_[23102]_ ;
  assign \new_[22935]_  = ~\new_[29611]_  & ~\new_[6186]_ ;
  assign \new_[22936]_  = ~\new_[30151]_  | ~\new_[6270]_ ;
  assign \new_[22937]_  = ~\new_[30138]_  & ~\new_[5995]_ ;
  assign \new_[22938]_  = ~\new_[24898]_  | ~\new_[30084]_ ;
  assign \new_[22939]_  = ~\new_[23093]_ ;
  assign \new_[22940]_  = ~\new_[30174]_  | ~\new_[6199]_ ;
  assign \new_[22941]_  = ~\new_[30024]_  | ~\new_[5927]_ ;
  assign \new_[22942]_  = ~\new_[29410]_  | ~\new_[29082]_ ;
  assign \new_[22943]_  = ~\new_[30033]_  | ~\new_[6057]_ ;
  assign \new_[22944]_  = ~\new_[30287]_  | ~\new_[6037]_ ;
  assign \new_[22945]_  = ~\new_[30344]_  & ~\new_[5980]_ ;
  assign \new_[22946]_  = ~\new_[29765]_  | ~\new_[5897]_ ;
  assign \new_[22947]_  = ~\new_[29853]_  | ~\new_[6174]_ ;
  assign \new_[22948]_  = ~\new_[30755]_  | ~\new_[31499]_ ;
  assign \new_[22949]_  = ~\new_[30287]_  | ~\new_[5910]_ ;
  assign \new_[22950]_  = ~\new_[29997]_  & ~\new_[30445]_ ;
  assign \new_[22951]_  = ~\new_[28806]_  | ~\new_[30432]_ ;
  assign \new_[22952]_  = ~\new_[28204]_  & ~\new_[29699]_ ;
  assign \new_[22953]_  = ~\new_[30309]_  | ~\new_[6270]_ ;
  assign \new_[22954]_  = ~\new_[30442]_  | ~\new_[31045]_ ;
  assign \new_[22955]_  = ~\new_[26736]_  | ~\new_[24607]_ ;
  assign \new_[22956]_  = ~\new_[28535]_  | ~\new_[5929]_ ;
  assign \new_[22957]_  = ~\new_[30109]_  & ~\new_[26563]_ ;
  assign \new_[22958]_  = ~\new_[29077]_  | ~\new_[6069]_ ;
  assign \new_[22959]_  = ~\new_[30333]_  & ~\new_[6088]_ ;
  assign \new_[22960]_  = ~\new_[24529]_ ;
  assign \new_[22961]_  = ~\new_[28397]_  & ~\new_[29909]_ ;
  assign \new_[22962]_  = ~\new_[29916]_  & ~\new_[24759]_ ;
  assign \new_[22963]_  = ~\new_[29055]_  & ~\new_[6037]_ ;
  assign \new_[22964]_  = ~\new_[28866]_  & ~\new_[5969]_ ;
  assign \new_[22965]_  = ~\new_[30375]_  | ~\new_[6069]_ ;
  assign \new_[22966]_  = ~\new_[30375]_  & ~\new_[30063]_ ;
  assign \new_[22967]_  = ~\new_[24388]_ ;
  assign \new_[22968]_  = ~\new_[29647]_  | ~\new_[6078]_ ;
  assign \new_[22969]_  = ~\new_[30629]_  & ~\new_[30747]_ ;
  assign \new_[22970]_  = ~\new_[29997]_  | ~\new_[5928]_ ;
  assign \new_[22971]_  = ~\new_[29589]_  | ~\new_[30158]_ ;
  assign \new_[22972]_  = ~\new_[29145]_  | ~\new_[29506]_ ;
  assign \new_[22973]_  = ~\new_[29810]_  & ~\new_[30109]_ ;
  assign \new_[22974]_  = ~\new_[30663]_  & ~\new_[28397]_ ;
  assign \new_[22975]_  = ~\new_[30063]_  | ~\new_[31400]_ ;
  assign \new_[22976]_  = ~\new_[30564]_  | ~\new_[6050]_ ;
  assign \new_[22977]_  = ~\new_[30176]_  | ~\new_[6062]_ ;
  assign \new_[22978]_  = ~\new_[24512]_ ;
  assign \new_[22979]_  = ~\new_[30399]_  | ~\new_[5907]_ ;
  assign \new_[22980]_  = ~\new_[24505]_ ;
  assign \new_[22981]_  = ~\new_[30579]_  | ~\new_[29210]_ ;
  assign \new_[22982]_  = ~\new_[28595]_  | ~\new_[30101]_ ;
  assign \new_[22983]_  = ~\new_[30542]_  | ~\new_[6049]_ ;
  assign \new_[22984]_  = ~\new_[29916]_  | ~\new_[5989]_ ;
  assign \new_[22985]_  = ~\new_[30053]_  | ~\new_[5902]_ ;
  assign \new_[22986]_  = ~\new_[29908]_  | ~\new_[5896]_ ;
  assign \new_[22987]_  = ~\new_[24413]_ ;
  assign \new_[22988]_  = ~\new_[28215]_  | ~\new_[30680]_ ;
  assign \new_[22989]_  = ~\new_[30620]_  | ~\new_[6078]_ ;
  assign \new_[22990]_  = ~\new_[30581]_  & ~\new_[30684]_ ;
  assign \new_[22991]_  = ~\new_[29889]_  | ~\new_[6050]_ ;
  assign \new_[22992]_  = ~\new_[29656]_  & ~\new_[5990]_ ;
  assign \new_[22993]_  = ~\new_[29940]_  | ~\new_[6062]_ ;
  assign \new_[22994]_  = ~\new_[29792]_  | ~\new_[5925]_ ;
  assign \new_[22995]_  = ~\new_[29889]_  & ~\new_[30564]_ ;
  assign \new_[22996]_  = ~\new_[28285]_  | ~\new_[29355]_ ;
  assign \new_[22997]_  = ~\new_[30148]_  | ~\new_[6091]_ ;
  assign \new_[22998]_  = ~\new_[24405]_ ;
  assign \new_[22999]_  = ~\new_[24408]_ ;
  assign \new_[23000]_  = ~\new_[30083]_  & ~\new_[6065]_ ;
  assign \new_[23001]_  = ~\new_[29623]_  | ~\new_[29061]_ ;
  assign \new_[23002]_  = ~\new_[30445]_  & ~\new_[29611]_ ;
  assign \new_[23003]_  = ~\new_[30062]_  | ~\new_[5904]_ ;
  assign \new_[23004]_  = ~\new_[24508]_ ;
  assign \new_[23005]_  = ~\new_[30542]_  | ~\new_[6050]_ ;
  assign \new_[23006]_  = ~\new_[30751]_  | ~\new_[28188]_ ;
  assign \new_[23007]_  = ~\new_[28877]_  | ~\new_[29171]_ ;
  assign \new_[23008]_  = ~\new_[29853]_  | ~\new_[6033]_ ;
  assign \new_[23009]_  = ~\new_[30099]_  | ~\new_[30295]_ ;
  assign \new_[23010]_  = ~\new_[30109]_  | ~\new_[6043]_ ;
  assign \new_[23011]_  = ~\new_[30048]_  | ~\new_[30636]_ ;
  assign \new_[23012]_  = ~\new_[29913]_  & ~\new_[6085]_ ;
  assign \new_[23013]_  = ~\new_[29907]_  | ~\new_[6040]_ ;
  assign \new_[23014]_  = ~\new_[30053]_  & ~\new_[30319]_ ;
  assign \new_[23015]_  = ~\new_[28894]_  | ~\new_[29219]_ ;
  assign \new_[23016]_  = ~\new_[24428]_ ;
  assign \new_[23017]_  = ~\new_[24430]_ ;
  assign \new_[23018]_  = ~\new_[30035]_  | ~\new_[30163]_ ;
  assign \new_[23019]_  = ~\new_[28317]_  | ~\new_[5970]_ ;
  assign \new_[23020]_  = ~\new_[30287]_  & ~\new_[29055]_ ;
  assign \new_[23021]_  = ~\new_[29853]_  | ~\new_[6034]_ ;
  assign \new_[23022]_  = ~\new_[30660]_  & ~\new_[30663]_ ;
  assign \new_[23023]_  = ~\new_[30126]_  & ~\new_[5998]_ ;
  assign \new_[23024]_  = ~\new_[24431]_ ;
  assign \new_[23025]_  = ~\new_[30185]_  | ~\new_[31422]_ ;
  assign \new_[23026]_  = ~\new_[28284]_  | ~\new_[6045]_ ;
  assign \new_[23027]_  = ~\new_[30399]_  | ~\new_[31648]_ ;
  assign \new_[23028]_  = ~\new_[29892]_  & ~\new_[6192]_ ;
  assign \new_[23029]_  = ~\new_[30755]_  | ~\new_[6215]_ ;
  assign \new_[23030]_  = ~\new_[30201]_  | ~\new_[6215]_ ;
  assign \new_[23031]_  = ~\new_[29569]_  | ~\new_[29563]_ ;
  assign \new_[23032]_  = ~\new_[24901]_  | ~\new_[26418]_ ;
  assign \new_[23033]_  = ~\new_[30267]_  | ~\new_[5905]_ ;
  assign \new_[23034]_  = ~\new_[30268]_  | ~\new_[5898]_ ;
  assign \new_[23035]_  = ~\new_[30294]_  & ~\new_[6060]_ ;
  assign \new_[23036]_  = ~\new_[30234]_  | ~\new_[5978]_ ;
  assign \new_[23037]_  = ~\new_[29893]_  | ~\new_[29912]_ ;
  assign \new_[23038]_  = ~\new_[29699]_  & ~\new_[6076]_ ;
  assign \new_[23039]_  = ~\new_[30225]_  | ~\new_[31499]_ ;
  assign \new_[23040]_  = ~\new_[24444]_ ;
  assign \new_[23041]_  = ~\new_[28031]_  | ~\new_[5926]_ ;
  assign \new_[23042]_  = ~\new_[30231]_  | ~\new_[6202]_ ;
  assign \new_[23043]_  = ~\new_[30326]_  | ~\new_[31157]_ ;
  assign \new_[23044]_  = ~\new_[28031]_  | ~\new_[5933]_ ;
  assign \new_[23045]_  = ~\new_[23547]_ ;
  assign \new_[23046]_  = ~\new_[23517]_ ;
  assign \new_[23047]_  = ~\new_[29940]_  | ~\new_[5983]_ ;
  assign \new_[23048]_  = ~\new_[24453]_ ;
  assign \new_[23049]_  = ~\new_[29940]_  | ~\new_[5901]_ ;
  assign \new_[23050]_  = ~\new_[27997]_  | ~\new_[29685]_ ;
  assign \new_[23051]_  = ~\new_[30743]_  | ~\new_[6034]_ ;
  assign \new_[23052]_  = ~\new_[28031]_  | ~\new_[6080]_ ;
  assign \new_[23053]_  = ~\new_[23245]_ ;
  assign \new_[23054]_  = ~\new_[29889]_  | ~\new_[31712]_ ;
  assign \new_[23055]_  = ~\new_[30618]_  & ~\new_[30632]_ ;
  assign \new_[23056]_  = ~\new_[29421]_  | ~\new_[29040]_ ;
  assign \new_[23057]_  = ~\new_[29931]_  | ~\new_[5898]_ ;
  assign \new_[23058]_  = ~\new_[29911]_  | ~\new_[30020]_ ;
  assign \new_[23059]_  = ~\new_[23185]_ ;
  assign \new_[23060]_  = ~\new_[24468]_ ;
  assign \new_[23061]_  = ~\new_[30212]_  | ~\new_[5903]_ ;
  assign \new_[23062]_  = ~\new_[28836]_  | ~\new_[29032]_ ;
  assign \new_[23063]_  = ~\new_[30743]_  | ~\new_[6174]_ ;
  assign \new_[23064]_  = ~\new_[24474]_ ;
  assign \new_[23065]_  = ~\new_[30442]_  | ~\new_[6093]_ ;
  assign \new_[23066]_  = ~\new_[29851]_  | ~\new_[28188]_ ;
  assign \new_[23067]_  = ~\new_[24492]_ ;
  assign \new_[23068]_  = ~\new_[29931]_  & ~\new_[30249]_ ;
  assign \new_[23069]_  = ~\new_[30564]_  | ~\new_[6049]_ ;
  assign \new_[23070]_  = (~\new_[30106]_  | ~\s14_data_i[13] ) & (~\new_[27347]_  | ~\s12_data_i[13] );
  assign \new_[23071]_  = ~\new_[23097]_ ;
  assign \new_[23072]_  = ~\new_[23176]_ ;
  assign \new_[23073]_  = ~\new_[30598]_  | ~\new_[6174]_ ;
  assign \new_[23074]_  = ~\new_[30336]_  & ~\new_[29251]_ ;
  assign \new_[23075]_  = ~\new_[25214]_  & ~\new_[30276]_ ;
  assign \new_[23076]_  = ~\new_[24378]_ ;
  assign \new_[23077]_  = ~\new_[29974]_  | ~\new_[28285]_ ;
  assign \new_[23078]_  = ~\new_[26321]_ ;
  assign \new_[23079]_  = ~\new_[28118]_  & ~\new_[27033]_ ;
  assign \new_[23080]_  = ~\new_[27601]_  | ~\new_[30410]_ ;
  assign \new_[23081]_  = ~\new_[29221]_  | ~\new_[28684]_ ;
  assign \new_[23082]_  = ~\new_[24541]_ ;
  assign \new_[23083]_  = ~\new_[27685]_  | ~\new_[28039]_ ;
  assign \new_[23084]_  = ~\new_[26316]_ ;
  assign \new_[23085]_  = ~\new_[30613]_  | ~\new_[30136]_ ;
  assign \new_[23086]_  = ~\new_[24554]_ ;
  assign \new_[23087]_  = ~\new_[26439]_ ;
  assign \new_[23088]_  = ~\new_[24561]_ ;
  assign \new_[23089]_  = ~\new_[24830]_ ;
  assign \new_[23090]_  = ~\new_[28918]_  | ~\new_[29501]_ ;
  assign \new_[23091]_  = ~\new_[26469]_ ;
  assign \new_[23092]_  = ~\new_[24568]_ ;
  assign \new_[23093]_  = ~\new_[30650]_  | ~\new_[26563]_ ;
  assign \new_[23094]_  = ~\new_[24573]_ ;
  assign \new_[23095]_  = ~\new_[30651]_  | ~\new_[6211]_ ;
  assign \new_[23096]_  = ~\new_[26310]_ ;
  assign \new_[23097]_  = ~\new_[27715]_  | ~\new_[30952]_ ;
  assign \new_[23098]_  = ~\new_[30445]_  | ~\new_[5928]_ ;
  assign \new_[23099]_  = ~\new_[26308]_ ;
  assign \new_[23100]_  = (~\new_[28223]_  | ~\s7_data_i[25] ) & (~\new_[28767]_  | ~\s6_data_i[25] );
  assign \new_[23101]_  = ~\new_[24598]_ ;
  assign \new_[23102]_  = ~\new_[29589]_  & ~\new_[29809]_ ;
  assign \new_[23103]_  = ~\new_[26647]_  | ~\new_[31423]_ ;
  assign \new_[23104]_  = ~\new_[29192]_  | ~\new_[28989]_ ;
  assign \new_[23105]_  = ~\new_[26251]_ ;
  assign \new_[23106]_  = \new_[29528]_  & \new_[30638]_ ;
  assign \new_[23107]_  = ~\new_[26259]_ ;
  assign \new_[23108]_  = ~\new_[27463]_  & ~\new_[30230]_ ;
  assign \new_[23109]_  = ~\new_[26465]_ ;
  assign \new_[23110]_  = ~\new_[28999]_  & ~\new_[28007]_ ;
  assign \new_[23111]_  = (~\new_[28392]_  | ~\s4_data_i[31] ) & (~\new_[29349]_  | ~\s0_data_i[31] );
  assign \new_[23112]_  = ~\new_[32161]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[23113]_  = ~\new_[26299]_ ;
  assign \new_[23114]_  = ~\new_[28188]_  | ~\new_[28935]_ ;
  assign \new_[23115]_  = ~\new_[24613]_ ;
  assign \new_[23116]_  = (~\new_[28714]_  | ~\s5_data_i[23] ) & (~\new_[30709]_  | ~\s3_data_i[23] );
  assign \new_[23117]_  = ~\new_[29042]_  | ~\new_[28926]_ ;
  assign \new_[23118]_  = ~\new_[29421]_  | ~\new_[29672]_ ;
  assign \new_[23119]_  = ~\new_[29865]_  | ~\new_[5978]_ ;
  assign \new_[23120]_  = ~\new_[26293]_ ;
  assign \new_[23121]_  = ~\new_[29020]_  | ~\new_[28232]_ ;
  assign \new_[23122]_  = ~\new_[26289]_ ;
  assign \new_[23123]_  = ~\new_[26285]_ ;
  assign \new_[23124]_  = ~\new_[30521]_  & ~\new_[30607]_ ;
  assign \new_[23125]_  = ~\new_[29772]_  | ~\new_[31648]_ ;
  assign \new_[23126]_  = ~\new_[30158]_  | ~\new_[28985]_ ;
  assign \new_[23127]_  = ~\new_[26277]_ ;
  assign \new_[23128]_  = ~\new_[30404]_  | ~\new_[5968]_ ;
  assign \new_[23129]_  = ~\new_[24653]_ ;
  assign \new_[23130]_  = (~\new_[28313]_  | ~\s7_data_i[20] ) & (~\new_[29707]_  | ~\s6_data_i[20] );
  assign \new_[23131]_  = ~\new_[28939]_  | ~\new_[29227]_ ;
  assign \new_[23132]_  = ~\new_[30038]_  | ~\new_[31440]_ ;
  assign \new_[23133]_  = (~\new_[28714]_  | ~\s5_data_i[12] ) & (~\new_[30709]_  | ~\s3_data_i[12] );
  assign \new_[23134]_  = ~\new_[25182]_ ;
  assign \new_[23135]_  = ~\new_[24662]_ ;
  assign \new_[23136]_  = ~\new_[29300]_  & ~\new_[29355]_ ;
  assign \new_[23137]_  = ~\new_[24661]_ ;
  assign \new_[23138]_  = ~\new_[24667]_ ;
  assign \new_[23139]_  = ~\new_[24677]_ ;
  assign \new_[23140]_  = ~\new_[26273]_ ;
  assign \new_[23141]_  = ~\new_[24668]_ ;
  assign \new_[23142]_  = ~\new_[29064]_  | ~\new_[5987]_ ;
  assign \new_[23143]_  = (~\new_[28768]_  | ~\s5_data_i[20] ) & (~\new_[30457]_  | ~\s3_data_i[20] );
  assign \new_[23144]_  = ~\new_[29997]_  & ~\new_[28001]_ ;
  assign \new_[23145]_  = ~\new_[29508]_  & ~\new_[30265]_ ;
  assign \new_[23146]_  = ~\new_[24674]_ ;
  assign \new_[23147]_  = (~\new_[28392]_  | ~\s4_data_i[0] ) & (~\new_[29349]_  | ~\s0_data_i[0] );
  assign \new_[23148]_  = ~\new_[28217]_  & ~\new_[27710]_ ;
  assign \new_[23149]_  = ~\new_[30409]_  | ~\new_[28786]_  | ~\new_[28138]_ ;
  assign \new_[23150]_  = (~\new_[28313]_  | ~\s7_data_i[16] ) & (~\new_[29707]_  | ~\s6_data_i[16] );
  assign n8084 = ~\new_[29554]_  | ~\new_[27026]_ ;
  assign \new_[23152]_  = ~\new_[29623]_  | ~\new_[29809]_ ;
  assign \new_[23153]_  = (~\new_[28223]_  | ~\s7_data_i[1] ) & (~\new_[28767]_  | ~\s6_data_i[1] );
  assign \new_[23154]_  = ~\new_[29381]_  & ~\new_[30327]_ ;
  assign \new_[23155]_  = ~\new_[26263]_ ;
  assign \new_[23156]_  = (~\new_[28223]_  | ~\s7_data_i[2] ) & (~\new_[28767]_  | ~\s6_data_i[2] );
  assign \new_[23157]_  = ~\new_[29229]_  | ~\new_[6075]_ ;
  assign \new_[23158]_  = ~\new_[30208]_  | ~\new_[31763]_ ;
  assign n8269 = ~\new_[29178]_  | ~\new_[26716]_ ;
  assign \new_[23160]_  = ~\new_[24709]_ ;
  assign n8169 = ~\new_[29484]_  | ~\new_[27023]_ ;
  assign \new_[23162]_  = ~\new_[26256]_ ;
  assign \new_[23163]_  = ~\new_[29290]_  & ~\new_[30034]_ ;
  assign \new_[23164]_  = ~\new_[24620]_ ;
  assign \new_[23165]_  = ~\new_[24710]_ ;
  assign \new_[23166]_  = ~\new_[26257]_ ;
  assign \new_[23167]_  = ~\new_[27570]_  & (~\new_[30242]_  | ~\new_[6053]_ );
  assign \new_[23168]_  = ~\new_[26254]_ ;
  assign \new_[23169]_  = ~\new_[30275]_  & (~\new_[28529]_  | ~\new_[29601]_ );
  assign \new_[23170]_  = ~\new_[27375]_  & ~\new_[29119]_ ;
  assign \new_[23171]_  = ~\new_[30115]_  | ~\new_[6079]_ ;
  assign \new_[23172]_  = ~\new_[30319]_  | ~\new_[5902]_ ;
  assign \new_[23173]_  = ~\new_[29831]_  | ~\new_[29233]_ ;
  assign \new_[23174]_  = ~\new_[26248]_ ;
  assign \new_[23175]_  = (~\new_[28136]_  | ~\s5_data_i[3] ) & (~\new_[29928]_  | ~\s3_data_i[3] );
  assign \new_[23176]_  = \new_[26647]_  & \new_[31690]_ ;
  assign \new_[23177]_  = (~\new_[28223]_  | ~\s7_data_i[29] ) & (~\new_[28767]_  | ~\s6_data_i[29] );
  assign \new_[23178]_  = ~\new_[30526]_  | ~\new_[6061]_ ;
  assign \new_[23179]_  = (~\new_[28392]_  | ~\s4_data_i[16] ) & (~\new_[29349]_  | ~\s0_data_i[16] );
  assign \new_[23180]_  = ~\new_[30423]_  | ~\new_[6194]_ ;
  assign \new_[23181]_  = ~\new_[29792]_  & ~\new_[28762]_ ;
  assign \new_[23182]_  = ~\new_[30243]_  | ~\new_[30595]_ ;
  assign \new_[23183]_  = ~\new_[30467]_  | ~\new_[30432]_ ;
  assign \new_[23184]_  = ~\new_[30185]_  & ~\new_[29598]_ ;
  assign \new_[23185]_  = ~\new_[30149]_  & ~\new_[27778]_ ;
  assign \new_[23186]_  = ~\new_[26227]_ ;
  assign \new_[23187]_  = ~\new_[25770]_ ;
  assign \new_[23188]_  = \new_[27476]_  & \new_[27406]_ ;
  assign \new_[23189]_  = ~\new_[27001]_  & ~\new_[30425]_ ;
  assign \new_[23190]_  = ~\new_[27003]_  & ~\new_[30289]_ ;
  assign \new_[23191]_  = \new_[27046]_  & \new_[27459]_ ;
  assign \new_[23192]_  = ~\new_[26955]_  & ~\new_[30038]_ ;
  assign \new_[23193]_  = \new_[26694]_  & \new_[27051]_ ;
  assign \new_[23194]_  = \new_[26868]_  | \new_[30145]_ ;
  assign \new_[23195]_  = \new_[26873]_  | \new_[26878]_ ;
  assign \new_[23196]_  = \new_[27408]_  & \new_[27820]_ ;
  assign \new_[23197]_  = \new_[27396]_  & \new_[27803]_ ;
  assign \new_[23198]_  = \new_[26884]_  | \new_[26887]_ ;
  assign \new_[23199]_  = \new_[27367]_  & \new_[27086]_ ;
  assign \new_[23200]_  = \new_[26882]_  | \new_[30375]_ ;
  assign \new_[23201]_  = \new_[27326]_  & \new_[27320]_ ;
  assign \new_[23202]_  = \new_[26932]_  | \new_[30038]_ ;
  assign \new_[23203]_  = ~\new_[26611]_  | ~\new_[30508]_ ;
  assign \new_[23204]_  = ~\new_[29959]_  | ~\new_[6208]_ ;
  assign \new_[23205]_  = \new_[27288]_  & \new_[27099]_ ;
  assign \new_[23206]_  = ~\new_[26893]_  & ~\new_[30629]_ ;
  assign \new_[23207]_  = \new_[26967]_  | \new_[30033]_ ;
  assign \new_[23208]_  = ~\new_[26513]_ ;
  assign \new_[23209]_  = ~\new_[27882]_  | ~\new_[30750]_ ;
  assign \new_[23210]_  = ~\new_[26960]_  & ~\new_[30642]_ ;
  assign \new_[23211]_  = \new_[26985]_  | \new_[27863]_ ;
  assign \new_[23212]_  = \new_[26914]_  | \new_[29889]_ ;
  assign \new_[23213]_  = ~\new_[26884]_  | ~\new_[26887]_ ;
  assign \new_[23214]_  = ~\new_[26932]_  & ~\new_[26955]_ ;
  assign \new_[23215]_  = ~\new_[26895]_  | ~\new_[26609]_ ;
  assign \new_[23216]_  = \new_[27180]_  & \new_[26818]_ ;
  assign \new_[23217]_  = ~\new_[27488]_  | ~\new_[30765]_ ;
  assign \new_[23218]_  = ~\new_[26985]_  | ~\new_[27863]_ ;
  assign \new_[23219]_  = \new_[26975]_  | \new_[30151]_ ;
  assign \new_[23220]_  = ~\new_[30069]_  | ~\new_[5903]_ ;
  assign \new_[23221]_  = \new_[26937]_  | \new_[26930]_ ;
  assign \new_[23222]_  = \new_[27527]_  | \new_[30029]_ ;
  assign \new_[23223]_  = \new_[27599]_  | \new_[30254]_ ;
  assign \new_[23224]_  = ~\new_[27072]_  | ~\new_[30574]_ ;
  assign \new_[23225]_  = \new_[26937]_  | \new_[30703]_ ;
  assign \new_[23226]_  = ~\new_[26942]_  | ~\new_[27510]_ ;
  assign \new_[23227]_  = ~\new_[27529]_  & ~\new_[28422]_ ;
  assign \new_[23228]_  = ~\new_[30042]_  | ~\new_[5894]_ ;
  assign \new_[23229]_  = \new_[26923]_  | \new_[29959]_ ;
  assign \new_[23230]_  = ~\new_[26984]_  | ~\new_[27696]_ ;
  assign \new_[23231]_  = \new_[29798]_  | \new_[31776]_ ;
  assign \new_[23232]_  = \new_[27309]_  & \new_[27094]_ ;
  assign \new_[23233]_  = ~\new_[30272]_  | ~\new_[5906]_ ;
  assign \new_[23234]_  = ~\new_[26975]_  & ~\new_[26976]_ ;
  assign \new_[23235]_  = ~\new_[26889]_  | ~\new_[28259]_ ;
  assign \new_[23236]_  = ~\new_[26981]_  | ~\new_[26760]_ ;
  assign \new_[23237]_  = ~\new_[26958]_  | ~\new_[30538]_ ;
  assign \new_[23238]_  = ~\new_[26906]_  | ~\new_[30721]_ ;
  assign \new_[23239]_  = ~\new_[26428]_ ;
  assign \new_[23240]_  = \new_[27668]_  & \new_[27348]_ ;
  assign \new_[23241]_  = \new_[26902]_  | \new_[29930]_ ;
  assign \new_[23242]_  = \new_[27460]_  & \new_[27461]_ ;
  assign \new_[23243]_  = \new_[27827]_  | \new_[30201]_ ;
  assign \new_[23244]_  = ~\new_[26934]_  & ~\new_[30201]_ ;
  assign \new_[23245]_  = ~\new_[30680]_  | ~\new_[24759]_ ;
  assign \new_[23246]_  = ~\new_[26969]_  & ~\new_[30033]_ ;
  assign \new_[23247]_  = ~\new_[26967]_  & ~\new_[26969]_ ;
  assign \new_[23248]_  = ~\new_[26971]_  | ~\new_[28395]_ ;
  assign \new_[23249]_  = ~\new_[26681]_  | ~\new_[27431]_ ;
  assign \new_[23250]_  = ~\new_[26876]_  | ~\new_[28395]_ ;
  assign \new_[23251]_  = \new_[26915]_  | \new_[26899]_ ;
  assign \new_[23252]_  = ~\new_[26921]_  | ~\new_[26922]_ ;
  assign \new_[23253]_  = ~\new_[26998]_  & ~\new_[30677]_ ;
  assign \new_[23254]_  = ~\new_[29174]_  & ~\new_[30087]_ ;
  assign \new_[23255]_  = ~\new_[26982]_  | ~\new_[30610]_ ;
  assign \new_[23256]_  = ~\new_[26983]_  & ~\new_[26910]_ ;
  assign \new_[23257]_  = (~\new_[28223]_  | ~\s7_data_i[8] ) & (~\new_[28767]_  | ~\s6_data_i[8] );
  assign \new_[23258]_  = ~\new_[29061]_  | ~\new_[28732]_ ;
  assign \new_[23259]_  = \new_[27127]_  & \new_[27123]_ ;
  assign \new_[23260]_  = \new_[27719]_  & \new_[27470]_ ;
  assign \new_[23261]_  = ~\new_[30038]_  | ~\new_[31422]_ ;
  assign \new_[23262]_  = ~\new_[26972]_  | ~\new_[27726]_ ;
  assign \new_[23263]_  = \new_[26916]_  & \new_[27763]_ ;
  assign \new_[23264]_  = \new_[26836]_  & \new_[27485]_ ;
  assign \new_[23265]_  = \new_[26736]_  | \new_[26867]_ ;
  assign \new_[23266]_  = ~\new_[30104]_  | ~\new_[28152]_  | ~\new_[28318]_ ;
  assign \new_[23267]_  = ~\new_[24555]_ ;
  assign \new_[23268]_  = ~\new_[24771]_ ;
  assign \new_[23269]_  = ~\new_[27775]_  | ~\new_[28144]_ ;
  assign \new_[23270]_  = ~\new_[30033]_  & (~\new_[28547]_  | ~\new_[29489]_ );
  assign \new_[23271]_  = ~\new_[29889]_  & (~\new_[28459]_  | ~\new_[29344]_ );
  assign \new_[23272]_  = ~\new_[27774]_  | ~\new_[28370]_ ;
  assign \new_[23273]_  = ~\new_[30693]_  | ~\new_[30107]_ ;
  assign \new_[23274]_  = \new_[26936]_  | \new_[28978]_ ;
  assign \new_[23275]_  = (~\new_[28768]_  | ~\s5_data_i[9] ) & (~\new_[30457]_  | ~\s3_data_i[9] );
  assign \new_[23276]_  = ~\new_[29810]_  & (~\new_[28458]_  | ~\new_[29294]_ );
  assign \new_[23277]_  = ~\new_[30192]_  | ~\new_[5897]_ ;
  assign \new_[23278]_  = ~\new_[30105]_  | ~\new_[28663]_  | ~\new_[28464]_ ;
  assign \new_[23279]_  = ~\new_[30151]_  & (~\new_[28174]_  | ~\new_[29390]_ );
  assign \new_[23280]_  = ~\new_[30201]_  & (~\new_[28436]_  | ~\new_[29577]_ );
  assign \new_[23281]_  = ~\new_[30326]_  & (~\new_[28457]_  | ~\new_[29461]_ );
  assign n8094 = ~\new_[29617]_  | ~\new_[27005]_ ;
  assign n8124 = ~\new_[29634]_  | ~\new_[27034]_ ;
  assign n8144 = ~\new_[28914]_  | ~\new_[27029]_ ;
  assign n8149 = ~\new_[28943]_  | ~\new_[27025]_ ;
  assign n8154 = ~\new_[28886]_  | ~\new_[27027]_ ;
  assign n8194 = ~\new_[29667]_  | ~\new_[27022]_ ;
  assign n8189 = ~\new_[28839]_  | ~\new_[27021]_ ;
  assign n8184 = ~\new_[29261]_  | ~\new_[27006]_ ;
  assign n8199 = ~\new_[29094]_  | ~\new_[27020]_ ;
  assign n8059 = ~\new_[29327]_  | ~\new_[27009]_ ;
  assign n8254 = ~\new_[29609]_  | ~\new_[27040]_ ;
  assign n8249 = ~\new_[29668]_  | ~\new_[27010]_ ;
  assign n8239 = ~\new_[29605]_  | ~\new_[26624]_ ;
  assign n8244 = ~\new_[28965]_  | ~\new_[27011]_ ;
  assign n8064 = ~\new_[29594]_  | ~\new_[27039]_ ;
  assign n8234 = ~\new_[29133]_  | ~\new_[26690]_ ;
  assign n8179 = ~\new_[29395]_  | ~\new_[27012]_ ;
  assign n8069 = ~\new_[29065]_  | ~\new_[27014]_ ;
  assign n8209 = ~\new_[29252]_  | ~\new_[27016]_ ;
  assign n8074 = ~\new_[28955]_  | ~\new_[27017]_ ;
  assign \new_[23302]_  = ~\new_[28766]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign n8264 = ~\new_[29693]_  | ~\new_[27019]_ ;
  assign n8204 = ~\new_[29107]_  | ~\new_[27018]_ ;
  assign n8079 = ~\new_[29614]_  | ~\new_[26697]_ ;
  assign \new_[23306]_  = ~\new_[30277]_  | ~\new_[5926]_ ;
  assign n8174 = ~\new_[28945]_  | ~\new_[26692]_ ;
  assign n8164 = ~\new_[29727]_  | ~\new_[27024]_ ;
  assign n8159 = ~\new_[29691]_  | ~\new_[26684]_ ;
  assign n8134 = ~\new_[29657]_  | ~\new_[27030]_ ;
  assign n8139 = ~\new_[29203]_  | ~\new_[27031]_ ;
  assign n8129 = ~\new_[28852]_  | ~\new_[26718]_ ;
  assign n8089 = ~\new_[29596]_  | ~\new_[27032]_ ;
  assign n8119 = ~\new_[29432]_  | ~\new_[27035]_ ;
  assign n8114 = ~\new_[29234]_  | ~\new_[27036]_ ;
  assign n8099 = ~\new_[29269]_  | ~\new_[26992]_ ;
  assign n8109 = ~\new_[29316]_  | ~\new_[27037]_ ;
  assign n8104 = ~\new_[28947]_  | ~\new_[26666]_ ;
  assign n8214 = ~\new_[29083]_  | ~\new_[27013]_ ;
  assign n8219 = ~\new_[29574]_  | ~\new_[26663]_ ;
  assign \new_[23321]_  = ~\new_[30145]_  & (~\new_[28469]_  | ~\new_[29500]_ );
  assign n8224 = ~\new_[29097]_  | ~\new_[27038]_ ;
  assign n8229 = ~\new_[29116]_  | ~\new_[26648]_ ;
  assign n8259 = ~\new_[28826]_  | ~\new_[27008]_ ;
  assign n8274 = ~\new_[29190]_  | ~\new_[27007]_ ;
  assign \new_[23326]_  = ~\new_[28503]_  & (~\new_[29431]_  | ~\new_[28045]_ );
  assign \new_[23327]_  = ~\new_[27643]_  & (~\new_[29380]_  | ~\new_[30367]_ );
  assign \new_[23328]_  = ~\new_[30467]_  | (~\new_[29482]_  & ~\new_[28745]_ );
  assign \new_[23329]_  = ~\new_[27616]_  & (~\new_[29176]_  | ~\new_[30290]_ );
  assign \new_[23330]_  = ~\new_[29994]_  | ~\new_[5901]_ ;
  assign \new_[23331]_  = ~\new_[26581]_  & ~\new_[28867]_ ;
  assign \new_[23332]_  = ~\new_[24795]_ ;
  assign \new_[23333]_  = ~\new_[27487]_  & ~\new_[29861]_ ;
  assign \new_[23334]_  = ~\new_[27544]_  | ~\new_[30150]_ ;
  assign \new_[23335]_  = ~\new_[26952]_  & ~\new_[30540]_ ;
  assign \new_[23336]_  = ~\new_[24798]_ ;
  assign \new_[23337]_  = \new_[26755]_  | \new_[29573]_ ;
  assign \new_[23338]_  = ~\new_[27329]_  & ~\new_[29578]_ ;
  assign \new_[23339]_  = ~\new_[26794]_  | ~\new_[30283]_ ;
  assign \new_[23340]_  = ~\new_[24803]_ ;
  assign \new_[23341]_  = \new_[28569]_  | \new_[29383]_ ;
  assign \new_[23342]_  = ~\new_[27437]_  | ~\new_[30221]_ ;
  assign \new_[23343]_  = ~\new_[27679]_  | ~\new_[30316]_ ;
  assign \new_[23344]_  = \new_[27761]_  | \new_[29784]_ ;
  assign \new_[23345]_  = ~\new_[24807]_ ;
  assign \new_[23346]_  = \new_[26745]_  & \new_[30544]_ ;
  assign \new_[23347]_  = ~\new_[28904]_  & ~\new_[26814]_ ;
  assign \new_[23348]_  = ~\new_[26686]_  | ~\new_[30617]_ ;
  assign \new_[23349]_  = ~\new_[24593]_ ;
  assign \new_[23350]_  = \new_[27750]_  | \new_[29784]_ ;
  assign \new_[23351]_  = \new_[26704]_  | \new_[29333]_ ;
  assign \new_[23352]_  = \new_[28522]_  | \new_[30044]_ ;
  assign \new_[23353]_  = ~\new_[27083]_  & ~\new_[30140]_ ;
  assign \new_[23354]_  = ~\new_[27431]_  & ~\new_[30845]_ ;
  assign \new_[23355]_  = ~\new_[24813]_ ;
  assign \new_[23356]_  = ~\new_[24814]_ ;
  assign \new_[23357]_  = ~\new_[5913]_  | ~\new_[28969]_  | ~\new_[28880]_ ;
  assign \new_[23358]_  = \new_[27904]_  & \new_[28069]_ ;
  assign \new_[23359]_  = ~\new_[26784]_  & ~\new_[30713]_ ;
  assign \new_[23360]_  = \new_[26822]_  | \new_[29839]_ ;
  assign \new_[23361]_  = ~\new_[26729]_  | ~\new_[29212]_ ;
  assign \new_[23362]_  = ~\new_[27371]_  & ~\new_[29195]_ ;
  assign \new_[23363]_  = ~\new_[28513]_  | ~\new_[27802]_ ;
  assign \new_[23364]_  = ~\new_[29475]_  | ~\new_[27845]_ ;
  assign \new_[23365]_  = ~\new_[24821]_ ;
  assign \new_[23366]_  = ~\new_[27898]_  | ~\new_[29527]_ ;
  assign \new_[23367]_  = \new_[27944]_  | \new_[29841]_ ;
  assign \new_[23368]_  = ~\new_[28414]_  | ~\new_[27577]_ ;
  assign \new_[23369]_  = (~\new_[28223]_  | ~\s7_data_i[10] ) & (~\new_[28767]_  | ~\s6_data_i[10] );
  assign \new_[23370]_  = ~\new_[27507]_  & ~\new_[30694]_ ;
  assign \new_[23371]_  = \new_[26847]_  | \new_[29648]_ ;
  assign \new_[23372]_  = ~\new_[27526]_  & ~\new_[30069]_ ;
  assign \new_[23373]_  = ~\new_[26775]_  | ~\new_[29079]_ ;
  assign \new_[23374]_  = \new_[27808]_  | \new_[29966]_ ;
  assign \new_[23375]_  = ~\new_[24832]_ ;
  assign \new_[23376]_  = \new_[27177]_  & \new_[29003]_ ;
  assign \new_[23377]_  = ~\new_[24833]_ ;
  assign \new_[23378]_  = \new_[27824]_  | \new_[29966]_ ;
  assign \new_[23379]_  = ~\new_[27542]_  & ~\new_[28027]_ ;
  assign \new_[23380]_  = ~\new_[27818]_  | ~\new_[30135]_ ;
  assign \new_[23381]_  = ~\new_[24544]_ ;
  assign \new_[23382]_  = \new_[29206]_  | \new_[29544]_ ;
  assign \new_[23383]_  = \new_[27678]_  | \new_[30425]_ ;
  assign \new_[23384]_  = \new_[27634]_  & \new_[30142]_ ;
  assign \new_[23385]_  = \new_[29447]_  & \new_[29159]_ ;
  assign \new_[23386]_  = ~\new_[27325]_  | ~\new_[29212]_ ;
  assign \new_[23387]_  = ~\new_[24838]_ ;
  assign \new_[23388]_  = \new_[27686]_  | \new_[30425]_ ;
  assign \new_[23389]_  = \new_[27503]_  | \new_[29181]_ ;
  assign \new_[23390]_  = \new_[26874]_  | \new_[29582]_ ;
  assign \new_[23391]_  = ~\new_[26653]_  | ~\new_[29813]_ ;
  assign \new_[23392]_  = \new_[27758]_  | \new_[30040]_ ;
  assign \new_[23393]_  = \new_[27758]_  & \new_[27942]_ ;
  assign \new_[23394]_  = ~\new_[28184]_  & ~\new_[30334]_ ;
  assign \new_[23395]_  = \new_[27561]_  & \new_[27802]_ ;
  assign \new_[23396]_  = ~\new_[28541]_  & ~\new_[30334]_ ;
  assign \new_[23397]_  = (~\new_[28392]_  | ~\s4_data_i[10] ) & (~\new_[29349]_  | ~\s0_data_i[10] );
  assign \new_[23398]_  = ~\new_[27231]_  | ~\new_[29320]_ ;
  assign \new_[23399]_  = ~\new_[26740]_  & ~\new_[30629]_ ;
  assign \new_[23400]_  = ~\new_[27298]_  & ~\new_[29815]_ ;
  assign \new_[23401]_  = ~\new_[26604]_  | ~\new_[29171]_ ;
  assign \new_[23402]_  = ~\new_[27298]_  & ~\new_[30575]_ ;
  assign \new_[23403]_  = ~\new_[28865]_  & ~\new_[29965]_ ;
  assign \new_[23404]_  = ~\new_[27674]_  & ~\new_[30109]_ ;
  assign \new_[23405]_  = ~\new_[24846]_ ;
  assign \new_[23406]_  = \new_[26779]_  | \new_[30400]_ ;
  assign \new_[23407]_  = \new_[29294]_  & \new_[29746]_ ;
  assign \new_[23408]_  = ~\new_[27516]_  & ~\new_[29930]_ ;
  assign \new_[23409]_  = ~\new_[24851]_ ;
  assign \new_[23410]_  = ~\new_[27530]_  | ~\new_[28866]_ ;
  assign \new_[23411]_  = ~\new_[5968]_  | ~\new_[30386]_  | ~\new_[29260]_ ;
  assign \new_[23412]_  = \new_[26901]_  | \new_[29736]_ ;
  assign \new_[23413]_  = ~\new_[24852]_ ;
  assign \new_[23414]_  = ~\new_[27773]_  | ~\new_[28989]_ ;
  assign \new_[23415]_  = \new_[27836]_  & \new_[29192]_ ;
  assign \new_[23416]_  = ~\new_[27836]_  | ~\new_[29983]_ ;
  assign \new_[23417]_  = ~\new_[29028]_  | ~\new_[30332]_ ;
  assign \new_[23418]_  = \new_[26592]_  | \new_[29736]_ ;
  assign \new_[23419]_  = ~\new_[26834]_  | ~\new_[29682]_ ;
  assign \new_[23420]_  = ~\new_[26609]_  | ~\new_[30604]_ ;
  assign \new_[23421]_  = \new_[29536]_  & \new_[30571]_ ;
  assign \new_[23422]_  = ~\new_[27896]_  | ~\new_[30665]_ ;
  assign \new_[23423]_  = ~\new_[27388]_  | ~\new_[30574]_ ;
  assign \new_[23424]_  = ~\new_[26597]_  | ~\new_[30550]_ ;
  assign \new_[23425]_  = ~\new_[29183]_  | ~\new_[27787]_ ;
  assign \new_[23426]_  = \new_[27736]_  & \new_[27787]_ ;
  assign \new_[23427]_  = ~\new_[29471]_  | ~\new_[27736]_ ;
  assign \new_[23428]_  = ~\new_[27511]_  & ~\new_[26857]_ ;
  assign \new_[23429]_  = \new_[26735]_  & \new_[26845]_ ;
  assign \new_[23430]_  = ~\new_[27541]_  | ~\new_[30022]_ ;
  assign \new_[23431]_  = \new_[27613]_  & \new_[27191]_ ;
  assign \new_[23432]_  = ~\new_[27499]_  & ~\new_[28833]_ ;
  assign \new_[23433]_  = ~\new_[27499]_  & ~\new_[30202]_ ;
  assign \new_[23434]_  = ~\new_[26803]_  | ~\new_[29228]_ ;
  assign \new_[23435]_  = \new_[27394]_  | \new_[30202]_ ;
  assign \new_[23436]_  = ~\new_[27887]_  & ~\new_[30785]_ ;
  assign \new_[23437]_  = ~\new_[26562]_ ;
  assign \new_[23438]_  = ~\new_[27516]_  & ~\new_[30769]_ ;
  assign \new_[23439]_  = ~\new_[26414]_ ;
  assign \new_[23440]_  = ~\new_[26953]_  & ~\new_[30319]_ ;
  assign \new_[23441]_  = ~\new_[24870]_ ;
  assign \new_[23442]_  = \new_[29351]_  & \new_[30686]_ ;
  assign \new_[23443]_  = \new_[27541]_  & \new_[30497]_ ;
  assign \new_[23444]_  = \new_[26710]_  | \new_[29767]_ ;
  assign \new_[23445]_  = ~\new_[26862]_  | ~\new_[28969]_ ;
  assign \new_[23446]_  = ~\new_[27532]_  & ~\new_[28678]_ ;
  assign \new_[23447]_  = ~\new_[26951]_  | ~\new_[29692]_ ;
  assign \new_[23448]_  = ~\new_[26815]_  | ~\new_[28837]_ ;
  assign \new_[23449]_  = ~\new_[27083]_  & ~\new_[29056]_ ;
  assign \new_[23450]_  = \new_[29601]_  & \new_[29299]_ ;
  assign \new_[23451]_  = \new_[29577]_  & \new_[30603]_ ;
  assign \new_[23452]_  = \new_[26614]_  | \new_[29827]_ ;
  assign \new_[23453]_  = ~\new_[24874]_ ;
  assign \new_[23454]_  = ~\new_[27442]_  | ~\new_[30294]_ ;
  assign \new_[23455]_  = \new_[27542]_  | \new_[29293]_ ;
  assign \new_[23456]_  = ~\new_[29569]_  & ~\new_[29672]_ ;
  assign \new_[23457]_  = ~\new_[27489]_  & ~\new_[30008]_ ;
  assign \new_[23458]_  = ~\new_[24880]_ ;
  assign \new_[23459]_  = \new_[27608]_  | \new_[30203]_ ;
  assign \new_[23460]_  = ~\new_[27602]_  & ~\new_[30192]_ ;
  assign \new_[23461]_  = ~\new_[30116]_  & ~\new_[26717]_ ;
  assign \new_[23462]_  = \new_[28482]_  | \new_[28899]_ ;
  assign \new_[23463]_  = ~\new_[28482]_  & ~\new_[30249]_ ;
  assign \new_[23464]_  = ~\new_[28510]_  & ~\new_[30249]_ ;
  assign \new_[23465]_  = ~\new_[26715]_  & ~\new_[30249]_ ;
  assign \new_[23466]_  = \new_[27498]_  | \new_[29931]_ ;
  assign \new_[23467]_  = ~\new_[28225]_  & ~\new_[30192]_ ;
  assign \new_[23468]_  = ~\new_[27744]_  | ~\new_[29139]_ ;
  assign \new_[23469]_  = ~\new_[26974]_  & ~\new_[30616]_ ;
  assign \new_[23470]_  = ~\new_[27310]_  & ~\new_[28998]_ ;
  assign \new_[23471]_  = ~\new_[24895]_ ;
  assign \new_[23472]_  = ~\new_[26517]_ ;
  assign \new_[23473]_  = ~\new_[5830]_  | ~\new_[29150]_  | ~\new_[29977]_ ;
  assign \new_[23474]_  = ~\new_[27536]_  & ~\new_[29013]_ ;
  assign \new_[23475]_  = ~\new_[28431]_  & ~\new_[29166]_ ;
  assign \new_[23476]_  = ~\new_[24898]_ ;
  assign \new_[23477]_  = \new_[26822]_  & \new_[27384]_ ;
  assign \new_[23478]_  = ~\new_[24899]_ ;
  assign \new_[23479]_  = \new_[27950]_  & \new_[28054]_ ;
  assign \new_[23480]_  = \new_[27556]_  | \new_[30389]_ ;
  assign \new_[23481]_  = ~\new_[26506]_ ;
  assign \new_[23482]_  = ~\new_[26743]_  | ~\new_[29922]_ ;
  assign \new_[23483]_  = \new_[28475]_  | \new_[29166]_ ;
  assign \new_[23484]_  = ~\new_[26502]_ ;
  assign \new_[23485]_  = ~\new_[24902]_ ;
  assign \new_[23486]_  = \new_[29474]_  & \new_[30846]_ ;
  assign \new_[23487]_  = \new_[29311]_  | \new_[29544]_ ;
  assign \new_[23488]_  = ~\new_[24907]_ ;
  assign \new_[23489]_  = \new_[29480]_  & \new_[30667]_ ;
  assign \new_[23490]_  = ~\new_[27723]_  | ~\new_[28732]_ ;
  assign \new_[23491]_  = ~\new_[27718]_  & ~\new_[30044]_ ;
  assign \new_[23492]_  = ~\new_[27403]_  & ~\new_[29062]_ ;
  assign \new_[23493]_  = \new_[27403]_  | \new_[29902]_ ;
  assign \new_[23494]_  = ~\new_[27687]_  | ~\new_[28121]_ ;
  assign \new_[23495]_  = ~\new_[28083]_  & ~\new_[27722]_ ;
  assign \new_[23496]_  = \new_[26607]_  | \new_[30443]_ ;
  assign \new_[23497]_  = ~\new_[24914]_ ;
  assign \new_[23498]_  = ~\new_[26616]_  & ~\new_[29959]_ ;
  assign \new_[23499]_  = \new_[27644]_  | \new_[30080]_ ;
  assign \new_[23500]_  = ~\new_[6031]_  | ~\new_[29922]_  | ~\new_[29782]_ ;
  assign \new_[23501]_  = \new_[27651]_  | \new_[29736]_ ;
  assign \new_[23502]_  = \new_[27687]_  & \new_[28877]_ ;
  assign \new_[23503]_  = ~\new_[27130]_  & ~\new_[29652]_ ;
  assign \new_[23504]_  = ~\new_[26950]_  & ~\new_[30637]_ ;
  assign \new_[23505]_  = ~\new_[29729]_  | ~\new_[27593]_ ;
  assign \new_[23506]_  = (~\new_[28392]_  | ~\s4_data_i[11] ) & (~\new_[29349]_  | ~\s0_data_i[11] );
  assign \new_[23507]_  = \new_[27642]_  | \new_[28402]_ ;
  assign \new_[23508]_  = ~\new_[26750]_  & ~\new_[29776]_ ;
  assign \new_[23509]_  = ~\new_[26834]_  | ~\new_[29233]_ ;
  assign \new_[23510]_  = ~\new_[26846]_  | ~\new_[30217]_ ;
  assign \new_[23511]_  = \new_[27648]_  | \new_[30240]_ ;
  assign \new_[23512]_  = ~\new_[29564]_  & ~\new_[29350]_ ;
  assign \new_[23513]_  = \new_[27656]_  | \new_[29222]_ ;
  assign \new_[23514]_  = \new_[28501]_  | \new_[29096]_ ;
  assign \new_[23515]_  = \new_[27646]_  | \new_[29222]_ ;
  assign \new_[23516]_  = ~\new_[24925]_ ;
  assign \new_[23517]_  = ~\new_[29792]_  & ~\new_[29324]_ ;
  assign \new_[23518]_  = ~\new_[26444]_ ;
  assign \new_[23519]_  = (~\new_[28392]_  | ~\s4_data_i[25] ) & (~\new_[29349]_  | ~\s0_data_i[25] );
  assign \new_[23520]_  = ~\new_[27504]_  & ~\new_[30443]_ ;
  assign \new_[23521]_  = ~\new_[27618]_  | ~\new_[30721]_ ;
  assign \new_[23522]_  = \new_[27950]_  | \new_[29089]_ ;
  assign \new_[23523]_  = \new_[27744]_  & \new_[29162]_ ;
  assign \new_[23524]_  = \new_[26675]_  | \new_[28899]_ ;
  assign \new_[23525]_  = (~\new_[28768]_  | ~\s5_data_i[12] ) & (~\new_[30457]_  | ~\s3_data_i[12] );
  assign \new_[23526]_  = ~\new_[27748]_  & ~\new_[28982]_ ;
  assign \new_[23527]_  = \new_[27707]_  & \new_[29441]_ ;
  assign \new_[23528]_  = ~\new_[24930]_ ;
  assign \new_[23529]_  = ~\new_[26413]_ ;
  assign \new_[23530]_  = ~\new_[27517]_  & ~\new_[28361]_ ;
  assign \new_[23531]_  = ~\new_[26702]_  & ~\new_[28909]_ ;
  assign \new_[23532]_  = ~\new_[26585]_  & ~\new_[30199]_ ;
  assign \new_[23533]_  = ~\new_[26991]_  & ~\new_[30688]_ ;
  assign \new_[23534]_  = ~\new_[26850]_  & ~\new_[29132]_ ;
  assign \new_[23535]_  = ~\new_[26991]_  | ~\new_[26708]_ ;
  assign \new_[23536]_  = ~\new_[27514]_  & ~\new_[30188]_ ;
  assign \new_[23537]_  = ~\new_[26384]_ ;
  assign \new_[23538]_  = ~\new_[26153]_ ;
  assign \new_[23539]_  = ~\new_[26980]_  & ~\new_[30301]_ ;
  assign \new_[23540]_  = ~\new_[26613]_  & ~\new_[30266]_ ;
  assign \new_[23541]_  = ~\new_[26885]_  | ~\new_[30344]_ ;
  assign \new_[23542]_  = ~\new_[26753]_  & ~\new_[29371]_ ;
  assign \new_[23543]_  = ~\new_[27610]_  | ~\new_[30246]_ ;
  assign \new_[23544]_  = ~\new_[24941]_ ;
  assign \new_[23545]_  = ~\new_[24942]_ ;
  assign \new_[23546]_  = \new_[26659]_  & \new_[29271]_ ;
  assign \new_[23547]_  = ~\new_[30136]_  | ~\new_[26638]_ ;
  assign \new_[23548]_  = ~\new_[24944]_ ;
  assign \new_[23549]_  = \new_[26685]_  | \new_[30407]_ ;
  assign \new_[23550]_  = ~\new_[6059]_  | ~\new_[30294]_  | ~\new_[29967]_ ;
  assign \new_[23551]_  = ~\new_[27311]_  & ~\new_[28797]_ ;
  assign \new_[23552]_  = ~\new_[26703]_  & ~\new_[28829]_ ;
  assign \new_[23553]_  = ~\new_[26602]_  | ~\new_[30117]_ ;
  assign \new_[23554]_  = \new_[29665]_  | \new_[29375]_ ;
  assign \new_[23555]_  = ~\new_[24948]_ ;
  assign \new_[23556]_  = ~\new_[24949]_ ;
  assign \new_[23557]_  = \new_[27579]_  & \new_[30627]_ ;
  assign \new_[23558]_  = ~\new_[5981]_  | ~\new_[29162]_  | ~\new_[30279]_ ;
  assign \new_[23559]_  = \new_[28942]_  | \new_[29375]_ ;
  assign \new_[23560]_  = \new_[28559]_  | \new_[29331]_ ;
  assign \new_[23561]_  = ~\new_[6071]_  | ~\new_[29892]_  | ~\new_[30600]_ ;
  assign \new_[23562]_  = \new_[26741]_  | \new_[29639]_ ;
  assign \new_[23563]_  = \new_[26741]_  & \new_[28641]_ ;
  assign \new_[23564]_  = ~\new_[24950]_ ;
  assign \new_[23565]_  = \new_[26724]_  & \new_[29817]_ ;
  assign \new_[23566]_  = ~\new_[26623]_  & ~\new_[29331]_ ;
  assign \new_[23567]_  = \new_[27801]_  & \new_[28828]_ ;
  assign \new_[23568]_  = \new_[27730]_  | \new_[30701]_ ;
  assign \new_[23569]_  = ~\new_[29151]_  | ~\new_[29789]_ ;
  assign \new_[23570]_  = ~\new_[24953]_ ;
  assign \new_[23571]_  = ~\new_[26809]_  & ~\new_[30302]_ ;
  assign \new_[23572]_  = ~\new_[26943]_  | ~\new_[30210]_ ;
  assign \new_[23573]_  = ~\new_[24955]_ ;
  assign \new_[23574]_  = ~\new_[28384]_  & ~\new_[29934]_ ;
  assign \new_[23575]_  = ~\new_[27704]_  | ~\new_[28050]_ ;
  assign \new_[23576]_  = ~\new_[27901]_  & ~\new_[30254]_ ;
  assign \new_[23577]_  = ~\new_[24956]_ ;
  assign \new_[23578]_  = ~\new_[27756]_  | ~\new_[29186]_ ;
  assign \new_[23579]_  = ~\new_[27558]_  | ~\new_[29162]_ ;
  assign \new_[23580]_  = ~\new_[5981]_  | ~\new_[30279]_  | ~\new_[29139]_ ;
  assign \new_[23581]_  = ~\new_[28554]_  & ~\new_[30319]_ ;
  assign \new_[23582]_  = \new_[26751]_  | \new_[29222]_ ;
  assign \new_[23583]_  = ~\new_[27098]_  & ~\new_[30209]_ ;
  assign \new_[23584]_  = ~\new_[26769]_  & ~\new_[29181]_ ;
  assign \new_[23585]_  = \new_[27756]_  & \new_[29397]_ ;
  assign \new_[23586]_  = ~\new_[27971]_  | ~\new_[30636]_ ;
  assign \new_[23587]_  = \new_[27685]_  & \new_[30329]_ ;
  assign \new_[23588]_  = \new_[27310]_  | \new_[30261]_ ;
  assign \new_[23589]_  = \new_[27620]_  | \new_[30068]_ ;
  assign \new_[23590]_  = ~\new_[28120]_  | ~\new_[29150]_ ;
  assign \new_[23591]_  = \new_[27845]_  & \new_[28039]_ ;
  assign \new_[23592]_  = \new_[29305]_  & \new_[30640]_ ;
  assign \new_[23593]_  = \new_[27621]_  | \new_[29833]_ ;
  assign \new_[23594]_  = ~\new_[30047]_  | ~\new_[6093]_ ;
  assign \new_[23595]_  = \new_[27632]_  & \new_[27285]_ ;
  assign \new_[23596]_  = ~\new_[27500]_  & ~\new_[26788]_ ;
  assign \new_[23597]_  = ~\new_[27986]_  | ~\new_[29064]_ ;
  assign \new_[23598]_  = ~\new_[27638]_  | ~\new_[29977]_ ;
  assign \new_[23599]_  = ~\new_[5985]_  | ~\new_[29506]_  | ~\new_[29887]_ ;
  assign \new_[23600]_  = ~\new_[27490]_  & ~\new_[30632]_ ;
  assign \new_[23601]_  = ~\new_[26941]_  & ~\new_[30746]_ ;
  assign \new_[23602]_  = ~\new_[27490]_  | ~\new_[27672]_ ;
  assign \new_[23603]_  = ~\new_[27671]_  & ~\new_[28021]_ ;
  assign \new_[23604]_  = ~\new_[24970]_ ;
  assign \new_[23605]_  = ~\new_[5968]_  | ~\new_[28866]_  | ~\new_[30386]_ ;
  assign \new_[23606]_  = ~\new_[5985]_  | ~\new_[29086]_  | ~\new_[29506]_ ;
  assign \new_[23607]_  = ~\new_[26578]_  | ~\new_[29086]_ ;
  assign \new_[23608]_  = ~\new_[27609]_  | ~\new_[29006]_ ;
  assign \new_[23609]_  = ~\new_[27753]_  & ~\new_[30168]_ ;
  assign \new_[23610]_  = \new_[27699]_  | \new_[30173]_ ;
  assign \new_[23611]_  = ~\new_[24977]_ ;
  assign \new_[23612]_  = (~\s7_data_i[28]  | ~\new_[27985]_ ) & (~\s6_data_i[28]  | ~\new_[29708]_ );
  assign \new_[23613]_  = \new_[27671]_  | \new_[29069]_ ;
  assign \new_[23614]_  = \new_[29415]_  | \new_[29544]_ ;
  assign \new_[23615]_  = ~\new_[24983]_ ;
  assign \new_[23616]_  = ~\new_[24986]_ ;
  assign \new_[23617]_  = \new_[27613]_  | \new_[30292]_ ;
  assign \new_[23618]_  = ~\new_[28453]_  & ~\new_[30008]_ ;
  assign \new_[23619]_  = ~\new_[28433]_  & ~\new_[30069]_ ;
  assign \new_[23620]_  = ~\new_[28186]_  & ~\new_[30069]_ ;
  assign \new_[23621]_  = ~\new_[29276]_  | ~\new_[29965]_ ;
  assign \new_[23622]_  = \new_[27608]_  & \new_[27826]_ ;
  assign \new_[23623]_  = ~\new_[26804]_  | ~\new_[30765]_ ;
  assign \new_[23624]_  = \new_[28441]_  | \new_[27591]_ ;
  assign \new_[23625]_  = ~\new_[24991]_ ;
  assign \new_[23626]_  = \new_[27951]_  | \new_[28857]_ ;
  assign \new_[23627]_  = \new_[27771]_  | \new_[29830]_ ;
  assign \new_[23628]_  = ~\new_[26767]_  | ~\new_[29974]_ ;
  assign \new_[23629]_  = ~\new_[26843]_  | ~\new_[28073]_ ;
  assign \new_[23630]_  = ~\new_[29248]_  | ~\new_[29663]_ ;
  assign \new_[23631]_  = ~\new_[24997]_ ;
  assign \new_[23632]_  = ~\new_[28449]_  & ~\new_[30319]_ ;
  assign \new_[23633]_  = ~\new_[26022]_ ;
  assign \new_[23634]_  = ~\new_[28578]_  | ~\new_[29590]_ ;
  assign \new_[23635]_  = \new_[27524]_  | \new_[30140]_ ;
  assign \new_[23636]_  = ~\new_[28061]_  | ~\new_[27561]_ ;
  assign \new_[23637]_  = \new_[27725]_  & \new_[29404]_ ;
  assign \new_[23638]_  = ~\new_[27666]_  | ~\new_[27635]_ ;
  assign \new_[23639]_  = ~\new_[25999]_ ;
  assign \new_[23640]_  = ~\new_[28153]_  & ~\new_[29595]_ ;
  assign \new_[23641]_  = \new_[27513]_  | \new_[29174]_ ;
  assign \new_[23642]_  = ~\new_[25001]_ ;
  assign \new_[23643]_  = \new_[28855]_  | \new_[29367]_ ;
  assign \new_[23644]_  = \new_[27495]_  | \new_[30415]_ ;
  assign \new_[23645]_  = ~\new_[28565]_  & ~\new_[30247]_ ;
  assign \new_[23646]_  = ~\new_[27514]_  & ~\new_[30661]_ ;
  assign \new_[23647]_  = \new_[27663]_  & \new_[30321]_ ;
  assign \new_[23648]_  = ~\new_[27640]_  & ~\new_[30093]_ ;
  assign \new_[23649]_  = ~\new_[27510]_  | ~\new_[30243]_ ;
  assign \new_[23650]_  = \new_[29449]_  | \new_[29367]_ ;
  assign \new_[23651]_  = (~\new_[27985]_  | ~\s7_data_i[31] ) & (~\new_[29708]_  | ~\s6_data_i[31] );
  assign \new_[23652]_  = ~\new_[27649]_  | ~\new_[30437]_ ;
  assign \new_[23653]_  = ~\new_[29487]_  & ~\new_[29750]_ ;
  assign \new_[23654]_  = ~\new_[27860]_  | ~\new_[30125]_ ;
  assign \new_[23655]_  = ~\new_[27923]_  | ~\new_[29225]_ ;
  assign \new_[23656]_  = \new_[27807]_  | \new_[30224]_ ;
  assign \new_[23657]_  = ~\new_[27571]_  | ~\new_[29032]_ ;
  assign \new_[23658]_  = ~\new_[27261]_  & ~\new_[30684]_ ;
  assign \new_[23659]_  = \new_[29390]_  & \new_[30635]_ ;
  assign \new_[23660]_  = ~\new_[28079]_  & ~\new_[29394]_ ;
  assign \new_[23661]_  = \new_[27596]_  & \new_[28640]_ ;
  assign \new_[23662]_  = ~\new_[26961]_  | ~\new_[29912]_ ;
  assign \new_[23663]_  = ~\new_[28251]_  | ~\new_[29560]_ ;
  assign \new_[23664]_  = ~\new_[25018]_ ;
  assign \new_[23665]_  = \new_[27632]_  | \new_[30043]_ ;
  assign \new_[23666]_  = ~\new_[27289]_  | ~\new_[28889]_ ;
  assign \new_[23667]_  = ~\new_[28291]_  & ~\new_[30008]_ ;
  assign \new_[23668]_  = ~\new_[25020]_ ;
  assign \new_[23669]_  = ~\new_[25100]_ ;
  assign \new_[23670]_  = ~\new_[25022]_ ;
  assign \new_[23671]_  = \new_[27515]_  & \new_[30505]_ ;
  assign \new_[23672]_  = ~\new_[29182]_  | ~\new_[27769]_ ;
  assign \new_[23673]_  = ~\new_[26950]_  | ~\new_[27682]_ ;
  assign \new_[23674]_  = ~\new_[25027]_ ;
  assign \new_[23675]_  = ~\new_[28335]_  | ~\new_[26940]_ ;
  assign \new_[23676]_  = ~\new_[27612]_  & ~\new_[30662]_ ;
  assign \new_[23677]_  = ~\new_[26733]_  | ~\new_[28878]_ ;
  assign \new_[23678]_  = ~\new_[5994]_  | ~\new_[30158]_  | ~\new_[30316]_ ;
  assign \new_[23679]_  = \new_[27093]_  | \new_[29100]_ ;
  assign \new_[23680]_  = ~\new_[25029]_ ;
  assign \new_[23681]_  = \new_[27769]_  & \new_[30491]_ ;
  assign \new_[23682]_  = ~\new_[25030]_ ;
  assign \new_[23683]_  = \new_[27410]_  | \new_[30173]_ ;
  assign \new_[23684]_  = \new_[29483]_  & \new_[30513]_ ;
  assign \new_[23685]_  = ~\new_[5919]_  | ~\new_[29175]_  | ~\new_[29974]_ ;
  assign \new_[23686]_  = \new_[26657]_  & \new_[5913]_ ;
  assign \new_[23687]_  = ~\new_[28446]_  & ~\new_[29331]_ ;
  assign \new_[23688]_  = ~\new_[28506]_  | ~\new_[27926]_ ;
  assign \new_[23689]_  = ~\new_[27177]_  | ~\new_[29969]_ ;
  assign \new_[23690]_  = \new_[28871]_  & \new_[30641]_ ;
  assign \new_[23691]_  = \new_[26940]_  & \new_[26655]_ ;
  assign \new_[23692]_  = ~\new_[27731]_  & ~\new_[28950]_ ;
  assign \new_[23693]_  = ~\new_[27695]_  & ~\new_[30174]_ ;
  assign \new_[23694]_  = ~\new_[25038]_ ;
  assign \new_[23695]_  = \new_[27723]_  & \new_[28985]_ ;
  assign \new_[23696]_  = ~\new_[29447]_  | ~\new_[29435]_ ;
  assign \new_[23697]_  = ~\new_[26837]_  & ~\new_[30066]_ ;
  assign \new_[23698]_  = ~\new_[27698]_  | ~\new_[29355]_ ;
  assign \new_[23699]_  = ~\new_[28747]_  | ~\new_[26745]_ ;
  assign \new_[23700]_  = \new_[27641]_  & \new_[26821]_ ;
  assign \new_[23701]_  = ~\new_[26590]_  & ~\new_[29773]_ ;
  assign \new_[23702]_  = ~\new_[26974]_  | ~\new_[27720]_ ;
  assign \new_[23703]_  = \new_[28449]_  | \new_[29573]_ ;
  assign \new_[23704]_  = ~\new_[28561]_  | ~\new_[27568]_ ;
  assign \new_[23705]_  = ~\new_[27562]_  | ~\new_[30508]_ ;
  assign \new_[23706]_  = ~\new_[5994]_  | ~\new_[28878]_  | ~\new_[30158]_ ;
  assign \new_[23707]_  = \new_[27621]_  & \new_[27915]_ ;
  assign \new_[23708]_  = ~\new_[25055]_ ;
  assign \new_[23709]_  = \new_[27464]_  | \new_[30114]_ ;
  assign \new_[23710]_  = \new_[27568]_  & \new_[30628]_ ;
  assign \new_[23711]_  = ~\new_[27567]_  & ~\new_[29758]_ ;
  assign \new_[23712]_  = \new_[26917]_  | \new_[30186]_ ;
  assign \new_[23713]_  = ~\new_[28294]_  & ~\new_[30272]_ ;
  assign \new_[23714]_  = ~\new_[30423]_  | ~\new_[5984]_ ;
  assign \new_[23715]_  = ~\new_[26864]_  & ~\new_[28166]_ ;
  assign \new_[23716]_  = ~\new_[27654]_  & ~\new_[30581]_ ;
  assign \new_[23717]_  = ~\new_[26844]_  & ~\new_[30093]_ ;
  assign \new_[23718]_  = \new_[26757]_  | \new_[30543]_ ;
  assign \new_[23719]_  = ~\new_[25061]_ ;
  assign \new_[23720]_  = \new_[26721]_  | \new_[30055]_ ;
  assign \new_[23721]_  = ~\new_[29964]_  | ~\new_[5995]_ ;
  assign \new_[23722]_  = ~\new_[26798]_  | ~\new_[28245]_ ;
  assign \new_[23723]_  = \new_[27694]_  | \new_[30055]_ ;
  assign \new_[23724]_  = \new_[26793]_  | \new_[30058]_ ;
  assign \new_[23725]_  = \new_[28048]_  | \new_[28982]_ ;
  assign \new_[23726]_  = ~\new_[25469]_ ;
  assign \new_[23727]_  = ~\new_[27534]_  | ~\new_[28007]_ ;
  assign \new_[23728]_  = ~\new_[27579]_  | ~\new_[30628]_ ;
  assign \new_[23729]_  = ~\new_[26746]_  & ~\new_[29916]_ ;
  assign \new_[23730]_  = \new_[26798]_  & \new_[28930]_ ;
  assign \new_[23731]_  = ~\new_[25068]_ ;
  assign \new_[23732]_  = ~\new_[27624]_  | ~\new_[29082]_ ;
  assign \new_[23733]_  = \new_[27512]_  & \new_[28762]_ ;
  assign \new_[23734]_  = ~\new_[27564]_  & ~\new_[29970]_ ;
  assign \new_[23735]_  = ~\new_[27689]_  | ~\new_[30147]_ ;
  assign \new_[23736]_  = ~\new_[27628]_  | ~\new_[30034]_ ;
  assign \new_[23737]_  = ~\new_[27518]_  | ~\new_[29219]_ ;
  assign \new_[23738]_  = ~\new_[27717]_  & ~\new_[30157]_ ;
  assign \new_[23739]_  = ~\new_[27548]_  | ~\new_[30352]_ ;
  assign \new_[23740]_  = \new_[26703]_  | \new_[29754]_ ;
  assign \new_[23741]_  = ~\new_[26629]_  | ~\new_[29887]_ ;
  assign \new_[23742]_  = \new_[29249]_  | \new_[29375]_ ;
  assign \new_[23743]_  = \new_[26602]_  & \new_[30411]_ ;
  assign \new_[23744]_  = \new_[26817]_  | \new_[28236]_ ;
  assign \new_[23745]_  = ~\new_[27604]_  | ~\new_[30160]_ ;
  assign \new_[23746]_  = \new_[26661]_  | \new_[29272]_ ;
  assign \new_[23747]_  = ~\new_[27703]_  | ~\new_[29456]_ ;
  assign \new_[23748]_  = ~\new_[25080]_ ;
  assign \new_[23749]_  = ~\new_[25082]_ ;
  assign \new_[23750]_  = ~\new_[27697]_  | ~\new_[28905]_ ;
  assign \new_[23751]_  = \new_[29156]_  | \new_[29367]_ ;
  assign \new_[23752]_  = ~\new_[27724]_  & ~\new_[30095]_ ;
  assign \new_[23753]_  = ~\new_[26933]_  & ~\new_[30762]_ ;
  assign \new_[23754]_  = ~\new_[25253]_ ;
  assign \new_[23755]_  = \new_[27635]_  & \new_[28684]_ ;
  assign \new_[23756]_  = \new_[26864]_  | \new_[29568]_ ;
  assign \new_[23757]_  = ~\new_[26659]_  | ~\new_[28684]_ ;
  assign \new_[23758]_  = ~\new_[27749]_  | ~\new_[28640]_ ;
  assign \new_[23759]_  = ~\new_[27507]_  & ~\new_[29909]_ ;
  assign \new_[23760]_  = ~\new_[27735]_  | ~\new_[27691]_ ;
  assign \new_[23761]_  = \new_[27690]_  & \new_[28898]_ ;
  assign \new_[23762]_  = \new_[27757]_  | \new_[30407]_ ;
  assign \new_[23763]_  = \new_[27966]_  | \new_[29629]_ ;
  assign \new_[23764]_  = ~\new_[27895]_  & ~\new_[30618]_ ;
  assign \new_[23765]_  = ~\new_[27371]_  & ~\new_[29841]_ ;
  assign \new_[23766]_  = \new_[27503]_  | \new_[30044]_ ;
  assign \new_[23767]_  = \new_[26753]_  | \new_[28966]_ ;
  assign \new_[23768]_  = ~\new_[27418]_  & ~\new_[30010]_ ;
  assign \new_[23769]_  = ~\new_[5979]_  | ~\new_[28870]_  | ~\new_[30246]_ ;
  assign \new_[23770]_  = \new_[27578]_  | \new_[28236]_ ;
  assign \new_[23771]_  = ~\new_[26839]_  & ~\new_[30285]_ ;
  assign \new_[23772]_  = ~\new_[28438]_  & ~\new_[30285]_ ;
  assign \new_[23773]_  = \new_[26664]_  | \new_[29855]_ ;
  assign \new_[23774]_  = \new_[26838]_  | \new_[29272]_ ;
  assign \new_[23775]_  = ~\new_[27525]_  & ~\new_[30199]_ ;
  assign \new_[23776]_  = ~\new_[28774]_  | ~\new_[27904]_ ;
  assign \new_[23777]_  = ~\new_[27158]_  & ~\new_[29181]_ ;
  assign \new_[23778]_  = ~\new_[27537]_  & ~\new_[30423]_ ;
  assign \new_[23779]_  = ~\new_[28363]_  & ~\new_[29663]_ ;
  assign \new_[23780]_  = ~\new_[26948]_  | ~\new_[30726]_ ;
  assign \new_[23781]_  = \new_[26861]_  & \new_[29455]_ ;
  assign \new_[23782]_  = ~\new_[25101]_ ;
  assign \new_[23783]_  = \new_[27546]_  & \new_[30735]_ ;
  assign \new_[23784]_  = \new_[28413]_  | \new_[28236]_ ;
  assign \new_[23785]_  = ~\new_[27961]_  & ~\new_[30568]_ ;
  assign \new_[23786]_  = ~\new_[24973]_ ;
  assign \new_[23787]_  = ~\new_[27629]_  | ~\new_[29040]_ ;
  assign \new_[23788]_  = ~\new_[28536]_  & ~\new_[29068]_ ;
  assign \new_[23789]_  = \new_[27594]_  & \new_[28355]_ ;
  assign \new_[23790]_  = \new_[27532]_  | \new_[30064]_ ;
  assign \new_[23791]_  = \new_[27641]_  | \new_[30307]_ ;
  assign \new_[23792]_  = ~\new_[26679]_  | ~\new_[29874]_ ;
  assign \new_[23793]_  = ~\new_[26522]_ ;
  assign \new_[23794]_  = \new_[27528]_  | \new_[30053]_ ;
  assign \new_[23795]_  = \new_[27492]_  | \new_[30212]_ ;
  assign \new_[23796]_  = \new_[27028]_  | \new_[29445]_ ;
  assign \new_[23797]_  = ~\new_[28788]_  | ~\new_[26655]_ ;
  assign \new_[23798]_  = ~\new_[26706]_  & ~\new_[29181]_ ;
  assign \new_[23799]_  = ~\new_[28177]_  & ~\new_[29934]_ ;
  assign \new_[23800]_  = ~\new_[27657]_  | ~\new_[27474]_ ;
  assign \new_[23801]_  = ~\new_[25108]_ ;
  assign \new_[23802]_  = ~\new_[29664]_  | ~\new_[29492]_  | ~\new_[29142]_  | ~\new_[30191]_ ;
  assign \new_[23803]_  = ~\new_[26917]_  & ~\new_[29359]_ ;
  assign \new_[23804]_  = \new_[27474]_  & \new_[29537]_ ;
  assign \new_[23805]_  = \new_[27749]_  & \new_[29608]_ ;
  assign \new_[23806]_  = ~\new_[26712]_  & ~\new_[30115]_ ;
  assign \new_[23807]_  = ~\new_[31900]_  | ~\new_[27474]_  | ~\new_[29537]_ ;
  assign \new_[23808]_  = \new_[27655]_  | \new_[30055]_ ;
  assign \new_[23809]_  = ~\new_[27136]_  & ~\new_[30501]_ ;
  assign \new_[23810]_  = ~\new_[27356]_  | ~\new_[30084]_ ;
  assign \new_[23811]_  = ~\new_[26859]_  & ~\new_[30677]_ ;
  assign \new_[23812]_  = ~\new_[29335]_  | ~\new_[29688]_  | ~\new_[29655]_  | ~\new_[30023]_ ;
  assign \new_[23813]_  = (~\new_[28313]_  | ~\s7_data_i[17] ) & (~\new_[29707]_  | ~\s6_data_i[17] );
  assign \new_[23814]_  = ~\new_[27136]_  & ~\new_[30115]_ ;
  assign \new_[23815]_  = ~\new_[27661]_  & ~\new_[29384]_ ;
  assign \new_[23816]_  = ~\new_[29581]_  | ~\new_[27848]_ ;
  assign \new_[23817]_  = ~\new_[25112]_ ;
  assign \new_[23818]_  = ~\new_[25113]_ ;
  assign \new_[23819]_  = ~\new_[26784]_  & ~\new_[30157]_ ;
  assign \new_[23820]_  = \new_[27661]_  | \new_[29398]_ ;
  assign \new_[23821]_  = ~\new_[5999]_  | ~\new_[29685]_  | ~\new_[30147]_ ;
  assign \new_[23822]_  = ~\new_[27261]_  | ~\new_[27383]_ ;
  assign \new_[23823]_  = \new_[26852]_  & \new_[28964]_ ;
  assign \new_[23824]_  = ~\new_[26866]_  & ~\new_[29277]_ ;
  assign \new_[23825]_  = ~\new_[5997]_  | ~\new_[28926]_  | ~\new_[30084]_ ;
  assign \new_[23826]_  = ~\new_[27267]_  | ~\new_[30126]_ ;
  assign \new_[23827]_  = ~\new_[26591]_  & ~\new_[29096]_ ;
  assign \new_[23828]_  = ~\new_[25119]_ ;
  assign \new_[23829]_  = ~\new_[26764]_  | ~\new_[27596]_ ;
  assign \new_[23830]_  = ~\new_[25122]_ ;
  assign \new_[23831]_  = ~\new_[26760]_  | ~\new_[30579]_ ;
  assign \new_[23832]_  = \new_[29536]_  & \new_[28001]_ ;
  assign \new_[23833]_  = ~\new_[27705]_  & ~\new_[30265]_ ;
  assign \new_[23834]_  = ~\new_[28432]_  & ~\new_[29096]_ ;
  assign \new_[23835]_  = ~\new_[27441]_  & ~\new_[26824]_ ;
  assign \new_[23836]_  = \new_[27644]_  & \new_[26596]_ ;
  assign \new_[23837]_  = ~\new_[25131]_ ;
  assign \new_[23838]_  = \new_[28305]_  | \new_[28950]_ ;
  assign \new_[23839]_  = ~\new_[27559]_  | ~\new_[30610]_ ;
  assign \new_[23840]_  = \new_[26704]_  & \new_[28307]_ ;
  assign \new_[23841]_  = ~\new_[27771]_  & ~\new_[28357]_ ;
  assign \new_[23842]_  = ~\new_[26782]_  & ~\new_[29166]_ ;
  assign \new_[23843]_  = \new_[27622]_  & \new_[29226]_ ;
  assign \new_[23844]_  = ~\new_[25135]_ ;
  assign \new_[23845]_  = ~\new_[28867]_  | ~\new_[6090]_ ;
  assign \new_[23846]_  = \new_[27497]_  | \new_[29564]_ ;
  assign \new_[23847]_  = \new_[26813]_  & \new_[29557]_ ;
  assign \new_[23848]_  = ~\new_[24610]_ ;
  assign \new_[23849]_  = ~\new_[27196]_  | ~\new_[29897]_ ;
  assign \new_[23850]_  = ~\new_[27637]_  | ~\new_[30218]_ ;
  assign \new_[23851]_  = \new_[26738]_  | \new_[29898]_ ;
  assign \new_[23852]_  = \new_[26709]_  | \new_[29827]_ ;
  assign \new_[23853]_  = \new_[27704]_  & \new_[29168]_ ;
  assign \new_[23854]_  = ~\new_[27198]_  & ~\new_[30047]_ ;
  assign \new_[23855]_  = ~\new_[27080]_  | ~\new_[28355]_ ;
  assign \new_[23856]_  = ~\new_[27493]_  & ~\new_[30607]_ ;
  assign \new_[23857]_  = ~\new_[27493]_  | ~\new_[26593]_ ;
  assign \new_[23858]_  = \new_[29601]_  & \new_[30494]_ ;
  assign \new_[23859]_  = ~\new_[24743]_ ;
  assign \new_[23860]_  = ~\new_[27700]_  | ~\new_[29061]_ ;
  assign \new_[23861]_  = ~\new_[26632]_  & ~\new_[30047]_ ;
  assign \new_[23862]_  = ~\new_[26900]_  | ~\new_[30025]_ ;
  assign \new_[23863]_  = ~\new_[27623]_  & ~\new_[30066]_ ;
  assign \new_[23864]_  = ~\new_[27555]_  | ~\new_[30021]_ ;
  assign \new_[23865]_  = \new_[27652]_  | \new_[29383]_ ;
  assign \new_[23866]_  = ~\new_[24738]_ ;
  assign \new_[23867]_  = ~\new_[24737]_ ;
  assign \new_[23868]_  = \new_[27080]_  & \new_[29455]_ ;
  assign \new_[23869]_  = \new_[27533]_  | \new_[29383]_ ;
  assign \new_[23870]_  = ~\new_[25141]_ ;
  assign \new_[23871]_  = ~\new_[27557]_  & ~\new_[30584]_ ;
  assign \new_[23872]_  = ~\new_[28410]_  & ~\new_[28982]_ ;
  assign \new_[23873]_  = \new_[26999]_  & \new_[30728]_ ;
  assign \new_[23874]_  = ~\new_[24732]_ ;
  assign \new_[23875]_  = \new_[29474]_  & \new_[28762]_ ;
  assign \new_[23876]_  = ~\new_[25146]_ ;
  assign \new_[23877]_  = ~\new_[25149]_ ;
  assign \new_[23878]_  = ~\new_[26695]_  | ~\new_[27546]_ ;
  assign \new_[23879]_  = ~\new_[27378]_  | ~\new_[29563]_ ;
  assign \new_[23880]_  = ~\new_[28785]_  & ~\new_[27783]_ ;
  assign \new_[23881]_  = ~\new_[27696]_  & ~\new_[30741]_ ;
  assign \new_[23882]_  = \new_[28740]_  | \new_[29119]_ ;
  assign \new_[23883]_  = ~\new_[28415]_  & ~\new_[29119]_ ;
  assign \new_[23884]_  = ~\new_[25151]_ ;
  assign \new_[23885]_  = ~\new_[28193]_  & ~\new_[28933]_ ;
  assign \new_[23886]_  = ~\new_[6033]_  | ~\new_[30283]_  | ~\new_[30416]_ ;
  assign \new_[23887]_  = ~\new_[27636]_  | ~\new_[26833]_ ;
  assign \new_[23888]_  = ~\new_[26668]_  & (~\new_[30097]_  | ~\new_[5895]_ );
  assign \new_[23889]_  = ~\new_[26725]_  & (~\new_[30599]_  | ~\new_[6273]_ );
  assign \new_[23890]_  = ~\new_[27518]_  & ~\new_[27088]_ ;
  assign \new_[23891]_  = ~\new_[27733]_  & (~\new_[30320]_  | ~\new_[5896]_ );
  assign \new_[23892]_  = ~\new_[6069]_  | ~\new_[29802]_  | ~\new_[30647]_ ;
  assign \new_[23893]_  = ~\new_[6032]_  | ~\new_[29975]_  | ~\new_[30676]_ ;
  assign \new_[23894]_  = ~\new_[27960]_  & (~\new_[30678]_  | ~\new_[6043]_ );
  assign \new_[23895]_  = ~\new_[27630]_  & (~\new_[30686]_  | ~\new_[6208]_ );
  assign \new_[23896]_  = ~\new_[6216]_  | ~\new_[29897]_  | ~\new_[30262]_ ;
  assign \new_[23897]_  = ~\new_[27626]_  & (~\new_[30172]_  | ~\new_[5897]_ );
  assign \new_[23898]_  = ~\new_[27060]_  & (~\new_[30640]_  | ~\new_[6199]_ );
  assign \new_[23899]_  = ~\new_[26913]_  & (~\new_[29888]_  | ~\new_[5903]_ );
  assign \new_[23900]_  = ~\new_[31232]_  | ~\new_[30409]_  | ~\new_[29929]_ ;
  assign \new_[23901]_  = ~\new_[27745]_  | ~\new_[26762]_ ;
  assign \new_[23902]_  = ~\new_[27664]_  & (~\new_[30061]_  | ~\new_[5905]_ );
  assign \new_[23903]_  = ~\new_[6084]_  | ~\new_[30142]_  | ~\new_[30725]_ ;
  assign \new_[23904]_  = ~\new_[6184]_  | ~\new_[30218]_  | ~\new_[30352]_ ;
  assign \new_[23905]_  = ~\new_[27619]_  | ~\new_[27795]_ ;
  assign \new_[23906]_  = ~\new_[27835]_  & (~\new_[30198]_  | ~\new_[6195]_ );
  assign \new_[23907]_  = ~\new_[6210]_  | ~\new_[29877]_  | ~\new_[30645]_ ;
  assign \new_[23908]_  = ~\new_[27773]_  & ~\new_[26855]_ ;
  assign \new_[23909]_  = ~\new_[31440]_  | ~\new_[30146]_  | ~\new_[30728]_ ;
  assign \new_[23910]_  = ~\new_[27667]_  & (~\new_[30159]_  | ~\new_[5906]_ );
  assign \new_[23911]_  = ~\new_[27624]_  & ~\new_[27290]_ ;
  assign \new_[23912]_  = ~\new_[27766]_  & (~\new_[30667]_  | ~\new_[6191]_ );
  assign \new_[23913]_  = ~\new_[27665]_  & (~\new_[29863]_  | ~\new_[5904]_ );
  assign \new_[23914]_  = ~\new_[27746]_  | ~\new_[27334]_ ;
  assign \new_[23915]_  = ~\new_[5924]_  | ~\new_[29979]_  | ~\new_[30563]_ ;
  assign \new_[23916]_  = ~\new_[27698]_  & ~\new_[27711]_ ;
  assign \new_[23917]_  = ~\new_[27680]_  & (~\new_[29868]_  | ~\new_[31235]_ );
  assign \new_[23918]_  = ~\new_[5926]_  | ~\new_[30105]_  | ~\new_[30009]_ ;
  assign \new_[23919]_  = ~\new_[27954]_  & (~\new_[30297]_  | ~\new_[6086]_ );
  assign \new_[23920]_  = ~\new_[28507]_  | ~\new_[27964]_ ;
  assign \new_[23921]_  = ~\new_[28081]_  & ~\new_[27714]_ ;
  assign \new_[23922]_  = ~\new_[28233]_  & ~\new_[27132]_ ;
  assign \new_[23923]_  = ~\new_[27752]_  & (~\new_[30092]_  | ~\new_[5902]_ );
  assign \new_[23924]_  = ~\new_[26403]_ ;
  assign \new_[23925]_  = ~\new_[26636]_  & (~\new_[29762]_  | ~\new_[5898]_ );
  assign \new_[23926]_  = ~\new_[31712]_  | ~\new_[30160]_  | ~\new_[30037]_ ;
  assign \new_[23927]_  = ~\new_[6072]_  | ~\new_[30180]_  | ~\new_[30321]_ ;
  assign \new_[23928]_  = ~\new_[27659]_  & (~\new_[30513]_  | ~\new_[6037]_ );
  assign \new_[23929]_  = ~\new_[6040]_  | ~\new_[30337]_  | ~\new_[30754]_ ;
  assign \new_[23930]_  = ~\new_[27754]_  & (~\new_[30603]_  | ~\new_[6089]_ );
  assign \new_[23931]_  = ~\new_[28392]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[23932]_  = ~\new_[28223]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[23933]_  = ~\new_[6196]_  | ~\new_[29870]_  | ~\new_[30752]_ ;
  assign \new_[23934]_  = ~\new_[28726]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[23935]_  = ~\new_[29043]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[23936]_  = ~\new_[27985]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[23937]_  = ~\new_[26401]_ ;
  assign \new_[23938]_  = ~\new_[28714]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[23939]_  = \new_[29483]_  & \new_[28183]_ ;
  assign \new_[23940]_  = ~\new_[29865]_  | ~\new_[5900]_ ;
  assign \new_[23941]_  = ~\new_[29660]_  | ~\new_[5922]_ ;
  assign \new_[23942]_  = ~\new_[28768]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[23943]_  = ~\new_[28767]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[23944]_  = ~\new_[28136]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[23945]_  = ~\new_[28313]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[23946]_  = ~\new_[30290]_  | ~\new_[30556]_ ;
  assign \new_[23947]_  = ~\new_[27762]_  | ~\new_[27392]_ ;
  assign \new_[23948]_  = ~\new_[6078]_  | ~\new_[29813]_  | ~\new_[30630]_ ;
  assign \new_[23949]_  = ~\new_[6066]_  | ~\new_[29867]_  | ~\new_[30814]_ ;
  assign \new_[23950]_  = ~\new_[26860]_  & (~\new_[30635]_  | ~\new_[6079]_ );
  assign \new_[23951]_  = ~\new_[27589]_  | ~\new_[27588]_ ;
  assign \new_[23952]_  = ~\new_[27575]_  & (~\new_[30494]_  | ~\new_[6073]_ );
  assign \new_[23953]_  = (~\new_[28768]_  | ~\s5_data_i[17] ) & (~\new_[30457]_  | ~\s3_data_i[17] );
  assign \new_[23954]_  = ~\new_[6094]_  | ~\new_[30104]_  | ~\new_[30150]_ ;
  assign \new_[23955]_  = ~\new_[27447]_  & (~\new_[28859]_  | ~\new_[29808]_ );
  assign \new_[23956]_  = ~\new_[27545]_  & (~\new_[28988]_  | ~\new_[30233]_ );
  assign \new_[23957]_  = (~\new_[28136]_  | ~\s5_data_i[6] ) & (~\new_[29928]_  | ~\s3_data_i[6] );
  assign \new_[23958]_  = (~\new_[28714]_  | ~\s5_data_i[24] ) & (~\new_[30709]_  | ~\s3_data_i[24] );
  assign \new_[23959]_  = (~\s7_data_i[16]  | ~\new_[27985]_ ) & (~\s6_data_i[16]  | ~\new_[29708]_ );
  assign \new_[23960]_  = (~\new_[28714]_  | ~\s5_data_i[19] ) & (~\new_[30709]_  | ~\s3_data_i[19] );
  assign \new_[23961]_  = (~\new_[28136]_  | ~\s5_data_i[12] ) & (~\new_[29928]_  | ~\s3_data_i[12] );
  assign \new_[23962]_  = \new_[26727]_  | \new_[29565]_ ;
  assign \new_[23963]_  = (~\new_[28714]_  | ~\s5_data_i[22] ) & (~\new_[30709]_  | ~\s3_data_i[22] );
  assign \new_[23964]_  = (~\new_[28136]_  | ~\s5_data_i[1] ) & (~\new_[29928]_  | ~\s3_data_i[1] );
  assign \new_[23965]_  = (~\new_[28136]_  | ~\s5_data_i[13] ) & (~\new_[29928]_  | ~\s3_data_i[13] );
  assign \new_[23966]_  = (~\new_[28714]_  | ~\s5_data_i[21] ) & (~\new_[30709]_  | ~\s3_data_i[21] );
  assign \new_[23967]_  = (~\new_[28313]_  | ~\s7_data_i[21] ) & (~\new_[29707]_  | ~\s6_data_i[21] );
  assign \new_[23968]_  = ~\new_[25602]_ ;
  assign \new_[23969]_  = (~\new_[28313]_  | ~\s7_data_i[24] ) & (~\new_[29707]_  | ~\s6_data_i[24] );
  assign \new_[23970]_  = (~\new_[28392]_  | ~\s4_data_i[30] ) & (~\new_[29349]_  | ~\s0_data_i[30] );
  assign \new_[23971]_  = (~\new_[28768]_  | ~\s5_data_i[5] ) & (~\new_[30457]_  | ~\s3_data_i[5] );
  assign \new_[23972]_  = (~\new_[28768]_  | ~\s5_data_i[26] ) & (~\new_[30457]_  | ~\s3_data_i[26] );
  assign \new_[23973]_  = (~\new_[28392]_  | ~\s4_data_i[5] ) & (~\new_[29349]_  | ~\s0_data_i[5] );
  assign \new_[23974]_  = (~\new_[28136]_  | ~\s5_data_i[14] ) & (~\new_[29928]_  | ~\s3_data_i[14] );
  assign \new_[23975]_  = (~\s7_data_i[15]  | ~\new_[27985]_ ) & (~\s6_data_i[15]  | ~\new_[29708]_ );
  assign \new_[23976]_  = (~\new_[28714]_  | ~\s5_data_i[16] ) & (~\new_[30709]_  | ~\s3_data_i[16] );
  assign \new_[23977]_  = (~\new_[28313]_  | ~\s7_data_i[12] ) & (~\new_[29707]_  | ~\s6_data_i[12] );
  assign \new_[23978]_  = (~\new_[28714]_  | ~\s5_data_i[15] ) & (~\new_[30709]_  | ~\s3_data_i[15] );
  assign \new_[23979]_  = (~\new_[28768]_  | ~\s5_data_i[6] ) & (~\new_[30457]_  | ~\s3_data_i[6] );
  assign \new_[23980]_  = (~\new_[28136]_  | ~\s5_data_i[8] ) & (~\new_[29928]_  | ~\s3_data_i[8] );
  assign \new_[23981]_  = (~\new_[28714]_  | ~\s5_data_i[14] ) & (~\new_[30709]_  | ~\s3_data_i[14] );
  assign \new_[23982]_  = (~\s7_data_i[9]  | ~\new_[27985]_ ) & (~\s6_data_i[9]  | ~\new_[29708]_ );
  assign \new_[23983]_  = (~\s7_data_i[2]  | ~\new_[27985]_ ) & (~\s6_data_i[2]  | ~\new_[29708]_ );
  assign \new_[23984]_  = ~\new_[28904]_  | ~\new_[6269]_ ;
  assign \new_[23985]_  = ~\new_[27623]_  & ~\new_[30780]_ ;
  assign \new_[23986]_  = (~\new_[28768]_  | ~\s5_data_i[8] ) & (~\new_[30457]_  | ~\s3_data_i[8] );
  assign \new_[23987]_  = (~\s7_data_i[10]  | ~\new_[27985]_ ) & (~\s6_data_i[10]  | ~\new_[29708]_ );
  assign \new_[23988]_  = \new_[29758]_  & \new_[5931]_ ;
  assign \new_[23989]_  = (~\new_[28714]_  | ~\s5_data_i[11] ) & (~\new_[30709]_  | ~\s3_data_i[11] );
  assign \new_[23990]_  = (~\new_[28768]_  | ~\s5_data_i[29] ) & (~\new_[30457]_  | ~\s3_data_i[29] );
  assign \new_[23991]_  = (~\new_[28768]_  | ~\s5_data_i[19] ) & (~\new_[30457]_  | ~\s3_data_i[19] );
  assign \new_[23992]_  = ~\new_[26391]_ ;
  assign \new_[23993]_  = (~\new_[28223]_  | ~\s7_data_i[20] ) & (~\new_[28767]_  | ~\s6_data_i[20] );
  assign \new_[23994]_  = (~\new_[28714]_  | ~\s5_data_i[20] ) & (~\new_[30709]_  | ~\s3_data_i[20] );
  assign \new_[23995]_  = (~\new_[28392]_  | ~\s4_data_i[9] ) & (~\new_[29349]_  | ~\s0_data_i[9] );
  assign \new_[23996]_  = (~\new_[28223]_  | ~\s7_data_i[11] ) & (~\new_[28767]_  | ~\s6_data_i[11] );
  assign \new_[23997]_  = ~\new_[26219]_ ;
  assign \new_[23998]_  = (~\new_[28223]_  | ~\s7_data_i[26] ) & (~\new_[28767]_  | ~\s6_data_i[26] );
  assign \new_[23999]_  = ~\new_[25466]_ ;
  assign \new_[24000]_  = (~\new_[28714]_  | ~\s5_data_i[6] ) & (~\new_[30709]_  | ~\s3_data_i[6] );
  assign \new_[24001]_  = (~\new_[28313]_  | ~\s7_data_i[1] ) & (~\new_[29707]_  | ~\s6_data_i[1] );
  assign \new_[24002]_  = ~\new_[25550]_ ;
  assign \new_[24003]_  = (~\new_[28223]_  | ~\s7_data_i[12] ) & (~\new_[28767]_  | ~\s6_data_i[12] );
  assign \new_[24004]_  = (~\new_[28313]_  | ~\s7_data_i[5] ) & (~\new_[29707]_  | ~\s6_data_i[5] );
  assign \new_[24005]_  = ~\new_[29754]_  | ~\new_[6195]_ ;
  assign \new_[24006]_  = ~\new_[28904]_  | ~\new_[6085]_ ;
  assign \new_[24007]_  = (~\new_[28714]_  | ~\s5_data_i[3] ) & (~\new_[30709]_  | ~\s3_data_i[3] );
  assign \new_[24008]_  = ~\new_[26389]_ ;
  assign \new_[24009]_  = (~\new_[28714]_  | ~\s5_data_i[2] ) & (~\new_[30709]_  | ~\s3_data_i[2] );
  assign \new_[24010]_  = (~\new_[28768]_  | ~\s5_data_i[28] ) & (~\new_[30457]_  | ~\s3_data_i[28] );
  assign \new_[24011]_  = (~\new_[28714]_  | ~\s5_data_i[10] ) & (~\new_[30709]_  | ~\s3_data_i[10] );
  assign \new_[24012]_  = (~\new_[28223]_  | ~\s7_data_i[13] ) & (~\new_[28767]_  | ~\s6_data_i[13] );
  assign \new_[24013]_  = (~\new_[28392]_  | ~\s4_data_i[13] ) & (~\new_[29349]_  | ~\s0_data_i[13] );
  assign \new_[24014]_  = (~\new_[28768]_  | ~\s5_data_i[14] ) & (~\new_[30457]_  | ~\s3_data_i[14] );
  assign \new_[24015]_  = (~\new_[28313]_  | ~\s7_data_i[31] ) & (~\new_[29707]_  | ~\s6_data_i[31] );
  assign \new_[24016]_  = ~\new_[28372]_  & ~\new_[30272]_ ;
  assign \new_[24017]_  = (~\new_[28223]_  | ~\s7_data_i[14] ) & (~\new_[28767]_  | ~\s6_data_i[14] );
  assign \new_[24018]_  = (~\s7_data_i[20]  | ~\new_[27985]_ ) & (~\s6_data_i[20]  | ~\new_[29708]_ );
  assign \new_[24019]_  = (~\new_[28313]_  | ~\s7_data_i[28] ) & (~\new_[29707]_  | ~\s6_data_i[28] );
  assign \new_[24020]_  = ~\new_[30116]_  | ~\new_[6214]_ ;
  assign \new_[24021]_  = ~\new_[26976]_  & ~\new_[30151]_ ;
  assign \new_[24022]_  = (~\new_[28313]_  | ~\s7_data_i[27] ) & (~\new_[29707]_  | ~\s6_data_i[27] );
  assign \new_[24023]_  = (~\new_[28313]_  | ~\s7_data_i[26] ) & (~\new_[29707]_  | ~\s6_data_i[26] );
  assign \new_[24024]_  = (~\new_[28392]_  | ~\s4_data_i[15] ) & (~\new_[29349]_  | ~\s0_data_i[15] );
  assign \new_[24025]_  = (~\new_[28768]_  | ~\s5_data_i[16] ) & (~\new_[30457]_  | ~\s3_data_i[16] );
  assign \new_[24026]_  = (~\new_[28223]_  | ~\s7_data_i[16] ) & (~\new_[28767]_  | ~\s6_data_i[16] );
  assign \new_[24027]_  = (~\new_[28223]_  | ~\s7_data_i[17] ) & (~\new_[28767]_  | ~\s6_data_i[17] );
  assign \new_[24028]_  = \new_[27560]_  | \new_[30400]_ ;
  assign \new_[24029]_  = (~\new_[28313]_  | ~\s7_data_i[14] ) & (~\new_[29707]_  | ~\s6_data_i[14] );
  assign \new_[24030]_  = (~\new_[28392]_  | ~\s4_data_i[18] ) & (~\new_[29349]_  | ~\s0_data_i[18] );
  assign \new_[24031]_  = (~\s7_data_i[24]  | ~\new_[27985]_ ) & (~\s6_data_i[24]  | ~\new_[29708]_ );
  assign \new_[24032]_  = (~\new_[28313]_  | ~\s7_data_i[9] ) & (~\new_[29707]_  | ~\s6_data_i[9] );
  assign \new_[24033]_  = (~\new_[28313]_  | ~\s7_data_i[4] ) & (~\new_[29707]_  | ~\s6_data_i[4] );
  assign \new_[24034]_  = (~\s7_data_i[25]  | ~\new_[27985]_ ) & (~\s6_data_i[25]  | ~\new_[29708]_ );
  assign \new_[24035]_  = ~\new_[30732]_  | ~\new_[6085]_ ;
  assign \new_[24036]_  = (~\new_[28392]_  | ~\s4_data_i[22] ) & (~\new_[29349]_  | ~\s0_data_i[22] );
  assign \new_[24037]_  = (~\new_[28313]_  | ~\s7_data_i[0] ) & (~\new_[29707]_  | ~\s6_data_i[0] );
  assign \new_[24038]_  = (~\new_[28313]_  | ~\s7_data_i[8] ) & (~\new_[29707]_  | ~\s6_data_i[8] );
  assign \new_[24039]_  = ~\new_[29435]_  | ~\new_[5966]_ ;
  assign \new_[24040]_  = (~\new_[28313]_  | ~\s7_data_i[23] ) & (~\new_[29707]_  | ~\s6_data_i[23] );
  assign \new_[24041]_  = (~\new_[28714]_  | ~\s5_data_i[18] ) & (~\new_[30709]_  | ~\s3_data_i[18] );
  assign \new_[24042]_  = (~\s7_data_i[12]  | ~\new_[27985]_ ) & (~\s6_data_i[12]  | ~\new_[29708]_ );
  assign \new_[24043]_  = ~\new_[26387]_ ;
  assign \new_[24044]_  = ~\new_[29003]_  | ~\new_[29219]_ ;
  assign \new_[24045]_  = (~\new_[28136]_  | ~\s5_data_i[23] ) & (~\new_[29928]_  | ~\s3_data_i[23] );
  assign \new_[24046]_  = (~\new_[28313]_  | ~\s7_data_i[25] ) & (~\new_[29707]_  | ~\s6_data_i[25] );
  assign \new_[24047]_  = (~\new_[28768]_  | ~\s5_data_i[23] ) & (~\new_[30457]_  | ~\s3_data_i[23] );
  assign \new_[24048]_  = (~\new_[28714]_  | ~\s5_data_i[13] ) & (~\new_[30709]_  | ~\s3_data_i[13] );
  assign \new_[24049]_  = (~\new_[28714]_  | ~\s5_data_i[8] ) & (~\new_[30709]_  | ~\s3_data_i[8] );
  assign \new_[24050]_  = (~\s7_data_i[6]  | ~\new_[27985]_ ) & (~\s6_data_i[6]  | ~\new_[29708]_ );
  assign \new_[24051]_  = (~\new_[28768]_  | ~\s5_data_i[24] ) & (~\new_[30457]_  | ~\s3_data_i[24] );
  assign \new_[24052]_  = ~\new_[29660]_  | ~\new_[5991]_ ;
  assign \new_[24053]_  = (~\s7_data_i[26]  | ~\new_[27985]_ ) & (~\s6_data_i[26]  | ~\new_[29708]_ );
  assign \new_[24054]_  = ~\new_[25674]_ ;
  assign \new_[24055]_  = (~\new_[28714]_  | ~\s5_data_i[5] ) & (~\new_[30709]_  | ~\s3_data_i[5] );
  assign \new_[24056]_  = (~\new_[28136]_  | ~\s5_data_i[24] ) & (~\new_[29928]_  | ~\s3_data_i[24] );
  assign \new_[24057]_  = (~\new_[28136]_  | ~\s5_data_i[30] ) & (~\new_[29928]_  | ~\s3_data_i[30] );
  assign \new_[24058]_  = (~\new_[28768]_  | ~\s5_data_i[30] ) & (~\new_[30457]_  | ~\s3_data_i[30] );
  assign \new_[24059]_  = (~\new_[28313]_  | ~\s7_data_i[10] ) & (~\new_[29707]_  | ~\s6_data_i[10] );
  assign \new_[24060]_  = ~\new_[30579]_  & ~\new_[31104]_ ;
  assign \new_[24061]_  = (~\new_[28313]_  | ~\s7_data_i[30] ) & (~\new_[29707]_  | ~\s6_data_i[30] );
  assign \new_[24062]_  = (~\s7_data_i[8]  | ~\new_[27985]_ ) & (~\s6_data_i[8]  | ~\new_[29708]_ );
  assign \new_[24063]_  = ~\new_[25715]_ ;
  assign \new_[24064]_  = (~\new_[28313]_  | ~\s7_data_i[29] ) & (~\new_[29707]_  | ~\s6_data_i[29] );
  assign \new_[24065]_  = ~\new_[29410]_  | ~\new_[30413]_ ;
  assign \new_[24066]_  = (~\new_[28392]_  | ~\s4_data_i[23] ) & (~\new_[29349]_  | ~\s0_data_i[23] );
  assign \new_[24067]_  = (~\new_[28392]_  | ~\s4_data_i[27] ) & (~\new_[29349]_  | ~\s0_data_i[27] );
  assign \new_[24068]_  = (~\new_[28313]_  | ~\s7_data_i[11] ) & (~\new_[29707]_  | ~\s6_data_i[11] );
  assign \new_[24069]_  = (~\new_[28136]_  | ~\s5_data_i[26] ) & (~\new_[29928]_  | ~\s3_data_i[26] );
  assign \new_[24070]_  = (~\new_[28768]_  | ~\s5_data_i[27] ) & (~\new_[30457]_  | ~\s3_data_i[27] );
  assign \new_[24071]_  = (~\s7_data_i[7]  | ~\new_[27985]_ ) & (~\s6_data_i[7]  | ~\new_[29708]_ );
  assign \new_[24072]_  = (~\new_[28392]_  | ~\s4_data_i[28] ) & (~\new_[29349]_  | ~\s0_data_i[28] );
  assign \new_[24073]_  = (~\new_[28136]_  | ~\s5_data_i[27] ) & (~\new_[29928]_  | ~\s3_data_i[27] );
  assign \new_[24074]_  = ~\new_[27509]_  & ~\new_[27959]_ ;
  assign \new_[24075]_  = (~\new_[28313]_  | ~\s7_data_i[7] ) & (~\new_[29707]_  | ~\s6_data_i[7] );
  assign \new_[24076]_  = (~\new_[28223]_  | ~\s7_data_i[27] ) & (~\new_[28767]_  | ~\s6_data_i[27] );
  assign \new_[24077]_  = (~\s7_data_i[5]  | ~\new_[27985]_ ) & (~\s6_data_i[5]  | ~\new_[29708]_ );
  assign \new_[24078]_  = (~\s7_data_i[14]  | ~\new_[27985]_ ) & (~\s6_data_i[14]  | ~\new_[29708]_ );
  assign \new_[24079]_  = ~\new_[30186]_  | ~\new_[6001]_ ;
  assign \new_[24080]_  = ~\new_[28985]_  | ~\new_[29061]_ ;
  assign \new_[24081]_  = ~\new_[26383]_ ;
  assign \new_[24082]_  = (~\new_[28313]_  | ~\s7_data_i[13] ) & (~\new_[29707]_  | ~\s6_data_i[13] );
  assign \new_[24083]_  = (~\s7_data_i[11]  | ~\new_[27985]_ ) & (~\s6_data_i[11]  | ~\new_[29708]_ );
  assign \new_[24084]_  = (~\new_[28768]_  | ~\s5_data_i[25] ) & (~\new_[30457]_  | ~\s3_data_i[25] );
  assign \new_[24085]_  = (~\s7_data_i[13]  | ~\new_[27985]_ ) & (~\s6_data_i[13]  | ~\new_[29708]_ );
  assign \new_[24086]_  = (~\new_[28136]_  | ~\s5_data_i[22] ) & (~\new_[29928]_  | ~\s3_data_i[22] );
  assign \new_[24087]_  = (~\s7_data_i[21]  | ~\new_[27985]_ ) & (~\s6_data_i[21]  | ~\new_[29708]_ );
  assign \new_[24088]_  = ~\new_[26549]_ ;
  assign \new_[24089]_  = (~\new_[28223]_  | ~\s7_data_i[28] ) & (~\new_[28767]_  | ~\s6_data_i[28] );
  assign \new_[24090]_  = (~\new_[28313]_  | ~\s7_data_i[6] ) & (~\new_[29707]_  | ~\s6_data_i[6] );
  assign \new_[24091]_  = ~\new_[29660]_  | ~\new_[5992]_ ;
  assign \new_[24092]_  = (~\new_[28392]_  | ~\s4_data_i[24] ) & (~\new_[29349]_  | ~\s0_data_i[24] );
  assign \new_[24093]_  = (~\new_[28223]_  | ~\s7_data_i[24] ) & (~\new_[28767]_  | ~\s6_data_i[24] );
  assign \new_[24094]_  = ~\new_[26381]_ ;
  assign \new_[24095]_  = (~\new_[28223]_  | ~\s7_data_i[23] ) & (~\new_[28767]_  | ~\s6_data_i[23] );
  assign \new_[24096]_  = (~\new_[28223]_  | ~\s7_data_i[22] ) & (~\new_[28767]_  | ~\s6_data_i[22] );
  assign \new_[24097]_  = ~\new_[28894]_  | ~\new_[29597]_ ;
  assign \new_[24098]_  = (~\new_[28768]_  | ~\s5_data_i[22] ) & (~\new_[30457]_  | ~\s3_data_i[22] );
  assign \new_[24099]_  = ~\new_[29540]_  | ~\new_[5987]_ ;
  assign \new_[24100]_  = (~\new_[28392]_  | ~\s4_data_i[21] ) & (~\new_[29349]_  | ~\s0_data_i[21] );
  assign \new_[24101]_  = (~\new_[28313]_  | ~\s7_data_i[15] ) & (~\new_[29707]_  | ~\s6_data_i[15] );
  assign \new_[24102]_  = (~\new_[28223]_  | ~\s7_data_i[21] ) & (~\new_[28767]_  | ~\s6_data_i[21] );
  assign \new_[24103]_  = (~\new_[28223]_  | ~\s7_data_i[31] ) & (~\new_[28767]_  | ~\s6_data_i[31] );
  assign \new_[24104]_  = (~\new_[28768]_  | ~\s5_data_i[21] ) & (~\new_[30457]_  | ~\s3_data_i[21] );
  assign \new_[24105]_  = (~\new_[28392]_  | ~\s4_data_i[20] ) & (~\new_[29349]_  | ~\s0_data_i[20] );
  assign \new_[24106]_  = ~\new_[26246]_ ;
  assign \new_[24107]_  = (~\s7_data_i[4]  | ~\new_[27985]_ ) & (~\s6_data_i[4]  | ~\new_[29708]_ );
  assign \new_[24108]_  = (~\new_[28392]_  | ~\s4_data_i[19] ) & (~\new_[29349]_  | ~\s0_data_i[19] );
  assign \new_[24109]_  = (~\new_[28223]_  | ~\s7_data_i[19] ) & (~\new_[28767]_  | ~\s6_data_i[19] );
  assign \new_[24110]_  = (~\s7_data_i[29]  | ~\new_[27985]_ ) & (~\s6_data_i[29]  | ~\new_[29708]_ );
  assign \new_[24111]_  = ~\new_[30228]_  | ~\new_[6192]_ ;
  assign \new_[24112]_  = (~\new_[28223]_  | ~\s7_data_i[18] ) & (~\new_[28767]_  | ~\s6_data_i[18] );
  assign \new_[24113]_  = ~\new_[30329]_  & ~\new_[31042]_ ;
  assign \new_[24114]_  = (~\s7_data_i[0]  | ~\new_[27985]_ ) & (~\s6_data_i[0]  | ~\new_[29708]_ );
  assign \new_[24115]_  = (~\new_[28768]_  | ~\s5_data_i[18] ) & (~\new_[30457]_  | ~\s3_data_i[18] );
  assign \new_[24116]_  = (~\new_[28392]_  | ~\s4_data_i[17] ) & (~\new_[29349]_  | ~\s0_data_i[17] );
  assign \new_[24117]_  = ~\new_[28824]_  | ~\new_[6052]_ ;
  assign \new_[24118]_  = (~\new_[28223]_  | ~\s7_data_i[15] ) & (~\new_[28767]_  | ~\s6_data_i[15] );
  assign \new_[24119]_  = (~\new_[28768]_  | ~\s5_data_i[15] ) & (~\new_[30457]_  | ~\s3_data_i[15] );
  assign \new_[24120]_  = (~\new_[28392]_  | ~\s4_data_i[14] ) & (~\new_[29349]_  | ~\s0_data_i[14] );
  assign \new_[24121]_  = (~\s7_data_i[3]  | ~\new_[27985]_ ) & (~\s6_data_i[3]  | ~\new_[29708]_ );
  assign \new_[24122]_  = (~\new_[28768]_  | ~\s5_data_i[13] ) & (~\new_[30457]_  | ~\s3_data_i[13] );
  assign \new_[24123]_  = ~\new_[29810]_  | ~\new_[5967]_ ;
  assign \new_[24124]_  = (~\new_[28392]_  | ~\s4_data_i[12] ) & (~\new_[29349]_  | ~\s0_data_i[12] );
  assign \new_[24125]_  = (~\new_[28714]_  | ~\s5_data_i[1] ) & (~\new_[30709]_  | ~\s3_data_i[1] );
  assign \new_[24126]_  = ~\new_[28393]_  | ~\new_[6039]_ ;
  assign \new_[24127]_  = (~\new_[28768]_  | ~\s5_data_i[11] ) & (~\new_[30457]_  | ~\s3_data_i[11] );
  assign \new_[24128]_  = (~\new_[28768]_  | ~\s5_data_i[10] ) & (~\new_[30457]_  | ~\s3_data_i[10] );
  assign \new_[24129]_  = (~\new_[28223]_  | ~\s7_data_i[9] ) & (~\new_[28767]_  | ~\s6_data_i[9] );
  assign \new_[24130]_  = (~\new_[28313]_  | ~\s7_data_i[18] ) & (~\new_[29707]_  | ~\s6_data_i[18] );
  assign \new_[24131]_  = (~\new_[28392]_  | ~\s4_data_i[8] ) & (~\new_[29349]_  | ~\s0_data_i[8] );
  assign \new_[24132]_  = (~\new_[28392]_  | ~\s4_data_i[7] ) & (~\new_[29349]_  | ~\s0_data_i[7] );
  assign \new_[24133]_  = (~\new_[28223]_  | ~\s7_data_i[7] ) & (~\new_[28767]_  | ~\s6_data_i[7] );
  assign \new_[24134]_  = (~\new_[28768]_  | ~\s5_data_i[7] ) & (~\new_[30457]_  | ~\s3_data_i[7] );
  assign \new_[24135]_  = \new_[26874]_  & \new_[28194]_ ;
  assign \new_[24136]_  = (~\new_[28392]_  | ~\s4_data_i[6] ) & (~\new_[29349]_  | ~\s0_data_i[6] );
  assign \new_[24137]_  = (~\new_[28223]_  | ~\s7_data_i[6] ) & (~\new_[28767]_  | ~\s6_data_i[6] );
  assign \new_[24138]_  = (~\new_[28136]_  | ~\s5_data_i[0] ) & (~\new_[29928]_  | ~\s3_data_i[0] );
  assign \new_[24139]_  = (~\new_[28223]_  | ~\s7_data_i[5] ) & (~\new_[28767]_  | ~\s6_data_i[5] );
  assign \new_[24140]_  = (~\new_[28392]_  | ~\s4_data_i[4] ) & (~\new_[29349]_  | ~\s0_data_i[4] );
  assign \new_[24141]_  = (~\new_[28223]_  | ~\s7_data_i[4] ) & (~\new_[28767]_  | ~\s6_data_i[4] );
  assign \new_[24142]_  = (~\new_[28768]_  | ~\s5_data_i[4] ) & (~\new_[30457]_  | ~\s3_data_i[4] );
  assign \new_[24143]_  = (~\new_[28313]_  | ~\s7_data_i[19] ) & (~\new_[29707]_  | ~\s6_data_i[19] );
  assign \new_[24144]_  = (~\new_[28392]_  | ~\s4_data_i[3] ) & (~\new_[29349]_  | ~\s0_data_i[3] );
  assign \new_[24145]_  = (~\new_[28223]_  | ~\s7_data_i[3] ) & (~\new_[28767]_  | ~\s6_data_i[3] );
  assign \new_[24146]_  = (~\new_[28768]_  | ~\s5_data_i[3] ) & (~\new_[30457]_  | ~\s3_data_i[3] );
  assign \new_[24147]_  = (~\new_[28392]_  | ~\s4_data_i[2] ) & (~\new_[29349]_  | ~\s0_data_i[2] );
  assign \new_[24148]_  = (~\s7_data_i[19]  | ~\new_[27985]_ ) & (~\s6_data_i[19]  | ~\new_[29708]_ );
  assign \new_[24149]_  = ~\new_[30275]_  & ~\new_[29299]_ ;
  assign \new_[24150]_  = (~\new_[28768]_  | ~\s5_data_i[2] ) & (~\new_[30457]_  | ~\s3_data_i[2] );
  assign \new_[24151]_  = (~\new_[28136]_  | ~\s5_data_i[9] ) & (~\new_[29928]_  | ~\s3_data_i[9] );
  assign \new_[24152]_  = (~\new_[28392]_  | ~\s4_data_i[1] ) & (~\new_[29349]_  | ~\s0_data_i[1] );
  assign \new_[24153]_  = ~\new_[26077]_ ;
  assign \new_[24154]_  = (~\new_[28768]_  | ~\s5_data_i[1] ) & (~\new_[30457]_  | ~\s3_data_i[1] );
  assign \new_[24155]_  = \new_[30205]_  | \new_[31900]_ ;
  assign \new_[24156]_  = (~\s7_data_i[1]  | ~\new_[27985]_ ) & (~\s6_data_i[1]  | ~\new_[29708]_ );
  assign \new_[24157]_  = ~\new_[29401]_  | ~\new_[29186]_ ;
  assign \new_[24158]_  = (~\new_[28768]_  | ~\s5_data_i[31] ) & (~\new_[30457]_  | ~\s3_data_i[31] );
  assign \new_[24159]_  = (~\s7_data_i[30]  | ~\new_[27985]_ ) & (~\s6_data_i[30]  | ~\new_[29708]_ );
  assign \new_[24160]_  = ~\new_[29540]_  | ~\new_[6213]_ ;
  assign \new_[24161]_  = (~\new_[28136]_  | ~\s5_data_i[31] ) & (~\new_[29928]_  | ~\s3_data_i[31] );
  assign \new_[24162]_  = ~\new_[26038]_ ;
  assign \new_[24163]_  = (~\new_[28136]_  | ~\s5_data_i[29] ) & (~\new_[29928]_  | ~\s3_data_i[29] );
  assign \new_[24164]_  = (~\s7_data_i[18]  | ~\new_[27985]_ ) & (~\s6_data_i[18]  | ~\new_[29708]_ );
  assign \new_[24165]_  = (~\new_[28136]_  | ~\s5_data_i[28] ) & (~\new_[29928]_  | ~\s3_data_i[28] );
  assign \new_[24166]_  = ~\new_[26930]_  & ~\new_[30703]_ ;
  assign \new_[24167]_  = (~\new_[28223]_  | ~\s7_data_i[30] ) & (~\new_[28767]_  | ~\s6_data_i[30] );
  assign \new_[24168]_  = (~\new_[28136]_  | ~\s5_data_i[4] ) & (~\new_[29928]_  | ~\s3_data_i[4] );
  assign \new_[24169]_  = (~\new_[28136]_  | ~\s5_data_i[25] ) & (~\new_[29928]_  | ~\s3_data_i[25] );
  assign \new_[24170]_  = ~\new_[26882]_  & ~\new_[26853]_ ;
  assign \new_[24171]_  = (~\new_[28392]_  | ~\s4_data_i[26] ) & (~\new_[29349]_  | ~\s0_data_i[26] );
  assign \new_[24172]_  = (~\s7_data_i[22]  | ~\new_[27985]_ ) & (~\s6_data_i[22]  | ~\new_[29708]_ );
  assign \new_[24173]_  = (~\new_[28136]_  | ~\s5_data_i[21] ) & (~\new_[29928]_  | ~\s3_data_i[21] );
  assign \new_[24174]_  = (~\new_[28136]_  | ~\s5_data_i[20] ) & (~\new_[29928]_  | ~\s3_data_i[20] );
  assign \new_[24175]_  = (~\new_[28714]_  | ~\s5_data_i[31] ) & (~\new_[30709]_  | ~\s3_data_i[31] );
  assign \new_[24176]_  = (~\new_[28768]_  | ~\s5_data_i[0] ) & (~\new_[30457]_  | ~\s3_data_i[0] );
  assign \new_[24177]_  = (~\new_[28136]_  | ~\s5_data_i[19] ) & (~\new_[29928]_  | ~\s3_data_i[19] );
  assign \new_[24178]_  = (~\new_[28714]_  | ~\s5_data_i[30] ) & (~\new_[30709]_  | ~\s3_data_i[30] );
  assign \new_[24179]_  = (~\new_[28136]_  | ~\s5_data_i[17] ) & (~\new_[29928]_  | ~\s3_data_i[17] );
  assign \new_[24180]_  = (~\new_[28136]_  | ~\s5_data_i[16] ) & (~\new_[29928]_  | ~\s3_data_i[16] );
  assign \new_[24181]_  = (~\new_[28714]_  | ~\s5_data_i[29] ) & (~\new_[30709]_  | ~\s3_data_i[29] );
  assign \new_[24182]_  = (~\new_[28136]_  | ~\s5_data_i[15] ) & (~\new_[29928]_  | ~\s3_data_i[15] );
  assign \new_[24183]_  = (~\new_[28714]_  | ~\s5_data_i[28] ) & (~\new_[30709]_  | ~\s3_data_i[28] );
  assign \new_[24184]_  = ~\new_[26132]_ ;
  assign \new_[24185]_  = (~\new_[28136]_  | ~\s5_data_i[10] ) & (~\new_[29928]_  | ~\s3_data_i[10] );
  assign \new_[24186]_  = \new_[26908]_  | \new_[26894]_ ;
  assign \new_[24187]_  = (~\s7_data_i[27]  | ~\new_[27985]_ ) & (~\s6_data_i[27]  | ~\new_[29708]_ );
  assign \new_[24188]_  = (~\new_[28714]_  | ~\s5_data_i[25] ) & (~\new_[30709]_  | ~\s3_data_i[25] );
  assign \new_[24189]_  = ~\new_[29991]_  | ~\new_[6203]_ ;
  assign \new_[24190]_  = (~\new_[28313]_  | ~\s7_data_i[22] ) & (~\new_[29707]_  | ~\s6_data_i[22] );
  assign \new_[24191]_  = ~\new_[29130]_  & ~\new_[31724]_ ;
  assign \new_[24192]_  = ~\new_[28953]_  | ~\new_[6245]_ ;
  assign \new_[24193]_  = ~\new_[29324]_  | ~\new_[5924]_ ;
  assign \new_[24194]_  = ~\new_[28953]_  | ~\new_[6203]_ ;
  assign \new_[24195]_  = ~\new_[29681]_  & ~\new_[30874]_ ;
  assign \new_[24196]_  = ~\new_[30835]_  | ~\new_[6210]_ ;
  assign \new_[24197]_  = ~\new_[30228]_  | ~\new_[6214]_ ;
  assign \new_[24198]_  = ~\new_[30074]_  | ~\new_[5982]_ ;
  assign \new_[24199]_  = ~\new_[28993]_  & ~\new_[30925]_ ;
  assign \new_[24200]_  = ~\new_[29743]_  | ~\new_[6041]_ ;
  assign \new_[24201]_  = ~\new_[27817]_  & ~\new_[31276]_ ;
  assign \new_[24202]_  = ~\new_[28934]_  & ~\new_[31844]_ ;
  assign \new_[24203]_  = ~\new_[30404]_  | ~\new_[5969]_ ;
  assign \new_[24204]_  = ~\new_[29199]_  | ~\new_[30511]_ ;
  assign \new_[24205]_  = ~\new_[29991]_  | ~\new_[6245]_ ;
  assign \new_[24206]_  = ~\new_[30644]_  | ~\new_[5987]_ ;
  assign \new_[24207]_  = ~\new_[28981]_  | ~\new_[6204]_ ;
  assign \new_[24208]_  = ~\new_[27892]_  | ~\new_[31033]_ ;
  assign \new_[24209]_  = ~\new_[30074]_  | ~\new_[6063]_ ;
  assign \new_[24210]_  = ~\new_[29199]_  | ~\new_[6046]_ ;
  assign \new_[24211]_  = ~\new_[29199]_  | ~\new_[31143]_ ;
  assign \new_[24212]_  = ~\new_[28981]_  | ~\new_[31143]_ ;
  assign \new_[24213]_  = ~\new_[26163]_ ;
  assign \new_[24214]_  = ~\new_[30186]_  | ~\new_[6086]_ ;
  assign \new_[24215]_  = ~\new_[28393]_  | ~\new_[6038]_ ;
  assign \new_[24216]_  = \new_[29306]_  & \new_[6204]_ ;
  assign \new_[24217]_  = ~\new_[28067]_  | ~\new_[5932]_ ;
  assign \new_[24218]_  = \new_[30340]_  | \new_[31406]_ ;
  assign \new_[24219]_  = ~\new_[30205]_  & ~\new_[31104]_ ;
  assign \new_[24220]_  = ~\new_[28867]_  | ~\new_[5930]_ ;
  assign \new_[24221]_  = \new_[28682]_  & \new_[5985]_ ;
  assign \new_[24222]_  = \new_[30644]_  & \new_[6212]_ ;
  assign \new_[24223]_  = ~\new_[29145]_  & ~\new_[30969]_ ;
  assign \new_[24224]_  = ~\new_[29754]_  | ~\new_[31176]_ ;
  assign \new_[24225]_  = \new_[29787]_  | \new_[31837]_ ;
  assign \new_[24226]_  = ~\new_[28981]_  | ~\new_[6046]_ ;
  assign \new_[24227]_  = ~\new_[29291]_  & ~\new_[31665]_ ;
  assign \new_[24228]_  = ~\new_[29540]_  | ~\new_[30848]_ ;
  assign \new_[24229]_  = ~\new_[29999]_  | ~\new_[5996]_ ;
  assign \new_[24230]_  = ~\new_[29964]_  | ~\new_[6268]_ ;
  assign \new_[24231]_  = ~\new_[28393]_  | ~\new_[5965]_ ;
  assign \new_[24232]_  = ~\new_[30074]_  | ~\new_[5981]_ ;
  assign \new_[24233]_  = ~\new_[30116]_  | ~\new_[6192]_ ;
  assign \new_[24234]_  = ~\new_[28824]_  | ~\new_[6053]_ ;
  assign \new_[24235]_  = ~\new_[29042]_  & ~\new_[31421]_ ;
  assign \new_[24236]_  = ~\new_[29743]_  | ~\new_[5966]_ ;
  assign \new_[24237]_  = ~\new_[29743]_  | ~\new_[6176]_ ;
  assign \new_[24238]_  = ~\new_[29754]_  | ~\new_[6060]_ ;
  assign \new_[24239]_  = ~\new_[28824]_  | ~\new_[6031]_ ;
  assign \new_[24240]_  = ~\new_[27883]_  | ~\new_[5910]_ ;
  assign \new_[24241]_  = ~\new_[30270]_  | ~\new_[31235]_ ;
  assign \new_[24242]_  = ~\new_[28953]_  | ~\new_[6246]_ ;
  assign \new_[24243]_  = ~\new_[30018]_  | ~\new_[6217]_ ;
  assign \new_[24244]_  = ~\new_[28067]_  | ~\new_[6005]_ ;
  assign \new_[24245]_  = ~\new_[28067]_  | ~\new_[6006]_ ;
  assign \new_[24246]_  = \new_[28409]_  & \new_[5964]_ ;
  assign \new_[24247]_  = ~\new_[30732]_  | ~\new_[6082]_ ;
  assign \new_[24248]_  = ~\new_[28904]_  | ~\new_[6082]_ ;
  assign \new_[24249]_  = ~\new_[30186]_  | ~\new_[5929]_ ;
  assign \new_[24250]_  = ~\new_[30116]_  | ~\new_[6071]_ ;
  assign \new_[24251]_  = ~\new_[29999]_  | ~\new_[6268]_ ;
  assign \new_[24252]_  = ~\new_[29999]_  | ~\new_[5995]_ ;
  assign \new_[24253]_  = ~\new_[30404]_  | ~\new_[6044]_ ;
  assign \new_[24254]_  = ~\new_[28867]_  | ~\new_[6183]_ ;
  assign \new_[24255]_  = ~\new_[26188]_ ;
  assign \new_[24256]_  = ~\new_[29700]_  & ~\new_[29445]_ ;
  assign \new_[24257]_  = ~\new_[24946]_ ;
  assign \new_[24258]_  = ~\new_[29058]_  | ~\new_[6051]_ ;
  assign \new_[24259]_  = ~\new_[30329]_  | ~\new_[28967]_ ;
  assign \new_[24260]_  = ~\new_[28934]_  | ~\new_[30386]_ ;
  assign \new_[24261]_  = ~\new_[29550]_  | ~\new_[30164]_ ;
  assign \new_[24262]_  = ~\new_[26531]_ ;
  assign \new_[24263]_  = ~\new_[29159]_  | ~\new_[30426]_ ;
  assign \new_[24264]_  = ~\new_[29219]_  | ~\new_[29969]_ ;
  assign \new_[24265]_  = ~\new_[29062]_  & ~\new_[31423]_ ;
  assign \new_[24266]_  = ~\new_[30221]_  & ~\new_[5963]_ ;
  assign \new_[24267]_  = ~\new_[29934]_  | ~\new_[5904]_ ;
  assign \new_[24268]_  = ~\new_[30033]_  & ~\new_[30515]_ ;
  assign \new_[24269]_  = ~\new_[29062]_  & ~\new_[29181]_ ;
  assign \new_[24270]_  = ~\new_[29115]_  | ~\new_[6193]_ ;
  assign \new_[24271]_  = ~\new_[30075]_  | ~\new_[6076]_ ;
  assign \new_[24272]_  = ~\new_[30202]_  & ~\new_[30192]_ ;
  assign \new_[24273]_  = ~\new_[30467]_  & ~\new_[29750]_ ;
  assign \new_[24274]_  = ~\new_[24787]_ ;
  assign \new_[24275]_  = ~\new_[24960]_ ;
  assign \new_[24276]_  = ~\new_[26214]_ ;
  assign \new_[24277]_  = ~\new_[29772]_  | ~\new_[5907]_ ;
  assign \new_[24278]_  = ~\new_[30515]_  | ~\new_[6197]_ ;
  assign \new_[24279]_  = ~\new_[30586]_  | ~\new_[30271]_ ;
  assign \new_[24280]_  = ~\new_[28870]_  | ~\new_[29271]_ ;
  assign \new_[24281]_  = ~\new_[25925]_ ;
  assign \new_[24282]_  = \new_[29861]_  | \new_[29119]_ ;
  assign \new_[24283]_  = ~\new_[26217]_ ;
  assign \new_[24284]_  = ~\new_[29817]_  | ~\new_[29701]_ ;
  assign \new_[24285]_  = (~\new_[28714]_  | ~\s5_data_i[26] ) & (~\new_[30709]_  | ~\s3_data_i[26] );
  assign \new_[24286]_  = ~\new_[29220]_  | ~\new_[29003]_ ;
  assign \new_[24287]_  = ~\new_[30140]_  & ~\new_[30272]_ ;
  assign \new_[24288]_  = ~\new_[29810]_  | ~\new_[6032]_ ;
  assign \new_[24289]_  = ~\new_[28924]_  | ~\new_[29068]_ ;
  assign \new_[24290]_  = ~\new_[26222]_ ;
  assign \new_[24291]_  = ~\new_[26223]_ ;
  assign \new_[24292]_  = ~\new_[29032]_  | ~\new_[28050]_ ;
  assign \new_[24293]_  = ~\new_[30411]_  | ~\new_[29040]_ ;
  assign \new_[24294]_  = ~\new_[26225]_ ;
  assign \new_[24295]_  = ~\new_[29157]_  & ~\new_[29174]_ ;
  assign \new_[24296]_  = ~\new_[30515]_  | ~\new_[6057]_ ;
  assign \new_[24297]_  = ~\new_[30188]_  | ~\new_[6073]_ ;
  assign \new_[24298]_  = ~\new_[30710]_  & ~\new_[30656]_ ;
  assign \new_[24299]_  = ~\new_[30277]_  | ~\new_[5933]_ ;
  assign \new_[24300]_  = ~\new_[28845]_  | ~\new_[29550]_ ;
  assign \new_[24301]_  = ~\new_[24961]_ ;
  assign \new_[24302]_  = ~\new_[29397]_  | ~\new_[29401]_ ;
  assign \new_[24303]_  = ~\new_[30410]_  | ~\new_[26655]_ ;
  assign \new_[24304]_  = ~\new_[30145]_  | ~\new_[6033]_ ;
  assign \new_[24305]_  = ~\new_[29291]_  | ~\new_[29220]_ ;
  assign \new_[24306]_  = ~\new_[30519]_  | ~\new_[30169]_ ;
  assign \new_[24307]_  = ~\new_[26345]_ ;
  assign \new_[24308]_  = ~\new_[29271]_  | ~\new_[29221]_ ;
  assign \new_[24309]_  = ~\new_[30066]_  | ~\new_[31400]_ ;
  assign \new_[24310]_  = ~\new_[26253]_ ;
  assign \new_[24311]_  = ~\new_[29355]_  | ~\new_[28073]_ ;
  assign \new_[24312]_  = ~\new_[29564]_  & ~\new_[30305]_ ;
  assign \new_[24313]_  = ~\new_[30415]_  & ~\new_[30334]_ ;
  assign \new_[24314]_  = ~\new_[24712]_ ;
  assign \new_[24315]_  = ~\new_[28017]_  | ~\new_[6215]_ ;
  assign \new_[24316]_  = ~\new_[29354]_  & ~\new_[29564]_ ;
  assign \new_[24317]_  = ~\new_[30649]_  & ~\new_[30616]_ ;
  assign \new_[24318]_  = ~\new_[26260]_ ;
  assign \new_[24319]_  = ~\new_[29841]_  & ~\new_[30285]_ ;
  assign \new_[24320]_  = ~\new_[30497]_  | ~\new_[28837]_ ;
  assign \new_[24321]_  = \new_[30167]_  & \new_[31406]_ ;
  assign \new_[24322]_  = ~\new_[24688]_ ;
  assign \new_[24323]_  = ~\new_[30157]_  | ~\new_[31499]_ ;
  assign \new_[24324]_  = ~\new_[30525]_  | ~\new_[30410]_ ;
  assign \new_[24325]_  = ~\new_[24675]_ ;
  assign \new_[24326]_  = ~\new_[30314]_  | ~\new_[5911]_ ;
  assign \new_[24327]_  = ~\new_[30285]_  | ~\new_[5895]_ ;
  assign \new_[24328]_  = ~\new_[30253]_  & ~\new_[29930]_ ;
  assign \new_[24329]_  = ~\new_[26272]_ ;
  assign \new_[24330]_  = ~\new_[29671]_  & ~\new_[29944]_ ;
  assign \new_[24331]_  = ~\new_[30550]_  | ~\new_[27787]_ ;
  assign \new_[24332]_  = ~\new_[30135]_  & ~\new_[5966]_ ;
  assign \new_[24333]_  = ~\new_[28887]_  | ~\new_[29578]_ ;
  assign \new_[24334]_  = ~\new_[26275]_ ;
  assign \new_[24335]_  = ~\new_[30367]_  | ~\new_[30559]_ ;
  assign \new_[24336]_  = ~\new_[30270]_  | ~\new_[31033]_ ;
  assign \new_[24337]_  = ~\new_[24656]_ ;
  assign \new_[24338]_  = ~\new_[30008]_  | ~\new_[5905]_ ;
  assign \new_[24339]_  = ~\new_[29050]_  | ~\new_[30670]_ ;
  assign \new_[24340]_  = ~\new_[24642]_ ;
  assign \new_[24341]_  = ~\new_[24633]_ ;
  assign \new_[24342]_  = \new_[29944]_  | \new_[28950]_ ;
  assign \new_[24343]_  = ~\new_[29445]_  & ~\new_[28962]_ ;
  assign \new_[24344]_  = ~\new_[30058]_  & ~\new_[29934]_ ;
  assign \new_[24345]_  = ~\new_[30297]_  | ~\new_[29701]_ ;
  assign \new_[24346]_  = ~\new_[24621]_ ;
  assign \new_[24347]_  = ~\new_[28944]_  & ~\new_[29959]_ ;
  assign \new_[24348]_  = ~\new_[24619]_ ;
  assign \new_[24349]_  = ~\new_[30199]_  | ~\new_[6197]_ ;
  assign \new_[24350]_  = ~\new_[30651]_  | ~\new_[6061]_ ;
  assign \new_[24351]_  = ~\new_[30242]_  | ~\new_[28837]_ ;
  assign \new_[24352]_  = ~\new_[24609]_ ;
  assign \new_[24353]_  = ~\new_[30334]_  | ~\new_[5896]_ ;
  assign \new_[24354]_  = ~\new_[24599]_ ;
  assign \new_[24355]_  = ~\new_[29785]_  & ~\new_[5922]_ ;
  assign \new_[24356]_  = ~\new_[24596]_ ;
  assign \new_[24357]_  = ~\new_[30651]_  & ~\new_[30835]_ ;
  assign \new_[24358]_  = ~\new_[30835]_  & ~\new_[6211]_ ;
  assign \new_[24359]_  = ~\new_[29174]_  & ~\new_[29202]_ ;
  assign \new_[24360]_  = ~\new_[29902]_  & ~\new_[30044]_ ;
  assign \new_[24361]_  = ~\new_[24586]_ ;
  assign \new_[24362]_  = ~\new_[29629]_  & ~\new_[29744]_ ;
  assign \new_[24363]_  = ~\new_[29886]_  & ~\new_[27778]_ ;
  assign \new_[24364]_  = ~\new_[24583]_ ;
  assign \new_[24365]_  = ~\new_[26307]_ ;
  assign \new_[24366]_  = ~\new_[30526]_  | ~\new_[6211]_ ;
  assign \new_[24367]_  = ~\new_[24570]_ ;
  assign \new_[24368]_  = ~\new_[30030]_  | ~\new_[29195]_ ;
  assign \new_[24369]_  = ~\new_[30208]_  | ~\new_[5908]_ ;
  assign \new_[24370]_  = ~\new_[29930]_  | ~\new_[6199]_ ;
  assign \new_[24371]_  = \new_[26983]_  & \new_[26910]_ ;
  assign \new_[24372]_  = ~\new_[30599]_  | ~\new_[28967]_ ;
  assign \new_[24373]_  = ~\new_[29254]_  | ~\new_[6067]_ ;
  assign \new_[24374]_  = ~\new_[29987]_  & ~\new_[28819]_ ;
  assign \new_[24375]_  = ~\new_[30265]_  | ~\new_[6186]_ ;
  assign \new_[24376]_  = ~\new_[26326]_ ;
  assign \new_[24377]_  = ~\new_[30731]_  | ~\new_[29971]_ ;
  assign \new_[24378]_  = ~\new_[28818]_  | ~\new_[29854]_ ;
  assign \new_[24379]_  = ~\new_[29748]_  & ~\new_[6202]_ ;
  assign \new_[24380]_  = ~\new_[29745]_  & ~\new_[6087]_ ;
  assign \new_[24381]_  = ~\new_[29815]_  | ~\new_[6043]_ ;
  assign \new_[24382]_  = ~\new_[29909]_  | ~\new_[6037]_ ;
  assign \new_[24383]_  = ~\new_[27802]_  | ~\new_[5922]_ ;
  assign \new_[24384]_  = ~\new_[30526]_  | ~\new_[30897]_ ;
  assign \new_[24385]_  = (~\new_[28136]_  | ~\s5_data_i[7] ) & (~\new_[29928]_  | ~\s3_data_i[7] );
  assign \new_[24386]_  = ~\new_[26548]_ ;
  assign \new_[24387]_  = ~\new_[29223]_  | ~\new_[30232]_ ;
  assign \new_[24388]_  = ~\new_[29907]_  & ~\new_[28183]_ ;
  assign \new_[24389]_  = ~\new_[26655]_  | ~\new_[6048]_ ;
  assign \new_[24390]_  = ~\new_[29082]_  | ~\new_[28245]_ ;
  assign \new_[24391]_  = ~\new_[29186]_  | ~\new_[5972]_ ;
  assign \new_[24392]_  = ~\new_[26453]_ ;
  assign \new_[24393]_  = ~\new_[30314]_  | ~\new_[6042]_ ;
  assign \new_[24394]_  = ~\new_[26921]_  & ~\new_[26922]_ ;
  assign \new_[24395]_  = ~\new_[26341]_ ;
  assign \new_[24396]_  = ~\new_[29455]_  | ~\new_[28850]_ ;
  assign \new_[24397]_  = ~\new_[30145]_  | ~\new_[6034]_ ;
  assign \new_[24398]_  = ~\new_[26470]_ ;
  assign \new_[24399]_  = ~\new_[26467]_ ;
  assign \new_[24400]_  = ~\new_[28930]_  | ~\new_[29082]_ ;
  assign \new_[24401]_  = ~\new_[28317]_  & ~\new_[30253]_ ;
  assign \new_[24402]_  = ~\new_[26350]_ ;
  assign \new_[24403]_  = ~\new_[29040]_  | ~\new_[30117]_ ;
  assign \new_[24404]_  = ~\new_[30042]_  | ~\new_[6094]_ ;
  assign \new_[24405]_  = ~\new_[28926]_  | ~\new_[29608]_ ;
  assign \new_[24406]_  = ~\new_[26354]_ ;
  assign \new_[24407]_  = ~\new_[28935]_  | ~\new_[5995]_ ;
  assign \new_[24408]_  = ~\new_[30386]_  | ~\new_[29192]_ ;
  assign \new_[24409]_  = ~\new_[30254]_  | ~\new_[6211]_ ;
  assign \new_[24410]_  = ~\new_[26356]_ ;
  assign \new_[24411]_  = ~\new_[26915]_  | ~\new_[26899]_ ;
  assign \new_[24412]_  = ~\new_[29238]_  & ~\new_[30188]_ ;
  assign \new_[24413]_  = ~\new_[30623]_  | ~\new_[26842]_ ;
  assign \new_[24414]_  = ~\new_[25330]_ ;
  assign \new_[24415]_  = ~\new_[30132]_  | ~\new_[30650]_ ;
  assign \new_[24416]_  = ~\new_[30656]_  & ~\new_[29238]_ ;
  assign \new_[24417]_  = ~\new_[24627]_ ;
  assign \new_[24418]_  = ~\new_[29168]_  | ~\new_[29032]_ ;
  assign \new_[24419]_  = ~\new_[28989]_  | ~\new_[29983]_ ;
  assign \new_[24420]_  = ~\new_[26209]_ ;
  assign \new_[24421]_  = ~\new_[29445]_  & ~\new_[30219]_ ;
  assign \new_[24422]_  = ~\new_[26560]_ ;
  assign \new_[24423]_  = ~\new_[30063]_  & ~\new_[29077]_ ;
  assign \new_[24424]_  = ~\new_[30627]_  | ~\new_[29015]_ ;
  assign \new_[24425]_  = ~\new_[30597]_  & ~\new_[28846]_ ;
  assign \new_[24426]_  = ~\new_[28017]_  | ~\new_[30998]_ ;
  assign \new_[24427]_  = ~\new_[30198]_  | ~\new_[29015]_ ;
  assign \new_[24428]_  = ~\new_[29685]_  | ~\new_[29571]_ ;
  assign \new_[24429]_  = ~\new_[25975]_ ;
  assign \new_[24430]_  = ~\new_[28595]_  & ~\new_[29595]_ ;
  assign \new_[24431]_  = ~\new_[30297]_  & ~\new_[28884]_ ;
  assign \new_[24432]_  = ~\new_[30515]_  & ~\new_[29452]_ ;
  assign \new_[24433]_  = ~\new_[30426]_  | ~\new_[29435]_ ;
  assign \new_[24434]_  = ~\new_[28979]_  & ~\new_[6056]_ ;
  assign \new_[24435]_  = ~\new_[25505]_ ;
  assign \new_[24436]_  = ~\new_[29212]_  | ~\new_[29593]_ ;
  assign \new_[24437]_  = ~\new_[25508]_ ;
  assign \new_[24438]_  = ~\new_[25460]_ ;
  assign \new_[24439]_  = ~\new_[29994]_  | ~\new_[5983]_ ;
  assign \new_[24440]_  = ~\new_[29047]_  & ~\new_[29629]_ ;
  assign \new_[24441]_  = ~\new_[26575]_ ;
  assign \new_[24442]_  = ~\new_[26398]_ ;
  assign \new_[24443]_  = ~\new_[25254]_ ;
  assign \new_[24444]_  = ~\new_[30297]_  | ~\new_[27778]_ ;
  assign \new_[24445]_  = ~\new_[29583]_  | ~\new_[30315]_ ;
  assign \new_[24446]_  = ~\new_[30642]_  & ~\new_[30557]_ ;
  assign \new_[24447]_  = ~\new_[29608]_  | ~\new_[29038]_ ;
  assign \new_[24448]_  = ~\new_[25006]_ ;
  assign \new_[24449]_  = ~\new_[30139]_  & ~\new_[6046]_ ;
  assign \new_[24450]_  = ~\new_[24760]_ ;
  assign \new_[24451]_  = ~\new_[30326]_  & ~\new_[30423]_ ;
  assign \new_[24452]_  = ~\new_[29038]_  | ~\new_[28640]_ ;
  assign \new_[24453]_  = ~\new_[29810]_  & ~\new_[29746]_ ;
  assign \new_[24454]_  = ~\new_[30010]_  | ~\new_[6194]_ ;
  assign \new_[24455]_  = ~\new_[24788]_ ;
  assign \new_[24456]_  = ~\new_[24783]_ ;
  assign \new_[24457]_  = ~\new_[28017]_  | ~\new_[31499]_ ;
  assign \new_[24458]_  = ~\new_[24776]_ ;
  assign \new_[24459]_  = ~\new_[28872]_  | ~\new_[29394]_ ;
  assign \new_[24460]_  = ~\new_[29978]_  | ~\new_[29064]_ ;
  assign \new_[24461]_  = ~\new_[26427]_ ;
  assign \new_[24462]_  = ~\new_[25775]_ ;
  assign \new_[24463]_  = (~\new_[28714]_  | ~\s5_data_i[17] ) & (~\new_[30709]_  | ~\s3_data_i[17] );
  assign \new_[24464]_  = ~\new_[26433]_ ;
  assign \new_[24465]_  = ~\new_[24758]_ ;
  assign \new_[24466]_  = ~\new_[29268]_  | ~\new_[29056]_ ;
  assign \new_[24467]_  = ~\new_[26543]_ ;
  assign \new_[24468]_  = ~\new_[29150]_  | ~\new_[29397]_ ;
  assign \new_[24469]_  = ~\new_[24751]_ ;
  assign \new_[24470]_  = ~\new_[28850]_  | ~\new_[28355]_ ;
  assign \new_[24471]_  = ~\new_[26440]_ ;
  assign \new_[24472]_  = ~\new_[30230]_  | ~\new_[6174]_ ;
  assign \new_[24473]_  = ~\new_[30249]_  | ~\new_[5898]_ ;
  assign \new_[24474]_  = ~\new_[29029]_  & ~\new_[30332]_ ;
  assign \new_[24475]_  = ~\new_[26353]_ ;
  assign \new_[24476]_  = ~\new_[27827]_  & ~\new_[26934]_ ;
  assign \new_[24477]_  = ~\new_[26452]_ ;
  assign \new_[24478]_  = ~\new_[26459]_ ;
  assign \new_[24479]_  = ~\new_[26455]_ ;
  assign \new_[24480]_  = ~\new_[26457]_ ;
  assign \new_[24481]_  = ~\new_[26460]_ ;
  assign \new_[24482]_  = ~\new_[24647]_ ;
  assign \new_[24483]_  = ~\new_[26912]_  | ~\new_[29831]_ ;
  assign \new_[24484]_  = ~\new_[27675]_  | ~\new_[29386]_ ;
  assign \new_[24485]_  = ~\new_[27458]_  | ~\new_[28542]_ ;
  assign \new_[24486]_  = (~\s7_data_i[23]  | ~\new_[27985]_ ) & (~\s6_data_i[23]  | ~\new_[29708]_ );
  assign \new_[24487]_  = ~\new_[28846]_  & ~\new_[28944]_ ;
  assign \new_[24488]_  = (~\new_[28714]_  | ~\s5_data_i[27] ) & (~\new_[30709]_  | ~\s3_data_i[27] );
  assign \new_[24489]_  = ~\new_[24538]_ ;
  assign \new_[24490]_  = ~\new_[27504]_  & ~\new_[29959]_ ;
  assign \new_[24491]_  = ~\new_[28836]_  | ~\new_[30327]_ ;
  assign \new_[24492]_  = ~\new_[27715]_  | ~\new_[31712]_ ;
  assign \new_[24493]_  = ~\new_[26482]_ ;
  assign \new_[24494]_  = ~\new_[26484]_ ;
  assign \new_[24495]_  = ~\new_[26510]_ ;
  assign \new_[24496]_  = ~\new_[26965]_  | ~\new_[27737]_ ;
  assign \new_[24497]_  = ~\new_[30093]_  | ~\new_[6049]_ ;
  assign \new_[24498]_  = ~\new_[30840]_  & ~\new_[29508]_ ;
  assign \new_[24499]_  = ~\new_[30309]_  & ~\new_[29647]_ ;
  assign \new_[24500]_  = ~\new_[26509]_ ;
  assign \new_[24501]_  = ~\new_[24660]_ ;
  assign \new_[24502]_  = (~\new_[28136]_  | ~\s5_data_i[2] ) & (~\new_[29928]_  | ~\s3_data_i[2] );
  assign \new_[24503]_  = (~\new_[28313]_  | ~\s7_data_i[2] ) & (~\new_[29707]_  | ~\s6_data_i[2] );
  assign \new_[24504]_  = (~\new_[28223]_  | ~\s7_data_i[0] ) & (~\new_[28767]_  | ~\s6_data_i[0] );
  assign \new_[24505]_  = ~\new_[29505]_  & ~\new_[30129]_ ;
  assign \new_[24506]_  = ~\new_[26995]_  & ~\new_[30204]_ ;
  assign \new_[24507]_  = ~\new_[29787]_  | ~\new_[30034]_ ;
  assign \new_[24508]_  = ~\new_[30232]_  | ~\new_[29159]_ ;
  assign \new_[24509]_  = ~\new_[26529]_ ;
  assign \new_[24510]_  = ~\new_[24754]_ ;
  assign \new_[24511]_  = ~\new_[26336]_ ;
  assign \new_[24512]_  = ~\new_[29907]_  | ~\new_[27883]_ ;
  assign \new_[24513]_  = ~\new_[27787]_  | ~\new_[6046]_ ;
  assign \new_[24514]_  = ~\new_[30057]_  | ~\new_[28833]_ ;
  assign \new_[24515]_  = ~\new_[30025]_  & ~\new_[6005]_ ;
  assign \new_[24516]_  = (~\s7_data_i[17]  | ~\new_[27985]_ ) & (~\s6_data_i[17]  | ~\new_[29708]_ );
  assign \new_[24517]_  = \new_[26888]_  | \new_[30325]_ ;
  assign \new_[24518]_  = (~\new_[28136]_  | ~\s5_data_i[18] ) & (~\new_[29928]_  | ~\s3_data_i[18] );
  assign \new_[24519]_  = (~\new_[28136]_  | ~\s5_data_i[5] ) & (~\new_[29928]_  | ~\s3_data_i[5] );
  assign \new_[24520]_  = ~\new_[29629]_  & ~\new_[30339]_ ;
  assign \new_[24521]_  = ~\new_[26551]_ ;
  assign \new_[24522]_  = \new_[27382]_  & \new_[26599]_ ;
  assign \new_[24523]_  = ~\new_[28883]_  | ~\new_[29465]_ ;
  assign \new_[24524]_  = \new_[27552]_  | \new_[29827]_ ;
  assign \new_[24525]_  = ~\new_[30210]_  | ~\new_[27802]_ ;
  assign \new_[24526]_  = ~\new_[26676]_  | ~\new_[30726]_ ;
  assign \new_[24527]_  = ~\new_[26474]_ ;
  assign \new_[24528]_  = ~\new_[26557]_ ;
  assign \new_[24529]_  = ~\new_[30279]_  | ~\new_[28877]_ ;
  assign \new_[24530]_  = \new_[27054]_  & \new_[27779]_ ;
  assign \new_[24531]_  = \new_[26735]_  | \new_[29899]_ ;
  assign \new_[24532]_  = ~\new_[30445]_  | ~\new_[6186]_ ;
  assign \new_[24533]_  = (~\new_[28392]_  | ~\s4_data_i[29] ) & (~\new_[29349]_  | ~\s0_data_i[29] );
  assign \new_[24534]_  = (~\new_[30200]_  | ~\s11_data_i[21] ) & (~\new_[29428]_  | ~\s8_data_i[21] );
  assign \new_[24535]_  = \new_[28187]_  | \new_[30342]_ ;
  assign \new_[24536]_  = (~\new_[30227]_  | ~\s10_data_i[16] ) & (~\new_[29706]_  | ~\s9_data_i[16] );
  assign \new_[24537]_  = \new_[29481]_  & \new_[28579]_ ;
  assign \new_[24538]_  = ~\new_[28197]_  | ~\new_[5927]_ ;
  assign \new_[24539]_  = (~\new_[29628]_  | ~\s4_data_i[21] ) & (~\new_[29258]_  | ~\s0_data_i[21] );
  assign \new_[24540]_  = (~\new_[30200]_  | ~\s11_data_i[14] ) & (~\new_[29428]_  | ~\s8_data_i[14] );
  assign \new_[24541]_  = ~\new_[30046]_  | ~\new_[29745]_ ;
  assign \new_[24542]_  = ~\new_[26591]_ ;
  assign \new_[24543]_  = ~\new_[26595]_ ;
  assign \new_[24544]_  = ~\new_[30196]_  | ~\new_[30032]_ ;
  assign \new_[24545]_  = (~\new_[30193]_  | ~\s7_data_i[23] ) & (~\new_[29298]_  | ~\s6_data_i[23] );
  assign \new_[24546]_  = (~\new_[29710]_  | ~\s10_data_i[1] ) & (~\new_[29024]_  | ~\s9_data_i[1] );
  assign \new_[24547]_  = ~\new_[27861]_ ;
  assign \new_[24548]_  = (~\new_[29149]_  | ~\s4_data_i[10] ) & (~\new_[29651]_  | ~\s0_data_i[10] );
  assign \new_[24549]_  = ~\new_[26611]_ ;
  assign \new_[24550]_  = ~\new_[26590]_ ;
  assign \new_[24551]_  = (~\new_[30060]_  | ~\s7_data_i[22] ) & (~\new_[29704]_  | ~\s6_data_i[22] );
  assign \new_[24552]_  = (~\new_[30260]_  | ~\s11_data_i[28] ) & (~\new_[29670]_  | ~\s8_data_i[28] );
  assign \new_[24553]_  = ~\new_[26612]_ ;
  assign \new_[24554]_  = ~\new_[28857]_  & ~\new_[28285]_ ;
  assign \new_[24555]_  = ~\new_[29889]_  & ~\new_[30011]_ ;
  assign \new_[24556]_  = (~\new_[29045]_  | ~\s10_data_i[4] ) & (~\new_[29951]_  | ~\s9_data_i[4] );
  assign \new_[24557]_  = ~\new_[26617]_ ;
  assign \new_[24558]_  = ~\new_[26585]_ ;
  assign \new_[24559]_  = (~\new_[29021]_  | ~\s10_data_i[23] ) & (~\new_[29709]_  | ~\s9_data_i[23] );
  assign \new_[24560]_  = (~\s14_data_i[28]  | ~\new_[30026]_ ) & (~\s12_data_i[28]  | ~\new_[29711]_ );
  assign \new_[24561]_  = ~\new_[29223]_  & ~\new_[28816]_ ;
  assign \new_[24562]_  = (~\new_[30311]_  | ~\s11_data_i[16] ) & (~\new_[29636]_  | ~\s8_data_i[16] );
  assign \new_[24563]_  = ~\new_[29869]_  | ~\new_[29978]_ ;
  assign \new_[24564]_  = ~\new_[30117]_  | ~\new_[6088]_ ;
  assign \new_[24565]_  = \new_[28586]_  | \new_[29966]_ ;
  assign \new_[24566]_  = ~\new_[30135]_  & ~\new_[28816]_ ;
  assign \new_[24567]_  = (~\new_[29149]_  | ~\s4_data_i[30] ) & (~\new_[29651]_  | ~\s0_data_i[30] );
  assign \new_[24568]_  = ~\new_[28770]_  | ~\new_[31479]_ ;
  assign \new_[24569]_  = ~\new_[26640]_ ;
  assign \new_[24570]_  = ~\new_[26657]_  & ~\new_[29692]_ ;
  assign \new_[24571]_  = ~\new_[32057]_ ;
  assign \new_[24572]_  = ~\new_[27798]_ ;
  assign \new_[24573]_  = ~\new_[28776]_  | ~\new_[31614]_ ;
  assign \new_[24574]_  = (~\new_[30311]_  | ~\s11_data_i[25] ) & (~\new_[29636]_  | ~\s8_data_i[25] );
  assign \new_[24575]_  = (~\new_[29025]_  | ~\s5_data_i[19] ) & (~\new_[30469]_  | ~\s3_data_i[19] );
  assign \new_[24576]_  = (~\new_[29705]_  | ~\s10_data_i[28] ) & (~\new_[30354]_  | ~\s9_data_i[28] );
  assign \new_[24577]_  = ~\new_[27649]_ ;
  assign \new_[24578]_  = ~\new_[28238]_  & (~\new_[30248]_  | ~\new_[6082]_ );
  assign \new_[24579]_  = (~\s10_data_i[12]  | ~\new_[29749]_ ) & (~\s9_data_i[12]  | ~\new_[29034]_ );
  assign \new_[24580]_  = ~\new_[26665]_ ;
  assign \new_[24581]_  = (~\new_[29976]_  | ~\s14_data_i[22] ) & (~\new_[28957]_  | ~\s12_data_i[22] );
  assign \new_[24582]_  = ~\new_[26669]_ ;
  assign \new_[24583]_  = ~\new_[30741]_  & ~\new_[27802]_ ;
  assign \new_[24584]_  = ~\new_[26672]_ ;
  assign \new_[24585]_  = ~\new_[26670]_ ;
  assign \new_[24586]_  = ~\new_[29151]_  & ~\new_[29885]_ ;
  assign \new_[24587]_  = (~\new_[30060]_  | ~\s7_data_i[25] ) & (~\new_[29704]_  | ~\s6_data_i[25] );
  assign \new_[24588]_  = (~\new_[29628]_  | ~\s4_data_i[25] ) & (~\new_[29258]_  | ~\s0_data_i[25] );
  assign \new_[24589]_  = ~\new_[29631]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[24590]_  = (~\new_[29976]_  | ~\s14_data_i[27] ) & (~\new_[28957]_  | ~\s12_data_i[27] );
  assign \new_[24591]_  = ~\new_[28280]_  | ~\new_[6000]_ ;
  assign \new_[24592]_  = (~\new_[30181]_  | ~\s14_data_i[26] ) & (~\new_[29640]_  | ~\s12_data_i[26] );
  assign \new_[24593]_  = \new_[28123]_  & \new_[29550]_ ;
  assign \new_[24594]_  = ~\new_[28306]_  & ~\new_[30225]_ ;
  assign \new_[24595]_  = ~\new_[26687]_ ;
  assign \new_[24596]_  = ~\new_[30206]_  & ~\new_[29401]_ ;
  assign \new_[24597]_  = (~\s11_data_i[23]  | ~\new_[29205]_ ) & (~\s8_data_i[23]  | ~\new_[29241]_ );
  assign \new_[24598]_  = ~\new_[28713]_  | ~\new_[5921]_ ;
  assign \new_[24599]_  = ~\new_[28110]_  & ~\new_[29854]_ ;
  assign \new_[24600]_  = ~\new_[28580]_  & (~\new_[30467]_  | ~\new_[6209]_ );
  assign \new_[24601]_  = ~\new_[28000]_  & ~\new_[30598]_ ;
  assign \new_[24602]_  = (~\new_[29710]_  | ~\s10_data_i[17] ) & (~\new_[29024]_  | ~\s9_data_i[17] );
  assign \new_[24603]_  = (~\new_[30227]_  | ~\s10_data_i[17] ) & (~\new_[29706]_  | ~\s9_data_i[17] );
  assign \new_[24604]_  = ~\new_[28154]_  & ~\new_[30445]_ ;
  assign \new_[24605]_  = ~\new_[28241]_  & ~\new_[30708]_ ;
  assign \new_[24606]_  = (~\s10_data_i[18]  | ~\new_[29749]_ ) & (~\s9_data_i[18]  | ~\new_[29034]_ );
  assign \new_[24607]_  = ~\new_[26867]_ ;
  assign \new_[24608]_  = (~\new_[30181]_  | ~\s14_data_i[27] ) & (~\new_[29640]_  | ~\s12_data_i[27] );
  assign \new_[24609]_  = ~\new_[30275]_  | ~\new_[28215]_ ;
  assign \new_[24610]_  = \new_[28596]_  & \new_[29180]_ ;
  assign \new_[24611]_  = (~\s11_data_i[21]  | ~\new_[29205]_ ) & (~\s8_data_i[21]  | ~\new_[29241]_ );
  assign \new_[24612]_  = ~\new_[30618]_  | ~\new_[28888]_ ;
  assign \new_[24613]_  = ~\new_[29869]_  | ~\new_[28609]_ ;
  assign \new_[24614]_  = (~\new_[30181]_  | ~\s14_data_i[28] ) & (~\new_[29640]_  | ~\s12_data_i[28] );
  assign \new_[24615]_  = ~\new_[27637]_ ;
  assign \new_[24616]_  = (~\new_[30311]_  | ~\s11_data_i[28] ) & (~\new_[29636]_  | ~\s8_data_i[28] );
  assign \new_[24617]_  = ~\new_[26707]_ ;
  assign \new_[24618]_  = (~\new_[29012]_  | ~\s10_data_i[22] ) & (~\new_[29185]_  | ~\s9_data_i[22] );
  assign \new_[24619]_  = ~\new_[29893]_  & ~\new_[28873]_ ;
  assign \new_[24620]_  = ~\new_[28227]_  | ~\new_[29118]_ ;
  assign \new_[24621]_  = \new_[28204]_  | \new_[28762]_ ;
  assign \new_[24622]_  = (~\s14_data_i[12]  | ~\new_[30026]_ ) & (~\s12_data_i[12]  | ~\new_[29711]_ );
  assign \new_[24623]_  = ~\new_[27085]_ ;
  assign \new_[24624]_  = ~\new_[30176]_  & ~\new_[6062]_ ;
  assign \new_[24625]_  = (~\new_[30311]_  | ~\s11_data_i[29] ) & (~\new_[29636]_  | ~\s8_data_i[29] );
  assign \new_[24626]_  = (~\new_[29045]_  | ~\s10_data_i[29] ) & (~\new_[29951]_  | ~\s9_data_i[29] );
  assign \new_[24627]_  = ~\new_[29825]_  & ~\new_[28052]_ ;
  assign \new_[24628]_  = ~\new_[26723]_ ;
  assign \new_[24629]_  = (~\new_[29628]_  | ~\s4_data_i[29] ) & (~\new_[29258]_  | ~\s0_data_i[29] );
  assign \new_[24630]_  = ~\new_[32135]_ ;
  assign \new_[24631]_  = ~\new_[29704]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[24632]_  = ~\new_[27630]_ ;
  assign \new_[24633]_  = \new_[30445]_  | \new_[28001]_ ;
  assign \new_[24634]_  = ~\new_[27251]_ ;
  assign \new_[24635]_  = ~\new_[5905]_  | ~\new_[30061]_  | ~\new_[29695]_ ;
  assign \new_[24636]_  = ~\new_[29817]_  | ~\new_[5929]_ ;
  assign \new_[24637]_  = (~\new_[29710]_  | ~\s10_data_i[31] ) & (~\new_[29024]_  | ~\s9_data_i[31] );
  assign \new_[24638]_  = (~\s4_data_i[12]  | ~\new_[30335]_ ) & (~\s0_data_i[12]  | ~\new_[29603]_ );
  assign \new_[24639]_  = (~\s11_data_i[27]  | ~\new_[29205]_ ) & (~\s8_data_i[27]  | ~\new_[29241]_ );
  assign \new_[24640]_  = ~\new_[28073]_  | ~\new_[5920]_ ;
  assign \new_[24641]_  = (~\new_[29953]_  | ~\s11_data_i[21] ) & (~\new_[29627]_  | ~\s8_data_i[21] );
  assign \new_[24642]_  = ~\new_[29197]_  & ~\new_[30331]_ ;
  assign \new_[24643]_  = (~\new_[28842]_  | ~\s4_data_i[1] ) & (~\new_[29434]_  | ~\s0_data_i[1] );
  assign \new_[24644]_  = ~\new_[26712]_ ;
  assign \new_[24645]_  = ~\new_[26739]_ ;
  assign \new_[24646]_  = ~\new_[29624]_  & (~\new_[29436]_  | ~\new_[29553]_ );
  assign \new_[24647]_  = ~\new_[28792]_  | ~\new_[6066]_ ;
  assign \new_[24648]_  = (~\new_[28842]_  | ~\s4_data_i[0] ) & (~\new_[29434]_  | ~\s0_data_i[0] );
  assign \new_[24649]_  = \new_[28150]_  & \new_[28275]_ ;
  assign \new_[24650]_  = (~\s11_data_i[18]  | ~\new_[29205]_ ) & (~\s8_data_i[18]  | ~\new_[29241]_ );
  assign \new_[24651]_  = (~\new_[29025]_  | ~\s5_data_i[1] ) & (~\new_[30469]_  | ~\s3_data_i[1] );
  assign \new_[24652]_  = ~\new_[28515]_  & (~\new_[30525]_  | ~\new_[6200]_ );
  assign \new_[24653]_  = \new_[28203]_  & \new_[31406]_ ;
  assign \new_[24654]_  = ~\new_[5901]_  | ~\new_[29404]_  | ~\new_[28828]_ ;
  assign \new_[24655]_  = (~\s11_data_i[1]  | ~\new_[29205]_ ) & (~\s8_data_i[1]  | ~\new_[29241]_ );
  assign \new_[24656]_  = ~\new_[30333]_  | ~\new_[28293]_ ;
  assign \new_[24657]_  = ~\new_[5896]_  | ~\new_[30320]_  | ~\new_[29320]_ ;
  assign \new_[24658]_  = (~\new_[30031]_  | ~\s7_data_i[10] ) & (~\new_[29052]_  | ~\s6_data_i[10] );
  assign \new_[24659]_  = (~\new_[30031]_  | ~\s7_data_i[1] ) & (~\new_[29052]_  | ~\s6_data_i[1] );
  assign \new_[24660]_  = ~\new_[28778]_  | ~\new_[31043]_ ;
  assign \new_[24661]_  = ~\new_[29573]_  & ~\new_[30092]_ ;
  assign \new_[24662]_  = ~\new_[29970]_  & ~\new_[28535]_ ;
  assign \new_[24663]_  = (~\new_[29705]_  | ~\s10_data_i[2] ) & (~\new_[30354]_  | ~\s9_data_i[2] );
  assign \new_[24664]_  = (~\new_[29705]_  | ~\s10_data_i[10] ) & (~\new_[30354]_  | ~\s9_data_i[10] );
  assign \new_[24665]_  = ~\new_[26733]_ ;
  assign \new_[24666]_  = (~\new_[30181]_  | ~\s14_data_i[15] ) & (~\new_[29640]_  | ~\s12_data_i[15] );
  assign \new_[24667]_  = ~\new_[28435]_  | ~\new_[30952]_ ;
  assign \new_[24668]_  = ~\new_[29276]_  & ~\new_[28020]_ ;
  assign \new_[24669]_  = (~\new_[30260]_  | ~\s11_data_i[26] ) & (~\new_[29670]_  | ~\s8_data_i[26] );
  assign \new_[24670]_  = \new_[28497]_  & \new_[28524]_ ;
  assign \new_[24671]_  = (~\new_[29534]_  | ~\s5_data_i[7] ) & (~\new_[29579]_  | ~\s3_data_i[7] );
  assign \new_[24672]_  = (~\new_[29628]_  | ~\s4_data_i[2] ) & (~\new_[29258]_  | ~\s0_data_i[2] );
  assign \new_[24673]_  = ~\new_[30348]_  & ~\new_[30066]_ ;
  assign \new_[24674]_  = ~\new_[28409]_  & ~\new_[29874]_ ;
  assign \new_[24675]_  = ~\new_[30337]_  | ~\new_[28397]_ ;
  assign \new_[24676]_  = (~\s14_data_i[2]  | ~\new_[30026]_ ) & (~\s12_data_i[2]  | ~\new_[29711]_ );
  assign \new_[24677]_  = ~\new_[29020]_  & ~\new_[30266]_ ;
  assign \new_[24678]_  = (~\s14_data_i[19]  | ~\new_[30026]_ ) & (~\s12_data_i[19]  | ~\new_[29711]_ );
  assign \new_[24679]_  = (~\new_[29641]_  | ~\s14_data_i[1] ) & (~\new_[29317]_  | ~\s12_data_i[1] );
  assign \new_[24680]_  = (~\new_[29710]_  | ~\s10_data_i[10] ) & (~\new_[29024]_  | ~\s9_data_i[10] );
  assign \new_[24681]_  = (~\new_[30031]_  | ~\s7_data_i[28] ) & (~\new_[29052]_  | ~\s6_data_i[28] );
  assign \new_[24682]_  = ~\new_[6036]_  | ~\new_[28650]_  | ~\new_[29841]_ ;
  assign \new_[24683]_  = ~\new_[26673]_ ;
  assign \new_[24684]_  = ~\new_[27610]_ ;
  assign \new_[24685]_  = ~\new_[28400]_  & (~\new_[30653]_  | ~\new_[6194]_ );
  assign \new_[24686]_  = (~\new_[30227]_  | ~\s10_data_i[18] ) & (~\new_[29706]_  | ~\s9_data_i[18] );
  assign \new_[24687]_  = ~\new_[6072]_  | ~\new_[30321]_  | ~\new_[30775]_ ;
  assign \new_[24688]_  = ~\new_[30837]_  | ~\new_[28762]_ ;
  assign \new_[24689]_  = \new_[28509]_  | \new_[30003]_ ;
  assign \new_[24690]_  = ~\new_[27167]_ ;
  assign \new_[24691]_  = ~\new_[28462]_  & (~\new_[30499]_  | ~\new_[6049]_ );
  assign \new_[24692]_  = ~\new_[26782]_ ;
  assign \new_[24693]_  = ~\new_[26765]_ ;
  assign \new_[24694]_  = ~\new_[27777]_ ;
  assign \new_[24695]_  = (~\new_[30200]_  | ~\s11_data_i[27] ) & (~\new_[29428]_  | ~\s8_data_i[27] );
  assign \new_[24696]_  = (~\new_[29953]_  | ~\s11_data_i[2] ) & (~\new_[29627]_  | ~\s8_data_i[2] );
  assign \new_[24697]_  = ~\new_[26785]_ ;
  assign n8294 = ~\new_[29697]_  | ~\new_[28349]_ ;
  assign \new_[24699]_  = ~\new_[26788]_ ;
  assign \new_[24700]_  = \new_[28405]_  | \new_[29508]_ ;
  assign \new_[24701]_  = (~\new_[30260]_  | ~\s11_data_i[16] ) & (~\new_[29670]_  | ~\s8_data_i[16] );
  assign \new_[24702]_  = (~\new_[29534]_  | ~\s5_data_i[13] ) & (~\new_[29579]_  | ~\s3_data_i[13] );
  assign \new_[24703]_  = (~\new_[30193]_  | ~\s7_data_i[0] ) & (~\new_[29298]_  | ~\s6_data_i[0] );
  assign \new_[24704]_  = ~\new_[30138]_  & ~\new_[28052]_ ;
  assign \new_[24705]_  = ~\new_[27604]_ ;
  assign \new_[24706]_  = (~\new_[28842]_  | ~\s4_data_i[23] ) & (~\new_[29434]_  | ~\s0_data_i[23] );
  assign \new_[24707]_  = (~\s11_data_i[9]  | ~\new_[29205]_ ) & (~\s8_data_i[9]  | ~\new_[29241]_ );
  assign \new_[24708]_  = (~\new_[29976]_  | ~\s14_data_i[4] ) & (~\new_[28957]_  | ~\s12_data_i[4] );
  assign \new_[24709]_  = ~\new_[30019]_  | ~\new_[29748]_ ;
  assign \new_[24710]_  = ~\new_[29855]_  & ~\new_[30097]_ ;
  assign \new_[24711]_  = (~\s2_data_i[2]  | ~\new_[29625]_ ) & (~\s1_data_i[2]  | ~\new_[29215]_ );
  assign \new_[24712]_  = ~\new_[29771]_  & ~\new_[29122]_ ;
  assign \new_[24713]_  = (~\new_[29628]_  | ~\s4_data_i[10] ) & (~\new_[29258]_  | ~\s0_data_i[10] );
  assign \new_[24714]_  = (~\s4_data_i[19]  | ~\new_[30335]_ ) & (~\s0_data_i[19]  | ~\new_[29603]_ );
  assign \new_[24715]_  = (~\new_[29012]_  | ~\s10_data_i[3] ) & (~\new_[29185]_  | ~\s9_data_i[3] );
  assign \new_[24716]_  = ~\new_[28182]_  | ~\new_[28412]_ ;
  assign \new_[24717]_  = (~\new_[29710]_  | ~\s10_data_i[29] ) & (~\new_[29024]_  | ~\s9_data_i[29] );
  assign \new_[24718]_  = ~\new_[5909]_  | ~\new_[28650]_  | ~\new_[29841]_ ;
  assign \new_[24719]_  = (~\new_[28842]_  | ~\s4_data_i[15] ) & (~\new_[29434]_  | ~\s0_data_i[15] );
  assign \new_[24720]_  = ~\new_[27597]_ ;
  assign \new_[24721]_  = ~\new_[30633]_  & ~\new_[29815]_ ;
  assign \new_[24722]_  = ~\new_[26804]_ ;
  assign \new_[24723]_  = (~\new_[29976]_  | ~\s14_data_i[10] ) & (~\new_[28957]_  | ~\s12_data_i[10] );
  assign \new_[24724]_  = \new_[28428]_  & \new_[30150]_ ;
  assign \new_[24725]_  = ~\new_[26988]_ ;
  assign \new_[24726]_  = \new_[28074]_  | \new_[29676]_ ;
  assign \new_[24727]_  = (~\new_[29953]_  | ~\s11_data_i[4] ) & (~\new_[29627]_  | ~\s8_data_i[4] );
  assign \new_[24728]_  = (~\s5_data_i[5]  | ~\new_[29649]_ ) & (~\s3_data_i[5]  | ~\new_[29035]_ );
  assign \new_[24729]_  = (~\new_[30031]_  | ~\s7_data_i[24] ) & (~\new_[29052]_  | ~\s6_data_i[24] );
  assign \new_[24730]_  = ~\new_[30649]_  | ~\new_[6050]_ ;
  assign \new_[24731]_  = (~\new_[30311]_  | ~\s11_data_i[8] ) & (~\new_[29636]_  | ~\s8_data_i[8] );
  assign \new_[24732]_  = ~\new_[26987]_ ;
  assign \new_[24733]_  = (~\new_[29534]_  | ~\s5_data_i[20] ) & (~\new_[29579]_  | ~\s3_data_i[20] );
  assign \new_[24734]_  = (~\new_[29021]_  | ~\s10_data_i[21] ) & (~\new_[29709]_  | ~\s9_data_i[21] );
  assign \new_[24735]_  = (~\new_[29036]_  | ~\s5_data_i[17] ) & (~\new_[30429]_  | ~\s3_data_i[17] );
  assign \new_[24736]_  = (~\s5_data_i[2]  | ~\new_[29649]_ ) & (~\s3_data_i[2]  | ~\new_[29035]_ );
  assign \new_[24737]_  = ~\new_[28118]_  | ~\new_[28850]_ ;
  assign \new_[24738]_  = ~\new_[28286]_  | ~\new_[28371]_ ;
  assign \new_[24739]_  = \new_[28201]_  & \new_[30025]_ ;
  assign \new_[24740]_  = ~\new_[26757]_ ;
  assign \new_[24741]_  = ~\new_[26756]_ ;
  assign \new_[24742]_  = ~\new_[28011]_  | ~\new_[31045]_ ;
  assign \new_[24743]_  = ~\new_[28369]_  | ~\new_[30432]_ ;
  assign \new_[24744]_  = ~\new_[26750]_ ;
  assign \new_[24745]_  = ~\new_[27766]_ ;
  assign \new_[24746]_  = ~\new_[29987]_  | ~\new_[30210]_ ;
  assign \new_[24747]_  = (~\new_[29025]_  | ~\s5_data_i[6] ) & (~\new_[30469]_  | ~\s3_data_i[6] );
  assign \new_[24748]_  = ~\new_[30350]_  & ~\new_[30010]_ ;
  assign \new_[24749]_  = \new_[27986]_  & \new_[30554]_ ;
  assign \new_[24750]_  = (~\new_[29628]_  | ~\s4_data_i[9] ) & (~\new_[29258]_  | ~\s0_data_i[9] );
  assign \new_[24751]_  = ~\new_[29943]_  | ~\new_[28979]_ ;
  assign \new_[24752]_  = ~\new_[28840]_  & ~\new_[28232]_ ;
  assign \new_[24753]_  = (~\s2_data_i[9]  | ~\new_[29625]_ ) & (~\s1_data_i[9]  | ~\new_[29215]_ );
  assign \new_[24754]_  = ~\new_[28682]_  & ~\new_[29887]_ ;
  assign \new_[24755]_  = (~\new_[29705]_  | ~\s10_data_i[6] ) & (~\new_[30354]_  | ~\s9_data_i[6] );
  assign \new_[24756]_  = ~\new_[26833]_ ;
  assign \new_[24757]_  = (~\s11_data_i[13]  | ~\new_[29205]_ ) & (~\s8_data_i[13]  | ~\new_[29241]_ );
  assign \new_[24758]_  = ~\new_[30145]_  & ~\new_[30152]_ ;
  assign \new_[24759]_  = ~\new_[29299]_ ;
  assign \new_[24760]_  = ~\new_[30236]_  & ~\new_[29032]_ ;
  assign \new_[24761]_  = ~\new_[27753]_ ;
  assign \new_[24762]_  = (~\s4_data_i[0]  | ~\new_[30335]_ ) & (~\s0_data_i[0]  | ~\new_[29603]_ );
  assign \new_[24763]_  = \new_[28429]_  & \new_[28663]_ ;
  assign \new_[24764]_  = ~\new_[30607]_  & ~\new_[30003]_ ;
  assign \new_[24765]_  = (~\new_[28842]_  | ~\s4_data_i[6] ) & (~\new_[29434]_  | ~\s0_data_i[6] );
  assign \new_[24766]_  = ~\new_[27622]_ ;
  assign \new_[24767]_  = (~\new_[29953]_  | ~\s11_data_i[8] ) & (~\new_[29627]_  | ~\s8_data_i[8] );
  assign \new_[24768]_  = ~\new_[26847]_ ;
  assign \new_[24769]_  = (~\s2_data_i[20]  | ~\new_[29625]_ ) & (~\s1_data_i[20]  | ~\new_[29215]_ );
  assign \new_[24770]_  = ~\new_[27748]_ ;
  assign \new_[24771]_  = ~\new_[28899]_  & ~\new_[29762]_ ;
  assign \new_[24772]_  = (~\s2_data_i[1]  | ~\new_[29625]_ ) & (~\s1_data_i[1]  | ~\new_[29215]_ );
  assign \new_[24773]_  = (~\new_[30193]_  | ~\s7_data_i[13] ) & (~\new_[29298]_  | ~\s6_data_i[13] );
  assign \new_[24774]_  = ~\new_[30164]_  | ~\new_[28114]_ ;
  assign \new_[24775]_  = (~\new_[29976]_  | ~\s14_data_i[7] ) & (~\new_[28957]_  | ~\s12_data_i[7] );
  assign \new_[24776]_  = ~\new_[29768]_  & ~\new_[29956]_ ;
  assign \new_[24777]_  = ~\new_[30038]_  & (~\new_[29244]_  | ~\new_[29351]_ );
  assign \new_[24778]_  = ~\new_[27558]_ ;
  assign \new_[24779]_  = (~\new_[29025]_  | ~\s5_data_i[0] ) & (~\new_[30469]_  | ~\s3_data_i[0] );
  assign \new_[24780]_  = ~\new_[27557]_ ;
  assign n8299 = ~\new_[28861]_  | ~\new_[28107]_ ;
  assign \new_[24782]_  = ~\new_[30068]_  & ~\new_[27892]_ ;
  assign \new_[24783]_  = ~\new_[29100]_  & ~\new_[30320]_ ;
  assign n8289 = ~\new_[29002]_  | ~\new_[28350]_ ;
  assign \new_[24785]_  = ~\new_[30043]_  & ~\new_[30267]_ ;
  assign n8279 = ~\new_[29702]_  | ~\new_[28351]_ ;
  assign \new_[24787]_  = ~\new_[28718]_  & ~\new_[29397]_ ;
  assign \new_[24788]_  = ~\new_[30217]_  | ~\new_[29831]_ ;
  assign n8284 = ~\new_[29369]_  | ~\new_[28080]_ ;
  assign \new_[24790]_  = \new_[28469]_  | \new_[29853]_ ;
  assign \new_[24791]_  = (~\new_[30031]_  | ~\s7_data_i[7] ) & (~\new_[29052]_  | ~\s6_data_i[7] );
  assign \new_[24792]_  = ~\new_[26860]_ ;
  assign \new_[24793]_  = (~\new_[28842]_  | ~\s4_data_i[7] ) & (~\new_[29434]_  | ~\s0_data_i[7] );
  assign \new_[24794]_  = \new_[28301]_  & \new_[30150]_ ;
  assign \new_[24795]_  = ~\new_[28545]_  | ~\new_[29900]_ ;
  assign \new_[24796]_  = \new_[28644]_  | \new_[30612]_ ;
  assign \new_[24797]_  = \new_[28555]_  | \new_[30566]_ ;
  assign \new_[24798]_  = ~\new_[28460]_  & ~\new_[30230]_ ;
  assign \new_[24799]_  = ~\new_[5932]_  | ~\new_[28371]_  | ~\new_[30021]_ ;
  assign \new_[24800]_  = \new_[28465]_  | \new_[28503]_ ;
  assign \new_[24801]_  = (~\new_[29953]_  | ~\s11_data_i[10] ) & (~\new_[29627]_  | ~\s8_data_i[10] );
  assign \new_[24802]_  = ~\new_[28201]_  | ~\new_[30021]_ ;
  assign \new_[24803]_  = ~\new_[28451]_  & ~\new_[30199]_ ;
  assign \new_[24804]_  = ~\new_[5964]_  | ~\new_[28845]_  | ~\new_[29874]_ ;
  assign \new_[24805]_  = \new_[28527]_  | \new_[29784]_ ;
  assign \new_[24806]_  = ~\new_[28269]_  | ~\new_[29874]_ ;
  assign \new_[24807]_  = ~\new_[28162]_  | ~\new_[30164]_ ;
  assign \new_[24808]_  = ~\new_[27987]_  | ~\new_[28114]_ ;
  assign \new_[24809]_  = ~\new_[28483]_  & ~\new_[29906]_ ;
  assign \new_[24810]_  = ~\new_[26878]_ ;
  assign \new_[24811]_  = ~\new_[28589]_  | ~\new_[29504]_ ;
  assign \new_[24812]_  = ~\new_[26675]_ ;
  assign \new_[24813]_  = ~\new_[28385]_  | ~\new_[30020]_ ;
  assign \new_[24814]_  = ~\new_[28495]_  | ~\new_[30296]_ ;
  assign \new_[24815]_  = ~\new_[28389]_  | ~\new_[28069]_ ;
  assign \new_[24816]_  = ~\new_[26676]_ ;
  assign \new_[24817]_  = ~\new_[26881]_ ;
  assign \new_[24818]_  = \new_[29344]_  & \new_[30499]_ ;
  assign \new_[24819]_  = \new_[29461]_  & \new_[30653]_ ;
  assign \new_[24820]_  = ~\new_[28182]_  & ~\new_[29855]_ ;
  assign \new_[24821]_  = ~\new_[28352]_  & ~\new_[28113]_ ;
  assign \new_[24822]_  = ~\new_[27978]_  | ~\new_[29260]_ ;
  assign \new_[24823]_  = ~\new_[28115]_  & ~\new_[30287]_ ;
  assign \new_[24824]_  = \new_[28532]_  | \new_[30663]_ ;
  assign \new_[24825]_  = ~\new_[26887]_ ;
  assign \new_[24826]_  = \new_[28394]_  | \new_[28397]_ ;
  assign \new_[24827]_  = \new_[28485]_  | \new_[30342]_ ;
  assign \new_[24828]_  = ~\new_[6038]_  | ~\new_[29079]_  | ~\new_[29220]_ ;
  assign \new_[24829]_  = ~\new_[28526]_  | ~\new_[30215]_ ;
  assign \new_[24830]_  = \new_[28591]_  & \new_[29412]_ ;
  assign \new_[24831]_  = ~\new_[28727]_  | ~\new_[30215]_ ;
  assign \new_[24832]_  = ~\new_[28473]_  | ~\new_[29220]_ ;
  assign \new_[24833]_  = \new_[28399]_  & \new_[29003]_ ;
  assign \new_[24834]_  = (~\s11_data_i[20]  | ~\new_[29205]_ ) & (~\s8_data_i[20]  | ~\new_[29241]_ );
  assign \new_[24835]_  = ~\new_[28259]_  & ~\new_[29743]_ ;
  assign \new_[24836]_  = \new_[28176]_  | \new_[30656]_ ;
  assign \new_[24837]_  = ~\new_[28219]_  | ~\new_[29411]_ ;
  assign \new_[24838]_  = ~\new_[29108]_  | ~\new_[28390]_ ;
  assign \new_[24839]_  = ~\new_[28704]_  & ~\new_[29100]_ ;
  assign \new_[24840]_  = \new_[28803]_  & \new_[29320]_ ;
  assign \new_[24841]_  = \new_[28803]_  | \new_[28329]_ ;
  assign \new_[24842]_  = \new_[28525]_  | \new_[30575]_ ;
  assign \new_[24843]_  = \new_[28722]_  | \new_[30747]_ ;
  assign \new_[24844]_  = ~\new_[28208]_  | ~\new_[30125]_ ;
  assign \new_[24845]_  = \new_[28733]_  & \new_[30842]_ ;
  assign \new_[24846]_  = ~\new_[28468]_  & ~\new_[30047]_ ;
  assign \new_[24847]_  = (~\s2_data_i[16]  | ~\new_[29625]_ ) & (~\s1_data_i[16]  | ~\new_[29215]_ );
  assign \new_[24848]_  = \new_[29444]_  & \new_[29746]_ ;
  assign \new_[24849]_  = \new_[28368]_  | \new_[30607]_ ;
  assign \new_[24850]_  = \new_[29480]_  & \new_[30572]_ ;
  assign \new_[24851]_  = ~\new_[28377]_  | ~\new_[29518]_ ;
  assign \new_[24852]_  = ~\new_[29848]_  & ~\new_[28989]_ ;
  assign \new_[24853]_  = ~\new_[28180]_  | ~\new_[29260]_ ;
  assign \new_[24854]_  = ~\new_[26581]_ ;
  assign \new_[24855]_  = \new_[28180]_  & \new_[28866]_ ;
  assign \new_[24856]_  = (~\s14_data_i[3]  | ~\new_[30026]_ ) & (~\s12_data_i[3]  | ~\new_[29711]_ );
  assign \new_[24857]_  = ~\new_[28519]_  & ~\new_[29199]_ ;
  assign \new_[24858]_  = ~\new_[28308]_  | ~\new_[30139]_ ;
  assign \new_[24859]_  = \new_[29454]_  | \new_[30289]_ ;
  assign \new_[24860]_  = ~\new_[26897]_ ;
  assign \new_[24861]_  = ~\new_[27537]_ ;
  assign \new_[24862]_  = \new_[28566]_  & \new_[30037]_ ;
  assign \new_[24863]_  = \new_[28130]_  | \new_[30289]_ ;
  assign \new_[24864]_  = \new_[28531]_  & \new_[29228]_ ;
  assign \new_[24865]_  = (~\new_[29976]_  | ~\s14_data_i[8] ) & (~\new_[28957]_  | ~\s12_data_i[8] );
  assign \new_[24866]_  = \new_[28551]_  | \new_[30769]_ ;
  assign \new_[24867]_  = \new_[28210]_  | \new_[28317]_ ;
  assign \new_[24868]_  = ~\new_[30293]_  | ~\new_[30617]_ ;
  assign \new_[24869]_  = \new_[28576]_  & \new_[30505]_ ;
  assign \new_[24870]_  = \new_[28597]_  & \new_[29462]_ ;
  assign \new_[24871]_  = \new_[28531]_  | \new_[28147]_ ;
  assign \new_[24872]_  = \new_[28634]_  | \new_[30342]_ ;
  assign \new_[24873]_  = ~\new_[6064]_  | ~\new_[30083]_  | ~\new_[30636]_ ;
  assign \new_[24874]_  = ~\new_[28403]_  | ~\new_[29524]_ ;
  assign \new_[24875]_  = ~\new_[6206]_  | ~\new_[29783]_  | ~\new_[30255]_ ;
  assign \new_[24876]_  = ~\new_[29761]_  | ~\new_[29783]_ ;
  assign \new_[24877]_  = \new_[28218]_  | \new_[30757]_ ;
  assign \new_[24878]_  = \new_[28147]_  & \new_[29228]_ ;
  assign \new_[24879]_  = ~\new_[28160]_  & ~\new_[29315]_ ;
  assign \new_[24880]_  = ~\new_[28489]_  | ~\new_[30255]_ ;
  assign \new_[24881]_  = ~\new_[28137]_  & ~\new_[30389]_ ;
  assign \new_[24882]_  = \new_[28788]_  & \new_[30446]_ ;
  assign \new_[24883]_  = ~\new_[26906]_ ;
  assign \new_[24884]_  = ~\new_[6001]_  | ~\new_[29886]_  | ~\new_[29386]_ ;
  assign \new_[24885]_  = ~\new_[28544]_  & ~\new_[28899]_ ;
  assign \new_[24886]_  = ~\new_[27882]_ ;
  assign \new_[24887]_  = ~\new_[26910]_ ;
  assign \new_[24888]_  = ~\new_[28585]_  & ~\new_[30598]_ ;
  assign \new_[24889]_  = \new_[28231]_  | \new_[30616]_ ;
  assign \new_[24890]_  = ~\new_[27863]_ ;
  assign \new_[24891]_  = \new_[28225]_  | \new_[30389]_ ;
  assign \new_[24892]_  = ~\new_[28150]_  & ~\new_[30564]_ ;
  assign \new_[24893]_  = ~\new_[28598]_  | ~\new_[28023]_ ;
  assign \new_[24894]_  = \new_[28445]_  | \new_[30616]_ ;
  assign \new_[24895]_  = ~\new_[28431]_  & ~\new_[30305]_ ;
  assign \new_[24896]_  = \new_[28459]_  | \new_[29935]_ ;
  assign \new_[24897]_  = \new_[28632]_  | \new_[29272]_ ;
  assign \new_[24898]_  = \new_[28518]_  & \new_[29608]_ ;
  assign \new_[24899]_  = ~\new_[28560]_  & ~\new_[28020]_ ;
  assign \new_[24900]_  = \new_[28442]_  | \new_[30348]_ ;
  assign \new_[24901]_  = ~\new_[6031]_  | ~\new_[29782]_  | ~\new_[30774]_ ;
  assign \new_[24902]_  = ~\new_[28799]_  | ~\new_[29782]_ ;
  assign \new_[24903]_  = \new_[29294]_  & \new_[30678]_ ;
  assign \new_[24904]_  = \new_[29413]_  | \new_[30162]_ ;
  assign \new_[24905]_  = \new_[28570]_  | \new_[29576]_ ;
  assign \new_[24906]_  = \new_[29351]_  & \new_[30697]_ ;
  assign \new_[24907]_  = ~\new_[26920]_ ;
  assign \new_[24908]_  = ~\new_[26939]_ ;
  assign \new_[24909]_  = \new_[28138]_  | \new_[29902]_ ;
  assign \new_[24910]_  = ~\new_[28772]_  & ~\new_[30185]_ ;
  assign \new_[24911]_  = \new_[28116]_  | \new_[30407]_ ;
  assign \new_[24912]_  = \new_[28496]_  | \new_[28846]_ ;
  assign \new_[24913]_  = \new_[29531]_  & \new_[29299]_ ;
  assign \new_[24914]_  = ~\new_[28432]_  & ~\new_[30339]_ ;
  assign \new_[24915]_  = ~\new_[27172]_ ;
  assign \new_[24916]_  = \new_[28498]_  | \new_[28846]_ ;
  assign \new_[24917]_  = \new_[28511]_  | \new_[28402]_ ;
  assign \new_[24918]_  = ~\new_[6190]_  | ~\new_[29225]_  | ~\new_[30125]_ ;
  assign \new_[24919]_  = ~\new_[28708]_  & ~\new_[29916]_ ;
  assign \new_[24920]_  = ~\new_[28481]_  & ~\new_[30174]_ ;
  assign \new_[24921]_  = ~\new_[31491]_  | ~\new_[30207]_  | ~\new_[30617]_ ;
  assign \new_[24922]_  = \new_[28144]_  | \new_[30224]_ ;
  assign \new_[24923]_  = ~\new_[27775]_ ;
  assign \new_[24924]_  = ~\new_[28213]_  | ~\new_[29392]_ ;
  assign \new_[24925]_  = ~\new_[28370]_  & ~\new_[30167]_ ;
  assign \new_[24926]_  = \new_[29183]_  & \new_[30000]_ ;
  assign \new_[24927]_  = \new_[28378]_  | \new_[30289]_ ;
  assign \new_[24928]_  = ~\new_[28437]_  & ~\new_[30219]_ ;
  assign \new_[24929]_  = ~\new_[30233]_  | ~\new_[29996]_ ;
  assign \new_[24930]_  = ~\new_[28621]_  | ~\new_[29904]_ ;
  assign \new_[24931]_  = \new_[28359]_  | \new_[30684]_ ;
  assign \new_[24932]_  = ~\new_[28164]_  & ~\new_[30515]_ ;
  assign \new_[24933]_  = \new_[28802]_  | \new_[30675]_ ;
  assign \new_[24934]_  = \new_[28540]_  | \new_[30273]_ ;
  assign \new_[24935]_  = ~\new_[5930]_  | ~\new_[29927]_  | ~\new_[30507]_ ;
  assign \new_[24936]_  = ~\new_[28451]_  & ~\new_[30675]_ ;
  assign \new_[24937]_  = \new_[28341]_  & \new_[29870]_ ;
  assign \new_[24938]_  = ~\new_[31491]_  | ~\new_[30617]_  | ~\new_[30434]_ ;
  assign \new_[24939]_  = ~\new_[5979]_  | ~\new_[30344]_  | ~\new_[28870]_ ;
  assign \new_[24940]_  = \new_[29558]_  | \new_[30014]_ ;
  assign \new_[24941]_  = ~\new_[28381]_  | ~\new_[28870]_ ;
  assign \new_[24942]_  = ~\new_[28274]_  | ~\new_[29221]_ ;
  assign \new_[24943]_  = ~\new_[6204]_  | ~\new_[30139]_  | ~\new_[30665]_ ;
  assign \new_[24944]_  = \new_[28543]_  & \new_[29271]_ ;
  assign \new_[24945]_  = \new_[27987]_  & \new_[29550]_ ;
  assign \new_[24946]_  = ~\new_[29506]_  | ~\new_[28930]_ ;
  assign \new_[24947]_  = ~\new_[28707]_  | ~\new_[30615]_ ;
  assign \new_[24948]_  = ~\new_[28287]_  | ~\new_[29967]_ ;
  assign \new_[24949]_  = ~\new_[28217]_  | ~\new_[29015]_ ;
  assign \new_[24950]_  = ~\new_[28446]_  & ~\new_[30087]_ ;
  assign \new_[24951]_  = \new_[28570]_  & \new_[28786]_ ;
  assign \new_[24952]_  = ~\new_[28382]_  & ~\new_[30087]_ ;
  assign \new_[24953]_  = ~\new_[28090]_  & ~\new_[28362]_ ;
  assign \new_[24954]_  = \new_[28416]_  | \new_[30028]_ ;
  assign \new_[24955]_  = ~\new_[28668]_  | ~\new_[30723]_ ;
  assign \new_[24956]_  = ~\new_[26931]_ ;
  assign \new_[24957]_  = ~\new_[28592]_  | ~\new_[29105]_ ;
  assign \new_[24958]_  = ~\new_[28472]_  | ~\new_[30083]_ ;
  assign \new_[24959]_  = ~\new_[26929]_ ;
  assign \new_[24960]_  = ~\new_[30325]_  & ~\new_[29798]_ ;
  assign \new_[24961]_  = ~\new_[28548]_  | ~\new_[28967]_ ;
  assign \new_[24962]_  = \new_[28185]_  | \new_[30028]_ ;
  assign \new_[24963]_  = ~\new_[28460]_  & ~\new_[30612]_ ;
  assign \new_[24964]_  = ~\new_[28336]_  & ~\new_[29573]_ ;
  assign \new_[24965]_  = ~\new_[27392]_ ;
  assign \new_[24966]_  = ~\new_[28556]_  & ~\new_[30423]_ ;
  assign \new_[24967]_  = ~\new_[27530]_ ;
  assign \new_[24968]_  = \new_[28743]_  | \new_[30696]_ ;
  assign \new_[24969]_  = \new_[28558]_  | \new_[28467]_ ;
  assign \new_[24970]_  = \new_[28582]_  & \new_[29817]_ ;
  assign \new_[24971]_  = \new_[28457]_  | \new_[30350]_ ;
  assign \new_[24972]_  = ~\new_[27976]_  | ~\new_[30432]_ ;
  assign \new_[24973]_  = ~\new_[28216]_  | ~\new_[30158]_ ;
  assign \new_[24974]_  = ~\new_[27437]_ ;
  assign \new_[24975]_  = ~\new_[6190]_  | ~\new_[29656]_  | ~\new_[29225]_ ;
  assign \new_[24976]_  = ~\new_[28497]_  & ~\new_[30651]_ ;
  assign \new_[24977]_  = \new_[28549]_  & \new_[28930]_ ;
  assign \new_[24978]_  = ~\new_[6212]_  | ~\new_[29891]_  | ~\new_[30595]_ ;
  assign \new_[24979]_  = \new_[29499]_  | \new_[30014]_ ;
  assign \new_[24980]_  = \new_[29469]_  | \new_[30014]_ ;
  assign \new_[24981]_  = \new_[28584]_  & \new_[29456]_ ;
  assign \new_[24982]_  = ~\new_[27488]_ ;
  assign \new_[24983]_  = ~\new_[28794]_  | ~\new_[30595]_ ;
  assign \new_[24984]_  = \new_[28584]_  | \new_[28339]_ ;
  assign \new_[24985]_  = \new_[28458]_  | \new_[30633]_ ;
  assign \new_[24986]_  = ~\new_[28196]_  & ~\new_[30254]_ ;
  assign \new_[24987]_  = \new_[28433]_  | \new_[29767]_ ;
  assign \new_[24988]_  = ~\new_[28440]_  & ~\new_[30478]_ ;
  assign \new_[24989]_  = ~\new_[28302]_  & ~\new_[29767]_ ;
  assign \new_[24990]_  = \new_[28604]_  | \new_[30780]_ ;
  assign \new_[24991]_  = ~\new_[28440]_  & ~\new_[30254]_ ;
  assign \new_[24992]_  = \new_[28441]_  & \new_[29975]_ ;
  assign \new_[24993]_  = ~\new_[27289]_ ;
  assign \new_[24994]_  = \new_[28465]_  & \new_[30283]_ ;
  assign \new_[24995]_  = \new_[28533]_  | \new_[30116]_ ;
  assign \new_[24996]_  = ~\new_[28550]_  & ~\new_[30651]_ ;
  assign \new_[24997]_  = ~\new_[28703]_  | ~\new_[30600]_ ;
  assign \new_[24998]_  = ~\new_[27431]_ ;
  assign \new_[24999]_  = ~\new_[28122]_  & ~\new_[30063]_ ;
  assign \new_[25000]_  = \new_[28340]_  & \new_[29006]_ ;
  assign \new_[25001]_  = ~\new_[28414]_  & ~\new_[30051]_ ;
  assign \new_[25002]_  = (~\s5_data_i[20]  | ~\new_[29649]_ ) & (~\s3_data_i[20]  | ~\new_[29035]_ );
  assign \new_[25003]_  = \new_[28139]_  | \new_[30837]_ ;
  assign \new_[25004]_  = \new_[28512]_  | \new_[29989]_ ;
  assign \new_[25005]_  = \new_[28562]_  | \new_[29540]_ ;
  assign \new_[25006]_  = ~\new_[30381]_  & ~\new_[30212]_ ;
  assign \new_[25007]_  = ~\new_[28376]_  | ~\new_[29656]_ ;
  assign \new_[25008]_  = ~\new_[28363]_  & ~\new_[30058]_ ;
  assign \new_[25009]_  = ~\new_[28079]_  & ~\new_[30415]_ ;
  assign \new_[25010]_  = \new_[28208]_  & \new_[29656]_ ;
  assign \new_[25011]_  = ~\new_[28800]_  | ~\new_[30789]_ ;
  assign \new_[25012]_  = \new_[28598]_  & \new_[29787]_ ;
  assign \new_[25013]_  = ~\new_[26948]_ ;
  assign \new_[25014]_  = \new_[28563]_  | \new_[30240]_ ;
  assign \new_[25015]_  = \new_[28436]_  | \new_[30755]_ ;
  assign \new_[25016]_  = ~\new_[28813]_  | ~\new_[29891]_ ;
  assign \new_[25017]_  = \new_[28329]_  & \new_[29320]_ ;
  assign \new_[25018]_  = \new_[28444]_  | \new_[30176]_ ;
  assign \new_[25019]_  = \new_[28453]_  | \new_[29565]_ ;
  assign \new_[25020]_  = ~\new_[28749]_  & ~\new_[30059]_ ;
  assign \new_[25021]_  = ~\new_[28798]_  & ~\new_[30569]_ ;
  assign \new_[25022]_  = \new_[28447]_  | \new_[29745]_ ;
  assign \new_[25023]_  = \new_[28184]_  | \new_[29100]_ ;
  assign \new_[25024]_  = ~\new_[26947]_ ;
  assign \new_[25025]_  = \new_[28784]_  & \new_[29979]_ ;
  assign \new_[25026]_  = \new_[27994]_  & \new_[29802]_ ;
  assign \new_[25027]_  = \new_[28220]_  & \new_[29787]_ ;
  assign \new_[25028]_  = ~\new_[28439]_  & ~\new_[30557]_ ;
  assign \new_[25029]_  = ~\new_[28383]_  | ~\new_[28926]_ ;
  assign \new_[25030]_  = \new_[28328]_  & \new_[29571]_ ;
  assign \new_[25031]_  = ~\new_[28811]_  & ~\new_[29648]_ ;
  assign \new_[25032]_  = (~\new_[29021]_  | ~\s10_data_i[7] ) & (~\new_[29709]_  | ~\s9_data_i[7] );
  assign \new_[25033]_  = (~\new_[30284]_  | ~\s11_data_i[15] ) & (~\new_[29420]_  | ~\s8_data_i[15] );
  assign \new_[25034]_  = ~\new_[28491]_  | ~\new_[30138]_ ;
  assign \new_[25035]_  = ~\new_[5996]_  | ~\new_[30702]_  | ~\new_[30610]_ ;
  assign \new_[25036]_  = \new_[28429]_  | \new_[29606]_ ;
  assign \new_[25037]_  = \new_[28177]_  | \new_[29648]_ ;
  assign \new_[25038]_  = \new_[28466]_  | \new_[30032]_ ;
  assign \new_[25039]_  = \new_[28464]_  | \new_[29944]_ ;
  assign \new_[25040]_  = ~\new_[28297]_  & ~\new_[30309]_ ;
  assign \new_[25041]_  = \new_[28230]_  | \new_[30501]_ ;
  assign \new_[25042]_  = \new_[28477]_  | \new_[30682]_ ;
  assign \new_[25043]_  = \new_[29489]_  & \new_[30691]_ ;
  assign \new_[25044]_  = ~\new_[28461]_  & ~\new_[30682]_ ;
  assign \new_[25045]_  = \new_[28174]_  | \new_[30620]_ ;
  assign \new_[25046]_  = ~\new_[30022]_  | ~\new_[6052]_ ;
  assign \new_[25047]_  = \new_[28523]_  | \new_[30400]_ ;
  assign \new_[25048]_  = ~\new_[28733]_  | ~\new_[30491]_ ;
  assign \new_[25049]_  = ~\new_[6269]_  | ~\new_[29913]_  | ~\new_[29210]_ ;
  assign \new_[25050]_  = \new_[28838]_  | \new_[30244]_ ;
  assign \new_[25051]_  = \new_[28529]_  | \new_[29238]_ ;
  assign \new_[25052]_  = \new_[28567]_  | \new_[30244]_ ;
  assign \new_[25053]_  = \new_[28471]_  & \new_[30205]_ ;
  assign \new_[25054]_  = \new_[29572]_  & \new_[29251]_ ;
  assign \new_[25055]_  = \new_[28539]_  & \new_[30205]_ ;
  assign \new_[25056]_  = \new_[28372]_  | \new_[29898]_ ;
  assign \new_[25057]_  = \new_[28339]_  & \new_[29456]_ ;
  assign \new_[25058]_  = ~\new_[28808]_  & ~\new_[29898]_ ;
  assign \new_[25059]_  = \new_[28564]_  | \new_[30637]_ ;
  assign \new_[25060]_  = \new_[28643]_  | \new_[30840]_ ;
  assign \new_[25061]_  = ~\new_[28455]_  & ~\new_[30265]_ ;
  assign \new_[25062]_  = \new_[29319]_  | \new_[30273]_ ;
  assign \new_[25063]_  = ~\new_[26956]_ ;
  assign \new_[25064]_  = ~\new_[28450]_  & ~\new_[30711]_ ;
  assign \new_[25065]_  = ~\new_[26973]_ ;
  assign \new_[25066]_  = \new_[28340]_  | \new_[28448]_ ;
  assign \new_[25067]_  = (~\s14_data_i[23]  | ~\new_[30026]_ ) & (~\s12_data_i[23]  | ~\new_[29711]_ );
  assign \new_[25068]_  = ~\new_[28450]_  & ~\new_[30093]_ ;
  assign \new_[25069]_  = \new_[29284]_  | \new_[30036]_ ;
  assign \new_[25070]_  = ~\new_[28311]_  | ~\new_[30552]_ ;
  assign \new_[25071]_  = ~\new_[28571]_  | ~\new_[29892]_ ;
  assign \new_[25072]_  = ~\new_[6071]_  | ~\new_[30600]_  | ~\new_[30538]_ ;
  assign \new_[25073]_  = ~\new_[28479]_  | ~\new_[30774]_ ;
  assign \new_[25074]_  = ~\new_[28439]_  | ~\new_[28072]_ ;
  assign \new_[25075]_  = \new_[28526]_  & \new_[29079]_ ;
  assign \new_[25076]_  = ~\new_[27072]_ ;
  assign \new_[25077]_  = ~\new_[6059]_  | ~\new_[29967]_  | ~\new_[30615]_ ;
  assign \new_[25078]_  = ~\new_[28167]_  & ~\new_[30564]_ ;
  assign \new_[25079]_  = ~\new_[27993]_  | ~\new_[30507]_ ;
  assign \new_[25080]_  = ~\new_[28240]_  | ~\new_[29927]_ ;
  assign \new_[25081]_  = ~\new_[6038]_  | ~\new_[29220]_  | ~\new_[30215]_ ;
  assign \new_[25082]_  = ~\new_[28561]_  & ~\new_[30286]_ ;
  assign \new_[25083]_  = ~\new_[6001]_  | ~\new_[29386]_  | ~\new_[30707]_ ;
  assign \new_[25084]_  = \new_[28484]_  | \new_[30244]_ ;
  assign \new_[25085]_  = \new_[29442]_  & \new_[28183]_ ;
  assign \new_[25086]_  = \new_[28480]_  | \new_[30173]_ ;
  assign \new_[25087]_  = \new_[28228]_  | \new_[28456]_ ;
  assign \new_[25088]_  = \new_[28228]_  & \new_[29527]_ ;
  assign \new_[25089]_  = \new_[28456]_  & \new_[29527]_ ;
  assign \new_[25090]_  = \new_[28452]_  | \new_[30557]_ ;
  assign \new_[25091]_  = \new_[28438]_  | \new_[29855]_ ;
  assign \new_[25092]_  = \new_[29489]_  & \new_[30717]_ ;
  assign \new_[25093]_  = \new_[29500]_  & \new_[30828]_ ;
  assign \new_[25094]_  = \new_[28547]_  | \new_[30070]_ ;
  assign \new_[25095]_  = \new_[28856]_  & \new_[6190]_ ;
  assign \new_[25096]_  = \new_[28434]_  | \new_[30688]_ ;
  assign \new_[25097]_  = \new_[28389]_  & \new_[30582]_ ;
  assign \new_[25098]_  = \new_[29451]_  & \new_[28888]_ ;
  assign \new_[25099]_  = \new_[28528]_  | \new_[30240]_ ;
  assign \new_[25100]_  = ~\new_[28096]_  | ~\new_[29022]_ ;
  assign \new_[25101]_  = ~\new_[28747]_  & ~\new_[29883]_ ;
  assign \new_[25102]_  = \new_[28221]_  & \new_[29867]_ ;
  assign \new_[25103]_  = ~\new_[28534]_  | ~\new_[30735]_ ;
  assign \new_[25104]_  = \new_[28269]_  & \new_[30221]_ ;
  assign \new_[25105]_  = ~\new_[28348]_  & ~\new_[30696]_ ;
  assign \new_[25106]_  = \new_[28674]_  | \new_[30632]_ ;
  assign \new_[25107]_  = ~\new_[28360]_  & ~\new_[30339]_ ;
  assign \new_[25108]_  = ~\new_[28348]_  & ~\new_[30010]_ ;
  assign \new_[25109]_  = \new_[28207]_  | \new_[28904]_ ;
  assign \new_[25110]_  = ~\new_[28455]_  & ~\new_[30543]_ ;
  assign \new_[25111]_  = ~\new_[28471]_  | ~\new_[29537]_ ;
  assign \new_[25112]_  = ~\new_[28233]_  | ~\new_[29972]_ ;
  assign \new_[25113]_  = \new_[28322]_  & \new_[29408]_ ;
  assign \new_[25114]_  = ~\new_[26849]_ ;
  assign \new_[25115]_  = ~\new_[26978]_ ;
  assign \new_[25116]_  = \new_[28687]_  & \new_[30283]_ ;
  assign \new_[25117]_  = ~\new_[28207]_  & ~\new_[28984]_ ;
  assign \new_[25118]_  = (~\new_[30284]_  | ~\s11_data_i[10] ) & (~\new_[29420]_  | ~\s8_data_i[10] );
  assign \new_[25119]_  = ~\new_[28593]_  | ~\new_[29201]_ ;
  assign \new_[25120]_  = ~\new_[28086]_  & ~\new_[29955]_ ;
  assign \new_[25121]_  = \new_[28587]_  | \new_[30557]_ ;
  assign \new_[25122]_  = ~\new_[28298]_  & ~\new_[30230]_ ;
  assign \new_[25123]_  = \new_[29414]_  | \new_[30162]_ ;
  assign \new_[25124]_  = ~\new_[28235]_  | ~\new_[29526]_ ;
  assign \new_[25125]_  = (~\new_[29631]_  | ~\s14_data_i[1] ) & (~\new_[29621]_  | ~\s12_data_i[1] );
  assign \new_[25126]_  = ~\new_[26982]_ ;
  assign \new_[25127]_  = ~\new_[26980]_ ;
  assign \new_[25128]_  = (~\s2_data_i[13]  | ~\new_[29625]_ ) & (~\s1_data_i[13]  | ~\new_[29215]_ );
  assign \new_[25129]_  = ~\new_[26846]_ ;
  assign \new_[25130]_  = \new_[28467]_  & \new_[30009]_ ;
  assign \new_[25131]_  = ~\new_[28583]_  | ~\new_[30702]_ ;
  assign \new_[25132]_  = \new_[29467]_  | \new_[30162]_ ;
  assign \new_[25133]_  = ~\new_[28169]_  | ~\new_[29913]_ ;
  assign \new_[25134]_  = ~\new_[28423]_  & ~\new_[30305]_ ;
  assign \new_[25135]_  = \new_[28404]_  | \new_[29774]_ ;
  assign \new_[25136]_  = ~\new_[28468]_  & ~\new_[30545]_ ;
  assign \new_[25137]_  = \new_[28454]_  & \new_[30262]_ ;
  assign \new_[25138]_  = ~\new_[28478]_  & ~\new_[30708]_ ;
  assign \new_[25139]_  = \new_[28318]_  | \new_[29861]_ ;
  assign \new_[25140]_  = \new_[28427]_  | \new_[30607]_ ;
  assign \new_[25141]_  = ~\new_[28410]_  & ~\new_[30219]_ ;
  assign \new_[25142]_  = \new_[28301]_  | \new_[28428]_ ;
  assign \new_[25143]_  = ~\new_[28099]_  | ~\new_[30724]_ ;
  assign \new_[25144]_  = \new_[28847]_  | \new_[30276]_ ;
  assign \new_[25145]_  = \new_[28534]_  & \new_[30764]_ ;
  assign \new_[25146]_  = \new_[28391]_  & \new_[30764]_ ;
  assign \new_[25147]_  = \new_[29009]_  | \new_[30276]_ ;
  assign \new_[25148]_  = (~\new_[29953]_  | ~\s11_data_i[5] ) & (~\new_[29627]_  | ~\s8_data_i[5] );
  assign \new_[25149]_  = ~\new_[28388]_  | ~\new_[29255]_ ;
  assign \new_[25150]_  = \new_[28074]_  & \new_[28152]_ ;
  assign \new_[25151]_  = ~\new_[28415]_  & ~\new_[28933]_ ;
  assign \new_[25152]_  = \new_[28000]_  & \new_[28127]_ ;
  assign \new_[25153]_  = ~\new_[28421]_  & (~\new_[30828]_  | ~\new_[6174]_ );
  assign \new_[25154]_  = ~\new_[5903]_  | ~\new_[29888]_  | ~\new_[29721]_ ;
  assign \new_[25155]_  = ~\new_[28614]_  & ~\new_[30577]_ ;
  assign \new_[25156]_  = ~\new_[5902]_  | ~\new_[30092]_  | ~\new_[28963]_ ;
  assign \new_[25157]_  = ~\new_[5895]_  | ~\new_[30097]_  | ~\new_[29527]_ ;
  assign \new_[25158]_  = ~\new_[27939]_ ;
  assign \new_[25159]_  = ~\new_[28302]_  | ~\new_[28575]_ ;
  assign \new_[25160]_  = ~\new_[5911]_  | ~\new_[28102]_  | ~\new_[30415]_ ;
  assign \new_[25161]_  = ~\new_[5898]_  | ~\new_[29762]_  | ~\new_[29103]_ ;
  assign \new_[25162]_  = ~\new_[6184]_  | ~\new_[30352]_  | ~\new_[30719]_ ;
  assign \new_[25163]_  = ~\new_[6216]_  | ~\new_[30262]_  | ~\new_[30799]_ ;
  assign \new_[25164]_  = ~\new_[28461]_  | ~\new_[28520]_ ;
  assign \new_[25165]_  = ~\new_[5912]_  | ~\new_[28015]_  | ~\new_[30202]_ ;
  assign \new_[25166]_  = \new_[29539]_  & \new_[27990]_ ;
  assign \new_[25167]_  = ~\new_[5897]_  | ~\new_[30172]_  | ~\new_[29228]_ ;
  assign \new_[25168]_  = ~\new_[28137]_  | ~\new_[28500]_ ;
  assign \new_[25169]_  = ~\new_[6096]_  | ~\new_[30505]_  | ~\new_[30573]_ ;
  assign \new_[25170]_  = ~\new_[28672]_  & (~\new_[30015]_  | ~\new_[6203]_ );
  assign \new_[25171]_  = ~\new_[6083]_  | ~\new_[28692]_  | ~\new_[30140]_ ;
  assign \new_[25172]_  = ~\new_[32134]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25173]_  = ~\new_[6045]_  | ~\new_[28015]_  | ~\new_[30202]_ ;
  assign \new_[25174]_  = (~\new_[29953]_  | ~\s11_data_i[15] ) & (~\new_[29627]_  | ~\s8_data_i[15] );
  assign \new_[25175]_  = ~\new_[31712]_  | ~\new_[30037]_  | ~\new_[30695]_ ;
  assign \new_[25176]_  = ~\new_[27165]_ ;
  assign \new_[25177]_  = ~\new_[31429]_  | ~\new_[29984]_  | ~\new_[29929]_ ;
  assign \new_[25178]_  = ~\new_[28369]_  & ~\new_[28504]_ ;
  assign \new_[25179]_  = ~\new_[28425]_  | ~\new_[28373]_ ;
  assign \new_[25180]_  = ~\new_[31440]_  | ~\new_[30728]_  | ~\new_[30555]_ ;
  assign \new_[25181]_  = ~\new_[5900]_  | ~\new_[29904]_  | ~\new_[29441]_ ;
  assign \new_[25182]_  = ~\new_[30375]_  & ~\new_[30572]_ ;
  assign \new_[25183]_  = ~\new_[5906]_  | ~\new_[30159]_  | ~\new_[29456]_ ;
  assign \new_[25184]_  = (~\new_[29012]_  | ~\s10_data_i[15] ) & (~\new_[29185]_  | ~\s9_data_i[15] );
  assign \new_[25185]_  = ~\new_[28725]_  & (~\new_[30638]_  | ~\new_[6211]_ );
  assign \new_[25186]_  = (~\new_[29631]_  | ~\s14_data_i[0] ) & (~\new_[29621]_  | ~\s12_data_i[0] );
  assign \new_[25187]_  = ~\new_[28808]_  | ~\new_[28108]_ ;
  assign \new_[25188]_  = ~\new_[28199]_  & (~\new_[30571]_  | ~\new_[6186]_ );
  assign \new_[25189]_  = ~\new_[5926]_  | ~\new_[28488]_  | ~\new_[29944]_ ;
  assign \new_[25190]_  = ~\new_[28336]_  | ~\new_[28631]_ ;
  assign \new_[25191]_  = ~\new_[5904]_  | ~\new_[29863]_  | ~\new_[29006]_ ;
  assign \new_[25192]_  = ~\new_[6074]_  | ~\new_[28649]_  | ~\new_[30058]_ ;
  assign \new_[25193]_  = ~\new_[6042]_  | ~\new_[28102]_  | ~\new_[30415]_ ;
  assign \new_[25194]_  = ~\new_[28655]_  & (~\new_[30693]_  | ~\new_[6214]_ );
  assign \new_[25195]_  = ~\new_[28704]_  | ~\new_[28222]_ ;
  assign \new_[25196]_  = ~\new_[5921]_  | ~\new_[28649]_  | ~\new_[30058]_ ;
  assign \new_[25197]_  = ~\new_[28103]_  & (~\new_[29987]_  | ~\new_[5992]_ );
  assign \new_[25198]_  = \new_[29551]_  & \new_[28178]_ ;
  assign \new_[25199]_  = ~\new_[31232]_  | ~\new_[28283]_  | ~\new_[30409]_ ;
  assign \new_[25200]_  = \new_[29098]_  & \new_[28411]_ ;
  assign \new_[25201]_  = \new_[28448]_  & \new_[29006]_ ;
  assign \new_[25202]_  = ~\new_[6096]_  | ~\new_[29780]_  | ~\new_[30505]_ ;
  assign \new_[25203]_  = ~\new_[5927]_  | ~\new_[28692]_  | ~\new_[30140]_ ;
  assign \new_[25204]_  = (~\new_[30200]_  | ~\s11_data_i[1] ) & (~\new_[29428]_  | ~\s8_data_i[1] );
  assign \new_[25205]_  = (~\new_[29036]_  | ~\s5_data_i[3] ) & (~\new_[30429]_  | ~\s3_data_i[3] );
  assign \new_[25206]_  = ~\new_[28811]_  | ~\new_[28474]_ ;
  assign \new_[25207]_  = ~\new_[28676]_  & (~\new_[30691]_  | ~\new_[6197]_ );
  assign \new_[25208]_  = ~\new_[6210]_  | ~\new_[30645]_  | ~\new_[30782]_ ;
  assign \new_[25209]_  = ~\new_[26728]_ ;
  assign \new_[25210]_  = ~\new_[29640]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[25211]_  = \new_[29289]_  & \new_[28276]_ ;
  assign \new_[25212]_  = (~\new_[29953]_  | ~\s11_data_i[16] ) & (~\new_[29627]_  | ~\s8_data_i[16] );
  assign \new_[25213]_  = ~\new_[27731]_ ;
  assign \new_[25214]_  = ~\new_[28407]_  & (~\new_[30233]_  | ~\new_[6095]_ );
  assign \new_[25215]_  = (~\new_[30227]_  | ~\s10_data_i[14] ) & (~\new_[29706]_  | ~\s9_data_i[14] );
  assign \new_[25216]_  = ~\new_[29749]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25217]_  = (~\new_[30284]_  | ~\s11_data_i[3] ) & (~\new_[29420]_  | ~\s8_data_i[3] );
  assign \new_[25218]_  = ~\new_[29205]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25219]_  = ~\new_[29711]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25220]_  = ~\new_[29625]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25221]_  = ~\new_[29035]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25222]_  = ~\new_[29649]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25223]_  = ~\new_[29708]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25224]_  = ~\new_[29241]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25225]_  = ~\new_[29034]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[25226]_  = ~\new_[28957]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25227]_  = ~\new_[32321]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25228]_  = ~\new_[29025]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25229]_  = ~\new_[29052]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25230]_  = ~\new_[29670]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25231]_  = ~\new_[29021]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[25232]_  = ~\new_[29709]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[25233]_  = (~\new_[29012]_  | ~\s10_data_i[16] ) & (~\new_[29185]_  | ~\s9_data_i[16] );
  assign \new_[25234]_  = ~\new_[29710]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[25235]_  = ~\new_[29428]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[25236]_  = ~\new_[29024]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[25237]_  = ~\new_[29012]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25238]_  = ~\new_[29317]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25239]_  = ~\new_[28132]_  & ~\m6_addr_i[28] ;
  assign \new_[25240]_  = ~\new_[28851]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25241]_  = ~\new_[29641]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25242]_  = ~\new_[29627]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25243]_  = ~\new_[29185]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[25244]_  = ~\new_[29045]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[25245]_  = ~\new_[32260]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[25246]_  = ~\new_[29628]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[25247]_  = ~\new_[29636]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[25248]_  = ~\new_[28801]_  | ~\new_[6048]_ ;
  assign \new_[25249]_  = ~\new_[29621]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25250]_  = ~\new_[29149]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25251]_  = (~\new_[29149]_  | ~\s4_data_i[3] ) & (~\new_[29651]_  | ~\s0_data_i[3] );
  assign \new_[25252]_  = ~\new_[29036]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25253]_  = ~\new_[28081]_  | ~\new_[29038]_ ;
  assign \new_[25254]_  = ~\new_[30243]_  & ~\new_[28609]_ ;
  assign \new_[25255]_  = ~\new_[29420]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25256]_  = ~\new_[29706]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[25257]_  = ~\new_[29604]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[25258]_  = ~\new_[29579]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[25259]_  = ~\new_[29534]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[25260]_  = ~\new_[29707]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[25261]_  = ~\new_[29298]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[25262]_  = ~\new_[28842]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25263]_  = ~\new_[29705]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[25264]_  = ~\new_[6080]_  | ~\new_[28488]_  | ~\new_[29944]_ ;
  assign \new_[25265]_  = ~\new_[28544]_  | ~\new_[28181]_ ;
  assign \new_[25266]_  = ~\new_[28568]_  & (~\new_[29869]_  | ~\new_[6213]_ );
  assign \new_[25267]_  = ~\new_[5907]_  | ~\new_[30016]_  | ~\new_[28898]_ ;
  assign \new_[25268]_  = ~\new_[5908]_  | ~\new_[29557]_  | ~\new_[29226]_ ;
  assign \new_[25269]_  = \new_[28478]_  & \new_[28128]_ ;
  assign \new_[25270]_  = ~\new_[28016]_  & (~\new_[30641]_  | ~\new_[6093]_ );
  assign \new_[25271]_  = ~\new_[5894]_  | ~\new_[29900]_  | ~\new_[30150]_ ;
  assign \new_[25272]_  = (~\new_[30060]_  | ~\s7_data_i[6] ) & (~\new_[29704]_  | ~\s6_data_i[6] );
  assign \new_[25273]_  = ~\new_[27048]_ ;
  assign \new_[25274]_  = (~\s4_data_i[16]  | ~\new_[30335]_ ) & (~\s0_data_i[16]  | ~\new_[29603]_ );
  assign \new_[25275]_  = (~\new_[30181]_  | ~\s14_data_i[5] ) & (~\new_[29640]_  | ~\s12_data_i[5] );
  assign \new_[25276]_  = (~\s10_data_i[29]  | ~\new_[29749]_ ) & (~\s9_data_i[29]  | ~\new_[29034]_ );
  assign \new_[25277]_  = (~\s5_data_i[8]  | ~\new_[29649]_ ) & (~\s3_data_i[8]  | ~\new_[29035]_ );
  assign \new_[25278]_  = (~\new_[29628]_  | ~\s4_data_i[4] ) & (~\new_[29258]_  | ~\s0_data_i[4] );
  assign \new_[25279]_  = (~\new_[29534]_  | ~\s5_data_i[6] ) & (~\new_[29579]_  | ~\s3_data_i[6] );
  assign \new_[25280]_  = (~\new_[30060]_  | ~\s7_data_i[4] ) & (~\new_[29704]_  | ~\s6_data_i[4] );
  assign \new_[25281]_  = (~\new_[30060]_  | ~\s7_data_i[12] ) & (~\new_[29704]_  | ~\s6_data_i[12] );
  assign \new_[25282]_  = (~\s14_data_i[22]  | ~\new_[30026]_ ) & (~\s12_data_i[22]  | ~\new_[29711]_ );
  assign \new_[25283]_  = (~\new_[29045]_  | ~\s10_data_i[3] ) & (~\new_[29951]_  | ~\s9_data_i[3] );
  assign \new_[25284]_  = (~\new_[29628]_  | ~\s4_data_i[12] ) & (~\new_[29258]_  | ~\s0_data_i[12] );
  assign \new_[25285]_  = (~\new_[29012]_  | ~\s10_data_i[17] ) & (~\new_[29185]_  | ~\s9_data_i[17] );
  assign \new_[25286]_  = (~\new_[30181]_  | ~\s14_data_i[3] ) & (~\new_[29640]_  | ~\s12_data_i[3] );
  assign \new_[25287]_  = (~\new_[30311]_  | ~\s11_data_i[1] ) & (~\new_[29636]_  | ~\s8_data_i[1] );
  assign \new_[25288]_  = (~\new_[30031]_  | ~\s7_data_i[15] ) & (~\new_[29052]_  | ~\s6_data_i[15] );
  assign \new_[25289]_  = (~\new_[29025]_  | ~\s5_data_i[4] ) & (~\new_[30469]_  | ~\s3_data_i[4] );
  assign \new_[25290]_  = (~\new_[29045]_  | ~\s10_data_i[2] ) & (~\new_[29951]_  | ~\s9_data_i[2] );
  assign \new_[25291]_  = (~\s5_data_i[23]  | ~\new_[29649]_ ) & (~\s3_data_i[23]  | ~\new_[29035]_ );
  assign \new_[25292]_  = (~\new_[30311]_  | ~\s11_data_i[2] ) & (~\new_[29636]_  | ~\s8_data_i[2] );
  assign \new_[25293]_  = (~\s10_data_i[16]  | ~\new_[29749]_ ) & (~\s9_data_i[16]  | ~\new_[29034]_ );
  assign \new_[25294]_  = (~\s5_data_i[16]  | ~\new_[29649]_ ) & (~\s3_data_i[16]  | ~\new_[29035]_ );
  assign \new_[25295]_  = (~\new_[30060]_  | ~\s7_data_i[1] ) & (~\new_[29704]_  | ~\s6_data_i[1] );
  assign \new_[25296]_  = (~\new_[29045]_  | ~\s10_data_i[1] ) & (~\new_[29951]_  | ~\s9_data_i[1] );
  assign \new_[25297]_  = (~\new_[30181]_  | ~\s14_data_i[1] ) & (~\new_[29640]_  | ~\s12_data_i[1] );
  assign \new_[25298]_  = (~\new_[29045]_  | ~\s10_data_i[0] ) & (~\new_[29951]_  | ~\s9_data_i[0] );
  assign \new_[25299]_  = ~\new_[27058]_ ;
  assign \new_[25300]_  = (~\new_[30311]_  | ~\s11_data_i[0] ) & (~\new_[29636]_  | ~\s8_data_i[0] );
  assign \new_[25301]_  = (~\s11_data_i[25]  | ~\new_[29205]_ ) & (~\s8_data_i[25]  | ~\new_[29241]_ );
  assign \new_[25302]_  = (~\new_[30311]_  | ~\s11_data_i[13] ) & (~\new_[29636]_  | ~\s8_data_i[13] );
  assign \new_[25303]_  = (~\s11_data_i[16]  | ~\new_[29205]_ ) & (~\s8_data_i[16]  | ~\new_[29241]_ );
  assign \new_[25304]_  = (~\s4_data_i[10]  | ~\new_[30335]_ ) & (~\s0_data_i[10]  | ~\new_[29603]_ );
  assign \new_[25305]_  = (~\new_[30260]_  | ~\s11_data_i[8] ) & (~\new_[29670]_  | ~\s8_data_i[8] );
  assign \new_[25306]_  = (~\new_[29534]_  | ~\s5_data_i[22] ) & (~\new_[29579]_  | ~\s3_data_i[22] );
  assign \new_[25307]_  = (~\new_[28842]_  | ~\s4_data_i[19] ) & (~\new_[29434]_  | ~\s0_data_i[19] );
  assign \new_[25308]_  = (~\s14_data_i[6]  | ~\new_[30026]_ ) & (~\s12_data_i[6]  | ~\new_[29711]_ );
  assign \new_[25309]_  = (~\new_[29631]_  | ~\s14_data_i[14] ) & (~\new_[29621]_  | ~\s12_data_i[14] );
  assign \new_[25310]_  = (~\s14_data_i[27]  | ~\new_[30026]_ ) & (~\s12_data_i[27]  | ~\new_[29711]_ );
  assign \new_[25311]_  = (~\new_[29705]_  | ~\s10_data_i[23] ) & (~\new_[30354]_  | ~\s9_data_i[23] );
  assign \new_[25312]_  = (~\new_[29976]_  | ~\s14_data_i[17] ) & (~\new_[28957]_  | ~\s12_data_i[17] );
  assign \new_[25313]_  = ~\new_[28801]_  | ~\new_[6200]_ ;
  assign \new_[25314]_  = (~\new_[30193]_  | ~\s7_data_i[25] ) & (~\new_[29298]_  | ~\s6_data_i[25] );
  assign \new_[25315]_  = ~\new_[27088]_ ;
  assign \new_[25316]_  = (~\new_[30200]_  | ~\s11_data_i[22] ) & (~\new_[29428]_  | ~\s8_data_i[22] );
  assign \new_[25317]_  = (~\new_[30200]_  | ~\s11_data_i[15] ) & (~\new_[29428]_  | ~\s8_data_i[15] );
  assign \new_[25318]_  = (~\new_[29025]_  | ~\s5_data_i[30] ) & (~\new_[30469]_  | ~\s3_data_i[30] );
  assign \new_[25319]_  = (~\s2_data_i[27]  | ~\new_[29625]_ ) & (~\s1_data_i[27]  | ~\new_[29215]_ );
  assign \new_[25320]_  = (~\s14_data_i[9]  | ~\new_[30026]_ ) & (~\s12_data_i[9]  | ~\new_[29711]_ );
  assign \new_[25321]_  = (~\new_[30227]_  | ~\s10_data_i[10] ) & (~\new_[29706]_  | ~\s9_data_i[10] );
  assign \new_[25322]_  = (~\new_[29149]_  | ~\s4_data_i[31] ) & (~\new_[29651]_  | ~\s0_data_i[31] );
  assign \new_[25323]_  = (~\new_[29021]_  | ~\s10_data_i[18] ) & (~\new_[29709]_  | ~\s9_data_i[18] );
  assign \new_[25324]_  = (~\new_[30227]_  | ~\s10_data_i[31] ) & (~\new_[29706]_  | ~\s9_data_i[31] );
  assign \new_[25325]_  = (~\s10_data_i[10]  | ~\new_[29749]_ ) & (~\s9_data_i[10]  | ~\new_[29034]_ );
  assign \new_[25326]_  = (~\s14_data_i[8]  | ~\new_[30026]_ ) & (~\s12_data_i[8]  | ~\new_[29711]_ );
  assign \new_[25327]_  = (~\new_[29710]_  | ~\s10_data_i[15] ) & (~\new_[29024]_  | ~\s9_data_i[15] );
  assign \new_[25328]_  = (~\new_[29631]_  | ~\s14_data_i[31] ) & (~\new_[29621]_  | ~\s12_data_i[31] );
  assign \new_[25329]_  = (~\s11_data_i[14]  | ~\new_[29205]_ ) & (~\s8_data_i[14]  | ~\new_[29241]_ );
  assign \new_[25330]_  = ~\new_[30543]_  | ~\new_[28001]_ ;
  assign \new_[25331]_  = (~\new_[29953]_  | ~\s11_data_i[18] ) & (~\new_[29627]_  | ~\s8_data_i[18] );
  assign \new_[25332]_  = (~\new_[30031]_  | ~\s7_data_i[22] ) & (~\new_[29052]_  | ~\s6_data_i[22] );
  assign \new_[25333]_  = (~\new_[30193]_  | ~\s7_data_i[17] ) & (~\new_[29298]_  | ~\s6_data_i[17] );
  assign \new_[25334]_  = (~\new_[30284]_  | ~\s11_data_i[30] ) & (~\new_[29420]_  | ~\s8_data_i[30] );
  assign \new_[25335]_  = (~\new_[30193]_  | ~\s7_data_i[7] ) & (~\new_[29298]_  | ~\s6_data_i[7] );
  assign \new_[25336]_  = (~\new_[29149]_  | ~\s4_data_i[7] ) & (~\new_[29651]_  | ~\s0_data_i[7] );
  assign \new_[25337]_  = (~\new_[30031]_  | ~\s7_data_i[31] ) & (~\new_[29052]_  | ~\s6_data_i[31] );
  assign \new_[25338]_  = (~\new_[29705]_  | ~\s10_data_i[18] ) & (~\new_[30354]_  | ~\s9_data_i[18] );
  assign \new_[25339]_  = (~\new_[30227]_  | ~\s10_data_i[29] ) & (~\new_[29706]_  | ~\s9_data_i[29] );
  assign \new_[25340]_  = (~\new_[30181]_  | ~\s14_data_i[14] ) & (~\new_[29640]_  | ~\s12_data_i[14] );
  assign \new_[25341]_  = ~\new_[27081]_ ;
  assign \new_[25342]_  = (~\s14_data_i[26]  | ~\new_[30026]_ ) & (~\s12_data_i[26]  | ~\new_[29711]_ );
  assign \new_[25343]_  = (~\new_[30026]_  | ~\s14_data_i[31] ) & (~\new_[29711]_  | ~\s12_data_i[31] );
  assign \new_[25344]_  = (~\new_[30227]_  | ~\s10_data_i[6] ) & (~\new_[29706]_  | ~\s9_data_i[6] );
  assign \new_[25345]_  = (~\new_[29036]_  | ~\s5_data_i[11] ) & (~\new_[30429]_  | ~\s3_data_i[11] );
  assign \new_[25346]_  = (~\new_[30284]_  | ~\s11_data_i[28] ) & (~\new_[29420]_  | ~\s8_data_i[28] );
  assign \new_[25347]_  = (~\new_[30031]_  | ~\s7_data_i[30] ) & (~\new_[29052]_  | ~\s6_data_i[30] );
  assign \new_[25348]_  = (~\new_[30311]_  | ~\s11_data_i[14] ) & (~\new_[29636]_  | ~\s8_data_i[14] );
  assign \new_[25349]_  = (~\new_[29045]_  | ~\s10_data_i[14] ) & (~\new_[29951]_  | ~\s9_data_i[14] );
  assign \new_[25350]_  = (~\new_[30227]_  | ~\s10_data_i[27] ) & (~\new_[29706]_  | ~\s9_data_i[27] );
  assign \new_[25351]_  = ~\new_[27093]_ ;
  assign \new_[25352]_  = (~\new_[29149]_  | ~\s4_data_i[26] ) & (~\new_[29651]_  | ~\s0_data_i[26] );
  assign \new_[25353]_  = (~\new_[29976]_  | ~\s14_data_i[29] ) & (~\new_[28957]_  | ~\s12_data_i[29] );
  assign \new_[25354]_  = (~\new_[30284]_  | ~\s11_data_i[26] ) & (~\new_[29420]_  | ~\s8_data_i[26] );
  assign \new_[25355]_  = (~\new_[29631]_  | ~\s14_data_i[26] ) & (~\new_[29621]_  | ~\s12_data_i[26] );
  assign \new_[25356]_  = (~\new_[29021]_  | ~\s10_data_i[15] ) & (~\new_[29709]_  | ~\s9_data_i[15] );
  assign \new_[25357]_  = ~\new_[30682]_  & ~\new_[30620]_ ;
  assign \new_[25358]_  = (~\new_[30060]_  | ~\s7_data_i[14] ) & (~\new_[29704]_  | ~\s6_data_i[14] );
  assign \new_[25359]_  = (~\new_[29012]_  | ~\s10_data_i[30] ) & (~\new_[29185]_  | ~\s9_data_i[30] );
  assign \new_[25360]_  = (~\new_[29012]_  | ~\s10_data_i[18] ) & (~\new_[29185]_  | ~\s9_data_i[18] );
  assign \new_[25361]_  = (~\new_[29149]_  | ~\s4_data_i[25] ) & (~\new_[29651]_  | ~\s0_data_i[25] );
  assign \new_[25362]_  = ~\new_[27095]_ ;
  assign \new_[25363]_  = (~\new_[29631]_  | ~\s14_data_i[25] ) & (~\new_[29621]_  | ~\s12_data_i[25] );
  assign \new_[25364]_  = (~\new_[30200]_  | ~\s11_data_i[17] ) & (~\new_[29428]_  | ~\s8_data_i[17] );
  assign \new_[25365]_  = (~\new_[29036]_  | ~\s5_data_i[25] ) & (~\new_[30429]_  | ~\s3_data_i[25] );
  assign \new_[25366]_  = (~\s10_data_i[5]  | ~\new_[29749]_ ) & (~\s9_data_i[5]  | ~\new_[29034]_ );
  assign \new_[25367]_  = (~\new_[29631]_  | ~\s14_data_i[6] ) & (~\new_[29621]_  | ~\s12_data_i[6] );
  assign \new_[25368]_  = (~\new_[29628]_  | ~\s4_data_i[14] ) & (~\new_[29258]_  | ~\s0_data_i[14] );
  assign \new_[25369]_  = (~\s5_data_i[13]  | ~\new_[29649]_ ) & (~\s3_data_i[13]  | ~\new_[29035]_ );
  assign \new_[25370]_  = (~\new_[29631]_  | ~\s14_data_i[24] ) & (~\new_[29621]_  | ~\s12_data_i[24] );
  assign \new_[25371]_  = (~\new_[29149]_  | ~\s4_data_i[23] ) & (~\new_[29651]_  | ~\s0_data_i[23] );
  assign \new_[25372]_  = (~\s11_data_i[15]  | ~\new_[29205]_ ) & (~\s8_data_i[15]  | ~\new_[29241]_ );
  assign \new_[25373]_  = (~\new_[29149]_  | ~\s4_data_i[11] ) & (~\new_[29651]_  | ~\s0_data_i[11] );
  assign \new_[25374]_  = (~\new_[30227]_  | ~\s10_data_i[23] ) & (~\new_[29706]_  | ~\s9_data_i[23] );
  assign \new_[25375]_  = (~\new_[30284]_  | ~\s11_data_i[23] ) & (~\new_[29420]_  | ~\s8_data_i[23] );
  assign \new_[25376]_  = (~\s4_data_i[22]  | ~\new_[30335]_ ) & (~\s0_data_i[22]  | ~\new_[29603]_ );
  assign \new_[25377]_  = (~\s5_data_i[14]  | ~\new_[29649]_ ) & (~\s3_data_i[14]  | ~\new_[29035]_ );
  assign \new_[25378]_  = (~\s14_data_i[15]  | ~\new_[30026]_ ) & (~\s12_data_i[15]  | ~\new_[29711]_ );
  assign \new_[25379]_  = (~\s10_data_i[23]  | ~\new_[29749]_ ) & (~\s9_data_i[23]  | ~\new_[29034]_ );
  assign \new_[25380]_  = ~\new_[26958]_ ;
  assign \new_[25381]_  = (~\new_[29631]_  | ~\s14_data_i[22] ) & (~\new_[29621]_  | ~\s12_data_i[22] );
  assign \new_[25382]_  = (~\new_[29036]_  | ~\s5_data_i[22] ) & (~\new_[30429]_  | ~\s3_data_i[22] );
  assign \new_[25383]_  = (~\s4_data_i[8]  | ~\new_[30335]_ ) & (~\s0_data_i[8]  | ~\new_[29603]_ );
  assign \new_[25384]_  = (~\new_[29012]_  | ~\s10_data_i[28] ) & (~\new_[29185]_  | ~\s9_data_i[28] );
  assign \new_[25385]_  = (~\new_[29149]_  | ~\s4_data_i[21] ) & (~\new_[29651]_  | ~\s0_data_i[21] );
  assign \new_[25386]_  = ~\new_[27564]_ ;
  assign \new_[25387]_  = (~\new_[29641]_  | ~\s14_data_i[26] ) & (~\new_[29317]_  | ~\s12_data_i[26] );
  assign \new_[25388]_  = (~\new_[30193]_  | ~\s7_data_i[5] ) & (~\new_[29298]_  | ~\s6_data_i[5] );
  assign \new_[25389]_  = (~\new_[30227]_  | ~\s10_data_i[21] ) & (~\new_[29706]_  | ~\s9_data_i[21] );
  assign \new_[25390]_  = (~\s2_data_i[30]  | ~\new_[29625]_ ) & (~\s1_data_i[30]  | ~\new_[29215]_ );
  assign \new_[25391]_  = (~\new_[29710]_  | ~\s10_data_i[20] ) & (~\new_[29024]_  | ~\s9_data_i[20] );
  assign \new_[25392]_  = (~\new_[29631]_  | ~\s14_data_i[12] ) & (~\new_[29621]_  | ~\s12_data_i[12] );
  assign \new_[25393]_  = (~\new_[30193]_  | ~\s7_data_i[12] ) & (~\new_[29298]_  | ~\s6_data_i[12] );
  assign \new_[25394]_  = (~\new_[30260]_  | ~\s11_data_i[19] ) & (~\new_[29670]_  | ~\s8_data_i[19] );
  assign \new_[25395]_  = (~\new_[29021]_  | ~\s10_data_i[12] ) & (~\new_[29709]_  | ~\s9_data_i[12] );
  assign \new_[25396]_  = (~\new_[30284]_  | ~\s11_data_i[20] ) & (~\new_[29420]_  | ~\s8_data_i[20] );
  assign \new_[25397]_  = (~\new_[29631]_  | ~\s14_data_i[20] ) & (~\new_[29621]_  | ~\s12_data_i[20] );
  assign \new_[25398]_  = (~\new_[29036]_  | ~\s5_data_i[20] ) & (~\new_[30429]_  | ~\s3_data_i[20] );
  assign \new_[25399]_  = (~\new_[29149]_  | ~\s4_data_i[19] ) & (~\new_[29651]_  | ~\s0_data_i[19] );
  assign \new_[25400]_  = (~\new_[30284]_  | ~\s11_data_i[19] ) & (~\new_[29420]_  | ~\s8_data_i[19] );
  assign \new_[25401]_  = (~\new_[29631]_  | ~\s14_data_i[19] ) & (~\new_[29621]_  | ~\s12_data_i[19] );
  assign \new_[25402]_  = (~\s11_data_i[8]  | ~\new_[29205]_ ) & (~\s8_data_i[8]  | ~\new_[29241]_ );
  assign \new_[25403]_  = (~\new_[29036]_  | ~\s5_data_i[19] ) & (~\new_[30429]_  | ~\s3_data_i[19] );
  assign \new_[25404]_  = (~\s4_data_i[5]  | ~\new_[30335]_ ) & (~\s0_data_i[5]  | ~\new_[29603]_ );
  assign \new_[25405]_  = (~\new_[30227]_  | ~\s10_data_i[4] ) & (~\new_[29706]_  | ~\s9_data_i[4] );
  assign \new_[25406]_  = (~\new_[29149]_  | ~\s4_data_i[18] ) & (~\new_[29651]_  | ~\s0_data_i[18] );
  assign \new_[25407]_  = (~\new_[30193]_  | ~\s7_data_i[11] ) & (~\new_[29298]_  | ~\s6_data_i[11] );
  assign \new_[25408]_  = (~\new_[29631]_  | ~\s14_data_i[18] ) & (~\new_[29621]_  | ~\s12_data_i[18] );
  assign \new_[25409]_  = ~\new_[27114]_ ;
  assign \new_[25410]_  = ~\new_[27115]_ ;
  assign \new_[25411]_  = (~\new_[28842]_  | ~\s4_data_i[26] ) & (~\new_[29434]_  | ~\s0_data_i[26] );
  assign \new_[25412]_  = (~\new_[29149]_  | ~\s4_data_i[17] ) & (~\new_[29651]_  | ~\s0_data_i[17] );
  assign \new_[25413]_  = ~\new_[29299]_  | ~\new_[5989]_ ;
  assign \new_[25414]_  = (~\s10_data_i[30]  | ~\new_[29749]_ ) & (~\s9_data_i[30]  | ~\new_[29034]_ );
  assign \new_[25415]_  = (~\new_[30060]_  | ~\s7_data_i[15] ) & (~\new_[29704]_  | ~\s6_data_i[15] );
  assign \new_[25416]_  = (~\new_[29631]_  | ~\s14_data_i[17] ) & (~\new_[29621]_  | ~\s12_data_i[17] );
  assign \new_[25417]_  = (~\s4_data_i[14]  | ~\new_[30335]_ ) & (~\s0_data_i[14]  | ~\new_[29603]_ );
  assign \new_[25418]_  = ~\new_[27120]_ ;
  assign \new_[25419]_  = (~\new_[29036]_  | ~\s5_data_i[16] ) & (~\new_[30429]_  | ~\s3_data_i[16] );
  assign \new_[25420]_  = (~\new_[29976]_  | ~\s14_data_i[24] ) & (~\new_[28957]_  | ~\s12_data_i[24] );
  assign \new_[25421]_  = (~\new_[29149]_  | ~\s4_data_i[15] ) & (~\new_[29651]_  | ~\s0_data_i[15] );
  assign \new_[25422]_  = (~\new_[29628]_  | ~\s4_data_i[15] ) & (~\new_[29258]_  | ~\s0_data_i[15] );
  assign \new_[25423]_  = (~\new_[30227]_  | ~\s10_data_i[15] ) & (~\new_[29706]_  | ~\s9_data_i[15] );
  assign \new_[25424]_  = (~\s11_data_i[26]  | ~\new_[29205]_ ) & (~\s8_data_i[26]  | ~\new_[29241]_ );
  assign \new_[25425]_  = (~\new_[30200]_  | ~\s11_data_i[18] ) & (~\new_[29428]_  | ~\s8_data_i[18] );
  assign \new_[25426]_  = (~\new_[29631]_  | ~\s14_data_i[15] ) & (~\new_[29621]_  | ~\s12_data_i[15] );
  assign \new_[25427]_  = (~\new_[30260]_  | ~\s11_data_i[30] ) & (~\new_[29670]_  | ~\s8_data_i[30] );
  assign \new_[25428]_  = (~\s10_data_i[14]  | ~\new_[29749]_ ) & (~\s9_data_i[14]  | ~\new_[29034]_ );
  assign \new_[25429]_  = (~\new_[30284]_  | ~\s11_data_i[14] ) & (~\new_[29420]_  | ~\s8_data_i[14] );
  assign \new_[25430]_  = (~\new_[29012]_  | ~\s10_data_i[27] ) & (~\new_[29185]_  | ~\s9_data_i[27] );
  assign \new_[25431]_  = (~\new_[29641]_  | ~\s14_data_i[9] ) & (~\new_[29317]_  | ~\s12_data_i[9] );
  assign \new_[25432]_  = (~\new_[30227]_  | ~\s10_data_i[13] ) & (~\new_[29706]_  | ~\s9_data_i[13] );
  assign \new_[25433]_  = (~\new_[30200]_  | ~\s11_data_i[16] ) & (~\new_[29428]_  | ~\s8_data_i[16] );
  assign \new_[25434]_  = (~\s14_data_i[29]  | ~\new_[30026]_ ) & (~\s12_data_i[29]  | ~\new_[29711]_ );
  assign \new_[25435]_  = (~\new_[30284]_  | ~\s11_data_i[13] ) & (~\new_[29420]_  | ~\s8_data_i[13] );
  assign \new_[25436]_  = (~\new_[29036]_  | ~\s5_data_i[13] ) & (~\new_[30429]_  | ~\s3_data_i[13] );
  assign \new_[25437]_  = (~\new_[29149]_  | ~\s4_data_i[12] ) & (~\new_[29651]_  | ~\s0_data_i[12] );
  assign \new_[25438]_  = (~\new_[30031]_  | ~\s7_data_i[16] ) & (~\new_[29052]_  | ~\s6_data_i[16] );
  assign \new_[25439]_  = ~\new_[27724]_ ;
  assign \new_[25440]_  = (~\new_[29036]_  | ~\s5_data_i[18] ) & (~\new_[30429]_  | ~\s3_data_i[18] );
  assign \new_[25441]_  = (~\new_[30227]_  | ~\s10_data_i[12] ) & (~\new_[29706]_  | ~\s9_data_i[12] );
  assign \new_[25442]_  = (~\new_[30193]_  | ~\s7_data_i[8] ) & (~\new_[29298]_  | ~\s6_data_i[8] );
  assign \new_[25443]_  = ~\new_[27133]_ ;
  assign \new_[25444]_  = (~\new_[29631]_  | ~\s14_data_i[13] ) & (~\new_[29621]_  | ~\s12_data_i[13] );
  assign \new_[25445]_  = (~\new_[30284]_  | ~\s11_data_i[2] ) & (~\new_[29420]_  | ~\s8_data_i[2] );
  assign \new_[25446]_  = (~\new_[29012]_  | ~\s10_data_i[19] ) & (~\new_[29185]_  | ~\s9_data_i[19] );
  assign \new_[25447]_  = ~\new_[27135]_ ;
  assign \new_[25448]_  = (~\new_[29012]_  | ~\s10_data_i[9] ) & (~\new_[29185]_  | ~\s9_data_i[9] );
  assign \new_[25449]_  = (~\new_[29021]_  | ~\s10_data_i[0] ) & (~\new_[29709]_  | ~\s9_data_i[0] );
  assign \new_[25450]_  = (~\new_[30227]_  | ~\s10_data_i[11] ) & (~\new_[29706]_  | ~\s9_data_i[11] );
  assign \new_[25451]_  = (~\new_[30284]_  | ~\s11_data_i[11] ) & (~\new_[29420]_  | ~\s8_data_i[11] );
  assign \new_[25452]_  = (~\new_[29705]_  | ~\s10_data_i[7] ) & (~\new_[30354]_  | ~\s9_data_i[7] );
  assign \new_[25453]_  = ~\new_[27815]_ ;
  assign \new_[25454]_  = (~\new_[30284]_  | ~\s11_data_i[6] ) & (~\new_[29420]_  | ~\s8_data_i[6] );
  assign \new_[25455]_  = (~\new_[29149]_  | ~\s4_data_i[8] ) & (~\new_[29651]_  | ~\s0_data_i[8] );
  assign \new_[25456]_  = ~\new_[27137]_ ;
  assign \new_[25457]_  = ~\new_[27103]_ ;
  assign \new_[25458]_  = (~\new_[29021]_  | ~\s10_data_i[20] ) & (~\new_[29709]_  | ~\s9_data_i[20] );
  assign \new_[25459]_  = ~\new_[27210]_ ;
  assign \new_[25460]_  = ~\new_[30762]_  & ~\new_[26655]_ ;
  assign \new_[25461]_  = (~\new_[29631]_  | ~\s14_data_i[10] ) & (~\new_[29621]_  | ~\s12_data_i[10] );
  assign \new_[25462]_  = (~\new_[29036]_  | ~\s5_data_i[10] ) & (~\new_[30429]_  | ~\s3_data_i[10] );
  assign \new_[25463]_  = \new_[29390]_  & \new_[30786]_ ;
  assign \new_[25464]_  = (~\s14_data_i[10]  | ~\new_[30026]_ ) & (~\s12_data_i[10]  | ~\new_[29711]_ );
  assign \new_[25465]_  = (~\s2_data_i[3]  | ~\new_[29625]_ ) & (~\s1_data_i[3]  | ~\new_[29215]_ );
  assign \new_[25466]_  = ~\new_[30258]_  & ~\new_[30053]_ ;
  assign \new_[25467]_  = (~\new_[30335]_  | ~\s4_data_i[31] ) & (~\new_[29603]_  | ~\s0_data_i[31] );
  assign \new_[25468]_  = (~\new_[30060]_  | ~\s7_data_i[16] ) & (~\new_[29704]_  | ~\s6_data_i[16] );
  assign \new_[25469]_  = ~\new_[28731]_  | ~\new_[29685]_ ;
  assign \new_[25470]_  = (~\new_[29149]_  | ~\s4_data_i[13] ) & (~\new_[29651]_  | ~\s0_data_i[13] );
  assign \new_[25471]_  = (~\s2_data_i[26]  | ~\new_[29625]_ ) & (~\s1_data_i[26]  | ~\new_[29215]_ );
  assign \new_[25472]_  = (~\new_[29534]_  | ~\s5_data_i[23] ) & (~\new_[29579]_  | ~\s3_data_i[23] );
  assign \new_[25473]_  = (~\new_[30193]_  | ~\s7_data_i[29] ) & (~\new_[29298]_  | ~\s6_data_i[29] );
  assign \new_[25474]_  = (~\new_[30284]_  | ~\s11_data_i[8] ) & (~\new_[29420]_  | ~\s8_data_i[8] );
  assign \new_[25475]_  = ~\new_[30616]_  & ~\new_[29935]_ ;
  assign \new_[25476]_  = (~\new_[29705]_  | ~\s10_data_i[25] ) & (~\new_[30354]_  | ~\s9_data_i[25] );
  assign \new_[25477]_  = (~\new_[29012]_  | ~\s10_data_i[10] ) & (~\new_[29185]_  | ~\s9_data_i[10] );
  assign \new_[25478]_  = (~\new_[30227]_  | ~\s10_data_i[7] ) & (~\new_[29706]_  | ~\s9_data_i[7] );
  assign \new_[25479]_  = (~\new_[29628]_  | ~\s4_data_i[16] ) & (~\new_[29258]_  | ~\s0_data_i[16] );
  assign \new_[25480]_  = (~\s14_data_i[16]  | ~\new_[30026]_ ) & (~\s12_data_i[16]  | ~\new_[29711]_ );
  assign \new_[25481]_  = (~\new_[29036]_  | ~\s5_data_i[14] ) & (~\new_[30429]_  | ~\s3_data_i[14] );
  assign \new_[25482]_  = (~\new_[29149]_  | ~\s4_data_i[6] ) & (~\new_[29651]_  | ~\s0_data_i[6] );
  assign \new_[25483]_  = ~\new_[28762]_  | ~\new_[5925]_ ;
  assign \new_[25484]_  = ~\new_[27152]_ ;
  assign \new_[25485]_  = (~\s5_data_i[9]  | ~\new_[29649]_ ) & (~\s3_data_i[9]  | ~\new_[29035]_ );
  assign \new_[25486]_  = (~\new_[30031]_  | ~\s7_data_i[12] ) & (~\new_[29052]_  | ~\s6_data_i[12] );
  assign \new_[25487]_  = ~\new_[27155]_ ;
  assign \new_[25488]_  = ~\new_[26844]_ ;
  assign \new_[25489]_  = (~\new_[29710]_  | ~\s10_data_i[6] ) & (~\new_[29024]_  | ~\s9_data_i[6] );
  assign \new_[25490]_  = (~\new_[30284]_  | ~\s11_data_i[5] ) & (~\new_[29420]_  | ~\s8_data_i[5] );
  assign \new_[25491]_  = (~\new_[29631]_  | ~\s14_data_i[5] ) & (~\new_[29621]_  | ~\s12_data_i[5] );
  assign \new_[25492]_  = (~\s10_data_i[0]  | ~\new_[29749]_ ) & (~\s9_data_i[0]  | ~\new_[29034]_ );
  assign \new_[25493]_  = (~\new_[29641]_  | ~\s14_data_i[11] ) & (~\new_[29317]_  | ~\s12_data_i[11] );
  assign \new_[25494]_  = ~\new_[27062]_ ;
  assign \new_[25495]_  = (~\s5_data_i[24]  | ~\new_[29649]_ ) & (~\s3_data_i[24]  | ~\new_[29035]_ );
  assign \new_[25496]_  = (~\s10_data_i[24]  | ~\new_[29749]_ ) & (~\s9_data_i[24]  | ~\new_[29034]_ );
  assign \new_[25497]_  = (~\new_[29149]_  | ~\s4_data_i[4] ) & (~\new_[29651]_  | ~\s0_data_i[4] );
  assign \new_[25498]_  = (~\new_[29953]_  | ~\s11_data_i[11] ) & (~\new_[29627]_  | ~\s8_data_i[11] );
  assign \new_[25499]_  = (~\new_[30200]_  | ~\s11_data_i[24] ) & (~\new_[29428]_  | ~\s8_data_i[24] );
  assign \new_[25500]_  = (~\new_[29012]_  | ~\s10_data_i[29] ) & (~\new_[29185]_  | ~\s9_data_i[29] );
  assign \new_[25501]_  = (~\new_[29021]_  | ~\s10_data_i[4] ) & (~\new_[29709]_  | ~\s9_data_i[4] );
  assign \new_[25502]_  = (~\new_[30311]_  | ~\s11_data_i[17] ) & (~\new_[29636]_  | ~\s8_data_i[17] );
  assign \new_[25503]_  = (~\new_[29149]_  | ~\s4_data_i[2] ) & (~\new_[29651]_  | ~\s0_data_i[2] );
  assign \new_[25504]_  = (~\new_[29710]_  | ~\s10_data_i[13] ) & (~\new_[29024]_  | ~\s9_data_i[13] );
  assign \new_[25505]_  = ~\new_[29851]_  | ~\new_[28052]_ ;
  assign \new_[25506]_  = (~\new_[29641]_  | ~\s14_data_i[28] ) & (~\new_[29317]_  | ~\s12_data_i[28] );
  assign \new_[25507]_  = (~\new_[29631]_  | ~\s14_data_i[3] ) & (~\new_[29621]_  | ~\s12_data_i[3] );
  assign \new_[25508]_  = ~\new_[30269]_  & ~\new_[29915]_ ;
  assign \new_[25509]_  = \new_[28463]_  | \new_[30566]_ ;
  assign \new_[25510]_  = (~\new_[29534]_  | ~\s5_data_i[18] ) & (~\new_[29579]_  | ~\s3_data_i[18] );
  assign \new_[25511]_  = (~\new_[29705]_  | ~\s10_data_i[8] ) & (~\new_[30354]_  | ~\s9_data_i[8] );
  assign \new_[25512]_  = (~\new_[30193]_  | ~\s7_data_i[3] ) & (~\new_[29298]_  | ~\s6_data_i[3] );
  assign \new_[25513]_  = (~\new_[30193]_  | ~\s7_data_i[9] ) & (~\new_[29298]_  | ~\s6_data_i[9] );
  assign \new_[25514]_  = (~\new_[29631]_  | ~\s14_data_i[2] ) & (~\new_[29621]_  | ~\s12_data_i[2] );
  assign \new_[25515]_  = (~\new_[30031]_  | ~\s7_data_i[8] ) & (~\new_[29052]_  | ~\s6_data_i[8] );
  assign \new_[25516]_  = (~\new_[29534]_  | ~\s5_data_i[25] ) & (~\new_[29579]_  | ~\s3_data_i[25] );
  assign \new_[25517]_  = (~\new_[30284]_  | ~\s11_data_i[1] ) & (~\new_[29420]_  | ~\s8_data_i[1] );
  assign \new_[25518]_  = (~\new_[30260]_  | ~\s11_data_i[17] ) & (~\new_[29670]_  | ~\s8_data_i[17] );
  assign \new_[25519]_  = (~\new_[29036]_  | ~\s5_data_i[1] ) & (~\new_[30429]_  | ~\s3_data_i[1] );
  assign \new_[25520]_  = (~\s10_data_i[13]  | ~\new_[29749]_ ) & (~\s9_data_i[13]  | ~\new_[29034]_ );
  assign \new_[25521]_  = (~\s4_data_i[25]  | ~\new_[30335]_ ) & (~\s0_data_i[25]  | ~\new_[29603]_ );
  assign \new_[25522]_  = (~\s10_data_i[3]  | ~\new_[29749]_ ) & (~\s9_data_i[3]  | ~\new_[29034]_ );
  assign \new_[25523]_  = (~\new_[28842]_  | ~\s4_data_i[29] ) & (~\new_[29434]_  | ~\s0_data_i[29] );
  assign \new_[25524]_  = (~\new_[29012]_  | ~\s10_data_i[20] ) & (~\new_[29185]_  | ~\s9_data_i[20] );
  assign \new_[25525]_  = (~\new_[29021]_  | ~\s10_data_i[9] ) & (~\new_[29709]_  | ~\s9_data_i[9] );
  assign \new_[25526]_  = (~\new_[30260]_  | ~\s11_data_i[9] ) & (~\new_[29670]_  | ~\s8_data_i[9] );
  assign \new_[25527]_  = (~\new_[29705]_  | ~\s10_data_i[17] ) & (~\new_[30354]_  | ~\s9_data_i[17] );
  assign \new_[25528]_  = (~\new_[29953]_  | ~\s11_data_i[13] ) & (~\new_[29627]_  | ~\s8_data_i[13] );
  assign \new_[25529]_  = (~\new_[29710]_  | ~\s10_data_i[24] ) & (~\new_[29024]_  | ~\s9_data_i[24] );
  assign \new_[25530]_  = (~\new_[29953]_  | ~\s11_data_i[25] ) & (~\new_[29627]_  | ~\s8_data_i[25] );
  assign \new_[25531]_  = (~\s5_data_i[30]  | ~\new_[29649]_ ) & (~\s3_data_i[30]  | ~\new_[29035]_ );
  assign \new_[25532]_  = (~\new_[29534]_  | ~\s5_data_i[16] ) & (~\new_[29579]_  | ~\s3_data_i[16] );
  assign \new_[25533]_  = (~\new_[29641]_  | ~\s14_data_i[14] ) & (~\new_[29317]_  | ~\s12_data_i[14] );
  assign \new_[25534]_  = (~\new_[29045]_  | ~\s10_data_i[16] ) & (~\new_[29951]_  | ~\s9_data_i[16] );
  assign \new_[25535]_  = (~\s4_data_i[30]  | ~\new_[30335]_ ) & (~\s0_data_i[30]  | ~\new_[29603]_ );
  assign \new_[25536]_  = (~\new_[29953]_  | ~\s11_data_i[14] ) & (~\new_[29627]_  | ~\s8_data_i[14] );
  assign \new_[25537]_  = (~\new_[29534]_  | ~\s5_data_i[31] ) & (~\new_[29579]_  | ~\s3_data_i[31] );
  assign \new_[25538]_  = (~\new_[29025]_  | ~\s5_data_i[29] ) & (~\new_[30469]_  | ~\s3_data_i[29] );
  assign \new_[25539]_  = (~\new_[30060]_  | ~\s7_data_i[18] ) & (~\new_[29704]_  | ~\s6_data_i[18] );
  assign \new_[25540]_  = (~\new_[29534]_  | ~\s5_data_i[30] ) & (~\new_[29579]_  | ~\s3_data_i[30] );
  assign \new_[25541]_  = (~\new_[30200]_  | ~\s11_data_i[30] ) & (~\new_[29428]_  | ~\s8_data_i[30] );
  assign \new_[25542]_  = (~\new_[30193]_  | ~\s7_data_i[19] ) & (~\new_[29298]_  | ~\s6_data_i[19] );
  assign \new_[25543]_  = (~\new_[29631]_  | ~\s14_data_i[16] ) & (~\new_[29621]_  | ~\s12_data_i[16] );
  assign \new_[25544]_  = ~\new_[27181]_ ;
  assign \new_[25545]_  = (~\new_[29628]_  | ~\s4_data_i[18] ) & (~\new_[29258]_  | ~\s0_data_i[18] );
  assign \new_[25546]_  = (~\new_[29025]_  | ~\s5_data_i[10] ) & (~\new_[30469]_  | ~\s3_data_i[10] );
  assign \new_[25547]_  = (~\s5_data_i[26]  | ~\new_[29649]_ ) & (~\s3_data_i[26]  | ~\new_[29035]_ );
  assign \new_[25548]_  = (~\new_[29705]_  | ~\s10_data_i[22] ) & (~\new_[30354]_  | ~\s9_data_i[22] );
  assign \new_[25549]_  = (~\new_[30260]_  | ~\s11_data_i[10] ) & (~\new_[29670]_  | ~\s8_data_i[10] );
  assign \new_[25550]_  = ~\new_[29997]_  | ~\new_[30099]_ ;
  assign \new_[25551]_  = (~\new_[29021]_  | ~\s10_data_i[10] ) & (~\new_[29709]_  | ~\s9_data_i[10] );
  assign \new_[25552]_  = (~\s2_data_i[7]  | ~\new_[29625]_ ) & (~\s1_data_i[7]  | ~\new_[29215]_ );
  assign \new_[25553]_  = (~\new_[30284]_  | ~\s11_data_i[16] ) & (~\new_[29420]_  | ~\s8_data_i[16] );
  assign \new_[25554]_  = (~\new_[29534]_  | ~\s5_data_i[27] ) & (~\new_[29579]_  | ~\s3_data_i[27] );
  assign \new_[25555]_  = (~\new_[30311]_  | ~\s11_data_i[19] ) & (~\new_[29636]_  | ~\s8_data_i[19] );
  assign \new_[25556]_  = (~\new_[30031]_  | ~\s7_data_i[17] ) & (~\new_[29052]_  | ~\s6_data_i[17] );
  assign \new_[25557]_  = (~\new_[30193]_  | ~\s7_data_i[10] ) & (~\new_[29298]_  | ~\s6_data_i[10] );
  assign \new_[25558]_  = ~\new_[27188]_ ;
  assign \new_[25559]_  = (~\new_[30200]_  | ~\s11_data_i[3] ) & (~\new_[29428]_  | ~\s8_data_i[3] );
  assign \new_[25560]_  = ~\new_[27947]_ ;
  assign \new_[25561]_  = (~\s5_data_i[29]  | ~\new_[29649]_ ) & (~\s3_data_i[29]  | ~\new_[29035]_ );
  assign \new_[25562]_  = (~\new_[29534]_  | ~\s5_data_i[24] ) & (~\new_[29579]_  | ~\s3_data_i[24] );
  assign \new_[25563]_  = (~\new_[29149]_  | ~\s4_data_i[16] ) & (~\new_[29651]_  | ~\s0_data_i[16] );
  assign \new_[25564]_  = ~\new_[27196]_ ;
  assign \new_[25565]_  = (~\new_[29705]_  | ~\s10_data_i[30] ) & (~\new_[30354]_  | ~\s9_data_i[30] );
  assign \new_[25566]_  = (~\new_[29021]_  | ~\s10_data_i[22] ) & (~\new_[29709]_  | ~\s9_data_i[22] );
  assign \new_[25567]_  = (~\s2_data_i[25]  | ~\new_[29625]_ ) & (~\s1_data_i[25]  | ~\new_[29215]_ );
  assign \new_[25568]_  = (~\new_[29534]_  | ~\s5_data_i[3] ) & (~\new_[29579]_  | ~\s3_data_i[3] );
  assign \new_[25569]_  = (~\new_[30060]_  | ~\s7_data_i[19] ) & (~\new_[29704]_  | ~\s6_data_i[19] );
  assign \new_[25570]_  = (~\new_[29045]_  | ~\s10_data_i[7] ) & (~\new_[29951]_  | ~\s9_data_i[7] );
  assign \new_[25571]_  = ~\new_[26820]_ ;
  assign \new_[25572]_  = (~\new_[29534]_  | ~\s5_data_i[21] ) & (~\new_[29579]_  | ~\s3_data_i[21] );
  assign \new_[25573]_  = ~\new_[27198]_ ;
  assign \new_[25574]_  = (~\new_[29628]_  | ~\s4_data_i[19] ) & (~\new_[29258]_  | ~\s0_data_i[19] );
  assign \new_[25575]_  = (~\new_[30227]_  | ~\s10_data_i[20] ) & (~\new_[29706]_  | ~\s9_data_i[20] );
  assign \new_[25576]_  = (~\s2_data_i[12]  | ~\new_[29625]_ ) & (~\s1_data_i[12]  | ~\new_[29215]_ );
  assign \new_[25577]_  = (~\new_[29628]_  | ~\s4_data_i[31] ) & (~\new_[29258]_  | ~\s0_data_i[31] );
  assign \new_[25578]_  = (~\new_[30200]_  | ~\s11_data_i[31] ) & (~\new_[29428]_  | ~\s8_data_i[31] );
  assign \new_[25579]_  = (~\s2_data_i[11]  | ~\new_[29625]_ ) & (~\s1_data_i[11]  | ~\new_[29215]_ );
  assign \new_[25580]_  = ~\new_[27206]_ ;
  assign \new_[25581]_  = (~\new_[29534]_  | ~\s5_data_i[17] ) & (~\new_[29579]_  | ~\s3_data_i[17] );
  assign \new_[25582]_  = (~\new_[30181]_  | ~\s14_data_i[20] ) & (~\new_[29640]_  | ~\s12_data_i[20] );
  assign \new_[25583]_  = (~\new_[29705]_  | ~\s10_data_i[11] ) & (~\new_[30354]_  | ~\s9_data_i[11] );
  assign \new_[25584]_  = (~\new_[30193]_  | ~\s7_data_i[6] ) & (~\new_[29298]_  | ~\s6_data_i[6] );
  assign \new_[25585]_  = (~\new_[29036]_  | ~\s5_data_i[6] ) & (~\new_[30429]_  | ~\s3_data_i[6] );
  assign \new_[25586]_  = (~\new_[29025]_  | ~\s5_data_i[23] ) & (~\new_[30469]_  | ~\s3_data_i[23] );
  assign \new_[25587]_  = (~\s4_data_i[11]  | ~\new_[30335]_ ) & (~\s0_data_i[11]  | ~\new_[29603]_ );
  assign \new_[25588]_  = (~\new_[29045]_  | ~\s10_data_i[20] ) & (~\new_[29951]_  | ~\s9_data_i[20] );
  assign \new_[25589]_  = (~\new_[30031]_  | ~\s7_data_i[13] ) & (~\new_[29052]_  | ~\s6_data_i[13] );
  assign \new_[25590]_  = ~\new_[28083]_  | ~\new_[6090]_ ;
  assign \new_[25591]_  = (~\new_[29036]_  | ~\s5_data_i[5] ) & (~\new_[30429]_  | ~\s3_data_i[5] );
  assign \new_[25592]_  = (~\new_[30200]_  | ~\s11_data_i[28] ) & (~\new_[29428]_  | ~\s8_data_i[28] );
  assign \new_[25593]_  = (~\new_[29749]_  | ~\s10_data_i[31] ) & (~\new_[29034]_  | ~\s9_data_i[31] );
  assign \new_[25594]_  = (~\new_[29012]_  | ~\s10_data_i[31] ) & (~\new_[29185]_  | ~\s9_data_i[31] );
  assign \new_[25595]_  = (~\new_[29021]_  | ~\s10_data_i[11] ) & (~\new_[29709]_  | ~\s9_data_i[11] );
  assign \new_[25596]_  = ~\new_[27224]_ ;
  assign \new_[25597]_  = (~\new_[29710]_  | ~\s10_data_i[27] ) & (~\new_[29024]_  | ~\s9_data_i[27] );
  assign \new_[25598]_  = ~\new_[30000]_  | ~\new_[30550]_ ;
  assign \new_[25599]_  = (~\new_[29012]_  | ~\s10_data_i[25] ) & (~\new_[29185]_  | ~\s9_data_i[25] );
  assign \new_[25600]_  = (~\new_[30260]_  | ~\s11_data_i[12] ) & (~\new_[29670]_  | ~\s8_data_i[12] );
  assign \new_[25601]_  = (~\new_[30031]_  | ~\s7_data_i[21] ) & (~\new_[29052]_  | ~\s6_data_i[21] );
  assign \new_[25602]_  = ~\new_[29767]_  & ~\new_[29888]_ ;
  assign \new_[25603]_  = (~\new_[29534]_  | ~\s5_data_i[10] ) & (~\new_[29579]_  | ~\s3_data_i[10] );
  assign \new_[25604]_  = (~\new_[29710]_  | ~\s10_data_i[26] ) & (~\new_[29024]_  | ~\s9_data_i[26] );
  assign \new_[25605]_  = (~\s11_data_i[11]  | ~\new_[29205]_ ) & (~\s8_data_i[11]  | ~\new_[29241]_ );
  assign \new_[25606]_  = (~\new_[30200]_  | ~\s11_data_i[26] ) & (~\new_[29428]_  | ~\s8_data_i[26] );
  assign \new_[25607]_  = ~\new_[26770]_ ;
  assign \new_[25608]_  = (~\new_[29036]_  | ~\s5_data_i[8] ) & (~\new_[30429]_  | ~\s3_data_i[8] );
  assign \new_[25609]_  = (~\new_[29710]_  | ~\s10_data_i[25] ) & (~\new_[29024]_  | ~\s9_data_i[25] );
  assign \new_[25610]_  = (~\new_[29953]_  | ~\s11_data_i[22] ) & (~\new_[29627]_  | ~\s8_data_i[22] );
  assign \new_[25611]_  = (~\new_[30200]_  | ~\s11_data_i[10] ) & (~\new_[29428]_  | ~\s8_data_i[10] );
  assign \new_[25612]_  = (~\new_[30200]_  | ~\s11_data_i[25] ) & (~\new_[29428]_  | ~\s8_data_i[25] );
  assign \new_[25613]_  = (~\new_[29641]_  | ~\s14_data_i[25] ) & (~\new_[29317]_  | ~\s12_data_i[25] );
  assign \new_[25614]_  = (~\new_[28842]_  | ~\s4_data_i[12] ) & (~\new_[29434]_  | ~\s0_data_i[12] );
  assign \new_[25615]_  = (~\new_[29534]_  | ~\s5_data_i[8] ) & (~\new_[29579]_  | ~\s3_data_i[8] );
  assign \new_[25616]_  = (~\new_[29641]_  | ~\s14_data_i[29] ) & (~\new_[29317]_  | ~\s12_data_i[29] );
  assign \new_[25617]_  = (~\new_[29953]_  | ~\s11_data_i[20] ) & (~\new_[29627]_  | ~\s8_data_i[20] );
  assign \new_[25618]_  = (~\new_[29628]_  | ~\s4_data_i[6] ) & (~\new_[29258]_  | ~\s0_data_i[6] );
  assign \new_[25619]_  = (~\new_[30200]_  | ~\s11_data_i[4] ) & (~\new_[29428]_  | ~\s8_data_i[4] );
  assign \new_[25620]_  = (~\s14_data_i[11]  | ~\new_[30026]_ ) & (~\s12_data_i[11]  | ~\new_[29711]_ );
  assign \new_[25621]_  = ~\new_[30542]_  | ~\new_[31712]_ ;
  assign \new_[25622]_  = (~\s2_data_i[22]  | ~\new_[29625]_ ) & (~\s1_data_i[22]  | ~\new_[29215]_ );
  assign \new_[25623]_  = (~\new_[29045]_  | ~\s10_data_i[21] ) & (~\new_[29951]_  | ~\s9_data_i[21] );
  assign \new_[25624]_  = (~\new_[29710]_  | ~\s10_data_i[23] ) & (~\new_[29024]_  | ~\s9_data_i[23] );
  assign \new_[25625]_  = (~\new_[30200]_  | ~\s11_data_i[23] ) & (~\new_[29428]_  | ~\s8_data_i[23] );
  assign \new_[25626]_  = (~\new_[30200]_  | ~\s11_data_i[5] ) & (~\new_[29428]_  | ~\s8_data_i[5] );
  assign \new_[25627]_  = ~\new_[27246]_ ;
  assign \new_[25628]_  = (~\new_[30227]_  | ~\s10_data_i[19] ) & (~\new_[29706]_  | ~\s9_data_i[19] );
  assign \new_[25629]_  = (~\s4_data_i[4]  | ~\new_[30335]_ ) & (~\s0_data_i[4]  | ~\new_[29603]_ );
  assign \new_[25630]_  = (~\new_[29534]_  | ~\s5_data_i[0] ) & (~\new_[29579]_  | ~\s3_data_i[0] );
  assign \new_[25631]_  = (~\new_[29012]_  | ~\s10_data_i[26] ) & (~\new_[29185]_  | ~\s9_data_i[26] );
  assign \new_[25632]_  = (~\new_[29710]_  | ~\s10_data_i[21] ) & (~\new_[29024]_  | ~\s9_data_i[21] );
  assign \new_[25633]_  = (~\new_[28842]_  | ~\s4_data_i[31] ) & (~\new_[29434]_  | ~\s0_data_i[31] );
  assign \new_[25634]_  = (~\s2_data_i[18]  | ~\new_[29625]_ ) & (~\s1_data_i[18]  | ~\new_[29215]_ );
  assign \new_[25635]_  = (~\new_[29710]_  | ~\s10_data_i[16] ) & (~\new_[29024]_  | ~\s9_data_i[16] );
  assign \new_[25636]_  = (~\new_[30200]_  | ~\s11_data_i[11] ) & (~\new_[29428]_  | ~\s8_data_i[11] );
  assign \new_[25637]_  = (~\new_[29534]_  | ~\s5_data_i[29] ) & (~\new_[29579]_  | ~\s3_data_i[29] );
  assign \new_[25638]_  = (~\new_[29025]_  | ~\s5_data_i[14] ) & (~\new_[30469]_  | ~\s3_data_i[14] );
  assign \new_[25639]_  = (~\s5_data_i[10]  | ~\new_[29649]_ ) & (~\s3_data_i[10]  | ~\new_[29035]_ );
  assign \new_[25640]_  = \new_[30286]_  & \new_[6059]_ ;
  assign \new_[25641]_  = (~\new_[28842]_  | ~\s4_data_i[13] ) & (~\new_[29434]_  | ~\s0_data_i[13] );
  assign \new_[25642]_  = (~\s14_data_i[30]  | ~\new_[30026]_ ) & (~\s12_data_i[30]  | ~\new_[29711]_ );
  assign \new_[25643]_  = (~\new_[29631]_  | ~\s14_data_i[8] ) & (~\new_[29621]_  | ~\s12_data_i[8] );
  assign \new_[25644]_  = (~\new_[30260]_  | ~\s11_data_i[14] ) & (~\new_[29670]_  | ~\s8_data_i[14] );
  assign \new_[25645]_  = (~\new_[29205]_  | ~\s11_data_i[31] ) & (~\new_[29241]_  | ~\s8_data_i[31] );
  assign \new_[25646]_  = (~\s5_data_i[0]  | ~\new_[29649]_ ) & (~\s3_data_i[0]  | ~\new_[29035]_ );
  assign \new_[25647]_  = (~\new_[29534]_  | ~\s5_data_i[9] ) & (~\new_[29579]_  | ~\s3_data_i[9] );
  assign \new_[25648]_  = (~\new_[29625]_  | ~\s2_data_i[31] ) & (~\new_[29215]_  | ~\s1_data_i[31] );
  assign \new_[25649]_  = (~\s2_data_i[10]  | ~\new_[29625]_ ) & (~\s1_data_i[10]  | ~\new_[29215]_ );
  assign \new_[25650]_  = (~\new_[29705]_  | ~\s10_data_i[16] ) & (~\new_[30354]_  | ~\s9_data_i[16] );
  assign \new_[25651]_  = (~\new_[29149]_  | ~\s4_data_i[20] ) & (~\new_[29651]_  | ~\s0_data_i[20] );
  assign \new_[25652]_  = (~\new_[30060]_  | ~\s7_data_i[30] ) & (~\new_[29704]_  | ~\s6_data_i[30] );
  assign \new_[25653]_  = (~\new_[29534]_  | ~\s5_data_i[4] ) & (~\new_[29579]_  | ~\s3_data_i[4] );
  assign \new_[25654]_  = (~\new_[30181]_  | ~\s14_data_i[23] ) & (~\new_[29640]_  | ~\s12_data_i[23] );
  assign \new_[25655]_  = (~\new_[29036]_  | ~\s5_data_i[21] ) & (~\new_[30429]_  | ~\s3_data_i[21] );
  assign \new_[25656]_  = (~\new_[29641]_  | ~\s14_data_i[23] ) & (~\new_[29317]_  | ~\s12_data_i[23] );
  assign \new_[25657]_  = (~\new_[30311]_  | ~\s11_data_i[23] ) & (~\new_[29636]_  | ~\s8_data_i[23] );
  assign \new_[25658]_  = ~\new_[28358]_  | ~\new_[6065]_ ;
  assign \new_[25659]_  = (~\new_[29036]_  | ~\s5_data_i[12] ) & (~\new_[30429]_  | ~\s3_data_i[12] );
  assign \new_[25660]_  = ~\new_[27290]_ ;
  assign \new_[25661]_  = (~\s2_data_i[23]  | ~\new_[29625]_ ) & (~\s1_data_i[23]  | ~\new_[29215]_ );
  assign \new_[25662]_  = (~\new_[29953]_  | ~\s11_data_i[29] ) & (~\new_[29627]_  | ~\s8_data_i[29] );
  assign \new_[25663]_  = (~\s4_data_i[29]  | ~\new_[30335]_ ) & (~\s0_data_i[29]  | ~\new_[29603]_ );
  assign \new_[25664]_  = (~\new_[30284]_  | ~\s11_data_i[21] ) & (~\new_[29420]_  | ~\s8_data_i[21] );
  assign \new_[25665]_  = (~\new_[29631]_  | ~\s14_data_i[21] ) & (~\new_[29621]_  | ~\s12_data_i[21] );
  assign \new_[25666]_  = (~\new_[29710]_  | ~\s10_data_i[18] ) & (~\new_[29024]_  | ~\s9_data_i[18] );
  assign \new_[25667]_  = (~\s2_data_i[15]  | ~\new_[29625]_ ) & (~\s1_data_i[15]  | ~\new_[29215]_ );
  assign \new_[25668]_  = (~\new_[29705]_  | ~\s10_data_i[26] ) & (~\new_[30354]_  | ~\s9_data_i[26] );
  assign \new_[25669]_  = (~\new_[29953]_  | ~\s11_data_i[23] ) & (~\new_[29627]_  | ~\s8_data_i[23] );
  assign \new_[25670]_  = ~\new_[26678]_ ;
  assign \new_[25671]_  = (~\new_[30060]_  | ~\s7_data_i[23] ) & (~\new_[29704]_  | ~\s6_data_i[23] );
  assign \new_[25672]_  = (~\new_[29705]_  | ~\s10_data_i[29] ) & (~\new_[30354]_  | ~\s9_data_i[29] );
  assign \new_[25673]_  = (~\s2_data_i[5]  | ~\new_[29625]_ ) & (~\s1_data_i[5]  | ~\new_[29215]_ );
  assign \new_[25674]_  = ~\new_[29623]_  & ~\new_[30059]_ ;
  assign \new_[25675]_  = ~\new_[26625]_ ;
  assign \new_[25676]_  = ~\new_[26622]_ ;
  assign \new_[25677]_  = (~\new_[29012]_  | ~\s10_data_i[24] ) & (~\new_[29185]_  | ~\s9_data_i[24] );
  assign \new_[25678]_  = (~\new_[29025]_  | ~\s5_data_i[15] ) & (~\new_[30469]_  | ~\s3_data_i[15] );
  assign \new_[25679]_  = (~\new_[30284]_  | ~\s11_data_i[22] ) & (~\new_[29420]_  | ~\s8_data_i[22] );
  assign \new_[25680]_  = (~\new_[30200]_  | ~\s11_data_i[12] ) & (~\new_[29428]_  | ~\s8_data_i[12] );
  assign \new_[25681]_  = (~\new_[30311]_  | ~\s11_data_i[24] ) & (~\new_[29636]_  | ~\s8_data_i[24] );
  assign \new_[25682]_  = (~\new_[29021]_  | ~\s10_data_i[13] ) & (~\new_[29709]_  | ~\s9_data_i[13] );
  assign \new_[25683]_  = (~\new_[30311]_  | ~\s11_data_i[21] ) & (~\new_[29636]_  | ~\s8_data_i[21] );
  assign \new_[25684]_  = (~\new_[30200]_  | ~\s11_data_i[13] ) & (~\new_[29428]_  | ~\s8_data_i[13] );
  assign \new_[25685]_  = (~\new_[30227]_  | ~\s10_data_i[22] ) & (~\new_[29706]_  | ~\s9_data_i[22] );
  assign \new_[25686]_  = (~\new_[29036]_  | ~\s5_data_i[0] ) & (~\new_[30429]_  | ~\s3_data_i[0] );
  assign \new_[25687]_  = ~\new_[26577]_ ;
  assign \new_[25688]_  = (~\new_[29710]_  | ~\s10_data_i[12] ) & (~\new_[29024]_  | ~\s9_data_i[12] );
  assign \new_[25689]_  = (~\new_[29045]_  | ~\s10_data_i[24] ) & (~\new_[29951]_  | ~\s9_data_i[24] );
  assign \new_[25690]_  = (~\new_[28842]_  | ~\s4_data_i[27] ) & (~\new_[29434]_  | ~\s0_data_i[27] );
  assign \new_[25691]_  = ~\new_[27277]_ ;
  assign \new_[25692]_  = (~\new_[30031]_  | ~\s7_data_i[27] ) & (~\new_[29052]_  | ~\s6_data_i[27] );
  assign \new_[25693]_  = (~\new_[29021]_  | ~\s10_data_i[17] ) & (~\new_[29709]_  | ~\s9_data_i[17] );
  assign \new_[25694]_  = (~\new_[30311]_  | ~\s11_data_i[4] ) & (~\new_[29636]_  | ~\s8_data_i[4] );
  assign \new_[25695]_  = ~\new_[27968]_ ;
  assign \new_[25696]_  = (~\s11_data_i[0]  | ~\new_[29205]_ ) & (~\s8_data_i[0]  | ~\new_[29241]_ );
  assign \new_[25697]_  = (~\new_[29631]_  | ~\s14_data_i[23] ) & (~\new_[29621]_  | ~\s12_data_i[23] );
  assign \new_[25698]_  = (~\s5_data_i[12]  | ~\new_[29649]_ ) & (~\s3_data_i[12]  | ~\new_[29035]_ );
  assign \new_[25699]_  = (~\new_[29021]_  | ~\s10_data_i[2] ) & (~\new_[29709]_  | ~\s9_data_i[2] );
  assign \new_[25700]_  = (~\new_[29953]_  | ~\s11_data_i[31] ) & (~\new_[29627]_  | ~\s8_data_i[31] );
  assign \new_[25701]_  = (~\s11_data_i[12]  | ~\new_[29205]_ ) & (~\s8_data_i[12]  | ~\new_[29241]_ );
  assign \new_[25702]_  = (~\new_[29036]_  | ~\s5_data_i[30] ) & (~\new_[30429]_  | ~\s3_data_i[30] );
  assign \new_[25703]_  = (~\new_[29036]_  | ~\s5_data_i[23] ) & (~\new_[30429]_  | ~\s3_data_i[23] );
  assign \new_[25704]_  = (~\s2_data_i[8]  | ~\new_[29625]_ ) & (~\s1_data_i[8]  | ~\new_[29215]_ );
  assign \new_[25705]_  = (~\new_[30193]_  | ~\s7_data_i[2] ) & (~\new_[29298]_  | ~\s6_data_i[2] );
  assign \new_[25706]_  = (~\new_[29976]_  | ~\s14_data_i[19] ) & (~\new_[28957]_  | ~\s12_data_i[19] );
  assign \new_[25707]_  = (~\new_[28842]_  | ~\s4_data_i[17] ) & (~\new_[29434]_  | ~\s0_data_i[17] );
  assign \new_[25708]_  = ~\new_[27267]_ ;
  assign \new_[25709]_  = (~\s2_data_i[14]  | ~\new_[29625]_ ) & (~\s1_data_i[14]  | ~\new_[29215]_ );
  assign \new_[25710]_  = (~\s11_data_i[24]  | ~\new_[29205]_ ) & (~\s8_data_i[24]  | ~\new_[29241]_ );
  assign \new_[25711]_  = ~\new_[30006]_  | ~\new_[5902]_ ;
  assign \new_[25712]_  = (~\new_[30031]_  | ~\s7_data_i[25] ) & (~\new_[29052]_  | ~\s6_data_i[25] );
  assign \new_[25713]_  = (~\new_[29036]_  | ~\s5_data_i[24] ) & (~\new_[30429]_  | ~\s3_data_i[24] );
  assign \new_[25714]_  = (~\s11_data_i[6]  | ~\new_[29205]_ ) & (~\s8_data_i[6]  | ~\new_[29241]_ );
  assign \new_[25715]_  = ~\new_[30038]_  | ~\new_[28057]_ ;
  assign \new_[25716]_  = (~\s4_data_i[21]  | ~\new_[30335]_ ) & (~\s0_data_i[21]  | ~\new_[29603]_ );
  assign \new_[25717]_  = (~\new_[29710]_  | ~\s10_data_i[9] ) & (~\new_[29024]_  | ~\s9_data_i[9] );
  assign \new_[25718]_  = (~\s5_data_i[11]  | ~\new_[29649]_ ) & (~\s3_data_i[11]  | ~\new_[29035]_ );
  assign \new_[25719]_  = (~\new_[29641]_  | ~\s14_data_i[27] ) & (~\new_[29317]_  | ~\s12_data_i[27] );
  assign \new_[25720]_  = (~\new_[30284]_  | ~\s11_data_i[24] ) & (~\new_[29420]_  | ~\s8_data_i[24] );
  assign \new_[25721]_  = (~\new_[30060]_  | ~\s7_data_i[29] ) & (~\new_[29704]_  | ~\s6_data_i[29] );
  assign \new_[25722]_  = (~\new_[30260]_  | ~\s11_data_i[25] ) & (~\new_[29670]_  | ~\s8_data_i[25] );
  assign \new_[25723]_  = (~\s4_data_i[26]  | ~\new_[30335]_ ) & (~\s0_data_i[26]  | ~\new_[29603]_ );
  assign \new_[25724]_  = (~\new_[29976]_  | ~\s14_data_i[25] ) & (~\new_[28957]_  | ~\s12_data_i[25] );
  assign \new_[25725]_  = (~\new_[29149]_  | ~\s4_data_i[29] ) & (~\new_[29651]_  | ~\s0_data_i[29] );
  assign \new_[25726]_  = (~\new_[30181]_  | ~\s14_data_i[7] ) & (~\new_[29640]_  | ~\s12_data_i[7] );
  assign \new_[25727]_  = (~\new_[30227]_  | ~\s10_data_i[24] ) & (~\new_[29706]_  | ~\s9_data_i[24] );
  assign \new_[25728]_  = ~\new_[27302]_ ;
  assign \new_[25729]_  = (~\new_[29710]_  | ~\s10_data_i[8] ) & (~\new_[29024]_  | ~\s9_data_i[8] );
  assign \new_[25730]_  = (~\new_[29534]_  | ~\s5_data_i[15] ) & (~\new_[29579]_  | ~\s3_data_i[15] );
  assign \new_[25731]_  = (~\new_[30227]_  | ~\s10_data_i[5] ) & (~\new_[29706]_  | ~\s9_data_i[5] );
  assign \new_[25732]_  = (~\s2_data_i[24]  | ~\new_[29625]_ ) & (~\s1_data_i[24]  | ~\new_[29215]_ );
  assign \new_[25733]_  = (~\new_[30311]_  | ~\s11_data_i[26] ) & (~\new_[29636]_  | ~\s8_data_i[26] );
  assign \new_[25734]_  = (~\new_[30260]_  | ~\s11_data_i[31] ) & (~\new_[29670]_  | ~\s8_data_i[31] );
  assign \new_[25735]_  = ~\new_[27793]_ ;
  assign \new_[25736]_  = (~\new_[29705]_  | ~\s10_data_i[27] ) & (~\new_[30354]_  | ~\s9_data_i[27] );
  assign \new_[25737]_  = (~\new_[29036]_  | ~\s5_data_i[29] ) & (~\new_[30429]_  | ~\s3_data_i[29] );
  assign \new_[25738]_  = (~\new_[29641]_  | ~\s14_data_i[24] ) & (~\new_[29317]_  | ~\s12_data_i[24] );
  assign \new_[25739]_  = (~\new_[30227]_  | ~\s10_data_i[25] ) & (~\new_[29706]_  | ~\s9_data_i[25] );
  assign \new_[25740]_  = (~\new_[29534]_  | ~\s5_data_i[28] ) & (~\new_[29579]_  | ~\s3_data_i[28] );
  assign \new_[25741]_  = (~\new_[29628]_  | ~\s4_data_i[26] ) & (~\new_[29258]_  | ~\s0_data_i[26] );
  assign \new_[25742]_  = (~\s10_data_i[11]  | ~\new_[29749]_ ) & (~\s9_data_i[11]  | ~\new_[29034]_ );
  assign \new_[25743]_  = (~\new_[29710]_  | ~\s10_data_i[22] ) & (~\new_[29024]_  | ~\s9_data_i[22] );
  assign \new_[25744]_  = (~\s4_data_i[7]  | ~\new_[30335]_ ) & (~\s0_data_i[7]  | ~\new_[29603]_ );
  assign \new_[25745]_  = (~\s5_data_i[15]  | ~\new_[29649]_ ) & (~\s3_data_i[15]  | ~\new_[29035]_ );
  assign \new_[25746]_  = (~\new_[28842]_  | ~\s4_data_i[22] ) & (~\new_[29434]_  | ~\s0_data_i[22] );
  assign \new_[25747]_  = (~\s5_data_i[6]  | ~\new_[29649]_ ) & (~\s3_data_i[6]  | ~\new_[29035]_ );
  assign \new_[25748]_  = (~\s4_data_i[9]  | ~\new_[30335]_ ) & (~\s0_data_i[9]  | ~\new_[29603]_ );
  assign \new_[25749]_  = (~\new_[29976]_  | ~\s14_data_i[31] ) & (~\new_[28957]_  | ~\s12_data_i[31] );
  assign \new_[25750]_  = (~\new_[30227]_  | ~\s10_data_i[26] ) & (~\new_[29706]_  | ~\s9_data_i[26] );
  assign \new_[25751]_  = (~\s11_data_i[30]  | ~\new_[29205]_ ) & (~\s8_data_i[30]  | ~\new_[29241]_ );
  assign \new_[25752]_  = (~\new_[29025]_  | ~\s5_data_i[31] ) & (~\new_[30469]_  | ~\s3_data_i[31] );
  assign \new_[25753]_  = ~\new_[27681]_ ;
  assign \new_[25754]_  = (~\s10_data_i[22]  | ~\new_[29749]_ ) & (~\s9_data_i[22]  | ~\new_[29034]_ );
  assign \new_[25755]_  = (~\new_[30260]_  | ~\s11_data_i[24] ) & (~\new_[29670]_  | ~\s8_data_i[24] );
  assign \new_[25756]_  = (~\new_[29036]_  | ~\s5_data_i[15] ) & (~\new_[30429]_  | ~\s3_data_i[15] );
  assign \new_[25757]_  = (~\new_[29036]_  | ~\s5_data_i[27] ) & (~\new_[30429]_  | ~\s3_data_i[27] );
  assign \new_[25758]_  = (~\new_[29631]_  | ~\s14_data_i[11] ) & (~\new_[29621]_  | ~\s12_data_i[11] );
  assign \new_[25759]_  = (~\new_[29628]_  | ~\s4_data_i[3] ) & (~\new_[29258]_  | ~\s0_data_i[3] );
  assign \new_[25760]_  = (~\s11_data_i[5]  | ~\new_[29205]_ ) & (~\s8_data_i[5]  | ~\new_[29241]_ );
  assign \new_[25761]_  = (~\new_[29631]_  | ~\s14_data_i[27] ) & (~\new_[29621]_  | ~\s12_data_i[27] );
  assign \new_[25762]_  = (~\new_[29149]_  | ~\s4_data_i[14] ) & (~\new_[29651]_  | ~\s0_data_i[14] );
  assign \new_[25763]_  = (~\new_[29710]_  | ~\s10_data_i[3] ) & (~\new_[29024]_  | ~\s9_data_i[3] );
  assign \new_[25764]_  = (~\new_[30031]_  | ~\s7_data_i[20] ) & (~\new_[29052]_  | ~\s6_data_i[20] );
  assign \new_[25765]_  = ~\new_[27322]_ ;
  assign \new_[25766]_  = (~\s5_data_i[25]  | ~\new_[29649]_ ) & (~\s3_data_i[25]  | ~\new_[29035]_ );
  assign \new_[25767]_  = ~\new_[28114]_  | ~\new_[5963]_ ;
  assign \new_[25768]_  = (~\new_[30200]_  | ~\s11_data_i[6] ) & (~\new_[29428]_  | ~\s8_data_i[6] );
  assign \new_[25769]_  = (~\new_[29534]_  | ~\s5_data_i[26] ) & (~\new_[29579]_  | ~\s3_data_i[26] );
  assign \new_[25770]_  = ~\new_[30038]_  & ~\new_[30697]_ ;
  assign \new_[25771]_  = ~\new_[27590]_ ;
  assign \new_[25772]_  = (~\new_[29025]_  | ~\s5_data_i[20] ) & (~\new_[30469]_  | ~\s3_data_i[20] );
  assign \new_[25773]_  = (~\new_[29149]_  | ~\s4_data_i[5] ) & (~\new_[29651]_  | ~\s0_data_i[5] );
  assign \new_[25774]_  = ~\new_[27323]_ ;
  assign \new_[25775]_  = ~\new_[30151]_  & ~\new_[30786]_ ;
  assign \new_[25776]_  = (~\new_[29534]_  | ~\s5_data_i[2] ) & (~\new_[29579]_  | ~\s3_data_i[2] );
  assign \new_[25777]_  = (~\new_[30227]_  | ~\s10_data_i[28] ) & (~\new_[29706]_  | ~\s9_data_i[28] );
  assign \new_[25778]_  = (~\new_[29149]_  | ~\s4_data_i[27] ) & (~\new_[29651]_  | ~\s0_data_i[27] );
  assign \new_[25779]_  = (~\new_[29705]_  | ~\s10_data_i[19] ) & (~\new_[30354]_  | ~\s9_data_i[19] );
  assign \new_[25780]_  = (~\new_[29534]_  | ~\s5_data_i[1] ) & (~\new_[29579]_  | ~\s3_data_i[1] );
  assign \new_[25781]_  = (~\new_[30260]_  | ~\s11_data_i[18] ) & (~\new_[29670]_  | ~\s8_data_i[18] );
  assign \new_[25782]_  = (~\new_[29036]_  | ~\s5_data_i[28] ) & (~\new_[30429]_  | ~\s3_data_i[28] );
  assign \new_[25783]_  = ~\new_[27105]_ ;
  assign \new_[25784]_  = (~\new_[29710]_  | ~\s10_data_i[5] ) & (~\new_[29024]_  | ~\s9_data_i[5] );
  assign \new_[25785]_  = (~\new_[29045]_  | ~\s10_data_i[28] ) & (~\new_[29951]_  | ~\s9_data_i[28] );
  assign \new_[25786]_  = (~\new_[30060]_  | ~\s7_data_i[3] ) & (~\new_[29704]_  | ~\s6_data_i[3] );
  assign \new_[25787]_  = (~\new_[29021]_  | ~\s10_data_i[5] ) & (~\new_[29709]_  | ~\s9_data_i[5] );
  assign \new_[25788]_  = (~\new_[29710]_  | ~\s10_data_i[28] ) & (~\new_[29024]_  | ~\s9_data_i[28] );
  assign \new_[25789]_  = (~\new_[30193]_  | ~\s7_data_i[16] ) & (~\new_[29298]_  | ~\s6_data_i[16] );
  assign \new_[25790]_  = (~\s14_data_i[13]  | ~\new_[30026]_ ) & (~\s12_data_i[13]  | ~\new_[29711]_ );
  assign \new_[25791]_  = (~\new_[29976]_  | ~\s14_data_i[23] ) & (~\new_[28957]_  | ~\s12_data_i[23] );
  assign \new_[25792]_  = (~\new_[30227]_  | ~\s10_data_i[30] ) & (~\new_[29706]_  | ~\s9_data_i[30] );
  assign \new_[25793]_  = (~\new_[30260]_  | ~\s11_data_i[20] ) & (~\new_[29670]_  | ~\s8_data_i[20] );
  assign \new_[25794]_  = (~\new_[29628]_  | ~\s4_data_i[28] ) & (~\new_[29258]_  | ~\s0_data_i[28] );
  assign \new_[25795]_  = (~\new_[30284]_  | ~\s11_data_i[17] ) & (~\new_[29420]_  | ~\s8_data_i[17] );
  assign \new_[25796]_  = (~\new_[29149]_  | ~\s4_data_i[1] ) & (~\new_[29651]_  | ~\s0_data_i[1] );
  assign \new_[25797]_  = (~\new_[30031]_  | ~\s7_data_i[19] ) & (~\new_[29052]_  | ~\s6_data_i[19] );
  assign \new_[25798]_  = (~\s11_data_i[10]  | ~\new_[29205]_ ) & (~\s8_data_i[10]  | ~\new_[29241]_ );
  assign \new_[25799]_  = (~\new_[29534]_  | ~\s5_data_i[14] ) & (~\new_[29579]_  | ~\s3_data_i[14] );
  assign \new_[25800]_  = ~\new_[27334]_ ;
  assign \new_[25801]_  = (~\new_[29641]_  | ~\s14_data_i[31] ) & (~\new_[29317]_  | ~\s12_data_i[31] );
  assign \new_[25802]_  = (~\new_[30260]_  | ~\s11_data_i[21] ) & (~\new_[29670]_  | ~\s8_data_i[21] );
  assign \new_[25803]_  = (~\new_[29149]_  | ~\s4_data_i[28] ) & (~\new_[29651]_  | ~\s0_data_i[28] );
  assign \new_[25804]_  = (~\new_[30260]_  | ~\s11_data_i[29] ) & (~\new_[29670]_  | ~\s8_data_i[29] );
  assign \new_[25805]_  = (~\new_[29021]_  | ~\s10_data_i[16] ) & (~\new_[29709]_  | ~\s9_data_i[16] );
  assign \new_[25806]_  = (~\new_[29036]_  | ~\s5_data_i[2] ) & (~\new_[30429]_  | ~\s3_data_i[2] );
  assign \new_[25807]_  = (~\s2_data_i[6]  | ~\new_[29625]_ ) & (~\s1_data_i[6]  | ~\new_[29215]_ );
  assign \new_[25808]_  = (~\new_[29976]_  | ~\s14_data_i[15] ) & (~\new_[28957]_  | ~\s12_data_i[15] );
  assign \new_[25809]_  = (~\new_[29025]_  | ~\s5_data_i[26] ) & (~\new_[30469]_  | ~\s3_data_i[26] );
  assign \new_[25810]_  = (~\new_[29710]_  | ~\s10_data_i[19] ) & (~\new_[29024]_  | ~\s9_data_i[19] );
  assign \new_[25811]_  = ~\new_[28183]_  | ~\new_[5910]_ ;
  assign \new_[25812]_  = (~\s4_data_i[6]  | ~\new_[30335]_ ) & (~\s0_data_i[6]  | ~\new_[29603]_ );
  assign \new_[25813]_  = (~\new_[30031]_  | ~\s7_data_i[26] ) & (~\new_[29052]_  | ~\s6_data_i[26] );
  assign \new_[25814]_  = (~\s4_data_i[15]  | ~\new_[30335]_ ) & (~\s0_data_i[15]  | ~\new_[29603]_ );
  assign \new_[25815]_  = (~\new_[29025]_  | ~\s5_data_i[18] ) & (~\new_[30469]_  | ~\s3_data_i[18] );
  assign \new_[25816]_  = (~\s4_data_i[24]  | ~\new_[30335]_ ) & (~\s0_data_i[24]  | ~\new_[29603]_ );
  assign \new_[25817]_  = (~\new_[30227]_  | ~\s10_data_i[1] ) & (~\new_[29706]_  | ~\s9_data_i[1] );
  assign \new_[25818]_  = ~\new_[27352]_ ;
  assign \new_[25819]_  = (~\new_[30311]_  | ~\s11_data_i[3] ) & (~\new_[29636]_  | ~\s8_data_i[3] );
  assign \new_[25820]_  = (~\new_[28842]_  | ~\s4_data_i[18] ) & (~\new_[29434]_  | ~\s0_data_i[18] );
  assign \new_[25821]_  = (~\new_[30200]_  | ~\s11_data_i[29] ) & (~\new_[29428]_  | ~\s8_data_i[29] );
  assign \new_[25822]_  = ~\new_[27343]_ ;
  assign \new_[25823]_  = (~\s11_data_i[22]  | ~\new_[29205]_ ) & (~\s8_data_i[22]  | ~\new_[29241]_ );
  assign \new_[25824]_  = \new_[28807]_  | \new_[30682]_ ;
  assign \new_[25825]_  = (~\s5_data_i[21]  | ~\new_[29649]_ ) & (~\s3_data_i[21]  | ~\new_[29035]_ );
  assign \new_[25826]_  = (~\s14_data_i[5]  | ~\new_[30026]_ ) & (~\s12_data_i[5]  | ~\new_[29711]_ );
  assign \new_[25827]_  = (~\new_[29953]_  | ~\s11_data_i[24] ) & (~\new_[29627]_  | ~\s8_data_i[24] );
  assign \new_[25828]_  = (~\new_[28842]_  | ~\s4_data_i[14] ) & (~\new_[29434]_  | ~\s0_data_i[14] );
  assign \new_[25829]_  = ~\new_[29171]_  | ~\new_[28121]_ ;
  assign \new_[25830]_  = (~\new_[30031]_  | ~\s7_data_i[14] ) & (~\new_[29052]_  | ~\s6_data_i[14] );
  assign \new_[25831]_  = (~\new_[29976]_  | ~\s14_data_i[30] ) & (~\new_[28957]_  | ~\s12_data_i[30] );
  assign \new_[25832]_  = (~\new_[29705]_  | ~\s10_data_i[14] ) & (~\new_[30354]_  | ~\s9_data_i[14] );
  assign \new_[25833]_  = (~\new_[29012]_  | ~\s10_data_i[23] ) & (~\new_[29185]_  | ~\s9_data_i[23] );
  assign \new_[25834]_  = ~\new_[27364]_ ;
  assign \new_[25835]_  = (~\new_[29036]_  | ~\s5_data_i[31] ) & (~\new_[30429]_  | ~\s3_data_i[31] );
  assign \new_[25836]_  = (~\new_[29976]_  | ~\s14_data_i[14] ) & (~\new_[28957]_  | ~\s12_data_i[14] );
  assign \new_[25837]_  = (~\new_[29025]_  | ~\s5_data_i[17] ) & (~\new_[30469]_  | ~\s3_data_i[17] );
  assign \new_[25838]_  = (~\s11_data_i[7]  | ~\new_[29205]_ ) & (~\s8_data_i[7]  | ~\new_[29241]_ );
  assign \new_[25839]_  = (~\new_[30284]_  | ~\s11_data_i[31] ) & (~\new_[29420]_  | ~\s8_data_i[31] );
  assign \new_[25840]_  = (~\s5_data_i[27]  | ~\new_[29649]_ ) & (~\s3_data_i[27]  | ~\new_[29035]_ );
  assign \new_[25841]_  = (~\s14_data_i[21]  | ~\new_[30026]_ ) & (~\s12_data_i[21]  | ~\new_[29711]_ );
  assign \new_[25842]_  = (~\new_[29641]_  | ~\s14_data_i[22] ) & (~\new_[29317]_  | ~\s12_data_i[22] );
  assign \new_[25843]_  = (~\new_[29705]_  | ~\s10_data_i[13] ) & (~\new_[30354]_  | ~\s9_data_i[13] );
  assign \new_[25844]_  = ~\new_[27369]_ ;
  assign \new_[25845]_  = (~\new_[29012]_  | ~\s10_data_i[21] ) & (~\new_[29185]_  | ~\s9_data_i[21] );
  assign \new_[25846]_  = ~\new_[30743]_  | ~\new_[6033]_ ;
  assign \new_[25847]_  = (~\new_[30260]_  | ~\s11_data_i[13] ) & (~\new_[29670]_  | ~\s8_data_i[13] );
  assign \new_[25848]_  = (~\new_[29641]_  | ~\s14_data_i[21] ) & (~\new_[29317]_  | ~\s12_data_i[21] );
  assign \new_[25849]_  = (~\new_[29976]_  | ~\s14_data_i[13] ) & (~\new_[28957]_  | ~\s12_data_i[13] );
  assign \new_[25850]_  = (~\new_[29025]_  | ~\s5_data_i[13] ) & (~\new_[30469]_  | ~\s3_data_i[13] );
  assign \new_[25851]_  = (~\new_[30181]_  | ~\s14_data_i[31] ) & (~\new_[29640]_  | ~\s12_data_i[31] );
  assign \new_[25852]_  = (~\s2_data_i[21]  | ~\new_[29625]_ ) & (~\s1_data_i[21]  | ~\new_[29215]_ );
  assign \new_[25853]_  = (~\new_[29641]_  | ~\s14_data_i[20] ) & (~\new_[29317]_  | ~\s12_data_i[20] );
  assign \new_[25854]_  = (~\new_[29641]_  | ~\s14_data_i[30] ) & (~\new_[29317]_  | ~\s12_data_i[30] );
  assign \new_[25855]_  = (~\new_[29705]_  | ~\s10_data_i[12] ) & (~\new_[30354]_  | ~\s9_data_i[12] );
  assign \new_[25856]_  = (~\s10_data_i[15]  | ~\new_[29749]_ ) & (~\s9_data_i[15]  | ~\new_[29034]_ );
  assign \new_[25857]_  = ~\new_[27373]_ ;
  assign \new_[25858]_  = (~\s10_data_i[4]  | ~\new_[29749]_ ) & (~\s9_data_i[4]  | ~\new_[29034]_ );
  assign \new_[25859]_  = (~\new_[29953]_  | ~\s11_data_i[19] ) & (~\new_[29627]_  | ~\s8_data_i[19] );
  assign \new_[25860]_  = (~\new_[30200]_  | ~\s11_data_i[20] ) & (~\new_[29428]_  | ~\s8_data_i[20] );
  assign \new_[25861]_  = ~\new_[29840]_  | ~\new_[5926]_ ;
  assign \new_[25862]_  = (~\new_[29976]_  | ~\s14_data_i[12] ) & (~\new_[28957]_  | ~\s12_data_i[12] );
  assign \new_[25863]_  = (~\s5_data_i[4]  | ~\new_[29649]_ ) & (~\s3_data_i[4]  | ~\new_[29035]_ );
  assign \new_[25864]_  = (~\new_[29025]_  | ~\s5_data_i[12] ) & (~\new_[30469]_  | ~\s3_data_i[12] );
  assign \new_[25865]_  = (~\new_[29045]_  | ~\s10_data_i[31] ) & (~\new_[29951]_  | ~\s9_data_i[31] );
  assign \new_[25866]_  = (~\new_[30227]_  | ~\s10_data_i[9] ) & (~\new_[29706]_  | ~\s9_data_i[9] );
  assign \new_[25867]_  = (~\new_[28842]_  | ~\s4_data_i[11] ) & (~\new_[29434]_  | ~\s0_data_i[11] );
  assign \new_[25868]_  = (~\s11_data_i[4]  | ~\new_[29205]_ ) & (~\s8_data_i[4]  | ~\new_[29241]_ );
  assign \new_[25869]_  = (~\new_[30031]_  | ~\s7_data_i[11] ) & (~\new_[29052]_  | ~\s6_data_i[11] );
  assign \new_[25870]_  = ~\new_[27056]_ ;
  assign \new_[25871]_  = (~\s14_data_i[4]  | ~\new_[30026]_ ) & (~\s12_data_i[4]  | ~\new_[29711]_ );
  assign \new_[25872]_  = (~\new_[29953]_  | ~\s11_data_i[17] ) & (~\new_[29627]_  | ~\s8_data_i[17] );
  assign \new_[25873]_  = (~\new_[29641]_  | ~\s14_data_i[17] ) & (~\new_[29317]_  | ~\s12_data_i[17] );
  assign \new_[25874]_  = (~\s2_data_i[4]  | ~\new_[29625]_ ) & (~\s1_data_i[4]  | ~\new_[29215]_ );
  assign \new_[25875]_  = (~\new_[29710]_  | ~\s10_data_i[0] ) & (~\new_[29024]_  | ~\s9_data_i[0] );
  assign \new_[25876]_  = (~\s4_data_i[20]  | ~\new_[30335]_ ) & (~\s0_data_i[20]  | ~\new_[29603]_ );
  assign \new_[25877]_  = (~\new_[29021]_  | ~\s10_data_i[19] ) & (~\new_[29709]_  | ~\s9_data_i[19] );
  assign \new_[25878]_  = (~\new_[28842]_  | ~\s4_data_i[10] ) & (~\new_[29434]_  | ~\s0_data_i[10] );
  assign \new_[25879]_  = (~\new_[29641]_  | ~\s14_data_i[16] ) & (~\new_[29317]_  | ~\s12_data_i[16] );
  assign \new_[25880]_  = ~\new_[26993]_ ;
  assign \new_[25881]_  = ~\new_[26777]_ ;
  assign \new_[25882]_  = (~\new_[29641]_  | ~\s14_data_i[15] ) & (~\new_[29317]_  | ~\s12_data_i[15] );
  assign \new_[25883]_  = (~\new_[29976]_  | ~\s14_data_i[0] ) & (~\new_[28957]_  | ~\s12_data_i[0] );
  assign \new_[25884]_  = (~\new_[29012]_  | ~\s10_data_i[14] ) & (~\new_[29185]_  | ~\s9_data_i[14] );
  assign \new_[25885]_  = (~\s4_data_i[3]  | ~\new_[30335]_ ) & (~\s0_data_i[3]  | ~\new_[29603]_ );
  assign \new_[25886]_  = (~\new_[28842]_  | ~\s4_data_i[9] ) & (~\new_[29434]_  | ~\s0_data_i[9] );
  assign \new_[25887]_  = (~\s10_data_i[20]  | ~\new_[29749]_ ) & (~\s9_data_i[20]  | ~\new_[29034]_ );
  assign \new_[25888]_  = (~\new_[30031]_  | ~\s7_data_i[9] ) & (~\new_[29052]_  | ~\s6_data_i[9] );
  assign \new_[25889]_  = (~\new_[29953]_  | ~\s11_data_i[30] ) & (~\new_[29627]_  | ~\s8_data_i[30] );
  assign \new_[25890]_  = (~\new_[29705]_  | ~\s10_data_i[9] ) & (~\new_[30354]_  | ~\s9_data_i[9] );
  assign \new_[25891]_  = (~\new_[29710]_  | ~\s10_data_i[7] ) & (~\new_[29024]_  | ~\s9_data_i[7] );
  assign \new_[25892]_  = ~\new_[27718]_ ;
  assign \new_[25893]_  = (~\new_[29012]_  | ~\s10_data_i[13] ) & (~\new_[29185]_  | ~\s9_data_i[13] );
  assign \new_[25894]_  = (~\new_[29641]_  | ~\s14_data_i[13] ) & (~\new_[29317]_  | ~\s12_data_i[13] );
  assign \new_[25895]_  = (~\new_[30260]_  | ~\s11_data_i[0] ) & (~\new_[29670]_  | ~\s8_data_i[0] );
  assign \new_[25896]_  = (~\new_[29976]_  | ~\s14_data_i[9] ) & (~\new_[28957]_  | ~\s12_data_i[9] );
  assign \new_[25897]_  = (~\s10_data_i[21]  | ~\new_[29749]_ ) & (~\s9_data_i[21]  | ~\new_[29034]_ );
  assign \new_[25898]_  = (~\new_[29012]_  | ~\s10_data_i[12] ) & (~\new_[29185]_  | ~\s9_data_i[12] );
  assign \new_[25899]_  = (~\new_[29710]_  | ~\s10_data_i[30] ) & (~\new_[29024]_  | ~\s9_data_i[30] );
  assign \new_[25900]_  = (~\s2_data_i[19]  | ~\new_[29625]_ ) & (~\s1_data_i[19]  | ~\new_[29215]_ );
  assign \new_[25901]_  = (~\s5_data_i[3]  | ~\new_[29649]_ ) & (~\s3_data_i[3]  | ~\new_[29035]_ );
  assign \new_[25902]_  = (~\new_[30200]_  | ~\s11_data_i[19] ) & (~\new_[29428]_  | ~\s8_data_i[19] );
  assign \new_[25903]_  = (~\new_[29953]_  | ~\s11_data_i[12] ) & (~\new_[29627]_  | ~\s8_data_i[12] );
  assign \new_[25904]_  = (~\new_[29641]_  | ~\s14_data_i[12] ) & (~\new_[29317]_  | ~\s12_data_i[12] );
  assign \new_[25905]_  = (~\new_[28842]_  | ~\s4_data_i[8] ) & (~\new_[29434]_  | ~\s0_data_i[8] );
  assign \new_[25906]_  = (~\new_[29705]_  | ~\s10_data_i[0] ) & (~\new_[30354]_  | ~\s9_data_i[0] );
  assign \new_[25907]_  = ~\new_[27393]_ ;
  assign \new_[25908]_  = (~\s11_data_i[3]  | ~\new_[29205]_ ) & (~\s8_data_i[3]  | ~\new_[29241]_ );
  assign \new_[25909]_  = (~\s11_data_i[29]  | ~\new_[29205]_ ) & (~\s8_data_i[29]  | ~\new_[29241]_ );
  assign \new_[25910]_  = (~\new_[29025]_  | ~\s5_data_i[8] ) & (~\new_[30469]_  | ~\s3_data_i[8] );
  assign \new_[25911]_  = (~\new_[29641]_  | ~\s14_data_i[10] ) & (~\new_[29317]_  | ~\s12_data_i[10] );
  assign \new_[25912]_  = (~\new_[30260]_  | ~\s11_data_i[27] ) & (~\new_[29670]_  | ~\s8_data_i[27] );
  assign \new_[25913]_  = (~\new_[29976]_  | ~\s14_data_i[16] ) & (~\new_[28957]_  | ~\s12_data_i[16] );
  assign \new_[25914]_  = (~\s14_data_i[20]  | ~\new_[30026]_ ) & (~\s12_data_i[20]  | ~\new_[29711]_ );
  assign \new_[25915]_  = (~\new_[30193]_  | ~\s7_data_i[4] ) & (~\new_[29298]_  | ~\s6_data_i[4] );
  assign \new_[25916]_  = ~\new_[27400]_ ;
  assign \new_[25917]_  = (~\new_[29649]_  | ~\s5_data_i[31] ) & (~\new_[29035]_  | ~\s3_data_i[31] );
  assign \new_[25918]_  = (~\new_[30193]_  | ~\s7_data_i[20] ) & (~\new_[29298]_  | ~\s6_data_i[20] );
  assign \new_[25919]_  = (~\new_[29953]_  | ~\s11_data_i[9] ) & (~\new_[29627]_  | ~\s8_data_i[9] );
  assign \new_[25920]_  = (~\new_[30260]_  | ~\s11_data_i[7] ) & (~\new_[29670]_  | ~\s8_data_i[7] );
  assign \new_[25921]_  = (~\new_[29021]_  | ~\s10_data_i[26] ) & (~\new_[29709]_  | ~\s9_data_i[26] );
  assign \new_[25922]_  = (~\new_[29025]_  | ~\s5_data_i[7] ) & (~\new_[30469]_  | ~\s3_data_i[7] );
  assign \new_[25923]_  = (~\new_[29012]_  | ~\s10_data_i[8] ) & (~\new_[29185]_  | ~\s9_data_i[8] );
  assign \new_[25924]_  = (~\new_[29631]_  | ~\s14_data_i[28] ) & (~\new_[29621]_  | ~\s12_data_i[28] );
  assign \new_[25925]_  = ~\new_[30389]_  & ~\new_[30172]_ ;
  assign \new_[25926]_  = (~\new_[29641]_  | ~\s14_data_i[8] ) & (~\new_[29317]_  | ~\s12_data_i[8] );
  assign \new_[25927]_  = (~\new_[30181]_  | ~\s14_data_i[9] ) & (~\new_[29640]_  | ~\s12_data_i[9] );
  assign \new_[25928]_  = (~\new_[29628]_  | ~\s4_data_i[1] ) & (~\new_[29258]_  | ~\s0_data_i[1] );
  assign \new_[25929]_  = (~\new_[30060]_  | ~\s7_data_i[9] ) & (~\new_[29704]_  | ~\s6_data_i[9] );
  assign \new_[25930]_  = (~\new_[28842]_  | ~\s4_data_i[25] ) & (~\new_[29434]_  | ~\s0_data_i[25] );
  assign \new_[25931]_  = ~\new_[27405]_ ;
  assign \new_[25932]_  = (~\new_[30260]_  | ~\s11_data_i[6] ) & (~\new_[29670]_  | ~\s8_data_i[6] );
  assign \new_[25933]_  = (~\new_[29953]_  | ~\s11_data_i[7] ) & (~\new_[29627]_  | ~\s8_data_i[7] );
  assign \new_[25934]_  = (~\s4_data_i[2]  | ~\new_[30335]_ ) & (~\s0_data_i[2]  | ~\new_[29603]_ );
  assign \new_[25935]_  = (~\new_[29641]_  | ~\s14_data_i[7] ) & (~\new_[29317]_  | ~\s12_data_i[7] );
  assign \new_[25936]_  = (~\new_[29534]_  | ~\s5_data_i[19] ) & (~\new_[29579]_  | ~\s3_data_i[19] );
  assign \new_[25937]_  = (~\new_[29976]_  | ~\s14_data_i[6] ) & (~\new_[28957]_  | ~\s12_data_i[6] );
  assign \new_[25938]_  = (~\s2_data_i[29]  | ~\new_[29625]_ ) & (~\s1_data_i[29]  | ~\new_[29215]_ );
  assign \new_[25939]_  = (~\new_[29012]_  | ~\s10_data_i[6] ) & (~\new_[29185]_  | ~\s9_data_i[6] );
  assign \new_[25940]_  = (~\new_[29025]_  | ~\s5_data_i[16] ) & (~\new_[30469]_  | ~\s3_data_i[16] );
  assign \new_[25941]_  = (~\s10_data_i[2]  | ~\new_[29749]_ ) & (~\s9_data_i[2]  | ~\new_[29034]_ );
  assign \new_[25942]_  = (~\new_[29705]_  | ~\s10_data_i[31] ) & (~\new_[30354]_  | ~\s9_data_i[31] );
  assign \new_[25943]_  = (~\new_[28842]_  | ~\s4_data_i[5] ) & (~\new_[29434]_  | ~\s0_data_i[5] );
  assign \new_[25944]_  = ~\new_[30743]_  & ~\new_[6174]_ ;
  assign \new_[25945]_  = (~\new_[29953]_  | ~\s11_data_i[6] ) & (~\new_[29627]_  | ~\s8_data_i[6] );
  assign \new_[25946]_  = (~\new_[30181]_  | ~\s14_data_i[10] ) & (~\new_[29640]_  | ~\s12_data_i[10] );
  assign \new_[25947]_  = \new_[29464]_  | \new_[30276]_ ;
  assign \new_[25948]_  = (~\new_[30031]_  | ~\s7_data_i[5] ) & (~\new_[29052]_  | ~\s6_data_i[5] );
  assign \new_[25949]_  = (~\new_[29705]_  | ~\s10_data_i[5] ) & (~\new_[30354]_  | ~\s9_data_i[5] );
  assign \new_[25950]_  = (~\new_[29953]_  | ~\s11_data_i[28] ) & (~\new_[29627]_  | ~\s8_data_i[28] );
  assign \new_[25951]_  = (~\new_[29012]_  | ~\s10_data_i[5] ) & (~\new_[29185]_  | ~\s9_data_i[5] );
  assign \new_[25952]_  = (~\new_[30181]_  | ~\s14_data_i[0] ) & (~\new_[29640]_  | ~\s12_data_i[0] );
  assign \new_[25953]_  = (~\new_[29641]_  | ~\s14_data_i[5] ) & (~\new_[29317]_  | ~\s12_data_i[5] );
  assign \new_[25954]_  = (~\new_[30031]_  | ~\s7_data_i[6] ) & (~\new_[29052]_  | ~\s6_data_i[6] );
  assign \new_[25955]_  = ~\new_[27414]_ ;
  assign \new_[25956]_  = (~\s11_data_i[2]  | ~\new_[29205]_ ) & (~\s8_data_i[2]  | ~\new_[29241]_ );
  assign \new_[25957]_  = (~\new_[29976]_  | ~\s14_data_i[18] ) & (~\new_[28957]_  | ~\s12_data_i[18] );
  assign \new_[25958]_  = (~\s4_data_i[23]  | ~\new_[30335]_ ) & (~\s0_data_i[23]  | ~\new_[29603]_ );
  assign \new_[25959]_  = (~\new_[30284]_  | ~\s11_data_i[29] ) & (~\new_[29420]_  | ~\s8_data_i[29] );
  assign \new_[25960]_  = (~\new_[28842]_  | ~\s4_data_i[16] ) & (~\new_[29434]_  | ~\s0_data_i[16] );
  assign \new_[25961]_  = (~\new_[29976]_  | ~\s14_data_i[1] ) & (~\new_[28957]_  | ~\s12_data_i[1] );
  assign \new_[25962]_  = (~\new_[30060]_  | ~\s7_data_i[0] ) & (~\new_[29704]_  | ~\s6_data_i[0] );
  assign \new_[25963]_  = (~\new_[29012]_  | ~\s10_data_i[4] ) & (~\new_[29185]_  | ~\s9_data_i[4] );
  assign \new_[25964]_  = (~\new_[29045]_  | ~\s10_data_i[8] ) & (~\new_[29951]_  | ~\s9_data_i[8] );
  assign \new_[25965]_  = (~\new_[29021]_  | ~\s10_data_i[25] ) & (~\new_[29709]_  | ~\s9_data_i[25] );
  assign \new_[25966]_  = ~\new_[27717]_ ;
  assign \new_[25967]_  = (~\new_[30193]_  | ~\s7_data_i[21] ) & (~\new_[29298]_  | ~\s6_data_i[21] );
  assign \new_[25968]_  = (~\new_[29045]_  | ~\s10_data_i[10] ) & (~\new_[29951]_  | ~\s9_data_i[10] );
  assign \new_[25969]_  = (~\new_[28842]_  | ~\s4_data_i[4] ) & (~\new_[29434]_  | ~\s0_data_i[4] );
  assign \new_[25970]_  = (~\new_[29641]_  | ~\s14_data_i[4] ) & (~\new_[29317]_  | ~\s12_data_i[4] );
  assign \new_[25971]_  = (~\new_[29628]_  | ~\s4_data_i[8] ) & (~\new_[29258]_  | ~\s0_data_i[8] );
  assign \new_[25972]_  = (~\new_[29628]_  | ~\s4_data_i[0] ) & (~\new_[29258]_  | ~\s0_data_i[0] );
  assign \new_[25973]_  = (~\new_[30031]_  | ~\s7_data_i[4] ) & (~\new_[29052]_  | ~\s6_data_i[4] );
  assign \new_[25974]_  = (~\new_[29705]_  | ~\s10_data_i[4] ) & (~\new_[30354]_  | ~\s9_data_i[4] );
  assign \new_[25975]_  = ~\new_[28836]_  & ~\new_[26657]_ ;
  assign \new_[25976]_  = ~\new_[26886]_ ;
  assign \new_[25977]_  = \new_[29566]_  & \new_[28001]_ ;
  assign \new_[25978]_  = (~\new_[29953]_  | ~\s11_data_i[3] ) & (~\new_[29627]_  | ~\s8_data_i[3] );
  assign \new_[25979]_  = (~\new_[30260]_  | ~\s11_data_i[4] ) & (~\new_[29670]_  | ~\s8_data_i[4] );
  assign \new_[25980]_  = (~\new_[29641]_  | ~\s14_data_i[3] ) & (~\new_[29317]_  | ~\s12_data_i[3] );
  assign \new_[25981]_  = (~\new_[30200]_  | ~\s11_data_i[8] ) & (~\new_[29428]_  | ~\s8_data_i[8] );
  assign \new_[25982]_  = (~\new_[29012]_  | ~\s10_data_i[2] ) & (~\new_[29185]_  | ~\s9_data_i[2] );
  assign \new_[25983]_  = (~\new_[29705]_  | ~\s10_data_i[24] ) & (~\new_[30354]_  | ~\s9_data_i[24] );
  assign \new_[25984]_  = (~\new_[29641]_  | ~\s14_data_i[2] ) & (~\new_[29317]_  | ~\s12_data_i[2] );
  assign \new_[25985]_  = (~\new_[29705]_  | ~\s10_data_i[15] ) & (~\new_[30354]_  | ~\s9_data_i[15] );
  assign \new_[25986]_  = (~\new_[30181]_  | ~\s14_data_i[6] ) & (~\new_[29640]_  | ~\s12_data_i[6] );
  assign \new_[25987]_  = ~\new_[26658]_ ;
  assign \new_[25988]_  = (~\s10_data_i[19]  | ~\new_[29749]_ ) & (~\s9_data_i[19]  | ~\new_[29034]_ );
  assign \new_[25989]_  = (~\new_[29012]_  | ~\s10_data_i[1] ) & (~\new_[29185]_  | ~\s9_data_i[1] );
  assign \new_[25990]_  = (~\s14_data_i[14]  | ~\new_[30026]_ ) & (~\s12_data_i[14]  | ~\new_[29711]_ );
  assign \new_[25991]_  = (~\new_[29953]_  | ~\s11_data_i[1] ) & (~\new_[29627]_  | ~\s8_data_i[1] );
  assign \new_[25992]_  = (~\s4_data_i[1]  | ~\new_[30335]_ ) & (~\s0_data_i[1]  | ~\new_[29603]_ );
  assign \new_[25993]_  = ~\new_[28492]_  & ~\new_[30109]_ ;
  assign \new_[25994]_  = (~\new_[30260]_  | ~\s11_data_i[3] ) & (~\new_[29670]_  | ~\s8_data_i[3] );
  assign \new_[25995]_  = (~\new_[30311]_  | ~\s11_data_i[9] ) & (~\new_[29636]_  | ~\s8_data_i[9] );
  assign \new_[25996]_  = ~\new_[27378]_ ;
  assign \new_[25997]_  = (~\new_[29976]_  | ~\s14_data_i[3] ) & (~\new_[28957]_  | ~\s12_data_i[3] );
  assign \new_[25998]_  = (~\new_[29025]_  | ~\s5_data_i[3] ) & (~\new_[30469]_  | ~\s3_data_i[3] );
  assign \new_[25999]_  = ~\new_[29230]_  | ~\new_[28594]_ ;
  assign \new_[26000]_  = (~\new_[30284]_  | ~\s11_data_i[12] ) & (~\new_[29420]_  | ~\s8_data_i[12] );
  assign \new_[26001]_  = (~\new_[29012]_  | ~\s10_data_i[0] ) & (~\new_[29185]_  | ~\s9_data_i[0] );
  assign \new_[26002]_  = (~\s10_data_i[26]  | ~\new_[29749]_ ) & (~\s9_data_i[26]  | ~\new_[29034]_ );
  assign \new_[26003]_  = ~\new_[27429]_ ;
  assign \new_[26004]_  = (~\new_[29021]_  | ~\s10_data_i[27] ) & (~\new_[29709]_  | ~\s9_data_i[27] );
  assign \new_[26005]_  = (~\new_[29953]_  | ~\s11_data_i[0] ) & (~\new_[29627]_  | ~\s8_data_i[0] );
  assign \new_[26006]_  = (~\new_[28842]_  | ~\s4_data_i[2] ) & (~\new_[29434]_  | ~\s0_data_i[2] );
  assign \new_[26007]_  = (~\new_[29641]_  | ~\s14_data_i[0] ) & (~\new_[29317]_  | ~\s12_data_i[0] );
  assign \new_[26008]_  = (~\new_[30060]_  | ~\s7_data_i[11] ) & (~\new_[29704]_  | ~\s6_data_i[11] );
  assign \new_[26009]_  = (~\s5_data_i[19]  | ~\new_[29649]_ ) & (~\s3_data_i[19]  | ~\new_[29035]_ );
  assign \new_[26010]_  = (~\new_[29641]_  | ~\s14_data_i[18] ) & (~\new_[29317]_  | ~\s12_data_i[18] );
  assign \new_[26011]_  = (~\new_[30260]_  | ~\s11_data_i[2] ) & (~\new_[29670]_  | ~\s8_data_i[2] );
  assign \new_[26012]_  = (~\new_[29025]_  | ~\s5_data_i[2] ) & (~\new_[30469]_  | ~\s3_data_i[2] );
  assign \new_[26013]_  = (~\new_[29976]_  | ~\s14_data_i[28] ) & (~\new_[28957]_  | ~\s12_data_i[28] );
  assign \new_[26014]_  = (~\new_[30193]_  | ~\s7_data_i[22] ) & (~\new_[29298]_  | ~\s6_data_i[22] );
  assign \new_[26015]_  = (~\s14_data_i[1]  | ~\new_[30026]_ ) & (~\s12_data_i[1]  | ~\new_[29711]_ );
  assign \new_[26016]_  = (~\new_[29705]_  | ~\s10_data_i[1] ) & (~\new_[30354]_  | ~\s9_data_i[1] );
  assign \new_[26017]_  = (~\new_[28842]_  | ~\s4_data_i[28] ) & (~\new_[29434]_  | ~\s0_data_i[28] );
  assign \new_[26018]_  = (~\new_[30260]_  | ~\s11_data_i[1] ) & (~\new_[29670]_  | ~\s8_data_i[1] );
  assign \new_[26019]_  = (~\new_[30031]_  | ~\s7_data_i[0] ) & (~\new_[29052]_  | ~\s6_data_i[0] );
  assign \new_[26020]_  = (~\new_[29025]_  | ~\s5_data_i[21] ) & (~\new_[30469]_  | ~\s3_data_i[21] );
  assign \new_[26021]_  = (~\s11_data_i[19]  | ~\new_[29205]_ ) & (~\s8_data_i[19]  | ~\new_[29241]_ );
  assign \new_[26022]_  = ~\new_[27991]_  | ~\new_[30107]_ ;
  assign \new_[26023]_  = (~\s10_data_i[28]  | ~\new_[29749]_ ) & (~\s9_data_i[28]  | ~\new_[29034]_ );
  assign \new_[26024]_  = (~\new_[30311]_  | ~\s11_data_i[31] ) & (~\new_[29636]_  | ~\s8_data_i[31] );
  assign \new_[26025]_  = ~\new_[27339]_ ;
  assign \new_[26026]_  = (~\s4_data_i[28]  | ~\new_[30335]_ ) & (~\s0_data_i[28]  | ~\new_[29603]_ );
  assign \new_[26027]_  = (~\new_[29021]_  | ~\s10_data_i[3] ) & (~\new_[29709]_  | ~\s9_data_i[3] );
  assign \new_[26028]_  = (~\new_[29628]_  | ~\s4_data_i[30] ) & (~\new_[29258]_  | ~\s0_data_i[30] );
  assign \new_[26029]_  = (~\new_[29045]_  | ~\s10_data_i[30] ) & (~\new_[29951]_  | ~\s9_data_i[30] );
  assign \new_[26030]_  = (~\new_[30311]_  | ~\s11_data_i[30] ) & (~\new_[29636]_  | ~\s8_data_i[30] );
  assign \new_[26031]_  = (~\new_[30181]_  | ~\s14_data_i[30] ) & (~\new_[29640]_  | ~\s12_data_i[30] );
  assign \new_[26032]_  = (~\new_[30031]_  | ~\s7_data_i[18] ) & (~\new_[29052]_  | ~\s6_data_i[18] );
  assign \new_[26033]_  = (~\new_[29976]_  | ~\s14_data_i[21] ) & (~\new_[28957]_  | ~\s12_data_i[21] );
  assign \new_[26034]_  = (~\s4_data_i[18]  | ~\new_[30335]_ ) & (~\s0_data_i[18]  | ~\new_[29603]_ );
  assign \new_[26035]_  = ~\new_[26720]_ ;
  assign \new_[26036]_  = (~\s14_data_i[7]  | ~\new_[30026]_ ) & (~\s12_data_i[7]  | ~\new_[29711]_ );
  assign \new_[26037]_  = (~\new_[30260]_  | ~\s11_data_i[15] ) & (~\new_[29670]_  | ~\s8_data_i[15] );
  assign \new_[26038]_  = ~\new_[29992]_  & ~\new_[30164]_ ;
  assign \new_[26039]_  = (~\s14_data_i[0]  | ~\new_[30026]_ ) & (~\s12_data_i[0]  | ~\new_[29711]_ );
  assign \new_[26040]_  = (~\new_[29045]_  | ~\s10_data_i[25] ) & (~\new_[29951]_  | ~\s9_data_i[25] );
  assign \new_[26041]_  = (~\s5_data_i[7]  | ~\new_[29649]_ ) & (~\s3_data_i[7]  | ~\new_[29035]_ );
  assign \new_[26042]_  = (~\new_[30181]_  | ~\s14_data_i[29] ) & (~\new_[29640]_  | ~\s12_data_i[29] );
  assign \new_[26043]_  = (~\s2_data_i[0]  | ~\new_[29625]_ ) & (~\s1_data_i[0]  | ~\new_[29215]_ );
  assign \new_[26044]_  = (~\new_[30060]_  | ~\s7_data_i[28] ) & (~\new_[29704]_  | ~\s6_data_i[28] );
  assign \new_[26045]_  = (~\new_[30227]_  | ~\s10_data_i[2] ) & (~\new_[29706]_  | ~\s9_data_i[2] );
  assign \new_[26046]_  = (~\new_[29641]_  | ~\s14_data_i[19] ) & (~\new_[29317]_  | ~\s12_data_i[19] );
  assign \new_[26047]_  = (~\s5_data_i[28]  | ~\new_[29649]_ ) & (~\s3_data_i[28]  | ~\new_[29035]_ );
  assign \new_[26048]_  = (~\new_[29705]_  | ~\s10_data_i[20] ) & (~\new_[30354]_  | ~\s9_data_i[20] );
  assign \new_[26049]_  = (~\new_[29025]_  | ~\s5_data_i[28] ) & (~\new_[30469]_  | ~\s3_data_i[28] );
  assign \new_[26050]_  = (~\new_[29628]_  | ~\s4_data_i[27] ) & (~\new_[29258]_  | ~\s0_data_i[27] );
  assign \new_[26051]_  = ~\new_[28562]_  & ~\new_[28960]_ ;
  assign \new_[26052]_  = (~\new_[29045]_  | ~\s10_data_i[27] ) & (~\new_[29951]_  | ~\s9_data_i[27] );
  assign \new_[26053]_  = ~\new_[26700]_ ;
  assign \new_[26054]_  = (~\new_[30311]_  | ~\s11_data_i[27] ) & (~\new_[29636]_  | ~\s8_data_i[27] );
  assign \new_[26055]_  = (~\new_[29976]_  | ~\s14_data_i[2] ) & (~\new_[28957]_  | ~\s12_data_i[2] );
  assign \new_[26056]_  = (~\new_[29025]_  | ~\s5_data_i[25] ) & (~\new_[30469]_  | ~\s3_data_i[25] );
  assign \new_[26057]_  = (~\new_[29045]_  | ~\s10_data_i[26] ) & (~\new_[29951]_  | ~\s9_data_i[26] );
  assign \new_[26058]_  = (~\s5_data_i[22]  | ~\new_[29649]_ ) & (~\s3_data_i[22]  | ~\new_[29035]_ );
  assign \new_[26059]_  = ~\new_[28111]_  | ~\new_[29877]_ ;
  assign \new_[26060]_  = (~\s5_data_i[1]  | ~\new_[29649]_ ) & (~\s3_data_i[1]  | ~\new_[29035]_ );
  assign \new_[26061]_  = (~\new_[30181]_  | ~\s14_data_i[25] ) & (~\new_[29640]_  | ~\s12_data_i[25] );
  assign \new_[26062]_  = (~\new_[28842]_  | ~\s4_data_i[20] ) & (~\new_[29434]_  | ~\s0_data_i[20] );
  assign \new_[26063]_  = (~\new_[30181]_  | ~\s14_data_i[4] ) & (~\new_[29640]_  | ~\s12_data_i[4] );
  assign \new_[26064]_  = (~\new_[29628]_  | ~\s4_data_i[24] ) & (~\new_[29258]_  | ~\s0_data_i[24] );
  assign \new_[26065]_  = (~\s11_data_i[28]  | ~\new_[29205]_ ) & (~\s8_data_i[28]  | ~\new_[29241]_ );
  assign \new_[26066]_  = (~\new_[30060]_  | ~\s7_data_i[24] ) & (~\new_[29704]_  | ~\s6_data_i[24] );
  assign \new_[26067]_  = (~\s10_data_i[7]  | ~\new_[29749]_ ) & (~\s9_data_i[7]  | ~\new_[29034]_ );
  assign \new_[26068]_  = (~\new_[30181]_  | ~\s14_data_i[24] ) & (~\new_[29640]_  | ~\s12_data_i[24] );
  assign \new_[26069]_  = ~\new_[27444]_ ;
  assign \new_[26070]_  = (~\new_[29705]_  | ~\s10_data_i[21] ) & (~\new_[30354]_  | ~\s9_data_i[21] );
  assign \new_[26071]_  = (~\new_[29628]_  | ~\s4_data_i[23] ) & (~\new_[29258]_  | ~\s0_data_i[23] );
  assign \new_[26072]_  = (~\new_[29045]_  | ~\s10_data_i[23] ) & (~\new_[29951]_  | ~\s9_data_i[23] );
  assign \new_[26073]_  = (~\s14_data_i[18]  | ~\new_[30026]_ ) & (~\s12_data_i[18]  | ~\new_[29711]_ );
  assign \new_[26074]_  = ~\new_[30842]_  & ~\new_[31180]_ ;
  assign \new_[26075]_  = (~\new_[28842]_  | ~\s4_data_i[21] ) & (~\new_[29434]_  | ~\s0_data_i[21] );
  assign \new_[26076]_  = (~\new_[30260]_  | ~\s11_data_i[22] ) & (~\new_[29670]_  | ~\s8_data_i[22] );
  assign \new_[26077]_  = ~\new_[30636]_  | ~\new_[30329]_ ;
  assign \new_[26078]_  = (~\new_[29628]_  | ~\s4_data_i[22] ) & (~\new_[29258]_  | ~\s0_data_i[22] );
  assign \new_[26079]_  = (~\new_[29045]_  | ~\s10_data_i[22] ) & (~\new_[29951]_  | ~\s9_data_i[22] );
  assign \new_[26080]_  = (~\s10_data_i[6]  | ~\new_[29749]_ ) & (~\s9_data_i[6]  | ~\new_[29034]_ );
  assign \new_[26081]_  = (~\new_[30311]_  | ~\s11_data_i[22] ) & (~\new_[29636]_  | ~\s8_data_i[22] );
  assign \new_[26082]_  = (~\new_[30181]_  | ~\s14_data_i[22] ) & (~\new_[29640]_  | ~\s12_data_i[22] );
  assign \new_[26083]_  = ~\new_[26627]_  & ~\new_[30067]_ ;
  assign \new_[26084]_  = (~\new_[30284]_  | ~\s11_data_i[0] ) & (~\new_[29420]_  | ~\s8_data_i[0] );
  assign \new_[26085]_  = ~\new_[27714]_ ;
  assign \new_[26086]_  = (~\new_[30193]_  | ~\s7_data_i[31] ) & (~\new_[29298]_  | ~\s6_data_i[31] );
  assign \new_[26087]_  = (~\new_[30060]_  | ~\s7_data_i[21] ) & (~\new_[29704]_  | ~\s6_data_i[21] );
  assign \new_[26088]_  = (~\s10_data_i[1]  | ~\new_[29749]_ ) & (~\s9_data_i[1]  | ~\new_[29034]_ );
  assign \new_[26089]_  = (~\new_[30181]_  | ~\s14_data_i[21] ) & (~\new_[29640]_  | ~\s12_data_i[21] );
  assign \new_[26090]_  = (~\new_[30200]_  | ~\s11_data_i[2] ) & (~\new_[29428]_  | ~\s8_data_i[2] );
  assign \new_[26091]_  = (~\new_[29953]_  | ~\s11_data_i[27] ) & (~\new_[29627]_  | ~\s8_data_i[27] );
  assign \new_[26092]_  = (~\new_[29628]_  | ~\s4_data_i[20] ) & (~\new_[29258]_  | ~\s0_data_i[20] );
  assign \new_[26093]_  = (~\new_[30031]_  | ~\s7_data_i[2] ) & (~\new_[29052]_  | ~\s6_data_i[2] );
  assign \new_[26094]_  = (~\new_[30060]_  | ~\s7_data_i[20] ) & (~\new_[29704]_  | ~\s6_data_i[20] );
  assign \new_[26095]_  = (~\new_[29021]_  | ~\s10_data_i[31] ) & (~\new_[29709]_  | ~\s9_data_i[31] );
  assign \new_[26096]_  = (~\new_[30311]_  | ~\s11_data_i[20] ) & (~\new_[29636]_  | ~\s8_data_i[20] );
  assign \new_[26097]_  = \new_[28097]_  | \new_[30684]_ ;
  assign \new_[26098]_  = (~\s2_data_i[28]  | ~\new_[29625]_ ) & (~\s1_data_i[28]  | ~\new_[29215]_ );
  assign \new_[26099]_  = (~\new_[29045]_  | ~\s10_data_i[19] ) & (~\new_[29951]_  | ~\s9_data_i[19] );
  assign \new_[26100]_  = (~\new_[30260]_  | ~\s11_data_i[23] ) & (~\new_[29670]_  | ~\s8_data_i[23] );
  assign \new_[26101]_  = (~\new_[30193]_  | ~\s7_data_i[30] ) & (~\new_[29298]_  | ~\s6_data_i[30] );
  assign \new_[26102]_  = (~\new_[30311]_  | ~\s11_data_i[5] ) & (~\new_[29636]_  | ~\s8_data_i[5] );
  assign \new_[26103]_  = ~\new_[27948]_ ;
  assign \new_[26104]_  = (~\new_[29021]_  | ~\s10_data_i[30] ) & (~\new_[29709]_  | ~\s9_data_i[30] );
  assign \new_[26105]_  = (~\new_[30181]_  | ~\s14_data_i[18] ) & (~\new_[29640]_  | ~\s12_data_i[18] );
  assign \new_[26106]_  = (~\new_[29628]_  | ~\s4_data_i[17] ) & (~\new_[29258]_  | ~\s0_data_i[17] );
  assign \new_[26107]_  = (~\s4_data_i[17]  | ~\new_[30335]_ ) & (~\s0_data_i[17]  | ~\new_[29603]_ );
  assign \new_[26108]_  = ~\new_[27462]_ ;
  assign \new_[26109]_  = (~\new_[29045]_  | ~\s10_data_i[17] ) & (~\new_[29951]_  | ~\s9_data_i[17] );
  assign \new_[26110]_  = (~\new_[29045]_  | ~\s10_data_i[11] ) & (~\new_[29951]_  | ~\s9_data_i[11] );
  assign \new_[26111]_  = (~\s14_data_i[25]  | ~\new_[30026]_ ) & (~\s12_data_i[25]  | ~\new_[29711]_ );
  assign \new_[26112]_  = (~\new_[29021]_  | ~\s10_data_i[14] ) & (~\new_[29709]_  | ~\s9_data_i[14] );
  assign \new_[26113]_  = (~\new_[29021]_  | ~\s10_data_i[29] ) & (~\new_[29709]_  | ~\s9_data_i[29] );
  assign \new_[26114]_  = (~\new_[30181]_  | ~\s14_data_i[16] ) & (~\new_[29640]_  | ~\s12_data_i[16] );
  assign \new_[26115]_  = (~\new_[29045]_  | ~\s10_data_i[15] ) & (~\new_[29951]_  | ~\s9_data_i[15] );
  assign \new_[26116]_  = (~\new_[30311]_  | ~\s11_data_i[15] ) & (~\new_[29636]_  | ~\s8_data_i[15] );
  assign \new_[26117]_  = ~\new_[29774]_  & ~\new_[6091]_ ;
  assign \new_[26118]_  = (~\s14_data_i[24]  | ~\new_[30026]_ ) & (~\s12_data_i[24]  | ~\new_[29711]_ );
  assign \new_[26119]_  = (~\new_[29021]_  | ~\s10_data_i[28] ) & (~\new_[29709]_  | ~\s9_data_i[28] );
  assign \new_[26120]_  = ~\new_[27562]_ ;
  assign \new_[26121]_  = ~\new_[28050]_  | ~\new_[5971]_ ;
  assign \new_[26122]_  = (~\new_[29628]_  | ~\s4_data_i[13] ) & (~\new_[29258]_  | ~\s0_data_i[13] );
  assign \new_[26123]_  = ~\new_[27472]_ ;
  assign \new_[26124]_  = (~\s5_data_i[17]  | ~\new_[29649]_ ) & (~\s3_data_i[17]  | ~\new_[29035]_ );
  assign \new_[26125]_  = (~\new_[30193]_  | ~\s7_data_i[28] ) & (~\new_[29298]_  | ~\s6_data_i[28] );
  assign \new_[26126]_  = (~\new_[28842]_  | ~\s4_data_i[30] ) & (~\new_[29434]_  | ~\s0_data_i[30] );
  assign \new_[26127]_  = (~\new_[30193]_  | ~\s7_data_i[27] ) & (~\new_[29298]_  | ~\s6_data_i[27] );
  assign \new_[26128]_  = ~\new_[27812]_ ;
  assign \new_[26129]_  = (~\s4_data_i[27]  | ~\new_[30335]_ ) & (~\s0_data_i[27]  | ~\new_[29603]_ );
  assign \new_[26130]_  = (~\new_[29628]_  | ~\s4_data_i[11] ) & (~\new_[29258]_  | ~\s0_data_i[11] );
  assign \new_[26131]_  = (~\s11_data_i[17]  | ~\new_[29205]_ ) & (~\s8_data_i[17]  | ~\new_[29241]_ );
  assign \new_[26132]_  = ~\new_[29782]_  | ~\new_[30497]_ ;
  assign \new_[26133]_  = (~\s4_data_i[13]  | ~\new_[30335]_ ) & (~\s0_data_i[13]  | ~\new_[29603]_ );
  assign \new_[26134]_  = (~\new_[30193]_  | ~\s7_data_i[26] ) & (~\new_[29298]_  | ~\s6_data_i[26] );
  assign \new_[26135]_  = (~\new_[30311]_  | ~\s11_data_i[6] ) & (~\new_[29636]_  | ~\s8_data_i[6] );
  assign \new_[26136]_  = ~\new_[27482]_ ;
  assign \new_[26137]_  = (~\new_[30311]_  | ~\s11_data_i[10] ) & (~\new_[29636]_  | ~\s8_data_i[10] );
  assign \new_[26138]_  = (~\s14_data_i[17]  | ~\new_[30026]_ ) & (~\s12_data_i[17]  | ~\new_[29711]_ );
  assign \new_[26139]_  = ~\new_[27770]_ ;
  assign \new_[26140]_  = (~\s10_data_i[9]  | ~\new_[29749]_ ) & (~\s9_data_i[9]  | ~\new_[29034]_ );
  assign \new_[26141]_  = (~\new_[30031]_  | ~\s7_data_i[29] ) & (~\new_[29052]_  | ~\s6_data_i[29] );
  assign \new_[26142]_  = ~\new_[27732]_ ;
  assign \new_[26143]_  = (~\new_[30060]_  | ~\s7_data_i[13] ) & (~\new_[29704]_  | ~\s6_data_i[13] );
  assign \new_[26144]_  = (~\new_[30060]_  | ~\s7_data_i[8] ) & (~\new_[29704]_  | ~\s6_data_i[8] );
  assign \new_[26145]_  = (~\new_[29045]_  | ~\s10_data_i[6] ) & (~\new_[29951]_  | ~\s9_data_i[6] );
  assign \new_[26146]_  = (~\new_[30227]_  | ~\s10_data_i[3] ) & (~\new_[29706]_  | ~\s9_data_i[3] );
  assign \new_[26147]_  = ~\new_[27708]_ ;
  assign \new_[26148]_  = (~\new_[30193]_  | ~\s7_data_i[24] ) & (~\new_[29298]_  | ~\s6_data_i[24] );
  assign \new_[26149]_  = (~\new_[29628]_  | ~\s4_data_i[7] ) & (~\new_[29258]_  | ~\s0_data_i[7] );
  assign \new_[26150]_  = ~\new_[27688]_ ;
  assign \new_[26151]_  = \new_[30051]_  & \new_[6031]_ ;
  assign \new_[26152]_  = ~\new_[30582]_  & ~\new_[31645]_ ;
  assign \new_[26153]_  = ~\new_[27997]_  & ~\new_[29918]_ ;
  assign \new_[26154]_  = (~\new_[29149]_  | ~\s4_data_i[22] ) & (~\new_[29651]_  | ~\s0_data_i[22] );
  assign \new_[26155]_  = ~\new_[28078]_  | ~\new_[6176]_ ;
  assign \new_[26156]_  = ~\new_[28601]_  & ~\new_[30957]_ ;
  assign \new_[26157]_  = \new_[29883]_  & \new_[5930]_ ;
  assign \new_[26158]_  = ~\new_[30099]_  | ~\new_[5928]_ ;
  assign \new_[26159]_  = ~\new_[28888]_  | ~\new_[5984]_ ;
  assign \new_[26160]_  = ~\new_[28801]_  | ~\new_[6206]_ ;
  assign \new_[26161]_  = ~\new_[28358]_  | ~\new_[6064]_ ;
  assign \new_[26162]_  = ~\new_[30312]_  | ~\new_[5898]_ ;
  assign \new_[26163]_  = ~\new_[30121]_  & ~\new_[29061]_ ;
  assign \new_[26164]_  = ~\new_[28129]_  & ~\m4_addr_i[28] ;
  assign \new_[26165]_  = ~\new_[28083]_  | ~\new_[6183]_ ;
  assign \new_[26166]_  = ~\new_[30751]_  & ~\new_[31108]_ ;
  assign \new_[26167]_  = ~\new_[29806]_  | ~\new_[6048]_ ;
  assign \new_[26168]_  = ~\new_[28001]_  | ~\new_[5928]_ ;
  assign \new_[26169]_  = ~\new_[27711]_ ;
  assign \new_[26170]_  = ~\new_[29746]_  | ~\new_[5967]_ ;
  assign \new_[26171]_  = \new_[29962]_  & \new_[6212]_ ;
  assign \new_[26172]_  = ~\new_[28215]_  | ~\new_[5989]_ ;
  assign \new_[26173]_  = ~\new_[28105]_  & ~\new_[31458]_ ;
  assign \new_[26174]_  = ~\new_[29806]_  | ~\new_[6200]_ ;
  assign \new_[26175]_  = ~\new_[28272]_  & ~\new_[31547]_ ;
  assign \new_[26176]_  = ~\new_[28344]_  | ~\new_[31121]_ ;
  assign \new_[26177]_  = (~\new_[30060]_  | ~\s7_data_i[26] ) & (~\new_[29704]_  | ~\s6_data_i[26] );
  assign \new_[26178]_  = \new_[29104]_  & \new_[31423]_ ;
  assign \new_[26179]_  = ~\new_[30764]_  & ~\new_[31855]_ ;
  assign \new_[26180]_  = ~\new_[26951]_ ;
  assign \new_[26181]_  = ~\new_[28083]_  | ~\new_[31132]_ ;
  assign \new_[26182]_  = (~\new_[29710]_  | ~\s10_data_i[2] ) & (~\new_[29024]_  | ~\s9_data_i[2] );
  assign \new_[26183]_  = ~\new_[28785]_  | ~\new_[6007]_ ;
  assign \new_[26184]_  = ~\new_[28785]_  | ~\new_[6217]_ ;
  assign \new_[26185]_  = ~\new_[28785]_  | ~\new_[6095]_ ;
  assign \new_[26186]_  = ~\new_[28078]_  | ~\new_[6041]_ ;
  assign \new_[26187]_  = ~\new_[29931]_  & ~\new_[28883]_ ;
  assign \new_[26188]_  = ~\new_[29386]_  | ~\new_[29817]_ ;
  assign \new_[26189]_  = ~\new_[28806]_  | ~\new_[5916]_ ;
  assign \new_[26190]_  = (~\new_[29021]_  | ~\s10_data_i[8] ) & (~\new_[29709]_  | ~\s9_data_i[8] );
  assign \new_[26191]_  = ~\new_[26905]_ ;
  assign \new_[26192]_  = ~\new_[29058]_  & ~\new_[29931]_ ;
  assign \new_[26193]_  = ~\new_[27536]_ ;
  assign \new_[26194]_  = ~\new_[26900]_ ;
  assign \new_[26195]_  = ~\new_[30114]_  & ~\new_[28924]_ ;
  assign \new_[26196]_  = (~\new_[30284]_  | ~\s11_data_i[25] ) & (~\new_[29420]_  | ~\s8_data_i[25] );
  assign \new_[26197]_  = ~\new_[26885]_ ;
  assign \new_[26198]_  = ~\new_[27710]_ ;
  assign \new_[26199]_  = ~\new_[26861]_ ;
  assign \new_[26200]_  = ~\new_[26710]_ ;
  assign \new_[26201]_  = ~\new_[26862]_ ;
  assign \new_[26202]_  = ~\new_[26730]_ ;
  assign \new_[26203]_  = ~\new_[27588]_ ;
  assign \new_[26204]_  = ~\new_[26755]_ ;
  assign \new_[26205]_  = ~\new_[27555]_ ;
  assign \new_[26206]_  = ~\new_[27556]_ ;
  assign \new_[26207]_  = (~\new_[29025]_  | ~\s5_data_i[22] ) & (~\new_[30469]_  | ~\s3_data_i[22] );
  assign \new_[26208]_  = ~\new_[30212]_  & ~\new_[28887]_ ;
  assign \new_[26209]_  = ~\new_[29410]_  & ~\new_[28682]_ ;
  assign \new_[26210]_  = ~\new_[27559]_ ;
  assign \new_[26211]_  = ~\new_[29229]_  & ~\new_[30114]_ ;
  assign \new_[26212]_  = ~\new_[30688]_  & ~\new_[30070]_ ;
  assign \new_[26213]_  = ~\new_[27060]_ ;
  assign \new_[26214]_  = ~\new_[30694]_  | ~\new_[28183]_ ;
  assign \new_[26215]_  = ~\new_[27566]_ ;
  assign \new_[26216]_  = ~\new_[28078]_  | ~\new_[5966]_ ;
  assign \new_[26217]_  = ~\new_[29911]_  & ~\new_[29880]_ ;
  assign \new_[26218]_  = ~\new_[28069]_  | ~\new_[6245]_ ;
  assign \new_[26219]_  = ~\new_[29656]_  | ~\new_[28610]_ ;
  assign \new_[26220]_  = ~\new_[27835]_ ;
  assign \new_[26221]_  = (~\new_[30181]_  | ~\s14_data_i[12] ) & (~\new_[29640]_  | ~\s12_data_i[12] );
  assign \new_[26222]_  = ~\new_[29968]_  & ~\new_[29038]_ ;
  assign \new_[26223]_  = ~\new_[30525]_  | ~\new_[29360]_ ;
  assign \new_[26224]_  = ~\new_[30015]_  | ~\new_[30296]_ ;
  assign \new_[26225]_  = ~\new_[30229]_  & ~\new_[28331]_ ;
  assign \new_[26226]_  = ~\new_[27575]_ ;
  assign \new_[26227]_  = ~\new_[29927]_  | ~\new_[30727]_ ;
  assign \new_[26228]_  = ~\new_[26708]_ ;
  assign \new_[26229]_  = ~\new_[26693]_ ;
  assign \new_[26230]_  = ~\new_[26835]_ ;
  assign \new_[26231]_  = ~\new_[26593]_ ;
  assign \new_[26232]_  = (~\new_[29641]_  | ~\s14_data_i[6] ) & (~\new_[29317]_  | ~\s12_data_i[6] );
  assign \new_[26233]_  = ~\new_[26727]_ ;
  assign \new_[26234]_  = ~\new_[28837]_  | ~\new_[30022]_ ;
  assign \new_[26235]_  = ~\new_[27580]_ ;
  assign \new_[26236]_  = ~\new_[26824]_ ;
  assign \new_[26237]_  = ~\new_[29251]_  | ~\new_[5970]_ ;
  assign \new_[26238]_  = ~\new_[28039]_  | ~\new_[6065]_ ;
  assign \new_[26239]_  = ~\new_[28357]_  & ~\new_[30390]_ ;
  assign \new_[26240]_  = \new_[30764]_  | \new_[31799]_ ;
  assign \new_[26241]_  = ~\new_[26857]_ ;
  assign \new_[26242]_  = ~\new_[30034]_  | ~\new_[28023]_ ;
  assign \new_[26243]_  = \new_[28639]_  & \new_[31276]_ ;
  assign \new_[26244]_  = ~\new_[30632]_  & ~\new_[30350]_ ;
  assign \new_[26245]_  = ~\new_[29989]_  & ~\new_[30075]_ ;
  assign \new_[26246]_  = ~\new_[30222]_  | ~\new_[29019]_ ;
  assign \new_[26247]_  = ~\new_[29254]_  & ~\new_[30053]_ ;
  assign \new_[26248]_  = ~\new_[30163]_  | ~\new_[30176]_ ;
  assign \new_[26249]_  = ~\new_[28358]_  | ~\new_[6273]_ ;
  assign \new_[26250]_  = ~\new_[26664]_ ;
  assign \new_[26251]_  = ~\new_[30229]_  | ~\new_[28816]_ ;
  assign \new_[26252]_  = ~\new_[26686]_ ;
  assign \new_[26253]_  = ~\new_[28880]_  | ~\new_[29168]_ ;
  assign \new_[26254]_  = ~\new_[30211]_  & ~\new_[30114]_ ;
  assign \new_[26255]_  = ~\new_[28684]_  | ~\new_[5980]_ ;
  assign \new_[26256]_  = ~\new_[28969]_  | ~\new_[28366]_ ;
  assign \new_[26257]_  = ~\new_[29648]_  & ~\new_[29863]_ ;
  assign \new_[26258]_  = ~\new_[28057]_  | ~\new_[31422]_ ;
  assign \new_[26259]_  = ~\new_[28781]_  & ~\new_[31045]_ ;
  assign \new_[26260]_  = ~\new_[30467]_  | ~\new_[30340]_ ;
  assign \new_[26261]_  = ~\new_[30292]_  & ~\new_[30304]_ ;
  assign \new_[26262]_  = ~\new_[29839]_  & ~\new_[30245]_ ;
  assign \new_[26263]_  = ~\new_[30328]_  & ~\new_[29221]_ ;
  assign \new_[26264]_  = (~\new_[30284]_  | ~\s11_data_i[27] ) & (~\new_[29420]_  | ~\s8_data_i[27] );
  assign \new_[26265]_  = ~\new_[30764]_  | ~\new_[29996]_ ;
  assign \new_[26266]_  = ~\new_[26767]_ ;
  assign \new_[26267]_  = ~\new_[28998]_  & ~\new_[28293]_ ;
  assign \new_[26268]_  = ~\new_[30724]_  & ~\new_[6217]_ ;
  assign \new_[26269]_  = ~\new_[26762]_ ;
  assign \new_[26270]_  = ~\new_[28806]_  | ~\new_[30434]_ ;
  assign \new_[26271]_  = ~\new_[27570]_ ;
  assign \new_[26272]_  = ~\new_[30036]_  & ~\new_[29817]_ ;
  assign \new_[26273]_  = ~\new_[30665]_  | ~\new_[30000]_ ;
  assign \new_[26274]_  = ~\new_[26855]_ ;
  assign \new_[26275]_  = ~\new_[29868]_  | ~\new_[30331]_ ;
  assign \new_[26276]_  = ~\new_[26746]_ ;
  assign \new_[26277]_  = ~\new_[30604]_  & ~\new_[29019]_ ;
  assign \new_[26278]_  = ~\new_[28466]_  & ~\new_[29944]_ ;
  assign \new_[26279]_  = ~\new_[26738]_ ;
  assign \new_[26280]_  = ~\new_[27084]_ ;
  assign \new_[26281]_  = ~\new_[30785]_  | ~\new_[29251]_ ;
  assign \new_[26282]_  = ~\new_[26732]_ ;
  assign \new_[26283]_  = ~\new_[26725]_ ;
  assign \new_[26284]_  = ~\new_[30003]_  & ~\new_[30047]_ ;
  assign \new_[26285]_  = ~\new_[29987]_  | ~\new_[28873]_ ;
  assign \new_[26286]_  = ~\new_[29008]_  | ~\new_[30312]_ ;
  assign \new_[26287]_  = ~\new_[28023]_  | ~\new_[5990]_ ;
  assign \new_[26288]_  = ~\new_[30554]_  | ~\new_[29978]_ ;
  assign \new_[26289]_  = ~\new_[30078]_  & ~\new_[29040]_ ;
  assign \new_[26290]_  = \new_[29528]_  & \new_[30213]_ ;
  assign \new_[26291]_  = ~\new_[28188]_  | ~\new_[5996]_ ;
  assign \new_[26292]_  = ~\new_[27427]_  & ~\new_[30214]_ ;
  assign \new_[26293]_  = ~\new_[30072]_  & ~\new_[28850]_ ;
  assign \new_[26294]_  = ~\new_[28967]_  | ~\new_[28039]_ ;
  assign \new_[26295]_  = ~\new_[26702]_ ;
  assign \new_[26296]_  = ~\new_[28285]_  | ~\new_[5920]_ ;
  assign \new_[26297]_  = ~\new_[29902]_  & ~\new_[29181]_ ;
  assign \new_[26298]_  = ~\new_[27638]_ ;
  assign \new_[26299]_  = \new_[30287]_  | \new_[28183]_ ;
  assign \new_[26300]_  = ~\new_[28678]_  & ~\new_[28366]_ ;
  assign \new_[26301]_  = (~\new_[28842]_  | ~\s4_data_i[24] ) & (~\new_[29434]_  | ~\s0_data_i[24] );
  assign \new_[26302]_  = ~\new_[30637]_  & ~\new_[29989]_ ;
  assign \new_[26303]_  = ~\new_[26679]_ ;
  assign \new_[26304]_  = ~\new_[29669]_  | ~\new_[30006]_ ;
  assign \new_[26305]_  = ~\new_[30629]_  | ~\new_[29746]_ ;
  assign \new_[26306]_  = (~\new_[29012]_  | ~\s10_data_i[7] ) & (~\new_[29185]_  | ~\s9_data_i[7] );
  assign \new_[26307]_  = ~\new_[30029]_  & ~\new_[30213]_ ;
  assign \new_[26308]_  = ~\new_[29583]_  & ~\new_[29799]_ ;
  assign \new_[26309]_  = ~\new_[28021]_  & ~\new_[29919]_ ;
  assign \new_[26310]_  = ~\new_[30466]_  & ~\new_[28188]_ ;
  assign \new_[26311]_  = ~\new_[29817]_  | ~\new_[30707]_ ;
  assign \new_[26312]_  = ~\new_[26629]_ ;
  assign \new_[26313]_  = ~\new_[26623]_ ;
  assign \new_[26314]_  = ~\new_[26616]_ ;
  assign \new_[26315]_  = ~\new_[28732]_  | ~\new_[5993]_ ;
  assign \new_[26316]_  = ~\new_[28993]_  & ~\new_[28232]_ ;
  assign \new_[26317]_  = ~\new_[26607]_ ;
  assign \new_[26318]_  = ~\new_[30225]_  & ~\new_[28017]_ ;
  assign \new_[26319]_  = ~\new_[26578]_ ;
  assign \new_[26320]_  = ~\new_[30660]_  | ~\new_[28183]_ ;
  assign \new_[26321]_  = ~\new_[30251]_  & ~\new_[29171]_ ;
  assign \new_[26322]_  = ~\new_[27659]_ ;
  assign \new_[26323]_  = ~\new_[27971]_ ;
  assign \new_[26324]_  = ~\new_[30070]_  & ~\new_[30199]_ ;
  assign \new_[26325]_  = ~\new_[28017]_  & ~\new_[31499]_ ;
  assign \new_[26326]_  = ~\new_[30048]_  & ~\new_[30235]_ ;
  assign \new_[26327]_  = (~\new_[29631]_  | ~\s14_data_i[29] ) & (~\new_[29621]_  | ~\s12_data_i[29] );
  assign \new_[26328]_  = ~\new_[27960]_ ;
  assign \new_[26329]_  = ~\new_[27959]_ ;
  assign \new_[26330]_  = ~\new_[28121]_  | ~\new_[5982]_ ;
  assign \new_[26331]_  = ~\new_[30437]_  & ~\new_[6090]_ ;
  assign \new_[26332]_  = ~\new_[28770]_  | ~\new_[30884]_ ;
  assign \new_[26333]_  = ~\new_[27897]_  & ~\new_[28610]_ ;
  assign \new_[26334]_  = ~\new_[27923]_ ;
  assign \new_[26335]_  = (~\new_[30060]_  | ~\s7_data_i[27] ) & (~\new_[29704]_  | ~\s6_data_i[27] );
  assign \new_[26336]_  = ~\new_[29162]_  | ~\new_[28012]_ ;
  assign \new_[26337]_  = ~\new_[30203]_  & ~\new_[30268]_ ;
  assign \new_[26338]_  = ~\new_[27860]_ ;
  assign \new_[26339]_  = ~\new_[28337]_  | ~\new_[5922]_ ;
  assign \new_[26340]_  = (~\new_[30193]_  | ~\s7_data_i[15] ) & (~\new_[29298]_  | ~\s6_data_i[15] );
  assign \new_[26341]_  = ~\new_[28278]_  & ~\new_[28856]_ ;
  assign \new_[26342]_  = ~\new_[29899]_  & ~\new_[29765]_ ;
  assign \new_[26343]_  = (~\new_[30311]_  | ~\s11_data_i[7] ) & (~\new_[29636]_  | ~\s8_data_i[7] );
  assign \new_[26344]_  = ~\new_[27818]_ ;
  assign \new_[26345]_  = ~\new_[29565]_  & ~\new_[30061]_ ;
  assign \new_[26346]_  = ~\new_[27689]_ ;
  assign \new_[26347]_  = ~\new_[26651]_  & ~\new_[28012]_ ;
  assign \new_[26348]_  = ~\new_[27801]_ ;
  assign \new_[26349]_  = ~\new_[27795]_ ;
  assign \new_[26350]_  = ~\new_[30600]_  | ~\new_[30842]_ ;
  assign \new_[26351]_  = ~\new_[28397]_  & ~\new_[30754]_ ;
  assign \new_[26352]_  = ~\new_[27695]_ ;
  assign \new_[26353]_  = ~\new_[29781]_  & ~\new_[30291]_ ;
  assign \new_[26354]_  = ~\new_[30617]_  | ~\new_[28806]_ ;
  assign \new_[26355]_  = ~\new_[27754]_ ;
  assign \new_[26356]_  = ~\new_[30033]_  & ~\new_[30717]_ ;
  assign \new_[26357]_  = \new_[28188]_  & \new_[5995]_ ;
  assign \new_[26358]_  = ~\new_[30080]_  & ~\new_[30024]_ ;
  assign \new_[26359]_  = ~\new_[27680]_ ;
  assign \new_[26360]_  = ~\new_[28166]_  & ~\new_[30239]_ ;
  assign \new_[26361]_  = ~\new_[29983]_  | ~\new_[5969]_ ;
  assign \new_[26362]_  = ~\new_[26729]_ ;
  assign \new_[26363]_  = ~\new_[26775]_ ;
  assign \new_[26364]_  = ~\new_[27707]_ ;
  assign \new_[26365]_  = ~\new_[30730]_  & ~\new_[6245]_ ;
  assign \new_[26366]_  = ~\new_[26706]_ ;
  assign \new_[26367]_  = ~\new_[30028]_  & ~\new_[30526]_ ;
  assign \new_[26368]_  = ~\new_[28640]_  | ~\new_[5998]_ ;
  assign \new_[26369]_  = ~\new_[30446]_  | ~\new_[30410]_ ;
  assign \new_[26370]_  = ~\new_[30842]_  | ~\new_[30107]_ ;
  assign \new_[26371]_  = (~\new_[29976]_  | ~\s14_data_i[26] ) & (~\new_[28957]_  | ~\s12_data_i[26] );
  assign \new_[26372]_  = ~\new_[27896]_ ;
  assign \new_[26373]_  = ~\new_[27442]_ ;
  assign \new_[26374]_  = ~\new_[28658]_  & ~\new_[28250]_ ;
  assign \new_[26375]_  = ~\new_[30130]_  & ~\new_[29902]_ ;
  assign \new_[26376]_  = (~\new_[30181]_  | ~\s14_data_i[8] ) & (~\new_[29640]_  | ~\s12_data_i[8] );
  assign \new_[26377]_  = ~\new_[28245]_  | ~\new_[5986]_ ;
  assign \new_[26378]_  = ~\new_[30432]_  | ~\new_[30552]_ ;
  assign \new_[26379]_  = ~\new_[27375]_ ;
  assign \new_[26380]_  = ~\new_[30248]_  | ~\new_[29972]_ ;
  assign \new_[26381]_  = ~\new_[29199]_  & ~\new_[27787]_ ;
  assign \new_[26382]_  = ~\new_[29868]_  | ~\new_[29212]_ ;
  assign \new_[26383]_  = ~\new_[30308]_  & ~\new_[29082]_ ;
  assign \new_[26384]_  = ~\new_[28590]_  | ~\new_[29510]_ ;
  assign \new_[26385]_  = ~\new_[27720]_ ;
  assign \new_[26386]_  = ~\new_[28045]_  | ~\new_[30322]_ ;
  assign \new_[26387]_  = ~\new_[28362]_  & ~\new_[29260]_ ;
  assign \new_[26388]_  = ~\new_[28337]_  | ~\new_[30784]_ ;
  assign \new_[26389]_  = ~\new_[30221]_  | ~\new_[28250]_ ;
  assign \new_[26390]_  = ~\new_[27132]_ ;
  assign \new_[26391]_  = ~\new_[28894]_  & ~\new_[30004]_ ;
  assign \new_[26392]_  = ~\new_[29833]_  & ~\new_[29914]_ ;
  assign \new_[26393]_  = ~\new_[27098]_ ;
  assign \new_[26394]_  = ~\new_[29891]_  & ~\new_[28609]_ ;
  assign \new_[26395]_  = ~\new_[28029]_  & ~\new_[29613]_ ;
  assign \new_[26396]_  = ~\new_[30684]_  & ~\new_[30348]_ ;
  assign \new_[26397]_  = ~\new_[29015]_  | ~\new_[30628]_ ;
  assign \new_[26398]_  = ~\new_[29563]_  | ~\new_[30411]_ ;
  assign \new_[26399]_  = ~\new_[29935]_  & ~\new_[30093]_ ;
  assign \new_[26400]_  = ~\new_[27033]_ ;
  assign \new_[26401]_  = ~\new_[29763]_  & ~\new_[29360]_ ;
  assign \new_[26402]_  = ~\new_[27728]_ ;
  assign \new_[26403]_  = ~\new_[28878]_  | ~\new_[28234]_ ;
  assign \new_[26404]_  = ~\new_[26961]_ ;
  assign \new_[26405]_  = ~\new_[26995]_ ;
  assign \new_[26406]_  = ~\new_[29969]_  | ~\new_[5965]_ ;
  assign \new_[26407]_  = (~\new_[29036]_  | ~\s5_data_i[26] ) & (~\new_[30429]_  | ~\s3_data_i[26] );
  assign \new_[26408]_  = \new_[28494]_  | \new_[30688]_ ;
  assign \new_[26409]_  = ~\new_[26933]_ ;
  assign \new_[26410]_  = ~\new_[30591]_  | ~\new_[28001]_ ;
  assign \new_[26411]_  = (~\new_[30284]_  | ~\s11_data_i[18] ) & (~\new_[29420]_  | ~\s8_data_i[18] );
  assign \new_[26412]_  = ~\new_[26912]_ ;
  assign \new_[26413]_  = ~\new_[28386]_  | ~\new_[29281]_ ;
  assign \new_[26414]_  = ~\new_[28675]_  & ~\new_[29995]_ ;
  assign \new_[26415]_  = ~\new_[30542]_  & ~\new_[6049]_ ;
  assign \new_[26416]_  = ~\new_[26866]_ ;
  assign \new_[26417]_  = (~\new_[30060]_  | ~\s7_data_i[7] ) & (~\new_[29704]_  | ~\s6_data_i[7] );
  assign \new_[26418]_  = ~\new_[26743]_ ;
  assign \new_[26419]_  = ~\new_[26795]_ ;
  assign \new_[26420]_  = ~\new_[30662]_  | ~\new_[28762]_ ;
  assign \new_[26421]_  = ~\new_[27383]_ ;
  assign \new_[26422]_  = ~\new_[28007]_  | ~\new_[5999]_ ;
  assign \new_[26423]_  = ~\new_[27388]_ ;
  assign \new_[26424]_  = ~\new_[27697]_ ;
  assign \new_[26425]_  = (~\s2_data_i[17]  | ~\new_[29625]_ ) & (~\s1_data_i[17]  | ~\new_[29215]_ );
  assign \new_[26426]_  = ~\new_[26941]_ ;
  assign \new_[26427]_  = ~\new_[30656]_  & ~\new_[28215]_ ;
  assign \new_[26428]_  = ~\new_[30161]_  | ~\new_[29774]_ ;
  assign \new_[26429]_  = (~\s10_data_i[8]  | ~\new_[29749]_ ) & (~\s9_data_i[8]  | ~\new_[29034]_ );
  assign \new_[26430]_  = ~\new_[30307]_  & ~\new_[30062]_ ;
  assign \new_[26431]_  = ~\new_[26837]_ ;
  assign \new_[26432]_  = ~\new_[28355]_  | ~\new_[6005]_ ;
  assign \new_[26433]_  = ~\new_[28236]_  & ~\new_[30411]_ ;
  assign \new_[26434]_  = ~\new_[27755]_ ;
  assign \new_[26435]_  = ~\new_[27356]_ ;
  assign \new_[26436]_  = (~\new_[29021]_  | ~\s10_data_i[24] ) & (~\new_[29709]_  | ~\s9_data_i[24] );
  assign \new_[26437]_  = ~\new_[29115]_  & ~\new_[30212]_ ;
  assign \new_[26438]_  = ~\new_[28285]_  | ~\new_[28905]_ ;
  assign \new_[26439]_  = ~\new_[29898]_  & ~\new_[30159]_ ;
  assign \new_[26440]_  = ~\new_[29826]_  & ~\new_[29219]_ ;
  assign \new_[26441]_  = (~\new_[30193]_  | ~\s7_data_i[18] ) & (~\new_[29298]_  | ~\s6_data_i[18] );
  assign \new_[26442]_  = ~\new_[30442]_  & ~\new_[6093]_ ;
  assign \new_[26443]_  = ~\new_[28027]_  & ~\new_[28234]_ ;
  assign \new_[26444]_  = \new_[29482]_  & \new_[28806]_ ;
  assign \new_[26445]_  = (~\s10_data_i[25]  | ~\new_[29749]_ ) & (~\s9_data_i[25]  | ~\new_[29034]_ );
  assign \new_[26446]_  = ~\new_[26925]_ ;
  assign \new_[26447]_  = ~\new_[27928]_ ;
  assign \new_[26448]_  = (~\new_[29534]_  | ~\s5_data_i[12] ) & (~\new_[29579]_  | ~\s3_data_i[12] );
  assign \new_[26449]_  = ~\new_[27772]_ ;
  assign \new_[26450]_  = ~\new_[27696]_ ;
  assign \new_[26451]_  = ~\new_[26799]_ ;
  assign \new_[26452]_  = ~\new_[28783]_  | ~\new_[5912]_ ;
  assign \new_[26453]_  = ~\new_[30094]_  & ~\new_[29931]_ ;
  assign \new_[26454]_  = ~\new_[26786]_ ;
  assign \new_[26455]_  = ~\new_[28125]_  & ~\new_[6066]_ ;
  assign \new_[26456]_  = ~\new_[26759]_ ;
  assign \new_[26457]_  = ~\new_[28793]_  | ~\new_[5918]_ ;
  assign \new_[26458]_  = (~\new_[29025]_  | ~\s5_data_i[9] ) & (~\new_[30469]_  | ~\s3_data_i[9] );
  assign \new_[26459]_  = ~\new_[29210]_  | ~\new_[30205]_ ;
  assign \new_[26460]_  = ~\new_[28149]_  | ~\new_[5911]_ ;
  assign \new_[26461]_  = (~\new_[30060]_  | ~\s7_data_i[10] ) & (~\new_[29704]_  | ~\s6_data_i[10] );
  assign \new_[26462]_  = ~\new_[26711]_ ;
  assign \new_[26463]_  = ~\new_[27792]_ ;
  assign \new_[26464]_  = ~\new_[27794]_ ;
  assign \new_[26465]_  = ~\new_[28516]_  & ~\new_[31423]_ ;
  assign \new_[26466]_  = ~\new_[26677]_ ;
  assign \new_[26467]_  = ~\new_[30201]_  & ~\new_[30444]_ ;
  assign \new_[26468]_  = \new_[28007]_  & \new_[6000]_ ;
  assign \new_[26469]_  = ~\new_[28791]_  | ~\new_[30884]_ ;
  assign \new_[26470]_  = ~\new_[29967]_  | ~\new_[30627]_ ;
  assign \new_[26471]_  = ~\new_[30205]_  | ~\new_[29972]_ ;
  assign \new_[26472]_  = (~\new_[29025]_  | ~\s5_data_i[24] ) & (~\new_[30469]_  | ~\s3_data_i[24] );
  assign \new_[26473]_  = (~\new_[30060]_  | ~\s7_data_i[31] ) & (~\new_[29704]_  | ~\s6_data_i[31] );
  assign \new_[26474]_  = ~\new_[28787]_  | ~\new_[31045]_ ;
  assign \new_[26475]_  = (~\new_[30311]_  | ~\s11_data_i[12] ) & (~\new_[29636]_  | ~\s8_data_i[12] );
  assign \new_[26476]_  = ~\new_[30032]_  & ~\new_[6080]_ ;
  assign \new_[26477]_  = ~\new_[27852]_ ;
  assign \new_[26478]_  = (~\new_[29045]_  | ~\s10_data_i[12] ) & (~\new_[29951]_  | ~\s9_data_i[12] );
  assign \new_[26479]_  = ~\new_[27690]_ ;
  assign \new_[26480]_  = ~\new_[27894]_ ;
  assign \new_[26481]_  = (~\new_[29149]_  | ~\s4_data_i[24] ) & (~\new_[29651]_  | ~\s0_data_i[24] );
  assign \new_[26482]_  = ~\new_[28705]_  | ~\new_[5909]_ ;
  assign \new_[26483]_  = (~\new_[29025]_  | ~\s5_data_i[27] ) & (~\new_[30469]_  | ~\s3_data_i[27] );
  assign \new_[26484]_  = ~\new_[28789]_  & ~\new_[31406]_ ;
  assign \new_[26485]_  = ~\new_[27816]_ ;
  assign \new_[26486]_  = ~\new_[26977]_ ;
  assign \new_[26487]_  = ~\new_[26921]_ ;
  assign \new_[26488]_  = \new_[28558]_  & \new_[30009]_ ;
  assign \new_[26489]_  = ~\new_[27821]_ ;
  assign \new_[26490]_  = (~\new_[30227]_  | ~\s10_data_i[8] ) & (~\new_[29706]_  | ~\s9_data_i[8] );
  assign \new_[26491]_  = ~\new_[26851]_ ;
  assign \new_[26492]_  = (~\new_[30181]_  | ~\s14_data_i[13] ) & (~\new_[29640]_  | ~\s12_data_i[13] );
  assign \new_[26493]_  = ~\new_[27372]_ ;
  assign \new_[26494]_  = ~\new_[30296]_  | ~\new_[28069]_ ;
  assign \new_[26495]_  = (~\new_[29021]_  | ~\s10_data_i[6] ) & (~\new_[29709]_  | ~\s9_data_i[6] );
  assign \new_[26496]_  = ~\new_[26582]_ ;
  assign \new_[26497]_  = (~\new_[29149]_  | ~\s4_data_i[9] ) & (~\new_[29651]_  | ~\s0_data_i[9] );
  assign \new_[26498]_  = ~\new_[27814]_ ;
  assign \new_[26499]_  = ~\new_[28776]_  | ~\new_[6208]_ ;
  assign \new_[26500]_  = (~\new_[29045]_  | ~\s10_data_i[13] ) & (~\new_[29951]_  | ~\s9_data_i[13] );
  assign \new_[26501]_  = ~\new_[28778]_  | ~\new_[6084]_ ;
  assign \new_[26502]_  = ~\new_[29400]_  | ~\new_[28664]_ ;
  assign \new_[26503]_  = ~\new_[27902]_ ;
  assign \new_[26504]_  = ~\new_[27682]_ ;
  assign \new_[26505]_  = (~\new_[30193]_  | ~\s7_data_i[14] ) & (~\new_[29298]_  | ~\s6_data_i[14] );
  assign \new_[26506]_  = ~\new_[29496]_  | ~\new_[28796]_ ;
  assign \new_[26507]_  = ~\new_[26781]_ ;
  assign \new_[26508]_  = ~\new_[28435]_  | ~\new_[31712]_ ;
  assign \new_[26509]_  = ~\new_[30438]_  & ~\new_[28337]_ ;
  assign \new_[26510]_  = ~\new_[28013]_  | ~\new_[5923]_ ;
  assign \new_[26511]_  = ~\new_[28533]_  & ~\new_[29370]_ ;
  assign \new_[26512]_  = (~\new_[30200]_  | ~\s11_data_i[0] ) & (~\new_[29428]_  | ~\s8_data_i[0] );
  assign \new_[26513]_  = ~\new_[29028]_  & ~\new_[28409]_ ;
  assign \new_[26514]_  = (~\new_[29976]_  | ~\s14_data_i[20] ) & (~\new_[28957]_  | ~\s12_data_i[20] );
  assign \new_[26515]_  = ~\new_[30040]_  & ~\new_[29908]_ ;
  assign \new_[26516]_  = (~\s10_data_i[17]  | ~\new_[29749]_ ) & (~\s9_data_i[17]  | ~\new_[29034]_ );
  assign \new_[26517]_  = ~\new_[29070]_  | ~\new_[28214]_ ;
  assign \new_[26518]_  = ~\new_[28425]_  & ~\new_[29565]_ ;
  assign \new_[26519]_  = (~\new_[30181]_  | ~\s14_data_i[2] ) & (~\new_[29640]_  | ~\s12_data_i[2] );
  assign \new_[26520]_  = ~\new_[27679]_ ;
  assign \new_[26521]_  = ~\new_[26850]_ ;
  assign \new_[26522]_  = ~\new_[28229]_  | ~\new_[29996]_ ;
  assign \new_[26523]_  = (~\new_[29012]_  | ~\s10_data_i[11] ) & (~\new_[29185]_  | ~\s9_data_i[11] );
  assign \new_[26524]_  = ~\new_[27857]_ ;
  assign \new_[26525]_  = ~\new_[32344]_ ;
  assign \new_[26526]_  = (~\new_[30060]_  | ~\s7_data_i[2] ) & (~\new_[29704]_  | ~\s6_data_i[2] );
  assign \new_[26527]_  = (~\s5_data_i[18]  | ~\new_[29649]_ ) & (~\s3_data_i[18]  | ~\new_[29035]_ );
  assign \new_[26528]_  = ~\new_[27871]_ ;
  assign \new_[26529]_  = ~\new_[28011]_  | ~\new_[31403]_ ;
  assign \new_[26530]_  = ~\new_[27701]_ ;
  assign \new_[26531]_  = ~\new_[28918]_  & ~\new_[28362]_ ;
  assign \new_[26532]_  = ~\new_[29553]_  | ~\new_[30081]_ ;
  assign \new_[26533]_  = ~\new_[26789]_ ;
  assign \new_[26534]_  = ~\new_[27925]_ ;
  assign \new_[26535]_  = ~\new_[27675]_ ;
  assign \new_[26536]_  = ~\new_[27910]_ ;
  assign \new_[26537]_  = (~\new_[30181]_  | ~\s14_data_i[17] ) & (~\new_[29640]_  | ~\s12_data_i[17] );
  assign \new_[26538]_  = ~\new_[30710]_  | ~\new_[29299]_ ;
  assign \new_[26539]_  = (~\new_[30060]_  | ~\s7_data_i[17] ) & (~\new_[29704]_  | ~\s6_data_i[17] );
  assign \new_[26540]_  = ~\new_[26608]_ ;
  assign \new_[26541]_  = ~\new_[27674]_ ;
  assign \new_[26542]_  = ~\new_[27957]_ ;
  assign \new_[26543]_  = ~\new_[28331]_  & ~\new_[30508]_ ;
  assign \new_[26544]_  = (~\new_[29710]_  | ~\s10_data_i[11] ) & (~\new_[29024]_  | ~\s9_data_i[11] );
  assign \new_[26545]_  = ~\new_[27291]_ ;
  assign \new_[26546]_  = (~\new_[30311]_  | ~\s11_data_i[18] ) & (~\new_[29636]_  | ~\s8_data_i[18] );
  assign \new_[26547]_  = ~\new_[27672]_ ;
  assign \new_[26548]_  = ~\new_[28020]_  & ~\new_[29139]_ ;
  assign \new_[26549]_  = \new_[28009]_  & \new_[31690]_ ;
  assign \new_[26550]_  = ~\new_[30566]_  & ~\new_[29853]_ ;
  assign \new_[26551]_  = \new_[28476]_  & \new_[29168]_ ;
  assign \new_[26552]_  = ~\new_[30640]_  & ~\new_[30253]_ ;
  assign \new_[26553]_  = ~\new_[28700]_  & ~\new_[30771]_ ;
  assign \new_[26554]_  = ~\new_[27940]_ ;
  assign \new_[26555]_  = (~\new_[29045]_  | ~\s10_data_i[18] ) & (~\new_[29951]_  | ~\s9_data_i[18] );
  assign \new_[26556]_  = ~\new_[30747]_  & ~\new_[30633]_ ;
  assign \new_[26557]_  = ~\new_[28470]_  & ~\new_[28815]_ ;
  assign \new_[26558]_  = (~\new_[30031]_  | ~\s7_data_i[23] ) & (~\new_[29052]_  | ~\s6_data_i[23] );
  assign \new_[26559]_  = (~\s10_data_i[27]  | ~\new_[29749]_ ) & (~\s9_data_i[27]  | ~\new_[29034]_ );
  assign \new_[26560]_  = ~\new_[28818]_  & ~\new_[29791]_ ;
  assign \new_[26561]_  = ~\new_[26809]_ ;
  assign \new_[26562]_  = \new_[29477]_  & \new_[28337]_ ;
  assign \new_[26563]_  = ~\new_[29746]_ ;
  assign \new_[26564]_  = ~\new_[26899]_ ;
  assign \new_[26565]_  = \new_[29128]_  | \new_[30273]_ ;
  assign \new_[26566]_  = (~\new_[29045]_  | ~\s10_data_i[9] ) & (~\new_[29951]_  | ~\s9_data_i[9] );
  assign \new_[26567]_  = (~\new_[29631]_  | ~\s14_data_i[30] ) & (~\new_[29621]_  | ~\s12_data_i[30] );
  assign \new_[26568]_  = ~\new_[30053]_  & ~\new_[28939]_ ;
  assign \new_[26569]_  = (~\new_[30181]_  | ~\s14_data_i[19] ) & (~\new_[29640]_  | ~\s12_data_i[19] );
  assign \new_[26570]_  = \new_[28009]_  & \new_[31423]_ ;
  assign \new_[26571]_  = ~\new_[27964]_ ;
  assign \new_[26572]_  = ~\new_[27954]_ ;
  assign \new_[26573]_  = ~\new_[30582]_  | ~\new_[30296]_ ;
  assign \new_[26574]_  = (~\new_[29953]_  | ~\s11_data_i[26] ) & (~\new_[29627]_  | ~\s8_data_i[26] );
  assign \new_[26575]_  = ~\new_[26660]_  & ~\new_[28121]_ ;
  assign \new_[26576]_  = ~\new_[26894]_ ;
  assign \new_[26577]_  = (~\new_[30085]_  | ~\s2_data_i[2] ) & (~\new_[30108]_  | ~\s1_data_i[2] );
  assign \new_[26578]_  = ~\new_[30173]_  & ~\new_[28930]_ ;
  assign \new_[26579]_  = (~\new_[29961]_  | ~\s4_data_i[26] ) & (~\new_[29819]_  | ~\s0_data_i[26] );
  assign \new_[26580]_  = ~\new_[27978]_ ;
  assign \new_[26581]_  = ~\new_[30437]_  | ~\new_[29184]_ ;
  assign \new_[26582]_  = ~\new_[29714]_  | ~\new_[5918]_ ;
  assign \new_[26583]_  = ~\new_[27981]_ ;
  assign \new_[26584]_  = (~\new_[30189]_  | ~\s2_data_i[22] ) & (~\new_[30195]_  | ~\s1_data_i[22] );
  assign \new_[26585]_  = ~\new_[30169]_  | ~\new_[29452]_ ;
  assign \new_[26586]_  = ~\new_[27988]_ ;
  assign \new_[26587]_  = ~\new_[27989]_ ;
  assign \new_[26588]_  = (~\new_[29961]_  | ~\s4_data_i[10] ) & (~\new_[29819]_  | ~\s0_data_i[10] );
  assign \new_[26589]_  = ~\new_[29368]_  & ~\new_[5918]_ ;
  assign \new_[26590]_  = ~\new_[29175]_  | ~\new_[30390]_ ;
  assign \new_[26591]_  = ~\new_[29582]_  | ~\new_[30016]_ ;
  assign \new_[26592]_  = ~\new_[29192]_  | ~\new_[29260]_ ;
  assign \new_[26593]_  = ~\new_[30325]_  | ~\new_[30586]_ ;
  assign \new_[26594]_  = ~\new_[27993]_ ;
  assign \new_[26595]_  = (~\new_[29788]_  | ~\s2_data_i[8] ) & (~\new_[30357]_  | ~\s1_data_i[8] );
  assign \new_[26596]_  = ~\new_[30024]_ ;
  assign \new_[26597]_  = ~\new_[30139]_  & ~\new_[29019]_ ;
  assign \new_[26598]_  = \new_[29742]_  | \new_[30952]_ ;
  assign \new_[26599]_  = (~\new_[29807]_  | ~\s14_data_i[19] ) & (~\new_[30626]_  | ~\s12_data_i[19] );
  assign \new_[26600]_  = \new_[28820]_  & \new_[30730]_ ;
  assign \new_[26601]_  = ~\new_[28690]_ ;
  assign \new_[26602]_  = \new_[29040]_  & \new_[6088]_ ;
  assign \new_[26603]_  = ~\new_[28314]_ ;
  assign \new_[26604]_  = ~\new_[29162]_  & ~\new_[29965]_ ;
  assign \new_[26605]_  = (~\new_[30189]_  | ~\s2_data_i[28] ) & (~\new_[30195]_  | ~\s1_data_i[28] );
  assign \new_[26606]_  = (~\new_[29948]_  | ~\s5_data_i[0] ) & (~\new_[29947]_  | ~\s3_data_i[0] );
  assign \new_[26607]_  = ~\new_[30728]_  | ~\new_[28944]_ ;
  assign \new_[26608]_  = ~\new_[29719]_  & ~\new_[5913]_ ;
  assign \new_[26609]_  = ~\new_[28308]_ ;
  assign \new_[26610]_  = ~\new_[28310]_ ;
  assign \new_[26611]_  = \new_[29158]_  & \new_[29159]_ ;
  assign \new_[26612]_  = \new_[29723]_  & \new_[6038]_ ;
  assign \new_[26613]_  = ~\new_[29150]_  | ~\new_[5973]_ ;
  assign \new_[26614]_  = ~\new_[29168]_  | ~\new_[29692]_ ;
  assign \new_[26615]_  = ~\new_[28202]_ ;
  assign \new_[26616]_  = ~\new_[30608]_  | ~\new_[29598]_ ;
  assign \new_[26617]_  = ~\new_[29421]_  & ~\new_[29758]_ ;
  assign \new_[26618]_  = ~\new_[29502]_  | ~\new_[30508]_ ;
  assign \new_[26619]_  = (~\new_[29949]_  | ~\s10_data_i[30] ) & (~\new_[29905]_  | ~\s9_data_i[30] );
  assign \new_[26620]_  = ~\new_[28006]_ ;
  assign \new_[26621]_  = ~\new_[28008]_ ;
  assign \new_[26622]_  = (~\new_[29788]_  | ~\s2_data_i[13] ) & (~\new_[30357]_  | ~\s1_data_i[13] );
  assign \new_[26623]_  = ~\new_[29639]_  | ~\new_[29404]_ ;
  assign \new_[26624]_  = ~\new_[30031]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[26625]_  = (~\new_[30013]_  | ~\s2_data_i[4] ) & (~\new_[29769]_  | ~\s1_data_i[4] );
  assign \new_[26626]_  = ~\new_[28010]_ ;
  assign \new_[26627]_  = ~\new_[28866]_ ;
  assign \new_[26628]_  = ~\new_[28688]_ ;
  assign \new_[26629]_  = ~\new_[30302]_  & ~\new_[28245]_ ;
  assign \new_[26630]_  = ~\new_[28014]_ ;
  assign \new_[26631]_  = ~\new_[28018]_ ;
  assign \new_[26632]_  = ~\new_[28016]_ ;
  assign \new_[26633]_  = ~\new_[28025]_ ;
  assign \new_[26634]_  = ~\new_[29039]_  | ~\new_[6066]_ ;
  assign \new_[26635]_  = ~\new_[28024]_ ;
  assign \new_[26636]_  = ~\new_[28544]_ ;
  assign \new_[26637]_  = ~\new_[28026]_ ;
  assign \new_[26638]_  = ~\new_[28888]_ ;
  assign \new_[26639]_  = ~\new_[29739]_  & ~\new_[5997]_ ;
  assign \new_[26640]_  = ~\new_[28900]_  | ~\new_[31043]_ ;
  assign \new_[26641]_  = ~\new_[32169]_ ;
  assign \new_[26642]_  = ~\new_[28863]_  | ~\new_[31406]_ ;
  assign \new_[26643]_  = ~\new_[28730]_ ;
  assign \new_[26644]_  = ~\new_[28040]_ ;
  assign \new_[26645]_  = \new_[29575]_  | \new_[31479]_ ;
  assign \new_[26646]_  = (~\new_[29788]_  | ~\s2_data_i[23] ) & (~\new_[30357]_  | ~\s1_data_i[23] );
  assign \new_[26647]_  = ~\new_[31232]_  & ~\new_[31906]_ ;
  assign \new_[26648]_  = ~\new_[29807]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[26649]_  = \new_[29396]_  | \new_[31043]_ ;
  assign \new_[26650]_  = ~\new_[28042]_ ;
  assign \new_[26651]_  = ~\new_[29162]_ ;
  assign \new_[26652]_  = ~\new_[28046]_ ;
  assign \new_[26653]_  = ~\new_[30620]_  & ~\new_[30115]_ ;
  assign \new_[26654]_  = ~\new_[28728]_ ;
  assign \new_[26655]_  = ~\new_[29360]_ ;
  assign \new_[26656]_  = (~\new_[30166]_  | ~\s14_data_i[14] ) & (~\new_[30298]_  | ~\s12_data_i[14] );
  assign \new_[26657]_  = ~\new_[29168]_ ;
  assign \new_[26658]_  = (~\new_[30189]_  | ~\s2_data_i[3] ) & (~\new_[30195]_  | ~\s1_data_i[3] );
  assign \new_[26659]_  = \new_[29221]_  & \new_[5980]_ ;
  assign \new_[26660]_  = ~\new_[29171]_ ;
  assign \new_[26661]_  = ~\new_[28985]_  | ~\new_[30316]_ ;
  assign \new_[26662]_  = ~\new_[28066]_ ;
  assign \new_[26663]_  = ~\new_[30193]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[26664]_  = ~\new_[28908]_  | ~\new_[30245]_ ;
  assign \new_[26665]_  = \new_[29191]_  | \new_[30884]_ ;
  assign \new_[26666]_  = ~\new_[30113]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[26667]_  = ~\new_[30491]_  | ~\new_[6192]_ ;
  assign \new_[26668]_  = ~\new_[28182]_ ;
  assign \new_[26669]_  = ~\new_[29725]_  | ~\new_[31539]_ ;
  assign \new_[26670]_  = ~\new_[28876]_  | ~\new_[5921]_ ;
  assign \new_[26671]_  = (~\new_[29949]_  | ~\s10_data_i[24] ) & (~\new_[29905]_  | ~\s9_data_i[24] );
  assign \new_[26672]_  = \new_[29723]_  & \new_[31665]_ ;
  assign \new_[26673]_  = ~\new_[30693]_  & ~\new_[30228]_ ;
  assign \new_[26674]_  = ~\new_[29861]_  & ~\new_[28933]_ ;
  assign \new_[26675]_  = ~\new_[28835]_  | ~\new_[30268]_ ;
  assign \new_[26676]_  = \new_[29458]_  & \new_[30582]_ ;
  assign \new_[26677]_  = ~\new_[28946]_  | ~\new_[6040]_ ;
  assign \new_[26678]_  = (~\new_[30113]_  | ~\s2_data_i[7] ) & (~\new_[30124]_  | ~\s1_data_i[7] );
  assign \new_[26679]_  = ~\new_[28270]_  & ~\new_[28114]_ ;
  assign \new_[26680]_  = ~\new_[28820]_  | ~\new_[30726]_ ;
  assign \new_[26681]_  = ~\new_[6246]_  | ~\new_[30730]_  | ~\new_[30020]_ ;
  assign \new_[26682]_  = ~\new_[28645]_ ;
  assign \new_[26683]_  = ~\new_[28082]_ ;
  assign \new_[26684]_  = ~\new_[32267]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[26685]_  = ~\new_[29271]_  | ~\new_[30246]_ ;
  assign \new_[26686]_  = ~\new_[29750]_  & ~\new_[30434]_ ;
  assign \new_[26687]_  = (~\new_[29846]_  | ~\s2_data_i[1] ) & (~\new_[30001]_  | ~\s1_data_i[1] );
  assign \new_[26688]_  = ~\new_[28085]_ ;
  assign \new_[26689]_  = \new_[29053]_  & \m6_addr_i[28] ;
  assign \new_[26690]_  = ~\new_[29788]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[26691]_  = (~\new_[29788]_  | ~\s2_data_i[25] ) & (~\new_[30357]_  | ~\s1_data_i[25] );
  assign \new_[26692]_  = ~\new_[30088]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[26693]_  = ~\new_[30242]_  | ~\new_[29122]_ ;
  assign \new_[26694]_  = (~\new_[29876]_  | ~\s11_data_i[23] ) & (~\new_[30341]_  | ~\s8_data_i[23] );
  assign \new_[26695]_  = ~\new_[28391]_ ;
  assign \new_[26696]_  = (~\new_[30166]_  | ~\s14_data_i[30] ) & (~\new_[30298]_  | ~\s12_data_i[30] );
  assign \new_[26697]_  = ~\new_[29961]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[26698]_  = ~\new_[28100]_ ;
  assign \new_[26699]_  = ~\new_[28723]_ ;
  assign \new_[26700]_  = (~\new_[30189]_  | ~\s2_data_i[15] ) & (~\new_[30195]_  | ~\s1_data_i[15] );
  assign \new_[26701]_  = ~\new_[28103]_ ;
  assign \new_[26702]_  = ~\new_[29212]_  | ~\new_[5976]_ ;
  assign \new_[26703]_  = ~\new_[29015]_  | ~\new_[6059]_ ;
  assign \new_[26704]_  = ~\new_[29564]_  | ~\new_[29226]_ ;
  assign \new_[26705]_  = ~\new_[28106]_ ;
  assign \new_[26706]_  = ~\new_[30130]_  | ~\new_[29602]_ ;
  assign \new_[26707]_  = ~\new_[30702]_  | ~\new_[30751]_ ;
  assign \new_[26708]_  = ~\new_[30033]_  | ~\new_[30519]_ ;
  assign \new_[26709]_  = ~\new_[29168]_  | ~\new_[5971]_ ;
  assign \new_[26710]_  = ~\new_[29633]_  | ~\new_[30304]_ ;
  assign \new_[26711]_  = ~\new_[29396]_  & ~\new_[6084]_ ;
  assign \new_[26712]_  = ~\new_[30556]_  | ~\new_[29647]_ ;
  assign \new_[26713]_  = ~\new_[28262]_ ;
  assign \new_[26714]_  = ~\new_[28282]_ ;
  assign \new_[26715]_  = ~\new_[29008]_  | ~\new_[5898]_ ;
  assign \new_[26716]_  = ~\new_[30026]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[26717]_  = ~\new_[30107]_  | ~\new_[30491]_ ;
  assign \new_[26718]_  = ~\new_[30284]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[26719]_  = ~\new_[28246]_ ;
  assign \new_[26720]_  = (~\new_[30013]_  | ~\s2_data_i[3] ) & (~\new_[29769]_  | ~\s1_data_i[3] );
  assign \new_[26721]_  = ~\new_[29571]_  | ~\new_[30147]_ ;
  assign \new_[26722]_  = (~\new_[29949]_  | ~\s10_data_i[25] ) & (~\new_[29905]_  | ~\s9_data_i[25] );
  assign \new_[26723]_  = \new_[29063]_  | \new_[6066]_ ;
  assign \new_[26724]_  = \new_[29701]_  & \new_[5929]_ ;
  assign \new_[26725]_  = ~\new_[30002]_  & ~\new_[28967]_ ;
  assign \new_[26726]_  = ~\new_[28120]_ ;
  assign \new_[26727]_  = ~\new_[28844]_  | ~\new_[30267]_ ;
  assign \new_[26728]_  = ~\new_[29118]_  | ~\new_[30764]_ ;
  assign \new_[26729]_  = ~\new_[30068]_  & ~\new_[29197]_ ;
  assign \new_[26730]_  = ~\new_[30248]_  & ~\new_[30715]_ ;
  assign \new_[26731]_  = ~\new_[28122]_ ;
  assign \new_[26732]_  = ~\new_[29868]_  & ~\new_[28909]_ ;
  assign \new_[26733]_  = ~\new_[29272]_  & ~\new_[28985]_ ;
  assign \new_[26734]_  = ~\new_[28306]_ ;
  assign \new_[26735]_  = ~\new_[30202]_  | ~\new_[29228]_ ;
  assign \new_[26736]_  = ~\new_[28976]_  | ~\new_[29425]_ ;
  assign \new_[26737]_  = (~\new_[29963]_  | ~\s4_data_i[3] ) & (~\new_[30481]_  | ~\s0_data_i[3] );
  assign \new_[26738]_  = ~\new_[29189]_  | ~\new_[30024]_ ;
  assign \new_[26739]_  = (~\new_[30113]_  | ~\s2_data_i[8] ) & (~\new_[30124]_  | ~\s1_data_i[8] );
  assign \new_[26740]_  = ~\new_[28525]_ ;
  assign \new_[26741]_  = ~\new_[29174]_  | ~\new_[28828]_ ;
  assign \new_[26742]_  = ~\new_[28135]_ ;
  assign \new_[26743]_  = ~\new_[29544]_  & ~\new_[30497]_ ;
  assign \new_[26744]_  = ~\new_[28583]_ ;
  assign \new_[26745]_  = ~\new_[28859]_  & ~\new_[29184]_ ;
  assign \new_[26746]_  = ~\new_[30661]_  | ~\new_[29299]_ ;
  assign \new_[26747]_  = (~\new_[29823]_  | ~\s7_data_i[31] ) & (~\new_[29954]_  | ~\s6_data_i[31] );
  assign \new_[26748]_  = ~\new_[28896]_  & ~\new_[5912]_ ;
  assign \new_[26749]_  = (~\new_[30088]_  | ~\s2_data_i[9] ) & (~\new_[29779]_  | ~\s1_data_i[9] );
  assign \new_[26750]_  = ~\new_[29922]_  | ~\new_[28834]_ ;
  assign \new_[26751]_  = ~\new_[28877]_  | ~\new_[29139]_ ;
  assign \new_[26752]_  = ~\new_[28483]_ ;
  assign \new_[26753]_  = ~\new_[29221]_  | ~\new_[5979]_ ;
  assign \new_[26754]_  = ~\new_[28161]_ ;
  assign \new_[26755]_  = ~\new_[28911]_  | ~\new_[29914]_ ;
  assign \new_[26756]_  = (~\new_[30189]_  | ~\s2_data_i[1] ) & (~\new_[30195]_  | ~\s1_data_i[1] );
  assign \new_[26757]_  = ~\new_[30142]_  | ~\new_[29508]_ ;
  assign \new_[26758]_  = (~\new_[30088]_  | ~\s2_data_i[0] ) & (~\new_[29779]_  | ~\s1_data_i[0] );
  assign \new_[26759]_  = \new_[28949]_  & \new_[31724]_ ;
  assign \new_[26760]_  = ~\new_[28169]_ ;
  assign \new_[26761]_  = ~\new_[28175]_ ;
  assign \new_[26762]_  = ~\new_[30044]_  | ~\new_[29104]_ ;
  assign \new_[26763]_  = ~\new_[28760]_ ;
  assign \new_[26764]_  = ~\new_[28518]_ ;
  assign \new_[26765]_  = ~\new_[29007]_  | ~\new_[5927]_ ;
  assign \new_[26766]_  = ~\new_[29645]_  & ~\new_[6038]_ ;
  assign \new_[26767]_  = ~\new_[29595]_  & ~\new_[28905]_ ;
  assign \new_[26768]_  = ~\new_[29994]_  | ~\new_[29404]_ ;
  assign \new_[26769]_  = ~\new_[29590]_  | ~\new_[30355]_ ;
  assign \new_[26770]_  = (~\new_[30113]_  | ~\s2_data_i[9] ) & (~\new_[30124]_  | ~\s1_data_i[9] );
  assign \new_[26771]_  = ~\new_[28292]_ ;
  assign \new_[26772]_  = (~\new_[30088]_  | ~\s2_data_i[19] ) & (~\new_[29779]_  | ~\s1_data_i[19] );
  assign \new_[26773]_  = (~\new_[30088]_  | ~\s2_data_i[1] ) & (~\new_[29779]_  | ~\s1_data_i[1] );
  assign \new_[26774]_  = ~\new_[28192]_ ;
  assign \new_[26775]_  = ~\new_[29966]_  & ~\new_[29003]_ ;
  assign \new_[26776]_  = ~\new_[28515]_ ;
  assign \new_[26777]_  = (~\new_[30189]_  | ~\s2_data_i[10] ) & (~\new_[30195]_  | ~\s1_data_i[10] );
  assign \new_[26778]_  = (~\new_[29846]_  | ~\s2_data_i[25] ) & (~\new_[30001]_  | ~\s1_data_i[25] );
  assign \new_[26779]_  = ~\new_[29608]_  | ~\new_[30084]_ ;
  assign \new_[26780]_  = (~\new_[30085]_  | ~\s2_data_i[18] ) & (~\new_[30108]_  | ~\s1_data_i[18] );
  assign \new_[26781]_  = ~\new_[29246]_  | ~\new_[31870]_ ;
  assign \new_[26782]_  = ~\new_[29333]_  | ~\new_[29557]_ ;
  assign \new_[26783]_  = (~\new_[30166]_  | ~\s14_data_i[27] ) & (~\new_[30298]_  | ~\s12_data_i[27] );
  assign \new_[26784]_  = ~\new_[30559]_  | ~\new_[6184]_ ;
  assign \new_[26785]_  = (~\new_[30085]_  | ~\s2_data_i[8] ) & (~\new_[30108]_  | ~\s1_data_i[8] );
  assign \new_[26786]_  = ~\new_[29737]_  & ~\new_[6040]_ ;
  assign \new_[26787]_  = (~\new_[29846]_  | ~\s2_data_i[31] ) & (~\new_[30001]_  | ~\s1_data_i[31] );
  assign \new_[26788]_  = \new_[29573]_  & \new_[28939]_ ;
  assign \new_[26789]_  = ~\new_[29134]_  & ~\new_[31406]_ ;
  assign \new_[26790]_  = ~\new_[30208]_  | ~\new_[29557]_ ;
  assign \new_[26791]_  = (~\new_[30189]_  | ~\s2_data_i[30] ) & (~\new_[30195]_  | ~\s1_data_i[30] );
  assign \new_[26792]_  = (~\new_[30088]_  | ~\s2_data_i[30] ) & (~\new_[29779]_  | ~\s1_data_i[30] );
  assign \new_[26793]_  = ~\new_[29006]_  | ~\new_[6074]_ ;
  assign \new_[26794]_  = ~\new_[29853]_  & ~\new_[30230]_ ;
  assign \new_[26795]_  = ~\new_[29212]_  | ~\new_[30331]_ ;
  assign \new_[26796]_  = (~\new_[29948]_  | ~\s5_data_i[29] ) & (~\new_[29947]_  | ~\s3_data_i[29] );
  assign \new_[26797]_  = (~\new_[30166]_  | ~\s14_data_i[18] ) & (~\new_[30298]_  | ~\s12_data_i[18] );
  assign \new_[26798]_  = \new_[29082]_  & \new_[5986]_ ;
  assign \new_[26799]_  = ~\new_[28952]_  | ~\new_[6208]_ ;
  assign \new_[26800]_  = ~\new_[28209]_ ;
  assign \new_[26801]_  = ~\new_[29725]_  | ~\new_[31148]_ ;
  assign \new_[26802]_  = (~\new_[30131]_  | ~\s7_data_i[27] ) & (~\new_[29939]_  | ~\s6_data_i[27] );
  assign \new_[26803]_  = ~\new_[29217]_  & ~\new_[30202]_ ;
  assign \new_[26804]_  = ~\new_[30569]_  & ~\new_[29064]_ ;
  assign \new_[26805]_  = (~\new_[29963]_  | ~\s4_data_i[29] ) & (~\new_[30481]_  | ~\s0_data_i[29] );
  assign \new_[26806]_  = ~\new_[28578]_ ;
  assign \new_[26807]_  = ~\new_[28227]_ ;
  assign \new_[26808]_  = (~\new_[29788]_  | ~\s2_data_i[30] ) & (~\new_[30357]_  | ~\s1_data_i[30] );
  assign \new_[26809]_  = ~\new_[29086]_  | ~\new_[30239]_ ;
  assign \new_[26810]_  = (~\new_[30085]_  | ~\s2_data_i[20] ) & (~\new_[30108]_  | ~\s1_data_i[20] );
  assign \new_[26811]_  = ~\new_[28672]_ ;
  assign \new_[26812]_  = ~\new_[30277]_  | ~\new_[28964]_ ;
  assign \new_[26813]_  = ~\new_[29333]_  & ~\new_[30208]_ ;
  assign \new_[26814]_  = ~\new_[29972]_  | ~\new_[29537]_ ;
  assign \new_[26815]_  = ~\new_[29922]_  & ~\new_[29122]_ ;
  assign \new_[26816]_  = ~\new_[28237]_ ;
  assign \new_[26817]_  = ~\new_[30411]_  | ~\new_[29560]_ ;
  assign \new_[26818]_  = (~\new_[29807]_  | ~\s14_data_i[31] ) & (~\new_[30626]_  | ~\s12_data_i[31] );
  assign \new_[26819]_  = ~\new_[28158]_ ;
  assign \new_[26820]_  = (~\new_[30113]_  | ~\s2_data_i[1] ) & (~\new_[30124]_  | ~\s1_data_i[1] );
  assign \new_[26821]_  = ~\new_[30062]_ ;
  assign \new_[26822]_  = ~\new_[29841]_  | ~\new_[29527]_ ;
  assign \new_[26823]_  = ~\new_[28882]_  & ~\new_[5921]_ ;
  assign \new_[26824]_  = \new_[29898]_  & \new_[29268]_ ;
  assign \new_[26825]_  = ~\new_[28196]_ ;
  assign \new_[26826]_  = ~\new_[28497]_ ;
  assign \new_[26827]_  = ~\new_[28673]_ ;
  assign \new_[26828]_  = ~\new_[28092]_ ;
  assign \new_[26829]_  = ~\new_[28086]_ ;
  assign \new_[26830]_  = (~\new_[30088]_  | ~\s2_data_i[26] ) & (~\new_[29779]_  | ~\s1_data_i[26] );
  assign \new_[26831]_  = ~\new_[28220]_ ;
  assign \new_[26832]_  = ~\new_[28708]_ ;
  assign \new_[26833]_  = ~\new_[29119]_  | ~\new_[29357]_ ;
  assign \new_[26834]_  = \new_[29212]_  & \new_[31394]_ ;
  assign \new_[26835]_  = ~\new_[30599]_  | ~\new_[30235]_ ;
  assign \new_[26836]_  = (~\new_[29876]_  | ~\s11_data_i[25] ) & (~\new_[30341]_  | ~\s8_data_i[25] );
  assign \new_[26837]_  = ~\new_[30670]_  | ~\new_[29077]_ ;
  assign \new_[26838]_  = ~\new_[28985]_  | ~\new_[5993]_ ;
  assign \new_[26839]_  = \new_[28992]_  | \new_[30030]_ ;
  assign \new_[26840]_  = \new_[29357]_  & \new_[6202]_ ;
  assign \new_[26841]_  = ~\new_[28585]_ ;
  assign \new_[26842]_  = ~\new_[29251]_ ;
  assign \new_[26843]_  = \new_[29355]_  & \new_[5920]_ ;
  assign \new_[26844]_  = ~\new_[29971]_  | ~\new_[30542]_ ;
  assign \new_[26845]_  = ~\new_[29765]_ ;
  assign \new_[26846]_  = ~\new_[28909]_  & ~\new_[29233]_ ;
  assign \new_[26847]_  = ~\new_[28864]_  | ~\new_[30062]_ ;
  assign \new_[26848]_  = (~\new_[30088]_  | ~\s2_data_i[8] ) & (~\new_[29779]_  | ~\s1_data_i[8] );
  assign \new_[26849]_  = \new_[29463]_  & \new_[29296]_ ;
  assign \new_[26850]_  = ~\new_[28967]_  | ~\new_[6064]_ ;
  assign \new_[26851]_  = ~\new_[29043]_ ;
  assign \new_[26852]_  = ~\new_[29606]_  & ~\new_[30277]_ ;
  assign \new_[26853]_  = ~\new_[29551]_  & ~\new_[30063]_ ;
  assign \new_[26854]_  = (~\new_[30189]_  | ~\s2_data_i[16] ) & (~\new_[30195]_  | ~\s1_data_i[16] );
  assign \new_[26855]_  = ~\new_[28934]_  & ~\new_[29501]_ ;
  assign \new_[26856]_  = \new_[29674]_  & \new_[30577]_ ;
  assign \new_[26857]_  = \new_[28899]_  & \new_[28883]_ ;
  assign \new_[26858]_  = ~\new_[28367]_ ;
  assign \new_[26859]_  = ~\new_[28230]_ ;
  assign \new_[26860]_  = ~\new_[30151]_  & ~\new_[30556]_ ;
  assign \new_[26861]_  = ~\new_[29383]_  & ~\new_[31683]_ ;
  assign \new_[26862]_  = ~\new_[29827]_  & ~\new_[29168]_ ;
  assign \new_[26863]_  = ~\new_[28287]_ ;
  assign \new_[26864]_  = ~\new_[29082]_  | ~\new_[5985]_ ;
  assign \new_[26865]_  = ~\new_[28479]_ ;
  assign \new_[26866]_  = ~\new_[28889]_  | ~\new_[29613]_ ;
  assign \new_[26867]_  = ~\new_[29587]_  | ~\new_[29511]_ ;
  assign \new_[26868]_  = \new_[29431]_  & \new_[30152]_ ;
  assign \new_[26869]_  = \new_[29500]_  & \new_[30152]_ ;
  assign \new_[26870]_  = (~\new_[30166]_  | ~\s14_data_i[0] ) & (~\new_[30298]_  | ~\s12_data_i[0] );
  assign \new_[26871]_  = ~\new_[28295]_ ;
  assign \new_[26872]_  = (~\new_[30088]_  | ~\s2_data_i[28] ) & (~\new_[29779]_  | ~\s1_data_i[28] );
  assign \new_[26873]_  = ~\new_[29513]_  | ~\new_[29517]_ ;
  assign \new_[26874]_  = ~\new_[29629]_  | ~\new_[28898]_ ;
  assign \new_[26875]_  = ~\new_[29211]_  | ~\new_[30730]_ ;
  assign \new_[26876]_  = ~\new_[6246]_  | ~\new_[30020]_  | ~\new_[30726]_ ;
  assign \new_[26877]_  = ~\new_[29014]_  | ~\new_[6066]_ ;
  assign \new_[26878]_  = ~\new_[29129]_  | ~\new_[29393]_ ;
  assign \new_[26879]_  = ~\new_[28297]_ ;
  assign \new_[26880]_  = \new_[29479]_  | \new_[30736]_ ;
  assign \new_[26881]_  = \new_[29388]_  & \new_[29473]_ ;
  assign \new_[26882]_  = \new_[29437]_  & \new_[30572]_ ;
  assign \new_[26883]_  = \new_[28871]_  & \new_[29798]_ ;
  assign \new_[26884]_  = ~\new_[29514]_  | ~\new_[28860]_ ;
  assign \new_[26885]_  = ~\new_[30407]_  & ~\new_[29271]_ ;
  assign \new_[26886]_  = (~\new_[30189]_  | ~\s2_data_i[4] ) & (~\new_[30195]_  | ~\s1_data_i[4] );
  assign \new_[26887]_  = ~\new_[29264]_  | ~\new_[29520]_ ;
  assign \new_[26888]_  = \new_[29457]_  & \new_[29798]_ ;
  assign \new_[26889]_  = ~\new_[6176]_  | ~\new_[30135]_  | ~\new_[30232]_ ;
  assign \new_[26890]_  = \new_[29026]_  | \new_[30425]_ ;
  assign \new_[26891]_  = \new_[29502]_  & \new_[30135]_ ;
  assign \new_[26892]_  = ~\new_[28002]_ ;
  assign \new_[26893]_  = \new_[29561]_  & \new_[29975]_ ;
  assign \new_[26894]_  = ~\new_[29521]_  | ~\new_[30256]_ ;
  assign \new_[26895]_  = ~\new_[6204]_  | ~\new_[30665]_  | ~\new_[30750]_ ;
  assign \new_[26896]_  = ~\new_[29490]_  | ~\new_[30750]_ ;
  assign \new_[26897]_  = ~\new_[29515]_  | ~\new_[29177]_ ;
  assign \new_[26898]_  = \new_[29490]_  & \new_[30139]_ ;
  assign \new_[26899]_  = \new_[29525]_  & \new_[29759]_ ;
  assign \new_[26900]_  = ~\new_[29383]_  & ~\new_[29455]_ ;
  assign \new_[26901]_  = ~\new_[29848]_  | ~\new_[29260]_ ;
  assign \new_[26902]_  = \new_[29478]_  | \new_[30253]_ ;
  assign \new_[26903]_  = ~\new_[29346]_  | ~\new_[30507]_ ;
  assign \new_[26904]_  = ~\new_[28777]_ ;
  assign \new_[26905]_  = ~\new_[30015]_  | ~\new_[29880]_ ;
  assign \new_[26906]_  = \new_[29498]_  & \new_[30446]_ ;
  assign \new_[26907]_  = \new_[29430]_  | \new_[30757]_ ;
  assign \new_[26908]_  = ~\new_[28823]_  | ~\new_[29507]_ ;
  assign \new_[26909]_  = \new_[29117]_  | \new_[30757]_ ;
  assign \new_[26910]_  = ~\new_[29530]_  | ~\new_[29426]_ ;
  assign \new_[26911]_  = ~\new_[29338]_  | ~\new_[30538]_ ;
  assign \new_[26912]_  = ~\new_[28402]_  & ~\new_[31870]_ ;
  assign \new_[26913]_  = ~\new_[28302]_ ;
  assign \new_[26914]_  = \new_[29440]_  & \new_[30011]_ ;
  assign \new_[26915]_  = ~\new_[29519]_  | ~\new_[29405]_ ;
  assign \new_[26916]_  = (~\new_[29876]_  | ~\s11_data_i[26] ) & (~\new_[30341]_  | ~\s8_data_i[26] );
  assign \new_[26917]_  = ~\new_[29701]_  | ~\new_[6001]_ ;
  assign \new_[26918]_  = \new_[29385]_  & \new_[30957]_ ;
  assign \new_[26919]_  = ~\new_[29485]_  | ~\new_[30544]_ ;
  assign \new_[26920]_  = ~\new_[29127]_  | ~\new_[29356]_ ;
  assign \new_[26921]_  = \new_[29403]_  & \new_[29529]_ ;
  assign \new_[26922]_  = ~\new_[29120]_  | ~\new_[29224]_ ;
  assign \new_[26923]_  = \new_[29244]_  | \new_[28944]_ ;
  assign \new_[26924]_  = ~\new_[28473]_ ;
  assign \new_[26925]_  = ~\new_[29712]_  | ~\new_[5912]_ ;
  assign \new_[26926]_  = (~\new_[30088]_  | ~\s2_data_i[7] ) & (~\new_[29779]_  | ~\s1_data_i[7] );
  assign \new_[26927]_  = \new_[29346]_  & \new_[30437]_ ;
  assign \new_[26928]_  = \new_[29577]_  & \new_[30444]_ ;
  assign \new_[26929]_  = (~\new_[30189]_  | ~\s2_data_i[0] ) & (~\new_[30195]_  | ~\s1_data_i[0] );
  assign \new_[26930]_  = \new_[28978]_  & \new_[30645]_ ;
  assign \new_[26931]_  = \new_[29512]_  & \new_[29522]_ ;
  assign \new_[26932]_  = \new_[29439]_  & \new_[30697]_ ;
  assign \new_[26933]_  = ~\new_[29783]_  | ~\new_[29347]_ ;
  assign \new_[26934]_  = ~\new_[29289]_  & ~\new_[30225]_ ;
  assign \new_[26935]_  = (~\new_[29807]_  | ~\s14_data_i[10] ) & (~\new_[30626]_  | ~\s12_data_i[10] );
  assign \new_[26936]_  = \new_[29286]_  | \new_[29624]_ ;
  assign \new_[26937]_  = \new_[29286]_  & \new_[30645]_ ;
  assign \new_[26938]_  = (~\new_[30088]_  | ~\s2_data_i[12] ) & (~\new_[29779]_  | ~\s1_data_i[12] );
  assign \new_[26939]_  = (~\new_[30189]_  | ~\s2_data_i[9] ) & (~\new_[30195]_  | ~\s1_data_i[9] );
  assign \new_[26940]_  = ~\new_[29315]_  & ~\new_[29347]_ ;
  assign \new_[26941]_  = ~\new_[29892]_  | ~\new_[29545]_ ;
  assign \new_[26942]_  = ~\new_[6212]_  | ~\new_[30595]_  | ~\new_[30765]_ ;
  assign \new_[26943]_  = ~\new_[29785]_  & ~\new_[28873]_ ;
  assign \new_[26944]_  = (~\new_[30131]_  | ~\s7_data_i[20] ) & (~\new_[29939]_  | ~\s6_data_i[20] );
  assign \new_[26945]_  = \new_[29387]_  & \new_[29785]_ ;
  assign \new_[26946]_  = ~\new_[28430]_ ;
  assign \new_[26947]_  = ~\new_[29438]_  | ~\new_[29509]_ ;
  assign \new_[26948]_  = ~\new_[30845]_  & ~\new_[28069]_ ;
  assign \new_[26949]_  = ~\new_[5991]_  | ~\new_[29912]_  | ~\new_[30784]_ ;
  assign \new_[26950]_  = ~\new_[30578]_  | ~\new_[5925]_ ;
  assign \new_[26951]_  = ~\new_[29952]_  & ~\new_[28050]_ ;
  assign \new_[26952]_  = ~\new_[28644]_ ;
  assign \new_[26953]_  = ~\new_[29669]_  | ~\new_[5902]_ ;
  assign \new_[26954]_  = ~\new_[28387]_ ;
  assign \new_[26955]_  = ~\new_[29481]_  & ~\new_[30185]_ ;
  assign \new_[26956]_  = ~\new_[29214]_  | ~\new_[29329]_ ;
  assign \new_[26957]_  = (~\new_[30088]_  | ~\s2_data_i[14] ) & (~\new_[29779]_  | ~\s1_data_i[14] );
  assign \new_[26958]_  = ~\new_[29182]_  & ~\new_[30228]_ ;
  assign \new_[26959]_  = \new_[29460]_  | \new_[30438]_ ;
  assign \new_[26960]_  = \new_[29468]_  & \new_[30352]_ ;
  assign \new_[26961]_  = ~\new_[28819]_  & ~\new_[30784]_ ;
  assign \new_[26962]_  = \new_[29485]_  & \new_[30727]_ ;
  assign \new_[26963]_  = (~\new_[29961]_  | ~\s4_data_i[3] ) & (~\new_[29819]_  | ~\s0_data_i[3] );
  assign \new_[26964]_  = ~\new_[28890]_  | ~\new_[5917]_ ;
  assign \new_[26965]_  = ~\new_[6064]_  | ~\new_[30636]_  | ~\new_[30574]_ ;
  assign \new_[26966]_  = ~\new_[28279]_ ;
  assign \new_[26967]_  = \new_[29443]_  & \new_[30717]_ ;
  assign \new_[26968]_  = \new_[29600]_  | \new_[30736]_ ;
  assign \new_[26969]_  = ~\new_[29539]_  & ~\new_[30515]_ ;
  assign \new_[26970]_  = ~\new_[28959]_  | ~\new_[30820]_ ;
  assign \new_[26971]_  = \new_[29448]_  | \new_[30736]_ ;
  assign \new_[26972]_  = ~\new_[6007]_  | ~\new_[29118]_  | ~\new_[30820]_ ;
  assign \new_[26973]_  = ~\new_[30138]_  | ~\new_[28891]_ ;
  assign \new_[26974]_  = ~\new_[30731]_  | ~\new_[6050]_ ;
  assign \new_[26975]_  = \new_[29176]_  & \new_[30786]_ ;
  assign \new_[26976]_  = ~\new_[29098]_  & ~\new_[30309]_ ;
  assign \new_[26977]_  = \new_[29741]_  & \new_[31421]_ ;
  assign \new_[26978]_  = ~\new_[29470]_  | ~\new_[29210]_ ;
  assign \new_[26979]_  = ~\new_[28370]_ ;
  assign \new_[26980]_  = ~\new_[30344]_  | ~\new_[29256]_ ;
  assign \new_[26981]_  = ~\new_[6269]_  | ~\new_[29210]_  | ~\new_[30789]_ ;
  assign \new_[26982]_  = ~\new_[29581]_  & ~\new_[29964]_ ;
  assign \new_[26983]_  = ~\new_[29402]_  | ~\new_[29242]_ ;
  assign \new_[26984]_  = ~\new_[5991]_  | ~\new_[29785]_  | ~\new_[29912]_ ;
  assign \new_[26985]_  = ~\new_[29208]_  | ~\new_[29516]_ ;
  assign \new_[26986]_  = ~\new_[29372]_  | ~\new_[30820]_ ;
  assign \new_[26987]_  = ~\new_[29173]_  | ~\new_[29523]_ ;
  assign \new_[26988]_  = (~\new_[30085]_  | ~\s2_data_i[1] ) & (~\new_[30108]_  | ~\s1_data_i[1] );
  assign \new_[26989]_  = ~\new_[6202]_  | ~\new_[29495]_  | ~\new_[29861]_ ;
  assign \new_[26990]_  = ~\new_[28330]_ ;
  assign \new_[26991]_  = ~\new_[30519]_  | ~\new_[6057]_ ;
  assign \new_[26992]_  = ~\new_[32338]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[26993]_  = (~\new_[29846]_  | ~\s2_data_i[0] ) & (~\new_[30001]_  | ~\s1_data_i[0] );
  assign \new_[26994]_  = ~\new_[29051]_  & (~\new_[29808]_  | ~\new_[6183]_ );
  assign \new_[26995]_  = ~\new_[28840]_  | ~\new_[29919]_ ;
  assign \new_[26996]_  = ~\new_[5933]_  | ~\new_[28964]_  | ~\new_[30009]_ ;
  assign \new_[26997]_  = (~\new_[29948]_  | ~\s5_data_i[2] ) & (~\new_[29947]_  | ~\s3_data_i[2] );
  assign \new_[26998]_  = \new_[29632]_  & \new_[29813]_ ;
  assign \new_[26999]_  = ~\new_[28944]_  & ~\new_[30555]_ ;
  assign \new_[27000]_  = ~\new_[29718]_  & ~\new_[5932]_ ;
  assign \new_[27001]_  = ~\new_[29450]_  & (~\new_[30229]_  | ~\new_[6041]_ );
  assign \new_[27002]_  = ~\new_[29537]_  | ~\new_[6085]_ ;
  assign \new_[27003]_  = ~\new_[29123]_  & (~\new_[30222]_  | ~\new_[6205]_ );
  assign \new_[27004]_  = ~\new_[29397]_  | ~\new_[5972]_ ;
  assign \new_[27005]_  = ~\new_[29905]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[27006]_  = ~\new_[29948]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27007]_  = ~\new_[30335]_  | ~\new_[31160]_  | ~m0_cyc_i;
  assign \new_[27008]_  = ~\new_[30260]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[27009]_  = ~\new_[32327]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[27010]_  = ~\new_[30189]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[27011]_  = ~\new_[30354]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[27012]_  = ~\new_[29963]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[27013]_  = ~\new_[30341]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[27014]_  = ~\new_[30200]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27015]_  = ~\new_[28502]_ ;
  assign \new_[27016]_  = ~\new_[30298]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27017]_  = ~\new_[32168]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27018]_  = ~\new_[30166]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27019]_  = ~\new_[29846]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27020]_  = ~\new_[29947]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27021]_  = ~\new_[29939]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27022]_  = ~\new_[30131]_  | ~\new_[31053]_  | ~m3_cyc_i;
  assign \new_[27023]_  = ~\new_[29953]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[27024]_  = ~\new_[30311]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27025]_  = ~\new_[30181]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27026]_  = ~\new_[30013]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27027]_  = ~\new_[29928]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27028]_  = ~\new_[29441]_  | ~\new_[6056]_ ;
  assign \new_[27029]_  = ~\new_[30060]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27030]_  = ~\new_[29951]_  | ~\new_[30918]_  | ~m5_cyc_i;
  assign \new_[27031]_  = ~\new_[30227]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[27032]_  = ~\new_[30085]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[27033]_  = ~\new_[29130]_  & ~\new_[29789]_ ;
  assign \new_[27034]_  = ~\new_[29954]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[27035]_  = ~\new_[29823]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[27036]_  = ~\new_[29949]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[27037]_  = ~\new_[30106]_  | ~\new_[31185]_  | ~m7_cyc_i;
  assign \new_[27038]_  = ~\new_[32056]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[27039]_  = ~\new_[29876]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[27040]_  = ~\new_[29976]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[27041]_  = ~\new_[6094]_  | ~\new_[29495]_  | ~\new_[29861]_ ;
  assign \new_[27042]_  = ~\new_[28058]_ ;
  assign \new_[27043]_  = (~\new_[29961]_  | ~\s4_data_i[12] ) & (~\new_[29819]_  | ~\s0_data_i[12] );
  assign \new_[27044]_  = (~\new_[29948]_  | ~\s5_data_i[11] ) & (~\new_[29947]_  | ~\s3_data_i[11] );
  assign \new_[27045]_  = (~\new_[29949]_  | ~\s10_data_i[0] ) & (~\new_[29905]_  | ~\s9_data_i[0] );
  assign \new_[27046]_  = (~\new_[29876]_  | ~\s11_data_i[24] ) & (~\new_[30341]_  | ~\s8_data_i[24] );
  assign \new_[27047]_  = (~\new_[29948]_  | ~\s5_data_i[8] ) & (~\new_[29947]_  | ~\s3_data_i[8] );
  assign \new_[27048]_  = (~\new_[30013]_  | ~\s2_data_i[5] ) & (~\new_[29769]_  | ~\s1_data_i[5] );
  assign \new_[27049]_  = (~\new_[30189]_  | ~\s2_data_i[26] ) & (~\new_[30195]_  | ~\s1_data_i[26] );
  assign \new_[27050]_  = (~\new_[29961]_  | ~\s4_data_i[16] ) & (~\new_[29819]_  | ~\s0_data_i[16] );
  assign \new_[27051]_  = (~\new_[29807]_  | ~\s14_data_i[23] ) & (~\new_[30626]_  | ~\s12_data_i[23] );
  assign \new_[27052]_  = (~\new_[29788]_  | ~\s2_data_i[22] ) & (~\new_[30357]_  | ~\s1_data_i[22] );
  assign \new_[27053]_  = (~\new_[30113]_  | ~\s2_data_i[24] ) & (~\new_[30124]_  | ~\s1_data_i[24] );
  assign \new_[27054]_  = (~\new_[29876]_  | ~\s11_data_i[22] ) & (~\new_[30341]_  | ~\s8_data_i[22] );
  assign \new_[27055]_  = \new_[29004]_  & \new_[31547]_ ;
  assign \new_[27056]_  = (~\new_[30113]_  | ~\s2_data_i[14] ) & (~\new_[30124]_  | ~\s1_data_i[14] );
  assign \new_[27057]_  = (~\new_[29961]_  | ~\s4_data_i[7] ) & (~\new_[29819]_  | ~\s0_data_i[7] );
  assign \new_[27058]_  = (~\new_[30013]_  | ~\s2_data_i[0] ) & (~\new_[29769]_  | ~\s1_data_i[0] );
  assign \new_[27059]_  = (~\new_[29948]_  | ~\s5_data_i[15] ) & (~\new_[29947]_  | ~\s3_data_i[15] );
  assign \new_[27060]_  = ~\new_[30336]_  & ~\new_[30623]_ ;
  assign \new_[27061]_  = (~\new_[29949]_  | ~\s10_data_i[29] ) & (~\new_[29905]_  | ~\s9_data_i[29] );
  assign \new_[27062]_  = (~\new_[30085]_  | ~\s2_data_i[6] ) & (~\new_[30108]_  | ~\s1_data_i[6] );
  assign \new_[27063]_  = (~\new_[29963]_  | ~\s4_data_i[20] ) & (~\new_[30481]_  | ~\s0_data_i[20] );
  assign \new_[27064]_  = (~\new_[29948]_  | ~\s5_data_i[17] ) & (~\new_[29947]_  | ~\s3_data_i[17] );
  assign \new_[27065]_  = (~\new_[30189]_  | ~\s2_data_i[24] ) & (~\new_[30195]_  | ~\s1_data_i[24] );
  assign \new_[27066]_  = (~\new_[30166]_  | ~\s14_data_i[13] ) & (~\new_[30298]_  | ~\s12_data_i[13] );
  assign \new_[27067]_  = (~\new_[30113]_  | ~\s2_data_i[23] ) & (~\new_[30124]_  | ~\s1_data_i[23] );
  assign \new_[27068]_  = (~\new_[29949]_  | ~\s10_data_i[7] ) & (~\new_[29905]_  | ~\s9_data_i[7] );
  assign \new_[27069]_  = (~\new_[29788]_  | ~\s2_data_i[18] ) & (~\new_[30357]_  | ~\s1_data_i[18] );
  assign \new_[27070]_  = (~\new_[30085]_  | ~\s2_data_i[31] ) & (~\new_[30108]_  | ~\s1_data_i[31] );
  assign \new_[27071]_  = (~\new_[30166]_  | ~\s14_data_i[16] ) & (~\new_[30298]_  | ~\s12_data_i[16] );
  assign \new_[27072]_  = ~\new_[29475]_  & ~\new_[29650]_ ;
  assign \new_[27073]_  = (~\new_[30166]_  | ~\s14_data_i[23] ) & (~\new_[30298]_  | ~\s12_data_i[23] );
  assign \new_[27074]_  = (~\new_[30085]_  | ~\s2_data_i[30] ) & (~\new_[30108]_  | ~\s1_data_i[30] );
  assign \new_[27075]_  = (~\new_[29788]_  | ~\s2_data_i[17] ) & (~\new_[30357]_  | ~\s1_data_i[17] );
  assign \new_[27076]_  = (~\new_[30131]_  | ~\s7_data_i[2] ) & (~\new_[29939]_  | ~\s6_data_i[2] );
  assign \new_[27077]_  = (~\new_[30088]_  | ~\s2_data_i[29] ) & (~\new_[29779]_  | ~\s1_data_i[29] );
  assign \new_[27078]_  = (~\new_[29961]_  | ~\s4_data_i[27] ) & (~\new_[29819]_  | ~\s0_data_i[27] );
  assign \new_[27079]_  = (~\new_[30085]_  | ~\s2_data_i[29] ) & (~\new_[30108]_  | ~\s1_data_i[29] );
  assign \new_[27080]_  = \new_[28850]_  & \new_[6005]_ ;
  assign \new_[27081]_  = (~\new_[29846]_  | ~\s2_data_i[8] ) & (~\new_[30001]_  | ~\s1_data_i[8] );
  assign \new_[27082]_  = (~\new_[30166]_  | ~\s14_data_i[17] ) & (~\new_[30298]_  | ~\s12_data_i[17] );
  assign \new_[27083]_  = ~\new_[28724]_  | ~\new_[5906]_ ;
  assign \new_[27084]_  = (~\new_[30013]_  | ~\s2_data_i[14] ) & (~\new_[29769]_  | ~\s1_data_i[14] );
  assign \new_[27085]_  = ~\new_[29735]_  & ~\new_[31148]_ ;
  assign \new_[27086]_  = (~\new_[29807]_  | ~\s14_data_i[18] ) & (~\new_[30626]_  | ~\s12_data_i[18] );
  assign \new_[27087]_  = (~\new_[30085]_  | ~\s2_data_i[27] ) & (~\new_[30108]_  | ~\s1_data_i[27] );
  assign \new_[27088]_  = ~\new_[29291]_  & ~\new_[29597]_ ;
  assign \new_[27089]_  = (~\new_[29788]_  | ~\s2_data_i[16] ) & (~\new_[30357]_  | ~\s1_data_i[16] );
  assign \new_[27090]_  = (~\new_[29823]_  | ~\s7_data_i[26] ) & (~\new_[29954]_  | ~\s6_data_i[26] );
  assign \new_[27091]_  = (~\new_[29963]_  | ~\s4_data_i[15] ) & (~\new_[30481]_  | ~\s0_data_i[15] );
  assign \new_[27092]_  = (~\new_[29823]_  | ~\s7_data_i[25] ) & (~\new_[29954]_  | ~\s6_data_i[25] );
  assign \new_[27093]_  = ~\new_[29112]_  | ~\new_[29908]_ ;
  assign \new_[27094]_  = (~\new_[29807]_  | ~\s14_data_i[15] ) & (~\new_[30626]_  | ~\s12_data_i[15] );
  assign \new_[27095]_  = (~\new_[29788]_  | ~\s2_data_i[10] ) & (~\new_[30357]_  | ~\s1_data_i[10] );
  assign \new_[27096]_  = (~\new_[30085]_  | ~\s2_data_i[25] ) & (~\new_[30108]_  | ~\s1_data_i[25] );
  assign \new_[27097]_  = (~\new_[30131]_  | ~\s7_data_i[23] ) & (~\new_[29939]_  | ~\s6_data_i[23] );
  assign \new_[27098]_  = ~\new_[30083]_  | ~\new_[29071]_ ;
  assign \new_[27099]_  = (~\new_[29807]_  | ~\s14_data_i[14] ) & (~\new_[30626]_  | ~\s12_data_i[14] );
  assign \new_[27100]_  = (~\new_[30088]_  | ~\s2_data_i[13] ) & (~\new_[29779]_  | ~\s1_data_i[13] );
  assign \new_[27101]_  = (~\new_[29823]_  | ~\s7_data_i[22] ) & (~\new_[29954]_  | ~\s6_data_i[22] );
  assign \new_[27102]_  = (~\new_[29963]_  | ~\s4_data_i[24] ) & (~\new_[30481]_  | ~\s0_data_i[24] );
  assign \new_[27103]_  = \new_[29741]_  & \new_[5997]_ ;
  assign \new_[27104]_  = (~\new_[29807]_  | ~\s14_data_i[13] ) & (~\new_[30626]_  | ~\s12_data_i[13] );
  assign \new_[27105]_  = (~\new_[29846]_  | ~\s2_data_i[10] ) & (~\new_[30001]_  | ~\s1_data_i[10] );
  assign \new_[27106]_  = (~\new_[30085]_  | ~\s2_data_i[21] ) & (~\new_[30108]_  | ~\s1_data_i[21] );
  assign \new_[27107]_  = (~\new_[29876]_  | ~\s11_data_i[12] ) & (~\new_[30341]_  | ~\s8_data_i[12] );
  assign \new_[27108]_  = (~\new_[29823]_  | ~\s7_data_i[19] ) & (~\new_[29954]_  | ~\s6_data_i[19] );
  assign \new_[27109]_  = (~\new_[29807]_  | ~\s14_data_i[12] ) & (~\new_[30626]_  | ~\s12_data_i[12] );
  assign \new_[27110]_  = (~\new_[30085]_  | ~\s2_data_i[19] ) & (~\new_[30108]_  | ~\s1_data_i[19] );
  assign \new_[27111]_  = (~\new_[29949]_  | ~\s10_data_i[4] ) & (~\new_[29905]_  | ~\s9_data_i[4] );
  assign \new_[27112]_  = (~\new_[29963]_  | ~\s4_data_i[11] ) & (~\new_[30481]_  | ~\s0_data_i[11] );
  assign \new_[27113]_  = (~\new_[29961]_  | ~\s4_data_i[24] ) & (~\new_[29819]_  | ~\s0_data_i[24] );
  assign \new_[27114]_  = (~\new_[29788]_  | ~\s2_data_i[11] ) & (~\new_[30357]_  | ~\s1_data_i[11] );
  assign \new_[27115]_  = (~\new_[30013]_  | ~\s2_data_i[15] ) & (~\new_[29769]_  | ~\s1_data_i[15] );
  assign \new_[27116]_  = (~\new_[29876]_  | ~\s11_data_i[11] ) & (~\new_[30341]_  | ~\s8_data_i[11] );
  assign \new_[27117]_  = (~\new_[29823]_  | ~\s7_data_i[17] ) & (~\new_[29954]_  | ~\s6_data_i[17] );
  assign \new_[27118]_  = (~\new_[29846]_  | ~\s2_data_i[17] ) & (~\new_[30001]_  | ~\s1_data_i[17] );
  assign \new_[27119]_  = (~\new_[29963]_  | ~\s4_data_i[10] ) & (~\new_[30481]_  | ~\s0_data_i[10] );
  assign \new_[27120]_  = (~\new_[30113]_  | ~\s2_data_i[0] ) & (~\new_[30124]_  | ~\s1_data_i[0] );
  assign \new_[27121]_  = (~\new_[29948]_  | ~\s5_data_i[6] ) & (~\new_[29947]_  | ~\s3_data_i[6] );
  assign \new_[27122]_  = (~\new_[29823]_  | ~\s7_data_i[15] ) & (~\new_[29954]_  | ~\s6_data_i[15] );
  assign \new_[27123]_  = (~\new_[29807]_  | ~\s14_data_i[29] ) & (~\new_[30626]_  | ~\s12_data_i[29] );
  assign \new_[27124]_  = (~\new_[30131]_  | ~\s7_data_i[11] ) & (~\new_[29939]_  | ~\s6_data_i[11] );
  assign \new_[27125]_  = (~\new_[29823]_  | ~\s7_data_i[14] ) & (~\new_[29954]_  | ~\s6_data_i[14] );
  assign \new_[27126]_  = (~\new_[30085]_  | ~\s2_data_i[14] ) & (~\new_[30108]_  | ~\s1_data_i[14] );
  assign \new_[27127]_  = (~\new_[29876]_  | ~\s11_data_i[29] ) & (~\new_[30341]_  | ~\s8_data_i[29] );
  assign \new_[27128]_  = (~\new_[29807]_  | ~\s14_data_i[6] ) & (~\new_[30626]_  | ~\s12_data_i[6] );
  assign \new_[27129]_  = (~\new_[30113]_  | ~\s2_data_i[29] ) & (~\new_[30124]_  | ~\s1_data_i[29] );
  assign \new_[27130]_  = \new_[29671]_  | \new_[30363]_ ;
  assign \new_[27131]_  = (~\new_[29963]_  | ~\s4_data_i[8] ) & (~\new_[30481]_  | ~\s0_data_i[8] );
  assign \new_[27132]_  = ~\new_[30579]_  & ~\new_[30732]_ ;
  assign \new_[27133]_  = (~\new_[30085]_  | ~\s2_data_i[12] ) & (~\new_[30108]_  | ~\s1_data_i[12] );
  assign \new_[27134]_  = (~\new_[29949]_  | ~\s10_data_i[18] ) & (~\new_[29905]_  | ~\s9_data_i[18] );
  assign \new_[27135]_  = (~\new_[29846]_  | ~\s2_data_i[13] ) & (~\new_[30001]_  | ~\s1_data_i[13] );
  assign \new_[27136]_  = ~\new_[30556]_  | ~\new_[6078]_ ;
  assign \new_[27137]_  = (~\new_[30085]_  | ~\s2_data_i[13] ) & (~\new_[30108]_  | ~\s1_data_i[13] );
  assign \new_[27138]_  = (~\new_[30013]_  | ~\s2_data_i[16] ) & (~\new_[29769]_  | ~\s1_data_i[16] );
  assign \new_[27139]_  = (~\new_[30166]_  | ~\s14_data_i[28] ) & (~\new_[30298]_  | ~\s12_data_i[28] );
  assign \new_[27140]_  = (~\new_[29963]_  | ~\s4_data_i[6] ) & (~\new_[30481]_  | ~\s0_data_i[6] );
  assign \new_[27141]_  = (~\new_[30131]_  | ~\s7_data_i[7] ) & (~\new_[29939]_  | ~\s6_data_i[7] );
  assign \new_[27142]_  = (~\new_[30088]_  | ~\s2_data_i[10] ) & (~\new_[29779]_  | ~\s1_data_i[10] );
  assign \new_[27143]_  = (~\new_[29963]_  | ~\s4_data_i[16] ) & (~\new_[30481]_  | ~\s0_data_i[16] );
  assign \new_[27144]_  = (~\new_[29876]_  | ~\s11_data_i[6] ) & (~\new_[30341]_  | ~\s8_data_i[6] );
  assign \new_[27145]_  = (~\new_[29823]_  | ~\s7_data_i[7] ) & (~\new_[29954]_  | ~\s6_data_i[7] );
  assign \new_[27146]_  = (~\new_[29961]_  | ~\s4_data_i[25] ) & (~\new_[29819]_  | ~\s0_data_i[25] );
  assign \new_[27147]_  = (~\new_[30131]_  | ~\s7_data_i[6] ) & (~\new_[29939]_  | ~\s6_data_i[6] );
  assign \new_[27148]_  = (~\new_[30113]_  | ~\s2_data_i[16] ) & (~\new_[30124]_  | ~\s1_data_i[16] );
  assign \new_[27149]_  = (~\new_[30088]_  | ~\s2_data_i[25] ) & (~\new_[29779]_  | ~\s1_data_i[25] );
  assign \new_[27150]_  = (~\new_[29823]_  | ~\s7_data_i[6] ) & (~\new_[29954]_  | ~\s6_data_i[6] );
  assign \new_[27151]_  = (~\new_[30166]_  | ~\s14_data_i[20] ) & (~\new_[30298]_  | ~\s12_data_i[20] );
  assign \new_[27152]_  = (~\new_[29788]_  | ~\s2_data_i[5] ) & (~\new_[30357]_  | ~\s1_data_i[5] );
  assign \new_[27153]_  = (~\new_[30131]_  | ~\s7_data_i[18] ) & (~\new_[29939]_  | ~\s6_data_i[18] );
  assign \new_[27154]_  = (~\new_[29823]_  | ~\s7_data_i[5] ) & (~\new_[29954]_  | ~\s6_data_i[5] );
  assign \new_[27155]_  = (~\new_[30085]_  | ~\s2_data_i[5] ) & (~\new_[30108]_  | ~\s1_data_i[5] );
  assign \new_[27156]_  = (~\new_[30166]_  | ~\s14_data_i[24] ) & (~\new_[30298]_  | ~\s12_data_i[24] );
  assign \new_[27157]_  = (~\new_[30166]_  | ~\s14_data_i[6] ) & (~\new_[30298]_  | ~\s12_data_i[6] );
  assign \new_[27158]_  = ~\new_[29602]_  | ~\new_[31429]_ ;
  assign \new_[27159]_  = (~\new_[29876]_  | ~\s11_data_i[1] ) & (~\new_[30341]_  | ~\s8_data_i[1] );
  assign \new_[27160]_  = (~\new_[29963]_  | ~\s4_data_i[4] ) & (~\new_[30481]_  | ~\s0_data_i[4] );
  assign \new_[27161]_  = (~\new_[29823]_  | ~\s7_data_i[4] ) & (~\new_[29954]_  | ~\s6_data_i[4] );
  assign \new_[27162]_  = (~\new_[30088]_  | ~\s2_data_i[11] ) & (~\new_[29779]_  | ~\s1_data_i[11] );
  assign \new_[27163]_  = (~\new_[29823]_  | ~\s7_data_i[2] ) & (~\new_[29954]_  | ~\s6_data_i[2] );
  assign \new_[27164]_  = (~\new_[29807]_  | ~\s14_data_i[8] ) & (~\new_[30626]_  | ~\s12_data_i[8] );
  assign \new_[27165]_  = (~\new_[29846]_  | ~\s2_data_i[4] ) & (~\new_[30001]_  | ~\s1_data_i[4] );
  assign \new_[27166]_  = (~\new_[30013]_  | ~\s2_data_i[17] ) & (~\new_[29769]_  | ~\s1_data_i[17] );
  assign \new_[27167]_  = (~\new_[29788]_  | ~\s2_data_i[3] ) & (~\new_[30357]_  | ~\s1_data_i[3] );
  assign \new_[27168]_  = (~\new_[29846]_  | ~\s2_data_i[24] ) & (~\new_[30001]_  | ~\s1_data_i[24] );
  assign \new_[27169]_  = (~\new_[29807]_  | ~\s14_data_i[3] ) & (~\new_[30626]_  | ~\s12_data_i[3] );
  assign \new_[27170]_  = ~\new_[6176]_  | ~\new_[30232]_  | ~\new_[30508]_ ;
  assign \new_[27171]_  = (~\new_[30088]_  | ~\s2_data_i[20] ) & (~\new_[29779]_  | ~\s1_data_i[20] );
  assign \new_[27172]_  = (~\new_[29788]_  | ~\s2_data_i[2] ) & (~\new_[30357]_  | ~\s1_data_i[2] );
  assign \new_[27173]_  = (~\new_[29949]_  | ~\s10_data_i[1] ) & (~\new_[29905]_  | ~\s9_data_i[1] );
  assign \new_[27174]_  = (~\new_[29949]_  | ~\s10_data_i[31] ) & (~\new_[29905]_  | ~\s9_data_i[31] );
  assign \new_[27175]_  = (~\new_[29876]_  | ~\s11_data_i[10] ) & (~\new_[30341]_  | ~\s8_data_i[10] );
  assign \new_[27176]_  = (~\new_[30113]_  | ~\s2_data_i[30] ) & (~\new_[30124]_  | ~\s1_data_i[30] );
  assign \new_[27177]_  = \new_[29219]_  & \new_[5965]_ ;
  assign \new_[27178]_  = (~\new_[30131]_  | ~\s7_data_i[13] ) & (~\new_[29939]_  | ~\s6_data_i[13] );
  assign \new_[27179]_  = (~\new_[29876]_  | ~\s11_data_i[5] ) & (~\new_[30341]_  | ~\s8_data_i[5] );
  assign \new_[27180]_  = (~\new_[29876]_  | ~\s11_data_i[31] ) & (~\new_[30341]_  | ~\s8_data_i[31] );
  assign \new_[27181]_  = (~\new_[30113]_  | ~\s2_data_i[6] ) & (~\new_[30124]_  | ~\s1_data_i[6] );
  assign \new_[27182]_  = (~\new_[30085]_  | ~\s2_data_i[16] ) & (~\new_[30108]_  | ~\s1_data_i[16] );
  assign \new_[27183]_  = (~\new_[30113]_  | ~\s2_data_i[28] ) & (~\new_[30124]_  | ~\s1_data_i[28] );
  assign \new_[27184]_  = (~\new_[29823]_  | ~\s7_data_i[12] ) & (~\new_[29954]_  | ~\s6_data_i[12] );
  assign \new_[27185]_  = (~\new_[30113]_  | ~\s2_data_i[17] ) & (~\new_[30124]_  | ~\s1_data_i[17] );
  assign \new_[27186]_  = (~\new_[29788]_  | ~\s2_data_i[19] ) & (~\new_[30357]_  | ~\s1_data_i[19] );
  assign \new_[27187]_  = (~\new_[29949]_  | ~\s10_data_i[26] ) & (~\new_[29905]_  | ~\s9_data_i[26] );
  assign \new_[27188]_  = (~\new_[29846]_  | ~\s2_data_i[6] ) & (~\new_[30001]_  | ~\s1_data_i[6] );
  assign \new_[27189]_  = (~\new_[29949]_  | ~\s10_data_i[5] ) & (~\new_[29905]_  | ~\s9_data_i[5] );
  assign \new_[27190]_  = (~\new_[29823]_  | ~\s7_data_i[16] ) & (~\new_[29954]_  | ~\s6_data_i[16] );
  assign \new_[27191]_  = ~\new_[30304]_ ;
  assign \new_[27192]_  = (~\new_[30088]_  | ~\s2_data_i[16] ) & (~\new_[29779]_  | ~\s1_data_i[16] );
  assign \new_[27193]_  = (~\new_[29961]_  | ~\s4_data_i[23] ) & (~\new_[29819]_  | ~\s0_data_i[23] );
  assign \new_[27194]_  = (~\new_[29823]_  | ~\s7_data_i[9] ) & (~\new_[29954]_  | ~\s6_data_i[9] );
  assign \new_[27195]_  = (~\new_[29949]_  | ~\s10_data_i[21] ) & (~\new_[29905]_  | ~\s9_data_i[21] );
  assign \new_[27196]_  = ~\new_[30607]_  & ~\new_[30586]_ ;
  assign \new_[27197]_  = (~\new_[30131]_  | ~\s7_data_i[31] ) & (~\new_[29939]_  | ~\s6_data_i[31] );
  assign \new_[27198]_  = ~\new_[30271]_  | ~\new_[30442]_ ;
  assign \new_[27199]_  = (~\new_[30166]_  | ~\s14_data_i[31] ) & (~\new_[30298]_  | ~\s12_data_i[31] );
  assign \new_[27200]_  = (~\new_[30113]_  | ~\s2_data_i[19] ) & (~\new_[30124]_  | ~\s1_data_i[19] );
  assign \new_[27201]_  = (~\new_[29949]_  | ~\s10_data_i[16] ) & (~\new_[29905]_  | ~\s9_data_i[16] );
  assign \new_[27202]_  = (~\new_[29948]_  | ~\s5_data_i[31] ) & (~\new_[29947]_  | ~\s3_data_i[31] );
  assign \new_[27203]_  = (~\new_[30113]_  | ~\s2_data_i[18] ) & (~\new_[30124]_  | ~\s1_data_i[18] );
  assign \new_[27204]_  = (~\new_[30085]_  | ~\s2_data_i[17] ) & (~\new_[30108]_  | ~\s1_data_i[17] );
  assign \new_[27205]_  = (~\new_[30131]_  | ~\s7_data_i[30] ) & (~\new_[29939]_  | ~\s6_data_i[30] );
  assign \new_[27206]_  = (~\new_[29788]_  | ~\s2_data_i[1] ) & (~\new_[30357]_  | ~\s1_data_i[1] );
  assign \new_[27207]_  = (~\new_[29846]_  | ~\s2_data_i[30] ) & (~\new_[30001]_  | ~\s1_data_i[30] );
  assign \new_[27208]_  = (~\new_[29949]_  | ~\s10_data_i[17] ) & (~\new_[29905]_  | ~\s9_data_i[17] );
  assign \new_[27209]_  = (~\new_[29948]_  | ~\s5_data_i[30] ) & (~\new_[29947]_  | ~\s3_data_i[30] );
  assign \new_[27210]_  = (~\new_[30085]_  | ~\s2_data_i[10] ) & (~\new_[30108]_  | ~\s1_data_i[10] );
  assign \new_[27211]_  = (~\new_[29807]_  | ~\s14_data_i[11] ) & (~\new_[30626]_  | ~\s12_data_i[11] );
  assign \new_[27212]_  = (~\new_[29961]_  | ~\s4_data_i[29] ) & (~\new_[29819]_  | ~\s0_data_i[29] );
  assign \new_[27213]_  = ~\new_[32343]_  | ~m7_stb_i;
  assign \new_[27214]_  = (~\new_[30131]_  | ~\s7_data_i[29] ) & (~\new_[29939]_  | ~\s6_data_i[29] );
  assign \new_[27215]_  = (~\new_[29961]_  | ~\s4_data_i[1] ) & (~\new_[29819]_  | ~\s0_data_i[1] );
  assign \new_[27216]_  = (~\new_[30166]_  | ~\s14_data_i[25] ) & (~\new_[30298]_  | ~\s12_data_i[25] );
  assign \new_[27217]_  = (~\new_[29823]_  | ~\s7_data_i[13] ) & (~\new_[29954]_  | ~\s6_data_i[13] );
  assign \new_[27218]_  = (~\new_[29963]_  | ~\s4_data_i[0] ) & (~\new_[30481]_  | ~\s0_data_i[0] );
  assign \new_[27219]_  = (~\new_[30131]_  | ~\s7_data_i[28] ) & (~\new_[29939]_  | ~\s6_data_i[28] );
  assign \new_[27220]_  = (~\new_[29949]_  | ~\s10_data_i[28] ) & (~\new_[29905]_  | ~\s9_data_i[28] );
  assign \new_[27221]_  = (~\new_[29788]_  | ~\s2_data_i[29] ) & (~\new_[30357]_  | ~\s1_data_i[29] );
  assign \new_[27222]_  = (~\new_[29823]_  | ~\s7_data_i[3] ) & (~\new_[29954]_  | ~\s6_data_i[3] );
  assign \new_[27223]_  = (~\new_[30131]_  | ~\s7_data_i[1] ) & (~\new_[29939]_  | ~\s6_data_i[1] );
  assign \new_[27224]_  = (~\new_[30113]_  | ~\s2_data_i[12] ) & (~\new_[30124]_  | ~\s1_data_i[12] );
  assign \new_[27225]_  = (~\new_[29961]_  | ~\s4_data_i[30] ) & (~\new_[29819]_  | ~\s0_data_i[30] );
  assign \new_[27226]_  = (~\new_[29788]_  | ~\s2_data_i[31] ) & (~\new_[30357]_  | ~\s1_data_i[31] );
  assign \new_[27227]_  = (~\new_[30131]_  | ~\s7_data_i[15] ) & (~\new_[29939]_  | ~\s6_data_i[15] );
  assign \new_[27228]_  = (~\new_[29961]_  | ~\s4_data_i[17] ) & (~\new_[29819]_  | ~\s0_data_i[17] );
  assign \new_[27229]_  = (~\new_[29823]_  | ~\s7_data_i[18] ) & (~\new_[29954]_  | ~\s6_data_i[18] );
  assign \new_[27230]_  = (~\new_[30131]_  | ~\s7_data_i[26] ) & (~\new_[29939]_  | ~\s6_data_i[26] );
  assign \new_[27231]_  = ~\new_[29541]_  & ~\new_[30415]_ ;
  assign \new_[27232]_  = ~\new_[28573]_ ;
  assign \new_[27233]_  = (~\new_[30166]_  | ~\s14_data_i[26] ) & (~\new_[30298]_  | ~\s12_data_i[26] );
  assign \new_[27234]_  = (~\new_[29949]_  | ~\s10_data_i[20] ) & (~\new_[29905]_  | ~\s9_data_i[20] );
  assign \new_[27235]_  = (~\new_[29949]_  | ~\s10_data_i[23] ) & (~\new_[29905]_  | ~\s9_data_i[23] );
  assign \new_[27236]_  = (~\new_[29846]_  | ~\s2_data_i[22] ) & (~\new_[30001]_  | ~\s1_data_i[22] );
  assign \new_[27237]_  = (~\new_[30131]_  | ~\s7_data_i[25] ) & (~\new_[29939]_  | ~\s6_data_i[25] );
  assign \new_[27238]_  = (~\new_[30166]_  | ~\s14_data_i[2] ) & (~\new_[30298]_  | ~\s12_data_i[2] );
  assign \new_[27239]_  = (~\new_[29948]_  | ~\s5_data_i[25] ) & (~\new_[29947]_  | ~\s3_data_i[25] );
  assign \new_[27240]_  = ~\new_[28345]_ ;
  assign \new_[27241]_  = ~\new_[28383]_ ;
  assign \new_[27242]_  = (~\new_[30131]_  | ~\s7_data_i[24] ) & (~\new_[29939]_  | ~\s6_data_i[24] );
  assign \new_[27243]_  = (~\new_[29948]_  | ~\s5_data_i[24] ) & (~\new_[29947]_  | ~\s3_data_i[24] );
  assign \new_[27244]_  = (~\new_[30113]_  | ~\s2_data_i[25] ) & (~\new_[30124]_  | ~\s1_data_i[25] );
  assign \new_[27245]_  = (~\new_[30166]_  | ~\s14_data_i[8] ) & (~\new_[30298]_  | ~\s12_data_i[8] );
  assign \new_[27246]_  = (~\new_[30113]_  | ~\s2_data_i[2] ) & (~\new_[30124]_  | ~\s1_data_i[2] );
  assign \new_[27247]_  = (~\new_[29949]_  | ~\s10_data_i[8] ) & (~\new_[29905]_  | ~\s9_data_i[8] );
  assign \new_[27248]_  = (~\new_[29823]_  | ~\s7_data_i[10] ) & (~\new_[29954]_  | ~\s6_data_i[10] );
  assign \new_[27249]_  = (~\new_[30166]_  | ~\s14_data_i[22] ) & (~\new_[30298]_  | ~\s12_data_i[22] );
  assign \new_[27250]_  = (~\new_[30189]_  | ~\s2_data_i[19] ) & (~\new_[30195]_  | ~\s1_data_i[19] );
  assign \new_[27251]_  = (~\new_[29788]_  | ~\s2_data_i[12] ) & (~\new_[30357]_  | ~\s1_data_i[12] );
  assign \new_[27252]_  = (~\new_[29807]_  | ~\s14_data_i[2] ) & (~\new_[30626]_  | ~\s12_data_i[2] );
  assign \new_[27253]_  = (~\new_[30131]_  | ~\s7_data_i[3] ) & (~\new_[29939]_  | ~\s6_data_i[3] );
  assign \new_[27254]_  = ~\new_[30727]_  | ~\new_[30723]_ ;
  assign \new_[27255]_  = (~\new_[29949]_  | ~\s10_data_i[9] ) & (~\new_[29905]_  | ~\s9_data_i[9] );
  assign \new_[27256]_  = (~\new_[29948]_  | ~\s5_data_i[26] ) & (~\new_[29947]_  | ~\s3_data_i[26] );
  assign \new_[27257]_  = (~\new_[29948]_  | ~\s5_data_i[19] ) & (~\new_[29947]_  | ~\s3_data_i[19] );
  assign \new_[27258]_  = (~\new_[29961]_  | ~\s4_data_i[18] ) & (~\new_[29819]_  | ~\s0_data_i[18] );
  assign \new_[27259]_  = (~\new_[29963]_  | ~\s4_data_i[12] ) & (~\new_[30481]_  | ~\s0_data_i[12] );
  assign \new_[27260]_  = (~\new_[29948]_  | ~\s5_data_i[14] ) & (~\new_[29947]_  | ~\s3_data_i[14] );
  assign \new_[27261]_  = ~\new_[29050]_  | ~\new_[6070]_ ;
  assign \new_[27262]_  = (~\new_[29876]_  | ~\s11_data_i[2] ) & (~\new_[30341]_  | ~\s8_data_i[2] );
  assign \new_[27263]_  = (~\new_[29846]_  | ~\s2_data_i[16] ) & (~\new_[30001]_  | ~\s1_data_i[16] );
  assign \new_[27264]_  = ~\new_[28385]_ ;
  assign \new_[27265]_  = (~\new_[29823]_  | ~\s7_data_i[21] ) & (~\new_[29954]_  | ~\s6_data_i[21] );
  assign \new_[27266]_  = (~\new_[29876]_  | ~\s11_data_i[13] ) & (~\new_[30341]_  | ~\s8_data_i[13] );
  assign \new_[27267]_  = ~\new_[30400]_  & ~\new_[29608]_ ;
  assign \new_[27268]_  = (~\new_[29961]_  | ~\s4_data_i[15] ) & (~\new_[29819]_  | ~\s0_data_i[15] );
  assign \new_[27269]_  = (~\new_[30088]_  | ~\s2_data_i[24] ) & (~\new_[29779]_  | ~\s1_data_i[24] );
  assign \new_[27270]_  = \new_[32127]_  & m6_stb_i;
  assign \new_[27271]_  = (~\new_[30085]_  | ~\s2_data_i[22] ) & (~\new_[30108]_  | ~\s1_data_i[22] );
  assign \new_[27272]_  = ~\new_[30628]_  | ~\new_[6060]_ ;
  assign \new_[27273]_  = (~\new_[29949]_  | ~\s10_data_i[27] ) & (~\new_[29905]_  | ~\s9_data_i[27] );
  assign \new_[27274]_  = (~\new_[30131]_  | ~\s7_data_i[17] ) & (~\new_[29939]_  | ~\s6_data_i[17] );
  assign \new_[27275]_  = (~\new_[30013]_  | ~\s2_data_i[24] ) & (~\new_[29769]_  | ~\s1_data_i[24] );
  assign \new_[27276]_  = (~\new_[29963]_  | ~\s4_data_i[13] ) & (~\new_[30481]_  | ~\s0_data_i[13] );
  assign \new_[27277]_  = (~\new_[29846]_  | ~\s2_data_i[12] ) & (~\new_[30001]_  | ~\s1_data_i[12] );
  assign \new_[27278]_  = (~\new_[29949]_  | ~\s10_data_i[15] ) & (~\new_[29905]_  | ~\s9_data_i[15] );
  assign \new_[27279]_  = (~\new_[30189]_  | ~\s2_data_i[29] ) & (~\new_[30195]_  | ~\s1_data_i[29] );
  assign \new_[27280]_  = (~\new_[30085]_  | ~\s2_data_i[23] ) & (~\new_[30108]_  | ~\s1_data_i[23] );
  assign \new_[27281]_  = \new_[29202]_  & \new_[6062]_ ;
  assign \new_[27282]_  = (~\new_[29949]_  | ~\s10_data_i[10] ) & (~\new_[29905]_  | ~\s9_data_i[10] );
  assign \new_[27283]_  = (~\new_[29846]_  | ~\s2_data_i[26] ) & (~\new_[30001]_  | ~\s1_data_i[26] );
  assign \new_[27284]_  = ~\new_[28399]_ ;
  assign \new_[27285]_  = ~\new_[30267]_ ;
  assign \new_[27286]_  = (~\new_[29823]_  | ~\s7_data_i[23] ) & (~\new_[29954]_  | ~\s6_data_i[23] );
  assign \new_[27287]_  = (~\new_[29948]_  | ~\s5_data_i[27] ) & (~\new_[29947]_  | ~\s3_data_i[27] );
  assign \new_[27288]_  = (~\new_[29876]_  | ~\s11_data_i[14] ) & (~\new_[30341]_  | ~\s8_data_i[14] );
  assign \new_[27289]_  = ~\new_[30055]_  & ~\new_[29571]_ ;
  assign \new_[27290]_  = ~\new_[29145]_  & ~\new_[30413]_ ;
  assign \new_[27291]_  = (~\new_[30085]_  | ~\s2_data_i[0] ) & (~\new_[30108]_  | ~\s1_data_i[0] );
  assign \new_[27292]_  = (~\new_[30013]_  | ~\s2_data_i[25] ) & (~\new_[29769]_  | ~\s1_data_i[25] );
  assign \new_[27293]_  = (~\new_[29788]_  | ~\s2_data_i[14] ) & (~\new_[30357]_  | ~\s1_data_i[14] );
  assign \new_[27294]_  = (~\new_[29963]_  | ~\s4_data_i[2] ) & (~\new_[30481]_  | ~\s0_data_i[2] );
  assign \new_[27295]_  = (~\new_[30166]_  | ~\s14_data_i[1] ) & (~\new_[30298]_  | ~\s12_data_i[1] );
  assign \new_[27296]_  = (~\new_[30166]_  | ~\s14_data_i[12] ) & (~\new_[30298]_  | ~\s12_data_i[12] );
  assign \new_[27297]_  = (~\new_[29963]_  | ~\s4_data_i[14] ) & (~\new_[30481]_  | ~\s0_data_i[14] );
  assign \new_[27298]_  = ~\new_[30650]_  | ~\new_[6032]_ ;
  assign \new_[27299]_  = (~\new_[30085]_  | ~\s2_data_i[24] ) & (~\new_[30108]_  | ~\s1_data_i[24] );
  assign \new_[27300]_  = (~\new_[29846]_  | ~\s2_data_i[23] ) & (~\new_[30001]_  | ~\s1_data_i[23] );
  assign \new_[27301]_  = (~\new_[29948]_  | ~\s5_data_i[10] ) & (~\new_[29947]_  | ~\s3_data_i[10] );
  assign \new_[27302]_  = (~\new_[29846]_  | ~\s2_data_i[14] ) & (~\new_[30001]_  | ~\s1_data_i[14] );
  assign \new_[27303]_  = (~\new_[30166]_  | ~\s14_data_i[5] ) & (~\new_[30298]_  | ~\s12_data_i[5] );
  assign \new_[27304]_  = (~\new_[29823]_  | ~\s7_data_i[29] ) & (~\new_[29954]_  | ~\s6_data_i[29] );
  assign \new_[27305]_  = (~\new_[29823]_  | ~\s7_data_i[11] ) & (~\new_[29954]_  | ~\s6_data_i[11] );
  assign \new_[27306]_  = (~\new_[30131]_  | ~\s7_data_i[16] ) & (~\new_[29939]_  | ~\s6_data_i[16] );
  assign \new_[27307]_  = (~\new_[29961]_  | ~\s4_data_i[19] ) & (~\new_[29819]_  | ~\s0_data_i[19] );
  assign \new_[27308]_  = (~\new_[29948]_  | ~\s5_data_i[4] ) & (~\new_[29947]_  | ~\s3_data_i[4] );
  assign \new_[27309]_  = (~\new_[29876]_  | ~\s11_data_i[15] ) & (~\new_[30341]_  | ~\s8_data_i[15] );
  assign \new_[27310]_  = ~\new_[29040]_  | ~\new_[5931]_ ;
  assign \new_[27311]_  = \new_[29248]_  & \new_[6074]_ ;
  assign \new_[27312]_  = (~\new_[30131]_  | ~\s7_data_i[5] ) & (~\new_[29939]_  | ~\s6_data_i[5] );
  assign \new_[27313]_  = (~\new_[29949]_  | ~\s10_data_i[12] ) & (~\new_[29905]_  | ~\s9_data_i[12] );
  assign \new_[27314]_  = (~\new_[29949]_  | ~\s10_data_i[14] ) & (~\new_[29905]_  | ~\s9_data_i[14] );
  assign \new_[27315]_  = (~\new_[30085]_  | ~\s2_data_i[26] ) & (~\new_[30108]_  | ~\s1_data_i[26] );
  assign \new_[27316]_  = (~\new_[29949]_  | ~\s10_data_i[13] ) & (~\new_[29905]_  | ~\s9_data_i[13] );
  assign \new_[27317]_  = (~\new_[30013]_  | ~\s2_data_i[27] ) & (~\new_[29769]_  | ~\s1_data_i[27] );
  assign \new_[27318]_  = (~\new_[29948]_  | ~\s5_data_i[28] ) & (~\new_[29947]_  | ~\s3_data_i[28] );
  assign \new_[27319]_  = (~\new_[29963]_  | ~\s4_data_i[18] ) & (~\new_[30481]_  | ~\s0_data_i[18] );
  assign \new_[27320]_  = (~\new_[29807]_  | ~\s14_data_i[16] ) & (~\new_[30626]_  | ~\s12_data_i[16] );
  assign \new_[27321]_  = (~\new_[29961]_  | ~\s4_data_i[11] ) & (~\new_[29819]_  | ~\s0_data_i[11] );
  assign \new_[27322]_  = (~\new_[30013]_  | ~\s2_data_i[1] ) & (~\new_[29769]_  | ~\s1_data_i[1] );
  assign \new_[27323]_  = (~\new_[30085]_  | ~\s2_data_i[15] ) & (~\new_[30108]_  | ~\s1_data_i[15] );
  assign \new_[27324]_  = (~\new_[29823]_  | ~\s7_data_i[27] ) & (~\new_[29954]_  | ~\s6_data_i[27] );
  assign \new_[27325]_  = ~\new_[29682]_  & ~\new_[30331]_ ;
  assign \new_[27326]_  = (~\new_[29876]_  | ~\s11_data_i[16] ) & (~\new_[30341]_  | ~\s8_data_i[16] );
  assign \new_[27327]_  = (~\new_[29948]_  | ~\s5_data_i[16] ) & (~\new_[29947]_  | ~\s3_data_i[16] );
  assign \new_[27328]_  = (~\new_[30013]_  | ~\s2_data_i[28] ) & (~\new_[29769]_  | ~\s1_data_i[28] );
  assign \new_[27329]_  = ~\new_[29619]_  | ~\new_[5903]_ ;
  assign \new_[27330]_  = (~\new_[30085]_  | ~\s2_data_i[28] ) & (~\new_[30108]_  | ~\s1_data_i[28] );
  assign \new_[27331]_  = (~\new_[29876]_  | ~\s11_data_i[3] ) & (~\new_[30341]_  | ~\s8_data_i[3] );
  assign \new_[27332]_  = (~\new_[29948]_  | ~\s5_data_i[21] ) & (~\new_[29947]_  | ~\s3_data_i[21] );
  assign \new_[27333]_  = (~\new_[29961]_  | ~\s4_data_i[6] ) & (~\new_[29819]_  | ~\s0_data_i[6] );
  assign \new_[27334]_  = ~\new_[29331]_  | ~\new_[29202]_ ;
  assign \new_[27335]_  = (~\new_[29823]_  | ~\s7_data_i[20] ) & (~\new_[29954]_  | ~\s6_data_i[20] );
  assign \new_[27336]_  = (~\new_[29823]_  | ~\s7_data_i[28] ) & (~\new_[29954]_  | ~\s6_data_i[28] );
  assign \new_[27337]_  = \new_[30510]_  & \new_[28974]_ ;
  assign \new_[27338]_  = (~\new_[29961]_  | ~\s4_data_i[28] ) & (~\new_[29819]_  | ~\s0_data_i[28] );
  assign \new_[27339]_  = (~\new_[30113]_  | ~\s2_data_i[3] ) & (~\new_[30124]_  | ~\s1_data_i[3] );
  assign \new_[27340]_  = (~\new_[30166]_  | ~\s14_data_i[15] ) & (~\new_[30298]_  | ~\s12_data_i[15] );
  assign \new_[27341]_  = \new_[30363]_  & \new_[6080]_ ;
  assign \new_[27342]_  = (~\new_[29807]_  | ~\s14_data_i[1] ) & (~\new_[30626]_  | ~\s12_data_i[1] );
  assign \new_[27343]_  = (~\new_[30113]_  | ~\s2_data_i[15] ) & (~\new_[30124]_  | ~\s1_data_i[15] );
  assign \new_[27344]_  = (~\new_[30189]_  | ~\s2_data_i[18] ) & (~\new_[30195]_  | ~\s1_data_i[18] );
  assign \new_[27345]_  = (~\new_[29846]_  | ~\s2_data_i[28] ) & (~\new_[30001]_  | ~\s1_data_i[28] );
  assign \new_[27346]_  = (~\new_[30013]_  | ~\s2_data_i[29] ) & (~\new_[29769]_  | ~\s1_data_i[29] );
  assign \new_[27347]_  = \new_[28974]_  & \new_[30990]_ ;
  assign \new_[27348]_  = (~\new_[29807]_  | ~\s14_data_i[17] ) & (~\new_[30626]_  | ~\s12_data_i[17] );
  assign \new_[27349]_  = (~\new_[29961]_  | ~\s4_data_i[8] ) & (~\new_[29819]_  | ~\s0_data_i[8] );
  assign \new_[27350]_  = (~\new_[30088]_  | ~\s2_data_i[27] ) & (~\new_[29779]_  | ~\s1_data_i[27] );
  assign \new_[27351]_  = (~\new_[30189]_  | ~\s2_data_i[17] ) & (~\new_[30195]_  | ~\s1_data_i[17] );
  assign \new_[27352]_  = (~\new_[29846]_  | ~\s2_data_i[15] ) & (~\new_[30001]_  | ~\s1_data_i[15] );
  assign \new_[27353]_  = ~\new_[29576]_  & ~\new_[29777]_ ;
  assign \new_[27354]_  = (~\new_[29963]_  | ~\s4_data_i[17] ) & (~\new_[30481]_  | ~\s0_data_i[17] );
  assign \new_[27355]_  = (~\new_[30131]_  | ~\s7_data_i[22] ) & (~\new_[29939]_  | ~\s6_data_i[22] );
  assign \new_[27356]_  = ~\new_[29955]_  & ~\new_[28640]_ ;
  assign \new_[27357]_  = (~\new_[29948]_  | ~\s5_data_i[20] ) & (~\new_[29947]_  | ~\s3_data_i[20] );
  assign \new_[27358]_  = (~\new_[30013]_  | ~\s2_data_i[30] ) & (~\new_[29769]_  | ~\s1_data_i[30] );
  assign \new_[27359]_  = ~\new_[28376]_ ;
  assign \new_[27360]_  = ~\new_[28703]_ ;
  assign \new_[27361]_  = (~\new_[29846]_  | ~\s2_data_i[29] ) & (~\new_[30001]_  | ~\s1_data_i[29] );
  assign \new_[27362]_  = (~\new_[30088]_  | ~\s2_data_i[23] ) & (~\new_[29779]_  | ~\s1_data_i[23] );
  assign \new_[27363]_  = ~\new_[29246]_  | ~\new_[31235]_ ;
  assign \new_[27364]_  = (~\new_[30189]_  | ~\s2_data_i[14] ) & (~\new_[30195]_  | ~\s1_data_i[14] );
  assign \new_[27365]_  = ~\new_[28572]_ ;
  assign \new_[27366]_  = (~\new_[30088]_  | ~\s2_data_i[22] ) & (~\new_[29779]_  | ~\s1_data_i[22] );
  assign \new_[27367]_  = (~\new_[29876]_  | ~\s11_data_i[18] ) & (~\new_[30341]_  | ~\s8_data_i[18] );
  assign \new_[27368]_  = (~\new_[29963]_  | ~\s4_data_i[7] ) & (~\new_[30481]_  | ~\s0_data_i[7] );
  assign \new_[27369]_  = (~\new_[30189]_  | ~\s2_data_i[13] ) & (~\new_[30195]_  | ~\s1_data_i[13] );
  assign \new_[27370]_  = (~\new_[30088]_  | ~\s2_data_i[21] ) & (~\new_[29779]_  | ~\s1_data_i[21] );
  assign \new_[27371]_  = ~\new_[28249]_  | ~\new_[5895]_ ;
  assign \new_[27372]_  = ~\new_[28821]_  | ~\new_[31423]_ ;
  assign \new_[27373]_  = (~\new_[30189]_  | ~\s2_data_i[12] ) & (~\new_[30195]_  | ~\s1_data_i[12] );
  assign \new_[27374]_  = (~\new_[30131]_  | ~\s7_data_i[0] ) & (~\new_[29939]_  | ~\s6_data_i[0] );
  assign \new_[27375]_  = ~\new_[29676]_  | ~\new_[29900]_ ;
  assign \new_[27376]_  = (~\new_[30088]_  | ~\s2_data_i[18] ) & (~\new_[29779]_  | ~\s1_data_i[18] );
  assign \new_[27377]_  = \new_[29344]_  & \new_[30011]_ ;
  assign \new_[27378]_  = ~\new_[29758]_  & ~\new_[29560]_ ;
  assign \new_[27379]_  = ~\new_[28321]_ ;
  assign \new_[27380]_  = (~\new_[30088]_  | ~\s2_data_i[17] ) & (~\new_[29779]_  | ~\s1_data_i[17] );
  assign \new_[27381]_  = (~\new_[30166]_  | ~\s14_data_i[4] ) & (~\new_[30298]_  | ~\s12_data_i[4] );
  assign \new_[27382]_  = (~\new_[29876]_  | ~\s11_data_i[19] ) & (~\new_[30341]_  | ~\s8_data_i[19] );
  assign \new_[27383]_  = ~\new_[30375]_  | ~\new_[29050]_ ;
  assign \new_[27384]_  = ~\new_[30245]_ ;
  assign \new_[27385]_  = (~\new_[30088]_  | ~\s2_data_i[15] ) & (~\new_[29779]_  | ~\s1_data_i[15] );
  assign \new_[27386]_  = (~\new_[29948]_  | ~\s5_data_i[5] ) & (~\new_[29947]_  | ~\s3_data_i[5] );
  assign \new_[27387]_  = (~\new_[29948]_  | ~\s5_data_i[23] ) & (~\new_[29947]_  | ~\s3_data_i[23] );
  assign \new_[27388]_  = ~\new_[30209]_  & ~\new_[28039]_ ;
  assign \new_[27389]_  = (~\new_[29963]_  | ~\s4_data_i[19] ) & (~\new_[30481]_  | ~\s0_data_i[19] );
  assign \new_[27390]_  = (~\new_[29846]_  | ~\s2_data_i[20] ) & (~\new_[30001]_  | ~\s1_data_i[20] );
  assign \new_[27391]_  = (~\new_[30166]_  | ~\s14_data_i[10] ) & (~\new_[30298]_  | ~\s12_data_i[10] );
  assign \new_[27392]_  = ~\new_[28982]_  | ~\new_[28962]_ ;
  assign \new_[27393]_  = (~\new_[30189]_  | ~\s2_data_i[8] ) & (~\new_[30195]_  | ~\s1_data_i[8] );
  assign \new_[27394]_  = ~\new_[29228]_  | ~\new_[6045]_ ;
  assign \new_[27395]_  = ~\new_[28753]_ ;
  assign \new_[27396]_  = (~\new_[29876]_  | ~\s11_data_i[20] ) & (~\new_[30341]_  | ~\s8_data_i[20] );
  assign \new_[27397]_  = (~\new_[30113]_  | ~\s2_data_i[31] ) & (~\new_[30124]_  | ~\s1_data_i[31] );
  assign \new_[27398]_  = (~\new_[29961]_  | ~\s4_data_i[20] ) & (~\new_[29819]_  | ~\s0_data_i[20] );
  assign \new_[27399]_  = (~\new_[29788]_  | ~\s2_data_i[20] ) & (~\new_[30357]_  | ~\s1_data_i[20] );
  assign \new_[27400]_  = (~\new_[30189]_  | ~\s2_data_i[7] ) & (~\new_[30195]_  | ~\s1_data_i[7] );
  assign \new_[27401]_  = ~\new_[28571]_ ;
  assign \new_[27402]_  = ~\new_[28849]_  | ~\new_[31406]_ ;
  assign \new_[27403]_  = ~\new_[28283]_  | ~\new_[31429]_ ;
  assign \new_[27404]_  = (~\new_[30113]_  | ~\s2_data_i[26] ) & (~\new_[30124]_  | ~\s1_data_i[26] );
  assign \new_[27405]_  = (~\new_[30189]_  | ~\s2_data_i[6] ) & (~\new_[30195]_  | ~\s1_data_i[6] );
  assign \new_[27406]_  = (~\new_[29807]_  | ~\s14_data_i[27] ) & (~\new_[30626]_  | ~\s12_data_i[27] );
  assign \new_[27407]_  = ~\new_[28216]_ ;
  assign \new_[27408]_  = (~\new_[29876]_  | ~\s11_data_i[21] ) & (~\new_[30341]_  | ~\s8_data_i[21] );
  assign \new_[27409]_  = (~\new_[30088]_  | ~\s2_data_i[6] ) & (~\new_[29779]_  | ~\s1_data_i[6] );
  assign \new_[27410]_  = ~\new_[28930]_  | ~\new_[29887]_ ;
  assign \new_[27411]_  = (~\new_[29948]_  | ~\s5_data_i[18] ) & (~\new_[29947]_  | ~\s3_data_i[18] );
  assign \new_[27412]_  = (~\new_[30088]_  | ~\s2_data_i[5] ) & (~\new_[29779]_  | ~\s1_data_i[5] );
  assign \new_[27413]_  = (~\new_[29788]_  | ~\s2_data_i[21] ) & (~\new_[30357]_  | ~\s1_data_i[21] );
  assign \new_[27414]_  = (~\new_[30013]_  | ~\s2_data_i[8] ) & (~\new_[29769]_  | ~\s1_data_i[8] );
  assign \new_[27415]_  = (~\new_[29963]_  | ~\s4_data_i[9] ) & (~\new_[30481]_  | ~\s0_data_i[9] );
  assign \new_[27416]_  = (~\new_[30088]_  | ~\s2_data_i[4] ) & (~\new_[29779]_  | ~\s1_data_i[4] );
  assign \new_[27417]_  = (~\new_[29949]_  | ~\s10_data_i[19] ) & (~\new_[29905]_  | ~\s9_data_i[19] );
  assign \new_[27418]_  = ~\new_[28400]_ ;
  assign \new_[27419]_  = (~\new_[29963]_  | ~\s4_data_i[21] ) & (~\new_[30481]_  | ~\s0_data_i[21] );
  assign \new_[27420]_  = (~\new_[30088]_  | ~\s2_data_i[3] ) & (~\new_[29779]_  | ~\s1_data_i[3] );
  assign \new_[27421]_  = (~\new_[29949]_  | ~\s10_data_i[6] ) & (~\new_[29905]_  | ~\s9_data_i[6] );
  assign \new_[27422]_  = (~\new_[30088]_  | ~\s2_data_i[2] ) & (~\new_[29779]_  | ~\s1_data_i[2] );
  assign \new_[27423]_  = (~\new_[29963]_  | ~\s4_data_i[25] ) & (~\new_[30481]_  | ~\s0_data_i[25] );
  assign \new_[27424]_  = (~\new_[30131]_  | ~\s7_data_i[21] ) & (~\new_[29939]_  | ~\s6_data_i[21] );
  assign \new_[27425]_  = ~\new_[28655]_ ;
  assign \new_[27426]_  = \new_[28959]_  & \new_[30724]_ ;
  assign \new_[27427]_  = ~\new_[29079]_ ;
  assign \new_[27428]_  = (~\new_[30088]_  | ~\s2_data_i[31] ) & (~\new_[29779]_  | ~\s1_data_i[31] );
  assign \new_[27429]_  = (~\new_[30013]_  | ~\s2_data_i[2] ) & (~\new_[29769]_  | ~\s1_data_i[2] );
  assign \new_[27430]_  = (~\new_[29949]_  | ~\s10_data_i[2] ) & (~\new_[29905]_  | ~\s9_data_i[2] );
  assign \new_[27431]_  = ~\new_[30730]_  | ~\new_[29722]_ ;
  assign \new_[27432]_  = (~\new_[30189]_  | ~\s2_data_i[23] ) & (~\new_[30195]_  | ~\s1_data_i[23] );
  assign \new_[27433]_  = (~\new_[30189]_  | ~\s2_data_i[25] ) & (~\new_[30195]_  | ~\s1_data_i[25] );
  assign \new_[27434]_  = (~\new_[30013]_  | ~\s2_data_i[31] ) & (~\new_[29769]_  | ~\s1_data_i[31] );
  assign \new_[27435]_  = (~\new_[30189]_  | ~\s2_data_i[20] ) & (~\new_[30195]_  | ~\s1_data_i[20] );
  assign \new_[27436]_  = (~\new_[29961]_  | ~\s4_data_i[0] ) & (~\new_[29819]_  | ~\s0_data_i[0] );
  assign \new_[27437]_  = ~\new_[29784]_  & ~\new_[29550]_ ;
  assign \new_[27438]_  = (~\new_[30113]_  | ~\s2_data_i[20] ) & (~\new_[30124]_  | ~\s1_data_i[20] );
  assign \new_[27439]_  = ~\new_[28260]_ ;
  assign \new_[27440]_  = (~\new_[30013]_  | ~\s2_data_i[26] ) & (~\new_[29769]_  | ~\s1_data_i[26] );
  assign \new_[27441]_  = \new_[29268]_  & \new_[6083]_ ;
  assign \new_[27442]_  = ~\new_[29375]_  & ~\new_[30627]_ ;
  assign \new_[27443]_  = (~\new_[30189]_  | ~\s2_data_i[21] ) & (~\new_[30195]_  | ~\s1_data_i[21] );
  assign \new_[27444]_  = (~\new_[30189]_  | ~\s2_data_i[2] ) & (~\new_[30195]_  | ~\s1_data_i[2] );
  assign \new_[27445]_  = (~\new_[30013]_  | ~\s2_data_i[23] ) & (~\new_[29769]_  | ~\s1_data_i[23] );
  assign \new_[27446]_  = (~\new_[29948]_  | ~\s5_data_i[22] ) & (~\new_[29947]_  | ~\s3_data_i[22] );
  assign \new_[27447]_  = ~\new_[28419]_ ;
  assign \new_[27448]_  = (~\new_[30113]_  | ~\s2_data_i[21] ) & (~\new_[30124]_  | ~\s1_data_i[21] );
  assign \new_[27449]_  = ~\new_[28805]_ ;
  assign \new_[27450]_  = (~\new_[30013]_  | ~\s2_data_i[22] ) & (~\new_[29769]_  | ~\s1_data_i[22] );
  assign \new_[27451]_  = (~\new_[29963]_  | ~\s4_data_i[31] ) & (~\new_[30481]_  | ~\s0_data_i[31] );
  assign \new_[27452]_  = (~\new_[29961]_  | ~\s4_data_i[2] ) & (~\new_[29819]_  | ~\s0_data_i[2] );
  assign \new_[27453]_  = (~\new_[29846]_  | ~\s2_data_i[21] ) & (~\new_[30001]_  | ~\s1_data_i[21] );
  assign \new_[27454]_  = (~\new_[30013]_  | ~\s2_data_i[21] ) & (~\new_[29769]_  | ~\s1_data_i[21] );
  assign \new_[27455]_  = (~\new_[30013]_  | ~\s2_data_i[20] ) & (~\new_[29769]_  | ~\s1_data_i[20] );
  assign \new_[27456]_  = (~\new_[29948]_  | ~\s5_data_i[3] ) & (~\new_[29947]_  | ~\s3_data_i[3] );
  assign \new_[27457]_  = (~\new_[30166]_  | ~\s14_data_i[3] ) & (~\new_[30298]_  | ~\s12_data_i[3] );
  assign \new_[27458]_  = ~\new_[6206]_  | ~\new_[30255]_  | ~\new_[30721]_ ;
  assign \new_[27459]_  = (~\new_[29807]_  | ~\s14_data_i[24] ) & (~\new_[30626]_  | ~\s12_data_i[24] );
  assign \new_[27460]_  = (~\new_[29876]_  | ~\s11_data_i[30] ) & (~\new_[30341]_  | ~\s8_data_i[30] );
  assign \new_[27461]_  = (~\new_[29807]_  | ~\s14_data_i[30] ) & (~\new_[30626]_  | ~\s12_data_i[30] );
  assign \new_[27462]_  = (~\new_[29846]_  | ~\s2_data_i[3] ) & (~\new_[30001]_  | ~\s1_data_i[3] );
  assign \new_[27463]_  = ~\new_[28421]_ ;
  assign \new_[27464]_  = ~\new_[29695]_  | ~\new_[6075]_ ;
  assign \new_[27465]_  = ~\new_[28422]_ ;
  assign \new_[27466]_  = ~\new_[28424]_ ;
  assign \new_[27467]_  = (~\new_[30131]_  | ~\s7_data_i[9] ) & (~\new_[29939]_  | ~\s6_data_i[9] );
  assign \new_[27468]_  = (~\new_[29788]_  | ~\s2_data_i[28] ) & (~\new_[30357]_  | ~\s1_data_i[28] );
  assign \new_[27469]_  = (~\new_[29961]_  | ~\s4_data_i[22] ) & (~\new_[29819]_  | ~\s0_data_i[22] );
  assign \new_[27470]_  = (~\new_[29807]_  | ~\s14_data_i[28] ) & (~\new_[30626]_  | ~\s12_data_i[28] );
  assign \new_[27471]_  = (~\new_[30131]_  | ~\s7_data_i[12] ) & (~\new_[29939]_  | ~\s6_data_i[12] );
  assign \new_[27472]_  = (~\new_[30013]_  | ~\s2_data_i[13] ) & (~\new_[29769]_  | ~\s1_data_i[13] );
  assign \new_[27473]_  = (~\new_[29963]_  | ~\s4_data_i[27] ) & (~\new_[30481]_  | ~\s0_data_i[27] );
  assign \new_[27474]_  = ~\new_[28984]_  & ~\new_[30170]_ ;
  assign \new_[27475]_  = (~\new_[29788]_  | ~\s2_data_i[27] ) & (~\new_[30357]_  | ~\s1_data_i[27] );
  assign \new_[27476]_  = (~\new_[29876]_  | ~\s11_data_i[27] ) & (~\new_[30341]_  | ~\s8_data_i[27] );
  assign \new_[27477]_  = (~\new_[30166]_  | ~\s14_data_i[11] ) & (~\new_[30298]_  | ~\s12_data_i[11] );
  assign \new_[27478]_  = (~\new_[29788]_  | ~\s2_data_i[24] ) & (~\new_[30357]_  | ~\s1_data_i[24] );
  assign \new_[27479]_  = (~\new_[29963]_  | ~\s4_data_i[26] ) & (~\new_[30481]_  | ~\s0_data_i[26] );
  assign \new_[27480]_  = (~\new_[30131]_  | ~\s7_data_i[19] ) & (~\new_[29939]_  | ~\s6_data_i[19] );
  assign \new_[27481]_  = ~\new_[28481]_ ;
  assign \new_[27482]_  = (~\new_[30013]_  | ~\s2_data_i[10] ) & (~\new_[29769]_  | ~\s1_data_i[10] );
  assign \new_[27483]_  = (~\new_[30113]_  | ~\s2_data_i[22] ) & (~\new_[30124]_  | ~\s1_data_i[22] );
  assign \new_[27484]_  = (~\new_[29949]_  | ~\s10_data_i[22] ) & (~\new_[29905]_  | ~\s9_data_i[22] );
  assign \new_[27485]_  = (~\new_[29807]_  | ~\s14_data_i[25] ) & (~\new_[30626]_  | ~\s12_data_i[25] );
  assign \new_[27486]_  = (~\new_[29948]_  | ~\s5_data_i[12] ) & (~\new_[29947]_  | ~\s3_data_i[12] );
  assign \new_[27487]_  = ~\new_[28545]_ ;
  assign \new_[27488]_  = ~\new_[29729]_  & ~\new_[29962]_ ;
  assign \new_[27489]_  = ~\new_[29235]_  | ~\new_[5905]_ ;
  assign \new_[27490]_  = ~\new_[30613]_  | ~\new_[5984]_ ;
  assign \new_[27491]_  = ~\new_[28849]_  | ~\new_[31121]_ ;
  assign \new_[27492]_  = ~\new_[29721]_  | ~\new_[6193]_ ;
  assign \new_[27493]_  = ~\new_[30586]_  | ~\new_[6092]_ ;
  assign \new_[27494]_  = \new_[29744]_  & \new_[6087]_ ;
  assign \new_[27495]_  = ~\new_[29320]_  | ~\new_[6042]_ ;
  assign \new_[27496]_  = \new_[29350]_  & \new_[6091]_ ;
  assign \new_[27497]_  = ~\new_[29226]_  | ~\new_[6091]_ ;
  assign \new_[27498]_  = ~\new_[29103]_  | ~\new_[6051]_ ;
  assign \new_[27499]_  = ~\new_[28070]_  | ~\new_[5897]_ ;
  assign \new_[27500]_  = \new_[28939]_  & \new_[6067]_ ;
  assign \new_[27501]_  = ~\new_[30446]_  & ~\new_[31165]_ ;
  assign \new_[27502]_  = ~\new_[29728]_  | ~\new_[5923]_ ;
  assign \new_[27503]_  = ~\new_[29590]_  | ~\new_[31232]_ ;
  assign \new_[27504]_  = ~\new_[30608]_  | ~\new_[31440]_ ;
  assign \new_[27505]_  = ~\new_[28621]_ ;
  assign \new_[27506]_  = ~\new_[30557]_  & ~\new_[30755]_ ;
  assign \new_[27507]_  = ~\new_[30763]_  | ~\new_[6040]_ ;
  assign \new_[27508]_  = ~\new_[28489]_ ;
  assign \new_[27509]_  = \new_[28887]_  & \new_[6193]_ ;
  assign \new_[27510]_  = ~\new_[28813]_ ;
  assign \new_[27511]_  = \new_[28883]_  & \new_[6051]_ ;
  assign \new_[27512]_  = \new_[29324]_  & \new_[5925]_ ;
  assign \new_[27513]_  = ~\new_[28828]_  | ~\new_[6062]_ ;
  assign \new_[27514]_  = ~\new_[30680]_  | ~\new_[6072]_ ;
  assign \new_[27515]_  = \new_[30767]_  & \new_[5970]_ ;
  assign \new_[27516]_  = ~\new_[30623]_  | ~\new_[6096]_ ;
  assign \new_[27517]_  = \new_[28924]_  & \new_[6075]_ ;
  assign \new_[27518]_  = ~\new_[29079]_  & ~\new_[29597]_ ;
  assign \new_[27519]_  = ~\new_[29342]_  & ~\m3_addr_i[28] ;
  assign \new_[27520]_  = (~\new_[29823]_  | ~\s7_data_i[1] ) & (~\new_[29954]_  | ~\s6_data_i[1] );
  assign \new_[27521]_  = \new_[28962]_  & \new_[6056]_ ;
  assign \new_[27522]_  = (~\new_[29823]_  | ~\s7_data_i[24] ) & (~\new_[29954]_  | ~\s6_data_i[24] );
  assign \new_[27523]_  = (~\new_[29788]_  | ~\s2_data_i[15] ) & (~\new_[30357]_  | ~\s1_data_i[15] );
  assign \new_[27524]_  = ~\new_[29456]_  | ~\new_[6083]_ ;
  assign \new_[27525]_  = ~\new_[28676]_ ;
  assign \new_[27526]_  = ~\new_[29588]_  | ~\new_[5903]_ ;
  assign \new_[27527]_  = \new_[29436]_  & \new_[30213]_ ;
  assign \new_[27528]_  = ~\new_[28963]_  | ~\new_[6067]_ ;
  assign \new_[27529]_  = \new_[28872]_  & \new_[6042]_ ;
  assign \new_[27530]_  = ~\new_[29736]_  & ~\new_[29192]_ ;
  assign \new_[27531]_  = ~\new_[30735]_  | ~\new_[6217]_ ;
  assign \new_[27532]_  = ~\new_[29032]_  | ~\new_[5913]_ ;
  assign \new_[27533]_  = ~\new_[29455]_  | ~\new_[30021]_ ;
  assign \new_[27534]_  = ~\new_[28889]_  & ~\new_[29918]_ ;
  assign \new_[27535]_  = \new_[32049]_  & m2_stb_i;
  assign \new_[27536]_  = ~\new_[28837]_  | ~\new_[6031]_ ;
  assign \new_[27537]_  = ~\new_[30696]_  | ~\new_[28888]_ ;
  assign \new_[27538]_  = \new_[29715]_  & \new_[31458]_ ;
  assign \new_[27539]_  = ~\new_[28476]_ ;
  assign \new_[27540]_  = ~\new_[28298]_ ;
  assign \new_[27541]_  = \new_[28837]_  & \new_[6052]_ ;
  assign \new_[27542]_  = ~\new_[29061]_  | ~\new_[5994]_ ;
  assign \new_[27543]_  = ~\new_[28478]_ ;
  assign \new_[27544]_  = ~\new_[29172]_  & ~\new_[29861]_ ;
  assign \new_[27545]_  = ~\new_[28289]_ ;
  assign \new_[27546]_  = ~\new_[28988]_  & ~\new_[28830]_ ;
  assign \new_[27547]_  = ~\new_[29387]_  | ~\new_[30784]_ ;
  assign \new_[27548]_  = ~\new_[30755]_  & ~\new_[30157]_ ;
  assign \new_[27549]_  = ~\new_[28115]_ ;
  assign \new_[27550]_  = ~\new_[28286]_ ;
  assign \new_[27551]_  = ~\new_[28123]_ ;
  assign \new_[27552]_  = ~\new_[30236]_  | ~\new_[29692]_ ;
  assign \new_[27553]_  = ~\new_[29582]_  & ~\new_[29772]_ ;
  assign \new_[27554]_  = (~\new_[30166]_  | ~\s14_data_i[29] ) & (~\new_[30298]_  | ~\s12_data_i[29] );
  assign \new_[27555]_  = ~\new_[29906]_  & ~\new_[28355]_ ;
  assign \new_[27556]_  = ~\new_[28968]_  | ~\new_[29765]_ ;
  assign \new_[27557]_  = ~\new_[30724]_  | ~\new_[28830]_ ;
  assign \new_[27558]_  = ~\new_[29222]_  & ~\new_[28877]_ ;
  assign \new_[27559]_  = ~\new_[29113]_  & ~\new_[28935]_ ;
  assign \new_[27560]_  = ~\new_[29608]_  | ~\new_[5998]_ ;
  assign \new_[27561]_  = ~\new_[28076]_  & ~\new_[28977]_ ;
  assign \new_[27562]_  = ~\new_[29743]_  & ~\new_[29435]_ ;
  assign \new_[27563]_  = \new_[30271]_  & \new_[29798]_ ;
  assign \new_[27564]_  = ~\new_[29886]_  | ~\new_[29266]_ ;
  assign \new_[27565]_  = ~\new_[29043]_  | ~m0_stb_i;
  assign \new_[27566]_  = ~\new_[29225]_  | ~\new_[29787]_ ;
  assign \new_[27567]_  = ~\new_[29563]_  | ~\new_[6003]_ ;
  assign \new_[27568]_  = ~\new_[28829]_  & ~\new_[30216]_ ;
  assign \new_[27569]_  = (~\new_[29961]_  | ~\s4_data_i[9] ) & (~\new_[29819]_  | ~\s0_data_i[9] );
  assign \new_[27570]_  = ~\new_[30733]_  & ~\new_[28837]_ ;
  assign \new_[27571]_  = ~\new_[28969]_  & ~\new_[30327]_ ;
  assign \new_[27572]_  = ~\new_[28259]_ ;
  assign \new_[27573]_  = \new_[30322]_  & \new_[30152]_ ;
  assign \new_[27574]_  = ~\new_[29397]_  | ~\new_[29977]_ ;
  assign \new_[27575]_  = ~\new_[30275]_  & ~\new_[30680]_ ;
  assign \new_[27576]_  = ~\new_[29602]_  | ~\new_[30355]_ ;
  assign \new_[27577]_  = ~\new_[29013]_  & ~\new_[28834]_ ;
  assign \new_[27578]_  = ~\new_[30078]_  | ~\new_[29560]_ ;
  assign \new_[27579]_  = \new_[29015]_  & \new_[6060]_ ;
  assign \new_[27580]_  = ~\new_[30599]_  & ~\new_[29650]_ ;
  assign \new_[27581]_  = ~\new_[28565]_ ;
  assign \new_[27582]_  = ~\new_[30058]_  & ~\new_[29248]_ ;
  assign \new_[27583]_  = ~\new_[28241]_ ;
  assign \new_[27584]_  = ~\new_[28240]_ ;
  assign \new_[27585]_  = ~\new_[29676]_  & ~\new_[30042]_ ;
  assign \new_[27586]_  = \new_[29046]_  & \m4_addr_i[28] ;
  assign \new_[27587]_  = ~\new_[28499]_ ;
  assign \new_[27588]_  = ~\new_[29166]_  | ~\new_[29350]_ ;
  assign \new_[27589]_  = ~\new_[29350]_  | ~\new_[29774]_ ;
  assign \new_[27590]_  = (~\new_[30113]_  | ~\s2_data_i[13] ) & (~\new_[30124]_  | ~\s1_data_i[13] );
  assign \new_[27591]_  = ~\new_[30678]_  & ~\new_[30633]_ ;
  assign \new_[27592]_  = ~\new_[28815]_ ;
  assign \new_[27593]_  = ~\new_[28960]_  & ~\new_[30644]_ ;
  assign \new_[27594]_  = ~\new_[28191]_  & ~\new_[29960]_ ;
  assign \new_[27595]_  = ~\new_[28113]_ ;
  assign \new_[27596]_  = ~\new_[29384]_  & ~\new_[29946]_ ;
  assign \new_[27597]_  = ~\new_[30525]_  & ~\new_[29806]_ ;
  assign \new_[27598]_  = (~\new_[29846]_  | ~\s2_data_i[18] ) & (~\new_[30001]_  | ~\s1_data_i[18] );
  assign \new_[27599]_  = \new_[29422]_  | \new_[30526]_ ;
  assign \new_[27600]_  = ~\new_[28398]_ ;
  assign \new_[27601]_  = ~\new_[29783]_  & ~\new_[29360]_ ;
  assign \new_[27602]_  = \new_[29217]_  | \new_[30057]_ ;
  assign \new_[27603]_  = (~\new_[30131]_  | ~\s7_data_i[8] ) & (~\new_[29939]_  | ~\s6_data_i[8] );
  assign \new_[27604]_  = ~\new_[30616]_  & ~\new_[30731]_ ;
  assign \new_[27605]_  = ~\new_[28514]_ ;
  assign \new_[27606]_  = ~\new_[28407]_ ;
  assign \new_[27607]_  = (~\new_[29846]_  | ~\s2_data_i[19] ) & (~\new_[30001]_  | ~\s1_data_i[19] );
  assign \new_[27608]_  = ~\new_[29931]_  | ~\new_[29103]_ ;
  assign \new_[27609]_  = ~\new_[29101]_  & ~\new_[30058]_ ;
  assign \new_[27610]_  = ~\new_[30301]_  & ~\new_[28684]_ ;
  assign \new_[27611]_  = ~\new_[30544]_  | ~\new_[6090]_ ;
  assign \new_[27612]_  = ~\new_[28139]_ ;
  assign \new_[27613]_  = ~\new_[30212]_  | ~\new_[29721]_ ;
  assign \new_[27614]_  = ~\new_[28167]_ ;
  assign \new_[27615]_  = ~\new_[28519]_ ;
  assign \new_[27616]_  = ~\new_[28520]_ ;
  assign \new_[27617]_  = ~\new_[28164]_ ;
  assign \new_[27618]_  = ~\new_[28160]_ ;
  assign \new_[27619]_  = ~\new_[29744]_  | ~\new_[29745]_ ;
  assign \new_[27620]_  = ~\new_[30217]_  | ~\new_[28909]_ ;
  assign \new_[27621]_  = ~\new_[30053]_  | ~\new_[28963]_ ;
  assign \new_[27622]_  = ~\new_[30299]_  & ~\new_[29564]_ ;
  assign \new_[27623]_  = ~\new_[30670]_  | ~\new_[6069]_ ;
  assign \new_[27624]_  = ~\new_[29086]_  & ~\new_[30413]_ ;
  assign \new_[27625]_  = ~\new_[28150]_ ;
  assign \new_[27626]_  = ~\new_[28137]_ ;
  assign \new_[27627]_  = ~\new_[28707]_ ;
  assign \new_[27628]_  = ~\new_[29656]_  & ~\new_[30129]_ ;
  assign \new_[27629]_  = ~\new_[30333]_  & ~\new_[29672]_ ;
  assign \new_[27630]_  = ~\new_[30038]_  & ~\new_[30608]_ ;
  assign \new_[27631]_  = \new_[30058]_  | \new_[29648]_ ;
  assign \new_[27632]_  = ~\new_[30114]_  | ~\new_[29695]_ ;
  assign \new_[27633]_  = ~\new_[28111]_ ;
  assign \new_[27634]_  = ~\new_[29508]_  & ~\new_[30725]_ ;
  assign \new_[27635]_  = ~\new_[29371]_  & ~\new_[29256]_ ;
  assign \new_[27636]_  = ~\new_[29357]_  | ~\new_[29748]_ ;
  assign \new_[27637]_  = ~\new_[30557]_  & ~\new_[30367]_ ;
  assign \new_[27638]_  = ~\new_[30204]_  & ~\new_[29186]_ ;
  assign \new_[27639]_  = ~\new_[29861]_  & ~\new_[29357]_ ;
  assign \new_[27640]_  = ~\new_[28462]_ ;
  assign \new_[27641]_  = ~\new_[30058]_  | ~\new_[29006]_ ;
  assign \new_[27642]_  = ~\new_[29169]_  | ~\new_[29233]_ ;
  assign \new_[27643]_  = ~\new_[28072]_ ;
  assign \new_[27644]_  = ~\new_[30140]_  | ~\new_[29456]_ ;
  assign \new_[27645]_  = (~\new_[30189]_  | ~\s2_data_i[31] ) & (~\new_[30195]_  | ~\s1_data_i[31] );
  assign \new_[27646]_  = ~\new_[30251]_  | ~\new_[29139]_ ;
  assign \new_[27647]_  = ~\new_[28065]_ ;
  assign \new_[27648]_  = ~\new_[29290]_  | ~\new_[30125]_ ;
  assign \new_[27649]_  = ~\new_[29367]_  & ~\new_[30727]_ ;
  assign \new_[27650]_  = ~\new_[28000]_ ;
  assign \new_[27651]_  = ~\new_[29192]_  | ~\new_[5969]_ ;
  assign \new_[27652]_  = ~\new_[29455]_  | ~\new_[6005]_ ;
  assign \new_[27653]_  = ~\new_[29808]_  | ~\new_[30723]_ ;
  assign \new_[27654]_  = ~\new_[28604]_ ;
  assign \new_[27655]_  = ~\new_[29571]_  | ~\new_[6000]_ ;
  assign \new_[27656]_  = ~\new_[28877]_  | ~\new_[5982]_ ;
  assign \new_[27657]_  = ~\new_[28539]_ ;
  assign \new_[27658]_  = ~\new_[28353]_ ;
  assign \new_[27659]_  = ~\new_[29907]_  & ~\new_[30763]_ ;
  assign \new_[27660]_  = ~\new_[29588]_  | ~\new_[29619]_ ;
  assign \new_[27661]_  = ~\new_[29038]_  | ~\new_[5997]_ ;
  assign \new_[27662]_  = ~\new_[27976]_ ;
  assign \new_[27663]_  = ~\new_[29238]_  & ~\new_[30775]_ ;
  assign \new_[27664]_  = ~\new_[28425]_ ;
  assign \new_[27665]_  = ~\new_[28811]_ ;
  assign \new_[27666]_  = ~\new_[28543]_ ;
  assign \new_[27667]_  = ~\new_[28808]_ ;
  assign \new_[27668]_  = (~\new_[29876]_  | ~\s11_data_i[17] ) & (~\new_[30341]_  | ~\s8_data_i[17] );
  assign \new_[27669]_  = ~\new_[28800]_ ;
  assign \new_[27670]_  = ~\new_[28797]_ ;
  assign \new_[27671]_  = ~\new_[29401]_  | ~\new_[5830]_ ;
  assign \new_[27672]_  = ~\new_[30326]_  | ~\new_[30613]_ ;
  assign \new_[27673]_  = ~\new_[28745]_ ;
  assign \new_[27674]_  = ~\new_[30575]_  | ~\new_[29746]_ ;
  assign \new_[27675]_  = ~\new_[28884]_  & ~\new_[30707]_ ;
  assign \new_[27676]_  = ~\new_[28727]_ ;
  assign \new_[27677]_  = ~\new_[28700]_ ;
  assign \new_[27678]_  = ~\new_[29159]_  | ~\new_[5966]_ ;
  assign \new_[27679]_  = ~\new_[30118]_  & ~\new_[28732]_ ;
  assign \new_[27680]_  = ~\new_[29169]_  & ~\new_[29212]_ ;
  assign \new_[27681]_  = (~\new_[29846]_  | ~\s2_data_i[5] ) & (~\new_[30001]_  | ~\s1_data_i[5] );
  assign \new_[27682]_  = ~\new_[29792]_  | ~\new_[30578]_ ;
  assign \new_[27683]_  = ~\new_[28654]_ ;
  assign \new_[27684]_  = (~\new_[29961]_  | ~\s4_data_i[31] ) & (~\new_[29819]_  | ~\s0_data_i[31] );
  assign \new_[27685]_  = \new_[28967]_  & \new_[6065]_ ;
  assign \new_[27686]_  = ~\new_[29159]_  | ~\new_[30508]_ ;
  assign \new_[27687]_  = \new_[29171]_  & \new_[5982]_ ;
  assign \new_[27688]_  = (~\new_[30013]_  | ~\s2_data_i[7] ) & (~\new_[29769]_  | ~\s1_data_i[7] );
  assign \new_[27689]_  = ~\new_[29277]_  & ~\new_[28280]_ ;
  assign \new_[27690]_  = ~\new_[30054]_  & ~\new_[29629]_ ;
  assign \new_[27691]_  = ~\new_[29359]_  & ~\new_[29266]_ ;
  assign \new_[27692]_  = ~\new_[30229]_  | ~\new_[30426]_ ;
  assign \new_[27693]_  = ~\new_[28546]_ ;
  assign \new_[27694]_  = ~\new_[28999]_  | ~\new_[30147]_ ;
  assign \new_[27695]_  = ~\new_[30769]_  | ~\new_[29251]_ ;
  assign \new_[27696]_  = ~\new_[29785]_  | ~\new_[28977]_ ;
  assign \new_[27697]_  = ~\new_[29773]_  & ~\new_[28073]_ ;
  assign \new_[27698]_  = ~\new_[29175]_  & ~\new_[30101]_ ;
  assign \new_[27699]_  = ~\new_[28930]_  | ~\new_[5986]_ ;
  assign \new_[27700]_  = ~\new_[28878]_  & ~\new_[29809]_ ;
  assign \new_[27701]_  = ~\new_[28903]_  | ~\new_[5923]_ ;
  assign \new_[27702]_  = ~\new_[28757]_ ;
  assign \new_[27703]_  = ~\new_[29167]_  & ~\new_[30140]_ ;
  assign \new_[27704]_  = \new_[29032]_  & \new_[5971]_ ;
  assign \new_[27705]_  = ~\new_[28199]_ ;
  assign \new_[27706]_  = ~\new_[28504]_ ;
  assign \new_[27707]_  = ~\new_[30183]_  & ~\new_[29445]_ ;
  assign \new_[27708]_  = (~\new_[30085]_  | ~\s2_data_i[3] ) & (~\new_[30108]_  | ~\s1_data_i[3] );
  assign \new_[27709]_  = ~\new_[28491]_ ;
  assign \new_[27710]_  = ~\new_[29332]_  & ~\new_[30250]_ ;
  assign \new_[27711]_  = ~\new_[29681]_  & ~\new_[30101]_ ;
  assign \new_[27712]_  = (~\new_[29948]_  | ~\s5_data_i[1] ) & (~\new_[29947]_  | ~\s3_data_i[1] );
  assign \new_[27713]_  = ~\new_[30591]_  | ~\new_[5928]_ ;
  assign \new_[27714]_  = ~\new_[29042]_  & ~\new_[30315]_ ;
  assign \new_[27715]_  = \new_[6050]_  & \new_[6049]_ ;
  assign \new_[27716]_  = (~\new_[30166]_  | ~\s14_data_i[19] ) & (~\new_[30298]_  | ~\s12_data_i[19] );
  assign \new_[27717]_  = ~\new_[30559]_  | ~\new_[28017]_ ;
  assign \new_[27718]_  = ~\new_[29576]_  | ~\new_[29984]_ ;
  assign \new_[27719]_  = (~\new_[29876]_  | ~\s11_data_i[28] ) & (~\new_[30341]_  | ~\s8_data_i[28] );
  assign \new_[27720]_  = ~\new_[29889]_  | ~\new_[30731]_ ;
  assign \new_[27721]_  = ~\new_[29089]_  & ~\new_[29865]_ ;
  assign \new_[27722]_  = ~\new_[30723]_  | ~\new_[30544]_ ;
  assign \new_[27723]_  = \new_[29061]_  & \new_[5993]_ ;
  assign \new_[27724]_  = ~\new_[29079]_  | ~\new_[30214]_ ;
  assign \new_[27725]_  = ~\new_[29639]_  & ~\new_[29994]_ ;
  assign \new_[27726]_  = ~\new_[28099]_ ;
  assign \new_[27727]_  = ~\new_[29944]_  & ~\new_[29652]_ ;
  assign \new_[27728]_  = ~\new_[30595]_  | ~\new_[30554]_ ;
  assign \new_[27729]_  = ~\new_[28328]_ ;
  assign \new_[27730]_  = ~\new_[30617]_  | ~\new_[29750]_ ;
  assign \new_[27731]_  = ~\new_[29606]_  | ~\new_[28964]_ ;
  assign \new_[27732]_  = (~\new_[30085]_  | ~\s2_data_i[11] ) & (~\new_[30108]_  | ~\s1_data_i[11] );
  assign \new_[27733]_  = ~\new_[28704]_ ;
  assign \new_[27734]_  = ~\new_[28154]_ ;
  assign \new_[27735]_  = ~\new_[28582]_ ;
  assign \new_[27736]_  = ~\new_[28685]_  & ~\new_[29950]_ ;
  assign \new_[27737]_  = ~\new_[28472]_ ;
  assign \new_[27738]_  = ~\new_[28581]_ ;
  assign \new_[27739]_  = \new_[30415]_  | \new_[29100]_ ;
  assign \new_[27740]_  = ~\new_[28406]_ ;
  assign \new_[27741]_  = ~\new_[28251]_ ;
  assign \new_[27742]_  = ~\new_[30568]_  | ~\new_[6057]_ ;
  assign \new_[27743]_  = ~\new_[30140]_  & ~\new_[29268]_ ;
  assign \new_[27744]_  = \new_[29171]_  & \new_[5981]_ ;
  assign \new_[27745]_  = ~\new_[29104]_  | ~\new_[29062]_ ;
  assign \new_[27746]_  = ~\new_[29202]_  | ~\new_[30176]_ ;
  assign \new_[27747]_  = (~\new_[29963]_  | ~\s4_data_i[5] ) & (~\new_[30481]_  | ~\s0_data_i[5] );
  assign \new_[27748]_  = ~\new_[29089]_  | ~\new_[29904]_ ;
  assign \new_[27749]_  = \new_[29038]_  & \new_[5998]_ ;
  assign \new_[27750]_  = ~\new_[29550]_  | ~\new_[29874]_ ;
  assign \new_[27751]_  = ~\new_[28556]_ ;
  assign \new_[27752]_  = ~\new_[28336]_ ;
  assign \new_[27753]_  = ~\new_[28866]_  | ~\new_[30067]_ ;
  assign \new_[27754]_  = ~\new_[30201]_  & ~\new_[30559]_ ;
  assign \new_[27755]_  = (~\new_[30013]_  | ~\s2_data_i[9] ) & (~\new_[29769]_  | ~\s1_data_i[9] );
  assign \new_[27756]_  = \new_[29401]_  & \new_[5972]_ ;
  assign \new_[27757]_  = ~\new_[29271]_  | ~\new_[5980]_ ;
  assign \new_[27758]_  = ~\new_[30415]_  | ~\new_[29320]_ ;
  assign \new_[27759]_  = ~\new_[28755]_ ;
  assign \new_[27760]_  = ~\new_[29472]_  | ~m4_stb_i;
  assign \new_[27761]_  = ~\new_[29550]_  | ~\new_[5963]_ ;
  assign \new_[27762]_  = ~\new_[28962]_  | ~\new_[28979]_ ;
  assign \new_[27763]_  = (~\new_[29807]_  | ~\s14_data_i[26] ) & (~\new_[30626]_  | ~\s12_data_i[26] );
  assign \new_[27764]_  = ~\new_[28588]_ ;
  assign \new_[27765]_  = ~\new_[29944]_  & ~\new_[30363]_ ;
  assign \new_[27766]_  = ~\new_[30375]_  & ~\new_[30670]_ ;
  assign \new_[27767]_  = ~\new_[29374]_  & ~\new_[5923]_ ;
  assign \new_[27768]_  = (~\new_[29961]_  | ~\s4_data_i[21] ) & (~\new_[29819]_  | ~\s0_data_i[21] );
  assign \new_[27769]_  = ~\new_[29370]_  & ~\new_[29545]_ ;
  assign \new_[27770]_  = (~\new_[30013]_  | ~\s2_data_i[6] ) & (~\new_[29769]_  | ~\s1_data_i[6] );
  assign \new_[27771]_  = ~\new_[29355]_  | ~\new_[5919]_ ;
  assign \new_[27772]_  = ~\new_[30693]_  | ~\new_[30291]_ ;
  assign \new_[27773]_  = ~\new_[28866]_  & ~\new_[29501]_ ;
  assign \new_[27774]_  = ~\new_[29466]_  | ~\new_[30207]_ ;
  assign \new_[27775]_  = ~\new_[29466]_  | ~\new_[30434]_ ;
  assign \new_[27776]_  = ~\new_[28374]_ ;
  assign \new_[27777]_  = ~\new_[29718]_  & ~\new_[31724]_ ;
  assign \new_[27778]_  = ~\new_[28535]_ ;
  assign \new_[27779]_  = (~\new_[29807]_  | ~\s14_data_i[22] ) & (~\new_[30626]_  | ~\s12_data_i[22] );
  assign \new_[27780]_  = ~\new_[28173]_ ;
  assign \new_[27781]_  = ~\new_[28171]_ ;
  assign \new_[27782]_  = ~\new_[28381]_ ;
  assign \new_[27783]_  = ~\new_[29996]_  | ~\new_[30735]_ ;
  assign \new_[27784]_  = ~\new_[28156]_ ;
  assign \new_[27785]_  = (~\new_[29788]_  | ~\s2_data_i[26] ) & (~\new_[30357]_  | ~\s1_data_i[26] );
  assign \new_[27786]_  = (~\new_[29823]_  | ~\s7_data_i[30] ) & (~\new_[29954]_  | ~\s6_data_i[30] );
  assign \new_[27787]_  = ~\new_[29019]_ ;
  assign \new_[27788]_  = ~\new_[28117]_ ;
  assign \new_[27789]_  = (~\new_[29823]_  | ~\s7_data_i[8] ) & (~\new_[29954]_  | ~\s6_data_i[8] );
  assign \new_[27790]_  = (~\new_[29961]_  | ~\s4_data_i[13] ) & (~\new_[29819]_  | ~\s0_data_i[13] );
  assign \new_[27791]_  = ~\new_[28361]_ ;
  assign \new_[27792]_  = ~\new_[28941]_  & ~\new_[6209]_ ;
  assign \new_[27793]_  = (~\new_[29846]_  | ~\s2_data_i[11] ) & (~\new_[30001]_  | ~\s1_data_i[11] );
  assign \new_[27794]_  = ~\new_[29717]_  | ~\new_[6078]_ ;
  assign \new_[27795]_  = ~\new_[29096]_  | ~\new_[29744]_ ;
  assign \new_[27796]_  = ~\new_[28084]_ ;
  assign \new_[27797]_  = ~\new_[28064]_ ;
  assign \new_[27798]_  = ~\new_[29739]_  & ~\new_[31421]_ ;
  assign \new_[27799]_  = ~\new_[28034]_ ;
  assign \new_[27800]_  = (~\new_[29846]_  | ~\s2_data_i[27] ) & (~\new_[30001]_  | ~\s1_data_i[27] );
  assign \new_[27801]_  = ~\new_[29941]_  & ~\new_[29174]_ ;
  assign \new_[27802]_  = ~\new_[28873]_ ;
  assign \new_[27803]_  = (~\new_[29807]_  | ~\s14_data_i[20] ) & (~\new_[30626]_  | ~\s12_data_i[20] );
  assign \new_[27804]_  = ~\new_[27999]_ ;
  assign \new_[27805]_  = ~\new_[29235]_  | ~\new_[30257]_ ;
  assign \new_[27806]_  = ~\new_[27977]_ ;
  assign \new_[27807]_  = ~\new_[30552]_  | ~\new_[5916]_ ;
  assign \new_[27808]_  = ~\new_[29003]_  | ~\new_[5965]_ ;
  assign \new_[27809]_  = ~\new_[28628]_ ;
  assign \new_[27810]_  = (~\new_[29961]_  | ~\s4_data_i[5] ) & (~\new_[29819]_  | ~\s0_data_i[5] );
  assign \new_[27811]_  = ~\new_[28334]_ ;
  assign \new_[27812]_  = (~\new_[30013]_  | ~\s2_data_i[12] ) & (~\new_[29769]_  | ~\s1_data_i[12] );
  assign \new_[27813]_  = ~\new_[28662]_ ;
  assign \new_[27814]_  = ~\new_[29575]_  & ~\new_[30884]_ ;
  assign \new_[27815]_  = (~\new_[30113]_  | ~\s2_data_i[4] ) & (~\new_[30124]_  | ~\s1_data_i[4] );
  assign \new_[27816]_  = ~\new_[29645]_  & ~\new_[31665]_ ;
  assign \new_[27817]_  = ~\new_[28639]_ ;
  assign \new_[27818]_  = ~\new_[30425]_  & ~\new_[29159]_ ;
  assign \new_[27819]_  = ~\new_[29099]_  & ~\new_[5927]_ ;
  assign \new_[27820]_  = (~\new_[29807]_  | ~\s14_data_i[21] ) & (~\new_[30626]_  | ~\s12_data_i[21] );
  assign \new_[27821]_  = ~\new_[30222]_  & ~\new_[29306]_ ;
  assign \new_[27822]_  = (~\new_[29949]_  | ~\s10_data_i[11] ) & (~\new_[29905]_  | ~\s9_data_i[11] );
  assign \new_[27823]_  = ~\new_[28907]_  | ~\new_[5909]_ ;
  assign \new_[27824]_  = ~\new_[29003]_  | ~\new_[30215]_ ;
  assign \new_[27825]_  = (~\new_[30131]_  | ~\s7_data_i[10] ) & (~\new_[29939]_  | ~\s6_data_i[10] );
  assign \new_[27826]_  = ~\new_[30268]_ ;
  assign \new_[27827]_  = \new_[29380]_  & \new_[30444]_ ;
  assign \new_[27828]_  = ~\new_[28653]_ ;
  assign \new_[27829]_  = ~\new_[28919]_  | ~\new_[5921]_ ;
  assign \new_[27830]_  = ~\new_[28143]_ ;
  assign \new_[27831]_  = ~\new_[28771]_ ;
  assign \new_[27832]_  = ~\new_[28656]_ ;
  assign \new_[27833]_  = ~\new_[28657]_ ;
  assign \new_[27834]_  = ~\new_[28364]_ ;
  assign \new_[27835]_  = ~\new_[30718]_  & ~\new_[29015]_ ;
  assign \new_[27836]_  = \new_[28989]_  & \new_[5969]_ ;
  assign \new_[27837]_  = ~\new_[28647]_ ;
  assign \new_[27838]_  = ~\new_[28814]_ ;
  assign \new_[27839]_  = ~\new_[28917]_  | ~\new_[5918]_ ;
  assign \new_[27840]_  = ~\new_[29755]_  | ~\new_[31406]_ ;
  assign \new_[27841]_  = ~\new_[28028]_ ;
  assign \new_[27842]_  = ~\new_[28670]_ ;
  assign \new_[27843]_  = ~\new_[28671]_ ;
  assign \new_[27844]_  = ~\new_[28151]_ ;
  assign \new_[27845]_  = ~\new_[29132]_  & ~\new_[29071]_ ;
  assign \new_[27846]_  = ~\new_[28568]_ ;
  assign \new_[27847]_  = ~\new_[28104]_ ;
  assign \new_[27848]_  = ~\new_[29165]_  & ~\new_[28891]_ ;
  assign \new_[27849]_  = ~\new_[28109]_ ;
  assign \new_[27850]_  = ~\new_[28071]_ ;
  assign \new_[27851]_  = ~\new_[28051]_ ;
  assign \new_[27852]_  = ~\new_[29742]_  & ~\new_[31712]_ ;
  assign \new_[27853]_  = ~\new_[28038]_ ;
  assign \new_[27854]_  = ~\new_[29593]_  | ~\new_[5976]_ ;
  assign \new_[27855]_  = \new_[28974]_  & \new_[31061]_ ;
  assign \new_[27856]_  = ~\new_[28689]_ ;
  assign \new_[27857]_  = ~\new_[28881]_  | ~\new_[5978]_ ;
  assign \new_[27858]_  = ~\new_[27996]_ ;
  assign \new_[27859]_  = (~\new_[29963]_  | ~\s4_data_i[28] ) & (~\new_[30481]_  | ~\s0_data_i[28] );
  assign \new_[27860]_  = ~\new_[28211]_  & ~\new_[28023]_ ;
  assign \new_[27861]_  = ~\new_[28972]_  | ~\new_[5926]_ ;
  assign \new_[27862]_  = ~\new_[27992]_ ;
  assign \new_[27863]_  = ~\new_[29389]_  | ~\new_[29406]_ ;
  assign \new_[27864]_  = ~\new_[28271]_ ;
  assign \new_[27865]_  = (~\new_[29876]_  | ~\s11_data_i[8] ) & (~\new_[30341]_  | ~\s8_data_i[8] );
  assign \new_[27866]_  = \new_[29738]_  | \new_[31614]_ ;
  assign \new_[27867]_  = ~\new_[28741]_ ;
  assign \new_[27868]_  = (~\new_[30113]_  | ~\s2_data_i[27] ) & (~\new_[30124]_  | ~\s1_data_i[27] );
  assign \new_[27869]_  = ~\new_[28224]_ ;
  assign \new_[27870]_  = ~\new_[28702]_ ;
  assign \new_[27871]_  = \new_[29427]_  | \new_[31045]_ ;
  assign \new_[27872]_  = (~\new_[30189]_  | ~\s2_data_i[27] ) & (~\new_[30195]_  | ~\s1_data_i[27] );
  assign \new_[27873]_  = ~\new_[28952]_  | ~\new_[31614]_ ;
  assign \new_[27874]_  = ~\new_[29546]_  | ~\new_[31045]_ ;
  assign \new_[27875]_  = ~\new_[28265]_ ;
  assign \new_[27876]_  = ~\new_[28862]_  & ~\new_[5909]_ ;
  assign \new_[27877]_  = ~\new_[28323]_ ;
  assign \new_[27878]_  = ~\new_[28247]_ ;
  assign \new_[27879]_  = \new_[28974]_  & \new_[31105]_ ;
  assign \new_[27880]_  = (~\new_[29963]_  | ~\s4_data_i[22] ) & (~\new_[30481]_  | ~\s0_data_i[22] );
  assign \new_[27881]_  = ~\new_[28751]_ ;
  assign \new_[27882]_  = ~\new_[29471]_  & ~\new_[29306]_ ;
  assign \new_[27883]_  = ~\new_[28397]_ ;
  assign \new_[27884]_  = ~\new_[28617]_ ;
  assign \new_[27885]_  = ~\new_[28679]_ ;
  assign \new_[27886]_  = ~\new_[28112]_ ;
  assign \new_[27887]_  = ~\new_[28551]_ ;
  assign \new_[27888]_  = ~\new_[28288]_ ;
  assign \new_[27889]_  = ~\new_[28717]_ ;
  assign \new_[27890]_  = ~\new_[28987]_  | ~\new_[5911]_ ;
  assign \new_[27891]_  = ~\new_[28243]_ ;
  assign \new_[27892]_  = ~\new_[29197]_ ;
  assign \new_[27893]_  = ~\new_[28148]_ ;
  assign \new_[27894]_  = ~\new_[29738]_  & ~\new_[31438]_ ;
  assign \new_[27895]_  = ~\new_[28743]_ ;
  assign \new_[27896]_  = ~\new_[29306]_  & ~\new_[30750]_ ;
  assign \new_[27897]_  = ~\new_[29656]_ ;
  assign \new_[27898]_  = ~\new_[28992]_  & ~\new_[29841]_ ;
  assign \new_[27899]_  = ~\new_[28343]_ ;
  assign \new_[27900]_  = ~\new_[28093]_ ;
  assign \new_[27901]_  = ~\new_[28725]_ ;
  assign \new_[27902]_  = \new_[28949]_  & \new_[5932]_ ;
  assign \new_[27903]_  = ~\new_[28055]_ ;
  assign \new_[27904]_  = ~\new_[29016]_  & ~\new_[29722]_ ;
  assign \new_[27905]_  = ~\new_[28550]_ ;
  assign \new_[27906]_  = ~\new_[28990]_  | ~\new_[5912]_ ;
  assign \new_[27907]_  = ~\new_[28238]_ ;
  assign \new_[27908]_  = ~\new_[28729]_ ;
  assign \new_[27909]_  = ~\new_[28731]_ ;
  assign \new_[27910]_  = ~\new_[28900]_  | ~\new_[6084]_ ;
  assign \new_[27911]_  = ~\new_[28549]_ ;
  assign \new_[27912]_  = (~\new_[29948]_  | ~\s5_data_i[13] ) & (~\new_[29947]_  | ~\s3_data_i[13] );
  assign \new_[27913]_  = ~\new_[28736]_ ;
  assign \new_[27914]_  = ~\new_[28580]_ ;
  assign \new_[27915]_  = ~\new_[29914]_ ;
  assign \new_[27916]_  = ~\new_[29726]_  | ~\new_[5926]_ ;
  assign \new_[27917]_  = ~\new_[28744]_ ;
  assign \new_[27918]_  = ~\new_[28492]_ ;
  assign \new_[27919]_  = ~\new_[28780]_ ;
  assign \new_[27920]_  = ~\new_[28775]_ ;
  assign \new_[27921]_  = ~\new_[28764]_ ;
  assign \new_[27922]_  = ~\new_[30521]_  | ~\new_[6092]_ ;
  assign \new_[27923]_  = ~\new_[28856]_  & ~\new_[30125]_ ;
  assign \new_[27924]_  = ~\new_[28738]_ ;
  assign \new_[27925]_  = ~\new_[28885]_  | ~\new_[5909]_ ;
  assign \new_[27926]_  = ~\new_[28686]_  & ~\new_[29981]_ ;
  assign \new_[27927]_  = (~\new_[29807]_  | ~\s14_data_i[5] ) & (~\new_[30626]_  | ~\s12_data_i[5] );
  assign \new_[27928]_  = ~\new_[28941]_  & ~\new_[31772]_ ;
  assign \new_[27929]_  = ~\new_[28242]_ ;
  assign \new_[27930]_  = ~\new_[28759]_ ;
  assign \new_[27931]_  = ~\new_[29720]_  | ~\new_[5927]_ ;
  assign \new_[27932]_  = ~\new_[28320]_ ;
  assign \new_[27933]_  = ~\new_[29067]_  & ~\new_[5911]_ ;
  assign \new_[27934]_  = ~\new_[28763]_ ;
  assign \new_[27935]_  = ~\new_[28332]_ ;
  assign \new_[27936]_  = (~\new_[30013]_  | ~\s2_data_i[18] ) & (~\new_[29769]_  | ~\s1_data_i[18] );
  assign \new_[27937]_  = ~\new_[28772]_ ;
  assign \new_[27938]_  = ~\new_[28629]_ ;
  assign \new_[27939]_  = ~\new_[29753]_  & ~\new_[6078]_ ;
  assign \new_[27940]_  = ~\new_[28958]_  | ~\new_[5911]_ ;
  assign \new_[27941]_  = ~\new_[28680]_ ;
  assign \new_[27942]_  = ~\new_[29908]_ ;
  assign \new_[27943]_  = ~\new_[28779]_ ;
  assign \new_[27944]_  = ~\new_[29527]_  | ~\new_[6036]_ ;
  assign \new_[27945]_  = ~\new_[28068]_ ;
  assign \new_[27946]_  = \new_[29971]_  & \new_[30011]_ ;
  assign \new_[27947]_  = (~\new_[29788]_  | ~\s2_data_i[6] ) & (~\new_[30357]_  | ~\s1_data_i[6] );
  assign \new_[27948]_  = (~\new_[29846]_  | ~\s2_data_i[2] ) & (~\new_[30001]_  | ~\s1_data_i[2] );
  assign \new_[27949]_  = ~\new_[29262]_  | ~\new_[5978]_ ;
  assign \new_[27950]_  = ~\new_[29445]_  | ~\new_[29441]_ ;
  assign \new_[27951]_  = ~\new_[29300]_  | ~\new_[28905]_ ;
  assign \new_[27952]_  = ~\new_[28799]_ ;
  assign \new_[27953]_  = ~\new_[28794]_ ;
  assign \new_[27954]_  = ~\new_[30652]_  & ~\new_[29701]_ ;
  assign \new_[27955]_  = (~\new_[29963]_  | ~\s4_data_i[30] ) & (~\new_[30481]_  | ~\s0_data_i[30] );
  assign \new_[27956]_  = ~\new_[28769]_ ;
  assign \new_[27957]_  = ~\new_[29724]_  & ~\new_[31176]_ ;
  assign \new_[27958]_  = ~\new_[30222]_  | ~\new_[30550]_ ;
  assign \new_[27959]_  = \new_[29767]_  & \new_[28887]_ ;
  assign \new_[27960]_  = ~\new_[29810]_  & ~\new_[30650]_ ;
  assign \new_[27961]_  = ~\new_[28802]_ ;
  assign \new_[27962]_  = ~\new_[30415]_  & ~\new_[28872]_ ;
  assign \new_[27963]_  = (~\new_[30013]_  | ~\s2_data_i[19] ) & (~\new_[29769]_  | ~\s1_data_i[19] );
  assign \new_[27964]_  = ~\new_[28950]_  | ~\new_[30363]_ ;
  assign \new_[27965]_  = ~\new_[28798]_ ;
  assign \new_[27966]_  = ~\new_[28898]_  | ~\new_[6087]_ ;
  assign \new_[27967]_  = ~\new_[28810]_ ;
  assign \new_[27968]_  = (~\new_[30113]_  | ~\s2_data_i[10] ) & (~\new_[30124]_  | ~\s1_data_i[10] );
  assign \new_[27969]_  = (~\new_[30166]_  | ~\s14_data_i[21] ) & (~\new_[30298]_  | ~\s12_data_i[21] );
  assign \new_[27970]_  = (~\new_[29963]_  | ~\s4_data_i[23] ) & (~\new_[30481]_  | ~\s0_data_i[23] );
  assign \new_[27971]_  = ~\new_[29650]_  & ~\new_[30574]_ ;
  assign \new_[27972]_  = ~\new_[28299]_ ;
  assign \new_[27973]_  = ~\new_[29123]_ ;
  assign \new_[27974]_  = ~\new_[28983]_ ;
  assign \new_[27975]_  = ~\new_[29000]_ ;
  assign \new_[27976]_  = ~\new_[30701]_  & ~\new_[30293]_ ;
  assign \new_[27977]_  = ~\new_[30395]_  | ~\new_[31148]_ ;
  assign \new_[27978]_  = ~\new_[30168]_  & ~\new_[29983]_ ;
  assign \new_[27979]_  = ~\new_[29481]_ ;
  assign \new_[27980]_  = ~\new_[29620]_ ;
  assign \new_[27981]_  = \new_[29796]_  & \new_[6059]_ ;
  assign \new_[27982]_  = ~\new_[30629]_  | ~\new_[5967]_ ;
  assign \new_[27983]_  = ~\new_[32161]_  | ~m3_stb_i;
  assign \new_[27984]_  = ~\new_[28832]_ ;
  assign \new_[27985]_  = \new_[30050]_  & \new_[30869]_ ;
  assign \new_[27986]_  = \new_[29978]_  & \new_[5987]_ ;
  assign \new_[27987]_  = \new_[30164]_  & \new_[5963]_ ;
  assign \new_[27988]_  = ~\new_[30359]_  | ~\new_[31411]_ ;
  assign \new_[27989]_  = ~\new_[30391]_  & ~\new_[31870]_ ;
  assign \new_[27990]_  = ~\new_[30568]_  | ~\new_[30717]_ ;
  assign \new_[27991]_  = ~\new_[29892]_  & ~\new_[30291]_ ;
  assign \new_[27992]_  = ~\new_[30353]_  & ~\new_[5923]_ ;
  assign \new_[27993]_  = ~\new_[28867]_  & ~\new_[30544]_ ;
  assign \new_[27994]_  = ~\new_[30348]_  & ~\new_[30647]_ ;
  assign \new_[27995]_  = ~\new_[29616]_ ;
  assign \new_[27996]_  = ~\new_[30137]_  & ~\new_[31416]_ ;
  assign \new_[27997]_  = ~\new_[29613]_ ;
  assign \new_[27998]_  = ~\new_[29292]_ ;
  assign \new_[27999]_  = ~\new_[30414]_  & ~\new_[6190]_ ;
  assign \new_[28000]_  = ~\new_[30612]_  | ~\new_[30152]_ ;
  assign \new_[28001]_  = ~\new_[29611]_ ;
  assign \new_[28002]_  = ~\new_[29884]_  & ~\new_[31645]_ ;
  assign \new_[28003]_  = ~\new_[29612]_ ;
  assign \new_[28004]_  = ~\new_[30030]_ ;
  assign \new_[28005]_  = ~\new_[29283]_ ;
  assign \new_[28006]_  = ~\new_[30382]_  | ~\new_[31648]_ ;
  assign \new_[28007]_  = ~\new_[29277]_ ;
  assign \new_[28008]_  = ~\new_[29844]_  & ~\new_[5979]_ ;
  assign \new_[28009]_  = ~\new_[31815]_  & ~\new_[31906]_ ;
  assign \new_[28010]_  = \new_[30324]_  & \new_[5964]_ ;
  assign \new_[28011]_  = ~\new_[6093]_  & ~\new_[31776]_ ;
  assign \new_[28012]_  = ~\new_[28865]_ ;
  assign \new_[28013]_  = ~\new_[29374]_ ;
  assign \new_[28014]_  = ~\new_[30391]_  & ~\new_[31235]_ ;
  assign \new_[28015]_  = ~\new_[29137]_ ;
  assign \new_[28016]_  = ~\new_[30325]_  & ~\new_[30271]_ ;
  assign \new_[28017]_  = ~\new_[30444]_ ;
  assign \new_[28018]_  = ~\new_[30383]_  | ~\new_[31014]_ ;
  assign \new_[28019]_  = ~\new_[28970]_ ;
  assign \new_[28020]_  = ~\new_[28877]_ ;
  assign \new_[28021]_  = ~\new_[28840]_ ;
  assign \new_[28022]_  = ~\new_[29766]_  | ~\new_[31235]_ ;
  assign \new_[28023]_  = ~\new_[30129]_ ;
  assign \new_[28024]_  = ~\new_[29836]_  | ~\new_[31433]_ ;
  assign \new_[28025]_  = ~\new_[30137]_  & ~\new_[6001]_ ;
  assign \new_[28026]_  = ~\new_[30017]_  | ~\new_[31442]_ ;
  assign \new_[28027]_  = ~\new_[28878]_ ;
  assign \new_[28028]_  = ~\new_[29811]_  | ~\new_[31165]_ ;
  assign \new_[28029]_  = ~\new_[28889]_ ;
  assign \new_[28030]_  = ~\new_[30689]_  & ~\new_[5991]_ ;
  assign \new_[28031]_  = ~\new_[30363]_ ;
  assign \new_[28032]_  = ~\new_[30377]_  | ~\new_[6078]_ ;
  assign \new_[28033]_  = ~\new_[28897]_ ;
  assign \new_[28034]_  = ~\new_[29998]_  & ~\new_[6176]_ ;
  assign \new_[28035]_  = ~\new_[28901]_ ;
  assign \new_[28036]_  = ~\new_[28910]_ ;
  assign \new_[28037]_  = ~\new_[29901]_  | ~\new_[31230]_ ;
  assign \new_[28038]_  = \new_[29896]_  | \new_[6038]_ ;
  assign \new_[28039]_  = ~\new_[30235]_ ;
  assign \new_[28040]_  = \new_[30338]_  & \new_[5985]_ ;
  assign \new_[28041]_  = ~\new_[28920]_ ;
  assign \new_[28042]_  = \new_[29938]_  & \new_[6246]_ ;
  assign \new_[28043]_  = ~\new_[29901]_  | ~\new_[6066]_ ;
  assign \new_[28044]_  = ~\new_[30380]_  | ~\new_[31403]_ ;
  assign \new_[28045]_  = ~\new_[29853]_ ;
  assign \new_[28046]_  = ~\new_[29896]_  & ~\new_[31665]_ ;
  assign \new_[28047]_  = ~\new_[29200]_ ;
  assign \new_[28048]_  = ~\new_[30005]_  | ~\new_[29865]_ ;
  assign \new_[28049]_  = ~\new_[30042]_  | ~\new_[29900]_ ;
  assign \new_[28050]_  = ~\new_[30327]_ ;
  assign \new_[28051]_  = ~\new_[29797]_  & ~\new_[6038]_ ;
  assign \new_[28052]_  = ~\new_[28935]_ ;
  assign \new_[28053]_  = ~\new_[28932]_ ;
  assign \new_[28054]_  = ~\new_[29865]_ ;
  assign \new_[28055]_  = ~\new_[29920]_  | ~\new_[30976]_ ;
  assign \new_[28056]_  = ~\new_[29170]_ ;
  assign \new_[28057]_  = ~\new_[28944]_ ;
  assign \new_[28058]_  = ~\new_[30396]_  & ~\new_[30998]_ ;
  assign \new_[28059]_  = ~\new_[29661]_ ;
  assign \new_[28060]_  = \new_[29957]_  | \new_[5923]_ ;
  assign \new_[28061]_  = ~\new_[29477]_ ;
  assign \new_[28062]_  = ~\new_[29362]_ ;
  assign \new_[28063]_  = ~\new_[29160]_ ;
  assign \new_[28064]_  = ~\new_[30065]_  & ~\new_[5964]_ ;
  assign \new_[28065]_  = ~\new_[30248]_  | ~\new_[30732]_ ;
  assign \new_[28066]_  = ~\new_[30112]_  | ~\new_[31855]_ ;
  assign \new_[28067]_  = ~\new_[30021]_ ;
  assign \new_[28068]_  = ~\new_[29829]_  | ~\new_[31464]_ ;
  assign \new_[28069]_  = ~\new_[29880]_ ;
  assign \new_[28070]_  = ~\new_[30389]_ ;
  assign \new_[28071]_  = \new_[29818]_  & \new_[6059]_ ;
  assign \new_[28072]_  = ~\new_[30201]_  | ~\new_[30367]_ ;
  assign \new_[28073]_  = ~\new_[30101]_ ;
  assign \new_[28074]_  = ~\new_[29861]_  | ~\new_[30150]_ ;
  assign \new_[28075]_  = ~\new_[30387]_  | ~\new_[6209]_ ;
  assign \new_[28076]_  = ~\new_[29785]_ ;
  assign \new_[28077]_  = ~\new_[30430]_  & ~\new_[5931]_ ;
  assign \new_[28078]_  = ~\new_[30508]_ ;
  assign \new_[28079]_  = ~\new_[30079]_  | ~\new_[5896]_ ;
  assign \new_[28080]_  = ~\new_[30429]_  | ~\new_[31047]_  | ~m6_cyc_i;
  assign \new_[28081]_  = ~\new_[30126]_  & ~\new_[30315]_ ;
  assign \new_[28082]_  = ~\new_[30379]_  & ~\new_[30969]_ ;
  assign \new_[28083]_  = ~\new_[30507]_ ;
  assign \new_[28084]_  = ~\new_[29875]_  | ~\new_[31648]_ ;
  assign \new_[28085]_  = ~\new_[30049]_  | ~\new_[5926]_ ;
  assign \new_[28086]_  = ~\new_[30126]_  | ~\new_[29946]_ ;
  assign \new_[28087]_  = \new_[30012]_  | \new_[5926]_ ;
  assign \new_[28088]_  = ~\new_[28980]_ ;
  assign \new_[28089]_  = ~\new_[30125]_ ;
  assign \new_[28090]_  = ~\new_[30386]_  | ~\new_[6044]_ ;
  assign \new_[28091]_  = ~\new_[30206]_  | ~\new_[29977]_ ;
  assign \new_[28092]_  = ~\new_[30233]_  & ~\new_[30018]_ ;
  assign \new_[28093]_  = \new_[29842]_  & \new_[5913]_ ;
  assign \new_[28094]_  = ~\new_[29894]_  | ~\new_[6094]_ ;
  assign \new_[28095]_  = \new_[29866]_  | \new_[31438]_ ;
  assign \new_[28096]_  = (~\new_[6083]_  | ~\new_[30489]_ ) & (~\new_[6186]_  | ~\new_[31094]_ );
  assign \new_[28097]_  = ~\new_[30375]_  | ~\new_[30647]_ ;
  assign \new_[28098]_  = ~\new_[30202]_  & ~\new_[30057]_ ;
  assign \new_[28099]_  = ~\new_[30276]_  & ~\new_[30764]_ ;
  assign \new_[28100]_  = ~\new_[29778]_  & ~\new_[6210]_ ;
  assign \new_[28101]_  = ~\new_[29552]_ ;
  assign \new_[28102]_  = ~\new_[28994]_ ;
  assign \new_[28103]_  = ~\new_[30788]_  & ~\new_[30210]_ ;
  assign \new_[28104]_  = ~\new_[29822]_  | ~\new_[31455]_ ;
  assign \new_[28105]_  = ~\new_[29715]_ ;
  assign \new_[28106]_  = ~\new_[30356]_  & ~\new_[5921]_ ;
  assign \new_[28107]_  = ~\new_[30469]_  | ~\new_[31162]_  | ~m1_cyc_i;
  assign \new_[28108]_  = ~\new_[30024]_  | ~\new_[30159]_ ;
  assign \new_[28109]_  = ~\new_[29845]_  & ~\new_[5918]_ ;
  assign \new_[28110]_  = ~\new_[29256]_ ;
  assign \new_[28111]_  = ~\new_[30028]_  & ~\new_[29553]_ ;
  assign \new_[28112]_  = ~\new_[30378]_  & ~\new_[6269]_ ;
  assign \new_[28113]_  = \new_[29855]_  & \new_[30030]_ ;
  assign \new_[28114]_  = ~\new_[30332]_ ;
  assign \new_[28115]_  = ~\new_[30111]_  | ~\new_[30660]_ ;
  assign \new_[28116]_  = ~\new_[30328]_  | ~\new_[30246]_ ;
  assign \new_[28117]_  = ~\new_[30313]_  & ~\new_[5924]_ ;
  assign \new_[28118]_  = ~\new_[30025]_  & ~\new_[29789]_ ;
  assign \new_[28119]_  = ~\new_[29662]_ ;
  assign \new_[28120]_  = ~\new_[30266]_  & ~\new_[29977]_ ;
  assign \new_[28121]_  = ~\new_[29965]_ ;
  assign \new_[28122]_  = ~\new_[30071]_  | ~\new_[30581]_ ;
  assign \new_[28123]_  = ~\new_[29784]_  & ~\new_[31669]_ ;
  assign \new_[28124]_  = ~\new_[30226]_  | ~\new_[31479]_ ;
  assign \new_[28125]_  = ~\new_[29039]_ ;
  assign \new_[28126]_  = ~\new_[29945]_  & ~\new_[5913]_ ;
  assign \new_[28127]_  = ~\new_[30540]_  | ~\new_[30152]_ ;
  assign \new_[28128]_  = ~\new_[30521]_  | ~\new_[29798]_ ;
  assign \new_[28129]_  = ~\new_[29046]_ ;
  assign \new_[28130]_  = ~\new_[30000]_  | ~\new_[30750]_ ;
  assign \new_[28131]_  = ~\new_[29535]_ ;
  assign \new_[28132]_  = ~\new_[29053]_ ;
  assign \new_[28133]_  = ~\new_[29051]_ ;
  assign \new_[28134]_  = ~\new_[29450]_ ;
  assign \new_[28135]_  = ~\new_[29851]_  & ~\new_[29964]_ ;
  assign \new_[28136]_  = ~\new_[30871]_  & ~\new_[30954]_ ;
  assign \new_[28137]_  = ~\new_[29899]_  | ~\new_[30172]_ ;
  assign \new_[28138]_  = ~\new_[29929]_  | ~\new_[31423]_ ;
  assign \new_[28139]_  = ~\new_[29979]_  | ~\new_[29989]_ ;
  assign \new_[28140]_  = ~\new_[29378]_ ;
  assign \new_[28141]_  = ~\new_[29570]_ ;
  assign \new_[28142]_  = ~\new_[29372]_ ;
  assign \new_[28143]_  = ~\new_[29824]_  & ~\new_[5917]_ ;
  assign \new_[28144]_  = ~\new_[29828]_  | ~\new_[30434]_ ;
  assign \new_[28145]_  = ~\new_[29379]_ ;
  assign \new_[28146]_  = ~\new_[29059]_ ;
  assign \new_[28147]_  = ~\new_[30202]_  & ~\new_[31569]_ ;
  assign \new_[28148]_  = ~\new_[29860]_  & ~\new_[5927]_ ;
  assign \new_[28149]_  = ~\new_[29067]_ ;
  assign \new_[28150]_  = ~\new_[30711]_  | ~\new_[30011]_ ;
  assign \new_[28151]_  = ~\new_[29835]_  & ~\new_[5911]_ ;
  assign \new_[28152]_  = ~\new_[30042]_ ;
  assign \new_[28153]_  = ~\new_[29974]_  | ~\new_[5988]_ ;
  assign \new_[28154]_  = ~\new_[30089]_  | ~\new_[30591]_ ;
  assign \new_[28155]_  = ~\new_[29073]_ ;
  assign \new_[28156]_  = ~\new_[29921]_  & ~\new_[5981]_ ;
  assign \new_[28157]_  = ~\new_[29076]_ ;
  assign \new_[28158]_  = ~\new_[29917]_  & ~\new_[31235]_ ;
  assign \new_[28159]_  = ~\new_[29257]_ ;
  assign \new_[28160]_  = ~\new_[30410]_  | ~\new_[6206]_ ;
  assign \new_[28161]_  = \new_[30383]_  & \new_[5979]_ ;
  assign \new_[28162]_  = ~\new_[30221]_  & ~\new_[30332]_ ;
  assign \new_[28163]_  = ~\new_[29049]_ ;
  assign \new_[28164]_  = ~\new_[30349]_  | ~\new_[30568]_ ;
  assign \new_[28165]_  = ~\new_[29085]_ ;
  assign \new_[28166]_  = ~\new_[29086]_ ;
  assign \new_[28167]_  = ~\new_[30160]_  | ~\new_[30649]_ ;
  assign \new_[28168]_  = ~\new_[29091]_ ;
  assign \new_[28169]_  = ~\new_[30244]_  & ~\new_[30205]_ ;
  assign \new_[28170]_  = ~\new_[29090]_ ;
  assign \new_[28171]_  = ~\new_[29472]_ ;
  assign \new_[28172]_  = ~\new_[29836]_  | ~\new_[6096]_ ;
  assign \new_[28173]_  = ~\new_[30384]_  | ~\new_[30897]_ ;
  assign \new_[28174]_  = ~\new_[29813]_  | ~\new_[6079]_ ;
  assign \new_[28175]_  = ~\new_[29879]_  | ~\new_[5978]_ ;
  assign \new_[28176]_  = ~\new_[30275]_  | ~\new_[30775]_ ;
  assign \new_[28177]_  = ~\new_[29881]_  | ~\new_[5921]_ ;
  assign \new_[28178]_  = ~\new_[30581]_  | ~\new_[30572]_ ;
  assign \new_[28179]_  = ~\new_[29694]_ ;
  assign \new_[28180]_  = ~\new_[30168]_  & ~\new_[31844]_ ;
  assign \new_[28181]_  = ~\new_[30268]_  | ~\new_[29762]_ ;
  assign \new_[28182]_  = ~\new_[29839]_  | ~\new_[30097]_ ;
  assign \new_[28183]_  = ~\new_[29055]_ ;
  assign \new_[28184]_  = ~\new_[30102]_  | ~\new_[5911]_ ;
  assign \new_[28185]_  = ~\new_[30213]_  | ~\new_[6061]_ ;
  assign \new_[28186]_  = ~\new_[30381]_  | ~\new_[30141]_ ;
  assign \new_[28187]_  = ~\new_[30329]_  | ~\new_[6065]_ ;
  assign \new_[28188]_  = ~\new_[29113]_ ;
  assign \new_[28189]_  = ~\new_[30041]_  | ~\new_[6040]_ ;
  assign \new_[28190]_  = ~\new_[29188]_ ;
  assign \new_[28191]_  = ~\new_[30025]_ ;
  assign \new_[28192]_  = \new_[29829]_  & \new_[6176]_ ;
  assign \new_[28193]_  = ~\new_[29873]_  | ~\new_[30231]_ ;
  assign \new_[28194]_  = ~\new_[29772]_ ;
  assign \new_[28195]_  = ~\new_[29121]_ ;
  assign \new_[28196]_  = \new_[30651]_  | \new_[30213]_ ;
  assign \new_[28197]_  = ~\new_[29099]_ ;
  assign \new_[28198]_  = ~\new_[30202]_  | ~\new_[5897]_ ;
  assign \new_[28199]_  = ~\new_[29997]_  & ~\new_[30295]_ ;
  assign \new_[28200]_  = ~\new_[30791]_  & ~\new_[31132]_ ;
  assign \new_[28201]_  = ~\new_[29906]_  & ~\new_[31724]_ ;
  assign \new_[28202]_  = \new_[29811]_  & \new_[6206]_ ;
  assign \new_[28203]_  = ~\new_[29134]_ ;
  assign \new_[28204]_  = ~\new_[29324]_ ;
  assign \new_[28205]_  = ~\new_[29204]_ ;
  assign \new_[28206]_  = ~\new_[29138]_ ;
  assign \new_[28207]_  = ~\new_[29972]_  | ~\new_[6269]_ ;
  assign \new_[28208]_  = \new_[30034]_  & \new_[6190]_ ;
  assign \new_[28209]_  = ~\new_[29895]_  & ~\new_[5911]_ ;
  assign \new_[28210]_  = ~\new_[30336]_  | ~\new_[30573]_ ;
  assign \new_[28211]_  = ~\new_[30034]_ ;
  assign \new_[28212]_  = ~\new_[29143]_ ;
  assign \new_[28213]_  = (~\new_[5898]_  | ~\new_[30587]_ ) & (~\new_[6050]_  | ~\new_[31212]_ );
  assign \new_[28214]_  = (~\new_[5923]_  | ~\new_[30704]_ ) & (~\new_[5996]_  | ~\new_[31339]_ );
  assign \new_[28215]_  = ~\new_[29238]_ ;
  assign \new_[28216]_  = ~\new_[30059]_  & ~\new_[30316]_ ;
  assign \new_[28217]_  = ~\new_[30294]_  & ~\new_[30250]_ ;
  assign \new_[28218]_  = ~\new_[29926]_  | ~\new_[30721]_ ;
  assign \new_[28219]_  = (~\new_[30625]_  | ~\new_[5897]_ ) & (~\new_[31211]_  | ~\new_[5971]_ );
  assign \new_[28220]_  = ~\new_[30240]_  & ~\new_[31837]_ ;
  assign \new_[28221]_  = ~\new_[30350]_  & ~\new_[30814]_ ;
  assign \new_[28222]_  = ~\new_[29908]_  | ~\new_[30320]_ ;
  assign \new_[28223]_  = \new_[29804]_  & \new_[31135]_ ;
  assign \new_[28224]_  = ~\new_[30362]_  & ~\new_[31140]_ ;
  assign \new_[28225]_  = ~\new_[30282]_  | ~\new_[5912]_ ;
  assign \new_[28226]_  = ~\new_[30370]_  | ~\new_[31648]_ ;
  assign \new_[28227]_  = ~\new_[30018]_  & ~\new_[30820]_ ;
  assign \new_[28228]_  = ~\new_[29924]_  & ~\new_[29841]_ ;
  assign \new_[28229]_  = ~\new_[30724]_  & ~\new_[29956]_ ;
  assign \new_[28230]_  = ~\new_[29813]_  | ~\new_[30620]_ ;
  assign \new_[28231]_  = ~\new_[29889]_  | ~\new_[30695]_ ;
  assign \new_[28232]_  = ~\new_[29186]_ ;
  assign \new_[28233]_  = ~\new_[29913]_  & ~\new_[30732]_ ;
  assign \new_[28234]_  = ~\new_[29589]_ ;
  assign \new_[28235]_  = (~\new_[6067]_  | ~\new_[30796]_ ) & (~\new_[6194]_  | ~\new_[30988]_ );
  assign \new_[28236]_  = ~\new_[29563]_ ;
  assign \new_[28237]_  = ~\new_[30366]_  & ~\new_[5991]_ ;
  assign \new_[28238]_  = ~\new_[30737]_  & ~\new_[29972]_ ;
  assign \new_[28239]_  = ~\new_[29821]_  | ~\new_[5977]_ ;
  assign \new_[28240]_  = ~\new_[29883]_  & ~\new_[30507]_ ;
  assign \new_[28241]_  = ~\new_[29897]_  | ~\new_[30521]_ ;
  assign \new_[28242]_  = \new_[30382]_  & \new_[31390]_ ;
  assign \new_[28243]_  = ~\new_[30366]_  & ~\new_[31787]_ ;
  assign \new_[28244]_  = ~\new_[29689]_ ;
  assign \new_[28245]_  = ~\new_[30413]_ ;
  assign \new_[28246]_  = ~\new_[29844]_  & ~\new_[31014]_ ;
  assign \new_[28247]_  = ~\new_[29852]_  & ~\new_[31419]_ ;
  assign \new_[28248]_  = ~\new_[29060]_ ;
  assign \new_[28249]_  = ~\new_[29855]_ ;
  assign \new_[28250]_  = ~\new_[29029]_ ;
  assign \new_[28251]_  = ~\new_[29985]_  & ~\new_[30117]_ ;
  assign \new_[28252]_  = ~\new_[30373]_  | ~\new_[6040]_ ;
  assign \new_[28253]_  = ~\new_[29470]_ ;
  assign \new_[28254]_  = ~\new_[29001]_ ;
  assign \new_[28255]_  = ~\new_[29011]_ ;
  assign \new_[28256]_  = ~\new_[29861]_  | ~\new_[5894]_ ;
  assign \new_[28257]_  = ~\new_[30401]_  | ~\new_[6078]_ ;
  assign \new_[28258]_  = ~\new_[29423]_ ;
  assign \new_[28259]_  = ~\new_[30135]_  | ~\new_[29981]_ ;
  assign \new_[28260]_  = ~\new_[29890]_  | ~\new_[31416]_ ;
  assign \new_[28261]_  = ~\new_[30179]_  & ~\new_[6190]_ ;
  assign \new_[28262]_  = ~\new_[29857]_  & ~\new_[31724]_ ;
  assign \new_[28263]_  = ~\new_[29775]_  | ~\new_[6040]_ ;
  assign \new_[28264]_  = ~\new_[29812]_  | ~\new_[30998]_ ;
  assign \new_[28265]_  = ~\new_[29816]_  & ~\new_[5909]_ ;
  assign \new_[28266]_  = ~\new_[30361]_  & ~\new_[31423]_ ;
  assign \new_[28267]_  = ~\new_[29696]_ ;
  assign \new_[28268]_  = ~\new_[29713]_ ;
  assign \new_[28269]_  = \new_[30164]_  & \new_[5964]_ ;
  assign \new_[28270]_  = ~\new_[30164]_ ;
  assign \new_[28271]_  = ~\new_[29820]_  & ~\new_[6094]_ ;
  assign \new_[28272]_  = ~\new_[29004]_ ;
  assign \new_[28273]_  = ~\new_[29321]_ ;
  assign \new_[28274]_  = ~\new_[30344]_  & ~\new_[29854]_ ;
  assign \new_[28275]_  = ~\new_[30649]_  | ~\new_[30011]_ ;
  assign \new_[28276]_  = ~\new_[30642]_  | ~\new_[30444]_ ;
  assign \new_[28277]_  = ~\new_[30618]_  | ~\new_[5984]_ ;
  assign \new_[28278]_  = ~\new_[29290]_ ;
  assign \new_[28279]_  = ~\new_[30368]_  & ~\new_[31464]_ ;
  assign \new_[28280]_  = ~\new_[29918]_ ;
  assign \new_[28281]_  = ~\new_[28996]_ ;
  assign \new_[28282]_  = \new_[29849]_  & \new_[5999]_ ;
  assign \new_[28283]_  = ~\new_[30044]_ ;
  assign \new_[28284]_  = ~\new_[30057]_ ;
  assign \new_[28285]_  = ~\new_[29595]_ ;
  assign \new_[28286]_  = ~\new_[29885]_  & ~\new_[30021]_ ;
  assign \new_[28287]_  = ~\new_[30286]_  & ~\new_[30615]_ ;
  assign \new_[28288]_  = \new_[29890]_  & \new_[6001]_ ;
  assign \new_[28289]_  = ~\new_[30233]_  | ~\new_[29956]_ ;
  assign \new_[28290]_  = ~\new_[29822]_  | ~\new_[6072]_ ;
  assign \new_[28291]_  = ~\new_[30211]_  | ~\new_[30076]_ ;
  assign \new_[28292]_  = \new_[29834]_  | \new_[6190]_ ;
  assign \new_[28293]_  = ~\new_[29569]_ ;
  assign \new_[28294]_  = ~\new_[30317]_  | ~\new_[29882]_ ;
  assign \new_[28295]_  = ~\new_[30379]_  & ~\new_[5985]_ ;
  assign \new_[28296]_  = ~\new_[29289]_ ;
  assign \new_[28297]_  = ~\new_[30278]_  | ~\new_[30677]_ ;
  assign \new_[28298]_  = \new_[30598]_  | \new_[30152]_ ;
  assign \new_[28299]_  = ~\new_[30385]_  & ~\new_[31724]_ ;
  assign \new_[28300]_  = ~\new_[29920]_  | ~\new_[6033]_ ;
  assign \new_[28301]_  = ~\new_[29873]_  & ~\new_[29861]_ ;
  assign \new_[28302]_  = ~\new_[30292]_  | ~\new_[29888]_ ;
  assign \new_[28303]_  = ~\new_[30226]_  | ~\new_[6196]_ ;
  assign \new_[28304]_  = ~\new_[29488]_ ;
  assign \new_[28305]_  = ~\new_[30105]_  | ~\new_[30277]_ ;
  assign \new_[28306]_  = ~\new_[30218]_  | ~\new_[30642]_ ;
  assign \new_[28307]_  = ~\new_[30208]_ ;
  assign \new_[28308]_  = ~\new_[30289]_  & ~\new_[30000]_ ;
  assign \new_[28309]_  = ~\new_[29131]_ ;
  assign \new_[28310]_  = ~\new_[30324]_  | ~\new_[31419]_ ;
  assign \new_[28311]_  = ~\new_[29487]_ ;
  assign \new_[28312]_  = ~\new_[29106]_ ;
  assign \new_[28313]_  = \new_[31061]_  & \new_[29990]_ ;
  assign \new_[28314]_  = ~\new_[30368]_  & ~\new_[6176]_ ;
  assign \new_[28315]_  = ~\new_[29031]_ ;
  assign \new_[28316]_  = \new_[30394]_  | \new_[5921]_ ;
  assign \new_[28317]_  = ~\new_[30505]_ ;
  assign \new_[28318]_  = ~\new_[30150]_  | ~\new_[6202]_ ;
  assign \new_[28319]_  = ~\new_[29179]_ ;
  assign \new_[28320]_  = ~\new_[30385]_  & ~\new_[5932]_ ;
  assign \new_[28321]_  = \new_[30392]_  | \new_[5926]_ ;
  assign \new_[28322]_  = (~\new_[5917]_  | ~\new_[30796]_ ) & (~\new_[6066]_  | ~\new_[30988]_ );
  assign \new_[28323]_  = ~\new_[30919]_  & ~\new_[5968]_ ;
  assign \new_[28324]_  = ~\new_[29338]_ ;
  assign \new_[28325]_  = \new_[29973]_  | \new_[5918]_ ;
  assign \new_[28326]_  = ~\new_[29580]_ ;
  assign \new_[28327]_  = \new_[29764]_  | \new_[5909]_ ;
  assign \new_[28328]_  = ~\new_[30055]_  & ~\new_[31862]_ ;
  assign \new_[28329]_  = ~\new_[30415]_  & ~\new_[31903]_ ;
  assign \new_[28330]_  = ~\new_[30039]_  & ~\new_[5927]_ ;
  assign \new_[28331]_  = ~\new_[29159]_ ;
  assign \new_[28332]_  = \new_[29766]_  & \new_[31870]_ ;
  assign \new_[28333]_  = ~\new_[29074]_ ;
  assign \new_[28334]_  = ~\new_[30017]_  | ~\new_[30998]_ ;
  assign \new_[28335]_  = ~\new_[29498]_ ;
  assign \new_[28336]_  = ~\new_[29833]_  | ~\new_[30092]_ ;
  assign \new_[28337]_  = ~\new_[28819]_ ;
  assign \new_[28338]_  = ~\new_[29547]_ ;
  assign \new_[28339]_  = ~\new_[30140]_  & ~\new_[31839]_ ;
  assign \new_[28340]_  = ~\new_[29881]_  & ~\new_[30058]_ ;
  assign \new_[28341]_  = ~\new_[30070]_  & ~\new_[30752]_ ;
  assign \new_[28342]_  = ~\new_[28827]_ ;
  assign \new_[28343]_  = ~\new_[29800]_  & ~\new_[6007]_ ;
  assign \new_[28344]_  = ~\new_[30293]_ ;
  assign \new_[28345]_  = ~\new_[29803]_  & ~\new_[31421]_ ;
  assign \new_[28346]_  = ~\new_[30299]_  | ~\new_[30148]_ ;
  assign \new_[28347]_  = ~\new_[28843]_ ;
  assign \new_[28348]_  = ~\new_[30136]_  | ~\new_[6066]_ ;
  assign \new_[28349]_  = ~\new_[30626]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[28350]_  = ~\new_[30709]_  | ~\new_[30968]_  | ~m2_cyc_i;
  assign \new_[28351]_  = ~\new_[30457]_  | ~\new_[31199]_  | ~m4_cyc_i;
  assign \new_[28352]_  = \new_[30030]_  & \new_[6036]_ ;
  assign \new_[28353]_  = ~\new_[30198]_  | ~\new_[30250]_ ;
  assign \new_[28354]_  = \new_[29988]_  | \new_[5911]_ ;
  assign \new_[28355]_  = ~\new_[29789]_ ;
  assign \new_[28356]_  = ~\new_[30241]_  | ~\new_[31148]_ ;
  assign \new_[28357]_  = ~\new_[29175]_ ;
  assign \new_[28358]_  = ~\new_[30574]_ ;
  assign \new_[28359]_  = ~\new_[30572]_  | ~\new_[6070]_ ;
  assign \new_[28360]_  = ~\new_[30103]_  | ~\new_[5907]_ ;
  assign \new_[28361]_  = ~\new_[30257]_  & ~\new_[30076]_ ;
  assign \new_[28362]_  = ~\new_[29192]_ ;
  assign \new_[28363]_  = ~\new_[29910]_  | ~\new_[5904]_ ;
  assign \new_[28364]_  = ~\new_[30699]_  & ~\new_[5931]_ ;
  assign \new_[28365]_  = ~\new_[29348]_ ;
  assign \new_[28366]_  = ~\new_[29381]_ ;
  assign \new_[28367]_  = ~\new_[30398]_  & ~\new_[6096]_ ;
  assign \new_[28368]_  = ~\new_[30325]_  | ~\new_[30799]_ ;
  assign \new_[28369]_  = ~\new_[30207]_  & ~\new_[30340]_ ;
  assign \new_[28370]_  = ~\new_[30432]_  | ~\new_[30340]_ ;
  assign \new_[28371]_  = ~\new_[29383]_ ;
  assign \new_[28372]_  = ~\new_[30317]_  | ~\new_[5927]_ ;
  assign \new_[28373]_  = ~\new_[30267]_  | ~\new_[30061]_ ;
  assign \new_[28374]_  = ~\new_[30153]_  | ~\new_[5917]_ ;
  assign \new_[28375]_  = ~\new_[29135]_ ;
  assign \new_[28376]_  = ~\new_[30240]_  & ~\new_[29787]_ ;
  assign \new_[28377]_  = (~\new_[30590]_  | ~\new_[5908]_ ) & (~\new_[30935]_  | ~\new_[6092]_ );
  assign \new_[28378]_  = ~\new_[30000]_  | ~\new_[6046]_ ;
  assign \new_[28379]_  = ~\new_[29278]_ ;
  assign \new_[28380]_  = ~\new_[29841]_  & ~\new_[30030]_ ;
  assign \new_[28381]_  = ~\new_[29791]_  & ~\new_[30246]_ ;
  assign \new_[28382]_  = ~\new_[30035]_  | ~\new_[5901]_ ;
  assign \new_[28383]_  = ~\new_[29799]_  & ~\new_[30084]_ ;
  assign \new_[28384]_  = ~\new_[29881]_  | ~\new_[30127]_ ;
  assign \new_[28385]_  = ~\new_[29991]_  & ~\new_[30726]_ ;
  assign \new_[28386]_  = (~\new_[5914]_  | ~\new_[30587]_ ) & (~\new_[6207]_  | ~\new_[31212]_ );
  assign \new_[28387]_  = ~\new_[30338]_  | ~\new_[30969]_ ;
  assign \new_[28388]_  = (~\new_[30738]_  | ~\new_[5907]_ ) & (~\new_[31187]_  | ~\new_[6215]_ );
  assign \new_[28389]_  = \new_[30296]_  & \new_[6245]_ ;
  assign \new_[28390]_  = (~\new_[6045]_  | ~\new_[30625]_ ) & (~\new_[6199]_  | ~\new_[30859]_ );
  assign \new_[28391]_  = ~\new_[30276]_  & ~\new_[31799]_ ;
  assign \new_[28392]_  = \new_[30562]_  & \new_[29804]_ ;
  assign \new_[28393]_  = ~\new_[30215]_ ;
  assign \new_[28394]_  = ~\new_[30337]_  | ~\new_[6037]_ ;
  assign \new_[28395]_  = ~\new_[29211]_ ;
  assign \new_[28396]_  = ~\new_[29364]_ ;
  assign \new_[28397]_  = ~\new_[30346]_  & ~\new_[4231]_ ;
  assign \new_[28398]_  = ~\new_[30015]_  & ~\new_[29991]_ ;
  assign \new_[28399]_  = ~\new_[29966]_  & ~\new_[31616]_ ;
  assign \new_[28400]_  = ~\new_[30326]_  & ~\new_[30136]_ ;
  assign \new_[28401]_  = \new_[29841]_  | \new_[29855]_ ;
  assign \new_[28402]_  = ~\new_[30217]_ ;
  assign \new_[28403]_  = (~\new_[6087]_  | ~\new_[30738]_ ) & (~\new_[6089]_  | ~\new_[31187]_ );
  assign \new_[28404]_  = ~\new_[30161]_  | ~\new_[5908]_ ;
  assign \new_[28405]_  = ~\new_[30142]_  | ~\new_[6186]_ ;
  assign \new_[28406]_  = ~\new_[30242]_  & ~\new_[30051]_ ;
  assign \new_[28407]_  = ~\new_[30706]_  & ~\new_[29996]_ ;
  assign \new_[28408]_  = ~\new_[29642]_ ;
  assign \new_[28409]_  = ~\new_[29550]_ ;
  assign \new_[28410]_  = ~\new_[30183]_  | ~\new_[5978]_ ;
  assign \new_[28411]_  = ~\new_[30677]_  | ~\new_[30786]_ ;
  assign \new_[28412]_  = ~\new_[30245]_  | ~\new_[30097]_ ;
  assign \new_[28413]_  = ~\new_[30411]_  | ~\new_[6088]_ ;
  assign \new_[28414]_  = ~\new_[29782]_  | ~\new_[6053]_ ;
  assign \new_[28415]_  = ~\new_[29873]_  | ~\new_[6094]_ ;
  assign \new_[28416]_  = ~\new_[30029]_  | ~\new_[30782]_ ;
  assign \new_[28417]_  = ~\new_[29551]_ ;
  assign \new_[28418]_  = ~\new_[30374]_  & ~\new_[5964]_ ;
  assign \new_[28419]_  = ~\new_[29808]_  | ~\new_[29915]_ ;
  assign \new_[28420]_  = ~\new_[30183]_  | ~\new_[30234]_ ;
  assign \new_[28421]_  = ~\new_[30145]_  & ~\new_[30322]_ ;
  assign \new_[28422]_  = ~\new_[30079]_  & ~\new_[30314]_ ;
  assign \new_[28423]_  = ~\new_[30128]_  | ~\new_[5908]_ ;
  assign \new_[28424]_  = ~\new_[30371]_  & ~\new_[5909]_ ;
  assign \new_[28425]_  = ~\new_[30043]_  | ~\new_[30061]_ ;
  assign \new_[28426]_  = ~\new_[29433]_ ;
  assign \new_[28427]_  = ~\new_[29798]_  | ~\new_[6092]_ ;
  assign \new_[28428]_  = ~\new_[29861]_  & ~\new_[31474]_ ;
  assign \new_[28429]_  = ~\new_[29944]_  | ~\new_[30009]_ ;
  assign \new_[28430]_  = \new_[29859]_  | \new_[6066]_ ;
  assign \new_[28431]_  = ~\new_[30299]_  | ~\new_[6004]_ ;
  assign \new_[28432]_  = ~\new_[30054]_  | ~\new_[6002]_ ;
  assign \new_[28433]_  = ~\new_[30381]_  | ~\new_[5918]_ ;
  assign \new_[28434]_  = ~\new_[30717]_  | ~\new_[6057]_ ;
  assign \new_[28435]_  = ~\new_[31741]_  & ~\new_[6049]_ ;
  assign \new_[28436]_  = ~\new_[30352]_  | ~\new_[6089]_ ;
  assign \new_[28437]_  = ~\new_[30223]_  | ~\new_[5900]_ ;
  assign \new_[28438]_  = ~\new_[29924]_  | ~\new_[5909]_ ;
  assign \new_[28439]_  = ~\new_[30367]_  | ~\new_[6215]_ ;
  assign \new_[28440]_  = ~\new_[30081]_  | ~\new_[6210]_ ;
  assign \new_[28441]_  = \new_[30132]_  & \new_[5967]_ ;
  assign \new_[28442]_  = ~\new_[29802]_  | ~\new_[6191]_ ;
  assign \new_[28443]_  = ~\new_[29837]_  | ~\new_[6078]_ ;
  assign \new_[28444]_  = ~\new_[30163]_  | ~\new_[5901]_ ;
  assign \new_[28445]_  = ~\new_[30011]_  | ~\new_[6050]_ ;
  assign \new_[28446]_  = ~\new_[29941]_  | ~\new_[5983]_ ;
  assign \new_[28447]_  = ~\new_[30046]_  | ~\new_[5907]_ ;
  assign \new_[28448]_  = ~\new_[30058]_  & ~\new_[31707]_ ;
  assign \new_[28449]_  = ~\new_[30258]_  | ~\new_[5917]_ ;
  assign \new_[28450]_  = ~\new_[29971]_  | ~\new_[6207]_ ;
  assign \new_[28451]_  = ~\new_[30169]_  | ~\new_[6196]_ ;
  assign \new_[28452]_  = ~\new_[30444]_  | ~\new_[6215]_ ;
  assign \new_[28453]_  = ~\new_[30211]_  | ~\new_[5923]_ ;
  assign \new_[28454]_  = ~\new_[30003]_  & ~\new_[30799]_ ;
  assign \new_[28455]_  = ~\new_[30295]_  | ~\new_[6084]_ ;
  assign \new_[28456]_  = ~\new_[29841]_  & ~\new_[31800]_ ;
  assign \new_[28457]_  = ~\new_[29867]_  | ~\new_[6194]_ ;
  assign \new_[28458]_  = ~\new_[29975]_  | ~\new_[6043]_ ;
  assign \new_[28459]_  = ~\new_[30037]_  | ~\new_[6049]_ ;
  assign \new_[28460]_  = ~\new_[30322]_  | ~\new_[6033]_ ;
  assign \new_[28461]_  = ~\new_[30290]_  | ~\new_[6270]_ ;
  assign \new_[28462]_  = ~\new_[29889]_  & ~\new_[29971]_ ;
  assign \new_[28463]_  = ~\new_[30152]_  | ~\new_[6034]_ ;
  assign \new_[28464]_  = ~\new_[30009]_  | ~\new_[6080]_ ;
  assign \new_[28465]_  = ~\new_[29853]_  & ~\new_[31593]_ ;
  assign \new_[28466]_  = ~\new_[30196]_  | ~\new_[5933]_ ;
  assign \new_[28467]_  = ~\new_[29944]_  & ~\new_[31765]_ ;
  assign \new_[28468]_  = ~\new_[30271]_  | ~\new_[6216]_ ;
  assign \new_[28469]_  = ~\new_[30283]_  | ~\new_[6174]_ ;
  assign \new_[28470]_  = \new_[30057]_  & \new_[6045]_ ;
  assign \new_[28471]_  = \new_[29972]_  & \new_[6085]_ ;
  assign \new_[28472]_  = ~\new_[30342]_  & ~\new_[30329]_ ;
  assign \new_[28473]_  = ~\new_[30004]_  & ~\new_[30215]_ ;
  assign \new_[28474]_  = ~\new_[30062]_  | ~\new_[29863]_ ;
  assign \new_[28475]_  = ~\new_[30123]_  | ~\new_[30208]_ ;
  assign \new_[28476]_  = ~\new_[29827]_  & ~\new_[31660]_ ;
  assign \new_[28477]_  = ~\new_[30151]_  | ~\new_[30630]_ ;
  assign \new_[28478]_  = ~\new_[30545]_  | ~\new_[29798]_ ;
  assign \new_[28479]_  = ~\new_[29776]_  & ~\new_[30022]_ ;
  assign \new_[28480]_  = ~\new_[30308]_  | ~\new_[29887]_ ;
  assign \new_[28481]_  = ~\new_[29780]_  | ~\new_[30785]_ ;
  assign \new_[28482]_  = ~\new_[30094]_  | ~\new_[5914]_ ;
  assign \new_[28483]_  = ~\new_[30025]_  | ~\new_[29960]_ ;
  assign \new_[28484]_  = ~\new_[30205]_  | ~\new_[30789]_ ;
  assign \new_[28485]_  = ~\new_[30329]_  | ~\new_[30574]_ ;
  assign \new_[28486]_  = ~\new_[29098]_ ;
  assign \new_[28487]_  = ~\new_[29635]_ ;
  assign \new_[28488]_  = ~\new_[29453]_ ;
  assign \new_[28489]_  = ~\new_[29806]_  & ~\new_[30721]_ ;
  assign \new_[28490]_  = ~\new_[29772]_  | ~\new_[30016]_ ;
  assign \new_[28491]_  = ~\new_[30162]_  & ~\new_[30751]_ ;
  assign \new_[28492]_  = ~\new_[30318]_  | ~\new_[30629]_ ;
  assign \new_[28493]_  = ~\new_[28951]_ ;
  assign \new_[28494]_  = ~\new_[30033]_  | ~\new_[30752]_ ;
  assign \new_[28495]_  = ~\new_[30730]_  & ~\new_[29880]_ ;
  assign \new_[28496]_  = ~\new_[30038]_  | ~\new_[30555]_ ;
  assign \new_[28497]_  = ~\new_[30478]_  | ~\new_[30213]_ ;
  assign \new_[28498]_  = ~\new_[30697]_  | ~\new_[31422]_ ;
  assign \new_[28499]_  = ~\new_[30020]_  | ~\new_[30582]_ ;
  assign \new_[28500]_  = ~\new_[29765]_  | ~\new_[30172]_ ;
  assign \new_[28501]_  = ~\new_[30280]_  | ~\new_[29772]_ ;
  assign \new_[28502]_  = \new_[30133]_  & \new_[6269]_ ;
  assign \new_[28503]_  = ~\new_[30828]_  & ~\new_[29853]_ ;
  assign \new_[28504]_  = ~\new_[30293]_  & ~\new_[30340]_ ;
  assign \new_[28505]_  = ~\new_[30415]_  | ~\new_[5896]_ ;
  assign \new_[28506]_  = ~\new_[29158]_ ;
  assign \new_[28507]_  = ~\new_[30363]_  | ~\new_[30032]_ ;
  assign \new_[28508]_  = ~\new_[29777]_  | ~\new_[29984]_ ;
  assign \new_[28509]_  = ~\new_[30262]_  | ~\new_[6093]_ ;
  assign \new_[28510]_  = ~\new_[30094]_  | ~\new_[29814]_ ;
  assign \new_[28511]_  = ~\new_[29831]_  | ~\new_[5976]_ ;
  assign \new_[28512]_  = ~\new_[29979]_  | ~\new_[6076]_ ;
  assign \new_[28513]_  = \new_[30210]_  & \new_[5922]_ ;
  assign \new_[28514]_  = ~\new_[30255]_  | ~\new_[30446]_ ;
  assign \new_[28515]_  = ~\new_[29926]_  & ~\new_[30410]_ ;
  assign \new_[28516]_  = ~\new_[28821]_ ;
  assign \new_[28517]_  = ~\new_[29841]_  | ~\new_[5895]_ ;
  assign \new_[28518]_  = ~\new_[30400]_  & ~\new_[31553]_ ;
  assign \new_[28519]_  = ~\new_[30139]_  | ~\new_[29950]_ ;
  assign \new_[28520]_  = ~\new_[30151]_  | ~\new_[30290]_ ;
  assign \new_[28521]_  = ~\new_[30140]_  | ~\new_[5906]_ ;
  assign \new_[28522]_  = ~\new_[30409]_  | ~\new_[29777]_ ;
  assign \new_[28523]_  = ~\new_[29968]_  | ~\new_[30084]_ ;
  assign \new_[28524]_  = ~\new_[30703]_  | ~\new_[30213]_ ;
  assign \new_[28525]_  = ~\new_[29975]_  | ~\new_[30633]_ ;
  assign \new_[28526]_  = ~\new_[30095]_  & ~\new_[31665]_ ;
  assign \new_[28527]_  = ~\new_[29992]_  | ~\new_[29874]_ ;
  assign \new_[28528]_  = ~\new_[29787]_  | ~\new_[5990]_ ;
  assign \new_[28529]_  = ~\new_[30321]_  | ~\new_[6073]_ ;
  assign \new_[28530]_  = ~\new_[29944]_  | ~\new_[5933]_ ;
  assign \new_[28531]_  = ~\new_[30282]_  & ~\new_[30202]_ ;
  assign \new_[28532]_  = ~\new_[29907]_  | ~\new_[30754]_ ;
  assign \new_[28533]_  = ~\new_[30107]_  | ~\new_[6071]_ ;
  assign \new_[28534]_  = \new_[29996]_  & \new_[6217]_ ;
  assign \new_[28535]_  = ~\new_[30098]_  | ~\new_[4440]_ ;
  assign \new_[28536]_  = ~\new_[30257]_  | ~\new_[5905]_ ;
  assign \new_[28537]_  = ~\new_[30597]_  | ~\new_[31440]_ ;
  assign \new_[28538]_  = ~\new_[29865]_  | ~\new_[29904]_ ;
  assign \new_[28539]_  = ~\new_[30244]_  & ~\new_[31900]_ ;
  assign \new_[28540]_  = ~\new_[29790]_  | ~\new_[30538]_ ;
  assign \new_[28541]_  = ~\new_[30102]_  | ~\new_[30314]_ ;
  assign \new_[28542]_  = ~\new_[29761]_ ;
  assign \new_[28543]_  = ~\new_[30407]_  & ~\new_[31608]_ ;
  assign \new_[28544]_  = ~\new_[30203]_  | ~\new_[29762]_ ;
  assign \new_[28545]_  = \new_[30019]_  & \new_[5894]_ ;
  assign \new_[28546]_  = ~\new_[29869]_  & ~\new_[29962]_ ;
  assign \new_[28547]_  = ~\new_[29870]_  | ~\new_[6197]_ ;
  assign \new_[28548]_  = ~\new_[30083]_  & ~\new_[30235]_ ;
  assign \new_[28549]_  = ~\new_[30173]_  & ~\new_[31643]_ ;
  assign \new_[28550]_  = ~\new_[29877]_  | ~\new_[30703]_ ;
  assign \new_[28551]_  = ~\new_[30505]_  | ~\new_[30253]_ ;
  assign \new_[28552]_  = ~\new_[28961]_ ;
  assign \new_[28553]_  = ~\new_[29555]_ ;
  assign \new_[28554]_  = ~\new_[30258]_  | ~\new_[30052]_ ;
  assign \new_[28555]_  = ~\new_[30145]_  | ~\new_[30416]_ ;
  assign \new_[28556]_  = ~\new_[30178]_  | ~\new_[30618]_ ;
  assign \new_[28557]_  = ~\new_[29494]_ ;
  assign \new_[28558]_  = ~\new_[29840]_  & ~\new_[29944]_ ;
  assign \new_[28559]_  = ~\new_[30086]_  | ~\new_[29994]_ ;
  assign \new_[28560]_  = ~\new_[30279]_  | ~\new_[6063]_ ;
  assign \new_[28561]_  = ~\new_[29967]_  | ~\new_[6195]_ ;
  assign \new_[28562]_  = ~\new_[29978]_  | ~\new_[6212]_ ;
  assign \new_[28563]_  = ~\new_[29787]_  | ~\new_[30125]_ ;
  assign \new_[28564]_  = ~\new_[29792]_  | ~\new_[30563]_ ;
  assign \new_[28565]_  = ~\new_[30294]_  | ~\new_[30216]_ ;
  assign \new_[28566]_  = ~\new_[29935]_  & ~\new_[30695]_ ;
  assign \new_[28567]_  = ~\new_[30205]_  | ~\new_[6085]_ ;
  assign \new_[28568]_  = ~\new_[30553]_  & ~\new_[29978]_ ;
  assign \new_[28569]_  = ~\new_[30072]_  | ~\new_[30021]_ ;
  assign \new_[28570]_  = ~\new_[29902]_  | ~\new_[29929]_ ;
  assign \new_[28571]_  = ~\new_[30273]_  & ~\new_[30842]_ ;
  assign \new_[28572]_  = ~\new_[30198]_  & ~\new_[30286]_ ;
  assign \new_[28573]_  = ~\new_[30343]_  | ~\new_[30662]_ ;
  assign \new_[28574]_  = ~\new_[29941]_  | ~\new_[29940]_ ;
  assign \new_[28575]_  = ~\new_[30304]_  | ~\new_[29888]_ ;
  assign \new_[28576]_  = ~\new_[30253]_  & ~\new_[30573]_ ;
  assign \new_[28577]_  = \new_[30140]_  | \new_[29898]_ ;
  assign \new_[28578]_  = ~\new_[30044]_  & ~\new_[29984]_ ;
  assign \new_[28579]_  = ~\new_[30597]_  | ~\new_[30697]_ ;
  assign \new_[28580]_  = ~\new_[29828]_  & ~\new_[30432]_ ;
  assign \new_[28581]_  = ~\new_[30133]_  | ~\new_[31104]_ ;
  assign \new_[28582]_  = ~\new_[30036]_  & ~\new_[31789]_ ;
  assign \new_[28583]_  = ~\new_[29964]_  & ~\new_[30610]_ ;
  assign \new_[28584]_  = ~\new_[30317]_  & ~\new_[30140]_ ;
  assign \new_[28585]_  = ~\new_[29794]_  | ~\new_[30540]_ ;
  assign \new_[28586]_  = ~\new_[29826]_  | ~\new_[30215]_ ;
  assign \new_[28587]_  = ~\new_[30201]_  | ~\new_[30719]_ ;
  assign \new_[28588]_  = ~\new_[30364]_  & ~\new_[5997]_ ;
  assign \new_[28589]_  = (~\new_[30489]_  | ~\new_[5906]_ ) & (~\new_[31094]_  | ~\new_[5928]_ );
  assign \new_[28590]_  = (~\new_[30587]_  | ~\new_[6051]_ ) & (~\new_[30877]_  | ~\new_[5973]_ );
  assign \new_[28591]_  = (~\new_[5912]_  | ~\new_[30625]_ ) & (~\new_[6096]_  | ~\new_[30859]_ );
  assign \new_[28592]_  = (~\new_[6091]_  | ~\new_[30590]_ ) & (~\new_[6093]_  | ~\new_[30935]_ );
  assign \new_[28593]_  = (~\new_[30796]_  | ~\new_[5902]_ ) & (~\new_[30988]_  | ~\new_[5984]_ );
  assign \new_[28594]_  = (~\new_[6004]_  | ~\new_[30590]_ ) & (~\new_[6216]_  | ~\new_[30935]_ );
  assign \new_[28595]_  = ~\new_[29300]_ ;
  assign \new_[28596]_  = (~\new_[5927]_  | ~\new_[30489]_ ) & (~\new_[6084]_  | ~\new_[31094]_ );
  assign \new_[28597]_  = (~\new_[6002]_  | ~\new_[30738]_ ) & (~\new_[6184]_  | ~\new_[31187]_ );
  assign \new_[28598]_  = \new_[30034]_  & \new_[5990]_ ;
  assign \new_[28599]_  = \new_[29770]_  | \new_[31648]_ ;
  assign \new_[28600]_  = ~\new_[29155]_ ;
  assign \new_[28601]_  = ~\new_[29385]_ ;
  assign \new_[28602]_  = ~\new_[29532]_ ;
  assign \new_[28603]_  = \new_[30402]_  | \new_[5912]_ ;
  assign \new_[28604]_  = ~\new_[29802]_  | ~\new_[30348]_ ;
  assign \new_[28605]_  = ~\new_[29110]_ ;
  assign \new_[28606]_  = ~\new_[30054]_  | ~\new_[30399]_ ;
  assign \new_[28607]_  = \new_[29872]_  | \new_[5983]_ ;
  assign \new_[28608]_  = ~\new_[29265]_ ;
  assign \new_[28609]_  = ~\new_[29064]_ ;
  assign \new_[28610]_  = ~\new_[29505]_ ;
  assign \new_[28611]_  = ~\new_[29310]_ ;
  assign \new_[28612]_  = ~\new_[29539]_ ;
  assign \new_[28613]_  = \new_[30096]_  | \new_[5978]_ ;
  assign \new_[28614]_  = ~\new_[29674]_ ;
  assign \new_[28615]_  = ~\new_[29675]_ ;
  assign \new_[28616]_  = ~\new_[29538]_ ;
  assign \new_[28617]_  = \new_[29862]_  | \new_[5913]_ ;
  assign \new_[28618]_  = ~\new_[29373]_ ;
  assign \new_[28619]_  = ~\new_[28971]_ ;
  assign \new_[28620]_  = \new_[30393]_  | \new_[5927]_ ;
  assign \new_[28621]_  = \new_[29943]_  & \new_[5900]_ ;
  assign \new_[28622]_  = ~\new_[29161]_ ;
  assign \new_[28623]_  = ~\new_[28922]_ ;
  assign \new_[28624]_  = ~\new_[29542]_ ;
  assign \new_[28625]_  = ~\new_[28986]_ ;
  assign \new_[28626]_  = ~\new_[28841]_ ;
  assign \new_[28627]_  = ~\new_[29358]_ ;
  assign \new_[28628]_  = ~\new_[30177]_  | ~\new_[5924]_ ;
  assign \new_[28629]_  = ~\new_[30274]_  & ~\new_[5913]_ ;
  assign \new_[28630]_  = ~\new_[30657]_  & ~\new_[5968]_ ;
  assign \new_[28631]_  = ~\new_[29914]_  | ~\new_[30092]_ ;
  assign \new_[28632]_  = ~\new_[30121]_  | ~\new_[30316]_ ;
  assign \new_[28633]_  = ~\new_[28975]_ ;
  assign \new_[28634]_  = ~\new_[30002]_  | ~\new_[30574]_ ;
  assign \new_[28635]_  = ~\new_[29337]_ ;
  assign \new_[28636]_  = ~\new_[29353]_ ;
  assign \new_[28637]_  = ~\new_[29010]_ ;
  assign \new_[28638]_  = ~\new_[29334]_ ;
  assign \new_[28639]_  = ~\new_[30922]_  & ~\new_[31407]_ ;
  assign \new_[28640]_  = ~\new_[30315]_ ;
  assign \new_[28641]_  = ~\new_[29994]_ ;
  assign \new_[28642]_  = ~\new_[29345]_ ;
  assign \new_[28643]_  = ~\new_[29997]_  | ~\new_[30725]_ ;
  assign \new_[28644]_  = ~\new_[30283]_  | ~\new_[29853]_ ;
  assign \new_[28645]_  = ~\new_[29884]_  & ~\new_[6246]_ ;
  assign \new_[28646]_  = ~\new_[29282]_ ;
  assign \new_[28647]_  = \new_[29795]_  | \new_[5978]_ ;
  assign \new_[28648]_  = ~\new_[29146]_ ;
  assign \new_[28649]_  = ~\new_[29325]_ ;
  assign \new_[28650]_  = ~\new_[29027]_ ;
  assign \new_[28651]_  = ~\new_[30351]_  | ~\new_[31712]_ ;
  assign \new_[28652]_  = ~\new_[29752]_ ;
  assign \new_[28653]_  = ~\new_[29832]_  | ~\new_[31787]_ ;
  assign \new_[28654]_  = ~\new_[29808]_  & ~\new_[29883]_ ;
  assign \new_[28655]_  = ~\new_[29790]_  & ~\new_[30107]_ ;
  assign \new_[28656]_  = ~\new_[30365]_  & ~\new_[5918]_ ;
  assign \new_[28657]_  = \new_[29803]_  | \new_[5997]_ ;
  assign \new_[28658]_  = ~\new_[30221]_ ;
  assign \new_[28659]_  = \new_[30202]_  | \new_[30389]_ ;
  assign \new_[28660]_  = ~\new_[29446]_ ;
  assign \new_[28661]_  = ~\new_[29416]_ ;
  assign \new_[28662]_  = ~\new_[30397]_  & ~\new_[6059]_ ;
  assign \new_[28663]_  = ~\new_[30277]_ ;
  assign \new_[28664]_  = (~\new_[6075]_  | ~\new_[30704]_ ) & (~\new_[6076]_  | ~\new_[31072]_ );
  assign \new_[28665]_  = ~\new_[29114]_ ;
  assign \new_[28666]_  = ~\new_[29584]_ ;
  assign \new_[28667]_  = ~\new_[29677]_ ;
  assign \new_[28668]_  = ~\new_[30437]_  & ~\new_[29915]_ ;
  assign \new_[28669]_  = ~\new_[29303]_ ;
  assign \new_[28670]_  = ~\new_[29797]_  & ~\new_[31665]_ ;
  assign \new_[28671]_  = \new_[30372]_  & \new_[6190]_ ;
  assign \new_[28672]_  = ~\new_[30541]_  & ~\new_[30296]_ ;
  assign \new_[28673]_  = \new_[29793]_  | \new_[5926]_ ;
  assign \new_[28674]_  = ~\new_[30326]_  | ~\new_[30814]_ ;
  assign \new_[28675]_  = ~\new_[28999]_ ;
  assign \new_[28676]_  = ~\new_[30033]_  & ~\new_[30169]_ ;
  assign \new_[28677]_  = ~\new_[30380]_  | ~\new_[6216]_ ;
  assign \new_[28678]_  = ~\new_[28969]_ ;
  assign \new_[28679]_  = ~\new_[30378]_  & ~\new_[31104]_ ;
  assign \new_[28680]_  = ~\new_[29938]_  | ~\new_[31645]_ ;
  assign \new_[28681]_  = ~\new_[30597]_  | ~\new_[31422]_ ;
  assign \new_[28682]_  = ~\new_[28930]_ ;
  assign \new_[28683]_  = ~\new_[28925]_ ;
  assign \new_[28684]_  = ~\new_[29854]_ ;
  assign \new_[28685]_  = ~\new_[30139]_ ;
  assign \new_[28686]_  = ~\new_[30135]_ ;
  assign \new_[28687]_  = ~\new_[29853]_  & ~\new_[30416]_ ;
  assign \new_[28688]_  = ~\new_[29864]_  & ~\new_[5912]_ ;
  assign \new_[28689]_  = ~\new_[30440]_  & ~\new_[31132]_ ;
  assign \new_[28690]_  = ~\new_[29850]_  & ~\new_[5921]_ ;
  assign \new_[28691]_  = ~\new_[29756]_ ;
  assign \new_[28692]_  = ~\new_[29486]_ ;
  assign \new_[28693]_  = ~\new_[30722]_  & ~\new_[6246]_ ;
  assign \new_[28694]_  = ~\new_[29250]_ ;
  assign \new_[28695]_  = ~\new_[32328]_ ;
  assign \new_[28696]_  = ~\new_[29730]_ ;
  assign \new_[28697]_  = ~\new_[29622]_ ;
  assign \new_[28698]_  = ~\new_[29243]_ ;
  assign \new_[28699]_  = ~\new_[29232]_ ;
  assign \new_[28700]_  = ~\new_[29913]_  | ~\new_[30170]_ ;
  assign \new_[28701]_  = ~\new_[30388]_  & ~\new_[6176]_ ;
  assign \new_[28702]_  = \new_[29832]_  & \new_[5991]_ ;
  assign \new_[28703]_  = ~\new_[30228]_  & ~\new_[30538]_ ;
  assign \new_[28704]_  = ~\new_[30040]_  | ~\new_[30320]_ ;
  assign \new_[28705]_  = ~\new_[28862]_ ;
  assign \new_[28706]_  = ~\new_[30359]_  | ~\new_[6210]_ ;
  assign \new_[28707]_  = ~\new_[30247]_  & ~\new_[30628]_ ;
  assign \new_[28708]_  = ~\new_[30180]_  | ~\new_[30710]_ ;
  assign \new_[28709]_  = ~\new_[28991]_ ;
  assign \new_[28710]_  = ~\new_[29933]_  | ~\new_[6208]_ ;
  assign \new_[28711]_  = ~\new_[29686]_ ;
  assign \new_[28712]_  = ~\new_[32268]_ ;
  assign \new_[28713]_  = ~\new_[28882]_ ;
  assign \new_[28714]_  = ~\new_[30867]_  & ~\new_[30778]_ ;
  assign \new_[28715]_  = ~\new_[29733]_ ;
  assign \new_[28716]_  = ~\new_[29194]_ ;
  assign \new_[28717]_  = ~\new_[29800]_  & ~\new_[31855]_ ;
  assign \new_[28718]_  = ~\new_[29150]_ ;
  assign \new_[28719]_  = ~\new_[29343]_ ;
  assign \new_[28720]_  = ~\new_[30360]_  | ~\new_[31043]_ ;
  assign \new_[28721]_  = ~\new_[29030]_ ;
  assign \new_[28722]_  = ~\new_[29810]_  | ~\new_[30676]_ ;
  assign \new_[28723]_  = ~\new_[29852]_  & ~\new_[5964]_ ;
  assign \new_[28724]_  = ~\new_[29898]_ ;
  assign \new_[28725]_  = ~\new_[30029]_  & ~\new_[30081]_ ;
  assign \new_[28726]_  = \new_[31152]_  & \new_[30050]_ ;
  assign \new_[28727]_  = ~\new_[30095]_  & ~\new_[29969]_ ;
  assign \new_[28728]_  = ~\new_[30364]_  & ~\new_[31421]_ ;
  assign \new_[28729]_  = \new_[30949]_  | \new_[5968]_ ;
  assign \new_[28730]_  = ~\new_[29917]_  & ~\new_[31870]_ ;
  assign \new_[28731]_  = ~\new_[29995]_  & ~\new_[30147]_ ;
  assign \new_[28732]_  = ~\new_[29809]_ ;
  assign \new_[28733]_  = \new_[30107]_  & \new_[6192]_ ;
  assign \new_[28734]_  = ~\new_[28875]_ ;
  assign \new_[28735]_  = ~\new_[30351]_  | ~\new_[30952]_ ;
  assign \new_[28736]_  = ~\new_[30405]_  & ~\new_[5923]_ ;
  assign \new_[28737]_  = ~\new_[29140]_ ;
  assign \new_[28738]_  = ~\new_[30370]_  | ~\new_[31390]_ ;
  assign \new_[28739]_  = ~\new_[28858]_ ;
  assign \new_[28740]_  = ~\new_[30104]_  | ~\new_[30042]_ ;
  assign \new_[28741]_  = ~\new_[29936]_  & ~\new_[31165]_ ;
  assign \new_[28742]_  = ~\new_[30154]_  & ~\new_[31406]_ ;
  assign \new_[28743]_  = ~\new_[29867]_  | ~\new_[30350]_ ;
  assign \new_[28744]_  = ~\new_[30264]_  & ~\new_[5912]_ ;
  assign \new_[28745]_  = ~\new_[30207]_  | ~\new_[30293]_ ;
  assign \new_[28746]_  = ~\new_[29716]_ ;
  assign \new_[28747]_  = ~\new_[29927]_  | ~\new_[6183]_ ;
  assign \new_[28748]_  = ~\new_[29874]_ ;
  assign \new_[28749]_  = ~\new_[30158]_  | ~\new_[6077]_ ;
  assign \new_[28750]_  = ~\new_[29638]_ ;
  assign \new_[28751]_  = ~\new_[29834]_  & ~\new_[31482]_ ;
  assign \new_[28752]_  = ~\new_[29078]_ ;
  assign \new_[28753]_  = ~\new_[29862]_  & ~\new_[31159]_ ;
  assign \new_[28754]_  = \new_[29866]_  | \new_[31614]_ ;
  assign \new_[28755]_  = \new_[29857]_  | \new_[5932]_ ;
  assign \new_[28756]_  = ~\new_[29126]_ ;
  assign \new_[28757]_  = \new_[30372]_  & \new_[31482]_ ;
  assign \new_[28758]_  = ~\new_[29878]_  & ~\new_[31176]_ ;
  assign \new_[28759]_  = ~\new_[29796]_  | ~\new_[31441]_ ;
  assign \new_[28760]_  = \new_[30112]_  & \new_[6007]_ ;
  assign \new_[28761]_  = ~\new_[29057]_ ;
  assign \new_[28762]_  = ~\new_[29699]_ ;
  assign \new_[28763]_  = \new_[29923]_  | \new_[6078]_ ;
  assign \new_[28764]_  = ~\new_[29936]_  & ~\new_[6206]_ ;
  assign \new_[28765]_  = ~\new_[29703]_ ;
  assign \new_[28766]_  = \new_[30376]_  & \m3_addr_i[28] ;
  assign \new_[28767]_  = \new_[29804]_  & \new_[31206]_ ;
  assign \new_[28768]_  = \new_[29804]_  & \new_[31155]_ ;
  assign \new_[28769]_  = ~\new_[29812]_  | ~\new_[31442]_ ;
  assign \new_[28770]_  = ~\new_[6197]_  & ~\new_[31596]_ ;
  assign \new_[28771]_  = ~\new_[30362]_  & ~\new_[5999]_ ;
  assign \new_[28772]_  = ~\new_[30146]_  | ~\new_[30597]_ ;
  assign \new_[28773]_  = ~\new_[29549]_ ;
  assign \new_[28774]_  = ~\new_[29458]_ ;
  assign \new_[28775]_  = \new_[30361]_  | \new_[31690]_ ;
  assign \new_[28776]_  = ~\new_[31440]_  & ~\new_[31588]_ ;
  assign \new_[28777]_  = \new_[29903]_  | \new_[5978]_ ;
  assign \new_[28778]_  = ~\new_[6186]_  & ~\new_[31901]_ ;
  assign \new_[28779]_  = ~\new_[30252]_  | ~\new_[5983]_ ;
  assign \new_[28780]_  = ~\new_[30395]_  | ~\new_[31539]_ ;
  assign \new_[28781]_  = ~\new_[29546]_ ;
  assign \new_[28782]_  = ~\new_[29731]_ ;
  assign \new_[28783]_  = ~\new_[28896]_ ;
  assign \new_[28784]_  = ~\new_[29989]_  & ~\new_[30563]_ ;
  assign \new_[28785]_  = ~\new_[30820]_ ;
  assign \new_[28786]_  = ~\new_[29777]_ ;
  assign \new_[28787]_  = ~\new_[29427]_ ;
  assign \new_[28788]_  = \new_[30410]_  & \new_[6048]_ ;
  assign \new_[28789]_  = ~\new_[29755]_ ;
  assign \new_[28790]_  = ~\new_[29548]_ ;
  assign \new_[28791]_  = ~\new_[29191]_ ;
  assign \new_[28792]_  = ~\new_[29063]_ ;
  assign \new_[28793]_  = ~\new_[29368]_ ;
  assign \new_[28794]_  = ~\new_[29962]_  & ~\new_[30765]_ ;
  assign \new_[28795]_  = ~\new_[29084]_ ;
  assign \new_[28796]_  = (~\new_[30704]_  | ~\new_[5905]_ ) & (~\new_[30974]_  | ~\new_[5993]_ );
  assign \new_[28797]_  = ~\new_[29910]_  & ~\new_[30127]_ ;
  assign \new_[28798]_  = ~\new_[29891]_  | ~\new_[30644]_ ;
  assign \new_[28799]_  = ~\new_[30051]_  & ~\new_[30774]_ ;
  assign \new_[28800]_  = ~\new_[30771]_  & ~\new_[29537]_ ;
  assign \new_[28801]_  = ~\new_[30721]_ ;
  assign \new_[28802]_  = ~\new_[29870]_  | ~\new_[30070]_ ;
  assign \new_[28803]_  = ~\new_[30102]_  & ~\new_[30415]_ ;
  assign \new_[28804]_  = ~\new_[30360]_  | ~\new_[6084]_ ;
  assign \new_[28805]_  = ~\new_[29849]_  | ~\new_[31140]_ ;
  assign \new_[28806]_  = ~\new_[29750]_ ;
  assign \new_[28807]_  = ~\new_[30786]_  | ~\new_[6270]_ ;
  assign \new_[28808]_  = ~\new_[30080]_  | ~\new_[30159]_ ;
  assign \new_[28809]_  = ~\new_[30058]_  | ~\new_[5904]_ ;
  assign \new_[28810]_  = ~\new_[30197]_  | ~\new_[5914]_ ;
  assign \new_[28811]_  = ~\new_[30307]_  | ~\new_[29863]_ ;
  assign \new_[28812]_  = ~\new_[29760]_ ;
  assign \new_[28813]_  = ~\new_[30014]_  & ~\new_[30554]_ ;
  assign \new_[28814]_  = \new_[30347]_  | \new_[6040]_ ;
  assign \new_[28815]_  = \new_[30389]_  & \new_[30057]_ ;
  assign \new_[28816]_  = ~\new_[29435]_ ;
  assign \new_[28817]_  = ~\new_[30526]_  & ~\new_[30254]_ ;
  assign \new_[28818]_  = ~\new_[30328]_ ;
  assign \new_[28819]_  = ~\new_[30692]_  & ~\new_[31774]_ ;
  assign \new_[28820]_  = ~\new_[30845]_  & ~\new_[31645]_ ;
  assign \new_[28821]_  = ~\new_[31232]_  & ~\new_[31429]_ ;
  assign \new_[28822]_  = ~\new_[30428]_  & ~\new_[5999]_ ;
  assign \new_[28823]_  = (~\new_[31497]_  | ~\new_[5896]_ ) & (~\new_[30986]_  | ~\new_[5967]_ );
  assign \new_[28824]_  = ~\new_[30774]_ ;
  assign \new_[28825]_  = ~\new_[30710]_  | ~\new_[6072]_ ;
  assign \new_[28826]_  = ~\new_[30468]_  | ~n8464;
  assign \new_[28827]_  = \new_[30826]_  & \new_[31039]_ ;
  assign \new_[28828]_  = ~\new_[30087]_ ;
  assign \new_[28829]_  = ~\new_[30294]_ ;
  assign \new_[28830]_  = ~\new_[29768]_ ;
  assign \new_[28831]_  = \new_[30655]_  | \new_[31148]_ ;
  assign \new_[28832]_  = ~\new_[30803]_  & ~\new_[30850]_ ;
  assign \new_[28833]_  = ~\new_[30172]_ ;
  assign \new_[28834]_  = ~\new_[29771]_ ;
  assign \new_[28835]_  = ~\new_[30203]_ ;
  assign \new_[28836]_  = ~\new_[30236]_ ;
  assign \new_[28837]_  = ~\new_[29776]_ ;
  assign \new_[28838]_  = ~\new_[30737]_  | ~\new_[30789]_ ;
  assign \new_[28839]_  = ~\new_[30658]_  | ~n8649;
  assign \new_[28840]_  = ~\new_[30524]_  | ~\new_[4086]_ ;
  assign \new_[28841]_  = ~\new_[30565]_  | ~\new_[6094]_ ;
  assign \new_[28842]_  = \new_[30422]_  & \new_[31082]_ ;
  assign \new_[28843]_  = \new_[30634]_  & \new_[5981]_ ;
  assign \new_[28844]_  = ~\new_[30043]_ ;
  assign \new_[28845]_  = ~\new_[29784]_ ;
  assign \new_[28846]_  = ~\new_[30728]_ ;
  assign \new_[28847]_  = ~\new_[30764]_  | ~\new_[6217]_ ;
  assign \new_[28848]_  = ~\new_[29786]_ ;
  assign \new_[28849]_  = ~\new_[30432]_ ;
  assign \new_[28850]_  = ~\new_[29906]_ ;
  assign \new_[28851]_  = \new_[31155]_  & \new_[30712]_ ;
  assign \new_[28852]_  = ~\new_[30619]_  | ~n8604;
  assign \new_[28853]_  = ~\new_[30581]_  | ~\new_[6070]_ ;
  assign \new_[28854]_  = ~\new_[30435]_  & ~\new_[6001]_ ;
  assign \new_[28855]_  = ~\new_[30727]_  | ~\new_[6090]_ ;
  assign \new_[28856]_  = ~\new_[29787]_ ;
  assign \new_[28857]_  = ~\new_[29974]_ ;
  assign \new_[28858]_  = ~\new_[30474]_  | ~\new_[5983]_ ;
  assign \new_[28859]_  = ~\new_[30437]_ ;
  assign \new_[28860]_  = (~\new_[30944]_  | ~\new_[5982]_ ) & (~\new_[31487]_  | ~\new_[6065]_ );
  assign \new_[28861]_  = ~\new_[30468]_  | ~n8509;
  assign \new_[28862]_  = ~\new_[6036]_  | ~\new_[5895]_ ;
  assign \new_[28863]_  = ~\new_[30154]_ ;
  assign \new_[28864]_  = ~\new_[30307]_ ;
  assign \new_[28865]_  = ~\new_[30779]_  | ~\new_[4123]_ ;
  assign \new_[28866]_  = ~\new_[30503]_  | ~\new_[4056]_ ;
  assign \new_[28867]_  = ~\new_[30723]_ ;
  assign \new_[28868]_  = ~\new_[30412]_ ;
  assign \new_[28869]_  = ~\new_[30408]_ ;
  assign \new_[28870]_  = ~\new_[30407]_ ;
  assign \new_[28871]_  = ~\new_[30545]_  & ~\new_[30521]_ ;
  assign \new_[28872]_  = ~\new_[30314]_ ;
  assign \new_[28873]_  = \new_[30739]_  & \new_[4151]_ ;
  assign \new_[28874]_  = \new_[30624]_  | \new_[31788]_ ;
  assign \new_[28875]_  = ~\new_[30773]_  | ~\new_[30976]_ ;
  assign \new_[28876]_  = ~\new_[30356]_ ;
  assign \new_[28877]_  = ~\new_[30705]_  | ~\new_[4126]_ ;
  assign \new_[28878]_  = ~\new_[30450]_  | ~\new_[4253]_ ;
  assign \new_[28879]_  = ~\new_[30836]_  & ~\new_[6031]_ ;
  assign \new_[28880]_  = ~\new_[29827]_ ;
  assign \new_[28881]_  = ~\new_[29903]_ ;
  assign \new_[28882]_  = ~\new_[6074]_  | ~\new_[5904]_ ;
  assign \new_[28883]_  = ~\new_[29814]_ ;
  assign \new_[28884]_  = ~\new_[29817]_ ;
  assign \new_[28885]_  = ~\new_[29816]_ ;
  assign \new_[28886]_  = ~\new_[30479]_  | ~n8329;
  assign \new_[28887]_  = ~\new_[30141]_ ;
  assign \new_[28888]_  = \new_[30716]_  | \new_[4135]_ ;
  assign \new_[28889]_  = ~\new_[30790]_  | ~\new_[4442]_ ;
  assign \new_[28890]_  = ~\new_[29824]_ ;
  assign \new_[28891]_  = ~\new_[29825]_ ;
  assign \new_[28892]_  = ~\new_[30611]_  | ~n8609;
  assign \new_[28893]_  = ~\new_[30147]_ ;
  assign \new_[28894]_  = ~\new_[29826]_ ;
  assign \new_[28895]_  = ~\new_[30110]_ ;
  assign \new_[28896]_  = ~\new_[6045]_  | ~\new_[5897]_ ;
  assign \new_[28897]_  = ~\new_[30843]_  & ~\new_[31165]_ ;
  assign \new_[28898]_  = ~\new_[30339]_ ;
  assign \new_[28899]_  = ~\new_[30312]_ ;
  assign \new_[28900]_  = \new_[6186]_  & \new_[5928]_ ;
  assign \new_[28901]_  = ~\new_[30567]_  & ~\new_[31855]_ ;
  assign \new_[28902]_  = ~\new_[30533]_  | ~n8904;
  assign \new_[28903]_  = ~\new_[30353]_ ;
  assign \new_[28904]_  = ~\new_[30789]_ ;
  assign \new_[28905]_  = ~\new_[29830]_ ;
  assign \new_[28906]_  = ~\new_[30619]_  | ~n8939;
  assign \new_[28907]_  = ~\new_[30371]_ ;
  assign \new_[28908]_  = ~\new_[29839]_ ;
  assign \new_[28909]_  = ~\new_[29831]_ ;
  assign \new_[28910]_  = ~\new_[30529]_  & ~\new_[30874]_ ;
  assign \new_[28911]_  = ~\new_[29833]_ ;
  assign \new_[28912]_  = ~\new_[30100]_ ;
  assign \new_[28913]_  = ~\new_[30714]_  | ~\new_[6096]_ ;
  assign \new_[28914]_  = ~\new_[30479]_  | ~n8839;
  assign \new_[28915]_  = ~\new_[29843]_ ;
  assign \new_[28916]_  = ~\new_[30479]_  | ~n8804;
  assign \new_[28917]_  = ~\new_[29845]_ ;
  assign \new_[28918]_  = ~\new_[29848]_ ;
  assign \new_[28919]_  = ~\new_[29850]_ ;
  assign \new_[28920]_  = ~\new_[30473]_  | ~\new_[31494]_ ;
  assign \new_[28921]_  = ~\new_[30690]_  | ~n8789;
  assign \new_[28922]_  = ~\new_[30622]_  | ~\new_[6096]_ ;
  assign \new_[28923]_  = ~\new_[30654]_  | ~n8404;
  assign \new_[28924]_  = ~\new_[30076]_ ;
  assign \new_[28925]_  = ~\new_[30800]_  | ~\new_[30925]_ ;
  assign \new_[28926]_  = ~\new_[30400]_ ;
  assign \new_[28927]_  = ~\new_[30631]_  | ~n8354;
  assign \new_[28928]_  = ~\new_[30619]_  | ~n8719;
  assign \new_[28929]_  = ~\new_[29856]_ ;
  assign \new_[28930]_  = ~\new_[30801]_  | ~\new_[4142]_ ;
  assign \new_[28931]_  = ~\new_[29858]_ ;
  assign \new_[28932]_  = \new_[30838]_  & \new_[5994]_ ;
  assign \new_[28933]_  = ~\new_[30150]_ ;
  assign \new_[28934]_  = ~\new_[30067]_ ;
  assign \new_[28935]_  = \new_[30427]_  | \new_[31299]_ ;
  assign \new_[28936]_  = \new_[30418]_  | \new_[30894]_ ;
  assign \new_[28937]_  = ~\new_[30658]_  | ~n8704;
  assign \new_[28938]_  = ~\new_[30567]_  & ~\new_[6007]_ ;
  assign \new_[28939]_  = ~\new_[30052]_ ;
  assign \new_[28940]_  = ~\new_[30581]_  | ~\new_[6069]_ ;
  assign \new_[28941]_  = ~\new_[31491]_  | ~\new_[31471]_ ;
  assign \new_[28942]_  = ~\new_[30627]_  | ~\new_[30615]_ ;
  assign \new_[28943]_  = ~\new_[30479]_  | ~n8434;
  assign \new_[28944]_  = ~\new_[30583]_  & ~\new_[3882]_ ;
  assign \new_[28945]_  = ~\new_[30611]_  | ~n8739;
  assign \new_[28946]_  = ~\new_[30347]_ ;
  assign \new_[28947]_  = ~\new_[30690]_  | ~n8674;
  assign \new_[28948]_  = ~\new_[29871]_ ;
  assign \new_[28949]_  = ~\new_[6006]_  & ~\new_[6005]_ ;
  assign \new_[28950]_  = ~\new_[30196]_ ;
  assign \new_[28951]_  = \new_[30668]_  & \new_[5919]_ ;
  assign \new_[28952]_  = ~\new_[31685]_  & ~\new_[31588]_ ;
  assign \new_[28953]_  = ~\new_[30726]_ ;
  assign \new_[28954]_  = ~\new_[30654]_  | ~n8614;
  assign \new_[28955]_  = ~\new_[30658]_  | ~n8534;
  assign \new_[28956]_  = ~\new_[30703]_  | ~\new_[6061]_ ;
  assign \new_[28957]_  = \new_[30422]_  & \new_[30947]_ ;
  assign \new_[28958]_  = ~\new_[29895]_ ;
  assign \new_[28959]_  = ~\new_[30584]_  & ~\new_[31855]_ ;
  assign \new_[28960]_  = ~\new_[29891]_ ;
  assign \new_[28961]_  = ~\new_[30919]_  & ~\new_[31844]_ ;
  assign \new_[28962]_  = ~\new_[30234]_ ;
  assign \new_[28963]_  = ~\new_[30319]_ ;
  assign \new_[28964]_  = ~\new_[30032]_ ;
  assign \new_[28965]_  = ~\new_[30468]_  | ~n8634;
  assign \new_[28966]_  = ~\new_[30246]_ ;
  assign \new_[28967]_  = ~\new_[30209]_ ;
  assign \new_[28968]_  = ~\new_[29899]_ ;
  assign \new_[28969]_  = ~\new_[30475]_  | ~\new_[4072]_ ;
  assign \new_[28970]_  = \new_[30520]_  & \new_[31416]_ ;
  assign \new_[28971]_  = \new_[30768]_  & \new_[31844]_ ;
  assign \new_[28972]_  = ~\new_[30392]_ ;
  assign \new_[28973]_  = ~\new_[30448]_  | ~\new_[5924]_ ;
  assign \new_[28974]_  = ~\m7_addr_i[29]  & ~\m7_addr_i[28] ;
  assign \new_[28975]_  = ~\new_[30534]_  | ~\new_[5983]_ ;
  assign \new_[28976]_  = (~\new_[31216]_  | ~\new_[5895]_ ) & (~\new_[31008]_  | ~\new_[5910]_ );
  assign \new_[28977]_  = ~\new_[29893]_ ;
  assign \new_[28978]_  = ~\new_[30526]_  & ~\new_[30782]_ ;
  assign \new_[28979]_  = ~\new_[29904]_ ;
  assign \new_[28980]_  = \new_[30547]_  & \new_[6059]_ ;
  assign \new_[28981]_  = ~\new_[30750]_ ;
  assign \new_[28982]_  = ~\new_[29943]_ ;
  assign \new_[28983]_  = \new_[30527]_  | \new_[31763]_ ;
  assign \new_[28984]_  = ~\new_[29913]_ ;
  assign \new_[28985]_  = ~\new_[30059]_ ;
  assign \new_[28986]_  = ~\new_[30576]_  & ~\new_[5931]_ ;
  assign \new_[28987]_  = ~\new_[29835]_ ;
  assign \new_[28988]_  = ~\new_[30724]_ ;
  assign \new_[28989]_  = ~\new_[30168]_ ;
  assign \new_[28990]_  = ~\new_[30264]_ ;
  assign \new_[28991]_  = \new_[30495]_  | \new_[30897]_ ;
  assign \new_[28992]_  = ~\new_[29924]_ ;
  assign \new_[28993]_  = ~\new_[29919]_ ;
  assign \new_[28994]_  = ~\new_[30551]_  | ~\new_[5911]_ ;
  assign \new_[28995]_  = ~\new_[29925]_ ;
  assign \new_[28996]_  = ~\new_[30431]_  | ~\new_[5978]_ ;
  assign \new_[28997]_  = ~\new_[30175]_ ;
  assign \new_[28998]_  = ~\new_[30333]_ ;
  assign \new_[28999]_  = \new_[30455]_  & \new_[4449]_ ;
  assign \new_[29000]_  = \new_[30500]_  & \new_[6176]_ ;
  assign \new_[29001]_  = ~\new_[30819]_  & ~\new_[30851]_ ;
  assign \new_[29002]_  = ~\new_[30654]_  | ~n8714;
  assign \new_[29003]_  = ~\new_[30004]_ ;
  assign \new_[29004]_  = ~\new_[31398]_  & ~\m2_addr_i[29] ;
  assign \new_[29005]_  = ~\new_[30194]_ ;
  assign \new_[29006]_  = ~\new_[29934]_ ;
  assign \new_[29007]_  = ~\new_[29860]_ ;
  assign \new_[29008]_  = ~\new_[29931]_ ;
  assign \new_[29009]_  = ~\new_[30764]_  | ~\new_[30820]_ ;
  assign \new_[29010]_  = ~\new_[30819]_  & ~\new_[30839]_ ;
  assign \new_[29011]_  = \new_[30826]_  & \new_[6031]_ ;
  assign \new_[29012]_  = \new_[30674]_  & \new_[31206]_ ;
  assign \new_[29013]_  = ~\new_[29922]_ ;
  assign \new_[29014]_  = ~\new_[29859]_ ;
  assign \new_[29015]_  = ~\new_[30247]_ ;
  assign \new_[29016]_  = ~\new_[30730]_ ;
  assign \new_[29017]_  = ~\new_[30073]_ ;
  assign \new_[29018]_  = ~\new_[30468]_  | ~n8384;
  assign \new_[29019]_  = ~\new_[30766]_  & ~\new_[31412]_ ;
  assign \new_[29020]_  = ~\new_[30206]_ ;
  assign \new_[29021]_  = \new_[30806]_  & \new_[31059]_ ;
  assign \new_[29022]_  = (~\new_[6185]_  | ~\new_[31119]_ ) & (~\new_[6086]_  | ~\new_[31221]_ );
  assign \new_[29023]_  = ~\new_[30654]_  | ~n8539;
  assign \new_[29024]_  = \new_[30816]_  & \new_[31145]_ ;
  assign \new_[29025]_  = ~\new_[30685]_  & ~\new_[30985]_ ;
  assign \new_[29026]_  = ~\new_[30420]_  | ~\new_[30508]_ ;
  assign \new_[29027]_  = ~\new_[30588]_  | ~\new_[5909]_ ;
  assign \new_[29028]_  = ~\new_[29992]_ ;
  assign \new_[29029]_  = ~\new_[30528]_  | ~\new_[4206]_ ;
  assign \new_[29030]_  = ~\new_[30720]_  | ~\new_[31648]_ ;
  assign \new_[29031]_  = ~\new_[30912]_  & ~\new_[6071]_ ;
  assign \new_[29032]_  = ~\new_[29952]_ ;
  assign \new_[29033]_  = ~\new_[29942]_ ;
  assign \new_[29034]_  = \new_[31152]_  & \new_[30536]_ ;
  assign \new_[29035]_  = \new_[30869]_  & \new_[30536]_ ;
  assign \new_[29036]_  = \new_[31065]_  & \new_[30744]_ ;
  assign \new_[29037]_  = ~\new_[30619]_  | ~n8849;
  assign \new_[29038]_  = ~\new_[29955]_ ;
  assign \new_[29039]_  = ~\new_[6194]_  & ~\new_[5984]_ ;
  assign \new_[29040]_  = ~\new_[29985]_ ;
  assign \new_[29041]_  = \new_[30866]_  & \new_[30851]_ ;
  assign \new_[29042]_  = ~\new_[29946]_ ;
  assign \new_[29043]_  = ~\new_[31138]_  & ~\new_[30823]_ ;
  assign \new_[29044]_  = ~\new_[30785]_  | ~\new_[6096]_ ;
  assign \new_[29045]_  = \new_[30506]_  & \new_[30818]_ ;
  assign \new_[29046]_  = ~\new_[31253]_  & ~\m4_addr_i[29] ;
  assign \new_[29047]_  = ~\new_[30054]_ ;
  assign \new_[29048]_  = ~\new_[30479]_  | ~n8869;
  assign \new_[29049]_  = ~\new_[30834]_  | ~\new_[5918]_ ;
  assign \new_[29050]_  = ~\new_[30348]_ ;
  assign \new_[29051]_  = ~\new_[30502]_  & ~\new_[30723]_ ;
  assign \new_[29052]_  = \new_[31082]_  & \new_[30802]_ ;
  assign \new_[29053]_  = ~\new_[31274]_  & ~\m6_addr_i[29] ;
  assign \new_[29054]_  = ~\new_[30220]_ ;
  assign \new_[29055]_  = ~\new_[30419]_  & ~\new_[4218]_ ;
  assign \new_[29056]_  = ~\new_[30159]_ ;
  assign \new_[29057]_  = ~\new_[30622]_  | ~\new_[31433]_ ;
  assign \new_[29058]_  = ~\new_[30094]_ ;
  assign \new_[29059]_  = ~\new_[30953]_  & ~\new_[6064]_ ;
  assign \new_[29060]_  = ~\new_[30449]_  | ~\new_[5917]_ ;
  assign \new_[29061]_  = ~\new_[30118]_ ;
  assign \new_[29062]_  = ~\new_[29984]_ ;
  assign \new_[29063]_  = ~\new_[6194]_  | ~\new_[5984]_ ;
  assign \new_[29064]_  = \new_[30716]_  | \new_[31417]_ ;
  assign \new_[29065]_  = ~\new_[30658]_  | ~n8564;
  assign \new_[29066]_  = ~\new_[30772]_  & ~\new_[5914]_ ;
  assign \new_[29067]_  = ~\new_[6042]_  | ~\new_[5896]_ ;
  assign \new_[29068]_  = ~\new_[30061]_ ;
  assign \new_[29069]_  = ~\new_[29977]_ ;
  assign \new_[29070]_  = (~\new_[5924]_  | ~\new_[31072]_ ) & (~\new_[5994]_  | ~\new_[30974]_ );
  assign \new_[29071]_  = ~\new_[30048]_ ;
  assign \new_[29072]_  = ~\new_[30654]_  | ~n8834;
  assign \new_[29073]_  = ~\new_[30734]_  & ~\new_[6072]_ ;
  assign \new_[29074]_  = ~\new_[30760]_  & ~\new_[31042]_ ;
  assign \new_[29075]_  = ~\new_[30611]_  | ~n8399;
  assign \new_[29076]_  = ~\new_[30480]_  | ~\new_[31340]_ ;
  assign \new_[29077]_  = ~\new_[30572]_ ;
  assign \new_[29078]_  = ~\new_[30440]_  & ~\new_[31259]_ ;
  assign \new_[29079]_  = ~\new_[30465]_  | ~\new_[4220]_ ;
  assign \new_[29080]_  = ~\new_[30533]_  | ~n8559;
  assign \new_[29081]_  = ~\new_[30533]_  | ~n8929;
  assign \new_[29082]_  = ~\new_[30302]_ ;
  assign \new_[29083]_  = ~\new_[30654]_  | ~n8314;
  assign \new_[29084]_  = ~\new_[30657]_  & ~\new_[31844]_ ;
  assign \new_[29085]_  = \new_[30671]_  & \new_[31787]_ ;
  assign \new_[29086]_  = ~\new_[30808]_  | ~\new_[4137]_ ;
  assign \new_[29087]_  = ~\new_[29993]_ ;
  assign \new_[29088]_  = ~\new_[30288]_ ;
  assign \new_[29089]_  = ~\new_[30005]_ ;
  assign \new_[29090]_  = ~\new_[30424]_  & ~\new_[6033]_ ;
  assign \new_[29091]_  = ~\new_[30673]_  & ~\new_[30993]_ ;
  assign \new_[29092]_  = ~\new_[30281]_ ;
  assign \new_[29093]_  = ~\new_[30690]_  | ~n8424;
  assign \new_[29094]_  = ~\new_[30658]_  | ~n8679;
  assign \new_[29095]_  = ~\new_[30027]_ ;
  assign \new_[29096]_  = ~\new_[30046]_ ;
  assign \new_[29097]_  = ~\new_[30654]_  | ~n8469;
  assign \new_[29098]_  = ~\new_[30501]_  | ~\new_[30786]_ ;
  assign \new_[29099]_  = ~\new_[6083]_  | ~\new_[5906]_ ;
  assign \new_[29100]_  = ~\new_[30079]_ ;
  assign \new_[29101]_  = ~\new_[29881]_ ;
  assign \new_[29102]_  = ~\new_[30330]_ ;
  assign \new_[29103]_  = ~\new_[30249]_ ;
  assign \new_[29104]_  = ~\new_[30355]_ ;
  assign \new_[29105]_  = (~\new_[6006]_  | ~\new_[30936]_ ) & (~\new_[6095]_  | ~\new_[31303]_ );
  assign \new_[29106]_  = \new_[30758]_  & \new_[6071]_ ;
  assign \new_[29107]_  = ~\new_[30658]_  | ~n8624;
  assign \new_[29108]_  = (~\new_[6047]_  | ~\new_[31211]_ ) & (~\new_[6200]_  | ~\new_[31337]_ );
  assign \new_[29109]_  = ~\new_[30690]_  | ~n8484;
  assign \new_[29110]_  = \new_[30829]_  & \new_[31042]_ ;
  assign \new_[29111]_  = ~\new_[30533]_  | ~n8684;
  assign \new_[29112]_  = ~\new_[30040]_ ;
  assign \new_[29113]_  = ~\new_[30841]_  & ~\new_[31754]_ ;
  assign \new_[29114]_  = ~\new_[30668]_  | ~\new_[30874]_ ;
  assign \new_[29115]_  = ~\new_[30381]_ ;
  assign \new_[29116]_  = ~\new_[30654]_  | ~n8824;
  assign \new_[29117]_  = ~\new_[30446]_  | ~\new_[6048]_ ;
  assign \new_[29118]_  = ~\new_[30276]_ ;
  assign \new_[29119]_  = ~\new_[30019]_ ;
  assign \new_[29120]_  = (~\new_[6080]_  | ~\new_[31543]_ ) & (~\new_[6079]_  | ~\new_[30908]_ );
  assign \new_[29121]_  = ~\new_[30602]_  & ~\new_[30850]_ ;
  assign \new_[29122]_  = ~\new_[30022]_ ;
  assign \new_[29123]_  = ~\new_[30648]_  & ~\new_[30550]_ ;
  assign \new_[29124]_  = ~\new_[30642]_  | ~\new_[6215]_ ;
  assign \new_[29125]_  = ~\new_[30517]_  | ~\new_[5924]_ ;
  assign \new_[29126]_  = ~\new_[30773]_  | ~\new_[6033]_ ;
  assign \new_[29127]_  = (~\new_[5926]_  | ~\new_[31543]_ ) & (~\new_[6078]_  | ~\new_[30908]_ );
  assign \new_[29128]_  = ~\new_[30842]_  | ~\new_[6192]_ ;
  assign \new_[29129]_  = (~\new_[6058]_  | ~\new_[30989]_ ) & (~\new_[6195]_  | ~\new_[31452]_ );
  assign \new_[29130]_  = ~\new_[29960]_ ;
  assign \new_[29131]_  = \new_[30461]_  & \new_[6059]_ ;
  assign \new_[29132]_  = ~\new_[30083]_ ;
  assign \new_[29133]_  = ~\new_[30654]_  | ~n8769;
  assign \new_[29134]_  = ~\new_[31491]_  | ~\new_[5916]_ ;
  assign \new_[29135]_  = ~\new_[30761]_  | ~\new_[31763]_ ;
  assign \new_[29136]_  = ~\new_[30677]_  | ~\new_[6078]_ ;
  assign \new_[29137]_  = ~\new_[30561]_  | ~\new_[5912]_ ;
  assign \new_[29138]_  = \new_[30646]_  | \new_[31648]_ ;
  assign \new_[29139]_  = ~\new_[30074]_ ;
  assign \new_[29140]_  = ~\new_[30523]_  & ~\new_[5981]_ ;
  assign \new_[29141]_  = ~\new_[30611]_  | ~n8359;
  assign \new_[29142]_  = \new_[31685]_  | \new_[30477]_ ;
  assign \new_[29143]_  = \new_[30815]_  & \new_[31108]_ ;
  assign \new_[29144]_  = ~\new_[30783]_  & ~\new_[5996]_ ;
  assign \new_[29145]_  = ~\new_[30239]_ ;
  assign \new_[29146]_  = \new_[30768]_  & \new_[5968]_ ;
  assign \new_[29147]_  = ~\new_[30539]_  | ~\new_[5983]_ ;
  assign \new_[29148]_  = ~\new_[30155]_ ;
  assign \new_[29149]_  = \new_[30745]_  & \new_[31065]_ ;
  assign \new_[29150]_  = ~\new_[30522]_  | ~\new_[4089]_ ;
  assign \new_[29151]_  = ~\new_[30072]_ ;
  assign \new_[29152]_  = ~\new_[30300]_ ;
  assign \new_[29153]_  = \new_[30485]_  & n8309;
  assign \new_[29154]_  = ~\new_[30045]_ ;
  assign \new_[29155]_  = \new_[30824]_  & \new_[31855]_ ;
  assign \new_[29156]_  = ~\new_[30727]_  | ~\new_[30507]_ ;
  assign \new_[29157]_  = ~\new_[29941]_ ;
  assign \new_[29158]_  = ~\new_[30425]_  & ~\new_[31617]_ ;
  assign \new_[29159]_  = ~\new_[30509]_  | ~\new_[4231]_ ;
  assign \new_[29160]_  = ~\new_[31163]_  & ~\new_[6212]_ ;
  assign \new_[29161]_  = \new_[30825]_  & \new_[5913]_ ;
  assign \new_[29162]_  = ~\new_[30666]_  | ~\new_[4121]_ ;
  assign \new_[29163]_  = ~\new_[30533]_  | ~n8414;
  assign \new_[29164]_  = ~\new_[30479]_  | ~n8374;
  assign \new_[29165]_  = ~\new_[30138]_ ;
  assign \new_[29166]_  = ~\new_[30161]_ ;
  assign \new_[29167]_  = ~\new_[30317]_ ;
  assign \new_[29168]_  = ~\new_[30464]_  | ~\new_[4098]_ ;
  assign \new_[29169]_  = ~\new_[29868]_ ;
  assign \new_[29170]_  = \new_[30776]_  & \new_[6206]_ ;
  assign \new_[29171]_  = ~\new_[30532]_  | ~\new_[4132]_ ;
  assign \new_[29172]_  = ~\new_[29873]_ ;
  assign \new_[29173]_  = (~\new_[5909]_  | ~\new_[31216]_ ) & (~\new_[6040]_  | ~\new_[31008]_ );
  assign \new_[29174]_  = ~\new_[30035]_ ;
  assign \new_[29175]_  = ~\new_[30452]_  | ~\new_[4237]_ ;
  assign \new_[29176]_  = \new_[30556]_  & \new_[6270]_ ;
  assign \new_[29177]_  = (~\new_[5919]_  | ~\new_[31075]_ ) & (~\new_[6071]_  | ~\new_[31228]_ );
  assign \new_[29178]_  = ~\new_[30533]_  | ~n8754;
  assign \new_[29179]_  = \new_[30639]_  & \new_[5964]_ ;
  assign \new_[29180]_  = (~\new_[5999]_  | ~\new_[31119]_ ) & (~\new_[6001]_  | ~\new_[31221]_ );
  assign \new_[29181]_  = ~\new_[29929]_ ;
  assign \new_[29182]_  = ~\new_[30600]_  | ~\new_[6214]_ ;
  assign \new_[29183]_  = \new_[30550]_  & \new_[6046]_ ;
  assign \new_[29184]_  = ~\new_[30269]_ ;
  assign \new_[29185]_  = \new_[30674]_  & \new_[31155]_ ;
  assign \new_[29186]_  = ~\new_[30804]_  | ~\new_[4084]_ ;
  assign \new_[29187]_  = ~\new_[31167]_  & ~\new_[5919]_ ;
  assign \new_[29188]_  = \new_[30643]_  & \new_[5999]_ ;
  assign \new_[29189]_  = ~\new_[30080]_ ;
  assign \new_[29190]_  = ~\new_[30533]_  | ~n8389;
  assign \new_[29191]_  = ~\new_[6197]_  | ~\new_[6057]_ ;
  assign \new_[29192]_  = ~\new_[30659]_  | ~\new_[4061]_ ;
  assign \new_[29193]_  = ~\new_[30417]_  & ~\new_[6071]_ ;
  assign \new_[29194]_  = \new_[30560]_  & \new_[6176]_ ;
  assign \new_[29195]_  = ~\new_[30097]_ ;
  assign \new_[29196]_  = ~\new_[30822]_  & ~\new_[5917]_ ;
  assign \new_[29197]_  = ~\new_[30687]_  | ~\new_[3879]_ ;
  assign \new_[29198]_  = ~\new_[30533]_  | ~n8794;
  assign \new_[29199]_  = ~\new_[30550]_ ;
  assign \new_[29200]_  = \new_[30781]_  | \new_[5924]_ ;
  assign \new_[29201]_  = (~\new_[31055]_  | ~\new_[5986]_ ) & (~\new_[31518]_  | ~\new_[5987]_ );
  assign \new_[29202]_  = ~\new_[29940]_ ;
  assign \new_[29203]_  = ~\new_[30619]_  | ~n8854;
  assign \new_[29204]_  = \new_[30824]_  & \new_[6007]_ ;
  assign \new_[29205]_  = \new_[30756]_  & \new_[30536]_ ;
  assign \new_[29206]_  = ~\new_[30497]_  | ~\new_[30774]_ ;
  assign \new_[29207]_  = ~\new_[30533]_  | ~n8494;
  assign \new_[29208]_  = (~\new_[30937]_  | ~\new_[5963]_ ) & (~\new_[31328]_  | ~\new_[6245]_ );
  assign \new_[29209]_  = ~\new_[30710]_  | ~\new_[5989]_ ;
  assign \new_[29210]_  = ~\new_[30244]_ ;
  assign \new_[29211]_  = ~\new_[30736]_  & ~\new_[30582]_ ;
  assign \new_[29212]_  = ~\new_[30270]_ ;
  assign \new_[29213]_  = ~\new_[30479]_  | ~n8344;
  assign \new_[29214]_  = (~\new_[5911]_  | ~\new_[31497]_ ) & (~\new_[6032]_  | ~\new_[30986]_ );
  assign \new_[29215]_  = \new_[30999]_  & \new_[30536]_ ;
  assign \new_[29216]_  = ~\new_[30690]_  | ~n8524;
  assign \new_[29217]_  = ~\new_[30282]_ ;
  assign \new_[29218]_  = \new_[30655]_  | \new_[31539]_ ;
  assign \new_[29219]_  = ~\new_[30095]_ ;
  assign \new_[29220]_  = ~\new_[29966]_ ;
  assign \new_[29221]_  = ~\new_[30301]_ ;
  assign \new_[29222]_  = ~\new_[30279]_ ;
  assign \new_[29223]_  = ~\new_[29981]_ ;
  assign \new_[29224]_  = (~\new_[6081]_  | ~\new_[30930]_ ) & (~\new_[6082]_  | ~\new_[31473]_ );
  assign \new_[29225]_  = ~\new_[30240]_ ;
  assign \new_[29226]_  = ~\new_[30305]_ ;
  assign \new_[29227]_  = ~\new_[30092]_ ;
  assign \new_[29228]_  = ~\new_[30192]_ ;
  assign \new_[29229]_  = ~\new_[30211]_ ;
  assign \new_[29230]_  = (~\new_[5932]_  | ~\new_[30936]_ ) & (~\new_[6007]_  | ~\new_[31303]_ );
  assign \new_[29231]_  = ~\new_[30619]_  | ~n8819;
  assign \new_[29232]_  = \new_[30605]_  | \new_[6204]_ ;
  assign \new_[29233]_  = ~\new_[30323]_ ;
  assign \new_[29234]_  = ~\new_[30690]_  | ~n8599;
  assign \new_[29235]_  = ~\new_[30114]_ ;
  assign \new_[29236]_  = \new_[30459]_  | \new_[6078]_ ;
  assign \new_[29237]_  = ~\new_[30498]_  & ~\new_[5979]_ ;
  assign \new_[29238]_  = ~\new_[30692]_  & ~\new_[4158]_ ;
  assign \new_[29239]_  = ~\new_[30611]_  | ~n8749;
  assign \new_[29240]_  = ~\new_[30533]_  | ~n8709;
  assign \new_[29241]_  = \new_[31152]_  & \new_[30827]_ ;
  assign \new_[29242]_  = (~\new_[30970]_  | ~\new_[5990]_ ) & (~\new_[31437]_  | ~\new_[5922]_ );
  assign \new_[29243]_  = ~\new_[30621]_  | ~\new_[31259]_ ;
  assign \new_[29244]_  = ~\new_[30728]_  | ~\new_[6208]_ ;
  assign \new_[29245]_  = ~\new_[30468]_  | ~n8334;
  assign \new_[29246]_  = ~\new_[31394]_  & ~\new_[31345]_ ;
  assign \new_[29247]_  = ~\new_[29980]_ ;
  assign \new_[29248]_  = ~\new_[30127]_ ;
  assign \new_[29249]_  = ~\new_[30718]_  | ~\new_[30615]_ ;
  assign \new_[29250]_  = ~\new_[30594]_  | ~\new_[31455]_ ;
  assign \new_[29251]_  = \new_[30530]_  | \new_[4070]_ ;
  assign \new_[29252]_  = ~\new_[30658]_  | ~n8544;
  assign \new_[29253]_  = ~\new_[30690]_  | ~n8934;
  assign \new_[29254]_  = ~\new_[30258]_ ;
  assign \new_[29255]_  = (~\new_[31136]_  | ~\new_[6088]_ ) & (~\new_[31263]_  | ~\new_[6090]_ );
  assign \new_[29256]_  = \new_[30797]_  & \new_[4107]_ ;
  assign \new_[29257]_  = \new_[30740]_  & \new_[5979]_ ;
  assign \new_[29258]_  = \new_[30844]_  & \new_[30471]_ ;
  assign \new_[29259]_  = ~\new_[30468]_  | ~n8879;
  assign \new_[29260]_  = ~\new_[30404]_ ;
  assign \new_[29261]_  = ~\new_[30658]_  | ~n8774;
  assign \new_[29262]_  = ~\new_[29795]_ ;
  assign \new_[29263]_  = ~\new_[30533]_  | ~n8699;
  assign \new_[29264]_  = (~\new_[6062]_  | ~\new_[31317]_ ) & (~\new_[6063]_  | ~\new_[30944]_ );
  assign \new_[29265]_  = ~\new_[30433]_  & ~\new_[5994]_ ;
  assign \new_[29266]_  = ~\new_[30149]_ ;
  assign \new_[29267]_  = ~\new_[30690]_  | ~n8689;
  assign \new_[29268]_  = ~\new_[29882]_ ;
  assign \new_[29269]_  = ~\new_[30690]_  | ~n8489;
  assign \new_[29270]_  = ~\new_[30468]_  | ~n8884;
  assign \new_[29271]_  = ~\new_[29791]_ ;
  assign \new_[29272]_  = ~\new_[30158]_ ;
  assign \new_[29273]_  = ~\new_[31194]_  & ~\new_[5830]_ ;
  assign \new_[29274]_  = ~\new_[29958]_ ;
  assign \new_[29275]_  = ~\new_[30619]_  | ~n8309;
  assign \new_[29276]_  = ~\new_[30251]_ ;
  assign \new_[29277]_  = \new_[30606]_  & \new_[4451]_ ;
  assign \new_[29278]_  = ~\new_[30810]_  | ~\new_[6094]_ ;
  assign \new_[29279]_  = ~\new_[30748]_  & ~\new_[5985]_ ;
  assign \new_[29280]_  = ~\new_[30654]_  | ~n8474;
  assign \new_[29281]_  = (~\new_[5830]_  | ~\new_[30877]_ ) & (~\new_[6031]_  | ~\new_[31434]_ );
  assign \new_[29282]_  = ~\new_[30451]_  | ~\new_[5923]_ ;
  assign \new_[29283]_  = ~\new_[30418]_  & ~\new_[6069]_ ;
  assign \new_[29284]_  = ~\new_[30652]_  | ~\new_[30707]_ ;
  assign \new_[29285]_  = ~\new_[30654]_  | ~n8594;
  assign \new_[29286]_  = ~\new_[30526]_  & ~\new_[31777]_ ;
  assign \new_[29287]_  = ~\new_[30263]_ ;
  assign \new_[29288]_  = ~\new_[30611]_  | ~n8914;
  assign \new_[29289]_  = ~\new_[30713]_  | ~\new_[30444]_ ;
  assign \new_[29290]_  = \new_[30458]_  & \new_[4162]_ ;
  assign \new_[29291]_  = ~\new_[30214]_ ;
  assign \new_[29292]_  = \new_[30698]_  & \new_[5985]_ ;
  assign \new_[29293]_  = ~\new_[30316]_ ;
  assign \new_[29294]_  = ~\new_[30575]_  & ~\new_[30629]_ ;
  assign \new_[29295]_  = ~\new_[30690]_  | ~n8419;
  assign \new_[29296]_  = (~\new_[5979]_  | ~\new_[30989]_ ) & (~\new_[6059]_  | ~\new_[31452]_ );
  assign \new_[29297]_  = ~\new_[30514]_  | ~\new_[30998]_ ;
  assign \new_[29298]_  = \new_[30439]_  & \new_[31059]_ ;
  assign \new_[29299]_  = ~\new_[30739]_  | ~\new_[31012]_ ;
  assign \new_[29300]_  = \new_[30482]_  & \new_[4244]_ ;
  assign \new_[29301]_  = ~\new_[30787]_  & ~\new_[30848]_ ;
  assign \new_[29302]_  = ~\new_[30568]_  | ~\new_[6196]_ ;
  assign \new_[29303]_  = ~\new_[30558]_  | ~\new_[6069]_ ;
  assign \new_[29304]_  = ~\new_[30345]_ ;
  assign \new_[29305]_  = ~\new_[30769]_  & ~\new_[30785]_ ;
  assign \new_[29306]_  = ~\new_[30000]_ ;
  assign \new_[29307]_  = ~\new_[30611]_  | ~n8664;
  assign \new_[29308]_  = ~\new_[30611]_  | ~n8479;
  assign \new_[29309]_  = ~\new_[30468]_  | ~n8349;
  assign \new_[29310]_  = ~\new_[30783]_  & ~\new_[31108]_ ;
  assign \new_[29311]_  = ~\new_[30733]_  | ~\new_[30774]_ ;
  assign \new_[29312]_  = ~\new_[30658]_  | ~n8354;
  assign \new_[29313]_  = ~\new_[30831]_  | ~\new_[5924]_ ;
  assign \new_[29314]_  = ~\new_[30171]_ ;
  assign \new_[29315]_  = ~\new_[29783]_ ;
  assign \new_[29316]_  = ~\new_[30690]_  | ~n8894;
  assign \new_[29317]_  = \new_[30562]_  & \new_[30712]_ ;
  assign \new_[29318]_  = ~\new_[30540]_  | ~\new_[6034]_ ;
  assign \new_[29319]_  = ~\new_[30842]_  | ~\new_[30538]_ ;
  assign \new_[29320]_  = ~\new_[30334]_ ;
  assign \new_[29321]_  = \new_[31011]_  | \new_[5981]_ ;
  assign \new_[29322]_  = ~\new_[30703]_  | ~\new_[30897]_ ;
  assign \new_[29323]_  = ~\new_[30611]_  | ~n8449;
  assign \new_[29324]_  = \new_[30841]_  | \new_[4262]_ ;
  assign \new_[29325]_  = ~\new_[30753]_  | ~\new_[5921]_ ;
  assign \new_[29326]_  = ~\new_[30479]_  | ~n8809;
  assign \new_[29327]_  = ~\new_[30468]_  | ~n8844;
  assign \new_[29328]_  = ~\new_[30690]_  | ~n8909;
  assign \new_[29329]_  = (~\new_[5968]_  | ~\new_[30882]_ ) & (~\new_[6204]_  | ~\new_[31393]_ );
  assign \new_[29330]_  = ~\new_[30306]_ ;
  assign \new_[29331]_  = ~\new_[30163]_ ;
  assign \new_[29332]_  = ~\new_[30216]_ ;
  assign \new_[29333]_  = ~\new_[30123]_ ;
  assign \new_[29334]_  = ~\new_[30417]_  & ~\new_[31180]_ ;
  assign \new_[29335]_  = \new_[31923]_  | \new_[30570]_ ;
  assign \new_[29336]_  = ~\new_[30642]_  | ~\new_[6184]_ ;
  assign \new_[29337]_  = ~\new_[30428]_  & ~\new_[31140]_ ;
  assign \new_[29338]_  = ~\new_[30746]_  & ~\new_[30491]_ ;
  assign \new_[29339]_  = ~\new_[30090]_ ;
  assign \new_[29340]_  = ~\new_[30658]_  | ~n8409;
  assign \new_[29341]_  = ~\new_[30479]_  | ~n8369;
  assign \new_[29342]_  = ~\new_[30376]_ ;
  assign \new_[29343]_  = ~\new_[30838]_  | ~\new_[30851]_ ;
  assign \new_[29344]_  = ~\new_[30711]_  & ~\new_[30649]_ ;
  assign \new_[29345]_  = ~\new_[30602]_  & ~\new_[6212]_ ;
  assign \new_[29346]_  = \new_[30723]_  & \new_[5930]_ ;
  assign \new_[29347]_  = ~\new_[29763]_ ;
  assign \new_[29348]_  = \new_[30698]_  & \new_[30969]_ ;
  assign \new_[29349]_  = \new_[30562]_  & \new_[30997]_ ;
  assign \new_[29350]_  = ~\new_[30148]_ ;
  assign \new_[29351]_  = ~\new_[30443]_  & ~\new_[30597]_ ;
  assign \new_[29352]_  = ~\new_[30785]_  | ~\new_[5970]_ ;
  assign \new_[29353]_  = \new_[30664]_  & \new_[31104]_ ;
  assign \new_[29354]_  = ~\new_[30299]_ ;
  assign \new_[29355]_  = ~\new_[29773]_ ;
  assign \new_[29356]_  = (~\new_[5997]_  | ~\new_[30930]_ ) & (~\new_[6269]_  | ~\new_[31473]_ );
  assign \new_[29357]_  = ~\new_[30231]_ ;
  assign \new_[29358]_  = \new_[30832]_  & \new_[6190]_ ;
  assign \new_[29359]_  = ~\new_[29886]_ ;
  assign \new_[29360]_  = ~\new_[30530]_  & ~\new_[31446]_ ;
  assign \new_[29361]_  = ~\new_[30082]_ ;
  assign \new_[29362]_  = \new_[30740]_  & \new_[31014]_ ;
  assign \new_[29363]_  = ~\new_[30237]_ ;
  assign \new_[29364]_  = \new_[30803]_  | \new_[30848]_ ;
  assign \new_[29365]_  = ~\new_[30540]_  | ~\new_[6033]_ ;
  assign \new_[29366]_  = ~\new_[30649]_  | ~\new_[31712]_ ;
  assign \new_[29367]_  = ~\new_[29927]_ ;
  assign \new_[29368]_  = ~\new_[6193]_  | ~\new_[5903]_ ;
  assign \new_[29369]_  = ~\new_[30619]_  | ~n8639;
  assign \new_[29370]_  = ~\new_[29892]_ ;
  assign \new_[29371]_  = ~\new_[30344]_ ;
  assign \new_[29372]_  = ~\new_[30584]_  & ~\new_[30735]_ ;
  assign \new_[29373]_  = \new_[30643]_  & \new_[31140]_ ;
  assign \new_[29374]_  = ~\new_[6075]_  | ~\new_[5905]_ ;
  assign \new_[29375]_  = ~\new_[29967]_ ;
  assign \new_[29376]_  = ~\new_[30479]_  | ~n8619;
  assign \new_[29377]_  = ~\new_[30658]_  | ~n8579;
  assign \new_[29378]_  = ~\new_[30689]_  & ~\new_[31787]_ ;
  assign \new_[29379]_  = \new_[30520]_  & \new_[6001]_ ;
  assign \new_[29380]_  = \new_[30559]_  & \new_[6215]_ ;
  assign \new_[29381]_  = ~\new_[30460]_  | ~\new_[4074]_ ;
  assign \new_[29382]_  = ~\new_[30660]_  | ~\new_[5910]_ ;
  assign \new_[29383]_  = \new_[30535]_  & \new_[4043]_ ;
  assign \new_[29384]_  = ~\new_[30126]_ ;
  assign \new_[29385]_  = ~\new_[31265]_  & ~\new_[31292]_ ;
  assign \new_[29386]_  = ~\new_[30036]_ ;
  assign \new_[29387]_  = ~\new_[30741]_  & ~\new_[31787]_ ;
  assign \new_[29388]_  = (~\new_[5983]_  | ~\new_[31317]_ ) & (~\new_[6210]_  | ~\new_[31158]_ );
  assign \new_[29389]_  = (~\new_[6035]_  | ~\new_[30937]_ ) & (~\new_[6203]_  | ~\new_[31328]_ );
  assign \new_[29390]_  = ~\new_[30501]_  & ~\new_[30677]_ ;
  assign \new_[29391]_  = ~\new_[30611]_  | ~n8454;
  assign \new_[29392]_  = (~\new_[5972]_  | ~\new_[30877]_ ) & (~\new_[6052]_  | ~\new_[31434]_ );
  assign \new_[29393]_  = (~\new_[6056]_  | ~\new_[31468]_ ) & (~\new_[6197]_  | ~\new_[31050]_ );
  assign \new_[29394]_  = ~\new_[30320]_ ;
  assign \new_[29395]_  = ~\new_[30654]_  | ~n8569;
  assign \new_[29396]_  = \new_[6186]_  | \new_[5928]_ ;
  assign \new_[29397]_  = ~\new_[30266]_ ;
  assign \new_[29398]_  = ~\new_[30084]_ ;
  assign \new_[29399]_  = ~\new_[30591]_  | ~\new_[6084]_ ;
  assign \new_[29400]_  = (~\new_[6077]_  | ~\new_[30974]_ ) & (~\new_[6268]_  | ~\new_[31339]_ );
  assign \new_[29401]_  = ~\new_[30204]_ ;
  assign \new_[29402]_  = (~\new_[31220]_  | ~\new_[5904]_ ) & (~\new_[30973]_  | ~\new_[5989]_ );
  assign \new_[29403]_  = (~\new_[30930]_  | ~\new_[5998]_ ) & (~\new_[31473]_  | ~\new_[6085]_ );
  assign \new_[29404]_  = ~\new_[30176]_ ;
  assign \new_[29405]_  = (~\new_[31075]_  | ~\new_[5920]_ ) & (~\new_[31228]_  | ~\new_[6192]_ );
  assign \new_[29406]_  = (~\new_[6202]_  | ~\new_[31495]_ ) & (~\new_[6174]_  | ~\new_[30978]_ );
  assign \new_[29407]_  = \new_[30734]_  | \new_[31455]_ ;
  assign \new_[29408]_  = (~\new_[5985]_  | ~\new_[31055]_ ) & (~\new_[6212]_  | ~\new_[31518]_ );
  assign \new_[29409]_  = ~\new_[30468]_  | ~n8589;
  assign \new_[29410]_  = ~\new_[30308]_ ;
  assign \new_[29411]_  = (~\new_[30859]_  | ~\new_[5970]_ ) & (~\new_[31337]_  | ~\new_[6048]_ );
  assign \new_[29412]_  = (~\new_[5913]_  | ~\new_[31211]_ ) & (~\new_[6206]_  | ~\new_[31337]_ );
  assign \new_[29413]_  = ~\new_[30466]_  | ~\new_[30610]_ ;
  assign \new_[29414]_  = ~\new_[30751]_  | ~\new_[30610]_ ;
  assign \new_[29415]_  = ~\new_[30497]_  | ~\new_[6052]_ ;
  assign \new_[29416]_  = ~\new_[30472]_  & ~\new_[5830]_ ;
  assign \new_[29417]_  = ~\new_[30468]_  | ~n8779;
  assign \new_[29418]_  = ~\new_[30619]_  | ~n8799;
  assign \new_[29419]_  = ~\new_[30660]_  | ~\new_[6040]_ ;
  assign \new_[29420]_  = \new_[31208]_  & \new_[30745]_ ;
  assign \new_[29421]_  = ~\new_[30078]_ ;
  assign \new_[29422]_  = ~\new_[30645]_  | ~\new_[6211]_ ;
  assign \new_[29423]_  = ~\new_[30673]_  & ~\new_[6204]_ ;
  assign \new_[29424]_  = \new_[30807]_  | \new_[6040]_ ;
  assign \new_[29425]_  = (~\new_[31022]_  | ~\new_[5965]_ ) & (~\new_[31550]_  | ~\new_[5966]_ );
  assign \new_[29426]_  = (~\new_[6189]_  | ~\new_[30970]_ ) & (~\new_[5992]_  | ~\new_[31437]_ );
  assign \new_[29427]_  = ~\new_[6093]_  | ~\new_[6092]_ ;
  assign \new_[29428]_  = \new_[30816]_  & \new_[31189]_ ;
  assign \new_[29429]_  = ~\new_[30479]_  | ~n8364;
  assign \new_[29430]_  = ~\new_[30446]_  | ~\new_[30721]_ ;
  assign \new_[29431]_  = ~\new_[30598]_  & ~\new_[31593]_ ;
  assign \new_[29432]_  = ~\new_[30619]_  | ~n8574;
  assign \new_[29433]_  = \new_[30473]_  & \new_[5931]_ ;
  assign \new_[29434]_  = \new_[30422]_  & \new_[31197]_ ;
  assign \new_[29435]_  = \new_[30419]_  | \new_[31413]_ ;
  assign \new_[29436]_  = ~\new_[30651]_  & ~\new_[31777]_ ;
  assign \new_[29437]_  = \new_[30670]_  & \new_[6070]_ ;
  assign \new_[29438]_  = (~\new_[5964]_  | ~\new_[30937]_ ) & (~\new_[6246]_  | ~\new_[31328]_ );
  assign \new_[29439]_  = \new_[30608]_  & \new_[31422]_ ;
  assign \new_[29440]_  = ~\new_[30564]_  & ~\new_[31741]_ ;
  assign \new_[29441]_  = ~\new_[30219]_ ;
  assign \new_[29442]_  = \new_[30763]_  & \new_[5910]_ ;
  assign \new_[29443]_  = ~\new_[30515]_  & ~\new_[31596]_ ;
  assign \new_[29444]_  = \new_[30650]_  & \new_[5967]_ ;
  assign \new_[29445]_  = ~\new_[30223]_ ;
  assign \new_[29446]_  = \new_[30770]_  | \new_[5983]_ ;
  assign \new_[29447]_  = \new_[30426]_  & \new_[5966]_ ;
  assign \new_[29448]_  = ~\new_[30541]_  | ~\new_[30726]_ ;
  assign \new_[29449]_  = ~\new_[30502]_  | ~\new_[30507]_ ;
  assign \new_[29450]_  = ~\new_[30420]_  & ~\new_[30426]_ ;
  assign \new_[29451]_  = ~\new_[30423]_  & ~\new_[31562]_ ;
  assign \new_[29452]_  = ~\new_[30717]_ ;
  assign \new_[29453]_  = ~\new_[30833]_  | ~\new_[5926]_ ;
  assign \new_[29454]_  = ~\new_[30648]_  | ~\new_[30750]_ ;
  assign \new_[29455]_  = ~\new_[29885]_ ;
  assign \new_[29456]_  = ~\new_[30272]_ ;
  assign \new_[29457]_  = ~\new_[30708]_  & ~\new_[31776]_ ;
  assign \new_[29458]_  = ~\new_[30736]_  & ~\new_[31915]_ ;
  assign \new_[29459]_  = ~\new_[30629]_  | ~\new_[6032]_ ;
  assign \new_[29460]_  = ~\new_[30788]_  | ~\new_[30784]_ ;
  assign \new_[29461]_  = ~\new_[30696]_  & ~\new_[30618]_ ;
  assign \new_[29462]_  = (~\new_[5931]_  | ~\new_[31136]_ ) & (~\new_[5930]_  | ~\new_[31263]_ );
  assign \new_[29463]_  = (~\new_[5978]_  | ~\new_[31468]_ ) & (~\new_[6196]_  | ~\new_[31050]_ );
  assign \new_[29464]_  = ~\new_[30706]_  | ~\new_[30820]_ ;
  assign \new_[29465]_  = ~\new_[29762]_ ;
  assign \new_[29466]_  = \new_[30432]_  & \new_[31491]_ ;
  assign \new_[29467]_  = ~\new_[30751]_  | ~\new_[5995]_ ;
  assign \new_[29468]_  = ~\new_[30755]_  & ~\new_[30719]_ ;
  assign \new_[29469]_  = ~\new_[30554]_  | ~\new_[5987]_ ;
  assign \new_[29470]_  = ~\new_[30715]_  & ~\new_[30789]_ ;
  assign \new_[29471]_  = ~\new_[30665]_  | ~\new_[6205]_ ;
  assign \new_[29472]_  = \new_[31135]_  & \new_[30712]_ ;
  assign \new_[29473]_  = (~\new_[5981]_  | ~\new_[30944]_ ) & (~\new_[6064]_  | ~\new_[31487]_ );
  assign \new_[29474]_  = ~\new_[30837]_  & ~\new_[30662]_ ;
  assign \new_[29475]_  = ~\new_[30636]_  | ~\new_[6273]_ ;
  assign \new_[29476]_  = ~\new_[32321]_  | ~m1_stb_i;
  assign \new_[29477]_  = ~\new_[30438]_  & ~\new_[31819]_ ;
  assign \new_[29478]_  = ~\new_[30505]_  | ~\new_[6199]_ ;
  assign \new_[29479]_  = ~\new_[30582]_  | ~\new_[30726]_ ;
  assign \new_[29480]_  = ~\new_[30780]_  & ~\new_[30581]_ ;
  assign \new_[29481]_  = ~\new_[30443]_  | ~\new_[30697]_ ;
  assign \new_[29482]_  = \new_[30617]_  & \new_[6209]_ ;
  assign \new_[29483]_  = ~\new_[30694]_  & ~\new_[30660]_ ;
  assign \new_[29484]_  = ~\new_[30611]_  | ~n8429;
  assign \new_[29485]_  = \new_[30723]_  & \new_[6090]_ ;
  assign \new_[29486]_  = ~\new_[30847]_  | ~\new_[5927]_ ;
  assign \new_[29487]_  = ~\new_[30432]_  | ~\new_[5916]_ ;
  assign \new_[29488]_  = ~\new_[30949]_  & ~\new_[31844]_ ;
  assign \new_[29489]_  = ~\new_[30675]_  & ~\new_[30568]_ ;
  assign \new_[29490]_  = \new_[30550]_  & \new_[6204]_ ;
  assign \new_[29491]_  = ~\new_[32260]_  | ~m5_stb_i;
  assign \new_[29492]_  = \new_[31652]_  | \new_[30570]_ ;
  assign \new_[29493]_  = ~\new_[30662]_  | ~\new_[5925]_ ;
  assign \new_[29494]_  = \new_[30671]_  & \new_[5991]_ ;
  assign \new_[29495]_  = ~\new_[30259]_ ;
  assign \new_[29496]_  = (~\new_[31072]_  | ~\new_[5925]_ ) & (~\new_[31339]_  | ~\new_[5995]_ );
  assign \new_[29497]_  = ~\new_[30611]_  | ~n8304;
  assign \new_[29498]_  = ~\new_[30757]_  & ~\new_[31928]_ ;
  assign \new_[29499]_  = ~\new_[30553]_  | ~\new_[30765]_ ;
  assign \new_[29500]_  = ~\new_[30612]_  & ~\new_[30540]_ ;
  assign \new_[29501]_  = ~\new_[29983]_ ;
  assign \new_[29502]_  = \new_[30426]_  & \new_[6176]_ ;
  assign \new_[29503]_  = ~\new_[30677]_  | ~\new_[6270]_ ;
  assign \new_[29504]_  = (~\new_[31119]_  | ~\new_[6000]_ ) & (~\new_[31221]_  | ~\new_[5929]_ );
  assign \new_[29505]_  = ~\new_[30531]_  | ~\new_[4155]_ ;
  assign \new_[29506]_  = ~\new_[30173]_ ;
  assign \new_[29507]_  = (~\new_[30882]_  | ~\new_[5969]_ ) & (~\new_[31393]_  | ~\new_[6046]_ );
  assign \new_[29508]_  = ~\new_[30099]_ ;
  assign \new_[29509]_  = (~\new_[6094]_  | ~\new_[31495]_ ) & (~\new_[6033]_  | ~\new_[30978]_ );
  assign \new_[29510]_  = (~\new_[31212]_  | ~\new_[6049]_ ) & (~\new_[31434]_  | ~\new_[6053]_ );
  assign \new_[29511]_  = (~\new_[6037]_  | ~\new_[31008]_ ) & (~\new_[6041]_  | ~\new_[31550]_ );
  assign \new_[29512]_  = (~\new_[5921]_  | ~\new_[31220]_ ) & (~\new_[6072]_  | ~\new_[30973]_ );
  assign \new_[29513]_  = (~\new_[31468]_  | ~\new_[5900]_ ) & (~\new_[31050]_  | ~\new_[6057]_ );
  assign \new_[29514]_  = (~\new_[31317]_  | ~\new_[5901]_ ) & (~\new_[31158]_  | ~\new_[6061]_ );
  assign \new_[29515]_  = (~\new_[5918]_  | ~\new_[31451]_ ) & (~\new_[6069]_  | ~\new_[30956]_ );
  assign \new_[29516]_  = (~\new_[31495]_  | ~\new_[5894]_ ) & (~\new_[30978]_  | ~\new_[6034]_ );
  assign \new_[29517]_  = (~\new_[30989]_  | ~\new_[5980]_ ) & (~\new_[31452]_  | ~\new_[6060]_ );
  assign \new_[29518]_  = (~\new_[30936]_  | ~\new_[6005]_ ) & (~\new_[31303]_  | ~\new_[6217]_ );
  assign \new_[29519]_  = (~\new_[31451]_  | ~\new_[5903]_ ) & (~\new_[30956]_  | ~\new_[6070]_ );
  assign \new_[29520]_  = (~\new_[6211]_  | ~\new_[31158]_ ) & (~\new_[6273]_  | ~\new_[31487]_ );
  assign \new_[29521]_  = (~\new_[6043]_  | ~\new_[30986]_ ) & (~\new_[6044]_  | ~\new_[30882]_ );
  assign \new_[29522]_  = (~\new_[6190]_  | ~\new_[30970]_ ) & (~\new_[5991]_  | ~\new_[31437]_ );
  assign \new_[29523]_  = (~\new_[6038]_  | ~\new_[31022]_ ) & (~\new_[6176]_  | ~\new_[31550]_ );
  assign \new_[29524]_  = (~\new_[6003]_  | ~\new_[31136]_ ) & (~\new_[6183]_  | ~\new_[31263]_ );
  assign \new_[29525]_  = (~\new_[5988]_  | ~\new_[31075]_ ) & (~\new_[6214]_  | ~\new_[31228]_ );
  assign \new_[29526]_  = (~\new_[6068]_  | ~\new_[31055]_ ) & (~\new_[6213]_  | ~\new_[31518]_ );
  assign \new_[29527]_  = ~\new_[30285]_ ;
  assign \new_[29528]_  = ~\new_[30478]_  & ~\new_[30703]_ ;
  assign \new_[29529]_  = (~\new_[31543]_  | ~\new_[5933]_ ) & (~\new_[30908]_  | ~\new_[6270]_ );
  assign \new_[29530]_  = (~\new_[6074]_  | ~\new_[31220]_ ) & (~\new_[6073]_  | ~\new_[30973]_ );
  assign \new_[29531]_  = \new_[30680]_  & \new_[5989]_ ;
  assign \new_[29532]_  = ~\new_[30836]_  & ~\new_[31039]_ ;
  assign \new_[29533]_  = \new_[30436]_  | \new_[6094]_ ;
  assign \new_[29534]_  = ~\new_[30749]_  & ~\new_[31141]_ ;
  assign \new_[29535]_  = ~\new_[30435]_  & ~\new_[31416]_ ;
  assign \new_[29536]_  = ~\new_[30543]_  & ~\new_[30591]_ ;
  assign \new_[29537]_  = ~\new_[30732]_ ;
  assign \new_[29538]_  = \new_[30758]_  & \new_[31180]_ ;
  assign \new_[29539]_  = ~\new_[30675]_  | ~\new_[30717]_ ;
  assign \new_[29540]_  = ~\new_[30765]_ ;
  assign \new_[29541]_  = ~\new_[30102]_ ;
  assign \new_[29542]_  = ~\new_[30593]_  & ~\new_[5930]_ ;
  assign \new_[29543]_  = ~\new_[30182]_ ;
  assign \new_[29544]_  = ~\new_[29782]_ ;
  assign \new_[29545]_  = ~\new_[29781]_ ;
  assign \new_[29546]_  = ~\new_[6093]_  & ~\new_[6092]_ ;
  assign \new_[29547]_  = \new_[30759]_  & \new_[31645]_ ;
  assign \new_[29548]_  = ~\new_[30421]_  & ~\new_[31104]_ ;
  assign \new_[29549]_  = \new_[30512]_  & \new_[5964]_ ;
  assign \new_[29550]_  = ~\new_[30504]_  | ~\new_[4209]_ ;
  assign \new_[29551]_  = ~\new_[30780]_  | ~\new_[30572]_ ;
  assign \new_[29552]_  = \new_[30456]_  | \new_[6078]_ ;
  assign \new_[29553]_  = ~\new_[30526]_ ;
  assign \new_[29554]_  = ~\new_[30479]_  | ~n8734;
  assign \new_[29555]_  = \new_[30441]_  | \new_[6094]_ ;
  assign \new_[29556]_  = ~\new_[30190]_ ;
  assign \new_[29557]_  = ~\new_[29774]_ ;
  assign \new_[29558]_  = ~\new_[30554]_  | ~\new_[30765]_ ;
  assign \new_[29559]_  = ~\new_[30611]_  | ~n8899;
  assign \new_[29560]_  = ~\new_[30261]_ ;
  assign \new_[29561]_  = ~\new_[30633]_  & ~\new_[30676]_ ;
  assign \new_[29562]_  = ~\new_[30468]_  | ~n8519;
  assign \new_[29563]_  = ~\new_[30470]_  | ~\new_[4272]_ ;
  assign \new_[29564]_  = ~\new_[30128]_ ;
  assign \new_[29565]_  = ~\new_[30257]_ ;
  assign \new_[29566]_  = ~\new_[30445]_  & ~\new_[31901]_ ;
  assign \new_[29567]_  = ~\new_[30406]_ ;
  assign \new_[29568]_  = ~\new_[29887]_ ;
  assign \new_[29569]_  = ~\new_[30729]_  | ~\new_[4271]_ ;
  assign \new_[29570]_  = \new_[30664]_  & \new_[6269]_ ;
  assign \new_[29571]_  = ~\new_[29995]_ ;
  assign \new_[29572]_  = \new_[30623]_  & \new_[5970]_ ;
  assign \new_[29573]_  = ~\new_[30006]_ ;
  assign \new_[29574]_  = ~\new_[30654]_  | ~n8499;
  assign \new_[29575]_  = \new_[6197]_  | \new_[6057]_ ;
  assign \new_[29576]_  = ~\new_[30409]_ ;
  assign \new_[29577]_  = ~\new_[30713]_  & ~\new_[30642]_ ;
  assign \new_[29578]_  = ~\new_[29888]_ ;
  assign \new_[29579]_  = ~\new_[31492]_  & ~\new_[30454]_ ;
  assign \new_[29580]_  = ~\new_[30498]_  & ~\new_[31014]_ ;
  assign \new_[29581]_  = ~\new_[30702]_  | ~\new_[6268]_ ;
  assign \new_[29582]_  = ~\new_[30280]_ ;
  assign \new_[29583]_  = ~\new_[29968]_ ;
  assign \new_[29584]_  = \new_[30821]_  | \new_[5978]_ ;
  assign \new_[29585]_  = ~\new_[30480]_  | ~\new_[31763]_ ;
  assign \new_[29586]_  = ~\new_[30760]_  & ~\new_[6064]_ ;
  assign \new_[29587]_  = (~\new_[6036]_  | ~\new_[31216]_ ) & (~\new_[6039]_  | ~\new_[31022]_ );
  assign \new_[29588]_  = ~\new_[30212]_ ;
  assign \new_[29589]_  = ~\new_[30476]_  | ~\new_[4255]_ ;
  assign \new_[29590]_  = ~\new_[30130]_ ;
  assign \new_[29591]_  = ~\new_[30619]_  | ~n8584;
  assign \new_[29592]_  = ~\new_[30619]_  | ~n8659;
  assign \new_[29593]_  = ~\new_[30331]_ ;
  assign \new_[29594]_  = ~\new_[30654]_  | ~n8529;
  assign \new_[29595]_  = \new_[30805]_  & \new_[4248]_ ;
  assign \new_[29596]_  = ~\new_[30619]_  | ~n8644;
  assign \new_[29597]_  = ~\new_[29969]_ ;
  assign \new_[29598]_  = ~\new_[30697]_ ;
  assign \new_[29599]_  = ~\new_[30463]_  | ~\new_[5914]_ ;
  assign \new_[29600]_  = ~\new_[30582]_  | ~\new_[6245]_ ;
  assign \new_[29601]_  = ~\new_[30661]_  & ~\new_[30710]_ ;
  assign \new_[29602]_  = ~\new_[29902]_ ;
  assign \new_[29603]_  = \new_[30827]_  & \new_[30999]_ ;
  assign \new_[29604]_  = ~\new_[31122]_  & ~\new_[30454]_ ;
  assign \new_[29605]_  = ~\new_[30468]_  | ~n8394;
  assign \new_[29606]_  = ~\new_[30105]_ ;
  assign \new_[29607]_  = ~\new_[30533]_  | ~n8729;
  assign \new_[29608]_  = ~\new_[29799]_ ;
  assign \new_[29609]_  = ~\new_[30468]_  | ~n8889;
  assign \new_[29610]_  = ~\new_[30658]_  | ~n8919;
  assign \new_[29611]_  = ~\new_[30580]_  & ~\new_[4440]_ ;
  assign \new_[29612]_  = \new_[30585]_  | \new_[5926]_ ;
  assign \new_[29613]_  = \new_[30679]_  & \new_[4444]_ ;
  assign \new_[29614]_  = ~\new_[30658]_  | ~n8829;
  assign \new_[29615]_  = ~\new_[30611]_  | ~n8859;
  assign \new_[29616]_  = ~\new_[30472]_  & ~\new_[30925]_ ;
  assign \new_[29617]_  = ~\new_[30690]_  | ~n8444;
  assign \new_[29618]_  = ~\new_[30654]_  | ~n8379;
  assign \new_[29619]_  = ~\new_[29767]_ ;
  assign \new_[29620]_  = \new_[30518]_  | \new_[6040]_ ;
  assign \new_[29621]_  = \new_[30745]_  & \new_[30592]_ ;
  assign \new_[29622]_  = \new_[30621]_  & \new_[5930]_ ;
  assign \new_[29623]_  = ~\new_[30121]_ ;
  assign \new_[29624]_  = ~\new_[30638]_  & ~\new_[30526]_ ;
  assign \new_[29625]_  = \new_[30827]_  & \new_[30869]_ ;
  assign \new_[29626]_  = ~\new_[30690]_  | ~n8814;
  assign \new_[29627]_  = \new_[30674]_  & \new_[30562]_ ;
  assign \new_[29628]_  = \new_[30844]_  & \new_[30681]_ ;
  assign \new_[29629]_  = ~\new_[30103]_ ;
  assign \new_[29630]_  = ~\new_[30421]_  & ~\new_[6269]_ ;
  assign \new_[29631]_  = \new_[31111]_  & \new_[30592]_ ;
  assign \new_[29632]_  = ~\new_[30620]_  & ~\new_[30630]_ ;
  assign \new_[29633]_  = ~\new_[30292]_ ;
  assign \new_[29634]_  = ~\new_[30619]_  | ~n8654;
  assign \new_[29635]_  = \new_[30601]_  & \new_[6190]_ ;
  assign \new_[29636]_  = \new_[30506]_  & \new_[30844]_ ;
  assign \new_[29637]_  = ~\new_[30187]_ ;
  assign \new_[29638]_  = \new_[31089]_  | \new_[6031]_ ;
  assign \new_[29639]_  = ~\new_[30086]_ ;
  assign \new_[29640]_  = \new_[30844]_  & \new_[31200]_ ;
  assign \new_[29641]_  = \new_[31206]_  & \new_[30712]_ ;
  assign \new_[29642]_  = ~\new_[30605]_  & ~\new_[30993]_ ;
  assign \new_[29643]_  = ~\new_[30156]_ ;
  assign \new_[29644]_  = ~\new_[30611]_  | ~n8759;
  assign \new_[29645]_  = ~\new_[6039]_  | ~\new_[5965]_ ;
  assign \new_[29646]_  = ~\new_[30493]_  | ~\new_[6210]_ ;
  assign \new_[29647]_  = ~\new_[30786]_ ;
  assign \new_[29648]_  = ~\new_[29910]_ ;
  assign \new_[29649]_  = ~\new_[30823]_  & ~\new_[31265]_ ;
  assign \new_[29650]_  = ~\new_[30329]_ ;
  assign \new_[29651]_  = \new_[30745]_  & \new_[31004]_ ;
  assign \new_[29652]_  = ~\new_[30009]_ ;
  assign \new_[29653]_  = ~\new_[30619]_  | ~n8744;
  assign \new_[29654]_  = ~\new_[30479]_  | ~n8319;
  assign \new_[29655]_  = \new_[31588]_  | \new_[30477]_ ;
  assign \new_[29656]_  = ~\new_[30811]_  | ~\new_[4153]_ ;
  assign \new_[29657]_  = ~\new_[30479]_  | ~n8924;
  assign \new_[29658]_  = ~\new_[30843]_  & ~\new_[6206]_ ;
  assign \new_[29659]_  = \new_[30424]_  | \new_[30976]_ ;
  assign \new_[29660]_  = ~\new_[30784]_ ;
  assign \new_[29661]_  = \new_[30492]_  & \new_[5981]_ ;
  assign \new_[29662]_  = ~\new_[30722]_  & ~\new_[31645]_ ;
  assign \new_[29663]_  = ~\new_[29863]_ ;
  assign \new_[29664]_  = \new_[31615]_  | \new_[30596]_ ;
  assign \new_[29665]_  = ~\new_[30627]_  | ~\new_[6060]_ ;
  assign \new_[29666]_  = ~\new_[29937]_ ;
  assign \new_[29667]_  = ~\new_[30658]_  | ~n8504;
  assign \new_[29668]_  = ~\new_[30468]_  | ~n8724;
  assign \new_[29669]_  = ~\new_[30053]_ ;
  assign \new_[29670]_  = \new_[30462]_  & \new_[30422]_ ;
  assign \new_[29671]_  = ~\new_[29840]_ ;
  assign \new_[29672]_  = ~\new_[30117]_ ;
  assign \new_[29673]_  = ~\new_[30369]_ ;
  assign \new_[29674]_  = ~\new_[31492]_  & ~\m7_addr_i[29] ;
  assign \new_[29675]_  = ~\new_[30594]_  | ~\new_[6072]_ ;
  assign \new_[29676]_  = ~\new_[30104]_ ;
  assign \new_[29677]_  = \new_[30815]_  & \new_[5996]_ ;
  assign \new_[29678]_  = \new_[30634]_  & \new_[31096]_ ;
  assign \new_[29679]_  = ~\new_[30403]_ ;
  assign \new_[29680]_  = ~\new_[30533]_  | ~n8514;
  assign \new_[29681]_  = ~\new_[30390]_ ;
  assign \new_[29682]_  = ~\new_[30068]_ ;
  assign \new_[29683]_  = ~\new_[30658]_  | ~n8864;
  assign \new_[29684]_  = ~\new_[30619]_  | ~n8549;
  assign \new_[29685]_  = ~\new_[30055]_ ;
  assign \new_[29686]_  = ~\new_[30699]_  & ~\new_[31494]_ ;
  assign \new_[29687]_  = ~\new_[30690]_  | ~n8694;
  assign \new_[29688]_  = \new_[31345]_  | \new_[30596]_ ;
  assign \new_[29689]_  = ~\new_[30809]_  | ~\new_[5914]_ ;
  assign \new_[29690]_  = ~\new_[30468]_  | ~n8874;
  assign \new_[29691]_  = ~\new_[30479]_  | ~n8324;
  assign \new_[29692]_  = ~\new_[30064]_ ;
  assign \new_[29693]_  = ~\new_[30658]_  | ~n8459;
  assign \new_[29694]_  = \new_[30759]_  & \new_[6246]_ ;
  assign \new_[29695]_  = ~\new_[30008]_ ;
  assign \new_[29696]_  = \new_[30829]_  & \new_[6064]_ ;
  assign \new_[29697]_  = ~\new_[30654]_  | ~n8629;
  assign \new_[29698]_  = ~\new_[30690]_  | ~n8554;
  assign \new_[29699]_  = ~\new_[30427]_  & ~\new_[4251]_ ;
  assign \new_[29700]_  = ~\new_[30183]_ ;
  assign \new_[29701]_  = ~\new_[29970]_ ;
  assign \new_[29702]_  = ~\new_[30611]_  | ~n8764;
  assign \new_[29703]_  = ~\new_[30529]_  & ~\new_[5919]_ ;
  assign \new_[29704]_  = \new_[30681]_  & \new_[30818]_ ;
  assign \new_[29705]_  = \new_[30462]_  & \new_[30802]_ ;
  assign \new_[29706]_  = \new_[31208]_  & \new_[30744]_ ;
  assign \new_[29707]_  = \new_[31061]_  & \new_[30537]_ ;
  assign \new_[29708]_  = \new_[30798]_  & \new_[30869]_ ;
  assign \new_[29709]_  = \new_[30806]_  & \new_[30924]_ ;
  assign \new_[29710]_  = \new_[30816]_  & \new_[31038]_ ;
  assign \new_[29711]_  = \new_[30798]_  & \new_[31152]_ ;
  assign \new_[29712]_  = ~\new_[29864]_ ;
  assign \new_[29713]_  = ~\new_[31182]_  & ~\new_[6031]_ ;
  assign \new_[29714]_  = ~\new_[30365]_ ;
  assign \new_[29715]_  = ~\new_[31312]_  & ~\new_[31538]_ ;
  assign \new_[29716]_  = ~\new_[30558]_  | ~\new_[30894]_ ;
  assign \new_[29717]_  = ~\new_[29923]_ ;
  assign \new_[29718]_  = ~\new_[6006]_  | ~\new_[6005]_ ;
  assign \new_[29719]_  = ~\new_[29842]_ ;
  assign \new_[29720]_  = ~\new_[30039]_ ;
  assign \new_[29721]_  = ~\new_[30069]_ ;
  assign \new_[29722]_  = ~\new_[29911]_ ;
  assign \new_[29723]_  = ~\new_[6039]_  & ~\new_[5965]_ ;
  assign \new_[29724]_  = ~\new_[29818]_ ;
  assign \new_[29725]_  = ~\new_[6043]_  & ~\new_[31397]_ ;
  assign \new_[29726]_  = ~\new_[29793]_ ;
  assign \new_[29727]_  = ~\new_[30479]_  | ~n8339;
  assign \new_[29728]_  = ~\new_[30405]_ ;
  assign \new_[29729]_  = ~\new_[30595]_  | ~\new_[6213]_ ;
  assign \new_[29730]_  = ~\new_[31021]_  & ~\new_[5996]_ ;
  assign \new_[29731]_  = ~\new_[30748]_  & ~\new_[30969]_ ;
  assign \new_[29732]_  = ~\new_[30533]_  | ~n8669;
  assign \new_[29733]_  = \new_[30609]_  & \new_[5913]_ ;
  assign \new_[29734]_  = ~\new_[30533]_  | ~n8439;
  assign \new_[29735]_  = ~\new_[30241]_ ;
  assign \new_[29736]_  = ~\new_[30386]_ ;
  assign \new_[29737]_  = ~\new_[29775]_ ;
  assign \new_[29738]_  = ~\new_[31685]_  | ~\new_[31588]_ ;
  assign \new_[29739]_  = ~\new_[6081]_  | ~\new_[5998]_ ;
  assign \new_[29740]_  = ~\new_[30662]_  | ~\new_[5924]_ ;
  assign \new_[29741]_  = ~\new_[6081]_  & ~\new_[5998]_ ;
  assign \new_[29742]_  = \new_[6050]_  | \new_[6049]_ ;
  assign \new_[29743]_  = ~\new_[30426]_ ;
  assign \new_[29744]_  = ~\new_[30399]_ ;
  assign \new_[29745]_  = ~\new_[30016]_ ;
  assign \new_[29746]_  = \new_[30766]_  | \new_[4054]_ ;
  assign \new_[29747]_  = ~\new_[30533]_  | ~n8784;
  assign \new_[29748]_  = ~\new_[29900]_ ;
  assign \new_[29749]_  = \new_[30756]_  & \new_[30827]_ ;
  assign \new_[29750]_  = ~\new_[30583]_  & ~\new_[31896]_ ;
  assign \new_[29751]_  = ~\new_[30521]_  | ~\new_[6216]_ ;
  assign \new_[29752]_  = \new_[30527]_  | \new_[31340]_ ;
  assign \new_[29753]_  = ~\new_[30401]_ ;
  assign \new_[29754]_  = ~\new_[30615]_ ;
  assign \new_[29755]_  = ~\new_[31491]_  & ~\new_[31121]_ ;
  assign \new_[29756]_  = \new_[30800]_  & \new_[5830]_ ;
  assign \new_[29757]_  = ~\new_[30618]_  | ~\new_[31157]_ ;
  assign \new_[29758]_  = ~\new_[30411]_ ;
  assign \new_[29759]_  = (~\new_[6193]_  | ~\new_[31451]_ ) & (~\new_[6191]_  | ~\new_[30956]_ );
  assign \new_[29760]_  = \new_[30776]_  & \new_[31165]_ ;
  assign \new_[29761]_  = ~\new_[30757]_  & ~\new_[30446]_ ;
  assign \new_[29762]_  = \new_[30901]_  | \new_[4084]_ ;
  assign \new_[29763]_  = ~\new_[31005]_  | ~\new_[4074]_ ;
  assign \new_[29764]_  = ~\new_[30588]_ ;
  assign \new_[29765]_  = ~\new_[30889]_  & ~\new_[4074]_ ;
  assign \new_[29766]_  = ~\new_[31394]_  & ~\new_[31033]_ ;
  assign \new_[29767]_  = ~\new_[30913]_  & ~\new_[4246]_ ;
  assign \new_[29768]_  = ~\new_[30943]_  | ~\new_[4042]_ ;
  assign \new_[29769]_  = ~\new_[30954]_  & ~\new_[30922]_ ;
  assign \new_[29770]_  = ~\new_[30720]_ ;
  assign \new_[29771]_  = ~\new_[31109]_  | ~\new_[4088]_ ;
  assign \new_[29772]_  = ~\new_[30865]_  & ~\new_[4271]_ ;
  assign \new_[29773]_  = ~\new_[30913]_  & ~\new_[31571]_ ;
  assign \new_[29774]_  = ~\new_[31170]_  & ~\new_[4038]_ ;
  assign \new_[29775]_  = ~\new_[6037]_  & ~\new_[5910]_ ;
  assign \new_[29776]_  = \new_[31006]_  & \new_[4096]_ ;
  assign \new_[29777]_  = ~\new_[30941]_  & ~\new_[3879]_ ;
  assign \new_[29778]_  = ~\new_[30493]_ ;
  assign \new_[29779]_  = \new_[31155]_  & \new_[30997]_ ;
  assign \new_[29780]_  = ~\new_[30769]_ ;
  assign \new_[29781]_  = ~\new_[31106]_  | ~\new_[4239]_ ;
  assign \new_[29782]_  = ~\new_[30927]_  | ~\new_[4089]_ ;
  assign \new_[29783]_  = ~\new_[31142]_  | ~\new_[4072]_ ;
  assign \new_[29784]_  = ~\new_[31077]_  & ~\new_[31556]_ ;
  assign \new_[29785]_  = ~\new_[31002]_  | ~\new_[4153]_ ;
  assign \new_[29786]_  = ~\new_[31011]_  & ~\new_[31096]_ ;
  assign \new_[29787]_  = \new_[31097]_  | \new_[31774]_ ;
  assign \new_[29788]_  = \new_[31059]_  & \new_[31210]_ ;
  assign \new_[29789]_  = ~\new_[31170]_  & ~\new_[31702]_ ;
  assign \new_[29790]_  = ~\new_[30693]_ ;
  assign \new_[29791]_  = \new_[30911]_  & \new_[4110]_ ;
  assign \new_[29792]_  = ~\new_[30846]_ ;
  assign \new_[29793]_  = \new_[6080]_  | \new_[31765]_ ;
  assign \new_[29794]_  = ~\new_[30612]_ ;
  assign \new_[29795]_  = \new_[6056]_  | \new_[31866]_ ;
  assign \new_[29796]_  = ~\new_[31725]_  & ~\new_[6060]_ ;
  assign \new_[29797]_  = ~\new_[31616]_  | ~\new_[5965]_ ;
  assign \new_[29798]_  = ~\new_[30442]_ ;
  assign \new_[29799]_  = ~\new_[31149]_  & ~\new_[31558]_ ;
  assign \new_[29800]_  = ~\new_[31799]_  | ~\new_[6217]_ ;
  assign \new_[29801]_  = ~\new_[30742]_ ;
  assign \new_[29802]_  = ~\new_[30684]_ ;
  assign \new_[29803]_  = \new_[31553]_  | \new_[5998]_ ;
  assign \new_[29804]_  = ~\m4_addr_i[31]  & ~\new_[31922]_ ;
  assign \new_[29805]_  = \new_[31118]_  | \new_[6210]_ ;
  assign \new_[29806]_  = ~\new_[30446]_ ;
  assign \new_[29807]_  = \new_[31059]_  & \new_[31017]_ ;
  assign \new_[29808]_  = ~\new_[30502]_ ;
  assign \new_[29809]_  = \new_[31201]_  & \new_[4251]_ ;
  assign \new_[29810]_  = ~\new_[30678]_ ;
  assign \new_[29811]_  = ~\new_[31928]_  & ~\new_[6048]_ ;
  assign \new_[29812]_  = \new_[31905]_  & \new_[6215]_ ;
  assign \new_[29813]_  = ~\new_[30682]_ ;
  assign \new_[29814]_  = ~\new_[31139]_  & ~\new_[4094]_ ;
  assign \new_[29815]_  = ~\new_[30676]_ ;
  assign \new_[29816]_  = ~\new_[6036]_  | ~\new_[31800]_ ;
  assign \new_[29817]_  = \new_[31026]_  | \new_[31682]_ ;
  assign \new_[29818]_  = \new_[31725]_  & \new_[6060]_ ;
  assign \new_[29819]_  = \new_[31189]_  & \new_[31333]_ ;
  assign \new_[29820]_  = ~\new_[30810]_ ;
  assign \new_[29821]_  = ~\new_[30596]_ ;
  assign \new_[29822]_  = ~\new_[6073]_  & ~\new_[31895]_ ;
  assign \new_[29823]_  = \new_[31065]_  & \new_[30939]_ ;
  assign \new_[29824]_  = ~\new_[31925]_  | ~\new_[5902]_ ;
  assign \new_[29825]_  = ~\new_[31054]_  | ~\new_[4255]_ ;
  assign \new_[29826]_  = ~\new_[31092]_  & ~\new_[31590]_ ;
  assign \new_[29827]_  = ~\new_[30857]_  & ~\new_[31823]_ ;
  assign \new_[29828]_  = ~\new_[30467]_ ;
  assign \new_[29829]_  = ~\new_[31617]_  & ~\new_[5966]_ ;
  assign \new_[29830]_  = ~\new_[31184]_  & ~\new_[31713]_ ;
  assign \new_[29831]_  = \new_[30895]_  | \new_[31896]_ ;
  assign \new_[29832]_  = ~\new_[31819]_  & ~\new_[5922]_ ;
  assign \new_[29833]_  = ~\new_[30887]_  & ~\new_[4137]_ ;
  assign \new_[29834]_  = \new_[31837]_  | \new_[5990]_ ;
  assign \new_[29835]_  = \new_[6042]_  | \new_[31903]_ ;
  assign \new_[29836]_  = ~\new_[6199]_  & ~\new_[31887]_ ;
  assign \new_[29837]_  = ~\new_[30459]_ ;
  assign \new_[29838]_  = ~\new_[31156]_  | ~\new_[31442]_ ;
  assign \new_[29839]_  = ~\new_[31168]_  & ~\new_[4220]_ ;
  assign \new_[29840]_  = ~\new_[30932]_  | ~\new_[31681]_ ;
  assign \new_[29841]_  = ~\new_[31093]_  & ~\new_[4231]_ ;
  assign \new_[29842]_  = \new_[31660]_  & \new_[5971]_ ;
  assign \new_[29843]_  = ~\new_[31179]_  | ~\new_[31180]_ ;
  assign \new_[29844]_  = ~\new_[31608]_  | ~\new_[5980]_ ;
  assign \new_[29845]_  = \new_[6193]_  | \new_[31686]_ ;
  assign \new_[29846]_  = \new_[31038]_  & \new_[31333]_ ;
  assign \new_[29847]_  = \new_[31088]_  | \new_[5914]_ ;
  assign \new_[29848]_  = ~\new_[31078]_  & ~\new_[31852]_ ;
  assign \new_[29849]_  = ~\new_[31862]_  & ~\new_[6000]_ ;
  assign \new_[29850]_  = \new_[6074]_  | \new_[31707]_ ;
  assign \new_[29851]_  = ~\new_[30466]_ ;
  assign \new_[29852]_  = ~\new_[31669]_  | ~\new_[5963]_ ;
  assign \new_[29853]_  = ~\new_[30994]_  & ~\new_[4209]_ ;
  assign \new_[29854]_  = \new_[30962]_  & \new_[4103]_ ;
  assign \new_[29855]_  = ~\new_[30959]_  & ~\new_[4229]_ ;
  assign \new_[29856]_  = \new_[31195]_  & \new_[5930]_ ;
  assign \new_[29857]_  = \new_[31683]_  | \new_[6005]_ ;
  assign \new_[29858]_  = \new_[30890]_  & \new_[5981]_ ;
  assign \new_[29859]_  = \new_[6194]_  | \new_[31562]_ ;
  assign \new_[29860]_  = ~\new_[6083]_  | ~\new_[31839]_ ;
  assign \new_[29861]_  = ~\new_[31087]_  & ~\new_[4209]_ ;
  assign \new_[29862]_  = \new_[31660]_  | \new_[5971]_ ;
  assign \new_[29863]_  = ~\new_[30958]_  | ~\new_[31012]_ ;
  assign \new_[29864]_  = ~\new_[6045]_  | ~\new_[31569]_ ;
  assign \new_[29865]_  = ~\new_[31113]_  & ~\new_[4107]_ ;
  assign \new_[29866]_  = ~\new_[31440]_  | ~\new_[31588]_ ;
  assign \new_[29867]_  = ~\new_[30632]_ ;
  assign \new_[29868]_  = ~\new_[31120]_  | ~\new_[3886]_ ;
  assign \new_[29869]_  = ~\new_[30553]_ ;
  assign \new_[29870]_  = ~\new_[30688]_ ;
  assign \new_[29871]_  = \new_[31085]_  & \new_[6204]_ ;
  assign \new_[29872]_  = ~\new_[30474]_ ;
  assign \new_[29873]_  = ~\new_[30929]_  | ~\new_[31710]_ ;
  assign \new_[29874]_  = ~\new_[30929]_  | ~\new_[4211]_ ;
  assign \new_[29875]_  = ~\new_[30646]_ ;
  assign \new_[29876]_  = ~\new_[30891]_  & ~\new_[31401]_ ;
  assign \new_[29877]_  = ~\new_[30478]_ ;
  assign \new_[29878]_  = ~\new_[30461]_ ;
  assign \new_[29879]_  = ~\new_[30821]_ ;
  assign \new_[29880]_  = \new_[30886]_  & \new_[4202]_ ;
  assign \new_[29881]_  = ~\new_[31066]_  | ~\new_[31604]_ ;
  assign \new_[29882]_  = ~\new_[30938]_  & ~\new_[4449]_ ;
  assign \new_[29883]_  = ~\new_[30727]_ ;
  assign \new_[29884]_  = ~\new_[31915]_  | ~\new_[6245]_ ;
  assign \new_[29885]_  = ~\new_[31016]_  & ~\new_[31768]_ ;
  assign \new_[29886]_  = ~\new_[30945]_  | ~\new_[4442]_ ;
  assign \new_[29887]_  = ~\new_[30940]_  | ~\new_[4144]_ ;
  assign \new_[29888]_  = \new_[31086]_  | \new_[4235]_ ;
  assign \new_[29889]_  = ~\new_[30499]_ ;
  assign \new_[29890]_  = ~\new_[31789]_  & ~\new_[5929]_ ;
  assign \new_[29891]_  = ~\new_[31027]_  | ~\new_[4137]_ ;
  assign \new_[29892]_  = ~\new_[31203]_  | ~\new_[4237]_ ;
  assign \new_[29893]_  = ~\new_[31007]_  | ~\new_[4155]_ ;
  assign \new_[29894]_  = ~\new_[30441]_ ;
  assign \new_[29895]_  = ~\new_[6042]_  | ~\new_[31903]_ ;
  assign \new_[29896]_  = \new_[31616]_  | \new_[5965]_ ;
  assign \new_[29897]_  = ~\new_[30545]_ ;
  assign \new_[29898]_  = ~\new_[30946]_  & ~\new_[4451]_ ;
  assign \new_[29899]_  = ~\new_[30980]_  & ~\new_[4072]_ ;
  assign \new_[29900]_  = ~\new_[31023]_  | ~\new_[31828]_ ;
  assign \new_[29901]_  = \new_[6194]_  & \new_[31562]_ ;
  assign \new_[29902]_  = ~\new_[30895]_  & ~\new_[3882]_ ;
  assign \new_[29903]_  = ~\new_[6056]_  | ~\new_[31866]_ ;
  assign \new_[29904]_  = ~\new_[30962]_  | ~\new_[31744]_ ;
  assign \new_[29905]_  = ~\new_[31122]_  & ~\new_[31141]_ ;
  assign \new_[29906]_  = \new_[30914]_  & \new_[4051]_ ;
  assign \new_[29907]_  = ~\new_[30513]_ ;
  assign \new_[29908]_  = ~\new_[31213]_  & ~\new_[4058]_ ;
  assign \new_[29909]_  = ~\new_[30754]_ ;
  assign \new_[29910]_  = ~\new_[30950]_  | ~\new_[31911]_ ;
  assign \new_[29911]_  = ~\new_[31204]_  | ~\new_[4206]_ ;
  assign \new_[29912]_  = ~\new_[30438]_ ;
  assign \new_[29913]_  = ~\new_[31198]_  | ~\new_[4170]_ ;
  assign \new_[29914]_  = ~\new_[31063]_  & ~\new_[4139]_ ;
  assign \new_[29915]_  = ~\new_[30544]_ ;
  assign \new_[29916]_  = ~\new_[30680]_ ;
  assign \new_[29917]_  = ~\new_[31394]_  | ~\new_[31345]_ ;
  assign \new_[29918]_  = \new_[31036]_  & \new_[4440]_ ;
  assign \new_[29919]_  = ~\new_[30967]_  & ~\new_[31716]_ ;
  assign \new_[29920]_  = ~\new_[6174]_  & ~\new_[31593]_ ;
  assign \new_[29921]_  = ~\new_[30492]_ ;
  assign \new_[29922]_  = ~\new_[30984]_  | ~\new_[4086]_ ;
  assign \new_[29923]_  = ~\new_[6079]_  | ~\new_[6270]_ ;
  assign \new_[29924]_  = ~\new_[30888]_  | ~\new_[31717]_ ;
  assign \new_[29925]_  = ~\new_[31089]_  & ~\new_[31039]_ ;
  assign \new_[29926]_  = ~\new_[30525]_ ;
  assign \new_[29927]_  = ~\new_[31144]_  | ~\new_[4272]_ ;
  assign \new_[29928]_  = ~\new_[30922]_  & ~\new_[31498]_ ;
  assign \new_[29929]_  = ~\new_[31051]_  | ~\new_[31867]_ ;
  assign \new_[29930]_  = ~\new_[30573]_ ;
  assign \new_[29931]_  = ~\new_[31171]_  & ~\new_[4090]_ ;
  assign \new_[29932]_  = \new_[30923]_  | \new_[31455]_ ;
  assign \new_[29933]_  = ~\new_[30477]_ ;
  assign \new_[29934]_  = ~\new_[31186]_  & ~\new_[4156]_ ;
  assign \new_[29935]_  = ~\new_[30731]_ ;
  assign \new_[29936]_  = ~\new_[31928]_  | ~\new_[6048]_ ;
  assign \new_[29937]_  = \new_[30860]_  & \new_[6212]_ ;
  assign \new_[29938]_  = ~\new_[31915]_  & ~\new_[6245]_ ;
  assign \new_[29939]_  = \new_[30934]_  & \new_[31038]_ ;
  assign \new_[29940]_  = ~\new_[31046]_  & ~\new_[4130]_ ;
  assign \new_[29941]_  = \new_[30902]_  | \new_[4128]_ ;
  assign \new_[29942]_  = \new_[30909]_  | \new_[5983]_ ;
  assign \new_[29943]_  = ~\new_[30870]_  | ~\new_[31570]_ ;
  assign \new_[29944]_  = ~\new_[31149]_  & ~\new_[4175]_ ;
  assign \new_[29945]_  = ~\new_[30825]_ ;
  assign \new_[29946]_  = ~\new_[31060]_  & ~\new_[31727]_ ;
  assign \new_[29947]_  = \new_[31333]_  & \new_[31013]_ ;
  assign \new_[29948]_  = \new_[30934]_  & \new_[31145]_ ;
  assign \new_[29949]_  = ~\new_[31122]_  & ~\new_[31146]_ ;
  assign \new_[29950]_  = ~\new_[30604]_ ;
  assign \new_[29951]_  = ~\new_[31207]_  & ~\new_[30954]_ ;
  assign \new_[29952]_  = ~\new_[30955]_  & ~\new_[31802]_ ;
  assign \new_[29953]_  = ~\new_[30951]_  & ~\new_[31490]_ ;
  assign \new_[29954]_  = \new_[31065]_  & \new_[31111]_ ;
  assign \new_[29955]_  = ~\new_[30963]_  & ~\new_[31605]_ ;
  assign \new_[29956]_  = ~\new_[30735]_ ;
  assign \new_[29957]_  = ~\new_[30451]_ ;
  assign \new_[29958]_  = ~\new_[31163]_  & ~\new_[30850]_ ;
  assign \new_[29959]_  = ~\new_[30555]_ ;
  assign \new_[29960]_  = ~\new_[30898]_  & ~\new_[31723]_ ;
  assign \new_[29961]_  = \new_[31189]_  & \new_[30934]_ ;
  assign \new_[29962]_  = ~\new_[30554]_ ;
  assign \new_[29963]_  = ~\new_[31280]_  & ~\new_[30867]_ ;
  assign \new_[29964]_  = ~\new_[30751]_ ;
  assign \new_[29965]_  = ~\new_[30975]_  & ~\new_[31607]_ ;
  assign \new_[29966]_  = ~\new_[31069]_  & ~\new_[31580]_ ;
  assign \new_[29967]_  = ~\new_[30858]_  | ~\new_[4108]_ ;
  assign \new_[29968]_  = ~\new_[31071]_  & ~\new_[31601]_ ;
  assign \new_[29969]_  = ~\new_[31019]_  | ~\new_[4218]_ ;
  assign \new_[29970]_  = \new_[31034]_  & \new_[4451]_ ;
  assign \new_[29971]_  = ~\new_[30564]_ ;
  assign \new_[29972]_  = ~\new_[30771]_ ;
  assign \new_[29973]_  = ~\new_[30834]_ ;
  assign \new_[29974]_  = ~\new_[30910]_  | ~\new_[4240]_ ;
  assign \new_[29975]_  = ~\new_[30747]_ ;
  assign \new_[29976]_  = ~\new_[31164]_  & ~\new_[31327]_ ;
  assign \new_[29977]_  = ~\new_[31099]_  | ~\new_[4092]_ ;
  assign \new_[29978]_  = ~\new_[30569]_ ;
  assign \new_[29979]_  = ~\new_[30637]_ ;
  assign \new_[29980]_  = \new_[30996]_  & \new_[5919]_ ;
  assign \new_[29981]_  = \new_[31010]_  & \new_[4222]_ ;
  assign \new_[29982]_  = ~\new_[31067]_  | ~\new_[31433]_ ;
  assign \new_[29983]_  = ~\new_[31174]_  | ~\new_[4054]_ ;
  assign \new_[29984]_  = \new_[31024]_  | \new_[3875]_ ;
  assign \new_[29985]_  = \new_[31030]_  & \new_[4280]_ ;
  assign \new_[29986]_  = \new_[31118]_  | \new_[31411]_ ;
  assign \new_[29987]_  = ~\new_[30788]_ ;
  assign \new_[29988]_  = ~\new_[30551]_ ;
  assign \new_[29989]_  = ~\new_[30578]_ ;
  assign \new_[29990]_  = ~\new_[30454]_ ;
  assign \new_[29991]_  = ~\new_[30582]_ ;
  assign \new_[29992]_  = ~\new_[31029]_  & ~\new_[31602]_ ;
  assign \new_[29993]_  = ~\new_[31194]_  & ~\new_[30925]_ ;
  assign \new_[29994]_  = ~\new_[30921]_  & ~\new_[4123]_ ;
  assign \new_[29995]_  = ~\new_[31123]_  & ~\new_[31682]_ ;
  assign \new_[29996]_  = ~\new_[30584]_ ;
  assign \new_[29997]_  = ~\new_[30571]_ ;
  assign \new_[29998]_  = ~\new_[30560]_ ;
  assign \new_[29999]_  = ~\new_[30610]_ ;
  assign \new_[30000]_  = ~\new_[31098]_  | ~\new_[4061]_ ;
  assign \new_[30001]_  = \new_[31145]_  & \new_[31333]_ ;
  assign \new_[30002]_  = ~\new_[30599]_ ;
  assign \new_[30003]_  = ~\new_[30586]_ ;
  assign \new_[30004]_  = ~\new_[31093]_  & ~\new_[31809]_ ;
  assign \new_[30005]_  = ~\new_[31181]_  | ~\new_[31826]_ ;
  assign \new_[30006]_  = \new_[31169]_  | \new_[4148]_ ;
  assign \new_[30007]_  = ~\new_[30948]_  | ~\new_[6069]_ ;
  assign \new_[30008]_  = \new_[31103]_  & \new_[31649]_ ;
  assign \new_[30009]_  = \new_[31127]_  | \new_[4173]_ ;
  assign \new_[30010]_  = ~\new_[30814]_ ;
  assign \new_[30011]_  = ~\new_[30542]_ ;
  assign \new_[30012]_  = ~\new_[30833]_ ;
  assign \new_[30013]_  = ~\new_[30862]_  & ~\new_[30922]_ ;
  assign \new_[30014]_  = ~\new_[30595]_ ;
  assign \new_[30015]_  = ~\new_[30541]_ ;
  assign \new_[30016]_  = ~\new_[31056]_  | ~\new_[31806]_ ;
  assign \new_[30017]_  = \new_[31499]_  & \new_[6215]_ ;
  assign \new_[30018]_  = ~\new_[30764]_ ;
  assign \new_[30019]_  = ~\new_[31074]_  | ~\new_[31850]_ ;
  assign \new_[30020]_  = ~\new_[30736]_ ;
  assign \new_[30021]_  = ~\new_[31150]_  | ~\new_[4047]_ ;
  assign \new_[30022]_  = ~\new_[30855]_  | ~\new_[4084]_ ;
  assign \new_[30023]_  = \new_[31906]_  | \new_[31102]_ ;
  assign \new_[30024]_  = ~\new_[31018]_  & ~\new_[4444]_ ;
  assign \new_[30025]_  = ~\new_[30899]_  | ~\new_[4040]_ ;
  assign \new_[30026]_  = ~\new_[30915]_  & ~\new_[31138]_ ;
  assign \new_[30027]_  = \new_[30991]_  & \new_[5930]_ ;
  assign \new_[30028]_  = ~\new_[30645]_ ;
  assign \new_[30029]_  = ~\new_[30638]_ ;
  assign \new_[30030]_  = \new_[31092]_  | \new_[4227]_ ;
  assign \new_[30031]_  = \new_[31082]_  & \new_[31191]_ ;
  assign \new_[30032]_  = ~\new_[31032]_  & ~\new_[4168]_ ;
  assign \new_[30033]_  = ~\new_[30691]_ ;
  assign \new_[30034]_  = ~\new_[30950]_  | ~\new_[4164]_ ;
  assign \new_[30035]_  = \new_[30853]_  | \new_[4126]_ ;
  assign \new_[30036]_  = \new_[30863]_  & \new_[4445]_ ;
  assign \new_[30037]_  = ~\new_[30616]_ ;
  assign \new_[30038]_  = ~\new_[30686]_ ;
  assign \new_[30039]_  = \new_[6083]_  | \new_[31839]_ ;
  assign \new_[30040]_  = ~\new_[31205]_  & ~\new_[4056]_ ;
  assign \new_[30041]_  = ~\new_[30807]_ ;
  assign \new_[30042]_  = ~\new_[31166]_  & ~\new_[4206]_ ;
  assign \new_[30043]_  = ~\new_[31003]_  & ~\new_[4253]_ ;
  assign \new_[30044]_  = ~\new_[30971]_  & ~\new_[3888]_ ;
  assign \new_[30045]_  = \new_[30872]_  & \new_[6064]_ ;
  assign \new_[30046]_  = ~\new_[31030]_  | ~\new_[31627]_ ;
  assign \new_[30047]_  = ~\new_[30799]_ ;
  assign \new_[30048]_  = ~\new_[30849]_  | ~\new_[4123]_ ;
  assign \new_[30049]_  = ~\new_[30585]_ ;
  assign \new_[30050]_  = ~\new_[30823]_ ;
  assign \new_[30051]_  = ~\new_[30497]_ ;
  assign \new_[30052]_  = ~\new_[31037]_  & ~\new_[4146]_ ;
  assign \new_[30053]_  = ~\new_[30906]_  & ~\new_[4142]_ ;
  assign \new_[30054]_  = \new_[31090]_  | \new_[4276]_ ;
  assign \new_[30055]_  = ~\new_[31125]_  & ~\new_[31628]_ ;
  assign \new_[30056]_  = \new_[30933]_  | \new_[5917]_ ;
  assign \new_[30057]_  = ~\new_[31172]_  | ~\new_[31679]_ ;
  assign \new_[30058]_  = ~\new_[31097]_  & ~\new_[4158]_ ;
  assign \new_[30059]_  = ~\new_[30896]_  & ~\new_[31656]_ ;
  assign \new_[30060]_  = ~\new_[30871]_  & ~\new_[31498]_ ;
  assign \new_[30061]_  = ~\new_[31201]_  | ~\new_[31299]_ ;
  assign \new_[30062]_  = ~\new_[30905]_  & ~\new_[4155]_ ;
  assign \new_[30063]_  = ~\new_[30670]_ ;
  assign \new_[30064]_  = \new_[31079]_  & \new_[4077]_ ;
  assign \new_[30065]_  = ~\new_[30639]_ ;
  assign \new_[30066]_  = ~\new_[30647]_ ;
  assign \new_[30067]_  = ~\new_[31213]_  & ~\new_[31838]_ ;
  assign \new_[30068]_  = \new_[31009]_  & \new_[3877]_ ;
  assign \new_[30069]_  = \new_[30910]_  & \new_[31916]_ ;
  assign \new_[30070]_  = ~\new_[30519]_ ;
  assign \new_[30071]_  = ~\new_[30780]_ ;
  assign \new_[30072]_  = ~\new_[30961]_  & ~\new_[31886]_ ;
  assign \new_[30073]_  = \new_[31196]_  | \new_[31763]_ ;
  assign \new_[30074]_  = ~\new_[30902]_  & ~\new_[31899]_ ;
  assign \new_[30075]_  = ~\new_[30563]_ ;
  assign \new_[30076]_  = ~\new_[30977]_  & ~\new_[4260]_ ;
  assign \new_[30077]_  = \new_[31085]_  & \new_[30993]_ ;
  assign \new_[30078]_  = ~\new_[30983]_  & ~\new_[31909]_ ;
  assign \new_[30079]_  = \new_[30979]_  | \new_[4067]_ ;
  assign \new_[30080]_  = ~\new_[31131]_  & ~\new_[4442]_ ;
  assign \new_[30081]_  = ~\new_[30651]_ ;
  assign \new_[30082]_  = \new_[31175]_  & \new_[5994]_ ;
  assign \new_[30083]_  = ~\new_[31188]_  | ~\new_[4121]_ ;
  assign \new_[30084]_  = ~\new_[30932]_  | ~\new_[4177]_ ;
  assign \new_[30085]_  = \new_[31111]_  & \new_[31004]_ ;
  assign \new_[30086]_  = \new_[31062]_  | \new_[4121]_ ;
  assign \new_[30087]_  = \new_[31031]_  & \new_[31587]_ ;
  assign \new_[30088]_  = \new_[31206]_  & \new_[30997]_ ;
  assign \new_[30089]_  = ~\new_[30543]_ ;
  assign \new_[30090]_  = ~\new_[31115]_  | ~\new_[31108]_ ;
  assign \new_[30091]_  = ~\new_[30447]_ ;
  assign \new_[30092]_  = ~\new_[31073]_  | ~\new_[31417]_ ;
  assign \new_[30093]_  = ~\new_[30695]_ ;
  assign \new_[30094]_  = ~\new_[31099]_  | ~\new_[31566]_ ;
  assign \new_[30095]_  = ~\new_[30959]_  & ~\new_[31918]_ ;
  assign \new_[30096]_  = ~\new_[30431]_ ;
  assign \new_[30097]_  = ~\new_[31019]_  | ~\new_[31413]_ ;
  assign \new_[30098]_  = ~\new_[30580]_ ;
  assign \new_[30099]_  = \new_[31026]_  | \new_[4453]_ ;
  assign \new_[30100]_  = \new_[30981]_  | \new_[31340]_ ;
  assign \new_[30101]_  = ~\new_[31086]_  & ~\new_[31932]_ ;
  assign \new_[30102]_  = \new_[30881]_  | \new_[4063]_ ;
  assign \new_[30103]_  = ~\new_[31080]_  | ~\new_[31811]_ ;
  assign \new_[30104]_  = ~\new_[31084]_  | ~\new_[31880]_ ;
  assign \new_[30105]_  = ~\new_[30873]_  | ~\new_[31711]_ ;
  assign \new_[30106]_  = ~\new_[31146]_  & ~\new_[31355]_ ;
  assign \new_[30107]_  = ~\new_[30746]_ ;
  assign \new_[30108]_  = ~\new_[31193]_  & ~\new_[31274]_ ;
  assign \new_[30109]_  = ~\new_[30650]_ ;
  assign \new_[30110]_  = \new_[31179]_  & \new_[6071]_ ;
  assign \new_[30111]_  = ~\new_[30694]_ ;
  assign \new_[30112]_  = ~\new_[31799]_  & ~\new_[6217]_ ;
  assign \new_[30113]_  = ~\new_[31146]_  & ~\new_[31492]_ ;
  assign \new_[30114]_  = ~\new_[30896]_  & ~\new_[4264]_ ;
  assign \new_[30115]_  = ~\new_[30630]_ ;
  assign \new_[30116]_  = ~\new_[30538]_ ;
  assign \new_[30117]_  = ~\new_[31056]_  | ~\new_[4267]_ ;
  assign \new_[30118]_  = \new_[30885]_  & \new_[4262]_ ;
  assign \new_[30119]_  = \new_[30923]_  | \new_[6072]_ ;
  assign \new_[30120]_  = \new_[31102]_  | \new_[31690]_ ;
  assign \new_[30121]_  = ~\new_[30977]_  & ~\new_[31666]_ ;
  assign \new_[30122]_  = ~\new_[31156]_  | ~\new_[6184]_ ;
  assign \new_[30123]_  = ~\new_[30899]_  | ~\new_[31769]_ ;
  assign \new_[30124]_  = ~\new_[31141]_  & ~\new_[31492]_ ;
  assign \new_[30125]_  = ~\new_[31066]_  | ~\new_[4160]_ ;
  assign \new_[30126]_  = ~\new_[30873]_  | ~\new_[4170]_ ;
  assign \new_[30127]_  = ~\new_[31058]_  & ~\new_[4162]_ ;
  assign \new_[30128]_  = \new_[31016]_  | \new_[4045]_ ;
  assign \new_[30129]_  = \new_[30958]_  & \new_[4151]_ ;
  assign \new_[30130]_  = ~\new_[30920]_  & ~\new_[3884]_ ;
  assign \new_[30131]_  = \new_[30934]_  & \new_[31013]_ ;
  assign \new_[30132]_  = ~\new_[30633]_ ;
  assign \new_[30133]_  = ~\new_[31900]_  & ~\new_[6085]_ ;
  assign \new_[30134]_  = ~\new_[31064]_  | ~\new_[30976]_ ;
  assign \new_[30135]_  = ~\new_[31107]_  | ~\new_[4220]_ ;
  assign \new_[30136]_  = ~\new_[30423]_ ;
  assign \new_[30137]_  = ~\new_[31789]_  | ~\new_[5929]_ ;
  assign \new_[30138]_  = ~\new_[31177]_  | ~\new_[4253]_ ;
  assign \new_[30139]_  = ~\new_[30856]_  | ~\new_[4056]_ ;
  assign \new_[30140]_  = ~\new_[31123]_  & ~\new_[4453]_ ;
  assign \new_[30141]_  = ~\new_[31035]_  & ~\new_[4244]_ ;
  assign \new_[30142]_  = ~\new_[30840]_ ;
  assign \new_[30143]_  = ~\new_[31025]_  | ~\new_[30894]_ ;
  assign \new_[30144]_  = ~\new_[31067]_  | ~\new_[6096]_ ;
  assign \new_[30145]_  = ~\new_[30828]_ ;
  assign \new_[30146]_  = ~\new_[30443]_ ;
  assign \new_[30147]_  = ~\new_[31015]_  | ~\new_[4447]_ ;
  assign \new_[30148]_  = ~\new_[30961]_  & ~\new_[4049]_ ;
  assign \new_[30149]_  = ~\new_[30852]_  | ~\new_[4444]_ ;
  assign \new_[30150]_  = \new_[31077]_  | \new_[4207]_ ;
  assign \new_[30151]_  = ~\new_[30635]_ ;
  assign \new_[30152]_  = ~\new_[30743]_ ;
  assign \new_[30153]_  = ~\new_[30822]_ ;
  assign \new_[30154]_  = ~\new_[31652]_  | ~\new_[31121]_ ;
  assign \new_[30155]_  = \new_[30854]_  & \new_[5931]_ ;
  assign \new_[30156]_  = ~\new_[31021]_  & ~\new_[31108]_ ;
  assign \new_[30157]_  = ~\new_[30719]_ ;
  assign \new_[30158]_  = ~\new_[31103]_  | ~\new_[4256]_ ;
  assign \new_[30159]_  = ~\new_[31036]_  | ~\new_[31914]_ ;
  assign \new_[30160]_  = ~\new_[30711]_ ;
  assign \new_[30161]_  = ~\new_[30914]_  | ~\new_[31620]_ ;
  assign \new_[30162]_  = ~\new_[30702]_ ;
  assign \new_[30163]_  = \new_[31041]_  | \new_[4132]_ ;
  assign \new_[30164]_  = ~\new_[31074]_  | ~\new_[4215]_ ;
  assign \new_[30165]_  = \new_[30981]_  | \new_[31763]_ ;
  assign \new_[30166]_  = \new_[31038]_  & \new_[31402]_ ;
  assign \new_[30167]_  = ~\new_[30434]_ ;
  assign \new_[30168]_  = ~\new_[30979]_  & ~\new_[31632]_ ;
  assign \new_[30169]_  = ~\new_[30515]_ ;
  assign \new_[30170]_  = ~\new_[30579]_ ;
  assign \new_[30171]_  = ~\new_[30872]_  | ~\new_[31042]_ ;
  assign \new_[30172]_  = ~\new_[30868]_  | ~\new_[31446]_ ;
  assign \new_[30173]_  = ~\new_[31068]_  & ~\new_[31659]_ ;
  assign \new_[30174]_  = ~\new_[30623]_ ;
  assign \new_[30175]_  = ~\new_[31167]_  & ~\new_[30874]_ ;
  assign \new_[30176]_  = ~\new_[30975]_  & ~\new_[4119]_ ;
  assign \new_[30177]_  = ~\new_[30781]_ ;
  assign \new_[30178]_  = ~\new_[30696]_ ;
  assign \new_[30179]_  = ~\new_[30832]_ ;
  assign \new_[30180]_  = ~\new_[30661]_ ;
  assign \new_[30181]_  = ~\new_[30862]_  & ~\new_[31552]_ ;
  assign \new_[30182]_  = ~\new_[30992]_  & ~\new_[6204]_ ;
  assign \new_[30183]_  = ~\new_[30960]_  | ~\new_[31672]_ ;
  assign \new_[30184]_  = ~\new_[31939]_  | ~\new_[31857]_  | ~\new_[31863]_ ;
  assign \new_[30185]_  = ~\new_[30608]_ ;
  assign \new_[30186]_  = ~\new_[30707]_ ;
  assign \new_[30187]_  = ~\new_[30948]_  | ~\new_[30894]_ ;
  assign \new_[30188]_  = ~\new_[30775]_ ;
  assign \new_[30189]_  = ~\new_[31164]_  & ~\new_[31312]_ ;
  assign \new_[30190]_  = \new_[30864]_  & \new_[5931]_ ;
  assign \new_[30191]_  = \new_[31815]_  | \new_[31102]_ ;
  assign \new_[30192]_  = ~\new_[30857]_  & ~\new_[4075]_ ;
  assign \new_[30193]_  = ~\new_[30867]_  & ~\new_[31401]_ ;
  assign \new_[30194]_  = ~\new_[31182]_  & ~\new_[31039]_ ;
  assign \new_[30195]_  = ~\new_[30985]_  & ~\new_[31312]_ ;
  assign \new_[30196]_  = \new_[30963]_  | \new_[4181]_ ;
  assign \new_[30197]_  = ~\new_[30772]_ ;
  assign \new_[30198]_  = ~\new_[30718]_ ;
  assign \new_[30199]_  = ~\new_[30752]_ ;
  assign \new_[30200]_  = ~\new_[30879]_  & ~\new_[31284]_ ;
  assign \new_[30201]_  = ~\new_[30603]_ ;
  assign \new_[30202]_  = ~\new_[30903]_  & ~\new_[4098]_ ;
  assign \new_[30203]_  = ~\new_[30892]_  & ~\new_[4086]_ ;
  assign \new_[30204]_  = \new_[31048]_  & \new_[4096]_ ;
  assign \new_[30205]_  = ~\new_[30715]_ ;
  assign \new_[30206]_  = ~\new_[31139]_  & ~\new_[31657]_ ;
  assign \new_[30207]_  = ~\new_[30701]_ ;
  assign \new_[30208]_  = ~\new_[30898]_  & ~\new_[4042]_ ;
  assign \new_[30209]_  = \new_[31114]_  & \new_[4132]_ ;
  assign \new_[30210]_  = ~\new_[30741]_ ;
  assign \new_[30211]_  = ~\new_[31083]_  | ~\new_[31748]_ ;
  assign \new_[30212]_  = ~\new_[30900]_  & ~\new_[4248]_ ;
  assign \new_[30213]_  = ~\new_[30835]_ ;
  assign \new_[30214]_  = ~\new_[30876]_  & ~\new_[31658]_ ;
  assign \new_[30215]_  = ~\new_[30888]_  | ~\new_[4225]_ ;
  assign \new_[30216]_  = \new_[30987]_  & \new_[4107]_ ;
  assign \new_[30217]_  = ~\new_[31051]_  | ~\new_[3880]_ ;
  assign \new_[30218]_  = ~\new_[30713]_ ;
  assign \new_[30219]_  = ~\new_[31137]_  & ~\new_[4108]_ ;
  assign \new_[30220]_  = \new_[31115]_  & \new_[5996]_ ;
  assign \new_[30221]_  = ~\new_[31084]_  | ~\new_[4204]_ ;
  assign \new_[30222]_  = ~\new_[30648]_ ;
  assign \new_[30223]_  = ~\new_[30911]_  | ~\new_[31876]_ ;
  assign \new_[30224]_  = ~\new_[30617]_ ;
  assign \new_[30225]_  = ~\new_[30559]_ ;
  assign \new_[30226]_  = \new_[6197]_  & \new_[31596]_ ;
  assign \new_[30227]_  = \new_[31208]_  & \new_[31111]_ ;
  assign \new_[30228]_  = ~\new_[30842]_ ;
  assign \new_[30229]_  = ~\new_[30420]_ ;
  assign \new_[30230]_  = ~\new_[30416]_ ;
  assign \new_[30231]_  = ~\new_[31029]_  & ~\new_[4213]_ ;
  assign \new_[30232]_  = ~\new_[30425]_ ;
  assign \new_[30233]_  = ~\new_[30706]_ ;
  assign \new_[30234]_  = ~\new_[31153]_  & ~\new_[4114]_ ;
  assign \new_[30235]_  = \new_[31133]_  & \new_[4119]_ ;
  assign \new_[30236]_  = \new_[31172]_  & \new_[4079]_ ;
  assign \new_[30237]_  = \new_[30942]_  & \new_[30925]_ ;
  assign \new_[30238]_  = ~\new_[31025]_  | ~\new_[6069]_ ;
  assign \new_[30239]_  = ~\new_[31063]_  & ~\new_[31696]_ ;
  assign \new_[30240]_  = ~\new_[31186]_  & ~\new_[31714]_ ;
  assign \new_[30241]_  = ~\new_[6043]_  & ~\new_[5967]_ ;
  assign \new_[30242]_  = ~\new_[30733]_ ;
  assign \new_[30243]_  = ~\new_[30644]_ ;
  assign \new_[30244]_  = \new_[31124]_  & \new_[4173]_ ;
  assign \new_[30245]_  = ~\new_[30876]_  & ~\new_[4222]_ ;
  assign \new_[30246]_  = ~\new_[30960]_  | ~\new_[4112]_ ;
  assign \new_[30247]_  = \new_[31112]_  & \new_[4116]_ ;
  assign \new_[30248]_  = ~\new_[30737]_ ;
  assign \new_[30249]_  = ~\new_[30964]_  & ~\new_[4089]_ ;
  assign \new_[30250]_  = ~\new_[30628]_ ;
  assign \new_[30251]_  = ~\new_[31046]_  & ~\new_[31889]_ ;
  assign \new_[30252]_  = ~\new_[30770]_ ;
  assign \new_[30253]_  = ~\new_[30767]_ ;
  assign \new_[30254]_  = ~\new_[30782]_ ;
  assign \new_[30255]_  = ~\new_[30757]_ ;
  assign \new_[30256]_  = (~\new_[6042]_  | ~\new_[31497]_ ) & (~\new_[6205]_  | ~\new_[31393]_ );
  assign \new_[30257]_  = ~\new_[30885]_  | ~\new_[31754]_ ;
  assign \new_[30258]_  = ~\new_[30940]_  | ~\new_[31708]_ ;
  assign \new_[30259]_  = ~\new_[31049]_  | ~\new_[6094]_ ;
  assign \new_[30260]_  = ~\new_[30966]_  & ~\new_[31467]_ ;
  assign \new_[30261]_  = ~\new_[31090]_  & ~\new_[31801]_ ;
  assign \new_[30262]_  = ~\new_[30607]_ ;
  assign \new_[30263]_  = ~\new_[30893]_  & ~\new_[5914]_ ;
  assign \new_[30264]_  = \new_[6045]_  | \new_[31569]_ ;
  assign \new_[30265]_  = ~\new_[30725]_ ;
  assign \new_[30266]_  = ~\new_[31171]_  & ~\new_[31731]_ ;
  assign \new_[30267]_  = ~\new_[31154]_  & ~\new_[4255]_ ;
  assign \new_[30268]_  = ~\new_[30967]_  & ~\new_[4088]_ ;
  assign \new_[30269]_  = ~\new_[31190]_  | ~\new_[4271]_ ;
  assign \new_[30270]_  = ~\new_[30971]_  & ~\new_[31743]_ ;
  assign \new_[30271]_  = ~\new_[30708]_ ;
  assign \new_[30272]_  = ~\new_[31125]_  & ~\new_[4445]_ ;
  assign \new_[30273]_  = ~\new_[30600]_ ;
  assign \new_[30274]_  = ~\new_[30609]_ ;
  assign \new_[30275]_  = ~\new_[30494]_ ;
  assign \new_[30276]_  = \new_[31192]_  & \new_[4043]_ ;
  assign \new_[30277]_  = ~\new_[31060]_  & ~\new_[4172]_ ;
  assign \new_[30278]_  = ~\new_[30501]_ ;
  assign \new_[30279]_  = ~\new_[31031]_  | ~\new_[4124]_ ;
  assign \new_[30280]_  = ~\new_[31116]_  | ~\new_[31755]_ ;
  assign \new_[30281]_  = \new_[30996]_  & \new_[30874]_ ;
  assign \new_[30282]_  = ~\new_[31079]_  | ~\new_[31792]_ ;
  assign \new_[30283]_  = ~\new_[30566]_ ;
  assign \new_[30284]_  = \new_[31208]_  & \new_[30939]_ ;
  assign \new_[30285]_  = ~\new_[31069]_  & ~\new_[4223]_ ;
  assign \new_[30286]_  = ~\new_[30627]_ ;
  assign \new_[30287]_  = ~\new_[30763]_ ;
  assign \new_[30288]_  = \new_[30866]_  & \new_[5994]_ ;
  assign \new_[30289]_  = ~\new_[30665]_ ;
  assign \new_[30290]_  = ~\new_[30620]_ ;
  assign \new_[30291]_  = ~\new_[30491]_ ;
  assign \new_[30292]_  = ~\new_[31070]_  & ~\new_[4237]_ ;
  assign \new_[30293]_  = ~\new_[30995]_  | ~\new_[3879]_ ;
  assign \new_[30294]_  = ~\new_[31110]_  | ~\new_[4105]_ ;
  assign \new_[30295]_  = ~\new_[30445]_ ;
  assign \new_[30296]_  = ~\new_[30845]_ ;
  assign \new_[30297]_  = ~\new_[30652]_ ;
  assign \new_[30298]_  = \new_[31189]_  & \new_[31402]_ ;
  assign \new_[30299]_  = ~\new_[31150]_  | ~\new_[31816]_ ;
  assign \new_[30300]_  = ~\new_[30912]_  & ~\new_[31180]_ ;
  assign \new_[30301]_  = \new_[30870]_  & \new_[4116]_ ;
  assign \new_[30302]_  = ~\new_[31169]_  & ~\new_[31771]_ ;
  assign \new_[30303]_  = ~\new_[31064]_  | ~\new_[6033]_ ;
  assign \new_[30304]_  = ~\new_[31052]_  & ~\new_[4239]_ ;
  assign \new_[30305]_  = ~\new_[31044]_  & ~\new_[4043]_ ;
  assign \new_[30306]_  = \new_[31161]_  | \new_[5983]_ ;
  assign \new_[30307]_  = ~\new_[31020]_  & ~\new_[4153]_ ;
  assign \new_[30308]_  = ~\new_[31037]_  & ~\new_[31904]_ ;
  assign \new_[30309]_  = ~\new_[30556]_ ;
  assign \new_[30310]_  = ~\new_[31326]_  | ~\new_[31857]_  | ~\new_[31863]_ ;
  assign \new_[30311]_  = ~\new_[31207]_  & ~\new_[31498]_ ;
  assign \new_[30312]_  = ~\new_[31048]_  | ~\new_[31937]_ ;
  assign \new_[30313]_  = ~\new_[30831]_ ;
  assign \new_[30314]_  = ~\new_[31078]_  & ~\new_[4065]_ ;
  assign \new_[30315]_  = ~\new_[31032]_  & ~\new_[31770]_ ;
  assign \new_[30316]_  = ~\new_[31083]_  | ~\new_[4258]_ ;
  assign \new_[30317]_  = ~\new_[31015]_  | ~\new_[31921]_ ;
  assign \new_[30318]_  = ~\new_[30575]_ ;
  assign \new_[30319]_  = ~\new_[31068]_  & ~\new_[4140]_ ;
  assign \new_[30320]_  = ~\new_[31174]_  | ~\new_[31412]_ ;
  assign \new_[30321]_  = ~\new_[30656]_ ;
  assign \new_[30322]_  = ~\new_[30598]_ ;
  assign \new_[30323]_  = ~\new_[30920]_  & ~\new_[31709]_ ;
  assign \new_[30324]_  = ~\new_[31669]_  & ~\new_[5963]_ ;
  assign \new_[30325]_  = ~\new_[30641]_ ;
  assign \new_[30326]_  = ~\new_[30653]_ ;
  assign \new_[30327]_  = \new_[30868]_  & \new_[4070]_ ;
  assign \new_[30328]_  = ~\new_[31153]_  & ~\new_[31841]_ ;
  assign \new_[30329]_  = ~\new_[30875]_  | ~\new_[4126]_ ;
  assign \new_[30330]_  = \new_[31081]_  | \new_[5924]_ ;
  assign \new_[30331]_  = ~\new_[31024]_  & ~\new_[31834]_ ;
  assign \new_[30332]_  = \new_[31023]_  & \new_[4202]_ ;
  assign \new_[30333]_  = ~\new_[31116]_  | ~\new_[4269]_ ;
  assign \new_[30334]_  = ~\new_[30972]_  & ~\new_[4059]_ ;
  assign \new_[30335]_  = ~\new_[30915]_  & ~\new_[31265]_ ;
  assign \new_[30336]_  = ~\new_[30640]_ ;
  assign \new_[30337]_  = ~\new_[30663]_ ;
  assign \new_[30338]_  = ~\new_[31643]_  & ~\new_[5986]_ ;
  assign \new_[30339]_  = ~\new_[30907]_  & ~\new_[4272]_ ;
  assign \new_[30340]_  = ~\new_[30552]_ ;
  assign \new_[30341]_  = ~\new_[30891]_  & ~\new_[31280]_ ;
  assign \new_[30342]_  = ~\new_[30636]_ ;
  assign \new_[30343]_  = ~\new_[30837]_ ;
  assign \new_[30344]_  = ~\new_[31181]_  | ~\new_[4105]_ ;
  assign \new_[30345]_  = ~\new_[31134]_  & ~\new_[5917]_ ;
  assign \new_[30346]_  = ~\new_[30509]_ ;
  assign \new_[30347]_  = ~\new_[6037]_  | ~\new_[5910]_ ;
  assign \new_[30348]_  = ~\new_[31178]_  & ~\new_[4248]_ ;
  assign \new_[30349]_  = ~\new_[30675]_ ;
  assign \new_[30350]_  = ~\new_[30613]_ ;
  assign \new_[30351]_  = \new_[31741]_  & \new_[6049]_ ;
  assign \new_[30352]_  = ~\new_[30557]_ ;
  assign \new_[30353]_  = ~\new_[6075]_  | ~\new_[31567]_ ;
  assign \new_[30354]_  = ~\new_[30966]_  & ~\new_[30985]_ ;
  assign \new_[30355]_  = \new_[31120]_  & \new_[31613]_ ;
  assign \new_[30356]_  = ~\new_[6074]_  | ~\new_[31707]_ ;
  assign \new_[30357]_  = \new_[30924]_  & \new_[31210]_ ;
  assign \new_[30358]_  = \new_[31126]_  | \new_[5924]_ ;
  assign \new_[30359]_  = ~\new_[6211]_  & ~\new_[31777]_ ;
  assign \new_[30360]_  = \new_[6186]_  & \new_[31901]_ ;
  assign \new_[30361]_  = ~\new_[31232]_  | ~\new_[31906]_ ;
  assign \new_[30362]_  = ~\new_[31862]_  | ~\new_[6000]_ ;
  assign \new_[30363]_  = \new_[31071]_  | \new_[4179]_ ;
  assign \new_[30364]_  = ~\new_[31553]_  | ~\new_[5998]_ ;
  assign \new_[30365]_  = ~\new_[6193]_  | ~\new_[31686]_ ;
  assign \new_[30366]_  = ~\new_[31819]_  | ~\new_[5922]_ ;
  assign \new_[30367]_  = ~\new_[30755]_ ;
  assign \new_[30368]_  = ~\new_[31617]_  | ~\new_[5966]_ ;
  assign \new_[30369]_  = ~\new_[30953]_  & ~\new_[31042]_ ;
  assign \new_[30370]_  = ~\new_[6087]_  & ~\new_[31128]_ ;
  assign \new_[30371]_  = \new_[6036]_  | \new_[31800]_ ;
  assign \new_[30372]_  = \new_[31837]_  & \new_[5990]_ ;
  assign \new_[30373]_  = ~\new_[30518]_ ;
  assign \new_[30374]_  = ~\new_[30512]_ ;
  assign \new_[30375]_  = ~\new_[30667]_ ;
  assign \new_[30376]_  = ~\new_[30861]_  & ~\m3_addr_i[29] ;
  assign \new_[30377]_  = ~\new_[30456]_ ;
  assign \new_[30378]_  = ~\new_[31900]_  | ~\new_[6085]_ ;
  assign \new_[30379]_  = ~\new_[31643]_  | ~\new_[5986]_ ;
  assign \new_[30380]_  = \new_[6093]_  & \new_[31776]_ ;
  assign \new_[30381]_  = \new_[31184]_  | \new_[4242]_ ;
  assign \new_[30382]_  = \new_[6087]_  & \new_[31128]_ ;
  assign \new_[30383]_  = ~\new_[31608]_  & ~\new_[5980]_ ;
  assign \new_[30384]_  = ~\new_[30495]_ ;
  assign \new_[30385]_  = ~\new_[31683]_  | ~\new_[6005]_ ;
  assign \new_[30386]_  = \new_[30972]_  | \new_[31646]_ ;
  assign \new_[30387]_  = ~\new_[30570]_ ;
  assign \new_[30388]_  = ~\new_[30500]_ ;
  assign \new_[30389]_  = ~\new_[30955]_  & ~\new_[4081]_ ;
  assign \new_[30390]_  = ~\new_[31052]_  & ~\new_[31898]_ ;
  assign \new_[30391]_  = ~\new_[31394]_  | ~\new_[5976]_ ;
  assign \new_[30392]_  = ~\new_[6080]_  | ~\new_[31765]_ ;
  assign \new_[30393]_  = ~\new_[30847]_ ;
  assign \new_[30394]_  = ~\new_[30753]_ ;
  assign \new_[30395]_  = \new_[6043]_  & \new_[5967]_ ;
  assign \new_[30396]_  = ~\new_[30514]_ ;
  assign \new_[30397]_  = ~\new_[30547]_ ;
  assign \new_[30398]_  = ~\new_[30714]_ ;
  assign \new_[30399]_  = ~\new_[30983]_  & ~\new_[4278]_ ;
  assign \new_[30400]_  = ~\new_[31127]_  & ~\new_[31813]_ ;
  assign \new_[30401]_  = ~\new_[6079]_  & ~\new_[6270]_ ;
  assign \new_[30402]_  = ~\new_[30561]_ ;
  assign \new_[30403]_  = ~\new_[30992]_  & ~\new_[30993]_ ;
  assign \new_[30404]_  = ~\new_[30881]_  & ~\new_[31891]_ ;
  assign \new_[30405]_  = \new_[6075]_  | \new_[31567]_ ;
  assign \new_[30406]_  = \new_[31202]_  | \new_[6094]_ ;
  assign \new_[30407]_  = ~\new_[31137]_  & ~\new_[31814]_ ;
  assign \new_[30408]_  = \new_[30942]_  & \new_[5830]_ ;
  assign \new_[30409]_  = ~\new_[31009]_  | ~\new_[31897]_ ;
  assign \new_[30410]_  = ~\new_[30762]_ ;
  assign \new_[30411]_  = ~\new_[31080]_  | ~\new_[4274]_ ;
  assign \new_[30412]_  = ~\new_[30883]_  & ~\new_[5914]_ ;
  assign \new_[30413]_  = \new_[31073]_  & \new_[4135]_ ;
  assign \new_[30414]_  = ~\new_[30601]_ ;
  assign \new_[30415]_  = ~\new_[31129]_  & ~\new_[4061]_ ;
  assign \new_[30416]_  = ~\new_[31480]_  | ~\new_[31710]_ ;
  assign \new_[30417]_  = ~\new_[6214]_  | ~\new_[6192]_ ;
  assign \new_[30418]_  = \new_[6191]_  | \new_[6070]_ ;
  assign \new_[30419]_  = ~\new_[4217]_  | ~n8339;
  assign \new_[30420]_  = \new_[31214]_  & \new_[4227]_ ;
  assign \new_[30421]_  = ~\new_[6082]_  | ~\new_[6085]_ ;
  assign \new_[30422]_  = ~\new_[31538]_  & ~\m1_addr_i[28] ;
  assign \new_[30423]_  = ~\new_[31311]_  & ~\new_[4148]_ ;
  assign \new_[30424]_  = \new_[6174]_  | \new_[6034]_ ;
  assign \new_[30425]_  = ~\new_[31418]_  & ~\new_[31580]_ ;
  assign \new_[30426]_  = \new_[31439]_  | \new_[31918]_ ;
  assign \new_[30427]_  = ~\new_[4250]_  | ~n8364;
  assign \new_[30428]_  = ~\new_[6185]_  | ~\new_[6000]_ ;
  assign \new_[30429]_  = ~\new_[31274]_  & ~\new_[31546]_ ;
  assign \new_[30430]_  = ~\new_[30864]_ ;
  assign \new_[30431]_  = ~\new_[6056]_  & ~\new_[5900]_ ;
  assign \new_[30432]_  = ~\new_[31507]_  | ~\new_[3888]_ ;
  assign \new_[30433]_  = ~\new_[31175]_ ;
  assign \new_[30434]_  = ~\new_[31324]_  | ~\new_[3884]_ ;
  assign \new_[30435]_  = ~\new_[6086]_  | ~\new_[5929]_ ;
  assign \new_[30436]_  = ~\new_[31049]_ ;
  assign \new_[30437]_  = \new_[31218]_  | \new_[31755]_ ;
  assign \new_[30438]_  = \new_[31449]_  & \new_[4156]_ ;
  assign \new_[30439]_  = ~\new_[30867]_ ;
  assign \new_[30440]_  = ~\new_[31362]_  | ~\new_[6090]_ ;
  assign \new_[30441]_  = \new_[6202]_  | \new_[31474]_ ;
  assign \new_[30442]_  = ~\new_[31436]_  & ~\new_[4038]_ ;
  assign \new_[30443]_  = \new_[31391]_  & \new_[31897]_ ;
  assign \new_[30444]_  = ~\new_[31338]_  | ~\new_[31806]_ ;
  assign \new_[30445]_  = ~\new_[31323]_  & ~\new_[4451]_ ;
  assign \new_[30446]_  = ~\new_[31500]_  | ~\new_[4098]_ ;
  assign \new_[30447]_  = ~\new_[31297]_  | ~\new_[5914]_ ;
  assign \new_[30448]_  = ~\new_[31081]_ ;
  assign \new_[30449]_  = ~\new_[31134]_ ;
  assign \new_[30450]_  = ~\new_[31003]_ ;
  assign \new_[30451]_  = ~\new_[6075]_  & ~\new_[5905]_ ;
  assign \new_[30452]_  = ~\new_[31070]_ ;
  assign \new_[30453]_  = ~\new_[31863]_  | ~\new_[6449]_ ;
  assign \new_[30454]_  = ~\m7_addr_i[29]  | ~\m7_addr_i[28] ;
  assign \new_[30455]_  = ~\new_[30938]_ ;
  assign \new_[30456]_  = \new_[6079]_  | \new_[31548]_ ;
  assign \new_[30457]_  = ~\new_[31253]_  & ~\new_[31490]_ ;
  assign \new_[30458]_  = ~\new_[31058]_ ;
  assign \new_[30459]_  = ~\new_[6079]_  | ~\new_[31548]_ ;
  assign \new_[30460]_  = ~\new_[30889]_ ;
  assign \new_[30461]_  = \new_[6195]_  & \new_[6060]_ ;
  assign \new_[30462]_  = ~\new_[30966]_ ;
  assign \new_[30463]_  = ~\new_[30893]_ ;
  assign \new_[30464]_  = ~\new_[30903]_ ;
  assign \new_[30465]_  = ~\new_[31168]_ ;
  assign \new_[30466]_  = \new_[31484]_  & \new_[4260]_ ;
  assign \new_[30467]_  = ~\new_[31470]_  | ~\new_[3886]_ ;
  assign \new_[30468]_  = ~\new_[31162]_ ;
  assign \new_[30469]_  = ~\new_[31312]_  & ~\new_[31467]_ ;
  assign \new_[30470]_  = ~\new_[30907]_ ;
  assign \new_[30471]_  = ~\new_[30922]_ ;
  assign \new_[30472]_  = ~\new_[5972]_  | ~\new_[31431]_ ;
  assign \new_[30473]_  = ~\new_[31521]_  & ~\new_[6088]_ ;
  assign \new_[30474]_  = ~\new_[6062]_  & ~\new_[5901]_ ;
  assign \new_[30475]_  = ~\new_[30980]_ ;
  assign \new_[30476]_  = ~\new_[31154]_ ;
  assign \new_[30477]_  = ~\new_[31940]_  | ~\new_[31326]_ ;
  assign \new_[30478]_  = ~\new_[31219]_  & ~\new_[4121]_ ;
  assign \new_[30479]_  = ~\new_[30918]_ ;
  assign \new_[30480]_  = ~\new_[6091]_  & ~\new_[31383]_ ;
  assign \new_[30481]_  = ~\new_[31280]_  & ~\new_[31398]_ ;
  assign \new_[30482]_  = ~\new_[31035]_ ;
  assign \new_[30483]_  = \new_[31231]_  & n8404;
  assign \new_[30484]_  = s6_m4_cyc_r_reg;
  assign \new_[30485]_  = s15_m6_cyc_r_reg;
  assign \new_[30486]_  = s8_m2_cyc_r_reg;
  assign \new_[30487]_  = s5_m5_cyc_r_reg;
  assign \new_[30488]_  = s13_m5_cyc_r_reg;
  assign \new_[30489]_  = ~\new_[6440]_  & ~\new_[6449]_ ;
  assign \new_[30490]_  = s3_m5_cyc_r_reg;
  assign \new_[30491]_  = ~\new_[31540]_  | ~\new_[4235]_ ;
  assign \new_[30492]_  = ~\new_[6063]_  & ~\new_[5982]_ ;
  assign \new_[30493]_  = ~\new_[6211]_  & ~\new_[6061]_ ;
  assign \new_[30494]_  = ~\new_[31269]_  | ~\new_[31641]_ ;
  assign \new_[30495]_  = ~\new_[6211]_  | ~\new_[6061]_ ;
  assign \new_[30496]_  = ~\new_[31863]_  | ~\new_[7224]_ ;
  assign \new_[30497]_  = \new_[31465]_  | \new_[31731]_ ;
  assign \new_[30498]_  = ~\new_[6058]_  | ~\new_[5980]_ ;
  assign \new_[30499]_  = \new_[31293]_  | \new_[4094]_ ;
  assign \new_[30500]_  = \new_[6041]_  & \new_[5966]_ ;
  assign \new_[30501]_  = ~\new_[31426]_  & ~\new_[4170]_ ;
  assign \new_[30502]_  = ~\new_[31331]_  & ~\new_[31909]_ ;
  assign \new_[30503]_  = ~\new_[31205]_ ;
  assign \new_[30504]_  = ~\new_[31087]_ ;
  assign \new_[30505]_  = \new_[31358]_  | \new_[4075]_ ;
  assign \new_[30506]_  = ~\new_[31207]_ ;
  assign \new_[30507]_  = \new_[31483]_  | \new_[31801]_ ;
  assign \new_[30508]_  = \new_[31245]_  | \new_[31717]_ ;
  assign \new_[30509]_  = \new_[4230]_  & n8464;
  assign \new_[30510]_  = ~\new_[31122]_ ;
  assign \new_[30511]_  = ~\new_[30993]_ ;
  assign \new_[30512]_  = \new_[6035]_  & \new_[5963]_ ;
  assign \new_[30513]_  = ~\new_[31214]_  | ~\new_[31590]_ ;
  assign \new_[30514]_  = ~\new_[31499]_  & ~\new_[6215]_ ;
  assign \new_[30515]_  = ~\new_[31341]_  & ~\new_[4116]_ ;
  assign \new_[30516]_  = ~\new_[31863]_  | ~\new_[7440]_ ;
  assign \new_[30517]_  = ~\new_[31126]_ ;
  assign \new_[30518]_  = \new_[6037]_  | \new_[31506]_ ;
  assign \new_[30519]_  = ~\new_[31476]_  | ~\new_[31876]_ ;
  assign \new_[30520]_  = ~\new_[6086]_  & ~\new_[5929]_ ;
  assign \new_[30521]_  = ~\new_[31549]_  & ~\new_[4042]_ ;
  assign \new_[30522]_  = ~\new_[30964]_ ;
  assign \new_[30523]_  = ~\new_[30890]_ ;
  assign \new_[30524]_  = ~\new_[30892]_ ;
  assign \new_[30525]_  = ~\new_[31404]_  | ~\new_[4079]_ ;
  assign \new_[30526]_  = ~\new_[31396]_  & ~\new_[4126]_ ;
  assign \new_[30527]_  = ~\new_[6091]_  | ~\new_[31383]_ ;
  assign \new_[30528]_  = ~\new_[31166]_ ;
  assign \new_[30529]_  = ~\new_[31408]_  | ~\new_[5920]_ ;
  assign \new_[30530]_  = ~\new_[4069]_  | ~n8324;
  assign \new_[30531]_  = ~\new_[30905]_ ;
  assign \new_[30532]_  = ~\new_[31041]_ ;
  assign \new_[30533]_  = ~\new_[31160]_ ;
  assign \new_[30534]_  = ~\new_[31161]_ ;
  assign \new_[30535]_  = ~\new_[31044]_ ;
  assign \new_[30536]_  = ~\new_[31292]_  & ~\new_[31485]_ ;
  assign \new_[30537]_  = ~\new_[31146]_ ;
  assign \new_[30538]_  = ~\new_[31541]_  | ~\new_[4242]_ ;
  assign \new_[30539]_  = ~\new_[30909]_ ;
  assign \new_[30540]_  = ~\new_[31414]_  & ~\new_[4206]_ ;
  assign \new_[30541]_  = \new_[31388]_  & \new_[4213]_ ;
  assign \new_[30542]_  = ~\new_[31405]_  & ~\new_[4084]_ ;
  assign \new_[30543]_  = ~\new_[31305]_  & ~\new_[4442]_ ;
  assign \new_[30544]_  = ~\new_[31338]_  | ~\new_[4267]_ ;
  assign \new_[30545]_  = \new_[31278]_  & \new_[31769]_ ;
  assign \new_[30546]_  = s1_m1_cyc_r_reg;
  assign \new_[30547]_  = ~\new_[6195]_  & ~\new_[6060]_ ;
  assign \new_[30548]_  = s11_m5_cyc_r_reg;
  assign \new_[30549]_  = s12_m5_cyc_r_reg;
  assign \new_[30550]_  = \new_[31215]_  | \new_[31632]_ ;
  assign \new_[30551]_  = ~\new_[6042]_  & ~\new_[5896]_ ;
  assign \new_[30552]_  = ~\new_[31271]_  | ~\new_[3875]_ ;
  assign \new_[30553]_  = ~\new_[31425]_  & ~\new_[31904]_ ;
  assign \new_[30554]_  = ~\new_[31430]_  | ~\new_[4142]_ ;
  assign \new_[30555]_  = ~\new_[31324]_  | ~\new_[31709]_ ;
  assign \new_[30556]_  = ~\new_[31266]_  | ~\new_[31605]_ ;
  assign \new_[30557]_  = ~\new_[31304]_  & ~\new_[4272]_ ;
  assign \new_[30558]_  = \new_[31400]_  & \new_[6070]_ ;
  assign \new_[30559]_  = \new_[31457]_  | \new_[4280]_ ;
  assign \new_[30560]_  = ~\new_[6041]_  & ~\new_[5966]_ ;
  assign \new_[30561]_  = ~\new_[6045]_  & ~\new_[5897]_ ;
  assign \new_[30562]_  = ~\m4_addr_i[29]  & ~\m4_addr_i[28] ;
  assign \new_[30563]_  = \new_[31257]_  | \new_[4258]_ ;
  assign \new_[30564]_  = ~\new_[31478]_  & ~\new_[4096]_ ;
  assign \new_[30565]_  = ~\new_[31202]_ ;
  assign \new_[30566]_  = \new_[31315]_  & \new_[31556]_ ;
  assign \new_[30567]_  = ~\new_[6095]_  | ~\new_[6217]_ ;
  assign \new_[30568]_  = ~\new_[31275]_  & ~\new_[4107]_ ;
  assign \new_[30569]_  = ~\new_[31311]_  & ~\new_[31771]_ ;
  assign \new_[30570]_  = ~\new_[31100]_ ;
  assign \new_[30571]_  = ~\new_[31310]_  | ~\new_[31856]_ ;
  assign \new_[30572]_  = ~\new_[31540]_  | ~\new_[31932]_ ;
  assign \new_[30573]_  = \new_[31332]_  | \new_[4077]_ ;
  assign \new_[30574]_  = ~\new_[31217]_  | ~\new_[4128]_ ;
  assign \new_[30575]_  = ~\new_[31512]_  & ~\new_[4056]_ ;
  assign \new_[30576]_  = ~\new_[30854]_ ;
  assign \new_[30577]_  = ~\new_[31894]_ ;
  assign \new_[30578]_  = ~\new_[31281]_  | ~\new_[31656]_ ;
  assign \new_[30579]_  = ~\new_[31270]_  | ~\new_[4172]_ ;
  assign \new_[30580]_  = ~\new_[4439]_  | ~n8369;
  assign \new_[30581]_  = ~\new_[31493]_  & ~\new_[4239]_ ;
  assign \new_[30582]_  = ~\new_[31225]_  | ~\new_[4209]_ ;
  assign \new_[30583]_  = ~\new_[3881]_  | ~n8349;
  assign \new_[30584]_  = ~\new_[31435]_  & ~\new_[31620]_ ;
  assign \new_[30585]_  = ~\new_[6080]_  | ~\new_[5933]_ ;
  assign \new_[30586]_  = \new_[31268]_  | \new_[4045]_ ;
  assign \new_[30587]_  = ~\new_[7222]_  & ~\new_[7917]_ ;
  assign \new_[30588]_  = ~\new_[6036]_  & ~\new_[5895]_ ;
  assign \new_[30589]_  = ~\new_[31384]_  | ~n8759;
  assign \new_[30590]_  = ~\new_[6784]_  & ~\new_[7440]_ ;
  assign \new_[30591]_  = ~\new_[31432]_  & ~\new_[4444]_ ;
  assign \new_[30592]_  = \m6_addr_i[31]  & \m6_addr_i[30] ;
  assign \new_[30593]_  = ~\new_[31195]_ ;
  assign \new_[30594]_  = \new_[6073]_  & \new_[5989]_ ;
  assign \new_[30595]_  = \new_[31267]_  | \new_[31659]_ ;
  assign \new_[30596]_  = ~\new_[31778]_  | ~\new_[31938]_ ;
  assign \new_[30597]_  = ~\new_[31444]_  & ~\new_[3879]_ ;
  assign \new_[30598]_  = \new_[31501]_  & \new_[31850]_ ;
  assign \new_[30599]_  = ~\new_[31250]_  | ~\new_[4130]_ ;
  assign \new_[30600]_  = \new_[31347]_  | \new_[31916]_ ;
  assign \new_[30601]_  = ~\new_[6189]_  & ~\new_[5990]_ ;
  assign \new_[30602]_  = ~\new_[31410]_  | ~\new_[5987]_ ;
  assign \new_[30603]_  = \new_[31331]_  | \new_[4278]_ ;
  assign \new_[30604]_  = ~\new_[31320]_  | ~\new_[4058]_ ;
  assign \new_[30605]_  = \new_[31551]_  | \new_[6046]_ ;
  assign \new_[30606]_  = ~\new_[30946]_ ;
  assign \new_[30607]_  = ~\new_[31273]_  & ~\new_[4043]_ ;
  assign \new_[30608]_  = ~\new_[31507]_  | ~\new_[31743]_ ;
  assign \new_[30609]_  = ~\new_[6047]_  & ~\new_[5971]_ ;
  assign \new_[30610]_  = \new_[31257]_  | \new_[31748]_ ;
  assign \new_[30611]_  = ~\new_[31199]_ ;
  assign \new_[30612]_  = \new_[31443]_  & \new_[31880]_ ;
  assign \new_[30613]_  = ~\new_[31430]_  | ~\new_[31629]_ ;
  assign \new_[30614]_  = ~\new_[31863]_  | ~\new_[6791]_ ;
  assign \new_[30615]_  = ~\new_[31415]_  | ~\new_[4112]_ ;
  assign \new_[30616]_  = ~\new_[31335]_  & ~\new_[4089]_ ;
  assign \new_[30617]_  = ~\new_[31505]_  | ~\new_[3880]_ ;
  assign \new_[30618]_  = \new_[31351]_  & \new_[31696]_ ;
  assign \new_[30619]_  = ~\new_[31047]_ ;
  assign \new_[30620]_  = ~\new_[31461]_  & ~\new_[4175]_ ;
  assign \new_[30621]_  = ~\new_[31362]_  & ~\new_[6090]_ ;
  assign \new_[30622]_  = \new_[6199]_  & \new_[5970]_ ;
  assign \new_[30623]_  = \new_[31309]_  | \new_[4081]_ ;
  assign \new_[30624]_  = ~s15_m1_cyc_r_reg;
  assign \new_[30625]_  = ~\new_[6375]_  & ~\new_[6791]_ ;
  assign \new_[30626]_  = ~\new_[31280]_  & ~\new_[31502]_ ;
  assign \new_[30627]_  = ~\new_[31476]_  | ~\new_[4110]_ ;
  assign \new_[30628]_  = ~\new_[31427]_  | ~\new_[4103]_ ;
  assign \new_[30629]_  = \new_[31320]_  & \new_[31838]_ ;
  assign \new_[30630]_  = ~\new_[31509]_  | ~\new_[31681]_ ;
  assign \new_[30631]_  = s15_m3_cyc_r_reg;
  assign \new_[30632]_  = ~\new_[31267]_  & ~\new_[4140]_ ;
  assign \new_[30633]_  = ~\new_[31445]_  & ~\new_[4061]_ ;
  assign \new_[30634]_  = \new_[6063]_  & \new_[5982]_ ;
  assign \new_[30635]_  = \new_[31409]_  | \new_[4179]_ ;
  assign \new_[30636]_  = ~\new_[31375]_  | ~\new_[4124]_ ;
  assign \new_[30637]_  = ~\new_[31302]_  & ~\new_[4256]_ ;
  assign \new_[30638]_  = ~\new_[31250]_  | ~\new_[31889]_ ;
  assign \new_[30639]_  = ~\new_[6035]_  & ~\new_[5963]_ ;
  assign \new_[30640]_  = ~\new_[31404]_  | ~\new_[31679]_ ;
  assign \new_[30641]_  = \new_[31301]_  | \new_[4049]_ ;
  assign \new_[30642]_  = ~\new_[31353]_  & ~\new_[4271]_ ;
  assign \new_[30643]_  = ~\new_[6185]_  & ~\new_[6000]_ ;
  assign \new_[30644]_  = \new_[31351]_  & \new_[4139]_ ;
  assign \new_[30645]_  = ~\new_[31375]_  | ~\new_[31587]_ ;
  assign \new_[30646]_  = ~\new_[6087]_  | ~\new_[5907]_ ;
  assign \new_[30647]_  = ~\new_[31541]_  | ~\new_[31713]_ ;
  assign \new_[30648]_  = \new_[31319]_  & \new_[4065]_ ;
  assign \new_[30649]_  = ~\new_[31475]_  & ~\new_[4088]_ ;
  assign \new_[30650]_  = \new_[31215]_  | \new_[4067]_ ;
  assign \new_[30651]_  = ~\new_[31545]_  & ~\new_[4132]_ ;
  assign \new_[30652]_  = \new_[31310]_  & \new_[4449]_ ;
  assign \new_[30653]_  = \new_[31425]_  | \new_[4146]_ ;
  assign \new_[30654]_  = ~\new_[30968]_ ;
  assign \new_[30655]_  = ~\new_[6043]_  | ~\new_[31397]_ ;
  assign \new_[30656]_  = \new_[31449]_  & \new_[31714]_ ;
  assign \new_[30657]_  = ~\new_[6044]_  | ~\new_[5969]_ ;
  assign \new_[30658]_  = ~\new_[31053]_ ;
  assign \new_[30659]_  = ~\new_[31129]_ ;
  assign \new_[30660]_  = ~\new_[31469]_  & ~\new_[4222]_ ;
  assign \new_[30661]_  = ~\new_[31536]_  & ~\new_[4153]_ ;
  assign \new_[30662]_  = ~\new_[31420]_  & ~\new_[4255]_ ;
  assign \new_[30663]_  = ~\new_[31418]_  & ~\new_[4223]_ ;
  assign \new_[30664]_  = ~\new_[6082]_  & ~\new_[6085]_ ;
  assign \new_[30665]_  = \new_[31424]_  | \new_[31646]_ ;
  assign \new_[30666]_  = ~\new_[31062]_ ;
  assign \new_[30667]_  = ~\new_[31306]_  | ~\new_[31854]_ ;
  assign \new_[30668]_  = ~\new_[31408]_  & ~\new_[5920]_ ;
  assign \new_[30669]_  = ~\new_[31863]_  | ~\new_[6782]_ ;
  assign \new_[30670]_  = ~\new_[31356]_  | ~\new_[31571]_ ;
  assign \new_[30671]_  = ~\new_[5992]_  & ~\new_[5922]_ ;
  assign \new_[30672]_  = \new_[31456]_  & n8809;
  assign \new_[30673]_  = ~\new_[31551]_  | ~\new_[6046]_ ;
  assign \new_[30674]_  = ~\new_[30951]_ ;
  assign \new_[30675]_  = ~\new_[31489]_  & ~\new_[4105]_ ;
  assign \new_[30676]_  = \new_[31260]_  | \new_[4063]_ ;
  assign \new_[30677]_  = \new_[31270]_  & \new_[31727]_ ;
  assign \new_[30678]_  = ~\new_[31319]_  | ~\new_[31852]_ ;
  assign \new_[30679]_  = ~\new_[31018]_ ;
  assign \new_[30680]_  = ~\new_[31256]_  | ~\new_[31911]_ ;
  assign \new_[30681]_  = ~\new_[30871]_ ;
  assign \new_[30682]_  = ~\new_[31254]_  & ~\new_[4173]_ ;
  assign \new_[30683]_  = ~\new_[31294]_  | ~n8554;
  assign \new_[30684]_  = ~\new_[31347]_  & ~\new_[4240]_ ;
  assign \new_[30685]_  = ~\new_[31082]_ ;
  assign \new_[30686]_  = ~\new_[31470]_  | ~\new_[31613]_ ;
  assign \new_[30687]_  = ~\new_[30941]_ ;
  assign \new_[30688]_  = ~\new_[31264]_  & ~\new_[4108]_ ;
  assign \new_[30689]_  = ~\new_[5992]_  | ~\new_[5922]_ ;
  assign \new_[30690]_  = ~\new_[31185]_ ;
  assign \new_[30691]_  = ~\new_[31378]_  | ~\new_[31841]_ ;
  assign \new_[30692]_  = ~\new_[4157]_  | ~n8874;
  assign \new_[30693]_  = ~\new_[31306]_  | ~\new_[4244]_ ;
  assign \new_[30694]_  = ~\new_[31272]_  & ~\new_[4220]_ ;
  assign \new_[30695]_  = ~\new_[31329]_  | ~\new_[31566]_ ;
  assign \new_[30696]_  = ~\new_[31350]_  & ~\new_[4137]_ ;
  assign \new_[30697]_  = ~\new_[31271]_  | ~\new_[31834]_ ;
  assign \new_[30698]_  = ~\new_[6068]_  & ~\new_[5986]_ ;
  assign \new_[30699]_  = ~\new_[31521]_  | ~\new_[6088]_ ;
  assign \new_[30700]_  = \new_[31240]_  & n8439;
  assign \new_[30701]_  = \new_[31391]_  & \new_[3877]_ ;
  assign \new_[30702]_  = \new_[31302]_  | \new_[31649]_ ;
  assign \new_[30703]_  = ~\new_[31226]_  & ~\new_[4123]_ ;
  assign \new_[30704]_  = ~\new_[6439]_  & ~\new_[6794]_ ;
  assign \new_[30705]_  = ~\new_[30853]_ ;
  assign \new_[30706]_  = ~\new_[31301]_  & ~\new_[31886]_ ;
  assign \new_[30707]_  = ~\new_[31454]_  | ~\new_[4447]_ ;
  assign \new_[30708]_  = ~\new_[31435]_  & ~\new_[4051]_ ;
  assign \new_[30709]_  = ~\new_[31398]_  & ~\new_[31401]_ ;
  assign \new_[30710]_  = ~\new_[31460]_  & ~\new_[4155]_ ;
  assign \new_[30711]_  = ~\new_[31514]_  & ~\new_[4086]_ ;
  assign \new_[30712]_  = \m4_addr_i[31]  & \m4_addr_i[30] ;
  assign \new_[30713]_  = ~\new_[31218]_  & ~\new_[4269]_ ;
  assign \new_[30714]_  = ~\new_[6199]_  & ~\new_[5970]_ ;
  assign \new_[30715]_  = ~\new_[31461]_  & ~\new_[31558]_ ;
  assign \new_[30716]_  = ~\new_[4134]_  | ~n8329;
  assign \new_[30717]_  = ~\new_[31427]_  | ~\new_[31744]_ ;
  assign \new_[30718]_  = \new_[31378]_  & \new_[4114]_ ;
  assign \new_[30719]_  = \new_[31483]_  | \new_[4276]_ ;
  assign \new_[30720]_  = ~\new_[6087]_  & ~\new_[5907]_ ;
  assign \new_[30721]_  = \new_[31332]_  | \new_[31792]_ ;
  assign \new_[30722]_  = ~\new_[6203]_  | ~\new_[6245]_ ;
  assign \new_[30723]_  = \new_[31457]_  | \new_[31627]_ ;
  assign \new_[30724]_  = ~\new_[31278]_  | ~\new_[4040]_ ;
  assign \new_[30725]_  = ~\new_[31454]_  | ~\new_[31921]_ ;
  assign \new_[30726]_  = ~\new_[31480]_  | ~\new_[4211]_ ;
  assign \new_[30727]_  = \new_[31252]_  | \new_[31811]_ ;
  assign \new_[30728]_  = ~\new_[31505]_  | ~\new_[31867]_ ;
  assign \new_[30729]_  = ~\new_[30865]_ ;
  assign \new_[30730]_  = ~\new_[31443]_  | ~\new_[4204]_ ;
  assign \new_[30731]_  = \new_[31465]_  | \new_[4090]_ ;
  assign \new_[30732]_  = \new_[31535]_  & \new_[4168]_ ;
  assign \new_[30733]_  = ~\new_[31293]_  & ~\new_[31657]_ ;
  assign \new_[30734]_  = \new_[6073]_  | \new_[5989]_ ;
  assign \new_[30735]_  = \new_[31436]_  | \new_[31702]_ ;
  assign \new_[30736]_  = \new_[31315]_  & \new_[4207]_ ;
  assign \new_[30737]_  = ~\new_[31409]_  & ~\new_[31601]_ ;
  assign \new_[30738]_  = ~\new_[6783]_  & ~\new_[7915]_ ;
  assign \new_[30739]_  = \new_[4150]_  & n8319;
  assign \new_[30740]_  = ~\new_[6058]_  & ~\new_[5980]_ ;
  assign \new_[30741]_  = \new_[31256]_  & \new_[4164]_ ;
  assign \new_[30742]_  = ~\new_[31227]_  | ~\new_[5917]_ ;
  assign \new_[30743]_  = ~\new_[31504]_  & ~\new_[4202]_ ;
  assign \new_[30744]_  = ~\new_[31193]_ ;
  assign \new_[30745]_  = ~\m6_addr_i[29]  & ~\m6_addr_i[28] ;
  assign \new_[30746]_  = \new_[31356]_  & \new_[4246]_ ;
  assign \new_[30747]_  = ~\new_[31424]_  & ~\new_[4059]_ ;
  assign \new_[30748]_  = ~\new_[6068]_  | ~\new_[5986]_ ;
  assign \new_[30749]_  = ~\new_[31061]_ ;
  assign \new_[30750]_  = \new_[31260]_  | \new_[31891]_ ;
  assign \new_[30751]_  = ~\new_[31281]_  | ~\new_[4264]_ ;
  assign \new_[30752]_  = ~\new_[31415]_  | ~\new_[31672]_ ;
  assign \new_[30753]_  = ~\new_[6074]_  & ~\new_[5904]_ ;
  assign \new_[30754]_  = \new_[31245]_  | \new_[4225]_ ;
  assign \new_[30755]_  = ~\new_[31252]_  & ~\new_[4274]_ ;
  assign \new_[30756]_  = ~\new_[31138]_ ;
  assign \new_[30757]_  = ~\new_[31358]_  & ~\new_[31823]_ ;
  assign \new_[30758]_  = ~\new_[6214]_  & ~\new_[6192]_ ;
  assign \new_[30759]_  = ~\new_[6203]_  & ~\new_[6245]_ ;
  assign \new_[30760]_  = ~\new_[6273]_  | ~\new_[6065]_ ;
  assign \new_[30761]_  = ~\new_[31196]_ ;
  assign \new_[30762]_  = ~\new_[31309]_  & ~\new_[31802]_ ;
  assign \new_[30763]_  = \new_[31439]_  | \new_[4229]_ ;
  assign \new_[30764]_  = \new_[31268]_  | \new_[31768]_ ;
  assign \new_[30765]_  = \new_[31488]_  | \new_[31708]_ ;
  assign \new_[30766]_  = ~\new_[4053]_  | ~n8344;
  assign \new_[30767]_  = ~\new_[31500]_  | ~\new_[31618]_ ;
  assign \new_[30768]_  = ~\new_[6044]_  & ~\new_[5969]_ ;
  assign \new_[30769]_  = ~\new_[31544]_  & ~\new_[4072]_ ;
  assign \new_[30770]_  = ~\new_[6062]_  | ~\new_[5901]_ ;
  assign \new_[30771]_  = \new_[31266]_  & \new_[4181]_ ;
  assign \new_[30772]_  = ~\new_[5898]_  | ~\new_[6051]_ ;
  assign \new_[30773]_  = \new_[6174]_  & \new_[6034]_ ;
  assign \new_[30774]_  = ~\new_[31329]_  | ~\new_[4092]_ ;
  assign \new_[30775]_  = ~\new_[31346]_  | ~\new_[31604]_ ;
  assign \new_[30776]_  = ~\new_[6200]_  & ~\new_[6048]_ ;
  assign \new_[30777]_  = s10_m4_cyc_r_reg;
  assign \new_[30778]_  = ~\new_[30924]_ ;
  assign \new_[30779]_  = ~\new_[30921]_ ;
  assign \new_[30780]_  = ~\new_[31300]_  & ~\new_[4237]_ ;
  assign \new_[30781]_  = ~\new_[6076]_  | ~\new_[5925]_ ;
  assign \new_[30782]_  = ~\new_[31217]_  | ~\new_[31899]_ ;
  assign \new_[30783]_  = ~\new_[6268]_  | ~\new_[5995]_ ;
  assign \new_[30784]_  = ~\new_[31346]_  | ~\new_[4160]_ ;
  assign \new_[30785]_  = ~\new_[31322]_  & ~\new_[4074]_ ;
  assign \new_[30786]_  = ~\new_[31535]_  | ~\new_[31770]_ ;
  assign \new_[30787]_  = ~\new_[30860]_ ;
  assign \new_[30788]_  = \new_[31269]_  & \new_[4162]_ ;
  assign \new_[30789]_  = ~\new_[31509]_  | ~\new_[4177]_ ;
  assign \new_[30790]_  = ~\new_[31131]_ ;
  assign \new_[30791]_  = ~\new_[30991]_ ;
  assign \new_[30792]_  = s6_m5_cyc_r_reg;
  assign \new_[30793]_  = s8_m5_cyc_r_reg;
  assign \new_[30794]_  = s10_m5_cyc_r_reg;
  assign \new_[30795]_  = s5_m2_cyc_r_reg;
  assign \new_[30796]_  = ~\new_[6376]_  & ~\new_[6792]_ ;
  assign \new_[30797]_  = ~\new_[31113]_ ;
  assign \new_[30798]_  = ~\new_[30915]_ ;
  assign \new_[30799]_  = \new_[31262]_  | \new_[4047]_ ;
  assign \new_[30800]_  = ~\new_[5972]_  & ~\new_[31431]_ ;
  assign \new_[30801]_  = ~\new_[30906]_ ;
  assign \new_[30802]_  = ~\new_[31164]_ ;
  assign \new_[30803]_  = \new_[31410]_  | \new_[5987]_ ;
  assign \new_[30804]_  = ~\new_[30901]_ ;
  assign \new_[30805]_  = ~\new_[30900]_ ;
  assign \new_[30806]_  = ~\new_[30891]_ ;
  assign \new_[30807]_  = ~\new_[6037]_  | ~\new_[31506]_ ;
  assign \new_[30808]_  = ~\new_[30887]_ ;
  assign \new_[30809]_  = ~\new_[30883]_ ;
  assign \new_[30810]_  = \new_[6202]_  & \new_[31474]_ ;
  assign \new_[30811]_  = ~\new_[31020]_ ;
  assign \new_[30812]_  = ~\new_[31863]_  | ~\new_[6376]_ ;
  assign \new_[30813]_  = ~\new_[31863]_  | ~\new_[7917]_ ;
  assign \new_[30814]_  = \new_[31488]_  | \new_[4144]_ ;
  assign \new_[30815]_  = ~\new_[6268]_  & ~\new_[5995]_ ;
  assign \new_[30816]_  = ~\new_[30879]_ ;
  assign \new_[30817]_  = ~\new_[31863]_  | ~\new_[6794]_ ;
  assign \new_[30818]_  = ~\new_[30862]_ ;
  assign \new_[30819]_  = ~\new_[31229]_  | ~\new_[5993]_ ;
  assign \new_[30820]_  = \new_[31262]_  | \new_[31816]_ ;
  assign \new_[30821]_  = ~\new_[6056]_  | ~\new_[5900]_ ;
  assign \new_[30822]_  = ~\new_[6067]_  | ~\new_[5902]_ ;
  assign \new_[30823]_  = ~\m0_addr_i[30]  | ~\m0_addr_i[28] ;
  assign \new_[30824]_  = ~\new_[6095]_  & ~\new_[6217]_ ;
  assign \new_[30825]_  = \new_[6047]_  & \new_[5971]_ ;
  assign \new_[30826]_  = ~\new_[6052]_  & ~\new_[6053]_ ;
  assign \new_[30827]_  = ~\new_[31292]_  & ~\m0_addr_i[28] ;
  assign \new_[30828]_  = ~\new_[31388]_  | ~\new_[31602]_ ;
  assign \new_[30829]_  = ~\new_[6273]_  & ~\new_[6065]_ ;
  assign \new_[30830]_  = ~\new_[31863]_  | ~\new_[7915]_ ;
  assign \new_[30831]_  = ~\new_[6076]_  & ~\new_[5925]_ ;
  assign \new_[30832]_  = \new_[6189]_  & \new_[5990]_ ;
  assign \new_[30833]_  = ~\new_[6080]_  & ~\new_[5933]_ ;
  assign \new_[30834]_  = ~\new_[6193]_  & ~\new_[5903]_ ;
  assign \new_[30835]_  = ~\new_[31510]_  & ~\new_[4119]_ ;
  assign \new_[30836]_  = ~\new_[6052]_  | ~\new_[6053]_ ;
  assign \new_[30837]_  = ~\new_[31529]_  & ~\new_[4253]_ ;
  assign \new_[30838]_  = ~\new_[31229]_  & ~\new_[5993]_ ;
  assign \new_[30839]_  = ~\new_[30851]_ ;
  assign \new_[30840]_  = ~\new_[31277]_  & ~\new_[4445]_ ;
  assign \new_[30841]_  = ~\new_[4261]_  | ~n8304;
  assign \new_[30842]_  = ~\new_[31321]_  | ~\new_[4248]_ ;
  assign \new_[30843]_  = ~\new_[6200]_  | ~\new_[6048]_ ;
  assign \new_[30844]_  = ~\new_[31407]_  & ~\m5_addr_i[28] ;
  assign \new_[30845]_  = \new_[31501]_  & \new_[4215]_ ;
  assign \new_[30846]_  = ~\new_[31484]_  | ~\new_[31666]_ ;
  assign \new_[30847]_  = ~\new_[6083]_  & ~\new_[5906]_ ;
  assign \new_[30848]_  = ~\new_[30850]_ ;
  assign \new_[30849]_  = ~\new_[31226]_ ;
  assign \new_[30850]_  = ~\new_[6212]_ ;
  assign \new_[30851]_  = ~\new_[5994]_ ;
  assign \new_[30852]_  = ~\new_[31432]_ ;
  assign \new_[30853]_  = ~\new_[31673]_  | ~n8724;
  assign \new_[30854]_  = ~\new_[6003]_  & ~\new_[6088]_ ;
  assign \new_[30855]_  = ~\new_[31405]_ ;
  assign \new_[30856]_  = ~\new_[31512]_ ;
  assign \new_[30857]_  = ~\new_[31633]_  | ~n8794;
  assign \new_[30858]_  = ~\new_[31264]_ ;
  assign \new_[30859]_  = \new_[6375]_  & \new_[31582]_ ;
  assign \new_[30860]_  = \new_[6213]_  & \new_[5987]_ ;
  assign \new_[30861]_  = ~\new_[31333]_ ;
  assign \new_[30862]_  = \new_[31797]_  | \m5_addr_i[28] ;
  assign \new_[30863]_  = ~\new_[31277]_ ;
  assign \new_[30864]_  = \new_[6003]_  & \new_[6088]_ ;
  assign \new_[30865]_  = ~\new_[31662]_  | ~n8444;
  assign \new_[30866]_  = \new_[6077]_  & \new_[5993]_ ;
  assign \new_[30867]_  = \m2_addr_i[31]  | \new_[31699]_ ;
  assign \new_[30868]_  = ~\new_[4069]_  & ~\new_[31803]_ ;
  assign \new_[30869]_  = \m0_addr_i[29]  & \new_[31764]_ ;
  assign \new_[30870]_  = ~\new_[4115]_  & ~\new_[31559]_ ;
  assign \new_[30871]_  = ~\new_[31892]_  | ~\m5_addr_i[30] ;
  assign \new_[30872]_  = ~\new_[31719]_  & ~\new_[6065]_ ;
  assign \new_[30873]_  = ~\new_[4169]_  & ~\new_[31568]_ ;
  assign \new_[30874]_  = ~\new_[5919]_ ;
  assign \new_[30875]_  = ~\new_[31396]_ ;
  assign \new_[30876]_  = ~\new_[31700]_  | ~n8934;
  assign \new_[30877]_  = ~\new_[7222]_  & ~\new_[31573]_ ;
  assign \new_[30878]_  = ~\new_[31863]_  | ~\new_[6781]_ ;
  assign \new_[30879]_  = ~\m3_addr_i[31]  | ~\new_[31594]_ ;
  assign \new_[30880]_  = ~\new_[31863]_  | ~\new_[6793]_ ;
  assign \new_[30881]_  = ~\new_[31600]_  | ~n8629;
  assign \new_[30882]_  = \new_[31775]_  & \new_[6790]_ ;
  assign \new_[30883]_  = \new_[5898]_  | \new_[31705]_ ;
  assign \new_[30884]_  = ~\new_[31479]_ ;
  assign \new_[30885]_  = ~\new_[4261]_  & ~\new_[31589]_ ;
  assign \new_[30886]_  = ~\new_[31504]_ ;
  assign \new_[30887]_  = ~\new_[31849]_  | ~n8639;
  assign \new_[30888]_  = \new_[31555]_  & n8529;
  assign \new_[30889]_  = ~\new_[31642]_  | ~n8489;
  assign \new_[30890]_  = \new_[31695]_  & \new_[5982]_ ;
  assign \new_[30891]_  = ~\m2_addr_i[31]  | ~\new_[31699]_ ;
  assign \new_[30892]_  = ~\new_[31827]_  | ~n8549;
  assign \new_[30893]_  = ~\new_[5898]_  | ~\new_[31705]_ ;
  assign \new_[30894]_  = ~\new_[6069]_ ;
  assign \new_[30895]_  = \new_[3881]_  | \new_[31788]_ ;
  assign \new_[30896]_  = ~\new_[31586]_  | ~n8879;
  assign \new_[30897]_  = ~\new_[31411]_ ;
  assign \new_[30898]_  = ~\new_[31653]_  | ~n8789;
  assign \new_[30899]_  = \new_[31912]_  & n8849;
  assign \new_[30900]_  = ~\new_[31729]_  | ~n8884;
  assign \new_[30901]_  = ~\new_[31637]_  | ~n8434;
  assign \new_[30902]_  = ~\new_[31581]_  | ~n8769;
  assign \new_[30903]_  = ~\new_[31878]_  | ~n8844;
  assign \new_[30904]_  = ~\new_[31863]_  | ~\new_[6439]_ ;
  assign \new_[30905]_  = ~\new_[31936]_  | ~n8419;
  assign \new_[30906]_  = ~\new_[31929]_  | ~n8509;
  assign \new_[30907]_  = ~\new_[31840]_  | ~n8514;
  assign \new_[30908]_  = ~\new_[31817]_  & ~\new_[7439]_ ;
  assign \new_[30909]_  = ~\new_[31634]_  | ~\new_[5901]_ ;
  assign \new_[30910]_  = ~\new_[4233]_  & ~\new_[31722]_ ;
  assign \new_[30911]_  = ~\new_[4109]_  & ~\new_[31554]_ ;
  assign \new_[30912]_  = ~\new_[31624]_  | ~\new_[6192]_ ;
  assign \new_[30913]_  = ~\new_[31825]_  | ~n8609;
  assign \new_[30914]_  = \new_[31858]_  & n8449;
  assign \new_[30915]_  = ~\m0_addr_i[30]  | ~\new_[31485]_ ;
  assign \new_[30916]_  = ~\new_[31863]_  | ~\new_[6440]_ ;
  assign \new_[30917]_  = ~\new_[31863]_  | ~\new_[6789]_ ;
  assign \new_[30918]_  = ~m5_cyc_i | ~\new_[31638]_ ;
  assign \new_[30919]_  = ~\new_[31751]_  | ~\new_[5969]_ ;
  assign \new_[30920]_  = ~\new_[31847]_  | ~n8404;
  assign \new_[30921]_  = ~\new_[31919]_  | ~n8674;
  assign \new_[30922]_  = \m5_addr_i[31]  | \m5_addr_i[30] ;
  assign \new_[30923]_  = ~\new_[6073]_  | ~\new_[31895]_ ;
  assign \new_[30924]_  = ~\m2_addr_i[29]  & ~\new_[31668]_ ;
  assign \new_[30925]_  = ~\new_[5830]_ ;
  assign \new_[30926]_  = s8_m1_cyc_r_reg;
  assign \new_[30927]_  = ~\new_[31335]_ ;
  assign \new_[30928]_  = ~\new_[31863]_  | ~\new_[6790]_ ;
  assign \new_[30929]_  = ~\new_[4210]_  & ~\new_[31687]_ ;
  assign \new_[30930]_  = \new_[31817]_  & \new_[7439]_ ;
  assign \new_[30931]_  = ~\new_[31863]_  | ~\new_[6436]_ ;
  assign \new_[30932]_  = ~\new_[4176]_  & ~\new_[31598]_ ;
  assign \new_[30933]_  = ~\new_[31227]_ ;
  assign \new_[30934]_  = ~\m3_addr_i[31]  & ~\new_[31594]_ ;
  assign \new_[30935]_  = \new_[6784]_  & \new_[31742]_ ;
  assign \new_[30936]_  = ~\new_[6784]_  & ~\new_[31742]_ ;
  assign \new_[30937]_  = \new_[31766]_  & \new_[7918]_ ;
  assign \new_[30938]_  = ~\new_[31882]_  | ~n8919;
  assign \new_[30939]_  = ~\new_[31546]_ ;
  assign \new_[30940]_  = \new_[31730]_  & n8714;
  assign \new_[30941]_  = ~\new_[31842]_  | ~n8554;
  assign \new_[30942]_  = ~\new_[5972]_  & ~\new_[5973]_ ;
  assign \new_[30943]_  = ~\new_[31549]_ ;
  assign \new_[30944]_  = \new_[31560]_  & \new_[7436]_ ;
  assign \new_[30945]_  = ~\new_[31305]_ ;
  assign \new_[30946]_  = ~\new_[31829]_  | ~n8859;
  assign \new_[30947]_  = ~\new_[31327]_ ;
  assign \new_[30948]_  = \new_[31795]_  & \new_[6070]_ ;
  assign \new_[30949]_  = \new_[31751]_  | \new_[5969]_ ;
  assign \new_[30950]_  = \new_[31630]_  & n8399;
  assign \new_[30951]_  = ~\m4_addr_i[31]  | ~\new_[31922]_ ;
  assign \new_[30952]_  = ~\new_[31712]_ ;
  assign \new_[30953]_  = ~\new_[31719]_  | ~\new_[6065]_ ;
  assign \new_[30954]_  = ~\new_[31797]_  | ~\m5_addr_i[28] ;
  assign \new_[30955]_  = ~\new_[31721]_  | ~n8454;
  assign \new_[30956]_  = ~\new_[31595]_  & ~\new_[7916]_ ;
  assign \new_[30957]_  = ~\new_[31485]_ ;
  assign \new_[30958]_  = ~\new_[4150]_  & ~\new_[31864]_ ;
  assign \new_[30959]_  = ~\new_[31820]_  | ~n8429;
  assign \new_[30960]_  = ~\new_[4111]_  & ~\new_[31574]_ ;
  assign \new_[30961]_  = ~\new_[31663]_  | ~n8864;
  assign \new_[30962]_  = ~\new_[4102]_  & ~\new_[31655]_ ;
  assign \new_[30963]_  = ~\new_[31680]_  | ~n8914;
  assign \new_[30964]_  = ~\new_[31752]_  | ~n8754;
  assign \new_[30965]_  = ~\new_[31863]_  | ~\new_[7439]_ ;
  assign \new_[30966]_  = ~\m1_addr_i[31]  | ~\new_[31893]_ ;
  assign \new_[30967]_  = ~\new_[31625]_  | ~n8894;
  assign \new_[30968]_  = ~m2_cyc_i | ~\new_[31639]_ ;
  assign \new_[30969]_  = ~\new_[5985]_ ;
  assign \new_[30970]_  = \new_[31934]_  & \new_[6793]_ ;
  assign \new_[30971]_  = ~\new_[31606]_  | ~n8759;
  assign \new_[30972]_  = ~\new_[31908]_  | ~n8684;
  assign \new_[30973]_  = ~\new_[31934]_  & ~\new_[6793]_ ;
  assign \new_[30974]_  = ~\new_[6439]_  & ~\new_[31835]_ ;
  assign \new_[30975]_  = ~\new_[31833]_  | ~n8734;
  assign \new_[30976]_  = ~\new_[6033]_ ;
  assign \new_[30977]_  = ~\new_[31879]_  | ~n8649;
  assign \new_[30978]_  = ~\new_[31766]_  & ~\new_[7918]_ ;
  assign \new_[30979]_  = ~\new_[31654]_  | ~n8899;
  assign \new_[30980]_  = ~\new_[31734]_  | ~n8719;
  assign \new_[30981]_  = \new_[6091]_  | \new_[5908]_ ;
  assign \new_[30982]_  = ~\new_[31863]_  | ~\new_[6438]_ ;
  assign \new_[30983]_  = ~\new_[31808]_  | ~n8579;
  assign \new_[30984]_  = ~\new_[31514]_ ;
  assign \new_[30985]_  = ~\new_[31845]_  | ~\m1_addr_i[28] ;
  assign \new_[30986]_  = ~\new_[31775]_  & ~\new_[6790]_ ;
  assign \new_[30987]_  = ~\new_[31275]_ ;
  assign \new_[30988]_  = ~\new_[31933]_  & ~\new_[6792]_ ;
  assign \new_[30989]_  = ~\new_[6781]_  & ~\new_[31674]_ ;
  assign \new_[30990]_  = ~\new_[31355]_ ;
  assign \new_[30991]_  = \new_[6183]_  & \new_[6090]_ ;
  assign \new_[30992]_  = \new_[6205]_  | \new_[6046]_ ;
  assign \new_[30993]_  = ~\new_[6204]_ ;
  assign \new_[30994]_  = ~\new_[31225]_ ;
  assign \new_[30995]_  = ~\new_[31444]_ ;
  assign \new_[30996]_  = ~\new_[5988]_  & ~\new_[5920]_ ;
  assign \new_[30997]_  = ~\new_[31253]_ ;
  assign \new_[30998]_  = ~\new_[31442]_ ;
  assign \new_[30999]_  = ~\new_[31265]_ ;
  assign \new_[31000]_  = ~\new_[31342]_ ;
  assign \new_[31001]_  = ~\new_[31892]_ ;
  assign \new_[31002]_  = ~\new_[31536]_ ;
  assign \new_[31003]_  = ~\new_[31805]_  | ~n8654;
  assign \new_[31004]_  = ~\new_[31274]_ ;
  assign \new_[31005]_  = ~\new_[31322]_ ;
  assign \new_[31006]_  = ~\new_[31478]_ ;
  assign \new_[31007]_  = ~\new_[31460]_ ;
  assign \new_[31008]_  = \new_[6436]_  & \new_[31910]_ ;
  assign \new_[31009]_  = ~\new_[3876]_  & ~\new_[31661]_ ;
  assign \new_[31010]_  = ~\new_[31469]_ ;
  assign \new_[31011]_  = \new_[31695]_  | \new_[5982]_ ;
  assign \new_[31012]_  = ~\new_[4151]_ ;
  assign \new_[31013]_  = ~\new_[31284]_ ;
  assign \new_[31014]_  = ~\new_[5979]_ ;
  assign \new_[31015]_  = ~\new_[4446]_  & ~\new_[31599]_ ;
  assign \new_[31016]_  = ~\new_[31735]_  | ~n8589;
  assign \new_[31017]_  = ~\new_[31502]_ ;
  assign \new_[31018]_  = ~\new_[31684]_  | ~n8694;
  assign \new_[31019]_  = ~\new_[4217]_  & ~\new_[31636]_ ;
  assign \new_[31020]_  = ~\new_[31737]_  | ~n8744;
  assign \new_[31021]_  = ~\new_[31890]_  | ~\new_[5995]_ ;
  assign \new_[31022]_  = ~\new_[6436]_  & ~\new_[31910]_ ;
  assign \new_[31023]_  = ~\new_[4201]_  & ~\new_[31871]_ ;
  assign \new_[31024]_  = ~\new_[31621]_  | ~n8809;
  assign \new_[31025]_  = ~\new_[31795]_  & ~\new_[6070]_ ;
  assign \new_[31026]_  = ~\new_[4452]_  | ~n8384;
  assign \new_[31027]_  = ~\new_[31350]_ ;
  assign \new_[31028]_  = ~\new_[31863]_  | ~\new_[6784]_ ;
  assign \new_[31029]_  = ~\new_[31622]_  | ~n8409;
  assign \new_[31030]_  = \new_[31761]_  & n8479;
  assign \new_[31031]_  = ~\new_[4117]_  & ~\new_[31868]_ ;
  assign \new_[31032]_  = ~\new_[31917]_  | ~n8839;
  assign \new_[31033]_  = ~\new_[31345]_ ;
  assign \new_[31034]_  = ~\new_[31323]_ ;
  assign \new_[31035]_  = ~\new_[31767]_  | ~n8829;
  assign \new_[31036]_  = ~\new_[4439]_  & ~\new_[31651]_ ;
  assign \new_[31037]_  = ~\new_[31749]_  | ~n8679;
  assign \new_[31038]_  = ~\new_[31757]_  & ~\m3_addr_i[28] ;
  assign \new_[31039]_  = ~\new_[6031]_ ;
  assign \new_[31040]_  = ~\new_[31863]_  | ~\new_[6792]_ ;
  assign \new_[31041]_  = ~\new_[31859]_  | ~n8739;
  assign \new_[31042]_  = ~\new_[6064]_ ;
  assign \new_[31043]_  = ~\new_[6084]_ ;
  assign \new_[31044]_  = ~\new_[31902]_  | ~n8414;
  assign \new_[31045]_  = ~\new_[31403]_ ;
  assign \new_[31046]_  = ~\new_[31675]_  | ~n8459;
  assign \new_[31047]_  = ~m6_cyc_i | ~\new_[31783]_ ;
  assign \new_[31048]_  = \new_[31926]_  & n8749;
  assign \new_[31049]_  = ~\new_[6202]_  & ~\new_[5894]_ ;
  assign \new_[31050]_  = \new_[6781]_  & \new_[31674]_ ;
  assign \new_[31051]_  = ~\new_[3873]_  & ~\new_[31869]_ ;
  assign \new_[31052]_  = ~\new_[31603]_  | ~n8484;
  assign \new_[31053]_  = ~m3_cyc_i | ~\new_[31920]_ ;
  assign \new_[31054]_  = ~\new_[31420]_ ;
  assign \new_[31055]_  = \new_[31933]_  & \new_[6792]_ ;
  assign \new_[31056]_  = ~\new_[4266]_  & ~\new_[31579]_ ;
  assign \new_[31057]_  = ~\new_[31863]_  | ~\new_[7918]_ ;
  assign \new_[31058]_  = ~\new_[31821]_  | ~n8774;
  assign \new_[31059]_  = \m2_addr_i[29]  & \new_[31668]_ ;
  assign \new_[31060]_  = ~\new_[31732]_  | ~n8424;
  assign \new_[31061]_  = ~\m7_addr_i[31]  & ~\new_[31704]_ ;
  assign \new_[31062]_  = ~\new_[31796]_  | ~n8644;
  assign \new_[31063]_  = ~\new_[31860]_  | ~n8814;
  assign \new_[31064]_  = \new_[6174]_  & \new_[31593]_ ;
  assign \new_[31065]_  = ~\m6_addr_i[31]  & ~\new_[31861]_ ;
  assign \new_[31066]_  = ~\new_[4159]_  & ~\new_[31591]_ ;
  assign \new_[31067]_  = \new_[6199]_  & \new_[31887]_ ;
  assign \new_[31068]_  = ~\new_[31807]_  | ~n8729;
  assign \new_[31069]_  = ~\new_[31822]_  | ~n8929;
  assign \new_[31070]_  = ~\new_[31843]_  | ~n8584;
  assign \new_[31071]_  = ~\new_[31756]_  | ~n8504;
  assign \new_[31072]_  = \new_[6439]_  & \new_[31835]_ ;
  assign \new_[31073]_  = ~\new_[4134]_  & ~\new_[31930]_ ;
  assign \new_[31074]_  = ~\new_[4214]_  & ~\new_[31791]_ ;
  assign \new_[31075]_  = \new_[31595]_  & \new_[7916]_ ;
  assign \new_[31076]_  = ~\new_[31863]_  | ~\new_[7222]_ ;
  assign \new_[31077]_  = ~\new_[31694]_  | ~n8559;
  assign \new_[31078]_  = ~\new_[31831]_  | ~n8544;
  assign \new_[31079]_  = \new_[31786]_  & n8469;
  assign \new_[31080]_  = ~\new_[4273]_  & ~\new_[31561]_ ;
  assign \new_[31081]_  = \new_[6076]_  | \new_[31836]_ ;
  assign \new_[31082]_  = ~\m1_addr_i[31]  & ~\new_[31893]_ ;
  assign \new_[31083]_  = \new_[31701]_  & n8834;
  assign \new_[31084]_  = ~\new_[4203]_  & ~\new_[31577]_ ;
  assign \new_[31085]_  = \new_[6205]_  & \new_[6046]_ ;
  assign \new_[31086]_  = ~\new_[31611]_  | ~n8869;
  assign \new_[31087]_  = ~\new_[31798]_  | ~n8519;
  assign \new_[31088]_  = ~\new_[31297]_ ;
  assign \new_[31089]_  = \new_[6052]_  | \new_[31733]_ ;
  assign \new_[31090]_  = ~\new_[31670]_  | ~n8614;
  assign \new_[31091]_  = ~\new_[31863]_  | ~\new_[6780]_ ;
  assign \new_[31092]_  = ~\new_[31851]_  | ~n8564;
  assign \new_[31093]_  = ~\new_[31784]_  | ~n8464;
  assign \new_[31094]_  = \new_[6440]_  & \new_[31692]_ ;
  assign \new_[31095]_  = ~\new_[31664]_ ;
  assign \new_[31096]_  = ~\new_[5981]_ ;
  assign \new_[31097]_  = ~\new_[31881]_  | ~n8874;
  assign \new_[31098]_  = ~\new_[31445]_ ;
  assign \new_[31099]_  = ~\new_[4091]_  & ~\new_[31583]_ ;
  assign \new_[31100]_  = ~\new_[31865]_  & ~\new_[31941]_ ;
  assign \new_[31101]_  = ~\new_[31863]_  | ~\new_[7916]_ ;
  assign \new_[31102]_  = ~\new_[31778]_  | ~\new_[31941]_ ;
  assign \new_[31103]_  = ~\new_[4249]_  & ~\new_[31740]_ ;
  assign \new_[31104]_  = ~\new_[6269]_ ;
  assign \new_[31105]_  = ~\new_[31492]_ ;
  assign \new_[31106]_  = ~\new_[31493]_ ;
  assign \new_[31107]_  = ~\new_[31272]_ ;
  assign \new_[31108]_  = ~\new_[5996]_ ;
  assign \new_[31109]_  = ~\new_[31475]_ ;
  assign \new_[31110]_  = ~\new_[31489]_ ;
  assign \new_[31111]_  = ~\new_[31873]_  & ~\m6_addr_i[28] ;
  assign \new_[31112]_  = ~\new_[31341]_ ;
  assign \new_[31113]_  = ~\new_[31824]_  | ~n8689;
  assign \new_[31114]_  = ~\new_[31545]_ ;
  assign \new_[31115]_  = ~\new_[31890]_  & ~\new_[5995]_ ;
  assign \new_[31116]_  = ~\new_[4268]_  & ~\new_[31720]_ ;
  assign \new_[31117]_  = ~\new_[31863]_  | ~\new_[7436]_ ;
  assign \new_[31118]_  = ~\new_[6211]_  | ~\new_[31777]_ ;
  assign \new_[31119]_  = ~\new_[6440]_  & ~\new_[31692]_ ;
  assign \new_[31120]_  = ~\new_[3885]_  & ~\new_[31779]_ ;
  assign \new_[31121]_  = ~\new_[31471]_ ;
  assign \new_[31122]_  = ~\m7_addr_i[31]  | ~\new_[31704]_ ;
  assign \new_[31123]_  = ~\new_[31746]_  | ~n8384;
  assign \new_[31124]_  = ~\new_[31254]_ ;
  assign \new_[31125]_  = ~\new_[31676]_  | ~n8494;
  assign \new_[31126]_  = ~\new_[6076]_  | ~\new_[31836]_ ;
  assign \new_[31127]_  = ~\new_[31693]_  | ~n8904;
  assign \new_[31128]_  = ~\new_[5907]_ ;
  assign \new_[31129]_  = ~\new_[31780]_  | ~n8779;
  assign \new_[31130]_  = ~\new_[31863]_  | ~\new_[7435]_ ;
  assign \new_[31131]_  = ~\new_[31697]_  | ~n8659;
  assign \new_[31132]_  = ~\new_[31259]_ ;
  assign \new_[31133]_  = ~\new_[31510]_ ;
  assign \new_[31134]_  = \new_[31925]_  | \new_[5902]_ ;
  assign \new_[31135]_  = ~\new_[31490]_ ;
  assign \new_[31136]_  = ~\new_[6783]_  & ~\new_[31753]_ ;
  assign \new_[31137]_  = ~\new_[31785]_  | ~n8709;
  assign \new_[31138]_  = ~\m0_addr_i[29]  | ~\m0_addr_i[31] ;
  assign \new_[31139]_  = ~\new_[31927]_  | ~n8624;
  assign \new_[31140]_  = ~\new_[5999]_ ;
  assign \new_[31141]_  = \m7_addr_i[29]  | \new_[31894]_ ;
  assign \new_[31142]_  = ~\new_[31544]_ ;
  assign \new_[31143]_  = ~\new_[31551]_ ;
  assign \new_[31144]_  = ~\new_[31304]_ ;
  assign \new_[31145]_  = \new_[31757]_  & \m3_addr_i[28] ;
  assign \new_[31146]_  = ~\m7_addr_i[29]  | ~\new_[31894]_ ;
  assign \new_[31147]_  = ~\new_[31428]_ ;
  assign \new_[31148]_  = ~\new_[31539]_ ;
  assign \new_[31149]_  = ~\new_[31738]_  | ~n8394;
  assign \new_[31150]_  = \new_[31557]_  & n8474;
  assign \new_[31151]_  = ~\new_[31863]_  | ~\new_[6783]_ ;
  assign \new_[31152]_  = ~\m0_addr_i[29]  & ~\new_[31764]_ ;
  assign \new_[31153]_  = ~\new_[31875]_  | ~n8704;
  assign \new_[31154]_  = ~\new_[31762]_  | ~n8524;
  assign \new_[31155]_  = ~\m4_addr_i[29]  & ~\new_[31565]_ ;
  assign \new_[31156]_  = ~\new_[31905]_  & ~\new_[6215]_ ;
  assign \new_[31157]_  = ~\new_[31230]_ ;
  assign \new_[31158]_  = ~\new_[31560]_  & ~\new_[7436]_ ;
  assign \new_[31159]_  = ~\new_[5913]_ ;
  assign \new_[31160]_  = ~m0_cyc_i | ~\new_[31578]_ ;
  assign \new_[31161]_  = \new_[31634]_  | \new_[5901]_ ;
  assign \new_[31162]_  = ~m1_cyc_i | ~\new_[31818]_ ;
  assign \new_[31163]_  = \new_[6213]_  | \new_[5987]_ ;
  assign \new_[31164]_  = \new_[31845]_  | \m1_addr_i[28] ;
  assign \new_[31165]_  = ~\new_[6206]_ ;
  assign \new_[31166]_  = ~\new_[31924]_  | ~n8599;
  assign \new_[31167]_  = ~\new_[5988]_  | ~\new_[5920]_ ;
  assign \new_[31168]_  = ~\new_[31635]_  | ~n8604;
  assign \new_[31169]_  = ~\new_[31706]_  | ~n8764;
  assign \new_[31170]_  = ~\new_[31689]_  | ~n8804;
  assign \new_[31171]_  = ~\new_[31758]_  | ~n8889;
  assign \new_[31172]_  = \new_[31877]_  & n8534;
  assign \new_[31173]_  = ~\new_[31863]_  | ~\new_[7437]_ ;
  assign \new_[31174]_  = ~\new_[4053]_  & ~\new_[31631]_ ;
  assign \new_[31175]_  = ~\new_[6077]_  & ~\new_[5993]_ ;
  assign \new_[31176]_  = ~\new_[31441]_ ;
  assign \new_[31177]_  = ~\new_[31529]_ ;
  assign \new_[31178]_  = ~\new_[31321]_ ;
  assign \new_[31179]_  = ~\new_[31624]_  & ~\new_[6192]_ ;
  assign \new_[31180]_  = ~\new_[6071]_ ;
  assign \new_[31181]_  = ~\new_[4104]_  & ~\new_[31650]_ ;
  assign \new_[31182]_  = ~\new_[6052]_  | ~\new_[31733]_ ;
  assign \new_[31183]_  = ~\new_[31863]_  | ~\new_[6375]_ ;
  assign \new_[31184]_  = ~\new_[31677]_  | ~n8569;
  assign \new_[31185]_  = ~m7_cyc_i | ~\new_[31883]_ ;
  assign \new_[31186]_  = ~\new_[31872]_  | ~n8784;
  assign \new_[31187]_  = \new_[6783]_  & \new_[31753]_ ;
  assign \new_[31188]_  = ~\new_[31219]_ ;
  assign \new_[31189]_  = ~\m3_addr_i[29]  & ~\m3_addr_i[28] ;
  assign \new_[31190]_  = ~\new_[31353]_ ;
  assign \new_[31191]_  = ~\new_[31467]_ ;
  assign \new_[31192]_  = ~\new_[31273]_ ;
  assign \new_[31193]_  = ~\new_[31873]_  | ~\m6_addr_i[28] ;
  assign \new_[31194]_  = ~\new_[5972]_  | ~\new_[5973]_ ;
  assign \new_[31195]_  = ~\new_[6183]_  & ~\new_[6090]_ ;
  assign \new_[31196]_  = ~\new_[6091]_  | ~\new_[5908]_ ;
  assign \new_[31197]_  = ~\new_[31312]_ ;
  assign \new_[31198]_  = ~\new_[31426]_ ;
  assign \new_[31199]_  = ~m4_cyc_i | ~\new_[31715]_ ;
  assign \new_[31200]_  = ~\new_[31552]_ ;
  assign \new_[31201]_  = ~\new_[4250]_  & ~\new_[31584]_ ;
  assign \new_[31202]_  = ~\new_[6202]_  | ~\new_[5894]_ ;
  assign \new_[31203]_  = ~\new_[31300]_ ;
  assign \new_[31204]_  = ~\new_[31414]_ ;
  assign \new_[31205]_  = ~\new_[31572]_  | ~n8939;
  assign \new_[31206]_  = \m4_addr_i[29]  & \new_[31565]_ ;
  assign \new_[31207]_  = \new_[31892]_  | \m5_addr_i[30] ;
  assign \new_[31208]_  = \m6_addr_i[31]  & \new_[31861]_ ;
  assign \new_[31209]_  = ~\new_[31863]_  | ~\new_[6437]_ ;
  assign \new_[31210]_  = ~\new_[31398]_ ;
  assign \new_[31211]_  = ~\new_[6375]_  & ~\new_[31582]_ ;
  assign \new_[31212]_  = \new_[7222]_  & \new_[31573]_ ;
  assign \new_[31213]_  = ~\new_[31728]_  | ~n8909;
  assign \new_[31214]_  = \new_[4226]_  & n8564;
  assign \new_[31215]_  = ~\new_[4066]_  | ~n8899;
  assign \new_[31216]_  = ~\new_[6436]_  & ~\new_[6789]_ ;
  assign \new_[31217]_  = \new_[4127]_  & n8769;
  assign \new_[31218]_  = ~\new_[4268]_  | ~n8819;
  assign \new_[31219]_  = ~\new_[4120]_  | ~n8644;
  assign \new_[31220]_  = ~\new_[6438]_  & ~\new_[6793]_ ;
  assign \new_[31221]_  = \new_[6440]_  & \new_[6449]_ ;
  assign \new_[31222]_  = s4_m0_cyc_r_reg;
  assign \new_[31223]_  = s7_m1_cyc_r_reg;
  assign \new_[31224]_  = s5_m4_cyc_r_reg;
  assign \new_[31225]_  = \new_[4208]_  & n8519;
  assign \new_[31226]_  = ~\new_[4122]_  | ~n8674;
  assign \new_[31227]_  = ~\new_[6067]_  & ~\new_[5902]_ ;
  assign \new_[31228]_  = \new_[7224]_  & \new_[7916]_ ;
  assign \new_[31229]_  = ~\new_[6077]_ ;
  assign \new_[31230]_  = ~\new_[6066]_ ;
  assign \new_[31231]_  = s15_m2_cyc_r_reg;
  assign \new_[31232]_  = ~\new_[31815]_ ;
  assign \new_[31233]_  = s10_m3_cyc_r_reg;
  assign \new_[31234]_  = s0_m0_cyc_r_reg;
  assign \new_[31235]_  = ~\new_[31870]_ ;
  assign \new_[31236]_  = s5_m7_cyc_r_reg;
  assign \new_[31237]_  = s7_m7_cyc_r_reg;
  assign \new_[31238]_  = s11_m4_cyc_r_reg;
  assign \new_[31239]_  = s14_m5_cyc_r_reg;
  assign \new_[31240]_  = s15_m0_cyc_r_reg;
  assign \new_[31241]_  = s9_m7_cyc_r_reg;
  assign \new_[31242]_  = s0_m4_cyc_r_reg;
  assign \new_[31243]_  = s13_m4_cyc_r_reg;
  assign \new_[31244]_  = s2_m3_cyc_r_reg;
  assign \new_[31245]_  = ~\new_[4224]_  | ~n8529;
  assign \new_[31246]_  = s11_m1_cyc_r_reg;
  assign \new_[31247]_  = s13_m2_cyc_r_reg;
  assign \new_[31248]_  = s0_m2_cyc_r_reg;
  assign \new_[31249]_  = s9_m4_cyc_r_reg;
  assign \new_[31250]_  = \new_[4129]_  & n8459;
  assign \new_[31251]_  = s4_m7_cyc_r_reg;
  assign \new_[31252]_  = ~\new_[4273]_  | ~n8634;
  assign \new_[31253]_  = \m4_addr_i[31]  | \m4_addr_i[30] ;
  assign \new_[31254]_  = ~\new_[4166]_  | ~n8904;
  assign \new_[31255]_  = s13_m7_cyc_r_reg;
  assign \new_[31256]_  = \new_[4163]_  & n8399;
  assign \new_[31257]_  = ~\new_[4257]_  | ~n8834;
  assign \new_[31258]_  = s8_m0_cyc_r_reg;
  assign \new_[31259]_  = ~\new_[5930]_ ;
  assign \new_[31260]_  = ~\new_[4062]_  | ~n8629;
  assign \new_[31261]_  = s7_m2_cyc_r_reg;
  assign \new_[31262]_  = ~\new_[4046]_  | ~n8474;
  assign \new_[31263]_  = \new_[6783]_  & \new_[7915]_ ;
  assign \new_[31264]_  = ~\new_[4101]_  | ~n8709;
  assign \new_[31265]_  = \m0_addr_i[29]  | \m0_addr_i[31] ;
  assign \new_[31266]_  = \new_[4180]_  & n8914;
  assign \new_[31267]_  = ~\new_[4133]_  | ~n8729;
  assign \new_[31268]_  = ~\new_[4044]_  | ~n8589;
  assign \new_[31269]_  = \new_[4161]_  & n8774;
  assign \new_[31270]_  = \new_[4171]_  & n8424;
  assign \new_[31271]_  = \new_[3874]_  & n8809;
  assign \new_[31272]_  = ~\new_[4219]_  | ~n8604;
  assign \new_[31273]_  = ~\new_[4036]_  | ~n8414;
  assign \new_[31274]_  = \m6_addr_i[31]  | \m6_addr_i[30] ;
  assign \new_[31275]_  = ~\new_[4106]_  | ~n8689;
  assign \new_[31276]_  = ~\new_[31832]_ ;
  assign \new_[31277]_  = ~\new_[4438]_  | ~n8494;
  assign \new_[31278]_  = \new_[4039]_  & n8849;
  assign \new_[31279]_  = s7_m3_cyc_r_reg;
  assign \new_[31280]_  = \m2_addr_i[29]  | \m2_addr_i[28] ;
  assign \new_[31281]_  = \new_[4263]_  & n8879;
  assign \new_[31282]_  = s3_m1_cyc_r_reg;
  assign \new_[31283]_  = s9_m0_cyc_r_reg;
  assign \new_[31284]_  = ~\m3_addr_i[29]  | ~\m3_addr_i[28] ;
  assign \new_[31285]_  = s10_m1_cyc_r_reg;
  assign \new_[31286]_  = s6_m7_cyc_r_reg;
  assign \new_[31287]_  = s11_m2_cyc_r_reg;
  assign \new_[31288]_  = s13_m3_cyc_r_reg;
  assign \new_[31289]_  = s10_m2_cyc_r_reg;
  assign \new_[31290]_  = s12_m3_cyc_r_reg;
  assign \new_[31291]_  = s14_m6_cyc_r_reg;
  assign \new_[31292]_  = ~\new_[31691]_ ;
  assign \new_[31293]_  = ~\new_[4093]_  | ~n8624;
  assign \new_[31294]_  = s15_m7_cyc_r_reg;
  assign \new_[31295]_  = s10_m0_cyc_r_reg;
  assign \new_[31296]_  = s11_m3_cyc_r_reg;
  assign \new_[31297]_  = ~\new_[5898]_  & ~\new_[6051]_ ;
  assign \new_[31298]_  = s4_m2_cyc_r_reg;
  assign \new_[31299]_  = ~\new_[4251]_ ;
  assign \new_[31300]_  = ~\new_[4236]_  | ~n8584;
  assign \new_[31301]_  = ~\new_[4048]_  | ~n8864;
  assign \new_[31302]_  = ~\new_[4249]_  | ~n8669;
  assign \new_[31303]_  = \new_[6784]_  & \new_[7440]_ ;
  assign \new_[31304]_  = ~\new_[4265]_  | ~n8514;
  assign \new_[31305]_  = ~\new_[4441]_  | ~n8659;
  assign \new_[31306]_  = \new_[4243]_  & n8829;
  assign \new_[31307]_  = s7_m6_cyc_r_reg;
  assign \new_[31308]_  = ~\new_[31893]_ ;
  assign \new_[31309]_  = ~\new_[4080]_  | ~n8454;
  assign \new_[31310]_  = \new_[4448]_  & n8919;
  assign \new_[31311]_  = ~\new_[4147]_  | ~n8764;
  assign \new_[31312]_  = \m1_addr_i[31]  | \m1_addr_i[30] ;
  assign \new_[31313]_  = s9_m3_cyc_r_reg;
  assign \new_[31314]_  = s4_m6_cyc_r_reg;
  assign \new_[31315]_  = \new_[4200]_  & n8559;
  assign \new_[31316]_  = s0_m1_cyc_r_reg;
  assign \new_[31317]_  = ~\new_[6780]_  & ~\new_[7436]_ ;
  assign \new_[31318]_  = s1_m2_cyc_r_reg;
  assign \new_[31319]_  = \new_[4064]_  & n8544;
  assign \new_[31320]_  = \new_[4057]_  & n8909;
  assign \new_[31321]_  = \new_[4247]_  & n8884;
  assign \new_[31322]_  = ~\new_[4073]_  | ~n8489;
  assign \new_[31323]_  = ~\new_[4450]_  | ~n8859;
  assign \new_[31324]_  = \new_[3883]_  & n8404;
  assign \new_[31325]_  = s10_m7_cyc_r_reg;
  assign \new_[31326]_  = ~\new_[31778]_ ;
  assign \new_[31327]_  = ~\m1_addr_i[31]  | ~\m1_addr_i[30] ;
  assign \new_[31328]_  = \new_[7435]_  & \new_[7918]_ ;
  assign \new_[31329]_  = \new_[4091]_  & n8824;
  assign \new_[31330]_  = s11_m6_cyc_r_reg;
  assign \new_[31331]_  = ~\new_[4277]_  | ~n8579;
  assign \new_[31332]_  = ~\new_[4076]_  | ~n8469;
  assign \new_[31333]_  = ~\m3_addr_i[31]  & ~\m3_addr_i[30] ;
  assign \new_[31334]_  = s4_m4_cyc_r_reg;
  assign \new_[31335]_  = ~\new_[4082]_  | ~n8754;
  assign \new_[31336]_  = s9_m2_cyc_r_reg;
  assign \new_[31337]_  = \new_[6375]_  & \new_[6791]_ ;
  assign \new_[31338]_  = \new_[4266]_  & n8924;
  assign \new_[31339]_  = \new_[6439]_  & \new_[6794]_ ;
  assign \new_[31340]_  = ~\new_[31763]_ ;
  assign \new_[31341]_  = ~\new_[4115]_  | ~n8664;
  assign \new_[31342]_  = ~\m2_addr_i[29] ;
  assign \new_[31343]_  = s1_m5_cyc_r_reg;
  assign \new_[31344]_  = s14_m3_cyc_r_reg;
  assign \new_[31345]_  = ~\new_[5976]_ ;
  assign \new_[31346]_  = \new_[4159]_  & n8379;
  assign \new_[31347]_  = ~\new_[4233]_  | ~n8389;
  assign \new_[31348]_  = s12_m2_cyc_r_reg;
  assign \new_[31349]_  = s9_m1_cyc_r_reg;
  assign \new_[31350]_  = ~\new_[4136]_  | ~n8639;
  assign \new_[31351]_  = \new_[4138]_  & n8814;
  assign \new_[31352]_  = s3_m6_cyc_r_reg;
  assign \new_[31353]_  = ~\new_[4270]_  | ~n8444;
  assign \new_[31354]_  = s2_m6_cyc_r_reg;
  assign \new_[31355]_  = ~\m7_addr_i[31]  | ~\m7_addr_i[30] ;
  assign \new_[31356]_  = \new_[4245]_  & n8609;
  assign \new_[31357]_  = s6_m3_cyc_r_reg;
  assign \new_[31358]_  = ~\new_[4068]_  | ~n8794;
  assign \new_[31359]_  = s6_m6_cyc_r_reg;
  assign \new_[31360]_  = s8_m6_cyc_r_reg;
  assign \new_[31361]_  = s1_m4_cyc_r_reg;
  assign \new_[31362]_  = ~\new_[6183]_ ;
  assign \new_[31363]_  = s6_m0_cyc_r_reg;
  assign \new_[31364]_  = s2_m7_cyc_r_reg;
  assign \new_[31365]_  = s3_m3_cyc_r_reg;
  assign \new_[31366]_  = s12_m0_cyc_r_reg;
  assign \new_[31367]_  = s1_m7_cyc_r_reg;
  assign \new_[31368]_  = s8_m7_cyc_r_reg;
  assign \new_[31369]_  = s2_m0_cyc_r_reg;
  assign \new_[31370]_  = s1_m3_cyc_r_reg;
  assign \new_[31371]_  = s1_m0_cyc_r_reg;
  assign \new_[31372]_  = s3_m2_cyc_r_reg;
  assign \new_[31373]_  = s13_m6_cyc_r_reg;
  assign \new_[31374]_  = s2_m1_cyc_r_reg;
  assign \new_[31375]_  = \new_[4117]_  & n8699;
  assign \new_[31376]_  = s3_m0_cyc_r_reg;
  assign \new_[31377]_  = s2_m5_cyc_r_reg;
  assign \new_[31378]_  = \new_[4113]_  & n8704;
  assign \new_[31379]_  = s2_m4_cyc_r_reg;
  assign \new_[31380]_  = s5_m6_cyc_r_reg;
  assign \new_[31381]_  = s14_m4_cyc_r_reg;
  assign \new_[31382]_  = s14_m0_cyc_r_reg;
  assign \new_[31383]_  = ~\new_[5908]_ ;
  assign \new_[31384]_  = s15_m4_cyc_r_reg;
  assign \new_[31385]_  = s3_m4_cyc_r_reg;
  assign \new_[31386]_  = s2_m2_cyc_r_reg;
  assign \new_[31387]_  = s5_m3_cyc_r_reg;
  assign \new_[31388]_  = \new_[4212]_  & n8409;
  assign \new_[31389]_  = s12_m1_cyc_r_reg;
  assign \new_[31390]_  = ~\new_[31648]_ ;
  assign \new_[31391]_  = \new_[3876]_  & n8309;
  assign \new_[31392]_  = s5_m0_cyc_r_reg;
  assign \new_[31393]_  = \new_[6437]_  & \new_[6790]_ ;
  assign \new_[31394]_  = ~\new_[31615]_ ;
  assign \new_[31395]_  = s0_m7_cyc_r_reg;
  assign \new_[31396]_  = ~\new_[4125]_  | ~n8724;
  assign \new_[31397]_  = ~\new_[5967]_ ;
  assign \new_[31398]_  = \m2_addr_i[31]  | \m2_addr_i[30] ;
  assign \new_[31399]_  = ~\new_[31736]_ ;
  assign \new_[31400]_  = ~\new_[31795]_ ;
  assign \new_[31401]_  = ~\m2_addr_i[29]  | ~\m2_addr_i[28] ;
  assign \new_[31402]_  = \m3_addr_i[31]  & \m3_addr_i[30] ;
  assign \new_[31403]_  = ~\new_[6216]_ ;
  assign \new_[31404]_  = \new_[4078]_  & n8534;
  assign \new_[31405]_  = ~\new_[4083]_  | ~n8434;
  assign \new_[31406]_  = ~\new_[31772]_ ;
  assign \new_[31407]_  = ~\new_[31797]_ ;
  assign \new_[31408]_  = ~\new_[5988]_ ;
  assign \new_[31409]_  = ~\new_[4178]_  | ~n8504;
  assign \new_[31410]_  = ~\new_[6213]_ ;
  assign \new_[31411]_  = ~\new_[6210]_ ;
  assign \new_[31412]_  = ~\new_[4054]_ ;
  assign \new_[31413]_  = ~\new_[4218]_ ;
  assign \new_[31414]_  = ~\new_[4205]_  | ~n8599;
  assign \new_[31415]_  = \new_[4111]_  & n8594;
  assign \new_[31416]_  = ~\new_[6001]_ ;
  assign \new_[31417]_  = ~\new_[4135]_ ;
  assign \new_[31418]_  = ~\new_[4216]_  | ~n8929;
  assign \new_[31419]_  = ~\new_[5964]_ ;
  assign \new_[31420]_  = ~\new_[4254]_  | ~n8524;
  assign \new_[31421]_  = ~\new_[5997]_ ;
  assign \new_[31422]_  = ~\new_[31588]_ ;
  assign \new_[31423]_  = ~\new_[31690]_ ;
  assign \new_[31424]_  = ~\new_[4052]_  | ~n8684;
  assign \new_[31425]_  = ~\new_[4145]_  | ~n8679;
  assign \new_[31426]_  = ~\new_[4169]_  | ~n8574;
  assign \new_[31427]_  = \new_[4102]_  & n8619;
  assign \new_[31428]_  = ~\m5_addr_i[30] ;
  assign \new_[31429]_  = ~\new_[31906]_ ;
  assign \new_[31430]_  = \new_[4141]_  & n8509;
  assign \new_[31431]_  = ~\new_[5973]_ ;
  assign \new_[31432]_  = ~\new_[4443]_  | ~n8694;
  assign \new_[31433]_  = ~\new_[6096]_ ;
  assign \new_[31434]_  = \new_[7222]_  & \new_[7917]_ ;
  assign \new_[31435]_  = ~\new_[4050]_  | ~n8449;
  assign \new_[31436]_  = ~\new_[4037]_  | ~n8804;
  assign \new_[31437]_  = \new_[6438]_  & \new_[6793]_ ;
  assign \new_[31438]_  = ~\new_[31614]_ ;
  assign \new_[31439]_  = ~\new_[4228]_  | ~n8429;
  assign \new_[31440]_  = ~\new_[31685]_ ;
  assign \new_[31441]_  = ~\new_[6059]_ ;
  assign \new_[31442]_  = ~\new_[6184]_ ;
  assign \new_[31443]_  = \new_[4203]_  & n8854;
  assign \new_[31444]_  = ~\new_[3878]_  | ~n8554;
  assign \new_[31445]_  = ~\new_[4060]_  | ~n8779;
  assign \new_[31446]_  = ~\new_[4070]_ ;
  assign \new_[31447]_  = ~\new_[31773]_ ;
  assign \new_[31448]_  = s13_m0_cyc_r_reg;
  assign \new_[31449]_  = \new_[4149]_  & n8784;
  assign \new_[31450]_  = s1_m6_cyc_r_reg;
  assign \new_[31451]_  = ~\new_[7224]_  & ~\new_[7916]_ ;
  assign \new_[31452]_  = \new_[6781]_  & \new_[7437]_ ;
  assign \new_[31453]_  = s0_m5_cyc_r_reg;
  assign \new_[31454]_  = \new_[4446]_  & n8314;
  assign \new_[31455]_  = ~\new_[6072]_ ;
  assign \new_[31456]_  = s15_m5_cyc_r_reg;
  assign \new_[31457]_  = ~\new_[4279]_  | ~n8479;
  assign \new_[31458]_  = ~\new_[31640]_ ;
  assign \new_[31459]_  = s3_m7_cyc_r_reg;
  assign \new_[31460]_  = ~\new_[4154]_  | ~n8419;
  assign \new_[31461]_  = ~\new_[4174]_  | ~n8394;
  assign \new_[31462]_  = s9_m6_cyc_r_reg;
  assign \new_[31463]_  = s14_m2_cyc_r_reg;
  assign \new_[31464]_  = ~\new_[6176]_ ;
  assign \new_[31465]_  = ~\new_[4099]_  | ~n8889;
  assign \new_[31466]_  = s4_m3_cyc_r_reg;
  assign \new_[31467]_  = ~\m1_addr_i[29]  | ~\m1_addr_i[28] ;
  assign \new_[31468]_  = ~\new_[6781]_  & ~\new_[7437]_ ;
  assign \new_[31469]_  = ~\new_[4221]_  | ~n8934;
  assign \new_[31470]_  = \new_[3885]_  & n8354;
  assign \new_[31471]_  = ~\new_[5916]_ ;
  assign \new_[31472]_  = s6_m2_cyc_r_reg;
  assign \new_[31473]_  = \new_[6782]_  & \new_[7439]_ ;
  assign \new_[31474]_  = ~\new_[5894]_ ;
  assign \new_[31475]_  = ~\new_[4087]_  | ~n8894;
  assign \new_[31476]_  = \new_[4109]_  & n8334;
  assign \new_[31477]_  = ~\new_[31760]_ ;
  assign \new_[31478]_  = ~\new_[4095]_  | ~n8749;
  assign \new_[31479]_  = ~\new_[6196]_ ;
  assign \new_[31480]_  = \new_[4210]_  & n8539;
  assign \new_[31481]_  = \m0_addr_i[29] ;
  assign \new_[31482]_  = ~\new_[6190]_ ;
  assign \new_[31483]_  = ~\new_[4275]_  | ~n8614;
  assign \new_[31484]_  = \new_[4259]_  & n8649;
  assign \new_[31485]_  = ~\m0_addr_i[28] ;
  assign \new_[31486]_  = ~\new_[31699]_ ;
  assign \new_[31487]_  = \new_[6780]_  & \new_[7436]_ ;
  assign \new_[31488]_  = ~\new_[4143]_  | ~n8714;
  assign \new_[31489]_  = ~\new_[4104]_  | ~n8799;
  assign \new_[31490]_  = ~\m4_addr_i[29]  | ~\m4_addr_i[28] ;
  assign \new_[31491]_  = ~\new_[31652]_ ;
  assign \new_[31492]_  = \m7_addr_i[31]  | \m7_addr_i[30] ;
  assign \new_[31493]_  = ~\new_[4238]_  | ~n8484;
  assign \new_[31494]_  = ~\new_[5931]_ ;
  assign \new_[31495]_  = ~\new_[7435]_  & ~\new_[7918]_ ;
  assign \new_[31496]_  = ~\new_[31610]_ ;
  assign \new_[31497]_  = ~\new_[6437]_  & ~\new_[6790]_ ;
  assign \new_[31498]_  = ~\m5_addr_i[29]  | ~\m5_addr_i[28] ;
  assign \new_[31499]_  = ~\new_[31905]_ ;
  assign \new_[31500]_  = \new_[4097]_  & n8844;
  assign \new_[31501]_  = \new_[4214]_  & n8359;
  assign \new_[31502]_  = ~\m2_addr_i[31]  | ~\m2_addr_i[30] ;
  assign \new_[31503]_  = s7_m5_cyc_r_reg;
  assign \new_[31504]_  = ~\new_[4201]_  | ~n8374;
  assign \new_[31505]_  = \new_[3873]_  & n8439;
  assign \new_[31506]_  = ~\new_[5910]_ ;
  assign \new_[31507]_  = \new_[3887]_  & n8759;
  assign \new_[31508]_  = s13_m1_cyc_r_reg;
  assign \new_[31509]_  = \new_[4176]_  & n8499;
  assign \new_[31510]_  = ~\new_[4118]_  | ~n8734;
  assign \new_[31511]_  = s0_m6_cyc_r_reg;
  assign \new_[31512]_  = ~\new_[4055]_  | ~n8939;
  assign \new_[31513]_  = s10_m6_cyc_r_reg;
  assign \new_[31514]_  = ~\new_[4085]_  | ~n8549;
  assign \new_[31515]_  = s8_m4_cyc_r_reg;
  assign \new_[31516]_  = s0_m3_cyc_r_reg;
  assign \new_[31517]_  = s4_m5_cyc_r_reg;
  assign \new_[31518]_  = \new_[6376]_  & \new_[6792]_ ;
  assign \new_[31519]_  = s5_m1_cyc_r_reg;
  assign \new_[31520]_  = s6_m1_cyc_r_reg;
  assign \new_[31521]_  = ~\new_[6003]_ ;
  assign \new_[31522]_  = s4_m1_cyc_r_reg;
  assign \new_[31523]_  = s14_m1_cyc_r_reg;
  assign \new_[31524]_  = s14_m7_cyc_r_reg;
  assign \new_[31525]_  = s12_m4_cyc_r_reg;
  assign \new_[31526]_  = s7_m0_cyc_r_reg;
  assign \new_[31527]_  = s12_m7_cyc_r_reg;
  assign \new_[31528]_  = s7_m4_cyc_r_reg;
  assign \new_[31529]_  = ~\new_[4252]_  | ~n8654;
  assign \new_[31530]_  = s8_m3_cyc_r_reg;
  assign \new_[31531]_  = \m7_addr_i[29] ;
  assign \new_[31532]_  = s9_m5_cyc_r_reg;
  assign \new_[31533]_  = s11_m0_cyc_r_reg;
  assign \new_[31534]_  = s11_m7_cyc_r_reg;
  assign \new_[31535]_  = \new_[4167]_  & n8839;
  assign \new_[31536]_  = ~\new_[4152]_  | ~n8744;
  assign \new_[31537]_  = ~\new_[31623]_ ;
  assign \new_[31538]_  = ~\new_[31845]_ ;
  assign \new_[31539]_  = ~\new_[6032]_ ;
  assign \new_[31540]_  = \new_[4234]_  & n8869;
  assign \new_[31541]_  = \new_[4241]_  & n8569;
  assign \new_[31542]_  = s12_m6_cyc_r_reg;
  assign \new_[31543]_  = ~\new_[6782]_  & ~\new_[7439]_ ;
  assign \new_[31544]_  = ~\new_[4071]_  | ~n8719;
  assign \new_[31545]_  = ~\new_[4131]_  | ~n8739;
  assign \new_[31546]_  = ~\m6_addr_i[29]  | ~\m6_addr_i[28] ;
  assign \new_[31547]_  = ~\new_[31668]_ ;
  assign \new_[31548]_  = ~\new_[6270]_ ;
  assign \new_[31549]_  = ~\new_[4041]_  | ~n8789;
  assign \new_[31550]_  = \new_[6436]_  & \new_[6789]_ ;
  assign \new_[31551]_  = ~\new_[6205]_ ;
  assign \new_[31552]_  = ~\m5_addr_i[31]  | ~\m5_addr_i[30] ;
  assign \new_[31553]_  = ~\new_[6081]_ ;
  assign \new_[31554]_  = ~n8334;
  assign \new_[31555]_  = ~\new_[4224]_ ;
  assign \new_[31556]_  = ~\new_[4207]_ ;
  assign \new_[31557]_  = ~\new_[4046]_ ;
  assign \new_[31558]_  = ~\new_[4175]_ ;
  assign \new_[31559]_  = ~n8664;
  assign \new_[31560]_  = ~\new_[6780]_ ;
  assign \new_[31561]_  = ~n8634;
  assign \new_[31562]_  = ~\new_[5984]_ ;
  assign \new_[31563]_  = ~\m5_addr_i[26] ;
  assign \new_[31564]_  = ~\new_[6785]_ ;
  assign \new_[31565]_  = ~\m4_addr_i[28] ;
  assign \new_[31566]_  = ~\new_[4092]_ ;
  assign \new_[31567]_  = ~\new_[5905]_ ;
  assign \new_[31568]_  = ~n8574;
  assign \new_[31569]_  = ~\new_[5897]_ ;
  assign \new_[31570]_  = ~\new_[4116]_ ;
  assign \new_[31571]_  = ~\new_[4246]_ ;
  assign \new_[31572]_  = ~\new_[4055]_ ;
  assign \new_[31573]_  = ~\new_[7917]_ ;
  assign \new_[31574]_  = ~n8594;
  assign \new_[31575]_  = ~\new_[6445]_ ;
  assign \new_[31576]_  = ~\new_[7919]_ ;
  assign \new_[31577]_  = ~n8854;
  assign \new_[31578]_  = ~m0_stb_i;
  assign \new_[31579]_  = ~n8924;
  assign \new_[31580]_  = ~\new_[4223]_ ;
  assign \new_[31581]_  = ~\new_[4127]_ ;
  assign \new_[31582]_  = ~\new_[6791]_ ;
  assign \new_[31583]_  = ~n8824;
  assign \new_[31584]_  = ~n8364;
  assign \new_[31585]_  = ~\m7_addr_i[2] ;
  assign \new_[31586]_  = ~\new_[4263]_ ;
  assign \new_[31587]_  = ~\new_[4124]_ ;
  assign \new_[31588]_  = ~\new_[5975]_ ;
  assign \new_[31589]_  = ~n8304;
  assign \new_[31590]_  = ~\new_[4227]_ ;
  assign \new_[31591]_  = ~n8379;
  assign \new_[31592]_  = ~\m2_addr_i[2] ;
  assign \new_[31593]_  = ~\new_[6034]_ ;
  assign \new_[31594]_  = ~\m3_addr_i[30] ;
  assign \new_[31595]_  = ~\new_[7224]_ ;
  assign \new_[31596]_  = ~\new_[6057]_ ;
  assign \new_[31597]_  = ~\new_[7221]_ ;
  assign \new_[31598]_  = ~n8499;
  assign \new_[31599]_  = ~n8314;
  assign \new_[31600]_  = ~\new_[4062]_ ;
  assign \new_[31601]_  = ~\new_[4179]_ ;
  assign \new_[31602]_  = ~\new_[4213]_ ;
  assign \new_[31603]_  = ~\new_[4238]_ ;
  assign \new_[31604]_  = ~\new_[4160]_ ;
  assign \new_[31605]_  = ~\new_[4181]_ ;
  assign \new_[31606]_  = ~\new_[3887]_ ;
  assign \new_[31607]_  = ~\new_[4119]_ ;
  assign \new_[31608]_  = ~\new_[6058]_ ;
  assign \new_[31609]_  = ~\m2_addr_i[26] ;
  assign \new_[31610]_  = ~\m7_addr_i[31] ;
  assign \new_[31611]_  = ~\new_[4234]_ ;
  assign \new_[31612]_  = ~\m6_addr_i[25] ;
  assign \new_[31613]_  = ~\new_[3886]_ ;
  assign \new_[31614]_  = ~\new_[6208]_ ;
  assign \new_[31615]_  = ~\new_[5915]_ ;
  assign \new_[31616]_  = ~\new_[6039]_ ;
  assign \new_[31617]_  = ~\new_[6041]_ ;
  assign \new_[31618]_  = ~\new_[4098]_ ;
  assign \new_[31619]_  = ~\m3_addr_i[24] ;
  assign \new_[31620]_  = ~\new_[4051]_ ;
  assign \new_[31621]_  = ~\new_[3874]_ ;
  assign \new_[31622]_  = ~\new_[4212]_ ;
  assign \new_[31623]_  = ~\m2_addr_i[31] ;
  assign \new_[31624]_  = ~\new_[6214]_ ;
  assign \new_[31625]_  = ~\new_[4087]_ ;
  assign \new_[31626]_  = ~\m5_addr_i[24] ;
  assign \new_[31627]_  = ~\new_[4280]_ ;
  assign \new_[31628]_  = ~\new_[4445]_ ;
  assign \new_[31629]_  = ~\new_[4142]_ ;
  assign \new_[31630]_  = ~\new_[4163]_ ;
  assign \new_[31631]_  = ~n8344;
  assign \new_[31632]_  = ~\new_[4067]_ ;
  assign \new_[31633]_  = ~\new_[4068]_ ;
  assign \new_[31634]_  = ~\new_[6062]_ ;
  assign \new_[31635]_  = ~\new_[4219]_ ;
  assign \new_[31636]_  = ~n8339;
  assign \new_[31637]_  = ~\new_[4083]_ ;
  assign \new_[31638]_  = ~m5_stb_i;
  assign \new_[31639]_  = ~m2_stb_i;
  assign \new_[31640]_  = ~\m1_addr_i[28] ;
  assign \new_[31641]_  = ~\new_[4162]_ ;
  assign \new_[31642]_  = ~\new_[4073]_ ;
  assign \new_[31643]_  = ~\new_[6068]_ ;
  assign \new_[31644]_  = ~\m6_addr_i[26] ;
  assign \new_[31645]_  = ~\new_[6246]_ ;
  assign \new_[31646]_  = ~\new_[4059]_ ;
  assign \new_[31647]_  = ~\m0_addr_i[4] ;
  assign \new_[31648]_  = \new_[6002]_ ;
  assign \new_[31649]_  = ~\new_[4256]_ ;
  assign \new_[31650]_  = ~n8799;
  assign \new_[31651]_  = ~n8369;
  assign \new_[31652]_  = ~\new_[6055]_ ;
  assign \new_[31653]_  = ~\new_[4041]_ ;
  assign \new_[31654]_  = ~\new_[4066]_ ;
  assign \new_[31655]_  = ~n8619;
  assign \new_[31656]_  = ~\new_[4264]_ ;
  assign \new_[31657]_  = ~\new_[4094]_ ;
  assign \new_[31658]_  = ~\new_[4222]_ ;
  assign \new_[31659]_  = ~\new_[4140]_ ;
  assign \new_[31660]_  = ~\new_[6047]_ ;
  assign \new_[31661]_  = ~n8309;
  assign \new_[31662]_  = ~\new_[4270]_ ;
  assign \new_[31663]_  = ~\new_[4048]_ ;
  assign \new_[31664]_  = ~\m2_addr_i[5] ;
  assign \new_[31665]_  = ~\new_[6038]_ ;
  assign \new_[31666]_  = ~\new_[4260]_ ;
  assign \new_[31667]_  = ~\m7_addr_i[24] ;
  assign \new_[31668]_  = ~\m2_addr_i[28] ;
  assign \new_[31669]_  = ~\new_[6035]_ ;
  assign \new_[31670]_  = ~\new_[4275]_ ;
  assign \new_[31671]_  = ~\m5_addr_i[4] ;
  assign \new_[31672]_  = ~\new_[4112]_ ;
  assign \new_[31673]_  = ~\new_[4125]_ ;
  assign \new_[31674]_  = ~\new_[7437]_ ;
  assign \new_[31675]_  = ~\new_[4129]_ ;
  assign \new_[31676]_  = ~\new_[4438]_ ;
  assign \new_[31677]_  = ~\new_[4241]_ ;
  assign \new_[31678]_  = ~\new_[6446]_ ;
  assign \new_[31679]_  = ~\new_[4079]_ ;
  assign \new_[31680]_  = ~\new_[4180]_ ;
  assign \new_[31681]_  = ~\new_[4177]_ ;
  assign \new_[31682]_  = ~\new_[4453]_ ;
  assign \new_[31683]_  = ~\new_[6006]_ ;
  assign \new_[31684]_  = ~\new_[4443]_ ;
  assign \new_[31685]_  = ~\new_[6054]_ ;
  assign \new_[31686]_  = ~\new_[5903]_ ;
  assign \new_[31687]_  = ~n8539;
  assign \new_[31688]_  = ~\m2_addr_i[25] ;
  assign \new_[31689]_  = ~\new_[4037]_ ;
  assign \new_[31690]_  = ~\new_[6271]_ ;
  assign \new_[31691]_  = ~\m0_addr_i[30] ;
  assign \new_[31692]_  = ~\new_[6449]_ ;
  assign \new_[31693]_  = ~\new_[4166]_ ;
  assign \new_[31694]_  = ~\new_[4200]_ ;
  assign \new_[31695]_  = ~\new_[6063]_ ;
  assign \new_[31696]_  = ~\new_[4139]_ ;
  assign \new_[31697]_  = ~\new_[4441]_ ;
  assign \new_[31698]_  = ~\new_[6788]_ ;
  assign \new_[31699]_  = ~\m2_addr_i[30] ;
  assign \new_[31700]_  = ~\new_[4221]_ ;
  assign \new_[31701]_  = ~\new_[4257]_ ;
  assign \new_[31702]_  = ~\new_[4038]_ ;
  assign \new_[31703]_  = ~\m2_addr_i[4] ;
  assign \new_[31704]_  = ~\m7_addr_i[30] ;
  assign \new_[31705]_  = ~\new_[6051]_ ;
  assign \new_[31706]_  = ~\new_[4147]_ ;
  assign \new_[31707]_  = ~\new_[5904]_ ;
  assign \new_[31708]_  = ~\new_[4144]_ ;
  assign \new_[31709]_  = ~\new_[3884]_ ;
  assign \new_[31710]_  = ~\new_[4211]_ ;
  assign \new_[31711]_  = ~\new_[4170]_ ;
  assign \new_[31712]_  = \new_[6207]_ ;
  assign \new_[31713]_  = ~\new_[4242]_ ;
  assign \new_[31714]_  = ~\new_[4156]_ ;
  assign \new_[31715]_  = ~m4_stb_i;
  assign \new_[31716]_  = ~\new_[4088]_ ;
  assign \new_[31717]_  = ~\new_[4225]_ ;
  assign \new_[31718]_  = ~\new_[6444]_ ;
  assign \new_[31719]_  = ~\new_[6273]_ ;
  assign \new_[31720]_  = ~n8819;
  assign \new_[31721]_  = ~\new_[4080]_ ;
  assign \new_[31722]_  = ~n8389;
  assign \new_[31723]_  = ~\new_[4042]_ ;
  assign \new_[31724]_  = ~\new_[5932]_ ;
  assign \new_[31725]_  = ~\new_[6195]_ ;
  assign \new_[31726]_  = \m7_addr_i[3] ;
  assign \new_[31727]_  = ~\new_[4172]_ ;
  assign \new_[31728]_  = ~\new_[4057]_ ;
  assign \new_[31729]_  = ~\new_[4247]_ ;
  assign \new_[31730]_  = ~\new_[4143]_ ;
  assign \new_[31731]_  = ~\new_[4090]_ ;
  assign \new_[31732]_  = ~\new_[4171]_ ;
  assign \new_[31733]_  = ~\new_[6053]_ ;
  assign \new_[31734]_  = ~\new_[4071]_ ;
  assign \new_[31735]_  = ~\new_[4044]_ ;
  assign \new_[31736]_  = ~\m2_addr_i[3] ;
  assign \new_[31737]_  = ~\new_[4152]_ ;
  assign \new_[31738]_  = ~\new_[4174]_ ;
  assign \new_[31739]_  = ~\m1_addr_i[26] ;
  assign \new_[31740]_  = ~n8669;
  assign \new_[31741]_  = ~\new_[6050]_ ;
  assign \new_[31742]_  = ~\new_[7440]_ ;
  assign \new_[31743]_  = ~\new_[3888]_ ;
  assign \new_[31744]_  = ~\new_[4103]_ ;
  assign \new_[31745]_  = ~\m6_addr_i[27] ;
  assign \new_[31746]_  = ~\new_[4452]_ ;
  assign \new_[31747]_  = ~\m5_addr_i[2] ;
  assign \new_[31748]_  = ~\new_[4258]_ ;
  assign \new_[31749]_  = ~\new_[4145]_ ;
  assign \new_[31750]_  = ~\m2_addr_i[27] ;
  assign \new_[31751]_  = ~\new_[6044]_ ;
  assign \new_[31752]_  = ~\new_[4082]_ ;
  assign \new_[31753]_  = ~\new_[7915]_ ;
  assign \new_[31754]_  = ~\new_[4262]_ ;
  assign \new_[31755]_  = ~\new_[4269]_ ;
  assign \new_[31756]_  = ~\new_[4178]_ ;
  assign \new_[31757]_  = ~\m3_addr_i[29] ;
  assign \new_[31758]_  = ~\new_[4099]_ ;
  assign \new_[31759]_  = ~\new_[6786]_ ;
  assign \new_[31760]_  = ~\m1_addr_i[2] ;
  assign \new_[31761]_  = ~\new_[4279]_ ;
  assign \new_[31762]_  = ~\new_[4254]_ ;
  assign \new_[31763]_  = \new_[6004]_ ;
  assign \new_[31764]_  = ~\m0_addr_i[31] ;
  assign \new_[31765]_  = ~\new_[5933]_ ;
  assign \new_[31766]_  = ~\new_[7435]_ ;
  assign \new_[31767]_  = ~\new_[4243]_ ;
  assign \new_[31768]_  = ~\new_[4045]_ ;
  assign \new_[31769]_  = ~\new_[4040]_ ;
  assign \new_[31770]_  = ~\new_[4168]_ ;
  assign \new_[31771]_  = ~\new_[4148]_ ;
  assign \new_[31772]_  = ~\new_[6209]_ ;
  assign \new_[31773]_  = ~\m1_addr_i[31] ;
  assign \new_[31774]_  = ~\new_[4158]_ ;
  assign \new_[31775]_  = ~\new_[6437]_ ;
  assign \new_[31776]_  = ~\new_[6092]_ ;
  assign \new_[31777]_  = ~\new_[6061]_ ;
  assign \new_[31778]_  = ~\new_[6779]_ ;
  assign \new_[31779]_  = ~n8354;
  assign \new_[31780]_  = ~\new_[4060]_ ;
  assign \new_[31781]_  = ~\new_[4455]_ ;
  assign \new_[31782]_  = ~\m7_addr_i[4] ;
  assign \new_[31783]_  = ~m6_stb_i;
  assign \new_[31784]_  = ~\new_[4230]_ ;
  assign \new_[31785]_  = ~\new_[4101]_ ;
  assign \new_[31786]_  = ~\new_[4076]_ ;
  assign \new_[31787]_  = ~\new_[5991]_ ;
  assign \new_[31788]_  = ~n8349;
  assign \new_[31789]_  = ~\new_[6086]_ ;
  assign \new_[31790]_  = ~\m1_addr_i[25] ;
  assign \new_[31791]_  = ~n8359;
  assign \new_[31792]_  = ~\new_[4077]_ ;
  assign \new_[31793]_  = ~\m5_addr_i[25] ;
  assign \new_[31794]_  = ~\m5_addr_i[27] ;
  assign \new_[31795]_  = ~\new_[6191]_ ;
  assign \new_[31796]_  = ~\new_[4120]_ ;
  assign \new_[31797]_  = ~\m5_addr_i[29] ;
  assign \new_[31798]_  = ~\new_[4208]_ ;
  assign \new_[31799]_  = ~\new_[6095]_ ;
  assign \new_[31800]_  = ~\new_[5895]_ ;
  assign \new_[31801]_  = ~\new_[4276]_ ;
  assign \new_[31802]_  = ~\new_[4081]_ ;
  assign \new_[31803]_  = ~n8324;
  assign \new_[31804]_  = ~\new_[6448]_ ;
  assign \new_[31805]_  = ~\new_[4252]_ ;
  assign \new_[31806]_  = ~\new_[4267]_ ;
  assign \new_[31807]_  = ~\new_[4133]_ ;
  assign \new_[31808]_  = ~\new_[4277]_ ;
  assign \new_[31809]_  = ~\new_[4231]_ ;
  assign \new_[31810]_  = ~\new_[6442]_ ;
  assign \new_[31811]_  = ~\new_[4274]_ ;
  assign \new_[31812]_  = ~\m0_addr_i[2] ;
  assign \new_[31813]_  = ~\new_[4173]_ ;
  assign \new_[31814]_  = ~\new_[4108]_ ;
  assign \new_[31815]_  = ~\new_[5974]_ ;
  assign \new_[31816]_  = ~\new_[4047]_ ;
  assign \new_[31817]_  = ~\new_[6782]_ ;
  assign \new_[31818]_  = ~m1_stb_i;
  assign \new_[31819]_  = ~\new_[5992]_ ;
  assign \new_[31820]_  = ~\new_[4228]_ ;
  assign \new_[31821]_  = ~\new_[4161]_ ;
  assign \new_[31822]_  = ~\new_[4216]_ ;
  assign \new_[31823]_  = ~\new_[4075]_ ;
  assign \new_[31824]_  = ~\new_[4106]_ ;
  assign \new_[31825]_  = ~\new_[4245]_ ;
  assign \new_[31826]_  = ~\new_[4105]_ ;
  assign \new_[31827]_  = ~\new_[4085]_ ;
  assign \new_[31828]_  = ~\new_[4202]_ ;
  assign \new_[31829]_  = ~\new_[4450]_ ;
  assign \new_[31830]_  = ~\new_[6787]_ ;
  assign \new_[31831]_  = ~\new_[4064]_ ;
  assign \new_[31832]_  = ~\m5_addr_i[28] ;
  assign \new_[31833]_  = ~\new_[4118]_ ;
  assign \new_[31834]_  = ~\new_[3875]_ ;
  assign \new_[31835]_  = ~\new_[6794]_ ;
  assign \new_[31836]_  = ~\new_[5925]_ ;
  assign \new_[31837]_  = ~\new_[6189]_ ;
  assign \new_[31838]_  = ~\new_[4058]_ ;
  assign \new_[31839]_  = ~\new_[5906]_ ;
  assign \new_[31840]_  = ~\new_[4265]_ ;
  assign \new_[31841]_  = ~\new_[4114]_ ;
  assign \new_[31842]_  = ~\new_[3878]_ ;
  assign \new_[31843]_  = ~\new_[4236]_ ;
  assign \new_[31844]_  = ~\new_[5968]_ ;
  assign \new_[31845]_  = ~\m1_addr_i[29] ;
  assign \new_[31846]_  = ~\new_[6441]_ ;
  assign \new_[31847]_  = ~\new_[3883]_ ;
  assign \new_[31848]_  = \m0_addr_i[5] ;
  assign \new_[31849]_  = ~\new_[4136]_ ;
  assign \new_[31850]_  = ~\new_[4215]_ ;
  assign \new_[31851]_  = ~\new_[4226]_ ;
  assign \new_[31852]_  = ~\new_[4065]_ ;
  assign \new_[31853]_  = ~\new_[7920]_ ;
  assign \new_[31854]_  = ~\new_[4244]_ ;
  assign \new_[31855]_  = ~\new_[6007]_ ;
  assign \new_[31856]_  = ~\new_[4449]_ ;
  assign \new_[31857]_  = ~\new_[6274]_ ;
  assign \new_[31858]_  = ~\new_[4050]_ ;
  assign \new_[31859]_  = ~\new_[4131]_ ;
  assign \new_[31860]_  = ~\new_[4138]_ ;
  assign \new_[31861]_  = ~\m6_addr_i[30] ;
  assign \new_[31862]_  = ~\new_[6185]_ ;
  assign \new_[31863]_  = ~rst_i;
  assign \new_[31864]_  = ~n8319;
  assign \new_[31865]_  = ~\new_[6779]_ ;
  assign \new_[31866]_  = ~\new_[5900]_ ;
  assign \new_[31867]_  = ~\new_[3880]_ ;
  assign \new_[31868]_  = ~n8699;
  assign \new_[31869]_  = ~n8439;
  assign \new_[31870]_  = ~\new_[5977]_ ;
  assign \new_[31871]_  = ~n8374;
  assign \new_[31872]_  = ~\new_[4149]_ ;
  assign \new_[31873]_  = ~\m6_addr_i[29] ;
  assign \new_[31874]_  = ~\m6_addr_i[3] ;
  assign \new_[31875]_  = ~\new_[4113]_ ;
  assign \new_[31876]_  = ~\new_[4110]_ ;
  assign \new_[31877]_  = ~\new_[4078]_ ;
  assign \new_[31878]_  = ~\new_[4097]_ ;
  assign \new_[31879]_  = ~\new_[4259]_ ;
  assign \new_[31880]_  = ~\new_[4204]_ ;
  assign \new_[31881]_  = ~\new_[4157]_ ;
  assign \new_[31882]_  = ~\new_[4448]_ ;
  assign \new_[31883]_  = ~m7_stb_i;
  assign \new_[31884]_  = \m0_addr_i[3] ;
  assign \new_[31885]_  = \m7_addr_i[30] ;
  assign \new_[31886]_  = ~\new_[4049]_ ;
  assign \new_[31887]_  = ~\new_[5970]_ ;
  assign \new_[31888]_  = ~\new_[6443]_ ;
  assign \new_[31889]_  = ~\new_[4130]_ ;
  assign \new_[31890]_  = ~\new_[6268]_ ;
  assign \new_[31891]_  = ~\new_[4063]_ ;
  assign \new_[31892]_  = ~\m5_addr_i[31] ;
  assign \new_[31893]_  = ~\m1_addr_i[30] ;
  assign \new_[31894]_  = ~\m7_addr_i[28] ;
  assign \new_[31895]_  = ~\new_[5989]_ ;
  assign \new_[31896]_  = ~\new_[3882]_ ;
  assign \new_[31897]_  = ~\new_[3877]_ ;
  assign \new_[31898]_  = ~\new_[4239]_ ;
  assign \new_[31899]_  = ~\new_[4128]_ ;
  assign \new_[31900]_  = ~\new_[6082]_ ;
  assign \new_[31901]_  = ~\new_[5928]_ ;
  assign \new_[31902]_  = ~\new_[4036]_ ;
  assign \new_[31903]_  = ~\new_[5896]_ ;
  assign \new_[31904]_  = ~\new_[4146]_ ;
  assign \new_[31905]_  = ~\new_[6089]_ ;
  assign \new_[31906]_  = ~\new_[5899]_ ;
  assign \new_[31907]_  = ~\m1_addr_i[24] ;
  assign \new_[31908]_  = ~\new_[4052]_ ;
  assign \new_[31909]_  = ~\new_[4278]_ ;
  assign \new_[31910]_  = ~\new_[6789]_ ;
  assign \new_[31911]_  = ~\new_[4164]_ ;
  assign \new_[31912]_  = ~\new_[4039]_ ;
  assign \new_[31913]_  = ~\m1_addr_i[27] ;
  assign \new_[31914]_  = ~\new_[4440]_ ;
  assign \new_[31915]_  = ~\new_[6203]_ ;
  assign \new_[31916]_  = ~\new_[4240]_ ;
  assign \new_[31917]_  = ~\new_[4167]_ ;
  assign \new_[31918]_  = ~\new_[4229]_ ;
  assign \new_[31919]_  = ~\new_[4122]_ ;
  assign \new_[31920]_  = ~m3_stb_i;
  assign \new_[31921]_  = ~\new_[4447]_ ;
  assign \new_[31922]_  = ~\m4_addr_i[30] ;
  assign \new_[31923]_  = ~\new_[5916]_ ;
  assign \new_[31924]_  = ~\new_[4205]_ ;
  assign \new_[31925]_  = ~\new_[6067]_ ;
  assign \new_[31926]_  = ~\new_[4095]_ ;
  assign \new_[31927]_  = ~\new_[4093]_ ;
  assign \new_[31928]_  = ~\new_[6200]_ ;
  assign \new_[31929]_  = ~\new_[4141]_ ;
  assign \new_[31930]_  = ~n8329;
  assign \new_[31931]_  = ~\new_[4454]_ ;
  assign \new_[31932]_  = ~\new_[4235]_ ;
  assign \new_[31933]_  = ~\new_[6376]_ ;
  assign \new_[31934]_  = ~\new_[6438]_ ;
  assign \new_[31935]_  = ~\new_[6447]_ ;
  assign \new_[31936]_  = ~\new_[4154]_ ;
  assign \new_[31937]_  = ~\new_[4096]_ ;
  assign \new_[31938]_  = ~\new_[31941]_ ;
  assign \new_[31939]_  = ~\new_[31940]_ ;
  assign \new_[31940]_  = \new_[31941]_ ;
  assign \new_[31941]_  = ~\new_[7434]_ ;
  assign n7424 = ~\new_[7218]_ ;
  assign \new_[31943]_  = ~\new_[31948]_  | ~\new_[5089]_  | ~\new_[31944]_ ;
  assign \new_[31944]_  = \new_[31945]_  & \new_[31946]_ ;
  assign \new_[31945]_  = \new_[14717]_  & \new_[14714]_ ;
  assign \new_[31946]_  = ~\new_[31947]_ ;
  assign \new_[31947]_  = ~\new_[16118]_  | ~\new_[16119]_  | ~\new_[14713]_ ;
  assign \new_[31948]_  = \new_[31949]_  & \new_[31953]_ ;
  assign \new_[31949]_  = ~\new_[31950]_ ;
  assign \new_[31950]_  = ~\new_[31952]_  | ~\new_[16951]_  | ~\new_[31951]_ ;
  assign \new_[31951]_  = ~s14_err_i | ~\new_[17272]_  | ~\new_[29641]_ ;
  assign \new_[31952]_  = ~s12_err_i | ~\new_[19615]_  | ~\new_[29317]_ ;
  assign \new_[31953]_  = ~\new_[31954]_ ;
  assign \new_[31954]_  = ~\new_[14715]_  | ~\new_[17813]_  | ~\new_[16954]_ ;
  assign \new_[31955]_  = ~\new_[31959]_  | ~\new_[5090]_  | ~\new_[31956]_ ;
  assign \new_[31956]_  = ~\new_[31957]_  & ~\new_[31958]_ ;
  assign \new_[31957]_  = ~\new_[16957]_  | ~\new_[16122]_  | ~\new_[13324]_ ;
  assign \new_[31958]_  = ~\new_[14725]_  | ~\new_[14721]_ ;
  assign \new_[31959]_  = \new_[31960]_  & \new_[31962]_ ;
  assign \new_[31960]_  = ~\new_[31961]_ ;
  assign \new_[31961]_  = ~\new_[14722]_  | ~\new_[17814]_  | ~\new_[14719]_ ;
  assign \new_[31962]_  = ~\new_[31963]_ ;
  assign \new_[31963]_  = ~\new_[31965]_  | ~\new_[16121]_  | ~\new_[31964]_ ;
  assign \new_[31964]_  = ~s14_rty_i | ~\new_[17272]_  | ~\new_[29641]_ ;
  assign \new_[31965]_  = ~s12_rty_i | ~\new_[19615]_  | ~\new_[29317]_ ;
  assign \new_[31966]_  = ~\new_[31973]_  | ~\new_[5091]_  | ~\new_[31967]_ ;
  assign \new_[31967]_  = \new_[31968]_  & \new_[31972]_ ;
  assign \new_[31968]_  = ~\new_[31970]_  & (~\new_[18015]_  | ~\new_[31969]_ );
  assign \new_[31969]_  = \new_[30311]_  & s11_err_i;
  assign \new_[31970]_  = ~\new_[16140]_  | ~\new_[31971]_ ;
  assign \new_[31971]_  = ~s8_err_i | ~\new_[18760]_  | ~\new_[29636]_ ;
  assign \new_[31972]_  = \new_[14754]_  & \new_[17020]_ ;
  assign \new_[31973]_  = \new_[31974]_  & \new_[31976]_ ;
  assign \new_[31974]_  = ~\new_[31975]_ ;
  assign \new_[31975]_  = ~\new_[13357]_  | ~\new_[18654]_  | ~\new_[17021]_ ;
  assign \new_[31976]_  = ~\new_[31977]_ ;
  assign \new_[31977]_  = ~\new_[18655]_  | ~\new_[17019]_  | ~\new_[17022]_ ;
  assign \new_[31978]_  = ~\new_[31984]_  | ~\new_[31983]_  | ~\new_[31979]_  | ~\new_[31982]_ ;
  assign \new_[31979]_  = ~\new_[32260]_  | ~\new_[31980]_  | ~\new_[31981]_ ;
  assign \new_[31980]_  = \new_[32278]_  & s15_rty_i;
  assign \new_[31981]_  = \new_[17367]_  & \new_[19372]_ ;
  assign \new_[31982]_  = ~s13_rty_i | ~\new_[17194]_  | ~\new_[32267]_ ;
  assign \new_[31983]_  = ~s6_rty_i | ~\new_[18742]_  | ~\new_[29704]_ ;
  assign \new_[31984]_  = ~s7_rty_i | ~\new_[20542]_  | ~\new_[30060]_ ;
  assign \new_[31985]_  = \new_[31980]_ ;
  assign \new_[31986]_  = ~\new_[31994]_  | ~\new_[31993]_  | ~\new_[31987]_  | ~\new_[31992]_ ;
  assign \new_[31987]_  = ~\new_[32343]_  | ~\new_[31988]_  | ~\new_[31989]_ ;
  assign \new_[31988]_  = \new_[32278]_  & s15_err_i;
  assign \new_[31989]_  = \new_[14830]_ ;
  assign \new_[31990]_  = \new_[31991]_ ;
  assign \new_[31991]_  = ~\new_[22413]_  | ~\new_[20813]_  | ~\new_[22102]_ ;
  assign \new_[31992]_  = ~s13_err_i | ~\new_[18114]_  | ~\new_[32338]_ ;
  assign \new_[31993]_  = ~s0_err_i | ~\new_[18826]_  | ~\new_[27879]_ ;
  assign \new_[31994]_  = ~s4_err_i | ~\new_[19584]_  | ~\new_[27855]_ ;
  assign \new_[31995]_  = ~\new_[31989]_ ;
  assign \new_[31996]_  = ~\new_[31991]_ ;
  assign \new_[31997]_  = \new_[31988]_ ;
  assign \new_[31998]_  = (~\s13_data_i[28]  | ~\new_[32327]_ ) & (~\new_[31999]_  | ~\new_[32321]_ );
  assign \new_[31999]_  = \new_[32278]_  & \s15_data_i[28] ;
  assign \new_[32000]_  = ~\new_[32001]_  | ~\new_[32301]_ ;
  assign \new_[32001]_  = ~\new_[32002]_  & ~\new_[32003]_ ;
  assign \new_[32002]_  = ~\new_[31860]_  & ~\new_[5891]_ ;
  assign \new_[32003]_  = ~\new_[5735]_  | ~\new_[5734]_ ;
  assign \new_[32004]_  = \new_[32005]_  & \new_[32007]_ ;
  assign \new_[32005]_  = ~\new_[32006]_  | ~\new_[32161]_ ;
  assign \new_[32006]_  = \new_[3819]_  ? \new_[32011]_  : \s15_data_i[15] ;
  assign \new_[32007]_  = ~\new_[32168]_  | ~\s13_data_i[15] ;
  assign \new_[32008]_  = \new_[32009]_  & \new_[32012]_ ;
  assign \new_[32009]_  = ~\new_[32010]_  | ~\new_[32127]_ ;
  assign \new_[32010]_  = \new_[3820]_  ? \new_[32011]_  : \s15_data_i[13] ;
  assign \new_[32011]_  = ~\new_[32315]_ ;
  assign \new_[32012]_  = ~\new_[32134]_  | ~\s13_data_i[13] ;
  assign \m2_data_o[9]  = ~\new_[3675]_  | ~\new_[32014]_ ;
  assign \new_[32014]_  = \new_[32015]_  & \new_[32016]_ ;
  assign \new_[32015]_  = \new_[27415]_  & \new_[25513]_ ;
  assign \new_[32016]_  = ~\new_[32017]_  & ~\new_[32022]_ ;
  assign \new_[32017]_  = ~\new_[32021]_  | ~\new_[32020]_  | ~\new_[32018]_  | ~\new_[32019]_ ;
  assign \new_[32018]_  = ~\new_[28714]_  | ~\s5_data_i[9] ;
  assign \new_[32019]_  = ~\new_[29807]_  | ~\s14_data_i[9] ;
  assign \new_[32020]_  = (~\s8_data_i[9]  | ~\new_[30341]_ ) & (~\new_[30709]_  | ~\s3_data_i[9] );
  assign \new_[32021]_  = (~\s11_data_i[9]  | ~\new_[29876]_ ) & (~\new_[30626]_  | ~\s12_data_i[9] );
  assign \new_[32022]_  = ~\new_[25525]_  | ~\new_[32023]_ ;
  assign \new_[32023]_  = (~\s1_data_i[9]  | ~\new_[30357]_ ) & (~\new_[29788]_  | ~\s2_data_i[9] );
  assign \m2_data_o[7]  = ~\new_[3739]_  | ~\new_[32025]_ ;
  assign \new_[32025]_  = \new_[32026]_  & \new_[32027]_ ;
  assign \new_[32026]_  = \new_[27368]_  & \new_[25335]_ ;
  assign \new_[32027]_  = ~\new_[32028]_  & ~\new_[32033]_ ;
  assign \new_[32028]_  = ~\new_[32032]_  | ~\new_[32031]_  | ~\new_[32029]_  | ~\new_[32030]_ ;
  assign \new_[32029]_  = ~\new_[28714]_  | ~\s5_data_i[7] ;
  assign \new_[32030]_  = ~\new_[29807]_  | ~\s14_data_i[7] ;
  assign \new_[32031]_  = (~\s8_data_i[7]  | ~\new_[30341]_ ) & (~\new_[30709]_  | ~\s3_data_i[7] );
  assign \new_[32032]_  = (~\s11_data_i[7]  | ~\new_[29876]_ ) & (~\new_[30626]_  | ~\s12_data_i[7] );
  assign \new_[32033]_  = ~\new_[25032]_  | ~\new_[32034]_ ;
  assign \new_[32034]_  = (~\s1_data_i[7]  | ~\new_[30357]_ ) & (~\new_[29788]_  | ~\s2_data_i[7] );
  assign \m2_data_o[4]  = ~\new_[3684]_  | ~\new_[32036]_ ;
  assign \new_[32036]_  = \new_[32037]_  & \new_[32038]_ ;
  assign \new_[32037]_  = \new_[27160]_  & \new_[25915]_ ;
  assign \new_[32038]_  = ~\new_[32039]_  & ~\new_[32044]_ ;
  assign \new_[32039]_  = ~\new_[32043]_  | ~\new_[32042]_  | ~\new_[32040]_  | ~\new_[32041]_ ;
  assign \new_[32040]_  = ~\new_[28714]_  | ~\s5_data_i[4] ;
  assign \new_[32041]_  = ~\new_[29807]_  | ~\s14_data_i[4] ;
  assign \new_[32042]_  = (~\s8_data_i[4]  | ~\new_[30341]_ ) & (~\new_[30709]_  | ~\s3_data_i[4] );
  assign \new_[32043]_  = (~\s11_data_i[4]  | ~\new_[29876]_ ) & (~\new_[30626]_  | ~\s12_data_i[4] );
  assign \new_[32044]_  = ~\new_[25501]_  | ~\new_[32045]_ ;
  assign \new_[32045]_  = (~\s1_data_i[4]  | ~\new_[30357]_ ) & (~\new_[29788]_  | ~\s2_data_i[4] );
  assign \new_[32046]_  = ~\new_[32055]_  | ~\new_[32047]_  | ~\new_[32050]_ ;
  assign \new_[32047]_  = ~\new_[32048]_  | ~\new_[32049]_ ;
  assign \new_[32048]_  = \new_[3812]_  ? \new_[32011]_  : \s15_data_i[1] ;
  assign \new_[32049]_  = ~\new_[31401]_  & ~\new_[31502]_ ;
  assign \new_[32050]_  = ~\new_[32051]_ ;
  assign \new_[32051]_  = ~\new_[32054]_  | ~\new_[32052]_  | ~\new_[32053]_ ;
  assign \new_[32052]_  = (~\s9_data_i[1]  | ~\new_[29709]_ ) & (~\new_[29021]_  | ~\s10_data_i[1] );
  assign \new_[32053]_  = (~\s6_data_i[1]  | ~\new_[29298]_ ) & (~\new_[30193]_  | ~\s7_data_i[1] );
  assign \new_[32054]_  = (~\s0_data_i[1]  | ~\new_[30481]_ ) & (~\new_[29963]_  | ~\s4_data_i[1] );
  assign \new_[32055]_  = ~\new_[32056]_  | ~\s13_data_i[1] ;
  assign \new_[32056]_  = \new_[30924]_  & \new_[31017]_ ;
  assign \new_[32057]_  = ~\new_[32049]_ ;
  assign \new_[32058]_  = ~\new_[5728]_  | ~\new_[5727]_ ;
  assign \new_[32059]_  = ~\new_[31417]_  & ~\new_[5891]_ ;
  assign \new_[32060]_  = ~\new_[32061]_  | ~\new_[32062]_ ;
  assign \new_[32061]_  = ~\new_[5943]_  | ~\new_[4084]_ ;
  assign \new_[32062]_  = ~\new_[32068]_  | ~\new_[4151]_ ;
  assign \new_[32063]_  = ~\new_[5943]_  | ~\new_[4093]_ ;
  assign \new_[32064]_  = ~\new_[32068]_  | ~\new_[4161]_ ;
  assign \new_[32065]_  = \new_[32066]_  & \new_[32067]_ ;
  assign \new_[32066]_  = ~\new_[4143]_  | ~\new_[32171]_ ;
  assign \new_[32067]_  = ~\new_[32068]_  | ~\new_[4159]_ ;
  assign \new_[32068]_  = ~\new_[32069]_ ;
  assign \new_[32069]_  = ~\new_[32070]_ ;
  assign \new_[32070]_  = \new_[6373]_  & \new_[6374]_ ;
  assign \m2_data_o[0]  = ~\new_[3746]_  | ~\new_[32072]_ ;
  assign \new_[32072]_  = \new_[32073]_  & \new_[32074]_ ;
  assign \new_[32073]_  = \new_[27218]_  & \new_[24703]_ ;
  assign \new_[32074]_  = ~\new_[32075]_  & ~\new_[32080]_ ;
  assign \new_[32075]_  = ~\new_[32079]_  | ~\new_[32078]_  | ~\new_[32076]_  | ~\new_[32077]_ ;
  assign \new_[32076]_  = ~\new_[28714]_  | ~\s5_data_i[0] ;
  assign \new_[32077]_  = ~\new_[29807]_  | ~\s14_data_i[0] ;
  assign \new_[32078]_  = (~\s8_data_i[0]  | ~\new_[30341]_ ) & (~\new_[30709]_  | ~\s3_data_i[0] );
  assign \new_[32079]_  = (~\s11_data_i[0]  | ~\new_[29876]_ ) & (~\new_[30626]_  | ~\s12_data_i[0] );
  assign \new_[32080]_  = ~\new_[25449]_  | ~\new_[32081]_ ;
  assign \new_[32081]_  = (~\s1_data_i[0]  | ~\new_[30357]_ ) & (~\new_[29788]_  | ~\s2_data_i[0] );
  assign \new_[32082]_  = ~\new_[32090]_  | ~\new_[32083]_  | ~\new_[32085]_ ;
  assign \new_[32083]_  = ~\new_[32084]_  | ~\new_[32161]_ ;
  assign \new_[32084]_  = \new_[3804]_  ? \new_[32011]_  : \s15_data_i[14] ;
  assign \new_[32085]_  = ~\new_[32086]_ ;
  assign \new_[32086]_  = ~\new_[32089]_  | ~\new_[32087]_  | ~\new_[32088]_ ;
  assign \new_[32087]_  = (~\s0_data_i[14]  | ~\new_[29819]_ ) & (~\new_[29961]_  | ~\s4_data_i[14] );
  assign \new_[32088]_  = (~\s9_data_i[14]  | ~\new_[29024]_ ) & (~\new_[29710]_  | ~\s10_data_i[14] );
  assign \new_[32089]_  = (~\s6_data_i[14]  | ~\new_[29939]_ ) & (~\new_[30131]_  | ~\s7_data_i[14] );
  assign \new_[32090]_  = ~\new_[32168]_  | ~\s13_data_i[14] ;
  assign \m6_data_o[9]  = ~\new_[3679]_  | ~\new_[32092]_ ;
  assign \new_[32092]_  = \new_[32093]_  & \new_[32094]_ ;
  assign \new_[32093]_  = \new_[26497]_  & \new_[27194]_ ;
  assign \new_[32094]_  = ~\new_[32095]_  & ~\new_[32100]_ ;
  assign \new_[32095]_  = ~\new_[32099]_  | ~\new_[32098]_  | ~\new_[32096]_  | ~\new_[32097]_ ;
  assign \new_[32096]_  = (~\s12_data_i[9]  | ~\new_[29621]_ ) & (~\new_[29631]_  | ~\s14_data_i[9] );
  assign \new_[32097]_  = (~\s8_data_i[9]  | ~\new_[29420]_ ) & (~\new_[30429]_  | ~\s3_data_i[9] );
  assign \new_[32098]_  = ~\new_[30284]_  | ~\s11_data_i[9] ;
  assign \new_[32099]_  = ~\new_[29036]_  | ~\s5_data_i[9] ;
  assign \new_[32100]_  = ~\new_[25866]_  | ~\new_[32101]_ ;
  assign \new_[32101]_  = (~\s1_data_i[9]  | ~\new_[30108]_ ) & (~\new_[30085]_  | ~\s2_data_i[9] );
  assign \m6_data_o[7]  = ~\new_[3742]_  | ~\new_[32103]_ ;
  assign \new_[32103]_  = \new_[32104]_  & \new_[32105]_ ;
  assign \new_[32104]_  = \new_[25336]_  & \new_[27145]_ ;
  assign \new_[32105]_  = ~\new_[32106]_  & ~\new_[32111]_ ;
  assign \new_[32106]_  = ~\new_[32110]_  | ~\new_[32109]_  | ~\new_[32107]_  | ~\new_[32108]_ ;
  assign \new_[32107]_  = (~\s12_data_i[7]  | ~\new_[29621]_ ) & (~\new_[29631]_  | ~\s14_data_i[7] );
  assign \new_[32108]_  = (~\s8_data_i[7]  | ~\new_[29420]_ ) & (~\new_[30429]_  | ~\s3_data_i[7] );
  assign \new_[32109]_  = ~\new_[30284]_  | ~\s11_data_i[7] ;
  assign \new_[32110]_  = ~\new_[29036]_  | ~\s5_data_i[7] ;
  assign \new_[32111]_  = ~\new_[25478]_  | ~\new_[32112]_ ;
  assign \new_[32112]_  = (~\s1_data_i[7]  | ~\new_[30108]_ ) & (~\new_[30085]_  | ~\s2_data_i[7] );
  assign \m6_data_o[4]  = ~\new_[3685]_  | ~\new_[32114]_ ;
  assign \new_[32114]_  = \new_[32115]_  & \new_[32116]_ ;
  assign \new_[32115]_  = \new_[25497]_  & \new_[27161]_ ;
  assign \new_[32116]_  = ~\new_[32117]_  & ~\new_[32122]_ ;
  assign \new_[32117]_  = ~\new_[32121]_  | ~\new_[32120]_  | ~\new_[32118]_  | ~\new_[32119]_ ;
  assign \new_[32118]_  = (~\s12_data_i[4]  | ~\new_[29621]_ ) & (~\new_[29631]_  | ~\s14_data_i[4] );
  assign \new_[32119]_  = (~\s8_data_i[4]  | ~\new_[29420]_ ) & (~\new_[30429]_  | ~\s3_data_i[4] );
  assign \new_[32120]_  = ~\new_[30284]_  | ~\s11_data_i[4] ;
  assign \new_[32121]_  = ~\new_[29036]_  | ~\s5_data_i[4] ;
  assign \new_[32122]_  = ~\new_[25405]_  | ~\new_[32123]_ ;
  assign \new_[32123]_  = (~\s1_data_i[4]  | ~\new_[30108]_ ) & (~\new_[30085]_  | ~\s2_data_i[4] );
  assign \new_[32124]_  = ~\new_[32133]_  | ~\new_[32125]_  | ~\new_[32128]_ ;
  assign \new_[32125]_  = ~\new_[32126]_  | ~\new_[32127]_ ;
  assign \new_[32126]_  = \new_[3825]_  ? \new_[5883]_  : \s15_data_i[0] ;
  assign \new_[32127]_  = \new_[30939]_  & \new_[30592]_ ;
  assign \new_[32128]_  = ~\new_[32129]_ ;
  assign \new_[32129]_  = ~\new_[32132]_  | ~\new_[32130]_  | ~\new_[32131]_ ;
  assign \new_[32130]_  = (~\s0_data_i[0]  | ~\new_[29651]_ ) & (~\new_[29149]_  | ~\s4_data_i[0] );
  assign \new_[32131]_  = (~\s6_data_i[0]  | ~\new_[29954]_ ) & (~\new_[29823]_  | ~\s7_data_i[0] );
  assign \new_[32132]_  = (~\s9_data_i[0]  | ~\new_[29706]_ ) & (~\new_[30227]_  | ~\s10_data_i[0] );
  assign \new_[32133]_  = ~\new_[32134]_  | ~\s13_data_i[0] ;
  assign \new_[32134]_  = \new_[30744]_  & \new_[30592]_ ;
  assign \new_[32135]_  = ~\new_[32127]_ ;
  assign \m3_data_o[9]  = ~\new_[3703]_  | ~\new_[32137]_ ;
  assign \new_[32137]_  = \new_[32138]_  & \new_[32145]_ ;
  assign \new_[32138]_  = ~\new_[32139]_  & ~\new_[32144]_ ;
  assign \new_[32139]_  = ~\new_[32143]_  | ~\new_[32142]_  | ~\new_[32140]_  | ~\new_[32141]_ ;
  assign \new_[32140]_  = (~\s8_data_i[9]  | ~\new_[29428]_ ) & (~\new_[29948]_  | ~\s5_data_i[9] );
  assign \new_[32141]_  = (~\s11_data_i[9]  | ~\new_[30200]_ ) & (~\new_[30166]_  | ~\s14_data_i[9] );
  assign \new_[32142]_  = ~\new_[29947]_  | ~\s3_data_i[9] ;
  assign \new_[32143]_  = ~\new_[30298]_  | ~\s12_data_i[9] ;
  assign \new_[32144]_  = ~\new_[27467]_  | ~\new_[27569]_ ;
  assign \new_[32145]_  = \new_[25717]_  & \new_[32146]_ ;
  assign \new_[32146]_  = (~\s1_data_i[9]  | ~\new_[30001]_ ) & (~\new_[29846]_  | ~\s2_data_i[9] );
  assign \m3_data_o[7]  = ~\new_[3758]_  | ~\new_[32148]_ ;
  assign \new_[32148]_  = \new_[32149]_  & \new_[32156]_ ;
  assign \new_[32149]_  = ~\new_[32150]_  & ~\new_[32155]_ ;
  assign \new_[32150]_  = ~\new_[32154]_  | ~\new_[32153]_  | ~\new_[32151]_  | ~\new_[32152]_ ;
  assign \new_[32151]_  = (~\s8_data_i[7]  | ~\new_[29428]_ ) & (~\new_[29948]_  | ~\s5_data_i[7] );
  assign \new_[32152]_  = (~\s11_data_i[7]  | ~\new_[30200]_ ) & (~\new_[30166]_  | ~\s14_data_i[7] );
  assign \new_[32153]_  = ~\new_[29947]_  | ~\s3_data_i[7] ;
  assign \new_[32154]_  = ~\new_[30298]_  | ~\s12_data_i[7] ;
  assign \new_[32155]_  = ~\new_[27141]_  | ~\new_[27057]_ ;
  assign \new_[32156]_  = \new_[25891]_  & \new_[32157]_ ;
  assign \new_[32157]_  = (~\s1_data_i[7]  | ~\new_[30001]_ ) & (~\new_[29846]_  | ~\s2_data_i[7] );
  assign \new_[32158]_  = ~\new_[32167]_  | ~\new_[32159]_  | ~\new_[32162]_ ;
  assign \new_[32159]_  = ~\new_[32160]_  | ~\new_[32161]_ ;
  assign \new_[32160]_  = \new_[3810]_  ? \new_[5883]_  : \s15_data_i[4] ;
  assign \new_[32161]_  = \new_[31013]_  & \new_[31402]_ ;
  assign \new_[32162]_  = ~\new_[32163]_ ;
  assign \new_[32163]_  = ~\new_[32166]_  | ~\new_[32164]_  | ~\new_[32165]_ ;
  assign \new_[32164]_  = (~\s0_data_i[4]  | ~\new_[29819]_ ) & (~\new_[29961]_  | ~\s4_data_i[4] );
  assign \new_[32165]_  = (~\s9_data_i[4]  | ~\new_[29024]_ ) & (~\new_[29710]_  | ~\s10_data_i[4] );
  assign \new_[32166]_  = (~\s6_data_i[4]  | ~\new_[29939]_ ) & (~\new_[30131]_  | ~\s7_data_i[4] );
  assign \new_[32167]_  = ~\new_[32168]_  | ~\s13_data_i[4] ;
  assign \new_[32168]_  = \new_[31145]_  & \new_[31402]_ ;
  assign \new_[32169]_  = ~\new_[32161]_ ;
  assign \new_[32170]_  = \new_[32171]_  & \new_[4136]_ ;
  assign \new_[32171]_  = ~\new_[32172]_ ;
  assign \new_[32172]_  = ~\new_[32173]_  | ~\new_[32330]_ ;
  assign \new_[32173]_  = ~\new_[32174]_ ;
  assign \new_[32174]_  = ~\new_[6600]_  | ~\new_[7922]_ ;
  assign \new_[32175]_  = ~\new_[32182]_  | ~\new_[32179]_  | ~\new_[32176]_  | ~\new_[32177]_ ;
  assign \new_[32176]_  = ~\new_[5593]_  & ~\new_[5819]_ ;
  assign \new_[32177]_  = ~\new_[32178]_  & ~\new_[5592]_ ;
  assign \new_[32178]_  = ~\new_[5717]_  | ~\new_[5876]_ ;
  assign \new_[32179]_  = ~\new_[32180]_  & ~\new_[32181]_ ;
  assign \new_[32180]_  = ~\new_[31622]_  & ~\new_[5956]_ ;
  assign \new_[32181]_  = ~\new_[5885]_  & ~\new_[31877]_ ;
  assign \new_[32182]_  = ~\new_[6021]_  | ~\new_[4448]_ ;
  assign \new_[32183]_  = ~\new_[32184]_  | ~\new_[32189]_ ;
  assign \new_[32184]_  = ~\new_[32185]_  & ~\new_[32186]_ ;
  assign \new_[32185]_  = ~\new_[5753]_  | ~\new_[5752]_ ;
  assign \new_[32186]_  = ~\new_[32187]_  | ~\new_[32063]_ ;
  assign \new_[32187]_  = ~\new_[32188]_  | ~\new_[4064]_ ;
  assign \new_[32188]_  = ~\new_[5940]_ ;
  assign \new_[32189]_  = ~\new_[32190]_  & (~\new_[32171]_  | ~\new_[4145]_ );
  assign \new_[32190]_  = ~\new_[32064]_ ;
  assign \new_[32191]_  = ~\new_[32192]_  | ~\new_[4454]_ ;
  assign \new_[32192]_  = ~\new_[32193]_ ;
  assign \new_[32193]_  = ~\new_[32289]_  | ~\new_[32287]_ ;
  assign \m7_data_o[11]  = ~\new_[32195]_  | ~\new_[3693]_ ;
  assign \new_[32195]_  = \new_[32196]_  & \new_[32203]_ ;
  assign \new_[32196]_  = ~\new_[32197]_  & ~\new_[32198]_ ;
  assign \new_[32197]_  = ~\new_[24068]_  | ~\new_[22672]_ ;
  assign \new_[32198]_  = ~\new_[32202]_  | ~\new_[32201]_  | ~\new_[32199]_  | ~\new_[32200]_ ;
  assign \new_[32199]_  = (~\s11_data_i[11]  | ~\new_[29604]_ ) & (~\new_[30106]_  | ~\s14_data_i[11] );
  assign \new_[32200]_  = ~\new_[27347]_  | ~\s12_data_i[11] ;
  assign \new_[32201]_  = ~\new_[27337]_  | ~\s8_data_i[11] ;
  assign \new_[32202]_  = (~\s3_data_i[11]  | ~\new_[29579]_ ) & (~\new_[29534]_  | ~\s5_data_i[11] );
  assign \new_[32203]_  = \new_[27822]_  & \new_[32204]_ ;
  assign \new_[32204]_  = (~\s1_data_i[11]  | ~\new_[30124]_ ) & (~\new_[30113]_  | ~\s2_data_i[11] );
  assign \m7_data_o[5]  = ~\new_[3696]_  | ~\new_[32206]_ ;
  assign \new_[32206]_  = \new_[32207]_  & \new_[32214]_ ;
  assign \new_[32207]_  = ~\new_[32208]_  & ~\new_[32209]_ ;
  assign \new_[32208]_  = ~\new_[24004]_  | ~\new_[22588]_ ;
  assign \new_[32209]_  = ~\new_[32213]_  | ~\new_[32212]_  | ~\new_[32210]_  | ~\new_[32211]_ ;
  assign \new_[32210]_  = (~\s11_data_i[5]  | ~\new_[29604]_ ) & (~\new_[30106]_  | ~\s14_data_i[5] );
  assign \new_[32211]_  = ~\new_[27347]_  | ~\s12_data_i[5] ;
  assign \new_[32212]_  = ~\new_[27337]_  | ~\s8_data_i[5] ;
  assign \new_[32213]_  = (~\s3_data_i[5]  | ~\new_[29579]_ ) & (~\s5_data_i[5]  | ~\new_[29534]_ );
  assign \new_[32214]_  = \new_[27189]_  & \new_[32215]_ ;
  assign \new_[32215]_  = (~\s1_data_i[5]  | ~\new_[30124]_ ) & (~\new_[30113]_  | ~\s2_data_i[5] );
  assign \new_[32216]_  = ~\new_[32223]_  | ~\new_[32217]_  | ~\new_[32218]_ ;
  assign \new_[32217]_  = ~\new_[32320]_  | ~\new_[32343]_ ;
  assign \new_[32218]_  = ~\new_[32219]_ ;
  assign \new_[32219]_  = ~\new_[32222]_  | ~\new_[32220]_  | ~\new_[32221]_ ;
  assign \new_[32220]_  = (~\s6_data_i[3]  | ~\new_[29707]_ ) & (~\new_[28313]_  | ~\s7_data_i[3] );
  assign \new_[32221]_  = (~\s0_data_i[3]  | ~\new_[27879]_ ) & (~\new_[27855]_  | ~\s4_data_i[3] );
  assign \new_[32222]_  = (~\s9_data_i[3]  | ~\new_[29905]_ ) & (~\new_[29949]_  | ~\s10_data_i[3] );
  assign \new_[32223]_  = ~\new_[32338]_  | ~\s13_data_i[3] ;
  assign \m1_data_o[11]  = ~\new_[3713]_  | ~\new_[32225]_ ;
  assign \new_[32225]_  = \new_[32226]_  & \new_[32228]_ ;
  assign \new_[32226]_  = \new_[25583]_  & \new_[32227]_ ;
  assign \new_[32227]_  = (~\s1_data_i[11]  | ~\new_[30195]_ ) & (~\new_[30189]_  | ~\s2_data_i[11] );
  assign \new_[32228]_  = ~\new_[32229]_  & ~\new_[32230]_ ;
  assign \new_[32229]_  = ~\new_[25869]_  | ~\new_[25867]_ ;
  assign \new_[32230]_  = ~\new_[32234]_  | ~\new_[32233]_  | ~\new_[32231]_  | ~\new_[32232]_ ;
  assign \new_[32231]_  = (~\s3_data_i[11]  | ~\new_[30469]_ ) & (~\new_[29025]_  | ~\s5_data_i[11] );
  assign \new_[32232]_  = (~\s11_data_i[11]  | ~\new_[30260]_ ) & (~\new_[29976]_  | ~\s14_data_i[11] );
  assign \new_[32233]_  = ~\new_[28957]_  | ~\s12_data_i[11] ;
  assign \new_[32234]_  = ~\new_[29670]_  | ~\s8_data_i[11] ;
  assign \m1_data_o[5]  = ~\new_[3654]_  | ~\new_[32236]_ ;
  assign \new_[32236]_  = \new_[32237]_  & \new_[32239]_ ;
  assign \new_[32237]_  = \new_[25949]_  & \new_[32238]_ ;
  assign \new_[32238]_  = (~\s1_data_i[5]  | ~\new_[30195]_ ) & (~\new_[30189]_  | ~\s2_data_i[5] );
  assign \new_[32239]_  = ~\new_[32240]_  & ~\new_[32241]_ ;
  assign \new_[32240]_  = ~\new_[25948]_  | ~\new_[25943]_ ;
  assign \new_[32241]_  = ~\new_[32245]_  | ~\new_[32244]_  | ~\new_[32242]_  | ~\new_[32243]_ ;
  assign \new_[32242]_  = (~\s3_data_i[5]  | ~\new_[30469]_ ) & (~\new_[29025]_  | ~\s5_data_i[5] );
  assign \new_[32243]_  = (~\s11_data_i[5]  | ~\new_[30260]_ ) & (~\new_[29976]_  | ~\s14_data_i[5] );
  assign \new_[32244]_  = ~\new_[28957]_  | ~\s12_data_i[5] ;
  assign \new_[32245]_  = ~\new_[29670]_  | ~\s8_data_i[5] ;
  assign \m5_data_o[11]  = ~\new_[32247]_  | ~\new_[3665]_ ;
  assign \new_[32247]_  = \new_[32248]_  & \new_[32250]_ ;
  assign \new_[32248]_  = \new_[26110]_  & \new_[32249]_ ;
  assign \new_[32249]_  = (~\s1_data_i[11]  | ~\new_[29769]_ ) & (~\new_[30013]_  | ~\s2_data_i[11] );
  assign \new_[32250]_  = ~\new_[32251]_  & ~\new_[32256]_ ;
  assign \new_[32251]_  = ~\new_[32255]_  | ~\new_[32254]_  | ~\new_[32252]_  | ~\new_[32253]_ ;
  assign \new_[32252]_  = (~\s8_data_i[11]  | ~\new_[29636]_ ) & (~\new_[29928]_  | ~\s3_data_i[11] );
  assign \new_[32253]_  = ~\new_[28136]_  | ~\s5_data_i[11] ;
  assign \new_[32254]_  = (~\s11_data_i[11]  | ~\new_[30311]_ ) & (~\new_[30181]_  | ~\s14_data_i[11] );
  assign \new_[32255]_  = ~\new_[29640]_  | ~\s12_data_i[11] ;
  assign \new_[32256]_  = ~\new_[26008]_  | ~\new_[26130]_ ;
  assign \new_[32257]_  = ~\new_[32266]_  | ~\new_[32258]_  | ~\new_[32261]_ ;
  assign \new_[32258]_  = ~\new_[32259]_  | ~\new_[32260]_ ;
  assign \new_[32259]_  = \new_[3809]_  ? \new_[5882]_  : \s15_data_i[5] ;
  assign \new_[32260]_  = ~\new_[31498]_  & ~\new_[31552]_ ;
  assign \new_[32261]_  = ~\new_[32262]_ ;
  assign \new_[32262]_  = ~\new_[32265]_  | ~\new_[32263]_  | ~\new_[32264]_ ;
  assign \new_[32263]_  = (~\s0_data_i[5]  | ~\new_[29258]_ ) & (~\new_[29628]_  | ~\s4_data_i[5] );
  assign \new_[32264]_  = (~\s6_data_i[5]  | ~\new_[29704]_ ) & (~\new_[30060]_  | ~\s7_data_i[5] );
  assign \new_[32265]_  = (~\s9_data_i[5]  | ~\new_[29951]_ ) & (~\new_[29045]_  | ~\s10_data_i[5] );
  assign \new_[32266]_  = ~\new_[32267]_  | ~\s13_data_i[5] ;
  assign \new_[32267]_  = ~\new_[31552]_  & ~\new_[30954]_ ;
  assign \new_[32268]_  = ~\new_[32260]_ ;
  assign \new_[32269]_  = ~\new_[32275]_  | (~\new_[32270]_  & ~\new_[32273]_ );
  assign \new_[32270]_  = ~\new_[4887]_  | ~\new_[32271]_  | ~\new_[32272]_ ;
  assign \new_[32271]_  = ~\new_[5785]_  & ~\new_[32060]_ ;
  assign \new_[32272]_  = ~\new_[32059]_  & ~\new_[32058]_ ;
  assign \new_[32273]_  = ~\new_[5554]_  | ~\new_[4739]_ ;
  assign \new_[32274]_  = \new_[32340]_ ;
  assign \new_[32275]_  = ~\new_[32274]_ ;
  assign \new_[32276]_  = (~\s13_data_i[29]  | ~\new_[32327]_ ) & (~\new_[32277]_  | ~\new_[32321]_ );
  assign \new_[32277]_  = \new_[32278]_  & \s15_data_i[29] ;
  assign \new_[32278]_  = \new_[32279]_ ;
  assign \new_[32279]_  = ~\new_[32280]_  | ~\new_[32281]_ ;
  assign \new_[32280]_  = ~\new_[32336]_ ;
  assign \new_[32281]_  = ~\new_[32335]_ ;
  assign \new_[32282]_  = ~\new_[32283]_ ;
  assign \new_[32283]_  = ~\new_[32280]_  | ~\new_[32281]_ ;
  assign \new_[32284]_  = ~\new_[32285]_  | ~\new_[4454]_ ;
  assign \new_[32285]_  = ~\new_[32286]_ ;
  assign \new_[32286]_  = ~\new_[32287]_  | ~\new_[32333]_ ;
  assign \new_[32287]_  = ~\new_[32293]_ ;
  assign \new_[32288]_  = \new_[32285]_ ;
  assign \new_[32289]_  = \new_[32291]_  & \s15_addr_o[4] ;
  assign \s15_addr_o[4]  = ~\new_[14457]_  | ~\new_[14459]_  | ~\new_[14456]_  | ~\new_[14460]_ ;
  assign \new_[32291]_  = ~\new_[32304]_ ;
  assign \s15_addr_o[5]  = ~\new_[32304]_ ;
  assign \new_[32293]_  = ~\s15_addr_o[3]  | ~\new_[32294]_ ;
  assign \new_[32294]_  = ~\s15_addr_o[2] ;
  assign \new_[32295]_  = ~\new_[15996]_  & ~\new_[15998]_ ;
  assign \new_[32296]_  = ~\new_[32297]_  & (~\new_[17312]_  | ~\m4_addr_i[2] );
  assign \new_[32297]_  = \new_[17341]_  & \m6_addr_i[2] ;
  assign \new_[32298]_  = ~\new_[15992]_  & ~\new_[15993]_ ;
  assign \new_[32299]_  = ~\new_[32300]_  & (~\new_[17256]_  | ~\m1_addr_i[2] );
  assign \new_[32300]_  = \new_[17226]_  & \m3_addr_i[2] ;
  assign \new_[32301]_  = ~\new_[32302]_  & (~\new_[4087]_  | ~\new_[5943]_ );
  assign \new_[32302]_  = ~\new_[32303]_  | (~\new_[5938]_  & ~\new_[31728]_ );
  assign \new_[32303]_  = ~\new_[32068]_  | ~\new_[4154]_ ;
  assign \new_[32304]_  = ~\new_[32305]_  & ~\new_[32306]_ ;
  assign \new_[32305]_  = ~\new_[15988]_  | ~\new_[15989]_  | ~\new_[14591]_  | ~\new_[14592]_ ;
  assign \new_[32306]_  = ~\new_[32312]_  | ~\new_[32311]_  | ~\new_[32307]_  | ~\new_[32310]_ ;
  assign \new_[32307]_  = ~\new_[32349]_  | ~\m0_addr_i[5] ;
  assign \new_[32308]_  = ~\new_[32309]_  | ~\new_[21244]_ ;
  assign \new_[32309]_  = \new_[21250]_  & \new_[22411]_ ;
  assign \new_[32310]_  = ~\new_[17257]_  | ~\m1_addr_i[5] ;
  assign \new_[32311]_  = ~\new_[17326]_  | ~\m2_addr_i[5] ;
  assign \new_[32312]_  = ~\m3_addr_i[5]  | ~\new_[21241]_  | ~\new_[19377]_  | ~\new_[21049]_ ;
  assign \new_[32313]_  = ~\new_[28075]_  | ~\new_[30120]_  | ~\new_[28710]_  | ~\new_[28239]_ ;
  assign \new_[32314]_  = ~\new_[28075]_  | ~\new_[30120]_  | ~\new_[28710]_  | ~\new_[28239]_ ;
  assign \new_[32315]_  = \new_[32342]_ ;
  assign \new_[32316]_  = ~\new_[6374]_  | ~\new_[32287]_ ;
  assign \new_[32317]_  = ~\new_[6374]_  | ~\new_[32287]_ ;
  assign \new_[32318]_  = ~\new_[32326]_  | ~\new_[32325]_  | ~\new_[32319]_  | ~\new_[32322]_ ;
  assign \new_[32319]_  = ~\new_[32320]_  | ~\new_[32321]_ ;
  assign \new_[32320]_  = \new_[3824]_  ? \new_[5882]_  : \s15_data_i[3] ;
  assign \new_[32321]_  = ~\new_[31467]_  & ~\new_[31327]_ ;
  assign \new_[32322]_  = \new_[32323]_  & \new_[32324]_ ;
  assign \new_[32323]_  = (~\s0_data_i[3]  | ~\new_[29434]_ ) & (~\new_[28842]_  | ~\s4_data_i[3] );
  assign \new_[32324]_  = (~\s6_data_i[3]  | ~\new_[29052]_ ) & (~\new_[30031]_  | ~\s7_data_i[3] );
  assign \new_[32325]_  = (~\s9_data_i[3]  | ~\new_[30354]_ ) & (~\new_[29705]_  | ~\s10_data_i[3] );
  assign \new_[32326]_  = ~\new_[32327]_  | ~\s13_data_i[3] ;
  assign \new_[32327]_  = ~\new_[30985]_  & ~\new_[31327]_ ;
  assign \new_[32328]_  = ~\new_[32321]_ ;
  assign \new_[32329]_  = ~\new_[32330]_  | ~\new_[32333]_ ;
  assign \new_[32330]_  = \new_[32331]_ ;
  assign \new_[32331]_  = ~\new_[32294]_  & (~\new_[9318]_  | ~\new_[8474]_ );
  assign \s15_addr_o[2]  = ~\new_[32299]_  | ~\new_[32298]_  | ~\new_[32296]_  | ~\new_[32295]_ ;
  assign \new_[32333]_  = \s15_addr_o[5]  & \new_[7921]_ ;
  assign \s15_addr_o[3]  = ~\new_[9318]_  | ~\new_[8474]_ ;
  assign \new_[32335]_  = ~\new_[7218]_  | ~s15_stb_o | ~\s15_addr_o[25] ;
  assign \new_[32336]_  = ~\s15_addr_o[24]  | ~\s15_addr_o[26]  | ~\s15_addr_o[27] ;
  assign \new_[32337]_  = (~\s13_data_i[31]  | ~\new_[32338]_ ) & (~\new_[32339]_  | ~\new_[32343]_ );
  assign \new_[32338]_  = ~\new_[31355]_  & ~\new_[31141]_ ;
  assign \new_[32339]_  = \new_[32340]_  & \s15_data_i[31] ;
  assign \new_[32340]_  = ~\new_[32341]_ ;
  assign \new_[32341]_  = \new_[32342]_ ;
  assign \new_[32342]_  = ~\new_[32335]_  & ~\new_[32336]_ ;
  assign \new_[32343]_  = ~\new_[31355]_  & ~\new_[30454]_ ;
  assign \new_[32344]_  = ~\new_[32343]_ ;
  assign \new_[32345]_  = ~\new_[32348]_ ;
  assign \new_[32346]_  = \new_[32347]_ ;
  assign \new_[32347]_  = \new_[32348]_ ;
  assign \new_[32348]_  = ~\new_[32308]_ ;
  assign \new_[32349]_  = ~\new_[32308]_ ;
  assign \new_[32350]_  = ~\new_[32351]_ ;
  assign \new_[32351]_  = ~\new_[18936]_ ;
  always @ (posedge clock) begin
    \\rf_rf_dout_reg[14]  <= n5094;
    \\rf_rf_dout_reg[12]  <= n5099;
    \\rf_rf_dout_reg[11]  <= n5104;
    \\rf_rf_dout_reg[9]  <= n5109;
    \\rf_rf_dout_reg[6]  <= n5114;
    \\rf_rf_dout_reg[5]  <= n5119;
    \\rf_rf_dout_reg[4]  <= n5124;
    \\rf_rf_dout_reg[2]  <= n5129;
    \\rf_rf_dout_reg[1]  <= n5134;
    \\rf_rf_dout_reg[15]  <= n5139;
    \\rf_rf_dout_reg[13]  <= n5144;
    \\rf_rf_dout_reg[10]  <= n5149;
    \\rf_rf_dout_reg[8]  <= n5154;
    \\rf_rf_dout_reg[7]  <= n5159;
    \\rf_rf_dout_reg[3]  <= n5164;
    \\rf_rf_dout_reg[0]  <= n5169;
    \\rf_conf15_reg[0]  <= n5174;
    \\rf_conf15_reg[10]  <= n5179;
    \\rf_conf15_reg[11]  <= n5184;
    \\rf_conf15_reg[12]  <= n5189;
    \\rf_conf15_reg[13]  <= n5194;
    \\rf_conf15_reg[14]  <= n5199;
    \\rf_conf15_reg[15]  <= n5204;
    \\rf_conf15_reg[1]  <= n5209;
    \\rf_conf15_reg[2]  <= n5214;
    \\rf_conf15_reg[3]  <= n5219;
    \\rf_conf15_reg[4]  <= n5224;
    \\rf_conf15_reg[5]  <= n5229;
    \\rf_conf15_reg[6]  <= n5234;
    \\rf_conf15_reg[7]  <= n5239;
    \\rf_conf15_reg[8]  <= n5244;
    \\rf_conf15_reg[9]  <= n5249;
    \\rf_conf0_reg[0]  <= n5254;
    \\rf_conf0_reg[10]  <= n5259;
    \\rf_conf0_reg[11]  <= n5264;
    \\rf_conf0_reg[12]  <= n5269;
    \\rf_conf0_reg[13]  <= n5274;
    \\rf_conf0_reg[14]  <= n5279;
    \\rf_conf0_reg[15]  <= n5284;
    \\rf_conf0_reg[1]  <= n5289;
    \\rf_conf0_reg[2]  <= n5294;
    \\rf_conf0_reg[3]  <= n5299;
    \\rf_conf0_reg[4]  <= n5304;
    \\rf_conf0_reg[5]  <= n5309;
    \\rf_conf0_reg[6]  <= n5314;
    \\rf_conf0_reg[7]  <= n5319;
    \\rf_conf0_reg[8]  <= n5324;
    \\rf_conf0_reg[9]  <= n5329;
    \\rf_conf12_reg[0]  <= n5334;
    \\rf_conf12_reg[10]  <= n5339;
    \\rf_conf12_reg[11]  <= n5344;
    \\rf_conf12_reg[12]  <= n5349;
    \\rf_conf12_reg[13]  <= n5354;
    \\rf_conf12_reg[14]  <= n5359;
    \\rf_conf12_reg[15]  <= n5364;
    \\rf_conf12_reg[1]  <= n5369;
    \\rf_conf12_reg[2]  <= n5374;
    \\rf_conf12_reg[3]  <= n5379;
    \\rf_conf12_reg[4]  <= n5384;
    \\rf_conf12_reg[5]  <= n5389;
    \\rf_conf12_reg[6]  <= n5394;
    \\rf_conf12_reg[7]  <= n5399;
    \\rf_conf12_reg[8]  <= n5404;
    \\rf_conf12_reg[9]  <= n5409;
    \\rf_conf13_reg[0]  <= n5414;
    \\rf_conf13_reg[10]  <= n5419;
    \\rf_conf13_reg[11]  <= n5424;
    \\rf_conf13_reg[12]  <= n5429;
    \\rf_conf13_reg[13]  <= n5434;
    \\rf_conf13_reg[14]  <= n5439;
    \\rf_conf13_reg[15]  <= n5444;
    \\rf_conf13_reg[1]  <= n5449;
    \\rf_conf13_reg[4]  <= n5454;
    \\rf_conf13_reg[5]  <= n5459;
    \\rf_conf13_reg[6]  <= n5464;
    \\rf_conf13_reg[7]  <= n5469;
    \\rf_conf13_reg[8]  <= n5474;
    \\rf_conf13_reg[9]  <= n5479;
    \\rf_conf14_reg[0]  <= n5484;
    \\rf_conf14_reg[10]  <= n5489;
    \\rf_conf14_reg[11]  <= n5494;
    \\rf_conf14_reg[12]  <= n5499;
    \\rf_conf14_reg[13]  <= n5504;
    \\rf_conf14_reg[14]  <= n5509;
    \\rf_conf14_reg[15]  <= n5514;
    \\rf_conf14_reg[1]  <= n5519;
    \\rf_conf14_reg[3]  <= n5524;
    \\rf_conf14_reg[4]  <= n5529;
    \\rf_conf14_reg[5]  <= n5534;
    \\rf_conf14_reg[6]  <= n5539;
    \\rf_conf14_reg[7]  <= n5544;
    \\rf_conf14_reg[8]  <= n5549;
    \\rf_conf14_reg[9]  <= n5554;
    \\rf_conf13_reg[2]  <= n5559;
    \\rf_conf13_reg[3]  <= n5564;
    \\rf_conf14_reg[2]  <= n5569;
    \\rf_conf1_reg[0]  <= n5574;
    \\rf_conf1_reg[10]  <= n5579;
    \\rf_conf1_reg[11]  <= n5584;
    \\rf_conf1_reg[12]  <= n5589;
    \\rf_conf1_reg[13]  <= n5594;
    \\rf_conf1_reg[14]  <= n5599;
    \\rf_conf1_reg[15]  <= n5604;
    \\rf_conf1_reg[1]  <= n5609;
    \\rf_conf1_reg[2]  <= n5614;
    \\rf_conf1_reg[3]  <= n5619;
    \\rf_conf1_reg[4]  <= n5624;
    \\rf_conf1_reg[5]  <= n5629;
    \\rf_conf1_reg[6]  <= n5634;
    \\rf_conf1_reg[7]  <= n5639;
    \\rf_conf1_reg[8]  <= n5644;
    \\rf_conf1_reg[9]  <= n5649;
    \\rf_conf2_reg[0]  <= n5654;
    \\rf_conf2_reg[10]  <= n5659;
    \\rf_conf2_reg[11]  <= n5664;
    \\rf_conf2_reg[12]  <= n5669;
    \\rf_conf2_reg[13]  <= n5674;
    \\rf_conf2_reg[14]  <= n5679;
    \\rf_conf2_reg[15]  <= n5684;
    \\rf_conf2_reg[1]  <= n5689;
    \\rf_conf2_reg[2]  <= n5694;
    \\rf_conf2_reg[3]  <= n5699;
    \\rf_conf2_reg[4]  <= n5704;
    \\rf_conf2_reg[5]  <= n5709;
    \\rf_conf2_reg[6]  <= n5714;
    \\rf_conf2_reg[7]  <= n5719;
    \\rf_conf2_reg[8]  <= n5724;
    \\rf_conf2_reg[9]  <= n5729;
    \\rf_conf3_reg[0]  <= n5734;
    \\rf_conf3_reg[10]  <= n5739;
    \\rf_conf3_reg[11]  <= n5744;
    \\rf_conf3_reg[12]  <= n5749;
    \\rf_conf3_reg[13]  <= n5754;
    \\rf_conf3_reg[14]  <= n5759;
    \\rf_conf3_reg[15]  <= n5764;
    \\rf_conf3_reg[1]  <= n5769;
    \\rf_conf3_reg[2]  <= n5774;
    \\rf_conf3_reg[3]  <= n5779;
    \\rf_conf3_reg[4]  <= n5784;
    \\rf_conf3_reg[5]  <= n5789;
    \\rf_conf3_reg[6]  <= n5794;
    \\rf_conf3_reg[7]  <= n5799;
    \\rf_conf3_reg[8]  <= n5804;
    \\rf_conf3_reg[9]  <= n5809;
    \\rf_conf5_reg[0]  <= n5814;
    \\rf_conf5_reg[10]  <= n5819;
    \\rf_conf5_reg[11]  <= n5824;
    \\rf_conf5_reg[12]  <= n5829;
    \\rf_conf5_reg[13]  <= n5834;
    \\rf_conf5_reg[14]  <= n5839;
    \\rf_conf5_reg[15]  <= n5844;
    \\rf_conf5_reg[1]  <= n5849;
    \\rf_conf5_reg[2]  <= n5854;
    \\rf_conf5_reg[3]  <= n5859;
    \\rf_conf5_reg[4]  <= n5864;
    \\rf_conf5_reg[5]  <= n5869;
    \\rf_conf5_reg[6]  <= n5874;
    \\rf_conf5_reg[7]  <= n5879;
    \\rf_conf5_reg[8]  <= n5884;
    \\rf_conf5_reg[9]  <= n5889;
    \\rf_conf7_reg[0]  <= n5894;
    \\rf_conf7_reg[10]  <= n5899;
    \\rf_conf7_reg[11]  <= n5904;
    \\rf_conf7_reg[12]  <= n5909;
    \\rf_conf7_reg[13]  <= n5914;
    \\rf_conf7_reg[14]  <= n5919;
    \\rf_conf7_reg[15]  <= n5924;
    \\rf_conf7_reg[1]  <= n5929;
    \\rf_conf7_reg[2]  <= n5934;
    \\rf_conf7_reg[3]  <= n5939;
    \\rf_conf7_reg[4]  <= n5944;
    \\rf_conf7_reg[5]  <= n5949;
    \\rf_conf7_reg[6]  <= n5954;
    \\rf_conf7_reg[7]  <= n5959;
    \\rf_conf7_reg[8]  <= n5964;
    \\rf_conf7_reg[9]  <= n5969;
    \\rf_conf10_reg[0]  <= n5974;
    \\rf_conf10_reg[10]  <= n5979;
    \\rf_conf10_reg[11]  <= n5984;
    \\rf_conf10_reg[12]  <= n5989;
    \\rf_conf10_reg[13]  <= n5994;
    \\rf_conf10_reg[14]  <= n5999;
    \\rf_conf10_reg[15]  <= n6004;
    \\rf_conf10_reg[1]  <= n6009;
    \\rf_conf10_reg[2]  <= n6014;
    \\rf_conf10_reg[3]  <= n6019;
    \\rf_conf10_reg[4]  <= n6024;
    \\rf_conf10_reg[5]  <= n6029;
    \\rf_conf10_reg[6]  <= n6034;
    \\rf_conf10_reg[7]  <= n6039;
    \\rf_conf10_reg[8]  <= n6044;
    \\rf_conf10_reg[9]  <= n6049;
    \\rf_conf11_reg[0]  <= n6054;
    \\rf_conf11_reg[10]  <= n6059;
    \\rf_conf11_reg[11]  <= n6064;
    \\rf_conf11_reg[12]  <= n6069;
    \\rf_conf11_reg[13]  <= n6074;
    \\rf_conf11_reg[14]  <= n6079;
    \\rf_conf11_reg[15]  <= n6084;
    \\rf_conf11_reg[1]  <= n6089;
    \\rf_conf11_reg[4]  <= n6094;
    \\rf_conf11_reg[5]  <= n6099;
    \\rf_conf11_reg[6]  <= n6104;
    \\rf_conf11_reg[7]  <= n6109;
    \\rf_conf11_reg[8]  <= n6114;
    \\rf_conf11_reg[9]  <= n6119;
    \\rf_conf11_reg[2]  <= n6124;
    \\rf_conf11_reg[3]  <= n6129;
    \\rf_conf4_reg[0]  <= n6134;
    \\rf_conf4_reg[10]  <= n6139;
    \\rf_conf4_reg[11]  <= n6144;
    \\rf_conf4_reg[12]  <= n6149;
    \\rf_conf4_reg[13]  <= n6154;
    \\rf_conf4_reg[14]  <= n6159;
    \\rf_conf4_reg[15]  <= n6164;
    \\rf_conf4_reg[1]  <= n6169;
    \\rf_conf4_reg[4]  <= n6174;
    \\rf_conf4_reg[5]  <= n6179;
    \\rf_conf4_reg[6]  <= n6184;
    \\rf_conf4_reg[7]  <= n6189;
    \\rf_conf4_reg[8]  <= n6194;
    \\rf_conf4_reg[9]  <= n6199;
    \\rf_conf4_reg[2]  <= n6204;
    \\rf_conf4_reg[3]  <= n6209;
    \\rf_conf6_reg[0]  <= n6214;
    \\rf_conf6_reg[10]  <= n6219;
    \\rf_conf6_reg[11]  <= n6224;
    \\rf_conf6_reg[12]  <= n6229;
    \\rf_conf6_reg[13]  <= n6234;
    \\rf_conf6_reg[14]  <= n6239;
    \\rf_conf6_reg[15]  <= n6244;
    \\rf_conf6_reg[1]  <= n6249;
    \\rf_conf6_reg[4]  <= n6254;
    \\rf_conf6_reg[5]  <= n6259;
    \\rf_conf6_reg[6]  <= n6264;
    \\rf_conf6_reg[7]  <= n6269;
    \\rf_conf6_reg[8]  <= n6274;
    \\rf_conf6_reg[9]  <= n6279;
    \\rf_conf6_reg[2]  <= n6284;
    \\rf_conf6_reg[3]  <= n6289;
    \\rf_conf9_reg[0]  <= n6294;
    \\rf_conf9_reg[10]  <= n6299;
    \\rf_conf9_reg[11]  <= n6304;
    \\rf_conf9_reg[12]  <= n6309;
    \\rf_conf9_reg[13]  <= n6314;
    \\rf_conf9_reg[14]  <= n6319;
    \\rf_conf9_reg[15]  <= n6324;
    \\rf_conf9_reg[1]  <= n6329;
    \\rf_conf9_reg[2]  <= n6334;
    \\rf_conf9_reg[3]  <= n6339;
    \\rf_conf9_reg[4]  <= n6344;
    \\rf_conf9_reg[5]  <= n6349;
    \\rf_conf9_reg[6]  <= n6354;
    \\rf_conf9_reg[7]  <= n6359;
    \\rf_conf9_reg[8]  <= n6364;
    \\rf_conf9_reg[9]  <= n6369;
    \\rf_conf8_reg[0]  <= n6374;
    \\rf_conf8_reg[10]  <= n6379;
    \\rf_conf8_reg[11]  <= n6384;
    \\rf_conf8_reg[12]  <= n6389;
    \\rf_conf8_reg[13]  <= n6394;
    \\rf_conf8_reg[14]  <= n6399;
    \\rf_conf8_reg[15]  <= n6404;
    \\rf_conf8_reg[1]  <= n6409;
    \\rf_conf8_reg[4]  <= n6414;
    \\rf_conf8_reg[5]  <= n6419;
    \\rf_conf8_reg[6]  <= n6424;
    \\rf_conf8_reg[7]  <= n6429;
    \\rf_conf8_reg[8]  <= n6434;
    \\rf_conf8_reg[9]  <= n6439;
    \\rf_conf8_reg[2]  <= n6444;
    \\rf_conf8_reg[3]  <= n6449;
    rf_rf_we_reg <= n6454;
    rf_rf_ack_reg <= n6459;
    \\s14_msel_arb2_state_reg[0]  <= n6464;
    \\s10_msel_arb0_state_reg[1]  <= n6469;
    \\s11_msel_arb0_state_reg[1]  <= n6474;
    \\s12_msel_arb0_state_reg[1]  <= n6479;
    \\s13_msel_arb0_state_reg[1]  <= n6484;
    \\s14_msel_arb0_state_reg[1]  <= n6489;
    \\s15_msel_arb0_state_reg[1]  <= n6494;
    \\s1_msel_arb0_state_reg[1]  <= n6499;
    \\s2_msel_arb0_state_reg[1]  <= n6504;
    \\s3_msel_arb0_state_reg[1]  <= n6509;
    \\s4_msel_arb0_state_reg[1]  <= n6514;
    \\s5_msel_arb0_state_reg[1]  <= n6519;
    \\s6_msel_arb0_state_reg[1]  <= n6524;
    \\s8_msel_arb0_state_reg[1]  <= n6529;
    \\s9_msel_arb0_state_reg[1]  <= n6534;
    \\s0_msel_arb0_state_reg[1]  <= n6539;
    \\s11_msel_arb0_state_reg[0]  <= n6544;
    \\s11_msel_arb1_state_reg[1]  <= n6549;
    \\s12_msel_arb0_state_reg[0]  <= n6554;
    \\s13_msel_arb0_state_reg[0]  <= n6559;
    \\s13_msel_arb2_state_reg[0]  <= n6564;
    \\s14_msel_arb0_state_reg[0]  <= n6569;
    \\s15_msel_arb2_state_reg[0]  <= n6574;
    \\s15_msel_arb3_state_reg[1]  <= n6579;
    \\s3_msel_arb0_state_reg[0]  <= n6584;
    \\s4_msel_arb0_state_reg[0]  <= n6589;
    \\s4_msel_arb2_state_reg[0]  <= n6594;
    \\s4_msel_arb2_state_reg[1]  <= n6599;
    \\s5_msel_arb0_state_reg[0]  <= n6604;
    \\s5_msel_arb3_state_reg[1]  <= n6609;
    \\s6_msel_arb0_state_reg[0]  <= n6614;
    \\s6_msel_arb1_state_reg[0]  <= n6619;
    \\s6_msel_arb1_state_reg[1]  <= n6624;
    \\s7_msel_arb0_state_reg[0]  <= n6629;
    \\s8_msel_arb0_state_reg[0]  <= n6634;
    \\s8_msel_arb1_state_reg[1]  <= n6639;
    \\s8_msel_arb3_state_reg[1]  <= n6644;
    \\s9_msel_arb3_state_reg[0]  <= n6649;
    \\s9_msel_arb2_state_reg[0]  <= n6654;
    \\s0_msel_arb2_state_reg[0]  <= n6659;
    \\s7_msel_arb0_state_reg[1]  <= n6664;
    \\s10_msel_arb2_state_reg[1]  <= n6669;
    \\s10_msel_arb2_state_reg[0]  <= n6674;
    \\s11_msel_arb2_state_reg[1]  <= n6679;
    \\s11_msel_arb3_state_reg[1]  <= n6684;
    \\s12_msel_arb1_state_reg[1]  <= n6689;
    \\s12_msel_arb2_state_reg[0]  <= n6694;
    \\s12_msel_arb2_state_reg[1]  <= n6699;
    \\s13_msel_arb1_state_reg[1]  <= n6704;
    \\s13_msel_arb2_state_reg[1]  <= n6709;
    \\s14_msel_arb2_state_reg[1]  <= n6714;
    \\s14_msel_arb2_state_reg[2]  <= n6719;
    \\s15_msel_arb0_state_reg[0]  <= n6724;
    \\s15_msel_arb1_state_reg[1]  <= n6729;
    \\s15_msel_arb2_state_reg[1]  <= n6734;
    \\s15_msel_arb2_state_reg[2]  <= n6739;
    \\s1_msel_arb0_state_reg[0]  <= n6744;
    \\s1_msel_arb2_state_reg[0]  <= n6749;
    \\s1_msel_arb2_state_reg[1]  <= n6754;
    \\s2_msel_arb2_state_reg[0]  <= n6759;
    \\s2_msel_arb2_state_reg[1]  <= n6764;
    \\s2_msel_arb0_state_reg[0]  <= n6769;
    \\s3_msel_arb1_state_reg[1]  <= n6774;
    \\s3_msel_arb2_state_reg[0]  <= n6779;
    \\s3_msel_arb2_state_reg[1]  <= n6784;
    \\s3_msel_arb3_state_reg[1]  <= n6789;
    \\s4_msel_arb2_state_reg[2]  <= n6794;
    \\s5_msel_arb1_state_reg[1]  <= n6799;
    \\s5_msel_arb2_state_reg[1]  <= n6804;
    \\s5_msel_arb3_state_reg[0]  <= n6809;
    \\s5_msel_arb3_state_reg[2]  <= n6814;
    \\s6_msel_arb2_state_reg[1]  <= n6819;
    \\s6_msel_arb2_state_reg[0]  <= n6824;
    \\s6_msel_arb3_state_reg[1]  <= n6829;
    \\s6_msel_arb3_state_reg[0]  <= n6834;
    \\s7_msel_arb2_state_reg[0]  <= n6839;
    \\s7_msel_arb2_state_reg[1]  <= n6844;
    \\s8_msel_arb2_state_reg[0]  <= n6849;
    \\s8_msel_arb2_state_reg[1]  <= n6854;
    \\s8_msel_arb3_state_reg[0]  <= n6859;
    \\s9_msel_arb0_state_reg[0]  <= n6864;
    \\s9_msel_arb2_state_reg[2]  <= n6869;
    \\s0_msel_arb0_state_reg[0]  <= n6874;
    \\s0_msel_arb2_state_reg[1]  <= n6879;
    \\s0_msel_arb2_state_reg[2]  <= n6884;
    \\s0_msel_arb3_state_reg[0]  <= n6889;
    \\s14_msel_arb3_state_reg[0]  <= n6894;
    \\s12_msel_arb1_state_reg[0]  <= n6899;
    \\s10_msel_arb1_state_reg[0]  <= n6904;
    \\s10_msel_arb1_state_reg[1]  <= n6909;
    \\s10_msel_arb2_state_reg[2]  <= n6914;
    \\s11_msel_arb0_state_reg[2]  <= n6919;
    \\s11_msel_arb1_state_reg[2]  <= n6924;
    \\s11_msel_arb2_state_reg[0]  <= n6929;
    \\s11_msel_arb2_state_reg[2]  <= n6934;
    \\s11_msel_arb1_state_reg[0]  <= n6939;
    \\s11_msel_arb3_state_reg[2]  <= n6944;
    \\s12_msel_arb0_state_reg[2]  <= n6949;
    \\s12_msel_arb1_state_reg[2]  <= n6954;
    \\s12_msel_arb2_state_reg[2]  <= n6959;
    \\s13_msel_arb0_state_reg[2]  <= n6964;
    \\s12_msel_arb3_state_reg[1]  <= n6969;
    \\s13_msel_arb2_state_reg[2]  <= n6974;
    \\s13_msel_arb3_state_reg[1]  <= n6979;
    \\s14_msel_arb1_state_reg[2]  <= n6984;
    \\s14_msel_arb1_state_reg[1]  <= n6989;
    \\s14_msel_arb0_state_reg[2]  <= n6994;
    \\s14_msel_arb3_state_reg[1]  <= n6999;
    \\s14_msel_arb3_state_reg[2]  <= n7004;
    \\s15_msel_arb1_state_reg[0]  <= n7009;
    \\s15_msel_arb3_state_reg[0]  <= n7014;
    \\s1_msel_arb0_state_reg[2]  <= n7019;
    \\s1_msel_arb1_state_reg[1]  <= n7024;
    \\s1_msel_arb2_state_reg[2]  <= n7029;
    \\s1_msel_arb3_state_reg[0]  <= n7034;
    \\s1_msel_arb3_state_reg[1]  <= n7039;
    \\s2_msel_arb1_state_reg[1]  <= n7044;
    \\s2_msel_arb0_state_reg[2]  <= n7049;
    \\s2_msel_arb2_state_reg[2]  <= n7054;
    \\s2_msel_arb3_state_reg[0]  <= n7059;
    \\s2_msel_arb3_state_reg[1]  <= n7064;
    \\s3_msel_arb1_state_reg[0]  <= n7069;
    \\s3_msel_arb0_state_reg[2]  <= n7074;
    \\s3_msel_arb2_state_reg[2]  <= n7079;
    \\s4_msel_arb1_state_reg[0]  <= n7084;
    \\s4_msel_arb1_state_reg[1]  <= n7089;
    \\s4_msel_arb3_state_reg[0]  <= n7094;
    \\s5_msel_arb1_state_reg[0]  <= n7099;
    \\s5_msel_arb1_state_reg[2]  <= n7104;
    \\s5_msel_arb0_state_reg[2]  <= n7109;
    \\s6_msel_arb0_state_reg[2]  <= n7114;
    \\s6_msel_arb1_state_reg[2]  <= n7119;
    \\s6_msel_arb2_state_reg[2]  <= n7124;
    \\s7_msel_arb1_state_reg[0]  <= n7129;
    \\s7_msel_arb1_state_reg[2]  <= n7134;
    \\s7_msel_arb0_state_reg[2]  <= n7139;
    \\s7_msel_arb2_state_reg[2]  <= n7144;
    \\s7_msel_arb3_state_reg[2]  <= n7149;
    \\s8_msel_arb0_state_reg[2]  <= n7154;
    \\s8_msel_arb1_state_reg[0]  <= n7159;
    \\s7_msel_arb3_state_reg[1]  <= n7164;
    \\s8_msel_arb3_state_reg[2]  <= n7169;
    \\s9_msel_arb0_state_reg[2]  <= n7174;
    \\s9_msel_arb2_state_reg[1]  <= n7179;
    \\s9_msel_arb1_state_reg[2]  <= n7184;
    \\s9_msel_arb3_state_reg[1]  <= n7189;
    \\s0_msel_arb0_state_reg[2]  <= n7194;
    \\s0_msel_arb1_state_reg[1]  <= n7199;
    \\s0_msel_arb1_state_reg[2]  <= n7204;
    \\s10_msel_arb0_state_reg[0]  <= n7209;
    \\s0_msel_arb3_state_reg[2]  <= n7214;
    \\s13_msel_arb1_state_reg[0]  <= n7219;
    \\s10_msel_arb1_state_reg[2]  <= n7224;
    \\s11_msel_arb3_state_reg[0]  <= n7229;
    \\s9_msel_arb3_state_reg[2]  <= n7234;
    \\s9_msel_arb1_state_reg[0]  <= n7239;
    \\s8_msel_arb2_state_reg[2]  <= n7244;
    \\s8_msel_arb1_state_reg[2]  <= n7249;
    \\s5_msel_arb2_state_reg[2]  <= n7254;
    \\s5_msel_arb2_state_reg[0]  <= n7259;
    \\s4_msel_arb1_state_reg[2]  <= n7264;
    \\s4_msel_arb3_state_reg[1]  <= n7269;
    \\s4_msel_arb0_state_reg[2]  <= n7274;
    \\s3_msel_arb1_state_reg[2]  <= n7279;
    \\s1_msel_arb3_state_reg[2]  <= n7284;
    \\s1_msel_arb1_state_reg[0]  <= n7289;
    \\s1_msel_arb1_state_reg[2]  <= n7294;
    \\s13_msel_arb1_state_reg[2]  <= n7299;
    \\s13_msel_arb3_state_reg[2]  <= n7304;
    \\s10_msel_arb0_state_reg[2]  <= n7309;
    \\s10_msel_arb3_state_reg[2]  <= n7314;
    \\s12_msel_arb3_state_reg[0]  <= n7319;
    \\s12_msel_arb3_state_reg[2]  <= n7324;
    \\s13_msel_arb3_state_reg[0]  <= n7329;
    \\s14_msel_arb1_state_reg[0]  <= n7334;
    \\s15_msel_arb1_state_reg[2]  <= n7339;
    \\s15_msel_arb3_state_reg[2]  <= n7344;
    \\s2_msel_arb1_state_reg[0]  <= n7349;
    \\s2_msel_arb1_state_reg[2]  <= n7354;
    \\s3_msel_arb3_state_reg[0]  <= n7359;
    \\s3_msel_arb3_state_reg[2]  <= n7364;
    \\s4_msel_arb3_state_reg[2]  <= n7369;
    \\s9_msel_arb1_state_reg[1]  <= n7374;
    \\s0_msel_arb1_state_reg[0]  <= n7379;
    \\s0_msel_arb3_state_reg[1]  <= n7384;
    \\s10_msel_arb3_state_reg[1]  <= n7389;
    \\s10_msel_arb3_state_reg[0]  <= n7394;
    \\s6_msel_arb3_state_reg[2]  <= n7399;
    \\s7_msel_arb3_state_reg[0]  <= n7404;
    \\s7_msel_arb1_state_reg[1]  <= n7409;
    \\s15_msel_arb0_state_reg[2]  <= n7414;
    \\s2_msel_arb3_state_reg[2]  <= n7419;
    s15_next_reg <= n7424;
    \\s13_msel_pri_out_reg[0]  <= n7429;
    \\s3_msel_pri_out_reg[0]  <= n7434;
    \\s11_msel_pri_out_reg[0]  <= n7439;
    \\s12_msel_pri_out_reg[0]  <= n7444;
    \\s5_msel_pri_out_reg[0]  <= n7449;
    \\s6_msel_pri_out_reg[0]  <= n7454;
    \\s8_msel_pri_out_reg[0]  <= n7459;
    s12_next_reg <= n7464;
    s13_next_reg <= n7469;
    s14_next_reg <= n7474;
    s3_next_reg <= n7479;
    s6_next_reg <= n7484;
    s9_next_reg <= n7489;
    s8_next_reg <= n7494;
    s0_next_reg <= n7499;
    \\s8_msel_pri_out_reg[1]  <= n7504;
    \\s15_msel_pri_out_reg[0]  <= n7509;
    \\s2_msel_pri_out_reg[0]  <= n7514;
    \\s1_msel_pri_out_reg[0]  <= n7519;
    \\s7_msel_pri_out_reg[0]  <= n7524;
    \\s9_msel_pri_out_reg[0]  <= n7529;
    \\s0_msel_pri_out_reg[0]  <= n7534;
    s11_next_reg <= n7539;
    s2_next_reg <= n7544;
    s4_next_reg <= n7549;
    s7_next_reg <= n7554;
    \\s11_msel_pri_out_reg[1]  <= n7559;
    \\s12_msel_pri_out_reg[1]  <= n7564;
    \\s13_msel_pri_out_reg[1]  <= n7569;
    \\s3_msel_pri_out_reg[1]  <= n7574;
    \\s5_msel_pri_out_reg[1]  <= n7579;
    \\s6_msel_pri_out_reg[1]  <= n7584;
    s5_next_reg <= n7589;
    \\s14_msel_pri_out_reg[0]  <= n7594;
    \\s4_msel_pri_out_reg[0]  <= n7599;
    \\s15_msel_pri_out_reg[1]  <= n7604;
    \\s10_msel_pri_out_reg[0]  <= n7609;
    \\s2_msel_pri_out_reg[1]  <= n7614;
    \\s1_msel_pri_out_reg[1]  <= n7619;
    \\s7_msel_pri_out_reg[1]  <= n7624;
    \\s0_msel_pri_out_reg[1]  <= n7629;
    \\s9_msel_pri_out_reg[1]  <= n7634;
    \\s4_msel_pri_out_reg[1]  <= n7639;
    \\s14_msel_pri_out_reg[1]  <= n7644;
    \\s10_msel_pri_out_reg[1]  <= n7649;
    s1_next_reg <= n7654;
    s10_next_reg <= n7659;
    m5_s0_cyc_o_reg <= n7664;
    m2_s0_cyc_o_reg <= n7669;
    m4_s0_cyc_o_reg <= n7674;
    m5_s1_cyc_o_reg <= n7679;
    m7_s0_cyc_o_reg <= n7684;
    m6_s0_cyc_o_reg <= n7689;
    m0_s0_cyc_o_reg <= n7694;
    m1_s0_cyc_o_reg <= n7699;
    m2_s1_cyc_o_reg <= n7704;
    m7_s1_cyc_o_reg <= n7709;
    m2_s15_cyc_o_reg <= n7714;
    m4_s15_cyc_o_reg <= n7719;
    m7_s12_cyc_o_reg <= n7724;
    m7_s8_cyc_o_reg <= n7729;
    m7_s4_cyc_o_reg <= n7734;
    m7_s15_cyc_o_reg <= n7739;
    m6_s15_cyc_o_reg <= n7744;
    m6_s1_cyc_o_reg <= n7749;
    m4_s1_cyc_o_reg <= n7754;
    m1_s1_cyc_o_reg <= n7759;
    m3_s0_cyc_o_reg <= n7764;
    m0_s1_cyc_o_reg <= n7769;
    m0_s13_cyc_o_reg <= n7774;
    m0_s15_cyc_o_reg <= n7779;
    m0_s7_cyc_o_reg <= n7784;
    m4_s6_cyc_o_reg <= n7789;
    m5_s5_cyc_o_reg <= n7794;
    m4_s4_cyc_o_reg <= n7799;
    m4_s5_cyc_o_reg <= n7804;
    m7_s7_cyc_o_reg <= n7809;
    m4_s7_cyc_o_reg <= n7814;
    m2_s5_cyc_o_reg <= n7819;
    m3_s15_cyc_o_reg <= n7824;
    m3_s1_cyc_o_reg <= n7829;
    m0_s2_cyc_o_reg <= n7834;
    m0_s6_cyc_o_reg <= n7839;
    m1_s15_cyc_o_reg <= n7844;
    m1_s4_cyc_o_reg <= n7849;
    m1_s8_cyc_o_reg <= n7854;
    m2_s10_cyc_o_reg <= n7859;
    m4_s10_cyc_o_reg <= n7864;
    m4_s12_cyc_o_reg <= n7869;
    m4_s8_cyc_o_reg <= n7874;
    m5_s10_cyc_o_reg <= n7879;
    m5_s12_cyc_o_reg <= n7884;
    m5_s15_cyc_o_reg <= n7889;
    m5_s8_cyc_o_reg <= n7894;
    m6_s12_cyc_o_reg <= n7899;
    m6_s4_cyc_o_reg <= n7904;
    m7_s11_cyc_o_reg <= n7909;
    m7_s5_cyc_o_reg <= n7914;
    m6_s14_cyc_o_reg <= n7919;
    m7_s6_cyc_o_reg <= n7924;
    m6_s8_cyc_o_reg <= n7929;
    m6_s9_cyc_o_reg <= n7934;
    m6_s5_cyc_o_reg <= n7939;
    m5_s4_cyc_o_reg <= n7944;
    m6_s13_cyc_o_reg <= n7949;
    m5_s6_cyc_o_reg <= n7954;
    m4_s9_cyc_o_reg <= n7959;
    m4_s13_cyc_o_reg <= n7964;
    m4_s14_cyc_o_reg <= n7969;
    m3_s9_cyc_o_reg <= n7974;
    m3_s8_cyc_o_reg <= n7979;
    m3_s10_cyc_o_reg <= n7984;
    m2_s6_cyc_o_reg <= n7989;
    m2_s9_cyc_o_reg <= n7994;
    m1_s6_cyc_o_reg <= n7999;
    m0_s8_cyc_o_reg <= n8004;
    m1_s5_cyc_o_reg <= n8009;
    m0_s9_cyc_o_reg <= n8014;
    m1_s12_cyc_o_reg <= n8019;
    m1_s10_cyc_o_reg <= n8024;
    m0_s3_cyc_o_reg <= n8029;
    m0_s5_cyc_o_reg <= n8034;
    m0_s12_cyc_o_reg <= n8039;
    m0_s11_cyc_o_reg <= n8044;
    m0_s10_cyc_o_reg <= n8049;
    m7_s3_cyc_o_reg <= n8054;
    m1_s13_cyc_o_reg <= n8059;
    m2_s11_cyc_o_reg <= n8064;
    m3_s11_cyc_o_reg <= n8069;
    m3_s13_cyc_o_reg <= n8074;
    m3_s4_cyc_o_reg <= n8079;
    m5_s2_cyc_o_reg <= n8084;
    m6_s2_cyc_o_reg <= n8089;
    m7_s9_cyc_o_reg <= n8094;
    m7_s13_cyc_o_reg <= n8099;
    m7_s2_cyc_o_reg <= n8104;
    m7_s14_cyc_o_reg <= n8109;
    m7_s10_cyc_o_reg <= n8114;
    m6_s7_cyc_o_reg <= n8119;
    m6_s6_cyc_o_reg <= n8124;
    m6_s11_cyc_o_reg <= n8129;
    m5_s9_cyc_o_reg <= n8134;
    m6_s10_cyc_o_reg <= n8139;
    m5_s7_cyc_o_reg <= n8144;
    m5_s14_cyc_o_reg <= n8149;
    m5_s3_cyc_o_reg <= n8154;
    m5_s13_cyc_o_reg <= n8159;
    m5_s11_cyc_o_reg <= n8164;
    m4_s11_cyc_o_reg <= n8169;
    m4_s2_cyc_o_reg <= n8174;
    m2_s4_cyc_o_reg <= n8179;
    m3_s5_cyc_o_reg <= n8184;
    m3_s6_cyc_o_reg <= n8189;
    m3_s7_cyc_o_reg <= n8194;
    m3_s3_cyc_o_reg <= n8199;
    m3_s14_cyc_o_reg <= n8204;
    m3_s12_cyc_o_reg <= n8209;
    m2_s8_cyc_o_reg <= n8214;
    m2_s7_cyc_o_reg <= n8219;
    m2_s13_cyc_o_reg <= n8224;
    m2_s14_cyc_o_reg <= n8229;
    m2_s2_cyc_o_reg <= n8234;
    m1_s7_cyc_o_reg <= n8239;
    m1_s9_cyc_o_reg <= n8244;
    m1_s2_cyc_o_reg <= n8249;
    m1_s14_cyc_o_reg <= n8254;
    m1_s11_cyc_o_reg <= n8259;
    m3_s2_cyc_o_reg <= n8264;
    m0_s14_cyc_o_reg <= n8269;
    m0_s4_cyc_o_reg <= n8274;
    m4_s3_cyc_o_reg <= n8279;
    m6_s3_cyc_o_reg <= n8284;
    m2_s3_cyc_o_reg <= n8289;
    m2_s12_cyc_o_reg <= n8294;
    m1_s3_cyc_o_reg <= n8299;
    s6_m4_cyc_r_reg <= n8304;
    s15_m6_cyc_r_reg <= n8309;
    s8_m2_cyc_r_reg <= n8314;
    s5_m5_cyc_r_reg <= n8319;
    s13_m5_cyc_r_reg <= n8324;
    s3_m5_cyc_r_reg <= n8329;
    s1_m1_cyc_r_reg <= n8334;
    s11_m5_cyc_r_reg <= n8339;
    s12_m5_cyc_r_reg <= n8344;
    s15_m1_cyc_r_reg <= n8349;
    s15_m3_cyc_r_reg <= n8354;
    s10_m4_cyc_r_reg <= n8359;
    s6_m5_cyc_r_reg <= n8364;
    s8_m5_cyc_r_reg <= n8369;
    s10_m5_cyc_r_reg <= n8374;
    s5_m2_cyc_r_reg <= n8379;
    s8_m1_cyc_r_reg <= n8384;
    s4_m0_cyc_r_reg <= n8389;
    s7_m1_cyc_r_reg <= n8394;
    s5_m4_cyc_r_reg <= n8399;
    s15_m2_cyc_r_reg <= n8404;
    s10_m3_cyc_r_reg <= n8409;
    s0_m0_cyc_r_reg <= n8414;
    s5_m7_cyc_r_reg <= n8419;
    s7_m7_cyc_r_reg <= n8424;
    s11_m4_cyc_r_reg <= n8429;
    s14_m5_cyc_r_reg <= n8434;
    s15_m0_cyc_r_reg <= n8439;
    s9_m7_cyc_r_reg <= n8444;
    s0_m4_cyc_r_reg <= n8449;
    s13_m4_cyc_r_reg <= n8454;
    s2_m3_cyc_r_reg <= n8459;
    s11_m1_cyc_r_reg <= n8464;
    s13_m2_cyc_r_reg <= n8469;
    s0_m2_cyc_r_reg <= n8474;
    s9_m4_cyc_r_reg <= n8479;
    s4_m7_cyc_r_reg <= n8484;
    s13_m7_cyc_r_reg <= n8489;
    s8_m0_cyc_r_reg <= n8494;
    s7_m2_cyc_r_reg <= n8499;
    s7_m3_cyc_r_reg <= n8504;
    s3_m1_cyc_r_reg <= n8509;
    s9_m0_cyc_r_reg <= n8514;
    s10_m1_cyc_r_reg <= n8519;
    s6_m7_cyc_r_reg <= n8524;
    s11_m2_cyc_r_reg <= n8529;
    s13_m3_cyc_r_reg <= n8534;
    s10_m2_cyc_r_reg <= n8539;
    s12_m3_cyc_r_reg <= n8544;
    s14_m6_cyc_r_reg <= n8549;
    s15_m7_cyc_r_reg <= n8554;
    s10_m0_cyc_r_reg <= n8559;
    s11_m3_cyc_r_reg <= n8564;
    s4_m2_cyc_r_reg <= n8569;
    s7_m6_cyc_r_reg <= n8574;
    s9_m3_cyc_r_reg <= n8579;
    s4_m6_cyc_r_reg <= n8584;
    s0_m1_cyc_r_reg <= n8589;
    s1_m2_cyc_r_reg <= n8594;
    s10_m7_cyc_r_reg <= n8599;
    s11_m6_cyc_r_reg <= n8604;
    s4_m4_cyc_r_reg <= n8609;
    s9_m2_cyc_r_reg <= n8614;
    s1_m5_cyc_r_reg <= n8619;
    s14_m3_cyc_r_reg <= n8624;
    s12_m2_cyc_r_reg <= n8629;
    s9_m1_cyc_r_reg <= n8634;
    s3_m6_cyc_r_reg <= n8639;
    s2_m6_cyc_r_reg <= n8644;
    s6_m3_cyc_r_reg <= n8649;
    s6_m6_cyc_r_reg <= n8654;
    s8_m6_cyc_r_reg <= n8659;
    s1_m4_cyc_r_reg <= n8664;
    s6_m0_cyc_r_reg <= n8669;
    s2_m7_cyc_r_reg <= n8674;
    s3_m3_cyc_r_reg <= n8679;
    s12_m0_cyc_r_reg <= n8684;
    s1_m7_cyc_r_reg <= n8689;
    s8_m7_cyc_r_reg <= n8694;
    s2_m0_cyc_r_reg <= n8699;
    s1_m3_cyc_r_reg <= n8704;
    s1_m0_cyc_r_reg <= n8709;
    s3_m2_cyc_r_reg <= n8714;
    s13_m6_cyc_r_reg <= n8719;
    s2_m1_cyc_r_reg <= n8724;
    s3_m0_cyc_r_reg <= n8729;
    s2_m5_cyc_r_reg <= n8734;
    s2_m4_cyc_r_reg <= n8739;
    s5_m6_cyc_r_reg <= n8744;
    s14_m4_cyc_r_reg <= n8749;
    s14_m0_cyc_r_reg <= n8754;
    s15_m4_cyc_r_reg <= n8759;
    s3_m4_cyc_r_reg <= n8764;
    s2_m2_cyc_r_reg <= n8769;
    s5_m3_cyc_r_reg <= n8774;
    s12_m1_cyc_r_reg <= n8779;
    s5_m0_cyc_r_reg <= n8784;
    s0_m7_cyc_r_reg <= n8789;
    s13_m0_cyc_r_reg <= n8794;
    s1_m6_cyc_r_reg <= n8799;
    s0_m5_cyc_r_reg <= n8804;
    s15_m5_cyc_r_reg <= n8809;
    s3_m7_cyc_r_reg <= n8814;
    s9_m6_cyc_r_reg <= n8819;
    s14_m2_cyc_r_reg <= n8824;
    s4_m3_cyc_r_reg <= n8829;
    s6_m2_cyc_r_reg <= n8834;
    s7_m5_cyc_r_reg <= n8839;
    s13_m1_cyc_r_reg <= n8844;
    s0_m6_cyc_r_reg <= n8849;
    s10_m6_cyc_r_reg <= n8854;
    s8_m4_cyc_r_reg <= n8859;
    s0_m3_cyc_r_reg <= n8864;
    s4_m5_cyc_r_reg <= n8869;
    s5_m1_cyc_r_reg <= n8874;
    s6_m1_cyc_r_reg <= n8879;
    s4_m1_cyc_r_reg <= n8884;
    s14_m1_cyc_r_reg <= n8889;
    s14_m7_cyc_r_reg <= n8894;
    s12_m4_cyc_r_reg <= n8899;
    s7_m0_cyc_r_reg <= n8904;
    s12_m7_cyc_r_reg <= n8909;
    s7_m4_cyc_r_reg <= n8914;
    s8_m3_cyc_r_reg <= n8919;
    s9_m5_cyc_r_reg <= n8924;
    s11_m0_cyc_r_reg <= n8929;
    s11_m7_cyc_r_reg <= n8934;
    s12_m6_cyc_r_reg <= n8939;
  end
  initial begin
    \\rf_conf15_reg[0]  <= 1'b0;
    \\rf_conf15_reg[10]  <= 1'b0;
    \\rf_conf15_reg[11]  <= 1'b0;
    \\rf_conf15_reg[12]  <= 1'b0;
    \\rf_conf15_reg[13]  <= 1'b0;
    \\rf_conf15_reg[14]  <= 1'b0;
    \\rf_conf15_reg[15]  <= 1'b0;
    \\rf_conf15_reg[1]  <= 1'b0;
    \\rf_conf15_reg[2]  <= 1'b0;
    \\rf_conf15_reg[3]  <= 1'b0;
    \\rf_conf15_reg[4]  <= 1'b0;
    \\rf_conf15_reg[5]  <= 1'b0;
    \\rf_conf15_reg[6]  <= 1'b0;
    \\rf_conf15_reg[7]  <= 1'b0;
    \\rf_conf15_reg[8]  <= 1'b0;
    \\rf_conf15_reg[9]  <= 1'b0;
    \\rf_conf0_reg[0]  <= 1'b0;
    \\rf_conf0_reg[10]  <= 1'b0;
    \\rf_conf0_reg[11]  <= 1'b0;
    \\rf_conf0_reg[12]  <= 1'b0;
    \\rf_conf0_reg[13]  <= 1'b0;
    \\rf_conf0_reg[14]  <= 1'b0;
    \\rf_conf0_reg[15]  <= 1'b0;
    \\rf_conf0_reg[1]  <= 1'b0;
    \\rf_conf0_reg[2]  <= 1'b0;
    \\rf_conf0_reg[3]  <= 1'b0;
    \\rf_conf0_reg[4]  <= 1'b0;
    \\rf_conf0_reg[5]  <= 1'b0;
    \\rf_conf0_reg[6]  <= 1'b0;
    \\rf_conf0_reg[7]  <= 1'b0;
    \\rf_conf0_reg[8]  <= 1'b0;
    \\rf_conf0_reg[9]  <= 1'b0;
    \\rf_conf12_reg[0]  <= 1'b0;
    \\rf_conf12_reg[10]  <= 1'b0;
    \\rf_conf12_reg[11]  <= 1'b0;
    \\rf_conf12_reg[12]  <= 1'b0;
    \\rf_conf12_reg[13]  <= 1'b0;
    \\rf_conf12_reg[14]  <= 1'b0;
    \\rf_conf12_reg[15]  <= 1'b0;
    \\rf_conf12_reg[1]  <= 1'b0;
    \\rf_conf12_reg[2]  <= 1'b0;
    \\rf_conf12_reg[3]  <= 1'b0;
    \\rf_conf12_reg[4]  <= 1'b0;
    \\rf_conf12_reg[5]  <= 1'b0;
    \\rf_conf12_reg[6]  <= 1'b0;
    \\rf_conf12_reg[7]  <= 1'b0;
    \\rf_conf12_reg[8]  <= 1'b0;
    \\rf_conf12_reg[9]  <= 1'b0;
    \\rf_conf13_reg[0]  <= 1'b0;
    \\rf_conf13_reg[10]  <= 1'b0;
    \\rf_conf13_reg[11]  <= 1'b0;
    \\rf_conf13_reg[12]  <= 1'b0;
    \\rf_conf13_reg[13]  <= 1'b0;
    \\rf_conf13_reg[14]  <= 1'b0;
    \\rf_conf13_reg[15]  <= 1'b0;
    \\rf_conf13_reg[1]  <= 1'b0;
    \\rf_conf13_reg[4]  <= 1'b0;
    \\rf_conf13_reg[5]  <= 1'b0;
    \\rf_conf13_reg[6]  <= 1'b0;
    \\rf_conf13_reg[7]  <= 1'b0;
    \\rf_conf13_reg[8]  <= 1'b0;
    \\rf_conf13_reg[9]  <= 1'b0;
    \\rf_conf14_reg[0]  <= 1'b0;
    \\rf_conf14_reg[10]  <= 1'b0;
    \\rf_conf14_reg[11]  <= 1'b0;
    \\rf_conf14_reg[12]  <= 1'b0;
    \\rf_conf14_reg[13]  <= 1'b0;
    \\rf_conf14_reg[14]  <= 1'b0;
    \\rf_conf14_reg[15]  <= 1'b0;
    \\rf_conf14_reg[1]  <= 1'b0;
    \\rf_conf14_reg[3]  <= 1'b0;
    \\rf_conf14_reg[4]  <= 1'b0;
    \\rf_conf14_reg[5]  <= 1'b0;
    \\rf_conf14_reg[6]  <= 1'b0;
    \\rf_conf14_reg[7]  <= 1'b0;
    \\rf_conf14_reg[8]  <= 1'b0;
    \\rf_conf14_reg[9]  <= 1'b0;
    \\rf_conf13_reg[2]  <= 1'b0;
    \\rf_conf13_reg[3]  <= 1'b0;
    \\rf_conf14_reg[2]  <= 1'b0;
    \\rf_conf1_reg[0]  <= 1'b0;
    \\rf_conf1_reg[10]  <= 1'b0;
    \\rf_conf1_reg[11]  <= 1'b0;
    \\rf_conf1_reg[12]  <= 1'b0;
    \\rf_conf1_reg[13]  <= 1'b0;
    \\rf_conf1_reg[14]  <= 1'b0;
    \\rf_conf1_reg[15]  <= 1'b0;
    \\rf_conf1_reg[1]  <= 1'b0;
    \\rf_conf1_reg[2]  <= 1'b0;
    \\rf_conf1_reg[3]  <= 1'b0;
    \\rf_conf1_reg[4]  <= 1'b0;
    \\rf_conf1_reg[5]  <= 1'b0;
    \\rf_conf1_reg[6]  <= 1'b0;
    \\rf_conf1_reg[7]  <= 1'b0;
    \\rf_conf1_reg[8]  <= 1'b0;
    \\rf_conf1_reg[9]  <= 1'b0;
    \\rf_conf2_reg[0]  <= 1'b0;
    \\rf_conf2_reg[10]  <= 1'b0;
    \\rf_conf2_reg[11]  <= 1'b0;
    \\rf_conf2_reg[12]  <= 1'b0;
    \\rf_conf2_reg[13]  <= 1'b0;
    \\rf_conf2_reg[14]  <= 1'b0;
    \\rf_conf2_reg[15]  <= 1'b0;
    \\rf_conf2_reg[1]  <= 1'b0;
    \\rf_conf2_reg[2]  <= 1'b0;
    \\rf_conf2_reg[3]  <= 1'b0;
    \\rf_conf2_reg[4]  <= 1'b0;
    \\rf_conf2_reg[5]  <= 1'b0;
    \\rf_conf2_reg[6]  <= 1'b0;
    \\rf_conf2_reg[7]  <= 1'b0;
    \\rf_conf2_reg[8]  <= 1'b0;
    \\rf_conf2_reg[9]  <= 1'b0;
    \\rf_conf3_reg[0]  <= 1'b0;
    \\rf_conf3_reg[10]  <= 1'b0;
    \\rf_conf3_reg[11]  <= 1'b0;
    \\rf_conf3_reg[12]  <= 1'b0;
    \\rf_conf3_reg[13]  <= 1'b0;
    \\rf_conf3_reg[14]  <= 1'b0;
    \\rf_conf3_reg[15]  <= 1'b0;
    \\rf_conf3_reg[1]  <= 1'b0;
    \\rf_conf3_reg[2]  <= 1'b0;
    \\rf_conf3_reg[3]  <= 1'b0;
    \\rf_conf3_reg[4]  <= 1'b0;
    \\rf_conf3_reg[5]  <= 1'b0;
    \\rf_conf3_reg[6]  <= 1'b0;
    \\rf_conf3_reg[7]  <= 1'b0;
    \\rf_conf3_reg[8]  <= 1'b0;
    \\rf_conf3_reg[9]  <= 1'b0;
    \\rf_conf5_reg[0]  <= 1'b0;
    \\rf_conf5_reg[10]  <= 1'b0;
    \\rf_conf5_reg[11]  <= 1'b0;
    \\rf_conf5_reg[12]  <= 1'b0;
    \\rf_conf5_reg[13]  <= 1'b0;
    \\rf_conf5_reg[14]  <= 1'b0;
    \\rf_conf5_reg[15]  <= 1'b0;
    \\rf_conf5_reg[1]  <= 1'b0;
    \\rf_conf5_reg[2]  <= 1'b0;
    \\rf_conf5_reg[3]  <= 1'b0;
    \\rf_conf5_reg[4]  <= 1'b0;
    \\rf_conf5_reg[5]  <= 1'b0;
    \\rf_conf5_reg[6]  <= 1'b0;
    \\rf_conf5_reg[7]  <= 1'b0;
    \\rf_conf5_reg[8]  <= 1'b0;
    \\rf_conf5_reg[9]  <= 1'b0;
    \\rf_conf7_reg[0]  <= 1'b0;
    \\rf_conf7_reg[10]  <= 1'b0;
    \\rf_conf7_reg[11]  <= 1'b0;
    \\rf_conf7_reg[12]  <= 1'b0;
    \\rf_conf7_reg[13]  <= 1'b0;
    \\rf_conf7_reg[14]  <= 1'b0;
    \\rf_conf7_reg[15]  <= 1'b0;
    \\rf_conf7_reg[1]  <= 1'b0;
    \\rf_conf7_reg[2]  <= 1'b0;
    \\rf_conf7_reg[3]  <= 1'b0;
    \\rf_conf7_reg[4]  <= 1'b0;
    \\rf_conf7_reg[5]  <= 1'b0;
    \\rf_conf7_reg[6]  <= 1'b0;
    \\rf_conf7_reg[7]  <= 1'b0;
    \\rf_conf7_reg[8]  <= 1'b0;
    \\rf_conf7_reg[9]  <= 1'b0;
    \\rf_conf10_reg[0]  <= 1'b0;
    \\rf_conf10_reg[10]  <= 1'b0;
    \\rf_conf10_reg[11]  <= 1'b0;
    \\rf_conf10_reg[12]  <= 1'b0;
    \\rf_conf10_reg[13]  <= 1'b0;
    \\rf_conf10_reg[14]  <= 1'b0;
    \\rf_conf10_reg[15]  <= 1'b0;
    \\rf_conf10_reg[1]  <= 1'b0;
    \\rf_conf10_reg[2]  <= 1'b0;
    \\rf_conf10_reg[3]  <= 1'b0;
    \\rf_conf10_reg[4]  <= 1'b0;
    \\rf_conf10_reg[5]  <= 1'b0;
    \\rf_conf10_reg[6]  <= 1'b0;
    \\rf_conf10_reg[7]  <= 1'b0;
    \\rf_conf10_reg[8]  <= 1'b0;
    \\rf_conf10_reg[9]  <= 1'b0;
    \\rf_conf11_reg[0]  <= 1'b0;
    \\rf_conf11_reg[10]  <= 1'b0;
    \\rf_conf11_reg[11]  <= 1'b0;
    \\rf_conf11_reg[12]  <= 1'b0;
    \\rf_conf11_reg[13]  <= 1'b0;
    \\rf_conf11_reg[14]  <= 1'b0;
    \\rf_conf11_reg[15]  <= 1'b0;
    \\rf_conf11_reg[1]  <= 1'b0;
    \\rf_conf11_reg[4]  <= 1'b0;
    \\rf_conf11_reg[5]  <= 1'b0;
    \\rf_conf11_reg[6]  <= 1'b0;
    \\rf_conf11_reg[7]  <= 1'b0;
    \\rf_conf11_reg[8]  <= 1'b0;
    \\rf_conf11_reg[9]  <= 1'b0;
    \\rf_conf11_reg[2]  <= 1'b0;
    \\rf_conf11_reg[3]  <= 1'b0;
    \\rf_conf4_reg[0]  <= 1'b0;
    \\rf_conf4_reg[10]  <= 1'b0;
    \\rf_conf4_reg[11]  <= 1'b0;
    \\rf_conf4_reg[12]  <= 1'b0;
    \\rf_conf4_reg[13]  <= 1'b0;
    \\rf_conf4_reg[14]  <= 1'b0;
    \\rf_conf4_reg[15]  <= 1'b0;
    \\rf_conf4_reg[1]  <= 1'b0;
    \\rf_conf4_reg[4]  <= 1'b0;
    \\rf_conf4_reg[5]  <= 1'b0;
    \\rf_conf4_reg[6]  <= 1'b0;
    \\rf_conf4_reg[7]  <= 1'b0;
    \\rf_conf4_reg[8]  <= 1'b0;
    \\rf_conf4_reg[9]  <= 1'b0;
    \\rf_conf4_reg[2]  <= 1'b0;
    \\rf_conf4_reg[3]  <= 1'b0;
    \\rf_conf6_reg[0]  <= 1'b0;
    \\rf_conf6_reg[10]  <= 1'b0;
    \\rf_conf6_reg[11]  <= 1'b0;
    \\rf_conf6_reg[12]  <= 1'b0;
    \\rf_conf6_reg[13]  <= 1'b0;
    \\rf_conf6_reg[14]  <= 1'b0;
    \\rf_conf6_reg[15]  <= 1'b0;
    \\rf_conf6_reg[1]  <= 1'b0;
    \\rf_conf6_reg[4]  <= 1'b0;
    \\rf_conf6_reg[5]  <= 1'b0;
    \\rf_conf6_reg[6]  <= 1'b0;
    \\rf_conf6_reg[7]  <= 1'b0;
    \\rf_conf6_reg[8]  <= 1'b0;
    \\rf_conf6_reg[9]  <= 1'b0;
    \\rf_conf6_reg[2]  <= 1'b0;
    \\rf_conf6_reg[3]  <= 1'b0;
    \\rf_conf9_reg[0]  <= 1'b0;
    \\rf_conf9_reg[10]  <= 1'b0;
    \\rf_conf9_reg[11]  <= 1'b0;
    \\rf_conf9_reg[12]  <= 1'b0;
    \\rf_conf9_reg[13]  <= 1'b0;
    \\rf_conf9_reg[14]  <= 1'b0;
    \\rf_conf9_reg[15]  <= 1'b0;
    \\rf_conf9_reg[1]  <= 1'b0;
    \\rf_conf9_reg[2]  <= 1'b0;
    \\rf_conf9_reg[3]  <= 1'b0;
    \\rf_conf9_reg[4]  <= 1'b0;
    \\rf_conf9_reg[5]  <= 1'b0;
    \\rf_conf9_reg[6]  <= 1'b0;
    \\rf_conf9_reg[7]  <= 1'b0;
    \\rf_conf9_reg[8]  <= 1'b0;
    \\rf_conf9_reg[9]  <= 1'b0;
    \\rf_conf8_reg[0]  <= 1'b0;
    \\rf_conf8_reg[10]  <= 1'b0;
    \\rf_conf8_reg[11]  <= 1'b0;
    \\rf_conf8_reg[12]  <= 1'b0;
    \\rf_conf8_reg[13]  <= 1'b0;
    \\rf_conf8_reg[14]  <= 1'b0;
    \\rf_conf8_reg[15]  <= 1'b0;
    \\rf_conf8_reg[1]  <= 1'b0;
    \\rf_conf8_reg[4]  <= 1'b0;
    \\rf_conf8_reg[5]  <= 1'b0;
    \\rf_conf8_reg[6]  <= 1'b0;
    \\rf_conf8_reg[7]  <= 1'b0;
    \\rf_conf8_reg[8]  <= 1'b0;
    \\rf_conf8_reg[9]  <= 1'b0;
    \\rf_conf8_reg[2]  <= 1'b0;
    \\rf_conf8_reg[3]  <= 1'b0;
    \\s14_msel_arb2_state_reg[0]  <= 1'b0;
    \\s10_msel_arb0_state_reg[1]  <= 1'b0;
    \\s11_msel_arb0_state_reg[1]  <= 1'b0;
    \\s12_msel_arb0_state_reg[1]  <= 1'b0;
    \\s13_msel_arb0_state_reg[1]  <= 1'b0;
    \\s14_msel_arb0_state_reg[1]  <= 1'b0;
    \\s15_msel_arb0_state_reg[1]  <= 1'b0;
    \\s1_msel_arb0_state_reg[1]  <= 1'b0;
    \\s2_msel_arb0_state_reg[1]  <= 1'b0;
    \\s3_msel_arb0_state_reg[1]  <= 1'b0;
    \\s4_msel_arb0_state_reg[1]  <= 1'b0;
    \\s5_msel_arb0_state_reg[1]  <= 1'b0;
    \\s6_msel_arb0_state_reg[1]  <= 1'b0;
    \\s8_msel_arb0_state_reg[1]  <= 1'b0;
    \\s9_msel_arb0_state_reg[1]  <= 1'b0;
    \\s0_msel_arb0_state_reg[1]  <= 1'b0;
    \\s11_msel_arb0_state_reg[0]  <= 1'b0;
    \\s11_msel_arb1_state_reg[1]  <= 1'b0;
    \\s12_msel_arb0_state_reg[0]  <= 1'b0;
    \\s13_msel_arb0_state_reg[0]  <= 1'b0;
    \\s13_msel_arb2_state_reg[0]  <= 1'b0;
    \\s14_msel_arb0_state_reg[0]  <= 1'b0;
    \\s15_msel_arb2_state_reg[0]  <= 1'b0;
    \\s15_msel_arb3_state_reg[1]  <= 1'b0;
    \\s3_msel_arb0_state_reg[0]  <= 1'b0;
    \\s4_msel_arb0_state_reg[0]  <= 1'b0;
    \\s4_msel_arb2_state_reg[0]  <= 1'b0;
    \\s4_msel_arb2_state_reg[1]  <= 1'b0;
    \\s5_msel_arb0_state_reg[0]  <= 1'b0;
    \\s5_msel_arb3_state_reg[1]  <= 1'b0;
    \\s6_msel_arb0_state_reg[0]  <= 1'b0;
    \\s6_msel_arb1_state_reg[0]  <= 1'b0;
    \\s6_msel_arb1_state_reg[1]  <= 1'b0;
    \\s7_msel_arb0_state_reg[0]  <= 1'b0;
    \\s8_msel_arb0_state_reg[0]  <= 1'b0;
    \\s8_msel_arb1_state_reg[1]  <= 1'b0;
    \\s8_msel_arb3_state_reg[1]  <= 1'b0;
    \\s9_msel_arb3_state_reg[0]  <= 1'b0;
    \\s9_msel_arb2_state_reg[0]  <= 1'b0;
    \\s0_msel_arb2_state_reg[0]  <= 1'b0;
    \\s7_msel_arb0_state_reg[1]  <= 1'b0;
    \\s10_msel_arb2_state_reg[1]  <= 1'b0;
    \\s10_msel_arb2_state_reg[0]  <= 1'b0;
    \\s11_msel_arb2_state_reg[1]  <= 1'b0;
    \\s11_msel_arb3_state_reg[1]  <= 1'b0;
    \\s12_msel_arb1_state_reg[1]  <= 1'b0;
    \\s12_msel_arb2_state_reg[0]  <= 1'b0;
    \\s12_msel_arb2_state_reg[1]  <= 1'b0;
    \\s13_msel_arb1_state_reg[1]  <= 1'b0;
    \\s13_msel_arb2_state_reg[1]  <= 1'b0;
    \\s14_msel_arb2_state_reg[1]  <= 1'b0;
    \\s14_msel_arb2_state_reg[2]  <= 1'b0;
    \\s15_msel_arb0_state_reg[0]  <= 1'b0;
    \\s15_msel_arb1_state_reg[1]  <= 1'b0;
    \\s15_msel_arb2_state_reg[1]  <= 1'b0;
    \\s15_msel_arb2_state_reg[2]  <= 1'b0;
    \\s1_msel_arb0_state_reg[0]  <= 1'b0;
    \\s1_msel_arb2_state_reg[0]  <= 1'b0;
    \\s1_msel_arb2_state_reg[1]  <= 1'b0;
    \\s2_msel_arb2_state_reg[0]  <= 1'b0;
    \\s2_msel_arb2_state_reg[1]  <= 1'b0;
    \\s2_msel_arb0_state_reg[0]  <= 1'b0;
    \\s3_msel_arb1_state_reg[1]  <= 1'b0;
    \\s3_msel_arb2_state_reg[0]  <= 1'b0;
    \\s3_msel_arb2_state_reg[1]  <= 1'b0;
    \\s3_msel_arb3_state_reg[1]  <= 1'b0;
    \\s4_msel_arb2_state_reg[2]  <= 1'b0;
    \\s5_msel_arb1_state_reg[1]  <= 1'b0;
    \\s5_msel_arb2_state_reg[1]  <= 1'b0;
    \\s5_msel_arb3_state_reg[0]  <= 1'b0;
    \\s5_msel_arb3_state_reg[2]  <= 1'b0;
    \\s6_msel_arb2_state_reg[1]  <= 1'b0;
    \\s6_msel_arb2_state_reg[0]  <= 1'b0;
    \\s6_msel_arb3_state_reg[1]  <= 1'b0;
    \\s6_msel_arb3_state_reg[0]  <= 1'b0;
    \\s7_msel_arb2_state_reg[0]  <= 1'b0;
    \\s7_msel_arb2_state_reg[1]  <= 1'b0;
    \\s8_msel_arb2_state_reg[0]  <= 1'b0;
    \\s8_msel_arb2_state_reg[1]  <= 1'b0;
    \\s8_msel_arb3_state_reg[0]  <= 1'b0;
    \\s9_msel_arb0_state_reg[0]  <= 1'b0;
    \\s9_msel_arb2_state_reg[2]  <= 1'b0;
    \\s0_msel_arb0_state_reg[0]  <= 1'b0;
    \\s0_msel_arb2_state_reg[1]  <= 1'b0;
    \\s0_msel_arb2_state_reg[2]  <= 1'b0;
    \\s0_msel_arb3_state_reg[0]  <= 1'b0;
    \\s14_msel_arb3_state_reg[0]  <= 1'b0;
    \\s12_msel_arb1_state_reg[0]  <= 1'b0;
    \\s10_msel_arb1_state_reg[0]  <= 1'b0;
    \\s10_msel_arb1_state_reg[1]  <= 1'b0;
    \\s10_msel_arb2_state_reg[2]  <= 1'b0;
    \\s11_msel_arb0_state_reg[2]  <= 1'b0;
    \\s11_msel_arb1_state_reg[2]  <= 1'b0;
    \\s11_msel_arb2_state_reg[0]  <= 1'b0;
    \\s11_msel_arb2_state_reg[2]  <= 1'b0;
    \\s11_msel_arb1_state_reg[0]  <= 1'b0;
    \\s11_msel_arb3_state_reg[2]  <= 1'b0;
    \\s12_msel_arb0_state_reg[2]  <= 1'b0;
    \\s12_msel_arb1_state_reg[2]  <= 1'b0;
    \\s12_msel_arb2_state_reg[2]  <= 1'b0;
    \\s13_msel_arb0_state_reg[2]  <= 1'b0;
    \\s12_msel_arb3_state_reg[1]  <= 1'b0;
    \\s13_msel_arb2_state_reg[2]  <= 1'b0;
    \\s13_msel_arb3_state_reg[1]  <= 1'b0;
    \\s14_msel_arb1_state_reg[2]  <= 1'b0;
    \\s14_msel_arb1_state_reg[1]  <= 1'b0;
    \\s14_msel_arb0_state_reg[2]  <= 1'b0;
    \\s14_msel_arb3_state_reg[1]  <= 1'b0;
    \\s14_msel_arb3_state_reg[2]  <= 1'b0;
    \\s15_msel_arb1_state_reg[0]  <= 1'b0;
    \\s15_msel_arb3_state_reg[0]  <= 1'b0;
    \\s1_msel_arb0_state_reg[2]  <= 1'b0;
    \\s1_msel_arb1_state_reg[1]  <= 1'b0;
    \\s1_msel_arb2_state_reg[2]  <= 1'b0;
    \\s1_msel_arb3_state_reg[0]  <= 1'b0;
    \\s1_msel_arb3_state_reg[1]  <= 1'b0;
    \\s2_msel_arb1_state_reg[1]  <= 1'b0;
    \\s2_msel_arb0_state_reg[2]  <= 1'b0;
    \\s2_msel_arb2_state_reg[2]  <= 1'b0;
    \\s2_msel_arb3_state_reg[0]  <= 1'b0;
    \\s2_msel_arb3_state_reg[1]  <= 1'b0;
    \\s3_msel_arb1_state_reg[0]  <= 1'b0;
    \\s3_msel_arb0_state_reg[2]  <= 1'b0;
    \\s3_msel_arb2_state_reg[2]  <= 1'b0;
    \\s4_msel_arb1_state_reg[0]  <= 1'b0;
    \\s4_msel_arb1_state_reg[1]  <= 1'b0;
    \\s4_msel_arb3_state_reg[0]  <= 1'b0;
    \\s5_msel_arb1_state_reg[0]  <= 1'b0;
    \\s5_msel_arb1_state_reg[2]  <= 1'b0;
    \\s5_msel_arb0_state_reg[2]  <= 1'b0;
    \\s6_msel_arb0_state_reg[2]  <= 1'b0;
    \\s6_msel_arb1_state_reg[2]  <= 1'b0;
    \\s6_msel_arb2_state_reg[2]  <= 1'b0;
    \\s7_msel_arb1_state_reg[0]  <= 1'b0;
    \\s7_msel_arb1_state_reg[2]  <= 1'b0;
    \\s7_msel_arb0_state_reg[2]  <= 1'b0;
    \\s7_msel_arb2_state_reg[2]  <= 1'b0;
    \\s7_msel_arb3_state_reg[2]  <= 1'b0;
    \\s8_msel_arb0_state_reg[2]  <= 1'b0;
    \\s8_msel_arb1_state_reg[0]  <= 1'b0;
    \\s7_msel_arb3_state_reg[1]  <= 1'b0;
    \\s8_msel_arb3_state_reg[2]  <= 1'b0;
    \\s9_msel_arb0_state_reg[2]  <= 1'b0;
    \\s9_msel_arb2_state_reg[1]  <= 1'b0;
    \\s9_msel_arb1_state_reg[2]  <= 1'b0;
    \\s9_msel_arb3_state_reg[1]  <= 1'b0;
    \\s0_msel_arb0_state_reg[2]  <= 1'b0;
    \\s0_msel_arb1_state_reg[1]  <= 1'b0;
    \\s0_msel_arb1_state_reg[2]  <= 1'b0;
    \\s10_msel_arb0_state_reg[0]  <= 1'b0;
    \\s0_msel_arb3_state_reg[2]  <= 1'b0;
    \\s13_msel_arb1_state_reg[0]  <= 1'b0;
    \\s10_msel_arb1_state_reg[2]  <= 1'b0;
    \\s11_msel_arb3_state_reg[0]  <= 1'b0;
    \\s9_msel_arb3_state_reg[2]  <= 1'b0;
    \\s9_msel_arb1_state_reg[0]  <= 1'b0;
    \\s8_msel_arb2_state_reg[2]  <= 1'b0;
    \\s8_msel_arb1_state_reg[2]  <= 1'b0;
    \\s5_msel_arb2_state_reg[2]  <= 1'b0;
    \\s5_msel_arb2_state_reg[0]  <= 1'b0;
    \\s4_msel_arb1_state_reg[2]  <= 1'b0;
    \\s4_msel_arb3_state_reg[1]  <= 1'b0;
    \\s4_msel_arb0_state_reg[2]  <= 1'b0;
    \\s3_msel_arb1_state_reg[2]  <= 1'b0;
    \\s1_msel_arb3_state_reg[2]  <= 1'b0;
    \\s1_msel_arb1_state_reg[0]  <= 1'b0;
    \\s1_msel_arb1_state_reg[2]  <= 1'b0;
    \\s13_msel_arb1_state_reg[2]  <= 1'b0;
    \\s13_msel_arb3_state_reg[2]  <= 1'b0;
    \\s10_msel_arb0_state_reg[2]  <= 1'b0;
    \\s10_msel_arb3_state_reg[2]  <= 1'b0;
    \\s12_msel_arb3_state_reg[0]  <= 1'b0;
    \\s12_msel_arb3_state_reg[2]  <= 1'b0;
    \\s13_msel_arb3_state_reg[0]  <= 1'b0;
    \\s14_msel_arb1_state_reg[0]  <= 1'b0;
    \\s15_msel_arb1_state_reg[2]  <= 1'b0;
    \\s15_msel_arb3_state_reg[2]  <= 1'b0;
    \\s2_msel_arb1_state_reg[0]  <= 1'b0;
    \\s2_msel_arb1_state_reg[2]  <= 1'b0;
    \\s3_msel_arb3_state_reg[0]  <= 1'b0;
    \\s3_msel_arb3_state_reg[2]  <= 1'b0;
    \\s4_msel_arb3_state_reg[2]  <= 1'b0;
    \\s9_msel_arb1_state_reg[1]  <= 1'b0;
    \\s0_msel_arb1_state_reg[0]  <= 1'b0;
    \\s0_msel_arb3_state_reg[1]  <= 1'b0;
    \\s10_msel_arb3_state_reg[1]  <= 1'b0;
    \\s10_msel_arb3_state_reg[0]  <= 1'b0;
    \\s6_msel_arb3_state_reg[2]  <= 1'b0;
    \\s7_msel_arb3_state_reg[0]  <= 1'b0;
    \\s7_msel_arb1_state_reg[1]  <= 1'b0;
    \\s15_msel_arb0_state_reg[2]  <= 1'b0;
    \\s2_msel_arb3_state_reg[2]  <= 1'b0;
    m5_s0_cyc_o_reg <= 1'b0;
    m2_s0_cyc_o_reg <= 1'b0;
    m4_s0_cyc_o_reg <= 1'b0;
    m5_s1_cyc_o_reg <= 1'b0;
    m7_s0_cyc_o_reg <= 1'b0;
    m6_s0_cyc_o_reg <= 1'b0;
    m0_s0_cyc_o_reg <= 1'b0;
    m1_s0_cyc_o_reg <= 1'b0;
    m2_s1_cyc_o_reg <= 1'b0;
    m7_s1_cyc_o_reg <= 1'b0;
    m2_s15_cyc_o_reg <= 1'b0;
    m4_s15_cyc_o_reg <= 1'b0;
    m7_s12_cyc_o_reg <= 1'b0;
    m7_s8_cyc_o_reg <= 1'b0;
    m7_s4_cyc_o_reg <= 1'b0;
    m7_s15_cyc_o_reg <= 1'b0;
    m6_s15_cyc_o_reg <= 1'b0;
    m6_s1_cyc_o_reg <= 1'b0;
    m4_s1_cyc_o_reg <= 1'b0;
    m1_s1_cyc_o_reg <= 1'b0;
    m3_s0_cyc_o_reg <= 1'b0;
    m0_s1_cyc_o_reg <= 1'b0;
    m0_s13_cyc_o_reg <= 1'b0;
    m0_s15_cyc_o_reg <= 1'b0;
    m0_s7_cyc_o_reg <= 1'b0;
    m4_s6_cyc_o_reg <= 1'b0;
    m5_s5_cyc_o_reg <= 1'b0;
    m4_s4_cyc_o_reg <= 1'b0;
    m4_s5_cyc_o_reg <= 1'b0;
    m7_s7_cyc_o_reg <= 1'b0;
    m4_s7_cyc_o_reg <= 1'b0;
    m2_s5_cyc_o_reg <= 1'b0;
    m3_s15_cyc_o_reg <= 1'b0;
    m3_s1_cyc_o_reg <= 1'b0;
    m0_s2_cyc_o_reg <= 1'b0;
    m0_s6_cyc_o_reg <= 1'b0;
    m1_s15_cyc_o_reg <= 1'b0;
    m1_s4_cyc_o_reg <= 1'b0;
    m1_s8_cyc_o_reg <= 1'b0;
    m2_s10_cyc_o_reg <= 1'b0;
    m4_s10_cyc_o_reg <= 1'b0;
    m4_s12_cyc_o_reg <= 1'b0;
    m4_s8_cyc_o_reg <= 1'b0;
    m5_s10_cyc_o_reg <= 1'b0;
    m5_s12_cyc_o_reg <= 1'b0;
    m5_s15_cyc_o_reg <= 1'b0;
    m5_s8_cyc_o_reg <= 1'b0;
    m6_s12_cyc_o_reg <= 1'b0;
    m6_s4_cyc_o_reg <= 1'b0;
    m7_s11_cyc_o_reg <= 1'b0;
    m7_s5_cyc_o_reg <= 1'b0;
    m6_s14_cyc_o_reg <= 1'b0;
    m7_s6_cyc_o_reg <= 1'b0;
    m6_s8_cyc_o_reg <= 1'b0;
    m6_s9_cyc_o_reg <= 1'b0;
    m6_s5_cyc_o_reg <= 1'b0;
    m5_s4_cyc_o_reg <= 1'b0;
    m6_s13_cyc_o_reg <= 1'b0;
    m5_s6_cyc_o_reg <= 1'b0;
    m4_s9_cyc_o_reg <= 1'b0;
    m4_s13_cyc_o_reg <= 1'b0;
    m4_s14_cyc_o_reg <= 1'b0;
    m3_s9_cyc_o_reg <= 1'b0;
    m3_s8_cyc_o_reg <= 1'b0;
    m3_s10_cyc_o_reg <= 1'b0;
    m2_s6_cyc_o_reg <= 1'b0;
    m2_s9_cyc_o_reg <= 1'b0;
    m1_s6_cyc_o_reg <= 1'b0;
    m0_s8_cyc_o_reg <= 1'b0;
    m1_s5_cyc_o_reg <= 1'b0;
    m0_s9_cyc_o_reg <= 1'b0;
    m1_s12_cyc_o_reg <= 1'b0;
    m1_s10_cyc_o_reg <= 1'b0;
    m0_s3_cyc_o_reg <= 1'b0;
    m0_s5_cyc_o_reg <= 1'b0;
    m0_s12_cyc_o_reg <= 1'b0;
    m0_s11_cyc_o_reg <= 1'b0;
    m0_s10_cyc_o_reg <= 1'b0;
    m7_s3_cyc_o_reg <= 1'b0;
    m1_s13_cyc_o_reg <= 1'b0;
    m2_s11_cyc_o_reg <= 1'b0;
    m3_s11_cyc_o_reg <= 1'b0;
    m3_s13_cyc_o_reg <= 1'b0;
    m3_s4_cyc_o_reg <= 1'b0;
    m5_s2_cyc_o_reg <= 1'b0;
    m6_s2_cyc_o_reg <= 1'b0;
    m7_s9_cyc_o_reg <= 1'b0;
    m7_s13_cyc_o_reg <= 1'b0;
    m7_s2_cyc_o_reg <= 1'b0;
    m7_s14_cyc_o_reg <= 1'b0;
    m7_s10_cyc_o_reg <= 1'b0;
    m6_s7_cyc_o_reg <= 1'b0;
    m6_s6_cyc_o_reg <= 1'b0;
    m6_s11_cyc_o_reg <= 1'b0;
    m5_s9_cyc_o_reg <= 1'b0;
    m6_s10_cyc_o_reg <= 1'b0;
    m5_s7_cyc_o_reg <= 1'b0;
    m5_s14_cyc_o_reg <= 1'b0;
    m5_s3_cyc_o_reg <= 1'b0;
    m5_s13_cyc_o_reg <= 1'b0;
    m5_s11_cyc_o_reg <= 1'b0;
    m4_s11_cyc_o_reg <= 1'b0;
    m4_s2_cyc_o_reg <= 1'b0;
    m2_s4_cyc_o_reg <= 1'b0;
    m3_s5_cyc_o_reg <= 1'b0;
    m3_s6_cyc_o_reg <= 1'b0;
    m3_s7_cyc_o_reg <= 1'b0;
    m3_s3_cyc_o_reg <= 1'b0;
    m3_s14_cyc_o_reg <= 1'b0;
    m3_s12_cyc_o_reg <= 1'b0;
    m2_s8_cyc_o_reg <= 1'b0;
    m2_s7_cyc_o_reg <= 1'b0;
    m2_s13_cyc_o_reg <= 1'b0;
    m2_s14_cyc_o_reg <= 1'b0;
    m2_s2_cyc_o_reg <= 1'b0;
    m1_s7_cyc_o_reg <= 1'b0;
    m1_s9_cyc_o_reg <= 1'b0;
    m1_s2_cyc_o_reg <= 1'b0;
    m1_s14_cyc_o_reg <= 1'b0;
    m1_s11_cyc_o_reg <= 1'b0;
    m3_s2_cyc_o_reg <= 1'b0;
    m0_s14_cyc_o_reg <= 1'b0;
    m0_s4_cyc_o_reg <= 1'b0;
    m4_s3_cyc_o_reg <= 1'b0;
    m6_s3_cyc_o_reg <= 1'b0;
    m2_s3_cyc_o_reg <= 1'b0;
    m2_s12_cyc_o_reg <= 1'b0;
    m1_s3_cyc_o_reg <= 1'b0;
  end
endmodule


