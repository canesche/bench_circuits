module top ( 
    pp, pq, pr, ps, pt, pu, pv, pw, px, py, pa, pb, pc, pe, pf, pg, ph, pi,
    pj, pk, pl, pm, pn, po,
    pa0, pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pz, pk0, pl0, pm0,
    pn0, po0, pp0, pq0, pr0, ps0, pt0  );
  input  pp, pq, pr, ps, pt, pu, pv, pw, px, py, pa, pb, pc, pe, pf, pg,
    ph, pi, pj, pk, pl, pm, pn, po;
  output pa0, pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pz, pk0, pl0, pm0,
    pn0, po0, pp0, pq0, pr0, ps0, pt0;
  wire new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n550_, new_n551_, new_n552_,
    new_n553_;
  assign new_n46_ = pq & pw;
  assign new_n47_ = pq & ~pv;
  assign new_n48_ = ~new_n46_ & ~new_n47_;
  assign new_n49_ = ~pv & ~py;
  assign new_n50_ = pw & new_n48_;
  assign new_n51_ = ~new_n49_ & new_n50_;
  assign new_n52_ = ps & ~pv;
  assign new_n53_ = ps & ~pf;
  assign new_n54_ = pt & ~pf;
  assign new_n55_ = ~pt & ~pu;
  assign new_n56_ = pt & new_n55_;
  assign new_n57_ = pt & ~pv;
  assign new_n58_ = ~pv & py;
  assign new_n59_ = pu & new_n58_;
  assign new_n60_ = ~pu & pv;
  assign new_n61_ = ~new_n59_ & ~new_n60_;
  assign new_n62_ = ~pf & new_n61_;
  assign new_n63_ = new_n55_ & new_n61_;
  assign new_n64_ = ps & new_n55_;
  assign new_n65_ = ~pv & new_n61_;
  assign new_n66_ = ~new_n64_ & ~new_n65_;
  assign new_n67_ = ~new_n62_ & ~new_n63_;
  assign new_n68_ = new_n66_ & new_n67_;
  assign new_n69_ = ~new_n56_ & ~new_n57_;
  assign new_n70_ = ~new_n52_ & ~new_n53_;
  assign new_n71_ = ~new_n54_ & new_n70_;
  assign new_n72_ = new_n69_ & new_n71_;
  assign new_n73_ = new_n68_ & new_n72_;
  assign new_n74_ = new_n48_ & new_n73_;
  assign new_n75_ = ~pu & new_n74_;
  assign new_n76_ = pt & new_n50_;
  assign new_n77_ = ~ps & new_n50_;
  assign new_n78_ = ~pu & new_n50_;
  assign new_n79_ = ~new_n49_ & new_n74_;
  assign new_n80_ = pt & new_n74_;
  assign new_n81_ = ~ps & new_n74_;
  assign new_n82_ = ~new_n51_ & ~new_n75_;
  assign new_n83_ = ~new_n76_ & ~new_n77_;
  assign new_n84_ = new_n82_ & new_n83_;
  assign new_n85_ = ~new_n80_ & ~new_n81_;
  assign new_n86_ = ~new_n78_ & ~new_n79_;
  assign new_n87_ = new_n85_ & new_n86_;
  assign pa0 = ~new_n84_ | ~new_n87_;
  assign new_n89_ = ~pt & py;
  assign new_n90_ = ~pv & new_n89_;
  assign new_n91_ = ~ps & new_n90_;
  assign new_n92_ = pv & ~pg;
  assign new_n93_ = ~pu & ~pv;
  assign new_n94_ = ~new_n91_ & ~new_n92_;
  assign new_n95_ = ~new_n55_ & ~new_n93_;
  assign new_n96_ = new_n94_ & new_n95_;
  assign new_n97_ = ~pt & ~py;
  assign new_n98_ = new_n52_ & new_n97_;
  assign new_n99_ = new_n96_ & new_n98_;
  assign new_n100_ = ~pw & new_n96_;
  assign pb0 = new_n99_ | new_n100_;
  assign new_n102_ = ~ps & new_n58_;
  assign new_n103_ = pq & new_n102_;
  assign new_n104_ = ~pt & new_n103_;
  assign new_n105_ = ~pw & new_n93_;
  assign new_n106_ = ~new_n104_ & ~new_n105_;
  assign new_n107_ = pw & new_n106_;
  assign new_n108_ = new_n98_ & new_n107_;
  assign new_n109_ = ~ps & new_n108_;
  assign new_n110_ = pt & new_n108_;
  assign new_n111_ = pt & new_n106_;
  assign new_n112_ = pw & new_n111_;
  assign new_n113_ = ~pq & new_n112_;
  assign new_n114_ = pu & new_n106_;
  assign new_n115_ = pw & new_n114_;
  assign new_n116_ = ~pq & new_n115_;
  assign new_n117_ = ~ps & new_n106_;
  assign new_n118_ = pw & new_n117_;
  assign new_n119_ = ~pq & new_n118_;
  assign new_n120_ = pt & pv;
  assign new_n121_ = pu & pv;
  assign new_n122_ = pt & ~pu;
  assign new_n123_ = ~new_n120_ & ~new_n121_;
  assign new_n124_ = ~new_n122_ & new_n123_;
  assign new_n125_ = new_n98_ & new_n106_;
  assign new_n126_ = new_n124_ & new_n125_;
  assign new_n127_ = pt & new_n126_;
  assign new_n128_ = ph & new_n125_;
  assign new_n129_ = pu & new_n128_;
  assign new_n130_ = ~ps & new_n126_;
  assign new_n131_ = ~pq & pw;
  assign new_n132_ = new_n106_ & new_n131_;
  assign new_n133_ = ph & new_n132_;
  assign new_n134_ = ~pq & new_n133_;
  assign new_n135_ = new_n124_ & new_n132_;
  assign new_n136_ = ~pq & new_n135_;
  assign new_n137_ = ~pw & new_n133_;
  assign new_n138_ = pu & new_n126_;
  assign new_n139_ = new_n98_ & new_n133_;
  assign new_n140_ = ~pw & new_n106_;
  assign new_n141_ = new_n124_ & new_n140_;
  assign new_n142_ = ~ps & new_n141_;
  assign new_n143_ = ph & new_n140_;
  assign new_n144_ = pt & new_n143_;
  assign new_n145_ = new_n114_ & new_n124_;
  assign new_n146_ = ~pq & new_n145_;
  assign new_n147_ = pu & new_n143_;
  assign new_n148_ = pu & new_n141_;
  assign new_n149_ = ~ps & new_n128_;
  assign new_n150_ = pt & new_n141_;
  assign new_n151_ = pt & new_n128_;
  assign new_n152_ = ~pw & new_n135_;
  assign new_n153_ = new_n98_ & new_n135_;
  assign new_n154_ = new_n111_ & new_n124_;
  assign new_n155_ = ~pq & new_n154_;
  assign new_n156_ = ph & new_n114_;
  assign new_n157_ = ~pq & new_n156_;
  assign new_n158_ = new_n117_ & new_n124_;
  assign new_n159_ = ~pq & new_n158_;
  assign new_n160_ = ~ps & new_n143_;
  assign new_n161_ = ph & new_n111_;
  assign new_n162_ = ~pq & new_n161_;
  assign new_n163_ = new_n125_ & new_n131_;
  assign new_n164_ = pw & new_n163_;
  assign new_n165_ = ph & new_n117_;
  assign new_n166_ = ~pq & new_n165_;
  assign new_n167_ = pu & new_n108_;
  assign new_n168_ = new_n107_ & new_n131_;
  assign new_n169_ = ~pq & new_n168_;
  assign new_n170_ = ~new_n144_ & ~new_n146_;
  assign new_n171_ = ~new_n139_ & ~new_n142_;
  assign new_n172_ = new_n170_ & new_n171_;
  assign new_n173_ = ~new_n137_ & ~new_n138_;
  assign new_n174_ = ~new_n134_ & ~new_n136_;
  assign new_n175_ = new_n173_ & new_n174_;
  assign new_n176_ = new_n172_ & new_n175_;
  assign new_n177_ = ~new_n109_ & ~new_n110_;
  assign new_n178_ = ~new_n113_ & ~new_n116_;
  assign new_n179_ = new_n177_ & new_n178_;
  assign new_n180_ = ~new_n129_ & ~new_n130_;
  assign new_n181_ = ~new_n119_ & ~new_n127_;
  assign new_n182_ = new_n180_ & new_n181_;
  assign new_n183_ = new_n179_ & new_n182_;
  assign new_n184_ = new_n176_ & new_n183_;
  assign new_n185_ = ~new_n167_ & ~new_n169_;
  assign new_n186_ = ~new_n164_ & ~new_n166_;
  assign new_n187_ = new_n185_ & new_n186_;
  assign new_n188_ = ~new_n160_ & ~new_n162_;
  assign new_n189_ = ~new_n157_ & ~new_n159_;
  assign new_n190_ = new_n188_ & new_n189_;
  assign new_n191_ = new_n187_ & new_n190_;
  assign new_n192_ = ~new_n153_ & ~new_n155_;
  assign new_n193_ = ~new_n151_ & ~new_n152_;
  assign new_n194_ = new_n192_ & new_n193_;
  assign new_n195_ = ~new_n147_ & ~new_n148_;
  assign new_n196_ = ~new_n149_ & ~new_n150_;
  assign new_n197_ = new_n195_ & new_n196_;
  assign new_n198_ = new_n194_ & new_n197_;
  assign new_n199_ = new_n191_ & new_n198_;
  assign pc0 = ~new_n184_ | ~new_n199_;
  assign new_n201_ = pu & ~pv;
  assign new_n202_ = pv & ~pi;
  assign new_n203_ = ~ps & ~pv;
  assign new_n204_ = ~new_n201_ & ~new_n202_;
  assign new_n205_ = ~new_n55_ & ~new_n203_;
  assign new_n206_ = new_n204_ & new_n205_;
  assign pd0 = ~pw & new_n206_;
  assign new_n208_ = ~pt & pv;
  assign new_n209_ = ~pu & new_n208_;
  assign new_n210_ = ~ps & new_n209_;
  assign new_n211_ = ~pj & new_n120_;
  assign new_n212_ = ps & new_n57_;
  assign new_n213_ = pu & ~pj;
  assign new_n214_ = ~new_n210_ & ~new_n211_;
  assign new_n215_ = ~new_n212_ & ~new_n213_;
  assign new_n216_ = new_n214_ & new_n215_;
  assign new_n217_ = ~pw & new_n216_;
  assign new_n218_ = ~pu & new_n217_;
  assign new_n219_ = pv & new_n217_;
  assign pe0 = new_n218_ | new_n219_;
  assign pf0 = ~pa & ~pk;
  assign new_n222_ = pk & pm;
  assign new_n223_ = ~pl & new_n222_;
  assign new_n224_ = ~pa & new_n223_;
  assign new_n225_ = pk & ~pn;
  assign new_n226_ = ~pl & new_n225_;
  assign new_n227_ = ~pa & new_n226_;
  assign new_n228_ = ~pk & pl;
  assign new_n229_ = ~pa & new_n228_;
  assign new_n230_ = ~new_n224_ & ~new_n227_;
  assign pg0 = new_n229_ | ~new_n230_;
  assign new_n232_ = ~pl & pm;
  assign new_n233_ = ~pa & new_n232_;
  assign new_n234_ = pk & ~pm;
  assign new_n235_ = pl & new_n234_;
  assign new_n236_ = ~pa & new_n235_;
  assign new_n237_ = ~pk & pm;
  assign new_n238_ = ~pa & new_n237_;
  assign new_n239_ = ~new_n233_ & ~new_n236_;
  assign ph0 = new_n238_ | ~new_n239_;
  assign new_n241_ = ~pl & ~pm;
  assign new_n242_ = pk & new_n241_;
  assign new_n243_ = pl & pn;
  assign new_n244_ = pm & new_n243_;
  assign new_n245_ = pk & new_n244_;
  assign new_n246_ = ~new_n242_ & ~new_n245_;
  assign new_n247_ = ~pa & new_n246_;
  assign new_n248_ = pk & pl;
  assign new_n249_ = pm & new_n248_;
  assign new_n250_ = new_n247_ & new_n249_;
  assign new_n251_ = pn & new_n247_;
  assign pi0 = new_n250_ | new_n251_;
  assign new_n253_ = ~pa & po;
  assign new_n254_ = ~px & new_n253_;
  assign new_n255_ = ~pk & new_n254_;
  assign new_n256_ = pl & new_n254_;
  assign new_n257_ = ~pa & ~po;
  assign new_n258_ = px & new_n257_;
  assign new_n259_ = pl & new_n258_;
  assign new_n260_ = pm & new_n258_;
  assign new_n261_ = ~pk & new_n258_;
  assign new_n262_ = ~pl & pn;
  assign new_n263_ = new_n234_ & new_n262_;
  assign new_n264_ = ~px & ~pa;
  assign new_n265_ = new_n263_ & new_n264_;
  assign new_n266_ = pl & new_n265_;
  assign new_n267_ = pm & new_n265_;
  assign new_n268_ = pn & po;
  assign new_n269_ = ~pa & ~new_n268_;
  assign new_n270_ = new_n263_ & new_n269_;
  assign new_n271_ = ~po & new_n270_;
  assign new_n272_ = ~px & new_n270_;
  assign new_n273_ = new_n257_ & new_n263_;
  assign new_n274_ = pm & new_n273_;
  assign new_n275_ = ~pk & new_n265_;
  assign new_n276_ = pl & new_n273_;
  assign new_n277_ = new_n264_ & ~new_n268_;
  assign new_n278_ = po & new_n277_;
  assign new_n279_ = ~pk & new_n273_;
  assign new_n280_ = pm & new_n254_;
  assign new_n281_ = px & ~pa;
  assign new_n282_ = ~new_n268_ & new_n281_;
  assign new_n283_ = ~po & new_n282_;
  assign new_n284_ = ~new_n280_ & ~new_n283_;
  assign new_n285_ = ~new_n278_ & ~new_n279_;
  assign new_n286_ = new_n284_ & new_n285_;
  assign new_n287_ = ~new_n275_ & ~new_n276_;
  assign new_n288_ = ~new_n272_ & ~new_n274_;
  assign new_n289_ = new_n287_ & new_n288_;
  assign new_n290_ = new_n286_ & new_n289_;
  assign new_n291_ = ~new_n255_ & ~new_n256_;
  assign new_n292_ = ~new_n259_ & ~new_n260_;
  assign new_n293_ = new_n291_ & new_n292_;
  assign new_n294_ = ~new_n267_ & ~new_n271_;
  assign new_n295_ = ~new_n261_ & ~new_n266_;
  assign new_n296_ = new_n294_ & new_n295_;
  assign new_n297_ = new_n293_ & new_n296_;
  assign pj0 = ~new_n290_ | ~new_n297_;
  assign new_n299_ = ~pe & new_n120_;
  assign new_n300_ = ~ps & pv;
  assign new_n301_ = ~pe & new_n300_;
  assign new_n302_ = pu & ~pe;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = ~new_n210_ & ~new_n299_;
  assign new_n305_ = ~new_n201_ & new_n304_;
  assign new_n306_ = new_n303_ & new_n305_;
  assign pz = ~pw & new_n306_;
  assign new_n308_ = ~pq & pr;
  assign new_n309_ = px & new_n308_;
  assign new_n310_ = po & new_n309_;
  assign new_n311_ = ~pp & ~po;
  assign new_n312_ = pp & px;
  assign new_n313_ = po & new_n312_;
  assign new_n314_ = ~new_n310_ & ~new_n311_;
  assign new_n315_ = ~pa & ~new_n313_;
  assign new_n316_ = new_n314_ & new_n315_;
  assign new_n317_ = ~pp & ~new_n308_;
  assign new_n318_ = px & new_n316_;
  assign new_n319_ = new_n317_ & new_n318_;
  assign new_n320_ = pp & new_n316_;
  assign new_n321_ = pl & new_n320_;
  assign new_n322_ = ~pk & new_n318_;
  assign new_n323_ = ~pm & pn;
  assign new_n324_ = po & new_n323_;
  assign new_n325_ = new_n318_ & ~new_n324_;
  assign new_n326_ = pl & new_n318_;
  assign new_n327_ = new_n263_ & new_n316_;
  assign new_n328_ = ~new_n324_ & new_n327_;
  assign new_n329_ = new_n317_ & new_n327_;
  assign new_n330_ = ~pk & new_n327_;
  assign new_n331_ = new_n317_ & new_n320_;
  assign new_n332_ = pl & new_n327_;
  assign new_n333_ = ~pk & new_n320_;
  assign new_n334_ = new_n320_ & ~new_n324_;
  assign new_n335_ = ~new_n332_ & ~new_n333_;
  assign new_n336_ = ~new_n334_ & new_n335_;
  assign new_n337_ = ~new_n329_ & ~new_n330_;
  assign new_n338_ = ~new_n331_ & new_n337_;
  assign new_n339_ = new_n336_ & new_n338_;
  assign new_n340_ = ~new_n319_ & ~new_n321_;
  assign new_n341_ = ~new_n322_ & new_n340_;
  assign new_n342_ = ~new_n325_ & ~new_n326_;
  assign new_n343_ = ~new_n328_ & new_n342_;
  assign new_n344_ = new_n341_ & new_n343_;
  assign pk0 = ~new_n339_ | ~new_n344_;
  assign new_n346_ = ~pq & ~po;
  assign new_n347_ = ~pp & ~pq;
  assign new_n348_ = ~new_n346_ & ~new_n347_;
  assign new_n349_ = ~pa & new_n348_;
  assign new_n350_ = px & new_n349_;
  assign new_n351_ = ~pp & new_n350_;
  assign new_n352_ = ~pq & new_n350_;
  assign new_n353_ = pq & new_n349_;
  assign new_n354_ = ~pp & new_n353_;
  assign new_n355_ = ~po & new_n350_;
  assign new_n356_ = ~po & new_n353_;
  assign new_n357_ = ~pm & new_n262_;
  assign new_n358_ = pk & new_n357_;
  assign new_n359_ = ~px & ~new_n358_;
  assign new_n360_ = new_n349_ & new_n359_;
  assign new_n361_ = new_n263_ & new_n360_;
  assign new_n362_ = px & new_n360_;
  assign new_n363_ = new_n263_ & new_n349_;
  assign new_n364_ = ~pq & new_n363_;
  assign new_n365_ = pq & new_n360_;
  assign new_n366_ = ~po & new_n363_;
  assign new_n367_ = ~pp & new_n363_;
  assign new_n368_ = ~new_n351_ & ~new_n352_;
  assign new_n369_ = ~new_n354_ & new_n368_;
  assign new_n370_ = ~new_n355_ & ~new_n356_;
  assign new_n371_ = ~new_n361_ & new_n370_;
  assign new_n372_ = new_n369_ & new_n371_;
  assign new_n373_ = ~new_n366_ & ~new_n367_;
  assign new_n374_ = ~new_n362_ & ~new_n364_;
  assign new_n375_ = ~new_n365_ & new_n374_;
  assign new_n376_ = new_n373_ & new_n375_;
  assign pl0 = ~new_n372_ | ~new_n376_;
  assign new_n378_ = ~pq & ~pr;
  assign new_n379_ = ~pr & ~po;
  assign new_n380_ = ~pp & ~pr;
  assign new_n381_ = ~new_n378_ & ~new_n379_;
  assign new_n382_ = ~pa & ~new_n380_;
  assign new_n383_ = new_n381_ & new_n382_;
  assign new_n384_ = ~po & new_n383_;
  assign new_n385_ = px & new_n384_;
  assign new_n386_ = ~pk & new_n385_;
  assign new_n387_ = pl & new_n385_;
  assign new_n388_ = pq & pr;
  assign new_n389_ = pp & new_n388_;
  assign new_n390_ = ~new_n347_ & ~new_n389_;
  assign new_n391_ = new_n383_ & new_n390_;
  assign new_n392_ = new_n263_ & new_n391_;
  assign new_n393_ = pr & new_n391_;
  assign new_n394_ = px & new_n391_;
  assign new_n395_ = ~new_n324_ & new_n383_;
  assign new_n396_ = pr & new_n395_;
  assign new_n397_ = ~po & new_n396_;
  assign new_n398_ = ~px & new_n396_;
  assign new_n399_ = pr & new_n384_;
  assign new_n400_ = ~pk & new_n399_;
  assign new_n401_ = pl & new_n399_;
  assign new_n402_ = ~px & new_n383_;
  assign new_n403_ = pr & new_n402_;
  assign new_n404_ = ~pk & new_n403_;
  assign new_n405_ = pl & new_n403_;
  assign new_n406_ = new_n263_ & new_n383_;
  assign new_n407_ = ~new_n324_ & new_n406_;
  assign new_n408_ = ~po & new_n407_;
  assign new_n409_ = ~px & new_n407_;
  assign new_n410_ = px & new_n383_;
  assign new_n411_ = ~new_n324_ & new_n410_;
  assign new_n412_ = ~po & new_n411_;
  assign new_n413_ = new_n263_ & new_n402_;
  assign new_n414_ = ~pk & new_n413_;
  assign new_n415_ = pl & new_n413_;
  assign new_n416_ = new_n263_ & new_n384_;
  assign new_n417_ = ~pk & new_n416_;
  assign new_n418_ = pl & new_n416_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = ~new_n414_ & ~new_n415_;
  assign new_n421_ = new_n419_ & new_n420_;
  assign new_n422_ = ~new_n409_ & ~new_n412_;
  assign new_n423_ = ~new_n404_ & ~new_n405_;
  assign new_n424_ = ~new_n408_ & new_n423_;
  assign new_n425_ = new_n422_ & new_n424_;
  assign new_n426_ = new_n421_ & new_n425_;
  assign new_n427_ = ~new_n400_ & ~new_n401_;
  assign new_n428_ = ~new_n397_ & ~new_n398_;
  assign new_n429_ = new_n427_ & new_n428_;
  assign new_n430_ = ~new_n393_ & ~new_n394_;
  assign new_n431_ = ~new_n386_ & ~new_n387_;
  assign new_n432_ = ~new_n392_ & new_n431_;
  assign new_n433_ = new_n430_ & new_n432_;
  assign new_n434_ = new_n429_ & new_n433_;
  assign pm0 = ~new_n426_ | ~new_n434_;
  assign new_n436_ = ps & ~pa;
  assign new_n437_ = new_n359_ & new_n436_;
  assign new_n438_ = po & ~new_n359_;
  assign new_n439_ = ~pp & new_n308_;
  assign new_n440_ = new_n438_ & new_n439_;
  assign new_n441_ = ~pa & new_n440_;
  assign new_n442_ = pp & new_n441_;
  assign new_n443_ = ~po & new_n436_;
  assign new_n444_ = ps & new_n308_;
  assign new_n445_ = new_n436_ & ~new_n444_;
  assign new_n446_ = pp & new_n436_;
  assign new_n447_ = new_n359_ & new_n441_;
  assign new_n448_ = ~po & new_n441_;
  assign new_n449_ = new_n441_ & ~new_n444_;
  assign new_n450_ = ~new_n437_ & ~new_n442_;
  assign new_n451_ = ~new_n443_ & ~new_n445_;
  assign new_n452_ = new_n450_ & new_n451_;
  assign new_n453_ = ~new_n448_ & ~new_n449_;
  assign new_n454_ = ~new_n446_ & ~new_n447_;
  assign new_n455_ = new_n453_ & new_n454_;
  assign pn0 = ~new_n452_ | ~new_n455_;
  assign new_n457_ = ~pl & new_n234_;
  assign new_n458_ = pn & new_n457_;
  assign new_n459_ = ~px & ~new_n458_;
  assign new_n460_ = ~new_n60_ & ~new_n459_;
  assign new_n461_ = ~pp & po;
  assign new_n462_ = ~pq & ps;
  assign new_n463_ = pr & ~pt;
  assign new_n464_ = new_n462_ & new_n463_;
  assign new_n465_ = new_n460_ & new_n461_;
  assign new_n466_ = new_n464_ & new_n465_;
  assign new_n467_ = ~pa & new_n466_;
  assign new_n468_ = pr & po;
  assign new_n469_ = new_n462_ & new_n468_;
  assign new_n470_ = ~pp & new_n469_;
  assign new_n471_ = new_n263_ & new_n470_;
  assign new_n472_ = px & new_n470_;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign new_n474_ = pt & new_n473_;
  assign new_n475_ = ~pa & new_n474_;
  assign po0 = new_n467_ | new_n475_;
  assign new_n477_ = ~px & ~pn;
  assign new_n478_ = ~px & pl;
  assign new_n479_ = ~px & pm;
  assign new_n480_ = ~px & ~pk;
  assign new_n481_ = ~new_n477_ & ~new_n478_;
  assign new_n482_ = ~new_n479_ & ~new_n480_;
  assign new_n483_ = new_n481_ & new_n482_;
  assign new_n484_ = ~pq & new_n461_;
  assign new_n485_ = pr & pt;
  assign new_n486_ = ps & ~pu;
  assign new_n487_ = new_n485_ & new_n486_;
  assign new_n488_ = new_n483_ & new_n484_;
  assign new_n489_ = new_n487_ & new_n488_;
  assign new_n490_ = ~pa & new_n489_;
  assign new_n491_ = ps & po;
  assign new_n492_ = new_n485_ & new_n491_;
  assign new_n493_ = ~pp & new_n492_;
  assign new_n494_ = ~pq & new_n493_;
  assign new_n495_ = new_n263_ & new_n494_;
  assign new_n496_ = px & new_n494_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = pu & new_n497_;
  assign new_n499_ = ~pa & new_n498_;
  assign pp0 = new_n490_ | new_n499_;
  assign new_n501_ = ps & pu;
  assign new_n502_ = new_n57_ & new_n501_;
  assign new_n503_ = ~pq & po;
  assign new_n504_ = ~pp & pr;
  assign new_n505_ = new_n503_ & new_n504_;
  assign new_n506_ = new_n483_ & new_n502_;
  assign new_n507_ = new_n505_ & new_n506_;
  assign new_n508_ = ~pa & new_n507_;
  assign new_n509_ = pr & ~pu;
  assign new_n510_ = ps & new_n509_;
  assign new_n511_ = ~pt & new_n510_;
  assign new_n512_ = pr & pu;
  assign new_n513_ = ps & new_n512_;
  assign new_n514_ = pt & new_n513_;
  assign new_n515_ = ~new_n511_ & ~new_n514_;
  assign new_n516_ = po & ~new_n515_;
  assign new_n517_ = ~pp & new_n516_;
  assign new_n518_ = ~pq & new_n517_;
  assign new_n519_ = new_n263_ & new_n518_;
  assign new_n520_ = px & new_n518_;
  assign new_n521_ = ~new_n519_ & ~new_n520_;
  assign new_n522_ = pv & new_n521_;
  assign new_n523_ = ~pa & new_n522_;
  assign pq0 = new_n508_ | new_n523_;
  assign new_n525_ = pw & ~pa;
  assign new_n526_ = ~new_n49_ & new_n525_;
  assign new_n527_ = ~pt & new_n58_;
  assign new_n528_ = ~ps & pu;
  assign new_n529_ = new_n527_ & new_n528_;
  assign new_n530_ = ~pa & new_n529_;
  assign new_n531_ = ~pu & new_n530_;
  assign new_n532_ = pt & new_n525_;
  assign new_n533_ = ~ps & new_n525_;
  assign new_n534_ = ~pu & new_n525_;
  assign new_n535_ = ~new_n49_ & new_n530_;
  assign new_n536_ = pt & new_n530_;
  assign new_n537_ = ~ps & new_n530_;
  assign new_n538_ = ~new_n526_ & ~new_n531_;
  assign new_n539_ = ~new_n532_ & ~new_n533_;
  assign new_n540_ = new_n538_ & new_n539_;
  assign new_n541_ = ~new_n536_ & ~new_n537_;
  assign new_n542_ = ~new_n534_ & ~new_n535_;
  assign new_n543_ = new_n541_ & new_n542_;
  assign pr0 = ~new_n540_ | ~new_n543_;
  assign new_n545_ = ~px & pb;
  assign new_n546_ = ~pa & new_n545_;
  assign new_n547_ = px & ~pb;
  assign new_n548_ = ~pa & new_n547_;
  assign ps0 = new_n546_ | new_n548_;
  assign new_n550_ = ~py & pc;
  assign new_n551_ = ~pa & new_n550_;
  assign new_n552_ = py & ~pc;
  assign new_n553_ = ~pa & new_n552_;
  assign pt0 = new_n551_ | new_n553_;
endmodule

