module i2 ( 
    \V62(1) , \V30(31) , \V30(29) , \V30(27) , \V30(25) , \V30(23) ,
    \V30(21) , \V30(19) , \V30(17) , \V30(15) , \V30(13) , \V30(11) ,
    \V30(9) , \V30(7) , \V30(5) , \V30(3) , \V30(2) , \V30(4) , \V30(6) ,
    \V30(8) , \V30(10) , \V30(12) , \V30(14) , \V30(16) , \V30(18) ,
    \V30(20) , \V30(22) , \V30(24) , \V30(26) , \V30(28) , \V30(30) ,
    \V62(0) , \V64(0) , \V62(31) , \V62(29) , \V62(27) , \V62(25) ,
    \V62(23) , \V62(21) , \V62(19) , \V62(17) , \V62(15) , \V62(13) ,
    \V62(11) , \V62(9) , \V62(7) , \V62(5) , \V62(3) , \V62(2) , \V62(4) ,
    \V62(6) , \V62(8) , \V62(10) , \V62(12) , \V62(14) , \V62(16) ,
    \V62(18) , \V62(20) , \V62(22) , \V62(24) , \V62(26) , \V62(28) ,
    \V62(30) , \V63(0) , \V126(1) , \V94(31) , \V94(29) , \V94(27) ,
    \V94(25) , \V94(23) , \V94(21) , \V94(19) , \V94(17) , \V94(15) ,
    \V94(13) , \V94(11) , \V94(9) , \V94(7) , \V94(5) , \V94(3) , \V94(2) ,
    \V94(4) , \V94(6) , \V94(8) , \V94(10) , \V94(12) , \V94(14) ,
    \V94(16) , \V94(18) , \V94(20) , \V94(22) , \V94(24) , \V94(26) ,
    \V94(28) , \V94(30) , \V126(0) , \V128(0) , \V126(31) , \V126(29) ,
    \V126(27) , \V126(25) , \V126(23) , \V126(21) , \V126(19) , \V126(17) ,
    \V126(15) , \V126(13) , \V126(11) , \V126(9) , \V126(7) , \V126(5) ,
    \V126(3) , \V126(2) , \V126(4) , \V126(6) , \V126(8) , \V126(10) ,
    \V126(12) , \V126(14) , \V126(16) , \V126(18) , \V126(20) , \V126(22) ,
    \V126(24) , \V126(26) , \V126(28) , \V126(30) , \V127(0) , \V201(0) ,
    \V129(0) , \V201(1) , \V130(0) , \V176(1) , \V144(31) , \V144(29) ,
    \V144(27) , \V144(25) , \V144(23) , \V144(21) , \V144(19) , \V144(18) ,
    \V144(20) , \V144(22) , \V144(24) , \V144(26) , \V144(28) , \V144(30) ,
    \V176(0) , \V176(17) , \V176(15) , \V176(13) , \V176(11) , \V176(9) ,
    \V176(7) , \V176(5) , \V176(3) , \V176(2) , \V176(4) , \V176(6) ,
    \V176(8) , \V176(10) , \V176(12) , \V176(14) , \V176(16) , \V178(1) ,
    \V176(31) , \V176(29) , \V176(27) , \V176(25) , \V176(23) , \V176(21) ,
    \V176(19) , \V176(18) , \V176(20) , \V176(22) , \V176(24) , \V176(26) ,
    \V176(28) , \V176(30) , \V178(0) , \V201(3) , \V201(2) , \V188(25) ,
    \V188(23) , \V188(22) , \V188(24) , \V188(29) , \V188(27) , \V188(26) ,
    \V188(28) , \V190(1) , \V188(31) , \V188(30) , \V190(0) , \V201(5) ,
    \V201(4) , \V201(7) , \V191(31) , \V201(6) , \V193(0) , \V193(1) ,
    \V202(0)   );
  input  \V62(1) , \V30(31) , \V30(29) , \V30(27) , \V30(25) , \V30(23) ,
    \V30(21) , \V30(19) , \V30(17) , \V30(15) , \V30(13) , \V30(11) ,
    \V30(9) , \V30(7) , \V30(5) , \V30(3) , \V30(2) , \V30(4) , \V30(6) ,
    \V30(8) , \V30(10) , \V30(12) , \V30(14) , \V30(16) , \V30(18) ,
    \V30(20) , \V30(22) , \V30(24) , \V30(26) , \V30(28) , \V30(30) ,
    \V62(0) , \V64(0) , \V62(31) , \V62(29) , \V62(27) , \V62(25) ,
    \V62(23) , \V62(21) , \V62(19) , \V62(17) , \V62(15) , \V62(13) ,
    \V62(11) , \V62(9) , \V62(7) , \V62(5) , \V62(3) , \V62(2) , \V62(4) ,
    \V62(6) , \V62(8) , \V62(10) , \V62(12) , \V62(14) , \V62(16) ,
    \V62(18) , \V62(20) , \V62(22) , \V62(24) , \V62(26) , \V62(28) ,
    \V62(30) , \V63(0) , \V126(1) , \V94(31) , \V94(29) , \V94(27) ,
    \V94(25) , \V94(23) , \V94(21) , \V94(19) , \V94(17) , \V94(15) ,
    \V94(13) , \V94(11) , \V94(9) , \V94(7) , \V94(5) , \V94(3) , \V94(2) ,
    \V94(4) , \V94(6) , \V94(8) , \V94(10) , \V94(12) , \V94(14) ,
    \V94(16) , \V94(18) , \V94(20) , \V94(22) , \V94(24) , \V94(26) ,
    \V94(28) , \V94(30) , \V126(0) , \V128(0) , \V126(31) , \V126(29) ,
    \V126(27) , \V126(25) , \V126(23) , \V126(21) , \V126(19) , \V126(17) ,
    \V126(15) , \V126(13) , \V126(11) , \V126(9) , \V126(7) , \V126(5) ,
    \V126(3) , \V126(2) , \V126(4) , \V126(6) , \V126(8) , \V126(10) ,
    \V126(12) , \V126(14) , \V126(16) , \V126(18) , \V126(20) , \V126(22) ,
    \V126(24) , \V126(26) , \V126(28) , \V126(30) , \V127(0) , \V201(0) ,
    \V129(0) , \V201(1) , \V130(0) , \V176(1) , \V144(31) , \V144(29) ,
    \V144(27) , \V144(25) , \V144(23) , \V144(21) , \V144(19) , \V144(18) ,
    \V144(20) , \V144(22) , \V144(24) , \V144(26) , \V144(28) , \V144(30) ,
    \V176(0) , \V176(17) , \V176(15) , \V176(13) , \V176(11) , \V176(9) ,
    \V176(7) , \V176(5) , \V176(3) , \V176(2) , \V176(4) , \V176(6) ,
    \V176(8) , \V176(10) , \V176(12) , \V176(14) , \V176(16) , \V178(1) ,
    \V176(31) , \V176(29) , \V176(27) , \V176(25) , \V176(23) , \V176(21) ,
    \V176(19) , \V176(18) , \V176(20) , \V176(22) , \V176(24) , \V176(26) ,
    \V176(28) , \V176(30) , \V178(0) , \V201(3) , \V201(2) , \V188(25) ,
    \V188(23) , \V188(22) , \V188(24) , \V188(29) , \V188(27) , \V188(26) ,
    \V188(28) , \V190(1) , \V188(31) , \V188(30) , \V190(0) , \V201(5) ,
    \V201(4) , \V201(7) , \V191(31) , \V201(6) , \V193(0) , \V193(1) ;
  output \V202(0) ;
  wire new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_;
  assign new_n203_ = \V201(7)  & \V193(1) ;
  assign new_n204_ = \V201(6)  & \V193(0) ;
  assign new_n205_ = \V201(7)  & new_n204_;
  assign new_n206_ = ~\V188(30)  & ~\V190(0) ;
  assign new_n207_ = ~\V190(1)  & ~\V188(31) ;
  assign new_n208_ = new_n206_ & new_n207_;
  assign new_n209_ = \V201(5)  & ~new_n208_;
  assign new_n210_ = ~\V188(26)  & ~\V188(28) ;
  assign new_n211_ = ~\V188(29)  & ~\V188(27) ;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_ = \V201(4)  & ~new_n212_;
  assign new_n214_ = \V201(5)  & new_n213_;
  assign new_n215_ = ~\V176(30)  & ~\V178(0) ;
  assign new_n216_ = ~\V176(26)  & ~\V176(28) ;
  assign new_n217_ = new_n215_ & new_n216_;
  assign new_n218_ = ~\V176(22)  & ~\V176(24) ;
  assign new_n219_ = ~\V176(18)  & ~\V176(20) ;
  assign new_n220_ = new_n218_ & new_n219_;
  assign new_n221_ = new_n217_ & new_n220_;
  assign new_n222_ = ~\V176(21)  & ~\V176(19) ;
  assign new_n223_ = ~\V176(25)  & ~\V176(23) ;
  assign new_n224_ = new_n222_ & new_n223_;
  assign new_n225_ = ~\V176(29)  & ~\V176(27) ;
  assign new_n226_ = ~\V178(1)  & ~\V176(31) ;
  assign new_n227_ = new_n225_ & new_n226_;
  assign new_n228_ = new_n224_ & new_n227_;
  assign new_n229_ = new_n221_ & new_n228_;
  assign new_n230_ = \V201(3)  & ~new_n229_;
  assign new_n231_ = ~\V176(14)  & ~\V176(16) ;
  assign new_n232_ = ~\V176(10)  & ~\V176(12) ;
  assign new_n233_ = new_n231_ & new_n232_;
  assign new_n234_ = ~\V176(6)  & ~\V176(8) ;
  assign new_n235_ = ~\V176(2)  & ~\V176(4) ;
  assign new_n236_ = new_n234_ & new_n235_;
  assign new_n237_ = new_n233_ & new_n236_;
  assign new_n238_ = ~\V176(5)  & ~\V176(3) ;
  assign new_n239_ = ~\V176(9)  & ~\V176(7) ;
  assign new_n240_ = new_n238_ & new_n239_;
  assign new_n241_ = ~\V176(13)  & ~\V176(11) ;
  assign new_n242_ = ~\V176(17)  & ~\V176(15) ;
  assign new_n243_ = new_n241_ & new_n242_;
  assign new_n244_ = new_n240_ & new_n243_;
  assign new_n245_ = new_n237_ & new_n244_;
  assign new_n246_ = \V201(2)  & ~new_n245_;
  assign new_n247_ = \V201(3)  & new_n246_;
  assign new_n248_ = ~\V126(30)  & ~\V127(0) ;
  assign new_n249_ = ~\V126(26)  & ~\V126(28) ;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = ~\V126(22)  & ~\V126(24) ;
  assign new_n252_ = ~\V126(18)  & ~\V126(20) ;
  assign new_n253_ = new_n251_ & new_n252_;
  assign new_n254_ = new_n250_ & new_n253_;
  assign new_n255_ = ~\V126(14)  & ~\V126(16) ;
  assign new_n256_ = ~\V126(10)  & ~\V126(12) ;
  assign new_n257_ = new_n255_ & new_n256_;
  assign new_n258_ = ~\V126(6)  & ~\V126(8) ;
  assign new_n259_ = ~\V126(2)  & ~\V126(4) ;
  assign new_n260_ = new_n258_ & new_n259_;
  assign new_n261_ = new_n257_ & new_n260_;
  assign new_n262_ = new_n254_ & new_n261_;
  assign new_n263_ = ~\V126(5)  & ~\V126(3) ;
  assign new_n264_ = ~\V126(9)  & ~\V126(7) ;
  assign new_n265_ = new_n263_ & new_n264_;
  assign new_n266_ = ~\V126(13)  & ~\V126(11) ;
  assign new_n267_ = ~\V126(17)  & ~\V126(15) ;
  assign new_n268_ = new_n266_ & new_n267_;
  assign new_n269_ = new_n265_ & new_n268_;
  assign new_n270_ = ~\V126(21)  & ~\V126(19) ;
  assign new_n271_ = ~\V126(25)  & ~\V126(23) ;
  assign new_n272_ = new_n270_ & new_n271_;
  assign new_n273_ = ~\V126(29)  & ~\V126(27) ;
  assign new_n274_ = ~\V128(0)  & ~\V126(31) ;
  assign new_n275_ = new_n273_ & new_n274_;
  assign new_n276_ = new_n272_ & new_n275_;
  assign new_n277_ = new_n269_ & new_n276_;
  assign new_n278_ = new_n262_ & new_n277_;
  assign new_n279_ = \V201(1)  & ~new_n278_;
  assign new_n280_ = \V201(0)  & new_n279_;
  assign new_n281_ = \V201(0)  & \V130(0) ;
  assign new_n282_ = ~\V30(30)  & ~\V62(0) ;
  assign new_n283_ = ~\V30(26)  & ~\V30(28) ;
  assign new_n284_ = new_n282_ & new_n283_;
  assign new_n285_ = ~\V30(22)  & ~\V30(24) ;
  assign new_n286_ = ~\V30(18)  & ~\V30(20) ;
  assign new_n287_ = new_n285_ & new_n286_;
  assign new_n288_ = new_n284_ & new_n287_;
  assign new_n289_ = ~\V30(14)  & ~\V30(16) ;
  assign new_n290_ = ~\V30(10)  & ~\V30(12) ;
  assign new_n291_ = new_n289_ & new_n290_;
  assign new_n292_ = ~\V30(6)  & ~\V30(8) ;
  assign new_n293_ = ~\V30(2)  & ~\V30(4) ;
  assign new_n294_ = new_n292_ & new_n293_;
  assign new_n295_ = new_n291_ & new_n294_;
  assign new_n296_ = new_n288_ & new_n295_;
  assign new_n297_ = ~\V30(5)  & ~\V30(3) ;
  assign new_n298_ = ~\V30(9)  & ~\V30(7) ;
  assign new_n299_ = new_n297_ & new_n298_;
  assign new_n300_ = ~\V30(13)  & ~\V30(11) ;
  assign new_n301_ = ~\V30(17)  & ~\V30(15) ;
  assign new_n302_ = new_n300_ & new_n301_;
  assign new_n303_ = new_n299_ & new_n302_;
  assign new_n304_ = ~\V30(21)  & ~\V30(19) ;
  assign new_n305_ = ~\V30(25)  & ~\V30(23) ;
  assign new_n306_ = new_n304_ & new_n305_;
  assign new_n307_ = ~\V30(29)  & ~\V30(27) ;
  assign new_n308_ = ~\V62(1)  & ~\V30(31) ;
  assign new_n309_ = new_n307_ & new_n308_;
  assign new_n310_ = new_n306_ & new_n309_;
  assign new_n311_ = new_n303_ & new_n310_;
  assign new_n312_ = new_n296_ & new_n311_;
  assign new_n313_ = \V201(1)  & ~new_n312_;
  assign new_n314_ = ~\V201(0)  & new_n313_;
  assign new_n315_ = ~\V201(0)  & \V129(0) ;
  assign new_n316_ = ~\V62(30)  & ~\V63(0) ;
  assign new_n317_ = ~\V62(26)  & ~\V62(28) ;
  assign new_n318_ = new_n316_ & new_n317_;
  assign new_n319_ = ~\V62(22)  & ~\V62(24) ;
  assign new_n320_ = ~\V62(18)  & ~\V62(20) ;
  assign new_n321_ = new_n319_ & new_n320_;
  assign new_n322_ = new_n318_ & new_n321_;
  assign new_n323_ = ~\V62(14)  & ~\V62(16) ;
  assign new_n324_ = ~\V62(10)  & ~\V62(12) ;
  assign new_n325_ = new_n323_ & new_n324_;
  assign new_n326_ = ~\V62(6)  & ~\V62(8) ;
  assign new_n327_ = ~\V62(2)  & ~\V62(4) ;
  assign new_n328_ = new_n326_ & new_n327_;
  assign new_n329_ = new_n325_ & new_n328_;
  assign new_n330_ = new_n322_ & new_n329_;
  assign new_n331_ = ~\V62(5)  & ~\V62(3) ;
  assign new_n332_ = ~\V62(9)  & ~\V62(7) ;
  assign new_n333_ = new_n331_ & new_n332_;
  assign new_n334_ = ~\V62(13)  & ~\V62(11) ;
  assign new_n335_ = ~\V62(17)  & ~\V62(15) ;
  assign new_n336_ = new_n334_ & new_n335_;
  assign new_n337_ = new_n333_ & new_n336_;
  assign new_n338_ = ~\V62(21)  & ~\V62(19) ;
  assign new_n339_ = ~\V62(25)  & ~\V62(23) ;
  assign new_n340_ = new_n338_ & new_n339_;
  assign new_n341_ = ~\V62(29)  & ~\V62(27) ;
  assign new_n342_ = ~\V64(0)  & ~\V62(31) ;
  assign new_n343_ = new_n341_ & new_n342_;
  assign new_n344_ = new_n340_ & new_n343_;
  assign new_n345_ = new_n337_ & new_n344_;
  assign new_n346_ = new_n330_ & new_n345_;
  assign new_n347_ = \V201(1)  & ~new_n346_;
  assign new_n348_ = ~\V201(0)  & new_n347_;
  assign new_n349_ = ~\V94(30)  & ~\V126(0) ;
  assign new_n350_ = ~\V94(26)  & ~\V94(28) ;
  assign new_n351_ = new_n349_ & new_n350_;
  assign new_n352_ = ~\V94(22)  & ~\V94(24) ;
  assign new_n353_ = ~\V94(18)  & ~\V94(20) ;
  assign new_n354_ = new_n352_ & new_n353_;
  assign new_n355_ = new_n351_ & new_n354_;
  assign new_n356_ = ~\V94(14)  & ~\V94(16) ;
  assign new_n357_ = ~\V94(10)  & ~\V94(12) ;
  assign new_n358_ = new_n356_ & new_n357_;
  assign new_n359_ = ~\V94(6)  & ~\V94(8) ;
  assign new_n360_ = ~\V94(2)  & ~\V94(4) ;
  assign new_n361_ = new_n359_ & new_n360_;
  assign new_n362_ = new_n358_ & new_n361_;
  assign new_n363_ = new_n355_ & new_n362_;
  assign new_n364_ = ~\V94(5)  & ~\V94(3) ;
  assign new_n365_ = ~\V94(9)  & ~\V94(7) ;
  assign new_n366_ = new_n364_ & new_n365_;
  assign new_n367_ = ~\V94(13)  & ~\V94(11) ;
  assign new_n368_ = ~\V94(17)  & ~\V94(15) ;
  assign new_n369_ = new_n367_ & new_n368_;
  assign new_n370_ = new_n366_ & new_n369_;
  assign new_n371_ = ~\V94(21)  & ~\V94(19) ;
  assign new_n372_ = ~\V94(25)  & ~\V94(23) ;
  assign new_n373_ = new_n371_ & new_n372_;
  assign new_n374_ = ~\V94(29)  & ~\V94(27) ;
  assign new_n375_ = ~\V126(1)  & ~\V94(31) ;
  assign new_n376_ = new_n374_ & new_n375_;
  assign new_n377_ = new_n373_ & new_n376_;
  assign new_n378_ = new_n370_ & new_n377_;
  assign new_n379_ = new_n363_ & new_n378_;
  assign new_n380_ = \V201(1)  & ~new_n379_;
  assign new_n381_ = \V201(0)  & new_n380_;
  assign new_n382_ = ~\V144(30)  & ~\V176(0) ;
  assign new_n383_ = ~\V144(26)  & ~\V144(28) ;
  assign new_n384_ = new_n382_ & new_n383_;
  assign new_n385_ = ~\V144(22)  & ~\V144(24) ;
  assign new_n386_ = ~\V144(18)  & ~\V144(20) ;
  assign new_n387_ = new_n385_ & new_n386_;
  assign new_n388_ = new_n384_ & new_n387_;
  assign new_n389_ = ~\V144(21)  & ~\V144(19) ;
  assign new_n390_ = ~\V144(25)  & ~\V144(23) ;
  assign new_n391_ = new_n389_ & new_n390_;
  assign new_n392_ = ~\V144(29)  & ~\V144(27) ;
  assign new_n393_ = ~\V176(1)  & ~\V144(31) ;
  assign new_n394_ = new_n392_ & new_n393_;
  assign new_n395_ = new_n391_ & new_n394_;
  assign new_n396_ = new_n388_ & new_n395_;
  assign new_n397_ = \V201(3)  & ~new_n396_;
  assign new_n398_ = \V201(2)  & new_n397_;
  assign new_n399_ = \V201(2)  & ~new_n229_;
  assign new_n400_ = \V201(3)  & new_n399_;
  assign new_n401_ = ~\V188(22)  & ~\V188(24) ;
  assign new_n402_ = ~\V188(25)  & ~\V188(23) ;
  assign new_n403_ = new_n401_ & new_n402_;
  assign new_n404_ = \V201(5)  & ~new_n403_;
  assign new_n405_ = \V201(4)  & new_n404_;
  assign new_n406_ = \V201(4)  & ~new_n208_;
  assign new_n407_ = \V201(5)  & new_n406_;
  assign new_n408_ = \V201(7)  & \V191(31) ;
  assign new_n409_ = \V201(6)  & new_n408_;
  assign new_n410_ = \V201(6)  & \V193(1) ;
  assign new_n411_ = \V201(7)  & new_n410_;
  assign new_n412_ = ~new_n409_ & ~new_n411_;
  assign new_n413_ = ~new_n410_ & new_n412_;
  assign new_n414_ = ~new_n405_ & ~new_n407_;
  assign new_n415_ = ~new_n406_ & new_n414_;
  assign new_n416_ = new_n413_ & new_n415_;
  assign new_n417_ = ~new_n398_ & ~new_n400_;
  assign new_n418_ = ~new_n399_ & new_n417_;
  assign new_n419_ = ~new_n315_ & ~new_n348_;
  assign new_n420_ = ~new_n381_ & new_n419_;
  assign new_n421_ = new_n418_ & new_n420_;
  assign new_n422_ = new_n416_ & new_n421_;
  assign new_n423_ = ~new_n280_ & ~new_n281_;
  assign new_n424_ = ~new_n314_ & new_n423_;
  assign new_n425_ = ~new_n230_ & ~new_n246_;
  assign new_n426_ = ~new_n247_ & new_n425_;
  assign new_n427_ = new_n424_ & new_n426_;
  assign new_n428_ = ~new_n209_ & ~new_n213_;
  assign new_n429_ = ~new_n214_ & new_n428_;
  assign new_n430_ = ~new_n203_ & ~new_n204_;
  assign new_n431_ = ~new_n205_ & new_n430_;
  assign new_n432_ = new_n429_ & new_n431_;
  assign new_n433_ = new_n427_ & new_n432_;
  assign \V202(0)  = ~new_n422_ | ~new_n433_;
endmodule

