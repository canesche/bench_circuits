module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3, pj0,
    pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4, pl1,
    pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0, pp0,
    pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3, pq2,
    pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2, pu3,
    pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0, pz3,
    pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po,
    pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3,
    pj0, pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4,
    pl1, pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0,
    pp0, pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3,
    pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2,
    pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0,
    pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po;
  output pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5;
  wire new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1516_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1562_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1706_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1879_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1919_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2081_;
  assign pe5 = pm0 & pn3;
  assign pf6 = ~pl4 | ~pk1;
  assign new_n285_ = ~pi1 & ~ph1;
  assign new_n286_ = ~pj1 & new_n285_;
  assign new_n287_ = ~pk1 & new_n286_;
  assign new_n288_ = ~pl1 & new_n287_;
  assign new_n289_ = ~pa4 & pz3;
  assign new_n290_ = ~px3 & new_n289_;
  assign new_n291_ = py3 & new_n290_;
  assign new_n292_ = ~pb4 & new_n291_;
  assign new_n293_ = ~pc4 & new_n292_;
  assign new_n294_ = pl4 & ~new_n293_;
  assign new_n295_ = ~new_n288_ & ~new_n294_;
  assign new_n296_ = ~px1 & new_n295_;
  assign new_n297_ = po0 & ~pq0;
  assign new_n298_ = pn0 & new_n297_;
  assign new_n299_ = ~new_n288_ & new_n297_;
  assign new_n300_ = pq & new_n297_;
  assign new_n301_ = ~new_n298_ & ~new_n299_;
  assign new_n302_ = ~new_n300_ & new_n301_;
  assign new_n303_ = ~new_n296_ & ~new_n302_;
  assign new_n304_ = ~pn0 & new_n303_;
  assign new_n305_ = new_n293_ & new_n304_;
  assign new_n306_ = pl4 & ~py1;
  assign new_n307_ = new_n304_ & ~new_n306_;
  assign new_n308_ = px1 & new_n303_;
  assign new_n309_ = ~new_n306_ & new_n308_;
  assign new_n310_ = ~pn0 & new_n288_;
  assign new_n311_ = new_n308_ & new_n310_;
  assign new_n312_ = new_n293_ & new_n308_;
  assign new_n313_ = new_n294_ & new_n303_;
  assign new_n314_ = ~new_n306_ & new_n313_;
  assign new_n315_ = new_n310_ & new_n313_;
  assign new_n316_ = new_n304_ & new_n310_;
  assign new_n317_ = new_n293_ & new_n313_;
  assign new_n318_ = ~new_n305_ & ~new_n307_;
  assign new_n319_ = ~new_n309_ & new_n318_;
  assign new_n320_ = ~new_n311_ & ~new_n312_;
  assign new_n321_ = new_n319_ & new_n320_;
  assign new_n322_ = ~new_n316_ & ~new_n317_;
  assign new_n323_ = ~new_n314_ & ~new_n315_;
  assign new_n324_ = new_n322_ & new_n323_;
  assign pg7 = ~new_n321_ | ~new_n324_;
  assign new_n326_ = pl4 & pz2;
  assign new_n327_ = ~pk0 & pl0;
  assign new_n328_ = pk0 & ~pl0;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = new_n288_ & new_n329_;
  assign new_n331_ = ~pm0 & new_n330_;
  assign new_n332_ = ~pn0 & new_n331_;
  assign new_n333_ = py2 & ~new_n332_;
  assign new_n334_ = ~pl4 & new_n333_;
  assign new_n335_ = ~pm0 & ~pn0;
  assign new_n336_ = new_n288_ & new_n335_;
  assign new_n337_ = new_n329_ & new_n336_;
  assign new_n338_ = po & new_n337_;
  assign new_n339_ = ~new_n334_ & ~new_n338_;
  assign new_n340_ = ~new_n326_ & new_n339_;
  assign new_n341_ = ~new_n293_ & new_n340_;
  assign new_n342_ = new_n293_ & new_n339_;
  assign new_n343_ = ~py2 & new_n342_;
  assign new_n344_ = ~py2 & new_n340_;
  assign new_n345_ = ~pl0 & new_n288_;
  assign new_n346_ = ~pk0 & new_n345_;
  assign new_n347_ = pl0 & new_n288_;
  assign new_n348_ = pk0 & new_n347_;
  assign new_n349_ = ~new_n346_ & ~new_n348_;
  assign new_n350_ = ~pm0 & ~new_n349_;
  assign new_n351_ = ~pn0 & new_n350_;
  assign new_n352_ = new_n339_ & new_n351_;
  assign new_n353_ = ~new_n341_ & ~new_n343_;
  assign new_n354_ = ~new_n344_ & ~new_n352_;
  assign new_n355_ = new_n353_ & new_n354_;
  assign new_n356_ = po0 & new_n355_;
  assign ph8 = ~pq0 & new_n356_;
  assign new_n358_ = ~px3 & ~new_n293_;
  assign new_n359_ = py3 & new_n358_;
  assign new_n360_ = ~pz3 & new_n359_;
  assign new_n361_ = pl4 & new_n360_;
  assign new_n362_ = ~pq0 & ~new_n361_;
  assign new_n363_ = pn0 & new_n362_;
  assign new_n364_ = ~new_n288_ & new_n362_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = pl4 & py3;
  assign new_n367_ = ~new_n293_ & new_n366_;
  assign new_n368_ = ~px3 & new_n367_;
  assign new_n369_ = pz3 & ~new_n368_;
  assign new_n370_ = ~new_n365_ & ~new_n369_;
  assign pi9 = ~po0 | ~new_n370_;
  assign pd5 = pm0 & pm3;
  assign new_n373_ = ~pw1 & new_n295_;
  assign new_n374_ = pl0 & new_n297_;
  assign new_n375_ = new_n301_ & ~new_n374_;
  assign new_n376_ = ~new_n373_ & ~new_n375_;
  assign new_n377_ = ~pn0 & new_n376_;
  assign new_n378_ = new_n293_ & new_n377_;
  assign new_n379_ = pl4 & ~px1;
  assign new_n380_ = new_n377_ & ~new_n379_;
  assign new_n381_ = pw1 & new_n376_;
  assign new_n382_ = ~new_n379_ & new_n381_;
  assign new_n383_ = new_n310_ & new_n381_;
  assign new_n384_ = new_n293_ & new_n381_;
  assign new_n385_ = new_n294_ & new_n376_;
  assign new_n386_ = ~new_n379_ & new_n385_;
  assign new_n387_ = new_n310_ & new_n385_;
  assign new_n388_ = new_n310_ & new_n377_;
  assign new_n389_ = new_n293_ & new_n385_;
  assign new_n390_ = ~new_n378_ & ~new_n380_;
  assign new_n391_ = ~new_n382_ & new_n390_;
  assign new_n392_ = ~new_n383_ & ~new_n384_;
  assign new_n393_ = new_n391_ & new_n392_;
  assign new_n394_ = ~new_n388_ & ~new_n389_;
  assign new_n395_ = ~new_n386_ & ~new_n387_;
  assign new_n396_ = new_n394_ & new_n395_;
  assign pf7 = ~new_n393_ | ~new_n396_;
  assign pg6 = ~pl4 | ~pl1;
  assign new_n399_ = ~py3 & new_n358_;
  assign new_n400_ = pl4 & new_n399_;
  assign new_n401_ = ~pq0 & ~new_n400_;
  assign new_n402_ = pn0 & new_n401_;
  assign new_n403_ = ~new_n288_ & new_n401_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = pl4 & new_n358_;
  assign new_n406_ = py3 & ~new_n405_;
  assign new_n407_ = ~new_n404_ & ~new_n406_;
  assign ph9 = ~po0 | ~new_n407_;
  assign new_n409_ = ~pq0 & pz2;
  assign new_n410_ = new_n310_ & new_n329_;
  assign new_n411_ = ~pm0 & new_n410_;
  assign new_n412_ = ~new_n294_ & ~new_n411_;
  assign new_n413_ = new_n409_ & new_n412_;
  assign new_n414_ = po0 & new_n413_;
  assign new_n415_ = new_n288_ & new_n297_;
  assign new_n416_ = pp & ~pm0;
  assign new_n417_ = ~pn0 & new_n416_;
  assign new_n418_ = new_n329_ & new_n415_;
  assign new_n419_ = new_n417_ & new_n418_;
  assign pi8 = new_n414_ | new_n419_;
  assign pd6 = ~pi1 | ~pl4;
  assign new_n422_ = ~pv1 & new_n295_;
  assign new_n423_ = pk0 & new_n297_;
  assign new_n424_ = new_n301_ & ~new_n423_;
  assign new_n425_ = ~new_n422_ & ~new_n424_;
  assign new_n426_ = ~pn0 & new_n425_;
  assign new_n427_ = new_n293_ & new_n426_;
  assign new_n428_ = pl4 & ~pw1;
  assign new_n429_ = new_n426_ & ~new_n428_;
  assign new_n430_ = pv1 & new_n425_;
  assign new_n431_ = ~new_n428_ & new_n430_;
  assign new_n432_ = new_n310_ & new_n430_;
  assign new_n433_ = new_n293_ & new_n430_;
  assign new_n434_ = new_n294_ & new_n425_;
  assign new_n435_ = ~new_n428_ & new_n434_;
  assign new_n436_ = new_n310_ & new_n434_;
  assign new_n437_ = new_n310_ & new_n426_;
  assign new_n438_ = new_n293_ & new_n434_;
  assign new_n439_ = ~new_n427_ & ~new_n429_;
  assign new_n440_ = ~new_n431_ & new_n439_;
  assign new_n441_ = ~new_n432_ & ~new_n433_;
  assign new_n442_ = new_n440_ & new_n441_;
  assign new_n443_ = ~new_n437_ & ~new_n438_;
  assign new_n444_ = ~new_n435_ & ~new_n436_;
  assign new_n445_ = new_n443_ & new_n444_;
  assign pe7 = ~new_n442_ | ~new_n445_;
  assign pg5 = pm0 & pp3;
  assign new_n448_ = pa3 & ~pq0;
  assign new_n449_ = ~pk1 & ~pj1;
  assign new_n450_ = ~pl1 & new_n449_;
  assign new_n451_ = pe4 & pf4;
  assign new_n452_ = ~pg4 & new_n451_;
  assign new_n453_ = ~ph4 & new_n452_;
  assign new_n454_ = pk1 & pj1;
  assign new_n455_ = ph1 & ~px0;
  assign new_n456_ = pi1 & ~py0;
  assign new_n457_ = pb1 & ~pk1;
  assign new_n458_ = ~pj1 & new_n457_;
  assign new_n459_ = pa1 & ~pl1;
  assign new_n460_ = pz0 & new_n459_;
  assign new_n461_ = pa1 & pb1;
  assign new_n462_ = ~pj1 & new_n461_;
  assign new_n463_ = pz0 & new_n457_;
  assign new_n464_ = pz0 & new_n461_;
  assign new_n465_ = ~pk1 & ~pl1;
  assign new_n466_ = ~pj1 & new_n465_;
  assign new_n467_ = ~pj1 & new_n459_;
  assign new_n468_ = pz0 & new_n465_;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = ~new_n464_ & ~new_n466_;
  assign new_n471_ = new_n469_ & new_n470_;
  assign new_n472_ = ~new_n458_ & ~new_n460_;
  assign new_n473_ = ~new_n462_ & ~new_n463_;
  assign new_n474_ = new_n472_ & new_n473_;
  assign new_n475_ = new_n471_ & new_n474_;
  assign new_n476_ = ~new_n455_ & ~new_n456_;
  assign new_n477_ = ~new_n475_ & new_n476_;
  assign new_n478_ = ~new_n288_ & ~new_n454_;
  assign new_n479_ = ~new_n477_ & new_n478_;
  assign new_n480_ = ~new_n453_ & new_n479_;
  assign new_n481_ = ~pj1 & new_n480_;
  assign new_n482_ = ~pl1 & new_n480_;
  assign new_n483_ = ~new_n481_ & ~new_n482_;
  assign new_n484_ = pk1 & pl1;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = pk4 & new_n485_;
  assign new_n487_ = ~pi1 & new_n465_;
  assign new_n488_ = ~pj1 & new_n487_;
  assign new_n489_ = new_n450_ & new_n486_;
  assign new_n490_ = new_n488_ & new_n489_;
  assign new_n491_ = ~pi1 & new_n486_;
  assign new_n492_ = new_n488_ & new_n491_;
  assign new_n493_ = ~ph1 & new_n489_;
  assign new_n494_ = ~ph1 & new_n491_;
  assign new_n495_ = ~new_n490_ & ~new_n492_;
  assign new_n496_ = ~new_n493_ & ~new_n494_;
  assign new_n497_ = new_n495_ & new_n496_;
  assign new_n498_ = new_n448_ & new_n497_;
  assign new_n499_ = po0 & new_n498_;
  assign new_n500_ = pb3 & ~new_n453_;
  assign new_n501_ = pk4 & new_n500_;
  assign new_n502_ = ph1 & ~new_n488_;
  assign new_n503_ = pi1 & ~new_n450_;
  assign new_n504_ = pj1 & pl1;
  assign new_n505_ = ~new_n484_ & ~new_n504_;
  assign new_n506_ = ~new_n454_ & new_n505_;
  assign new_n507_ = ph1 & new_n506_;
  assign new_n508_ = ~new_n450_ & new_n506_;
  assign new_n509_ = pi1 & new_n506_;
  assign new_n510_ = ~new_n507_ & ~new_n508_;
  assign new_n511_ = ~new_n509_ & new_n510_;
  assign new_n512_ = ~new_n502_ & ~new_n503_;
  assign new_n513_ = ~new_n511_ & new_n512_;
  assign new_n514_ = new_n297_ & ~new_n477_;
  assign new_n515_ = new_n501_ & new_n513_;
  assign new_n516_ = new_n514_ & new_n515_;
  assign pj8 = new_n499_ | new_n516_;
  assign new_n518_ = ~pq0 & ~new_n293_;
  assign new_n519_ = ~px3 & new_n518_;
  assign new_n520_ = pz3 & py3;
  assign new_n521_ = ~pa4 & ~pb4;
  assign new_n522_ = pl4 & new_n521_;
  assign new_n523_ = new_n520_ & new_n522_;
  assign new_n524_ = po0 & new_n523_;
  assign new_n525_ = ~new_n310_ & new_n519_;
  assign new_n526_ = new_n524_ & new_n525_;
  assign new_n527_ = pb4 & ~pq0;
  assign new_n528_ = py3 & ~px3;
  assign new_n529_ = pl4 & new_n289_;
  assign new_n530_ = new_n528_ & new_n529_;
  assign new_n531_ = ~new_n293_ & new_n530_;
  assign new_n532_ = ~new_n310_ & ~new_n531_;
  assign new_n533_ = new_n527_ & new_n532_;
  assign new_n534_ = po0 & new_n533_;
  assign new_n535_ = pm0 & ~pn0;
  assign new_n536_ = po0 & new_n535_;
  assign new_n537_ = ~pq0 & new_n536_;
  assign new_n538_ = new_n288_ & new_n537_;
  assign new_n539_ = ~new_n526_ & ~new_n534_;
  assign pk9 = new_n538_ | ~new_n539_;
  assign new_n541_ = ~pu1 & new_n295_;
  assign new_n542_ = pm0 & new_n297_;
  assign new_n543_ = new_n301_ & ~new_n542_;
  assign new_n544_ = ~new_n541_ & ~new_n543_;
  assign new_n545_ = ~pn0 & new_n544_;
  assign new_n546_ = new_n293_ & new_n545_;
  assign new_n547_ = pl4 & ~pv1;
  assign new_n548_ = new_n545_ & ~new_n547_;
  assign new_n549_ = pu1 & new_n544_;
  assign new_n550_ = ~new_n547_ & new_n549_;
  assign new_n551_ = new_n310_ & new_n549_;
  assign new_n552_ = new_n293_ & new_n549_;
  assign new_n553_ = new_n294_ & new_n544_;
  assign new_n554_ = ~new_n547_ & new_n553_;
  assign new_n555_ = new_n310_ & new_n553_;
  assign new_n556_ = new_n310_ & new_n545_;
  assign new_n557_ = new_n293_ & new_n553_;
  assign new_n558_ = ~new_n546_ & ~new_n548_;
  assign new_n559_ = ~new_n550_ & new_n558_;
  assign new_n560_ = ~new_n551_ & ~new_n552_;
  assign new_n561_ = new_n559_ & new_n560_;
  assign new_n562_ = ~new_n556_ & ~new_n557_;
  assign new_n563_ = ~new_n554_ & ~new_n555_;
  assign new_n564_ = new_n562_ & new_n563_;
  assign pd7 = ~new_n561_ | ~new_n564_;
  assign pe6 = ~pl4 | ~pj1;
  assign pf5 = po3 & pm0;
  assign new_n568_ = pl4 & new_n520_;
  assign new_n569_ = new_n358_ & new_n568_;
  assign new_n570_ = ~new_n288_ & new_n569_;
  assign new_n571_ = pn0 & new_n288_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = new_n329_ & new_n572_;
  assign new_n574_ = pa4 & new_n573_;
  assign new_n575_ = new_n288_ & new_n573_;
  assign new_n576_ = new_n288_ & new_n572_;
  assign new_n577_ = pm0 & new_n576_;
  assign new_n578_ = ~new_n288_ & new_n572_;
  assign new_n579_ = pa4 & new_n578_;
  assign new_n580_ = pa4 & new_n572_;
  assign new_n581_ = pm0 & new_n580_;
  assign new_n582_ = ~new_n574_ & ~new_n575_;
  assign new_n583_ = ~new_n577_ & new_n582_;
  assign new_n584_ = ~new_n579_ & ~new_n581_;
  assign new_n585_ = new_n583_ & new_n584_;
  assign new_n586_ = ~pn0 & new_n585_;
  assign new_n587_ = ~new_n359_ & new_n586_;
  assign new_n588_ = ~new_n529_ & new_n586_;
  assign new_n589_ = ~pa4 & new_n585_;
  assign new_n590_ = ~new_n529_ & new_n589_;
  assign new_n591_ = new_n310_ & new_n589_;
  assign new_n592_ = ~new_n359_ & new_n589_;
  assign new_n593_ = ~new_n293_ & new_n568_;
  assign new_n594_ = ~px3 & new_n593_;
  assign new_n595_ = new_n585_ & new_n594_;
  assign new_n596_ = ~new_n529_ & new_n595_;
  assign new_n597_ = new_n310_ & new_n595_;
  assign new_n598_ = new_n310_ & new_n586_;
  assign new_n599_ = ~new_n359_ & new_n595_;
  assign new_n600_ = ~new_n587_ & ~new_n588_;
  assign new_n601_ = ~new_n590_ & new_n600_;
  assign new_n602_ = ~new_n591_ & ~new_n592_;
  assign new_n603_ = new_n601_ & new_n602_;
  assign new_n604_ = ~new_n598_ & ~new_n599_;
  assign new_n605_ = ~new_n596_ & ~new_n597_;
  assign new_n606_ = new_n604_ & new_n605_;
  assign new_n607_ = new_n603_ & new_n606_;
  assign new_n608_ = po0 & new_n607_;
  assign pj9 = ~pq0 & new_n608_;
  assign new_n610_ = pb3 & ~pq0;
  assign new_n611_ = new_n497_ & new_n610_;
  assign new_n612_ = po0 & new_n611_;
  assign new_n613_ = pc3 & ~new_n453_;
  assign new_n614_ = pk4 & new_n613_;
  assign new_n615_ = new_n513_ & new_n614_;
  assign new_n616_ = new_n514_ & new_n615_;
  assign pk8 = new_n612_ | new_n616_;
  assign new_n618_ = ~pj3 & pl0;
  assign new_n619_ = pk0 & new_n618_;
  assign new_n620_ = ~pj3 & ~pl0;
  assign new_n621_ = ~pk0 & new_n620_;
  assign new_n622_ = ~new_n619_ & ~new_n621_;
  assign new_n623_ = pm0 & new_n622_;
  assign new_n624_ = pl0 & new_n623_;
  assign new_n625_ = pk0 & new_n624_;
  assign new_n626_ = ~pl0 & new_n623_;
  assign new_n627_ = ~pk0 & new_n626_;
  assign new_n628_ = pr3 & new_n623_;
  assign new_n629_ = ~new_n625_ & ~new_n627_;
  assign pa5 = new_n628_ | ~new_n629_;
  assign new_n631_ = pm1 & pl1;
  assign pb6 = pk4 | ~new_n631_;
  assign new_n633_ = ~pt1 & new_n295_;
  assign new_n634_ = pd0 & new_n297_;
  assign new_n635_ = new_n301_ & ~new_n634_;
  assign new_n636_ = ~new_n633_ & ~new_n635_;
  assign new_n637_ = ~pn0 & new_n636_;
  assign new_n638_ = new_n293_ & new_n637_;
  assign new_n639_ = pl4 & ~pu1;
  assign new_n640_ = new_n637_ & ~new_n639_;
  assign new_n641_ = pt1 & new_n636_;
  assign new_n642_ = ~new_n639_ & new_n641_;
  assign new_n643_ = new_n310_ & new_n641_;
  assign new_n644_ = new_n293_ & new_n641_;
  assign new_n645_ = new_n294_ & new_n636_;
  assign new_n646_ = ~new_n639_ & new_n645_;
  assign new_n647_ = new_n310_ & new_n645_;
  assign new_n648_ = new_n310_ & new_n637_;
  assign new_n649_ = new_n293_ & new_n645_;
  assign new_n650_ = ~new_n638_ & ~new_n640_;
  assign new_n651_ = ~new_n642_ & new_n650_;
  assign new_n652_ = ~new_n643_ & ~new_n644_;
  assign new_n653_ = new_n651_ & new_n652_;
  assign new_n654_ = ~new_n648_ & ~new_n649_;
  assign new_n655_ = ~new_n646_ & ~new_n647_;
  assign new_n656_ = new_n654_ & new_n655_;
  assign pc7 = ~new_n653_ | ~new_n656_;
  assign new_n658_ = pc3 & ~pq0;
  assign new_n659_ = new_n497_ & new_n658_;
  assign new_n660_ = po0 & new_n659_;
  assign new_n661_ = pd3 & ~new_n453_;
  assign new_n662_ = pk4 & new_n661_;
  assign new_n663_ = new_n513_ & new_n662_;
  assign new_n664_ = new_n514_ & new_n663_;
  assign pl8 = new_n660_ | new_n664_;
  assign new_n666_ = ~pq0 & new_n288_;
  assign new_n667_ = po0 & new_n666_;
  assign new_n668_ = ~pn0 & new_n667_;
  assign new_n669_ = ~pg1 & ~pq0;
  assign new_n670_ = pd4 & pk4;
  assign new_n671_ = ~new_n477_ & new_n670_;
  assign new_n672_ = ~new_n453_ & new_n671_;
  assign new_n673_ = ~new_n453_ & ~new_n477_;
  assign new_n674_ = pk4 & new_n673_;
  assign new_n675_ = ~pd4 & ~new_n674_;
  assign new_n676_ = ~new_n672_ & ~new_n675_;
  assign new_n677_ = new_n669_ & new_n676_;
  assign new_n678_ = po0 & new_n677_;
  assign pm9 = new_n668_ | new_n678_;
  assign new_n680_ = ~ps1 & new_n295_;
  assign new_n681_ = pe0 & new_n297_;
  assign new_n682_ = new_n301_ & ~new_n681_;
  assign new_n683_ = ~new_n680_ & ~new_n682_;
  assign new_n684_ = ~pn0 & new_n683_;
  assign new_n685_ = new_n293_ & new_n684_;
  assign new_n686_ = pl4 & ~pt1;
  assign new_n687_ = new_n684_ & ~new_n686_;
  assign new_n688_ = ps1 & new_n683_;
  assign new_n689_ = ~new_n686_ & new_n688_;
  assign new_n690_ = new_n310_ & new_n688_;
  assign new_n691_ = new_n293_ & new_n688_;
  assign new_n692_ = new_n294_ & new_n683_;
  assign new_n693_ = ~new_n686_ & new_n692_;
  assign new_n694_ = new_n310_ & new_n692_;
  assign new_n695_ = new_n310_ & new_n684_;
  assign new_n696_ = new_n293_ & new_n692_;
  assign new_n697_ = ~new_n685_ & ~new_n687_;
  assign new_n698_ = ~new_n689_ & new_n697_;
  assign new_n699_ = ~new_n690_ & ~new_n691_;
  assign new_n700_ = new_n698_ & new_n699_;
  assign new_n701_ = ~new_n695_ & ~new_n696_;
  assign new_n702_ = ~new_n693_ & ~new_n694_;
  assign new_n703_ = new_n701_ & new_n702_;
  assign pb7 = ~new_n700_ | ~new_n703_;
  assign pc6 = ~pl4 | ~ph1;
  assign new_n706_ = ~pa4 & new_n520_;
  assign new_n707_ = ~pb4 & ~pc4;
  assign new_n708_ = pl4 & new_n707_;
  assign new_n709_ = new_n706_ & new_n708_;
  assign new_n710_ = po0 & new_n709_;
  assign new_n711_ = new_n525_ & new_n710_;
  assign new_n712_ = pc4 & ~pq0;
  assign new_n713_ = pz3 & new_n528_;
  assign new_n714_ = new_n522_ & new_n713_;
  assign new_n715_ = ~new_n293_ & new_n714_;
  assign new_n716_ = ~new_n310_ & ~new_n715_;
  assign new_n717_ = new_n712_ & new_n716_;
  assign new_n718_ = po0 & new_n717_;
  assign new_n719_ = po0 & new_n335_;
  assign new_n720_ = ~pq0 & new_n719_;
  assign new_n721_ = new_n288_ & new_n720_;
  assign new_n722_ = ~new_n711_ & ~new_n718_;
  assign pl9 = new_n721_ | ~new_n722_;
  assign new_n724_ = pd3 & ~pq0;
  assign new_n725_ = new_n497_ & new_n724_;
  assign new_n726_ = po0 & new_n725_;
  assign new_n727_ = pe3 & ~new_n453_;
  assign new_n728_ = pk4 & new_n727_;
  assign new_n729_ = new_n513_ & new_n728_;
  assign new_n730_ = new_n514_ & new_n729_;
  assign pm8 = new_n726_ | new_n730_;
  assign new_n732_ = ~pr1 & new_n295_;
  assign new_n733_ = pf0 & new_n297_;
  assign new_n734_ = new_n301_ & ~new_n733_;
  assign new_n735_ = ~new_n732_ & ~new_n734_;
  assign new_n736_ = ~pn0 & new_n735_;
  assign new_n737_ = new_n293_ & new_n736_;
  assign new_n738_ = pl4 & ~ps1;
  assign new_n739_ = new_n736_ & ~new_n738_;
  assign new_n740_ = pr1 & new_n735_;
  assign new_n741_ = ~new_n738_ & new_n740_;
  assign new_n742_ = new_n310_ & new_n740_;
  assign new_n743_ = new_n293_ & new_n740_;
  assign new_n744_ = new_n294_ & new_n735_;
  assign new_n745_ = ~new_n738_ & new_n744_;
  assign new_n746_ = new_n310_ & new_n744_;
  assign new_n747_ = new_n310_ & new_n736_;
  assign new_n748_ = new_n293_ & new_n744_;
  assign new_n749_ = ~new_n737_ & ~new_n739_;
  assign new_n750_ = ~new_n741_ & new_n749_;
  assign new_n751_ = ~new_n742_ & ~new_n743_;
  assign new_n752_ = new_n750_ & new_n751_;
  assign new_n753_ = ~new_n747_ & ~new_n748_;
  assign new_n754_ = ~new_n745_ & ~new_n746_;
  assign new_n755_ = new_n753_ & new_n754_;
  assign pa7 = ~new_n752_ | ~new_n755_;
  assign new_n757_ = pl0 & ~pl3;
  assign new_n758_ = pk0 & new_n757_;
  assign new_n759_ = ~pl0 & ~pl3;
  assign new_n760_ = ~pk0 & new_n759_;
  assign new_n761_ = ~new_n758_ & ~new_n760_;
  assign new_n762_ = pm0 & new_n761_;
  assign new_n763_ = pl0 & new_n762_;
  assign new_n764_ = pk0 & new_n763_;
  assign new_n765_ = ~pl0 & new_n762_;
  assign new_n766_ = ~pk0 & new_n765_;
  assign new_n767_ = pt3 & new_n762_;
  assign new_n768_ = ~new_n764_ & ~new_n766_;
  assign pc5 = new_n767_ | ~new_n768_;
  assign new_n770_ = pe3 & ~pq0;
  assign new_n771_ = new_n497_ & new_n770_;
  assign new_n772_ = po0 & new_n771_;
  assign new_n773_ = pf3 & ~new_n453_;
  assign new_n774_ = pk4 & new_n773_;
  assign new_n775_ = new_n513_ & new_n774_;
  assign new_n776_ = new_n514_ & new_n775_;
  assign pn8 = new_n772_ | new_n776_;
  assign new_n778_ = ~pd4 & ~new_n453_;
  assign new_n779_ = pe4 & ~pf4;
  assign new_n780_ = pk4 & new_n779_;
  assign new_n781_ = new_n778_ & new_n780_;
  assign new_n782_ = ~new_n477_ & new_n781_;
  assign new_n783_ = ~new_n310_ & ~new_n782_;
  assign new_n784_ = ~pg1 & new_n783_;
  assign new_n785_ = ~pq0 & new_n784_;
  assign new_n786_ = ~pd4 & pe4;
  assign new_n787_ = pk4 & new_n786_;
  assign new_n788_ = ~new_n477_ & new_n787_;
  assign new_n789_ = ~new_n453_ & new_n788_;
  assign new_n790_ = pf4 & ~new_n789_;
  assign new_n791_ = new_n785_ & ~new_n790_;
  assign po9 = ~po0 | ~new_n791_;
  assign new_n793_ = pk1 & pm1;
  assign pa6 = pk4 | ~new_n793_;
  assign new_n795_ = ~pk3 & pl0;
  assign new_n796_ = pk0 & new_n795_;
  assign new_n797_ = ~pk3 & ~pl0;
  assign new_n798_ = ~pk0 & new_n797_;
  assign new_n799_ = ~new_n796_ & ~new_n798_;
  assign new_n800_ = pm0 & new_n799_;
  assign new_n801_ = pl0 & new_n800_;
  assign new_n802_ = pk0 & new_n801_;
  assign new_n803_ = ~pl0 & new_n800_;
  assign new_n804_ = ~pk0 & new_n803_;
  assign new_n805_ = ps3 & new_n800_;
  assign new_n806_ = ~new_n802_ & ~new_n804_;
  assign pb5 = new_n805_ | ~new_n806_;
  assign new_n808_ = ~pd4 & ~pe4;
  assign new_n809_ = pk4 & new_n808_;
  assign new_n810_ = ~new_n477_ & new_n809_;
  assign new_n811_ = ~new_n453_ & new_n810_;
  assign new_n812_ = ~new_n310_ & ~new_n811_;
  assign new_n813_ = ~pg1 & new_n812_;
  assign new_n814_ = ~pq0 & new_n813_;
  assign new_n815_ = ~pd4 & pk4;
  assign new_n816_ = ~new_n477_ & new_n815_;
  assign new_n817_ = ~new_n453_ & new_n816_;
  assign new_n818_ = pe4 & ~new_n817_;
  assign new_n819_ = new_n814_ & ~new_n818_;
  assign pn9 = ~po0 | ~new_n819_;
  assign new_n821_ = pf3 & ~pq0;
  assign new_n822_ = new_n497_ & new_n821_;
  assign new_n823_ = po0 & new_n822_;
  assign new_n824_ = pg3 & ~new_n453_;
  assign new_n825_ = pk4 & new_n824_;
  assign new_n826_ = new_n513_ & new_n825_;
  assign new_n827_ = new_n514_ & new_n826_;
  assign po8 = new_n823_ | new_n827_;
  assign new_n829_ = ~pq0 & pr3;
  assign new_n830_ = new_n497_ & new_n829_;
  assign new_n831_ = po0 & new_n830_;
  assign new_n832_ = ps3 & ~new_n453_;
  assign new_n833_ = pk4 & new_n832_;
  assign new_n834_ = new_n513_ & new_n833_;
  assign new_n835_ = new_n514_ & new_n834_;
  assign pa9 = new_n831_ | new_n835_;
  assign new_n837_ = ~pf1 & ~pi4;
  assign new_n838_ = pf1 & pi4;
  assign pn6 = new_n837_ | new_n838_;
  assign new_n840_ = ~pf2 & new_n295_;
  assign new_n841_ = py & new_n297_;
  assign new_n842_ = new_n301_ & ~new_n841_;
  assign new_n843_ = ~new_n840_ & ~new_n842_;
  assign new_n844_ = ~pn0 & new_n843_;
  assign new_n845_ = new_n293_ & new_n844_;
  assign new_n846_ = ~pg2 & pl4;
  assign new_n847_ = new_n844_ & ~new_n846_;
  assign new_n848_ = pf2 & new_n843_;
  assign new_n849_ = ~new_n846_ & new_n848_;
  assign new_n850_ = new_n310_ & new_n848_;
  assign new_n851_ = new_n293_ & new_n848_;
  assign new_n852_ = new_n294_ & new_n843_;
  assign new_n853_ = ~new_n846_ & new_n852_;
  assign new_n854_ = new_n310_ & new_n852_;
  assign new_n855_ = new_n310_ & new_n844_;
  assign new_n856_ = new_n293_ & new_n852_;
  assign new_n857_ = ~new_n845_ & ~new_n847_;
  assign new_n858_ = ~new_n849_ & new_n857_;
  assign new_n859_ = ~new_n850_ & ~new_n851_;
  assign new_n860_ = new_n858_ & new_n859_;
  assign new_n861_ = ~new_n855_ & ~new_n856_;
  assign new_n862_ = ~new_n853_ & ~new_n854_;
  assign new_n863_ = new_n861_ & new_n862_;
  assign po7 = ~new_n860_ | ~new_n863_;
  assign new_n865_ = pl0 & ph;
  assign new_n866_ = pp & ~pl0;
  assign new_n867_ = pk0 & new_n866_;
  assign new_n868_ = ~pk0 & ph;
  assign new_n869_ = ~new_n865_ & ~new_n867_;
  assign new_n870_ = ~new_n868_ & new_n869_;
  assign new_n871_ = new_n310_ & new_n870_;
  assign new_n872_ = ~pm0 & new_n871_;
  assign new_n873_ = pl4 & ~ps2;
  assign new_n874_ = ~new_n336_ & new_n873_;
  assign new_n875_ = ~new_n293_ & new_n874_;
  assign new_n876_ = ~pm0 & new_n310_;
  assign new_n877_ = ~new_n294_ & ~new_n876_;
  assign new_n878_ = ~pr2 & new_n877_;
  assign new_n879_ = ~new_n872_ & ~new_n875_;
  assign new_n880_ = ~new_n878_ & new_n879_;
  assign new_n881_ = po0 & new_n880_;
  assign pa8 = ~pq0 & new_n881_;
  assign pl5 = pg1 & ~pj4;
  assign new_n884_ = ~pe2 & new_n295_;
  assign new_n885_ = px & new_n297_;
  assign new_n886_ = new_n301_ & ~new_n885_;
  assign new_n887_ = ~new_n884_ & ~new_n886_;
  assign new_n888_ = ~pn0 & new_n887_;
  assign new_n889_ = new_n293_ & new_n888_;
  assign new_n890_ = ~pf2 & pl4;
  assign new_n891_ = new_n888_ & ~new_n890_;
  assign new_n892_ = pe2 & new_n887_;
  assign new_n893_ = ~new_n890_ & new_n892_;
  assign new_n894_ = new_n310_ & new_n892_;
  assign new_n895_ = new_n293_ & new_n892_;
  assign new_n896_ = new_n294_ & new_n887_;
  assign new_n897_ = ~new_n890_ & new_n896_;
  assign new_n898_ = new_n310_ & new_n896_;
  assign new_n899_ = new_n310_ & new_n888_;
  assign new_n900_ = new_n293_ & new_n896_;
  assign new_n901_ = ~new_n889_ & ~new_n891_;
  assign new_n902_ = ~new_n893_ & new_n901_;
  assign new_n903_ = ~new_n894_ & ~new_n895_;
  assign new_n904_ = new_n902_ & new_n903_;
  assign new_n905_ = ~new_n899_ & ~new_n900_;
  assign new_n906_ = ~new_n897_ & ~new_n898_;
  assign new_n907_ = new_n905_ & new_n906_;
  assign pn7 = ~new_n904_ | ~new_n907_;
  assign new_n909_ = px3 & new_n289_;
  assign new_n910_ = py3 & new_n909_;
  assign new_n911_ = ~pb4 & new_n910_;
  assign po6 = ~pc4 & new_n911_;
  assign new_n913_ = pl4 & pt2;
  assign new_n914_ = ps2 & ~new_n332_;
  assign new_n915_ = ~pl4 & new_n914_;
  assign new_n916_ = pi & new_n337_;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = ~new_n913_ & new_n917_;
  assign new_n919_ = ~new_n293_ & new_n918_;
  assign new_n920_ = new_n293_ & new_n917_;
  assign new_n921_ = ~ps2 & new_n920_;
  assign new_n922_ = ~ps2 & new_n918_;
  assign new_n923_ = new_n351_ & new_n917_;
  assign new_n924_ = ~new_n919_ & ~new_n921_;
  assign new_n925_ = ~new_n922_ & ~new_n923_;
  assign new_n926_ = new_n924_ & new_n925_;
  assign new_n927_ = po0 & new_n926_;
  assign pb8 = ~pq0 & new_n927_;
  assign new_n929_ = ~pq0 & pt3;
  assign new_n930_ = new_n497_ & new_n929_;
  assign new_n931_ = po0 & new_n930_;
  assign new_n932_ = pu3 & ~new_n453_;
  assign new_n933_ = pk4 & new_n932_;
  assign new_n934_ = new_n513_ & new_n933_;
  assign new_n935_ = new_n514_ & new_n934_;
  assign pc9 = new_n931_ | new_n935_;
  assign new_n937_ = ~pd2 & new_n295_;
  assign new_n938_ = pw & new_n297_;
  assign new_n939_ = new_n301_ & ~new_n938_;
  assign new_n940_ = ~new_n937_ & ~new_n939_;
  assign new_n941_ = ~pn0 & new_n940_;
  assign new_n942_ = new_n293_ & new_n941_;
  assign new_n943_ = ~pe2 & pl4;
  assign new_n944_ = new_n941_ & ~new_n943_;
  assign new_n945_ = pd2 & new_n940_;
  assign new_n946_ = ~new_n943_ & new_n945_;
  assign new_n947_ = new_n310_ & new_n945_;
  assign new_n948_ = new_n293_ & new_n945_;
  assign new_n949_ = new_n294_ & new_n940_;
  assign new_n950_ = ~new_n943_ & new_n949_;
  assign new_n951_ = new_n310_ & new_n949_;
  assign new_n952_ = new_n310_ & new_n941_;
  assign new_n953_ = new_n293_ & new_n949_;
  assign new_n954_ = ~new_n942_ & ~new_n944_;
  assign new_n955_ = ~new_n946_ & new_n954_;
  assign new_n956_ = ~new_n947_ & ~new_n948_;
  assign new_n957_ = new_n955_ & new_n956_;
  assign new_n958_ = ~new_n952_ & ~new_n953_;
  assign new_n959_ = ~new_n950_ & ~new_n951_;
  assign new_n960_ = new_n958_ & new_n959_;
  assign pm7 = ~new_n957_ | ~new_n960_;
  assign new_n962_ = pi1 & ~pn0;
  assign po5 = pk4 | ~new_n962_;
  assign new_n964_ = ps3 & ~pq0;
  assign new_n965_ = new_n497_ & new_n964_;
  assign new_n966_ = po0 & new_n965_;
  assign new_n967_ = pt3 & ~new_n453_;
  assign new_n968_ = pk4 & new_n967_;
  assign new_n969_ = new_n513_ & new_n968_;
  assign new_n970_ = new_n514_ & new_n969_;
  assign pb9 = new_n966_ | new_n970_;
  assign new_n972_ = pl4 & pu2;
  assign new_n973_ = pt2 & ~new_n332_;
  assign new_n974_ = ~pl4 & new_n973_;
  assign new_n975_ = pj & new_n337_;
  assign new_n976_ = ~new_n974_ & ~new_n975_;
  assign new_n977_ = ~new_n972_ & new_n976_;
  assign new_n978_ = ~new_n293_ & new_n977_;
  assign new_n979_ = new_n293_ & new_n976_;
  assign new_n980_ = ~pt2 & new_n979_;
  assign new_n981_ = ~pt2 & new_n977_;
  assign new_n982_ = new_n351_ & new_n976_;
  assign new_n983_ = ~new_n978_ & ~new_n980_;
  assign new_n984_ = ~new_n981_ & ~new_n982_;
  assign new_n985_ = new_n983_ & new_n984_;
  assign new_n986_ = po0 & new_n985_;
  assign pc8 = ~pq0 & new_n986_;
  assign new_n988_ = ~pc2 & new_n295_;
  assign new_n989_ = pv & new_n297_;
  assign new_n990_ = new_n301_ & ~new_n989_;
  assign new_n991_ = ~new_n988_ & ~new_n990_;
  assign new_n992_ = ~pn0 & new_n991_;
  assign new_n993_ = new_n293_ & new_n992_;
  assign new_n994_ = ~pd2 & pl4;
  assign new_n995_ = new_n992_ & ~new_n994_;
  assign new_n996_ = pc2 & new_n991_;
  assign new_n997_ = ~new_n994_ & new_n996_;
  assign new_n998_ = new_n310_ & new_n996_;
  assign new_n999_ = new_n293_ & new_n996_;
  assign new_n1000_ = new_n294_ & new_n991_;
  assign new_n1001_ = ~new_n994_ & new_n1000_;
  assign new_n1002_ = new_n310_ & new_n1000_;
  assign new_n1003_ = new_n310_ & new_n992_;
  assign new_n1004_ = new_n293_ & new_n1000_;
  assign new_n1005_ = ~new_n993_ & ~new_n995_;
  assign new_n1006_ = ~new_n997_ & new_n1005_;
  assign new_n1007_ = ~new_n998_ & ~new_n999_;
  assign new_n1008_ = new_n1006_ & new_n1007_;
  assign new_n1009_ = ~new_n1003_ & ~new_n1004_;
  assign new_n1010_ = ~new_n1001_ & ~new_n1002_;
  assign new_n1011_ = new_n1009_ & new_n1010_;
  assign pl7 = ~new_n1008_ | ~new_n1011_;
  assign new_n1013_ = ph1 & ~pn0;
  assign pn5 = pk4 | ~new_n1013_;
  assign new_n1015_ = pl4 & pv2;
  assign new_n1016_ = pu2 & ~new_n332_;
  assign new_n1017_ = ~pl4 & new_n1016_;
  assign new_n1018_ = pk & new_n337_;
  assign new_n1019_ = ~new_n1017_ & ~new_n1018_;
  assign new_n1020_ = ~new_n1015_ & new_n1019_;
  assign new_n1021_ = ~new_n293_ & new_n1020_;
  assign new_n1022_ = new_n293_ & new_n1019_;
  assign new_n1023_ = ~pu2 & new_n1022_;
  assign new_n1024_ = ~pu2 & new_n1020_;
  assign new_n1025_ = new_n351_ & new_n1019_;
  assign new_n1026_ = ~new_n1021_ & ~new_n1023_;
  assign new_n1027_ = ~new_n1024_ & ~new_n1025_;
  assign new_n1028_ = new_n1026_ & new_n1027_;
  assign new_n1029_ = po0 & new_n1028_;
  assign pd8 = ~pq0 & new_n1029_;
  assign new_n1031_ = ~pq0 & pv3;
  assign new_n1032_ = new_n497_ & new_n1031_;
  assign new_n1033_ = po0 & new_n1032_;
  assign new_n1034_ = pw3 & ~new_n453_;
  assign new_n1035_ = pk4 & new_n1034_;
  assign new_n1036_ = new_n513_ & new_n1035_;
  assign new_n1037_ = new_n514_ & new_n1036_;
  assign pe9 = new_n1033_ | new_n1037_;
  assign pi5 = pm0 & pr3;
  assign new_n1040_ = ~pb2 & new_n295_;
  assign new_n1041_ = pu & new_n297_;
  assign new_n1042_ = new_n301_ & ~new_n1041_;
  assign new_n1043_ = ~new_n1040_ & ~new_n1042_;
  assign new_n1044_ = ~pn0 & new_n1043_;
  assign new_n1045_ = new_n293_ & new_n1044_;
  assign new_n1046_ = ~pc2 & pl4;
  assign new_n1047_ = new_n1044_ & ~new_n1046_;
  assign new_n1048_ = pb2 & new_n1043_;
  assign new_n1049_ = ~new_n1046_ & new_n1048_;
  assign new_n1050_ = new_n310_ & new_n1048_;
  assign new_n1051_ = new_n293_ & new_n1048_;
  assign new_n1052_ = new_n294_ & new_n1043_;
  assign new_n1053_ = ~new_n1046_ & new_n1052_;
  assign new_n1054_ = new_n310_ & new_n1052_;
  assign new_n1055_ = new_n310_ & new_n1044_;
  assign new_n1056_ = new_n293_ & new_n1052_;
  assign new_n1057_ = ~new_n1045_ & ~new_n1047_;
  assign new_n1058_ = ~new_n1049_ & new_n1057_;
  assign new_n1059_ = ~new_n1050_ & ~new_n1051_;
  assign new_n1060_ = new_n1058_ & new_n1059_;
  assign new_n1061_ = ~new_n1055_ & ~new_n1056_;
  assign new_n1062_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1063_ = new_n1061_ & new_n1062_;
  assign pk7 = ~new_n1060_ | ~new_n1063_;
  assign new_n1065_ = ~pq0 & pu3;
  assign new_n1066_ = new_n497_ & new_n1065_;
  assign new_n1067_ = po0 & new_n1066_;
  assign new_n1068_ = pv3 & ~new_n453_;
  assign new_n1069_ = pk4 & new_n1068_;
  assign new_n1070_ = new_n513_ & new_n1069_;
  assign new_n1071_ = new_n514_ & new_n1070_;
  assign pd9 = new_n1067_ | new_n1071_;
  assign new_n1073_ = pl4 & pw2;
  assign new_n1074_ = pv2 & ~new_n332_;
  assign new_n1075_ = ~pl4 & new_n1074_;
  assign new_n1076_ = pl & new_n337_;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1073_ & new_n1077_;
  assign new_n1079_ = ~new_n293_ & new_n1078_;
  assign new_n1080_ = new_n293_ & new_n1077_;
  assign new_n1081_ = ~pv2 & new_n1080_;
  assign new_n1082_ = ~pv2 & new_n1078_;
  assign new_n1083_ = new_n351_ & new_n1077_;
  assign new_n1084_ = ~new_n1079_ & ~new_n1081_;
  assign new_n1085_ = ~new_n1082_ & ~new_n1083_;
  assign new_n1086_ = new_n1084_ & new_n1085_;
  assign new_n1087_ = po0 & new_n1086_;
  assign pe8 = ~pq0 & new_n1087_;
  assign ph5 = pm0 & pq3;
  assign new_n1090_ = ~pa2 & new_n295_;
  assign new_n1091_ = pt & new_n297_;
  assign new_n1092_ = new_n301_ & ~new_n1091_;
  assign new_n1093_ = ~new_n1090_ & ~new_n1092_;
  assign new_n1094_ = ~pn0 & new_n1093_;
  assign new_n1095_ = new_n293_ & new_n1094_;
  assign new_n1096_ = ~pb2 & pl4;
  assign new_n1097_ = new_n1094_ & ~new_n1096_;
  assign new_n1098_ = pa2 & new_n1093_;
  assign new_n1099_ = ~new_n1096_ & new_n1098_;
  assign new_n1100_ = new_n310_ & new_n1098_;
  assign new_n1101_ = new_n293_ & new_n1098_;
  assign new_n1102_ = new_n294_ & new_n1093_;
  assign new_n1103_ = ~new_n1096_ & new_n1102_;
  assign new_n1104_ = new_n310_ & new_n1102_;
  assign new_n1105_ = new_n310_ & new_n1094_;
  assign new_n1106_ = new_n293_ & new_n1102_;
  assign new_n1107_ = ~new_n1095_ & ~new_n1097_;
  assign new_n1108_ = ~new_n1099_ & new_n1107_;
  assign new_n1109_ = ~new_n1100_ & ~new_n1101_;
  assign new_n1110_ = new_n1108_ & new_n1109_;
  assign new_n1111_ = ~new_n1105_ & ~new_n1106_;
  assign new_n1112_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1113_ = new_n1111_ & new_n1112_;
  assign pj7 = ~new_n1110_ | ~new_n1113_;
  assign new_n1115_ = pl4 & px2;
  assign new_n1116_ = pw2 & ~new_n332_;
  assign new_n1117_ = ~pl4 & new_n1116_;
  assign new_n1118_ = pm & new_n337_;
  assign new_n1119_ = ~new_n1117_ & ~new_n1118_;
  assign new_n1120_ = ~new_n1115_ & new_n1119_;
  assign new_n1121_ = ~new_n293_ & new_n1120_;
  assign new_n1122_ = new_n293_ & new_n1119_;
  assign new_n1123_ = ~pw2 & new_n1122_;
  assign new_n1124_ = ~pw2 & new_n1120_;
  assign new_n1125_ = new_n351_ & new_n1119_;
  assign new_n1126_ = ~new_n1121_ & ~new_n1123_;
  assign new_n1127_ = ~new_n1124_ & ~new_n1125_;
  assign new_n1128_ = new_n1126_ & new_n1127_;
  assign new_n1129_ = po0 & new_n1128_;
  assign pf8 = ~pq0 & new_n1129_;
  assign new_n1131_ = px3 & ~new_n293_;
  assign new_n1132_ = pl4 & new_n1131_;
  assign new_n1133_ = ~new_n301_ & ~new_n1132_;
  assign new_n1134_ = ~new_n293_ & new_n1133_;
  assign new_n1135_ = pl4 & new_n1134_;
  assign new_n1136_ = px3 & new_n1133_;
  assign pg9 = new_n1135_ | new_n1136_;
  assign new_n1138_ = ~pz1 & new_n295_;
  assign new_n1139_ = ps & new_n297_;
  assign new_n1140_ = new_n301_ & ~new_n1139_;
  assign new_n1141_ = ~new_n1138_ & ~new_n1140_;
  assign new_n1142_ = ~pn0 & new_n1141_;
  assign new_n1143_ = new_n293_ & new_n1142_;
  assign new_n1144_ = ~pa2 & pl4;
  assign new_n1145_ = new_n1142_ & ~new_n1144_;
  assign new_n1146_ = pz1 & new_n1141_;
  assign new_n1147_ = ~new_n1144_ & new_n1146_;
  assign new_n1148_ = new_n310_ & new_n1146_;
  assign new_n1149_ = new_n293_ & new_n1146_;
  assign new_n1150_ = new_n294_ & new_n1141_;
  assign new_n1151_ = ~new_n1144_ & new_n1150_;
  assign new_n1152_ = new_n310_ & new_n1150_;
  assign new_n1153_ = new_n310_ & new_n1142_;
  assign new_n1154_ = new_n293_ & new_n1150_;
  assign new_n1155_ = ~new_n1143_ & ~new_n1145_;
  assign new_n1156_ = ~new_n1147_ & new_n1155_;
  assign new_n1157_ = ~new_n1148_ & ~new_n1149_;
  assign new_n1158_ = new_n1156_ & new_n1157_;
  assign new_n1159_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1160_ = ~new_n1151_ & ~new_n1152_;
  assign new_n1161_ = new_n1159_ & new_n1160_;
  assign pi7 = ~new_n1158_ | ~new_n1161_;
  assign pk5 = pm0 & pt3;
  assign new_n1164_ = ~pq0 & pw3;
  assign new_n1165_ = ~ph1 & new_n450_;
  assign new_n1166_ = ~pi1 & new_n1165_;
  assign new_n1167_ = pj1 & ~new_n465_;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = ~new_n477_ & new_n1168_;
  assign new_n1170_ = ~pk1 & new_n1169_;
  assign new_n1171_ = ~pl1 & new_n1169_;
  assign new_n1172_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = ~new_n453_ & ~new_n1172_;
  assign new_n1174_ = pk4 & new_n1173_;
  assign new_n1175_ = new_n450_ & new_n1174_;
  assign new_n1176_ = new_n488_ & new_n1175_;
  assign new_n1177_ = ~pi1 & new_n1174_;
  assign new_n1178_ = new_n488_ & new_n1177_;
  assign new_n1179_ = ~ph1 & new_n1175_;
  assign new_n1180_ = ~ph1 & new_n1177_;
  assign new_n1181_ = ~new_n1176_ & ~new_n1178_;
  assign new_n1182_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1183_ = new_n1181_ & new_n1182_;
  assign new_n1184_ = new_n1164_ & new_n1183_;
  assign new_n1185_ = po0 & new_n1184_;
  assign new_n1186_ = pt0 & new_n450_;
  assign new_n1187_ = pi1 & new_n1186_;
  assign new_n1188_ = ~pj1 & pv0;
  assign new_n1189_ = pk1 & new_n1188_;
  assign new_n1190_ = ~pl1 & new_n1189_;
  assign new_n1191_ = ~new_n465_ & ~new_n1190_;
  assign new_n1192_ = ~pw0 & new_n1191_;
  assign new_n1193_ = pj1 & new_n1191_;
  assign new_n1194_ = pj1 & ~new_n1190_;
  assign new_n1195_ = ~pu0 & new_n1194_;
  assign new_n1196_ = ~pj1 & ~new_n1190_;
  assign new_n1197_ = ~pw0 & new_n1196_;
  assign new_n1198_ = ~pw0 & ~new_n1190_;
  assign new_n1199_ = ~pu0 & new_n1198_;
  assign new_n1200_ = ~pk1 & pl1;
  assign new_n1201_ = ~new_n1190_ & ~new_n1200_;
  assign new_n1202_ = ~new_n465_ & new_n1201_;
  assign new_n1203_ = ~pu0 & new_n1201_;
  assign new_n1204_ = ~pj1 & new_n1201_;
  assign new_n1205_ = ~new_n1203_ & ~new_n1204_;
  assign new_n1206_ = ~new_n1199_ & ~new_n1202_;
  assign new_n1207_ = new_n1205_ & new_n1206_;
  assign new_n1208_ = ~new_n1192_ & ~new_n1193_;
  assign new_n1209_ = ~new_n1195_ & ~new_n1197_;
  assign new_n1210_ = new_n1208_ & new_n1209_;
  assign new_n1211_ = new_n1207_ & new_n1210_;
  assign new_n1212_ = ~pi1 & new_n1211_;
  assign new_n1213_ = ~new_n1187_ & ~new_n1212_;
  assign new_n1214_ = ~ps0 & new_n1213_;
  assign new_n1215_ = ~pi1 & ph1;
  assign new_n1216_ = new_n1213_ & ~new_n1215_;
  assign new_n1217_ = ph1 & ~new_n1215_;
  assign new_n1218_ = ph1 & ~new_n450_;
  assign new_n1219_ = ph1 & ~ps0;
  assign new_n1220_ = ~new_n450_ & new_n1213_;
  assign new_n1221_ = ~new_n1214_ & ~new_n1216_;
  assign new_n1222_ = ~new_n1217_ & new_n1221_;
  assign new_n1223_ = ~new_n1218_ & ~new_n1219_;
  assign new_n1224_ = ~new_n1220_ & new_n1223_;
  assign new_n1225_ = new_n1222_ & new_n1224_;
  assign new_n1226_ = new_n674_ & new_n1225_;
  assign new_n1227_ = new_n297_ & new_n1226_;
  assign pf9 = new_n1185_ | new_n1227_;
  assign new_n1229_ = pl4 & py2;
  assign new_n1230_ = px2 & ~new_n332_;
  assign new_n1231_ = ~pl4 & new_n1230_;
  assign new_n1232_ = pn & new_n337_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = ~new_n1229_ & new_n1233_;
  assign new_n1235_ = ~new_n293_ & new_n1234_;
  assign new_n1236_ = new_n293_ & new_n1233_;
  assign new_n1237_ = ~px2 & new_n1236_;
  assign new_n1238_ = ~px2 & new_n1234_;
  assign new_n1239_ = new_n351_ & new_n1233_;
  assign new_n1240_ = ~new_n1235_ & ~new_n1237_;
  assign new_n1241_ = ~new_n1238_ & ~new_n1239_;
  assign new_n1242_ = new_n1240_ & new_n1241_;
  assign new_n1243_ = po0 & new_n1242_;
  assign pg8 = ~pq0 & new_n1243_;
  assign new_n1245_ = ~py1 & new_n295_;
  assign new_n1246_ = pr & new_n297_;
  assign new_n1247_ = new_n301_ & ~new_n1246_;
  assign new_n1248_ = ~new_n1245_ & ~new_n1247_;
  assign new_n1249_ = ~pn0 & new_n1248_;
  assign new_n1250_ = new_n293_ & new_n1249_;
  assign new_n1251_ = pl4 & ~pz1;
  assign new_n1252_ = new_n1249_ & ~new_n1251_;
  assign new_n1253_ = py1 & new_n1248_;
  assign new_n1254_ = ~new_n1251_ & new_n1253_;
  assign new_n1255_ = new_n310_ & new_n1253_;
  assign new_n1256_ = new_n293_ & new_n1253_;
  assign new_n1257_ = new_n294_ & new_n1248_;
  assign new_n1258_ = ~new_n1251_ & new_n1257_;
  assign new_n1259_ = new_n310_ & new_n1257_;
  assign new_n1260_ = new_n310_ & new_n1249_;
  assign new_n1261_ = new_n293_ & new_n1257_;
  assign new_n1262_ = ~new_n1250_ & ~new_n1252_;
  assign new_n1263_ = ~new_n1254_ & new_n1262_;
  assign new_n1264_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1265_ = new_n1263_ & new_n1264_;
  assign new_n1266_ = ~new_n1260_ & ~new_n1261_;
  assign new_n1267_ = ~new_n1258_ & ~new_n1259_;
  assign new_n1268_ = new_n1266_ & new_n1267_;
  assign ph7 = ~new_n1265_ | ~new_n1268_;
  assign pj5 = pm0 & ps3;
  assign new_n1271_ = ~pc4 & new_n521_;
  assign new_n1272_ = py3 & new_n1271_;
  assign new_n1273_ = pz3 & new_n1272_;
  assign new_n1274_ = ~new_n520_ & new_n1273_;
  assign new_n1275_ = ~new_n1271_ & new_n1273_;
  assign new_n1276_ = pn1 & ~new_n1271_;
  assign new_n1277_ = pf1 & ~pi4;
  assign new_n1278_ = ~pf1 & pi4;
  assign new_n1279_ = ~new_n1277_ & ~new_n1278_;
  assign new_n1280_ = pn1 & new_n1279_;
  assign new_n1281_ = pn1 & ~new_n520_;
  assign new_n1282_ = new_n1273_ & new_n1279_;
  assign new_n1283_ = ~new_n1274_ & ~new_n1275_;
  assign new_n1284_ = ~new_n1276_ & new_n1283_;
  assign new_n1285_ = ~new_n1280_ & ~new_n1281_;
  assign new_n1286_ = ~new_n1282_ & new_n1285_;
  assign pu5 = ~new_n1284_ | ~new_n1286_;
  assign new_n1288_ = ~pg4 & ~ph4;
  assign new_n1289_ = pe4 & new_n1288_;
  assign new_n1290_ = pf4 & new_n1289_;
  assign new_n1291_ = ph1 & ~new_n1290_;
  assign new_n1292_ = ~px0 & new_n1291_;
  assign new_n1293_ = pi1 & ~new_n1290_;
  assign new_n1294_ = ~py0 & new_n1293_;
  assign new_n1295_ = ~pg1 & new_n451_;
  assign new_n1296_ = pd4 & new_n1295_;
  assign new_n1297_ = ~pg4 & new_n1296_;
  assign new_n1298_ = ~ph4 & new_n1297_;
  assign new_n1299_ = new_n1290_ & ~new_n1298_;
  assign new_n1300_ = pl1 & ~new_n1298_;
  assign new_n1301_ = ~pb1 & new_n1300_;
  assign new_n1302_ = ~pn4 & ~new_n1298_;
  assign new_n1303_ = ~new_n1299_ & ~new_n1301_;
  assign new_n1304_ = ~new_n1302_ & new_n1303_;
  assign new_n1305_ = pa1 & new_n1304_;
  assign new_n1306_ = ~pj1 & new_n1305_;
  assign new_n1307_ = pz0 & new_n1305_;
  assign new_n1308_ = ~pk1 & new_n1304_;
  assign new_n1309_ = ~pj1 & new_n1308_;
  assign new_n1310_ = pz0 & new_n1304_;
  assign new_n1311_ = ~pk1 & new_n1310_;
  assign new_n1312_ = new_n1290_ & new_n1304_;
  assign new_n1313_ = ~new_n1306_ & ~new_n1307_;
  assign new_n1314_ = ~new_n1309_ & new_n1313_;
  assign new_n1315_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1316_ = new_n1314_ & new_n1315_;
  assign new_n1317_ = ~new_n1292_ & ~new_n1294_;
  assign new_n1318_ = ~new_n1316_ & new_n1317_;
  assign new_n1319_ = pm1 & new_n1318_;
  assign new_n1320_ = po0 & ~new_n1319_;
  assign new_n1321_ = ~pq0 & new_n1320_;
  assign new_n1322_ = pp0 & new_n1321_;
  assign new_n1323_ = ~pn0 & new_n1322_;
  assign new_n1324_ = pm1 & new_n1321_;
  assign pv6 = new_n1323_ | new_n1324_;
  assign new_n1326_ = pl0 & pd;
  assign new_n1327_ = ~pl0 & pl;
  assign new_n1328_ = pk0 & new_n1327_;
  assign new_n1329_ = ~pk0 & pd;
  assign new_n1330_ = ~new_n1326_ & ~new_n1328_;
  assign new_n1331_ = ~new_n1329_ & new_n1330_;
  assign new_n1332_ = new_n310_ & new_n1331_;
  assign new_n1333_ = ~pm0 & new_n1332_;
  assign new_n1334_ = pl4 & ~po2;
  assign new_n1335_ = ~new_n336_ & new_n1334_;
  assign new_n1336_ = ~new_n293_ & new_n1335_;
  assign new_n1337_ = ~pn2 & new_n877_;
  assign new_n1338_ = ~new_n1333_ & ~new_n1336_;
  assign new_n1339_ = ~new_n1337_ & new_n1338_;
  assign new_n1340_ = po0 & new_n1339_;
  assign pw7 = ~pq0 & new_n1340_;
  assign new_n1342_ = po3 & ~pq0;
  assign new_n1343_ = new_n497_ & new_n1342_;
  assign new_n1344_ = po0 & new_n1343_;
  assign new_n1345_ = pp3 & ~new_n453_;
  assign new_n1346_ = pk4 & new_n1345_;
  assign new_n1347_ = new_n513_ & new_n1346_;
  assign new_n1348_ = new_n514_ & new_n1347_;
  assign px8 = new_n1344_ | new_n1348_;
  assign new_n1350_ = pl0 & pc;
  assign new_n1351_ = ~pl0 & pk;
  assign new_n1352_ = pk0 & new_n1351_;
  assign new_n1353_ = ~pk0 & pc;
  assign new_n1354_ = ~new_n1350_ & ~new_n1352_;
  assign new_n1355_ = ~new_n1353_ & new_n1354_;
  assign new_n1356_ = new_n310_ & new_n1355_;
  assign new_n1357_ = ~pm0 & new_n1356_;
  assign new_n1358_ = pl4 & ~pn2;
  assign new_n1359_ = ~new_n336_ & new_n1358_;
  assign new_n1360_ = ~new_n293_ & new_n1359_;
  assign new_n1361_ = ~pm2 & new_n877_;
  assign new_n1362_ = ~new_n1357_ & ~new_n1360_;
  assign new_n1363_ = ~new_n1361_ & new_n1362_;
  assign new_n1364_ = po0 & new_n1363_;
  assign pv7 = ~pq0 & new_n1364_;
  assign new_n1366_ = ~pn1 & new_n295_;
  assign new_n1367_ = pj0 & new_n297_;
  assign new_n1368_ = new_n301_ & ~new_n1367_;
  assign new_n1369_ = ~new_n1366_ & ~new_n1368_;
  assign new_n1370_ = ~pn0 & new_n1369_;
  assign new_n1371_ = new_n293_ & new_n1370_;
  assign new_n1372_ = pl4 & ~po1;
  assign new_n1373_ = new_n1370_ & ~new_n1372_;
  assign new_n1374_ = pn1 & new_n1369_;
  assign new_n1375_ = ~new_n1372_ & new_n1374_;
  assign new_n1376_ = new_n310_ & new_n1374_;
  assign new_n1377_ = new_n293_ & new_n1374_;
  assign new_n1378_ = new_n294_ & new_n1369_;
  assign new_n1379_ = ~new_n1372_ & new_n1378_;
  assign new_n1380_ = new_n310_ & new_n1378_;
  assign new_n1381_ = new_n310_ & new_n1370_;
  assign new_n1382_ = new_n293_ & new_n1378_;
  assign new_n1383_ = ~new_n1371_ & ~new_n1373_;
  assign new_n1384_ = ~new_n1375_ & new_n1383_;
  assign new_n1385_ = ~new_n1376_ & ~new_n1377_;
  assign new_n1386_ = new_n1384_ & new_n1385_;
  assign new_n1387_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1388_ = ~new_n1379_ & ~new_n1380_;
  assign new_n1389_ = new_n1387_ & new_n1388_;
  assign pw6 = ~new_n1386_ | ~new_n1389_;
  assign new_n1391_ = ~pq0 & pp3;
  assign new_n1392_ = new_n497_ & new_n1391_;
  assign new_n1393_ = po0 & new_n1392_;
  assign new_n1394_ = pq3 & ~new_n453_;
  assign new_n1395_ = pk4 & new_n1394_;
  assign new_n1396_ = new_n513_ & new_n1395_;
  assign new_n1397_ = new_n514_ & new_n1396_;
  assign py8 = new_n1393_ | new_n1397_;
  assign new_n1399_ = ~pe1 & ~pn0;
  assign new_n1400_ = new_n288_ & new_n1399_;
  assign new_n1401_ = ~pe1 & new_n288_;
  assign new_n1402_ = ~pn0 & new_n1401_;
  assign new_n1403_ = ~pk1 & ~new_n1402_;
  assign new_n1404_ = po0 & ~new_n1403_;
  assign new_n1405_ = ~pq0 & new_n1404_;
  assign new_n1406_ = new_n1400_ & new_n1405_;
  assign new_n1407_ = ~new_n288_ & new_n1406_;
  assign new_n1408_ = pn0 & new_n1406_;
  assign new_n1409_ = ~pg1 & new_n1405_;
  assign new_n1410_ = pn0 & new_n1409_;
  assign new_n1411_ = ~pc1 & ~pe1;
  assign new_n1412_ = ~pe1 & ~pd1;
  assign new_n1413_ = ~pc1 & ~pd1;
  assign new_n1414_ = ~new_n1411_ & ~new_n1412_;
  assign new_n1415_ = ~new_n1413_ & new_n1414_;
  assign new_n1416_ = new_n1409_ & new_n1415_;
  assign new_n1417_ = ~new_n288_ & new_n1409_;
  assign new_n1418_ = new_n1406_ & new_n1415_;
  assign new_n1419_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1420_ = ~new_n1410_ & new_n1419_;
  assign new_n1421_ = ~new_n1416_ & ~new_n1417_;
  assign new_n1422_ = ~new_n1418_ & new_n1421_;
  assign pt6 = ~new_n1420_ | ~new_n1422_;
  assign new_n1424_ = pl0 & pb;
  assign new_n1425_ = ~pl0 & pj;
  assign new_n1426_ = pk0 & new_n1425_;
  assign new_n1427_ = ~pk0 & pb;
  assign new_n1428_ = ~new_n1424_ & ~new_n1426_;
  assign new_n1429_ = ~new_n1427_ & new_n1428_;
  assign new_n1430_ = new_n310_ & new_n1429_;
  assign new_n1431_ = ~pm0 & new_n1430_;
  assign new_n1432_ = pl4 & ~pm2;
  assign new_n1433_ = ~new_n336_ & new_n1432_;
  assign new_n1434_ = ~new_n293_ & new_n1433_;
  assign new_n1435_ = ~pl2 & new_n877_;
  assign new_n1436_ = ~new_n1431_ & ~new_n1434_;
  assign new_n1437_ = ~new_n1435_ & new_n1436_;
  assign new_n1438_ = po0 & new_n1437_;
  assign pu7 = ~pq0 & new_n1438_;
  assign new_n1440_ = ~pe3 & pl0;
  assign new_n1441_ = pk0 & new_n1440_;
  assign new_n1442_ = ~pe3 & ~pl0;
  assign new_n1443_ = ~pk0 & new_n1442_;
  assign new_n1444_ = ~new_n1441_ & ~new_n1443_;
  assign new_n1445_ = pm0 & new_n1444_;
  assign new_n1446_ = pl0 & new_n1445_;
  assign new_n1447_ = pk0 & new_n1446_;
  assign new_n1448_ = ~pl0 & new_n1445_;
  assign new_n1449_ = ~pk0 & new_n1448_;
  assign new_n1450_ = pm3 & new_n1445_;
  assign new_n1451_ = ~new_n1447_ & ~new_n1449_;
  assign pv4 = new_n1450_ | ~new_n1451_;
  assign new_n1453_ = ~pq0 & pq3;
  assign new_n1454_ = new_n497_ & new_n1453_;
  assign new_n1455_ = po0 & new_n1454_;
  assign new_n1456_ = pr3 & ~new_n453_;
  assign new_n1457_ = pk4 & new_n1456_;
  assign new_n1458_ = new_n513_ & new_n1457_;
  assign new_n1459_ = new_n514_ & new_n1458_;
  assign pz8 = new_n1455_ | new_n1459_;
  assign new_n1461_ = pl0 & pa;
  assign new_n1462_ = ~pl0 & pi;
  assign new_n1463_ = pk0 & new_n1462_;
  assign new_n1464_ = ~pk0 & pa;
  assign new_n1465_ = ~new_n1461_ & ~new_n1463_;
  assign new_n1466_ = ~new_n1464_ & new_n1465_;
  assign new_n1467_ = new_n310_ & new_n1466_;
  assign new_n1468_ = ~pm0 & new_n1467_;
  assign new_n1469_ = pl4 & ~pl2;
  assign new_n1470_ = ~new_n336_ & new_n1469_;
  assign new_n1471_ = ~new_n293_ & new_n1470_;
  assign new_n1472_ = ~pk2 & new_n877_;
  assign new_n1473_ = ~new_n1468_ & ~new_n1471_;
  assign new_n1474_ = ~new_n1472_ & new_n1473_;
  assign new_n1475_ = po0 & new_n1474_;
  assign pt7 = ~pq0 & new_n1475_;
  assign new_n1477_ = po0 & ~new_n1402_;
  assign new_n1478_ = ~pq0 & new_n1477_;
  assign new_n1479_ = pl1 & new_n1478_;
  assign new_n1480_ = ~pg1 & new_n1479_;
  assign new_n1481_ = ~pd1 & new_n288_;
  assign new_n1482_ = ~pn0 & new_n1481_;
  assign new_n1483_ = ~pc1 & new_n1482_;
  assign new_n1484_ = new_n1478_ & new_n1483_;
  assign pu6 = new_n1480_ | new_n1484_;
  assign new_n1486_ = ~pf3 & pl0;
  assign new_n1487_ = pk0 & new_n1486_;
  assign new_n1488_ = ~pf3 & ~pl0;
  assign new_n1489_ = ~pk0 & new_n1488_;
  assign new_n1490_ = ~new_n1487_ & ~new_n1489_;
  assign new_n1491_ = pm0 & new_n1490_;
  assign new_n1492_ = pl0 & new_n1491_;
  assign new_n1493_ = pk0 & new_n1492_;
  assign new_n1494_ = ~pl0 & new_n1491_;
  assign new_n1495_ = ~pk0 & new_n1494_;
  assign new_n1496_ = pn3 & new_n1491_;
  assign new_n1497_ = ~new_n1493_ & ~new_n1495_;
  assign pw4 = new_n1496_ | ~new_n1497_;
  assign new_n1499_ = ~pd3 & ~pl3;
  assign new_n1500_ = ~pd3 & pl0;
  assign new_n1501_ = ~new_n759_ & ~new_n1499_;
  assign new_n1502_ = ~new_n1500_ & new_n1501_;
  assign new_n1503_ = ~pm0 & ~pt3;
  assign new_n1504_ = ~pd3 & ~pl0;
  assign new_n1505_ = ~new_n757_ & ~new_n1499_;
  assign new_n1506_ = ~new_n1504_ & new_n1505_;
  assign new_n1507_ = new_n1502_ & ~new_n1503_;
  assign new_n1508_ = new_n1506_ & new_n1507_;
  assign new_n1509_ = ~new_n1503_ & new_n1506_;
  assign new_n1510_ = ~pk0 & new_n1509_;
  assign new_n1511_ = pk0 & new_n1507_;
  assign new_n1512_ = ~pm0 & ~new_n1503_;
  assign new_n1513_ = ~new_n1508_ & ~new_n1510_;
  assign new_n1514_ = ~new_n1511_ & ~new_n1512_;
  assign pp4 = ~new_n1513_ | ~new_n1514_;
  assign new_n1516_ = pk1 & ~pn0;
  assign pq5 = pk4 | ~new_n1516_;
  assign new_n1518_ = ~pi1 & ~new_n1402_;
  assign new_n1519_ = po0 & ~new_n1518_;
  assign new_n1520_ = ~pq0 & new_n1519_;
  assign new_n1521_ = new_n1400_ & new_n1520_;
  assign new_n1522_ = ~new_n288_ & new_n1521_;
  assign new_n1523_ = pn0 & new_n1521_;
  assign new_n1524_ = ~pg1 & new_n1520_;
  assign new_n1525_ = pn0 & new_n1524_;
  assign new_n1526_ = ~pe1 & pd1;
  assign new_n1527_ = ~new_n1411_ & ~new_n1526_;
  assign new_n1528_ = ~new_n1413_ & new_n1527_;
  assign new_n1529_ = new_n1524_ & new_n1528_;
  assign new_n1530_ = ~new_n288_ & new_n1524_;
  assign new_n1531_ = new_n1521_ & new_n1528_;
  assign new_n1532_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1533_ = ~new_n1525_ & new_n1532_;
  assign new_n1534_ = ~new_n1529_ & ~new_n1530_;
  assign new_n1535_ = ~new_n1531_ & new_n1534_;
  assign pr6 = ~new_n1533_ | ~new_n1535_;
  assign new_n1537_ = ~pj2 & new_n295_;
  assign new_n1538_ = pc0 & new_n297_;
  assign new_n1539_ = new_n301_ & ~new_n1538_;
  assign new_n1540_ = ~new_n1537_ & ~new_n1539_;
  assign new_n1541_ = ~pn0 & new_n1540_;
  assign new_n1542_ = new_n293_ & new_n1541_;
  assign new_n1543_ = pl4 & ~pk2;
  assign new_n1544_ = new_n1541_ & ~new_n1543_;
  assign new_n1545_ = pj2 & new_n1540_;
  assign new_n1546_ = ~new_n1543_ & new_n1545_;
  assign new_n1547_ = new_n310_ & new_n1545_;
  assign new_n1548_ = new_n293_ & new_n1545_;
  assign new_n1549_ = new_n294_ & new_n1540_;
  assign new_n1550_ = ~new_n1543_ & new_n1549_;
  assign new_n1551_ = new_n310_ & new_n1549_;
  assign new_n1552_ = new_n310_ & new_n1541_;
  assign new_n1553_ = new_n293_ & new_n1549_;
  assign new_n1554_ = ~new_n1542_ & ~new_n1544_;
  assign new_n1555_ = ~new_n1546_ & new_n1554_;
  assign new_n1556_ = ~new_n1547_ & ~new_n1548_;
  assign new_n1557_ = new_n1555_ & new_n1556_;
  assign new_n1558_ = ~new_n1552_ & ~new_n1553_;
  assign new_n1559_ = ~new_n1550_ & ~new_n1551_;
  assign new_n1560_ = new_n1558_ & new_n1559_;
  assign ps7 = ~new_n1557_ | ~new_n1560_;
  assign new_n1562_ = pj1 & ~pn0;
  assign pp5 = pk4 | ~new_n1562_;
  assign new_n1564_ = ~pc3 & ~pk3;
  assign new_n1565_ = ~pc3 & pl0;
  assign new_n1566_ = ~new_n797_ & ~new_n1564_;
  assign new_n1567_ = ~new_n1565_ & new_n1566_;
  assign new_n1568_ = ~pm0 & ~ps3;
  assign new_n1569_ = ~pc3 & ~pl0;
  assign new_n1570_ = ~new_n795_ & ~new_n1564_;
  assign new_n1571_ = ~new_n1569_ & new_n1570_;
  assign new_n1572_ = new_n1567_ & ~new_n1568_;
  assign new_n1573_ = new_n1571_ & new_n1572_;
  assign new_n1574_ = ~new_n1568_ & new_n1571_;
  assign new_n1575_ = ~pk0 & new_n1574_;
  assign new_n1576_ = pk0 & new_n1572_;
  assign new_n1577_ = ~pm0 & ~new_n1568_;
  assign new_n1578_ = ~new_n1573_ & ~new_n1575_;
  assign new_n1579_ = ~new_n1576_ & ~new_n1577_;
  assign pq4 = ~new_n1578_ | ~new_n1579_;
  assign new_n1581_ = ~pi2 & new_n295_;
  assign new_n1582_ = pb0 & new_n297_;
  assign new_n1583_ = new_n301_ & ~new_n1582_;
  assign new_n1584_ = ~new_n1581_ & ~new_n1583_;
  assign new_n1585_ = ~pn0 & new_n1584_;
  assign new_n1586_ = new_n293_ & new_n1585_;
  assign new_n1587_ = ~pj2 & pl4;
  assign new_n1588_ = new_n1585_ & ~new_n1587_;
  assign new_n1589_ = pi2 & new_n1584_;
  assign new_n1590_ = ~new_n1587_ & new_n1589_;
  assign new_n1591_ = new_n310_ & new_n1589_;
  assign new_n1592_ = new_n293_ & new_n1589_;
  assign new_n1593_ = new_n294_ & new_n1584_;
  assign new_n1594_ = ~new_n1587_ & new_n1593_;
  assign new_n1595_ = new_n310_ & new_n1593_;
  assign new_n1596_ = new_n310_ & new_n1585_;
  assign new_n1597_ = new_n293_ & new_n1593_;
  assign new_n1598_ = ~new_n1586_ & ~new_n1588_;
  assign new_n1599_ = ~new_n1590_ & new_n1598_;
  assign new_n1600_ = ~new_n1591_ & ~new_n1592_;
  assign new_n1601_ = new_n1599_ & new_n1600_;
  assign new_n1602_ = ~new_n1596_ & ~new_n1597_;
  assign new_n1603_ = ~new_n1594_ & ~new_n1595_;
  assign new_n1604_ = new_n1602_ & new_n1603_;
  assign pr7 = ~new_n1601_ | ~new_n1604_;
  assign new_n1606_ = ~pj1 & ~new_n1402_;
  assign new_n1607_ = po0 & ~new_n1606_;
  assign new_n1608_ = ~pq0 & new_n1607_;
  assign new_n1609_ = new_n1400_ & new_n1608_;
  assign new_n1610_ = ~new_n288_ & new_n1609_;
  assign new_n1611_ = pn0 & new_n1609_;
  assign new_n1612_ = ~pg1 & new_n1608_;
  assign new_n1613_ = pn0 & new_n1612_;
  assign new_n1614_ = pc1 & ~pe1;
  assign new_n1615_ = ~new_n1412_ & ~new_n1614_;
  assign new_n1616_ = ~new_n1413_ & new_n1615_;
  assign new_n1617_ = new_n1612_ & new_n1616_;
  assign new_n1618_ = ~new_n288_ & new_n1612_;
  assign new_n1619_ = new_n1609_ & new_n1616_;
  assign new_n1620_ = ~new_n1610_ & ~new_n1611_;
  assign new_n1621_ = ~new_n1613_ & new_n1620_;
  assign new_n1622_ = ~new_n1617_ & ~new_n1618_;
  assign new_n1623_ = ~new_n1619_ & new_n1622_;
  assign ps6 = ~new_n1621_ | ~new_n1623_;
  assign pp6 = new_n297_ & new_n1318_;
  assign new_n1626_ = ~ph2 & new_n295_;
  assign new_n1627_ = pa0 & new_n297_;
  assign new_n1628_ = new_n301_ & ~new_n1627_;
  assign new_n1629_ = ~new_n1626_ & ~new_n1628_;
  assign new_n1630_ = ~pn0 & new_n1629_;
  assign new_n1631_ = new_n293_ & new_n1630_;
  assign new_n1632_ = pl4 & ~pi2;
  assign new_n1633_ = new_n1630_ & ~new_n1632_;
  assign new_n1634_ = ph2 & new_n1629_;
  assign new_n1635_ = ~new_n1632_ & new_n1634_;
  assign new_n1636_ = new_n310_ & new_n1634_;
  assign new_n1637_ = new_n293_ & new_n1634_;
  assign new_n1638_ = new_n294_ & new_n1629_;
  assign new_n1639_ = ~new_n1632_ & new_n1638_;
  assign new_n1640_ = new_n310_ & new_n1638_;
  assign new_n1641_ = new_n310_ & new_n1630_;
  assign new_n1642_ = new_n293_ & new_n1638_;
  assign new_n1643_ = ~new_n1631_ & ~new_n1633_;
  assign new_n1644_ = ~new_n1635_ & new_n1643_;
  assign new_n1645_ = ~new_n1636_ & ~new_n1637_;
  assign new_n1646_ = new_n1644_ & new_n1645_;
  assign new_n1647_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1648_ = ~new_n1639_ & ~new_n1640_;
  assign new_n1649_ = new_n1647_ & new_n1648_;
  assign pq7 = ~new_n1646_ | ~new_n1649_;
  assign new_n1651_ = ~pb3 & ~pj3;
  assign new_n1652_ = ~pb3 & pl0;
  assign new_n1653_ = ~new_n620_ & ~new_n1651_;
  assign new_n1654_ = ~new_n1652_ & new_n1653_;
  assign new_n1655_ = ~pm0 & ~pr3;
  assign new_n1656_ = ~pb3 & ~pl0;
  assign new_n1657_ = ~new_n618_ & ~new_n1651_;
  assign new_n1658_ = ~new_n1656_ & new_n1657_;
  assign new_n1659_ = new_n1654_ & ~new_n1655_;
  assign new_n1660_ = new_n1658_ & new_n1659_;
  assign new_n1661_ = ~new_n1655_ & new_n1658_;
  assign new_n1662_ = ~pk0 & new_n1661_;
  assign new_n1663_ = pk0 & new_n1659_;
  assign new_n1664_ = ~pm0 & ~new_n1655_;
  assign new_n1665_ = ~new_n1660_ & ~new_n1662_;
  assign new_n1666_ = ~new_n1663_ & ~new_n1664_;
  assign pr4 = ~new_n1665_ | ~new_n1666_;
  assign new_n1668_ = ~pg2 & new_n295_;
  assign new_n1669_ = pz & new_n297_;
  assign new_n1670_ = new_n301_ & ~new_n1669_;
  assign new_n1671_ = ~new_n1668_ & ~new_n1670_;
  assign new_n1672_ = ~pn0 & new_n1671_;
  assign new_n1673_ = new_n293_ & new_n1672_;
  assign new_n1674_ = pl4 & ~ph2;
  assign new_n1675_ = new_n1672_ & ~new_n1674_;
  assign new_n1676_ = pg2 & new_n1671_;
  assign new_n1677_ = ~new_n1674_ & new_n1676_;
  assign new_n1678_ = new_n310_ & new_n1676_;
  assign new_n1679_ = new_n293_ & new_n1676_;
  assign new_n1680_ = new_n294_ & new_n1671_;
  assign new_n1681_ = ~new_n1674_ & new_n1680_;
  assign new_n1682_ = new_n310_ & new_n1680_;
  assign new_n1683_ = new_n310_ & new_n1672_;
  assign new_n1684_ = new_n293_ & new_n1680_;
  assign new_n1685_ = ~new_n1673_ & ~new_n1675_;
  assign new_n1686_ = ~new_n1677_ & new_n1685_;
  assign new_n1687_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1688_ = new_n1686_ & new_n1687_;
  assign new_n1689_ = ~new_n1683_ & ~new_n1684_;
  assign new_n1690_ = ~new_n1681_ & ~new_n1682_;
  assign new_n1691_ = new_n1689_ & new_n1690_;
  assign pp7 = ~new_n1688_ | ~new_n1691_;
  assign new_n1693_ = ph1 & new_n669_;
  assign new_n1694_ = pc1 & pe1;
  assign new_n1695_ = pe1 & pd1;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = ~pn0 & new_n1696_;
  assign new_n1698_ = new_n288_ & new_n1697_;
  assign new_n1699_ = new_n1693_ & ~new_n1698_;
  assign new_n1700_ = po0 & new_n1699_;
  assign new_n1701_ = ~pc1 & new_n297_;
  assign new_n1702_ = new_n288_ & new_n1412_;
  assign new_n1703_ = new_n1701_ & new_n1702_;
  assign new_n1704_ = ~pn0 & new_n1703_;
  assign pq6 = new_n1700_ | new_n1704_;
  assign new_n1706_ = pl1 & ~pn0;
  assign pr5 = pk4 | ~new_n1706_;
  assign new_n1708_ = ~pi3 & ~pl0;
  assign new_n1709_ = ~pa3 & ~pi3;
  assign new_n1710_ = ~pa3 & pl0;
  assign new_n1711_ = ~new_n1708_ & ~new_n1709_;
  assign new_n1712_ = ~new_n1710_ & new_n1711_;
  assign new_n1713_ = ~pm0 & ~pq3;
  assign new_n1714_ = ~pi3 & pl0;
  assign new_n1715_ = ~pa3 & ~pl0;
  assign new_n1716_ = ~new_n1709_ & ~new_n1714_;
  assign new_n1717_ = ~new_n1715_ & new_n1716_;
  assign new_n1718_ = new_n1712_ & ~new_n1713_;
  assign new_n1719_ = new_n1717_ & new_n1718_;
  assign new_n1720_ = ~new_n1713_ & new_n1717_;
  assign new_n1721_ = ~pk0 & new_n1720_;
  assign new_n1722_ = pk0 & new_n1718_;
  assign new_n1723_ = ~pm0 & ~new_n1713_;
  assign new_n1724_ = ~new_n1719_ & ~new_n1721_;
  assign new_n1725_ = ~new_n1722_ & ~new_n1723_;
  assign ps4 = ~new_n1724_ | ~new_n1725_;
  assign new_n1727_ = pg3 & ~pq0;
  assign new_n1728_ = new_n497_ & new_n1727_;
  assign new_n1729_ = po0 & new_n1728_;
  assign new_n1730_ = ph3 & ~new_n453_;
  assign new_n1731_ = pk4 & new_n1730_;
  assign new_n1732_ = new_n513_ & new_n1731_;
  assign new_n1733_ = new_n514_ & new_n1732_;
  assign pp8 = new_n1729_ | new_n1733_;
  assign new_n1735_ = pf4 & new_n786_;
  assign new_n1736_ = pk4 & new_n1288_;
  assign new_n1737_ = ~pg1 & ~new_n453_;
  assign new_n1738_ = new_n1735_ & new_n1736_;
  assign new_n1739_ = new_n1737_ & new_n1738_;
  assign new_n1740_ = ~new_n310_ & new_n514_;
  assign new_n1741_ = new_n1739_ & new_n1740_;
  assign new_n1742_ = ph4 & new_n669_;
  assign new_n1743_ = pe4 & new_n778_;
  assign new_n1744_ = pf4 & ~pg4;
  assign new_n1745_ = pk4 & new_n1744_;
  assign new_n1746_ = new_n1743_ & new_n1745_;
  assign new_n1747_ = ~new_n477_ & new_n1746_;
  assign new_n1748_ = ~new_n310_ & ~new_n1747_;
  assign new_n1749_ = new_n1742_ & new_n1748_;
  assign new_n1750_ = po0 & new_n1749_;
  assign new_n1751_ = ~new_n1741_ & ~new_n1750_;
  assign pq9 = new_n538_ | ~new_n1751_;
  assign new_n1753_ = ~pq0 & ~new_n477_;
  assign new_n1754_ = ~new_n453_ & new_n1753_;
  assign new_n1755_ = ~pd4 & ~pg1;
  assign new_n1756_ = pe4 & new_n1755_;
  assign new_n1757_ = new_n1745_ & new_n1756_;
  assign new_n1758_ = po0 & new_n1757_;
  assign new_n1759_ = ~new_n310_ & new_n1754_;
  assign new_n1760_ = new_n1758_ & new_n1759_;
  assign new_n1761_ = pg4 & new_n669_;
  assign new_n1762_ = pk4 & new_n451_;
  assign new_n1763_ = new_n778_ & new_n1762_;
  assign new_n1764_ = ~new_n477_ & new_n1763_;
  assign new_n1765_ = ~new_n310_ & ~new_n1764_;
  assign new_n1766_ = new_n1761_ & new_n1765_;
  assign new_n1767_ = po0 & new_n1766_;
  assign new_n1768_ = pl0 & pm0;
  assign new_n1769_ = ~pk0 & new_n1768_;
  assign new_n1770_ = ~pl0 & pm0;
  assign new_n1771_ = pk0 & new_n1770_;
  assign new_n1772_ = ~new_n1769_ & ~new_n1771_;
  assign new_n1773_ = ~pn0 & new_n1772_;
  assign new_n1774_ = po0 & new_n1773_;
  assign new_n1775_ = ~pq0 & new_n1774_;
  assign new_n1776_ = new_n288_ & new_n1775_;
  assign new_n1777_ = ~new_n1760_ & ~new_n1767_;
  assign pp9 = new_n1776_ | ~new_n1777_;
  assign new_n1779_ = ph3 & ~pq0;
  assign new_n1780_ = new_n497_ & new_n1779_;
  assign new_n1781_ = po0 & new_n1780_;
  assign new_n1782_ = pi3 & ~new_n453_;
  assign new_n1783_ = pk4 & new_n1782_;
  assign new_n1784_ = new_n513_ & new_n1783_;
  assign new_n1785_ = new_n514_ & new_n1784_;
  assign pq8 = new_n1781_ | new_n1785_;
  assign new_n1787_ = pi3 & ~pq0;
  assign new_n1788_ = new_n497_ & new_n1787_;
  assign new_n1789_ = po0 & new_n1788_;
  assign new_n1790_ = pj3 & ~new_n453_;
  assign new_n1791_ = pk4 & new_n1790_;
  assign new_n1792_ = new_n513_ & new_n1791_;
  assign new_n1793_ = new_n514_ & new_n1792_;
  assign pr8 = new_n1789_ | new_n1793_;
  assign new_n1795_ = pj4 & new_n669_;
  assign new_n1796_ = ps0 & new_n450_;
  assign new_n1797_ = ~pi1 & new_n1796_;
  assign new_n1798_ = pt0 & new_n465_;
  assign new_n1799_ = ~pj1 & new_n1798_;
  assign new_n1800_ = pi1 & ~new_n1799_;
  assign new_n1801_ = ~pi1 & ~pk1;
  assign new_n1802_ = ~pl1 & new_n1801_;
  assign new_n1803_ = ~pu0 & new_n1802_;
  assign new_n1804_ = ~ph1 & new_n1803_;
  assign new_n1805_ = ~pl1 & ~new_n453_;
  assign new_n1806_ = ~pk1 & new_n1805_;
  assign new_n1807_ = ~pj1 & ~new_n453_;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_ = ~new_n484_ & ~new_n1808_;
  assign new_n1810_ = ~new_n477_ & new_n1809_;
  assign new_n1811_ = pk4 & new_n1810_;
  assign new_n1812_ = pn4 & new_n1811_;
  assign new_n1813_ = ~new_n1800_ & ~new_n1804_;
  assign new_n1814_ = new_n1812_ & new_n1813_;
  assign new_n1815_ = ~pi1 & ~pj1;
  assign new_n1816_ = new_n1797_ & new_n1814_;
  assign new_n1817_ = ~new_n1815_ & new_n1816_;
  assign new_n1818_ = ~pl1 & ~pv0;
  assign new_n1819_ = ~pk1 & ~pw0;
  assign new_n1820_ = ~new_n465_ & ~new_n1818_;
  assign new_n1821_ = ~new_n1819_ & new_n1820_;
  assign new_n1822_ = new_n1816_ & new_n1821_;
  assign new_n1823_ = new_n1814_ & new_n1821_;
  assign new_n1824_ = ~ph1 & new_n1823_;
  assign new_n1825_ = ph1 & new_n1816_;
  assign new_n1826_ = new_n1814_ & ~new_n1815_;
  assign new_n1827_ = ~ph1 & new_n1826_;
  assign new_n1828_ = ~new_n1817_ & ~new_n1822_;
  assign new_n1829_ = ~new_n1824_ & new_n1828_;
  assign new_n1830_ = ~new_n1825_ & ~new_n1827_;
  assign new_n1831_ = new_n1829_ & new_n1830_;
  assign new_n1832_ = new_n1795_ & new_n1831_;
  assign new_n1833_ = po0 & new_n1832_;
  assign new_n1834_ = ~pg1 & new_n673_;
  assign new_n1835_ = ~pj4 & pk4;
  assign new_n1836_ = pn4 & new_n1835_;
  assign new_n1837_ = po0 & new_n1836_;
  assign new_n1838_ = ~pq0 & new_n1837_;
  assign new_n1839_ = new_n1225_ & new_n1834_;
  assign new_n1840_ = new_n1838_ & new_n1839_;
  assign ps9 = new_n1833_ | new_n1840_;
  assign new_n1842_ = pi4 & pn1;
  assign new_n1843_ = ~new_n293_ & new_n297_;
  assign new_n1844_ = ~new_n1842_ & new_n1843_;
  assign new_n1845_ = pl4 & new_n1844_;
  assign new_n1846_ = pn1 & new_n1845_;
  assign new_n1847_ = pi4 & new_n1845_;
  assign pr9 = new_n1846_ | new_n1847_;
  assign new_n1849_ = pj3 & ~pq0;
  assign new_n1850_ = new_n497_ & new_n1849_;
  assign new_n1851_ = po0 & new_n1850_;
  assign new_n1852_ = pk3 & ~new_n453_;
  assign new_n1853_ = pk4 & new_n1852_;
  assign new_n1854_ = new_n513_ & new_n1853_;
  assign new_n1855_ = new_n514_ & new_n1854_;
  assign ps8 = new_n1851_ | new_n1855_;
  assign new_n1857_ = pk3 & ~pq0;
  assign new_n1858_ = new_n497_ & new_n1857_;
  assign new_n1859_ = po0 & new_n1858_;
  assign new_n1860_ = pl3 & ~new_n453_;
  assign new_n1861_ = pk4 & new_n1860_;
  assign new_n1862_ = new_n513_ & new_n1861_;
  assign new_n1863_ = new_n514_ & new_n1862_;
  assign pt8 = new_n1859_ | new_n1863_;
  assign pu9 = pm1 & new_n1843_;
  assign new_n1866_ = ~pg3 & pl0;
  assign new_n1867_ = pk0 & new_n1866_;
  assign new_n1868_ = ~pg3 & ~pl0;
  assign new_n1869_ = ~pk0 & new_n1868_;
  assign new_n1870_ = ~new_n1867_ & ~new_n1869_;
  assign new_n1871_ = pm0 & new_n1870_;
  assign new_n1872_ = pl0 & new_n1871_;
  assign new_n1873_ = pk0 & new_n1872_;
  assign new_n1874_ = ~pl0 & new_n1871_;
  assign new_n1875_ = ~pk0 & new_n1874_;
  assign new_n1876_ = po3 & new_n1871_;
  assign new_n1877_ = ~new_n1873_ & ~new_n1875_;
  assign px4 = new_n1876_ | ~new_n1877_;
  assign new_n1879_ = pi1 & pm1;
  assign py5 = pk4 | ~new_n1879_;
  assign new_n1881_ = ~pq1 & new_n295_;
  assign new_n1882_ = pg0 & new_n297_;
  assign new_n1883_ = new_n301_ & ~new_n1882_;
  assign new_n1884_ = ~new_n1881_ & ~new_n1883_;
  assign new_n1885_ = ~pn0 & new_n1884_;
  assign new_n1886_ = new_n293_ & new_n1885_;
  assign new_n1887_ = pl4 & ~pr1;
  assign new_n1888_ = new_n1885_ & ~new_n1887_;
  assign new_n1889_ = pq1 & new_n1884_;
  assign new_n1890_ = ~new_n1887_ & new_n1889_;
  assign new_n1891_ = new_n310_ & new_n1889_;
  assign new_n1892_ = new_n293_ & new_n1889_;
  assign new_n1893_ = new_n294_ & new_n1884_;
  assign new_n1894_ = ~new_n1887_ & new_n1893_;
  assign new_n1895_ = new_n310_ & new_n1893_;
  assign new_n1896_ = new_n310_ & new_n1885_;
  assign new_n1897_ = new_n293_ & new_n1893_;
  assign new_n1898_ = ~new_n1886_ & ~new_n1888_;
  assign new_n1899_ = ~new_n1890_ & new_n1898_;
  assign new_n1900_ = ~new_n1891_ & ~new_n1892_;
  assign new_n1901_ = new_n1899_ & new_n1900_;
  assign new_n1902_ = ~new_n1896_ & ~new_n1897_;
  assign new_n1903_ = ~new_n1894_ & ~new_n1895_;
  assign new_n1904_ = new_n1902_ & new_n1903_;
  assign pz6 = ~new_n1901_ | ~new_n1904_;
  assign new_n1906_ = pm1 & ~pq0;
  assign new_n1907_ = new_n706_ & new_n1906_;
  assign new_n1908_ = po0 & new_n1907_;
  assign new_n1909_ = ~pb4 & new_n1908_;
  assign pt9 = ~pc4 & new_n1909_;
  assign new_n1911_ = pl3 & ~pq0;
  assign new_n1912_ = new_n497_ & new_n1911_;
  assign new_n1913_ = po0 & new_n1912_;
  assign new_n1914_ = pm3 & ~new_n453_;
  assign new_n1915_ = pk4 & new_n1914_;
  assign new_n1916_ = new_n513_ & new_n1915_;
  assign new_n1917_ = new_n514_ & new_n1916_;
  assign pu8 = new_n1913_ | new_n1917_;
  assign new_n1919_ = ph1 & pm1;
  assign px5 = pk4 | ~new_n1919_;
  assign new_n1921_ = ~ph3 & pl0;
  assign new_n1922_ = pk0 & new_n1921_;
  assign new_n1923_ = ~ph3 & ~pl0;
  assign new_n1924_ = ~pk0 & new_n1923_;
  assign new_n1925_ = ~new_n1922_ & ~new_n1924_;
  assign new_n1926_ = pm0 & new_n1925_;
  assign new_n1927_ = pl0 & new_n1926_;
  assign new_n1928_ = pk0 & new_n1927_;
  assign new_n1929_ = ~pl0 & new_n1926_;
  assign new_n1930_ = ~pk0 & new_n1929_;
  assign new_n1931_ = pp3 & new_n1926_;
  assign new_n1932_ = ~new_n1928_ & ~new_n1930_;
  assign py4 = new_n1931_ | ~new_n1932_;
  assign new_n1934_ = pl0 & pg;
  assign new_n1935_ = ~pl0 & po;
  assign new_n1936_ = pk0 & new_n1935_;
  assign new_n1937_ = ~pk0 & pg;
  assign new_n1938_ = ~new_n1934_ & ~new_n1936_;
  assign new_n1939_ = ~new_n1937_ & new_n1938_;
  assign new_n1940_ = new_n310_ & new_n1939_;
  assign new_n1941_ = ~pm0 & new_n1940_;
  assign new_n1942_ = pl4 & ~pr2;
  assign new_n1943_ = ~new_n336_ & new_n1942_;
  assign new_n1944_ = ~new_n293_ & new_n1943_;
  assign new_n1945_ = ~pq2 & new_n877_;
  assign new_n1946_ = ~new_n1941_ & ~new_n1944_;
  assign new_n1947_ = ~new_n1945_ & new_n1946_;
  assign new_n1948_ = po0 & new_n1947_;
  assign pz7 = ~pq0 & new_n1948_;
  assign new_n1950_ = pm3 & ~pq0;
  assign new_n1951_ = new_n497_ & new_n1950_;
  assign new_n1952_ = po0 & new_n1951_;
  assign new_n1953_ = pn3 & ~new_n453_;
  assign new_n1954_ = pk4 & new_n1953_;
  assign new_n1955_ = new_n513_ & new_n1954_;
  assign new_n1956_ = new_n514_ & new_n1955_;
  assign pv8 = new_n1952_ | new_n1956_;
  assign pw9 = pk4 & new_n514_;
  assign new_n1959_ = ~po1 & new_n295_;
  assign new_n1960_ = pi0 & new_n297_;
  assign new_n1961_ = new_n301_ & ~new_n1960_;
  assign new_n1962_ = ~new_n1959_ & ~new_n1961_;
  assign new_n1963_ = ~pn0 & new_n1962_;
  assign new_n1964_ = new_n293_ & new_n1963_;
  assign new_n1965_ = pl4 & ~pp1;
  assign new_n1966_ = new_n1963_ & ~new_n1965_;
  assign new_n1967_ = po1 & new_n1962_;
  assign new_n1968_ = ~new_n1965_ & new_n1967_;
  assign new_n1969_ = new_n310_ & new_n1967_;
  assign new_n1970_ = new_n293_ & new_n1967_;
  assign new_n1971_ = new_n294_ & new_n1962_;
  assign new_n1972_ = ~new_n1965_ & new_n1971_;
  assign new_n1973_ = new_n310_ & new_n1971_;
  assign new_n1974_ = new_n310_ & new_n1963_;
  assign new_n1975_ = new_n293_ & new_n1971_;
  assign new_n1976_ = ~new_n1964_ & ~new_n1966_;
  assign new_n1977_ = ~new_n1968_ & new_n1976_;
  assign new_n1978_ = ~new_n1969_ & ~new_n1970_;
  assign new_n1979_ = new_n1977_ & new_n1978_;
  assign new_n1980_ = ~new_n1974_ & ~new_n1975_;
  assign new_n1981_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1982_ = new_n1980_ & new_n1981_;
  assign px6 = ~new_n1979_ | ~new_n1982_;
  assign new_n1984_ = pl0 & pf;
  assign new_n1985_ = ~pl0 & pn;
  assign new_n1986_ = pk0 & new_n1985_;
  assign new_n1987_ = ~pk0 & pf;
  assign new_n1988_ = ~new_n1984_ & ~new_n1986_;
  assign new_n1989_ = ~new_n1987_ & new_n1988_;
  assign new_n1990_ = new_n310_ & new_n1989_;
  assign new_n1991_ = ~pm0 & new_n1990_;
  assign new_n1992_ = pl4 & ~pq2;
  assign new_n1993_ = ~new_n336_ & new_n1992_;
  assign new_n1994_ = ~new_n293_ & new_n1993_;
  assign new_n1995_ = ~pp2 & new_n877_;
  assign new_n1996_ = ~new_n1991_ & ~new_n1994_;
  assign new_n1997_ = ~new_n1995_ & new_n1996_;
  assign new_n1998_ = po0 & new_n1997_;
  assign py7 = ~pq0 & new_n1998_;
  assign new_n2000_ = pk0 & new_n1714_;
  assign new_n2001_ = ~pk0 & new_n1708_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = pm0 & new_n2002_;
  assign new_n2004_ = pl0 & new_n2003_;
  assign new_n2005_ = pk0 & new_n2004_;
  assign new_n2006_ = ~pl0 & new_n2003_;
  assign new_n2007_ = ~pk0 & new_n2006_;
  assign new_n2008_ = pq3 & new_n2003_;
  assign new_n2009_ = ~new_n2005_ & ~new_n2007_;
  assign pz4 = new_n2008_ | ~new_n2009_;
  assign new_n2011_ = ~pa1 & pk1;
  assign new_n2012_ = ~pb1 & pl1;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = ~new_n453_ & new_n2013_;
  assign new_n2015_ = pz0 & new_n2014_;
  assign new_n2016_ = py0 & new_n2015_;
  assign new_n2017_ = ~pj1 & new_n2014_;
  assign new_n2018_ = py0 & new_n2017_;
  assign new_n2019_ = ~pi1 & new_n2015_;
  assign new_n2020_ = ~pi1 & new_n2017_;
  assign new_n2021_ = ~new_n2016_ & ~new_n2018_;
  assign new_n2022_ = ~new_n2019_ & ~new_n2020_;
  assign new_n2023_ = new_n2021_ & new_n2022_;
  assign new_n2024_ = ~new_n455_ & ~new_n2023_;
  assign new_n2025_ = pn4 & new_n2024_;
  assign new_n2026_ = new_n477_ & ~new_n2025_;
  assign new_n2027_ = po0 & ~new_n2026_;
  assign new_n2028_ = ~pq0 & new_n2027_;
  assign new_n2029_ = new_n2025_ & new_n2028_;
  assign new_n2030_ = new_n1318_ & new_n2028_;
  assign pv9 = new_n2029_ | new_n2030_;
  assign new_n2032_ = pn3 & ~pq0;
  assign new_n2033_ = new_n497_ & new_n2032_;
  assign new_n2034_ = po0 & new_n2033_;
  assign new_n2035_ = po3 & ~new_n453_;
  assign new_n2036_ = pk4 & new_n2035_;
  assign new_n2037_ = new_n513_ & new_n2036_;
  assign new_n2038_ = new_n514_ & new_n2037_;
  assign pw8 = new_n2034_ | new_n2038_;
  assign new_n2040_ = pl0 & pe;
  assign new_n2041_ = ~pl0 & pm;
  assign new_n2042_ = pk0 & new_n2041_;
  assign new_n2043_ = ~pk0 & pe;
  assign new_n2044_ = ~new_n2040_ & ~new_n2042_;
  assign new_n2045_ = ~new_n2043_ & new_n2044_;
  assign new_n2046_ = new_n310_ & new_n2045_;
  assign new_n2047_ = ~pm0 & new_n2046_;
  assign new_n2048_ = pl4 & ~pp2;
  assign new_n2049_ = ~new_n336_ & new_n2048_;
  assign new_n2050_ = ~new_n293_ & new_n2049_;
  assign new_n2051_ = ~po2 & new_n877_;
  assign new_n2052_ = ~new_n2047_ & ~new_n2050_;
  assign new_n2053_ = ~new_n2051_ & new_n2052_;
  assign new_n2054_ = po0 & new_n2053_;
  assign px7 = ~pq0 & new_n2054_;
  assign new_n2056_ = ~pp1 & new_n295_;
  assign new_n2057_ = ph0 & new_n297_;
  assign new_n2058_ = new_n301_ & ~new_n2057_;
  assign new_n2059_ = ~new_n2056_ & ~new_n2058_;
  assign new_n2060_ = ~pn0 & new_n2059_;
  assign new_n2061_ = new_n293_ & new_n2060_;
  assign new_n2062_ = pl4 & ~pq1;
  assign new_n2063_ = new_n2060_ & ~new_n2062_;
  assign new_n2064_ = pp1 & new_n2059_;
  assign new_n2065_ = ~new_n2062_ & new_n2064_;
  assign new_n2066_ = new_n310_ & new_n2064_;
  assign new_n2067_ = new_n293_ & new_n2064_;
  assign new_n2068_ = new_n294_ & new_n2059_;
  assign new_n2069_ = ~new_n2062_ & new_n2068_;
  assign new_n2070_ = new_n310_ & new_n2068_;
  assign new_n2071_ = new_n310_ & new_n2060_;
  assign new_n2072_ = new_n293_ & new_n2068_;
  assign new_n2073_ = ~new_n2061_ & ~new_n2063_;
  assign new_n2074_ = ~new_n2065_ & new_n2073_;
  assign new_n2075_ = ~new_n2066_ & ~new_n2067_;
  assign new_n2076_ = new_n2074_ & new_n2075_;
  assign new_n2077_ = ~new_n2071_ & ~new_n2072_;
  assign new_n2078_ = ~new_n2069_ & ~new_n2070_;
  assign new_n2079_ = new_n2077_ & new_n2078_;
  assign py6 = ~new_n2076_ | ~new_n2079_;
  assign new_n2081_ = pj1 & pm1;
  assign pz5 = pk4 | ~new_n2081_;
  assign pl6 = ~pl1;
  assign po4 = ~pg1;
  assign pj6 = ~pj1;
  assign pk6 = ~pk1;
  assign ph6 = ~ph1;
  assign pi6 = ~pi1;
  assign pm5 = pm4;
  assign pm6 = pk4;
  assign pt4 = pu3;
  assign pt5 = pu5;
  assign pu4 = pv3;
  assign pw5 = pu5;
  assign pv5 = pu5;
  assign ps5 = pu5;
endmodule

