// Benchmark "testing" written by ABC on Thu Oct  8 22:16:37 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A7  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A7;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2311]_ , \new_[2312]_ ,
    \new_[2313]_ , \new_[2314]_ , \new_[2315]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2385]_ , \new_[2386]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2389]_ , \new_[2390]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2395]_ , \new_[2396]_ ,
    \new_[2397]_ , \new_[2398]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2570]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2574]_ , \new_[2575]_ , \new_[2576]_ ,
    \new_[2577]_ , \new_[2578]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2602]_ , \new_[2603]_ , \new_[2604]_ ,
    \new_[2605]_ , \new_[2606]_ , \new_[2607]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2610]_ , \new_[2611]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2614]_ , \new_[2615]_ , \new_[2616]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2619]_ , \new_[2620]_ ,
    \new_[2621]_ , \new_[2622]_ , \new_[2623]_ , \new_[2624]_ ,
    \new_[2625]_ , \new_[2626]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2630]_ , \new_[2631]_ , \new_[2632]_ ,
    \new_[2633]_ , \new_[2634]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2637]_ , \new_[2638]_ , \new_[2639]_ , \new_[2640]_ ,
    \new_[2641]_ , \new_[2642]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2646]_ , \new_[2647]_ , \new_[2648]_ ,
    \new_[2649]_ , \new_[2650]_ , \new_[2651]_ , \new_[2652]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2657]_ , \new_[2658]_ , \new_[2659]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2724]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2728]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2778]_ , \new_[2779]_ , \new_[2780]_ ,
    \new_[2781]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2843]_ , \new_[2844]_ ,
    \new_[2845]_ , \new_[2846]_ , \new_[2847]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2851]_ , \new_[2852]_ ,
    \new_[2853]_ , \new_[2854]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2862]_ , \new_[2863]_ , \new_[2864]_ ,
    \new_[2865]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2872]_ ,
    \new_[2873]_ , \new_[2874]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2880]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2885]_ , \new_[2886]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2893]_ , \new_[2894]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2902]_ , \new_[2903]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2908]_ ,
    \new_[2909]_ , \new_[2910]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2946]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2949]_ , \new_[2950]_ , \new_[2951]_ , \new_[2952]_ ,
    \new_[2953]_ , \new_[2954]_ , \new_[2955]_ , \new_[2956]_ ,
    \new_[2957]_ , \new_[2958]_ , \new_[2959]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2963]_ , \new_[2964]_ ,
    \new_[2965]_ , \new_[2966]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2970]_ , \new_[2971]_ , \new_[2972]_ ,
    \new_[2973]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2978]_ , \new_[2979]_ , \new_[2980]_ ,
    \new_[2981]_ , \new_[2982]_ , \new_[2983]_ , \new_[2984]_ ,
    \new_[2985]_ , \new_[2986]_ , \new_[2987]_ , \new_[2988]_ ,
    \new_[2989]_ , \new_[2990]_ , \new_[2991]_ , \new_[2992]_ ,
    \new_[2993]_ , \new_[2994]_ , \new_[2995]_ , \new_[2996]_ ,
    \new_[2997]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3004]_ ,
    \new_[3005]_ , \new_[3006]_ , \new_[3007]_ , \new_[3008]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3011]_ , \new_[3012]_ ,
    \new_[3013]_ , \new_[3014]_ , \new_[3015]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3020]_ ,
    \new_[3021]_ , \new_[3022]_ , \new_[3023]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3027]_ , \new_[3028]_ ,
    \new_[3029]_ , \new_[3030]_ , \new_[3031]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3034]_ , \new_[3035]_ , \new_[3036]_ ,
    \new_[3037]_ , \new_[3038]_ , \new_[3039]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3042]_ , \new_[3043]_ , \new_[3044]_ ,
    \new_[3045]_ , \new_[3046]_ , \new_[3047]_ , \new_[3048]_ ,
    \new_[3049]_ , \new_[3050]_ , \new_[3051]_ , \new_[3052]_ ,
    \new_[3053]_ , \new_[3054]_ , \new_[3055]_ , \new_[3056]_ ,
    \new_[3057]_ , \new_[3058]_ , \new_[3059]_ , \new_[3060]_ ,
    \new_[3061]_ , \new_[3062]_ , \new_[3063]_ , \new_[3064]_ ,
    \new_[3065]_ , \new_[3066]_ , \new_[3067]_ , \new_[3068]_ ,
    \new_[3069]_ , \new_[3070]_ , \new_[3071]_ , \new_[3072]_ ,
    \new_[3073]_ , \new_[3074]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3078]_ , \new_[3079]_ , \new_[3080]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3083]_ , \new_[3084]_ ,
    \new_[3085]_ , \new_[3086]_ , \new_[3087]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3091]_ , \new_[3092]_ ,
    \new_[3093]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3109]_ , \new_[3110]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3177]_ , \new_[3178]_ , \new_[3179]_ , \new_[3180]_ ,
    \new_[3181]_ , \new_[3182]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3186]_ , \new_[3187]_ , \new_[3188]_ ,
    \new_[3189]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3198]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3229]_ , \new_[3230]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3233]_ , \new_[3234]_ , \new_[3235]_ , \new_[3236]_ ,
    \new_[3237]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3247]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3252]_ ,
    \new_[3253]_ , \new_[3254]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3258]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3261]_ , \new_[3262]_ , \new_[3263]_ , \new_[3264]_ ,
    \new_[3265]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3269]_ , \new_[3270]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3300]_ ,
    \new_[3301]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3335]_ , \new_[3336]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3341]_ , \new_[3342]_ , \new_[3343]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3526]_ , \new_[3527]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3531]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3534]_ , \new_[3535]_ , \new_[3536]_ ,
    \new_[3537]_ , \new_[3538]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3542]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3546]_ , \new_[3547]_ , \new_[3548]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3557]_ , \new_[3558]_ , \new_[3559]_ , \new_[3560]_ ,
    \new_[3561]_ , \new_[3562]_ , \new_[3563]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3596]_ ,
    \new_[3597]_ , \new_[3598]_ , \new_[3599]_ , \new_[3600]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3604]_ ,
    \new_[3605]_ , \new_[3606]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3610]_ , \new_[3611]_ , \new_[3612]_ ,
    \new_[3613]_ , \new_[3614]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3618]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3622]_ , \new_[3623]_ , \new_[3624]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3629]_ , \new_[3630]_ , \new_[3631]_ , \new_[3632]_ ,
    \new_[3633]_ , \new_[3634]_ , \new_[3635]_ , \new_[3636]_ ,
    \new_[3637]_ , \new_[3638]_ , \new_[3639]_ , \new_[3640]_ ,
    \new_[3641]_ , \new_[3642]_ , \new_[3643]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3654]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3661]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3666]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3669]_ , \new_[3670]_ , \new_[3671]_ , \new_[3672]_ ,
    \new_[3673]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3677]_ , \new_[3678]_ , \new_[3679]_ , \new_[3680]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3683]_ , \new_[3684]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3692]_ ,
    \new_[3693]_ , \new_[3694]_ , \new_[3695]_ , \new_[3696]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3701]_ , \new_[3702]_ , \new_[3703]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3706]_ , \new_[3707]_ , \new_[3708]_ ,
    \new_[3709]_ , \new_[3710]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3716]_ ,
    \new_[3717]_ , \new_[3718]_ , \new_[3719]_ , \new_[3720]_ ,
    \new_[3721]_ , \new_[3722]_ , \new_[3723]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3729]_ , \new_[3730]_ , \new_[3731]_ , \new_[3732]_ ,
    \new_[3733]_ , \new_[3734]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3737]_ , \new_[3738]_ , \new_[3739]_ , \new_[3740]_ ,
    \new_[3741]_ , \new_[3742]_ , \new_[3743]_ , \new_[3744]_ ,
    \new_[3745]_ , \new_[3746]_ , \new_[3747]_ , \new_[3748]_ ,
    \new_[3749]_ , \new_[3750]_ , \new_[3751]_ , \new_[3752]_ ,
    \new_[3753]_ , \new_[3754]_ , \new_[3755]_ , \new_[3756]_ ,
    \new_[3757]_ , \new_[3758]_ , \new_[3759]_ , \new_[3760]_ ,
    \new_[3761]_ , \new_[3762]_ , \new_[3763]_ , \new_[3764]_ ,
    \new_[3765]_ , \new_[3766]_ , \new_[3767]_ , \new_[3768]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3773]_ , \new_[3774]_ , \new_[3775]_ , \new_[3776]_ ,
    \new_[3777]_ , \new_[3778]_ , \new_[3779]_ , \new_[3780]_ ,
    \new_[3781]_ , \new_[3782]_ , \new_[3783]_ , \new_[3784]_ ,
    \new_[3785]_ , \new_[3786]_ , \new_[3787]_ , \new_[3788]_ ,
    \new_[3789]_ , \new_[3790]_ , \new_[3791]_ , \new_[3792]_ ,
    \new_[3793]_ , \new_[3794]_ , \new_[3795]_ , \new_[3796]_ ,
    \new_[3797]_ , \new_[3798]_ , \new_[3799]_ , \new_[3800]_ ,
    \new_[3801]_ , \new_[3802]_ , \new_[3803]_ , \new_[3804]_ ,
    \new_[3805]_ , \new_[3806]_ , \new_[3807]_ , \new_[3808]_ ,
    \new_[3809]_ , \new_[3810]_ , \new_[3811]_ , \new_[3812]_ ,
    \new_[3813]_ , \new_[3814]_ , \new_[3815]_ , \new_[3816]_ ,
    \new_[3817]_ , \new_[3818]_ , \new_[3819]_ , \new_[3820]_ ,
    \new_[3821]_ , \new_[3822]_ , \new_[3823]_ , \new_[3824]_ ,
    \new_[3825]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3829]_ , \new_[3830]_ , \new_[3831]_ , \new_[3832]_ ,
    \new_[3833]_ , \new_[3834]_ , \new_[3835]_ , \new_[3836]_ ,
    \new_[3837]_ , \new_[3838]_ , \new_[3842]_ , \new_[3843]_ ,
    \new_[3846]_ , \new_[3849]_ , \new_[3850]_ , \new_[3851]_ ,
    \new_[3855]_ , \new_[3856]_ , \new_[3859]_ , \new_[3862]_ ,
    \new_[3863]_ , \new_[3864]_ , \new_[3865]_ , \new_[3869]_ ,
    \new_[3870]_ , \new_[3873]_ , \new_[3876]_ , \new_[3877]_ ,
    \new_[3878]_ , \new_[3881]_ , \new_[3884]_ , \new_[3885]_ ,
    \new_[3888]_ , \new_[3891]_ , \new_[3892]_ , \new_[3893]_ ,
    \new_[3894]_ , \new_[3895]_ , \new_[3899]_ , \new_[3900]_ ,
    \new_[3903]_ , \new_[3906]_ , \new_[3907]_ , \new_[3908]_ ,
    \new_[3911]_ , \new_[3914]_ , \new_[3915]_ , \new_[3918]_ ,
    \new_[3921]_ , \new_[3922]_ , \new_[3923]_ , \new_[3924]_ ,
    \new_[3928]_ , \new_[3929]_ , \new_[3932]_ , \new_[3935]_ ,
    \new_[3936]_ , \new_[3937]_ , \new_[3940]_ , \new_[3943]_ ,
    \new_[3944]_ , \new_[3947]_ , \new_[3950]_ , \new_[3951]_ ,
    \new_[3952]_ , \new_[3953]_ , \new_[3954]_ , \new_[3955]_ ,
    \new_[3959]_ , \new_[3960]_ , \new_[3963]_ , \new_[3966]_ ,
    \new_[3967]_ , \new_[3968]_ , \new_[3971]_ , \new_[3974]_ ,
    \new_[3975]_ , \new_[3978]_ , \new_[3981]_ , \new_[3982]_ ,
    \new_[3983]_ , \new_[3984]_ , \new_[3988]_ , \new_[3989]_ ,
    \new_[3992]_ , \new_[3995]_ , \new_[3996]_ , \new_[3997]_ ,
    \new_[4000]_ , \new_[4003]_ , \new_[4004]_ , \new_[4007]_ ,
    \new_[4010]_ , \new_[4011]_ , \new_[4012]_ , \new_[4013]_ ,
    \new_[4014]_ , \new_[4018]_ , \new_[4019]_ , \new_[4022]_ ,
    \new_[4025]_ , \new_[4026]_ , \new_[4027]_ , \new_[4030]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4037]_ , \new_[4040]_ ,
    \new_[4041]_ , \new_[4042]_ , \new_[4043]_ , \new_[4047]_ ,
    \new_[4048]_ , \new_[4051]_ , \new_[4054]_ , \new_[4055]_ ,
    \new_[4056]_ , \new_[4059]_ , \new_[4062]_ , \new_[4063]_ ,
    \new_[4066]_ , \new_[4069]_ , \new_[4070]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4074]_ , \new_[4075]_ ,
    \new_[4079]_ , \new_[4080]_ , \new_[4083]_ , \new_[4086]_ ,
    \new_[4087]_ , \new_[4088]_ , \new_[4091]_ , \new_[4094]_ ,
    \new_[4095]_ , \new_[4098]_ , \new_[4101]_ , \new_[4102]_ ,
    \new_[4103]_ , \new_[4104]_ , \new_[4108]_ , \new_[4109]_ ,
    \new_[4112]_ , \new_[4115]_ , \new_[4116]_ , \new_[4117]_ ,
    \new_[4120]_ , \new_[4123]_ , \new_[4124]_ , \new_[4127]_ ,
    \new_[4130]_ , \new_[4131]_ , \new_[4132]_ , \new_[4133]_ ,
    \new_[4134]_ , \new_[4138]_ , \new_[4139]_ , \new_[4142]_ ,
    \new_[4145]_ , \new_[4146]_ , \new_[4147]_ , \new_[4150]_ ,
    \new_[4153]_ , \new_[4154]_ , \new_[4157]_ , \new_[4160]_ ,
    \new_[4161]_ , \new_[4162]_ , \new_[4163]_ , \new_[4167]_ ,
    \new_[4168]_ , \new_[4171]_ , \new_[4174]_ , \new_[4175]_ ,
    \new_[4176]_ , \new_[4179]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4186]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4192]_ , \new_[4193]_ , \new_[4194]_ , \new_[4198]_ ,
    \new_[4199]_ , \new_[4202]_ , \new_[4205]_ , \new_[4206]_ ,
    \new_[4207]_ , \new_[4210]_ , \new_[4213]_ , \new_[4214]_ ,
    \new_[4217]_ , \new_[4220]_ , \new_[4221]_ , \new_[4222]_ ,
    \new_[4223]_ , \new_[4227]_ , \new_[4228]_ , \new_[4231]_ ,
    \new_[4234]_ , \new_[4235]_ , \new_[4236]_ , \new_[4239]_ ,
    \new_[4242]_ , \new_[4243]_ , \new_[4246]_ , \new_[4249]_ ,
    \new_[4250]_ , \new_[4251]_ , \new_[4252]_ , \new_[4253]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4261]_ , \new_[4264]_ ,
    \new_[4265]_ , \new_[4266]_ , \new_[4269]_ , \new_[4272]_ ,
    \new_[4273]_ , \new_[4276]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4286]_ , \new_[4287]_ ,
    \new_[4290]_ , \new_[4293]_ , \new_[4294]_ , \new_[4295]_ ,
    \new_[4298]_ , \new_[4301]_ , \new_[4302]_ , \new_[4305]_ ,
    \new_[4308]_ , \new_[4309]_ , \new_[4310]_ , \new_[4311]_ ,
    \new_[4312]_ , \new_[4313]_ , \new_[4314]_ , \new_[4315]_ ,
    \new_[4319]_ , \new_[4320]_ , \new_[4323]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4328]_ , \new_[4331]_ , \new_[4334]_ ,
    \new_[4335]_ , \new_[4338]_ , \new_[4341]_ , \new_[4342]_ ,
    \new_[4343]_ , \new_[4344]_ , \new_[4348]_ , \new_[4349]_ ,
    \new_[4352]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4360]_ , \new_[4363]_ , \new_[4364]_ , \new_[4367]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4372]_ , \new_[4373]_ ,
    \new_[4374]_ , \new_[4378]_ , \new_[4379]_ , \new_[4382]_ ,
    \new_[4385]_ , \new_[4386]_ , \new_[4387]_ , \new_[4390]_ ,
    \new_[4393]_ , \new_[4394]_ , \new_[4397]_ , \new_[4400]_ ,
    \new_[4401]_ , \new_[4402]_ , \new_[4403]_ , \new_[4407]_ ,
    \new_[4408]_ , \new_[4411]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4416]_ , \new_[4419]_ , \new_[4422]_ , \new_[4423]_ ,
    \new_[4426]_ , \new_[4429]_ , \new_[4430]_ , \new_[4431]_ ,
    \new_[4432]_ , \new_[4433]_ , \new_[4434]_ , \new_[4438]_ ,
    \new_[4439]_ , \new_[4442]_ , \new_[4445]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4450]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4457]_ , \new_[4460]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4467]_ , \new_[4468]_ , \new_[4471]_ ,
    \new_[4474]_ , \new_[4475]_ , \new_[4476]_ , \new_[4479]_ ,
    \new_[4482]_ , \new_[4483]_ , \new_[4486]_ , \new_[4489]_ ,
    \new_[4490]_ , \new_[4491]_ , \new_[4492]_ , \new_[4493]_ ,
    \new_[4497]_ , \new_[4498]_ , \new_[4501]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4509]_ , \new_[4512]_ ,
    \new_[4513]_ , \new_[4516]_ , \new_[4519]_ , \new_[4520]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4526]_ , \new_[4527]_ ,
    \new_[4530]_ , \new_[4533]_ , \new_[4534]_ , \new_[4535]_ ,
    \new_[4538]_ , \new_[4541]_ , \new_[4542]_ , \new_[4545]_ ,
    \new_[4548]_ , \new_[4549]_ , \new_[4550]_ , \new_[4551]_ ,
    \new_[4552]_ , \new_[4553]_ , \new_[4554]_ , \new_[4558]_ ,
    \new_[4559]_ , \new_[4562]_ , \new_[4565]_ , \new_[4566]_ ,
    \new_[4567]_ , \new_[4570]_ , \new_[4573]_ , \new_[4574]_ ,
    \new_[4577]_ , \new_[4580]_ , \new_[4581]_ , \new_[4582]_ ,
    \new_[4583]_ , \new_[4587]_ , \new_[4588]_ , \new_[4591]_ ,
    \new_[4594]_ , \new_[4595]_ , \new_[4596]_ , \new_[4599]_ ,
    \new_[4602]_ , \new_[4603]_ , \new_[4606]_ , \new_[4609]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4612]_ , \new_[4613]_ ,
    \new_[4617]_ , \new_[4618]_ , \new_[4621]_ , \new_[4624]_ ,
    \new_[4625]_ , \new_[4626]_ , \new_[4629]_ , \new_[4632]_ ,
    \new_[4633]_ , \new_[4636]_ , \new_[4639]_ , \new_[4640]_ ,
    \new_[4641]_ , \new_[4642]_ , \new_[4646]_ , \new_[4647]_ ,
    \new_[4650]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4658]_ , \new_[4661]_ , \new_[4662]_ , \new_[4665]_ ,
    \new_[4668]_ , \new_[4669]_ , \new_[4670]_ , \new_[4671]_ ,
    \new_[4672]_ , \new_[4673]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4681]_ , \new_[4684]_ , \new_[4685]_ , \new_[4686]_ ,
    \new_[4689]_ , \new_[4692]_ , \new_[4693]_ , \new_[4696]_ ,
    \new_[4699]_ , \new_[4700]_ , \new_[4701]_ , \new_[4702]_ ,
    \new_[4706]_ , \new_[4707]_ , \new_[4710]_ , \new_[4713]_ ,
    \new_[4714]_ , \new_[4715]_ , \new_[4718]_ , \new_[4721]_ ,
    \new_[4722]_ , \new_[4725]_ , \new_[4728]_ , \new_[4729]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4732]_ , \new_[4736]_ ,
    \new_[4737]_ , \new_[4740]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4748]_ , \new_[4751]_ , \new_[4752]_ ,
    \new_[4755]_ , \new_[4758]_ , \new_[4759]_ , \new_[4760]_ ,
    \new_[4761]_ , \new_[4765]_ , \new_[4766]_ , \new_[4769]_ ,
    \new_[4772]_ , \new_[4773]_ , \new_[4774]_ , \new_[4777]_ ,
    \new_[4780]_ , \new_[4781]_ , \new_[4784]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4789]_ , \new_[4790]_ , \new_[4791]_ ,
    \new_[4792]_ , \new_[4793]_ , \new_[4794]_ , \new_[4795]_ ,
    \new_[4799]_ , \new_[4800]_ , \new_[4803]_ , \new_[4806]_ ,
    \new_[4807]_ , \new_[4808]_ , \new_[4811]_ , \new_[4814]_ ,
    \new_[4815]_ , \new_[4818]_ , \new_[4821]_ , \new_[4822]_ ,
    \new_[4823]_ , \new_[4824]_ , \new_[4828]_ , \new_[4829]_ ,
    \new_[4832]_ , \new_[4835]_ , \new_[4836]_ , \new_[4837]_ ,
    \new_[4840]_ , \new_[4843]_ , \new_[4844]_ , \new_[4847]_ ,
    \new_[4850]_ , \new_[4851]_ , \new_[4852]_ , \new_[4853]_ ,
    \new_[4854]_ , \new_[4858]_ , \new_[4859]_ , \new_[4862]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4870]_ ,
    \new_[4873]_ , \new_[4874]_ , \new_[4877]_ , \new_[4880]_ ,
    \new_[4881]_ , \new_[4882]_ , \new_[4883]_ , \new_[4887]_ ,
    \new_[4888]_ , \new_[4891]_ , \new_[4894]_ , \new_[4895]_ ,
    \new_[4896]_ , \new_[4899]_ , \new_[4902]_ , \new_[4903]_ ,
    \new_[4906]_ , \new_[4909]_ , \new_[4910]_ , \new_[4911]_ ,
    \new_[4912]_ , \new_[4913]_ , \new_[4914]_ , \new_[4918]_ ,
    \new_[4919]_ , \new_[4922]_ , \new_[4925]_ , \new_[4926]_ ,
    \new_[4927]_ , \new_[4930]_ , \new_[4933]_ , \new_[4934]_ ,
    \new_[4937]_ , \new_[4940]_ , \new_[4941]_ , \new_[4942]_ ,
    \new_[4943]_ , \new_[4947]_ , \new_[4948]_ , \new_[4951]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4956]_ , \new_[4959]_ ,
    \new_[4962]_ , \new_[4963]_ , \new_[4966]_ , \new_[4969]_ ,
    \new_[4970]_ , \new_[4971]_ , \new_[4972]_ , \new_[4973]_ ,
    \new_[4977]_ , \new_[4978]_ , \new_[4981]_ , \new_[4984]_ ,
    \new_[4985]_ , \new_[4986]_ , \new_[4989]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4996]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5006]_ , \new_[5007]_ ,
    \new_[5010]_ , \new_[5013]_ , \new_[5014]_ , \new_[5015]_ ,
    \new_[5018]_ , \new_[5021]_ , \new_[5022]_ , \new_[5025]_ ,
    \new_[5028]_ , \new_[5029]_ , \new_[5030]_ , \new_[5031]_ ,
    \new_[5032]_ , \new_[5033]_ , \new_[5034]_ , \new_[5038]_ ,
    \new_[5039]_ , \new_[5042]_ , \new_[5045]_ , \new_[5046]_ ,
    \new_[5047]_ , \new_[5050]_ , \new_[5053]_ , \new_[5054]_ ,
    \new_[5057]_ , \new_[5060]_ , \new_[5061]_ , \new_[5062]_ ,
    \new_[5063]_ , \new_[5067]_ , \new_[5068]_ , \new_[5071]_ ,
    \new_[5074]_ , \new_[5075]_ , \new_[5076]_ , \new_[5079]_ ,
    \new_[5082]_ , \new_[5083]_ , \new_[5086]_ , \new_[5089]_ ,
    \new_[5090]_ , \new_[5091]_ , \new_[5092]_ , \new_[5093]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5101]_ , \new_[5104]_ ,
    \new_[5105]_ , \new_[5106]_ , \new_[5109]_ , \new_[5112]_ ,
    \new_[5113]_ , \new_[5116]_ , \new_[5119]_ , \new_[5120]_ ,
    \new_[5121]_ , \new_[5122]_ , \new_[5126]_ , \new_[5127]_ ,
    \new_[5130]_ , \new_[5133]_ , \new_[5134]_ , \new_[5135]_ ,
    \new_[5138]_ , \new_[5141]_ , \new_[5142]_ , \new_[5145]_ ,
    \new_[5148]_ , \new_[5149]_ , \new_[5150]_ , \new_[5151]_ ,
    \new_[5152]_ , \new_[5153]_ , \new_[5157]_ , \new_[5158]_ ,
    \new_[5161]_ , \new_[5164]_ , \new_[5165]_ , \new_[5166]_ ,
    \new_[5169]_ , \new_[5172]_ , \new_[5173]_ , \new_[5176]_ ,
    \new_[5179]_ , \new_[5180]_ , \new_[5181]_ , \new_[5182]_ ,
    \new_[5186]_ , \new_[5187]_ , \new_[5190]_ , \new_[5193]_ ,
    \new_[5194]_ , \new_[5195]_ , \new_[5198]_ , \new_[5201]_ ,
    \new_[5202]_ , \new_[5205]_ , \new_[5208]_ , \new_[5209]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5212]_ , \new_[5216]_ ,
    \new_[5217]_ , \new_[5220]_ , \new_[5223]_ , \new_[5224]_ ,
    \new_[5225]_ , \new_[5228]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5235]_ , \new_[5238]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5245]_ , \new_[5246]_ , \new_[5249]_ ,
    \new_[5252]_ , \new_[5253]_ , \new_[5254]_ , \new_[5257]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5264]_ , \new_[5267]_ ,
    \new_[5268]_ , \new_[5269]_ , \new_[5270]_ , \new_[5271]_ ,
    \new_[5272]_ , \new_[5273]_ , \new_[5274]_ , \new_[5278]_ ,
    \new_[5279]_ , \new_[5282]_ , \new_[5285]_ , \new_[5286]_ ,
    \new_[5287]_ , \new_[5290]_ , \new_[5293]_ , \new_[5294]_ ,
    \new_[5297]_ , \new_[5300]_ , \new_[5301]_ , \new_[5302]_ ,
    \new_[5303]_ , \new_[5307]_ , \new_[5308]_ , \new_[5311]_ ,
    \new_[5314]_ , \new_[5315]_ , \new_[5316]_ , \new_[5319]_ ,
    \new_[5322]_ , \new_[5323]_ , \new_[5326]_ , \new_[5329]_ ,
    \new_[5330]_ , \new_[5331]_ , \new_[5332]_ , \new_[5333]_ ,
    \new_[5337]_ , \new_[5338]_ , \new_[5341]_ , \new_[5344]_ ,
    \new_[5345]_ , \new_[5346]_ , \new_[5349]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5356]_ , \new_[5359]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5362]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5370]_ , \new_[5373]_ , \new_[5374]_ , \new_[5375]_ ,
    \new_[5378]_ , \new_[5381]_ , \new_[5382]_ , \new_[5385]_ ,
    \new_[5388]_ , \new_[5389]_ , \new_[5390]_ , \new_[5391]_ ,
    \new_[5392]_ , \new_[5393]_ , \new_[5397]_ , \new_[5398]_ ,
    \new_[5401]_ , \new_[5404]_ , \new_[5405]_ , \new_[5406]_ ,
    \new_[5409]_ , \new_[5412]_ , \new_[5413]_ , \new_[5416]_ ,
    \new_[5419]_ , \new_[5420]_ , \new_[5421]_ , \new_[5422]_ ,
    \new_[5426]_ , \new_[5427]_ , \new_[5430]_ , \new_[5433]_ ,
    \new_[5434]_ , \new_[5435]_ , \new_[5438]_ , \new_[5441]_ ,
    \new_[5442]_ , \new_[5445]_ , \new_[5448]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5451]_ , \new_[5452]_ , \new_[5456]_ ,
    \new_[5457]_ , \new_[5460]_ , \new_[5463]_ , \new_[5464]_ ,
    \new_[5465]_ , \new_[5468]_ , \new_[5471]_ , \new_[5472]_ ,
    \new_[5475]_ , \new_[5478]_ , \new_[5479]_ , \new_[5480]_ ,
    \new_[5481]_ , \new_[5485]_ , \new_[5486]_ , \new_[5489]_ ,
    \new_[5492]_ , \new_[5493]_ , \new_[5494]_ , \new_[5497]_ ,
    \new_[5500]_ , \new_[5501]_ , \new_[5504]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5513]_ , \new_[5517]_ , \new_[5518]_ ,
    \new_[5521]_ , \new_[5524]_ , \new_[5525]_ , \new_[5526]_ ,
    \new_[5529]_ , \new_[5532]_ , \new_[5533]_ , \new_[5536]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5541]_ , \new_[5542]_ ,
    \new_[5546]_ , \new_[5547]_ , \new_[5550]_ , \new_[5553]_ ,
    \new_[5554]_ , \new_[5555]_ , \new_[5558]_ , \new_[5561]_ ,
    \new_[5562]_ , \new_[5565]_ , \new_[5568]_ , \new_[5569]_ ,
    \new_[5570]_ , \new_[5571]_ , \new_[5572]_ , \new_[5576]_ ,
    \new_[5577]_ , \new_[5580]_ , \new_[5583]_ , \new_[5584]_ ,
    \new_[5585]_ , \new_[5588]_ , \new_[5591]_ , \new_[5592]_ ,
    \new_[5595]_ , \new_[5598]_ , \new_[5599]_ , \new_[5600]_ ,
    \new_[5601]_ , \new_[5605]_ , \new_[5606]_ , \new_[5609]_ ,
    \new_[5612]_ , \new_[5613]_ , \new_[5614]_ , \new_[5617]_ ,
    \new_[5620]_ , \new_[5621]_ , \new_[5624]_ , \new_[5627]_ ,
    \new_[5628]_ , \new_[5629]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5632]_ , \new_[5636]_ , \new_[5637]_ , \new_[5640]_ ,
    \new_[5643]_ , \new_[5644]_ , \new_[5645]_ , \new_[5648]_ ,
    \new_[5651]_ , \new_[5652]_ , \new_[5655]_ , \new_[5658]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5661]_ , \new_[5665]_ ,
    \new_[5666]_ , \new_[5669]_ , \new_[5672]_ , \new_[5673]_ ,
    \new_[5674]_ , \new_[5677]_ , \new_[5680]_ , \new_[5681]_ ,
    \new_[5684]_ , \new_[5687]_ , \new_[5688]_ , \new_[5689]_ ,
    \new_[5690]_ , \new_[5691]_ , \new_[5695]_ , \new_[5696]_ ,
    \new_[5699]_ , \new_[5702]_ , \new_[5703]_ , \new_[5704]_ ,
    \new_[5707]_ , \new_[5710]_ , \new_[5711]_ , \new_[5714]_ ,
    \new_[5717]_ , \new_[5718]_ , \new_[5719]_ , \new_[5720]_ ,
    \new_[5724]_ , \new_[5725]_ , \new_[5728]_ , \new_[5731]_ ,
    \new_[5732]_ , \new_[5733]_ , \new_[5736]_ , \new_[5739]_ ,
    \new_[5740]_ , \new_[5743]_ , \new_[5746]_ , \new_[5747]_ ,
    \new_[5748]_ , \new_[5749]_ , \new_[5750]_ , \new_[5751]_ ,
    \new_[5752]_ , \new_[5753]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5759]_ , \new_[5760]_ , \new_[5763]_ , \new_[5766]_ ,
    \new_[5767]_ , \new_[5768]_ , \new_[5771]_ , \new_[5774]_ ,
    \new_[5775]_ , \new_[5778]_ , \new_[5781]_ , \new_[5782]_ ,
    \new_[5783]_ , \new_[5784]_ , \new_[5788]_ , \new_[5789]_ ,
    \new_[5792]_ , \new_[5795]_ , \new_[5796]_ , \new_[5797]_ ,
    \new_[5800]_ , \new_[5803]_ , \new_[5804]_ , \new_[5807]_ ,
    \new_[5810]_ , \new_[5811]_ , \new_[5812]_ , \new_[5813]_ ,
    \new_[5814]_ , \new_[5818]_ , \new_[5819]_ , \new_[5822]_ ,
    \new_[5825]_ , \new_[5826]_ , \new_[5827]_ , \new_[5830]_ ,
    \new_[5833]_ , \new_[5834]_ , \new_[5837]_ , \new_[5840]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5843]_ , \new_[5847]_ ,
    \new_[5848]_ , \new_[5851]_ , \new_[5854]_ , \new_[5855]_ ,
    \new_[5856]_ , \new_[5859]_ , \new_[5862]_ , \new_[5863]_ ,
    \new_[5866]_ , \new_[5869]_ , \new_[5870]_ , \new_[5871]_ ,
    \new_[5872]_ , \new_[5873]_ , \new_[5874]_ , \new_[5878]_ ,
    \new_[5879]_ , \new_[5882]_ , \new_[5885]_ , \new_[5886]_ ,
    \new_[5887]_ , \new_[5890]_ , \new_[5893]_ , \new_[5894]_ ,
    \new_[5897]_ , \new_[5900]_ , \new_[5901]_ , \new_[5902]_ ,
    \new_[5903]_ , \new_[5907]_ , \new_[5908]_ , \new_[5911]_ ,
    \new_[5914]_ , \new_[5915]_ , \new_[5916]_ , \new_[5919]_ ,
    \new_[5922]_ , \new_[5923]_ , \new_[5926]_ , \new_[5929]_ ,
    \new_[5930]_ , \new_[5931]_ , \new_[5932]_ , \new_[5933]_ ,
    \new_[5937]_ , \new_[5938]_ , \new_[5941]_ , \new_[5944]_ ,
    \new_[5945]_ , \new_[5946]_ , \new_[5949]_ , \new_[5952]_ ,
    \new_[5953]_ , \new_[5956]_ , \new_[5959]_ , \new_[5960]_ ,
    \new_[5961]_ , \new_[5962]_ , \new_[5966]_ , \new_[5967]_ ,
    \new_[5970]_ , \new_[5973]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5978]_ , \new_[5981]_ , \new_[5982]_ , \new_[5985]_ ,
    \new_[5988]_ , \new_[5989]_ , \new_[5990]_ , \new_[5991]_ ,
    \new_[5992]_ , \new_[5993]_ , \new_[5994]_ , \new_[5998]_ ,
    \new_[5999]_ , \new_[6002]_ , \new_[6005]_ , \new_[6006]_ ,
    \new_[6007]_ , \new_[6010]_ , \new_[6013]_ , \new_[6014]_ ,
    \new_[6017]_ , \new_[6020]_ , \new_[6021]_ , \new_[6022]_ ,
    \new_[6023]_ , \new_[6027]_ , \new_[6028]_ , \new_[6031]_ ,
    \new_[6034]_ , \new_[6035]_ , \new_[6036]_ , \new_[6039]_ ,
    \new_[6042]_ , \new_[6043]_ , \new_[6046]_ , \new_[6049]_ ,
    \new_[6050]_ , \new_[6051]_ , \new_[6052]_ , \new_[6053]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6061]_ , \new_[6064]_ ,
    \new_[6065]_ , \new_[6066]_ , \new_[6069]_ , \new_[6072]_ ,
    \new_[6073]_ , \new_[6076]_ , \new_[6079]_ , \new_[6080]_ ,
    \new_[6081]_ , \new_[6082]_ , \new_[6086]_ , \new_[6087]_ ,
    \new_[6090]_ , \new_[6093]_ , \new_[6094]_ , \new_[6095]_ ,
    \new_[6098]_ , \new_[6101]_ , \new_[6102]_ , \new_[6105]_ ,
    \new_[6108]_ , \new_[6109]_ , \new_[6110]_ , \new_[6111]_ ,
    \new_[6112]_ , \new_[6113]_ , \new_[6117]_ , \new_[6118]_ ,
    \new_[6121]_ , \new_[6124]_ , \new_[6125]_ , \new_[6126]_ ,
    \new_[6129]_ , \new_[6132]_ , \new_[6133]_ , \new_[6136]_ ,
    \new_[6139]_ , \new_[6140]_ , \new_[6141]_ , \new_[6142]_ ,
    \new_[6146]_ , \new_[6147]_ , \new_[6150]_ , \new_[6153]_ ,
    \new_[6154]_ , \new_[6155]_ , \new_[6158]_ , \new_[6161]_ ,
    \new_[6162]_ , \new_[6165]_ , \new_[6168]_ , \new_[6169]_ ,
    \new_[6170]_ , \new_[6171]_ , \new_[6172]_ , \new_[6176]_ ,
    \new_[6177]_ , \new_[6180]_ , \new_[6183]_ , \new_[6184]_ ,
    \new_[6185]_ , \new_[6188]_ , \new_[6191]_ , \new_[6192]_ ,
    \new_[6195]_ , \new_[6198]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6201]_ , \new_[6205]_ , \new_[6206]_ , \new_[6209]_ ,
    \new_[6212]_ , \new_[6213]_ , \new_[6214]_ , \new_[6217]_ ,
    \new_[6220]_ , \new_[6221]_ , \new_[6224]_ , \new_[6227]_ ,
    \new_[6228]_ , \new_[6229]_ , \new_[6230]_ , \new_[6231]_ ,
    \new_[6232]_ , \new_[6233]_ , \new_[6234]_ , \new_[6238]_ ,
    \new_[6239]_ , \new_[6242]_ , \new_[6245]_ , \new_[6246]_ ,
    \new_[6247]_ , \new_[6250]_ , \new_[6253]_ , \new_[6254]_ ,
    \new_[6257]_ , \new_[6260]_ , \new_[6261]_ , \new_[6262]_ ,
    \new_[6263]_ , \new_[6267]_ , \new_[6268]_ , \new_[6271]_ ,
    \new_[6274]_ , \new_[6275]_ , \new_[6276]_ , \new_[6279]_ ,
    \new_[6282]_ , \new_[6283]_ , \new_[6286]_ , \new_[6289]_ ,
    \new_[6290]_ , \new_[6291]_ , \new_[6292]_ , \new_[6293]_ ,
    \new_[6297]_ , \new_[6298]_ , \new_[6301]_ , \new_[6304]_ ,
    \new_[6305]_ , \new_[6306]_ , \new_[6309]_ , \new_[6312]_ ,
    \new_[6313]_ , \new_[6316]_ , \new_[6319]_ , \new_[6320]_ ,
    \new_[6321]_ , \new_[6322]_ , \new_[6326]_ , \new_[6327]_ ,
    \new_[6330]_ , \new_[6333]_ , \new_[6334]_ , \new_[6335]_ ,
    \new_[6338]_ , \new_[6341]_ , \new_[6342]_ , \new_[6345]_ ,
    \new_[6348]_ , \new_[6349]_ , \new_[6350]_ , \new_[6351]_ ,
    \new_[6352]_ , \new_[6353]_ , \new_[6357]_ , \new_[6358]_ ,
    \new_[6361]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6369]_ , \new_[6372]_ , \new_[6373]_ , \new_[6376]_ ,
    \new_[6379]_ , \new_[6380]_ , \new_[6381]_ , \new_[6382]_ ,
    \new_[6386]_ , \new_[6387]_ , \new_[6390]_ , \new_[6393]_ ,
    \new_[6394]_ , \new_[6395]_ , \new_[6398]_ , \new_[6401]_ ,
    \new_[6402]_ , \new_[6405]_ , \new_[6408]_ , \new_[6409]_ ,
    \new_[6410]_ , \new_[6411]_ , \new_[6412]_ , \new_[6416]_ ,
    \new_[6417]_ , \new_[6420]_ , \new_[6423]_ , \new_[6424]_ ,
    \new_[6425]_ , \new_[6428]_ , \new_[6431]_ , \new_[6432]_ ,
    \new_[6435]_ , \new_[6438]_ , \new_[6439]_ , \new_[6440]_ ,
    \new_[6441]_ , \new_[6445]_ , \new_[6446]_ , \new_[6449]_ ,
    \new_[6452]_ , \new_[6453]_ , \new_[6454]_ , \new_[6457]_ ,
    \new_[6460]_ , \new_[6461]_ , \new_[6464]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6470]_ , \new_[6471]_ ,
    \new_[6472]_ , \new_[6473]_ , \new_[6477]_ , \new_[6478]_ ,
    \new_[6481]_ , \new_[6484]_ , \new_[6485]_ , \new_[6486]_ ,
    \new_[6489]_ , \new_[6492]_ , \new_[6493]_ , \new_[6496]_ ,
    \new_[6499]_ , \new_[6500]_ , \new_[6501]_ , \new_[6502]_ ,
    \new_[6506]_ , \new_[6507]_ , \new_[6510]_ , \new_[6513]_ ,
    \new_[6514]_ , \new_[6515]_ , \new_[6518]_ , \new_[6521]_ ,
    \new_[6522]_ , \new_[6525]_ , \new_[6528]_ , \new_[6529]_ ,
    \new_[6530]_ , \new_[6531]_ , \new_[6532]_ , \new_[6536]_ ,
    \new_[6537]_ , \new_[6540]_ , \new_[6543]_ , \new_[6544]_ ,
    \new_[6545]_ , \new_[6548]_ , \new_[6551]_ , \new_[6552]_ ,
    \new_[6555]_ , \new_[6558]_ , \new_[6559]_ , \new_[6560]_ ,
    \new_[6561]_ , \new_[6565]_ , \new_[6566]_ , \new_[6569]_ ,
    \new_[6572]_ , \new_[6573]_ , \new_[6574]_ , \new_[6577]_ ,
    \new_[6580]_ , \new_[6581]_ , \new_[6584]_ , \new_[6587]_ ,
    \new_[6588]_ , \new_[6589]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6592]_ , \new_[6596]_ , \new_[6597]_ , \new_[6600]_ ,
    \new_[6603]_ , \new_[6604]_ , \new_[6605]_ , \new_[6608]_ ,
    \new_[6611]_ , \new_[6612]_ , \new_[6615]_ , \new_[6618]_ ,
    \new_[6619]_ , \new_[6620]_ , \new_[6621]_ , \new_[6625]_ ,
    \new_[6626]_ , \new_[6629]_ , \new_[6632]_ , \new_[6633]_ ,
    \new_[6634]_ , \new_[6637]_ , \new_[6640]_ , \new_[6641]_ ,
    \new_[6644]_ , \new_[6647]_ , \new_[6648]_ , \new_[6649]_ ,
    \new_[6650]_ , \new_[6651]_ , \new_[6655]_ , \new_[6656]_ ,
    \new_[6659]_ , \new_[6662]_ , \new_[6663]_ , \new_[6664]_ ,
    \new_[6667]_ , \new_[6670]_ , \new_[6671]_ , \new_[6674]_ ,
    \new_[6677]_ , \new_[6678]_ , \new_[6679]_ , \new_[6680]_ ,
    \new_[6684]_ , \new_[6685]_ , \new_[6688]_ , \new_[6691]_ ,
    \new_[6692]_ , \new_[6693]_ , \new_[6696]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6703]_ , \new_[6706]_ , \new_[6707]_ ,
    \new_[6708]_ , \new_[6709]_ , \new_[6710]_ , \new_[6711]_ ,
    \new_[6712]_ , \new_[6713]_ , \new_[6714]_ , \new_[6718]_ ,
    \new_[6719]_ , \new_[6722]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6727]_ , \new_[6730]_ , \new_[6733]_ , \new_[6734]_ ,
    \new_[6737]_ , \new_[6740]_ , \new_[6741]_ , \new_[6742]_ ,
    \new_[6743]_ , \new_[6747]_ , \new_[6748]_ , \new_[6751]_ ,
    \new_[6754]_ , \new_[6755]_ , \new_[6756]_ , \new_[6759]_ ,
    \new_[6762]_ , \new_[6763]_ , \new_[6766]_ , \new_[6769]_ ,
    \new_[6770]_ , \new_[6771]_ , \new_[6772]_ , \new_[6773]_ ,
    \new_[6777]_ , \new_[6778]_ , \new_[6781]_ , \new_[6784]_ ,
    \new_[6785]_ , \new_[6786]_ , \new_[6789]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6796]_ , \new_[6799]_ , \new_[6800]_ ,
    \new_[6801]_ , \new_[6802]_ , \new_[6806]_ , \new_[6807]_ ,
    \new_[6810]_ , \new_[6813]_ , \new_[6814]_ , \new_[6815]_ ,
    \new_[6818]_ , \new_[6821]_ , \new_[6822]_ , \new_[6825]_ ,
    \new_[6828]_ , \new_[6829]_ , \new_[6830]_ , \new_[6831]_ ,
    \new_[6832]_ , \new_[6833]_ , \new_[6837]_ , \new_[6838]_ ,
    \new_[6841]_ , \new_[6844]_ , \new_[6845]_ , \new_[6846]_ ,
    \new_[6849]_ , \new_[6852]_ , \new_[6853]_ , \new_[6856]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6861]_ , \new_[6862]_ ,
    \new_[6866]_ , \new_[6867]_ , \new_[6870]_ , \new_[6873]_ ,
    \new_[6874]_ , \new_[6875]_ , \new_[6878]_ , \new_[6881]_ ,
    \new_[6882]_ , \new_[6885]_ , \new_[6888]_ , \new_[6889]_ ,
    \new_[6890]_ , \new_[6891]_ , \new_[6892]_ , \new_[6896]_ ,
    \new_[6897]_ , \new_[6900]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6905]_ , \new_[6908]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6915]_ , \new_[6918]_ , \new_[6919]_ , \new_[6920]_ ,
    \new_[6921]_ , \new_[6925]_ , \new_[6926]_ , \new_[6929]_ ,
    \new_[6932]_ , \new_[6933]_ , \new_[6934]_ , \new_[6937]_ ,
    \new_[6940]_ , \new_[6941]_ , \new_[6944]_ , \new_[6947]_ ,
    \new_[6948]_ , \new_[6949]_ , \new_[6950]_ , \new_[6951]_ ,
    \new_[6952]_ , \new_[6953]_ , \new_[6957]_ , \new_[6958]_ ,
    \new_[6961]_ , \new_[6964]_ , \new_[6965]_ , \new_[6966]_ ,
    \new_[6969]_ , \new_[6972]_ , \new_[6973]_ , \new_[6976]_ ,
    \new_[6979]_ , \new_[6980]_ , \new_[6981]_ , \new_[6982]_ ,
    \new_[6986]_ , \new_[6987]_ , \new_[6990]_ , \new_[6993]_ ,
    \new_[6994]_ , \new_[6995]_ , \new_[6998]_ , \new_[7001]_ ,
    \new_[7002]_ , \new_[7005]_ , \new_[7008]_ , \new_[7009]_ ,
    \new_[7010]_ , \new_[7011]_ , \new_[7012]_ , \new_[7016]_ ,
    \new_[7017]_ , \new_[7020]_ , \new_[7023]_ , \new_[7024]_ ,
    \new_[7025]_ , \new_[7028]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7035]_ , \new_[7038]_ , \new_[7039]_ , \new_[7040]_ ,
    \new_[7041]_ , \new_[7045]_ , \new_[7046]_ , \new_[7049]_ ,
    \new_[7052]_ , \new_[7053]_ , \new_[7054]_ , \new_[7057]_ ,
    \new_[7060]_ , \new_[7061]_ , \new_[7064]_ , \new_[7067]_ ,
    \new_[7068]_ , \new_[7069]_ , \new_[7070]_ , \new_[7071]_ ,
    \new_[7072]_ , \new_[7076]_ , \new_[7077]_ , \new_[7080]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7085]_ , \new_[7088]_ ,
    \new_[7091]_ , \new_[7092]_ , \new_[7095]_ , \new_[7098]_ ,
    \new_[7099]_ , \new_[7100]_ , \new_[7101]_ , \new_[7105]_ ,
    \new_[7106]_ , \new_[7109]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7114]_ , \new_[7117]_ , \new_[7120]_ , \new_[7121]_ ,
    \new_[7124]_ , \new_[7127]_ , \new_[7128]_ , \new_[7129]_ ,
    \new_[7130]_ , \new_[7131]_ , \new_[7135]_ , \new_[7136]_ ,
    \new_[7139]_ , \new_[7142]_ , \new_[7143]_ , \new_[7144]_ ,
    \new_[7147]_ , \new_[7150]_ , \new_[7151]_ , \new_[7154]_ ,
    \new_[7157]_ , \new_[7158]_ , \new_[7159]_ , \new_[7160]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7168]_ , \new_[7171]_ ,
    \new_[7172]_ , \new_[7173]_ , \new_[7176]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7183]_ , \new_[7186]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7192]_ , \new_[7193]_ , \new_[7197]_ , \new_[7198]_ ,
    \new_[7201]_ , \new_[7204]_ , \new_[7205]_ , \new_[7206]_ ,
    \new_[7209]_ , \new_[7212]_ , \new_[7213]_ , \new_[7216]_ ,
    \new_[7219]_ , \new_[7220]_ , \new_[7221]_ , \new_[7222]_ ,
    \new_[7226]_ , \new_[7227]_ , \new_[7230]_ , \new_[7233]_ ,
    \new_[7234]_ , \new_[7235]_ , \new_[7238]_ , \new_[7241]_ ,
    \new_[7242]_ , \new_[7245]_ , \new_[7248]_ , \new_[7249]_ ,
    \new_[7250]_ , \new_[7251]_ , \new_[7252]_ , \new_[7256]_ ,
    \new_[7257]_ , \new_[7260]_ , \new_[7263]_ , \new_[7264]_ ,
    \new_[7265]_ , \new_[7268]_ , \new_[7271]_ , \new_[7272]_ ,
    \new_[7275]_ , \new_[7278]_ , \new_[7279]_ , \new_[7280]_ ,
    \new_[7281]_ , \new_[7285]_ , \new_[7286]_ , \new_[7289]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7294]_ , \new_[7297]_ ,
    \new_[7300]_ , \new_[7301]_ , \new_[7304]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7312]_ , \new_[7316]_ , \new_[7317]_ , \new_[7320]_ ,
    \new_[7323]_ , \new_[7324]_ , \new_[7325]_ , \new_[7328]_ ,
    \new_[7331]_ , \new_[7332]_ , \new_[7335]_ , \new_[7338]_ ,
    \new_[7339]_ , \new_[7340]_ , \new_[7341]_ , \new_[7345]_ ,
    \new_[7346]_ , \new_[7349]_ , \new_[7352]_ , \new_[7353]_ ,
    \new_[7354]_ , \new_[7357]_ , \new_[7360]_ , \new_[7361]_ ,
    \new_[7364]_ , \new_[7367]_ , \new_[7368]_ , \new_[7369]_ ,
    \new_[7370]_ , \new_[7371]_ , \new_[7375]_ , \new_[7376]_ ,
    \new_[7379]_ , \new_[7382]_ , \new_[7383]_ , \new_[7384]_ ,
    \new_[7387]_ , \new_[7390]_ , \new_[7391]_ , \new_[7394]_ ,
    \new_[7397]_ , \new_[7398]_ , \new_[7399]_ , \new_[7400]_ ,
    \new_[7404]_ , \new_[7405]_ , \new_[7408]_ , \new_[7411]_ ,
    \new_[7412]_ , \new_[7413]_ , \new_[7416]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7423]_ , \new_[7426]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7429]_ , \new_[7430]_ , \new_[7431]_ ,
    \new_[7432]_ , \new_[7436]_ , \new_[7437]_ , \new_[7440]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7448]_ ,
    \new_[7451]_ , \new_[7452]_ , \new_[7455]_ , \new_[7458]_ ,
    \new_[7459]_ , \new_[7460]_ , \new_[7461]_ , \new_[7465]_ ,
    \new_[7466]_ , \new_[7469]_ , \new_[7472]_ , \new_[7473]_ ,
    \new_[7474]_ , \new_[7477]_ , \new_[7480]_ , \new_[7481]_ ,
    \new_[7484]_ , \new_[7487]_ , \new_[7488]_ , \new_[7489]_ ,
    \new_[7490]_ , \new_[7491]_ , \new_[7495]_ , \new_[7496]_ ,
    \new_[7499]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7507]_ , \new_[7510]_ , \new_[7511]_ , \new_[7514]_ ,
    \new_[7517]_ , \new_[7518]_ , \new_[7519]_ , \new_[7520]_ ,
    \new_[7524]_ , \new_[7525]_ , \new_[7528]_ , \new_[7531]_ ,
    \new_[7532]_ , \new_[7533]_ , \new_[7536]_ , \new_[7539]_ ,
    \new_[7540]_ , \new_[7543]_ , \new_[7546]_ , \new_[7547]_ ,
    \new_[7548]_ , \new_[7549]_ , \new_[7550]_ , \new_[7551]_ ,
    \new_[7555]_ , \new_[7556]_ , \new_[7559]_ , \new_[7562]_ ,
    \new_[7563]_ , \new_[7564]_ , \new_[7567]_ , \new_[7570]_ ,
    \new_[7571]_ , \new_[7574]_ , \new_[7577]_ , \new_[7578]_ ,
    \new_[7579]_ , \new_[7580]_ , \new_[7584]_ , \new_[7585]_ ,
    \new_[7588]_ , \new_[7591]_ , \new_[7592]_ , \new_[7593]_ ,
    \new_[7596]_ , \new_[7599]_ , \new_[7600]_ , \new_[7603]_ ,
    \new_[7606]_ , \new_[7607]_ , \new_[7608]_ , \new_[7609]_ ,
    \new_[7610]_ , \new_[7614]_ , \new_[7615]_ , \new_[7618]_ ,
    \new_[7621]_ , \new_[7622]_ , \new_[7623]_ , \new_[7626]_ ,
    \new_[7629]_ , \new_[7630]_ , \new_[7633]_ , \new_[7636]_ ,
    \new_[7637]_ , \new_[7638]_ , \new_[7639]_ , \new_[7643]_ ,
    \new_[7644]_ , \new_[7647]_ , \new_[7650]_ , \new_[7651]_ ,
    \new_[7652]_ , \new_[7655]_ , \new_[7658]_ , \new_[7659]_ ,
    \new_[7662]_ , \new_[7665]_ , \new_[7666]_ , \new_[7667]_ ,
    \new_[7668]_ , \new_[7669]_ , \new_[7670]_ , \new_[7671]_ ,
    \new_[7672]_ , \new_[7673]_ , \new_[7674]_ , \new_[7675]_ ,
    \new_[7679]_ , \new_[7680]_ , \new_[7683]_ , \new_[7686]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7692]_ , \new_[7693]_ ,
    \new_[7696]_ , \new_[7699]_ , \new_[7700]_ , \new_[7701]_ ,
    \new_[7702]_ , \new_[7706]_ , \new_[7707]_ , \new_[7710]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7715]_ , \new_[7718]_ ,
    \new_[7721]_ , \new_[7722]_ , \new_[7725]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7736]_ , \new_[7737]_ , \new_[7740]_ , \new_[7743]_ ,
    \new_[7744]_ , \new_[7745]_ , \new_[7748]_ , \new_[7751]_ ,
    \new_[7752]_ , \new_[7755]_ , \new_[7758]_ , \new_[7759]_ ,
    \new_[7760]_ , \new_[7761]_ , \new_[7765]_ , \new_[7766]_ ,
    \new_[7769]_ , \new_[7772]_ , \new_[7773]_ , \new_[7774]_ ,
    \new_[7777]_ , \new_[7780]_ , \new_[7781]_ , \new_[7784]_ ,
    \new_[7787]_ , \new_[7788]_ , \new_[7789]_ , \new_[7790]_ ,
    \new_[7791]_ , \new_[7792]_ , \new_[7796]_ , \new_[7797]_ ,
    \new_[7800]_ , \new_[7803]_ , \new_[7804]_ , \new_[7805]_ ,
    \new_[7808]_ , \new_[7811]_ , \new_[7812]_ , \new_[7815]_ ,
    \new_[7818]_ , \new_[7819]_ , \new_[7820]_ , \new_[7821]_ ,
    \new_[7825]_ , \new_[7826]_ , \new_[7829]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7834]_ , \new_[7837]_ , \new_[7840]_ ,
    \new_[7841]_ , \new_[7844]_ , \new_[7847]_ , \new_[7848]_ ,
    \new_[7849]_ , \new_[7850]_ , \new_[7851]_ , \new_[7855]_ ,
    \new_[7856]_ , \new_[7859]_ , \new_[7862]_ , \new_[7863]_ ,
    \new_[7864]_ , \new_[7867]_ , \new_[7870]_ , \new_[7871]_ ,
    \new_[7874]_ , \new_[7877]_ , \new_[7878]_ , \new_[7879]_ ,
    \new_[7880]_ , \new_[7884]_ , \new_[7885]_ , \new_[7888]_ ,
    \new_[7891]_ , \new_[7892]_ , \new_[7893]_ , \new_[7896]_ ,
    \new_[7899]_ , \new_[7900]_ , \new_[7903]_ , \new_[7906]_ ,
    \new_[7907]_ , \new_[7908]_ , \new_[7909]_ , \new_[7910]_ ,
    \new_[7911]_ , \new_[7912]_ , \new_[7916]_ , \new_[7917]_ ,
    \new_[7920]_ , \new_[7923]_ , \new_[7924]_ , \new_[7925]_ ,
    \new_[7928]_ , \new_[7931]_ , \new_[7932]_ , \new_[7935]_ ,
    \new_[7938]_ , \new_[7939]_ , \new_[7940]_ , \new_[7941]_ ,
    \new_[7945]_ , \new_[7946]_ , \new_[7949]_ , \new_[7952]_ ,
    \new_[7953]_ , \new_[7954]_ , \new_[7957]_ , \new_[7960]_ ,
    \new_[7961]_ , \new_[7964]_ , \new_[7967]_ , \new_[7968]_ ,
    \new_[7969]_ , \new_[7970]_ , \new_[7971]_ , \new_[7975]_ ,
    \new_[7976]_ , \new_[7979]_ , \new_[7982]_ , \new_[7983]_ ,
    \new_[7984]_ , \new_[7987]_ , \new_[7990]_ , \new_[7991]_ ,
    \new_[7994]_ , \new_[7997]_ , \new_[7998]_ , \new_[7999]_ ,
    \new_[8000]_ , \new_[8004]_ , \new_[8005]_ , \new_[8008]_ ,
    \new_[8011]_ , \new_[8012]_ , \new_[8013]_ , \new_[8016]_ ,
    \new_[8019]_ , \new_[8020]_ , \new_[8023]_ , \new_[8026]_ ,
    \new_[8027]_ , \new_[8028]_ , \new_[8029]_ , \new_[8030]_ ,
    \new_[8031]_ , \new_[8035]_ , \new_[8036]_ , \new_[8039]_ ,
    \new_[8042]_ , \new_[8043]_ , \new_[8044]_ , \new_[8047]_ ,
    \new_[8050]_ , \new_[8051]_ , \new_[8054]_ , \new_[8057]_ ,
    \new_[8058]_ , \new_[8059]_ , \new_[8060]_ , \new_[8064]_ ,
    \new_[8065]_ , \new_[8068]_ , \new_[8071]_ , \new_[8072]_ ,
    \new_[8073]_ , \new_[8076]_ , \new_[8079]_ , \new_[8080]_ ,
    \new_[8083]_ , \new_[8086]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8089]_ , \new_[8090]_ , \new_[8094]_ , \new_[8095]_ ,
    \new_[8098]_ , \new_[8101]_ , \new_[8102]_ , \new_[8103]_ ,
    \new_[8106]_ , \new_[8109]_ , \new_[8110]_ , \new_[8113]_ ,
    \new_[8116]_ , \new_[8117]_ , \new_[8118]_ , \new_[8119]_ ,
    \new_[8123]_ , \new_[8124]_ , \new_[8127]_ , \new_[8130]_ ,
    \new_[8131]_ , \new_[8132]_ , \new_[8135]_ , \new_[8138]_ ,
    \new_[8139]_ , \new_[8142]_ , \new_[8145]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8148]_ , \new_[8149]_ , \new_[8150]_ ,
    \new_[8151]_ , \new_[8152]_ , \new_[8156]_ , \new_[8157]_ ,
    \new_[8160]_ , \new_[8163]_ , \new_[8164]_ , \new_[8165]_ ,
    \new_[8168]_ , \new_[8171]_ , \new_[8172]_ , \new_[8175]_ ,
    \new_[8178]_ , \new_[8179]_ , \new_[8180]_ , \new_[8181]_ ,
    \new_[8185]_ , \new_[8186]_ , \new_[8189]_ , \new_[8192]_ ,
    \new_[8193]_ , \new_[8194]_ , \new_[8197]_ , \new_[8200]_ ,
    \new_[8201]_ , \new_[8204]_ , \new_[8207]_ , \new_[8208]_ ,
    \new_[8209]_ , \new_[8210]_ , \new_[8211]_ , \new_[8215]_ ,
    \new_[8216]_ , \new_[8219]_ , \new_[8222]_ , \new_[8223]_ ,
    \new_[8224]_ , \new_[8227]_ , \new_[8230]_ , \new_[8231]_ ,
    \new_[8234]_ , \new_[8237]_ , \new_[8238]_ , \new_[8239]_ ,
    \new_[8240]_ , \new_[8244]_ , \new_[8245]_ , \new_[8248]_ ,
    \new_[8251]_ , \new_[8252]_ , \new_[8253]_ , \new_[8256]_ ,
    \new_[8259]_ , \new_[8260]_ , \new_[8263]_ , \new_[8266]_ ,
    \new_[8267]_ , \new_[8268]_ , \new_[8269]_ , \new_[8270]_ ,
    \new_[8271]_ , \new_[8275]_ , \new_[8276]_ , \new_[8279]_ ,
    \new_[8282]_ , \new_[8283]_ , \new_[8284]_ , \new_[8287]_ ,
    \new_[8290]_ , \new_[8291]_ , \new_[8294]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8304]_ ,
    \new_[8305]_ , \new_[8308]_ , \new_[8311]_ , \new_[8312]_ ,
    \new_[8313]_ , \new_[8316]_ , \new_[8319]_ , \new_[8320]_ ,
    \new_[8323]_ , \new_[8326]_ , \new_[8327]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8330]_ , \new_[8334]_ , \new_[8335]_ ,
    \new_[8338]_ , \new_[8341]_ , \new_[8342]_ , \new_[8343]_ ,
    \new_[8346]_ , \new_[8349]_ , \new_[8350]_ , \new_[8353]_ ,
    \new_[8356]_ , \new_[8357]_ , \new_[8358]_ , \new_[8359]_ ,
    \new_[8363]_ , \new_[8364]_ , \new_[8367]_ , \new_[8370]_ ,
    \new_[8371]_ , \new_[8372]_ , \new_[8375]_ , \new_[8378]_ ,
    \new_[8379]_ , \new_[8382]_ , \new_[8385]_ , \new_[8386]_ ,
    \new_[8387]_ , \new_[8388]_ , \new_[8389]_ , \new_[8390]_ ,
    \new_[8391]_ , \new_[8395]_ , \new_[8396]_ , \new_[8399]_ ,
    \new_[8402]_ , \new_[8403]_ , \new_[8404]_ , \new_[8407]_ ,
    \new_[8410]_ , \new_[8411]_ , \new_[8414]_ , \new_[8417]_ ,
    \new_[8418]_ , \new_[8419]_ , \new_[8420]_ , \new_[8424]_ ,
    \new_[8425]_ , \new_[8428]_ , \new_[8431]_ , \new_[8432]_ ,
    \new_[8433]_ , \new_[8436]_ , \new_[8439]_ , \new_[8440]_ ,
    \new_[8443]_ , \new_[8446]_ , \new_[8447]_ , \new_[8448]_ ,
    \new_[8449]_ , \new_[8450]_ , \new_[8454]_ , \new_[8455]_ ,
    \new_[8458]_ , \new_[8461]_ , \new_[8462]_ , \new_[8463]_ ,
    \new_[8466]_ , \new_[8469]_ , \new_[8470]_ , \new_[8473]_ ,
    \new_[8476]_ , \new_[8477]_ , \new_[8478]_ , \new_[8479]_ ,
    \new_[8483]_ , \new_[8484]_ , \new_[8487]_ , \new_[8490]_ ,
    \new_[8491]_ , \new_[8492]_ , \new_[8495]_ , \new_[8498]_ ,
    \new_[8499]_ , \new_[8502]_ , \new_[8505]_ , \new_[8506]_ ,
    \new_[8507]_ , \new_[8508]_ , \new_[8509]_ , \new_[8510]_ ,
    \new_[8514]_ , \new_[8515]_ , \new_[8518]_ , \new_[8521]_ ,
    \new_[8522]_ , \new_[8523]_ , \new_[8526]_ , \new_[8529]_ ,
    \new_[8530]_ , \new_[8533]_ , \new_[8536]_ , \new_[8537]_ ,
    \new_[8538]_ , \new_[8539]_ , \new_[8543]_ , \new_[8544]_ ,
    \new_[8547]_ , \new_[8550]_ , \new_[8551]_ , \new_[8552]_ ,
    \new_[8555]_ , \new_[8558]_ , \new_[8559]_ , \new_[8562]_ ,
    \new_[8565]_ , \new_[8566]_ , \new_[8567]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8573]_ , \new_[8574]_ , \new_[8577]_ ,
    \new_[8580]_ , \new_[8581]_ , \new_[8582]_ , \new_[8585]_ ,
    \new_[8588]_ , \new_[8589]_ , \new_[8592]_ , \new_[8595]_ ,
    \new_[8596]_ , \new_[8597]_ , \new_[8598]_ , \new_[8602]_ ,
    \new_[8603]_ , \new_[8606]_ , \new_[8609]_ , \new_[8610]_ ,
    \new_[8611]_ , \new_[8614]_ , \new_[8617]_ , \new_[8618]_ ,
    \new_[8621]_ , \new_[8624]_ , \new_[8625]_ , \new_[8626]_ ,
    \new_[8627]_ , \new_[8628]_ , \new_[8629]_ , \new_[8630]_ ,
    \new_[8631]_ , \new_[8632]_ , \new_[8636]_ , \new_[8637]_ ,
    \new_[8640]_ , \new_[8643]_ , \new_[8644]_ , \new_[8645]_ ,
    \new_[8648]_ , \new_[8651]_ , \new_[8652]_ , \new_[8655]_ ,
    \new_[8658]_ , \new_[8659]_ , \new_[8660]_ , \new_[8661]_ ,
    \new_[8665]_ , \new_[8666]_ , \new_[8669]_ , \new_[8672]_ ,
    \new_[8673]_ , \new_[8674]_ , \new_[8677]_ , \new_[8680]_ ,
    \new_[8681]_ , \new_[8684]_ , \new_[8687]_ , \new_[8688]_ ,
    \new_[8689]_ , \new_[8690]_ , \new_[8691]_ , \new_[8695]_ ,
    \new_[8696]_ , \new_[8699]_ , \new_[8702]_ , \new_[8703]_ ,
    \new_[8704]_ , \new_[8707]_ , \new_[8710]_ , \new_[8711]_ ,
    \new_[8714]_ , \new_[8717]_ , \new_[8718]_ , \new_[8719]_ ,
    \new_[8720]_ , \new_[8724]_ , \new_[8725]_ , \new_[8728]_ ,
    \new_[8731]_ , \new_[8732]_ , \new_[8733]_ , \new_[8736]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8743]_ , \new_[8746]_ ,
    \new_[8747]_ , \new_[8748]_ , \new_[8749]_ , \new_[8750]_ ,
    \new_[8751]_ , \new_[8755]_ , \new_[8756]_ , \new_[8759]_ ,
    \new_[8762]_ , \new_[8763]_ , \new_[8764]_ , \new_[8767]_ ,
    \new_[8770]_ , \new_[8771]_ , \new_[8774]_ , \new_[8777]_ ,
    \new_[8778]_ , \new_[8779]_ , \new_[8780]_ , \new_[8784]_ ,
    \new_[8785]_ , \new_[8788]_ , \new_[8791]_ , \new_[8792]_ ,
    \new_[8793]_ , \new_[8796]_ , \new_[8799]_ , \new_[8800]_ ,
    \new_[8803]_ , \new_[8806]_ , \new_[8807]_ , \new_[8808]_ ,
    \new_[8809]_ , \new_[8810]_ , \new_[8814]_ , \new_[8815]_ ,
    \new_[8818]_ , \new_[8821]_ , \new_[8822]_ , \new_[8823]_ ,
    \new_[8826]_ , \new_[8829]_ , \new_[8830]_ , \new_[8833]_ ,
    \new_[8836]_ , \new_[8837]_ , \new_[8838]_ , \new_[8839]_ ,
    \new_[8843]_ , \new_[8844]_ , \new_[8847]_ , \new_[8850]_ ,
    \new_[8851]_ , \new_[8852]_ , \new_[8855]_ , \new_[8858]_ ,
    \new_[8859]_ , \new_[8862]_ , \new_[8865]_ , \new_[8866]_ ,
    \new_[8867]_ , \new_[8868]_ , \new_[8869]_ , \new_[8870]_ ,
    \new_[8871]_ , \new_[8875]_ , \new_[8876]_ , \new_[8879]_ ,
    \new_[8882]_ , \new_[8883]_ , \new_[8884]_ , \new_[8887]_ ,
    \new_[8890]_ , \new_[8891]_ , \new_[8894]_ , \new_[8897]_ ,
    \new_[8898]_ , \new_[8899]_ , \new_[8900]_ , \new_[8904]_ ,
    \new_[8905]_ , \new_[8908]_ , \new_[8911]_ , \new_[8912]_ ,
    \new_[8913]_ , \new_[8916]_ , \new_[8919]_ , \new_[8920]_ ,
    \new_[8923]_ , \new_[8926]_ , \new_[8927]_ , \new_[8928]_ ,
    \new_[8929]_ , \new_[8930]_ , \new_[8934]_ , \new_[8935]_ ,
    \new_[8938]_ , \new_[8941]_ , \new_[8942]_ , \new_[8943]_ ,
    \new_[8946]_ , \new_[8949]_ , \new_[8950]_ , \new_[8953]_ ,
    \new_[8956]_ , \new_[8957]_ , \new_[8958]_ , \new_[8959]_ ,
    \new_[8963]_ , \new_[8964]_ , \new_[8967]_ , \new_[8970]_ ,
    \new_[8971]_ , \new_[8972]_ , \new_[8975]_ , \new_[8978]_ ,
    \new_[8979]_ , \new_[8982]_ , \new_[8985]_ , \new_[8986]_ ,
    \new_[8987]_ , \new_[8988]_ , \new_[8989]_ , \new_[8990]_ ,
    \new_[8994]_ , \new_[8995]_ , \new_[8998]_ , \new_[9001]_ ,
    \new_[9002]_ , \new_[9003]_ , \new_[9006]_ , \new_[9009]_ ,
    \new_[9010]_ , \new_[9013]_ , \new_[9016]_ , \new_[9017]_ ,
    \new_[9018]_ , \new_[9019]_ , \new_[9023]_ , \new_[9024]_ ,
    \new_[9027]_ , \new_[9030]_ , \new_[9031]_ , \new_[9032]_ ,
    \new_[9035]_ , \new_[9038]_ , \new_[9039]_ , \new_[9042]_ ,
    \new_[9045]_ , \new_[9046]_ , \new_[9047]_ , \new_[9048]_ ,
    \new_[9049]_ , \new_[9053]_ , \new_[9054]_ , \new_[9057]_ ,
    \new_[9060]_ , \new_[9061]_ , \new_[9062]_ , \new_[9065]_ ,
    \new_[9068]_ , \new_[9069]_ , \new_[9072]_ , \new_[9075]_ ,
    \new_[9076]_ , \new_[9077]_ , \new_[9078]_ , \new_[9082]_ ,
    \new_[9083]_ , \new_[9086]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9091]_ , \new_[9094]_ , \new_[9097]_ , \new_[9098]_ ,
    \new_[9101]_ , \new_[9104]_ , \new_[9105]_ , \new_[9106]_ ,
    \new_[9107]_ , \new_[9108]_ , \new_[9109]_ , \new_[9110]_ ,
    \new_[9111]_ , \new_[9115]_ , \new_[9116]_ , \new_[9119]_ ,
    \new_[9122]_ , \new_[9123]_ , \new_[9124]_ , \new_[9127]_ ,
    \new_[9130]_ , \new_[9131]_ , \new_[9134]_ , \new_[9137]_ ,
    \new_[9138]_ , \new_[9139]_ , \new_[9140]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9148]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9156]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9163]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9174]_ , \new_[9175]_ ,
    \new_[9178]_ , \new_[9181]_ , \new_[9182]_ , \new_[9183]_ ,
    \new_[9186]_ , \new_[9189]_ , \new_[9190]_ , \new_[9193]_ ,
    \new_[9196]_ , \new_[9197]_ , \new_[9198]_ , \new_[9199]_ ,
    \new_[9203]_ , \new_[9204]_ , \new_[9207]_ , \new_[9210]_ ,
    \new_[9211]_ , \new_[9212]_ , \new_[9215]_ , \new_[9218]_ ,
    \new_[9219]_ , \new_[9222]_ , \new_[9225]_ , \new_[9226]_ ,
    \new_[9227]_ , \new_[9228]_ , \new_[9229]_ , \new_[9230]_ ,
    \new_[9234]_ , \new_[9235]_ , \new_[9238]_ , \new_[9241]_ ,
    \new_[9242]_ , \new_[9243]_ , \new_[9246]_ , \new_[9249]_ ,
    \new_[9250]_ , \new_[9253]_ , \new_[9256]_ , \new_[9257]_ ,
    \new_[9258]_ , \new_[9259]_ , \new_[9263]_ , \new_[9264]_ ,
    \new_[9267]_ , \new_[9270]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9275]_ , \new_[9278]_ , \new_[9279]_ , \new_[9282]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9293]_ , \new_[9294]_ , \new_[9297]_ ,
    \new_[9300]_ , \new_[9301]_ , \new_[9302]_ , \new_[9305]_ ,
    \new_[9308]_ , \new_[9309]_ , \new_[9312]_ , \new_[9315]_ ,
    \new_[9316]_ , \new_[9317]_ , \new_[9318]_ , \new_[9322]_ ,
    \new_[9323]_ , \new_[9326]_ , \new_[9329]_ , \new_[9330]_ ,
    \new_[9331]_ , \new_[9334]_ , \new_[9337]_ , \new_[9338]_ ,
    \new_[9341]_ , \new_[9344]_ , \new_[9345]_ , \new_[9346]_ ,
    \new_[9347]_ , \new_[9348]_ , \new_[9349]_ , \new_[9350]_ ,
    \new_[9354]_ , \new_[9355]_ , \new_[9358]_ , \new_[9361]_ ,
    \new_[9362]_ , \new_[9363]_ , \new_[9366]_ , \new_[9369]_ ,
    \new_[9370]_ , \new_[9373]_ , \new_[9376]_ , \new_[9377]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9383]_ , \new_[9384]_ ,
    \new_[9387]_ , \new_[9390]_ , \new_[9391]_ , \new_[9392]_ ,
    \new_[9395]_ , \new_[9398]_ , \new_[9399]_ , \new_[9402]_ ,
    \new_[9405]_ , \new_[9406]_ , \new_[9407]_ , \new_[9408]_ ,
    \new_[9409]_ , \new_[9413]_ , \new_[9414]_ , \new_[9417]_ ,
    \new_[9420]_ , \new_[9421]_ , \new_[9422]_ , \new_[9425]_ ,
    \new_[9428]_ , \new_[9429]_ , \new_[9432]_ , \new_[9435]_ ,
    \new_[9436]_ , \new_[9437]_ , \new_[9438]_ , \new_[9442]_ ,
    \new_[9443]_ , \new_[9446]_ , \new_[9449]_ , \new_[9450]_ ,
    \new_[9451]_ , \new_[9454]_ , \new_[9457]_ , \new_[9458]_ ,
    \new_[9461]_ , \new_[9464]_ , \new_[9465]_ , \new_[9466]_ ,
    \new_[9467]_ , \new_[9468]_ , \new_[9469]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9477]_ , \new_[9480]_ , \new_[9481]_ ,
    \new_[9482]_ , \new_[9485]_ , \new_[9488]_ , \new_[9489]_ ,
    \new_[9492]_ , \new_[9495]_ , \new_[9496]_ , \new_[9497]_ ,
    \new_[9498]_ , \new_[9502]_ , \new_[9503]_ , \new_[9506]_ ,
    \new_[9509]_ , \new_[9510]_ , \new_[9511]_ , \new_[9514]_ ,
    \new_[9517]_ , \new_[9518]_ , \new_[9521]_ , \new_[9524]_ ,
    \new_[9525]_ , \new_[9526]_ , \new_[9527]_ , \new_[9528]_ ,
    \new_[9532]_ , \new_[9533]_ , \new_[9536]_ , \new_[9539]_ ,
    \new_[9540]_ , \new_[9541]_ , \new_[9544]_ , \new_[9547]_ ,
    \new_[9548]_ , \new_[9551]_ , \new_[9554]_ , \new_[9555]_ ,
    \new_[9556]_ , \new_[9557]_ , \new_[9561]_ , \new_[9562]_ ,
    \new_[9565]_ , \new_[9568]_ , \new_[9569]_ , \new_[9570]_ ,
    \new_[9573]_ , \new_[9576]_ , \new_[9577]_ , \new_[9580]_ ,
    \new_[9583]_ , \new_[9584]_ , \new_[9585]_ , \new_[9586]_ ,
    \new_[9587]_ , \new_[9588]_ , \new_[9589]_ , \new_[9590]_ ,
    \new_[9591]_ , \new_[9592]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9600]_ , \new_[9603]_ , \new_[9604]_ , \new_[9605]_ ,
    \new_[9608]_ , \new_[9611]_ , \new_[9612]_ , \new_[9615]_ ,
    \new_[9618]_ , \new_[9619]_ , \new_[9620]_ , \new_[9621]_ ,
    \new_[9625]_ , \new_[9626]_ , \new_[9629]_ , \new_[9632]_ ,
    \new_[9633]_ , \new_[9634]_ , \new_[9637]_ , \new_[9640]_ ,
    \new_[9641]_ , \new_[9644]_ , \new_[9647]_ , \new_[9648]_ ,
    \new_[9649]_ , \new_[9650]_ , \new_[9651]_ , \new_[9655]_ ,
    \new_[9656]_ , \new_[9659]_ , \new_[9662]_ , \new_[9663]_ ,
    \new_[9664]_ , \new_[9667]_ , \new_[9670]_ , \new_[9671]_ ,
    \new_[9674]_ , \new_[9677]_ , \new_[9678]_ , \new_[9679]_ ,
    \new_[9680]_ , \new_[9684]_ , \new_[9685]_ , \new_[9688]_ ,
    \new_[9691]_ , \new_[9692]_ , \new_[9693]_ , \new_[9696]_ ,
    \new_[9699]_ , \new_[9700]_ , \new_[9703]_ , \new_[9706]_ ,
    \new_[9707]_ , \new_[9708]_ , \new_[9709]_ , \new_[9710]_ ,
    \new_[9711]_ , \new_[9715]_ , \new_[9716]_ , \new_[9719]_ ,
    \new_[9722]_ , \new_[9723]_ , \new_[9724]_ , \new_[9727]_ ,
    \new_[9730]_ , \new_[9731]_ , \new_[9734]_ , \new_[9737]_ ,
    \new_[9738]_ , \new_[9739]_ , \new_[9740]_ , \new_[9744]_ ,
    \new_[9745]_ , \new_[9748]_ , \new_[9751]_ , \new_[9752]_ ,
    \new_[9753]_ , \new_[9756]_ , \new_[9759]_ , \new_[9760]_ ,
    \new_[9763]_ , \new_[9766]_ , \new_[9767]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9770]_ , \new_[9774]_ , \new_[9775]_ ,
    \new_[9778]_ , \new_[9781]_ , \new_[9782]_ , \new_[9783]_ ,
    \new_[9786]_ , \new_[9789]_ , \new_[9790]_ , \new_[9793]_ ,
    \new_[9796]_ , \new_[9797]_ , \new_[9798]_ , \new_[9799]_ ,
    \new_[9803]_ , \new_[9804]_ , \new_[9807]_ , \new_[9810]_ ,
    \new_[9811]_ , \new_[9812]_ , \new_[9815]_ , \new_[9818]_ ,
    \new_[9819]_ , \new_[9822]_ , \new_[9825]_ , \new_[9826]_ ,
    \new_[9827]_ , \new_[9828]_ , \new_[9829]_ , \new_[9830]_ ,
    \new_[9831]_ , \new_[9835]_ , \new_[9836]_ , \new_[9839]_ ,
    \new_[9842]_ , \new_[9843]_ , \new_[9844]_ , \new_[9847]_ ,
    \new_[9850]_ , \new_[9851]_ , \new_[9854]_ , \new_[9857]_ ,
    \new_[9858]_ , \new_[9859]_ , \new_[9860]_ , \new_[9864]_ ,
    \new_[9865]_ , \new_[9868]_ , \new_[9871]_ , \new_[9872]_ ,
    \new_[9873]_ , \new_[9876]_ , \new_[9879]_ , \new_[9880]_ ,
    \new_[9883]_ , \new_[9886]_ , \new_[9887]_ , \new_[9888]_ ,
    \new_[9889]_ , \new_[9890]_ , \new_[9894]_ , \new_[9895]_ ,
    \new_[9898]_ , \new_[9901]_ , \new_[9902]_ , \new_[9903]_ ,
    \new_[9906]_ , \new_[9909]_ , \new_[9910]_ , \new_[9913]_ ,
    \new_[9916]_ , \new_[9917]_ , \new_[9918]_ , \new_[9919]_ ,
    \new_[9923]_ , \new_[9924]_ , \new_[9927]_ , \new_[9930]_ ,
    \new_[9931]_ , \new_[9932]_ , \new_[9935]_ , \new_[9938]_ ,
    \new_[9939]_ , \new_[9942]_ , \new_[9945]_ , \new_[9946]_ ,
    \new_[9947]_ , \new_[9948]_ , \new_[9949]_ , \new_[9950]_ ,
    \new_[9954]_ , \new_[9955]_ , \new_[9958]_ , \new_[9961]_ ,
    \new_[9962]_ , \new_[9963]_ , \new_[9966]_ , \new_[9969]_ ,
    \new_[9970]_ , \new_[9973]_ , \new_[9976]_ , \new_[9977]_ ,
    \new_[9978]_ , \new_[9979]_ , \new_[9983]_ , \new_[9984]_ ,
    \new_[9987]_ , \new_[9990]_ , \new_[9991]_ , \new_[9992]_ ,
    \new_[9995]_ , \new_[9998]_ , \new_[9999]_ , \new_[10002]_ ,
    \new_[10005]_ , \new_[10006]_ , \new_[10007]_ , \new_[10008]_ ,
    \new_[10009]_ , \new_[10013]_ , \new_[10014]_ , \new_[10017]_ ,
    \new_[10020]_ , \new_[10021]_ , \new_[10022]_ , \new_[10025]_ ,
    \new_[10028]_ , \new_[10029]_ , \new_[10032]_ , \new_[10035]_ ,
    \new_[10036]_ , \new_[10037]_ , \new_[10038]_ , \new_[10042]_ ,
    \new_[10043]_ , \new_[10046]_ , \new_[10049]_ , \new_[10050]_ ,
    \new_[10051]_ , \new_[10054]_ , \new_[10057]_ , \new_[10058]_ ,
    \new_[10061]_ , \new_[10064]_ , \new_[10065]_ , \new_[10066]_ ,
    \new_[10067]_ , \new_[10068]_ , \new_[10069]_ , \new_[10070]_ ,
    \new_[10071]_ , \new_[10075]_ , \new_[10076]_ , \new_[10079]_ ,
    \new_[10082]_ , \new_[10083]_ , \new_[10084]_ , \new_[10087]_ ,
    \new_[10090]_ , \new_[10091]_ , \new_[10094]_ , \new_[10097]_ ,
    \new_[10098]_ , \new_[10099]_ , \new_[10100]_ , \new_[10104]_ ,
    \new_[10105]_ , \new_[10108]_ , \new_[10111]_ , \new_[10112]_ ,
    \new_[10113]_ , \new_[10116]_ , \new_[10119]_ , \new_[10120]_ ,
    \new_[10123]_ , \new_[10126]_ , \new_[10127]_ , \new_[10128]_ ,
    \new_[10129]_ , \new_[10130]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10138]_ , \new_[10141]_ , \new_[10142]_ , \new_[10143]_ ,
    \new_[10146]_ , \new_[10149]_ , \new_[10150]_ , \new_[10153]_ ,
    \new_[10156]_ , \new_[10157]_ , \new_[10158]_ , \new_[10159]_ ,
    \new_[10163]_ , \new_[10164]_ , \new_[10167]_ , \new_[10170]_ ,
    \new_[10171]_ , \new_[10172]_ , \new_[10175]_ , \new_[10178]_ ,
    \new_[10179]_ , \new_[10182]_ , \new_[10185]_ , \new_[10186]_ ,
    \new_[10187]_ , \new_[10188]_ , \new_[10189]_ , \new_[10190]_ ,
    \new_[10194]_ , \new_[10195]_ , \new_[10198]_ , \new_[10201]_ ,
    \new_[10202]_ , \new_[10203]_ , \new_[10206]_ , \new_[10209]_ ,
    \new_[10210]_ , \new_[10213]_ , \new_[10216]_ , \new_[10217]_ ,
    \new_[10218]_ , \new_[10219]_ , \new_[10223]_ , \new_[10224]_ ,
    \new_[10227]_ , \new_[10230]_ , \new_[10231]_ , \new_[10232]_ ,
    \new_[10235]_ , \new_[10238]_ , \new_[10239]_ , \new_[10242]_ ,
    \new_[10245]_ , \new_[10246]_ , \new_[10247]_ , \new_[10248]_ ,
    \new_[10249]_ , \new_[10253]_ , \new_[10254]_ , \new_[10257]_ ,
    \new_[10260]_ , \new_[10261]_ , \new_[10262]_ , \new_[10265]_ ,
    \new_[10268]_ , \new_[10269]_ , \new_[10272]_ , \new_[10275]_ ,
    \new_[10276]_ , \new_[10277]_ , \new_[10278]_ , \new_[10282]_ ,
    \new_[10283]_ , \new_[10286]_ , \new_[10289]_ , \new_[10290]_ ,
    \new_[10291]_ , \new_[10294]_ , \new_[10297]_ , \new_[10298]_ ,
    \new_[10301]_ , \new_[10304]_ , \new_[10305]_ , \new_[10306]_ ,
    \new_[10307]_ , \new_[10308]_ , \new_[10309]_ , \new_[10310]_ ,
    \new_[10314]_ , \new_[10315]_ , \new_[10318]_ , \new_[10321]_ ,
    \new_[10322]_ , \new_[10323]_ , \new_[10326]_ , \new_[10329]_ ,
    \new_[10330]_ , \new_[10333]_ , \new_[10336]_ , \new_[10337]_ ,
    \new_[10338]_ , \new_[10339]_ , \new_[10343]_ , \new_[10344]_ ,
    \new_[10347]_ , \new_[10350]_ , \new_[10351]_ , \new_[10352]_ ,
    \new_[10355]_ , \new_[10358]_ , \new_[10359]_ , \new_[10362]_ ,
    \new_[10365]_ , \new_[10366]_ , \new_[10367]_ , \new_[10368]_ ,
    \new_[10369]_ , \new_[10373]_ , \new_[10374]_ , \new_[10377]_ ,
    \new_[10380]_ , \new_[10381]_ , \new_[10382]_ , \new_[10385]_ ,
    \new_[10388]_ , \new_[10389]_ , \new_[10392]_ , \new_[10395]_ ,
    \new_[10396]_ , \new_[10397]_ , \new_[10398]_ , \new_[10402]_ ,
    \new_[10403]_ , \new_[10406]_ , \new_[10409]_ , \new_[10410]_ ,
    \new_[10411]_ , \new_[10414]_ , \new_[10417]_ , \new_[10418]_ ,
    \new_[10421]_ , \new_[10424]_ , \new_[10425]_ , \new_[10426]_ ,
    \new_[10427]_ , \new_[10428]_ , \new_[10429]_ , \new_[10433]_ ,
    \new_[10434]_ , \new_[10437]_ , \new_[10440]_ , \new_[10441]_ ,
    \new_[10442]_ , \new_[10445]_ , \new_[10448]_ , \new_[10449]_ ,
    \new_[10452]_ , \new_[10455]_ , \new_[10456]_ , \new_[10457]_ ,
    \new_[10458]_ , \new_[10462]_ , \new_[10463]_ , \new_[10466]_ ,
    \new_[10469]_ , \new_[10470]_ , \new_[10471]_ , \new_[10474]_ ,
    \new_[10477]_ , \new_[10478]_ , \new_[10481]_ , \new_[10484]_ ,
    \new_[10485]_ , \new_[10486]_ , \new_[10487]_ , \new_[10488]_ ,
    \new_[10492]_ , \new_[10493]_ , \new_[10496]_ , \new_[10499]_ ,
    \new_[10500]_ , \new_[10501]_ , \new_[10504]_ , \new_[10507]_ ,
    \new_[10508]_ , \new_[10511]_ , \new_[10514]_ , \new_[10515]_ ,
    \new_[10516]_ , \new_[10517]_ , \new_[10521]_ , \new_[10522]_ ,
    \new_[10525]_ , \new_[10528]_ , \new_[10529]_ , \new_[10530]_ ,
    \new_[10533]_ , \new_[10536]_ , \new_[10537]_ , \new_[10540]_ ,
    \new_[10543]_ , \new_[10544]_ , \new_[10545]_ , \new_[10546]_ ,
    \new_[10547]_ , \new_[10548]_ , \new_[10549]_ , \new_[10550]_ ,
    \new_[10551]_ , \new_[10555]_ , \new_[10556]_ , \new_[10559]_ ,
    \new_[10562]_ , \new_[10563]_ , \new_[10564]_ , \new_[10567]_ ,
    \new_[10570]_ , \new_[10571]_ , \new_[10574]_ , \new_[10577]_ ,
    \new_[10578]_ , \new_[10579]_ , \new_[10580]_ , \new_[10584]_ ,
    \new_[10585]_ , \new_[10588]_ , \new_[10591]_ , \new_[10592]_ ,
    \new_[10593]_ , \new_[10596]_ , \new_[10599]_ , \new_[10600]_ ,
    \new_[10603]_ , \new_[10606]_ , \new_[10607]_ , \new_[10608]_ ,
    \new_[10609]_ , \new_[10610]_ , \new_[10614]_ , \new_[10615]_ ,
    \new_[10618]_ , \new_[10621]_ , \new_[10622]_ , \new_[10623]_ ,
    \new_[10626]_ , \new_[10629]_ , \new_[10630]_ , \new_[10633]_ ,
    \new_[10636]_ , \new_[10637]_ , \new_[10638]_ , \new_[10639]_ ,
    \new_[10643]_ , \new_[10644]_ , \new_[10647]_ , \new_[10650]_ ,
    \new_[10651]_ , \new_[10652]_ , \new_[10655]_ , \new_[10658]_ ,
    \new_[10659]_ , \new_[10662]_ , \new_[10665]_ , \new_[10666]_ ,
    \new_[10667]_ , \new_[10668]_ , \new_[10669]_ , \new_[10670]_ ,
    \new_[10674]_ , \new_[10675]_ , \new_[10678]_ , \new_[10681]_ ,
    \new_[10682]_ , \new_[10683]_ , \new_[10686]_ , \new_[10689]_ ,
    \new_[10690]_ , \new_[10693]_ , \new_[10696]_ , \new_[10697]_ ,
    \new_[10698]_ , \new_[10699]_ , \new_[10703]_ , \new_[10704]_ ,
    \new_[10707]_ , \new_[10710]_ , \new_[10711]_ , \new_[10712]_ ,
    \new_[10715]_ , \new_[10718]_ , \new_[10719]_ , \new_[10722]_ ,
    \new_[10725]_ , \new_[10726]_ , \new_[10727]_ , \new_[10728]_ ,
    \new_[10729]_ , \new_[10733]_ , \new_[10734]_ , \new_[10737]_ ,
    \new_[10740]_ , \new_[10741]_ , \new_[10742]_ , \new_[10745]_ ,
    \new_[10748]_ , \new_[10749]_ , \new_[10752]_ , \new_[10755]_ ,
    \new_[10756]_ , \new_[10757]_ , \new_[10758]_ , \new_[10762]_ ,
    \new_[10763]_ , \new_[10766]_ , \new_[10769]_ , \new_[10770]_ ,
    \new_[10771]_ , \new_[10774]_ , \new_[10777]_ , \new_[10778]_ ,
    \new_[10781]_ , \new_[10784]_ , \new_[10785]_ , \new_[10786]_ ,
    \new_[10787]_ , \new_[10788]_ , \new_[10789]_ , \new_[10790]_ ,
    \new_[10794]_ , \new_[10795]_ , \new_[10798]_ , \new_[10801]_ ,
    \new_[10802]_ , \new_[10803]_ , \new_[10806]_ , \new_[10809]_ ,
    \new_[10810]_ , \new_[10813]_ , \new_[10816]_ , \new_[10817]_ ,
    \new_[10818]_ , \new_[10819]_ , \new_[10823]_ , \new_[10824]_ ,
    \new_[10827]_ , \new_[10830]_ , \new_[10831]_ , \new_[10832]_ ,
    \new_[10835]_ , \new_[10838]_ , \new_[10839]_ , \new_[10842]_ ,
    \new_[10845]_ , \new_[10846]_ , \new_[10847]_ , \new_[10848]_ ,
    \new_[10849]_ , \new_[10853]_ , \new_[10854]_ , \new_[10857]_ ,
    \new_[10860]_ , \new_[10861]_ , \new_[10862]_ , \new_[10865]_ ,
    \new_[10868]_ , \new_[10869]_ , \new_[10872]_ , \new_[10875]_ ,
    \new_[10876]_ , \new_[10877]_ , \new_[10878]_ , \new_[10882]_ ,
    \new_[10883]_ , \new_[10886]_ , \new_[10889]_ , \new_[10890]_ ,
    \new_[10891]_ , \new_[10894]_ , \new_[10897]_ , \new_[10898]_ ,
    \new_[10901]_ , \new_[10904]_ , \new_[10905]_ , \new_[10906]_ ,
    \new_[10907]_ , \new_[10908]_ , \new_[10909]_ , \new_[10913]_ ,
    \new_[10914]_ , \new_[10917]_ , \new_[10920]_ , \new_[10921]_ ,
    \new_[10922]_ , \new_[10925]_ , \new_[10928]_ , \new_[10929]_ ,
    \new_[10932]_ , \new_[10935]_ , \new_[10936]_ , \new_[10937]_ ,
    \new_[10938]_ , \new_[10942]_ , \new_[10943]_ , \new_[10946]_ ,
    \new_[10949]_ , \new_[10950]_ , \new_[10951]_ , \new_[10954]_ ,
    \new_[10957]_ , \new_[10958]_ , \new_[10961]_ , \new_[10964]_ ,
    \new_[10965]_ , \new_[10966]_ , \new_[10967]_ , \new_[10968]_ ,
    \new_[10972]_ , \new_[10973]_ , \new_[10976]_ , \new_[10979]_ ,
    \new_[10980]_ , \new_[10981]_ , \new_[10984]_ , \new_[10987]_ ,
    \new_[10988]_ , \new_[10991]_ , \new_[10994]_ , \new_[10995]_ ,
    \new_[10996]_ , \new_[10997]_ , \new_[11001]_ , \new_[11002]_ ,
    \new_[11005]_ , \new_[11008]_ , \new_[11009]_ , \new_[11010]_ ,
    \new_[11013]_ , \new_[11016]_ , \new_[11017]_ , \new_[11020]_ ,
    \new_[11023]_ , \new_[11024]_ , \new_[11025]_ , \new_[11026]_ ,
    \new_[11027]_ , \new_[11028]_ , \new_[11029]_ , \new_[11030]_ ,
    \new_[11034]_ , \new_[11035]_ , \new_[11038]_ , \new_[11041]_ ,
    \new_[11042]_ , \new_[11043]_ , \new_[11046]_ , \new_[11049]_ ,
    \new_[11050]_ , \new_[11053]_ , \new_[11056]_ , \new_[11057]_ ,
    \new_[11058]_ , \new_[11059]_ , \new_[11063]_ , \new_[11064]_ ,
    \new_[11067]_ , \new_[11070]_ , \new_[11071]_ , \new_[11072]_ ,
    \new_[11075]_ , \new_[11078]_ , \new_[11079]_ , \new_[11082]_ ,
    \new_[11085]_ , \new_[11086]_ , \new_[11087]_ , \new_[11088]_ ,
    \new_[11089]_ , \new_[11093]_ , \new_[11094]_ , \new_[11097]_ ,
    \new_[11100]_ , \new_[11101]_ , \new_[11102]_ , \new_[11105]_ ,
    \new_[11108]_ , \new_[11109]_ , \new_[11112]_ , \new_[11115]_ ,
    \new_[11116]_ , \new_[11117]_ , \new_[11118]_ , \new_[11122]_ ,
    \new_[11123]_ , \new_[11126]_ , \new_[11129]_ , \new_[11130]_ ,
    \new_[11131]_ , \new_[11134]_ , \new_[11137]_ , \new_[11138]_ ,
    \new_[11141]_ , \new_[11144]_ , \new_[11145]_ , \new_[11146]_ ,
    \new_[11147]_ , \new_[11148]_ , \new_[11149]_ , \new_[11153]_ ,
    \new_[11154]_ , \new_[11157]_ , \new_[11160]_ , \new_[11161]_ ,
    \new_[11162]_ , \new_[11165]_ , \new_[11168]_ , \new_[11169]_ ,
    \new_[11172]_ , \new_[11175]_ , \new_[11176]_ , \new_[11177]_ ,
    \new_[11178]_ , \new_[11182]_ , \new_[11183]_ , \new_[11186]_ ,
    \new_[11189]_ , \new_[11190]_ , \new_[11191]_ , \new_[11194]_ ,
    \new_[11197]_ , \new_[11198]_ , \new_[11201]_ , \new_[11204]_ ,
    \new_[11205]_ , \new_[11206]_ , \new_[11207]_ , \new_[11208]_ ,
    \new_[11212]_ , \new_[11213]_ , \new_[11216]_ , \new_[11219]_ ,
    \new_[11220]_ , \new_[11221]_ , \new_[11224]_ , \new_[11227]_ ,
    \new_[11228]_ , \new_[11231]_ , \new_[11234]_ , \new_[11235]_ ,
    \new_[11236]_ , \new_[11237]_ , \new_[11241]_ , \new_[11242]_ ,
    \new_[11245]_ , \new_[11248]_ , \new_[11249]_ , \new_[11250]_ ,
    \new_[11253]_ , \new_[11256]_ , \new_[11257]_ , \new_[11260]_ ,
    \new_[11263]_ , \new_[11264]_ , \new_[11265]_ , \new_[11266]_ ,
    \new_[11267]_ , \new_[11268]_ , \new_[11269]_ , \new_[11273]_ ,
    \new_[11274]_ , \new_[11277]_ , \new_[11280]_ , \new_[11281]_ ,
    \new_[11282]_ , \new_[11285]_ , \new_[11288]_ , \new_[11289]_ ,
    \new_[11292]_ , \new_[11295]_ , \new_[11296]_ , \new_[11297]_ ,
    \new_[11298]_ , \new_[11302]_ , \new_[11303]_ , \new_[11306]_ ,
    \new_[11309]_ , \new_[11310]_ , \new_[11311]_ , \new_[11314]_ ,
    \new_[11317]_ , \new_[11318]_ , \new_[11321]_ , \new_[11324]_ ,
    \new_[11325]_ , \new_[11326]_ , \new_[11327]_ , \new_[11328]_ ,
    \new_[11332]_ , \new_[11333]_ , \new_[11336]_ , \new_[11339]_ ,
    \new_[11340]_ , \new_[11341]_ , \new_[11344]_ , \new_[11347]_ ,
    \new_[11348]_ , \new_[11351]_ , \new_[11354]_ , \new_[11355]_ ,
    \new_[11356]_ , \new_[11357]_ , \new_[11361]_ , \new_[11362]_ ,
    \new_[11365]_ , \new_[11368]_ , \new_[11369]_ , \new_[11370]_ ,
    \new_[11373]_ , \new_[11376]_ , \new_[11377]_ , \new_[11380]_ ,
    \new_[11383]_ , \new_[11384]_ , \new_[11385]_ , \new_[11386]_ ,
    \new_[11387]_ , \new_[11388]_ , \new_[11392]_ , \new_[11393]_ ,
    \new_[11396]_ , \new_[11399]_ , \new_[11400]_ , \new_[11401]_ ,
    \new_[11404]_ , \new_[11407]_ , \new_[11408]_ , \new_[11411]_ ,
    \new_[11414]_ , \new_[11415]_ , \new_[11416]_ , \new_[11417]_ ,
    \new_[11421]_ , \new_[11422]_ , \new_[11425]_ , \new_[11428]_ ,
    \new_[11429]_ , \new_[11430]_ , \new_[11433]_ , \new_[11436]_ ,
    \new_[11437]_ , \new_[11440]_ , \new_[11443]_ , \new_[11444]_ ,
    \new_[11445]_ , \new_[11446]_ , \new_[11447]_ , \new_[11451]_ ,
    \new_[11452]_ , \new_[11455]_ , \new_[11458]_ , \new_[11459]_ ,
    \new_[11460]_ , \new_[11463]_ , \new_[11466]_ , \new_[11467]_ ,
    \new_[11470]_ , \new_[11473]_ , \new_[11474]_ , \new_[11475]_ ,
    \new_[11476]_ , \new_[11480]_ , \new_[11481]_ , \new_[11484]_ ,
    \new_[11487]_ , \new_[11488]_ , \new_[11489]_ , \new_[11492]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11499]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11507]_ , \new_[11508]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11511]_ , \new_[11512]_ , \new_[11515]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11522]_ , \new_[11525]_ , \new_[11526]_ ,
    \new_[11529]_ , \new_[11532]_ , \new_[11533]_ , \new_[11536]_ ,
    \new_[11539]_ , \new_[11540]_ , \new_[11543]_ , \new_[11546]_ ,
    \new_[11547]_ , \new_[11550]_ , \new_[11553]_ , \new_[11554]_ ,
    \new_[11557]_ , \new_[11560]_ , \new_[11561]_ , \new_[11564]_ ,
    \new_[11567]_ , \new_[11568]_ , \new_[11571]_ , \new_[11574]_ ,
    \new_[11575]_ , \new_[11578]_ , \new_[11581]_ , \new_[11582]_ ,
    \new_[11585]_ , \new_[11588]_ , \new_[11589]_ , \new_[11592]_ ,
    \new_[11595]_ , \new_[11596]_ , \new_[11599]_ , \new_[11602]_ ,
    \new_[11603]_ , \new_[11606]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11613]_ , \new_[11616]_ , \new_[11617]_ , \new_[11620]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11627]_ , \new_[11630]_ ,
    \new_[11631]_ , \new_[11634]_ , \new_[11637]_ , \new_[11638]_ ,
    \new_[11641]_ , \new_[11644]_ , \new_[11645]_ , \new_[11648]_ ,
    \new_[11651]_ , \new_[11652]_ , \new_[11655]_ , \new_[11658]_ ,
    \new_[11659]_ , \new_[11662]_ , \new_[11665]_ , \new_[11666]_ ,
    \new_[11669]_ , \new_[11672]_ , \new_[11673]_ , \new_[11676]_ ,
    \new_[11679]_ , \new_[11680]_ , \new_[11683]_ , \new_[11686]_ ,
    \new_[11687]_ , \new_[11690]_ , \new_[11693]_ , \new_[11694]_ ,
    \new_[11697]_ , \new_[11700]_ , \new_[11701]_ , \new_[11704]_ ,
    \new_[11707]_ , \new_[11708]_ , \new_[11711]_ , \new_[11714]_ ,
    \new_[11715]_ , \new_[11718]_ , \new_[11721]_ , \new_[11722]_ ,
    \new_[11725]_ , \new_[11728]_ , \new_[11729]_ , \new_[11732]_ ,
    \new_[11735]_ , \new_[11736]_ , \new_[11739]_ , \new_[11742]_ ,
    \new_[11743]_ , \new_[11746]_ , \new_[11749]_ , \new_[11750]_ ,
    \new_[11753]_ , \new_[11756]_ , \new_[11757]_ , \new_[11760]_ ,
    \new_[11763]_ , \new_[11764]_ , \new_[11767]_ , \new_[11770]_ ,
    \new_[11771]_ , \new_[11774]_ , \new_[11777]_ , \new_[11778]_ ,
    \new_[11781]_ , \new_[11784]_ , \new_[11785]_ , \new_[11788]_ ,
    \new_[11791]_ , \new_[11792]_ , \new_[11795]_ , \new_[11798]_ ,
    \new_[11799]_ , \new_[11802]_ , \new_[11805]_ , \new_[11806]_ ,
    \new_[11809]_ , \new_[11812]_ , \new_[11813]_ , \new_[11816]_ ,
    \new_[11819]_ , \new_[11820]_ , \new_[11823]_ , \new_[11826]_ ,
    \new_[11827]_ , \new_[11830]_ , \new_[11833]_ , \new_[11834]_ ,
    \new_[11837]_ , \new_[11840]_ , \new_[11841]_ , \new_[11844]_ ,
    \new_[11847]_ , \new_[11848]_ , \new_[11851]_ , \new_[11854]_ ,
    \new_[11855]_ , \new_[11858]_ , \new_[11861]_ , \new_[11862]_ ,
    \new_[11865]_ , \new_[11868]_ , \new_[11869]_ , \new_[11872]_ ,
    \new_[11875]_ , \new_[11876]_ , \new_[11879]_ , \new_[11882]_ ,
    \new_[11883]_ , \new_[11886]_ , \new_[11889]_ , \new_[11890]_ ,
    \new_[11893]_ , \new_[11896]_ , \new_[11897]_ , \new_[11900]_ ,
    \new_[11903]_ , \new_[11904]_ , \new_[11907]_ , \new_[11910]_ ,
    \new_[11911]_ , \new_[11914]_ , \new_[11917]_ , \new_[11918]_ ,
    \new_[11921]_ , \new_[11924]_ , \new_[11925]_ , \new_[11928]_ ,
    \new_[11931]_ , \new_[11932]_ , \new_[11935]_ , \new_[11938]_ ,
    \new_[11939]_ , \new_[11942]_ , \new_[11945]_ , \new_[11946]_ ,
    \new_[11949]_ , \new_[11952]_ , \new_[11953]_ , \new_[11956]_ ,
    \new_[11959]_ , \new_[11960]_ , \new_[11963]_ , \new_[11966]_ ,
    \new_[11967]_ , \new_[11970]_ , \new_[11974]_ , \new_[11975]_ ,
    \new_[11976]_ , \new_[11979]_ , \new_[11982]_ , \new_[11983]_ ,
    \new_[11986]_ , \new_[11990]_ , \new_[11991]_ , \new_[11992]_ ,
    \new_[11995]_ , \new_[11998]_ , \new_[11999]_ , \new_[12002]_ ,
    \new_[12006]_ , \new_[12007]_ , \new_[12008]_ , \new_[12011]_ ,
    \new_[12014]_ , \new_[12015]_ , \new_[12018]_ , \new_[12022]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12027]_ , \new_[12030]_ ,
    \new_[12031]_ , \new_[12034]_ , \new_[12038]_ , \new_[12039]_ ,
    \new_[12040]_ , \new_[12043]_ , \new_[12046]_ , \new_[12047]_ ,
    \new_[12050]_ , \new_[12054]_ , \new_[12055]_ , \new_[12056]_ ,
    \new_[12059]_ , \new_[12062]_ , \new_[12063]_ , \new_[12066]_ ,
    \new_[12070]_ , \new_[12071]_ , \new_[12072]_ , \new_[12075]_ ,
    \new_[12078]_ , \new_[12079]_ , \new_[12082]_ , \new_[12086]_ ,
    \new_[12087]_ , \new_[12088]_ , \new_[12091]_ , \new_[12094]_ ,
    \new_[12095]_ , \new_[12098]_ , \new_[12102]_ , \new_[12103]_ ,
    \new_[12104]_ , \new_[12107]_ , \new_[12110]_ , \new_[12111]_ ,
    \new_[12114]_ , \new_[12118]_ , \new_[12119]_ , \new_[12120]_ ,
    \new_[12123]_ , \new_[12126]_ , \new_[12127]_ , \new_[12130]_ ,
    \new_[12134]_ , \new_[12135]_ , \new_[12136]_ , \new_[12139]_ ,
    \new_[12142]_ , \new_[12143]_ , \new_[12146]_ , \new_[12150]_ ,
    \new_[12151]_ , \new_[12152]_ , \new_[12155]_ , \new_[12158]_ ,
    \new_[12159]_ , \new_[12162]_ , \new_[12166]_ , \new_[12167]_ ,
    \new_[12168]_ , \new_[12171]_ , \new_[12174]_ , \new_[12175]_ ,
    \new_[12178]_ , \new_[12182]_ , \new_[12183]_ , \new_[12184]_ ,
    \new_[12187]_ , \new_[12190]_ , \new_[12191]_ , \new_[12194]_ ,
    \new_[12198]_ , \new_[12199]_ , \new_[12200]_ , \new_[12203]_ ,
    \new_[12206]_ , \new_[12207]_ , \new_[12210]_ , \new_[12214]_ ,
    \new_[12215]_ , \new_[12216]_ , \new_[12219]_ , \new_[12222]_ ,
    \new_[12223]_ , \new_[12226]_ , \new_[12230]_ , \new_[12231]_ ,
    \new_[12232]_ , \new_[12235]_ , \new_[12238]_ , \new_[12239]_ ,
    \new_[12242]_ , \new_[12246]_ , \new_[12247]_ , \new_[12248]_ ,
    \new_[12251]_ , \new_[12254]_ , \new_[12255]_ , \new_[12258]_ ,
    \new_[12262]_ , \new_[12263]_ , \new_[12264]_ , \new_[12267]_ ,
    \new_[12270]_ , \new_[12271]_ , \new_[12274]_ , \new_[12278]_ ,
    \new_[12279]_ , \new_[12280]_ , \new_[12283]_ , \new_[12286]_ ,
    \new_[12287]_ , \new_[12290]_ , \new_[12294]_ , \new_[12295]_ ,
    \new_[12296]_ , \new_[12299]_ , \new_[12302]_ , \new_[12303]_ ,
    \new_[12306]_ , \new_[12310]_ , \new_[12311]_ , \new_[12312]_ ,
    \new_[12315]_ , \new_[12318]_ , \new_[12319]_ , \new_[12322]_ ,
    \new_[12326]_ , \new_[12327]_ , \new_[12328]_ , \new_[12331]_ ,
    \new_[12334]_ , \new_[12335]_ , \new_[12338]_ , \new_[12342]_ ,
    \new_[12343]_ , \new_[12344]_ , \new_[12347]_ , \new_[12351]_ ,
    \new_[12352]_ , \new_[12353]_ , \new_[12356]_ , \new_[12360]_ ,
    \new_[12361]_ , \new_[12362]_ , \new_[12365]_ , \new_[12369]_ ,
    \new_[12370]_ , \new_[12371]_ , \new_[12374]_ , \new_[12378]_ ,
    \new_[12379]_ , \new_[12380]_ , \new_[12383]_ , \new_[12387]_ ,
    \new_[12388]_ , \new_[12389]_ , \new_[12392]_ , \new_[12396]_ ,
    \new_[12397]_ , \new_[12398]_ , \new_[12401]_ , \new_[12405]_ ,
    \new_[12406]_ , \new_[12407]_ , \new_[12410]_ , \new_[12414]_ ,
    \new_[12415]_ , \new_[12416]_ , \new_[12419]_ , \new_[12423]_ ,
    \new_[12424]_ , \new_[12425]_ , \new_[12428]_ , \new_[12432]_ ,
    \new_[12433]_ , \new_[12434]_ , \new_[12437]_ , \new_[12441]_ ,
    \new_[12442]_ , \new_[12443]_ , \new_[12446]_ , \new_[12450]_ ,
    \new_[12451]_ , \new_[12452]_ , \new_[12455]_ , \new_[12459]_ ,
    \new_[12460]_ , \new_[12461]_ , \new_[12464]_ , \new_[12468]_ ,
    \new_[12469]_ , \new_[12470]_ , \new_[12473]_ , \new_[12477]_ ,
    \new_[12478]_ , \new_[12479]_ , \new_[12482]_ , \new_[12486]_ ,
    \new_[12487]_ , \new_[12488]_ , \new_[12491]_ , \new_[12495]_ ,
    \new_[12496]_ , \new_[12497]_ , \new_[12500]_ , \new_[12504]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12509]_ , \new_[12513]_ ,
    \new_[12514]_ , \new_[12515]_ , \new_[12518]_ , \new_[12522]_ ,
    \new_[12523]_ , \new_[12524]_ , \new_[12527]_ , \new_[12531]_ ,
    \new_[12532]_ , \new_[12533]_ , \new_[12536]_ , \new_[12540]_ ,
    \new_[12541]_ , \new_[12542]_ , \new_[12545]_ , \new_[12549]_ ,
    \new_[12550]_ , \new_[12551]_ , \new_[12554]_ , \new_[12558]_ ,
    \new_[12559]_ , \new_[12560]_ , \new_[12563]_ , \new_[12567]_ ,
    \new_[12568]_ , \new_[12569]_ , \new_[12572]_ , \new_[12576]_ ,
    \new_[12577]_ , \new_[12578]_ , \new_[12581]_ , \new_[12585]_ ,
    \new_[12586]_ , \new_[12587]_ , \new_[12590]_ , \new_[12594]_ ,
    \new_[12595]_ , \new_[12596]_ , \new_[12599]_ , \new_[12603]_ ,
    \new_[12604]_ , \new_[12605]_ , \new_[12608]_ , \new_[12612]_ ,
    \new_[12613]_ , \new_[12614]_ , \new_[12617]_ , \new_[12621]_ ,
    \new_[12622]_ , \new_[12623]_ , \new_[12626]_ , \new_[12630]_ ,
    \new_[12631]_ , \new_[12632]_ , \new_[12635]_ , \new_[12639]_ ,
    \new_[12640]_ , \new_[12641]_ , \new_[12644]_ , \new_[12648]_ ,
    \new_[12649]_ , \new_[12650]_ , \new_[12653]_ , \new_[12657]_ ,
    \new_[12658]_ , \new_[12659]_ , \new_[12662]_ , \new_[12666]_ ,
    \new_[12667]_ , \new_[12668]_ , \new_[12671]_ , \new_[12675]_ ,
    \new_[12676]_ , \new_[12677]_ , \new_[12680]_ , \new_[12684]_ ,
    \new_[12685]_ , \new_[12686]_ , \new_[12689]_ , \new_[12693]_ ,
    \new_[12694]_ , \new_[12695]_ , \new_[12698]_ , \new_[12702]_ ,
    \new_[12703]_ , \new_[12704]_ , \new_[12707]_ , \new_[12711]_ ,
    \new_[12712]_ , \new_[12713]_ , \new_[12716]_ , \new_[12720]_ ,
    \new_[12721]_ , \new_[12722]_ , \new_[12725]_ , \new_[12729]_ ,
    \new_[12730]_ , \new_[12731]_ , \new_[12734]_ , \new_[12738]_ ,
    \new_[12739]_ , \new_[12740]_ , \new_[12743]_ , \new_[12747]_ ,
    \new_[12748]_ , \new_[12749]_ , \new_[12752]_ , \new_[12756]_ ,
    \new_[12757]_ , \new_[12758]_ , \new_[12761]_ , \new_[12765]_ ,
    \new_[12766]_ , \new_[12767]_ , \new_[12770]_ , \new_[12774]_ ,
    \new_[12775]_ , \new_[12776]_ , \new_[12779]_ , \new_[12783]_ ,
    \new_[12784]_ , \new_[12785]_ , \new_[12788]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12794]_ , \new_[12797]_ , \new_[12801]_ ,
    \new_[12802]_ , \new_[12803]_ , \new_[12806]_ , \new_[12810]_ ,
    \new_[12811]_ , \new_[12812]_ , \new_[12815]_ , \new_[12819]_ ,
    \new_[12820]_ , \new_[12821]_ , \new_[12824]_ , \new_[12828]_ ,
    \new_[12829]_ , \new_[12830]_ , \new_[12833]_ , \new_[12837]_ ,
    \new_[12838]_ , \new_[12839]_ , \new_[12842]_ , \new_[12846]_ ,
    \new_[12847]_ , \new_[12848]_ , \new_[12851]_ , \new_[12855]_ ,
    \new_[12856]_ , \new_[12857]_ , \new_[12860]_ , \new_[12864]_ ,
    \new_[12865]_ , \new_[12866]_ , \new_[12869]_ , \new_[12873]_ ,
    \new_[12874]_ , \new_[12875]_ , \new_[12878]_ , \new_[12882]_ ,
    \new_[12883]_ , \new_[12884]_ , \new_[12887]_ , \new_[12891]_ ,
    \new_[12892]_ , \new_[12893]_ , \new_[12896]_ , \new_[12900]_ ,
    \new_[12901]_ , \new_[12902]_ , \new_[12905]_ , \new_[12909]_ ,
    \new_[12910]_ , \new_[12911]_ , \new_[12914]_ , \new_[12918]_ ,
    \new_[12919]_ , \new_[12920]_ , \new_[12923]_ , \new_[12927]_ ,
    \new_[12928]_ , \new_[12929]_ , \new_[12932]_ , \new_[12936]_ ,
    \new_[12937]_ , \new_[12938]_ , \new_[12941]_ , \new_[12945]_ ,
    \new_[12946]_ , \new_[12947]_ , \new_[12950]_ , \new_[12954]_ ,
    \new_[12955]_ , \new_[12956]_ , \new_[12959]_ , \new_[12963]_ ,
    \new_[12964]_ , \new_[12965]_ , \new_[12968]_ , \new_[12972]_ ,
    \new_[12973]_ , \new_[12974]_ , \new_[12977]_ , \new_[12981]_ ,
    \new_[12982]_ , \new_[12983]_ , \new_[12986]_ , \new_[12990]_ ,
    \new_[12991]_ , \new_[12992]_ , \new_[12995]_ , \new_[12999]_ ,
    \new_[13000]_ , \new_[13001]_ , \new_[13004]_ , \new_[13008]_ ,
    \new_[13009]_ , \new_[13010]_ , \new_[13013]_ , \new_[13017]_ ,
    \new_[13018]_ , \new_[13019]_ , \new_[13022]_ , \new_[13026]_ ,
    \new_[13027]_ , \new_[13028]_ , \new_[13031]_ , \new_[13035]_ ,
    \new_[13036]_ , \new_[13037]_ , \new_[13040]_ , \new_[13044]_ ,
    \new_[13045]_ , \new_[13046]_ , \new_[13049]_ , \new_[13053]_ ,
    \new_[13054]_ , \new_[13055]_ , \new_[13058]_ , \new_[13062]_ ,
    \new_[13063]_ , \new_[13064]_ , \new_[13067]_ , \new_[13071]_ ,
    \new_[13072]_ , \new_[13073]_ , \new_[13076]_ , \new_[13080]_ ,
    \new_[13081]_ , \new_[13082]_ , \new_[13085]_ , \new_[13089]_ ,
    \new_[13090]_ , \new_[13091]_ , \new_[13094]_ , \new_[13098]_ ,
    \new_[13099]_ , \new_[13100]_ , \new_[13103]_ , \new_[13107]_ ,
    \new_[13108]_ , \new_[13109]_ , \new_[13112]_ , \new_[13116]_ ,
    \new_[13117]_ , \new_[13118]_ , \new_[13121]_ , \new_[13125]_ ,
    \new_[13126]_ , \new_[13127]_ , \new_[13130]_ , \new_[13134]_ ,
    \new_[13135]_ , \new_[13136]_ , \new_[13139]_ , \new_[13143]_ ,
    \new_[13144]_ , \new_[13145]_ , \new_[13148]_ , \new_[13152]_ ,
    \new_[13153]_ , \new_[13154]_ , \new_[13157]_ , \new_[13161]_ ,
    \new_[13162]_ , \new_[13163]_ , \new_[13166]_ , \new_[13170]_ ,
    \new_[13171]_ , \new_[13172]_ , \new_[13175]_ , \new_[13179]_ ,
    \new_[13180]_ , \new_[13181]_ , \new_[13184]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13190]_ , \new_[13193]_ , \new_[13197]_ ,
    \new_[13198]_ , \new_[13199]_ , \new_[13202]_ , \new_[13206]_ ,
    \new_[13207]_ , \new_[13208]_ , \new_[13211]_ , \new_[13215]_ ,
    \new_[13216]_ , \new_[13217]_ , \new_[13220]_ , \new_[13224]_ ,
    \new_[13225]_ , \new_[13226]_ , \new_[13229]_ , \new_[13233]_ ,
    \new_[13234]_ , \new_[13235]_ , \new_[13238]_ , \new_[13242]_ ,
    \new_[13243]_ , \new_[13244]_ , \new_[13247]_ , \new_[13251]_ ,
    \new_[13252]_ , \new_[13253]_ , \new_[13256]_ , \new_[13260]_ ,
    \new_[13261]_ , \new_[13262]_ , \new_[13265]_ , \new_[13269]_ ,
    \new_[13270]_ , \new_[13271]_ , \new_[13274]_ , \new_[13278]_ ,
    \new_[13279]_ , \new_[13280]_ , \new_[13283]_ , \new_[13287]_ ,
    \new_[13288]_ , \new_[13289]_ , \new_[13292]_ , \new_[13296]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13301]_ , \new_[13305]_ ,
    \new_[13306]_ , \new_[13307]_ , \new_[13310]_ , \new_[13314]_ ,
    \new_[13315]_ , \new_[13316]_ , \new_[13319]_ , \new_[13323]_ ,
    \new_[13324]_ , \new_[13325]_ , \new_[13328]_ , \new_[13332]_ ,
    \new_[13333]_ , \new_[13334]_ , \new_[13337]_ , \new_[13341]_ ,
    \new_[13342]_ , \new_[13343]_ , \new_[13346]_ , \new_[13350]_ ,
    \new_[13351]_ , \new_[13352]_ , \new_[13355]_ , \new_[13359]_ ,
    \new_[13360]_ , \new_[13361]_ , \new_[13364]_ , \new_[13368]_ ,
    \new_[13369]_ , \new_[13370]_ , \new_[13373]_ , \new_[13377]_ ,
    \new_[13378]_ , \new_[13379]_ , \new_[13382]_ , \new_[13386]_ ,
    \new_[13387]_ , \new_[13388]_ , \new_[13391]_ , \new_[13395]_ ,
    \new_[13396]_ , \new_[13397]_ , \new_[13400]_ , \new_[13404]_ ,
    \new_[13405]_ , \new_[13406]_ , \new_[13409]_ , \new_[13413]_ ,
    \new_[13414]_ , \new_[13415]_ , \new_[13418]_ , \new_[13422]_ ,
    \new_[13423]_ , \new_[13424]_ , \new_[13427]_ , \new_[13431]_ ,
    \new_[13432]_ , \new_[13433]_ , \new_[13436]_ , \new_[13440]_ ,
    \new_[13441]_ , \new_[13442]_ , \new_[13445]_ , \new_[13449]_ ,
    \new_[13450]_ , \new_[13451]_ , \new_[13454]_ , \new_[13458]_ ,
    \new_[13459]_ , \new_[13460]_ , \new_[13463]_ , \new_[13467]_ ,
    \new_[13468]_ , \new_[13469]_ , \new_[13472]_ , \new_[13476]_ ,
    \new_[13477]_ , \new_[13478]_ , \new_[13481]_ , \new_[13485]_ ,
    \new_[13486]_ , \new_[13487]_ , \new_[13490]_ , \new_[13494]_ ,
    \new_[13495]_ , \new_[13496]_ , \new_[13499]_ , \new_[13503]_ ,
    \new_[13504]_ , \new_[13505]_ , \new_[13508]_ , \new_[13512]_ ,
    \new_[13513]_ , \new_[13514]_ , \new_[13517]_ , \new_[13521]_ ,
    \new_[13522]_ , \new_[13523]_ , \new_[13526]_ , \new_[13530]_ ,
    \new_[13531]_ , \new_[13532]_ , \new_[13535]_ , \new_[13539]_ ,
    \new_[13540]_ , \new_[13541]_ , \new_[13544]_ , \new_[13548]_ ,
    \new_[13549]_ , \new_[13550]_ , \new_[13553]_ , \new_[13557]_ ,
    \new_[13558]_ , \new_[13559]_ , \new_[13562]_ , \new_[13566]_ ,
    \new_[13567]_ , \new_[13568]_ , \new_[13571]_ , \new_[13575]_ ,
    \new_[13576]_ , \new_[13577]_ , \new_[13580]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13586]_ , \new_[13589]_ , \new_[13593]_ ,
    \new_[13594]_ , \new_[13595]_ , \new_[13598]_ , \new_[13602]_ ,
    \new_[13603]_ , \new_[13604]_ , \new_[13607]_ , \new_[13611]_ ,
    \new_[13612]_ , \new_[13613]_ , \new_[13616]_ , \new_[13620]_ ,
    \new_[13621]_ , \new_[13622]_ , \new_[13625]_ , \new_[13629]_ ,
    \new_[13630]_ , \new_[13631]_ , \new_[13634]_ , \new_[13638]_ ,
    \new_[13639]_ , \new_[13640]_ , \new_[13643]_ , \new_[13647]_ ,
    \new_[13648]_ , \new_[13649]_ , \new_[13652]_ , \new_[13656]_ ,
    \new_[13657]_ , \new_[13658]_ , \new_[13661]_ , \new_[13665]_ ,
    \new_[13666]_ , \new_[13667]_ , \new_[13670]_ , \new_[13674]_ ,
    \new_[13675]_ , \new_[13676]_ , \new_[13679]_ , \new_[13683]_ ,
    \new_[13684]_ , \new_[13685]_ , \new_[13688]_ , \new_[13692]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13697]_ , \new_[13701]_ ,
    \new_[13702]_ , \new_[13703]_ , \new_[13706]_ , \new_[13710]_ ,
    \new_[13711]_ , \new_[13712]_ , \new_[13715]_ , \new_[13719]_ ,
    \new_[13720]_ , \new_[13721]_ , \new_[13724]_ , \new_[13728]_ ,
    \new_[13729]_ , \new_[13730]_ , \new_[13733]_ , \new_[13737]_ ,
    \new_[13738]_ , \new_[13739]_ , \new_[13742]_ , \new_[13746]_ ,
    \new_[13747]_ , \new_[13748]_ , \new_[13751]_ , \new_[13755]_ ,
    \new_[13756]_ , \new_[13757]_ , \new_[13760]_ , \new_[13764]_ ,
    \new_[13765]_ , \new_[13766]_ , \new_[13769]_ , \new_[13773]_ ,
    \new_[13774]_ , \new_[13775]_ , \new_[13778]_ , \new_[13782]_ ,
    \new_[13783]_ , \new_[13784]_ , \new_[13787]_ , \new_[13791]_ ,
    \new_[13792]_ , \new_[13793]_ , \new_[13796]_ , \new_[13800]_ ,
    \new_[13801]_ , \new_[13802]_ , \new_[13805]_ , \new_[13809]_ ,
    \new_[13810]_ , \new_[13811]_ , \new_[13814]_ , \new_[13818]_ ,
    \new_[13819]_ , \new_[13820]_ , \new_[13823]_ , \new_[13827]_ ,
    \new_[13828]_ , \new_[13829]_ , \new_[13832]_ , \new_[13836]_ ,
    \new_[13837]_ , \new_[13838]_ , \new_[13841]_ , \new_[13845]_ ,
    \new_[13846]_ , \new_[13847]_ , \new_[13850]_ , \new_[13854]_ ,
    \new_[13855]_ , \new_[13856]_ , \new_[13859]_ , \new_[13863]_ ,
    \new_[13864]_ , \new_[13865]_ , \new_[13868]_ , \new_[13872]_ ,
    \new_[13873]_ , \new_[13874]_ , \new_[13877]_ , \new_[13881]_ ,
    \new_[13882]_ , \new_[13883]_ , \new_[13886]_ , \new_[13890]_ ,
    \new_[13891]_ , \new_[13892]_ , \new_[13895]_ , \new_[13899]_ ,
    \new_[13900]_ , \new_[13901]_ , \new_[13904]_ , \new_[13908]_ ,
    \new_[13909]_ , \new_[13910]_ , \new_[13913]_ , \new_[13917]_ ,
    \new_[13918]_ , \new_[13919]_ , \new_[13922]_ , \new_[13926]_ ,
    \new_[13927]_ , \new_[13928]_ , \new_[13931]_ , \new_[13935]_ ,
    \new_[13936]_ , \new_[13937]_ , \new_[13940]_ , \new_[13944]_ ,
    \new_[13945]_ , \new_[13946]_ , \new_[13949]_ , \new_[13953]_ ,
    \new_[13954]_ , \new_[13955]_ , \new_[13958]_ , \new_[13962]_ ,
    \new_[13963]_ , \new_[13964]_ , \new_[13967]_ , \new_[13971]_ ,
    \new_[13972]_ , \new_[13973]_ , \new_[13976]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13982]_ , \new_[13985]_ , \new_[13989]_ ,
    \new_[13990]_ , \new_[13991]_ , \new_[13994]_ , \new_[13998]_ ,
    \new_[13999]_ , \new_[14000]_ , \new_[14003]_ , \new_[14007]_ ,
    \new_[14008]_ , \new_[14009]_ , \new_[14012]_ , \new_[14016]_ ,
    \new_[14017]_ , \new_[14018]_ , \new_[14021]_ , \new_[14025]_ ,
    \new_[14026]_ , \new_[14027]_ , \new_[14030]_ , \new_[14034]_ ,
    \new_[14035]_ , \new_[14036]_ , \new_[14039]_ , \new_[14043]_ ,
    \new_[14044]_ , \new_[14045]_ , \new_[14048]_ , \new_[14052]_ ,
    \new_[14053]_ , \new_[14054]_ , \new_[14057]_ , \new_[14061]_ ,
    \new_[14062]_ , \new_[14063]_ , \new_[14066]_ , \new_[14070]_ ,
    \new_[14071]_ , \new_[14072]_ , \new_[14075]_ , \new_[14079]_ ,
    \new_[14080]_ , \new_[14081]_ , \new_[14084]_ , \new_[14088]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14093]_ , \new_[14097]_ ,
    \new_[14098]_ , \new_[14099]_ , \new_[14102]_ , \new_[14106]_ ,
    \new_[14107]_ , \new_[14108]_ , \new_[14111]_ , \new_[14115]_ ,
    \new_[14116]_ , \new_[14117]_ , \new_[14120]_ , \new_[14124]_ ,
    \new_[14125]_ , \new_[14126]_ , \new_[14129]_ , \new_[14133]_ ,
    \new_[14134]_ , \new_[14135]_ , \new_[14138]_ , \new_[14142]_ ,
    \new_[14143]_ , \new_[14144]_ , \new_[14147]_ , \new_[14151]_ ,
    \new_[14152]_ , \new_[14153]_ , \new_[14156]_ , \new_[14160]_ ,
    \new_[14161]_ , \new_[14162]_ , \new_[14165]_ , \new_[14169]_ ,
    \new_[14170]_ , \new_[14171]_ , \new_[14174]_ , \new_[14178]_ ,
    \new_[14179]_ , \new_[14180]_ , \new_[14183]_ , \new_[14187]_ ,
    \new_[14188]_ , \new_[14189]_ , \new_[14192]_ , \new_[14196]_ ,
    \new_[14197]_ , \new_[14198]_ , \new_[14201]_ , \new_[14205]_ ,
    \new_[14206]_ , \new_[14207]_ , \new_[14210]_ , \new_[14214]_ ,
    \new_[14215]_ , \new_[14216]_ , \new_[14219]_ , \new_[14223]_ ,
    \new_[14224]_ , \new_[14225]_ , \new_[14228]_ , \new_[14232]_ ,
    \new_[14233]_ , \new_[14234]_ , \new_[14237]_ , \new_[14241]_ ,
    \new_[14242]_ , \new_[14243]_ , \new_[14246]_ , \new_[14250]_ ,
    \new_[14251]_ , \new_[14252]_ , \new_[14255]_ , \new_[14259]_ ,
    \new_[14260]_ , \new_[14261]_ , \new_[14264]_ , \new_[14268]_ ,
    \new_[14269]_ , \new_[14270]_ , \new_[14273]_ , \new_[14277]_ ,
    \new_[14278]_ , \new_[14279]_ , \new_[14282]_ , \new_[14286]_ ,
    \new_[14287]_ , \new_[14288]_ , \new_[14291]_ , \new_[14295]_ ,
    \new_[14296]_ , \new_[14297]_ , \new_[14300]_ , \new_[14304]_ ,
    \new_[14305]_ , \new_[14306]_ , \new_[14309]_ , \new_[14313]_ ,
    \new_[14314]_ , \new_[14315]_ , \new_[14318]_ , \new_[14322]_ ,
    \new_[14323]_ , \new_[14324]_ , \new_[14327]_ , \new_[14331]_ ,
    \new_[14332]_ , \new_[14333]_ , \new_[14336]_ , \new_[14340]_ ,
    \new_[14341]_ , \new_[14342]_ , \new_[14345]_ , \new_[14349]_ ,
    \new_[14350]_ , \new_[14351]_ , \new_[14354]_ , \new_[14358]_ ,
    \new_[14359]_ , \new_[14360]_ , \new_[14363]_ , \new_[14367]_ ,
    \new_[14368]_ , \new_[14369]_ , \new_[14372]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14378]_ , \new_[14381]_ , \new_[14385]_ ,
    \new_[14386]_ , \new_[14387]_ , \new_[14390]_ , \new_[14394]_ ,
    \new_[14395]_ , \new_[14396]_ , \new_[14399]_ , \new_[14403]_ ,
    \new_[14404]_ , \new_[14405]_ , \new_[14408]_ , \new_[14412]_ ,
    \new_[14413]_ , \new_[14414]_ , \new_[14417]_ , \new_[14421]_ ,
    \new_[14422]_ , \new_[14423]_ , \new_[14426]_ , \new_[14430]_ ,
    \new_[14431]_ , \new_[14432]_ , \new_[14435]_ , \new_[14439]_ ,
    \new_[14440]_ , \new_[14441]_ , \new_[14444]_ , \new_[14448]_ ,
    \new_[14449]_ , \new_[14450]_ , \new_[14453]_ , \new_[14457]_ ,
    \new_[14458]_ , \new_[14459]_ , \new_[14462]_ , \new_[14466]_ ,
    \new_[14467]_ , \new_[14468]_ , \new_[14471]_ , \new_[14475]_ ,
    \new_[14476]_ , \new_[14477]_ , \new_[14480]_ , \new_[14484]_ ,
    \new_[14485]_ , \new_[14486]_ , \new_[14489]_ , \new_[14493]_ ,
    \new_[14494]_ , \new_[14495]_ , \new_[14498]_ , \new_[14502]_ ,
    \new_[14503]_ , \new_[14504]_ , \new_[14507]_ , \new_[14511]_ ,
    \new_[14512]_ , \new_[14513]_ , \new_[14516]_ , \new_[14520]_ ,
    \new_[14521]_ , \new_[14522]_ , \new_[14525]_ , \new_[14529]_ ,
    \new_[14530]_ , \new_[14531]_ , \new_[14534]_ , \new_[14538]_ ,
    \new_[14539]_ , \new_[14540]_ , \new_[14543]_ , \new_[14547]_ ,
    \new_[14548]_ , \new_[14549]_ , \new_[14552]_ , \new_[14556]_ ,
    \new_[14557]_ , \new_[14558]_ , \new_[14561]_ , \new_[14565]_ ,
    \new_[14566]_ , \new_[14567]_ , \new_[14570]_ , \new_[14574]_ ,
    \new_[14575]_ , \new_[14576]_ , \new_[14579]_ , \new_[14583]_ ,
    \new_[14584]_ , \new_[14585]_ , \new_[14588]_ , \new_[14592]_ ,
    \new_[14593]_ , \new_[14594]_ , \new_[14597]_ , \new_[14601]_ ,
    \new_[14602]_ , \new_[14603]_ , \new_[14606]_ , \new_[14610]_ ,
    \new_[14611]_ , \new_[14612]_ , \new_[14615]_ , \new_[14619]_ ,
    \new_[14620]_ , \new_[14621]_ , \new_[14624]_ , \new_[14628]_ ,
    \new_[14629]_ , \new_[14630]_ , \new_[14633]_ , \new_[14637]_ ,
    \new_[14638]_ , \new_[14639]_ , \new_[14642]_ , \new_[14646]_ ,
    \new_[14647]_ , \new_[14648]_ , \new_[14651]_ , \new_[14655]_ ,
    \new_[14656]_ , \new_[14657]_ , \new_[14660]_ , \new_[14664]_ ,
    \new_[14665]_ , \new_[14666]_ , \new_[14669]_ , \new_[14673]_ ,
    \new_[14674]_ , \new_[14675]_ , \new_[14678]_ , \new_[14682]_ ,
    \new_[14683]_ , \new_[14684]_ , \new_[14687]_ , \new_[14691]_ ,
    \new_[14692]_ , \new_[14693]_ , \new_[14696]_ , \new_[14700]_ ,
    \new_[14701]_ , \new_[14702]_ , \new_[14705]_ , \new_[14709]_ ,
    \new_[14710]_ , \new_[14711]_ , \new_[14714]_ , \new_[14718]_ ,
    \new_[14719]_ , \new_[14720]_ , \new_[14723]_ , \new_[14727]_ ,
    \new_[14728]_ , \new_[14729]_ , \new_[14732]_ , \new_[14736]_ ,
    \new_[14737]_ , \new_[14738]_ , \new_[14741]_ , \new_[14745]_ ,
    \new_[14746]_ , \new_[14747]_ , \new_[14750]_ , \new_[14754]_ ,
    \new_[14755]_ , \new_[14756]_ , \new_[14759]_ , \new_[14763]_ ,
    \new_[14764]_ , \new_[14765]_ , \new_[14768]_ , \new_[14772]_ ,
    \new_[14773]_ , \new_[14774]_ , \new_[14777]_ , \new_[14781]_ ,
    \new_[14782]_ , \new_[14783]_ , \new_[14786]_ , \new_[14790]_ ,
    \new_[14791]_ , \new_[14792]_ , \new_[14795]_ , \new_[14799]_ ,
    \new_[14800]_ , \new_[14801]_ , \new_[14804]_ , \new_[14808]_ ,
    \new_[14809]_ , \new_[14810]_ , \new_[14813]_ , \new_[14817]_ ,
    \new_[14818]_ , \new_[14819]_ , \new_[14822]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14831]_ , \new_[14835]_ ,
    \new_[14836]_ , \new_[14837]_ , \new_[14840]_ , \new_[14844]_ ,
    \new_[14845]_ , \new_[14846]_ , \new_[14849]_ , \new_[14853]_ ,
    \new_[14854]_ , \new_[14855]_ , \new_[14858]_ , \new_[14862]_ ,
    \new_[14863]_ , \new_[14864]_ , \new_[14867]_ , \new_[14871]_ ,
    \new_[14872]_ , \new_[14873]_ , \new_[14876]_ , \new_[14880]_ ,
    \new_[14881]_ , \new_[14882]_ , \new_[14885]_ , \new_[14889]_ ,
    \new_[14890]_ , \new_[14891]_ , \new_[14894]_ , \new_[14898]_ ,
    \new_[14899]_ , \new_[14900]_ , \new_[14903]_ , \new_[14907]_ ,
    \new_[14908]_ , \new_[14909]_ , \new_[14912]_ , \new_[14916]_ ,
    \new_[14917]_ , \new_[14918]_ , \new_[14921]_ , \new_[14925]_ ,
    \new_[14926]_ , \new_[14927]_ , \new_[14930]_ , \new_[14934]_ ,
    \new_[14935]_ , \new_[14936]_ , \new_[14939]_ , \new_[14943]_ ,
    \new_[14944]_ , \new_[14945]_ , \new_[14948]_ , \new_[14952]_ ,
    \new_[14953]_ , \new_[14954]_ , \new_[14957]_ , \new_[14961]_ ,
    \new_[14962]_ , \new_[14963]_ , \new_[14966]_ , \new_[14970]_ ,
    \new_[14971]_ , \new_[14972]_ , \new_[14975]_ , \new_[14979]_ ,
    \new_[14980]_ , \new_[14981]_ , \new_[14984]_ , \new_[14988]_ ,
    \new_[14989]_ , \new_[14990]_ , \new_[14993]_ , \new_[14997]_ ,
    \new_[14998]_ , \new_[14999]_ , \new_[15002]_ , \new_[15006]_ ,
    \new_[15007]_ , \new_[15008]_ , \new_[15011]_ , \new_[15015]_ ,
    \new_[15016]_ , \new_[15017]_ , \new_[15020]_ , \new_[15024]_ ,
    \new_[15025]_ , \new_[15026]_ , \new_[15029]_ , \new_[15033]_ ,
    \new_[15034]_ , \new_[15035]_ , \new_[15038]_ , \new_[15042]_ ,
    \new_[15043]_ , \new_[15044]_ , \new_[15047]_ , \new_[15051]_ ,
    \new_[15052]_ , \new_[15053]_ , \new_[15056]_ , \new_[15060]_ ,
    \new_[15061]_ , \new_[15062]_ , \new_[15065]_ , \new_[15069]_ ,
    \new_[15070]_ , \new_[15071]_ , \new_[15074]_ , \new_[15078]_ ,
    \new_[15079]_ , \new_[15080]_ , \new_[15083]_ , \new_[15087]_ ,
    \new_[15088]_ , \new_[15089]_ , \new_[15092]_ , \new_[15096]_ ,
    \new_[15097]_ , \new_[15098]_ , \new_[15101]_ , \new_[15105]_ ,
    \new_[15106]_ , \new_[15107]_ , \new_[15110]_ , \new_[15114]_ ,
    \new_[15115]_ , \new_[15116]_ , \new_[15119]_ , \new_[15123]_ ,
    \new_[15124]_ , \new_[15125]_ , \new_[15128]_ , \new_[15132]_ ,
    \new_[15133]_ , \new_[15134]_ , \new_[15137]_ , \new_[15141]_ ,
    \new_[15142]_ , \new_[15143]_ , \new_[15146]_ , \new_[15150]_ ,
    \new_[15151]_ , \new_[15152]_ , \new_[15155]_ , \new_[15159]_ ,
    \new_[15160]_ , \new_[15161]_ , \new_[15164]_ , \new_[15168]_ ,
    \new_[15169]_ , \new_[15170]_ , \new_[15173]_ , \new_[15177]_ ,
    \new_[15178]_ , \new_[15179]_ , \new_[15182]_ , \new_[15186]_ ,
    \new_[15187]_ , \new_[15188]_ , \new_[15191]_ , \new_[15195]_ ,
    \new_[15196]_ , \new_[15197]_ , \new_[15200]_ , \new_[15204]_ ,
    \new_[15205]_ , \new_[15206]_ , \new_[15209]_ , \new_[15213]_ ,
    \new_[15214]_ , \new_[15215]_ , \new_[15218]_ , \new_[15222]_ ,
    \new_[15223]_ , \new_[15224]_ , \new_[15227]_ , \new_[15231]_ ,
    \new_[15232]_ , \new_[15233]_ , \new_[15236]_ , \new_[15240]_ ,
    \new_[15241]_ , \new_[15242]_ , \new_[15245]_ , \new_[15249]_ ,
    \new_[15250]_ , \new_[15251]_ , \new_[15254]_ , \new_[15258]_ ,
    \new_[15259]_ , \new_[15260]_ , \new_[15263]_ , \new_[15267]_ ,
    \new_[15268]_ , \new_[15269]_ , \new_[15272]_ , \new_[15276]_ ,
    \new_[15277]_ , \new_[15278]_ , \new_[15281]_ , \new_[15285]_ ,
    \new_[15286]_ , \new_[15287]_ , \new_[15290]_ , \new_[15294]_ ,
    \new_[15295]_ , \new_[15296]_ , \new_[15299]_ , \new_[15303]_ ,
    \new_[15304]_ , \new_[15305]_ , \new_[15308]_ , \new_[15312]_ ,
    \new_[15313]_ , \new_[15314]_ , \new_[15317]_ , \new_[15321]_ ,
    \new_[15322]_ , \new_[15323]_ , \new_[15326]_ , \new_[15330]_ ,
    \new_[15331]_ , \new_[15332]_ , \new_[15335]_ , \new_[15339]_ ,
    \new_[15340]_ , \new_[15341]_ , \new_[15344]_ , \new_[15348]_ ,
    \new_[15349]_ , \new_[15350]_ , \new_[15353]_ , \new_[15357]_ ,
    \new_[15358]_ , \new_[15359]_ , \new_[15362]_ , \new_[15366]_ ,
    \new_[15367]_ , \new_[15368]_ , \new_[15371]_ , \new_[15375]_ ,
    \new_[15376]_ , \new_[15377]_ , \new_[15380]_ , \new_[15384]_ ,
    \new_[15385]_ , \new_[15386]_ , \new_[15389]_ , \new_[15393]_ ,
    \new_[15394]_ , \new_[15395]_ , \new_[15398]_ , \new_[15402]_ ,
    \new_[15403]_ , \new_[15404]_ , \new_[15407]_ , \new_[15411]_ ,
    \new_[15412]_ , \new_[15413]_ , \new_[15416]_ , \new_[15420]_ ,
    \new_[15421]_ , \new_[15422]_ , \new_[15425]_ , \new_[15429]_ ,
    \new_[15430]_ , \new_[15431]_ , \new_[15434]_ , \new_[15438]_ ,
    \new_[15439]_ , \new_[15440]_ , \new_[15443]_ , \new_[15447]_ ,
    \new_[15448]_ , \new_[15449]_ , \new_[15452]_ , \new_[15456]_ ,
    \new_[15457]_ , \new_[15458]_ , \new_[15461]_ , \new_[15465]_ ,
    \new_[15466]_ , \new_[15467]_ , \new_[15470]_ , \new_[15474]_ ,
    \new_[15475]_ , \new_[15476]_ , \new_[15479]_ , \new_[15483]_ ,
    \new_[15484]_ , \new_[15485]_ , \new_[15488]_ , \new_[15492]_ ,
    \new_[15493]_ , \new_[15494]_ , \new_[15497]_ , \new_[15501]_ ,
    \new_[15502]_ , \new_[15503]_ , \new_[15506]_ , \new_[15510]_ ,
    \new_[15511]_ , \new_[15512]_ , \new_[15515]_ , \new_[15519]_ ,
    \new_[15520]_ , \new_[15521]_ , \new_[15524]_ , \new_[15528]_ ,
    \new_[15529]_ , \new_[15530]_ , \new_[15533]_ , \new_[15537]_ ,
    \new_[15538]_ , \new_[15539]_ , \new_[15542]_ , \new_[15546]_ ,
    \new_[15547]_ , \new_[15548]_ , \new_[15551]_ , \new_[15555]_ ,
    \new_[15556]_ , \new_[15557]_ , \new_[15560]_ , \new_[15564]_ ,
    \new_[15565]_ , \new_[15566]_ , \new_[15569]_ , \new_[15573]_ ,
    \new_[15574]_ , \new_[15575]_ , \new_[15578]_ , \new_[15582]_ ,
    \new_[15583]_ , \new_[15584]_ , \new_[15587]_ , \new_[15591]_ ,
    \new_[15592]_ , \new_[15593]_ , \new_[15596]_ , \new_[15600]_ ,
    \new_[15601]_ , \new_[15602]_ , \new_[15605]_ , \new_[15609]_ ,
    \new_[15610]_ , \new_[15611]_ , \new_[15614]_ , \new_[15618]_ ,
    \new_[15619]_ , \new_[15620]_ , \new_[15623]_ , \new_[15627]_ ,
    \new_[15628]_ , \new_[15629]_ , \new_[15632]_ , \new_[15636]_ ,
    \new_[15637]_ , \new_[15638]_ , \new_[15641]_ , \new_[15645]_ ,
    \new_[15646]_ , \new_[15647]_ , \new_[15650]_ , \new_[15654]_ ,
    \new_[15655]_ , \new_[15656]_ , \new_[15659]_ , \new_[15663]_ ,
    \new_[15664]_ , \new_[15665]_ , \new_[15668]_ , \new_[15672]_ ,
    \new_[15673]_ , \new_[15674]_ , \new_[15677]_ , \new_[15681]_ ,
    \new_[15682]_ , \new_[15683]_ , \new_[15686]_ , \new_[15690]_ ,
    \new_[15691]_ , \new_[15692]_ , \new_[15695]_ , \new_[15699]_ ,
    \new_[15700]_ , \new_[15701]_ , \new_[15704]_ , \new_[15708]_ ,
    \new_[15709]_ , \new_[15710]_ , \new_[15713]_ , \new_[15717]_ ,
    \new_[15718]_ , \new_[15719]_ , \new_[15722]_ , \new_[15726]_ ,
    \new_[15727]_ , \new_[15728]_ , \new_[15731]_ , \new_[15735]_ ,
    \new_[15736]_ , \new_[15737]_ , \new_[15740]_ , \new_[15744]_ ,
    \new_[15745]_ , \new_[15746]_ , \new_[15749]_ , \new_[15753]_ ,
    \new_[15754]_ , \new_[15755]_ , \new_[15758]_ , \new_[15762]_ ,
    \new_[15763]_ , \new_[15764]_ , \new_[15767]_ , \new_[15771]_ ,
    \new_[15772]_ , \new_[15773]_ , \new_[15776]_ , \new_[15780]_ ,
    \new_[15781]_ , \new_[15782]_ , \new_[15785]_ , \new_[15789]_ ,
    \new_[15790]_ , \new_[15791]_ , \new_[15794]_ , \new_[15798]_ ,
    \new_[15799]_ , \new_[15800]_ , \new_[15803]_ , \new_[15807]_ ,
    \new_[15808]_ , \new_[15809]_ , \new_[15812]_ , \new_[15816]_ ,
    \new_[15817]_ , \new_[15818]_ , \new_[15821]_ , \new_[15825]_ ,
    \new_[15826]_ , \new_[15827]_ , \new_[15830]_ , \new_[15834]_ ,
    \new_[15835]_ , \new_[15836]_ , \new_[15839]_ , \new_[15843]_ ,
    \new_[15844]_ , \new_[15845]_ , \new_[15848]_ , \new_[15852]_ ,
    \new_[15853]_ , \new_[15854]_ , \new_[15857]_ , \new_[15861]_ ,
    \new_[15862]_ , \new_[15863]_ , \new_[15866]_ , \new_[15870]_ ,
    \new_[15871]_ , \new_[15872]_ , \new_[15875]_ , \new_[15879]_ ,
    \new_[15880]_ , \new_[15881]_ , \new_[15884]_ , \new_[15888]_ ,
    \new_[15889]_ , \new_[15890]_ , \new_[15893]_ , \new_[15897]_ ,
    \new_[15898]_ , \new_[15899]_ , \new_[15902]_ , \new_[15906]_ ,
    \new_[15907]_ , \new_[15908]_ , \new_[15911]_ , \new_[15915]_ ,
    \new_[15916]_ , \new_[15917]_ , \new_[15920]_ , \new_[15924]_ ,
    \new_[15925]_ , \new_[15926]_ , \new_[15929]_ , \new_[15933]_ ,
    \new_[15934]_ , \new_[15935]_ , \new_[15938]_ , \new_[15942]_ ,
    \new_[15943]_ , \new_[15944]_ , \new_[15947]_ , \new_[15951]_ ,
    \new_[15952]_ , \new_[15953]_ , \new_[15956]_ , \new_[15960]_ ,
    \new_[15961]_ , \new_[15962]_ , \new_[15965]_ , \new_[15969]_ ,
    \new_[15970]_ , \new_[15971]_ , \new_[15974]_ , \new_[15978]_ ,
    \new_[15979]_ , \new_[15980]_ , \new_[15983]_ , \new_[15987]_ ,
    \new_[15988]_ , \new_[15989]_ , \new_[15992]_ , \new_[15996]_ ,
    \new_[15997]_ , \new_[15998]_ , \new_[16001]_ , \new_[16005]_ ,
    \new_[16006]_ , \new_[16007]_ , \new_[16010]_ , \new_[16014]_ ,
    \new_[16015]_ , \new_[16016]_ , \new_[16019]_ , \new_[16023]_ ,
    \new_[16024]_ , \new_[16025]_ , \new_[16028]_ , \new_[16032]_ ,
    \new_[16033]_ , \new_[16034]_ , \new_[16037]_ , \new_[16041]_ ,
    \new_[16042]_ , \new_[16043]_ , \new_[16046]_ , \new_[16050]_ ,
    \new_[16051]_ , \new_[16052]_ , \new_[16055]_ , \new_[16059]_ ,
    \new_[16060]_ , \new_[16061]_ , \new_[16064]_ , \new_[16068]_ ,
    \new_[16069]_ , \new_[16070]_ , \new_[16073]_ , \new_[16077]_ ,
    \new_[16078]_ , \new_[16079]_ , \new_[16082]_ , \new_[16086]_ ,
    \new_[16087]_ , \new_[16088]_ , \new_[16091]_ , \new_[16095]_ ,
    \new_[16096]_ , \new_[16097]_ , \new_[16100]_ , \new_[16104]_ ,
    \new_[16105]_ , \new_[16106]_ , \new_[16109]_ , \new_[16113]_ ,
    \new_[16114]_ , \new_[16115]_ , \new_[16118]_ , \new_[16122]_ ,
    \new_[16123]_ , \new_[16124]_ , \new_[16127]_ , \new_[16131]_ ,
    \new_[16132]_ , \new_[16133]_ , \new_[16136]_ , \new_[16140]_ ,
    \new_[16141]_ , \new_[16142]_ , \new_[16145]_ , \new_[16149]_ ,
    \new_[16150]_ , \new_[16151]_ , \new_[16154]_ , \new_[16158]_ ,
    \new_[16159]_ , \new_[16160]_ , \new_[16163]_ , \new_[16167]_ ,
    \new_[16168]_ , \new_[16169]_ , \new_[16172]_ , \new_[16176]_ ,
    \new_[16177]_ , \new_[16178]_ , \new_[16181]_ , \new_[16185]_ ,
    \new_[16186]_ , \new_[16187]_ , \new_[16190]_ , \new_[16194]_ ,
    \new_[16195]_ , \new_[16196]_ , \new_[16199]_ , \new_[16203]_ ,
    \new_[16204]_ , \new_[16205]_ , \new_[16208]_ , \new_[16212]_ ,
    \new_[16213]_ , \new_[16214]_ , \new_[16217]_ , \new_[16221]_ ,
    \new_[16222]_ , \new_[16223]_ , \new_[16226]_ , \new_[16230]_ ,
    \new_[16231]_ , \new_[16232]_ , \new_[16235]_ , \new_[16239]_ ,
    \new_[16240]_ , \new_[16241]_ , \new_[16244]_ , \new_[16248]_ ,
    \new_[16249]_ , \new_[16250]_ , \new_[16253]_ , \new_[16257]_ ,
    \new_[16258]_ , \new_[16259]_ , \new_[16262]_ , \new_[16266]_ ,
    \new_[16267]_ , \new_[16268]_ , \new_[16271]_ , \new_[16275]_ ,
    \new_[16276]_ , \new_[16277]_ , \new_[16280]_ , \new_[16284]_ ,
    \new_[16285]_ , \new_[16286]_ , \new_[16289]_ , \new_[16293]_ ,
    \new_[16294]_ , \new_[16295]_ , \new_[16298]_ , \new_[16302]_ ,
    \new_[16303]_ , \new_[16304]_ , \new_[16307]_ , \new_[16311]_ ,
    \new_[16312]_ , \new_[16313]_ , \new_[16316]_ , \new_[16320]_ ,
    \new_[16321]_ , \new_[16322]_ , \new_[16325]_ , \new_[16329]_ ,
    \new_[16330]_ , \new_[16331]_ , \new_[16334]_ , \new_[16338]_ ,
    \new_[16339]_ , \new_[16340]_ , \new_[16343]_ , \new_[16347]_ ,
    \new_[16348]_ , \new_[16349]_ , \new_[16352]_ , \new_[16356]_ ,
    \new_[16357]_ , \new_[16358]_ , \new_[16361]_ , \new_[16365]_ ,
    \new_[16366]_ , \new_[16367]_ , \new_[16370]_ , \new_[16374]_ ,
    \new_[16375]_ , \new_[16376]_ , \new_[16379]_ , \new_[16383]_ ,
    \new_[16384]_ , \new_[16385]_ , \new_[16388]_ , \new_[16392]_ ,
    \new_[16393]_ , \new_[16394]_ , \new_[16397]_ , \new_[16401]_ ,
    \new_[16402]_ , \new_[16403]_ , \new_[16406]_ , \new_[16410]_ ,
    \new_[16411]_ , \new_[16412]_ , \new_[16415]_ , \new_[16419]_ ,
    \new_[16420]_ , \new_[16421]_ , \new_[16424]_ , \new_[16428]_ ,
    \new_[16429]_ , \new_[16430]_ , \new_[16433]_ , \new_[16437]_ ,
    \new_[16438]_ , \new_[16439]_ , \new_[16442]_ , \new_[16446]_ ,
    \new_[16447]_ , \new_[16448]_ , \new_[16451]_ , \new_[16455]_ ,
    \new_[16456]_ , \new_[16457]_ , \new_[16460]_ , \new_[16464]_ ,
    \new_[16465]_ , \new_[16466]_ , \new_[16469]_ , \new_[16473]_ ,
    \new_[16474]_ , \new_[16475]_ , \new_[16478]_ , \new_[16482]_ ,
    \new_[16483]_ , \new_[16484]_ , \new_[16487]_ , \new_[16491]_ ,
    \new_[16492]_ , \new_[16493]_ , \new_[16496]_ , \new_[16500]_ ,
    \new_[16501]_ , \new_[16502]_ , \new_[16505]_ , \new_[16509]_ ,
    \new_[16510]_ , \new_[16511]_ , \new_[16514]_ , \new_[16518]_ ,
    \new_[16519]_ , \new_[16520]_ , \new_[16523]_ , \new_[16527]_ ,
    \new_[16528]_ , \new_[16529]_ , \new_[16532]_ , \new_[16536]_ ,
    \new_[16537]_ , \new_[16538]_ , \new_[16541]_ , \new_[16545]_ ,
    \new_[16546]_ , \new_[16547]_ , \new_[16550]_ , \new_[16554]_ ,
    \new_[16555]_ , \new_[16556]_ , \new_[16559]_ , \new_[16563]_ ,
    \new_[16564]_ , \new_[16565]_ , \new_[16568]_ , \new_[16572]_ ,
    \new_[16573]_ , \new_[16574]_ , \new_[16577]_ , \new_[16581]_ ,
    \new_[16582]_ , \new_[16583]_ , \new_[16586]_ , \new_[16590]_ ,
    \new_[16591]_ , \new_[16592]_ , \new_[16595]_ , \new_[16599]_ ,
    \new_[16600]_ , \new_[16601]_ , \new_[16604]_ , \new_[16608]_ ,
    \new_[16609]_ , \new_[16610]_ , \new_[16613]_ , \new_[16617]_ ,
    \new_[16618]_ , \new_[16619]_ , \new_[16622]_ , \new_[16626]_ ,
    \new_[16627]_ , \new_[16628]_ , \new_[16631]_ , \new_[16635]_ ,
    \new_[16636]_ , \new_[16637]_ , \new_[16640]_ , \new_[16644]_ ,
    \new_[16645]_ , \new_[16646]_ , \new_[16649]_ , \new_[16653]_ ,
    \new_[16654]_ , \new_[16655]_ , \new_[16658]_ , \new_[16662]_ ,
    \new_[16663]_ , \new_[16664]_ , \new_[16667]_ , \new_[16671]_ ,
    \new_[16672]_ , \new_[16673]_ , \new_[16676]_ , \new_[16680]_ ,
    \new_[16681]_ , \new_[16682]_ , \new_[16685]_ , \new_[16689]_ ,
    \new_[16690]_ , \new_[16691]_ , \new_[16694]_ , \new_[16698]_ ,
    \new_[16699]_ , \new_[16700]_ , \new_[16703]_ , \new_[16707]_ ,
    \new_[16708]_ , \new_[16709]_ , \new_[16712]_ , \new_[16716]_ ,
    \new_[16717]_ , \new_[16718]_ , \new_[16721]_ , \new_[16725]_ ,
    \new_[16726]_ , \new_[16727]_ , \new_[16730]_ , \new_[16734]_ ,
    \new_[16735]_ , \new_[16736]_ , \new_[16739]_ , \new_[16743]_ ,
    \new_[16744]_ , \new_[16745]_ , \new_[16748]_ , \new_[16752]_ ,
    \new_[16753]_ , \new_[16754]_ , \new_[16757]_ , \new_[16761]_ ,
    \new_[16762]_ , \new_[16763]_ , \new_[16766]_ , \new_[16770]_ ,
    \new_[16771]_ , \new_[16772]_ , \new_[16775]_ , \new_[16779]_ ,
    \new_[16780]_ , \new_[16781]_ , \new_[16784]_ , \new_[16788]_ ,
    \new_[16789]_ , \new_[16790]_ , \new_[16793]_ , \new_[16797]_ ,
    \new_[16798]_ , \new_[16799]_ , \new_[16802]_ , \new_[16806]_ ,
    \new_[16807]_ , \new_[16808]_ , \new_[16811]_ , \new_[16815]_ ,
    \new_[16816]_ , \new_[16817]_ , \new_[16820]_ , \new_[16824]_ ,
    \new_[16825]_ , \new_[16826]_ , \new_[16829]_ , \new_[16833]_ ,
    \new_[16834]_ , \new_[16835]_ , \new_[16838]_ , \new_[16842]_ ,
    \new_[16843]_ , \new_[16844]_ , \new_[16847]_ , \new_[16851]_ ,
    \new_[16852]_ , \new_[16853]_ , \new_[16856]_ , \new_[16860]_ ,
    \new_[16861]_ , \new_[16862]_ , \new_[16865]_ , \new_[16869]_ ,
    \new_[16870]_ , \new_[16871]_ , \new_[16874]_ , \new_[16878]_ ,
    \new_[16879]_ , \new_[16880]_ , \new_[16883]_ , \new_[16887]_ ,
    \new_[16888]_ , \new_[16889]_ , \new_[16892]_ , \new_[16896]_ ,
    \new_[16897]_ , \new_[16898]_ , \new_[16901]_ , \new_[16905]_ ,
    \new_[16906]_ , \new_[16907]_ , \new_[16910]_ , \new_[16914]_ ,
    \new_[16915]_ , \new_[16916]_ , \new_[16919]_ , \new_[16923]_ ,
    \new_[16924]_ , \new_[16925]_ , \new_[16928]_ , \new_[16932]_ ,
    \new_[16933]_ , \new_[16934]_ , \new_[16937]_ , \new_[16941]_ ,
    \new_[16942]_ , \new_[16943]_ , \new_[16946]_ , \new_[16950]_ ,
    \new_[16951]_ , \new_[16952]_ , \new_[16955]_ , \new_[16959]_ ,
    \new_[16960]_ , \new_[16961]_ , \new_[16964]_ , \new_[16968]_ ,
    \new_[16969]_ , \new_[16970]_ , \new_[16973]_ , \new_[16977]_ ,
    \new_[16978]_ , \new_[16979]_ , \new_[16982]_ , \new_[16986]_ ,
    \new_[16987]_ , \new_[16988]_ , \new_[16991]_ , \new_[16995]_ ,
    \new_[16996]_ , \new_[16997]_ , \new_[17000]_ , \new_[17004]_ ,
    \new_[17005]_ , \new_[17006]_ , \new_[17009]_ , \new_[17013]_ ,
    \new_[17014]_ , \new_[17015]_ , \new_[17018]_ , \new_[17022]_ ,
    \new_[17023]_ , \new_[17024]_ , \new_[17027]_ , \new_[17031]_ ,
    \new_[17032]_ , \new_[17033]_ , \new_[17036]_ , \new_[17040]_ ,
    \new_[17041]_ , \new_[17042]_ , \new_[17045]_ , \new_[17049]_ ,
    \new_[17050]_ , \new_[17051]_ , \new_[17054]_ , \new_[17058]_ ,
    \new_[17059]_ , \new_[17060]_ , \new_[17063]_ , \new_[17067]_ ,
    \new_[17068]_ , \new_[17069]_ , \new_[17072]_ , \new_[17076]_ ,
    \new_[17077]_ , \new_[17078]_ , \new_[17081]_ , \new_[17085]_ ,
    \new_[17086]_ , \new_[17087]_ , \new_[17090]_ , \new_[17094]_ ,
    \new_[17095]_ , \new_[17096]_ , \new_[17099]_ , \new_[17103]_ ,
    \new_[17104]_ , \new_[17105]_ , \new_[17108]_ , \new_[17112]_ ,
    \new_[17113]_ , \new_[17114]_ , \new_[17117]_ , \new_[17121]_ ,
    \new_[17122]_ , \new_[17123]_ , \new_[17126]_ , \new_[17130]_ ,
    \new_[17131]_ , \new_[17132]_ , \new_[17135]_ , \new_[17139]_ ,
    \new_[17140]_ , \new_[17141]_ , \new_[17144]_ , \new_[17148]_ ,
    \new_[17149]_ , \new_[17150]_ , \new_[17153]_ , \new_[17157]_ ,
    \new_[17158]_ , \new_[17159]_ , \new_[17162]_ , \new_[17166]_ ,
    \new_[17167]_ , \new_[17168]_ , \new_[17171]_ , \new_[17175]_ ,
    \new_[17176]_ , \new_[17177]_ , \new_[17180]_ , \new_[17184]_ ,
    \new_[17185]_ , \new_[17186]_ , \new_[17189]_ , \new_[17193]_ ,
    \new_[17194]_ , \new_[17195]_ , \new_[17198]_ , \new_[17202]_ ,
    \new_[17203]_ , \new_[17204]_ , \new_[17207]_ , \new_[17211]_ ,
    \new_[17212]_ , \new_[17213]_ , \new_[17216]_ , \new_[17220]_ ,
    \new_[17221]_ , \new_[17222]_ , \new_[17225]_ , \new_[17229]_ ,
    \new_[17230]_ , \new_[17231]_ , \new_[17234]_ , \new_[17238]_ ,
    \new_[17239]_ , \new_[17240]_ , \new_[17243]_ , \new_[17247]_ ,
    \new_[17248]_ , \new_[17249]_ , \new_[17252]_ , \new_[17256]_ ,
    \new_[17257]_ , \new_[17258]_ , \new_[17261]_ , \new_[17265]_ ,
    \new_[17266]_ , \new_[17267]_ , \new_[17270]_ , \new_[17274]_ ,
    \new_[17275]_ , \new_[17276]_ , \new_[17279]_ , \new_[17283]_ ,
    \new_[17284]_ , \new_[17285]_ , \new_[17288]_ , \new_[17292]_ ,
    \new_[17293]_ , \new_[17294]_ , \new_[17297]_ , \new_[17301]_ ,
    \new_[17302]_ , \new_[17303]_ , \new_[17306]_ , \new_[17310]_ ,
    \new_[17311]_ , \new_[17312]_ , \new_[17315]_ , \new_[17319]_ ,
    \new_[17320]_ , \new_[17321]_ , \new_[17324]_ , \new_[17328]_ ,
    \new_[17329]_ , \new_[17330]_ , \new_[17333]_ , \new_[17337]_ ,
    \new_[17338]_ , \new_[17339]_ , \new_[17342]_ , \new_[17346]_ ,
    \new_[17347]_ , \new_[17348]_ , \new_[17351]_ , \new_[17355]_ ,
    \new_[17356]_ , \new_[17357]_ , \new_[17360]_ , \new_[17364]_ ,
    \new_[17365]_ , \new_[17366]_ , \new_[17369]_ , \new_[17373]_ ,
    \new_[17374]_ , \new_[17375]_ , \new_[17378]_ , \new_[17382]_ ,
    \new_[17383]_ , \new_[17384]_ , \new_[17387]_ , \new_[17391]_ ,
    \new_[17392]_ , \new_[17393]_ , \new_[17396]_ , \new_[17400]_ ,
    \new_[17401]_ , \new_[17402]_ , \new_[17405]_ , \new_[17409]_ ,
    \new_[17410]_ , \new_[17411]_ , \new_[17414]_ , \new_[17418]_ ,
    \new_[17419]_ , \new_[17420]_ , \new_[17423]_ , \new_[17427]_ ,
    \new_[17428]_ , \new_[17429]_ , \new_[17432]_ , \new_[17436]_ ,
    \new_[17437]_ , \new_[17438]_ , \new_[17441]_ , \new_[17445]_ ,
    \new_[17446]_ , \new_[17447]_ , \new_[17450]_ , \new_[17454]_ ,
    \new_[17455]_ , \new_[17456]_ , \new_[17459]_ , \new_[17463]_ ,
    \new_[17464]_ , \new_[17465]_ , \new_[17469]_ , \new_[17470]_ ,
    \new_[17474]_ , \new_[17475]_ , \new_[17476]_ , \new_[17479]_ ,
    \new_[17483]_ , \new_[17484]_ , \new_[17485]_ , \new_[17489]_ ,
    \new_[17490]_ , \new_[17494]_ , \new_[17495]_ , \new_[17496]_ ,
    \new_[17499]_ , \new_[17503]_ , \new_[17504]_ , \new_[17505]_ ,
    \new_[17509]_ , \new_[17510]_ , \new_[17514]_ , \new_[17515]_ ,
    \new_[17516]_ , \new_[17519]_ , \new_[17523]_ , \new_[17524]_ ,
    \new_[17525]_ , \new_[17529]_ , \new_[17530]_ , \new_[17534]_ ,
    \new_[17535]_ , \new_[17536]_ , \new_[17539]_ , \new_[17543]_ ,
    \new_[17544]_ , \new_[17545]_ , \new_[17549]_ , \new_[17550]_ ,
    \new_[17554]_ , \new_[17555]_ , \new_[17556]_ , \new_[17559]_ ,
    \new_[17563]_ , \new_[17564]_ , \new_[17565]_ , \new_[17569]_ ,
    \new_[17570]_ , \new_[17574]_ , \new_[17575]_ , \new_[17576]_ ,
    \new_[17579]_ , \new_[17583]_ , \new_[17584]_ , \new_[17585]_ ,
    \new_[17589]_ , \new_[17590]_ , \new_[17594]_ , \new_[17595]_ ,
    \new_[17596]_ , \new_[17599]_ , \new_[17603]_ , \new_[17604]_ ,
    \new_[17605]_ , \new_[17609]_ , \new_[17610]_ , \new_[17614]_ ,
    \new_[17615]_ , \new_[17616]_ , \new_[17619]_ , \new_[17623]_ ,
    \new_[17624]_ , \new_[17625]_ , \new_[17629]_ , \new_[17630]_ ,
    \new_[17634]_ , \new_[17635]_ , \new_[17636]_ , \new_[17639]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17645]_ , \new_[17649]_ ,
    \new_[17650]_ , \new_[17654]_ , \new_[17655]_ , \new_[17656]_ ,
    \new_[17659]_ , \new_[17663]_ , \new_[17664]_ , \new_[17665]_ ,
    \new_[17669]_ , \new_[17670]_ , \new_[17674]_ , \new_[17675]_ ,
    \new_[17676]_ , \new_[17679]_ , \new_[17683]_ , \new_[17684]_ ,
    \new_[17685]_ , \new_[17689]_ , \new_[17690]_ , \new_[17694]_ ,
    \new_[17695]_ , \new_[17696]_ , \new_[17699]_ , \new_[17703]_ ,
    \new_[17704]_ , \new_[17705]_ , \new_[17709]_ , \new_[17710]_ ,
    \new_[17714]_ , \new_[17715]_ , \new_[17716]_ , \new_[17719]_ ,
    \new_[17723]_ , \new_[17724]_ , \new_[17725]_ , \new_[17729]_ ,
    \new_[17730]_ , \new_[17734]_ , \new_[17735]_ , \new_[17736]_ ,
    \new_[17739]_ , \new_[17743]_ , \new_[17744]_ , \new_[17745]_ ,
    \new_[17749]_ , \new_[17750]_ , \new_[17754]_ , \new_[17755]_ ,
    \new_[17756]_ , \new_[17759]_ , \new_[17763]_ , \new_[17764]_ ,
    \new_[17765]_ , \new_[17769]_ , \new_[17770]_ , \new_[17774]_ ,
    \new_[17775]_ , \new_[17776]_ , \new_[17779]_ , \new_[17783]_ ,
    \new_[17784]_ , \new_[17785]_ , \new_[17789]_ , \new_[17790]_ ,
    \new_[17794]_ , \new_[17795]_ , \new_[17796]_ , \new_[17799]_ ,
    \new_[17803]_ , \new_[17804]_ , \new_[17805]_ , \new_[17809]_ ,
    \new_[17810]_ , \new_[17814]_ , \new_[17815]_ , \new_[17816]_ ,
    \new_[17819]_ , \new_[17823]_ , \new_[17824]_ , \new_[17825]_ ,
    \new_[17829]_ , \new_[17830]_ , \new_[17834]_ , \new_[17835]_ ,
    \new_[17836]_ , \new_[17839]_ , \new_[17843]_ , \new_[17844]_ ,
    \new_[17845]_ , \new_[17849]_ , \new_[17850]_ , \new_[17854]_ ,
    \new_[17855]_ , \new_[17856]_ , \new_[17859]_ , \new_[17863]_ ,
    \new_[17864]_ , \new_[17865]_ , \new_[17869]_ , \new_[17870]_ ,
    \new_[17874]_ , \new_[17875]_ , \new_[17876]_ , \new_[17879]_ ,
    \new_[17883]_ , \new_[17884]_ , \new_[17885]_ , \new_[17889]_ ,
    \new_[17890]_ , \new_[17894]_ , \new_[17895]_ , \new_[17896]_ ,
    \new_[17899]_ , \new_[17903]_ , \new_[17904]_ , \new_[17905]_ ,
    \new_[17909]_ , \new_[17910]_ , \new_[17914]_ , \new_[17915]_ ,
    \new_[17916]_ , \new_[17919]_ , \new_[17923]_ , \new_[17924]_ ,
    \new_[17925]_ , \new_[17929]_ , \new_[17930]_ , \new_[17934]_ ,
    \new_[17935]_ , \new_[17936]_ , \new_[17939]_ , \new_[17943]_ ,
    \new_[17944]_ , \new_[17945]_ , \new_[17949]_ , \new_[17950]_ ,
    \new_[17954]_ , \new_[17955]_ , \new_[17956]_ , \new_[17959]_ ,
    \new_[17963]_ , \new_[17964]_ , \new_[17965]_ , \new_[17969]_ ,
    \new_[17970]_ , \new_[17974]_ , \new_[17975]_ , \new_[17976]_ ,
    \new_[17979]_ , \new_[17983]_ , \new_[17984]_ , \new_[17985]_ ,
    \new_[17989]_ , \new_[17990]_ , \new_[17994]_ , \new_[17995]_ ,
    \new_[17996]_ , \new_[17999]_ , \new_[18003]_ , \new_[18004]_ ,
    \new_[18005]_ , \new_[18009]_ , \new_[18010]_ , \new_[18014]_ ,
    \new_[18015]_ , \new_[18016]_ , \new_[18019]_ , \new_[18023]_ ,
    \new_[18024]_ , \new_[18025]_ , \new_[18029]_ , \new_[18030]_ ,
    \new_[18034]_ , \new_[18035]_ , \new_[18036]_ , \new_[18039]_ ,
    \new_[18043]_ , \new_[18044]_ , \new_[18045]_ , \new_[18049]_ ,
    \new_[18050]_ , \new_[18054]_ , \new_[18055]_ , \new_[18056]_ ,
    \new_[18059]_ , \new_[18063]_ , \new_[18064]_ , \new_[18065]_ ,
    \new_[18069]_ , \new_[18070]_ , \new_[18074]_ , \new_[18075]_ ,
    \new_[18076]_ , \new_[18079]_ , \new_[18083]_ , \new_[18084]_ ,
    \new_[18085]_ , \new_[18089]_ , \new_[18090]_ , \new_[18094]_ ,
    \new_[18095]_ , \new_[18096]_ , \new_[18099]_ , \new_[18103]_ ,
    \new_[18104]_ , \new_[18105]_ , \new_[18109]_ , \new_[18110]_ ,
    \new_[18114]_ , \new_[18115]_ , \new_[18116]_ , \new_[18119]_ ,
    \new_[18123]_ , \new_[18124]_ , \new_[18125]_ , \new_[18129]_ ,
    \new_[18130]_ , \new_[18134]_ , \new_[18135]_ , \new_[18136]_ ,
    \new_[18139]_ , \new_[18143]_ , \new_[18144]_ , \new_[18145]_ ,
    \new_[18149]_ , \new_[18150]_ , \new_[18154]_ , \new_[18155]_ ,
    \new_[18156]_ , \new_[18159]_ , \new_[18163]_ , \new_[18164]_ ,
    \new_[18165]_ , \new_[18169]_ , \new_[18170]_ , \new_[18174]_ ,
    \new_[18175]_ , \new_[18176]_ , \new_[18179]_ , \new_[18183]_ ,
    \new_[18184]_ , \new_[18185]_ , \new_[18189]_ , \new_[18190]_ ,
    \new_[18194]_ , \new_[18195]_ , \new_[18196]_ , \new_[18199]_ ,
    \new_[18203]_ , \new_[18204]_ , \new_[18205]_ , \new_[18209]_ ,
    \new_[18210]_ , \new_[18214]_ , \new_[18215]_ , \new_[18216]_ ,
    \new_[18219]_ , \new_[18223]_ , \new_[18224]_ , \new_[18225]_ ,
    \new_[18229]_ , \new_[18230]_ , \new_[18234]_ , \new_[18235]_ ,
    \new_[18236]_ , \new_[18239]_ , \new_[18243]_ , \new_[18244]_ ,
    \new_[18245]_ , \new_[18249]_ , \new_[18250]_ , \new_[18254]_ ,
    \new_[18255]_ , \new_[18256]_ , \new_[18259]_ , \new_[18263]_ ,
    \new_[18264]_ , \new_[18265]_ , \new_[18269]_ , \new_[18270]_ ,
    \new_[18274]_ , \new_[18275]_ , \new_[18276]_ , \new_[18279]_ ,
    \new_[18283]_ , \new_[18284]_ , \new_[18285]_ , \new_[18289]_ ,
    \new_[18290]_ , \new_[18294]_ , \new_[18295]_ , \new_[18296]_ ,
    \new_[18299]_ , \new_[18303]_ , \new_[18304]_ , \new_[18305]_ ,
    \new_[18309]_ , \new_[18310]_ , \new_[18314]_ , \new_[18315]_ ,
    \new_[18316]_ , \new_[18319]_ , \new_[18323]_ , \new_[18324]_ ,
    \new_[18325]_ , \new_[18329]_ , \new_[18330]_ , \new_[18334]_ ,
    \new_[18335]_ , \new_[18336]_ , \new_[18339]_ , \new_[18343]_ ,
    \new_[18344]_ , \new_[18345]_ , \new_[18349]_ , \new_[18350]_ ,
    \new_[18354]_ , \new_[18355]_ , \new_[18356]_ , \new_[18359]_ ,
    \new_[18363]_ , \new_[18364]_ , \new_[18365]_ , \new_[18369]_ ,
    \new_[18370]_ , \new_[18374]_ , \new_[18375]_ , \new_[18376]_ ,
    \new_[18379]_ , \new_[18383]_ , \new_[18384]_ , \new_[18385]_ ,
    \new_[18389]_ , \new_[18390]_ , \new_[18394]_ , \new_[18395]_ ,
    \new_[18396]_ , \new_[18399]_ , \new_[18403]_ , \new_[18404]_ ,
    \new_[18405]_ , \new_[18409]_ , \new_[18410]_ , \new_[18414]_ ,
    \new_[18415]_ , \new_[18416]_ , \new_[18419]_ , \new_[18423]_ ,
    \new_[18424]_ , \new_[18425]_ , \new_[18429]_ , \new_[18430]_ ,
    \new_[18434]_ , \new_[18435]_ , \new_[18436]_ , \new_[18439]_ ,
    \new_[18443]_ , \new_[18444]_ , \new_[18445]_ , \new_[18449]_ ,
    \new_[18450]_ , \new_[18454]_ , \new_[18455]_ , \new_[18456]_ ,
    \new_[18459]_ , \new_[18463]_ , \new_[18464]_ , \new_[18465]_ ,
    \new_[18469]_ , \new_[18470]_ , \new_[18474]_ , \new_[18475]_ ,
    \new_[18476]_ , \new_[18479]_ , \new_[18483]_ , \new_[18484]_ ,
    \new_[18485]_ , \new_[18489]_ , \new_[18490]_ , \new_[18494]_ ,
    \new_[18495]_ , \new_[18496]_ , \new_[18499]_ , \new_[18503]_ ,
    \new_[18504]_ , \new_[18505]_ , \new_[18509]_ , \new_[18510]_ ,
    \new_[18514]_ , \new_[18515]_ , \new_[18516]_ , \new_[18519]_ ,
    \new_[18523]_ , \new_[18524]_ , \new_[18525]_ , \new_[18529]_ ,
    \new_[18530]_ , \new_[18534]_ , \new_[18535]_ , \new_[18536]_ ,
    \new_[18539]_ , \new_[18543]_ , \new_[18544]_ , \new_[18545]_ ,
    \new_[18549]_ , \new_[18550]_ , \new_[18554]_ , \new_[18555]_ ,
    \new_[18556]_ , \new_[18559]_ , \new_[18563]_ , \new_[18564]_ ,
    \new_[18565]_ , \new_[18569]_ , \new_[18570]_ , \new_[18574]_ ,
    \new_[18575]_ , \new_[18576]_ , \new_[18579]_ , \new_[18583]_ ,
    \new_[18584]_ , \new_[18585]_ , \new_[18589]_ , \new_[18590]_ ,
    \new_[18594]_ , \new_[18595]_ , \new_[18596]_ , \new_[18599]_ ,
    \new_[18603]_ , \new_[18604]_ , \new_[18605]_ , \new_[18609]_ ,
    \new_[18610]_ , \new_[18614]_ , \new_[18615]_ , \new_[18616]_ ,
    \new_[18619]_ , \new_[18623]_ , \new_[18624]_ , \new_[18625]_ ,
    \new_[18629]_ , \new_[18630]_ , \new_[18634]_ , \new_[18635]_ ,
    \new_[18636]_ , \new_[18639]_ , \new_[18643]_ , \new_[18644]_ ,
    \new_[18645]_ , \new_[18649]_ , \new_[18650]_ , \new_[18654]_ ,
    \new_[18655]_ , \new_[18656]_ , \new_[18659]_ , \new_[18663]_ ,
    \new_[18664]_ , \new_[18665]_ , \new_[18669]_ , \new_[18670]_ ,
    \new_[18674]_ , \new_[18675]_ , \new_[18676]_ , \new_[18679]_ ,
    \new_[18683]_ , \new_[18684]_ , \new_[18685]_ , \new_[18689]_ ,
    \new_[18690]_ , \new_[18694]_ , \new_[18695]_ , \new_[18696]_ ,
    \new_[18699]_ , \new_[18703]_ , \new_[18704]_ , \new_[18705]_ ,
    \new_[18709]_ , \new_[18710]_ , \new_[18714]_ , \new_[18715]_ ,
    \new_[18716]_ , \new_[18719]_ , \new_[18723]_ , \new_[18724]_ ,
    \new_[18725]_ , \new_[18729]_ , \new_[18730]_ , \new_[18734]_ ,
    \new_[18735]_ , \new_[18736]_ , \new_[18739]_ , \new_[18743]_ ,
    \new_[18744]_ , \new_[18745]_ , \new_[18749]_ , \new_[18750]_ ,
    \new_[18754]_ , \new_[18755]_ , \new_[18756]_ , \new_[18759]_ ,
    \new_[18763]_ , \new_[18764]_ , \new_[18765]_ , \new_[18769]_ ,
    \new_[18770]_ , \new_[18774]_ , \new_[18775]_ , \new_[18776]_ ,
    \new_[18779]_ , \new_[18783]_ , \new_[18784]_ , \new_[18785]_ ,
    \new_[18789]_ , \new_[18790]_ , \new_[18794]_ , \new_[18795]_ ,
    \new_[18796]_ , \new_[18799]_ , \new_[18803]_ , \new_[18804]_ ,
    \new_[18805]_ , \new_[18809]_ , \new_[18810]_ , \new_[18814]_ ,
    \new_[18815]_ , \new_[18816]_ , \new_[18819]_ , \new_[18823]_ ,
    \new_[18824]_ , \new_[18825]_ , \new_[18829]_ , \new_[18830]_ ,
    \new_[18834]_ , \new_[18835]_ , \new_[18836]_ , \new_[18839]_ ,
    \new_[18843]_ , \new_[18844]_ , \new_[18845]_ , \new_[18849]_ ,
    \new_[18850]_ , \new_[18854]_ , \new_[18855]_ , \new_[18856]_ ,
    \new_[18859]_ , \new_[18863]_ , \new_[18864]_ , \new_[18865]_ ,
    \new_[18869]_ , \new_[18870]_ , \new_[18874]_ , \new_[18875]_ ,
    \new_[18876]_ , \new_[18879]_ , \new_[18883]_ , \new_[18884]_ ,
    \new_[18885]_ , \new_[18889]_ , \new_[18890]_ , \new_[18894]_ ,
    \new_[18895]_ , \new_[18896]_ , \new_[18899]_ , \new_[18903]_ ,
    \new_[18904]_ , \new_[18905]_ , \new_[18909]_ , \new_[18910]_ ,
    \new_[18914]_ , \new_[18915]_ , \new_[18916]_ , \new_[18919]_ ,
    \new_[18923]_ , \new_[18924]_ , \new_[18925]_ , \new_[18929]_ ,
    \new_[18930]_ , \new_[18934]_ , \new_[18935]_ , \new_[18936]_ ,
    \new_[18939]_ , \new_[18943]_ , \new_[18944]_ , \new_[18945]_ ,
    \new_[18949]_ , \new_[18950]_ , \new_[18954]_ , \new_[18955]_ ,
    \new_[18956]_ , \new_[18959]_ , \new_[18963]_ , \new_[18964]_ ,
    \new_[18965]_ , \new_[18969]_ , \new_[18970]_ , \new_[18974]_ ,
    \new_[18975]_ , \new_[18976]_ , \new_[18979]_ , \new_[18983]_ ,
    \new_[18984]_ , \new_[18985]_ , \new_[18989]_ , \new_[18990]_ ,
    \new_[18994]_ , \new_[18995]_ , \new_[18996]_ , \new_[18999]_ ,
    \new_[19003]_ , \new_[19004]_ , \new_[19005]_ , \new_[19009]_ ,
    \new_[19010]_ , \new_[19014]_ , \new_[19015]_ , \new_[19016]_ ,
    \new_[19019]_ , \new_[19023]_ , \new_[19024]_ , \new_[19025]_ ,
    \new_[19029]_ , \new_[19030]_ , \new_[19034]_ , \new_[19035]_ ,
    \new_[19036]_ , \new_[19039]_ , \new_[19043]_ , \new_[19044]_ ,
    \new_[19045]_ , \new_[19049]_ , \new_[19050]_ , \new_[19054]_ ,
    \new_[19055]_ , \new_[19056]_ , \new_[19059]_ , \new_[19063]_ ,
    \new_[19064]_ , \new_[19065]_ , \new_[19069]_ , \new_[19070]_ ,
    \new_[19074]_ , \new_[19075]_ , \new_[19076]_ , \new_[19079]_ ,
    \new_[19083]_ , \new_[19084]_ , \new_[19085]_ , \new_[19089]_ ,
    \new_[19090]_ , \new_[19094]_ , \new_[19095]_ , \new_[19096]_ ,
    \new_[19099]_ , \new_[19103]_ , \new_[19104]_ , \new_[19105]_ ,
    \new_[19109]_ , \new_[19110]_ , \new_[19114]_ , \new_[19115]_ ,
    \new_[19116]_ , \new_[19119]_ , \new_[19123]_ , \new_[19124]_ ,
    \new_[19125]_ , \new_[19129]_ , \new_[19130]_ , \new_[19134]_ ,
    \new_[19135]_ , \new_[19136]_ , \new_[19139]_ , \new_[19143]_ ,
    \new_[19144]_ , \new_[19145]_ , \new_[19149]_ , \new_[19150]_ ,
    \new_[19154]_ , \new_[19155]_ , \new_[19156]_ , \new_[19159]_ ,
    \new_[19163]_ , \new_[19164]_ , \new_[19165]_ , \new_[19169]_ ,
    \new_[19170]_ , \new_[19174]_ , \new_[19175]_ , \new_[19176]_ ,
    \new_[19179]_ , \new_[19183]_ , \new_[19184]_ , \new_[19185]_ ,
    \new_[19189]_ , \new_[19190]_ , \new_[19194]_ , \new_[19195]_ ,
    \new_[19196]_ , \new_[19199]_ , \new_[19203]_ , \new_[19204]_ ,
    \new_[19205]_ , \new_[19209]_ , \new_[19210]_ , \new_[19214]_ ,
    \new_[19215]_ , \new_[19216]_ , \new_[19219]_ , \new_[19223]_ ,
    \new_[19224]_ , \new_[19225]_ , \new_[19229]_ , \new_[19230]_ ,
    \new_[19234]_ , \new_[19235]_ , \new_[19236]_ , \new_[19239]_ ,
    \new_[19243]_ , \new_[19244]_ , \new_[19245]_ , \new_[19249]_ ,
    \new_[19250]_ , \new_[19254]_ , \new_[19255]_ , \new_[19256]_ ,
    \new_[19259]_ , \new_[19263]_ , \new_[19264]_ , \new_[19265]_ ,
    \new_[19269]_ , \new_[19270]_ , \new_[19274]_ , \new_[19275]_ ,
    \new_[19276]_ , \new_[19279]_ , \new_[19283]_ , \new_[19284]_ ,
    \new_[19285]_ , \new_[19289]_ , \new_[19290]_ , \new_[19294]_ ,
    \new_[19295]_ , \new_[19296]_ , \new_[19299]_ , \new_[19303]_ ,
    \new_[19304]_ , \new_[19305]_ , \new_[19309]_ , \new_[19310]_ ,
    \new_[19314]_ , \new_[19315]_ , \new_[19316]_ , \new_[19319]_ ,
    \new_[19323]_ , \new_[19324]_ , \new_[19325]_ , \new_[19329]_ ,
    \new_[19330]_ , \new_[19334]_ , \new_[19335]_ , \new_[19336]_ ,
    \new_[19339]_ , \new_[19343]_ , \new_[19344]_ , \new_[19345]_ ,
    \new_[19349]_ , \new_[19350]_ , \new_[19354]_ , \new_[19355]_ ,
    \new_[19356]_ , \new_[19359]_ , \new_[19363]_ , \new_[19364]_ ,
    \new_[19365]_ , \new_[19369]_ , \new_[19370]_ , \new_[19374]_ ,
    \new_[19375]_ , \new_[19376]_ , \new_[19379]_ , \new_[19383]_ ,
    \new_[19384]_ , \new_[19385]_ , \new_[19389]_ , \new_[19390]_ ,
    \new_[19394]_ , \new_[19395]_ , \new_[19396]_ , \new_[19399]_ ,
    \new_[19403]_ , \new_[19404]_ , \new_[19405]_ , \new_[19409]_ ,
    \new_[19410]_ , \new_[19414]_ , \new_[19415]_ , \new_[19416]_ ,
    \new_[19419]_ , \new_[19423]_ , \new_[19424]_ , \new_[19425]_ ,
    \new_[19429]_ , \new_[19430]_ , \new_[19434]_ , \new_[19435]_ ,
    \new_[19436]_ , \new_[19439]_ , \new_[19443]_ , \new_[19444]_ ,
    \new_[19445]_ , \new_[19449]_ , \new_[19450]_ , \new_[19454]_ ,
    \new_[19455]_ , \new_[19456]_ , \new_[19459]_ , \new_[19463]_ ,
    \new_[19464]_ , \new_[19465]_ , \new_[19469]_ , \new_[19470]_ ,
    \new_[19474]_ , \new_[19475]_ , \new_[19476]_ , \new_[19479]_ ,
    \new_[19483]_ , \new_[19484]_ , \new_[19485]_ , \new_[19489]_ ,
    \new_[19490]_ , \new_[19494]_ , \new_[19495]_ , \new_[19496]_ ,
    \new_[19499]_ , \new_[19503]_ , \new_[19504]_ , \new_[19505]_ ,
    \new_[19509]_ , \new_[19510]_ , \new_[19514]_ , \new_[19515]_ ,
    \new_[19516]_ , \new_[19519]_ , \new_[19523]_ , \new_[19524]_ ,
    \new_[19525]_ , \new_[19529]_ , \new_[19530]_ , \new_[19534]_ ,
    \new_[19535]_ , \new_[19536]_ , \new_[19539]_ , \new_[19543]_ ,
    \new_[19544]_ , \new_[19545]_ , \new_[19549]_ , \new_[19550]_ ,
    \new_[19554]_ , \new_[19555]_ , \new_[19556]_ , \new_[19559]_ ,
    \new_[19563]_ , \new_[19564]_ , \new_[19565]_ , \new_[19569]_ ,
    \new_[19570]_ , \new_[19574]_ , \new_[19575]_ , \new_[19576]_ ,
    \new_[19579]_ , \new_[19583]_ , \new_[19584]_ , \new_[19585]_ ,
    \new_[19589]_ , \new_[19590]_ , \new_[19594]_ , \new_[19595]_ ,
    \new_[19596]_ , \new_[19599]_ , \new_[19603]_ , \new_[19604]_ ,
    \new_[19605]_ , \new_[19609]_ , \new_[19610]_ , \new_[19614]_ ,
    \new_[19615]_ , \new_[19616]_ , \new_[19619]_ , \new_[19623]_ ,
    \new_[19624]_ , \new_[19625]_ , \new_[19629]_ , \new_[19630]_ ,
    \new_[19634]_ , \new_[19635]_ , \new_[19636]_ , \new_[19639]_ ,
    \new_[19643]_ , \new_[19644]_ , \new_[19645]_ , \new_[19649]_ ,
    \new_[19650]_ , \new_[19654]_ , \new_[19655]_ , \new_[19656]_ ,
    \new_[19659]_ , \new_[19663]_ , \new_[19664]_ , \new_[19665]_ ,
    \new_[19669]_ , \new_[19670]_ , \new_[19674]_ , \new_[19675]_ ,
    \new_[19676]_ , \new_[19679]_ , \new_[19683]_ , \new_[19684]_ ,
    \new_[19685]_ , \new_[19689]_ , \new_[19690]_ , \new_[19694]_ ,
    \new_[19695]_ , \new_[19696]_ , \new_[19699]_ , \new_[19703]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19709]_ , \new_[19710]_ ,
    \new_[19714]_ , \new_[19715]_ , \new_[19716]_ , \new_[19719]_ ,
    \new_[19723]_ , \new_[19724]_ , \new_[19725]_ , \new_[19729]_ ,
    \new_[19730]_ , \new_[19734]_ , \new_[19735]_ , \new_[19736]_ ,
    \new_[19739]_ , \new_[19743]_ , \new_[19744]_ , \new_[19745]_ ,
    \new_[19749]_ , \new_[19750]_ , \new_[19754]_ , \new_[19755]_ ,
    \new_[19756]_ , \new_[19759]_ , \new_[19763]_ , \new_[19764]_ ,
    \new_[19765]_ , \new_[19769]_ , \new_[19770]_ , \new_[19774]_ ,
    \new_[19775]_ , \new_[19776]_ , \new_[19779]_ , \new_[19783]_ ,
    \new_[19784]_ , \new_[19785]_ , \new_[19789]_ , \new_[19790]_ ,
    \new_[19794]_ , \new_[19795]_ , \new_[19796]_ , \new_[19799]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19805]_ , \new_[19809]_ ,
    \new_[19810]_ , \new_[19814]_ , \new_[19815]_ , \new_[19816]_ ,
    \new_[19819]_ , \new_[19823]_ , \new_[19824]_ , \new_[19825]_ ,
    \new_[19829]_ , \new_[19830]_ , \new_[19834]_ , \new_[19835]_ ,
    \new_[19836]_ , \new_[19839]_ , \new_[19843]_ , \new_[19844]_ ,
    \new_[19845]_ , \new_[19849]_ , \new_[19850]_ , \new_[19854]_ ,
    \new_[19855]_ , \new_[19856]_ , \new_[19859]_ , \new_[19863]_ ,
    \new_[19864]_ , \new_[19865]_ , \new_[19869]_ , \new_[19870]_ ,
    \new_[19874]_ , \new_[19875]_ , \new_[19876]_ , \new_[19879]_ ,
    \new_[19883]_ , \new_[19884]_ , \new_[19885]_ , \new_[19889]_ ,
    \new_[19890]_ , \new_[19894]_ , \new_[19895]_ , \new_[19896]_ ,
    \new_[19899]_ , \new_[19903]_ , \new_[19904]_ , \new_[19905]_ ,
    \new_[19909]_ , \new_[19910]_ , \new_[19914]_ , \new_[19915]_ ,
    \new_[19916]_ , \new_[19919]_ , \new_[19923]_ , \new_[19924]_ ,
    \new_[19925]_ , \new_[19929]_ , \new_[19930]_ , \new_[19934]_ ,
    \new_[19935]_ , \new_[19936]_ , \new_[19939]_ , \new_[19943]_ ,
    \new_[19944]_ , \new_[19945]_ , \new_[19949]_ , \new_[19950]_ ,
    \new_[19954]_ , \new_[19955]_ , \new_[19956]_ , \new_[19959]_ ,
    \new_[19963]_ , \new_[19964]_ , \new_[19965]_ , \new_[19969]_ ,
    \new_[19970]_ , \new_[19974]_ , \new_[19975]_ , \new_[19976]_ ,
    \new_[19979]_ , \new_[19983]_ , \new_[19984]_ , \new_[19985]_ ,
    \new_[19989]_ , \new_[19990]_ , \new_[19994]_ , \new_[19995]_ ,
    \new_[19996]_ , \new_[19999]_ , \new_[20003]_ , \new_[20004]_ ,
    \new_[20005]_ , \new_[20009]_ , \new_[20010]_ , \new_[20014]_ ,
    \new_[20015]_ , \new_[20016]_ , \new_[20019]_ , \new_[20023]_ ,
    \new_[20024]_ , \new_[20025]_ , \new_[20029]_ , \new_[20030]_ ,
    \new_[20034]_ , \new_[20035]_ , \new_[20036]_ , \new_[20039]_ ,
    \new_[20043]_ , \new_[20044]_ , \new_[20045]_ , \new_[20049]_ ,
    \new_[20050]_ , \new_[20054]_ , \new_[20055]_ , \new_[20056]_ ,
    \new_[20059]_ , \new_[20063]_ , \new_[20064]_ , \new_[20065]_ ,
    \new_[20069]_ , \new_[20070]_ , \new_[20074]_ , \new_[20075]_ ,
    \new_[20076]_ , \new_[20079]_ , \new_[20083]_ , \new_[20084]_ ,
    \new_[20085]_ , \new_[20089]_ , \new_[20090]_ , \new_[20094]_ ,
    \new_[20095]_ , \new_[20096]_ , \new_[20099]_ , \new_[20103]_ ,
    \new_[20104]_ , \new_[20105]_ , \new_[20109]_ , \new_[20110]_ ,
    \new_[20114]_ , \new_[20115]_ , \new_[20116]_ , \new_[20119]_ ,
    \new_[20123]_ , \new_[20124]_ , \new_[20125]_ , \new_[20129]_ ,
    \new_[20130]_ , \new_[20134]_ , \new_[20135]_ , \new_[20136]_ ,
    \new_[20139]_ , \new_[20143]_ , \new_[20144]_ , \new_[20145]_ ,
    \new_[20149]_ , \new_[20150]_ , \new_[20154]_ , \new_[20155]_ ,
    \new_[20156]_ , \new_[20159]_ , \new_[20163]_ , \new_[20164]_ ,
    \new_[20165]_ , \new_[20169]_ , \new_[20170]_ , \new_[20174]_ ,
    \new_[20175]_ , \new_[20176]_ , \new_[20179]_ , \new_[20183]_ ,
    \new_[20184]_ , \new_[20185]_ , \new_[20189]_ , \new_[20190]_ ,
    \new_[20194]_ , \new_[20195]_ , \new_[20196]_ , \new_[20199]_ ,
    \new_[20203]_ , \new_[20204]_ , \new_[20205]_ , \new_[20209]_ ,
    \new_[20210]_ , \new_[20214]_ , \new_[20215]_ , \new_[20216]_ ,
    \new_[20219]_ , \new_[20223]_ , \new_[20224]_ , \new_[20225]_ ,
    \new_[20229]_ , \new_[20230]_ , \new_[20234]_ , \new_[20235]_ ,
    \new_[20236]_ , \new_[20239]_ , \new_[20243]_ , \new_[20244]_ ,
    \new_[20245]_ , \new_[20249]_ , \new_[20250]_ , \new_[20254]_ ,
    \new_[20255]_ , \new_[20256]_ , \new_[20259]_ , \new_[20263]_ ,
    \new_[20264]_ , \new_[20265]_ , \new_[20269]_ , \new_[20270]_ ,
    \new_[20274]_ , \new_[20275]_ , \new_[20276]_ , \new_[20279]_ ,
    \new_[20283]_ , \new_[20284]_ , \new_[20285]_ , \new_[20289]_ ,
    \new_[20290]_ , \new_[20294]_ , \new_[20295]_ , \new_[20296]_ ,
    \new_[20299]_ , \new_[20303]_ , \new_[20304]_ , \new_[20305]_ ,
    \new_[20309]_ , \new_[20310]_ , \new_[20314]_ , \new_[20315]_ ,
    \new_[20316]_ , \new_[20319]_ , \new_[20323]_ , \new_[20324]_ ,
    \new_[20325]_ , \new_[20329]_ , \new_[20330]_ , \new_[20334]_ ,
    \new_[20335]_ , \new_[20336]_ , \new_[20339]_ , \new_[20343]_ ,
    \new_[20344]_ , \new_[20345]_ , \new_[20349]_ , \new_[20350]_ ,
    \new_[20354]_ , \new_[20355]_ , \new_[20356]_ , \new_[20359]_ ,
    \new_[20363]_ , \new_[20364]_ , \new_[20365]_ , \new_[20369]_ ,
    \new_[20370]_ , \new_[20374]_ , \new_[20375]_ , \new_[20376]_ ,
    \new_[20379]_ , \new_[20383]_ , \new_[20384]_ , \new_[20385]_ ,
    \new_[20389]_ , \new_[20390]_ , \new_[20394]_ , \new_[20395]_ ,
    \new_[20396]_ , \new_[20399]_ , \new_[20403]_ , \new_[20404]_ ,
    \new_[20405]_ , \new_[20409]_ , \new_[20410]_ , \new_[20414]_ ,
    \new_[20415]_ , \new_[20416]_ , \new_[20419]_ , \new_[20423]_ ,
    \new_[20424]_ , \new_[20425]_ , \new_[20429]_ , \new_[20430]_ ,
    \new_[20434]_ , \new_[20435]_ , \new_[20436]_ , \new_[20439]_ ,
    \new_[20443]_ , \new_[20444]_ , \new_[20445]_ , \new_[20449]_ ,
    \new_[20450]_ , \new_[20454]_ , \new_[20455]_ , \new_[20456]_ ,
    \new_[20459]_ , \new_[20463]_ , \new_[20464]_ , \new_[20465]_ ,
    \new_[20469]_ , \new_[20470]_ , \new_[20474]_ , \new_[20475]_ ,
    \new_[20476]_ , \new_[20479]_ , \new_[20483]_ , \new_[20484]_ ,
    \new_[20485]_ , \new_[20489]_ , \new_[20490]_ , \new_[20494]_ ,
    \new_[20495]_ , \new_[20496]_ , \new_[20499]_ , \new_[20503]_ ,
    \new_[20504]_ , \new_[20505]_ , \new_[20509]_ , \new_[20510]_ ,
    \new_[20514]_ , \new_[20515]_ , \new_[20516]_ , \new_[20519]_ ,
    \new_[20523]_ , \new_[20524]_ , \new_[20525]_ , \new_[20529]_ ,
    \new_[20530]_ , \new_[20534]_ , \new_[20535]_ , \new_[20536]_ ,
    \new_[20539]_ , \new_[20543]_ , \new_[20544]_ , \new_[20545]_ ,
    \new_[20549]_ , \new_[20550]_ , \new_[20554]_ , \new_[20555]_ ,
    \new_[20556]_ , \new_[20559]_ , \new_[20563]_ , \new_[20564]_ ,
    \new_[20565]_ , \new_[20569]_ , \new_[20570]_ , \new_[20574]_ ,
    \new_[20575]_ , \new_[20576]_ , \new_[20579]_ , \new_[20583]_ ,
    \new_[20584]_ , \new_[20585]_ , \new_[20589]_ , \new_[20590]_ ,
    \new_[20594]_ , \new_[20595]_ , \new_[20596]_ , \new_[20599]_ ,
    \new_[20603]_ , \new_[20604]_ , \new_[20605]_ , \new_[20609]_ ,
    \new_[20610]_ , \new_[20614]_ , \new_[20615]_ , \new_[20616]_ ,
    \new_[20619]_ , \new_[20623]_ , \new_[20624]_ , \new_[20625]_ ,
    \new_[20629]_ , \new_[20630]_ , \new_[20634]_ , \new_[20635]_ ,
    \new_[20636]_ , \new_[20639]_ , \new_[20643]_ , \new_[20644]_ ,
    \new_[20645]_ , \new_[20649]_ , \new_[20650]_ , \new_[20654]_ ,
    \new_[20655]_ , \new_[20656]_ , \new_[20659]_ , \new_[20663]_ ,
    \new_[20664]_ , \new_[20665]_ , \new_[20669]_ , \new_[20670]_ ,
    \new_[20674]_ , \new_[20675]_ , \new_[20676]_ , \new_[20679]_ ,
    \new_[20683]_ , \new_[20684]_ , \new_[20685]_ , \new_[20689]_ ,
    \new_[20690]_ , \new_[20694]_ , \new_[20695]_ , \new_[20696]_ ,
    \new_[20699]_ , \new_[20703]_ , \new_[20704]_ , \new_[20705]_ ,
    \new_[20709]_ , \new_[20710]_ , \new_[20714]_ , \new_[20715]_ ,
    \new_[20716]_ , \new_[20719]_ , \new_[20723]_ , \new_[20724]_ ,
    \new_[20725]_ , \new_[20729]_ , \new_[20730]_ , \new_[20734]_ ,
    \new_[20735]_ , \new_[20736]_ , \new_[20739]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20745]_ , \new_[20749]_ , \new_[20750]_ ,
    \new_[20754]_ , \new_[20755]_ , \new_[20756]_ , \new_[20759]_ ,
    \new_[20763]_ , \new_[20764]_ , \new_[20765]_ , \new_[20769]_ ,
    \new_[20770]_ , \new_[20774]_ , \new_[20775]_ , \new_[20776]_ ,
    \new_[20779]_ , \new_[20783]_ , \new_[20784]_ , \new_[20785]_ ,
    \new_[20789]_ , \new_[20790]_ , \new_[20794]_ , \new_[20795]_ ,
    \new_[20796]_ , \new_[20799]_ , \new_[20803]_ , \new_[20804]_ ,
    \new_[20805]_ , \new_[20809]_ , \new_[20810]_ , \new_[20814]_ ,
    \new_[20815]_ , \new_[20816]_ , \new_[20819]_ , \new_[20823]_ ,
    \new_[20824]_ , \new_[20825]_ , \new_[20829]_ , \new_[20830]_ ,
    \new_[20834]_ , \new_[20835]_ , \new_[20836]_ , \new_[20839]_ ,
    \new_[20843]_ , \new_[20844]_ , \new_[20845]_ , \new_[20849]_ ,
    \new_[20850]_ , \new_[20854]_ , \new_[20855]_ , \new_[20856]_ ,
    \new_[20859]_ , \new_[20863]_ , \new_[20864]_ , \new_[20865]_ ,
    \new_[20869]_ , \new_[20870]_ , \new_[20874]_ , \new_[20875]_ ,
    \new_[20876]_ , \new_[20879]_ , \new_[20883]_ , \new_[20884]_ ,
    \new_[20885]_ , \new_[20889]_ , \new_[20890]_ , \new_[20894]_ ,
    \new_[20895]_ , \new_[20896]_ , \new_[20899]_ , \new_[20903]_ ,
    \new_[20904]_ , \new_[20905]_ , \new_[20909]_ , \new_[20910]_ ,
    \new_[20914]_ , \new_[20915]_ , \new_[20916]_ , \new_[20919]_ ,
    \new_[20923]_ , \new_[20924]_ , \new_[20925]_ , \new_[20929]_ ,
    \new_[20930]_ , \new_[20934]_ , \new_[20935]_ , \new_[20936]_ ,
    \new_[20939]_ , \new_[20943]_ , \new_[20944]_ , \new_[20945]_ ,
    \new_[20949]_ , \new_[20950]_ , \new_[20954]_ , \new_[20955]_ ,
    \new_[20956]_ , \new_[20959]_ , \new_[20963]_ , \new_[20964]_ ,
    \new_[20965]_ , \new_[20969]_ , \new_[20970]_ , \new_[20974]_ ,
    \new_[20975]_ , \new_[20976]_ , \new_[20979]_ , \new_[20983]_ ,
    \new_[20984]_ , \new_[20985]_ , \new_[20989]_ , \new_[20990]_ ,
    \new_[20994]_ , \new_[20995]_ , \new_[20996]_ , \new_[20999]_ ,
    \new_[21003]_ , \new_[21004]_ , \new_[21005]_ , \new_[21009]_ ,
    \new_[21010]_ , \new_[21014]_ , \new_[21015]_ , \new_[21016]_ ,
    \new_[21019]_ , \new_[21023]_ , \new_[21024]_ , \new_[21025]_ ,
    \new_[21029]_ , \new_[21030]_ , \new_[21034]_ , \new_[21035]_ ,
    \new_[21036]_ , \new_[21039]_ , \new_[21043]_ , \new_[21044]_ ,
    \new_[21045]_ , \new_[21049]_ , \new_[21050]_ , \new_[21054]_ ,
    \new_[21055]_ , \new_[21056]_ , \new_[21059]_ , \new_[21063]_ ,
    \new_[21064]_ , \new_[21065]_ , \new_[21069]_ , \new_[21070]_ ,
    \new_[21074]_ , \new_[21075]_ , \new_[21076]_ , \new_[21079]_ ,
    \new_[21083]_ , \new_[21084]_ , \new_[21085]_ , \new_[21089]_ ,
    \new_[21090]_ , \new_[21094]_ , \new_[21095]_ , \new_[21096]_ ,
    \new_[21099]_ , \new_[21103]_ , \new_[21104]_ , \new_[21105]_ ,
    \new_[21109]_ , \new_[21110]_ , \new_[21114]_ , \new_[21115]_ ,
    \new_[21116]_ , \new_[21119]_ , \new_[21123]_ , \new_[21124]_ ,
    \new_[21125]_ , \new_[21129]_ , \new_[21130]_ , \new_[21134]_ ,
    \new_[21135]_ , \new_[21136]_ , \new_[21139]_ , \new_[21143]_ ,
    \new_[21144]_ , \new_[21145]_ , \new_[21149]_ , \new_[21150]_ ,
    \new_[21154]_ , \new_[21155]_ , \new_[21156]_ , \new_[21159]_ ,
    \new_[21163]_ , \new_[21164]_ , \new_[21165]_ , \new_[21169]_ ,
    \new_[21170]_ , \new_[21174]_ , \new_[21175]_ , \new_[21176]_ ,
    \new_[21179]_ , \new_[21183]_ , \new_[21184]_ , \new_[21185]_ ,
    \new_[21189]_ , \new_[21190]_ , \new_[21194]_ , \new_[21195]_ ,
    \new_[21196]_ , \new_[21199]_ , \new_[21203]_ , \new_[21204]_ ,
    \new_[21205]_ , \new_[21209]_ , \new_[21210]_ , \new_[21214]_ ,
    \new_[21215]_ , \new_[21216]_ , \new_[21219]_ , \new_[21223]_ ,
    \new_[21224]_ , \new_[21225]_ , \new_[21229]_ , \new_[21230]_ ,
    \new_[21234]_ , \new_[21235]_ , \new_[21236]_ , \new_[21239]_ ,
    \new_[21243]_ , \new_[21244]_ , \new_[21245]_ , \new_[21249]_ ,
    \new_[21250]_ , \new_[21254]_ , \new_[21255]_ , \new_[21256]_ ,
    \new_[21259]_ , \new_[21263]_ , \new_[21264]_ , \new_[21265]_ ,
    \new_[21269]_ , \new_[21270]_ , \new_[21274]_ , \new_[21275]_ ,
    \new_[21276]_ , \new_[21279]_ , \new_[21283]_ , \new_[21284]_ ,
    \new_[21285]_ , \new_[21289]_ , \new_[21290]_ , \new_[21294]_ ,
    \new_[21295]_ , \new_[21296]_ , \new_[21299]_ , \new_[21303]_ ,
    \new_[21304]_ , \new_[21305]_ , \new_[21309]_ , \new_[21310]_ ,
    \new_[21314]_ , \new_[21315]_ , \new_[21316]_ , \new_[21319]_ ,
    \new_[21323]_ , \new_[21324]_ , \new_[21325]_ , \new_[21329]_ ,
    \new_[21330]_ , \new_[21334]_ , \new_[21335]_ , \new_[21336]_ ,
    \new_[21339]_ , \new_[21343]_ , \new_[21344]_ , \new_[21345]_ ,
    \new_[21349]_ , \new_[21350]_ , \new_[21354]_ , \new_[21355]_ ,
    \new_[21356]_ , \new_[21359]_ , \new_[21363]_ , \new_[21364]_ ,
    \new_[21365]_ , \new_[21369]_ , \new_[21370]_ , \new_[21374]_ ,
    \new_[21375]_ , \new_[21376]_ , \new_[21379]_ , \new_[21383]_ ,
    \new_[21384]_ , \new_[21385]_ , \new_[21389]_ , \new_[21390]_ ,
    \new_[21394]_ , \new_[21395]_ , \new_[21396]_ , \new_[21399]_ ,
    \new_[21403]_ , \new_[21404]_ , \new_[21405]_ , \new_[21409]_ ,
    \new_[21410]_ , \new_[21414]_ , \new_[21415]_ , \new_[21416]_ ,
    \new_[21419]_ , \new_[21423]_ , \new_[21424]_ , \new_[21425]_ ,
    \new_[21429]_ , \new_[21430]_ , \new_[21434]_ , \new_[21435]_ ,
    \new_[21436]_ , \new_[21439]_ , \new_[21443]_ , \new_[21444]_ ,
    \new_[21445]_ , \new_[21449]_ , \new_[21450]_ , \new_[21454]_ ,
    \new_[21455]_ , \new_[21456]_ , \new_[21459]_ , \new_[21463]_ ,
    \new_[21464]_ , \new_[21465]_ , \new_[21469]_ , \new_[21470]_ ,
    \new_[21474]_ , \new_[21475]_ , \new_[21476]_ , \new_[21479]_ ,
    \new_[21483]_ , \new_[21484]_ , \new_[21485]_ , \new_[21489]_ ,
    \new_[21490]_ , \new_[21494]_ , \new_[21495]_ , \new_[21496]_ ,
    \new_[21499]_ , \new_[21503]_ , \new_[21504]_ , \new_[21505]_ ,
    \new_[21509]_ , \new_[21510]_ , \new_[21514]_ , \new_[21515]_ ,
    \new_[21516]_ , \new_[21519]_ , \new_[21523]_ , \new_[21524]_ ,
    \new_[21525]_ , \new_[21529]_ , \new_[21530]_ , \new_[21534]_ ,
    \new_[21535]_ , \new_[21536]_ , \new_[21539]_ , \new_[21543]_ ,
    \new_[21544]_ , \new_[21545]_ , \new_[21549]_ , \new_[21550]_ ,
    \new_[21554]_ , \new_[21555]_ , \new_[21556]_ , \new_[21559]_ ,
    \new_[21563]_ , \new_[21564]_ , \new_[21565]_ , \new_[21569]_ ,
    \new_[21570]_ , \new_[21574]_ , \new_[21575]_ , \new_[21576]_ ,
    \new_[21579]_ , \new_[21583]_ , \new_[21584]_ , \new_[21585]_ ,
    \new_[21589]_ , \new_[21590]_ , \new_[21594]_ , \new_[21595]_ ,
    \new_[21596]_ , \new_[21599]_ , \new_[21603]_ , \new_[21604]_ ,
    \new_[21605]_ , \new_[21609]_ , \new_[21610]_ , \new_[21614]_ ,
    \new_[21615]_ , \new_[21616]_ , \new_[21619]_ , \new_[21623]_ ,
    \new_[21624]_ , \new_[21625]_ , \new_[21629]_ , \new_[21630]_ ,
    \new_[21634]_ , \new_[21635]_ , \new_[21636]_ , \new_[21639]_ ,
    \new_[21643]_ , \new_[21644]_ , \new_[21645]_ , \new_[21649]_ ,
    \new_[21650]_ , \new_[21654]_ , \new_[21655]_ , \new_[21656]_ ,
    \new_[21659]_ , \new_[21663]_ , \new_[21664]_ , \new_[21665]_ ,
    \new_[21669]_ , \new_[21670]_ , \new_[21674]_ , \new_[21675]_ ,
    \new_[21676]_ , \new_[21679]_ , \new_[21683]_ , \new_[21684]_ ,
    \new_[21685]_ , \new_[21689]_ , \new_[21690]_ , \new_[21694]_ ,
    \new_[21695]_ , \new_[21696]_ , \new_[21699]_ , \new_[21703]_ ,
    \new_[21704]_ , \new_[21705]_ , \new_[21709]_ , \new_[21710]_ ,
    \new_[21714]_ , \new_[21715]_ , \new_[21716]_ , \new_[21719]_ ,
    \new_[21723]_ , \new_[21724]_ , \new_[21725]_ , \new_[21729]_ ,
    \new_[21730]_ , \new_[21734]_ , \new_[21735]_ , \new_[21736]_ ,
    \new_[21739]_ , \new_[21743]_ , \new_[21744]_ , \new_[21745]_ ,
    \new_[21749]_ , \new_[21750]_ , \new_[21754]_ , \new_[21755]_ ,
    \new_[21756]_ , \new_[21759]_ , \new_[21763]_ , \new_[21764]_ ,
    \new_[21765]_ , \new_[21769]_ , \new_[21770]_ , \new_[21774]_ ,
    \new_[21775]_ , \new_[21776]_ , \new_[21779]_ , \new_[21783]_ ,
    \new_[21784]_ , \new_[21785]_ , \new_[21789]_ , \new_[21790]_ ,
    \new_[21794]_ , \new_[21795]_ , \new_[21796]_ , \new_[21799]_ ,
    \new_[21803]_ , \new_[21804]_ , \new_[21805]_ , \new_[21809]_ ,
    \new_[21810]_ , \new_[21814]_ , \new_[21815]_ , \new_[21816]_ ,
    \new_[21819]_ , \new_[21823]_ , \new_[21824]_ , \new_[21825]_ ,
    \new_[21829]_ , \new_[21830]_ , \new_[21834]_ , \new_[21835]_ ,
    \new_[21836]_ , \new_[21839]_ , \new_[21843]_ , \new_[21844]_ ,
    \new_[21845]_ , \new_[21849]_ , \new_[21850]_ , \new_[21854]_ ,
    \new_[21855]_ , \new_[21856]_ , \new_[21859]_ , \new_[21863]_ ,
    \new_[21864]_ , \new_[21865]_ , \new_[21869]_ , \new_[21870]_ ,
    \new_[21874]_ , \new_[21875]_ , \new_[21876]_ , \new_[21879]_ ,
    \new_[21883]_ , \new_[21884]_ , \new_[21885]_ , \new_[21889]_ ,
    \new_[21890]_ , \new_[21894]_ , \new_[21895]_ , \new_[21896]_ ,
    \new_[21899]_ , \new_[21903]_ , \new_[21904]_ , \new_[21905]_ ,
    \new_[21909]_ , \new_[21910]_ , \new_[21914]_ , \new_[21915]_ ,
    \new_[21916]_ , \new_[21919]_ , \new_[21923]_ , \new_[21924]_ ,
    \new_[21925]_ , \new_[21929]_ , \new_[21930]_ , \new_[21934]_ ,
    \new_[21935]_ , \new_[21936]_ , \new_[21939]_ , \new_[21943]_ ,
    \new_[21944]_ , \new_[21945]_ , \new_[21949]_ , \new_[21950]_ ,
    \new_[21954]_ , \new_[21955]_ , \new_[21956]_ , \new_[21959]_ ,
    \new_[21963]_ , \new_[21964]_ , \new_[21965]_ , \new_[21969]_ ,
    \new_[21970]_ , \new_[21974]_ , \new_[21975]_ , \new_[21976]_ ,
    \new_[21979]_ , \new_[21983]_ , \new_[21984]_ , \new_[21985]_ ,
    \new_[21989]_ , \new_[21990]_ , \new_[21994]_ , \new_[21995]_ ,
    \new_[21996]_ , \new_[21999]_ , \new_[22003]_ , \new_[22004]_ ,
    \new_[22005]_ , \new_[22009]_ , \new_[22010]_ , \new_[22014]_ ,
    \new_[22015]_ , \new_[22016]_ , \new_[22019]_ , \new_[22023]_ ,
    \new_[22024]_ , \new_[22025]_ , \new_[22029]_ , \new_[22030]_ ,
    \new_[22034]_ , \new_[22035]_ , \new_[22036]_ , \new_[22039]_ ,
    \new_[22043]_ , \new_[22044]_ , \new_[22045]_ , \new_[22049]_ ,
    \new_[22050]_ , \new_[22054]_ , \new_[22055]_ , \new_[22056]_ ,
    \new_[22059]_ , \new_[22063]_ , \new_[22064]_ , \new_[22065]_ ,
    \new_[22069]_ , \new_[22070]_ , \new_[22074]_ , \new_[22075]_ ,
    \new_[22076]_ , \new_[22079]_ , \new_[22083]_ , \new_[22084]_ ,
    \new_[22085]_ , \new_[22089]_ , \new_[22090]_ , \new_[22094]_ ,
    \new_[22095]_ , \new_[22096]_ , \new_[22099]_ , \new_[22103]_ ,
    \new_[22104]_ , \new_[22105]_ , \new_[22109]_ , \new_[22110]_ ,
    \new_[22114]_ , \new_[22115]_ , \new_[22116]_ , \new_[22119]_ ,
    \new_[22123]_ , \new_[22124]_ , \new_[22125]_ , \new_[22129]_ ,
    \new_[22130]_ , \new_[22134]_ , \new_[22135]_ , \new_[22136]_ ,
    \new_[22139]_ , \new_[22143]_ , \new_[22144]_ , \new_[22145]_ ,
    \new_[22149]_ , \new_[22150]_ , \new_[22154]_ , \new_[22155]_ ,
    \new_[22156]_ , \new_[22159]_ , \new_[22163]_ , \new_[22164]_ ,
    \new_[22165]_ , \new_[22169]_ , \new_[22170]_ , \new_[22174]_ ,
    \new_[22175]_ , \new_[22176]_ , \new_[22179]_ , \new_[22183]_ ,
    \new_[22184]_ , \new_[22185]_ , \new_[22189]_ , \new_[22190]_ ,
    \new_[22194]_ , \new_[22195]_ , \new_[22196]_ , \new_[22199]_ ,
    \new_[22203]_ , \new_[22204]_ , \new_[22205]_ , \new_[22209]_ ,
    \new_[22210]_ , \new_[22214]_ , \new_[22215]_ , \new_[22216]_ ,
    \new_[22219]_ , \new_[22223]_ , \new_[22224]_ , \new_[22225]_ ,
    \new_[22229]_ , \new_[22230]_ , \new_[22234]_ , \new_[22235]_ ,
    \new_[22236]_ , \new_[22239]_ , \new_[22243]_ , \new_[22244]_ ,
    \new_[22245]_ , \new_[22249]_ , \new_[22250]_ , \new_[22254]_ ,
    \new_[22255]_ , \new_[22256]_ , \new_[22259]_ , \new_[22263]_ ,
    \new_[22264]_ , \new_[22265]_ , \new_[22269]_ , \new_[22270]_ ,
    \new_[22274]_ , \new_[22275]_ , \new_[22276]_ , \new_[22279]_ ,
    \new_[22283]_ , \new_[22284]_ , \new_[22285]_ , \new_[22289]_ ,
    \new_[22290]_ , \new_[22294]_ , \new_[22295]_ , \new_[22296]_ ,
    \new_[22299]_ , \new_[22303]_ , \new_[22304]_ , \new_[22305]_ ,
    \new_[22309]_ , \new_[22310]_ , \new_[22314]_ , \new_[22315]_ ,
    \new_[22316]_ , \new_[22319]_ , \new_[22323]_ , \new_[22324]_ ,
    \new_[22325]_ , \new_[22329]_ , \new_[22330]_ , \new_[22334]_ ,
    \new_[22335]_ , \new_[22336]_ , \new_[22339]_ , \new_[22343]_ ,
    \new_[22344]_ , \new_[22345]_ , \new_[22349]_ , \new_[22350]_ ,
    \new_[22354]_ , \new_[22355]_ , \new_[22356]_ , \new_[22359]_ ,
    \new_[22363]_ , \new_[22364]_ , \new_[22365]_ , \new_[22369]_ ,
    \new_[22370]_ , \new_[22374]_ , \new_[22375]_ , \new_[22376]_ ,
    \new_[22379]_ , \new_[22383]_ , \new_[22384]_ , \new_[22385]_ ,
    \new_[22389]_ , \new_[22390]_ , \new_[22394]_ , \new_[22395]_ ,
    \new_[22396]_ , \new_[22399]_ , \new_[22403]_ , \new_[22404]_ ,
    \new_[22405]_ , \new_[22409]_ , \new_[22410]_ , \new_[22414]_ ,
    \new_[22415]_ , \new_[22416]_ , \new_[22419]_ , \new_[22423]_ ,
    \new_[22424]_ , \new_[22425]_ , \new_[22429]_ , \new_[22430]_ ,
    \new_[22434]_ , \new_[22435]_ , \new_[22436]_ , \new_[22439]_ ,
    \new_[22443]_ , \new_[22444]_ , \new_[22445]_ , \new_[22449]_ ,
    \new_[22450]_ , \new_[22454]_ , \new_[22455]_ , \new_[22456]_ ,
    \new_[22459]_ , \new_[22463]_ , \new_[22464]_ , \new_[22465]_ ,
    \new_[22469]_ , \new_[22470]_ , \new_[22474]_ , \new_[22475]_ ,
    \new_[22476]_ , \new_[22479]_ , \new_[22483]_ , \new_[22484]_ ,
    \new_[22485]_ , \new_[22489]_ , \new_[22490]_ , \new_[22494]_ ,
    \new_[22495]_ , \new_[22496]_ , \new_[22499]_ , \new_[22503]_ ,
    \new_[22504]_ , \new_[22505]_ , \new_[22509]_ , \new_[22510]_ ,
    \new_[22514]_ , \new_[22515]_ , \new_[22516]_ , \new_[22519]_ ,
    \new_[22523]_ , \new_[22524]_ , \new_[22525]_ , \new_[22529]_ ,
    \new_[22530]_ , \new_[22534]_ , \new_[22535]_ , \new_[22536]_ ,
    \new_[22539]_ , \new_[22543]_ , \new_[22544]_ , \new_[22545]_ ,
    \new_[22549]_ , \new_[22550]_ , \new_[22554]_ , \new_[22555]_ ,
    \new_[22556]_ , \new_[22559]_ , \new_[22563]_ , \new_[22564]_ ,
    \new_[22565]_ , \new_[22569]_ , \new_[22570]_ , \new_[22574]_ ,
    \new_[22575]_ , \new_[22576]_ , \new_[22579]_ , \new_[22583]_ ,
    \new_[22584]_ , \new_[22585]_ , \new_[22589]_ , \new_[22590]_ ,
    \new_[22594]_ , \new_[22595]_ , \new_[22596]_ , \new_[22599]_ ,
    \new_[22603]_ , \new_[22604]_ , \new_[22605]_ , \new_[22609]_ ,
    \new_[22610]_ , \new_[22614]_ , \new_[22615]_ , \new_[22616]_ ,
    \new_[22619]_ , \new_[22623]_ , \new_[22624]_ , \new_[22625]_ ,
    \new_[22629]_ , \new_[22630]_ , \new_[22634]_ , \new_[22635]_ ,
    \new_[22636]_ , \new_[22639]_ , \new_[22643]_ , \new_[22644]_ ,
    \new_[22645]_ , \new_[22649]_ , \new_[22650]_ , \new_[22654]_ ,
    \new_[22655]_ , \new_[22656]_ , \new_[22659]_ , \new_[22663]_ ,
    \new_[22664]_ , \new_[22665]_ , \new_[22669]_ , \new_[22670]_ ,
    \new_[22674]_ , \new_[22675]_ , \new_[22676]_ , \new_[22679]_ ,
    \new_[22683]_ , \new_[22684]_ , \new_[22685]_ , \new_[22689]_ ,
    \new_[22690]_ , \new_[22694]_ , \new_[22695]_ , \new_[22696]_ ,
    \new_[22699]_ , \new_[22703]_ , \new_[22704]_ , \new_[22705]_ ,
    \new_[22709]_ , \new_[22710]_ , \new_[22714]_ , \new_[22715]_ ,
    \new_[22716]_ , \new_[22719]_ , \new_[22723]_ , \new_[22724]_ ,
    \new_[22725]_ , \new_[22729]_ , \new_[22730]_ , \new_[22734]_ ,
    \new_[22735]_ , \new_[22736]_ , \new_[22739]_ , \new_[22743]_ ,
    \new_[22744]_ , \new_[22745]_ , \new_[22749]_ , \new_[22750]_ ,
    \new_[22754]_ , \new_[22755]_ , \new_[22756]_ , \new_[22759]_ ,
    \new_[22763]_ , \new_[22764]_ , \new_[22765]_ , \new_[22769]_ ,
    \new_[22770]_ , \new_[22774]_ , \new_[22775]_ , \new_[22776]_ ,
    \new_[22779]_ , \new_[22783]_ , \new_[22784]_ , \new_[22785]_ ,
    \new_[22789]_ , \new_[22790]_ , \new_[22794]_ , \new_[22795]_ ,
    \new_[22796]_ , \new_[22799]_ , \new_[22803]_ , \new_[22804]_ ,
    \new_[22805]_ , \new_[22809]_ , \new_[22810]_ , \new_[22814]_ ,
    \new_[22815]_ , \new_[22816]_ , \new_[22819]_ , \new_[22823]_ ,
    \new_[22824]_ , \new_[22825]_ , \new_[22829]_ , \new_[22830]_ ,
    \new_[22834]_ , \new_[22835]_ , \new_[22836]_ , \new_[22839]_ ,
    \new_[22843]_ , \new_[22844]_ , \new_[22845]_ , \new_[22849]_ ,
    \new_[22850]_ , \new_[22854]_ , \new_[22855]_ , \new_[22856]_ ,
    \new_[22859]_ , \new_[22863]_ , \new_[22864]_ , \new_[22865]_ ,
    \new_[22869]_ , \new_[22870]_ , \new_[22874]_ , \new_[22875]_ ,
    \new_[22876]_ , \new_[22879]_ , \new_[22883]_ , \new_[22884]_ ,
    \new_[22885]_ , \new_[22889]_ , \new_[22890]_ , \new_[22894]_ ,
    \new_[22895]_ , \new_[22896]_ , \new_[22899]_ , \new_[22903]_ ,
    \new_[22904]_ , \new_[22905]_ , \new_[22909]_ , \new_[22910]_ ,
    \new_[22914]_ , \new_[22915]_ , \new_[22916]_ , \new_[22919]_ ,
    \new_[22923]_ , \new_[22924]_ , \new_[22925]_ , \new_[22929]_ ,
    \new_[22930]_ , \new_[22934]_ , \new_[22935]_ , \new_[22936]_ ,
    \new_[22939]_ , \new_[22943]_ , \new_[22944]_ , \new_[22945]_ ,
    \new_[22949]_ , \new_[22950]_ , \new_[22954]_ , \new_[22955]_ ,
    \new_[22956]_ , \new_[22959]_ , \new_[22963]_ , \new_[22964]_ ,
    \new_[22965]_ , \new_[22969]_ , \new_[22970]_ , \new_[22974]_ ,
    \new_[22975]_ , \new_[22976]_ , \new_[22979]_ , \new_[22983]_ ,
    \new_[22984]_ , \new_[22985]_ , \new_[22989]_ , \new_[22990]_ ,
    \new_[22994]_ , \new_[22995]_ , \new_[22996]_ , \new_[22999]_ ,
    \new_[23003]_ , \new_[23004]_ , \new_[23005]_ , \new_[23009]_ ,
    \new_[23010]_ , \new_[23014]_ , \new_[23015]_ , \new_[23016]_ ,
    \new_[23019]_ , \new_[23023]_ , \new_[23024]_ , \new_[23025]_ ,
    \new_[23029]_ , \new_[23030]_ , \new_[23034]_ , \new_[23035]_ ,
    \new_[23036]_ , \new_[23039]_ , \new_[23043]_ , \new_[23044]_ ,
    \new_[23045]_ , \new_[23049]_ , \new_[23050]_ , \new_[23054]_ ,
    \new_[23055]_ , \new_[23056]_ , \new_[23059]_ , \new_[23063]_ ,
    \new_[23064]_ , \new_[23065]_ , \new_[23069]_ , \new_[23070]_ ,
    \new_[23074]_ , \new_[23075]_ , \new_[23076]_ , \new_[23079]_ ,
    \new_[23083]_ , \new_[23084]_ , \new_[23085]_ , \new_[23089]_ ,
    \new_[23090]_ , \new_[23094]_ , \new_[23095]_ , \new_[23096]_ ,
    \new_[23099]_ , \new_[23103]_ , \new_[23104]_ , \new_[23105]_ ,
    \new_[23109]_ , \new_[23110]_ , \new_[23114]_ , \new_[23115]_ ,
    \new_[23116]_ , \new_[23119]_ , \new_[23123]_ , \new_[23124]_ ,
    \new_[23125]_ , \new_[23129]_ , \new_[23130]_ , \new_[23134]_ ,
    \new_[23135]_ , \new_[23136]_ , \new_[23139]_ , \new_[23143]_ ,
    \new_[23144]_ , \new_[23145]_ , \new_[23149]_ , \new_[23150]_ ,
    \new_[23154]_ , \new_[23155]_ , \new_[23156]_ , \new_[23159]_ ,
    \new_[23163]_ , \new_[23164]_ , \new_[23165]_ , \new_[23169]_ ,
    \new_[23170]_ , \new_[23174]_ , \new_[23175]_ , \new_[23176]_ ,
    \new_[23179]_ , \new_[23183]_ , \new_[23184]_ , \new_[23185]_ ,
    \new_[23189]_ , \new_[23190]_ , \new_[23194]_ , \new_[23195]_ ,
    \new_[23196]_ , \new_[23199]_ , \new_[23203]_ , \new_[23204]_ ,
    \new_[23205]_ , \new_[23209]_ , \new_[23210]_ , \new_[23214]_ ,
    \new_[23215]_ , \new_[23216]_ , \new_[23219]_ , \new_[23223]_ ,
    \new_[23224]_ , \new_[23225]_ , \new_[23229]_ , \new_[23230]_ ,
    \new_[23234]_ , \new_[23235]_ , \new_[23236]_ , \new_[23239]_ ,
    \new_[23243]_ , \new_[23244]_ , \new_[23245]_ , \new_[23249]_ ,
    \new_[23250]_ , \new_[23254]_ , \new_[23255]_ , \new_[23256]_ ,
    \new_[23259]_ , \new_[23263]_ , \new_[23264]_ , \new_[23265]_ ,
    \new_[23269]_ , \new_[23270]_ , \new_[23274]_ , \new_[23275]_ ,
    \new_[23276]_ , \new_[23279]_ , \new_[23283]_ , \new_[23284]_ ,
    \new_[23285]_ , \new_[23289]_ , \new_[23290]_ , \new_[23294]_ ,
    \new_[23295]_ , \new_[23296]_ , \new_[23299]_ , \new_[23303]_ ,
    \new_[23304]_ , \new_[23305]_ , \new_[23309]_ , \new_[23310]_ ,
    \new_[23314]_ , \new_[23315]_ , \new_[23316]_ , \new_[23319]_ ,
    \new_[23323]_ , \new_[23324]_ , \new_[23325]_ , \new_[23329]_ ,
    \new_[23330]_ , \new_[23334]_ , \new_[23335]_ , \new_[23336]_ ,
    \new_[23339]_ , \new_[23343]_ , \new_[23344]_ , \new_[23345]_ ,
    \new_[23349]_ , \new_[23350]_ , \new_[23354]_ , \new_[23355]_ ,
    \new_[23356]_ , \new_[23359]_ , \new_[23363]_ , \new_[23364]_ ,
    \new_[23365]_ , \new_[23369]_ , \new_[23370]_ , \new_[23374]_ ,
    \new_[23375]_ , \new_[23376]_ , \new_[23379]_ , \new_[23383]_ ,
    \new_[23384]_ , \new_[23385]_ , \new_[23389]_ , \new_[23390]_ ,
    \new_[23394]_ , \new_[23395]_ , \new_[23396]_ , \new_[23399]_ ,
    \new_[23403]_ , \new_[23404]_ , \new_[23405]_ , \new_[23409]_ ,
    \new_[23410]_ , \new_[23414]_ , \new_[23415]_ , \new_[23416]_ ,
    \new_[23419]_ , \new_[23423]_ , \new_[23424]_ , \new_[23425]_ ,
    \new_[23429]_ , \new_[23430]_ , \new_[23434]_ , \new_[23435]_ ,
    \new_[23436]_ , \new_[23439]_ , \new_[23443]_ , \new_[23444]_ ,
    \new_[23445]_ , \new_[23449]_ , \new_[23450]_ , \new_[23454]_ ,
    \new_[23455]_ , \new_[23456]_ , \new_[23459]_ , \new_[23463]_ ,
    \new_[23464]_ , \new_[23465]_ , \new_[23469]_ , \new_[23470]_ ,
    \new_[23474]_ , \new_[23475]_ , \new_[23476]_ , \new_[23479]_ ,
    \new_[23483]_ , \new_[23484]_ , \new_[23485]_ , \new_[23489]_ ,
    \new_[23490]_ , \new_[23494]_ , \new_[23495]_ , \new_[23496]_ ,
    \new_[23499]_ , \new_[23503]_ , \new_[23504]_ , \new_[23505]_ ,
    \new_[23509]_ , \new_[23510]_ , \new_[23514]_ , \new_[23515]_ ,
    \new_[23516]_ , \new_[23519]_ , \new_[23523]_ , \new_[23524]_ ,
    \new_[23525]_ , \new_[23529]_ , \new_[23530]_ , \new_[23534]_ ,
    \new_[23535]_ , \new_[23536]_ , \new_[23539]_ , \new_[23543]_ ,
    \new_[23544]_ , \new_[23545]_ , \new_[23549]_ , \new_[23550]_ ,
    \new_[23554]_ , \new_[23555]_ , \new_[23556]_ , \new_[23559]_ ,
    \new_[23563]_ , \new_[23564]_ , \new_[23565]_ , \new_[23569]_ ,
    \new_[23570]_ , \new_[23574]_ , \new_[23575]_ , \new_[23576]_ ,
    \new_[23579]_ , \new_[23583]_ , \new_[23584]_ , \new_[23585]_ ,
    \new_[23589]_ , \new_[23590]_ , \new_[23594]_ , \new_[23595]_ ,
    \new_[23596]_ , \new_[23599]_ , \new_[23603]_ , \new_[23604]_ ,
    \new_[23605]_ , \new_[23609]_ , \new_[23610]_ , \new_[23614]_ ,
    \new_[23615]_ , \new_[23616]_ , \new_[23619]_ , \new_[23623]_ ,
    \new_[23624]_ , \new_[23625]_ , \new_[23629]_ , \new_[23630]_ ,
    \new_[23634]_ , \new_[23635]_ , \new_[23636]_ , \new_[23639]_ ,
    \new_[23643]_ , \new_[23644]_ , \new_[23645]_ , \new_[23649]_ ,
    \new_[23650]_ , \new_[23654]_ , \new_[23655]_ , \new_[23656]_ ,
    \new_[23659]_ , \new_[23663]_ , \new_[23664]_ , \new_[23665]_ ,
    \new_[23669]_ , \new_[23670]_ , \new_[23674]_ , \new_[23675]_ ,
    \new_[23676]_ , \new_[23679]_ , \new_[23683]_ , \new_[23684]_ ,
    \new_[23685]_ , \new_[23689]_ , \new_[23690]_ , \new_[23694]_ ,
    \new_[23695]_ , \new_[23696]_ , \new_[23699]_ , \new_[23703]_ ,
    \new_[23704]_ , \new_[23705]_ , \new_[23709]_ , \new_[23710]_ ,
    \new_[23714]_ , \new_[23715]_ , \new_[23716]_ , \new_[23719]_ ,
    \new_[23723]_ , \new_[23724]_ , \new_[23725]_ , \new_[23729]_ ,
    \new_[23730]_ , \new_[23734]_ , \new_[23735]_ , \new_[23736]_ ,
    \new_[23739]_ , \new_[23743]_ , \new_[23744]_ , \new_[23745]_ ,
    \new_[23749]_ , \new_[23750]_ , \new_[23754]_ , \new_[23755]_ ,
    \new_[23756]_ , \new_[23759]_ , \new_[23763]_ , \new_[23764]_ ,
    \new_[23765]_ , \new_[23769]_ , \new_[23770]_ , \new_[23774]_ ,
    \new_[23775]_ , \new_[23776]_ , \new_[23779]_ , \new_[23783]_ ,
    \new_[23784]_ , \new_[23785]_ , \new_[23789]_ , \new_[23790]_ ,
    \new_[23794]_ , \new_[23795]_ , \new_[23796]_ , \new_[23799]_ ,
    \new_[23803]_ , \new_[23804]_ , \new_[23805]_ , \new_[23809]_ ,
    \new_[23810]_ , \new_[23814]_ , \new_[23815]_ , \new_[23816]_ ,
    \new_[23819]_ , \new_[23823]_ , \new_[23824]_ , \new_[23825]_ ,
    \new_[23829]_ , \new_[23830]_ , \new_[23834]_ , \new_[23835]_ ,
    \new_[23836]_ , \new_[23839]_ , \new_[23843]_ , \new_[23844]_ ,
    \new_[23845]_ , \new_[23849]_ , \new_[23850]_ , \new_[23854]_ ,
    \new_[23855]_ , \new_[23856]_ , \new_[23859]_ , \new_[23863]_ ,
    \new_[23864]_ , \new_[23865]_ , \new_[23869]_ , \new_[23870]_ ,
    \new_[23874]_ , \new_[23875]_ , \new_[23876]_ , \new_[23879]_ ,
    \new_[23883]_ , \new_[23884]_ , \new_[23885]_ , \new_[23889]_ ,
    \new_[23890]_ , \new_[23894]_ , \new_[23895]_ , \new_[23896]_ ,
    \new_[23899]_ , \new_[23903]_ , \new_[23904]_ , \new_[23905]_ ,
    \new_[23909]_ , \new_[23910]_ , \new_[23914]_ , \new_[23915]_ ,
    \new_[23916]_ , \new_[23919]_ , \new_[23923]_ , \new_[23924]_ ,
    \new_[23925]_ , \new_[23929]_ , \new_[23930]_ , \new_[23934]_ ,
    \new_[23935]_ , \new_[23936]_ , \new_[23939]_ , \new_[23943]_ ,
    \new_[23944]_ , \new_[23945]_ , \new_[23949]_ , \new_[23950]_ ,
    \new_[23954]_ , \new_[23955]_ , \new_[23956]_ , \new_[23959]_ ,
    \new_[23963]_ , \new_[23964]_ , \new_[23965]_ , \new_[23969]_ ,
    \new_[23970]_ , \new_[23974]_ , \new_[23975]_ , \new_[23976]_ ,
    \new_[23979]_ , \new_[23983]_ , \new_[23984]_ , \new_[23985]_ ,
    \new_[23989]_ , \new_[23990]_ , \new_[23994]_ , \new_[23995]_ ,
    \new_[23996]_ , \new_[23999]_ , \new_[24003]_ , \new_[24004]_ ,
    \new_[24005]_ , \new_[24009]_ , \new_[24010]_ , \new_[24014]_ ,
    \new_[24015]_ , \new_[24016]_ , \new_[24019]_ , \new_[24023]_ ,
    \new_[24024]_ , \new_[24025]_ , \new_[24029]_ , \new_[24030]_ ,
    \new_[24034]_ , \new_[24035]_ , \new_[24036]_ , \new_[24039]_ ,
    \new_[24043]_ , \new_[24044]_ , \new_[24045]_ , \new_[24049]_ ,
    \new_[24050]_ , \new_[24054]_ , \new_[24055]_ , \new_[24056]_ ,
    \new_[24059]_ , \new_[24063]_ , \new_[24064]_ , \new_[24065]_ ,
    \new_[24069]_ , \new_[24070]_ , \new_[24074]_ , \new_[24075]_ ,
    \new_[24076]_ , \new_[24079]_ , \new_[24083]_ , \new_[24084]_ ,
    \new_[24085]_ , \new_[24089]_ , \new_[24090]_ , \new_[24094]_ ,
    \new_[24095]_ , \new_[24096]_ , \new_[24099]_ , \new_[24103]_ ,
    \new_[24104]_ , \new_[24105]_ , \new_[24109]_ , \new_[24110]_ ,
    \new_[24114]_ , \new_[24115]_ , \new_[24116]_ , \new_[24119]_ ,
    \new_[24123]_ , \new_[24124]_ , \new_[24125]_ , \new_[24129]_ ,
    \new_[24130]_ , \new_[24134]_ , \new_[24135]_ , \new_[24136]_ ,
    \new_[24139]_ , \new_[24143]_ , \new_[24144]_ , \new_[24145]_ ,
    \new_[24149]_ , \new_[24150]_ , \new_[24154]_ , \new_[24155]_ ,
    \new_[24156]_ , \new_[24159]_ , \new_[24163]_ , \new_[24164]_ ,
    \new_[24165]_ , \new_[24169]_ , \new_[24170]_ , \new_[24174]_ ,
    \new_[24175]_ , \new_[24176]_ , \new_[24179]_ , \new_[24183]_ ,
    \new_[24184]_ , \new_[24185]_ , \new_[24189]_ , \new_[24190]_ ,
    \new_[24194]_ , \new_[24195]_ , \new_[24196]_ , \new_[24199]_ ,
    \new_[24203]_ , \new_[24204]_ , \new_[24205]_ , \new_[24209]_ ,
    \new_[24210]_ , \new_[24214]_ , \new_[24215]_ , \new_[24216]_ ,
    \new_[24219]_ , \new_[24223]_ , \new_[24224]_ , \new_[24225]_ ,
    \new_[24229]_ , \new_[24230]_ , \new_[24234]_ , \new_[24235]_ ,
    \new_[24236]_ , \new_[24239]_ , \new_[24243]_ , \new_[24244]_ ,
    \new_[24245]_ , \new_[24249]_ , \new_[24250]_ , \new_[24254]_ ,
    \new_[24255]_ , \new_[24256]_ , \new_[24259]_ , \new_[24263]_ ,
    \new_[24264]_ , \new_[24265]_ , \new_[24269]_ , \new_[24270]_ ,
    \new_[24274]_ , \new_[24275]_ , \new_[24276]_ , \new_[24279]_ ,
    \new_[24283]_ , \new_[24284]_ , \new_[24285]_ , \new_[24289]_ ,
    \new_[24290]_ , \new_[24294]_ , \new_[24295]_ , \new_[24296]_ ,
    \new_[24299]_ , \new_[24303]_ , \new_[24304]_ , \new_[24305]_ ,
    \new_[24309]_ , \new_[24310]_ , \new_[24314]_ , \new_[24315]_ ,
    \new_[24316]_ , \new_[24319]_ , \new_[24323]_ , \new_[24324]_ ,
    \new_[24325]_ , \new_[24329]_ , \new_[24330]_ , \new_[24334]_ ,
    \new_[24335]_ , \new_[24336]_ , \new_[24339]_ , \new_[24343]_ ,
    \new_[24344]_ , \new_[24345]_ , \new_[24349]_ , \new_[24350]_ ,
    \new_[24354]_ , \new_[24355]_ , \new_[24356]_ , \new_[24359]_ ,
    \new_[24363]_ , \new_[24364]_ , \new_[24365]_ , \new_[24369]_ ,
    \new_[24370]_ , \new_[24374]_ , \new_[24375]_ , \new_[24376]_ ,
    \new_[24379]_ , \new_[24383]_ , \new_[24384]_ , \new_[24385]_ ,
    \new_[24389]_ , \new_[24390]_ , \new_[24394]_ , \new_[24395]_ ,
    \new_[24396]_ , \new_[24399]_ , \new_[24403]_ , \new_[24404]_ ,
    \new_[24405]_ , \new_[24409]_ , \new_[24410]_ , \new_[24414]_ ,
    \new_[24415]_ , \new_[24416]_ , \new_[24419]_ , \new_[24423]_ ,
    \new_[24424]_ , \new_[24425]_ , \new_[24429]_ , \new_[24430]_ ,
    \new_[24434]_ , \new_[24435]_ , \new_[24436]_ , \new_[24439]_ ,
    \new_[24443]_ , \new_[24444]_ , \new_[24445]_ , \new_[24449]_ ,
    \new_[24450]_ , \new_[24454]_ , \new_[24455]_ , \new_[24456]_ ,
    \new_[24459]_ , \new_[24463]_ , \new_[24464]_ , \new_[24465]_ ,
    \new_[24469]_ , \new_[24470]_ , \new_[24474]_ , \new_[24475]_ ,
    \new_[24476]_ , \new_[24479]_ , \new_[24483]_ , \new_[24484]_ ,
    \new_[24485]_ , \new_[24489]_ , \new_[24490]_ , \new_[24494]_ ,
    \new_[24495]_ , \new_[24496]_ , \new_[24500]_ , \new_[24501]_ ,
    \new_[24505]_ , \new_[24506]_ , \new_[24507]_ , \new_[24511]_ ,
    \new_[24512]_ , \new_[24516]_ , \new_[24517]_ , \new_[24518]_ ,
    \new_[24522]_ , \new_[24523]_ , \new_[24527]_ , \new_[24528]_ ,
    \new_[24529]_ , \new_[24533]_ , \new_[24534]_ , \new_[24538]_ ,
    \new_[24539]_ , \new_[24540]_ , \new_[24544]_ , \new_[24545]_ ,
    \new_[24549]_ , \new_[24550]_ , \new_[24551]_ , \new_[24555]_ ,
    \new_[24556]_ , \new_[24560]_ , \new_[24561]_ , \new_[24562]_ ,
    \new_[24566]_ , \new_[24567]_ , \new_[24571]_ , \new_[24572]_ ,
    \new_[24573]_ , \new_[24577]_ , \new_[24578]_ , \new_[24582]_ ,
    \new_[24583]_ , \new_[24584]_ , \new_[24588]_ , \new_[24589]_ ,
    \new_[24593]_ , \new_[24594]_ , \new_[24595]_ , \new_[24599]_ ,
    \new_[24600]_ , \new_[24604]_ , \new_[24605]_ , \new_[24606]_ ,
    \new_[24610]_ , \new_[24611]_ , \new_[24615]_ , \new_[24616]_ ,
    \new_[24617]_ , \new_[24621]_ , \new_[24622]_ , \new_[24626]_ ,
    \new_[24627]_ , \new_[24628]_ , \new_[24632]_ , \new_[24633]_ ,
    \new_[24637]_ , \new_[24638]_ , \new_[24639]_ , \new_[24643]_ ,
    \new_[24644]_ , \new_[24648]_ , \new_[24649]_ , \new_[24650]_ ,
    \new_[24654]_ , \new_[24655]_ , \new_[24659]_ , \new_[24660]_ ,
    \new_[24661]_ , \new_[24665]_ , \new_[24666]_ , \new_[24670]_ ,
    \new_[24671]_ , \new_[24672]_ , \new_[24676]_ , \new_[24677]_ ,
    \new_[24681]_ , \new_[24682]_ , \new_[24683]_ , \new_[24687]_ ,
    \new_[24688]_ , \new_[24692]_ , \new_[24693]_ , \new_[24694]_ ,
    \new_[24698]_ , \new_[24699]_ , \new_[24703]_ , \new_[24704]_ ,
    \new_[24705]_ , \new_[24709]_ , \new_[24710]_ , \new_[24714]_ ,
    \new_[24715]_ , \new_[24716]_ , \new_[24720]_ , \new_[24721]_ ,
    \new_[24725]_ , \new_[24726]_ , \new_[24727]_ , \new_[24731]_ ,
    \new_[24732]_ , \new_[24736]_ , \new_[24737]_ , \new_[24738]_ ,
    \new_[24742]_ , \new_[24743]_ , \new_[24747]_ , \new_[24748]_ ,
    \new_[24749]_ , \new_[24753]_ , \new_[24754]_ , \new_[24758]_ ,
    \new_[24759]_ , \new_[24760]_ , \new_[24764]_ , \new_[24765]_ ,
    \new_[24769]_ , \new_[24770]_ , \new_[24771]_ , \new_[24775]_ ,
    \new_[24776]_ , \new_[24780]_ , \new_[24781]_ , \new_[24782]_ ,
    \new_[24786]_ , \new_[24787]_ , \new_[24791]_ , \new_[24792]_ ,
    \new_[24793]_ , \new_[24797]_ , \new_[24798]_ , \new_[24802]_ ,
    \new_[24803]_ , \new_[24804]_ , \new_[24808]_ , \new_[24809]_ ,
    \new_[24813]_ , \new_[24814]_ , \new_[24815]_ , \new_[24819]_ ,
    \new_[24820]_ , \new_[24824]_ , \new_[24825]_ , \new_[24826]_ ,
    \new_[24830]_ , \new_[24831]_ , \new_[24835]_ , \new_[24836]_ ,
    \new_[24837]_ , \new_[24841]_ , \new_[24842]_ , \new_[24846]_ ,
    \new_[24847]_ , \new_[24848]_ , \new_[24852]_ , \new_[24853]_ ,
    \new_[24857]_ , \new_[24858]_ , \new_[24859]_ , \new_[24863]_ ,
    \new_[24864]_ , \new_[24868]_ , \new_[24869]_ , \new_[24870]_ ,
    \new_[24874]_ , \new_[24875]_ , \new_[24879]_ , \new_[24880]_ ,
    \new_[24881]_ , \new_[24885]_ , \new_[24886]_ , \new_[24890]_ ,
    \new_[24891]_ , \new_[24892]_ , \new_[24896]_ , \new_[24897]_ ,
    \new_[24901]_ , \new_[24902]_ , \new_[24903]_ , \new_[24907]_ ,
    \new_[24908]_ , \new_[24912]_ , \new_[24913]_ , \new_[24914]_ ,
    \new_[24918]_ , \new_[24919]_ , \new_[24923]_ , \new_[24924]_ ,
    \new_[24925]_ , \new_[24929]_ , \new_[24930]_ , \new_[24934]_ ,
    \new_[24935]_ , \new_[24936]_ , \new_[24940]_ , \new_[24941]_ ,
    \new_[24945]_ , \new_[24946]_ , \new_[24947]_ , \new_[24951]_ ,
    \new_[24952]_ , \new_[24956]_ , \new_[24957]_ , \new_[24958]_ ,
    \new_[24962]_ , \new_[24963]_ , \new_[24967]_ , \new_[24968]_ ,
    \new_[24969]_ , \new_[24973]_ , \new_[24974]_ , \new_[24978]_ ,
    \new_[24979]_ , \new_[24980]_ , \new_[24984]_ , \new_[24985]_ ,
    \new_[24989]_ , \new_[24990]_ , \new_[24991]_ , \new_[24995]_ ,
    \new_[24996]_ , \new_[25000]_ , \new_[25001]_ , \new_[25002]_ ,
    \new_[25006]_ , \new_[25007]_ , \new_[25011]_ , \new_[25012]_ ,
    \new_[25013]_ , \new_[25017]_ , \new_[25018]_ , \new_[25022]_ ,
    \new_[25023]_ , \new_[25024]_ , \new_[25028]_ , \new_[25029]_ ,
    \new_[25033]_ , \new_[25034]_ , \new_[25035]_ , \new_[25039]_ ,
    \new_[25040]_ , \new_[25044]_ , \new_[25045]_ , \new_[25046]_ ,
    \new_[25050]_ , \new_[25051]_ , \new_[25055]_ , \new_[25056]_ ,
    \new_[25057]_ , \new_[25061]_ , \new_[25062]_ , \new_[25066]_ ,
    \new_[25067]_ , \new_[25068]_ , \new_[25072]_ , \new_[25073]_ ,
    \new_[25077]_ , \new_[25078]_ , \new_[25079]_ , \new_[25083]_ ,
    \new_[25084]_ , \new_[25088]_ , \new_[25089]_ , \new_[25090]_ ,
    \new_[25094]_ , \new_[25095]_ , \new_[25099]_ , \new_[25100]_ ,
    \new_[25101]_ , \new_[25105]_ , \new_[25106]_ , \new_[25110]_ ,
    \new_[25111]_ , \new_[25112]_ , \new_[25116]_ , \new_[25117]_ ,
    \new_[25121]_ , \new_[25122]_ , \new_[25123]_ , \new_[25127]_ ,
    \new_[25128]_ , \new_[25132]_ , \new_[25133]_ , \new_[25134]_ ,
    \new_[25138]_ , \new_[25139]_ , \new_[25143]_ , \new_[25144]_ ,
    \new_[25145]_ , \new_[25149]_ , \new_[25150]_ , \new_[25154]_ ,
    \new_[25155]_ , \new_[25156]_ , \new_[25160]_ , \new_[25161]_ ,
    \new_[25165]_ , \new_[25166]_ , \new_[25167]_ , \new_[25171]_ ,
    \new_[25172]_ , \new_[25176]_ , \new_[25177]_ , \new_[25178]_ ,
    \new_[25182]_ , \new_[25183]_ , \new_[25187]_ , \new_[25188]_ ,
    \new_[25189]_ , \new_[25193]_ , \new_[25194]_ , \new_[25198]_ ,
    \new_[25199]_ , \new_[25200]_ , \new_[25204]_ , \new_[25205]_ ,
    \new_[25209]_ , \new_[25210]_ , \new_[25211]_ , \new_[25215]_ ,
    \new_[25216]_ , \new_[25220]_ , \new_[25221]_ , \new_[25222]_ ,
    \new_[25226]_ , \new_[25227]_ , \new_[25231]_ , \new_[25232]_ ,
    \new_[25233]_ , \new_[25237]_ , \new_[25238]_ , \new_[25242]_ ,
    \new_[25243]_ , \new_[25244]_ , \new_[25248]_ , \new_[25249]_ ,
    \new_[25253]_ , \new_[25254]_ , \new_[25255]_ , \new_[25259]_ ,
    \new_[25260]_ , \new_[25264]_ , \new_[25265]_ , \new_[25266]_ ,
    \new_[25270]_ , \new_[25271]_ , \new_[25275]_ , \new_[25276]_ ,
    \new_[25277]_ , \new_[25281]_ , \new_[25282]_ , \new_[25286]_ ,
    \new_[25287]_ , \new_[25288]_ , \new_[25292]_ , \new_[25293]_ ,
    \new_[25297]_ , \new_[25298]_ , \new_[25299]_ , \new_[25303]_ ,
    \new_[25304]_ , \new_[25308]_ , \new_[25309]_ , \new_[25310]_ ,
    \new_[25314]_ , \new_[25315]_ , \new_[25319]_ , \new_[25320]_ ,
    \new_[25321]_ , \new_[25325]_ , \new_[25326]_ , \new_[25330]_ ,
    \new_[25331]_ , \new_[25332]_ , \new_[25336]_ , \new_[25337]_ ,
    \new_[25341]_ , \new_[25342]_ , \new_[25343]_ , \new_[25347]_ ,
    \new_[25348]_ , \new_[25352]_ , \new_[25353]_ , \new_[25354]_ ,
    \new_[25358]_ , \new_[25359]_ , \new_[25363]_ , \new_[25364]_ ,
    \new_[25365]_ , \new_[25369]_ , \new_[25370]_ , \new_[25374]_ ,
    \new_[25375]_ , \new_[25376]_ , \new_[25380]_ , \new_[25381]_ ,
    \new_[25385]_ , \new_[25386]_ , \new_[25387]_ , \new_[25391]_ ,
    \new_[25392]_ , \new_[25396]_ , \new_[25397]_ , \new_[25398]_ ,
    \new_[25402]_ , \new_[25403]_ , \new_[25407]_ , \new_[25408]_ ,
    \new_[25409]_ , \new_[25413]_ , \new_[25414]_ , \new_[25418]_ ,
    \new_[25419]_ , \new_[25420]_ , \new_[25424]_ , \new_[25425]_ ,
    \new_[25429]_ , \new_[25430]_ , \new_[25431]_ , \new_[25435]_ ,
    \new_[25436]_ , \new_[25440]_ , \new_[25441]_ , \new_[25442]_ ,
    \new_[25446]_ , \new_[25447]_ , \new_[25451]_ , \new_[25452]_ ,
    \new_[25453]_ , \new_[25457]_ , \new_[25458]_ , \new_[25462]_ ,
    \new_[25463]_ , \new_[25464]_ , \new_[25468]_ , \new_[25469]_ ,
    \new_[25473]_ , \new_[25474]_ , \new_[25475]_ , \new_[25479]_ ,
    \new_[25480]_ , \new_[25484]_ , \new_[25485]_ , \new_[25486]_ ,
    \new_[25490]_ , \new_[25491]_ , \new_[25495]_ , \new_[25496]_ ,
    \new_[25497]_ , \new_[25501]_ , \new_[25502]_ , \new_[25506]_ ,
    \new_[25507]_ , \new_[25508]_ , \new_[25512]_ , \new_[25513]_ ,
    \new_[25517]_ , \new_[25518]_ , \new_[25519]_ , \new_[25523]_ ,
    \new_[25524]_ , \new_[25528]_ , \new_[25529]_ , \new_[25530]_ ,
    \new_[25534]_ , \new_[25535]_ , \new_[25539]_ , \new_[25540]_ ,
    \new_[25541]_ , \new_[25545]_ , \new_[25546]_ , \new_[25550]_ ,
    \new_[25551]_ , \new_[25552]_ , \new_[25556]_ , \new_[25557]_ ,
    \new_[25561]_ , \new_[25562]_ , \new_[25563]_ , \new_[25567]_ ,
    \new_[25568]_ , \new_[25572]_ , \new_[25573]_ , \new_[25574]_ ,
    \new_[25578]_ , \new_[25579]_ , \new_[25583]_ , \new_[25584]_ ,
    \new_[25585]_ , \new_[25589]_ , \new_[25590]_ , \new_[25594]_ ,
    \new_[25595]_ , \new_[25596]_ , \new_[25600]_ , \new_[25601]_ ,
    \new_[25605]_ , \new_[25606]_ , \new_[25607]_ , \new_[25611]_ ,
    \new_[25612]_ , \new_[25616]_ , \new_[25617]_ , \new_[25618]_ ,
    \new_[25622]_ , \new_[25623]_ , \new_[25627]_ , \new_[25628]_ ,
    \new_[25629]_ , \new_[25633]_ , \new_[25634]_ , \new_[25638]_ ,
    \new_[25639]_ , \new_[25640]_ , \new_[25644]_ , \new_[25645]_ ,
    \new_[25649]_ , \new_[25650]_ , \new_[25651]_ , \new_[25655]_ ,
    \new_[25656]_ , \new_[25660]_ , \new_[25661]_ , \new_[25662]_ ,
    \new_[25666]_ , \new_[25667]_ , \new_[25671]_ , \new_[25672]_ ,
    \new_[25673]_ , \new_[25677]_ , \new_[25678]_ , \new_[25682]_ ,
    \new_[25683]_ , \new_[25684]_ , \new_[25688]_ , \new_[25689]_ ,
    \new_[25693]_ , \new_[25694]_ , \new_[25695]_ , \new_[25699]_ ,
    \new_[25700]_ , \new_[25704]_ , \new_[25705]_ , \new_[25706]_ ,
    \new_[25710]_ , \new_[25711]_ , \new_[25715]_ , \new_[25716]_ ,
    \new_[25717]_ , \new_[25721]_ , \new_[25722]_ , \new_[25726]_ ,
    \new_[25727]_ , \new_[25728]_ , \new_[25732]_ , \new_[25733]_ ,
    \new_[25737]_ , \new_[25738]_ , \new_[25739]_ , \new_[25743]_ ,
    \new_[25744]_ , \new_[25748]_ , \new_[25749]_ , \new_[25750]_ ,
    \new_[25754]_ , \new_[25755]_ , \new_[25759]_ , \new_[25760]_ ,
    \new_[25761]_ , \new_[25765]_ , \new_[25766]_ , \new_[25770]_ ,
    \new_[25771]_ , \new_[25772]_ , \new_[25776]_ , \new_[25777]_ ,
    \new_[25781]_ , \new_[25782]_ , \new_[25783]_ , \new_[25787]_ ,
    \new_[25788]_ , \new_[25792]_ , \new_[25793]_ , \new_[25794]_ ,
    \new_[25798]_ , \new_[25799]_ , \new_[25803]_ , \new_[25804]_ ,
    \new_[25805]_ , \new_[25809]_ , \new_[25810]_ , \new_[25814]_ ,
    \new_[25815]_ , \new_[25816]_ , \new_[25820]_ , \new_[25821]_ ,
    \new_[25825]_ , \new_[25826]_ , \new_[25827]_ , \new_[25831]_ ,
    \new_[25832]_ , \new_[25836]_ , \new_[25837]_ , \new_[25838]_ ,
    \new_[25842]_ , \new_[25843]_ , \new_[25847]_ , \new_[25848]_ ,
    \new_[25849]_ , \new_[25853]_ , \new_[25854]_ , \new_[25858]_ ,
    \new_[25859]_ , \new_[25860]_ , \new_[25864]_ , \new_[25865]_ ,
    \new_[25869]_ , \new_[25870]_ , \new_[25871]_ , \new_[25875]_ ,
    \new_[25876]_ , \new_[25880]_ , \new_[25881]_ , \new_[25882]_ ,
    \new_[25886]_ , \new_[25887]_ , \new_[25891]_ , \new_[25892]_ ,
    \new_[25893]_ , \new_[25897]_ , \new_[25898]_ , \new_[25902]_ ,
    \new_[25903]_ , \new_[25904]_ , \new_[25908]_ , \new_[25909]_ ,
    \new_[25913]_ , \new_[25914]_ , \new_[25915]_ , \new_[25919]_ ,
    \new_[25920]_ , \new_[25924]_ , \new_[25925]_ , \new_[25926]_ ,
    \new_[25930]_ , \new_[25931]_ , \new_[25935]_ , \new_[25936]_ ,
    \new_[25937]_ , \new_[25941]_ , \new_[25942]_ , \new_[25946]_ ,
    \new_[25947]_ , \new_[25948]_ , \new_[25952]_ , \new_[25953]_ ,
    \new_[25957]_ , \new_[25958]_ , \new_[25959]_ , \new_[25963]_ ,
    \new_[25964]_ , \new_[25968]_ , \new_[25969]_ , \new_[25970]_ ,
    \new_[25974]_ , \new_[25975]_ , \new_[25979]_ , \new_[25980]_ ,
    \new_[25981]_ , \new_[25985]_ , \new_[25986]_ , \new_[25990]_ ,
    \new_[25991]_ , \new_[25992]_ , \new_[25996]_ , \new_[25997]_ ,
    \new_[26001]_ , \new_[26002]_ , \new_[26003]_ , \new_[26007]_ ,
    \new_[26008]_ , \new_[26012]_ , \new_[26013]_ , \new_[26014]_ ,
    \new_[26018]_ , \new_[26019]_ , \new_[26023]_ , \new_[26024]_ ,
    \new_[26025]_ , \new_[26029]_ , \new_[26030]_ , \new_[26034]_ ,
    \new_[26035]_ , \new_[26036]_ , \new_[26040]_ , \new_[26041]_ ,
    \new_[26045]_ , \new_[26046]_ , \new_[26047]_ , \new_[26051]_ ,
    \new_[26052]_ , \new_[26056]_ , \new_[26057]_ , \new_[26058]_ ,
    \new_[26062]_ , \new_[26063]_ , \new_[26067]_ , \new_[26068]_ ,
    \new_[26069]_ , \new_[26073]_ , \new_[26074]_ , \new_[26078]_ ,
    \new_[26079]_ , \new_[26080]_ , \new_[26084]_ , \new_[26085]_ ,
    \new_[26089]_ , \new_[26090]_ , \new_[26091]_ , \new_[26095]_ ,
    \new_[26096]_ , \new_[26100]_ , \new_[26101]_ , \new_[26102]_ ,
    \new_[26106]_ , \new_[26107]_ , \new_[26111]_ , \new_[26112]_ ,
    \new_[26113]_ , \new_[26117]_ , \new_[26118]_ , \new_[26122]_ ,
    \new_[26123]_ , \new_[26124]_ , \new_[26128]_ , \new_[26129]_ ,
    \new_[26133]_ , \new_[26134]_ , \new_[26135]_ , \new_[26139]_ ,
    \new_[26140]_ , \new_[26144]_ , \new_[26145]_ , \new_[26146]_ ,
    \new_[26150]_ , \new_[26151]_ , \new_[26155]_ , \new_[26156]_ ,
    \new_[26157]_ , \new_[26161]_ , \new_[26162]_ , \new_[26166]_ ,
    \new_[26167]_ , \new_[26168]_ , \new_[26172]_ , \new_[26173]_ ,
    \new_[26177]_ , \new_[26178]_ , \new_[26179]_ , \new_[26183]_ ,
    \new_[26184]_ , \new_[26188]_ , \new_[26189]_ , \new_[26190]_ ,
    \new_[26194]_ , \new_[26195]_ , \new_[26199]_ , \new_[26200]_ ,
    \new_[26201]_ , \new_[26205]_ , \new_[26206]_ , \new_[26210]_ ,
    \new_[26211]_ , \new_[26212]_ , \new_[26216]_ , \new_[26217]_ ,
    \new_[26221]_ , \new_[26222]_ , \new_[26223]_ , \new_[26227]_ ,
    \new_[26228]_ , \new_[26232]_ , \new_[26233]_ , \new_[26234]_ ,
    \new_[26238]_ , \new_[26239]_ , \new_[26243]_ , \new_[26244]_ ,
    \new_[26245]_ , \new_[26249]_ , \new_[26250]_ , \new_[26254]_ ,
    \new_[26255]_ , \new_[26256]_ , \new_[26260]_ , \new_[26261]_ ,
    \new_[26265]_ , \new_[26266]_ , \new_[26267]_ , \new_[26271]_ ,
    \new_[26272]_ , \new_[26276]_ , \new_[26277]_ , \new_[26278]_ ,
    \new_[26282]_ , \new_[26283]_ , \new_[26287]_ , \new_[26288]_ ,
    \new_[26289]_ , \new_[26293]_ , \new_[26294]_ , \new_[26298]_ ,
    \new_[26299]_ , \new_[26300]_ , \new_[26304]_ , \new_[26305]_ ,
    \new_[26309]_ , \new_[26310]_ , \new_[26311]_ , \new_[26315]_ ,
    \new_[26316]_ , \new_[26320]_ , \new_[26321]_ , \new_[26322]_ ,
    \new_[26326]_ , \new_[26327]_ , \new_[26331]_ , \new_[26332]_ ,
    \new_[26333]_ , \new_[26337]_ , \new_[26338]_ , \new_[26342]_ ,
    \new_[26343]_ , \new_[26344]_ , \new_[26348]_ , \new_[26349]_ ,
    \new_[26353]_ , \new_[26354]_ , \new_[26355]_ , \new_[26359]_ ,
    \new_[26360]_ , \new_[26364]_ , \new_[26365]_ , \new_[26366]_ ,
    \new_[26370]_ , \new_[26371]_ , \new_[26375]_ , \new_[26376]_ ,
    \new_[26377]_ , \new_[26381]_ , \new_[26382]_ , \new_[26386]_ ,
    \new_[26387]_ , \new_[26388]_ , \new_[26392]_ , \new_[26393]_ ,
    \new_[26397]_ , \new_[26398]_ , \new_[26399]_ , \new_[26403]_ ,
    \new_[26404]_ , \new_[26408]_ , \new_[26409]_ , \new_[26410]_ ,
    \new_[26414]_ , \new_[26415]_ , \new_[26419]_ , \new_[26420]_ ,
    \new_[26421]_ , \new_[26425]_ , \new_[26426]_ , \new_[26430]_ ,
    \new_[26431]_ , \new_[26432]_ , \new_[26436]_ , \new_[26437]_ ,
    \new_[26441]_ , \new_[26442]_ , \new_[26443]_ , \new_[26447]_ ,
    \new_[26448]_ , \new_[26452]_ , \new_[26453]_ , \new_[26454]_ ,
    \new_[26458]_ , \new_[26459]_ , \new_[26463]_ , \new_[26464]_ ,
    \new_[26465]_ , \new_[26469]_ , \new_[26470]_ , \new_[26474]_ ,
    \new_[26475]_ , \new_[26476]_ , \new_[26480]_ , \new_[26481]_ ,
    \new_[26485]_ , \new_[26486]_ , \new_[26487]_ , \new_[26491]_ ,
    \new_[26492]_ , \new_[26496]_ , \new_[26497]_ , \new_[26498]_ ,
    \new_[26502]_ , \new_[26503]_ , \new_[26507]_ , \new_[26508]_ ,
    \new_[26509]_ , \new_[26513]_ , \new_[26514]_ , \new_[26518]_ ,
    \new_[26519]_ , \new_[26520]_ , \new_[26524]_ , \new_[26525]_ ,
    \new_[26529]_ , \new_[26530]_ , \new_[26531]_ , \new_[26535]_ ,
    \new_[26536]_ , \new_[26540]_ , \new_[26541]_ , \new_[26542]_ ,
    \new_[26546]_ , \new_[26547]_ , \new_[26551]_ , \new_[26552]_ ,
    \new_[26553]_ , \new_[26557]_ , \new_[26558]_ , \new_[26562]_ ,
    \new_[26563]_ , \new_[26564]_ , \new_[26568]_ , \new_[26569]_ ,
    \new_[26573]_ , \new_[26574]_ , \new_[26575]_ , \new_[26579]_ ,
    \new_[26580]_ , \new_[26584]_ , \new_[26585]_ , \new_[26586]_ ,
    \new_[26590]_ , \new_[26591]_ , \new_[26595]_ , \new_[26596]_ ,
    \new_[26597]_ , \new_[26601]_ , \new_[26602]_ , \new_[26606]_ ,
    \new_[26607]_ , \new_[26608]_ , \new_[26612]_ , \new_[26613]_ ,
    \new_[26617]_ , \new_[26618]_ , \new_[26619]_ , \new_[26623]_ ,
    \new_[26624]_ , \new_[26628]_ , \new_[26629]_ , \new_[26630]_ ,
    \new_[26634]_ , \new_[26635]_ , \new_[26639]_ , \new_[26640]_ ,
    \new_[26641]_ , \new_[26645]_ , \new_[26646]_ , \new_[26650]_ ,
    \new_[26651]_ , \new_[26652]_ , \new_[26656]_ , \new_[26657]_ ,
    \new_[26661]_ , \new_[26662]_ , \new_[26663]_ , \new_[26667]_ ,
    \new_[26668]_ , \new_[26672]_ , \new_[26673]_ , \new_[26674]_ ,
    \new_[26678]_ , \new_[26679]_ , \new_[26683]_ , \new_[26684]_ ,
    \new_[26685]_ , \new_[26689]_ , \new_[26690]_ , \new_[26694]_ ,
    \new_[26695]_ , \new_[26696]_ , \new_[26700]_ , \new_[26701]_ ,
    \new_[26705]_ , \new_[26706]_ , \new_[26707]_ , \new_[26711]_ ,
    \new_[26712]_ , \new_[26716]_ , \new_[26717]_ , \new_[26718]_ ,
    \new_[26722]_ , \new_[26723]_ , \new_[26727]_ , \new_[26728]_ ,
    \new_[26729]_ , \new_[26733]_ , \new_[26734]_ , \new_[26738]_ ,
    \new_[26739]_ , \new_[26740]_ , \new_[26744]_ , \new_[26745]_ ,
    \new_[26749]_ , \new_[26750]_ , \new_[26751]_ , \new_[26755]_ ,
    \new_[26756]_ , \new_[26760]_ , \new_[26761]_ , \new_[26762]_ ,
    \new_[26766]_ , \new_[26767]_ , \new_[26771]_ , \new_[26772]_ ,
    \new_[26773]_ , \new_[26777]_ , \new_[26778]_ , \new_[26782]_ ,
    \new_[26783]_ , \new_[26784]_ , \new_[26788]_ , \new_[26789]_ ,
    \new_[26793]_ , \new_[26794]_ , \new_[26795]_ , \new_[26799]_ ,
    \new_[26800]_ , \new_[26804]_ , \new_[26805]_ , \new_[26806]_ ,
    \new_[26810]_ , \new_[26811]_ , \new_[26815]_ , \new_[26816]_ ,
    \new_[26817]_ , \new_[26821]_ , \new_[26822]_ , \new_[26826]_ ,
    \new_[26827]_ , \new_[26828]_ , \new_[26832]_ , \new_[26833]_ ,
    \new_[26837]_ , \new_[26838]_ , \new_[26839]_ , \new_[26843]_ ,
    \new_[26844]_ , \new_[26848]_ , \new_[26849]_ , \new_[26850]_ ,
    \new_[26854]_ , \new_[26855]_ , \new_[26859]_ , \new_[26860]_ ,
    \new_[26861]_ , \new_[26865]_ , \new_[26866]_ , \new_[26870]_ ,
    \new_[26871]_ , \new_[26872]_ , \new_[26876]_ , \new_[26877]_ ,
    \new_[26881]_ , \new_[26882]_ , \new_[26883]_ , \new_[26887]_ ,
    \new_[26888]_ , \new_[26892]_ , \new_[26893]_ , \new_[26894]_ ,
    \new_[26898]_ , \new_[26899]_ , \new_[26903]_ , \new_[26904]_ ,
    \new_[26905]_ , \new_[26909]_ , \new_[26910]_ , \new_[26914]_ ,
    \new_[26915]_ , \new_[26916]_ , \new_[26920]_ , \new_[26921]_ ,
    \new_[26925]_ , \new_[26926]_ , \new_[26927]_ , \new_[26931]_ ,
    \new_[26932]_ , \new_[26936]_ , \new_[26937]_ , \new_[26938]_ ,
    \new_[26942]_ , \new_[26943]_ , \new_[26947]_ , \new_[26948]_ ,
    \new_[26949]_ , \new_[26953]_ , \new_[26954]_ , \new_[26958]_ ,
    \new_[26959]_ , \new_[26960]_ , \new_[26964]_ , \new_[26965]_ ,
    \new_[26969]_ , \new_[26970]_ , \new_[26971]_ , \new_[26975]_ ,
    \new_[26976]_ , \new_[26980]_ , \new_[26981]_ , \new_[26982]_ ,
    \new_[26986]_ , \new_[26987]_ , \new_[26991]_ , \new_[26992]_ ,
    \new_[26993]_ , \new_[26997]_ , \new_[26998]_ , \new_[27002]_ ,
    \new_[27003]_ , \new_[27004]_ , \new_[27008]_ , \new_[27009]_ ,
    \new_[27013]_ , \new_[27014]_ , \new_[27015]_ , \new_[27019]_ ,
    \new_[27020]_ , \new_[27024]_ , \new_[27025]_ , \new_[27026]_ ,
    \new_[27030]_ , \new_[27031]_ , \new_[27035]_ , \new_[27036]_ ,
    \new_[27037]_ , \new_[27041]_ , \new_[27042]_ , \new_[27046]_ ,
    \new_[27047]_ , \new_[27048]_ , \new_[27052]_ , \new_[27053]_ ,
    \new_[27057]_ , \new_[27058]_ , \new_[27059]_ , \new_[27063]_ ,
    \new_[27064]_ , \new_[27068]_ , \new_[27069]_ , \new_[27070]_ ,
    \new_[27074]_ , \new_[27075]_ , \new_[27079]_ , \new_[27080]_ ,
    \new_[27081]_ , \new_[27085]_ , \new_[27086]_ , \new_[27090]_ ,
    \new_[27091]_ , \new_[27092]_ , \new_[27096]_ , \new_[27097]_ ,
    \new_[27101]_ , \new_[27102]_ , \new_[27103]_ , \new_[27107]_ ,
    \new_[27108]_ , \new_[27112]_ , \new_[27113]_ , \new_[27114]_ ,
    \new_[27118]_ , \new_[27119]_ , \new_[27123]_ , \new_[27124]_ ,
    \new_[27125]_ , \new_[27129]_ , \new_[27130]_ , \new_[27134]_ ,
    \new_[27135]_ , \new_[27136]_ , \new_[27140]_ , \new_[27141]_ ,
    \new_[27145]_ , \new_[27146]_ , \new_[27147]_ , \new_[27151]_ ,
    \new_[27152]_ , \new_[27156]_ , \new_[27157]_ , \new_[27158]_ ,
    \new_[27162]_ , \new_[27163]_ , \new_[27167]_ , \new_[27168]_ ,
    \new_[27169]_ , \new_[27173]_ , \new_[27174]_ , \new_[27178]_ ,
    \new_[27179]_ , \new_[27180]_ , \new_[27184]_ , \new_[27185]_ ,
    \new_[27189]_ , \new_[27190]_ , \new_[27191]_ , \new_[27195]_ ,
    \new_[27196]_ , \new_[27200]_ , \new_[27201]_ , \new_[27202]_ ,
    \new_[27206]_ , \new_[27207]_ , \new_[27211]_ , \new_[27212]_ ,
    \new_[27213]_ , \new_[27217]_ , \new_[27218]_ , \new_[27222]_ ,
    \new_[27223]_ , \new_[27224]_ , \new_[27228]_ , \new_[27229]_ ,
    \new_[27233]_ , \new_[27234]_ , \new_[27235]_ , \new_[27239]_ ,
    \new_[27240]_ , \new_[27244]_ , \new_[27245]_ , \new_[27246]_ ,
    \new_[27250]_ , \new_[27251]_ , \new_[27255]_ , \new_[27256]_ ,
    \new_[27257]_ , \new_[27261]_ , \new_[27262]_ , \new_[27266]_ ,
    \new_[27267]_ , \new_[27268]_ , \new_[27272]_ , \new_[27273]_ ,
    \new_[27277]_ , \new_[27278]_ , \new_[27279]_ , \new_[27283]_ ,
    \new_[27284]_ , \new_[27288]_ , \new_[27289]_ , \new_[27290]_ ,
    \new_[27294]_ , \new_[27295]_ , \new_[27299]_ , \new_[27300]_ ,
    \new_[27301]_ , \new_[27305]_ , \new_[27306]_ , \new_[27310]_ ,
    \new_[27311]_ , \new_[27312]_ , \new_[27316]_ , \new_[27317]_ ,
    \new_[27321]_ , \new_[27322]_ , \new_[27323]_ , \new_[27327]_ ,
    \new_[27328]_ , \new_[27332]_ , \new_[27333]_ , \new_[27334]_ ,
    \new_[27338]_ , \new_[27339]_ , \new_[27343]_ , \new_[27344]_ ,
    \new_[27345]_ , \new_[27349]_ , \new_[27350]_ , \new_[27354]_ ,
    \new_[27355]_ , \new_[27356]_ , \new_[27360]_ , \new_[27361]_ ,
    \new_[27365]_ , \new_[27366]_ , \new_[27367]_ , \new_[27371]_ ,
    \new_[27372]_ , \new_[27376]_ , \new_[27377]_ , \new_[27378]_ ,
    \new_[27382]_ , \new_[27383]_ , \new_[27387]_ , \new_[27388]_ ,
    \new_[27389]_ , \new_[27393]_ , \new_[27394]_ , \new_[27398]_ ,
    \new_[27399]_ , \new_[27400]_ , \new_[27404]_ , \new_[27405]_ ,
    \new_[27409]_ , \new_[27410]_ , \new_[27411]_ , \new_[27415]_ ,
    \new_[27416]_ , \new_[27420]_ , \new_[27421]_ , \new_[27422]_ ,
    \new_[27426]_ , \new_[27427]_ , \new_[27431]_ , \new_[27432]_ ,
    \new_[27433]_ , \new_[27437]_ , \new_[27438]_ , \new_[27442]_ ,
    \new_[27443]_ , \new_[27444]_ , \new_[27448]_ , \new_[27449]_ ,
    \new_[27453]_ , \new_[27454]_ , \new_[27455]_ , \new_[27459]_ ,
    \new_[27460]_ , \new_[27464]_ , \new_[27465]_ , \new_[27466]_ ,
    \new_[27470]_ , \new_[27471]_ , \new_[27475]_ , \new_[27476]_ ,
    \new_[27477]_ , \new_[27481]_ , \new_[27482]_ , \new_[27486]_ ,
    \new_[27487]_ , \new_[27488]_ , \new_[27492]_ , \new_[27493]_ ,
    \new_[27497]_ , \new_[27498]_ , \new_[27499]_ , \new_[27503]_ ,
    \new_[27504]_ , \new_[27508]_ , \new_[27509]_ , \new_[27510]_ ,
    \new_[27514]_ , \new_[27515]_ , \new_[27519]_ , \new_[27520]_ ,
    \new_[27521]_ , \new_[27525]_ , \new_[27526]_ , \new_[27530]_ ,
    \new_[27531]_ , \new_[27532]_ , \new_[27536]_ , \new_[27537]_ ,
    \new_[27541]_ , \new_[27542]_ , \new_[27543]_ , \new_[27547]_ ,
    \new_[27548]_ , \new_[27552]_ , \new_[27553]_ , \new_[27554]_ ,
    \new_[27558]_ , \new_[27559]_ , \new_[27563]_ , \new_[27564]_ ,
    \new_[27565]_ , \new_[27569]_ , \new_[27570]_ , \new_[27574]_ ,
    \new_[27575]_ , \new_[27576]_ , \new_[27580]_ , \new_[27581]_ ,
    \new_[27585]_ , \new_[27586]_ , \new_[27587]_ , \new_[27591]_ ,
    \new_[27592]_ , \new_[27596]_ , \new_[27597]_ , \new_[27598]_ ,
    \new_[27602]_ , \new_[27603]_ , \new_[27607]_ , \new_[27608]_ ,
    \new_[27609]_ , \new_[27613]_ , \new_[27614]_ , \new_[27618]_ ,
    \new_[27619]_ , \new_[27620]_ , \new_[27624]_ , \new_[27625]_ ,
    \new_[27629]_ , \new_[27630]_ , \new_[27631]_ , \new_[27635]_ ,
    \new_[27636]_ , \new_[27640]_ , \new_[27641]_ , \new_[27642]_ ,
    \new_[27646]_ , \new_[27647]_ , \new_[27651]_ , \new_[27652]_ ,
    \new_[27653]_ , \new_[27657]_ , \new_[27658]_ , \new_[27662]_ ,
    \new_[27663]_ , \new_[27664]_ , \new_[27668]_ , \new_[27669]_ ,
    \new_[27673]_ , \new_[27674]_ , \new_[27675]_ , \new_[27679]_ ,
    \new_[27680]_ , \new_[27684]_ , \new_[27685]_ , \new_[27686]_ ,
    \new_[27690]_ , \new_[27691]_ , \new_[27695]_ , \new_[27696]_ ,
    \new_[27697]_ , \new_[27701]_ , \new_[27702]_ , \new_[27706]_ ,
    \new_[27707]_ , \new_[27708]_ , \new_[27712]_ , \new_[27713]_ ,
    \new_[27717]_ , \new_[27718]_ , \new_[27719]_ , \new_[27723]_ ,
    \new_[27724]_ , \new_[27728]_ , \new_[27729]_ , \new_[27730]_ ,
    \new_[27734]_ , \new_[27735]_ , \new_[27739]_ , \new_[27740]_ ,
    \new_[27741]_ , \new_[27745]_ , \new_[27746]_ , \new_[27750]_ ,
    \new_[27751]_ , \new_[27752]_ , \new_[27756]_ , \new_[27757]_ ,
    \new_[27761]_ , \new_[27762]_ , \new_[27763]_ , \new_[27767]_ ,
    \new_[27768]_ , \new_[27772]_ , \new_[27773]_ , \new_[27774]_ ,
    \new_[27778]_ , \new_[27779]_ , \new_[27783]_ , \new_[27784]_ ,
    \new_[27785]_ , \new_[27789]_ , \new_[27790]_ , \new_[27794]_ ,
    \new_[27795]_ , \new_[27796]_ , \new_[27800]_ , \new_[27801]_ ,
    \new_[27805]_ , \new_[27806]_ , \new_[27807]_ , \new_[27811]_ ,
    \new_[27812]_ , \new_[27816]_ , \new_[27817]_ , \new_[27818]_ ,
    \new_[27822]_ , \new_[27823]_ , \new_[27827]_ , \new_[27828]_ ,
    \new_[27829]_ , \new_[27833]_ , \new_[27834]_ , \new_[27838]_ ,
    \new_[27839]_ , \new_[27840]_ , \new_[27844]_ , \new_[27845]_ ,
    \new_[27849]_ , \new_[27850]_ , \new_[27851]_ , \new_[27855]_ ,
    \new_[27856]_ , \new_[27860]_ , \new_[27861]_ , \new_[27862]_ ,
    \new_[27866]_ , \new_[27867]_ , \new_[27871]_ , \new_[27872]_ ,
    \new_[27873]_ , \new_[27877]_ , \new_[27878]_ , \new_[27882]_ ,
    \new_[27883]_ , \new_[27884]_ , \new_[27888]_ , \new_[27889]_ ,
    \new_[27893]_ , \new_[27894]_ , \new_[27895]_ , \new_[27899]_ ,
    \new_[27900]_ , \new_[27904]_ , \new_[27905]_ , \new_[27906]_ ,
    \new_[27910]_ , \new_[27911]_ , \new_[27915]_ , \new_[27916]_ ,
    \new_[27917]_ , \new_[27921]_ , \new_[27922]_ , \new_[27926]_ ,
    \new_[27927]_ , \new_[27928]_ , \new_[27932]_ , \new_[27933]_ ,
    \new_[27937]_ , \new_[27938]_ , \new_[27939]_ , \new_[27943]_ ,
    \new_[27944]_ , \new_[27948]_ , \new_[27949]_ , \new_[27950]_ ,
    \new_[27954]_ , \new_[27955]_ , \new_[27959]_ , \new_[27960]_ ,
    \new_[27961]_ , \new_[27965]_ , \new_[27966]_ , \new_[27970]_ ,
    \new_[27971]_ , \new_[27972]_ , \new_[27976]_ , \new_[27977]_ ,
    \new_[27981]_ , \new_[27982]_ , \new_[27983]_ , \new_[27987]_ ,
    \new_[27988]_ , \new_[27992]_ , \new_[27993]_ , \new_[27994]_ ,
    \new_[27998]_ , \new_[27999]_ , \new_[28003]_ , \new_[28004]_ ,
    \new_[28005]_ , \new_[28009]_ , \new_[28010]_ , \new_[28014]_ ,
    \new_[28015]_ , \new_[28016]_ , \new_[28020]_ , \new_[28021]_ ,
    \new_[28025]_ , \new_[28026]_ , \new_[28027]_ , \new_[28031]_ ,
    \new_[28032]_ , \new_[28036]_ , \new_[28037]_ , \new_[28038]_ ,
    \new_[28042]_ , \new_[28043]_ , \new_[28047]_ , \new_[28048]_ ,
    \new_[28049]_ , \new_[28053]_ , \new_[28054]_ , \new_[28058]_ ,
    \new_[28059]_ , \new_[28060]_ , \new_[28064]_ , \new_[28065]_ ,
    \new_[28069]_ , \new_[28070]_ , \new_[28071]_ , \new_[28075]_ ,
    \new_[28076]_ , \new_[28080]_ , \new_[28081]_ , \new_[28082]_ ,
    \new_[28086]_ , \new_[28087]_ , \new_[28091]_ , \new_[28092]_ ,
    \new_[28093]_ , \new_[28097]_ , \new_[28098]_ , \new_[28102]_ ,
    \new_[28103]_ , \new_[28104]_ , \new_[28108]_ , \new_[28109]_ ,
    \new_[28113]_ , \new_[28114]_ , \new_[28115]_ , \new_[28119]_ ,
    \new_[28120]_ , \new_[28124]_ , \new_[28125]_ , \new_[28126]_ ,
    \new_[28130]_ , \new_[28131]_ , \new_[28135]_ , \new_[28136]_ ,
    \new_[28137]_ , \new_[28141]_ , \new_[28142]_ , \new_[28146]_ ,
    \new_[28147]_ , \new_[28148]_ , \new_[28152]_ , \new_[28153]_ ,
    \new_[28157]_ , \new_[28158]_ , \new_[28159]_ , \new_[28163]_ ,
    \new_[28164]_ , \new_[28168]_ , \new_[28169]_ , \new_[28170]_ ,
    \new_[28174]_ , \new_[28175]_ , \new_[28179]_ , \new_[28180]_ ,
    \new_[28181]_ , \new_[28185]_ , \new_[28186]_ , \new_[28190]_ ,
    \new_[28191]_ , \new_[28192]_ , \new_[28196]_ , \new_[28197]_ ,
    \new_[28201]_ , \new_[28202]_ , \new_[28203]_ , \new_[28207]_ ,
    \new_[28208]_ , \new_[28212]_ , \new_[28213]_ , \new_[28214]_ ,
    \new_[28218]_ , \new_[28219]_ , \new_[28223]_ , \new_[28224]_ ,
    \new_[28225]_ , \new_[28229]_ , \new_[28230]_ , \new_[28234]_ ,
    \new_[28235]_ , \new_[28236]_ , \new_[28240]_ , \new_[28241]_ ,
    \new_[28245]_ , \new_[28246]_ , \new_[28247]_ , \new_[28251]_ ,
    \new_[28252]_ , \new_[28256]_ , \new_[28257]_ , \new_[28258]_ ,
    \new_[28262]_ , \new_[28263]_ , \new_[28267]_ , \new_[28268]_ ,
    \new_[28269]_ , \new_[28273]_ , \new_[28274]_ , \new_[28278]_ ,
    \new_[28279]_ , \new_[28280]_ , \new_[28284]_ , \new_[28285]_ ,
    \new_[28289]_ , \new_[28290]_ , \new_[28291]_ , \new_[28295]_ ,
    \new_[28296]_ , \new_[28300]_ , \new_[28301]_ , \new_[28302]_ ,
    \new_[28306]_ , \new_[28307]_ , \new_[28311]_ , \new_[28312]_ ,
    \new_[28313]_ , \new_[28317]_ , \new_[28318]_ , \new_[28322]_ ,
    \new_[28323]_ , \new_[28324]_ , \new_[28328]_ , \new_[28329]_ ,
    \new_[28333]_ , \new_[28334]_ , \new_[28335]_ , \new_[28339]_ ,
    \new_[28340]_ , \new_[28344]_ , \new_[28345]_ , \new_[28346]_ ,
    \new_[28350]_ , \new_[28351]_ , \new_[28355]_ , \new_[28356]_ ,
    \new_[28357]_ , \new_[28361]_ , \new_[28362]_ , \new_[28366]_ ,
    \new_[28367]_ , \new_[28368]_ , \new_[28372]_ , \new_[28373]_ ,
    \new_[28377]_ , \new_[28378]_ , \new_[28379]_ , \new_[28383]_ ,
    \new_[28384]_ , \new_[28388]_ , \new_[28389]_ , \new_[28390]_ ,
    \new_[28394]_ , \new_[28395]_ , \new_[28399]_ , \new_[28400]_ ,
    \new_[28401]_ , \new_[28405]_ , \new_[28406]_ , \new_[28410]_ ,
    \new_[28411]_ , \new_[28412]_ , \new_[28416]_ , \new_[28417]_ ,
    \new_[28421]_ , \new_[28422]_ , \new_[28423]_ , \new_[28427]_ ,
    \new_[28428]_ , \new_[28432]_ , \new_[28433]_ , \new_[28434]_ ,
    \new_[28438]_ , \new_[28439]_ , \new_[28443]_ , \new_[28444]_ ,
    \new_[28445]_ , \new_[28449]_ , \new_[28450]_ , \new_[28454]_ ,
    \new_[28455]_ , \new_[28456]_ , \new_[28460]_ , \new_[28461]_ ,
    \new_[28465]_ , \new_[28466]_ , \new_[28467]_ , \new_[28471]_ ,
    \new_[28472]_ , \new_[28476]_ , \new_[28477]_ , \new_[28478]_ ,
    \new_[28482]_ , \new_[28483]_ , \new_[28487]_ , \new_[28488]_ ,
    \new_[28489]_ , \new_[28493]_ , \new_[28494]_ , \new_[28498]_ ,
    \new_[28499]_ , \new_[28500]_ , \new_[28504]_ , \new_[28505]_ ,
    \new_[28509]_ , \new_[28510]_ , \new_[28511]_ , \new_[28515]_ ,
    \new_[28516]_ , \new_[28520]_ , \new_[28521]_ , \new_[28522]_ ,
    \new_[28526]_ , \new_[28527]_ , \new_[28531]_ , \new_[28532]_ ,
    \new_[28533]_ , \new_[28537]_ , \new_[28538]_ , \new_[28542]_ ,
    \new_[28543]_ , \new_[28544]_ , \new_[28548]_ , \new_[28549]_ ,
    \new_[28553]_ , \new_[28554]_ , \new_[28555]_ , \new_[28559]_ ,
    \new_[28560]_ , \new_[28564]_ , \new_[28565]_ , \new_[28566]_ ,
    \new_[28570]_ , \new_[28571]_ , \new_[28575]_ , \new_[28576]_ ,
    \new_[28577]_ , \new_[28581]_ , \new_[28582]_ , \new_[28586]_ ,
    \new_[28587]_ , \new_[28588]_ , \new_[28592]_ , \new_[28593]_ ,
    \new_[28597]_ , \new_[28598]_ , \new_[28599]_ , \new_[28603]_ ,
    \new_[28604]_ , \new_[28608]_ , \new_[28609]_ , \new_[28610]_ ,
    \new_[28614]_ , \new_[28615]_ , \new_[28619]_ , \new_[28620]_ ,
    \new_[28621]_ , \new_[28625]_ , \new_[28626]_ , \new_[28630]_ ,
    \new_[28631]_ , \new_[28632]_ , \new_[28636]_ , \new_[28637]_ ,
    \new_[28641]_ , \new_[28642]_ , \new_[28643]_ , \new_[28647]_ ,
    \new_[28648]_ , \new_[28652]_ , \new_[28653]_ , \new_[28654]_ ,
    \new_[28658]_ , \new_[28659]_ , \new_[28663]_ , \new_[28664]_ ,
    \new_[28665]_ , \new_[28669]_ , \new_[28670]_ , \new_[28674]_ ,
    \new_[28675]_ , \new_[28676]_ , \new_[28680]_ , \new_[28681]_ ,
    \new_[28685]_ , \new_[28686]_ , \new_[28687]_ , \new_[28691]_ ,
    \new_[28692]_ , \new_[28696]_ , \new_[28697]_ , \new_[28698]_ ,
    \new_[28702]_ , \new_[28703]_ , \new_[28707]_ , \new_[28708]_ ,
    \new_[28709]_ , \new_[28713]_ , \new_[28714]_ , \new_[28718]_ ,
    \new_[28719]_ , \new_[28720]_ , \new_[28724]_ , \new_[28725]_ ,
    \new_[28729]_ , \new_[28730]_ , \new_[28731]_ , \new_[28735]_ ,
    \new_[28736]_ , \new_[28740]_ , \new_[28741]_ , \new_[28742]_ ,
    \new_[28746]_ , \new_[28747]_ , \new_[28751]_ , \new_[28752]_ ,
    \new_[28753]_ , \new_[28757]_ , \new_[28758]_ , \new_[28762]_ ,
    \new_[28763]_ , \new_[28764]_ , \new_[28768]_ , \new_[28769]_ ,
    \new_[28773]_ , \new_[28774]_ , \new_[28775]_ , \new_[28779]_ ,
    \new_[28780]_ , \new_[28784]_ , \new_[28785]_ , \new_[28786]_ ,
    \new_[28790]_ , \new_[28791]_ , \new_[28795]_ , \new_[28796]_ ,
    \new_[28797]_ , \new_[28801]_ , \new_[28802]_ , \new_[28806]_ ,
    \new_[28807]_ , \new_[28808]_ , \new_[28812]_ , \new_[28813]_ ,
    \new_[28817]_ , \new_[28818]_ , \new_[28819]_ , \new_[28823]_ ,
    \new_[28824]_ , \new_[28828]_ , \new_[28829]_ , \new_[28830]_ ,
    \new_[28834]_ , \new_[28835]_ , \new_[28839]_ , \new_[28840]_ ,
    \new_[28841]_ , \new_[28845]_ , \new_[28846]_ , \new_[28850]_ ,
    \new_[28851]_ , \new_[28852]_ , \new_[28856]_ , \new_[28857]_ ,
    \new_[28861]_ , \new_[28862]_ , \new_[28863]_ , \new_[28867]_ ,
    \new_[28868]_ , \new_[28872]_ , \new_[28873]_ , \new_[28874]_ ,
    \new_[28878]_ , \new_[28879]_ , \new_[28883]_ , \new_[28884]_ ,
    \new_[28885]_ , \new_[28889]_ , \new_[28890]_ , \new_[28894]_ ,
    \new_[28895]_ , \new_[28896]_ , \new_[28900]_ , \new_[28901]_ ,
    \new_[28905]_ , \new_[28906]_ , \new_[28907]_ , \new_[28911]_ ,
    \new_[28912]_ , \new_[28916]_ , \new_[28917]_ , \new_[28918]_ ,
    \new_[28922]_ , \new_[28923]_ , \new_[28927]_ , \new_[28928]_ ,
    \new_[28929]_ , \new_[28933]_ , \new_[28934]_ , \new_[28938]_ ,
    \new_[28939]_ , \new_[28940]_ , \new_[28944]_ , \new_[28945]_ ,
    \new_[28949]_ , \new_[28950]_ , \new_[28951]_ , \new_[28955]_ ,
    \new_[28956]_ , \new_[28960]_ , \new_[28961]_ , \new_[28962]_ ,
    \new_[28966]_ , \new_[28967]_ , \new_[28971]_ , \new_[28972]_ ,
    \new_[28973]_ , \new_[28977]_ , \new_[28978]_ , \new_[28982]_ ,
    \new_[28983]_ , \new_[28984]_ , \new_[28988]_ , \new_[28989]_ ,
    \new_[28993]_ , \new_[28994]_ , \new_[28995]_ , \new_[28999]_ ,
    \new_[29000]_ , \new_[29004]_ , \new_[29005]_ , \new_[29006]_ ,
    \new_[29010]_ , \new_[29011]_ , \new_[29015]_ , \new_[29016]_ ,
    \new_[29017]_ , \new_[29021]_ , \new_[29022]_ , \new_[29026]_ ,
    \new_[29027]_ , \new_[29028]_ , \new_[29032]_ , \new_[29033]_ ,
    \new_[29037]_ , \new_[29038]_ , \new_[29039]_ , \new_[29043]_ ,
    \new_[29044]_ , \new_[29048]_ , \new_[29049]_ , \new_[29050]_ ,
    \new_[29054]_ , \new_[29055]_ , \new_[29059]_ , \new_[29060]_ ,
    \new_[29061]_ , \new_[29065]_ , \new_[29066]_ , \new_[29070]_ ,
    \new_[29071]_ , \new_[29072]_ , \new_[29076]_ , \new_[29077]_ ,
    \new_[29081]_ , \new_[29082]_ , \new_[29083]_ , \new_[29087]_ ,
    \new_[29088]_ , \new_[29092]_ , \new_[29093]_ , \new_[29094]_ ,
    \new_[29098]_ , \new_[29099]_ , \new_[29103]_ , \new_[29104]_ ,
    \new_[29105]_ , \new_[29109]_ , \new_[29110]_ , \new_[29114]_ ,
    \new_[29115]_ , \new_[29116]_ , \new_[29120]_ , \new_[29121]_ ,
    \new_[29125]_ , \new_[29126]_ , \new_[29127]_ , \new_[29131]_ ,
    \new_[29132]_ , \new_[29136]_ , \new_[29137]_ , \new_[29138]_ ,
    \new_[29142]_ , \new_[29143]_ , \new_[29147]_ , \new_[29148]_ ,
    \new_[29149]_ , \new_[29153]_ , \new_[29154]_ , \new_[29158]_ ,
    \new_[29159]_ , \new_[29160]_ , \new_[29164]_ , \new_[29165]_ ,
    \new_[29169]_ , \new_[29170]_ , \new_[29171]_ , \new_[29175]_ ,
    \new_[29176]_ , \new_[29180]_ , \new_[29181]_ , \new_[29182]_ ,
    \new_[29186]_ , \new_[29187]_ , \new_[29191]_ , \new_[29192]_ ,
    \new_[29193]_ , \new_[29197]_ , \new_[29198]_ , \new_[29202]_ ,
    \new_[29203]_ , \new_[29204]_ , \new_[29208]_ , \new_[29209]_ ,
    \new_[29213]_ , \new_[29214]_ , \new_[29215]_ , \new_[29219]_ ,
    \new_[29220]_ , \new_[29224]_ , \new_[29225]_ , \new_[29226]_ ,
    \new_[29230]_ , \new_[29231]_ , \new_[29235]_ , \new_[29236]_ ,
    \new_[29237]_ , \new_[29241]_ , \new_[29242]_ , \new_[29246]_ ,
    \new_[29247]_ , \new_[29248]_ , \new_[29252]_ , \new_[29253]_ ,
    \new_[29257]_ , \new_[29258]_ , \new_[29259]_ , \new_[29263]_ ,
    \new_[29264]_ , \new_[29268]_ , \new_[29269]_ , \new_[29270]_ ,
    \new_[29274]_ , \new_[29275]_ , \new_[29279]_ , \new_[29280]_ ,
    \new_[29281]_ , \new_[29285]_ , \new_[29286]_ , \new_[29290]_ ,
    \new_[29291]_ , \new_[29292]_ , \new_[29296]_ , \new_[29297]_ ,
    \new_[29301]_ , \new_[29302]_ , \new_[29303]_ , \new_[29307]_ ,
    \new_[29308]_ , \new_[29312]_ , \new_[29313]_ , \new_[29314]_ ,
    \new_[29318]_ , \new_[29319]_ , \new_[29323]_ , \new_[29324]_ ,
    \new_[29325]_ , \new_[29329]_ , \new_[29330]_ , \new_[29334]_ ,
    \new_[29335]_ , \new_[29336]_ , \new_[29340]_ , \new_[29341]_ ,
    \new_[29345]_ , \new_[29346]_ , \new_[29347]_ , \new_[29351]_ ,
    \new_[29352]_ , \new_[29356]_ , \new_[29357]_ , \new_[29358]_ ,
    \new_[29362]_ , \new_[29363]_ , \new_[29367]_ , \new_[29368]_ ,
    \new_[29369]_ , \new_[29373]_ , \new_[29374]_ , \new_[29378]_ ,
    \new_[29379]_ , \new_[29380]_ , \new_[29384]_ , \new_[29385]_ ,
    \new_[29389]_ , \new_[29390]_ , \new_[29391]_ , \new_[29395]_ ,
    \new_[29396]_ , \new_[29400]_ , \new_[29401]_ , \new_[29402]_ ,
    \new_[29406]_ , \new_[29407]_ , \new_[29411]_ , \new_[29412]_ ,
    \new_[29413]_ , \new_[29417]_ , \new_[29418]_ , \new_[29422]_ ,
    \new_[29423]_ , \new_[29424]_ , \new_[29428]_ , \new_[29429]_ ,
    \new_[29433]_ , \new_[29434]_ , \new_[29435]_ , \new_[29439]_ ,
    \new_[29440]_ , \new_[29444]_ , \new_[29445]_ , \new_[29446]_ ,
    \new_[29450]_ , \new_[29451]_ , \new_[29455]_ , \new_[29456]_ ,
    \new_[29457]_ , \new_[29461]_ , \new_[29462]_ , \new_[29466]_ ,
    \new_[29467]_ , \new_[29468]_ , \new_[29472]_ , \new_[29473]_ ,
    \new_[29477]_ , \new_[29478]_ , \new_[29479]_ , \new_[29483]_ ,
    \new_[29484]_ , \new_[29488]_ , \new_[29489]_ , \new_[29490]_ ,
    \new_[29494]_ , \new_[29495]_ , \new_[29499]_ , \new_[29500]_ ,
    \new_[29501]_ , \new_[29505]_ , \new_[29506]_ , \new_[29510]_ ,
    \new_[29511]_ , \new_[29512]_ , \new_[29516]_ , \new_[29517]_ ,
    \new_[29521]_ , \new_[29522]_ , \new_[29523]_ , \new_[29527]_ ,
    \new_[29528]_ , \new_[29532]_ , \new_[29533]_ , \new_[29534]_ ,
    \new_[29538]_ , \new_[29539]_ , \new_[29543]_ , \new_[29544]_ ,
    \new_[29545]_ , \new_[29549]_ , \new_[29550]_ , \new_[29554]_ ,
    \new_[29555]_ , \new_[29556]_ , \new_[29560]_ , \new_[29561]_ ,
    \new_[29565]_ , \new_[29566]_ , \new_[29567]_ , \new_[29571]_ ,
    \new_[29572]_ , \new_[29576]_ , \new_[29577]_ , \new_[29578]_ ,
    \new_[29582]_ , \new_[29583]_ , \new_[29587]_ , \new_[29588]_ ,
    \new_[29589]_ , \new_[29593]_ , \new_[29594]_ , \new_[29598]_ ,
    \new_[29599]_ , \new_[29600]_ , \new_[29604]_ , \new_[29605]_ ,
    \new_[29609]_ , \new_[29610]_ , \new_[29611]_ , \new_[29615]_ ,
    \new_[29616]_ , \new_[29620]_ , \new_[29621]_ , \new_[29622]_ ,
    \new_[29626]_ , \new_[29627]_ , \new_[29631]_ , \new_[29632]_ ,
    \new_[29633]_ , \new_[29637]_ , \new_[29638]_ , \new_[29642]_ ,
    \new_[29643]_ , \new_[29644]_ , \new_[29648]_ , \new_[29649]_ ,
    \new_[29653]_ , \new_[29654]_ , \new_[29655]_ , \new_[29659]_ ,
    \new_[29660]_ , \new_[29664]_ , \new_[29665]_ , \new_[29666]_ ,
    \new_[29670]_ , \new_[29671]_ , \new_[29675]_ , \new_[29676]_ ,
    \new_[29677]_ , \new_[29681]_ , \new_[29682]_ , \new_[29686]_ ,
    \new_[29687]_ , \new_[29688]_ , \new_[29692]_ , \new_[29693]_ ,
    \new_[29697]_ , \new_[29698]_ , \new_[29699]_ , \new_[29703]_ ,
    \new_[29704]_ , \new_[29708]_ , \new_[29709]_ , \new_[29710]_ ,
    \new_[29714]_ , \new_[29715]_ , \new_[29719]_ , \new_[29720]_ ,
    \new_[29721]_ , \new_[29725]_ , \new_[29726]_ , \new_[29730]_ ,
    \new_[29731]_ , \new_[29732]_ , \new_[29736]_ , \new_[29737]_ ,
    \new_[29741]_ , \new_[29742]_ , \new_[29743]_ , \new_[29747]_ ,
    \new_[29748]_ , \new_[29752]_ , \new_[29753]_ , \new_[29754]_ ,
    \new_[29758]_ , \new_[29759]_ , \new_[29763]_ , \new_[29764]_ ,
    \new_[29765]_ , \new_[29769]_ , \new_[29770]_ , \new_[29774]_ ,
    \new_[29775]_ , \new_[29776]_ , \new_[29780]_ , \new_[29781]_ ,
    \new_[29785]_ , \new_[29786]_ , \new_[29787]_ , \new_[29791]_ ,
    \new_[29792]_ , \new_[29796]_ , \new_[29797]_ , \new_[29798]_ ,
    \new_[29802]_ , \new_[29803]_ , \new_[29807]_ , \new_[29808]_ ,
    \new_[29809]_ , \new_[29813]_ , \new_[29814]_ , \new_[29818]_ ,
    \new_[29819]_ , \new_[29820]_ , \new_[29824]_ , \new_[29825]_ ,
    \new_[29829]_ , \new_[29830]_ , \new_[29831]_ , \new_[29835]_ ,
    \new_[29836]_ , \new_[29840]_ , \new_[29841]_ , \new_[29842]_ ,
    \new_[29846]_ , \new_[29847]_ , \new_[29851]_ , \new_[29852]_ ,
    \new_[29853]_ , \new_[29857]_ , \new_[29858]_ , \new_[29862]_ ,
    \new_[29863]_ , \new_[29864]_ , \new_[29868]_ , \new_[29869]_ ,
    \new_[29873]_ , \new_[29874]_ , \new_[29875]_ , \new_[29879]_ ,
    \new_[29880]_ , \new_[29884]_ , \new_[29885]_ , \new_[29886]_ ,
    \new_[29890]_ , \new_[29891]_ , \new_[29895]_ , \new_[29896]_ ,
    \new_[29897]_ , \new_[29901]_ , \new_[29902]_ , \new_[29906]_ ,
    \new_[29907]_ , \new_[29908]_ , \new_[29912]_ , \new_[29913]_ ,
    \new_[29917]_ , \new_[29918]_ , \new_[29919]_ , \new_[29923]_ ,
    \new_[29924]_ , \new_[29928]_ , \new_[29929]_ , \new_[29930]_ ,
    \new_[29934]_ , \new_[29935]_ , \new_[29939]_ , \new_[29940]_ ,
    \new_[29941]_ , \new_[29945]_ , \new_[29946]_ , \new_[29950]_ ,
    \new_[29951]_ , \new_[29952]_ , \new_[29956]_ , \new_[29957]_ ,
    \new_[29961]_ , \new_[29962]_ , \new_[29963]_ , \new_[29967]_ ,
    \new_[29968]_ , \new_[29972]_ , \new_[29973]_ , \new_[29974]_ ,
    \new_[29978]_ , \new_[29979]_ , \new_[29983]_ , \new_[29984]_ ,
    \new_[29985]_ , \new_[29989]_ , \new_[29990]_ , \new_[29994]_ ,
    \new_[29995]_ , \new_[29996]_ , \new_[30000]_ , \new_[30001]_ ,
    \new_[30005]_ , \new_[30006]_ , \new_[30007]_ , \new_[30011]_ ,
    \new_[30012]_ , \new_[30016]_ , \new_[30017]_ , \new_[30018]_ ,
    \new_[30022]_ , \new_[30023]_ , \new_[30027]_ , \new_[30028]_ ,
    \new_[30029]_ , \new_[30033]_ , \new_[30034]_ , \new_[30038]_ ,
    \new_[30039]_ , \new_[30040]_ , \new_[30044]_ , \new_[30045]_ ,
    \new_[30049]_ , \new_[30050]_ , \new_[30051]_ , \new_[30055]_ ,
    \new_[30056]_ , \new_[30060]_ , \new_[30061]_ , \new_[30062]_ ,
    \new_[30066]_ , \new_[30067]_ , \new_[30071]_ , \new_[30072]_ ,
    \new_[30073]_ , \new_[30077]_ , \new_[30078]_ , \new_[30082]_ ,
    \new_[30083]_ , \new_[30084]_ , \new_[30088]_ , \new_[30089]_ ,
    \new_[30093]_ , \new_[30094]_ , \new_[30095]_ , \new_[30099]_ ,
    \new_[30100]_ , \new_[30104]_ , \new_[30105]_ , \new_[30106]_ ,
    \new_[30110]_ , \new_[30111]_ , \new_[30115]_ , \new_[30116]_ ,
    \new_[30117]_ , \new_[30121]_ , \new_[30122]_ , \new_[30126]_ ,
    \new_[30127]_ , \new_[30128]_ , \new_[30132]_ , \new_[30133]_ ,
    \new_[30137]_ , \new_[30138]_ , \new_[30139]_ , \new_[30143]_ ,
    \new_[30144]_ , \new_[30148]_ , \new_[30149]_ , \new_[30150]_ ,
    \new_[30154]_ , \new_[30155]_ , \new_[30159]_ , \new_[30160]_ ,
    \new_[30161]_ , \new_[30165]_ , \new_[30166]_ , \new_[30170]_ ,
    \new_[30171]_ , \new_[30172]_ , \new_[30176]_ , \new_[30177]_ ,
    \new_[30181]_ , \new_[30182]_ , \new_[30183]_ , \new_[30187]_ ,
    \new_[30188]_ , \new_[30192]_ , \new_[30193]_ , \new_[30194]_ ,
    \new_[30198]_ , \new_[30199]_ , \new_[30203]_ , \new_[30204]_ ,
    \new_[30205]_ , \new_[30209]_ , \new_[30210]_ , \new_[30214]_ ,
    \new_[30215]_ , \new_[30216]_ , \new_[30220]_ , \new_[30221]_ ,
    \new_[30225]_ , \new_[30226]_ , \new_[30227]_ , \new_[30231]_ ,
    \new_[30232]_ , \new_[30236]_ , \new_[30237]_ , \new_[30238]_ ,
    \new_[30242]_ , \new_[30243]_ , \new_[30247]_ , \new_[30248]_ ,
    \new_[30249]_ , \new_[30253]_ , \new_[30254]_ , \new_[30258]_ ,
    \new_[30259]_ , \new_[30260]_ , \new_[30264]_ , \new_[30265]_ ,
    \new_[30269]_ , \new_[30270]_ , \new_[30271]_ , \new_[30275]_ ,
    \new_[30276]_ , \new_[30280]_ , \new_[30281]_ , \new_[30282]_ ,
    \new_[30286]_ , \new_[30287]_ , \new_[30291]_ , \new_[30292]_ ,
    \new_[30293]_ , \new_[30297]_ , \new_[30298]_ , \new_[30302]_ ,
    \new_[30303]_ , \new_[30304]_ , \new_[30308]_ , \new_[30309]_ ,
    \new_[30313]_ , \new_[30314]_ , \new_[30315]_ , \new_[30319]_ ,
    \new_[30320]_ , \new_[30324]_ , \new_[30325]_ , \new_[30326]_ ,
    \new_[30330]_ , \new_[30331]_ , \new_[30335]_ , \new_[30336]_ ,
    \new_[30337]_ , \new_[30341]_ , \new_[30342]_ , \new_[30346]_ ,
    \new_[30347]_ , \new_[30348]_ , \new_[30352]_ , \new_[30353]_ ,
    \new_[30357]_ , \new_[30358]_ , \new_[30359]_ , \new_[30363]_ ,
    \new_[30364]_ , \new_[30368]_ , \new_[30369]_ , \new_[30370]_ ,
    \new_[30374]_ , \new_[30375]_ , \new_[30379]_ , \new_[30380]_ ,
    \new_[30381]_ , \new_[30385]_ , \new_[30386]_ , \new_[30390]_ ,
    \new_[30391]_ , \new_[30392]_ , \new_[30396]_ , \new_[30397]_ ,
    \new_[30401]_ , \new_[30402]_ , \new_[30403]_ , \new_[30407]_ ,
    \new_[30408]_ , \new_[30412]_ , \new_[30413]_ , \new_[30414]_ ,
    \new_[30418]_ , \new_[30419]_ , \new_[30423]_ , \new_[30424]_ ,
    \new_[30425]_ , \new_[30429]_ , \new_[30430]_ , \new_[30434]_ ,
    \new_[30435]_ , \new_[30436]_ , \new_[30440]_ , \new_[30441]_ ,
    \new_[30445]_ , \new_[30446]_ , \new_[30447]_ , \new_[30451]_ ,
    \new_[30452]_ , \new_[30456]_ , \new_[30457]_ , \new_[30458]_ ,
    \new_[30462]_ , \new_[30463]_ , \new_[30467]_ , \new_[30468]_ ,
    \new_[30469]_ , \new_[30473]_ , \new_[30474]_ , \new_[30478]_ ,
    \new_[30479]_ , \new_[30480]_ , \new_[30484]_ , \new_[30485]_ ,
    \new_[30489]_ , \new_[30490]_ , \new_[30491]_ , \new_[30495]_ ,
    \new_[30496]_ , \new_[30500]_ , \new_[30501]_ , \new_[30502]_ ,
    \new_[30506]_ , \new_[30507]_ , \new_[30511]_ , \new_[30512]_ ,
    \new_[30513]_ , \new_[30517]_ , \new_[30518]_ , \new_[30522]_ ,
    \new_[30523]_ , \new_[30524]_ , \new_[30528]_ , \new_[30529]_ ,
    \new_[30533]_ , \new_[30534]_ , \new_[30535]_ , \new_[30539]_ ,
    \new_[30540]_ , \new_[30544]_ , \new_[30545]_ , \new_[30546]_ ,
    \new_[30550]_ , \new_[30551]_ , \new_[30555]_ , \new_[30556]_ ,
    \new_[30557]_ , \new_[30561]_ , \new_[30562]_ , \new_[30566]_ ,
    \new_[30567]_ , \new_[30568]_ , \new_[30572]_ , \new_[30573]_ ,
    \new_[30577]_ , \new_[30578]_ , \new_[30579]_ , \new_[30583]_ ,
    \new_[30584]_ , \new_[30588]_ , \new_[30589]_ , \new_[30590]_ ,
    \new_[30594]_ , \new_[30595]_ , \new_[30599]_ , \new_[30600]_ ,
    \new_[30601]_ , \new_[30605]_ , \new_[30606]_ , \new_[30610]_ ,
    \new_[30611]_ , \new_[30612]_ , \new_[30616]_ , \new_[30617]_ ,
    \new_[30621]_ , \new_[30622]_ , \new_[30623]_ , \new_[30627]_ ,
    \new_[30628]_ , \new_[30632]_ , \new_[30633]_ , \new_[30634]_ ,
    \new_[30638]_ , \new_[30639]_ , \new_[30643]_ , \new_[30644]_ ,
    \new_[30645]_ , \new_[30649]_ , \new_[30650]_ , \new_[30654]_ ,
    \new_[30655]_ , \new_[30656]_ , \new_[30660]_ , \new_[30661]_ ,
    \new_[30665]_ , \new_[30666]_ , \new_[30667]_ , \new_[30671]_ ,
    \new_[30672]_ , \new_[30676]_ , \new_[30677]_ , \new_[30678]_ ,
    \new_[30682]_ , \new_[30683]_ , \new_[30687]_ , \new_[30688]_ ,
    \new_[30689]_ , \new_[30693]_ , \new_[30694]_ , \new_[30698]_ ,
    \new_[30699]_ , \new_[30700]_ , \new_[30704]_ , \new_[30705]_ ,
    \new_[30709]_ , \new_[30710]_ , \new_[30711]_ , \new_[30715]_ ,
    \new_[30716]_ , \new_[30720]_ , \new_[30721]_ , \new_[30722]_ ,
    \new_[30726]_ , \new_[30727]_ , \new_[30731]_ , \new_[30732]_ ,
    \new_[30733]_ , \new_[30737]_ , \new_[30738]_ , \new_[30742]_ ,
    \new_[30743]_ , \new_[30744]_ , \new_[30748]_ , \new_[30749]_ ,
    \new_[30753]_ , \new_[30754]_ , \new_[30755]_ , \new_[30759]_ ,
    \new_[30760]_ , \new_[30764]_ , \new_[30765]_ , \new_[30766]_ ,
    \new_[30770]_ , \new_[30771]_ , \new_[30775]_ , \new_[30776]_ ,
    \new_[30777]_ , \new_[30781]_ , \new_[30782]_ , \new_[30786]_ ,
    \new_[30787]_ , \new_[30788]_ , \new_[30792]_ , \new_[30793]_ ,
    \new_[30797]_ , \new_[30798]_ , \new_[30799]_ , \new_[30803]_ ,
    \new_[30804]_ , \new_[30808]_ , \new_[30809]_ , \new_[30810]_ ,
    \new_[30814]_ , \new_[30815]_ , \new_[30819]_ , \new_[30820]_ ,
    \new_[30821]_ , \new_[30825]_ , \new_[30826]_ , \new_[30830]_ ,
    \new_[30831]_ , \new_[30832]_ , \new_[30836]_ , \new_[30837]_ ,
    \new_[30841]_ , \new_[30842]_ , \new_[30843]_ , \new_[30847]_ ,
    \new_[30848]_ , \new_[30852]_ , \new_[30853]_ , \new_[30854]_ ,
    \new_[30858]_ , \new_[30859]_ , \new_[30863]_ , \new_[30864]_ ,
    \new_[30865]_ , \new_[30869]_ , \new_[30870]_ , \new_[30874]_ ,
    \new_[30875]_ , \new_[30876]_ , \new_[30880]_ , \new_[30881]_ ,
    \new_[30885]_ , \new_[30886]_ , \new_[30887]_ , \new_[30891]_ ,
    \new_[30892]_ , \new_[30896]_ , \new_[30897]_ , \new_[30898]_ ,
    \new_[30902]_ , \new_[30903]_ , \new_[30907]_ , \new_[30908]_ ,
    \new_[30909]_ , \new_[30913]_ , \new_[30914]_ , \new_[30918]_ ,
    \new_[30919]_ , \new_[30920]_ , \new_[30924]_ , \new_[30925]_ ,
    \new_[30929]_ , \new_[30930]_ , \new_[30931]_ , \new_[30935]_ ,
    \new_[30936]_ , \new_[30940]_ , \new_[30941]_ , \new_[30942]_ ,
    \new_[30946]_ , \new_[30947]_ , \new_[30951]_ , \new_[30952]_ ,
    \new_[30953]_ , \new_[30957]_ , \new_[30958]_ , \new_[30962]_ ,
    \new_[30963]_ , \new_[30964]_ , \new_[30968]_ , \new_[30969]_ ,
    \new_[30973]_ , \new_[30974]_ , \new_[30975]_ , \new_[30979]_ ,
    \new_[30980]_ , \new_[30984]_ , \new_[30985]_ , \new_[30986]_ ,
    \new_[30990]_ , \new_[30991]_ , \new_[30995]_ , \new_[30996]_ ,
    \new_[30997]_ , \new_[31001]_ , \new_[31002]_ , \new_[31006]_ ,
    \new_[31007]_ , \new_[31008]_ , \new_[31012]_ , \new_[31013]_ ,
    \new_[31017]_ , \new_[31018]_ , \new_[31019]_ , \new_[31023]_ ,
    \new_[31024]_ , \new_[31028]_ , \new_[31029]_ , \new_[31030]_ ,
    \new_[31034]_ , \new_[31035]_ , \new_[31039]_ , \new_[31040]_ ,
    \new_[31041]_ , \new_[31045]_ , \new_[31046]_ , \new_[31050]_ ,
    \new_[31051]_ , \new_[31052]_ , \new_[31056]_ , \new_[31057]_ ,
    \new_[31061]_ , \new_[31062]_ , \new_[31063]_ , \new_[31067]_ ,
    \new_[31068]_ , \new_[31072]_ , \new_[31073]_ , \new_[31074]_ ,
    \new_[31078]_ , \new_[31079]_ , \new_[31083]_ , \new_[31084]_ ,
    \new_[31085]_ , \new_[31089]_ , \new_[31090]_ , \new_[31094]_ ,
    \new_[31095]_ , \new_[31096]_ , \new_[31100]_ , \new_[31101]_ ,
    \new_[31105]_ , \new_[31106]_ , \new_[31107]_ , \new_[31111]_ ,
    \new_[31112]_ , \new_[31116]_ , \new_[31117]_ , \new_[31118]_ ,
    \new_[31122]_ , \new_[31123]_ , \new_[31127]_ , \new_[31128]_ ,
    \new_[31129]_ , \new_[31133]_ , \new_[31134]_ , \new_[31138]_ ,
    \new_[31139]_ , \new_[31140]_ , \new_[31144]_ , \new_[31145]_ ,
    \new_[31149]_ , \new_[31150]_ , \new_[31151]_ , \new_[31155]_ ,
    \new_[31156]_ , \new_[31160]_ , \new_[31161]_ , \new_[31162]_ ,
    \new_[31166]_ , \new_[31167]_ , \new_[31171]_ , \new_[31172]_ ,
    \new_[31173]_ , \new_[31177]_ , \new_[31178]_ , \new_[31182]_ ,
    \new_[31183]_ , \new_[31184]_ , \new_[31188]_ , \new_[31189]_ ,
    \new_[31193]_ , \new_[31194]_ , \new_[31195]_ , \new_[31199]_ ,
    \new_[31200]_ , \new_[31204]_ , \new_[31205]_ , \new_[31206]_ ,
    \new_[31210]_ , \new_[31211]_ , \new_[31215]_ , \new_[31216]_ ,
    \new_[31217]_ , \new_[31221]_ , \new_[31222]_ , \new_[31226]_ ,
    \new_[31227]_ , \new_[31228]_ , \new_[31232]_ , \new_[31233]_ ,
    \new_[31237]_ , \new_[31238]_ , \new_[31239]_ , \new_[31243]_ ,
    \new_[31244]_ , \new_[31248]_ , \new_[31249]_ , \new_[31250]_ ,
    \new_[31254]_ , \new_[31255]_ , \new_[31259]_ , \new_[31260]_ ,
    \new_[31261]_ , \new_[31265]_ , \new_[31266]_ , \new_[31270]_ ,
    \new_[31271]_ , \new_[31272]_ , \new_[31276]_ , \new_[31277]_ ,
    \new_[31281]_ , \new_[31282]_ , \new_[31283]_ , \new_[31287]_ ,
    \new_[31288]_ , \new_[31292]_ , \new_[31293]_ , \new_[31294]_ ,
    \new_[31298]_ , \new_[31299]_ , \new_[31303]_ , \new_[31304]_ ,
    \new_[31305]_ , \new_[31309]_ , \new_[31310]_ , \new_[31314]_ ,
    \new_[31315]_ , \new_[31316]_ , \new_[31320]_ , \new_[31321]_ ,
    \new_[31325]_ , \new_[31326]_ , \new_[31327]_ , \new_[31331]_ ,
    \new_[31332]_ , \new_[31336]_ , \new_[31337]_ , \new_[31338]_ ,
    \new_[31342]_ , \new_[31343]_ , \new_[31347]_ , \new_[31348]_ ,
    \new_[31349]_ , \new_[31353]_ , \new_[31354]_ , \new_[31358]_ ,
    \new_[31359]_ , \new_[31360]_ , \new_[31364]_ , \new_[31365]_ ,
    \new_[31369]_ , \new_[31370]_ , \new_[31371]_ , \new_[31375]_ ,
    \new_[31376]_ , \new_[31380]_ , \new_[31381]_ , \new_[31382]_ ,
    \new_[31386]_ , \new_[31387]_ , \new_[31391]_ , \new_[31392]_ ,
    \new_[31393]_ , \new_[31397]_ , \new_[31398]_ , \new_[31402]_ ,
    \new_[31403]_ , \new_[31404]_ , \new_[31408]_ , \new_[31409]_ ,
    \new_[31413]_ , \new_[31414]_ , \new_[31415]_ , \new_[31419]_ ,
    \new_[31420]_ , \new_[31424]_ , \new_[31425]_ , \new_[31426]_ ,
    \new_[31430]_ , \new_[31431]_ , \new_[31435]_ , \new_[31436]_ ,
    \new_[31437]_ , \new_[31441]_ , \new_[31442]_ , \new_[31446]_ ,
    \new_[31447]_ , \new_[31448]_ , \new_[31452]_ , \new_[31453]_ ,
    \new_[31457]_ , \new_[31458]_ , \new_[31459]_ , \new_[31463]_ ,
    \new_[31464]_ , \new_[31468]_ , \new_[31469]_ , \new_[31470]_ ,
    \new_[31474]_ , \new_[31475]_ , \new_[31479]_ , \new_[31480]_ ,
    \new_[31481]_ , \new_[31485]_ , \new_[31486]_ , \new_[31490]_ ,
    \new_[31491]_ , \new_[31492]_ , \new_[31496]_ , \new_[31497]_ ,
    \new_[31501]_ , \new_[31502]_ , \new_[31503]_ , \new_[31507]_ ,
    \new_[31508]_ , \new_[31512]_ , \new_[31513]_ , \new_[31514]_ ,
    \new_[31518]_ , \new_[31519]_ , \new_[31523]_ , \new_[31524]_ ,
    \new_[31525]_ , \new_[31529]_ , \new_[31530]_ , \new_[31534]_ ,
    \new_[31535]_ , \new_[31536]_ , \new_[31540]_ , \new_[31541]_ ,
    \new_[31545]_ , \new_[31546]_ , \new_[31547]_ , \new_[31551]_ ,
    \new_[31552]_ , \new_[31556]_ , \new_[31557]_ , \new_[31558]_ ,
    \new_[31562]_ , \new_[31563]_ , \new_[31567]_ , \new_[31568]_ ,
    \new_[31569]_ , \new_[31573]_ , \new_[31574]_ , \new_[31578]_ ,
    \new_[31579]_ , \new_[31580]_ , \new_[31584]_ , \new_[31585]_ ,
    \new_[31589]_ , \new_[31590]_ , \new_[31591]_ , \new_[31595]_ ,
    \new_[31596]_ , \new_[31600]_ , \new_[31601]_ , \new_[31602]_ ,
    \new_[31606]_ , \new_[31607]_ , \new_[31611]_ , \new_[31612]_ ,
    \new_[31613]_ , \new_[31617]_ , \new_[31618]_ , \new_[31622]_ ,
    \new_[31623]_ , \new_[31624]_ , \new_[31628]_ , \new_[31629]_ ,
    \new_[31633]_ , \new_[31634]_ , \new_[31635]_ , \new_[31639]_ ,
    \new_[31640]_ , \new_[31644]_ , \new_[31645]_ , \new_[31646]_ ,
    \new_[31650]_ , \new_[31651]_ , \new_[31655]_ , \new_[31656]_ ,
    \new_[31657]_ , \new_[31661]_ , \new_[31662]_ , \new_[31666]_ ,
    \new_[31667]_ , \new_[31668]_ , \new_[31672]_ , \new_[31673]_ ,
    \new_[31677]_ , \new_[31678]_ , \new_[31679]_ , \new_[31683]_ ,
    \new_[31684]_ , \new_[31688]_ , \new_[31689]_ , \new_[31690]_ ,
    \new_[31694]_ , \new_[31695]_ , \new_[31699]_ , \new_[31700]_ ,
    \new_[31701]_ , \new_[31705]_ , \new_[31706]_ , \new_[31710]_ ,
    \new_[31711]_ , \new_[31712]_ , \new_[31716]_ , \new_[31717]_ ,
    \new_[31721]_ , \new_[31722]_ , \new_[31723]_ , \new_[31727]_ ,
    \new_[31728]_ , \new_[31732]_ , \new_[31733]_ , \new_[31734]_ ,
    \new_[31738]_ , \new_[31739]_ , \new_[31743]_ , \new_[31744]_ ,
    \new_[31745]_ , \new_[31749]_ , \new_[31750]_ , \new_[31754]_ ,
    \new_[31755]_ , \new_[31756]_ , \new_[31760]_ , \new_[31761]_ ,
    \new_[31765]_ , \new_[31766]_ , \new_[31767]_ , \new_[31771]_ ,
    \new_[31772]_ , \new_[31776]_ , \new_[31777]_ , \new_[31778]_ ,
    \new_[31782]_ , \new_[31783]_ , \new_[31787]_ , \new_[31788]_ ,
    \new_[31789]_ , \new_[31793]_ , \new_[31794]_ , \new_[31798]_ ,
    \new_[31799]_ , \new_[31800]_ , \new_[31804]_ , \new_[31805]_ ,
    \new_[31809]_ , \new_[31810]_ , \new_[31811]_ , \new_[31815]_ ,
    \new_[31816]_ , \new_[31820]_ , \new_[31821]_ , \new_[31822]_ ,
    \new_[31826]_ , \new_[31827]_ , \new_[31831]_ , \new_[31832]_ ,
    \new_[31833]_ , \new_[31837]_ , \new_[31838]_ , \new_[31842]_ ,
    \new_[31843]_ , \new_[31844]_ , \new_[31848]_ , \new_[31849]_ ,
    \new_[31853]_ , \new_[31854]_ , \new_[31855]_ , \new_[31859]_ ,
    \new_[31860]_ , \new_[31864]_ , \new_[31865]_ , \new_[31866]_ ,
    \new_[31870]_ , \new_[31871]_ , \new_[31875]_ , \new_[31876]_ ,
    \new_[31877]_ , \new_[31881]_ , \new_[31882]_ , \new_[31886]_ ,
    \new_[31887]_ , \new_[31888]_ , \new_[31892]_ , \new_[31893]_ ,
    \new_[31897]_ , \new_[31898]_ , \new_[31899]_ , \new_[31903]_ ,
    \new_[31904]_ , \new_[31908]_ , \new_[31909]_ , \new_[31910]_ ,
    \new_[31914]_ , \new_[31915]_ , \new_[31919]_ , \new_[31920]_ ,
    \new_[31921]_ , \new_[31925]_ , \new_[31926]_ , \new_[31930]_ ,
    \new_[31931]_ , \new_[31932]_ , \new_[31936]_ , \new_[31937]_ ,
    \new_[31941]_ , \new_[31942]_ , \new_[31943]_ , \new_[31947]_ ,
    \new_[31948]_ , \new_[31952]_ , \new_[31953]_ , \new_[31954]_ ,
    \new_[31958]_ , \new_[31959]_ , \new_[31963]_ , \new_[31964]_ ,
    \new_[31965]_ , \new_[31969]_ , \new_[31970]_ , \new_[31974]_ ,
    \new_[31975]_ , \new_[31976]_ , \new_[31980]_ , \new_[31981]_ ,
    \new_[31985]_ , \new_[31986]_ , \new_[31987]_ , \new_[31991]_ ,
    \new_[31992]_ , \new_[31996]_ , \new_[31997]_ , \new_[31998]_ ,
    \new_[32002]_ , \new_[32003]_ , \new_[32007]_ , \new_[32008]_ ,
    \new_[32009]_ , \new_[32013]_ , \new_[32014]_ , \new_[32018]_ ,
    \new_[32019]_ , \new_[32020]_ , \new_[32024]_ , \new_[32025]_ ,
    \new_[32029]_ , \new_[32030]_ , \new_[32031]_ , \new_[32035]_ ,
    \new_[32036]_ , \new_[32040]_ , \new_[32041]_ , \new_[32042]_ ,
    \new_[32046]_ , \new_[32047]_ , \new_[32051]_ , \new_[32052]_ ,
    \new_[32053]_ , \new_[32057]_ , \new_[32058]_ , \new_[32062]_ ,
    \new_[32063]_ , \new_[32064]_ , \new_[32068]_ , \new_[32069]_ ,
    \new_[32073]_ , \new_[32074]_ , \new_[32075]_ , \new_[32079]_ ,
    \new_[32080]_ , \new_[32084]_ , \new_[32085]_ , \new_[32086]_ ,
    \new_[32090]_ , \new_[32091]_ , \new_[32095]_ , \new_[32096]_ ,
    \new_[32097]_ , \new_[32101]_ , \new_[32102]_ , \new_[32106]_ ,
    \new_[32107]_ , \new_[32108]_ , \new_[32112]_ , \new_[32113]_ ,
    \new_[32117]_ , \new_[32118]_ , \new_[32119]_ , \new_[32123]_ ,
    \new_[32124]_ , \new_[32128]_ , \new_[32129]_ , \new_[32130]_ ,
    \new_[32134]_ , \new_[32135]_ , \new_[32139]_ , \new_[32140]_ ,
    \new_[32141]_ , \new_[32145]_ , \new_[32146]_ , \new_[32150]_ ,
    \new_[32151]_ , \new_[32152]_ , \new_[32156]_ , \new_[32157]_ ,
    \new_[32161]_ , \new_[32162]_ , \new_[32163]_ , \new_[32167]_ ,
    \new_[32168]_ , \new_[32172]_ , \new_[32173]_ , \new_[32174]_ ,
    \new_[32178]_ , \new_[32179]_ , \new_[32183]_ , \new_[32184]_ ,
    \new_[32185]_ , \new_[32189]_ , \new_[32190]_ , \new_[32194]_ ,
    \new_[32195]_ , \new_[32196]_ , \new_[32200]_ , \new_[32201]_ ,
    \new_[32205]_ , \new_[32206]_ , \new_[32207]_ , \new_[32211]_ ,
    \new_[32212]_ , \new_[32216]_ , \new_[32217]_ , \new_[32218]_ ,
    \new_[32222]_ , \new_[32223]_ , \new_[32227]_ , \new_[32228]_ ,
    \new_[32229]_ , \new_[32233]_ , \new_[32234]_ , \new_[32238]_ ,
    \new_[32239]_ , \new_[32240]_ , \new_[32244]_ , \new_[32245]_ ,
    \new_[32249]_ , \new_[32250]_ , \new_[32251]_ , \new_[32255]_ ,
    \new_[32256]_ , \new_[32260]_ , \new_[32261]_ , \new_[32262]_ ,
    \new_[32266]_ , \new_[32267]_ , \new_[32271]_ , \new_[32272]_ ,
    \new_[32273]_ , \new_[32277]_ , \new_[32278]_ , \new_[32282]_ ,
    \new_[32283]_ , \new_[32284]_ , \new_[32288]_ , \new_[32289]_ ,
    \new_[32293]_ , \new_[32294]_ , \new_[32295]_ , \new_[32299]_ ,
    \new_[32300]_ , \new_[32304]_ , \new_[32305]_ , \new_[32306]_ ,
    \new_[32310]_ , \new_[32311]_ , \new_[32315]_ , \new_[32316]_ ,
    \new_[32317]_ , \new_[32321]_ , \new_[32322]_ , \new_[32326]_ ,
    \new_[32327]_ , \new_[32328]_ , \new_[32332]_ , \new_[32333]_ ,
    \new_[32337]_ , \new_[32338]_ , \new_[32339]_ , \new_[32343]_ ,
    \new_[32344]_ , \new_[32348]_ , \new_[32349]_ , \new_[32350]_ ,
    \new_[32354]_ , \new_[32355]_ , \new_[32359]_ , \new_[32360]_ ,
    \new_[32361]_ , \new_[32365]_ , \new_[32366]_ , \new_[32370]_ ,
    \new_[32371]_ , \new_[32372]_ , \new_[32376]_ , \new_[32377]_ ,
    \new_[32381]_ , \new_[32382]_ , \new_[32383]_ , \new_[32387]_ ,
    \new_[32388]_ , \new_[32392]_ , \new_[32393]_ , \new_[32394]_ ,
    \new_[32398]_ , \new_[32399]_ , \new_[32403]_ , \new_[32404]_ ,
    \new_[32405]_ , \new_[32409]_ , \new_[32410]_ , \new_[32414]_ ,
    \new_[32415]_ , \new_[32416]_ , \new_[32420]_ , \new_[32421]_ ,
    \new_[32425]_ , \new_[32426]_ , \new_[32427]_ , \new_[32431]_ ,
    \new_[32432]_ , \new_[32436]_ , \new_[32437]_ , \new_[32438]_ ,
    \new_[32442]_ , \new_[32443]_ , \new_[32447]_ , \new_[32448]_ ,
    \new_[32449]_ , \new_[32453]_ , \new_[32454]_ , \new_[32458]_ ,
    \new_[32459]_ , \new_[32460]_ , \new_[32464]_ , \new_[32465]_ ,
    \new_[32469]_ , \new_[32470]_ , \new_[32471]_ , \new_[32475]_ ,
    \new_[32476]_ , \new_[32480]_ , \new_[32481]_ , \new_[32482]_ ,
    \new_[32486]_ , \new_[32487]_ , \new_[32491]_ , \new_[32492]_ ,
    \new_[32493]_ , \new_[32497]_ , \new_[32498]_ , \new_[32502]_ ,
    \new_[32503]_ , \new_[32504]_ , \new_[32508]_ , \new_[32509]_ ,
    \new_[32513]_ , \new_[32514]_ , \new_[32515]_ , \new_[32519]_ ,
    \new_[32520]_ , \new_[32524]_ , \new_[32525]_ , \new_[32526]_ ,
    \new_[32530]_ , \new_[32531]_ , \new_[32535]_ , \new_[32536]_ ,
    \new_[32537]_ , \new_[32541]_ , \new_[32542]_ , \new_[32546]_ ,
    \new_[32547]_ , \new_[32548]_ , \new_[32552]_ , \new_[32553]_ ,
    \new_[32557]_ , \new_[32558]_ , \new_[32559]_ , \new_[32563]_ ,
    \new_[32564]_ , \new_[32568]_ , \new_[32569]_ , \new_[32570]_ ,
    \new_[32574]_ , \new_[32575]_ , \new_[32579]_ , \new_[32580]_ ,
    \new_[32581]_ , \new_[32585]_ , \new_[32586]_ , \new_[32590]_ ,
    \new_[32591]_ , \new_[32592]_ , \new_[32596]_ , \new_[32597]_ ,
    \new_[32601]_ , \new_[32602]_ , \new_[32603]_ , \new_[32607]_ ,
    \new_[32608]_ , \new_[32612]_ , \new_[32613]_ , \new_[32614]_ ,
    \new_[32618]_ , \new_[32619]_ , \new_[32623]_ , \new_[32624]_ ,
    \new_[32625]_ , \new_[32629]_ , \new_[32630]_ , \new_[32634]_ ,
    \new_[32635]_ , \new_[32636]_ , \new_[32640]_ , \new_[32641]_ ,
    \new_[32645]_ , \new_[32646]_ , \new_[32647]_ , \new_[32651]_ ,
    \new_[32652]_ , \new_[32656]_ , \new_[32657]_ , \new_[32658]_ ,
    \new_[32662]_ , \new_[32663]_ , \new_[32667]_ , \new_[32668]_ ,
    \new_[32669]_ , \new_[32673]_ , \new_[32674]_ , \new_[32678]_ ,
    \new_[32679]_ , \new_[32680]_ , \new_[32684]_ , \new_[32685]_ ,
    \new_[32689]_ , \new_[32690]_ , \new_[32691]_ , \new_[32695]_ ,
    \new_[32696]_ , \new_[32700]_ , \new_[32701]_ , \new_[32702]_ ,
    \new_[32706]_ , \new_[32707]_ , \new_[32711]_ , \new_[32712]_ ,
    \new_[32713]_ , \new_[32717]_ , \new_[32718]_ , \new_[32722]_ ,
    \new_[32723]_ , \new_[32724]_ , \new_[32728]_ , \new_[32729]_ ,
    \new_[32733]_ , \new_[32734]_ , \new_[32735]_ , \new_[32739]_ ,
    \new_[32740]_ , \new_[32744]_ , \new_[32745]_ , \new_[32746]_ ,
    \new_[32750]_ , \new_[32751]_ , \new_[32755]_ , \new_[32756]_ ,
    \new_[32757]_ , \new_[32761]_ , \new_[32762]_ , \new_[32766]_ ,
    \new_[32767]_ , \new_[32768]_ , \new_[32772]_ , \new_[32773]_ ,
    \new_[32777]_ , \new_[32778]_ , \new_[32779]_ , \new_[32783]_ ,
    \new_[32784]_ , \new_[32788]_ , \new_[32789]_ , \new_[32790]_ ,
    \new_[32794]_ , \new_[32795]_ , \new_[32799]_ , \new_[32800]_ ,
    \new_[32801]_ , \new_[32805]_ , \new_[32806]_ , \new_[32810]_ ,
    \new_[32811]_ , \new_[32812]_ , \new_[32816]_ , \new_[32817]_ ,
    \new_[32821]_ , \new_[32822]_ , \new_[32823]_ , \new_[32827]_ ,
    \new_[32828]_ , \new_[32832]_ , \new_[32833]_ , \new_[32834]_ ,
    \new_[32838]_ , \new_[32839]_ , \new_[32843]_ , \new_[32844]_ ,
    \new_[32845]_ , \new_[32849]_ , \new_[32850]_ , \new_[32854]_ ,
    \new_[32855]_ , \new_[32856]_ , \new_[32860]_ , \new_[32861]_ ,
    \new_[32865]_ , \new_[32866]_ , \new_[32867]_ , \new_[32871]_ ,
    \new_[32872]_ , \new_[32876]_ , \new_[32877]_ , \new_[32878]_ ,
    \new_[32882]_ , \new_[32883]_ , \new_[32887]_ , \new_[32888]_ ,
    \new_[32889]_ , \new_[32893]_ , \new_[32894]_ , \new_[32898]_ ,
    \new_[32899]_ , \new_[32900]_ , \new_[32904]_ , \new_[32905]_ ,
    \new_[32909]_ , \new_[32910]_ , \new_[32911]_ , \new_[32915]_ ,
    \new_[32916]_ , \new_[32920]_ , \new_[32921]_ , \new_[32922]_ ,
    \new_[32926]_ , \new_[32927]_ , \new_[32931]_ , \new_[32932]_ ,
    \new_[32933]_ , \new_[32937]_ , \new_[32938]_ , \new_[32942]_ ,
    \new_[32943]_ , \new_[32944]_ , \new_[32948]_ , \new_[32949]_ ,
    \new_[32953]_ , \new_[32954]_ , \new_[32955]_ , \new_[32959]_ ,
    \new_[32960]_ , \new_[32964]_ , \new_[32965]_ , \new_[32966]_ ,
    \new_[32970]_ , \new_[32971]_ , \new_[32975]_ , \new_[32976]_ ,
    \new_[32977]_ , \new_[32981]_ , \new_[32982]_ , \new_[32986]_ ,
    \new_[32987]_ , \new_[32988]_ , \new_[32992]_ , \new_[32993]_ ,
    \new_[32997]_ , \new_[32998]_ , \new_[32999]_ , \new_[33003]_ ,
    \new_[33004]_ , \new_[33008]_ , \new_[33009]_ , \new_[33010]_ ,
    \new_[33014]_ , \new_[33015]_ , \new_[33019]_ , \new_[33020]_ ,
    \new_[33021]_ , \new_[33025]_ , \new_[33026]_ , \new_[33030]_ ,
    \new_[33031]_ , \new_[33032]_ , \new_[33036]_ , \new_[33037]_ ,
    \new_[33041]_ , \new_[33042]_ , \new_[33043]_ , \new_[33047]_ ,
    \new_[33048]_ , \new_[33052]_ , \new_[33053]_ , \new_[33054]_ ,
    \new_[33058]_ , \new_[33059]_ , \new_[33063]_ , \new_[33064]_ ,
    \new_[33065]_ , \new_[33069]_ , \new_[33070]_ , \new_[33074]_ ,
    \new_[33075]_ , \new_[33076]_ , \new_[33080]_ , \new_[33081]_ ,
    \new_[33085]_ , \new_[33086]_ , \new_[33087]_ , \new_[33091]_ ,
    \new_[33092]_ , \new_[33096]_ , \new_[33097]_ , \new_[33098]_ ,
    \new_[33102]_ , \new_[33103]_ , \new_[33107]_ , \new_[33108]_ ,
    \new_[33109]_ , \new_[33113]_ , \new_[33114]_ , \new_[33118]_ ,
    \new_[33119]_ , \new_[33120]_ , \new_[33124]_ , \new_[33125]_ ,
    \new_[33129]_ , \new_[33130]_ , \new_[33131]_ , \new_[33135]_ ,
    \new_[33136]_ , \new_[33140]_ , \new_[33141]_ , \new_[33142]_ ,
    \new_[33146]_ , \new_[33147]_ , \new_[33151]_ , \new_[33152]_ ,
    \new_[33153]_ , \new_[33157]_ , \new_[33158]_ , \new_[33162]_ ,
    \new_[33163]_ , \new_[33164]_ , \new_[33168]_ , \new_[33169]_ ,
    \new_[33173]_ , \new_[33174]_ , \new_[33175]_ , \new_[33179]_ ,
    \new_[33180]_ , \new_[33184]_ , \new_[33185]_ , \new_[33186]_ ,
    \new_[33190]_ , \new_[33191]_ , \new_[33195]_ , \new_[33196]_ ,
    \new_[33197]_ , \new_[33201]_ , \new_[33202]_ , \new_[33206]_ ,
    \new_[33207]_ , \new_[33208]_ , \new_[33212]_ , \new_[33213]_ ,
    \new_[33217]_ , \new_[33218]_ , \new_[33219]_ , \new_[33223]_ ,
    \new_[33224]_ , \new_[33228]_ , \new_[33229]_ , \new_[33230]_ ,
    \new_[33234]_ , \new_[33235]_ , \new_[33239]_ , \new_[33240]_ ,
    \new_[33241]_ , \new_[33245]_ , \new_[33246]_ , \new_[33250]_ ,
    \new_[33251]_ , \new_[33252]_ , \new_[33256]_ , \new_[33257]_ ,
    \new_[33261]_ , \new_[33262]_ , \new_[33263]_ , \new_[33267]_ ,
    \new_[33268]_ , \new_[33272]_ , \new_[33273]_ , \new_[33274]_ ,
    \new_[33278]_ , \new_[33279]_ , \new_[33283]_ , \new_[33284]_ ,
    \new_[33285]_ , \new_[33289]_ , \new_[33290]_ , \new_[33294]_ ,
    \new_[33295]_ , \new_[33296]_ , \new_[33300]_ , \new_[33301]_ ,
    \new_[33305]_ , \new_[33306]_ , \new_[33307]_ , \new_[33311]_ ,
    \new_[33312]_ , \new_[33316]_ , \new_[33317]_ , \new_[33318]_ ,
    \new_[33322]_ , \new_[33323]_ , \new_[33327]_ , \new_[33328]_ ,
    \new_[33329]_ , \new_[33333]_ , \new_[33334]_ , \new_[33338]_ ,
    \new_[33339]_ , \new_[33340]_ , \new_[33344]_ , \new_[33345]_ ,
    \new_[33349]_ , \new_[33350]_ , \new_[33351]_ , \new_[33355]_ ,
    \new_[33356]_ , \new_[33360]_ , \new_[33361]_ , \new_[33362]_ ,
    \new_[33366]_ , \new_[33367]_ , \new_[33371]_ , \new_[33372]_ ,
    \new_[33373]_ , \new_[33377]_ , \new_[33378]_ , \new_[33382]_ ,
    \new_[33383]_ , \new_[33384]_ , \new_[33388]_ , \new_[33389]_ ,
    \new_[33393]_ , \new_[33394]_ , \new_[33395]_ , \new_[33399]_ ,
    \new_[33400]_ , \new_[33404]_ , \new_[33405]_ , \new_[33406]_ ,
    \new_[33410]_ , \new_[33411]_ , \new_[33415]_ , \new_[33416]_ ,
    \new_[33417]_ , \new_[33421]_ , \new_[33422]_ , \new_[33426]_ ,
    \new_[33427]_ , \new_[33428]_ , \new_[33432]_ , \new_[33433]_ ,
    \new_[33437]_ , \new_[33438]_ , \new_[33439]_ , \new_[33443]_ ,
    \new_[33444]_ , \new_[33448]_ , \new_[33449]_ , \new_[33450]_ ,
    \new_[33454]_ , \new_[33455]_ , \new_[33459]_ , \new_[33460]_ ,
    \new_[33461]_ , \new_[33465]_ , \new_[33466]_ , \new_[33470]_ ,
    \new_[33471]_ , \new_[33472]_ , \new_[33476]_ , \new_[33477]_ ,
    \new_[33481]_ , \new_[33482]_ , \new_[33483]_ , \new_[33487]_ ,
    \new_[33488]_ , \new_[33492]_ , \new_[33493]_ , \new_[33494]_ ,
    \new_[33498]_ , \new_[33499]_ , \new_[33503]_ , \new_[33504]_ ,
    \new_[33505]_ , \new_[33509]_ , \new_[33510]_ , \new_[33514]_ ,
    \new_[33515]_ , \new_[33516]_ , \new_[33520]_ , \new_[33521]_ ,
    \new_[33525]_ , \new_[33526]_ , \new_[33527]_ , \new_[33531]_ ,
    \new_[33532]_ , \new_[33536]_ , \new_[33537]_ , \new_[33538]_ ,
    \new_[33542]_ , \new_[33543]_ , \new_[33547]_ , \new_[33548]_ ,
    \new_[33549]_ , \new_[33553]_ , \new_[33554]_ , \new_[33558]_ ,
    \new_[33559]_ , \new_[33560]_ , \new_[33564]_ , \new_[33565]_ ,
    \new_[33569]_ , \new_[33570]_ , \new_[33571]_ , \new_[33575]_ ,
    \new_[33576]_ , \new_[33580]_ , \new_[33581]_ , \new_[33582]_ ,
    \new_[33586]_ , \new_[33587]_ , \new_[33591]_ , \new_[33592]_ ,
    \new_[33593]_ , \new_[33597]_ , \new_[33598]_ , \new_[33602]_ ,
    \new_[33603]_ , \new_[33604]_ , \new_[33608]_ , \new_[33609]_ ,
    \new_[33613]_ , \new_[33614]_ , \new_[33615]_ , \new_[33619]_ ,
    \new_[33620]_ , \new_[33624]_ , \new_[33625]_ , \new_[33626]_ ,
    \new_[33630]_ , \new_[33631]_ , \new_[33635]_ , \new_[33636]_ ,
    \new_[33637]_ , \new_[33641]_ , \new_[33642]_ , \new_[33646]_ ,
    \new_[33647]_ , \new_[33648]_ , \new_[33652]_ , \new_[33653]_ ,
    \new_[33657]_ , \new_[33658]_ , \new_[33659]_ , \new_[33663]_ ,
    \new_[33664]_ , \new_[33668]_ , \new_[33669]_ , \new_[33670]_ ,
    \new_[33674]_ , \new_[33675]_ , \new_[33679]_ , \new_[33680]_ ,
    \new_[33681]_ , \new_[33685]_ , \new_[33686]_ , \new_[33690]_ ,
    \new_[33691]_ , \new_[33692]_ , \new_[33696]_ , \new_[33697]_ ,
    \new_[33701]_ , \new_[33702]_ , \new_[33703]_ , \new_[33707]_ ,
    \new_[33708]_ , \new_[33712]_ , \new_[33713]_ , \new_[33714]_ ,
    \new_[33718]_ , \new_[33719]_ , \new_[33723]_ , \new_[33724]_ ,
    \new_[33725]_ , \new_[33729]_ , \new_[33730]_ , \new_[33734]_ ,
    \new_[33735]_ , \new_[33736]_ , \new_[33740]_ , \new_[33741]_ ,
    \new_[33745]_ , \new_[33746]_ , \new_[33747]_ , \new_[33751]_ ,
    \new_[33752]_ , \new_[33756]_ , \new_[33757]_ , \new_[33758]_ ,
    \new_[33762]_ , \new_[33763]_ , \new_[33767]_ , \new_[33768]_ ,
    \new_[33769]_ , \new_[33773]_ , \new_[33774]_ , \new_[33778]_ ,
    \new_[33779]_ , \new_[33780]_ , \new_[33784]_ , \new_[33785]_ ,
    \new_[33789]_ , \new_[33790]_ , \new_[33791]_ , \new_[33795]_ ,
    \new_[33796]_ , \new_[33800]_ , \new_[33801]_ , \new_[33802]_ ,
    \new_[33806]_ , \new_[33807]_ , \new_[33811]_ , \new_[33812]_ ,
    \new_[33813]_ , \new_[33817]_ , \new_[33818]_ , \new_[33822]_ ,
    \new_[33823]_ , \new_[33824]_ , \new_[33828]_ , \new_[33829]_ ,
    \new_[33833]_ , \new_[33834]_ , \new_[33835]_ , \new_[33839]_ ,
    \new_[33840]_ , \new_[33844]_ , \new_[33845]_ , \new_[33846]_ ,
    \new_[33850]_ , \new_[33851]_ , \new_[33855]_ , \new_[33856]_ ,
    \new_[33857]_ , \new_[33861]_ , \new_[33862]_ , \new_[33866]_ ,
    \new_[33867]_ , \new_[33868]_ , \new_[33872]_ , \new_[33873]_ ,
    \new_[33877]_ , \new_[33878]_ , \new_[33879]_ , \new_[33883]_ ,
    \new_[33884]_ , \new_[33888]_ , \new_[33889]_ , \new_[33890]_ ,
    \new_[33894]_ , \new_[33895]_ , \new_[33899]_ , \new_[33900]_ ,
    \new_[33901]_ , \new_[33905]_ , \new_[33906]_ , \new_[33910]_ ,
    \new_[33911]_ , \new_[33912]_ , \new_[33916]_ , \new_[33917]_ ,
    \new_[33921]_ , \new_[33922]_ , \new_[33923]_ , \new_[33927]_ ,
    \new_[33928]_ , \new_[33932]_ , \new_[33933]_ , \new_[33934]_ ,
    \new_[33938]_ , \new_[33939]_ , \new_[33943]_ , \new_[33944]_ ,
    \new_[33945]_ , \new_[33949]_ , \new_[33950]_ , \new_[33954]_ ,
    \new_[33955]_ , \new_[33956]_ , \new_[33960]_ , \new_[33961]_ ,
    \new_[33965]_ , \new_[33966]_ , \new_[33967]_ , \new_[33971]_ ,
    \new_[33972]_ , \new_[33976]_ , \new_[33977]_ , \new_[33978]_ ,
    \new_[33982]_ , \new_[33983]_ , \new_[33987]_ , \new_[33988]_ ,
    \new_[33989]_ , \new_[33993]_ , \new_[33994]_ , \new_[33998]_ ,
    \new_[33999]_ , \new_[34000]_ , \new_[34004]_ , \new_[34005]_ ,
    \new_[34009]_ , \new_[34010]_ , \new_[34011]_ , \new_[34015]_ ,
    \new_[34016]_ , \new_[34020]_ , \new_[34021]_ , \new_[34022]_ ,
    \new_[34026]_ , \new_[34027]_ , \new_[34031]_ , \new_[34032]_ ,
    \new_[34033]_ , \new_[34037]_ , \new_[34038]_ , \new_[34042]_ ,
    \new_[34043]_ , \new_[34044]_ , \new_[34048]_ , \new_[34049]_ ,
    \new_[34053]_ , \new_[34054]_ , \new_[34055]_ , \new_[34059]_ ,
    \new_[34060]_ , \new_[34064]_ , \new_[34065]_ , \new_[34066]_ ,
    \new_[34070]_ , \new_[34071]_ , \new_[34075]_ , \new_[34076]_ ,
    \new_[34077]_ , \new_[34081]_ , \new_[34082]_ , \new_[34086]_ ,
    \new_[34087]_ , \new_[34088]_ , \new_[34092]_ , \new_[34093]_ ,
    \new_[34097]_ , \new_[34098]_ , \new_[34099]_ , \new_[34103]_ ,
    \new_[34104]_ , \new_[34108]_ , \new_[34109]_ , \new_[34110]_ ,
    \new_[34114]_ , \new_[34115]_ , \new_[34119]_ , \new_[34120]_ ,
    \new_[34121]_ , \new_[34125]_ , \new_[34126]_ , \new_[34130]_ ,
    \new_[34131]_ , \new_[34132]_ , \new_[34136]_ , \new_[34137]_ ,
    \new_[34141]_ , \new_[34142]_ , \new_[34143]_ , \new_[34147]_ ,
    \new_[34148]_ , \new_[34152]_ , \new_[34153]_ , \new_[34154]_ ,
    \new_[34158]_ , \new_[34159]_ , \new_[34163]_ , \new_[34164]_ ,
    \new_[34165]_ , \new_[34169]_ , \new_[34170]_ , \new_[34174]_ ,
    \new_[34175]_ , \new_[34176]_ , \new_[34180]_ , \new_[34181]_ ,
    \new_[34185]_ , \new_[34186]_ , \new_[34187]_ , \new_[34191]_ ,
    \new_[34192]_ , \new_[34196]_ , \new_[34197]_ , \new_[34198]_ ,
    \new_[34202]_ , \new_[34203]_ , \new_[34207]_ , \new_[34208]_ ,
    \new_[34209]_ , \new_[34213]_ , \new_[34214]_ , \new_[34218]_ ,
    \new_[34219]_ , \new_[34220]_ , \new_[34224]_ , \new_[34225]_ ,
    \new_[34229]_ , \new_[34230]_ , \new_[34231]_ , \new_[34235]_ ,
    \new_[34236]_ , \new_[34240]_ , \new_[34241]_ , \new_[34242]_ ,
    \new_[34246]_ , \new_[34247]_ , \new_[34251]_ , \new_[34252]_ ,
    \new_[34253]_ , \new_[34257]_ , \new_[34258]_ , \new_[34262]_ ,
    \new_[34263]_ , \new_[34264]_ , \new_[34268]_ , \new_[34269]_ ,
    \new_[34273]_ , \new_[34274]_ , \new_[34275]_ , \new_[34279]_ ,
    \new_[34280]_ , \new_[34284]_ , \new_[34285]_ , \new_[34286]_ ,
    \new_[34290]_ , \new_[34291]_ , \new_[34295]_ , \new_[34296]_ ,
    \new_[34297]_ , \new_[34301]_ , \new_[34302]_ , \new_[34306]_ ,
    \new_[34307]_ , \new_[34308]_ , \new_[34312]_ , \new_[34313]_ ,
    \new_[34317]_ , \new_[34318]_ , \new_[34319]_ , \new_[34323]_ ,
    \new_[34324]_ , \new_[34328]_ , \new_[34329]_ , \new_[34330]_ ,
    \new_[34334]_ , \new_[34335]_ , \new_[34339]_ , \new_[34340]_ ,
    \new_[34341]_ , \new_[34345]_ , \new_[34346]_ , \new_[34350]_ ,
    \new_[34351]_ , \new_[34352]_ , \new_[34356]_ , \new_[34357]_ ,
    \new_[34361]_ , \new_[34362]_ , \new_[34363]_ , \new_[34367]_ ,
    \new_[34368]_ , \new_[34372]_ , \new_[34373]_ , \new_[34374]_ ,
    \new_[34378]_ , \new_[34379]_ , \new_[34383]_ , \new_[34384]_ ,
    \new_[34385]_ , \new_[34389]_ , \new_[34390]_ , \new_[34394]_ ,
    \new_[34395]_ , \new_[34396]_ , \new_[34400]_ , \new_[34401]_ ,
    \new_[34405]_ , \new_[34406]_ , \new_[34407]_ , \new_[34411]_ ,
    \new_[34412]_ , \new_[34416]_ , \new_[34417]_ , \new_[34418]_ ,
    \new_[34422]_ , \new_[34423]_ , \new_[34427]_ , \new_[34428]_ ,
    \new_[34429]_ , \new_[34433]_ , \new_[34434]_ , \new_[34438]_ ,
    \new_[34439]_ , \new_[34440]_ , \new_[34444]_ , \new_[34445]_ ,
    \new_[34449]_ , \new_[34450]_ , \new_[34451]_ , \new_[34455]_ ,
    \new_[34456]_ , \new_[34460]_ , \new_[34461]_ , \new_[34462]_ ,
    \new_[34466]_ , \new_[34467]_ , \new_[34471]_ , \new_[34472]_ ,
    \new_[34473]_ , \new_[34477]_ , \new_[34478]_ , \new_[34482]_ ,
    \new_[34483]_ , \new_[34484]_ , \new_[34488]_ , \new_[34489]_ ,
    \new_[34493]_ , \new_[34494]_ , \new_[34495]_ , \new_[34499]_ ,
    \new_[34500]_ , \new_[34504]_ , \new_[34505]_ , \new_[34506]_ ,
    \new_[34510]_ , \new_[34511]_ , \new_[34515]_ , \new_[34516]_ ,
    \new_[34517]_ , \new_[34521]_ , \new_[34522]_ , \new_[34526]_ ,
    \new_[34527]_ , \new_[34528]_ , \new_[34532]_ , \new_[34533]_ ,
    \new_[34537]_ , \new_[34538]_ , \new_[34539]_ , \new_[34543]_ ,
    \new_[34544]_ , \new_[34548]_ , \new_[34549]_ , \new_[34550]_ ,
    \new_[34554]_ , \new_[34555]_ , \new_[34559]_ , \new_[34560]_ ,
    \new_[34561]_ , \new_[34565]_ , \new_[34566]_ , \new_[34570]_ ,
    \new_[34571]_ , \new_[34572]_ , \new_[34576]_ , \new_[34577]_ ,
    \new_[34581]_ , \new_[34582]_ , \new_[34583]_ , \new_[34587]_ ,
    \new_[34588]_ , \new_[34592]_ , \new_[34593]_ , \new_[34594]_ ,
    \new_[34598]_ , \new_[34599]_ , \new_[34603]_ , \new_[34604]_ ,
    \new_[34605]_ , \new_[34609]_ , \new_[34610]_ , \new_[34614]_ ,
    \new_[34615]_ , \new_[34616]_ , \new_[34620]_ , \new_[34621]_ ,
    \new_[34625]_ , \new_[34626]_ , \new_[34627]_ , \new_[34631]_ ,
    \new_[34632]_ , \new_[34636]_ , \new_[34637]_ , \new_[34638]_ ,
    \new_[34642]_ , \new_[34643]_ , \new_[34647]_ , \new_[34648]_ ,
    \new_[34649]_ , \new_[34653]_ , \new_[34654]_ , \new_[34658]_ ,
    \new_[34659]_ , \new_[34660]_ , \new_[34664]_ , \new_[34665]_ ,
    \new_[34669]_ , \new_[34670]_ , \new_[34671]_ , \new_[34675]_ ,
    \new_[34676]_ , \new_[34680]_ , \new_[34681]_ , \new_[34682]_ ,
    \new_[34686]_ , \new_[34687]_ , \new_[34691]_ , \new_[34692]_ ,
    \new_[34693]_ , \new_[34697]_ , \new_[34698]_ , \new_[34702]_ ,
    \new_[34703]_ , \new_[34704]_ , \new_[34708]_ , \new_[34709]_ ,
    \new_[34713]_ , \new_[34714]_ , \new_[34715]_ , \new_[34719]_ ,
    \new_[34720]_ , \new_[34724]_ , \new_[34725]_ , \new_[34726]_ ,
    \new_[34730]_ , \new_[34731]_ , \new_[34735]_ , \new_[34736]_ ,
    \new_[34737]_ , \new_[34741]_ , \new_[34742]_ , \new_[34746]_ ,
    \new_[34747]_ , \new_[34748]_ , \new_[34752]_ , \new_[34753]_ ,
    \new_[34757]_ , \new_[34758]_ , \new_[34759]_ , \new_[34763]_ ,
    \new_[34764]_ , \new_[34768]_ , \new_[34769]_ , \new_[34770]_ ,
    \new_[34774]_ , \new_[34775]_ , \new_[34779]_ , \new_[34780]_ ,
    \new_[34781]_ , \new_[34785]_ , \new_[34786]_ , \new_[34790]_ ,
    \new_[34791]_ , \new_[34792]_ , \new_[34796]_ , \new_[34797]_ ,
    \new_[34801]_ , \new_[34802]_ , \new_[34803]_ , \new_[34807]_ ,
    \new_[34808]_ , \new_[34812]_ , \new_[34813]_ , \new_[34814]_ ,
    \new_[34818]_ , \new_[34819]_ , \new_[34823]_ , \new_[34824]_ ,
    \new_[34825]_ , \new_[34829]_ , \new_[34830]_ , \new_[34834]_ ,
    \new_[34835]_ , \new_[34836]_ , \new_[34840]_ , \new_[34841]_ ,
    \new_[34845]_ , \new_[34846]_ , \new_[34847]_ , \new_[34851]_ ,
    \new_[34852]_ , \new_[34856]_ , \new_[34857]_ , \new_[34858]_ ,
    \new_[34862]_ , \new_[34863]_ , \new_[34867]_ , \new_[34868]_ ,
    \new_[34869]_ , \new_[34873]_ , \new_[34874]_ , \new_[34878]_ ,
    \new_[34879]_ , \new_[34880]_ , \new_[34884]_ , \new_[34885]_ ,
    \new_[34889]_ , \new_[34890]_ , \new_[34891]_ , \new_[34895]_ ,
    \new_[34896]_ , \new_[34900]_ , \new_[34901]_ , \new_[34902]_ ,
    \new_[34906]_ , \new_[34907]_ , \new_[34911]_ , \new_[34912]_ ,
    \new_[34913]_ , \new_[34917]_ , \new_[34918]_ , \new_[34922]_ ,
    \new_[34923]_ , \new_[34924]_ , \new_[34928]_ , \new_[34929]_ ,
    \new_[34933]_ , \new_[34934]_ , \new_[34935]_ , \new_[34939]_ ,
    \new_[34940]_ , \new_[34944]_ , \new_[34945]_ , \new_[34946]_ ,
    \new_[34950]_ , \new_[34951]_ , \new_[34955]_ , \new_[34956]_ ,
    \new_[34957]_ , \new_[34961]_ , \new_[34962]_ , \new_[34966]_ ,
    \new_[34967]_ , \new_[34968]_ , \new_[34972]_ , \new_[34973]_ ,
    \new_[34977]_ , \new_[34978]_ , \new_[34979]_ , \new_[34983]_ ,
    \new_[34984]_ , \new_[34988]_ , \new_[34989]_ , \new_[34990]_ ,
    \new_[34994]_ , \new_[34995]_ , \new_[34999]_ , \new_[35000]_ ,
    \new_[35001]_ , \new_[35005]_ , \new_[35006]_ , \new_[35010]_ ,
    \new_[35011]_ , \new_[35012]_ , \new_[35016]_ , \new_[35017]_ ,
    \new_[35021]_ , \new_[35022]_ , \new_[35023]_ , \new_[35027]_ ,
    \new_[35028]_ , \new_[35032]_ , \new_[35033]_ , \new_[35034]_ ,
    \new_[35038]_ , \new_[35039]_ , \new_[35043]_ , \new_[35044]_ ,
    \new_[35045]_ , \new_[35049]_ , \new_[35050]_ , \new_[35054]_ ,
    \new_[35055]_ , \new_[35056]_ , \new_[35060]_ , \new_[35061]_ ,
    \new_[35065]_ , \new_[35066]_ , \new_[35067]_ , \new_[35071]_ ,
    \new_[35072]_ , \new_[35076]_ , \new_[35077]_ , \new_[35078]_ ,
    \new_[35082]_ , \new_[35083]_ , \new_[35087]_ , \new_[35088]_ ,
    \new_[35089]_ , \new_[35093]_ , \new_[35094]_ , \new_[35098]_ ,
    \new_[35099]_ , \new_[35100]_ , \new_[35104]_ , \new_[35105]_ ,
    \new_[35109]_ , \new_[35110]_ , \new_[35111]_ , \new_[35115]_ ,
    \new_[35116]_ , \new_[35120]_ , \new_[35121]_ , \new_[35122]_ ,
    \new_[35126]_ , \new_[35127]_ , \new_[35131]_ , \new_[35132]_ ,
    \new_[35133]_ , \new_[35137]_ , \new_[35138]_ , \new_[35142]_ ,
    \new_[35143]_ , \new_[35144]_ , \new_[35148]_ , \new_[35149]_ ,
    \new_[35153]_ , \new_[35154]_ , \new_[35155]_ , \new_[35159]_ ,
    \new_[35160]_ , \new_[35164]_ , \new_[35165]_ , \new_[35166]_ ,
    \new_[35170]_ , \new_[35171]_ , \new_[35175]_ , \new_[35176]_ ,
    \new_[35177]_ , \new_[35181]_ , \new_[35182]_ , \new_[35186]_ ,
    \new_[35187]_ , \new_[35188]_ , \new_[35192]_ , \new_[35193]_ ,
    \new_[35197]_ , \new_[35198]_ , \new_[35199]_ , \new_[35203]_ ,
    \new_[35204]_ , \new_[35208]_ , \new_[35209]_ , \new_[35210]_ ,
    \new_[35214]_ , \new_[35215]_ , \new_[35219]_ , \new_[35220]_ ,
    \new_[35221]_ , \new_[35225]_ , \new_[35226]_ , \new_[35230]_ ,
    \new_[35231]_ , \new_[35232]_ , \new_[35236]_ , \new_[35237]_ ,
    \new_[35241]_ , \new_[35242]_ , \new_[35243]_ , \new_[35247]_ ,
    \new_[35248]_ , \new_[35252]_ , \new_[35253]_ , \new_[35254]_ ,
    \new_[35258]_ , \new_[35259]_ , \new_[35263]_ , \new_[35264]_ ,
    \new_[35265]_ , \new_[35269]_ , \new_[35270]_ , \new_[35274]_ ,
    \new_[35275]_ , \new_[35276]_ , \new_[35280]_ , \new_[35281]_ ,
    \new_[35285]_ , \new_[35286]_ , \new_[35287]_ , \new_[35291]_ ,
    \new_[35292]_ , \new_[35296]_ , \new_[35297]_ , \new_[35298]_ ,
    \new_[35302]_ , \new_[35303]_ , \new_[35307]_ , \new_[35308]_ ,
    \new_[35309]_ , \new_[35313]_ , \new_[35314]_ , \new_[35318]_ ,
    \new_[35319]_ , \new_[35320]_ , \new_[35324]_ , \new_[35325]_ ,
    \new_[35329]_ , \new_[35330]_ , \new_[35331]_ , \new_[35335]_ ,
    \new_[35336]_ , \new_[35340]_ , \new_[35341]_ , \new_[35342]_ ,
    \new_[35346]_ , \new_[35347]_ , \new_[35351]_ , \new_[35352]_ ,
    \new_[35353]_ , \new_[35357]_ , \new_[35358]_ , \new_[35362]_ ,
    \new_[35363]_ , \new_[35364]_ , \new_[35368]_ , \new_[35369]_ ,
    \new_[35373]_ , \new_[35374]_ , \new_[35375]_ , \new_[35379]_ ,
    \new_[35380]_ , \new_[35384]_ , \new_[35385]_ , \new_[35386]_ ,
    \new_[35390]_ , \new_[35391]_ , \new_[35395]_ , \new_[35396]_ ,
    \new_[35397]_ , \new_[35401]_ , \new_[35402]_ , \new_[35406]_ ,
    \new_[35407]_ , \new_[35408]_ , \new_[35412]_ , \new_[35413]_ ,
    \new_[35417]_ , \new_[35418]_ , \new_[35419]_ , \new_[35423]_ ,
    \new_[35424]_ , \new_[35428]_ , \new_[35429]_ , \new_[35430]_ ,
    \new_[35434]_ , \new_[35435]_ , \new_[35439]_ , \new_[35440]_ ,
    \new_[35441]_ , \new_[35445]_ , \new_[35446]_ , \new_[35450]_ ,
    \new_[35451]_ , \new_[35452]_ , \new_[35456]_ , \new_[35457]_ ,
    \new_[35461]_ , \new_[35462]_ , \new_[35463]_ , \new_[35467]_ ,
    \new_[35468]_ , \new_[35472]_ , \new_[35473]_ , \new_[35474]_ ,
    \new_[35478]_ , \new_[35479]_ , \new_[35483]_ , \new_[35484]_ ,
    \new_[35485]_ , \new_[35489]_ , \new_[35490]_ , \new_[35494]_ ,
    \new_[35495]_ , \new_[35496]_ , \new_[35500]_ , \new_[35501]_ ,
    \new_[35505]_ , \new_[35506]_ , \new_[35507]_ , \new_[35511]_ ,
    \new_[35512]_ , \new_[35516]_ , \new_[35517]_ , \new_[35518]_ ,
    \new_[35522]_ , \new_[35523]_ , \new_[35527]_ , \new_[35528]_ ,
    \new_[35529]_ , \new_[35533]_ , \new_[35534]_ , \new_[35538]_ ,
    \new_[35539]_ , \new_[35540]_ , \new_[35544]_ , \new_[35545]_ ,
    \new_[35549]_ , \new_[35550]_ , \new_[35551]_ , \new_[35555]_ ,
    \new_[35556]_ , \new_[35560]_ , \new_[35561]_ , \new_[35562]_ ,
    \new_[35566]_ , \new_[35567]_ , \new_[35571]_ , \new_[35572]_ ,
    \new_[35573]_ , \new_[35577]_ , \new_[35578]_ , \new_[35582]_ ,
    \new_[35583]_ , \new_[35584]_ , \new_[35588]_ , \new_[35589]_ ,
    \new_[35593]_ , \new_[35594]_ , \new_[35595]_ , \new_[35599]_ ,
    \new_[35600]_ , \new_[35604]_ , \new_[35605]_ , \new_[35606]_ ,
    \new_[35610]_ , \new_[35611]_ , \new_[35615]_ , \new_[35616]_ ,
    \new_[35617]_ , \new_[35621]_ , \new_[35622]_ , \new_[35626]_ ,
    \new_[35627]_ , \new_[35628]_ , \new_[35632]_ , \new_[35633]_ ,
    \new_[35637]_ , \new_[35638]_ , \new_[35639]_ , \new_[35643]_ ,
    \new_[35644]_ , \new_[35648]_ , \new_[35649]_ , \new_[35650]_ ,
    \new_[35654]_ , \new_[35655]_ , \new_[35659]_ , \new_[35660]_ ,
    \new_[35661]_ , \new_[35665]_ , \new_[35666]_ , \new_[35670]_ ,
    \new_[35671]_ , \new_[35672]_ , \new_[35676]_ , \new_[35677]_ ,
    \new_[35681]_ , \new_[35682]_ , \new_[35683]_ , \new_[35687]_ ,
    \new_[35688]_ , \new_[35692]_ , \new_[35693]_ , \new_[35694]_ ,
    \new_[35698]_ , \new_[35699]_ , \new_[35703]_ , \new_[35704]_ ,
    \new_[35705]_ , \new_[35709]_ , \new_[35710]_ , \new_[35714]_ ,
    \new_[35715]_ , \new_[35716]_ , \new_[35720]_ , \new_[35721]_ ,
    \new_[35725]_ , \new_[35726]_ , \new_[35727]_ , \new_[35731]_ ,
    \new_[35732]_ , \new_[35736]_ , \new_[35737]_ , \new_[35738]_ ,
    \new_[35742]_ , \new_[35743]_ , \new_[35747]_ , \new_[35748]_ ,
    \new_[35749]_ , \new_[35753]_ , \new_[35754]_ , \new_[35758]_ ,
    \new_[35759]_ , \new_[35760]_ , \new_[35764]_ , \new_[35765]_ ,
    \new_[35769]_ , \new_[35770]_ , \new_[35771]_ , \new_[35775]_ ,
    \new_[35776]_ , \new_[35780]_ , \new_[35781]_ , \new_[35782]_ ,
    \new_[35786]_ , \new_[35787]_ , \new_[35791]_ , \new_[35792]_ ,
    \new_[35793]_ , \new_[35797]_ , \new_[35798]_ , \new_[35802]_ ,
    \new_[35803]_ , \new_[35804]_ , \new_[35808]_ , \new_[35809]_ ,
    \new_[35813]_ , \new_[35814]_ , \new_[35815]_ , \new_[35819]_ ,
    \new_[35820]_ , \new_[35824]_ , \new_[35825]_ , \new_[35826]_ ,
    \new_[35830]_ , \new_[35831]_ , \new_[35835]_ , \new_[35836]_ ,
    \new_[35837]_ , \new_[35841]_ , \new_[35842]_ , \new_[35846]_ ,
    \new_[35847]_ , \new_[35848]_ , \new_[35852]_ , \new_[35853]_ ,
    \new_[35857]_ , \new_[35858]_ , \new_[35859]_ , \new_[35863]_ ,
    \new_[35864]_ , \new_[35868]_ , \new_[35869]_ , \new_[35870]_ ,
    \new_[35874]_ , \new_[35875]_ , \new_[35879]_ , \new_[35880]_ ,
    \new_[35881]_ , \new_[35885]_ , \new_[35886]_ , \new_[35890]_ ,
    \new_[35891]_ , \new_[35892]_ , \new_[35896]_ , \new_[35897]_ ,
    \new_[35901]_ , \new_[35902]_ , \new_[35903]_ , \new_[35907]_ ,
    \new_[35908]_ , \new_[35912]_ , \new_[35913]_ , \new_[35914]_ ,
    \new_[35918]_ , \new_[35919]_ , \new_[35923]_ , \new_[35924]_ ,
    \new_[35925]_ , \new_[35929]_ , \new_[35930]_ , \new_[35934]_ ,
    \new_[35935]_ , \new_[35936]_ , \new_[35940]_ , \new_[35941]_ ,
    \new_[35945]_ , \new_[35946]_ , \new_[35947]_ , \new_[35951]_ ,
    \new_[35952]_ , \new_[35956]_ , \new_[35957]_ , \new_[35958]_ ,
    \new_[35962]_ , \new_[35963]_ , \new_[35967]_ , \new_[35968]_ ,
    \new_[35969]_ , \new_[35973]_ , \new_[35974]_ , \new_[35978]_ ,
    \new_[35979]_ , \new_[35980]_ , \new_[35984]_ , \new_[35985]_ ,
    \new_[35989]_ , \new_[35990]_ , \new_[35991]_ , \new_[35995]_ ,
    \new_[35996]_ , \new_[36000]_ , \new_[36001]_ , \new_[36002]_ ,
    \new_[36006]_ , \new_[36007]_ , \new_[36011]_ , \new_[36012]_ ,
    \new_[36013]_ , \new_[36017]_ , \new_[36018]_ , \new_[36022]_ ,
    \new_[36023]_ , \new_[36024]_ , \new_[36028]_ , \new_[36029]_ ,
    \new_[36033]_ , \new_[36034]_ , \new_[36035]_ , \new_[36039]_ ,
    \new_[36040]_ , \new_[36044]_ , \new_[36045]_ , \new_[36046]_ ,
    \new_[36050]_ , \new_[36051]_ , \new_[36055]_ , \new_[36056]_ ,
    \new_[36057]_ , \new_[36061]_ , \new_[36062]_ , \new_[36066]_ ,
    \new_[36067]_ , \new_[36068]_ , \new_[36072]_ , \new_[36073]_ ,
    \new_[36077]_ , \new_[36078]_ , \new_[36079]_ , \new_[36083]_ ,
    \new_[36084]_ , \new_[36088]_ , \new_[36089]_ , \new_[36090]_ ,
    \new_[36094]_ , \new_[36095]_ , \new_[36099]_ , \new_[36100]_ ,
    \new_[36101]_ , \new_[36105]_ , \new_[36106]_ , \new_[36110]_ ,
    \new_[36111]_ , \new_[36112]_ , \new_[36116]_ , \new_[36117]_ ,
    \new_[36121]_ , \new_[36122]_ , \new_[36123]_ , \new_[36127]_ ,
    \new_[36128]_ , \new_[36132]_ , \new_[36133]_ , \new_[36134]_ ,
    \new_[36138]_ , \new_[36139]_ , \new_[36143]_ , \new_[36144]_ ,
    \new_[36145]_ , \new_[36149]_ , \new_[36150]_ , \new_[36154]_ ,
    \new_[36155]_ , \new_[36156]_ , \new_[36160]_ , \new_[36161]_ ,
    \new_[36165]_ , \new_[36166]_ , \new_[36167]_ , \new_[36171]_ ,
    \new_[36172]_ , \new_[36176]_ , \new_[36177]_ , \new_[36178]_ ,
    \new_[36182]_ , \new_[36183]_ , \new_[36187]_ , \new_[36188]_ ,
    \new_[36189]_ , \new_[36193]_ , \new_[36194]_ , \new_[36198]_ ,
    \new_[36199]_ , \new_[36200]_ , \new_[36204]_ , \new_[36205]_ ,
    \new_[36209]_ , \new_[36210]_ , \new_[36211]_ , \new_[36215]_ ,
    \new_[36216]_ , \new_[36220]_ , \new_[36221]_ , \new_[36222]_ ,
    \new_[36226]_ , \new_[36227]_ , \new_[36231]_ , \new_[36232]_ ,
    \new_[36233]_ , \new_[36237]_ , \new_[36238]_ , \new_[36242]_ ,
    \new_[36243]_ , \new_[36244]_ , \new_[36248]_ , \new_[36249]_ ,
    \new_[36253]_ , \new_[36254]_ , \new_[36255]_ , \new_[36259]_ ,
    \new_[36260]_ , \new_[36264]_ , \new_[36265]_ , \new_[36266]_ ,
    \new_[36270]_ , \new_[36271]_ , \new_[36275]_ , \new_[36276]_ ,
    \new_[36277]_ , \new_[36281]_ , \new_[36282]_ , \new_[36286]_ ,
    \new_[36287]_ , \new_[36288]_ , \new_[36292]_ , \new_[36293]_ ,
    \new_[36297]_ , \new_[36298]_ , \new_[36299]_ , \new_[36303]_ ,
    \new_[36304]_ , \new_[36308]_ , \new_[36309]_ , \new_[36310]_ ,
    \new_[36314]_ , \new_[36315]_ , \new_[36319]_ , \new_[36320]_ ,
    \new_[36321]_ , \new_[36325]_ , \new_[36326]_ , \new_[36330]_ ,
    \new_[36331]_ , \new_[36332]_ , \new_[36336]_ , \new_[36337]_ ,
    \new_[36341]_ , \new_[36342]_ , \new_[36343]_ , \new_[36347]_ ,
    \new_[36348]_ , \new_[36352]_ , \new_[36353]_ , \new_[36354]_ ,
    \new_[36358]_ , \new_[36359]_ , \new_[36363]_ , \new_[36364]_ ,
    \new_[36365]_ , \new_[36369]_ , \new_[36370]_ , \new_[36374]_ ,
    \new_[36375]_ , \new_[36376]_ , \new_[36380]_ , \new_[36381]_ ,
    \new_[36385]_ , \new_[36386]_ , \new_[36387]_ , \new_[36391]_ ,
    \new_[36392]_ , \new_[36396]_ , \new_[36397]_ , \new_[36398]_ ,
    \new_[36402]_ , \new_[36403]_ , \new_[36407]_ , \new_[36408]_ ,
    \new_[36409]_ , \new_[36413]_ , \new_[36414]_ , \new_[36418]_ ,
    \new_[36419]_ , \new_[36420]_ , \new_[36424]_ , \new_[36425]_ ,
    \new_[36429]_ , \new_[36430]_ , \new_[36431]_ , \new_[36435]_ ,
    \new_[36436]_ , \new_[36440]_ , \new_[36441]_ , \new_[36442]_ ,
    \new_[36446]_ , \new_[36447]_ , \new_[36451]_ , \new_[36452]_ ,
    \new_[36453]_ , \new_[36457]_ , \new_[36458]_ , \new_[36462]_ ,
    \new_[36463]_ , \new_[36464]_ , \new_[36468]_ , \new_[36469]_ ,
    \new_[36473]_ , \new_[36474]_ , \new_[36475]_ , \new_[36479]_ ,
    \new_[36480]_ , \new_[36484]_ , \new_[36485]_ , \new_[36486]_ ,
    \new_[36490]_ , \new_[36491]_ , \new_[36495]_ , \new_[36496]_ ,
    \new_[36497]_ , \new_[36501]_ , \new_[36502]_ , \new_[36506]_ ,
    \new_[36507]_ , \new_[36508]_ , \new_[36512]_ , \new_[36513]_ ,
    \new_[36517]_ , \new_[36518]_ , \new_[36519]_ , \new_[36523]_ ,
    \new_[36524]_ , \new_[36528]_ , \new_[36529]_ , \new_[36530]_ ,
    \new_[36534]_ , \new_[36535]_ , \new_[36539]_ , \new_[36540]_ ,
    \new_[36541]_ , \new_[36545]_ , \new_[36546]_ , \new_[36550]_ ,
    \new_[36551]_ , \new_[36552]_ , \new_[36556]_ , \new_[36557]_ ,
    \new_[36561]_ , \new_[36562]_ , \new_[36563]_ , \new_[36567]_ ,
    \new_[36568]_ , \new_[36572]_ , \new_[36573]_ , \new_[36574]_ ,
    \new_[36578]_ , \new_[36579]_ , \new_[36583]_ , \new_[36584]_ ,
    \new_[36585]_ , \new_[36589]_ , \new_[36590]_ , \new_[36594]_ ,
    \new_[36595]_ , \new_[36596]_ , \new_[36600]_ , \new_[36601]_ ,
    \new_[36605]_ , \new_[36606]_ , \new_[36607]_ , \new_[36611]_ ,
    \new_[36612]_ , \new_[36616]_ , \new_[36617]_ , \new_[36618]_ ,
    \new_[36622]_ , \new_[36623]_ , \new_[36627]_ , \new_[36628]_ ,
    \new_[36629]_ , \new_[36633]_ , \new_[36634]_ , \new_[36638]_ ,
    \new_[36639]_ , \new_[36640]_ , \new_[36644]_ , \new_[36645]_ ,
    \new_[36649]_ , \new_[36650]_ , \new_[36651]_ , \new_[36655]_ ,
    \new_[36656]_ , \new_[36660]_ , \new_[36661]_ , \new_[36662]_ ,
    \new_[36666]_ , \new_[36667]_ , \new_[36671]_ , \new_[36672]_ ,
    \new_[36673]_ , \new_[36677]_ , \new_[36678]_ , \new_[36682]_ ,
    \new_[36683]_ , \new_[36684]_ , \new_[36688]_ , \new_[36689]_ ,
    \new_[36693]_ , \new_[36694]_ , \new_[36695]_ , \new_[36699]_ ,
    \new_[36700]_ , \new_[36704]_ , \new_[36705]_ , \new_[36706]_ ,
    \new_[36710]_ , \new_[36711]_ , \new_[36715]_ , \new_[36716]_ ,
    \new_[36717]_ , \new_[36721]_ , \new_[36722]_ , \new_[36726]_ ,
    \new_[36727]_ , \new_[36728]_ , \new_[36732]_ , \new_[36733]_ ,
    \new_[36737]_ , \new_[36738]_ , \new_[36739]_ , \new_[36743]_ ,
    \new_[36744]_ , \new_[36748]_ , \new_[36749]_ , \new_[36750]_ ,
    \new_[36754]_ , \new_[36755]_ , \new_[36759]_ , \new_[36760]_ ,
    \new_[36761]_ , \new_[36765]_ , \new_[36766]_ , \new_[36770]_ ,
    \new_[36771]_ , \new_[36772]_ , \new_[36776]_ , \new_[36777]_ ,
    \new_[36781]_ , \new_[36782]_ , \new_[36783]_ , \new_[36787]_ ,
    \new_[36788]_ , \new_[36792]_ , \new_[36793]_ , \new_[36794]_ ,
    \new_[36798]_ , \new_[36799]_ , \new_[36803]_ , \new_[36804]_ ,
    \new_[36805]_ , \new_[36809]_ , \new_[36810]_ , \new_[36814]_ ,
    \new_[36815]_ , \new_[36816]_ , \new_[36820]_ , \new_[36821]_ ,
    \new_[36825]_ , \new_[36826]_ , \new_[36827]_ , \new_[36831]_ ,
    \new_[36832]_ , \new_[36836]_ , \new_[36837]_ , \new_[36838]_ ,
    \new_[36842]_ , \new_[36843]_ , \new_[36847]_ , \new_[36848]_ ,
    \new_[36849]_ , \new_[36853]_ , \new_[36854]_ , \new_[36858]_ ,
    \new_[36859]_ , \new_[36860]_ , \new_[36864]_ , \new_[36865]_ ,
    \new_[36869]_ , \new_[36870]_ , \new_[36871]_ , \new_[36875]_ ,
    \new_[36876]_ , \new_[36880]_ , \new_[36881]_ , \new_[36882]_ ,
    \new_[36886]_ , \new_[36887]_ , \new_[36891]_ , \new_[36892]_ ,
    \new_[36893]_ , \new_[36897]_ , \new_[36898]_ , \new_[36902]_ ,
    \new_[36903]_ , \new_[36904]_ , \new_[36908]_ , \new_[36909]_ ,
    \new_[36913]_ , \new_[36914]_ , \new_[36915]_ , \new_[36919]_ ,
    \new_[36920]_ , \new_[36924]_ , \new_[36925]_ , \new_[36926]_ ,
    \new_[36930]_ , \new_[36931]_ , \new_[36935]_ , \new_[36936]_ ,
    \new_[36937]_ , \new_[36941]_ , \new_[36942]_ , \new_[36946]_ ,
    \new_[36947]_ , \new_[36948]_ , \new_[36952]_ , \new_[36953]_ ,
    \new_[36957]_ , \new_[36958]_ , \new_[36959]_ , \new_[36963]_ ,
    \new_[36964]_ , \new_[36968]_ , \new_[36969]_ , \new_[36970]_ ,
    \new_[36974]_ , \new_[36975]_ , \new_[36979]_ , \new_[36980]_ ,
    \new_[36981]_ , \new_[36985]_ , \new_[36986]_ , \new_[36990]_ ,
    \new_[36991]_ , \new_[36992]_ , \new_[36996]_ , \new_[36997]_ ,
    \new_[37001]_ , \new_[37002]_ , \new_[37003]_ , \new_[37007]_ ,
    \new_[37008]_ , \new_[37012]_ , \new_[37013]_ , \new_[37014]_ ,
    \new_[37018]_ , \new_[37019]_ , \new_[37023]_ , \new_[37024]_ ,
    \new_[37025]_ , \new_[37029]_ , \new_[37030]_ , \new_[37034]_ ,
    \new_[37035]_ , \new_[37036]_ , \new_[37040]_ , \new_[37041]_ ,
    \new_[37045]_ , \new_[37046]_ , \new_[37047]_ , \new_[37051]_ ,
    \new_[37052]_ , \new_[37056]_ , \new_[37057]_ , \new_[37058]_ ,
    \new_[37062]_ , \new_[37063]_ , \new_[37067]_ , \new_[37068]_ ,
    \new_[37069]_ , \new_[37073]_ , \new_[37074]_ , \new_[37078]_ ,
    \new_[37079]_ , \new_[37080]_ , \new_[37084]_ , \new_[37085]_ ,
    \new_[37089]_ , \new_[37090]_ , \new_[37091]_ , \new_[37095]_ ,
    \new_[37096]_ , \new_[37100]_ , \new_[37101]_ , \new_[37102]_ ,
    \new_[37106]_ , \new_[37107]_ , \new_[37111]_ , \new_[37112]_ ,
    \new_[37113]_ , \new_[37117]_ , \new_[37118]_ , \new_[37122]_ ,
    \new_[37123]_ , \new_[37124]_ , \new_[37128]_ , \new_[37129]_ ,
    \new_[37133]_ , \new_[37134]_ , \new_[37135]_ , \new_[37139]_ ,
    \new_[37140]_ , \new_[37144]_ , \new_[37145]_ , \new_[37146]_ ,
    \new_[37150]_ , \new_[37151]_ , \new_[37155]_ , \new_[37156]_ ,
    \new_[37157]_ , \new_[37161]_ , \new_[37162]_ , \new_[37166]_ ,
    \new_[37167]_ , \new_[37168]_ , \new_[37172]_ , \new_[37173]_ ,
    \new_[37177]_ , \new_[37178]_ , \new_[37179]_ , \new_[37183]_ ,
    \new_[37184]_ , \new_[37188]_ , \new_[37189]_ , \new_[37190]_ ,
    \new_[37194]_ , \new_[37195]_ , \new_[37199]_ , \new_[37200]_ ,
    \new_[37201]_ , \new_[37205]_ , \new_[37206]_ , \new_[37210]_ ,
    \new_[37211]_ , \new_[37212]_ , \new_[37216]_ , \new_[37217]_ ,
    \new_[37221]_ , \new_[37222]_ , \new_[37223]_ , \new_[37227]_ ,
    \new_[37228]_ , \new_[37232]_ , \new_[37233]_ , \new_[37234]_ ,
    \new_[37238]_ , \new_[37239]_ , \new_[37243]_ , \new_[37244]_ ,
    \new_[37245]_ , \new_[37249]_ , \new_[37250]_ , \new_[37254]_ ,
    \new_[37255]_ , \new_[37256]_ , \new_[37260]_ , \new_[37261]_ ,
    \new_[37265]_ , \new_[37266]_ , \new_[37267]_ , \new_[37271]_ ,
    \new_[37272]_ , \new_[37276]_ , \new_[37277]_ , \new_[37278]_ ,
    \new_[37282]_ , \new_[37283]_ , \new_[37287]_ , \new_[37288]_ ,
    \new_[37289]_ , \new_[37293]_ , \new_[37294]_ , \new_[37298]_ ,
    \new_[37299]_ , \new_[37300]_ , \new_[37304]_ , \new_[37305]_ ,
    \new_[37309]_ , \new_[37310]_ , \new_[37311]_ , \new_[37315]_ ,
    \new_[37316]_ , \new_[37320]_ , \new_[37321]_ , \new_[37322]_ ,
    \new_[37326]_ , \new_[37327]_ , \new_[37331]_ , \new_[37332]_ ,
    \new_[37333]_ , \new_[37337]_ , \new_[37338]_ , \new_[37342]_ ,
    \new_[37343]_ , \new_[37344]_ , \new_[37348]_ , \new_[37349]_ ,
    \new_[37353]_ , \new_[37354]_ , \new_[37355]_ , \new_[37359]_ ,
    \new_[37360]_ , \new_[37364]_ , \new_[37365]_ , \new_[37366]_ ,
    \new_[37370]_ , \new_[37371]_ , \new_[37375]_ , \new_[37376]_ ,
    \new_[37377]_ , \new_[37381]_ , \new_[37382]_ , \new_[37386]_ ,
    \new_[37387]_ , \new_[37388]_ , \new_[37392]_ , \new_[37393]_ ,
    \new_[37397]_ , \new_[37398]_ , \new_[37399]_ , \new_[37403]_ ,
    \new_[37404]_ , \new_[37408]_ , \new_[37409]_ , \new_[37410]_ ,
    \new_[37414]_ , \new_[37415]_ , \new_[37419]_ , \new_[37420]_ ,
    \new_[37421]_ , \new_[37425]_ , \new_[37426]_ , \new_[37430]_ ,
    \new_[37431]_ , \new_[37432]_ , \new_[37436]_ , \new_[37437]_ ,
    \new_[37441]_ , \new_[37442]_ , \new_[37443]_ , \new_[37447]_ ,
    \new_[37448]_ , \new_[37452]_ , \new_[37453]_ , \new_[37454]_ ,
    \new_[37458]_ , \new_[37459]_ , \new_[37463]_ , \new_[37464]_ ,
    \new_[37465]_ , \new_[37469]_ , \new_[37470]_ , \new_[37474]_ ,
    \new_[37475]_ , \new_[37476]_ , \new_[37480]_ , \new_[37481]_ ,
    \new_[37485]_ , \new_[37486]_ , \new_[37487]_ , \new_[37491]_ ,
    \new_[37492]_ , \new_[37496]_ , \new_[37497]_ , \new_[37498]_ ,
    \new_[37502]_ , \new_[37503]_ , \new_[37507]_ , \new_[37508]_ ,
    \new_[37509]_ , \new_[37513]_ , \new_[37514]_ , \new_[37518]_ ,
    \new_[37519]_ , \new_[37520]_ , \new_[37524]_ , \new_[37525]_ ,
    \new_[37529]_ , \new_[37530]_ , \new_[37531]_ , \new_[37535]_ ,
    \new_[37536]_ , \new_[37540]_ , \new_[37541]_ , \new_[37542]_ ,
    \new_[37546]_ , \new_[37547]_ , \new_[37551]_ , \new_[37552]_ ,
    \new_[37553]_ , \new_[37557]_ , \new_[37558]_ , \new_[37562]_ ,
    \new_[37563]_ , \new_[37564]_ , \new_[37568]_ , \new_[37569]_ ,
    \new_[37573]_ , \new_[37574]_ , \new_[37575]_ , \new_[37579]_ ,
    \new_[37580]_ , \new_[37584]_ , \new_[37585]_ , \new_[37586]_ ,
    \new_[37590]_ , \new_[37591]_ , \new_[37595]_ , \new_[37596]_ ,
    \new_[37597]_ , \new_[37601]_ , \new_[37602]_ , \new_[37606]_ ,
    \new_[37607]_ , \new_[37608]_ , \new_[37612]_ , \new_[37613]_ ,
    \new_[37617]_ , \new_[37618]_ , \new_[37619]_ , \new_[37623]_ ,
    \new_[37624]_ , \new_[37628]_ , \new_[37629]_ , \new_[37630]_ ,
    \new_[37634]_ , \new_[37635]_ , \new_[37639]_ , \new_[37640]_ ,
    \new_[37641]_ , \new_[37645]_ , \new_[37646]_ , \new_[37650]_ ,
    \new_[37651]_ , \new_[37652]_ , \new_[37656]_ , \new_[37657]_ ,
    \new_[37661]_ , \new_[37662]_ , \new_[37663]_ , \new_[37667]_ ,
    \new_[37668]_ , \new_[37672]_ , \new_[37673]_ , \new_[37674]_ ,
    \new_[37678]_ , \new_[37679]_ , \new_[37683]_ , \new_[37684]_ ,
    \new_[37685]_ , \new_[37689]_ , \new_[37690]_ , \new_[37694]_ ,
    \new_[37695]_ , \new_[37696]_ , \new_[37700]_ , \new_[37701]_ ,
    \new_[37705]_ , \new_[37706]_ , \new_[37707]_ , \new_[37711]_ ,
    \new_[37712]_ , \new_[37716]_ , \new_[37717]_ , \new_[37718]_ ,
    \new_[37722]_ , \new_[37723]_ , \new_[37727]_ , \new_[37728]_ ,
    \new_[37729]_ , \new_[37733]_ , \new_[37734]_ , \new_[37738]_ ,
    \new_[37739]_ , \new_[37740]_ , \new_[37744]_ , \new_[37745]_ ,
    \new_[37749]_ , \new_[37750]_ , \new_[37751]_ , \new_[37755]_ ,
    \new_[37756]_ , \new_[37760]_ , \new_[37761]_ , \new_[37762]_ ,
    \new_[37766]_ , \new_[37767]_ , \new_[37771]_ , \new_[37772]_ ,
    \new_[37773]_ , \new_[37777]_ , \new_[37778]_ , \new_[37782]_ ,
    \new_[37783]_ , \new_[37784]_ , \new_[37788]_ , \new_[37789]_ ,
    \new_[37793]_ , \new_[37794]_ , \new_[37795]_ , \new_[37799]_ ,
    \new_[37800]_ , \new_[37804]_ , \new_[37805]_ , \new_[37806]_ ,
    \new_[37810]_ , \new_[37811]_ , \new_[37815]_ , \new_[37816]_ ,
    \new_[37817]_ , \new_[37821]_ , \new_[37822]_ , \new_[37826]_ ,
    \new_[37827]_ , \new_[37828]_ , \new_[37832]_ , \new_[37833]_ ,
    \new_[37837]_ , \new_[37838]_ , \new_[37839]_ , \new_[37843]_ ,
    \new_[37844]_ , \new_[37848]_ , \new_[37849]_ , \new_[37850]_ ,
    \new_[37854]_ , \new_[37855]_ , \new_[37859]_ , \new_[37860]_ ,
    \new_[37861]_ , \new_[37865]_ , \new_[37866]_ , \new_[37870]_ ,
    \new_[37871]_ , \new_[37872]_ , \new_[37876]_ , \new_[37877]_ ,
    \new_[37881]_ , \new_[37882]_ , \new_[37883]_ , \new_[37887]_ ,
    \new_[37888]_ , \new_[37892]_ , \new_[37893]_ , \new_[37894]_ ,
    \new_[37898]_ , \new_[37899]_ , \new_[37903]_ , \new_[37904]_ ,
    \new_[37905]_ , \new_[37909]_ , \new_[37910]_ , \new_[37914]_ ,
    \new_[37915]_ , \new_[37916]_ , \new_[37920]_ , \new_[37921]_ ,
    \new_[37925]_ , \new_[37926]_ , \new_[37927]_ , \new_[37931]_ ,
    \new_[37932]_ , \new_[37936]_ , \new_[37937]_ , \new_[37938]_ ,
    \new_[37942]_ , \new_[37943]_ , \new_[37947]_ , \new_[37948]_ ,
    \new_[37949]_ , \new_[37953]_ , \new_[37954]_ , \new_[37958]_ ,
    \new_[37959]_ , \new_[37960]_ , \new_[37964]_ , \new_[37965]_ ,
    \new_[37969]_ , \new_[37970]_ , \new_[37971]_ , \new_[37975]_ ,
    \new_[37976]_ , \new_[37980]_ , \new_[37981]_ , \new_[37982]_ ,
    \new_[37986]_ , \new_[37987]_ , \new_[37991]_ , \new_[37992]_ ,
    \new_[37993]_ , \new_[37997]_ , \new_[37998]_ , \new_[38002]_ ,
    \new_[38003]_ , \new_[38004]_ , \new_[38008]_ , \new_[38009]_ ,
    \new_[38013]_ , \new_[38014]_ , \new_[38015]_ , \new_[38019]_ ,
    \new_[38020]_ , \new_[38024]_ , \new_[38025]_ , \new_[38026]_ ,
    \new_[38030]_ , \new_[38031]_ , \new_[38035]_ , \new_[38036]_ ,
    \new_[38037]_ , \new_[38041]_ , \new_[38042]_ , \new_[38046]_ ,
    \new_[38047]_ , \new_[38048]_ , \new_[38052]_ , \new_[38053]_ ,
    \new_[38057]_ , \new_[38058]_ , \new_[38059]_ , \new_[38063]_ ,
    \new_[38064]_ , \new_[38068]_ , \new_[38069]_ , \new_[38070]_ ,
    \new_[38074]_ , \new_[38075]_ , \new_[38079]_ , \new_[38080]_ ,
    \new_[38081]_ , \new_[38085]_ , \new_[38086]_ , \new_[38090]_ ,
    \new_[38091]_ , \new_[38092]_ , \new_[38096]_ , \new_[38097]_ ,
    \new_[38101]_ , \new_[38102]_ , \new_[38103]_ , \new_[38107]_ ,
    \new_[38108]_ , \new_[38112]_ , \new_[38113]_ , \new_[38114]_ ,
    \new_[38118]_ , \new_[38119]_ , \new_[38123]_ , \new_[38124]_ ,
    \new_[38125]_ , \new_[38129]_ , \new_[38130]_ , \new_[38134]_ ,
    \new_[38135]_ , \new_[38136]_ , \new_[38140]_ , \new_[38141]_ ,
    \new_[38145]_ , \new_[38146]_ , \new_[38147]_ , \new_[38151]_ ,
    \new_[38152]_ , \new_[38156]_ , \new_[38157]_ , \new_[38158]_ ,
    \new_[38162]_ , \new_[38163]_ , \new_[38167]_ , \new_[38168]_ ,
    \new_[38169]_ , \new_[38173]_ , \new_[38174]_ , \new_[38178]_ ,
    \new_[38179]_ , \new_[38180]_ , \new_[38184]_ , \new_[38185]_ ,
    \new_[38189]_ , \new_[38190]_ , \new_[38191]_ , \new_[38195]_ ,
    \new_[38196]_ , \new_[38200]_ , \new_[38201]_ , \new_[38202]_ ,
    \new_[38206]_ , \new_[38207]_ , \new_[38211]_ , \new_[38212]_ ,
    \new_[38213]_ , \new_[38217]_ , \new_[38218]_ , \new_[38222]_ ,
    \new_[38223]_ , \new_[38224]_ , \new_[38228]_ , \new_[38229]_ ,
    \new_[38233]_ , \new_[38234]_ , \new_[38235]_ , \new_[38239]_ ,
    \new_[38240]_ , \new_[38244]_ , \new_[38245]_ , \new_[38246]_ ,
    \new_[38250]_ , \new_[38251]_ , \new_[38255]_ , \new_[38256]_ ,
    \new_[38257]_ , \new_[38261]_ , \new_[38262]_ , \new_[38266]_ ,
    \new_[38267]_ , \new_[38268]_ , \new_[38272]_ , \new_[38273]_ ,
    \new_[38277]_ , \new_[38278]_ , \new_[38279]_ , \new_[38283]_ ,
    \new_[38284]_ , \new_[38288]_ , \new_[38289]_ , \new_[38290]_ ,
    \new_[38294]_ , \new_[38295]_ , \new_[38299]_ , \new_[38300]_ ,
    \new_[38301]_ , \new_[38305]_ , \new_[38306]_ , \new_[38310]_ ,
    \new_[38311]_ , \new_[38312]_ , \new_[38316]_ , \new_[38317]_ ,
    \new_[38321]_ , \new_[38322]_ , \new_[38323]_ , \new_[38327]_ ,
    \new_[38328]_ , \new_[38332]_ , \new_[38333]_ , \new_[38334]_ ,
    \new_[38338]_ , \new_[38339]_ , \new_[38343]_ , \new_[38344]_ ,
    \new_[38345]_ , \new_[38349]_ , \new_[38350]_ , \new_[38354]_ ,
    \new_[38355]_ , \new_[38356]_ , \new_[38360]_ , \new_[38361]_ ,
    \new_[38365]_ , \new_[38366]_ , \new_[38367]_ , \new_[38371]_ ,
    \new_[38372]_ , \new_[38376]_ , \new_[38377]_ , \new_[38378]_ ,
    \new_[38382]_ , \new_[38383]_ , \new_[38387]_ , \new_[38388]_ ,
    \new_[38389]_ , \new_[38393]_ , \new_[38394]_ , \new_[38398]_ ,
    \new_[38399]_ , \new_[38400]_ , \new_[38404]_ , \new_[38405]_ ,
    \new_[38409]_ , \new_[38410]_ , \new_[38411]_ , \new_[38415]_ ,
    \new_[38416]_ , \new_[38420]_ , \new_[38421]_ , \new_[38422]_ ,
    \new_[38426]_ , \new_[38427]_ , \new_[38431]_ , \new_[38432]_ ,
    \new_[38433]_ , \new_[38437]_ , \new_[38438]_ , \new_[38442]_ ,
    \new_[38443]_ , \new_[38444]_ , \new_[38448]_ , \new_[38449]_ ,
    \new_[38453]_ , \new_[38454]_ , \new_[38455]_ , \new_[38459]_ ,
    \new_[38460]_ , \new_[38464]_ , \new_[38465]_ , \new_[38466]_ ,
    \new_[38470]_ , \new_[38471]_ , \new_[38475]_ , \new_[38476]_ ,
    \new_[38477]_ , \new_[38481]_ , \new_[38482]_ , \new_[38486]_ ,
    \new_[38487]_ , \new_[38488]_ , \new_[38492]_ , \new_[38493]_ ,
    \new_[38497]_ , \new_[38498]_ , \new_[38499]_ , \new_[38503]_ ,
    \new_[38504]_ , \new_[38508]_ , \new_[38509]_ , \new_[38510]_ ,
    \new_[38514]_ , \new_[38515]_ , \new_[38519]_ , \new_[38520]_ ,
    \new_[38521]_ , \new_[38525]_ , \new_[38526]_ , \new_[38530]_ ,
    \new_[38531]_ , \new_[38532]_ , \new_[38536]_ , \new_[38537]_ ,
    \new_[38541]_ , \new_[38542]_ , \new_[38543]_ , \new_[38547]_ ,
    \new_[38548]_ , \new_[38552]_ , \new_[38553]_ , \new_[38554]_ ,
    \new_[38558]_ , \new_[38559]_ , \new_[38563]_ , \new_[38564]_ ,
    \new_[38565]_ , \new_[38569]_ , \new_[38570]_ , \new_[38574]_ ,
    \new_[38575]_ , \new_[38576]_ , \new_[38580]_ , \new_[38581]_ ,
    \new_[38585]_ , \new_[38586]_ , \new_[38587]_ , \new_[38591]_ ,
    \new_[38592]_ , \new_[38596]_ , \new_[38597]_ , \new_[38598]_ ,
    \new_[38602]_ , \new_[38603]_ , \new_[38607]_ , \new_[38608]_ ,
    \new_[38609]_ , \new_[38613]_ , \new_[38614]_ , \new_[38618]_ ,
    \new_[38619]_ , \new_[38620]_ , \new_[38624]_ , \new_[38625]_ ,
    \new_[38629]_ , \new_[38630]_ , \new_[38631]_ , \new_[38635]_ ,
    \new_[38636]_ , \new_[38640]_ , \new_[38641]_ , \new_[38642]_ ,
    \new_[38646]_ , \new_[38647]_ , \new_[38651]_ , \new_[38652]_ ,
    \new_[38653]_ , \new_[38657]_ , \new_[38658]_ , \new_[38662]_ ,
    \new_[38663]_ , \new_[38664]_ , \new_[38668]_ , \new_[38669]_ ,
    \new_[38673]_ , \new_[38674]_ , \new_[38675]_ , \new_[38679]_ ,
    \new_[38680]_ , \new_[38684]_ , \new_[38685]_ , \new_[38686]_ ,
    \new_[38690]_ , \new_[38691]_ , \new_[38695]_ , \new_[38696]_ ,
    \new_[38697]_ , \new_[38701]_ , \new_[38702]_ , \new_[38706]_ ,
    \new_[38707]_ , \new_[38708]_ , \new_[38712]_ , \new_[38713]_ ,
    \new_[38717]_ , \new_[38718]_ , \new_[38719]_ , \new_[38723]_ ,
    \new_[38724]_ , \new_[38728]_ , \new_[38729]_ , \new_[38730]_ ,
    \new_[38734]_ , \new_[38735]_ , \new_[38739]_ , \new_[38740]_ ,
    \new_[38741]_ , \new_[38745]_ , \new_[38746]_ , \new_[38750]_ ,
    \new_[38751]_ , \new_[38752]_ , \new_[38756]_ , \new_[38757]_ ,
    \new_[38761]_ , \new_[38762]_ , \new_[38763]_ , \new_[38767]_ ,
    \new_[38768]_ , \new_[38772]_ , \new_[38773]_ , \new_[38774]_ ,
    \new_[38778]_ , \new_[38779]_ , \new_[38783]_ , \new_[38784]_ ,
    \new_[38785]_ , \new_[38789]_ , \new_[38790]_ , \new_[38794]_ ,
    \new_[38795]_ , \new_[38796]_ , \new_[38800]_ , \new_[38801]_ ,
    \new_[38805]_ , \new_[38806]_ , \new_[38807]_ , \new_[38811]_ ,
    \new_[38812]_ , \new_[38816]_ , \new_[38817]_ , \new_[38818]_ ,
    \new_[38822]_ , \new_[38823]_ , \new_[38827]_ , \new_[38828]_ ,
    \new_[38829]_ , \new_[38833]_ , \new_[38834]_ , \new_[38838]_ ,
    \new_[38839]_ , \new_[38840]_ , \new_[38844]_ , \new_[38845]_ ,
    \new_[38849]_ , \new_[38850]_ , \new_[38851]_ , \new_[38855]_ ,
    \new_[38856]_ , \new_[38860]_ , \new_[38861]_ , \new_[38862]_ ,
    \new_[38866]_ , \new_[38867]_ , \new_[38871]_ , \new_[38872]_ ,
    \new_[38873]_ , \new_[38877]_ , \new_[38878]_ , \new_[38882]_ ,
    \new_[38883]_ , \new_[38884]_ , \new_[38888]_ , \new_[38889]_ ,
    \new_[38893]_ , \new_[38894]_ , \new_[38895]_ , \new_[38899]_ ,
    \new_[38900]_ , \new_[38904]_ , \new_[38905]_ , \new_[38906]_ ,
    \new_[38910]_ , \new_[38911]_ , \new_[38915]_ , \new_[38916]_ ,
    \new_[38917]_ , \new_[38921]_ , \new_[38922]_ , \new_[38926]_ ,
    \new_[38927]_ , \new_[38928]_ , \new_[38932]_ , \new_[38933]_ ,
    \new_[38937]_ , \new_[38938]_ , \new_[38939]_ , \new_[38943]_ ,
    \new_[38944]_ , \new_[38948]_ , \new_[38949]_ , \new_[38950]_ ,
    \new_[38954]_ , \new_[38955]_ , \new_[38959]_ , \new_[38960]_ ,
    \new_[38961]_ , \new_[38965]_ , \new_[38966]_ , \new_[38970]_ ,
    \new_[38971]_ , \new_[38972]_ , \new_[38976]_ , \new_[38977]_ ,
    \new_[38981]_ , \new_[38982]_ , \new_[38983]_ , \new_[38987]_ ,
    \new_[38988]_ , \new_[38992]_ , \new_[38993]_ , \new_[38994]_ ,
    \new_[38998]_ , \new_[38999]_ , \new_[39003]_ , \new_[39004]_ ,
    \new_[39005]_ , \new_[39009]_ , \new_[39010]_ , \new_[39014]_ ,
    \new_[39015]_ , \new_[39016]_ , \new_[39020]_ , \new_[39021]_ ,
    \new_[39025]_ , \new_[39026]_ , \new_[39027]_ , \new_[39031]_ ,
    \new_[39032]_ , \new_[39036]_ , \new_[39037]_ , \new_[39038]_ ,
    \new_[39042]_ , \new_[39043]_ , \new_[39047]_ , \new_[39048]_ ,
    \new_[39049]_ , \new_[39053]_ , \new_[39054]_ , \new_[39058]_ ,
    \new_[39059]_ , \new_[39060]_ , \new_[39064]_ , \new_[39065]_ ,
    \new_[39069]_ , \new_[39070]_ , \new_[39071]_ , \new_[39075]_ ,
    \new_[39076]_ , \new_[39080]_ , \new_[39081]_ , \new_[39082]_ ,
    \new_[39086]_ , \new_[39087]_ , \new_[39091]_ , \new_[39092]_ ,
    \new_[39093]_ , \new_[39097]_ , \new_[39098]_ , \new_[39102]_ ,
    \new_[39103]_ , \new_[39104]_ , \new_[39108]_ , \new_[39109]_ ,
    \new_[39113]_ , \new_[39114]_ , \new_[39115]_ , \new_[39119]_ ,
    \new_[39120]_ , \new_[39124]_ , \new_[39125]_ , \new_[39126]_ ,
    \new_[39130]_ , \new_[39131]_ , \new_[39135]_ , \new_[39136]_ ,
    \new_[39137]_ , \new_[39141]_ , \new_[39142]_ , \new_[39146]_ ,
    \new_[39147]_ , \new_[39148]_ , \new_[39152]_ , \new_[39153]_ ,
    \new_[39157]_ , \new_[39158]_ , \new_[39159]_ , \new_[39163]_ ,
    \new_[39164]_ , \new_[39168]_ , \new_[39169]_ , \new_[39170]_ ,
    \new_[39174]_ , \new_[39175]_ , \new_[39179]_ , \new_[39180]_ ,
    \new_[39181]_ , \new_[39185]_ , \new_[39186]_ , \new_[39190]_ ,
    \new_[39191]_ , \new_[39192]_ , \new_[39196]_ , \new_[39197]_ ,
    \new_[39201]_ , \new_[39202]_ , \new_[39203]_ , \new_[39207]_ ,
    \new_[39208]_ , \new_[39212]_ , \new_[39213]_ , \new_[39214]_ ,
    \new_[39218]_ , \new_[39219]_ , \new_[39223]_ , \new_[39224]_ ,
    \new_[39225]_ , \new_[39229]_ , \new_[39230]_ , \new_[39234]_ ,
    \new_[39235]_ , \new_[39236]_ , \new_[39240]_ , \new_[39241]_ ,
    \new_[39245]_ , \new_[39246]_ , \new_[39247]_ , \new_[39251]_ ,
    \new_[39252]_ , \new_[39256]_ , \new_[39257]_ , \new_[39258]_ ,
    \new_[39262]_ , \new_[39263]_ , \new_[39267]_ , \new_[39268]_ ,
    \new_[39269]_ , \new_[39273]_ , \new_[39274]_ , \new_[39278]_ ,
    \new_[39279]_ , \new_[39280]_ , \new_[39284]_ , \new_[39285]_ ,
    \new_[39289]_ , \new_[39290]_ , \new_[39291]_ , \new_[39295]_ ,
    \new_[39296]_ , \new_[39300]_ , \new_[39301]_ , \new_[39302]_ ,
    \new_[39306]_ , \new_[39307]_ , \new_[39311]_ , \new_[39312]_ ,
    \new_[39313]_ , \new_[39317]_ , \new_[39318]_ , \new_[39322]_ ,
    \new_[39323]_ , \new_[39324]_ , \new_[39328]_ , \new_[39329]_ ,
    \new_[39333]_ , \new_[39334]_ , \new_[39335]_ , \new_[39339]_ ,
    \new_[39340]_ , \new_[39344]_ , \new_[39345]_ , \new_[39346]_ ,
    \new_[39350]_ , \new_[39351]_ , \new_[39355]_ , \new_[39356]_ ,
    \new_[39357]_ , \new_[39361]_ , \new_[39362]_ , \new_[39366]_ ,
    \new_[39367]_ , \new_[39368]_ , \new_[39372]_ , \new_[39373]_ ,
    \new_[39377]_ , \new_[39378]_ , \new_[39379]_ , \new_[39383]_ ,
    \new_[39384]_ , \new_[39388]_ , \new_[39389]_ , \new_[39390]_ ,
    \new_[39394]_ , \new_[39395]_ , \new_[39399]_ , \new_[39400]_ ,
    \new_[39401]_ , \new_[39405]_ , \new_[39406]_ , \new_[39410]_ ,
    \new_[39411]_ , \new_[39412]_ , \new_[39416]_ , \new_[39417]_ ,
    \new_[39421]_ , \new_[39422]_ , \new_[39423]_ , \new_[39427]_ ,
    \new_[39428]_ , \new_[39432]_ , \new_[39433]_ , \new_[39434]_ ,
    \new_[39438]_ , \new_[39439]_ , \new_[39443]_ , \new_[39444]_ ,
    \new_[39445]_ , \new_[39449]_ , \new_[39450]_ , \new_[39454]_ ,
    \new_[39455]_ , \new_[39456]_ , \new_[39460]_ , \new_[39461]_ ,
    \new_[39465]_ , \new_[39466]_ , \new_[39467]_ , \new_[39471]_ ,
    \new_[39472]_ , \new_[39476]_ , \new_[39477]_ , \new_[39478]_ ,
    \new_[39482]_ , \new_[39483]_ , \new_[39487]_ , \new_[39488]_ ,
    \new_[39489]_ , \new_[39493]_ , \new_[39494]_ , \new_[39498]_ ,
    \new_[39499]_ , \new_[39500]_ , \new_[39504]_ , \new_[39505]_ ,
    \new_[39509]_ , \new_[39510]_ , \new_[39511]_ , \new_[39515]_ ,
    \new_[39516]_ , \new_[39520]_ , \new_[39521]_ , \new_[39522]_ ,
    \new_[39526]_ , \new_[39527]_ , \new_[39531]_ , \new_[39532]_ ,
    \new_[39533]_ , \new_[39537]_ , \new_[39538]_ , \new_[39542]_ ,
    \new_[39543]_ , \new_[39544]_ , \new_[39548]_ , \new_[39549]_ ,
    \new_[39553]_ , \new_[39554]_ , \new_[39555]_ , \new_[39559]_ ,
    \new_[39560]_ , \new_[39564]_ , \new_[39565]_ , \new_[39566]_ ,
    \new_[39570]_ , \new_[39571]_ , \new_[39575]_ , \new_[39576]_ ,
    \new_[39577]_ , \new_[39581]_ , \new_[39582]_ , \new_[39586]_ ,
    \new_[39587]_ , \new_[39588]_ , \new_[39592]_ , \new_[39593]_ ,
    \new_[39597]_ , \new_[39598]_ , \new_[39599]_ , \new_[39603]_ ,
    \new_[39604]_ , \new_[39608]_ , \new_[39609]_ , \new_[39610]_ ,
    \new_[39614]_ , \new_[39615]_ , \new_[39619]_ , \new_[39620]_ ,
    \new_[39621]_ , \new_[39625]_ , \new_[39626]_ , \new_[39630]_ ,
    \new_[39631]_ , \new_[39632]_ , \new_[39636]_ , \new_[39637]_ ,
    \new_[39641]_ , \new_[39642]_ , \new_[39643]_ , \new_[39647]_ ,
    \new_[39648]_ , \new_[39652]_ , \new_[39653]_ , \new_[39654]_ ,
    \new_[39658]_ , \new_[39659]_ , \new_[39663]_ , \new_[39664]_ ,
    \new_[39665]_ , \new_[39669]_ , \new_[39670]_ , \new_[39674]_ ,
    \new_[39675]_ , \new_[39676]_ , \new_[39680]_ , \new_[39681]_ ,
    \new_[39685]_ , \new_[39686]_ , \new_[39687]_ , \new_[39691]_ ,
    \new_[39692]_ , \new_[39696]_ , \new_[39697]_ , \new_[39698]_ ,
    \new_[39702]_ , \new_[39703]_ , \new_[39707]_ , \new_[39708]_ ,
    \new_[39709]_ , \new_[39713]_ , \new_[39714]_ , \new_[39718]_ ,
    \new_[39719]_ , \new_[39720]_ , \new_[39724]_ , \new_[39725]_ ,
    \new_[39729]_ , \new_[39730]_ , \new_[39731]_ , \new_[39735]_ ,
    \new_[39736]_ , \new_[39740]_ , \new_[39741]_ , \new_[39742]_ ,
    \new_[39746]_ , \new_[39747]_ , \new_[39751]_ , \new_[39752]_ ,
    \new_[39753]_ , \new_[39757]_ , \new_[39758]_ , \new_[39762]_ ,
    \new_[39763]_ , \new_[39764]_ , \new_[39768]_ , \new_[39769]_ ,
    \new_[39773]_ , \new_[39774]_ , \new_[39775]_ , \new_[39779]_ ,
    \new_[39780]_ , \new_[39784]_ , \new_[39785]_ , \new_[39786]_ ,
    \new_[39790]_ , \new_[39791]_ , \new_[39795]_ , \new_[39796]_ ,
    \new_[39797]_ , \new_[39801]_ , \new_[39802]_ , \new_[39806]_ ,
    \new_[39807]_ , \new_[39808]_ , \new_[39812]_ , \new_[39813]_ ,
    \new_[39817]_ , \new_[39818]_ , \new_[39819]_ , \new_[39823]_ ,
    \new_[39824]_ , \new_[39828]_ , \new_[39829]_ , \new_[39830]_ ,
    \new_[39834]_ , \new_[39835]_ , \new_[39839]_ , \new_[39840]_ ,
    \new_[39841]_ , \new_[39845]_ , \new_[39846]_ , \new_[39850]_ ,
    \new_[39851]_ , \new_[39852]_ , \new_[39856]_ , \new_[39857]_ ,
    \new_[39861]_ , \new_[39862]_ , \new_[39863]_ , \new_[39867]_ ,
    \new_[39868]_ , \new_[39872]_ , \new_[39873]_ , \new_[39874]_ ,
    \new_[39878]_ , \new_[39879]_ , \new_[39883]_ , \new_[39884]_ ,
    \new_[39885]_ , \new_[39889]_ , \new_[39890]_ , \new_[39894]_ ,
    \new_[39895]_ , \new_[39896]_ , \new_[39900]_ , \new_[39901]_ ,
    \new_[39905]_ , \new_[39906]_ , \new_[39907]_ , \new_[39911]_ ,
    \new_[39912]_ , \new_[39916]_ , \new_[39917]_ , \new_[39918]_ ,
    \new_[39922]_ , \new_[39923]_ , \new_[39927]_ , \new_[39928]_ ,
    \new_[39929]_ , \new_[39933]_ , \new_[39934]_ , \new_[39938]_ ,
    \new_[39939]_ , \new_[39940]_ , \new_[39944]_ , \new_[39945]_ ,
    \new_[39949]_ , \new_[39950]_ , \new_[39951]_ , \new_[39955]_ ,
    \new_[39956]_ , \new_[39960]_ , \new_[39961]_ , \new_[39962]_ ,
    \new_[39966]_ , \new_[39967]_ , \new_[39971]_ , \new_[39972]_ ,
    \new_[39973]_ , \new_[39977]_ , \new_[39978]_ , \new_[39982]_ ,
    \new_[39983]_ , \new_[39984]_ , \new_[39988]_ , \new_[39989]_ ,
    \new_[39993]_ , \new_[39994]_ , \new_[39995]_ , \new_[39999]_ ,
    \new_[40000]_ , \new_[40004]_ , \new_[40005]_ , \new_[40006]_ ,
    \new_[40010]_ , \new_[40011]_ , \new_[40015]_ , \new_[40016]_ ,
    \new_[40017]_ , \new_[40021]_ , \new_[40022]_ , \new_[40026]_ ,
    \new_[40027]_ , \new_[40028]_ , \new_[40032]_ , \new_[40033]_ ,
    \new_[40037]_ , \new_[40038]_ , \new_[40039]_ , \new_[40043]_ ,
    \new_[40044]_ , \new_[40048]_ , \new_[40049]_ , \new_[40050]_ ,
    \new_[40054]_ , \new_[40055]_ , \new_[40059]_ , \new_[40060]_ ,
    \new_[40061]_ , \new_[40065]_ , \new_[40066]_ , \new_[40070]_ ,
    \new_[40071]_ , \new_[40072]_ , \new_[40076]_ , \new_[40077]_ ,
    \new_[40081]_ , \new_[40082]_ , \new_[40083]_ , \new_[40087]_ ,
    \new_[40088]_ , \new_[40092]_ , \new_[40093]_ , \new_[40094]_ ,
    \new_[40098]_ , \new_[40099]_ , \new_[40103]_ , \new_[40104]_ ,
    \new_[40105]_ , \new_[40109]_ , \new_[40110]_ , \new_[40114]_ ,
    \new_[40115]_ , \new_[40116]_ , \new_[40120]_ , \new_[40121]_ ,
    \new_[40125]_ , \new_[40126]_ , \new_[40127]_ , \new_[40131]_ ,
    \new_[40132]_ , \new_[40136]_ , \new_[40137]_ , \new_[40138]_ ,
    \new_[40142]_ , \new_[40143]_ , \new_[40147]_ , \new_[40148]_ ,
    \new_[40149]_ , \new_[40153]_ , \new_[40154]_ , \new_[40158]_ ,
    \new_[40159]_ , \new_[40160]_ , \new_[40164]_ , \new_[40165]_ ,
    \new_[40169]_ , \new_[40170]_ , \new_[40171]_ , \new_[40175]_ ,
    \new_[40176]_ , \new_[40180]_ , \new_[40181]_ , \new_[40182]_ ,
    \new_[40186]_ , \new_[40187]_ , \new_[40191]_ , \new_[40192]_ ,
    \new_[40193]_ , \new_[40197]_ , \new_[40198]_ , \new_[40202]_ ,
    \new_[40203]_ , \new_[40204]_ , \new_[40208]_ , \new_[40209]_ ,
    \new_[40213]_ , \new_[40214]_ , \new_[40215]_ , \new_[40219]_ ,
    \new_[40220]_ , \new_[40224]_ , \new_[40225]_ , \new_[40226]_ ,
    \new_[40230]_ , \new_[40231]_ , \new_[40235]_ , \new_[40236]_ ,
    \new_[40237]_ , \new_[40241]_ , \new_[40242]_ , \new_[40246]_ ,
    \new_[40247]_ , \new_[40248]_ , \new_[40252]_ , \new_[40253]_ ,
    \new_[40257]_ , \new_[40258]_ , \new_[40259]_ , \new_[40263]_ ,
    \new_[40264]_ , \new_[40268]_ , \new_[40269]_ , \new_[40270]_ ,
    \new_[40274]_ , \new_[40275]_ , \new_[40279]_ , \new_[40280]_ ,
    \new_[40281]_ , \new_[40285]_ , \new_[40286]_ , \new_[40290]_ ,
    \new_[40291]_ , \new_[40292]_ , \new_[40296]_ , \new_[40297]_ ,
    \new_[40301]_ , \new_[40302]_ , \new_[40303]_ , \new_[40307]_ ,
    \new_[40308]_ , \new_[40312]_ , \new_[40313]_ , \new_[40314]_ ,
    \new_[40318]_ , \new_[40319]_ , \new_[40323]_ , \new_[40324]_ ,
    \new_[40325]_ , \new_[40329]_ , \new_[40330]_ , \new_[40334]_ ,
    \new_[40335]_ , \new_[40336]_ , \new_[40340]_ , \new_[40341]_ ,
    \new_[40345]_ , \new_[40346]_ , \new_[40347]_ , \new_[40351]_ ,
    \new_[40352]_ , \new_[40355]_ , \new_[40358]_ , \new_[40359]_ ,
    \new_[40360]_ , \new_[40364]_ , \new_[40365]_ , \new_[40369]_ ,
    \new_[40370]_ , \new_[40371]_ , \new_[40375]_ , \new_[40376]_ ,
    \new_[40379]_ , \new_[40382]_ , \new_[40383]_ , \new_[40384]_ ,
    \new_[40388]_ , \new_[40389]_ , \new_[40393]_ , \new_[40394]_ ,
    \new_[40395]_ , \new_[40399]_ , \new_[40400]_ , \new_[40403]_ ,
    \new_[40406]_ , \new_[40407]_ , \new_[40408]_ , \new_[40412]_ ,
    \new_[40413]_ , \new_[40417]_ , \new_[40418]_ , \new_[40419]_ ,
    \new_[40423]_ , \new_[40424]_ , \new_[40427]_ , \new_[40430]_ ,
    \new_[40431]_ , \new_[40432]_ , \new_[40436]_ , \new_[40437]_ ,
    \new_[40441]_ , \new_[40442]_ , \new_[40443]_ , \new_[40447]_ ,
    \new_[40448]_ , \new_[40451]_ , \new_[40454]_ , \new_[40455]_ ,
    \new_[40456]_ , \new_[40460]_ , \new_[40461]_ , \new_[40465]_ ,
    \new_[40466]_ , \new_[40467]_ , \new_[40471]_ , \new_[40472]_ ,
    \new_[40475]_ , \new_[40478]_ , \new_[40479]_ , \new_[40480]_ ,
    \new_[40484]_ , \new_[40485]_ , \new_[40489]_ , \new_[40490]_ ,
    \new_[40491]_ , \new_[40495]_ , \new_[40496]_ , \new_[40499]_ ,
    \new_[40502]_ , \new_[40503]_ , \new_[40504]_ , \new_[40508]_ ,
    \new_[40509]_ , \new_[40513]_ , \new_[40514]_ , \new_[40515]_ ,
    \new_[40519]_ , \new_[40520]_ , \new_[40523]_ , \new_[40526]_ ,
    \new_[40527]_ , \new_[40528]_ , \new_[40532]_ , \new_[40533]_ ,
    \new_[40537]_ , \new_[40538]_ , \new_[40539]_ , \new_[40543]_ ,
    \new_[40544]_ , \new_[40547]_ , \new_[40550]_ , \new_[40551]_ ,
    \new_[40552]_ , \new_[40556]_ , \new_[40557]_ , \new_[40561]_ ,
    \new_[40562]_ , \new_[40563]_ , \new_[40567]_ , \new_[40568]_ ,
    \new_[40571]_ , \new_[40574]_ , \new_[40575]_ , \new_[40576]_ ,
    \new_[40580]_ , \new_[40581]_ , \new_[40585]_ , \new_[40586]_ ,
    \new_[40587]_ , \new_[40591]_ , \new_[40592]_ , \new_[40595]_ ,
    \new_[40598]_ , \new_[40599]_ , \new_[40600]_ , \new_[40604]_ ,
    \new_[40605]_ , \new_[40609]_ , \new_[40610]_ , \new_[40611]_ ,
    \new_[40615]_ , \new_[40616]_ , \new_[40619]_ , \new_[40622]_ ,
    \new_[40623]_ , \new_[40624]_ , \new_[40628]_ , \new_[40629]_ ,
    \new_[40633]_ , \new_[40634]_ , \new_[40635]_ , \new_[40639]_ ,
    \new_[40640]_ , \new_[40643]_ , \new_[40646]_ , \new_[40647]_ ,
    \new_[40648]_ , \new_[40652]_ , \new_[40653]_ , \new_[40657]_ ,
    \new_[40658]_ , \new_[40659]_ , \new_[40663]_ , \new_[40664]_ ,
    \new_[40667]_ , \new_[40670]_ , \new_[40671]_ , \new_[40672]_ ,
    \new_[40676]_ , \new_[40677]_ , \new_[40681]_ , \new_[40682]_ ,
    \new_[40683]_ , \new_[40687]_ , \new_[40688]_ , \new_[40691]_ ,
    \new_[40694]_ , \new_[40695]_ , \new_[40696]_ , \new_[40700]_ ,
    \new_[40701]_ , \new_[40705]_ , \new_[40706]_ , \new_[40707]_ ,
    \new_[40711]_ , \new_[40712]_ , \new_[40715]_ , \new_[40718]_ ,
    \new_[40719]_ , \new_[40720]_ , \new_[40724]_ , \new_[40725]_ ,
    \new_[40729]_ , \new_[40730]_ , \new_[40731]_ , \new_[40735]_ ,
    \new_[40736]_ , \new_[40739]_ , \new_[40742]_ , \new_[40743]_ ,
    \new_[40744]_ , \new_[40748]_ , \new_[40749]_ , \new_[40753]_ ,
    \new_[40754]_ , \new_[40755]_ , \new_[40759]_ , \new_[40760]_ ,
    \new_[40763]_ , \new_[40766]_ , \new_[40767]_ , \new_[40768]_ ,
    \new_[40772]_ , \new_[40773]_ , \new_[40777]_ , \new_[40778]_ ,
    \new_[40779]_ , \new_[40783]_ , \new_[40784]_ , \new_[40787]_ ,
    \new_[40790]_ , \new_[40791]_ , \new_[40792]_ , \new_[40796]_ ,
    \new_[40797]_ , \new_[40801]_ , \new_[40802]_ , \new_[40803]_ ,
    \new_[40807]_ , \new_[40808]_ , \new_[40811]_ , \new_[40814]_ ,
    \new_[40815]_ , \new_[40816]_ , \new_[40820]_ , \new_[40821]_ ,
    \new_[40825]_ , \new_[40826]_ , \new_[40827]_ , \new_[40831]_ ,
    \new_[40832]_ , \new_[40835]_ , \new_[40838]_ , \new_[40839]_ ,
    \new_[40840]_ , \new_[40844]_ , \new_[40845]_ , \new_[40849]_ ,
    \new_[40850]_ , \new_[40851]_ , \new_[40855]_ , \new_[40856]_ ,
    \new_[40859]_ , \new_[40862]_ , \new_[40863]_ , \new_[40864]_ ,
    \new_[40868]_ , \new_[40869]_ , \new_[40873]_ , \new_[40874]_ ,
    \new_[40875]_ , \new_[40879]_ , \new_[40880]_ , \new_[40883]_ ,
    \new_[40886]_ , \new_[40887]_ , \new_[40888]_ , \new_[40892]_ ,
    \new_[40893]_ , \new_[40897]_ , \new_[40898]_ , \new_[40899]_ ,
    \new_[40903]_ , \new_[40904]_ , \new_[40907]_ , \new_[40910]_ ,
    \new_[40911]_ , \new_[40912]_ , \new_[40916]_ , \new_[40917]_ ,
    \new_[40921]_ , \new_[40922]_ , \new_[40923]_ , \new_[40927]_ ,
    \new_[40928]_ , \new_[40931]_ , \new_[40934]_ , \new_[40935]_ ,
    \new_[40936]_ , \new_[40940]_ , \new_[40941]_ , \new_[40945]_ ,
    \new_[40946]_ , \new_[40947]_ , \new_[40951]_ , \new_[40952]_ ,
    \new_[40955]_ , \new_[40958]_ , \new_[40959]_ , \new_[40960]_ ,
    \new_[40964]_ , \new_[40965]_ , \new_[40969]_ , \new_[40970]_ ,
    \new_[40971]_ , \new_[40975]_ , \new_[40976]_ , \new_[40979]_ ,
    \new_[40982]_ , \new_[40983]_ , \new_[40984]_ , \new_[40988]_ ,
    \new_[40989]_ , \new_[40993]_ , \new_[40994]_ , \new_[40995]_ ,
    \new_[40999]_ , \new_[41000]_ , \new_[41003]_ , \new_[41006]_ ,
    \new_[41007]_ , \new_[41008]_ , \new_[41012]_ , \new_[41013]_ ,
    \new_[41017]_ , \new_[41018]_ , \new_[41019]_ , \new_[41023]_ ,
    \new_[41024]_ , \new_[41027]_ , \new_[41030]_ , \new_[41031]_ ,
    \new_[41032]_ , \new_[41036]_ , \new_[41037]_ , \new_[41041]_ ,
    \new_[41042]_ , \new_[41043]_ , \new_[41047]_ , \new_[41048]_ ,
    \new_[41051]_ , \new_[41054]_ , \new_[41055]_ , \new_[41056]_ ,
    \new_[41060]_ , \new_[41061]_ , \new_[41065]_ , \new_[41066]_ ,
    \new_[41067]_ , \new_[41071]_ , \new_[41072]_ , \new_[41075]_ ,
    \new_[41078]_ , \new_[41079]_ , \new_[41080]_ , \new_[41084]_ ,
    \new_[41085]_ , \new_[41089]_ , \new_[41090]_ , \new_[41091]_ ,
    \new_[41095]_ , \new_[41096]_ , \new_[41099]_ , \new_[41102]_ ,
    \new_[41103]_ , \new_[41104]_ , \new_[41108]_ , \new_[41109]_ ,
    \new_[41113]_ , \new_[41114]_ , \new_[41115]_ , \new_[41119]_ ,
    \new_[41120]_ , \new_[41123]_ , \new_[41126]_ , \new_[41127]_ ,
    \new_[41128]_ , \new_[41132]_ , \new_[41133]_ , \new_[41137]_ ,
    \new_[41138]_ , \new_[41139]_ , \new_[41143]_ , \new_[41144]_ ,
    \new_[41147]_ , \new_[41150]_ , \new_[41151]_ , \new_[41152]_ ,
    \new_[41156]_ , \new_[41157]_ , \new_[41161]_ , \new_[41162]_ ,
    \new_[41163]_ , \new_[41167]_ , \new_[41168]_ , \new_[41171]_ ,
    \new_[41174]_ , \new_[41175]_ , \new_[41176]_ , \new_[41180]_ ,
    \new_[41181]_ , \new_[41185]_ , \new_[41186]_ , \new_[41187]_ ,
    \new_[41191]_ , \new_[41192]_ , \new_[41195]_ , \new_[41198]_ ,
    \new_[41199]_ , \new_[41200]_ , \new_[41204]_ , \new_[41205]_ ,
    \new_[41209]_ , \new_[41210]_ , \new_[41211]_ , \new_[41215]_ ,
    \new_[41216]_ , \new_[41219]_ , \new_[41222]_ , \new_[41223]_ ,
    \new_[41224]_ , \new_[41228]_ , \new_[41229]_ , \new_[41233]_ ,
    \new_[41234]_ , \new_[41235]_ , \new_[41239]_ , \new_[41240]_ ,
    \new_[41243]_ , \new_[41246]_ , \new_[41247]_ , \new_[41248]_ ,
    \new_[41252]_ , \new_[41253]_ , \new_[41257]_ , \new_[41258]_ ,
    \new_[41259]_ , \new_[41263]_ , \new_[41264]_ , \new_[41267]_ ,
    \new_[41270]_ , \new_[41271]_ , \new_[41272]_ , \new_[41276]_ ,
    \new_[41277]_ , \new_[41281]_ , \new_[41282]_ , \new_[41283]_ ,
    \new_[41287]_ , \new_[41288]_ , \new_[41291]_ , \new_[41294]_ ,
    \new_[41295]_ , \new_[41296]_ , \new_[41300]_ , \new_[41301]_ ,
    \new_[41305]_ , \new_[41306]_ , \new_[41307]_ , \new_[41311]_ ,
    \new_[41312]_ , \new_[41315]_ , \new_[41318]_ , \new_[41319]_ ,
    \new_[41320]_ , \new_[41324]_ , \new_[41325]_ , \new_[41329]_ ,
    \new_[41330]_ , \new_[41331]_ , \new_[41335]_ , \new_[41336]_ ,
    \new_[41339]_ , \new_[41342]_ , \new_[41343]_ , \new_[41344]_ ,
    \new_[41348]_ , \new_[41349]_ , \new_[41353]_ , \new_[41354]_ ,
    \new_[41355]_ , \new_[41359]_ , \new_[41360]_ , \new_[41363]_ ,
    \new_[41366]_ , \new_[41367]_ , \new_[41368]_ , \new_[41372]_ ,
    \new_[41373]_ , \new_[41377]_ , \new_[41378]_ , \new_[41379]_ ,
    \new_[41383]_ , \new_[41384]_ , \new_[41387]_ , \new_[41390]_ ,
    \new_[41391]_ , \new_[41392]_ , \new_[41396]_ , \new_[41397]_ ,
    \new_[41401]_ , \new_[41402]_ , \new_[41403]_ , \new_[41407]_ ,
    \new_[41408]_ , \new_[41411]_ , \new_[41414]_ , \new_[41415]_ ,
    \new_[41416]_ , \new_[41420]_ , \new_[41421]_ , \new_[41425]_ ,
    \new_[41426]_ , \new_[41427]_ , \new_[41431]_ , \new_[41432]_ ,
    \new_[41435]_ , \new_[41438]_ , \new_[41439]_ , \new_[41440]_ ,
    \new_[41444]_ , \new_[41445]_ , \new_[41449]_ , \new_[41450]_ ,
    \new_[41451]_ , \new_[41455]_ , \new_[41456]_ , \new_[41459]_ ,
    \new_[41462]_ , \new_[41463]_ , \new_[41464]_ , \new_[41468]_ ,
    \new_[41469]_ , \new_[41473]_ , \new_[41474]_ , \new_[41475]_ ,
    \new_[41479]_ , \new_[41480]_ , \new_[41483]_ , \new_[41486]_ ,
    \new_[41487]_ , \new_[41488]_ , \new_[41492]_ , \new_[41493]_ ,
    \new_[41497]_ , \new_[41498]_ , \new_[41499]_ , \new_[41503]_ ,
    \new_[41504]_ , \new_[41507]_ , \new_[41510]_ , \new_[41511]_ ,
    \new_[41512]_ , \new_[41516]_ , \new_[41517]_ , \new_[41521]_ ,
    \new_[41522]_ , \new_[41523]_ , \new_[41527]_ , \new_[41528]_ ,
    \new_[41531]_ , \new_[41534]_ , \new_[41535]_ , \new_[41536]_ ,
    \new_[41540]_ , \new_[41541]_ , \new_[41545]_ , \new_[41546]_ ,
    \new_[41547]_ , \new_[41551]_ , \new_[41552]_ , \new_[41555]_ ,
    \new_[41558]_ , \new_[41559]_ , \new_[41560]_ , \new_[41564]_ ,
    \new_[41565]_ , \new_[41569]_ , \new_[41570]_ , \new_[41571]_ ,
    \new_[41575]_ , \new_[41576]_ , \new_[41579]_ , \new_[41582]_ ,
    \new_[41583]_ , \new_[41584]_ , \new_[41588]_ , \new_[41589]_ ,
    \new_[41593]_ , \new_[41594]_ , \new_[41595]_ , \new_[41599]_ ,
    \new_[41600]_ , \new_[41603]_ , \new_[41606]_ , \new_[41607]_ ,
    \new_[41608]_ , \new_[41612]_ , \new_[41613]_ , \new_[41617]_ ,
    \new_[41618]_ , \new_[41619]_ , \new_[41623]_ , \new_[41624]_ ,
    \new_[41627]_ , \new_[41630]_ , \new_[41631]_ , \new_[41632]_ ,
    \new_[41636]_ , \new_[41637]_ , \new_[41641]_ , \new_[41642]_ ,
    \new_[41643]_ , \new_[41647]_ , \new_[41648]_ , \new_[41651]_ ,
    \new_[41654]_ , \new_[41655]_ , \new_[41656]_ , \new_[41660]_ ,
    \new_[41661]_ , \new_[41665]_ , \new_[41666]_ , \new_[41667]_ ,
    \new_[41671]_ , \new_[41672]_ , \new_[41675]_ , \new_[41678]_ ,
    \new_[41679]_ , \new_[41680]_ , \new_[41684]_ , \new_[41685]_ ,
    \new_[41689]_ , \new_[41690]_ , \new_[41691]_ , \new_[41695]_ ,
    \new_[41696]_ , \new_[41699]_ , \new_[41702]_ , \new_[41703]_ ,
    \new_[41704]_ , \new_[41708]_ , \new_[41709]_ , \new_[41713]_ ,
    \new_[41714]_ , \new_[41715]_ , \new_[41719]_ , \new_[41720]_ ,
    \new_[41723]_ , \new_[41726]_ , \new_[41727]_ , \new_[41728]_ ,
    \new_[41732]_ , \new_[41733]_ , \new_[41737]_ , \new_[41738]_ ,
    \new_[41739]_ , \new_[41743]_ , \new_[41744]_ , \new_[41747]_ ,
    \new_[41750]_ , \new_[41751]_ , \new_[41752]_ , \new_[41756]_ ,
    \new_[41757]_ , \new_[41761]_ , \new_[41762]_ , \new_[41763]_ ,
    \new_[41767]_ , \new_[41768]_ , \new_[41771]_ , \new_[41774]_ ,
    \new_[41775]_ , \new_[41776]_ , \new_[41780]_ , \new_[41781]_ ,
    \new_[41785]_ , \new_[41786]_ , \new_[41787]_ , \new_[41791]_ ,
    \new_[41792]_ , \new_[41795]_ , \new_[41798]_ , \new_[41799]_ ,
    \new_[41800]_ , \new_[41804]_ , \new_[41805]_ , \new_[41809]_ ,
    \new_[41810]_ , \new_[41811]_ , \new_[41815]_ , \new_[41816]_ ,
    \new_[41819]_ , \new_[41822]_ , \new_[41823]_ , \new_[41824]_ ,
    \new_[41828]_ , \new_[41829]_ , \new_[41833]_ , \new_[41834]_ ,
    \new_[41835]_ , \new_[41839]_ , \new_[41840]_ , \new_[41843]_ ,
    \new_[41846]_ , \new_[41847]_ , \new_[41848]_ , \new_[41852]_ ,
    \new_[41853]_ , \new_[41857]_ , \new_[41858]_ , \new_[41859]_ ,
    \new_[41863]_ , \new_[41864]_ , \new_[41867]_ , \new_[41870]_ ,
    \new_[41871]_ , \new_[41872]_ , \new_[41876]_ , \new_[41877]_ ,
    \new_[41881]_ , \new_[41882]_ , \new_[41883]_ , \new_[41887]_ ,
    \new_[41888]_ , \new_[41891]_ , \new_[41894]_ , \new_[41895]_ ,
    \new_[41896]_ , \new_[41900]_ , \new_[41901]_ , \new_[41905]_ ,
    \new_[41906]_ , \new_[41907]_ , \new_[41911]_ , \new_[41912]_ ,
    \new_[41915]_ , \new_[41918]_ , \new_[41919]_ , \new_[41920]_ ,
    \new_[41924]_ , \new_[41925]_ , \new_[41929]_ , \new_[41930]_ ,
    \new_[41931]_ , \new_[41935]_ , \new_[41936]_ , \new_[41939]_ ,
    \new_[41942]_ , \new_[41943]_ , \new_[41944]_ , \new_[41948]_ ,
    \new_[41949]_ , \new_[41953]_ , \new_[41954]_ , \new_[41955]_ ,
    \new_[41959]_ , \new_[41960]_ , \new_[41963]_ , \new_[41966]_ ,
    \new_[41967]_ , \new_[41968]_ , \new_[41972]_ , \new_[41973]_ ,
    \new_[41977]_ , \new_[41978]_ , \new_[41979]_ , \new_[41983]_ ,
    \new_[41984]_ , \new_[41987]_ , \new_[41990]_ , \new_[41991]_ ,
    \new_[41992]_ , \new_[41996]_ , \new_[41997]_ , \new_[42001]_ ,
    \new_[42002]_ , \new_[42003]_ , \new_[42007]_ , \new_[42008]_ ,
    \new_[42011]_ , \new_[42014]_ , \new_[42015]_ , \new_[42016]_ ,
    \new_[42020]_ , \new_[42021]_ , \new_[42025]_ , \new_[42026]_ ,
    \new_[42027]_ , \new_[42031]_ , \new_[42032]_ , \new_[42035]_ ,
    \new_[42038]_ , \new_[42039]_ , \new_[42040]_ , \new_[42044]_ ,
    \new_[42045]_ , \new_[42049]_ , \new_[42050]_ , \new_[42051]_ ,
    \new_[42055]_ , \new_[42056]_ , \new_[42059]_ , \new_[42062]_ ,
    \new_[42063]_ , \new_[42064]_ , \new_[42068]_ , \new_[42069]_ ,
    \new_[42073]_ , \new_[42074]_ , \new_[42075]_ , \new_[42079]_ ,
    \new_[42080]_ , \new_[42083]_ , \new_[42086]_ , \new_[42087]_ ,
    \new_[42088]_ , \new_[42092]_ , \new_[42093]_ , \new_[42097]_ ,
    \new_[42098]_ , \new_[42099]_ , \new_[42103]_ , \new_[42104]_ ,
    \new_[42107]_ , \new_[42110]_ , \new_[42111]_ , \new_[42112]_ ,
    \new_[42116]_ , \new_[42117]_ , \new_[42121]_ , \new_[42122]_ ,
    \new_[42123]_ , \new_[42127]_ , \new_[42128]_ , \new_[42131]_ ,
    \new_[42134]_ , \new_[42135]_ , \new_[42136]_ , \new_[42140]_ ,
    \new_[42141]_ , \new_[42145]_ , \new_[42146]_ , \new_[42147]_ ,
    \new_[42151]_ , \new_[42152]_ , \new_[42155]_ , \new_[42158]_ ,
    \new_[42159]_ , \new_[42160]_ , \new_[42164]_ , \new_[42165]_ ,
    \new_[42169]_ , \new_[42170]_ , \new_[42171]_ , \new_[42175]_ ,
    \new_[42176]_ , \new_[42179]_ , \new_[42182]_ , \new_[42183]_ ,
    \new_[42184]_ , \new_[42188]_ , \new_[42189]_ , \new_[42193]_ ,
    \new_[42194]_ , \new_[42195]_ , \new_[42199]_ , \new_[42200]_ ,
    \new_[42203]_ , \new_[42206]_ , \new_[42207]_ , \new_[42208]_ ,
    \new_[42212]_ , \new_[42213]_ , \new_[42217]_ , \new_[42218]_ ,
    \new_[42219]_ , \new_[42223]_ , \new_[42224]_ , \new_[42227]_ ,
    \new_[42230]_ , \new_[42231]_ , \new_[42232]_ , \new_[42236]_ ,
    \new_[42237]_ , \new_[42241]_ , \new_[42242]_ , \new_[42243]_ ,
    \new_[42247]_ , \new_[42248]_ , \new_[42251]_ , \new_[42254]_ ,
    \new_[42255]_ , \new_[42256]_ , \new_[42260]_ , \new_[42261]_ ,
    \new_[42265]_ , \new_[42266]_ , \new_[42267]_ , \new_[42271]_ ,
    \new_[42272]_ , \new_[42275]_ , \new_[42278]_ , \new_[42279]_ ,
    \new_[42280]_ , \new_[42284]_ , \new_[42285]_ , \new_[42289]_ ,
    \new_[42290]_ , \new_[42291]_ , \new_[42295]_ , \new_[42296]_ ,
    \new_[42299]_ , \new_[42302]_ , \new_[42303]_ , \new_[42304]_ ,
    \new_[42308]_ , \new_[42309]_ , \new_[42313]_ , \new_[42314]_ ,
    \new_[42315]_ , \new_[42319]_ , \new_[42320]_ , \new_[42323]_ ,
    \new_[42326]_ , \new_[42327]_ , \new_[42328]_ , \new_[42332]_ ,
    \new_[42333]_ , \new_[42337]_ , \new_[42338]_ , \new_[42339]_ ,
    \new_[42343]_ , \new_[42344]_ , \new_[42347]_ , \new_[42350]_ ,
    \new_[42351]_ , \new_[42352]_ , \new_[42356]_ , \new_[42357]_ ,
    \new_[42361]_ , \new_[42362]_ , \new_[42363]_ , \new_[42367]_ ,
    \new_[42368]_ , \new_[42371]_ , \new_[42374]_ , \new_[42375]_ ,
    \new_[42376]_ , \new_[42380]_ , \new_[42381]_ , \new_[42385]_ ,
    \new_[42386]_ , \new_[42387]_ , \new_[42391]_ , \new_[42392]_ ,
    \new_[42395]_ , \new_[42398]_ , \new_[42399]_ , \new_[42400]_ ,
    \new_[42404]_ , \new_[42405]_ , \new_[42409]_ , \new_[42410]_ ,
    \new_[42411]_ , \new_[42415]_ , \new_[42416]_ , \new_[42419]_ ,
    \new_[42422]_ , \new_[42423]_ , \new_[42424]_ , \new_[42428]_ ,
    \new_[42429]_ , \new_[42433]_ , \new_[42434]_ , \new_[42435]_ ,
    \new_[42439]_ , \new_[42440]_ , \new_[42443]_ , \new_[42446]_ ,
    \new_[42447]_ , \new_[42448]_ , \new_[42452]_ , \new_[42453]_ ,
    \new_[42457]_ , \new_[42458]_ , \new_[42459]_ , \new_[42463]_ ,
    \new_[42464]_ , \new_[42467]_ , \new_[42470]_ , \new_[42471]_ ,
    \new_[42472]_ , \new_[42476]_ , \new_[42477]_ , \new_[42481]_ ,
    \new_[42482]_ , \new_[42483]_ , \new_[42487]_ , \new_[42488]_ ,
    \new_[42491]_ , \new_[42494]_ , \new_[42495]_ , \new_[42496]_ ,
    \new_[42500]_ , \new_[42501]_ , \new_[42505]_ , \new_[42506]_ ,
    \new_[42507]_ , \new_[42511]_ , \new_[42512]_ , \new_[42515]_ ,
    \new_[42518]_ , \new_[42519]_ , \new_[42520]_ , \new_[42524]_ ,
    \new_[42525]_ , \new_[42529]_ , \new_[42530]_ , \new_[42531]_ ,
    \new_[42535]_ , \new_[42536]_ , \new_[42539]_ , \new_[42542]_ ,
    \new_[42543]_ , \new_[42544]_ , \new_[42548]_ , \new_[42549]_ ,
    \new_[42553]_ , \new_[42554]_ , \new_[42555]_ , \new_[42559]_ ,
    \new_[42560]_ , \new_[42563]_ , \new_[42566]_ , \new_[42567]_ ,
    \new_[42568]_ , \new_[42572]_ , \new_[42573]_ , \new_[42577]_ ,
    \new_[42578]_ , \new_[42579]_ , \new_[42583]_ , \new_[42584]_ ,
    \new_[42587]_ , \new_[42590]_ , \new_[42591]_ , \new_[42592]_ ,
    \new_[42596]_ , \new_[42597]_ , \new_[42601]_ , \new_[42602]_ ,
    \new_[42603]_ , \new_[42607]_ , \new_[42608]_ , \new_[42611]_ ,
    \new_[42614]_ , \new_[42615]_ , \new_[42616]_ , \new_[42620]_ ,
    \new_[42621]_ , \new_[42625]_ , \new_[42626]_ , \new_[42627]_ ,
    \new_[42631]_ , \new_[42632]_ , \new_[42635]_ , \new_[42638]_ ,
    \new_[42639]_ , \new_[42640]_ , \new_[42644]_ , \new_[42645]_ ,
    \new_[42649]_ , \new_[42650]_ , \new_[42651]_ , \new_[42655]_ ,
    \new_[42656]_ , \new_[42659]_ , \new_[42662]_ , \new_[42663]_ ,
    \new_[42664]_ , \new_[42668]_ , \new_[42669]_ , \new_[42673]_ ,
    \new_[42674]_ , \new_[42675]_ , \new_[42679]_ , \new_[42680]_ ,
    \new_[42683]_ , \new_[42686]_ , \new_[42687]_ , \new_[42688]_ ,
    \new_[42692]_ , \new_[42693]_ , \new_[42697]_ , \new_[42698]_ ,
    \new_[42699]_ , \new_[42703]_ , \new_[42704]_ , \new_[42707]_ ,
    \new_[42710]_ , \new_[42711]_ , \new_[42712]_ , \new_[42716]_ ,
    \new_[42717]_ , \new_[42721]_ , \new_[42722]_ , \new_[42723]_ ,
    \new_[42727]_ , \new_[42728]_ , \new_[42731]_ , \new_[42734]_ ,
    \new_[42735]_ , \new_[42736]_ , \new_[42740]_ , \new_[42741]_ ,
    \new_[42745]_ , \new_[42746]_ , \new_[42747]_ , \new_[42751]_ ,
    \new_[42752]_ , \new_[42755]_ , \new_[42758]_ , \new_[42759]_ ,
    \new_[42760]_ , \new_[42764]_ , \new_[42765]_ , \new_[42769]_ ,
    \new_[42770]_ , \new_[42771]_ , \new_[42775]_ , \new_[42776]_ ,
    \new_[42779]_ , \new_[42782]_ , \new_[42783]_ , \new_[42784]_ ,
    \new_[42788]_ , \new_[42789]_ , \new_[42793]_ , \new_[42794]_ ,
    \new_[42795]_ , \new_[42799]_ , \new_[42800]_ , \new_[42803]_ ,
    \new_[42806]_ , \new_[42807]_ , \new_[42808]_ , \new_[42812]_ ,
    \new_[42813]_ , \new_[42817]_ , \new_[42818]_ , \new_[42819]_ ,
    \new_[42823]_ , \new_[42824]_ , \new_[42827]_ , \new_[42830]_ ,
    \new_[42831]_ , \new_[42832]_ , \new_[42836]_ , \new_[42837]_ ,
    \new_[42841]_ , \new_[42842]_ , \new_[42843]_ , \new_[42847]_ ,
    \new_[42848]_ , \new_[42851]_ , \new_[42854]_ , \new_[42855]_ ,
    \new_[42856]_ , \new_[42860]_ , \new_[42861]_ , \new_[42865]_ ,
    \new_[42866]_ , \new_[42867]_ , \new_[42871]_ , \new_[42872]_ ,
    \new_[42875]_ , \new_[42878]_ , \new_[42879]_ , \new_[42880]_ ,
    \new_[42884]_ , \new_[42885]_ , \new_[42889]_ , \new_[42890]_ ,
    \new_[42891]_ , \new_[42895]_ , \new_[42896]_ , \new_[42899]_ ,
    \new_[42902]_ , \new_[42903]_ , \new_[42904]_ , \new_[42908]_ ,
    \new_[42909]_ , \new_[42913]_ , \new_[42914]_ , \new_[42915]_ ,
    \new_[42919]_ , \new_[42920]_ , \new_[42923]_ , \new_[42926]_ ,
    \new_[42927]_ , \new_[42928]_ , \new_[42932]_ , \new_[42933]_ ,
    \new_[42937]_ , \new_[42938]_ , \new_[42939]_ , \new_[42943]_ ,
    \new_[42944]_ , \new_[42947]_ , \new_[42950]_ , \new_[42951]_ ,
    \new_[42952]_ , \new_[42956]_ , \new_[42957]_ , \new_[42961]_ ,
    \new_[42962]_ , \new_[42963]_ , \new_[42967]_ , \new_[42968]_ ,
    \new_[42971]_ , \new_[42974]_ , \new_[42975]_ , \new_[42976]_ ,
    \new_[42980]_ , \new_[42981]_ , \new_[42985]_ , \new_[42986]_ ,
    \new_[42987]_ , \new_[42991]_ , \new_[42992]_ , \new_[42995]_ ,
    \new_[42998]_ , \new_[42999]_ , \new_[43000]_ , \new_[43004]_ ,
    \new_[43005]_ , \new_[43009]_ , \new_[43010]_ , \new_[43011]_ ,
    \new_[43015]_ , \new_[43016]_ , \new_[43019]_ , \new_[43022]_ ,
    \new_[43023]_ , \new_[43024]_ , \new_[43028]_ , \new_[43029]_ ,
    \new_[43033]_ , \new_[43034]_ , \new_[43035]_ , \new_[43039]_ ,
    \new_[43040]_ , \new_[43043]_ , \new_[43046]_ , \new_[43047]_ ,
    \new_[43048]_ , \new_[43052]_ , \new_[43053]_ , \new_[43057]_ ,
    \new_[43058]_ , \new_[43059]_ , \new_[43063]_ , \new_[43064]_ ,
    \new_[43067]_ , \new_[43070]_ , \new_[43071]_ , \new_[43072]_ ,
    \new_[43076]_ , \new_[43077]_ , \new_[43081]_ , \new_[43082]_ ,
    \new_[43083]_ , \new_[43087]_ , \new_[43088]_ , \new_[43091]_ ,
    \new_[43094]_ , \new_[43095]_ , \new_[43096]_ , \new_[43100]_ ,
    \new_[43101]_ , \new_[43105]_ , \new_[43106]_ , \new_[43107]_ ,
    \new_[43111]_ , \new_[43112]_ , \new_[43115]_ , \new_[43118]_ ,
    \new_[43119]_ , \new_[43120]_ , \new_[43124]_ , \new_[43125]_ ,
    \new_[43129]_ , \new_[43130]_ , \new_[43131]_ , \new_[43135]_ ,
    \new_[43136]_ , \new_[43139]_ , \new_[43142]_ , \new_[43143]_ ,
    \new_[43144]_ , \new_[43148]_ , \new_[43149]_ , \new_[43153]_ ,
    \new_[43154]_ , \new_[43155]_ , \new_[43159]_ , \new_[43160]_ ,
    \new_[43163]_ , \new_[43166]_ , \new_[43167]_ , \new_[43168]_ ,
    \new_[43172]_ , \new_[43173]_ , \new_[43177]_ , \new_[43178]_ ,
    \new_[43179]_ , \new_[43183]_ , \new_[43184]_ , \new_[43187]_ ,
    \new_[43190]_ , \new_[43191]_ , \new_[43192]_ , \new_[43196]_ ,
    \new_[43197]_ , \new_[43201]_ , \new_[43202]_ , \new_[43203]_ ,
    \new_[43207]_ , \new_[43208]_ , \new_[43211]_ , \new_[43214]_ ,
    \new_[43215]_ , \new_[43216]_ , \new_[43220]_ , \new_[43221]_ ,
    \new_[43225]_ , \new_[43226]_ , \new_[43227]_ , \new_[43231]_ ,
    \new_[43232]_ , \new_[43235]_ , \new_[43238]_ , \new_[43239]_ ,
    \new_[43240]_ , \new_[43244]_ , \new_[43245]_ , \new_[43249]_ ,
    \new_[43250]_ , \new_[43251]_ , \new_[43255]_ , \new_[43256]_ ,
    \new_[43259]_ , \new_[43262]_ , \new_[43263]_ , \new_[43264]_ ,
    \new_[43268]_ , \new_[43269]_ , \new_[43273]_ , \new_[43274]_ ,
    \new_[43275]_ , \new_[43279]_ , \new_[43280]_ , \new_[43283]_ ,
    \new_[43286]_ , \new_[43287]_ , \new_[43288]_ , \new_[43292]_ ,
    \new_[43293]_ , \new_[43297]_ , \new_[43298]_ , \new_[43299]_ ,
    \new_[43303]_ , \new_[43304]_ , \new_[43307]_ , \new_[43310]_ ,
    \new_[43311]_ , \new_[43312]_ , \new_[43316]_ , \new_[43317]_ ,
    \new_[43321]_ , \new_[43322]_ , \new_[43323]_ , \new_[43327]_ ,
    \new_[43328]_ , \new_[43331]_ , \new_[43334]_ , \new_[43335]_ ,
    \new_[43336]_ , \new_[43340]_ , \new_[43341]_ , \new_[43345]_ ,
    \new_[43346]_ , \new_[43347]_ , \new_[43351]_ , \new_[43352]_ ,
    \new_[43355]_ , \new_[43358]_ , \new_[43359]_ , \new_[43360]_ ,
    \new_[43364]_ , \new_[43365]_ , \new_[43369]_ , \new_[43370]_ ,
    \new_[43371]_ , \new_[43375]_ , \new_[43376]_ , \new_[43379]_ ,
    \new_[43382]_ , \new_[43383]_ , \new_[43384]_ , \new_[43388]_ ,
    \new_[43389]_ , \new_[43393]_ , \new_[43394]_ , \new_[43395]_ ,
    \new_[43399]_ , \new_[43400]_ , \new_[43403]_ , \new_[43406]_ ,
    \new_[43407]_ , \new_[43408]_ , \new_[43412]_ , \new_[43413]_ ,
    \new_[43417]_ , \new_[43418]_ , \new_[43419]_ , \new_[43423]_ ,
    \new_[43424]_ , \new_[43427]_ , \new_[43430]_ , \new_[43431]_ ,
    \new_[43432]_ , \new_[43436]_ , \new_[43437]_ , \new_[43441]_ ,
    \new_[43442]_ , \new_[43443]_ , \new_[43447]_ , \new_[43448]_ ,
    \new_[43451]_ , \new_[43454]_ , \new_[43455]_ , \new_[43456]_ ,
    \new_[43460]_ , \new_[43461]_ , \new_[43465]_ , \new_[43466]_ ,
    \new_[43467]_ , \new_[43471]_ , \new_[43472]_ , \new_[43475]_ ,
    \new_[43478]_ , \new_[43479]_ , \new_[43480]_ , \new_[43484]_ ,
    \new_[43485]_ , \new_[43489]_ , \new_[43490]_ , \new_[43491]_ ,
    \new_[43495]_ , \new_[43496]_ , \new_[43499]_ , \new_[43502]_ ,
    \new_[43503]_ , \new_[43504]_ , \new_[43508]_ , \new_[43509]_ ,
    \new_[43513]_ , \new_[43514]_ , \new_[43515]_ , \new_[43519]_ ,
    \new_[43520]_ , \new_[43523]_ , \new_[43526]_ , \new_[43527]_ ,
    \new_[43528]_ , \new_[43532]_ , \new_[43533]_ , \new_[43537]_ ,
    \new_[43538]_ , \new_[43539]_ , \new_[43543]_ , \new_[43544]_ ,
    \new_[43547]_ , \new_[43550]_ , \new_[43551]_ , \new_[43552]_ ,
    \new_[43556]_ , \new_[43557]_ , \new_[43561]_ , \new_[43562]_ ,
    \new_[43563]_ , \new_[43567]_ , \new_[43568]_ , \new_[43571]_ ,
    \new_[43574]_ , \new_[43575]_ , \new_[43576]_ , \new_[43580]_ ,
    \new_[43581]_ , \new_[43585]_ , \new_[43586]_ , \new_[43587]_ ,
    \new_[43591]_ , \new_[43592]_ , \new_[43595]_ , \new_[43598]_ ,
    \new_[43599]_ , \new_[43600]_ , \new_[43604]_ , \new_[43605]_ ,
    \new_[43609]_ , \new_[43610]_ , \new_[43611]_ , \new_[43615]_ ,
    \new_[43616]_ , \new_[43619]_ , \new_[43622]_ , \new_[43623]_ ,
    \new_[43624]_ , \new_[43628]_ , \new_[43629]_ , \new_[43633]_ ,
    \new_[43634]_ , \new_[43635]_ , \new_[43639]_ , \new_[43640]_ ,
    \new_[43643]_ , \new_[43646]_ , \new_[43647]_ , \new_[43648]_ ,
    \new_[43652]_ , \new_[43653]_ , \new_[43657]_ , \new_[43658]_ ,
    \new_[43659]_ , \new_[43663]_ , \new_[43664]_ , \new_[43667]_ ,
    \new_[43670]_ , \new_[43671]_ , \new_[43672]_ , \new_[43676]_ ,
    \new_[43677]_ , \new_[43681]_ , \new_[43682]_ , \new_[43683]_ ,
    \new_[43687]_ , \new_[43688]_ , \new_[43691]_ , \new_[43694]_ ,
    \new_[43695]_ , \new_[43696]_ , \new_[43700]_ , \new_[43701]_ ,
    \new_[43705]_ , \new_[43706]_ , \new_[43707]_ , \new_[43711]_ ,
    \new_[43712]_ , \new_[43715]_ , \new_[43718]_ , \new_[43719]_ ,
    \new_[43720]_ , \new_[43724]_ , \new_[43725]_ , \new_[43729]_ ,
    \new_[43730]_ , \new_[43731]_ , \new_[43735]_ , \new_[43736]_ ,
    \new_[43739]_ , \new_[43742]_ , \new_[43743]_ , \new_[43744]_ ,
    \new_[43748]_ , \new_[43749]_ , \new_[43753]_ , \new_[43754]_ ,
    \new_[43755]_ , \new_[43759]_ , \new_[43760]_ , \new_[43763]_ ,
    \new_[43766]_ , \new_[43767]_ , \new_[43768]_ , \new_[43772]_ ,
    \new_[43773]_ , \new_[43777]_ , \new_[43778]_ , \new_[43779]_ ,
    \new_[43783]_ , \new_[43784]_ , \new_[43787]_ , \new_[43790]_ ,
    \new_[43791]_ , \new_[43792]_ , \new_[43796]_ , \new_[43797]_ ,
    \new_[43801]_ , \new_[43802]_ , \new_[43803]_ , \new_[43807]_ ,
    \new_[43808]_ , \new_[43811]_ , \new_[43814]_ , \new_[43815]_ ,
    \new_[43816]_ , \new_[43820]_ , \new_[43821]_ , \new_[43825]_ ,
    \new_[43826]_ , \new_[43827]_ , \new_[43831]_ , \new_[43832]_ ,
    \new_[43835]_ , \new_[43838]_ , \new_[43839]_ , \new_[43840]_ ,
    \new_[43844]_ , \new_[43845]_ , \new_[43849]_ , \new_[43850]_ ,
    \new_[43851]_ , \new_[43855]_ , \new_[43856]_ , \new_[43859]_ ,
    \new_[43862]_ , \new_[43863]_ , \new_[43864]_ , \new_[43868]_ ,
    \new_[43869]_ , \new_[43873]_ , \new_[43874]_ , \new_[43875]_ ,
    \new_[43879]_ , \new_[43880]_ , \new_[43883]_ , \new_[43886]_ ,
    \new_[43887]_ , \new_[43888]_ , \new_[43892]_ , \new_[43893]_ ,
    \new_[43897]_ , \new_[43898]_ , \new_[43899]_ , \new_[43903]_ ,
    \new_[43904]_ , \new_[43907]_ , \new_[43910]_ , \new_[43911]_ ,
    \new_[43912]_ , \new_[43916]_ , \new_[43917]_ , \new_[43921]_ ,
    \new_[43922]_ , \new_[43923]_ , \new_[43927]_ , \new_[43928]_ ,
    \new_[43931]_ , \new_[43934]_ , \new_[43935]_ , \new_[43936]_ ,
    \new_[43940]_ , \new_[43941]_ , \new_[43945]_ , \new_[43946]_ ,
    \new_[43947]_ , \new_[43951]_ , \new_[43952]_ , \new_[43955]_ ,
    \new_[43958]_ , \new_[43959]_ , \new_[43960]_ , \new_[43964]_ ,
    \new_[43965]_ , \new_[43969]_ , \new_[43970]_ , \new_[43971]_ ,
    \new_[43975]_ , \new_[43976]_ , \new_[43979]_ , \new_[43982]_ ,
    \new_[43983]_ , \new_[43984]_ , \new_[43988]_ , \new_[43989]_ ,
    \new_[43993]_ , \new_[43994]_ , \new_[43995]_ , \new_[43999]_ ,
    \new_[44000]_ , \new_[44003]_ , \new_[44006]_ , \new_[44007]_ ,
    \new_[44008]_ , \new_[44012]_ , \new_[44013]_ , \new_[44017]_ ,
    \new_[44018]_ , \new_[44019]_ , \new_[44023]_ , \new_[44024]_ ,
    \new_[44027]_ , \new_[44030]_ , \new_[44031]_ , \new_[44032]_ ,
    \new_[44036]_ , \new_[44037]_ , \new_[44041]_ , \new_[44042]_ ,
    \new_[44043]_ , \new_[44047]_ , \new_[44048]_ , \new_[44051]_ ,
    \new_[44054]_ , \new_[44055]_ , \new_[44056]_ , \new_[44060]_ ,
    \new_[44061]_ , \new_[44065]_ , \new_[44066]_ , \new_[44067]_ ,
    \new_[44071]_ , \new_[44072]_ , \new_[44075]_ , \new_[44078]_ ,
    \new_[44079]_ , \new_[44080]_ , \new_[44084]_ , \new_[44085]_ ,
    \new_[44089]_ , \new_[44090]_ , \new_[44091]_ , \new_[44095]_ ,
    \new_[44096]_ , \new_[44099]_ , \new_[44102]_ , \new_[44103]_ ,
    \new_[44104]_ , \new_[44108]_ , \new_[44109]_ , \new_[44113]_ ,
    \new_[44114]_ , \new_[44115]_ , \new_[44119]_ , \new_[44120]_ ,
    \new_[44123]_ , \new_[44126]_ , \new_[44127]_ , \new_[44128]_ ,
    \new_[44132]_ , \new_[44133]_ , \new_[44137]_ , \new_[44138]_ ,
    \new_[44139]_ , \new_[44143]_ , \new_[44144]_ , \new_[44147]_ ,
    \new_[44150]_ , \new_[44151]_ , \new_[44152]_ , \new_[44156]_ ,
    \new_[44157]_ , \new_[44161]_ , \new_[44162]_ , \new_[44163]_ ,
    \new_[44167]_ , \new_[44168]_ , \new_[44171]_ , \new_[44174]_ ,
    \new_[44175]_ , \new_[44176]_ , \new_[44180]_ , \new_[44181]_ ,
    \new_[44185]_ , \new_[44186]_ , \new_[44187]_ , \new_[44191]_ ,
    \new_[44192]_ , \new_[44195]_ , \new_[44198]_ , \new_[44199]_ ,
    \new_[44200]_ , \new_[44204]_ , \new_[44205]_ , \new_[44209]_ ,
    \new_[44210]_ , \new_[44211]_ , \new_[44215]_ , \new_[44216]_ ,
    \new_[44219]_ , \new_[44222]_ , \new_[44223]_ , \new_[44224]_ ,
    \new_[44228]_ , \new_[44229]_ , \new_[44233]_ , \new_[44234]_ ,
    \new_[44235]_ , \new_[44239]_ , \new_[44240]_ , \new_[44243]_ ,
    \new_[44246]_ , \new_[44247]_ , \new_[44248]_ , \new_[44252]_ ,
    \new_[44253]_ , \new_[44257]_ , \new_[44258]_ , \new_[44259]_ ,
    \new_[44263]_ , \new_[44264]_ , \new_[44267]_ , \new_[44270]_ ,
    \new_[44271]_ , \new_[44272]_ , \new_[44276]_ , \new_[44277]_ ,
    \new_[44281]_ , \new_[44282]_ , \new_[44283]_ , \new_[44287]_ ,
    \new_[44288]_ , \new_[44291]_ , \new_[44294]_ , \new_[44295]_ ,
    \new_[44296]_ , \new_[44300]_ , \new_[44301]_ , \new_[44305]_ ,
    \new_[44306]_ , \new_[44307]_ , \new_[44311]_ , \new_[44312]_ ,
    \new_[44315]_ , \new_[44318]_ , \new_[44319]_ , \new_[44320]_ ,
    \new_[44324]_ , \new_[44325]_ , \new_[44329]_ , \new_[44330]_ ,
    \new_[44331]_ , \new_[44335]_ , \new_[44336]_ , \new_[44339]_ ,
    \new_[44342]_ , \new_[44343]_ , \new_[44344]_ , \new_[44348]_ ,
    \new_[44349]_ , \new_[44353]_ , \new_[44354]_ , \new_[44355]_ ,
    \new_[44359]_ , \new_[44360]_ , \new_[44363]_ , \new_[44366]_ ,
    \new_[44367]_ , \new_[44368]_ , \new_[44372]_ , \new_[44373]_ ,
    \new_[44377]_ , \new_[44378]_ , \new_[44379]_ , \new_[44383]_ ,
    \new_[44384]_ , \new_[44387]_ , \new_[44390]_ , \new_[44391]_ ,
    \new_[44392]_ , \new_[44396]_ , \new_[44397]_ , \new_[44401]_ ,
    \new_[44402]_ , \new_[44403]_ , \new_[44407]_ , \new_[44408]_ ,
    \new_[44411]_ , \new_[44414]_ , \new_[44415]_ , \new_[44416]_ ,
    \new_[44420]_ , \new_[44421]_ , \new_[44425]_ , \new_[44426]_ ,
    \new_[44427]_ , \new_[44431]_ , \new_[44432]_ , \new_[44435]_ ,
    \new_[44438]_ , \new_[44439]_ , \new_[44440]_ , \new_[44444]_ ,
    \new_[44445]_ , \new_[44449]_ , \new_[44450]_ , \new_[44451]_ ,
    \new_[44455]_ , \new_[44456]_ , \new_[44459]_ , \new_[44462]_ ,
    \new_[44463]_ , \new_[44464]_ , \new_[44468]_ , \new_[44469]_ ,
    \new_[44473]_ , \new_[44474]_ , \new_[44475]_ , \new_[44479]_ ,
    \new_[44480]_ , \new_[44483]_ , \new_[44486]_ , \new_[44487]_ ,
    \new_[44488]_ , \new_[44492]_ , \new_[44493]_ , \new_[44497]_ ,
    \new_[44498]_ , \new_[44499]_ , \new_[44503]_ , \new_[44504]_ ,
    \new_[44507]_ , \new_[44510]_ , \new_[44511]_ , \new_[44512]_ ,
    \new_[44516]_ , \new_[44517]_ , \new_[44521]_ , \new_[44522]_ ,
    \new_[44523]_ , \new_[44527]_ , \new_[44528]_ , \new_[44531]_ ,
    \new_[44534]_ , \new_[44535]_ , \new_[44536]_ , \new_[44540]_ ,
    \new_[44541]_ , \new_[44545]_ , \new_[44546]_ , \new_[44547]_ ,
    \new_[44551]_ , \new_[44552]_ , \new_[44555]_ , \new_[44558]_ ,
    \new_[44559]_ , \new_[44560]_ , \new_[44564]_ , \new_[44565]_ ,
    \new_[44569]_ , \new_[44570]_ , \new_[44571]_ , \new_[44575]_ ,
    \new_[44576]_ , \new_[44579]_ , \new_[44582]_ , \new_[44583]_ ,
    \new_[44584]_ , \new_[44588]_ , \new_[44589]_ , \new_[44593]_ ,
    \new_[44594]_ , \new_[44595]_ , \new_[44599]_ , \new_[44600]_ ,
    \new_[44603]_ , \new_[44606]_ , \new_[44607]_ , \new_[44608]_ ,
    \new_[44612]_ , \new_[44613]_ , \new_[44617]_ , \new_[44618]_ ,
    \new_[44619]_ , \new_[44623]_ , \new_[44624]_ , \new_[44627]_ ,
    \new_[44630]_ , \new_[44631]_ , \new_[44632]_ , \new_[44636]_ ,
    \new_[44637]_ , \new_[44641]_ , \new_[44642]_ , \new_[44643]_ ,
    \new_[44647]_ , \new_[44648]_ , \new_[44651]_ , \new_[44654]_ ,
    \new_[44655]_ , \new_[44656]_ , \new_[44660]_ , \new_[44661]_ ,
    \new_[44665]_ , \new_[44666]_ , \new_[44667]_ , \new_[44671]_ ,
    \new_[44672]_ , \new_[44675]_ , \new_[44678]_ , \new_[44679]_ ,
    \new_[44680]_ , \new_[44684]_ , \new_[44685]_ , \new_[44689]_ ,
    \new_[44690]_ , \new_[44691]_ , \new_[44695]_ , \new_[44696]_ ,
    \new_[44699]_ , \new_[44702]_ , \new_[44703]_ , \new_[44704]_ ,
    \new_[44708]_ , \new_[44709]_ , \new_[44713]_ , \new_[44714]_ ,
    \new_[44715]_ , \new_[44719]_ , \new_[44720]_ , \new_[44723]_ ,
    \new_[44726]_ , \new_[44727]_ , \new_[44728]_ , \new_[44732]_ ,
    \new_[44733]_ , \new_[44737]_ , \new_[44738]_ , \new_[44739]_ ,
    \new_[44743]_ , \new_[44744]_ , \new_[44747]_ , \new_[44750]_ ,
    \new_[44751]_ , \new_[44752]_ , \new_[44756]_ , \new_[44757]_ ,
    \new_[44761]_ , \new_[44762]_ , \new_[44763]_ , \new_[44767]_ ,
    \new_[44768]_ , \new_[44771]_ , \new_[44774]_ , \new_[44775]_ ,
    \new_[44776]_ , \new_[44780]_ , \new_[44781]_ , \new_[44785]_ ,
    \new_[44786]_ , \new_[44787]_ , \new_[44791]_ , \new_[44792]_ ,
    \new_[44795]_ , \new_[44798]_ , \new_[44799]_ , \new_[44800]_ ,
    \new_[44804]_ , \new_[44805]_ , \new_[44809]_ , \new_[44810]_ ,
    \new_[44811]_ , \new_[44815]_ , \new_[44816]_ , \new_[44819]_ ,
    \new_[44822]_ , \new_[44823]_ , \new_[44824]_ , \new_[44828]_ ,
    \new_[44829]_ , \new_[44833]_ , \new_[44834]_ , \new_[44835]_ ,
    \new_[44839]_ , \new_[44840]_ , \new_[44843]_ , \new_[44846]_ ,
    \new_[44847]_ , \new_[44848]_ , \new_[44852]_ , \new_[44853]_ ,
    \new_[44857]_ , \new_[44858]_ , \new_[44859]_ , \new_[44863]_ ,
    \new_[44864]_ , \new_[44867]_ , \new_[44870]_ , \new_[44871]_ ,
    \new_[44872]_ , \new_[44876]_ , \new_[44877]_ , \new_[44881]_ ,
    \new_[44882]_ , \new_[44883]_ , \new_[44887]_ , \new_[44888]_ ,
    \new_[44891]_ , \new_[44894]_ , \new_[44895]_ , \new_[44896]_ ,
    \new_[44900]_ , \new_[44901]_ , \new_[44905]_ , \new_[44906]_ ,
    \new_[44907]_ , \new_[44911]_ , \new_[44912]_ , \new_[44915]_ ,
    \new_[44918]_ , \new_[44919]_ , \new_[44920]_ , \new_[44924]_ ,
    \new_[44925]_ , \new_[44929]_ , \new_[44930]_ , \new_[44931]_ ,
    \new_[44935]_ , \new_[44936]_ , \new_[44939]_ , \new_[44942]_ ,
    \new_[44943]_ , \new_[44944]_ , \new_[44948]_ , \new_[44949]_ ,
    \new_[44953]_ , \new_[44954]_ , \new_[44955]_ , \new_[44959]_ ,
    \new_[44960]_ , \new_[44963]_ , \new_[44966]_ , \new_[44967]_ ,
    \new_[44968]_ , \new_[44972]_ , \new_[44973]_ , \new_[44977]_ ,
    \new_[44978]_ , \new_[44979]_ , \new_[44983]_ , \new_[44984]_ ,
    \new_[44987]_ , \new_[44990]_ , \new_[44991]_ , \new_[44992]_ ,
    \new_[44996]_ , \new_[44997]_ , \new_[45001]_ , \new_[45002]_ ,
    \new_[45003]_ , \new_[45007]_ , \new_[45008]_ , \new_[45011]_ ,
    \new_[45014]_ , \new_[45015]_ , \new_[45016]_ , \new_[45020]_ ,
    \new_[45021]_ , \new_[45025]_ , \new_[45026]_ , \new_[45027]_ ,
    \new_[45031]_ , \new_[45032]_ , \new_[45035]_ , \new_[45038]_ ,
    \new_[45039]_ , \new_[45040]_ , \new_[45044]_ , \new_[45045]_ ,
    \new_[45049]_ , \new_[45050]_ , \new_[45051]_ , \new_[45055]_ ,
    \new_[45056]_ , \new_[45059]_ , \new_[45062]_ , \new_[45063]_ ,
    \new_[45064]_ , \new_[45068]_ , \new_[45069]_ , \new_[45073]_ ,
    \new_[45074]_ , \new_[45075]_ , \new_[45079]_ , \new_[45080]_ ,
    \new_[45083]_ , \new_[45086]_ , \new_[45087]_ , \new_[45088]_ ,
    \new_[45092]_ , \new_[45093]_ , \new_[45097]_ , \new_[45098]_ ,
    \new_[45099]_ , \new_[45103]_ , \new_[45104]_ , \new_[45107]_ ,
    \new_[45110]_ , \new_[45111]_ , \new_[45112]_ , \new_[45116]_ ,
    \new_[45117]_ , \new_[45121]_ , \new_[45122]_ , \new_[45123]_ ,
    \new_[45127]_ , \new_[45128]_ , \new_[45131]_ , \new_[45134]_ ,
    \new_[45135]_ , \new_[45136]_ , \new_[45140]_ , \new_[45141]_ ,
    \new_[45145]_ , \new_[45146]_ , \new_[45147]_ , \new_[45151]_ ,
    \new_[45152]_ , \new_[45155]_ , \new_[45158]_ , \new_[45159]_ ,
    \new_[45160]_ , \new_[45164]_ , \new_[45165]_ , \new_[45169]_ ,
    \new_[45170]_ , \new_[45171]_ , \new_[45175]_ , \new_[45176]_ ,
    \new_[45179]_ , \new_[45182]_ , \new_[45183]_ , \new_[45184]_ ,
    \new_[45188]_ , \new_[45189]_ , \new_[45193]_ , \new_[45194]_ ,
    \new_[45195]_ , \new_[45199]_ , \new_[45200]_ , \new_[45203]_ ,
    \new_[45206]_ , \new_[45207]_ , \new_[45208]_ , \new_[45212]_ ,
    \new_[45213]_ , \new_[45217]_ , \new_[45218]_ , \new_[45219]_ ,
    \new_[45223]_ , \new_[45224]_ , \new_[45227]_ , \new_[45230]_ ,
    \new_[45231]_ , \new_[45232]_ , \new_[45236]_ , \new_[45237]_ ,
    \new_[45241]_ , \new_[45242]_ , \new_[45243]_ , \new_[45247]_ ,
    \new_[45248]_ , \new_[45251]_ , \new_[45254]_ , \new_[45255]_ ,
    \new_[45256]_ , \new_[45260]_ , \new_[45261]_ , \new_[45265]_ ,
    \new_[45266]_ , \new_[45267]_ , \new_[45271]_ , \new_[45272]_ ,
    \new_[45275]_ , \new_[45278]_ , \new_[45279]_ , \new_[45280]_ ,
    \new_[45284]_ , \new_[45285]_ , \new_[45289]_ , \new_[45290]_ ,
    \new_[45291]_ , \new_[45295]_ , \new_[45296]_ , \new_[45299]_ ,
    \new_[45302]_ , \new_[45303]_ , \new_[45304]_ , \new_[45308]_ ,
    \new_[45309]_ , \new_[45313]_ , \new_[45314]_ , \new_[45315]_ ,
    \new_[45319]_ , \new_[45320]_ , \new_[45323]_ , \new_[45326]_ ,
    \new_[45327]_ , \new_[45328]_ , \new_[45332]_ , \new_[45333]_ ,
    \new_[45337]_ , \new_[45338]_ , \new_[45339]_ , \new_[45343]_ ,
    \new_[45344]_ , \new_[45347]_ , \new_[45350]_ , \new_[45351]_ ,
    \new_[45352]_ , \new_[45356]_ , \new_[45357]_ , \new_[45361]_ ,
    \new_[45362]_ , \new_[45363]_ , \new_[45367]_ , \new_[45368]_ ,
    \new_[45371]_ , \new_[45374]_ , \new_[45375]_ , \new_[45376]_ ,
    \new_[45380]_ , \new_[45381]_ , \new_[45385]_ , \new_[45386]_ ,
    \new_[45387]_ , \new_[45391]_ , \new_[45392]_ , \new_[45395]_ ,
    \new_[45398]_ , \new_[45399]_ , \new_[45400]_ , \new_[45404]_ ,
    \new_[45405]_ , \new_[45409]_ , \new_[45410]_ , \new_[45411]_ ,
    \new_[45415]_ , \new_[45416]_ , \new_[45419]_ , \new_[45422]_ ,
    \new_[45423]_ , \new_[45424]_ , \new_[45428]_ , \new_[45429]_ ,
    \new_[45433]_ , \new_[45434]_ , \new_[45435]_ , \new_[45439]_ ,
    \new_[45440]_ , \new_[45443]_ , \new_[45446]_ , \new_[45447]_ ,
    \new_[45448]_ , \new_[45452]_ , \new_[45453]_ , \new_[45457]_ ,
    \new_[45458]_ , \new_[45459]_ , \new_[45463]_ , \new_[45464]_ ,
    \new_[45467]_ , \new_[45470]_ , \new_[45471]_ , \new_[45472]_ ,
    \new_[45476]_ , \new_[45477]_ , \new_[45481]_ , \new_[45482]_ ,
    \new_[45483]_ , \new_[45487]_ , \new_[45488]_ , \new_[45491]_ ,
    \new_[45494]_ , \new_[45495]_ , \new_[45496]_ , \new_[45500]_ ,
    \new_[45501]_ , \new_[45505]_ , \new_[45506]_ , \new_[45507]_ ,
    \new_[45511]_ , \new_[45512]_ , \new_[45515]_ , \new_[45518]_ ,
    \new_[45519]_ , \new_[45520]_ , \new_[45524]_ , \new_[45525]_ ,
    \new_[45529]_ , \new_[45530]_ , \new_[45531]_ , \new_[45535]_ ,
    \new_[45536]_ , \new_[45539]_ , \new_[45542]_ , \new_[45543]_ ,
    \new_[45544]_ , \new_[45548]_ , \new_[45549]_ , \new_[45553]_ ,
    \new_[45554]_ , \new_[45555]_ , \new_[45559]_ , \new_[45560]_ ,
    \new_[45563]_ , \new_[45566]_ , \new_[45567]_ , \new_[45568]_ ,
    \new_[45572]_ , \new_[45573]_ , \new_[45577]_ , \new_[45578]_ ,
    \new_[45579]_ , \new_[45583]_ , \new_[45584]_ , \new_[45587]_ ,
    \new_[45590]_ , \new_[45591]_ , \new_[45592]_ , \new_[45596]_ ,
    \new_[45597]_ , \new_[45601]_ , \new_[45602]_ , \new_[45603]_ ,
    \new_[45607]_ , \new_[45608]_ , \new_[45611]_ , \new_[45614]_ ,
    \new_[45615]_ , \new_[45616]_ , \new_[45620]_ , \new_[45621]_ ,
    \new_[45625]_ , \new_[45626]_ , \new_[45627]_ , \new_[45631]_ ,
    \new_[45632]_ , \new_[45635]_ , \new_[45638]_ , \new_[45639]_ ,
    \new_[45640]_ , \new_[45644]_ , \new_[45645]_ , \new_[45649]_ ,
    \new_[45650]_ , \new_[45651]_ , \new_[45655]_ , \new_[45656]_ ,
    \new_[45659]_ , \new_[45662]_ , \new_[45663]_ , \new_[45664]_ ,
    \new_[45668]_ , \new_[45669]_ , \new_[45673]_ , \new_[45674]_ ,
    \new_[45675]_ , \new_[45679]_ , \new_[45680]_ , \new_[45683]_ ,
    \new_[45686]_ , \new_[45687]_ , \new_[45688]_ , \new_[45692]_ ,
    \new_[45693]_ , \new_[45697]_ , \new_[45698]_ , \new_[45699]_ ,
    \new_[45703]_ , \new_[45704]_ , \new_[45707]_ , \new_[45710]_ ,
    \new_[45711]_ , \new_[45712]_ , \new_[45716]_ , \new_[45717]_ ,
    \new_[45721]_ , \new_[45722]_ , \new_[45723]_ , \new_[45727]_ ,
    \new_[45728]_ , \new_[45731]_ , \new_[45734]_ , \new_[45735]_ ,
    \new_[45736]_ , \new_[45740]_ , \new_[45741]_ , \new_[45745]_ ,
    \new_[45746]_ , \new_[45747]_ , \new_[45751]_ , \new_[45752]_ ,
    \new_[45755]_ , \new_[45758]_ , \new_[45759]_ , \new_[45760]_ ,
    \new_[45764]_ , \new_[45765]_ , \new_[45769]_ , \new_[45770]_ ,
    \new_[45771]_ , \new_[45775]_ , \new_[45776]_ , \new_[45779]_ ,
    \new_[45782]_ , \new_[45783]_ , \new_[45784]_ , \new_[45788]_ ,
    \new_[45789]_ , \new_[45793]_ , \new_[45794]_ , \new_[45795]_ ,
    \new_[45799]_ , \new_[45800]_ , \new_[45803]_ , \new_[45806]_ ,
    \new_[45807]_ , \new_[45808]_ , \new_[45812]_ , \new_[45813]_ ,
    \new_[45817]_ , \new_[45818]_ , \new_[45819]_ , \new_[45823]_ ,
    \new_[45824]_ , \new_[45827]_ , \new_[45830]_ , \new_[45831]_ ,
    \new_[45832]_ , \new_[45836]_ , \new_[45837]_ , \new_[45841]_ ,
    \new_[45842]_ , \new_[45843]_ , \new_[45847]_ , \new_[45848]_ ,
    \new_[45851]_ , \new_[45854]_ , \new_[45855]_ , \new_[45856]_ ,
    \new_[45860]_ , \new_[45861]_ , \new_[45865]_ , \new_[45866]_ ,
    \new_[45867]_ , \new_[45871]_ , \new_[45872]_ , \new_[45875]_ ,
    \new_[45878]_ , \new_[45879]_ , \new_[45880]_ , \new_[45884]_ ,
    \new_[45885]_ , \new_[45889]_ , \new_[45890]_ , \new_[45891]_ ,
    \new_[45895]_ , \new_[45896]_ , \new_[45899]_ , \new_[45902]_ ,
    \new_[45903]_ , \new_[45904]_ , \new_[45908]_ , \new_[45909]_ ,
    \new_[45913]_ , \new_[45914]_ , \new_[45915]_ , \new_[45919]_ ,
    \new_[45920]_ , \new_[45923]_ , \new_[45926]_ , \new_[45927]_ ,
    \new_[45928]_ , \new_[45932]_ , \new_[45933]_ , \new_[45937]_ ,
    \new_[45938]_ , \new_[45939]_ , \new_[45943]_ , \new_[45944]_ ,
    \new_[45947]_ , \new_[45950]_ , \new_[45951]_ , \new_[45952]_ ,
    \new_[45956]_ , \new_[45957]_ , \new_[45961]_ , \new_[45962]_ ,
    \new_[45963]_ , \new_[45967]_ , \new_[45968]_ , \new_[45971]_ ,
    \new_[45974]_ , \new_[45975]_ , \new_[45976]_ , \new_[45980]_ ,
    \new_[45981]_ , \new_[45985]_ , \new_[45986]_ , \new_[45987]_ ,
    \new_[45991]_ , \new_[45992]_ , \new_[45995]_ , \new_[45998]_ ,
    \new_[45999]_ , \new_[46000]_ , \new_[46004]_ , \new_[46005]_ ,
    \new_[46009]_ , \new_[46010]_ , \new_[46011]_ , \new_[46015]_ ,
    \new_[46016]_ , \new_[46019]_ , \new_[46022]_ , \new_[46023]_ ,
    \new_[46024]_ , \new_[46028]_ , \new_[46029]_ , \new_[46033]_ ,
    \new_[46034]_ , \new_[46035]_ , \new_[46039]_ , \new_[46040]_ ,
    \new_[46043]_ , \new_[46046]_ , \new_[46047]_ , \new_[46048]_ ,
    \new_[46052]_ , \new_[46053]_ , \new_[46057]_ , \new_[46058]_ ,
    \new_[46059]_ , \new_[46063]_ , \new_[46064]_ , \new_[46067]_ ,
    \new_[46070]_ , \new_[46071]_ , \new_[46072]_ , \new_[46076]_ ,
    \new_[46077]_ , \new_[46081]_ , \new_[46082]_ , \new_[46083]_ ,
    \new_[46087]_ , \new_[46088]_ , \new_[46091]_ , \new_[46094]_ ,
    \new_[46095]_ , \new_[46096]_ , \new_[46100]_ , \new_[46101]_ ,
    \new_[46105]_ , \new_[46106]_ , \new_[46107]_ , \new_[46111]_ ,
    \new_[46112]_ , \new_[46115]_ , \new_[46118]_ , \new_[46119]_ ,
    \new_[46120]_ , \new_[46124]_ , \new_[46125]_ , \new_[46129]_ ,
    \new_[46130]_ , \new_[46131]_ , \new_[46135]_ , \new_[46136]_ ,
    \new_[46139]_ , \new_[46142]_ , \new_[46143]_ , \new_[46144]_ ,
    \new_[46148]_ , \new_[46149]_ , \new_[46153]_ , \new_[46154]_ ,
    \new_[46155]_ , \new_[46159]_ , \new_[46160]_ , \new_[46163]_ ,
    \new_[46166]_ , \new_[46167]_ , \new_[46168]_ , \new_[46172]_ ,
    \new_[46173]_ , \new_[46177]_ , \new_[46178]_ , \new_[46179]_ ,
    \new_[46183]_ , \new_[46184]_ , \new_[46187]_ , \new_[46190]_ ,
    \new_[46191]_ , \new_[46192]_ , \new_[46196]_ , \new_[46197]_ ,
    \new_[46201]_ , \new_[46202]_ , \new_[46203]_ , \new_[46207]_ ,
    \new_[46208]_ , \new_[46211]_ , \new_[46214]_ , \new_[46215]_ ,
    \new_[46216]_ , \new_[46220]_ , \new_[46221]_ , \new_[46225]_ ,
    \new_[46226]_ , \new_[46227]_ , \new_[46231]_ , \new_[46232]_ ,
    \new_[46235]_ , \new_[46238]_ , \new_[46239]_ , \new_[46240]_ ,
    \new_[46244]_ , \new_[46245]_ , \new_[46249]_ , \new_[46250]_ ,
    \new_[46251]_ , \new_[46255]_ , \new_[46256]_ , \new_[46259]_ ,
    \new_[46262]_ , \new_[46263]_ , \new_[46264]_ , \new_[46268]_ ,
    \new_[46269]_ , \new_[46273]_ , \new_[46274]_ , \new_[46275]_ ,
    \new_[46279]_ , \new_[46280]_ , \new_[46283]_ , \new_[46286]_ ,
    \new_[46287]_ , \new_[46288]_ , \new_[46292]_ , \new_[46293]_ ,
    \new_[46297]_ , \new_[46298]_ , \new_[46299]_ , \new_[46303]_ ,
    \new_[46304]_ , \new_[46307]_ , \new_[46310]_ , \new_[46311]_ ,
    \new_[46312]_ , \new_[46316]_ , \new_[46317]_ , \new_[46321]_ ,
    \new_[46322]_ , \new_[46323]_ , \new_[46327]_ , \new_[46328]_ ,
    \new_[46331]_ , \new_[46334]_ , \new_[46335]_ , \new_[46336]_ ,
    \new_[46340]_ , \new_[46341]_ , \new_[46345]_ , \new_[46346]_ ,
    \new_[46347]_ , \new_[46351]_ , \new_[46352]_ , \new_[46355]_ ,
    \new_[46358]_ , \new_[46359]_ , \new_[46360]_ , \new_[46364]_ ,
    \new_[46365]_ , \new_[46369]_ , \new_[46370]_ , \new_[46371]_ ,
    \new_[46375]_ , \new_[46376]_ , \new_[46379]_ , \new_[46382]_ ,
    \new_[46383]_ , \new_[46384]_ , \new_[46388]_ , \new_[46389]_ ,
    \new_[46393]_ , \new_[46394]_ , \new_[46395]_ , \new_[46399]_ ,
    \new_[46400]_ , \new_[46403]_ , \new_[46406]_ , \new_[46407]_ ,
    \new_[46408]_ , \new_[46412]_ , \new_[46413]_ , \new_[46417]_ ,
    \new_[46418]_ , \new_[46419]_ , \new_[46423]_ , \new_[46424]_ ,
    \new_[46427]_ , \new_[46430]_ , \new_[46431]_ , \new_[46432]_ ,
    \new_[46436]_ , \new_[46437]_ , \new_[46441]_ , \new_[46442]_ ,
    \new_[46443]_ , \new_[46447]_ , \new_[46448]_ , \new_[46451]_ ,
    \new_[46454]_ , \new_[46455]_ , \new_[46456]_ , \new_[46460]_ ,
    \new_[46461]_ , \new_[46465]_ , \new_[46466]_ , \new_[46467]_ ,
    \new_[46471]_ , \new_[46472]_ , \new_[46475]_ , \new_[46478]_ ,
    \new_[46479]_ , \new_[46480]_ , \new_[46484]_ , \new_[46485]_ ,
    \new_[46489]_ , \new_[46490]_ , \new_[46491]_ , \new_[46495]_ ,
    \new_[46496]_ , \new_[46499]_ , \new_[46502]_ , \new_[46503]_ ,
    \new_[46504]_ , \new_[46508]_ , \new_[46509]_ , \new_[46513]_ ,
    \new_[46514]_ , \new_[46515]_ , \new_[46519]_ , \new_[46520]_ ,
    \new_[46523]_ , \new_[46526]_ , \new_[46527]_ , \new_[46528]_ ,
    \new_[46532]_ , \new_[46533]_ , \new_[46537]_ , \new_[46538]_ ,
    \new_[46539]_ , \new_[46543]_ , \new_[46544]_ , \new_[46547]_ ,
    \new_[46550]_ , \new_[46551]_ , \new_[46552]_ , \new_[46556]_ ,
    \new_[46557]_ , \new_[46561]_ , \new_[46562]_ , \new_[46563]_ ,
    \new_[46567]_ , \new_[46568]_ , \new_[46571]_ , \new_[46574]_ ,
    \new_[46575]_ , \new_[46576]_ , \new_[46580]_ , \new_[46581]_ ,
    \new_[46585]_ , \new_[46586]_ , \new_[46587]_ , \new_[46591]_ ,
    \new_[46592]_ , \new_[46595]_ , \new_[46598]_ , \new_[46599]_ ,
    \new_[46600]_ , \new_[46604]_ , \new_[46605]_ , \new_[46609]_ ,
    \new_[46610]_ , \new_[46611]_ , \new_[46615]_ , \new_[46616]_ ,
    \new_[46619]_ , \new_[46622]_ , \new_[46623]_ , \new_[46624]_ ,
    \new_[46628]_ , \new_[46629]_ , \new_[46633]_ , \new_[46634]_ ,
    \new_[46635]_ , \new_[46639]_ , \new_[46640]_ , \new_[46643]_ ,
    \new_[46646]_ , \new_[46647]_ , \new_[46648]_ , \new_[46652]_ ,
    \new_[46653]_ , \new_[46657]_ , \new_[46658]_ , \new_[46659]_ ,
    \new_[46663]_ , \new_[46664]_ , \new_[46667]_ , \new_[46670]_ ,
    \new_[46671]_ , \new_[46672]_ , \new_[46676]_ , \new_[46677]_ ,
    \new_[46681]_ , \new_[46682]_ , \new_[46683]_ , \new_[46687]_ ,
    \new_[46688]_ , \new_[46691]_ , \new_[46694]_ , \new_[46695]_ ,
    \new_[46696]_ , \new_[46700]_ , \new_[46701]_ , \new_[46705]_ ,
    \new_[46706]_ , \new_[46707]_ , \new_[46711]_ , \new_[46712]_ ,
    \new_[46715]_ , \new_[46718]_ , \new_[46719]_ , \new_[46720]_ ,
    \new_[46724]_ , \new_[46725]_ , \new_[46729]_ , \new_[46730]_ ,
    \new_[46731]_ , \new_[46735]_ , \new_[46736]_ , \new_[46739]_ ,
    \new_[46742]_ , \new_[46743]_ , \new_[46744]_ , \new_[46748]_ ,
    \new_[46749]_ , \new_[46753]_ , \new_[46754]_ , \new_[46755]_ ,
    \new_[46759]_ , \new_[46760]_ , \new_[46763]_ , \new_[46766]_ ,
    \new_[46767]_ , \new_[46768]_ , \new_[46772]_ , \new_[46773]_ ,
    \new_[46777]_ , \new_[46778]_ , \new_[46779]_ , \new_[46783]_ ,
    \new_[46784]_ , \new_[46787]_ , \new_[46790]_ , \new_[46791]_ ,
    \new_[46792]_ , \new_[46796]_ , \new_[46797]_ , \new_[46801]_ ,
    \new_[46802]_ , \new_[46803]_ , \new_[46807]_ , \new_[46808]_ ,
    \new_[46811]_ , \new_[46814]_ , \new_[46815]_ , \new_[46816]_ ,
    \new_[46820]_ , \new_[46821]_ , \new_[46825]_ , \new_[46826]_ ,
    \new_[46827]_ , \new_[46831]_ , \new_[46832]_ , \new_[46835]_ ,
    \new_[46838]_ , \new_[46839]_ , \new_[46840]_ , \new_[46844]_ ,
    \new_[46845]_ , \new_[46849]_ , \new_[46850]_ , \new_[46851]_ ,
    \new_[46855]_ , \new_[46856]_ , \new_[46859]_ , \new_[46862]_ ,
    \new_[46863]_ , \new_[46864]_ , \new_[46868]_ , \new_[46869]_ ,
    \new_[46873]_ , \new_[46874]_ , \new_[46875]_ , \new_[46879]_ ,
    \new_[46880]_ , \new_[46883]_ , \new_[46886]_ , \new_[46887]_ ,
    \new_[46888]_ , \new_[46892]_ , \new_[46893]_ , \new_[46897]_ ,
    \new_[46898]_ , \new_[46899]_ , \new_[46903]_ , \new_[46904]_ ,
    \new_[46907]_ , \new_[46910]_ , \new_[46911]_ , \new_[46912]_ ,
    \new_[46916]_ , \new_[46917]_ , \new_[46921]_ , \new_[46922]_ ,
    \new_[46923]_ , \new_[46927]_ , \new_[46928]_ , \new_[46931]_ ,
    \new_[46934]_ , \new_[46935]_ , \new_[46936]_ , \new_[46940]_ ,
    \new_[46941]_ , \new_[46945]_ , \new_[46946]_ , \new_[46947]_ ,
    \new_[46951]_ , \new_[46952]_ , \new_[46955]_ , \new_[46958]_ ,
    \new_[46959]_ , \new_[46960]_ , \new_[46964]_ , \new_[46965]_ ,
    \new_[46969]_ , \new_[46970]_ , \new_[46971]_ , \new_[46975]_ ,
    \new_[46976]_ , \new_[46979]_ , \new_[46982]_ , \new_[46983]_ ,
    \new_[46984]_ , \new_[46988]_ , \new_[46989]_ , \new_[46993]_ ,
    \new_[46994]_ , \new_[46995]_ , \new_[46999]_ , \new_[47000]_ ,
    \new_[47003]_ , \new_[47006]_ , \new_[47007]_ , \new_[47008]_ ,
    \new_[47012]_ , \new_[47013]_ , \new_[47017]_ , \new_[47018]_ ,
    \new_[47019]_ , \new_[47023]_ , \new_[47024]_ , \new_[47027]_ ,
    \new_[47030]_ , \new_[47031]_ , \new_[47032]_ , \new_[47036]_ ,
    \new_[47037]_ , \new_[47041]_ , \new_[47042]_ , \new_[47043]_ ,
    \new_[47047]_ , \new_[47048]_ , \new_[47051]_ , \new_[47054]_ ,
    \new_[47055]_ , \new_[47056]_ , \new_[47060]_ , \new_[47061]_ ,
    \new_[47065]_ , \new_[47066]_ , \new_[47067]_ , \new_[47071]_ ,
    \new_[47072]_ , \new_[47075]_ , \new_[47078]_ , \new_[47079]_ ,
    \new_[47080]_ , \new_[47084]_ , \new_[47085]_ , \new_[47089]_ ,
    \new_[47090]_ , \new_[47091]_ , \new_[47095]_ , \new_[47096]_ ,
    \new_[47099]_ , \new_[47102]_ , \new_[47103]_ , \new_[47104]_ ,
    \new_[47108]_ , \new_[47109]_ , \new_[47113]_ , \new_[47114]_ ,
    \new_[47115]_ , \new_[47119]_ , \new_[47120]_ , \new_[47123]_ ,
    \new_[47126]_ , \new_[47127]_ , \new_[47128]_ , \new_[47132]_ ,
    \new_[47133]_ , \new_[47137]_ , \new_[47138]_ , \new_[47139]_ ,
    \new_[47143]_ , \new_[47144]_ , \new_[47147]_ , \new_[47150]_ ,
    \new_[47151]_ , \new_[47152]_ , \new_[47156]_ , \new_[47157]_ ,
    \new_[47161]_ , \new_[47162]_ , \new_[47163]_ , \new_[47167]_ ,
    \new_[47168]_ , \new_[47171]_ , \new_[47174]_ , \new_[47175]_ ,
    \new_[47176]_ , \new_[47180]_ , \new_[47181]_ , \new_[47185]_ ,
    \new_[47186]_ , \new_[47187]_ , \new_[47191]_ , \new_[47192]_ ,
    \new_[47195]_ , \new_[47198]_ , \new_[47199]_ , \new_[47200]_ ,
    \new_[47204]_ , \new_[47205]_ , \new_[47209]_ , \new_[47210]_ ,
    \new_[47211]_ , \new_[47215]_ , \new_[47216]_ , \new_[47219]_ ,
    \new_[47222]_ , \new_[47223]_ , \new_[47224]_ , \new_[47228]_ ,
    \new_[47229]_ , \new_[47233]_ , \new_[47234]_ , \new_[47235]_ ,
    \new_[47239]_ , \new_[47240]_ , \new_[47243]_ , \new_[47246]_ ,
    \new_[47247]_ , \new_[47248]_ , \new_[47252]_ , \new_[47253]_ ,
    \new_[47257]_ , \new_[47258]_ , \new_[47259]_ , \new_[47263]_ ,
    \new_[47264]_ , \new_[47267]_ , \new_[47270]_ , \new_[47271]_ ,
    \new_[47272]_ , \new_[47276]_ , \new_[47277]_ , \new_[47281]_ ,
    \new_[47282]_ , \new_[47283]_ , \new_[47287]_ , \new_[47288]_ ,
    \new_[47291]_ , \new_[47294]_ , \new_[47295]_ , \new_[47296]_ ,
    \new_[47300]_ , \new_[47301]_ , \new_[47305]_ , \new_[47306]_ ,
    \new_[47307]_ , \new_[47311]_ , \new_[47312]_ , \new_[47315]_ ,
    \new_[47318]_ , \new_[47319]_ , \new_[47320]_ , \new_[47324]_ ,
    \new_[47325]_ , \new_[47329]_ , \new_[47330]_ , \new_[47331]_ ,
    \new_[47335]_ , \new_[47336]_ , \new_[47339]_ , \new_[47342]_ ,
    \new_[47343]_ , \new_[47344]_ , \new_[47348]_ , \new_[47349]_ ,
    \new_[47353]_ , \new_[47354]_ , \new_[47355]_ , \new_[47359]_ ,
    \new_[47360]_ , \new_[47363]_ , \new_[47366]_ , \new_[47367]_ ,
    \new_[47368]_ , \new_[47372]_ , \new_[47373]_ , \new_[47377]_ ,
    \new_[47378]_ , \new_[47379]_ , \new_[47383]_ , \new_[47384]_ ,
    \new_[47387]_ , \new_[47390]_ , \new_[47391]_ , \new_[47392]_ ,
    \new_[47396]_ , \new_[47397]_ , \new_[47401]_ , \new_[47402]_ ,
    \new_[47403]_ , \new_[47407]_ , \new_[47408]_ , \new_[47411]_ ,
    \new_[47414]_ , \new_[47415]_ , \new_[47416]_ , \new_[47420]_ ,
    \new_[47421]_ , \new_[47425]_ , \new_[47426]_ , \new_[47427]_ ,
    \new_[47431]_ , \new_[47432]_ , \new_[47435]_ , \new_[47438]_ ,
    \new_[47439]_ , \new_[47440]_ , \new_[47444]_ , \new_[47445]_ ,
    \new_[47449]_ , \new_[47450]_ , \new_[47451]_ , \new_[47455]_ ,
    \new_[47456]_ , \new_[47459]_ , \new_[47462]_ , \new_[47463]_ ,
    \new_[47464]_ , \new_[47468]_ , \new_[47469]_ , \new_[47473]_ ,
    \new_[47474]_ , \new_[47475]_ , \new_[47479]_ , \new_[47480]_ ,
    \new_[47483]_ , \new_[47486]_ , \new_[47487]_ , \new_[47488]_ ,
    \new_[47492]_ , \new_[47493]_ , \new_[47497]_ , \new_[47498]_ ,
    \new_[47499]_ , \new_[47503]_ , \new_[47504]_ , \new_[47507]_ ,
    \new_[47510]_ , \new_[47511]_ , \new_[47512]_ , \new_[47516]_ ,
    \new_[47517]_ , \new_[47521]_ , \new_[47522]_ , \new_[47523]_ ,
    \new_[47527]_ , \new_[47528]_ , \new_[47531]_ , \new_[47534]_ ,
    \new_[47535]_ , \new_[47536]_ , \new_[47540]_ , \new_[47541]_ ,
    \new_[47545]_ , \new_[47546]_ , \new_[47547]_ , \new_[47551]_ ,
    \new_[47552]_ , \new_[47555]_ , \new_[47558]_ , \new_[47559]_ ,
    \new_[47560]_ , \new_[47564]_ , \new_[47565]_ , \new_[47569]_ ,
    \new_[47570]_ , \new_[47571]_ , \new_[47575]_ , \new_[47576]_ ,
    \new_[47579]_ , \new_[47582]_ , \new_[47583]_ , \new_[47584]_ ,
    \new_[47588]_ , \new_[47589]_ , \new_[47593]_ , \new_[47594]_ ,
    \new_[47595]_ , \new_[47599]_ , \new_[47600]_ , \new_[47603]_ ,
    \new_[47606]_ , \new_[47607]_ , \new_[47608]_ , \new_[47612]_ ,
    \new_[47613]_ , \new_[47617]_ , \new_[47618]_ , \new_[47619]_ ,
    \new_[47623]_ , \new_[47624]_ , \new_[47627]_ , \new_[47630]_ ,
    \new_[47631]_ , \new_[47632]_ , \new_[47636]_ , \new_[47637]_ ,
    \new_[47641]_ , \new_[47642]_ , \new_[47643]_ , \new_[47647]_ ,
    \new_[47648]_ , \new_[47651]_ , \new_[47654]_ , \new_[47655]_ ,
    \new_[47656]_ , \new_[47660]_ , \new_[47661]_ , \new_[47665]_ ,
    \new_[47666]_ , \new_[47667]_ , \new_[47671]_ , \new_[47672]_ ,
    \new_[47675]_ , \new_[47678]_ , \new_[47679]_ , \new_[47680]_ ,
    \new_[47684]_ , \new_[47685]_ , \new_[47689]_ , \new_[47690]_ ,
    \new_[47691]_ , \new_[47695]_ , \new_[47696]_ , \new_[47699]_ ,
    \new_[47702]_ , \new_[47703]_ , \new_[47704]_ , \new_[47708]_ ,
    \new_[47709]_ , \new_[47713]_ , \new_[47714]_ , \new_[47715]_ ,
    \new_[47719]_ , \new_[47720]_ , \new_[47723]_ , \new_[47726]_ ,
    \new_[47727]_ , \new_[47728]_ , \new_[47732]_ , \new_[47733]_ ,
    \new_[47737]_ , \new_[47738]_ , \new_[47739]_ , \new_[47743]_ ,
    \new_[47744]_ , \new_[47747]_ , \new_[47750]_ , \new_[47751]_ ,
    \new_[47752]_ , \new_[47756]_ , \new_[47757]_ , \new_[47761]_ ,
    \new_[47762]_ , \new_[47763]_ , \new_[47767]_ , \new_[47768]_ ,
    \new_[47771]_ , \new_[47774]_ , \new_[47775]_ , \new_[47776]_ ,
    \new_[47780]_ , \new_[47781]_ , \new_[47785]_ , \new_[47786]_ ,
    \new_[47787]_ , \new_[47791]_ , \new_[47792]_ , \new_[47795]_ ,
    \new_[47798]_ , \new_[47799]_ , \new_[47800]_ , \new_[47804]_ ,
    \new_[47805]_ , \new_[47809]_ , \new_[47810]_ , \new_[47811]_ ,
    \new_[47815]_ , \new_[47816]_ , \new_[47819]_ , \new_[47822]_ ,
    \new_[47823]_ , \new_[47824]_ , \new_[47828]_ , \new_[47829]_ ,
    \new_[47833]_ , \new_[47834]_ , \new_[47835]_ , \new_[47839]_ ,
    \new_[47840]_ , \new_[47843]_ , \new_[47846]_ , \new_[47847]_ ,
    \new_[47848]_ , \new_[47852]_ , \new_[47853]_ , \new_[47857]_ ,
    \new_[47858]_ , \new_[47859]_ , \new_[47863]_ , \new_[47864]_ ,
    \new_[47867]_ , \new_[47870]_ , \new_[47871]_ , \new_[47872]_ ,
    \new_[47876]_ , \new_[47877]_ , \new_[47881]_ , \new_[47882]_ ,
    \new_[47883]_ , \new_[47887]_ , \new_[47888]_ , \new_[47891]_ ,
    \new_[47894]_ , \new_[47895]_ , \new_[47896]_ , \new_[47900]_ ,
    \new_[47901]_ , \new_[47905]_ , \new_[47906]_ , \new_[47907]_ ,
    \new_[47911]_ , \new_[47912]_ , \new_[47915]_ , \new_[47918]_ ,
    \new_[47919]_ , \new_[47920]_ , \new_[47924]_ , \new_[47925]_ ,
    \new_[47929]_ , \new_[47930]_ , \new_[47931]_ , \new_[47935]_ ,
    \new_[47936]_ , \new_[47939]_ , \new_[47942]_ , \new_[47943]_ ,
    \new_[47944]_ , \new_[47948]_ , \new_[47949]_ , \new_[47953]_ ,
    \new_[47954]_ , \new_[47955]_ , \new_[47959]_ , \new_[47960]_ ,
    \new_[47963]_ , \new_[47966]_ , \new_[47967]_ , \new_[47968]_ ,
    \new_[47972]_ , \new_[47973]_ , \new_[47977]_ , \new_[47978]_ ,
    \new_[47979]_ , \new_[47983]_ , \new_[47984]_ , \new_[47987]_ ,
    \new_[47990]_ , \new_[47991]_ , \new_[47992]_ , \new_[47996]_ ,
    \new_[47997]_ , \new_[48001]_ , \new_[48002]_ , \new_[48003]_ ,
    \new_[48007]_ , \new_[48008]_ , \new_[48011]_ , \new_[48014]_ ,
    \new_[48015]_ , \new_[48016]_ , \new_[48020]_ , \new_[48021]_ ,
    \new_[48025]_ , \new_[48026]_ , \new_[48027]_ , \new_[48031]_ ,
    \new_[48032]_ , \new_[48035]_ , \new_[48038]_ , \new_[48039]_ ,
    \new_[48040]_ , \new_[48044]_ , \new_[48045]_ , \new_[48049]_ ,
    \new_[48050]_ , \new_[48051]_ , \new_[48055]_ , \new_[48056]_ ,
    \new_[48059]_ , \new_[48062]_ , \new_[48063]_ , \new_[48064]_ ,
    \new_[48068]_ , \new_[48069]_ , \new_[48073]_ , \new_[48074]_ ,
    \new_[48075]_ , \new_[48079]_ , \new_[48080]_ , \new_[48083]_ ,
    \new_[48086]_ , \new_[48087]_ , \new_[48088]_ , \new_[48092]_ ,
    \new_[48093]_ , \new_[48097]_ , \new_[48098]_ , \new_[48099]_ ,
    \new_[48103]_ , \new_[48104]_ , \new_[48107]_ , \new_[48110]_ ,
    \new_[48111]_ , \new_[48112]_ , \new_[48116]_ , \new_[48117]_ ,
    \new_[48121]_ , \new_[48122]_ , \new_[48123]_ , \new_[48127]_ ,
    \new_[48128]_ , \new_[48131]_ , \new_[48134]_ , \new_[48135]_ ,
    \new_[48136]_ , \new_[48140]_ , \new_[48141]_ , \new_[48145]_ ,
    \new_[48146]_ , \new_[48147]_ , \new_[48151]_ , \new_[48152]_ ,
    \new_[48155]_ , \new_[48158]_ , \new_[48159]_ , \new_[48160]_ ,
    \new_[48164]_ , \new_[48165]_ , \new_[48169]_ , \new_[48170]_ ,
    \new_[48171]_ , \new_[48175]_ , \new_[48176]_ , \new_[48179]_ ,
    \new_[48182]_ , \new_[48183]_ , \new_[48184]_ , \new_[48188]_ ,
    \new_[48189]_ , \new_[48193]_ , \new_[48194]_ , \new_[48195]_ ,
    \new_[48199]_ , \new_[48200]_ , \new_[48203]_ , \new_[48206]_ ,
    \new_[48207]_ , \new_[48208]_ , \new_[48212]_ , \new_[48213]_ ,
    \new_[48217]_ , \new_[48218]_ , \new_[48219]_ , \new_[48223]_ ,
    \new_[48224]_ , \new_[48227]_ , \new_[48230]_ , \new_[48231]_ ,
    \new_[48232]_ , \new_[48236]_ , \new_[48237]_ , \new_[48241]_ ,
    \new_[48242]_ , \new_[48243]_ , \new_[48247]_ , \new_[48248]_ ,
    \new_[48251]_ , \new_[48254]_ , \new_[48255]_ , \new_[48256]_ ,
    \new_[48260]_ , \new_[48261]_ , \new_[48265]_ , \new_[48266]_ ,
    \new_[48267]_ , \new_[48271]_ , \new_[48272]_ , \new_[48275]_ ,
    \new_[48278]_ , \new_[48279]_ , \new_[48280]_ , \new_[48284]_ ,
    \new_[48285]_ , \new_[48289]_ , \new_[48290]_ , \new_[48291]_ ,
    \new_[48295]_ , \new_[48296]_ , \new_[48299]_ , \new_[48302]_ ,
    \new_[48303]_ , \new_[48304]_ , \new_[48308]_ , \new_[48309]_ ,
    \new_[48313]_ , \new_[48314]_ , \new_[48315]_ , \new_[48319]_ ,
    \new_[48320]_ , \new_[48323]_ , \new_[48326]_ , \new_[48327]_ ,
    \new_[48328]_ , \new_[48332]_ , \new_[48333]_ , \new_[48337]_ ,
    \new_[48338]_ , \new_[48339]_ , \new_[48343]_ , \new_[48344]_ ,
    \new_[48347]_ , \new_[48350]_ , \new_[48351]_ , \new_[48352]_ ,
    \new_[48356]_ , \new_[48357]_ , \new_[48361]_ , \new_[48362]_ ,
    \new_[48363]_ , \new_[48367]_ , \new_[48368]_ , \new_[48371]_ ,
    \new_[48374]_ , \new_[48375]_ , \new_[48376]_ , \new_[48380]_ ,
    \new_[48381]_ , \new_[48385]_ , \new_[48386]_ , \new_[48387]_ ,
    \new_[48391]_ , \new_[48392]_ , \new_[48395]_ , \new_[48398]_ ,
    \new_[48399]_ , \new_[48400]_ , \new_[48404]_ , \new_[48405]_ ,
    \new_[48409]_ , \new_[48410]_ , \new_[48411]_ , \new_[48415]_ ,
    \new_[48416]_ , \new_[48419]_ , \new_[48422]_ , \new_[48423]_ ,
    \new_[48424]_ , \new_[48428]_ , \new_[48429]_ , \new_[48433]_ ,
    \new_[48434]_ , \new_[48435]_ , \new_[48439]_ , \new_[48440]_ ,
    \new_[48443]_ , \new_[48446]_ , \new_[48447]_ , \new_[48448]_ ,
    \new_[48452]_ , \new_[48453]_ , \new_[48457]_ , \new_[48458]_ ,
    \new_[48459]_ , \new_[48463]_ , \new_[48464]_ , \new_[48467]_ ,
    \new_[48470]_ , \new_[48471]_ , \new_[48472]_ , \new_[48476]_ ,
    \new_[48477]_ , \new_[48481]_ , \new_[48482]_ , \new_[48483]_ ,
    \new_[48487]_ , \new_[48488]_ , \new_[48491]_ , \new_[48494]_ ,
    \new_[48495]_ , \new_[48496]_ , \new_[48500]_ , \new_[48501]_ ,
    \new_[48505]_ , \new_[48506]_ , \new_[48507]_ , \new_[48511]_ ,
    \new_[48512]_ , \new_[48515]_ , \new_[48518]_ , \new_[48519]_ ,
    \new_[48520]_ , \new_[48524]_ , \new_[48525]_ , \new_[48529]_ ,
    \new_[48530]_ , \new_[48531]_ , \new_[48535]_ , \new_[48536]_ ,
    \new_[48539]_ , \new_[48542]_ , \new_[48543]_ , \new_[48544]_ ,
    \new_[48548]_ , \new_[48549]_ , \new_[48553]_ , \new_[48554]_ ,
    \new_[48555]_ , \new_[48559]_ , \new_[48560]_ , \new_[48563]_ ,
    \new_[48566]_ , \new_[48567]_ , \new_[48568]_ , \new_[48572]_ ,
    \new_[48573]_ , \new_[48577]_ , \new_[48578]_ , \new_[48579]_ ,
    \new_[48583]_ , \new_[48584]_ , \new_[48587]_ , \new_[48590]_ ,
    \new_[48591]_ , \new_[48592]_ , \new_[48596]_ , \new_[48597]_ ,
    \new_[48601]_ , \new_[48602]_ , \new_[48603]_ , \new_[48607]_ ,
    \new_[48608]_ , \new_[48611]_ , \new_[48614]_ , \new_[48615]_ ,
    \new_[48616]_ , \new_[48620]_ , \new_[48621]_ , \new_[48625]_ ,
    \new_[48626]_ , \new_[48627]_ , \new_[48631]_ , \new_[48632]_ ,
    \new_[48635]_ , \new_[48638]_ , \new_[48639]_ , \new_[48640]_ ,
    \new_[48644]_ , \new_[48645]_ , \new_[48649]_ , \new_[48650]_ ,
    \new_[48651]_ , \new_[48655]_ , \new_[48656]_ , \new_[48659]_ ,
    \new_[48662]_ , \new_[48663]_ , \new_[48664]_ , \new_[48668]_ ,
    \new_[48669]_ , \new_[48673]_ , \new_[48674]_ , \new_[48675]_ ,
    \new_[48679]_ , \new_[48680]_ , \new_[48683]_ , \new_[48686]_ ,
    \new_[48687]_ , \new_[48688]_ , \new_[48692]_ , \new_[48693]_ ,
    \new_[48697]_ , \new_[48698]_ , \new_[48699]_ , \new_[48703]_ ,
    \new_[48704]_ , \new_[48707]_ , \new_[48710]_ , \new_[48711]_ ,
    \new_[48712]_ , \new_[48716]_ , \new_[48717]_ , \new_[48721]_ ,
    \new_[48722]_ , \new_[48723]_ , \new_[48727]_ , \new_[48728]_ ,
    \new_[48731]_ , \new_[48734]_ , \new_[48735]_ , \new_[48736]_ ,
    \new_[48740]_ , \new_[48741]_ , \new_[48745]_ , \new_[48746]_ ,
    \new_[48747]_ , \new_[48751]_ , \new_[48752]_ , \new_[48755]_ ,
    \new_[48758]_ , \new_[48759]_ , \new_[48760]_ , \new_[48764]_ ,
    \new_[48765]_ , \new_[48769]_ , \new_[48770]_ , \new_[48771]_ ,
    \new_[48775]_ , \new_[48776]_ , \new_[48779]_ , \new_[48782]_ ,
    \new_[48783]_ , \new_[48784]_ , \new_[48788]_ , \new_[48789]_ ,
    \new_[48793]_ , \new_[48794]_ , \new_[48795]_ , \new_[48799]_ ,
    \new_[48800]_ , \new_[48803]_ , \new_[48806]_ , \new_[48807]_ ,
    \new_[48808]_ , \new_[48812]_ , \new_[48813]_ , \new_[48817]_ ,
    \new_[48818]_ , \new_[48819]_ , \new_[48823]_ , \new_[48824]_ ,
    \new_[48827]_ , \new_[48830]_ , \new_[48831]_ , \new_[48832]_ ,
    \new_[48836]_ , \new_[48837]_ , \new_[48841]_ , \new_[48842]_ ,
    \new_[48843]_ , \new_[48847]_ , \new_[48848]_ , \new_[48851]_ ,
    \new_[48854]_ , \new_[48855]_ , \new_[48856]_ , \new_[48860]_ ,
    \new_[48861]_ , \new_[48865]_ , \new_[48866]_ , \new_[48867]_ ,
    \new_[48871]_ , \new_[48872]_ , \new_[48875]_ , \new_[48878]_ ,
    \new_[48879]_ , \new_[48880]_ , \new_[48884]_ , \new_[48885]_ ,
    \new_[48889]_ , \new_[48890]_ , \new_[48891]_ , \new_[48895]_ ,
    \new_[48896]_ , \new_[48899]_ , \new_[48902]_ , \new_[48903]_ ,
    \new_[48904]_ , \new_[48908]_ , \new_[48909]_ , \new_[48913]_ ,
    \new_[48914]_ , \new_[48915]_ , \new_[48919]_ , \new_[48920]_ ,
    \new_[48923]_ , \new_[48926]_ , \new_[48927]_ , \new_[48928]_ ,
    \new_[48932]_ , \new_[48933]_ , \new_[48937]_ , \new_[48938]_ ,
    \new_[48939]_ , \new_[48943]_ , \new_[48944]_ , \new_[48947]_ ,
    \new_[48950]_ , \new_[48951]_ , \new_[48952]_ , \new_[48956]_ ,
    \new_[48957]_ , \new_[48961]_ , \new_[48962]_ , \new_[48963]_ ,
    \new_[48967]_ , \new_[48968]_ , \new_[48971]_ , \new_[48974]_ ,
    \new_[48975]_ , \new_[48976]_ , \new_[48980]_ , \new_[48981]_ ,
    \new_[48985]_ , \new_[48986]_ , \new_[48987]_ , \new_[48991]_ ,
    \new_[48992]_ , \new_[48995]_ , \new_[48998]_ , \new_[48999]_ ,
    \new_[49000]_ , \new_[49004]_ , \new_[49005]_ , \new_[49009]_ ,
    \new_[49010]_ , \new_[49011]_ , \new_[49015]_ , \new_[49016]_ ,
    \new_[49019]_ , \new_[49022]_ , \new_[49023]_ , \new_[49024]_ ,
    \new_[49028]_ , \new_[49029]_ , \new_[49033]_ , \new_[49034]_ ,
    \new_[49035]_ , \new_[49039]_ , \new_[49040]_ , \new_[49043]_ ,
    \new_[49046]_ , \new_[49047]_ , \new_[49048]_ , \new_[49052]_ ,
    \new_[49053]_ , \new_[49057]_ , \new_[49058]_ , \new_[49059]_ ,
    \new_[49063]_ , \new_[49064]_ , \new_[49067]_ , \new_[49070]_ ,
    \new_[49071]_ , \new_[49072]_ , \new_[49076]_ , \new_[49077]_ ,
    \new_[49081]_ , \new_[49082]_ , \new_[49083]_ , \new_[49087]_ ,
    \new_[49088]_ , \new_[49091]_ , \new_[49094]_ , \new_[49095]_ ,
    \new_[49096]_ , \new_[49100]_ , \new_[49101]_ , \new_[49105]_ ,
    \new_[49106]_ , \new_[49107]_ , \new_[49111]_ , \new_[49112]_ ,
    \new_[49115]_ , \new_[49118]_ , \new_[49119]_ , \new_[49120]_ ,
    \new_[49124]_ , \new_[49125]_ , \new_[49129]_ , \new_[49130]_ ,
    \new_[49131]_ , \new_[49135]_ , \new_[49136]_ , \new_[49139]_ ,
    \new_[49142]_ , \new_[49143]_ , \new_[49144]_ , \new_[49148]_ ,
    \new_[49149]_ , \new_[49153]_ , \new_[49154]_ , \new_[49155]_ ,
    \new_[49159]_ , \new_[49160]_ , \new_[49163]_ , \new_[49166]_ ,
    \new_[49167]_ , \new_[49168]_ , \new_[49172]_ , \new_[49173]_ ,
    \new_[49177]_ , \new_[49178]_ , \new_[49179]_ , \new_[49183]_ ,
    \new_[49184]_ , \new_[49187]_ , \new_[49190]_ , \new_[49191]_ ,
    \new_[49192]_ , \new_[49196]_ , \new_[49197]_ , \new_[49201]_ ,
    \new_[49202]_ , \new_[49203]_ , \new_[49207]_ , \new_[49208]_ ,
    \new_[49211]_ , \new_[49214]_ , \new_[49215]_ , \new_[49216]_ ,
    \new_[49220]_ , \new_[49221]_ , \new_[49225]_ , \new_[49226]_ ,
    \new_[49227]_ , \new_[49231]_ , \new_[49232]_ , \new_[49235]_ ,
    \new_[49238]_ , \new_[49239]_ , \new_[49240]_ , \new_[49244]_ ,
    \new_[49245]_ , \new_[49249]_ , \new_[49250]_ , \new_[49251]_ ,
    \new_[49255]_ , \new_[49256]_ , \new_[49259]_ , \new_[49262]_ ,
    \new_[49263]_ , \new_[49264]_ , \new_[49268]_ , \new_[49269]_ ,
    \new_[49273]_ , \new_[49274]_ , \new_[49275]_ , \new_[49279]_ ,
    \new_[49280]_ , \new_[49283]_ , \new_[49286]_ , \new_[49287]_ ,
    \new_[49288]_ , \new_[49292]_ , \new_[49293]_ , \new_[49297]_ ,
    \new_[49298]_ , \new_[49299]_ , \new_[49303]_ , \new_[49304]_ ,
    \new_[49307]_ , \new_[49310]_ , \new_[49311]_ , \new_[49312]_ ,
    \new_[49316]_ , \new_[49317]_ , \new_[49321]_ , \new_[49322]_ ,
    \new_[49323]_ , \new_[49327]_ , \new_[49328]_ , \new_[49331]_ ,
    \new_[49334]_ , \new_[49335]_ , \new_[49336]_ , \new_[49340]_ ,
    \new_[49341]_ , \new_[49345]_ , \new_[49346]_ , \new_[49347]_ ,
    \new_[49351]_ , \new_[49352]_ , \new_[49355]_ , \new_[49358]_ ,
    \new_[49359]_ , \new_[49360]_ , \new_[49364]_ , \new_[49365]_ ,
    \new_[49369]_ , \new_[49370]_ , \new_[49371]_ , \new_[49375]_ ,
    \new_[49376]_ , \new_[49379]_ , \new_[49382]_ , \new_[49383]_ ,
    \new_[49384]_ , \new_[49388]_ , \new_[49389]_ , \new_[49393]_ ,
    \new_[49394]_ , \new_[49395]_ , \new_[49399]_ , \new_[49400]_ ,
    \new_[49403]_ , \new_[49406]_ , \new_[49407]_ , \new_[49408]_ ,
    \new_[49412]_ , \new_[49413]_ , \new_[49417]_ , \new_[49418]_ ,
    \new_[49419]_ , \new_[49423]_ , \new_[49424]_ , \new_[49427]_ ,
    \new_[49430]_ , \new_[49431]_ , \new_[49432]_ , \new_[49436]_ ,
    \new_[49437]_ , \new_[49441]_ , \new_[49442]_ , \new_[49443]_ ,
    \new_[49447]_ , \new_[49448]_ , \new_[49451]_ , \new_[49454]_ ,
    \new_[49455]_ , \new_[49456]_ , \new_[49460]_ , \new_[49461]_ ,
    \new_[49465]_ , \new_[49466]_ , \new_[49467]_ , \new_[49471]_ ,
    \new_[49472]_ , \new_[49475]_ , \new_[49478]_ , \new_[49479]_ ,
    \new_[49480]_ , \new_[49484]_ , \new_[49485]_ , \new_[49489]_ ,
    \new_[49490]_ , \new_[49491]_ , \new_[49495]_ , \new_[49496]_ ,
    \new_[49499]_ , \new_[49502]_ , \new_[49503]_ , \new_[49504]_ ,
    \new_[49508]_ , \new_[49509]_ , \new_[49513]_ , \new_[49514]_ ,
    \new_[49515]_ , \new_[49519]_ , \new_[49520]_ , \new_[49523]_ ,
    \new_[49526]_ , \new_[49527]_ , \new_[49528]_ , \new_[49532]_ ,
    \new_[49533]_ , \new_[49537]_ , \new_[49538]_ , \new_[49539]_ ,
    \new_[49543]_ , \new_[49544]_ , \new_[49547]_ , \new_[49550]_ ,
    \new_[49551]_ , \new_[49552]_ , \new_[49556]_ , \new_[49557]_ ,
    \new_[49561]_ , \new_[49562]_ , \new_[49563]_ , \new_[49567]_ ,
    \new_[49568]_ , \new_[49571]_ , \new_[49574]_ , \new_[49575]_ ,
    \new_[49576]_ , \new_[49580]_ , \new_[49581]_ , \new_[49585]_ ,
    \new_[49586]_ , \new_[49587]_ , \new_[49591]_ , \new_[49592]_ ,
    \new_[49595]_ , \new_[49598]_ , \new_[49599]_ , \new_[49600]_ ,
    \new_[49604]_ , \new_[49605]_ , \new_[49609]_ , \new_[49610]_ ,
    \new_[49611]_ , \new_[49615]_ , \new_[49616]_ , \new_[49619]_ ,
    \new_[49622]_ , \new_[49623]_ , \new_[49624]_ , \new_[49628]_ ,
    \new_[49629]_ , \new_[49633]_ , \new_[49634]_ , \new_[49635]_ ,
    \new_[49639]_ , \new_[49640]_ , \new_[49643]_ , \new_[49646]_ ,
    \new_[49647]_ , \new_[49648]_ , \new_[49652]_ , \new_[49653]_ ,
    \new_[49657]_ , \new_[49658]_ , \new_[49659]_ , \new_[49663]_ ,
    \new_[49664]_ , \new_[49667]_ , \new_[49670]_ , \new_[49671]_ ,
    \new_[49672]_ , \new_[49676]_ , \new_[49677]_ , \new_[49681]_ ,
    \new_[49682]_ , \new_[49683]_ , \new_[49687]_ , \new_[49688]_ ,
    \new_[49691]_ , \new_[49694]_ , \new_[49695]_ , \new_[49696]_ ,
    \new_[49700]_ , \new_[49701]_ , \new_[49705]_ , \new_[49706]_ ,
    \new_[49707]_ , \new_[49711]_ , \new_[49712]_ , \new_[49715]_ ,
    \new_[49718]_ , \new_[49719]_ , \new_[49720]_ , \new_[49724]_ ,
    \new_[49725]_ , \new_[49729]_ , \new_[49730]_ , \new_[49731]_ ,
    \new_[49735]_ , \new_[49736]_ , \new_[49739]_ , \new_[49742]_ ,
    \new_[49743]_ , \new_[49744]_ , \new_[49748]_ , \new_[49749]_ ,
    \new_[49753]_ , \new_[49754]_ , \new_[49755]_ , \new_[49759]_ ,
    \new_[49760]_ , \new_[49763]_ , \new_[49766]_ , \new_[49767]_ ,
    \new_[49768]_ , \new_[49772]_ , \new_[49773]_ , \new_[49777]_ ,
    \new_[49778]_ , \new_[49779]_ , \new_[49783]_ , \new_[49784]_ ,
    \new_[49787]_ , \new_[49790]_ , \new_[49791]_ , \new_[49792]_ ,
    \new_[49796]_ , \new_[49797]_ , \new_[49801]_ , \new_[49802]_ ,
    \new_[49803]_ , \new_[49807]_ , \new_[49808]_ , \new_[49811]_ ,
    \new_[49814]_ , \new_[49815]_ , \new_[49816]_ , \new_[49820]_ ,
    \new_[49821]_ , \new_[49825]_ , \new_[49826]_ , \new_[49827]_ ,
    \new_[49831]_ , \new_[49832]_ , \new_[49835]_ , \new_[49838]_ ,
    \new_[49839]_ , \new_[49840]_ , \new_[49844]_ , \new_[49845]_ ,
    \new_[49849]_ , \new_[49850]_ , \new_[49851]_ , \new_[49855]_ ,
    \new_[49856]_ , \new_[49859]_ , \new_[49862]_ , \new_[49863]_ ,
    \new_[49864]_ , \new_[49868]_ , \new_[49869]_ , \new_[49873]_ ,
    \new_[49874]_ , \new_[49875]_ , \new_[49879]_ , \new_[49880]_ ,
    \new_[49883]_ , \new_[49886]_ , \new_[49887]_ , \new_[49888]_ ,
    \new_[49892]_ , \new_[49893]_ , \new_[49897]_ , \new_[49898]_ ,
    \new_[49899]_ , \new_[49903]_ , \new_[49904]_ , \new_[49907]_ ,
    \new_[49910]_ , \new_[49911]_ , \new_[49912]_ , \new_[49916]_ ,
    \new_[49917]_ , \new_[49921]_ , \new_[49922]_ , \new_[49923]_ ,
    \new_[49927]_ , \new_[49928]_ , \new_[49931]_ , \new_[49934]_ ,
    \new_[49935]_ , \new_[49936]_ , \new_[49940]_ , \new_[49941]_ ,
    \new_[49945]_ , \new_[49946]_ , \new_[49947]_ , \new_[49951]_ ,
    \new_[49952]_ , \new_[49955]_ , \new_[49958]_ , \new_[49959]_ ,
    \new_[49960]_ , \new_[49964]_ , \new_[49965]_ , \new_[49969]_ ,
    \new_[49970]_ , \new_[49971]_ , \new_[49975]_ , \new_[49976]_ ,
    \new_[49979]_ , \new_[49982]_ , \new_[49983]_ , \new_[49984]_ ,
    \new_[49988]_ , \new_[49989]_ , \new_[49993]_ , \new_[49994]_ ,
    \new_[49995]_ , \new_[49999]_ , \new_[50000]_ , \new_[50003]_ ,
    \new_[50006]_ , \new_[50007]_ , \new_[50008]_ , \new_[50012]_ ,
    \new_[50013]_ , \new_[50017]_ , \new_[50018]_ , \new_[50019]_ ,
    \new_[50023]_ , \new_[50024]_ , \new_[50027]_ , \new_[50030]_ ,
    \new_[50031]_ , \new_[50032]_ , \new_[50036]_ , \new_[50037]_ ,
    \new_[50041]_ , \new_[50042]_ , \new_[50043]_ , \new_[50047]_ ,
    \new_[50048]_ , \new_[50051]_ , \new_[50054]_ , \new_[50055]_ ,
    \new_[50056]_ , \new_[50060]_ , \new_[50061]_ , \new_[50065]_ ,
    \new_[50066]_ , \new_[50067]_ , \new_[50071]_ , \new_[50072]_ ,
    \new_[50075]_ , \new_[50078]_ , \new_[50079]_ , \new_[50080]_ ,
    \new_[50084]_ , \new_[50085]_ , \new_[50089]_ , \new_[50090]_ ,
    \new_[50091]_ , \new_[50095]_ , \new_[50096]_ , \new_[50099]_ ,
    \new_[50102]_ , \new_[50103]_ , \new_[50104]_ , \new_[50108]_ ,
    \new_[50109]_ , \new_[50113]_ , \new_[50114]_ , \new_[50115]_ ,
    \new_[50119]_ , \new_[50120]_ , \new_[50123]_ , \new_[50126]_ ,
    \new_[50127]_ , \new_[50128]_ , \new_[50132]_ , \new_[50133]_ ,
    \new_[50137]_ , \new_[50138]_ , \new_[50139]_ , \new_[50143]_ ,
    \new_[50144]_ , \new_[50147]_ , \new_[50150]_ , \new_[50151]_ ,
    \new_[50152]_ , \new_[50156]_ , \new_[50157]_ , \new_[50161]_ ,
    \new_[50162]_ , \new_[50163]_ , \new_[50167]_ , \new_[50168]_ ,
    \new_[50171]_ , \new_[50174]_ , \new_[50175]_ , \new_[50176]_ ,
    \new_[50180]_ , \new_[50181]_ , \new_[50185]_ , \new_[50186]_ ,
    \new_[50187]_ , \new_[50191]_ , \new_[50192]_ , \new_[50195]_ ,
    \new_[50198]_ , \new_[50199]_ , \new_[50200]_ , \new_[50204]_ ,
    \new_[50205]_ , \new_[50209]_ , \new_[50210]_ , \new_[50211]_ ,
    \new_[50215]_ , \new_[50216]_ , \new_[50219]_ , \new_[50222]_ ,
    \new_[50223]_ , \new_[50224]_ , \new_[50228]_ , \new_[50229]_ ,
    \new_[50233]_ , \new_[50234]_ , \new_[50235]_ , \new_[50239]_ ,
    \new_[50240]_ , \new_[50243]_ , \new_[50246]_ , \new_[50247]_ ,
    \new_[50248]_ , \new_[50252]_ , \new_[50253]_ , \new_[50257]_ ,
    \new_[50258]_ , \new_[50259]_ , \new_[50263]_ , \new_[50264]_ ,
    \new_[50267]_ , \new_[50270]_ , \new_[50271]_ , \new_[50272]_ ,
    \new_[50276]_ , \new_[50277]_ , \new_[50281]_ , \new_[50282]_ ,
    \new_[50283]_ , \new_[50287]_ , \new_[50288]_ , \new_[50291]_ ,
    \new_[50294]_ , \new_[50295]_ , \new_[50296]_ , \new_[50300]_ ,
    \new_[50301]_ , \new_[50305]_ , \new_[50306]_ , \new_[50307]_ ,
    \new_[50311]_ , \new_[50312]_ , \new_[50315]_ , \new_[50318]_ ,
    \new_[50319]_ , \new_[50320]_ , \new_[50324]_ , \new_[50325]_ ,
    \new_[50329]_ , \new_[50330]_ , \new_[50331]_ , \new_[50335]_ ,
    \new_[50336]_ , \new_[50339]_ , \new_[50342]_ , \new_[50343]_ ,
    \new_[50344]_ , \new_[50348]_ , \new_[50349]_ , \new_[50353]_ ,
    \new_[50354]_ , \new_[50355]_ , \new_[50359]_ , \new_[50360]_ ,
    \new_[50363]_ , \new_[50366]_ , \new_[50367]_ , \new_[50368]_ ,
    \new_[50372]_ , \new_[50373]_ , \new_[50377]_ , \new_[50378]_ ,
    \new_[50379]_ , \new_[50383]_ , \new_[50384]_ , \new_[50387]_ ,
    \new_[50390]_ , \new_[50391]_ , \new_[50392]_ , \new_[50396]_ ,
    \new_[50397]_ , \new_[50401]_ , \new_[50402]_ , \new_[50403]_ ,
    \new_[50407]_ , \new_[50408]_ , \new_[50411]_ , \new_[50414]_ ,
    \new_[50415]_ , \new_[50416]_ , \new_[50420]_ , \new_[50421]_ ,
    \new_[50425]_ , \new_[50426]_ , \new_[50427]_ , \new_[50431]_ ,
    \new_[50432]_ , \new_[50435]_ , \new_[50438]_ , \new_[50439]_ ,
    \new_[50440]_ , \new_[50444]_ , \new_[50445]_ , \new_[50449]_ ,
    \new_[50450]_ , \new_[50451]_ , \new_[50455]_ , \new_[50456]_ ,
    \new_[50459]_ , \new_[50462]_ , \new_[50463]_ , \new_[50464]_ ,
    \new_[50468]_ , \new_[50469]_ , \new_[50473]_ , \new_[50474]_ ,
    \new_[50475]_ , \new_[50479]_ , \new_[50480]_ , \new_[50483]_ ,
    \new_[50486]_ , \new_[50487]_ , \new_[50488]_ , \new_[50492]_ ,
    \new_[50493]_ , \new_[50497]_ , \new_[50498]_ , \new_[50499]_ ,
    \new_[50503]_ , \new_[50504]_ , \new_[50507]_ , \new_[50510]_ ,
    \new_[50511]_ , \new_[50512]_ , \new_[50516]_ , \new_[50517]_ ,
    \new_[50521]_ , \new_[50522]_ , \new_[50523]_ , \new_[50527]_ ,
    \new_[50528]_ , \new_[50531]_ , \new_[50534]_ , \new_[50535]_ ,
    \new_[50536]_ , \new_[50540]_ , \new_[50541]_ , \new_[50545]_ ,
    \new_[50546]_ , \new_[50547]_ , \new_[50551]_ , \new_[50552]_ ,
    \new_[50555]_ , \new_[50558]_ , \new_[50559]_ , \new_[50560]_ ,
    \new_[50564]_ , \new_[50565]_ , \new_[50569]_ , \new_[50570]_ ,
    \new_[50571]_ , \new_[50575]_ , \new_[50576]_ , \new_[50579]_ ,
    \new_[50582]_ , \new_[50583]_ , \new_[50584]_ , \new_[50588]_ ,
    \new_[50589]_ , \new_[50593]_ , \new_[50594]_ , \new_[50595]_ ,
    \new_[50599]_ , \new_[50600]_ , \new_[50603]_ , \new_[50606]_ ,
    \new_[50607]_ , \new_[50608]_ , \new_[50612]_ , \new_[50613]_ ,
    \new_[50617]_ , \new_[50618]_ , \new_[50619]_ , \new_[50623]_ ,
    \new_[50624]_ , \new_[50627]_ , \new_[50630]_ , \new_[50631]_ ,
    \new_[50632]_ , \new_[50636]_ , \new_[50637]_ , \new_[50641]_ ,
    \new_[50642]_ , \new_[50643]_ , \new_[50647]_ , \new_[50648]_ ,
    \new_[50651]_ , \new_[50654]_ , \new_[50655]_ , \new_[50656]_ ,
    \new_[50660]_ , \new_[50661]_ , \new_[50665]_ , \new_[50666]_ ,
    \new_[50667]_ , \new_[50671]_ , \new_[50672]_ , \new_[50675]_ ,
    \new_[50678]_ , \new_[50679]_ , \new_[50680]_ , \new_[50684]_ ,
    \new_[50685]_ , \new_[50689]_ , \new_[50690]_ , \new_[50691]_ ,
    \new_[50695]_ , \new_[50696]_ , \new_[50699]_ , \new_[50702]_ ,
    \new_[50703]_ , \new_[50704]_ , \new_[50708]_ , \new_[50709]_ ,
    \new_[50713]_ , \new_[50714]_ , \new_[50715]_ , \new_[50719]_ ,
    \new_[50720]_ , \new_[50723]_ , \new_[50726]_ , \new_[50727]_ ,
    \new_[50728]_ , \new_[50732]_ , \new_[50733]_ , \new_[50737]_ ,
    \new_[50738]_ , \new_[50739]_ , \new_[50743]_ , \new_[50744]_ ,
    \new_[50747]_ , \new_[50750]_ , \new_[50751]_ , \new_[50752]_ ,
    \new_[50756]_ , \new_[50757]_ , \new_[50761]_ , \new_[50762]_ ,
    \new_[50763]_ , \new_[50767]_ , \new_[50768]_ , \new_[50771]_ ,
    \new_[50774]_ , \new_[50775]_ , \new_[50776]_ , \new_[50780]_ ,
    \new_[50781]_ , \new_[50785]_ , \new_[50786]_ , \new_[50787]_ ,
    \new_[50791]_ , \new_[50792]_ , \new_[50795]_ , \new_[50798]_ ,
    \new_[50799]_ , \new_[50800]_ , \new_[50804]_ , \new_[50805]_ ,
    \new_[50809]_ , \new_[50810]_ , \new_[50811]_ , \new_[50815]_ ,
    \new_[50816]_ , \new_[50819]_ , \new_[50822]_ , \new_[50823]_ ,
    \new_[50824]_ , \new_[50828]_ , \new_[50829]_ , \new_[50833]_ ,
    \new_[50834]_ , \new_[50835]_ , \new_[50839]_ , \new_[50840]_ ,
    \new_[50843]_ , \new_[50846]_ , \new_[50847]_ , \new_[50848]_ ,
    \new_[50852]_ , \new_[50853]_ , \new_[50857]_ , \new_[50858]_ ,
    \new_[50859]_ , \new_[50863]_ , \new_[50864]_ , \new_[50867]_ ,
    \new_[50870]_ , \new_[50871]_ , \new_[50872]_ , \new_[50876]_ ,
    \new_[50877]_ , \new_[50881]_ , \new_[50882]_ , \new_[50883]_ ,
    \new_[50887]_ , \new_[50888]_ , \new_[50891]_ , \new_[50894]_ ,
    \new_[50895]_ , \new_[50896]_ , \new_[50900]_ , \new_[50901]_ ,
    \new_[50905]_ , \new_[50906]_ , \new_[50907]_ , \new_[50911]_ ,
    \new_[50912]_ , \new_[50915]_ , \new_[50918]_ , \new_[50919]_ ,
    \new_[50920]_ , \new_[50924]_ , \new_[50925]_ , \new_[50929]_ ,
    \new_[50930]_ , \new_[50931]_ , \new_[50935]_ , \new_[50936]_ ,
    \new_[50939]_ , \new_[50942]_ , \new_[50943]_ , \new_[50944]_ ,
    \new_[50948]_ , \new_[50949]_ , \new_[50953]_ , \new_[50954]_ ,
    \new_[50955]_ , \new_[50959]_ , \new_[50960]_ , \new_[50963]_ ,
    \new_[50966]_ , \new_[50967]_ , \new_[50968]_ , \new_[50972]_ ,
    \new_[50973]_ , \new_[50977]_ , \new_[50978]_ , \new_[50979]_ ,
    \new_[50983]_ , \new_[50984]_ , \new_[50987]_ , \new_[50990]_ ,
    \new_[50991]_ , \new_[50992]_ , \new_[50996]_ , \new_[50997]_ ,
    \new_[51001]_ , \new_[51002]_ , \new_[51003]_ , \new_[51007]_ ,
    \new_[51008]_ , \new_[51011]_ , \new_[51014]_ , \new_[51015]_ ,
    \new_[51016]_ , \new_[51020]_ , \new_[51021]_ , \new_[51025]_ ,
    \new_[51026]_ , \new_[51027]_ , \new_[51031]_ , \new_[51032]_ ,
    \new_[51035]_ , \new_[51038]_ , \new_[51039]_ , \new_[51040]_ ,
    \new_[51044]_ , \new_[51045]_ , \new_[51049]_ , \new_[51050]_ ,
    \new_[51051]_ , \new_[51055]_ , \new_[51056]_ , \new_[51059]_ ,
    \new_[51062]_ , \new_[51063]_ , \new_[51064]_ , \new_[51068]_ ,
    \new_[51069]_ , \new_[51073]_ , \new_[51074]_ , \new_[51075]_ ,
    \new_[51079]_ , \new_[51080]_ , \new_[51083]_ , \new_[51086]_ ,
    \new_[51087]_ , \new_[51088]_ , \new_[51092]_ , \new_[51093]_ ,
    \new_[51097]_ , \new_[51098]_ , \new_[51099]_ , \new_[51103]_ ,
    \new_[51104]_ , \new_[51107]_ , \new_[51110]_ , \new_[51111]_ ,
    \new_[51112]_ , \new_[51116]_ , \new_[51117]_ , \new_[51121]_ ,
    \new_[51122]_ , \new_[51123]_ , \new_[51127]_ , \new_[51128]_ ,
    \new_[51131]_ , \new_[51134]_ , \new_[51135]_ , \new_[51136]_ ,
    \new_[51140]_ , \new_[51141]_ , \new_[51145]_ , \new_[51146]_ ,
    \new_[51147]_ , \new_[51151]_ , \new_[51152]_ , \new_[51155]_ ,
    \new_[51158]_ , \new_[51159]_ , \new_[51160]_ , \new_[51164]_ ,
    \new_[51165]_ , \new_[51169]_ , \new_[51170]_ , \new_[51171]_ ,
    \new_[51175]_ , \new_[51176]_ , \new_[51179]_ , \new_[51182]_ ,
    \new_[51183]_ , \new_[51184]_ , \new_[51188]_ , \new_[51189]_ ,
    \new_[51193]_ , \new_[51194]_ , \new_[51195]_ , \new_[51199]_ ,
    \new_[51200]_ , \new_[51203]_ , \new_[51206]_ , \new_[51207]_ ,
    \new_[51208]_ , \new_[51212]_ , \new_[51213]_ , \new_[51217]_ ,
    \new_[51218]_ , \new_[51219]_ , \new_[51223]_ , \new_[51224]_ ,
    \new_[51227]_ , \new_[51230]_ , \new_[51231]_ , \new_[51232]_ ,
    \new_[51236]_ , \new_[51237]_ , \new_[51241]_ , \new_[51242]_ ,
    \new_[51243]_ , \new_[51247]_ , \new_[51248]_ , \new_[51251]_ ,
    \new_[51254]_ , \new_[51255]_ , \new_[51256]_ , \new_[51260]_ ,
    \new_[51261]_ , \new_[51265]_ , \new_[51266]_ , \new_[51267]_ ,
    \new_[51271]_ , \new_[51272]_ , \new_[51275]_ , \new_[51278]_ ,
    \new_[51279]_ , \new_[51280]_ , \new_[51284]_ , \new_[51285]_ ,
    \new_[51289]_ , \new_[51290]_ , \new_[51291]_ , \new_[51295]_ ,
    \new_[51296]_ , \new_[51299]_ , \new_[51302]_ , \new_[51303]_ ,
    \new_[51304]_ , \new_[51308]_ , \new_[51309]_ , \new_[51313]_ ,
    \new_[51314]_ , \new_[51315]_ , \new_[51319]_ , \new_[51320]_ ,
    \new_[51323]_ , \new_[51326]_ , \new_[51327]_ , \new_[51328]_ ,
    \new_[51332]_ , \new_[51333]_ , \new_[51337]_ , \new_[51338]_ ,
    \new_[51339]_ , \new_[51343]_ , \new_[51344]_ , \new_[51347]_ ,
    \new_[51350]_ , \new_[51351]_ , \new_[51352]_ , \new_[51356]_ ,
    \new_[51357]_ , \new_[51361]_ , \new_[51362]_ , \new_[51363]_ ,
    \new_[51367]_ , \new_[51368]_ , \new_[51371]_ , \new_[51374]_ ,
    \new_[51375]_ , \new_[51376]_ , \new_[51380]_ , \new_[51381]_ ,
    \new_[51385]_ , \new_[51386]_ , \new_[51387]_ , \new_[51391]_ ,
    \new_[51392]_ , \new_[51395]_ , \new_[51398]_ , \new_[51399]_ ,
    \new_[51400]_ , \new_[51404]_ , \new_[51405]_ , \new_[51409]_ ,
    \new_[51410]_ , \new_[51411]_ , \new_[51415]_ , \new_[51416]_ ,
    \new_[51419]_ , \new_[51422]_ , \new_[51423]_ , \new_[51424]_ ,
    \new_[51428]_ , \new_[51429]_ , \new_[51433]_ , \new_[51434]_ ,
    \new_[51435]_ , \new_[51439]_ , \new_[51440]_ , \new_[51443]_ ,
    \new_[51446]_ , \new_[51447]_ , \new_[51448]_ , \new_[51452]_ ,
    \new_[51453]_ , \new_[51457]_ , \new_[51458]_ , \new_[51459]_ ,
    \new_[51463]_ , \new_[51464]_ , \new_[51467]_ , \new_[51470]_ ,
    \new_[51471]_ , \new_[51472]_ , \new_[51476]_ , \new_[51477]_ ,
    \new_[51481]_ , \new_[51482]_ , \new_[51483]_ , \new_[51487]_ ,
    \new_[51488]_ , \new_[51491]_ , \new_[51494]_ , \new_[51495]_ ,
    \new_[51496]_ , \new_[51500]_ , \new_[51501]_ , \new_[51505]_ ,
    \new_[51506]_ , \new_[51507]_ , \new_[51511]_ , \new_[51512]_ ,
    \new_[51515]_ , \new_[51518]_ , \new_[51519]_ , \new_[51520]_ ,
    \new_[51524]_ , \new_[51525]_ , \new_[51529]_ , \new_[51530]_ ,
    \new_[51531]_ , \new_[51535]_ , \new_[51536]_ , \new_[51539]_ ,
    \new_[51542]_ , \new_[51543]_ , \new_[51544]_ , \new_[51548]_ ,
    \new_[51549]_ , \new_[51553]_ , \new_[51554]_ , \new_[51555]_ ,
    \new_[51559]_ , \new_[51560]_ , \new_[51563]_ , \new_[51566]_ ,
    \new_[51567]_ , \new_[51568]_ , \new_[51572]_ , \new_[51573]_ ,
    \new_[51577]_ , \new_[51578]_ , \new_[51579]_ , \new_[51583]_ ,
    \new_[51584]_ , \new_[51587]_ , \new_[51590]_ , \new_[51591]_ ,
    \new_[51592]_ , \new_[51596]_ , \new_[51597]_ , \new_[51601]_ ,
    \new_[51602]_ , \new_[51603]_ , \new_[51607]_ , \new_[51608]_ ,
    \new_[51611]_ , \new_[51614]_ , \new_[51615]_ , \new_[51616]_ ,
    \new_[51620]_ , \new_[51621]_ , \new_[51625]_ , \new_[51626]_ ,
    \new_[51627]_ , \new_[51631]_ , \new_[51632]_ , \new_[51635]_ ,
    \new_[51638]_ , \new_[51639]_ , \new_[51640]_ , \new_[51644]_ ,
    \new_[51645]_ , \new_[51649]_ , \new_[51650]_ , \new_[51651]_ ,
    \new_[51655]_ , \new_[51656]_ , \new_[51659]_ , \new_[51662]_ ,
    \new_[51663]_ , \new_[51664]_ , \new_[51668]_ , \new_[51669]_ ,
    \new_[51673]_ , \new_[51674]_ , \new_[51675]_ , \new_[51679]_ ,
    \new_[51680]_ , \new_[51683]_ , \new_[51686]_ , \new_[51687]_ ,
    \new_[51688]_ , \new_[51692]_ , \new_[51693]_ , \new_[51697]_ ,
    \new_[51698]_ , \new_[51699]_ , \new_[51703]_ , \new_[51704]_ ,
    \new_[51707]_ , \new_[51710]_ , \new_[51711]_ , \new_[51712]_ ,
    \new_[51716]_ , \new_[51717]_ , \new_[51721]_ , \new_[51722]_ ,
    \new_[51723]_ , \new_[51727]_ , \new_[51728]_ , \new_[51731]_ ,
    \new_[51734]_ , \new_[51735]_ , \new_[51736]_ , \new_[51740]_ ,
    \new_[51741]_ , \new_[51745]_ , \new_[51746]_ , \new_[51747]_ ,
    \new_[51751]_ , \new_[51752]_ , \new_[51755]_ , \new_[51758]_ ,
    \new_[51759]_ , \new_[51760]_ , \new_[51764]_ , \new_[51765]_ ,
    \new_[51769]_ , \new_[51770]_ , \new_[51771]_ , \new_[51775]_ ,
    \new_[51776]_ , \new_[51779]_ , \new_[51782]_ , \new_[51783]_ ,
    \new_[51784]_ , \new_[51788]_ , \new_[51789]_ , \new_[51793]_ ,
    \new_[51794]_ , \new_[51795]_ , \new_[51799]_ , \new_[51800]_ ,
    \new_[51803]_ , \new_[51806]_ , \new_[51807]_ , \new_[51808]_ ,
    \new_[51812]_ , \new_[51813]_ , \new_[51817]_ , \new_[51818]_ ,
    \new_[51819]_ , \new_[51823]_ , \new_[51824]_ , \new_[51827]_ ,
    \new_[51830]_ , \new_[51831]_ , \new_[51832]_ , \new_[51836]_ ,
    \new_[51837]_ , \new_[51841]_ , \new_[51842]_ , \new_[51843]_ ,
    \new_[51847]_ , \new_[51848]_ , \new_[51851]_ , \new_[51854]_ ,
    \new_[51855]_ , \new_[51856]_ , \new_[51860]_ , \new_[51861]_ ,
    \new_[51865]_ , \new_[51866]_ , \new_[51867]_ , \new_[51871]_ ,
    \new_[51872]_ , \new_[51875]_ , \new_[51878]_ , \new_[51879]_ ,
    \new_[51880]_ , \new_[51884]_ , \new_[51885]_ , \new_[51889]_ ,
    \new_[51890]_ , \new_[51891]_ , \new_[51895]_ , \new_[51896]_ ,
    \new_[51899]_ , \new_[51902]_ , \new_[51903]_ , \new_[51904]_ ,
    \new_[51908]_ , \new_[51909]_ , \new_[51913]_ , \new_[51914]_ ,
    \new_[51915]_ , \new_[51919]_ , \new_[51920]_ , \new_[51923]_ ,
    \new_[51926]_ , \new_[51927]_ , \new_[51928]_ , \new_[51932]_ ,
    \new_[51933]_ , \new_[51937]_ , \new_[51938]_ , \new_[51939]_ ,
    \new_[51943]_ , \new_[51944]_ , \new_[51947]_ , \new_[51950]_ ,
    \new_[51951]_ , \new_[51952]_ , \new_[51956]_ , \new_[51957]_ ,
    \new_[51961]_ , \new_[51962]_ , \new_[51963]_ , \new_[51967]_ ,
    \new_[51968]_ , \new_[51971]_ , \new_[51974]_ , \new_[51975]_ ,
    \new_[51976]_ , \new_[51980]_ , \new_[51981]_ , \new_[51985]_ ,
    \new_[51986]_ , \new_[51987]_ , \new_[51991]_ , \new_[51992]_ ,
    \new_[51995]_ , \new_[51998]_ , \new_[51999]_ , \new_[52000]_ ,
    \new_[52004]_ , \new_[52005]_ , \new_[52009]_ , \new_[52010]_ ,
    \new_[52011]_ , \new_[52015]_ , \new_[52016]_ , \new_[52019]_ ,
    \new_[52022]_ , \new_[52023]_ , \new_[52024]_ , \new_[52028]_ ,
    \new_[52029]_ , \new_[52033]_ , \new_[52034]_ , \new_[52035]_ ,
    \new_[52039]_ , \new_[52040]_ , \new_[52043]_ , \new_[52046]_ ,
    \new_[52047]_ , \new_[52048]_ , \new_[52052]_ , \new_[52053]_ ,
    \new_[52057]_ , \new_[52058]_ , \new_[52059]_ , \new_[52063]_ ,
    \new_[52064]_ , \new_[52067]_ , \new_[52070]_ , \new_[52071]_ ,
    \new_[52072]_ , \new_[52076]_ , \new_[52077]_ , \new_[52081]_ ,
    \new_[52082]_ , \new_[52083]_ , \new_[52087]_ , \new_[52088]_ ,
    \new_[52091]_ , \new_[52094]_ , \new_[52095]_ , \new_[52096]_ ,
    \new_[52100]_ , \new_[52101]_ , \new_[52105]_ , \new_[52106]_ ,
    \new_[52107]_ , \new_[52111]_ , \new_[52112]_ , \new_[52115]_ ,
    \new_[52118]_ , \new_[52119]_ , \new_[52120]_ , \new_[52124]_ ,
    \new_[52125]_ , \new_[52129]_ , \new_[52130]_ , \new_[52131]_ ,
    \new_[52135]_ , \new_[52136]_ , \new_[52139]_ , \new_[52142]_ ,
    \new_[52143]_ , \new_[52144]_ , \new_[52148]_ , \new_[52149]_ ,
    \new_[52153]_ , \new_[52154]_ , \new_[52155]_ , \new_[52159]_ ,
    \new_[52160]_ , \new_[52163]_ , \new_[52166]_ , \new_[52167]_ ,
    \new_[52168]_ , \new_[52172]_ , \new_[52173]_ , \new_[52177]_ ,
    \new_[52178]_ , \new_[52179]_ , \new_[52183]_ , \new_[52184]_ ,
    \new_[52187]_ , \new_[52190]_ , \new_[52191]_ , \new_[52192]_ ,
    \new_[52196]_ , \new_[52197]_ , \new_[52201]_ , \new_[52202]_ ,
    \new_[52203]_ , \new_[52207]_ , \new_[52208]_ , \new_[52211]_ ,
    \new_[52214]_ , \new_[52215]_ , \new_[52216]_ , \new_[52220]_ ,
    \new_[52221]_ , \new_[52225]_ , \new_[52226]_ , \new_[52227]_ ,
    \new_[52231]_ , \new_[52232]_ , \new_[52235]_ , \new_[52238]_ ,
    \new_[52239]_ , \new_[52240]_ , \new_[52244]_ , \new_[52245]_ ,
    \new_[52249]_ , \new_[52250]_ , \new_[52251]_ , \new_[52255]_ ,
    \new_[52256]_ , \new_[52259]_ , \new_[52262]_ , \new_[52263]_ ,
    \new_[52264]_ , \new_[52268]_ , \new_[52269]_ , \new_[52273]_ ,
    \new_[52274]_ , \new_[52275]_ , \new_[52279]_ , \new_[52280]_ ,
    \new_[52283]_ , \new_[52286]_ , \new_[52287]_ , \new_[52288]_ ,
    \new_[52292]_ , \new_[52293]_ , \new_[52297]_ , \new_[52298]_ ,
    \new_[52299]_ , \new_[52303]_ , \new_[52304]_ , \new_[52307]_ ,
    \new_[52310]_ , \new_[52311]_ , \new_[52312]_ , \new_[52316]_ ,
    \new_[52317]_ , \new_[52321]_ , \new_[52322]_ , \new_[52323]_ ,
    \new_[52327]_ , \new_[52328]_ , \new_[52331]_ , \new_[52334]_ ,
    \new_[52335]_ , \new_[52336]_ , \new_[52340]_ , \new_[52341]_ ,
    \new_[52345]_ , \new_[52346]_ , \new_[52347]_ , \new_[52351]_ ,
    \new_[52352]_ , \new_[52355]_ , \new_[52358]_ , \new_[52359]_ ,
    \new_[52360]_ , \new_[52364]_ , \new_[52365]_ , \new_[52369]_ ,
    \new_[52370]_ , \new_[52371]_ , \new_[52375]_ , \new_[52376]_ ,
    \new_[52379]_ , \new_[52382]_ , \new_[52383]_ , \new_[52384]_ ,
    \new_[52388]_ , \new_[52389]_ , \new_[52393]_ , \new_[52394]_ ,
    \new_[52395]_ , \new_[52399]_ , \new_[52400]_ , \new_[52403]_ ,
    \new_[52406]_ , \new_[52407]_ , \new_[52408]_ , \new_[52412]_ ,
    \new_[52413]_ , \new_[52417]_ , \new_[52418]_ , \new_[52419]_ ,
    \new_[52423]_ , \new_[52424]_ , \new_[52427]_ , \new_[52430]_ ,
    \new_[52431]_ , \new_[52432]_ , \new_[52436]_ , \new_[52437]_ ,
    \new_[52441]_ , \new_[52442]_ , \new_[52443]_ , \new_[52447]_ ,
    \new_[52448]_ , \new_[52451]_ , \new_[52454]_ , \new_[52455]_ ,
    \new_[52456]_ , \new_[52460]_ , \new_[52461]_ , \new_[52465]_ ,
    \new_[52466]_ , \new_[52467]_ , \new_[52471]_ , \new_[52472]_ ,
    \new_[52475]_ , \new_[52478]_ , \new_[52479]_ , \new_[52480]_ ,
    \new_[52484]_ , \new_[52485]_ , \new_[52489]_ , \new_[52490]_ ,
    \new_[52491]_ , \new_[52495]_ , \new_[52496]_ , \new_[52499]_ ,
    \new_[52502]_ , \new_[52503]_ , \new_[52504]_ , \new_[52508]_ ,
    \new_[52509]_ , \new_[52513]_ , \new_[52514]_ , \new_[52515]_ ,
    \new_[52519]_ , \new_[52520]_ , \new_[52523]_ , \new_[52526]_ ,
    \new_[52527]_ , \new_[52528]_ , \new_[52532]_ , \new_[52533]_ ,
    \new_[52537]_ , \new_[52538]_ , \new_[52539]_ , \new_[52543]_ ,
    \new_[52544]_ , \new_[52547]_ , \new_[52550]_ , \new_[52551]_ ,
    \new_[52552]_ , \new_[52556]_ , \new_[52557]_ , \new_[52561]_ ,
    \new_[52562]_ , \new_[52563]_ , \new_[52567]_ , \new_[52568]_ ,
    \new_[52571]_ , \new_[52574]_ , \new_[52575]_ , \new_[52576]_ ,
    \new_[52580]_ , \new_[52581]_ , \new_[52585]_ , \new_[52586]_ ,
    \new_[52587]_ , \new_[52591]_ , \new_[52592]_ , \new_[52595]_ ,
    \new_[52598]_ , \new_[52599]_ , \new_[52600]_ , \new_[52604]_ ,
    \new_[52605]_ , \new_[52609]_ , \new_[52610]_ , \new_[52611]_ ,
    \new_[52615]_ , \new_[52616]_ , \new_[52619]_ , \new_[52622]_ ,
    \new_[52623]_ , \new_[52624]_ , \new_[52628]_ , \new_[52629]_ ,
    \new_[52633]_ , \new_[52634]_ , \new_[52635]_ , \new_[52639]_ ,
    \new_[52640]_ , \new_[52643]_ , \new_[52646]_ , \new_[52647]_ ,
    \new_[52648]_ , \new_[52652]_ , \new_[52653]_ , \new_[52657]_ ,
    \new_[52658]_ , \new_[52659]_ , \new_[52663]_ , \new_[52664]_ ,
    \new_[52667]_ , \new_[52670]_ , \new_[52671]_ , \new_[52672]_ ,
    \new_[52676]_ , \new_[52677]_ , \new_[52681]_ , \new_[52682]_ ,
    \new_[52683]_ , \new_[52687]_ , \new_[52688]_ , \new_[52691]_ ,
    \new_[52694]_ , \new_[52695]_ , \new_[52696]_ , \new_[52700]_ ,
    \new_[52701]_ , \new_[52705]_ , \new_[52706]_ , \new_[52707]_ ,
    \new_[52711]_ , \new_[52712]_ , \new_[52715]_ , \new_[52718]_ ,
    \new_[52719]_ , \new_[52720]_ , \new_[52724]_ , \new_[52725]_ ,
    \new_[52729]_ , \new_[52730]_ , \new_[52731]_ , \new_[52735]_ ,
    \new_[52736]_ , \new_[52739]_ , \new_[52742]_ , \new_[52743]_ ,
    \new_[52744]_ , \new_[52748]_ , \new_[52749]_ , \new_[52753]_ ,
    \new_[52754]_ , \new_[52755]_ , \new_[52759]_ , \new_[52760]_ ,
    \new_[52763]_ , \new_[52766]_ , \new_[52767]_ , \new_[52768]_ ,
    \new_[52772]_ , \new_[52773]_ , \new_[52777]_ , \new_[52778]_ ,
    \new_[52779]_ , \new_[52783]_ , \new_[52784]_ , \new_[52787]_ ,
    \new_[52790]_ , \new_[52791]_ , \new_[52792]_ , \new_[52796]_ ,
    \new_[52797]_ , \new_[52801]_ , \new_[52802]_ , \new_[52803]_ ,
    \new_[52807]_ , \new_[52808]_ , \new_[52811]_ , \new_[52814]_ ,
    \new_[52815]_ , \new_[52816]_ , \new_[52820]_ , \new_[52821]_ ,
    \new_[52825]_ , \new_[52826]_ , \new_[52827]_ , \new_[52831]_ ,
    \new_[52832]_ , \new_[52835]_ , \new_[52838]_ , \new_[52839]_ ,
    \new_[52840]_ , \new_[52844]_ , \new_[52845]_ , \new_[52849]_ ,
    \new_[52850]_ , \new_[52851]_ , \new_[52855]_ , \new_[52856]_ ,
    \new_[52859]_ , \new_[52862]_ , \new_[52863]_ , \new_[52864]_ ,
    \new_[52868]_ , \new_[52869]_ , \new_[52873]_ , \new_[52874]_ ,
    \new_[52875]_ , \new_[52879]_ , \new_[52880]_ , \new_[52883]_ ,
    \new_[52886]_ , \new_[52887]_ , \new_[52888]_ , \new_[52892]_ ,
    \new_[52893]_ , \new_[52897]_ , \new_[52898]_ , \new_[52899]_ ,
    \new_[52903]_ , \new_[52904]_ , \new_[52907]_ , \new_[52910]_ ,
    \new_[52911]_ , \new_[52912]_ , \new_[52916]_ , \new_[52917]_ ,
    \new_[52921]_ , \new_[52922]_ , \new_[52923]_ , \new_[52927]_ ,
    \new_[52928]_ , \new_[52931]_ , \new_[52934]_ , \new_[52935]_ ,
    \new_[52936]_ , \new_[52940]_ , \new_[52941]_ , \new_[52945]_ ,
    \new_[52946]_ , \new_[52947]_ , \new_[52951]_ , \new_[52952]_ ,
    \new_[52955]_ , \new_[52958]_ , \new_[52959]_ , \new_[52960]_ ,
    \new_[52964]_ , \new_[52965]_ , \new_[52969]_ , \new_[52970]_ ,
    \new_[52971]_ , \new_[52975]_ , \new_[52976]_ , \new_[52979]_ ,
    \new_[52982]_ , \new_[52983]_ , \new_[52984]_ , \new_[52988]_ ,
    \new_[52989]_ , \new_[52993]_ , \new_[52994]_ , \new_[52995]_ ,
    \new_[52999]_ , \new_[53000]_ , \new_[53003]_ , \new_[53006]_ ,
    \new_[53007]_ , \new_[53008]_ , \new_[53012]_ , \new_[53013]_ ,
    \new_[53017]_ , \new_[53018]_ , \new_[53019]_ , \new_[53023]_ ,
    \new_[53024]_ , \new_[53027]_ , \new_[53030]_ , \new_[53031]_ ,
    \new_[53032]_ , \new_[53036]_ , \new_[53037]_ , \new_[53041]_ ,
    \new_[53042]_ , \new_[53043]_ , \new_[53047]_ , \new_[53048]_ ,
    \new_[53051]_ , \new_[53054]_ , \new_[53055]_ , \new_[53056]_ ,
    \new_[53060]_ , \new_[53061]_ , \new_[53065]_ , \new_[53066]_ ,
    \new_[53067]_ , \new_[53071]_ , \new_[53072]_ , \new_[53075]_ ,
    \new_[53078]_ , \new_[53079]_ , \new_[53080]_ , \new_[53084]_ ,
    \new_[53085]_ , \new_[53089]_ , \new_[53090]_ , \new_[53091]_ ,
    \new_[53095]_ , \new_[53096]_ , \new_[53099]_ , \new_[53102]_ ,
    \new_[53103]_ , \new_[53104]_ , \new_[53108]_ , \new_[53109]_ ,
    \new_[53113]_ , \new_[53114]_ , \new_[53115]_ , \new_[53119]_ ,
    \new_[53120]_ , \new_[53123]_ , \new_[53126]_ , \new_[53127]_ ,
    \new_[53128]_ , \new_[53132]_ , \new_[53133]_ , \new_[53137]_ ,
    \new_[53138]_ , \new_[53139]_ , \new_[53143]_ , \new_[53144]_ ,
    \new_[53147]_ , \new_[53150]_ , \new_[53151]_ , \new_[53152]_ ,
    \new_[53156]_ , \new_[53157]_ , \new_[53161]_ , \new_[53162]_ ,
    \new_[53163]_ , \new_[53167]_ , \new_[53168]_ , \new_[53171]_ ,
    \new_[53174]_ , \new_[53175]_ , \new_[53176]_ , \new_[53180]_ ,
    \new_[53181]_ , \new_[53185]_ , \new_[53186]_ , \new_[53187]_ ,
    \new_[53191]_ , \new_[53192]_ , \new_[53195]_ , \new_[53198]_ ,
    \new_[53199]_ , \new_[53200]_ , \new_[53204]_ , \new_[53205]_ ,
    \new_[53209]_ , \new_[53210]_ , \new_[53211]_ , \new_[53215]_ ,
    \new_[53216]_ , \new_[53219]_ , \new_[53222]_ , \new_[53223]_ ,
    \new_[53224]_ , \new_[53228]_ , \new_[53229]_ , \new_[53233]_ ,
    \new_[53234]_ , \new_[53235]_ , \new_[53239]_ , \new_[53240]_ ,
    \new_[53243]_ , \new_[53246]_ , \new_[53247]_ , \new_[53248]_ ,
    \new_[53252]_ , \new_[53253]_ , \new_[53257]_ , \new_[53258]_ ,
    \new_[53259]_ , \new_[53263]_ , \new_[53264]_ , \new_[53267]_ ,
    \new_[53270]_ , \new_[53271]_ , \new_[53272]_ , \new_[53276]_ ,
    \new_[53277]_ , \new_[53281]_ , \new_[53282]_ , \new_[53283]_ ,
    \new_[53287]_ , \new_[53288]_ , \new_[53291]_ , \new_[53294]_ ,
    \new_[53295]_ , \new_[53296]_ , \new_[53300]_ , \new_[53301]_ ,
    \new_[53305]_ , \new_[53306]_ , \new_[53307]_ , \new_[53311]_ ,
    \new_[53312]_ , \new_[53315]_ , \new_[53318]_ , \new_[53319]_ ,
    \new_[53320]_ , \new_[53324]_ , \new_[53325]_ , \new_[53329]_ ,
    \new_[53330]_ , \new_[53331]_ , \new_[53335]_ , \new_[53336]_ ,
    \new_[53339]_ , \new_[53342]_ , \new_[53343]_ , \new_[53344]_ ,
    \new_[53348]_ , \new_[53349]_ , \new_[53353]_ , \new_[53354]_ ,
    \new_[53355]_ , \new_[53359]_ , \new_[53360]_ , \new_[53363]_ ,
    \new_[53366]_ , \new_[53367]_ , \new_[53368]_ , \new_[53372]_ ,
    \new_[53373]_ , \new_[53377]_ , \new_[53378]_ , \new_[53379]_ ,
    \new_[53383]_ , \new_[53384]_ , \new_[53387]_ , \new_[53390]_ ,
    \new_[53391]_ , \new_[53392]_ , \new_[53396]_ , \new_[53397]_ ,
    \new_[53401]_ , \new_[53402]_ , \new_[53403]_ , \new_[53407]_ ,
    \new_[53408]_ , \new_[53411]_ , \new_[53414]_ , \new_[53415]_ ,
    \new_[53416]_ , \new_[53420]_ , \new_[53421]_ , \new_[53425]_ ,
    \new_[53426]_ , \new_[53427]_ , \new_[53431]_ , \new_[53432]_ ,
    \new_[53435]_ , \new_[53438]_ , \new_[53439]_ , \new_[53440]_ ,
    \new_[53444]_ , \new_[53445]_ , \new_[53449]_ , \new_[53450]_ ,
    \new_[53451]_ , \new_[53455]_ , \new_[53456]_ , \new_[53459]_ ,
    \new_[53462]_ , \new_[53463]_ , \new_[53464]_ , \new_[53468]_ ,
    \new_[53469]_ , \new_[53473]_ , \new_[53474]_ , \new_[53475]_ ,
    \new_[53479]_ , \new_[53480]_ , \new_[53483]_ , \new_[53486]_ ,
    \new_[53487]_ , \new_[53488]_ , \new_[53492]_ , \new_[53493]_ ,
    \new_[53497]_ , \new_[53498]_ , \new_[53499]_ , \new_[53503]_ ,
    \new_[53504]_ , \new_[53507]_ , \new_[53510]_ , \new_[53511]_ ,
    \new_[53512]_ , \new_[53516]_ , \new_[53517]_ , \new_[53521]_ ,
    \new_[53522]_ , \new_[53523]_ , \new_[53527]_ , \new_[53528]_ ,
    \new_[53531]_ , \new_[53534]_ , \new_[53535]_ , \new_[53536]_ ,
    \new_[53540]_ , \new_[53541]_ , \new_[53545]_ , \new_[53546]_ ,
    \new_[53547]_ , \new_[53551]_ , \new_[53552]_ , \new_[53555]_ ,
    \new_[53558]_ , \new_[53559]_ , \new_[53560]_ , \new_[53564]_ ,
    \new_[53565]_ , \new_[53569]_ , \new_[53570]_ , \new_[53571]_ ,
    \new_[53575]_ , \new_[53576]_ , \new_[53579]_ , \new_[53582]_ ,
    \new_[53583]_ , \new_[53584]_ , \new_[53588]_ , \new_[53589]_ ,
    \new_[53593]_ , \new_[53594]_ , \new_[53595]_ , \new_[53599]_ ,
    \new_[53600]_ , \new_[53603]_ , \new_[53606]_ , \new_[53607]_ ,
    \new_[53608]_ , \new_[53612]_ , \new_[53613]_ , \new_[53617]_ ,
    \new_[53618]_ , \new_[53619]_ , \new_[53623]_ , \new_[53624]_ ,
    \new_[53627]_ , \new_[53630]_ , \new_[53631]_ , \new_[53632]_ ,
    \new_[53636]_ , \new_[53637]_ , \new_[53641]_ , \new_[53642]_ ,
    \new_[53643]_ , \new_[53647]_ , \new_[53648]_ , \new_[53651]_ ,
    \new_[53654]_ , \new_[53655]_ , \new_[53656]_ , \new_[53660]_ ,
    \new_[53661]_ , \new_[53665]_ , \new_[53666]_ , \new_[53667]_ ,
    \new_[53671]_ , \new_[53672]_ , \new_[53675]_ , \new_[53678]_ ,
    \new_[53679]_ , \new_[53680]_ , \new_[53684]_ , \new_[53685]_ ,
    \new_[53689]_ , \new_[53690]_ , \new_[53691]_ , \new_[53695]_ ,
    \new_[53696]_ , \new_[53699]_ , \new_[53702]_ , \new_[53703]_ ,
    \new_[53704]_ , \new_[53708]_ , \new_[53709]_ , \new_[53713]_ ,
    \new_[53714]_ , \new_[53715]_ , \new_[53719]_ , \new_[53720]_ ,
    \new_[53723]_ , \new_[53726]_ , \new_[53727]_ , \new_[53728]_ ,
    \new_[53732]_ , \new_[53733]_ , \new_[53737]_ , \new_[53738]_ ,
    \new_[53739]_ , \new_[53743]_ , \new_[53744]_ , \new_[53747]_ ,
    \new_[53750]_ , \new_[53751]_ , \new_[53752]_ , \new_[53756]_ ,
    \new_[53757]_ , \new_[53761]_ , \new_[53762]_ , \new_[53763]_ ,
    \new_[53767]_ , \new_[53768]_ , \new_[53771]_ , \new_[53774]_ ,
    \new_[53775]_ , \new_[53776]_ , \new_[53780]_ , \new_[53781]_ ,
    \new_[53785]_ , \new_[53786]_ , \new_[53787]_ , \new_[53791]_ ,
    \new_[53792]_ , \new_[53795]_ , \new_[53798]_ , \new_[53799]_ ,
    \new_[53800]_ , \new_[53804]_ , \new_[53805]_ , \new_[53809]_ ,
    \new_[53810]_ , \new_[53811]_ , \new_[53815]_ , \new_[53816]_ ,
    \new_[53819]_ , \new_[53822]_ , \new_[53823]_ , \new_[53824]_ ,
    \new_[53828]_ , \new_[53829]_ , \new_[53833]_ , \new_[53834]_ ,
    \new_[53835]_ , \new_[53839]_ , \new_[53840]_ , \new_[53843]_ ,
    \new_[53846]_ , \new_[53847]_ , \new_[53848]_ , \new_[53852]_ ,
    \new_[53853]_ , \new_[53857]_ , \new_[53858]_ , \new_[53859]_ ,
    \new_[53863]_ , \new_[53864]_ , \new_[53867]_ , \new_[53870]_ ,
    \new_[53871]_ , \new_[53872]_ , \new_[53876]_ , \new_[53877]_ ,
    \new_[53881]_ , \new_[53882]_ , \new_[53883]_ , \new_[53887]_ ,
    \new_[53888]_ , \new_[53891]_ , \new_[53894]_ , \new_[53895]_ ,
    \new_[53896]_ , \new_[53900]_ , \new_[53901]_ , \new_[53905]_ ,
    \new_[53906]_ , \new_[53907]_ , \new_[53911]_ , \new_[53912]_ ,
    \new_[53915]_ , \new_[53918]_ , \new_[53919]_ , \new_[53920]_ ,
    \new_[53924]_ , \new_[53925]_ , \new_[53929]_ , \new_[53930]_ ,
    \new_[53931]_ , \new_[53935]_ , \new_[53936]_ , \new_[53939]_ ,
    \new_[53942]_ , \new_[53943]_ , \new_[53944]_ , \new_[53948]_ ,
    \new_[53949]_ , \new_[53953]_ , \new_[53954]_ , \new_[53955]_ ,
    \new_[53959]_ , \new_[53960]_ , \new_[53963]_ , \new_[53966]_ ,
    \new_[53967]_ , \new_[53968]_ , \new_[53972]_ , \new_[53973]_ ,
    \new_[53977]_ , \new_[53978]_ , \new_[53979]_ , \new_[53983]_ ,
    \new_[53984]_ , \new_[53987]_ , \new_[53990]_ , \new_[53991]_ ,
    \new_[53992]_ , \new_[53996]_ , \new_[53997]_ , \new_[54001]_ ,
    \new_[54002]_ , \new_[54003]_ , \new_[54007]_ , \new_[54008]_ ,
    \new_[54011]_ , \new_[54014]_ , \new_[54015]_ , \new_[54016]_ ,
    \new_[54020]_ , \new_[54021]_ , \new_[54025]_ , \new_[54026]_ ,
    \new_[54027]_ , \new_[54031]_ , \new_[54032]_ , \new_[54035]_ ,
    \new_[54038]_ , \new_[54039]_ , \new_[54040]_ , \new_[54044]_ ,
    \new_[54045]_ , \new_[54049]_ , \new_[54050]_ , \new_[54051]_ ,
    \new_[54055]_ , \new_[54056]_ , \new_[54059]_ , \new_[54062]_ ,
    \new_[54063]_ , \new_[54064]_ , \new_[54068]_ , \new_[54069]_ ,
    \new_[54073]_ , \new_[54074]_ , \new_[54075]_ , \new_[54079]_ ,
    \new_[54080]_ , \new_[54083]_ , \new_[54086]_ , \new_[54087]_ ,
    \new_[54088]_ , \new_[54092]_ , \new_[54093]_ , \new_[54097]_ ,
    \new_[54098]_ , \new_[54099]_ , \new_[54103]_ , \new_[54104]_ ,
    \new_[54107]_ , \new_[54110]_ , \new_[54111]_ , \new_[54112]_ ,
    \new_[54116]_ , \new_[54117]_ , \new_[54121]_ , \new_[54122]_ ,
    \new_[54123]_ , \new_[54127]_ , \new_[54128]_ , \new_[54131]_ ,
    \new_[54134]_ , \new_[54135]_ , \new_[54136]_ , \new_[54140]_ ,
    \new_[54141]_ , \new_[54145]_ , \new_[54146]_ , \new_[54147]_ ,
    \new_[54151]_ , \new_[54152]_ , \new_[54155]_ , \new_[54158]_ ,
    \new_[54159]_ , \new_[54160]_ , \new_[54164]_ , \new_[54165]_ ,
    \new_[54169]_ , \new_[54170]_ , \new_[54171]_ , \new_[54175]_ ,
    \new_[54176]_ , \new_[54179]_ , \new_[54182]_ , \new_[54183]_ ,
    \new_[54184]_ , \new_[54188]_ , \new_[54189]_ , \new_[54193]_ ,
    \new_[54194]_ , \new_[54195]_ , \new_[54199]_ , \new_[54200]_ ,
    \new_[54203]_ , \new_[54206]_ , \new_[54207]_ , \new_[54208]_ ,
    \new_[54212]_ , \new_[54213]_ , \new_[54217]_ , \new_[54218]_ ,
    \new_[54219]_ , \new_[54223]_ , \new_[54224]_ , \new_[54227]_ ,
    \new_[54230]_ , \new_[54231]_ , \new_[54232]_ , \new_[54236]_ ,
    \new_[54237]_ , \new_[54241]_ , \new_[54242]_ , \new_[54243]_ ,
    \new_[54247]_ , \new_[54248]_ , \new_[54251]_ , \new_[54254]_ ,
    \new_[54255]_ , \new_[54256]_ , \new_[54260]_ , \new_[54261]_ ,
    \new_[54265]_ , \new_[54266]_ , \new_[54267]_ , \new_[54271]_ ,
    \new_[54272]_ , \new_[54275]_ , \new_[54278]_ , \new_[54279]_ ,
    \new_[54280]_ , \new_[54284]_ , \new_[54285]_ , \new_[54289]_ ,
    \new_[54290]_ , \new_[54291]_ , \new_[54295]_ , \new_[54296]_ ,
    \new_[54299]_ , \new_[54302]_ , \new_[54303]_ , \new_[54304]_ ,
    \new_[54308]_ , \new_[54309]_ , \new_[54313]_ , \new_[54314]_ ,
    \new_[54315]_ , \new_[54319]_ , \new_[54320]_ , \new_[54323]_ ,
    \new_[54326]_ , \new_[54327]_ , \new_[54328]_ , \new_[54332]_ ,
    \new_[54333]_ , \new_[54337]_ , \new_[54338]_ , \new_[54339]_ ,
    \new_[54343]_ , \new_[54344]_ , \new_[54347]_ , \new_[54350]_ ,
    \new_[54351]_ , \new_[54352]_ , \new_[54356]_ , \new_[54357]_ ,
    \new_[54361]_ , \new_[54362]_ , \new_[54363]_ , \new_[54367]_ ,
    \new_[54368]_ , \new_[54371]_ , \new_[54374]_ , \new_[54375]_ ,
    \new_[54376]_ , \new_[54380]_ , \new_[54381]_ , \new_[54385]_ ,
    \new_[54386]_ , \new_[54387]_ , \new_[54391]_ , \new_[54392]_ ,
    \new_[54395]_ , \new_[54398]_ , \new_[54399]_ , \new_[54400]_ ,
    \new_[54404]_ , \new_[54405]_ , \new_[54409]_ , \new_[54410]_ ,
    \new_[54411]_ , \new_[54415]_ , \new_[54416]_ , \new_[54419]_ ,
    \new_[54422]_ , \new_[54423]_ , \new_[54424]_ , \new_[54428]_ ,
    \new_[54429]_ , \new_[54433]_ , \new_[54434]_ , \new_[54435]_ ,
    \new_[54439]_ , \new_[54440]_ , \new_[54443]_ , \new_[54446]_ ,
    \new_[54447]_ , \new_[54448]_ , \new_[54452]_ , \new_[54453]_ ,
    \new_[54457]_ , \new_[54458]_ , \new_[54459]_ , \new_[54463]_ ,
    \new_[54464]_ , \new_[54467]_ , \new_[54470]_ , \new_[54471]_ ,
    \new_[54472]_ , \new_[54476]_ , \new_[54477]_ , \new_[54481]_ ,
    \new_[54482]_ , \new_[54483]_ , \new_[54487]_ , \new_[54488]_ ,
    \new_[54491]_ , \new_[54494]_ , \new_[54495]_ , \new_[54496]_ ,
    \new_[54500]_ , \new_[54501]_ , \new_[54505]_ , \new_[54506]_ ,
    \new_[54507]_ , \new_[54511]_ , \new_[54512]_ , \new_[54515]_ ,
    \new_[54518]_ , \new_[54519]_ , \new_[54520]_ , \new_[54524]_ ,
    \new_[54525]_ , \new_[54529]_ , \new_[54530]_ , \new_[54531]_ ,
    \new_[54535]_ , \new_[54536]_ , \new_[54539]_ , \new_[54542]_ ,
    \new_[54543]_ , \new_[54544]_ , \new_[54548]_ , \new_[54549]_ ,
    \new_[54553]_ , \new_[54554]_ , \new_[54555]_ , \new_[54559]_ ,
    \new_[54560]_ , \new_[54563]_ , \new_[54566]_ , \new_[54567]_ ,
    \new_[54568]_ , \new_[54572]_ , \new_[54573]_ , \new_[54577]_ ,
    \new_[54578]_ , \new_[54579]_ , \new_[54583]_ , \new_[54584]_ ,
    \new_[54587]_ , \new_[54590]_ , \new_[54591]_ , \new_[54592]_ ,
    \new_[54596]_ , \new_[54597]_ , \new_[54601]_ , \new_[54602]_ ,
    \new_[54603]_ , \new_[54607]_ , \new_[54608]_ , \new_[54611]_ ,
    \new_[54614]_ , \new_[54615]_ , \new_[54616]_ , \new_[54620]_ ,
    \new_[54621]_ , \new_[54625]_ , \new_[54626]_ , \new_[54627]_ ,
    \new_[54631]_ , \new_[54632]_ , \new_[54635]_ , \new_[54638]_ ,
    \new_[54639]_ , \new_[54640]_ , \new_[54644]_ , \new_[54645]_ ,
    \new_[54649]_ , \new_[54650]_ , \new_[54651]_ , \new_[54655]_ ,
    \new_[54656]_ , \new_[54659]_ , \new_[54662]_ , \new_[54663]_ ,
    \new_[54664]_ , \new_[54668]_ , \new_[54669]_ , \new_[54673]_ ,
    \new_[54674]_ , \new_[54675]_ , \new_[54679]_ , \new_[54680]_ ,
    \new_[54683]_ , \new_[54686]_ , \new_[54687]_ , \new_[54688]_ ,
    \new_[54692]_ , \new_[54693]_ , \new_[54697]_ , \new_[54698]_ ,
    \new_[54699]_ , \new_[54703]_ , \new_[54704]_ , \new_[54707]_ ,
    \new_[54710]_ , \new_[54711]_ , \new_[54712]_ , \new_[54716]_ ,
    \new_[54717]_ , \new_[54721]_ , \new_[54722]_ , \new_[54723]_ ,
    \new_[54727]_ , \new_[54728]_ , \new_[54731]_ , \new_[54734]_ ,
    \new_[54735]_ , \new_[54736]_ , \new_[54740]_ , \new_[54741]_ ,
    \new_[54745]_ , \new_[54746]_ , \new_[54747]_ , \new_[54751]_ ,
    \new_[54752]_ , \new_[54755]_ , \new_[54758]_ , \new_[54759]_ ,
    \new_[54760]_ , \new_[54764]_ , \new_[54765]_ , \new_[54769]_ ,
    \new_[54770]_ , \new_[54771]_ , \new_[54775]_ , \new_[54776]_ ,
    \new_[54779]_ , \new_[54782]_ , \new_[54783]_ , \new_[54784]_ ,
    \new_[54788]_ , \new_[54789]_ , \new_[54793]_ , \new_[54794]_ ,
    \new_[54795]_ , \new_[54799]_ , \new_[54800]_ , \new_[54803]_ ,
    \new_[54806]_ , \new_[54807]_ , \new_[54808]_ , \new_[54812]_ ,
    \new_[54813]_ , \new_[54817]_ , \new_[54818]_ , \new_[54819]_ ,
    \new_[54823]_ , \new_[54824]_ , \new_[54827]_ , \new_[54830]_ ,
    \new_[54831]_ , \new_[54832]_ , \new_[54836]_ , \new_[54837]_ ,
    \new_[54841]_ , \new_[54842]_ , \new_[54843]_ , \new_[54847]_ ,
    \new_[54848]_ , \new_[54851]_ , \new_[54854]_ , \new_[54855]_ ,
    \new_[54856]_ , \new_[54860]_ , \new_[54861]_ , \new_[54865]_ ,
    \new_[54866]_ , \new_[54867]_ , \new_[54871]_ , \new_[54872]_ ,
    \new_[54875]_ , \new_[54878]_ , \new_[54879]_ , \new_[54880]_ ,
    \new_[54884]_ , \new_[54885]_ , \new_[54889]_ , \new_[54890]_ ,
    \new_[54891]_ , \new_[54895]_ , \new_[54896]_ , \new_[54899]_ ,
    \new_[54902]_ , \new_[54903]_ , \new_[54904]_ , \new_[54908]_ ,
    \new_[54909]_ , \new_[54913]_ , \new_[54914]_ , \new_[54915]_ ,
    \new_[54919]_ , \new_[54920]_ , \new_[54923]_ , \new_[54926]_ ,
    \new_[54927]_ , \new_[54928]_ , \new_[54932]_ , \new_[54933]_ ,
    \new_[54937]_ , \new_[54938]_ , \new_[54939]_ , \new_[54943]_ ,
    \new_[54944]_ , \new_[54947]_ , \new_[54950]_ , \new_[54951]_ ,
    \new_[54952]_ , \new_[54956]_ , \new_[54957]_ , \new_[54961]_ ,
    \new_[54962]_ , \new_[54963]_ , \new_[54967]_ , \new_[54968]_ ,
    \new_[54971]_ , \new_[54974]_ , \new_[54975]_ , \new_[54976]_ ,
    \new_[54980]_ , \new_[54981]_ , \new_[54985]_ , \new_[54986]_ ,
    \new_[54987]_ , \new_[54991]_ , \new_[54992]_ , \new_[54995]_ ,
    \new_[54998]_ , \new_[54999]_ , \new_[55000]_ , \new_[55004]_ ,
    \new_[55005]_ , \new_[55009]_ , \new_[55010]_ , \new_[55011]_ ,
    \new_[55015]_ , \new_[55016]_ , \new_[55019]_ , \new_[55022]_ ,
    \new_[55023]_ , \new_[55024]_ , \new_[55028]_ , \new_[55029]_ ,
    \new_[55033]_ , \new_[55034]_ , \new_[55035]_ , \new_[55039]_ ,
    \new_[55040]_ , \new_[55043]_ , \new_[55046]_ , \new_[55047]_ ,
    \new_[55048]_ , \new_[55052]_ , \new_[55053]_ , \new_[55057]_ ,
    \new_[55058]_ , \new_[55059]_ , \new_[55063]_ , \new_[55064]_ ,
    \new_[55067]_ , \new_[55070]_ , \new_[55071]_ , \new_[55072]_ ,
    \new_[55076]_ , \new_[55077]_ , \new_[55081]_ , \new_[55082]_ ,
    \new_[55083]_ , \new_[55087]_ , \new_[55088]_ , \new_[55091]_ ,
    \new_[55094]_ , \new_[55095]_ , \new_[55096]_ , \new_[55100]_ ,
    \new_[55101]_ , \new_[55105]_ , \new_[55106]_ , \new_[55107]_ ,
    \new_[55111]_ , \new_[55112]_ , \new_[55115]_ , \new_[55118]_ ,
    \new_[55119]_ , \new_[55120]_ , \new_[55124]_ , \new_[55125]_ ,
    \new_[55129]_ , \new_[55130]_ , \new_[55131]_ , \new_[55135]_ ,
    \new_[55136]_ , \new_[55139]_ , \new_[55142]_ , \new_[55143]_ ,
    \new_[55144]_ , \new_[55148]_ , \new_[55149]_ , \new_[55153]_ ,
    \new_[55154]_ , \new_[55155]_ , \new_[55159]_ , \new_[55160]_ ,
    \new_[55163]_ , \new_[55166]_ , \new_[55167]_ , \new_[55168]_ ,
    \new_[55172]_ , \new_[55173]_ , \new_[55177]_ , \new_[55178]_ ,
    \new_[55179]_ , \new_[55183]_ , \new_[55184]_ , \new_[55187]_ ,
    \new_[55190]_ , \new_[55191]_ , \new_[55192]_ , \new_[55196]_ ,
    \new_[55197]_ , \new_[55201]_ , \new_[55202]_ , \new_[55203]_ ,
    \new_[55207]_ , \new_[55208]_ , \new_[55211]_ , \new_[55214]_ ,
    \new_[55215]_ , \new_[55216]_ , \new_[55220]_ , \new_[55221]_ ,
    \new_[55225]_ , \new_[55226]_ , \new_[55227]_ , \new_[55231]_ ,
    \new_[55232]_ , \new_[55235]_ , \new_[55238]_ , \new_[55239]_ ,
    \new_[55240]_ , \new_[55244]_ , \new_[55245]_ , \new_[55249]_ ,
    \new_[55250]_ , \new_[55251]_ , \new_[55255]_ , \new_[55256]_ ,
    \new_[55259]_ , \new_[55262]_ , \new_[55263]_ , \new_[55264]_ ,
    \new_[55268]_ , \new_[55269]_ , \new_[55273]_ , \new_[55274]_ ,
    \new_[55275]_ , \new_[55279]_ , \new_[55280]_ , \new_[55283]_ ,
    \new_[55286]_ , \new_[55287]_ , \new_[55288]_ , \new_[55292]_ ,
    \new_[55293]_ , \new_[55297]_ , \new_[55298]_ , \new_[55299]_ ,
    \new_[55303]_ , \new_[55304]_ , \new_[55307]_ , \new_[55310]_ ,
    \new_[55311]_ , \new_[55312]_ , \new_[55316]_ , \new_[55317]_ ,
    \new_[55321]_ , \new_[55322]_ , \new_[55323]_ , \new_[55327]_ ,
    \new_[55328]_ , \new_[55331]_ , \new_[55334]_ , \new_[55335]_ ,
    \new_[55336]_ , \new_[55340]_ , \new_[55341]_ , \new_[55345]_ ,
    \new_[55346]_ , \new_[55347]_ , \new_[55351]_ , \new_[55352]_ ,
    \new_[55355]_ , \new_[55358]_ , \new_[55359]_ , \new_[55360]_ ,
    \new_[55364]_ , \new_[55365]_ , \new_[55369]_ , \new_[55370]_ ,
    \new_[55371]_ , \new_[55375]_ , \new_[55376]_ , \new_[55379]_ ,
    \new_[55382]_ , \new_[55383]_ , \new_[55384]_ , \new_[55388]_ ,
    \new_[55389]_ , \new_[55393]_ , \new_[55394]_ , \new_[55395]_ ,
    \new_[55399]_ , \new_[55400]_ , \new_[55403]_ , \new_[55406]_ ,
    \new_[55407]_ , \new_[55408]_ , \new_[55412]_ , \new_[55413]_ ,
    \new_[55417]_ , \new_[55418]_ , \new_[55419]_ , \new_[55423]_ ,
    \new_[55424]_ , \new_[55427]_ , \new_[55430]_ , \new_[55431]_ ,
    \new_[55432]_ , \new_[55436]_ , \new_[55437]_ , \new_[55441]_ ,
    \new_[55442]_ , \new_[55443]_ , \new_[55447]_ , \new_[55448]_ ,
    \new_[55451]_ , \new_[55454]_ , \new_[55455]_ , \new_[55456]_ ,
    \new_[55460]_ , \new_[55461]_ , \new_[55465]_ , \new_[55466]_ ,
    \new_[55467]_ , \new_[55471]_ , \new_[55472]_ , \new_[55475]_ ,
    \new_[55478]_ , \new_[55479]_ , \new_[55480]_ , \new_[55484]_ ,
    \new_[55485]_ , \new_[55489]_ , \new_[55490]_ , \new_[55491]_ ,
    \new_[55495]_ , \new_[55496]_ , \new_[55499]_ , \new_[55502]_ ,
    \new_[55503]_ , \new_[55504]_ , \new_[55508]_ , \new_[55509]_ ,
    \new_[55513]_ , \new_[55514]_ , \new_[55515]_ , \new_[55519]_ ,
    \new_[55520]_ , \new_[55523]_ , \new_[55526]_ , \new_[55527]_ ,
    \new_[55528]_ , \new_[55532]_ , \new_[55533]_ , \new_[55537]_ ,
    \new_[55538]_ , \new_[55539]_ , \new_[55543]_ , \new_[55544]_ ,
    \new_[55547]_ , \new_[55550]_ , \new_[55551]_ , \new_[55552]_ ,
    \new_[55556]_ , \new_[55557]_ , \new_[55561]_ , \new_[55562]_ ,
    \new_[55563]_ , \new_[55567]_ , \new_[55568]_ , \new_[55571]_ ,
    \new_[55574]_ , \new_[55575]_ , \new_[55576]_ , \new_[55580]_ ,
    \new_[55581]_ , \new_[55585]_ , \new_[55586]_ , \new_[55587]_ ,
    \new_[55591]_ , \new_[55592]_ , \new_[55595]_ , \new_[55598]_ ,
    \new_[55599]_ , \new_[55600]_ , \new_[55604]_ , \new_[55605]_ ,
    \new_[55609]_ , \new_[55610]_ , \new_[55611]_ , \new_[55615]_ ,
    \new_[55616]_ , \new_[55619]_ , \new_[55622]_ , \new_[55623]_ ,
    \new_[55624]_ , \new_[55628]_ , \new_[55629]_ , \new_[55633]_ ,
    \new_[55634]_ , \new_[55635]_ , \new_[55639]_ , \new_[55640]_ ,
    \new_[55643]_ , \new_[55646]_ , \new_[55647]_ , \new_[55648]_ ,
    \new_[55652]_ , \new_[55653]_ , \new_[55657]_ , \new_[55658]_ ,
    \new_[55659]_ , \new_[55663]_ , \new_[55664]_ , \new_[55667]_ ,
    \new_[55670]_ , \new_[55671]_ , \new_[55672]_ , \new_[55676]_ ,
    \new_[55677]_ , \new_[55681]_ , \new_[55682]_ , \new_[55683]_ ,
    \new_[55687]_ , \new_[55688]_ , \new_[55691]_ , \new_[55694]_ ,
    \new_[55695]_ , \new_[55696]_ , \new_[55700]_ , \new_[55701]_ ,
    \new_[55705]_ , \new_[55706]_ , \new_[55707]_ , \new_[55711]_ ,
    \new_[55712]_ , \new_[55715]_ , \new_[55718]_ , \new_[55719]_ ,
    \new_[55720]_ , \new_[55724]_ , \new_[55725]_ , \new_[55729]_ ,
    \new_[55730]_ , \new_[55731]_ , \new_[55735]_ , \new_[55736]_ ,
    \new_[55739]_ , \new_[55742]_ , \new_[55743]_ , \new_[55744]_ ,
    \new_[55748]_ , \new_[55749]_ , \new_[55753]_ , \new_[55754]_ ,
    \new_[55755]_ , \new_[55759]_ , \new_[55760]_ , \new_[55763]_ ,
    \new_[55766]_ , \new_[55767]_ , \new_[55768]_ , \new_[55772]_ ,
    \new_[55773]_ , \new_[55777]_ , \new_[55778]_ , \new_[55779]_ ,
    \new_[55783]_ , \new_[55784]_ , \new_[55787]_ , \new_[55790]_ ,
    \new_[55791]_ , \new_[55792]_ , \new_[55796]_ , \new_[55797]_ ,
    \new_[55801]_ , \new_[55802]_ , \new_[55803]_ , \new_[55807]_ ,
    \new_[55808]_ , \new_[55811]_ , \new_[55814]_ , \new_[55815]_ ,
    \new_[55816]_ , \new_[55820]_ , \new_[55821]_ , \new_[55825]_ ,
    \new_[55826]_ , \new_[55827]_ , \new_[55831]_ , \new_[55832]_ ,
    \new_[55835]_ , \new_[55838]_ , \new_[55839]_ , \new_[55840]_ ,
    \new_[55844]_ , \new_[55845]_ , \new_[55849]_ , \new_[55850]_ ,
    \new_[55851]_ , \new_[55855]_ , \new_[55856]_ , \new_[55859]_ ,
    \new_[55862]_ , \new_[55863]_ , \new_[55864]_ , \new_[55868]_ ,
    \new_[55869]_ , \new_[55873]_ , \new_[55874]_ , \new_[55875]_ ,
    \new_[55879]_ , \new_[55880]_ , \new_[55883]_ , \new_[55886]_ ,
    \new_[55887]_ , \new_[55888]_ , \new_[55892]_ , \new_[55893]_ ,
    \new_[55897]_ , \new_[55898]_ , \new_[55899]_ , \new_[55903]_ ,
    \new_[55904]_ , \new_[55907]_ , \new_[55910]_ , \new_[55911]_ ,
    \new_[55912]_ , \new_[55916]_ , \new_[55917]_ , \new_[55921]_ ,
    \new_[55922]_ , \new_[55923]_ , \new_[55927]_ , \new_[55928]_ ,
    \new_[55931]_ , \new_[55934]_ , \new_[55935]_ , \new_[55936]_ ,
    \new_[55940]_ , \new_[55941]_ , \new_[55945]_ , \new_[55946]_ ,
    \new_[55947]_ , \new_[55951]_ , \new_[55952]_ , \new_[55955]_ ,
    \new_[55958]_ , \new_[55959]_ , \new_[55960]_ , \new_[55964]_ ,
    \new_[55965]_ , \new_[55969]_ , \new_[55970]_ , \new_[55971]_ ,
    \new_[55975]_ , \new_[55976]_ , \new_[55979]_ , \new_[55982]_ ,
    \new_[55983]_ , \new_[55984]_ , \new_[55988]_ , \new_[55989]_ ,
    \new_[55993]_ , \new_[55994]_ , \new_[55995]_ , \new_[55999]_ ,
    \new_[56000]_ , \new_[56003]_ , \new_[56006]_ , \new_[56007]_ ,
    \new_[56008]_ , \new_[56012]_ , \new_[56013]_ , \new_[56017]_ ,
    \new_[56018]_ , \new_[56019]_ , \new_[56023]_ , \new_[56024]_ ,
    \new_[56027]_ , \new_[56030]_ , \new_[56031]_ , \new_[56032]_ ,
    \new_[56036]_ , \new_[56037]_ , \new_[56041]_ , \new_[56042]_ ,
    \new_[56043]_ , \new_[56047]_ , \new_[56048]_ , \new_[56051]_ ,
    \new_[56054]_ , \new_[56055]_ , \new_[56056]_ , \new_[56060]_ ,
    \new_[56061]_ , \new_[56065]_ , \new_[56066]_ , \new_[56067]_ ,
    \new_[56071]_ , \new_[56072]_ , \new_[56075]_ , \new_[56078]_ ,
    \new_[56079]_ , \new_[56080]_ , \new_[56084]_ , \new_[56085]_ ,
    \new_[56089]_ , \new_[56090]_ , \new_[56091]_ , \new_[56095]_ ,
    \new_[56096]_ , \new_[56099]_ , \new_[56102]_ , \new_[56103]_ ,
    \new_[56104]_ , \new_[56108]_ , \new_[56109]_ , \new_[56113]_ ,
    \new_[56114]_ , \new_[56115]_ , \new_[56119]_ , \new_[56120]_ ,
    \new_[56123]_ , \new_[56126]_ , \new_[56127]_ , \new_[56128]_ ,
    \new_[56132]_ , \new_[56133]_ , \new_[56137]_ , \new_[56138]_ ,
    \new_[56139]_ , \new_[56143]_ , \new_[56144]_ , \new_[56147]_ ,
    \new_[56150]_ , \new_[56151]_ , \new_[56152]_ , \new_[56156]_ ,
    \new_[56157]_ , \new_[56161]_ , \new_[56162]_ , \new_[56163]_ ,
    \new_[56167]_ , \new_[56168]_ , \new_[56171]_ , \new_[56174]_ ,
    \new_[56175]_ , \new_[56176]_ , \new_[56180]_ , \new_[56181]_ ,
    \new_[56185]_ , \new_[56186]_ , \new_[56187]_ , \new_[56191]_ ,
    \new_[56192]_ , \new_[56195]_ , \new_[56198]_ , \new_[56199]_ ,
    \new_[56200]_ , \new_[56204]_ , \new_[56205]_ , \new_[56209]_ ,
    \new_[56210]_ , \new_[56211]_ , \new_[56215]_ , \new_[56216]_ ,
    \new_[56219]_ , \new_[56222]_ , \new_[56223]_ , \new_[56224]_ ,
    \new_[56228]_ , \new_[56229]_ , \new_[56233]_ , \new_[56234]_ ,
    \new_[56235]_ , \new_[56239]_ , \new_[56240]_ , \new_[56243]_ ,
    \new_[56246]_ , \new_[56247]_ , \new_[56248]_ , \new_[56252]_ ,
    \new_[56253]_ , \new_[56257]_ , \new_[56258]_ , \new_[56259]_ ,
    \new_[56263]_ , \new_[56264]_ , \new_[56267]_ , \new_[56270]_ ,
    \new_[56271]_ , \new_[56272]_ , \new_[56276]_ , \new_[56277]_ ,
    \new_[56281]_ , \new_[56282]_ , \new_[56283]_ , \new_[56287]_ ,
    \new_[56288]_ , \new_[56291]_ , \new_[56294]_ , \new_[56295]_ ,
    \new_[56296]_ , \new_[56300]_ , \new_[56301]_ , \new_[56305]_ ,
    \new_[56306]_ , \new_[56307]_ , \new_[56311]_ , \new_[56312]_ ,
    \new_[56315]_ , \new_[56318]_ , \new_[56319]_ , \new_[56320]_ ,
    \new_[56324]_ , \new_[56325]_ , \new_[56329]_ , \new_[56330]_ ,
    \new_[56331]_ , \new_[56335]_ , \new_[56336]_ , \new_[56339]_ ,
    \new_[56342]_ , \new_[56343]_ , \new_[56344]_ , \new_[56348]_ ,
    \new_[56349]_ , \new_[56353]_ , \new_[56354]_ , \new_[56355]_ ,
    \new_[56359]_ , \new_[56360]_ , \new_[56363]_ , \new_[56366]_ ,
    \new_[56367]_ , \new_[56368]_ , \new_[56372]_ , \new_[56373]_ ,
    \new_[56377]_ , \new_[56378]_ , \new_[56379]_ , \new_[56383]_ ,
    \new_[56384]_ , \new_[56387]_ , \new_[56390]_ , \new_[56391]_ ,
    \new_[56392]_ , \new_[56396]_ , \new_[56397]_ , \new_[56401]_ ,
    \new_[56402]_ , \new_[56403]_ , \new_[56407]_ , \new_[56408]_ ,
    \new_[56411]_ , \new_[56414]_ , \new_[56415]_ , \new_[56416]_ ,
    \new_[56420]_ , \new_[56421]_ , \new_[56425]_ , \new_[56426]_ ,
    \new_[56427]_ , \new_[56431]_ , \new_[56432]_ , \new_[56435]_ ,
    \new_[56438]_ , \new_[56439]_ , \new_[56440]_ , \new_[56444]_ ,
    \new_[56445]_ , \new_[56449]_ , \new_[56450]_ , \new_[56451]_ ,
    \new_[56455]_ , \new_[56456]_ , \new_[56459]_ , \new_[56462]_ ,
    \new_[56463]_ , \new_[56464]_ , \new_[56468]_ , \new_[56469]_ ,
    \new_[56473]_ , \new_[56474]_ , \new_[56475]_ , \new_[56479]_ ,
    \new_[56480]_ , \new_[56483]_ , \new_[56486]_ , \new_[56487]_ ,
    \new_[56488]_ , \new_[56492]_ , \new_[56493]_ , \new_[56497]_ ,
    \new_[56498]_ , \new_[56499]_ , \new_[56503]_ , \new_[56504]_ ,
    \new_[56507]_ , \new_[56510]_ , \new_[56511]_ , \new_[56512]_ ,
    \new_[56516]_ , \new_[56517]_ , \new_[56521]_ , \new_[56522]_ ,
    \new_[56523]_ , \new_[56527]_ , \new_[56528]_ , \new_[56531]_ ,
    \new_[56534]_ , \new_[56535]_ , \new_[56536]_ , \new_[56540]_ ,
    \new_[56541]_ , \new_[56545]_ , \new_[56546]_ , \new_[56547]_ ,
    \new_[56551]_ , \new_[56552]_ , \new_[56555]_ , \new_[56558]_ ,
    \new_[56559]_ , \new_[56560]_ , \new_[56564]_ , \new_[56565]_ ,
    \new_[56569]_ , \new_[56570]_ , \new_[56571]_ , \new_[56575]_ ,
    \new_[56576]_ , \new_[56579]_ , \new_[56582]_ , \new_[56583]_ ,
    \new_[56584]_ , \new_[56588]_ , \new_[56589]_ , \new_[56593]_ ,
    \new_[56594]_ , \new_[56595]_ , \new_[56599]_ , \new_[56600]_ ,
    \new_[56603]_ , \new_[56606]_ , \new_[56607]_ , \new_[56608]_ ,
    \new_[56612]_ , \new_[56613]_ , \new_[56617]_ , \new_[56618]_ ,
    \new_[56619]_ , \new_[56623]_ , \new_[56624]_ , \new_[56627]_ ,
    \new_[56630]_ , \new_[56631]_ , \new_[56632]_ , \new_[56636]_ ,
    \new_[56637]_ , \new_[56641]_ , \new_[56642]_ , \new_[56643]_ ,
    \new_[56647]_ , \new_[56648]_ , \new_[56651]_ , \new_[56654]_ ,
    \new_[56655]_ , \new_[56656]_ , \new_[56660]_ , \new_[56661]_ ,
    \new_[56665]_ , \new_[56666]_ , \new_[56667]_ , \new_[56671]_ ,
    \new_[56672]_ , \new_[56675]_ , \new_[56678]_ , \new_[56679]_ ,
    \new_[56680]_ , \new_[56684]_ , \new_[56685]_ , \new_[56689]_ ,
    \new_[56690]_ , \new_[56691]_ , \new_[56695]_ , \new_[56696]_ ,
    \new_[56699]_ , \new_[56702]_ , \new_[56703]_ , \new_[56704]_ ,
    \new_[56708]_ , \new_[56709]_ , \new_[56713]_ , \new_[56714]_ ,
    \new_[56715]_ , \new_[56719]_ , \new_[56720]_ , \new_[56723]_ ,
    \new_[56726]_ , \new_[56727]_ , \new_[56728]_ , \new_[56732]_ ,
    \new_[56733]_ , \new_[56737]_ , \new_[56738]_ , \new_[56739]_ ,
    \new_[56743]_ , \new_[56744]_ , \new_[56747]_ , \new_[56750]_ ,
    \new_[56751]_ , \new_[56752]_ , \new_[56756]_ , \new_[56757]_ ,
    \new_[56761]_ , \new_[56762]_ , \new_[56763]_ , \new_[56767]_ ,
    \new_[56768]_ , \new_[56771]_ , \new_[56774]_ , \new_[56775]_ ,
    \new_[56776]_ , \new_[56780]_ , \new_[56781]_ , \new_[56785]_ ,
    \new_[56786]_ , \new_[56787]_ , \new_[56791]_ , \new_[56792]_ ,
    \new_[56795]_ , \new_[56798]_ , \new_[56799]_ , \new_[56800]_ ,
    \new_[56804]_ , \new_[56805]_ , \new_[56809]_ , \new_[56810]_ ,
    \new_[56811]_ , \new_[56815]_ , \new_[56816]_ , \new_[56819]_ ,
    \new_[56822]_ , \new_[56823]_ , \new_[56824]_ , \new_[56828]_ ,
    \new_[56829]_ , \new_[56833]_ , \new_[56834]_ , \new_[56835]_ ,
    \new_[56839]_ , \new_[56840]_ , \new_[56843]_ , \new_[56846]_ ,
    \new_[56847]_ , \new_[56848]_ , \new_[56852]_ , \new_[56853]_ ,
    \new_[56857]_ , \new_[56858]_ , \new_[56859]_ , \new_[56863]_ ,
    \new_[56864]_ , \new_[56867]_ , \new_[56870]_ , \new_[56871]_ ,
    \new_[56872]_ , \new_[56876]_ , \new_[56877]_ , \new_[56881]_ ,
    \new_[56882]_ , \new_[56883]_ , \new_[56887]_ , \new_[56888]_ ,
    \new_[56891]_ , \new_[56894]_ , \new_[56895]_ , \new_[56896]_ ,
    \new_[56900]_ , \new_[56901]_ , \new_[56905]_ , \new_[56906]_ ,
    \new_[56907]_ , \new_[56911]_ , \new_[56912]_ , \new_[56915]_ ,
    \new_[56918]_ , \new_[56919]_ , \new_[56920]_ , \new_[56924]_ ,
    \new_[56925]_ , \new_[56929]_ , \new_[56930]_ , \new_[56931]_ ,
    \new_[56935]_ , \new_[56936]_ , \new_[56939]_ , \new_[56942]_ ,
    \new_[56943]_ , \new_[56944]_ , \new_[56948]_ , \new_[56949]_ ,
    \new_[56953]_ , \new_[56954]_ , \new_[56955]_ , \new_[56959]_ ,
    \new_[56960]_ , \new_[56963]_ , \new_[56966]_ , \new_[56967]_ ,
    \new_[56968]_ , \new_[56972]_ , \new_[56973]_ , \new_[56977]_ ,
    \new_[56978]_ , \new_[56979]_ , \new_[56983]_ , \new_[56984]_ ,
    \new_[56987]_ , \new_[56990]_ , \new_[56991]_ , \new_[56992]_ ,
    \new_[56996]_ , \new_[56997]_ , \new_[57001]_ , \new_[57002]_ ,
    \new_[57003]_ , \new_[57007]_ , \new_[57008]_ , \new_[57011]_ ,
    \new_[57014]_ , \new_[57015]_ , \new_[57016]_ , \new_[57020]_ ,
    \new_[57021]_ , \new_[57025]_ , \new_[57026]_ , \new_[57027]_ ,
    \new_[57031]_ , \new_[57032]_ , \new_[57035]_ , \new_[57038]_ ,
    \new_[57039]_ , \new_[57040]_ , \new_[57044]_ , \new_[57045]_ ,
    \new_[57049]_ , \new_[57050]_ , \new_[57051]_ , \new_[57055]_ ,
    \new_[57056]_ , \new_[57059]_ , \new_[57062]_ , \new_[57063]_ ,
    \new_[57064]_ , \new_[57068]_ , \new_[57069]_ , \new_[57073]_ ,
    \new_[57074]_ , \new_[57075]_ , \new_[57079]_ , \new_[57080]_ ,
    \new_[57083]_ , \new_[57086]_ , \new_[57087]_ , \new_[57088]_ ,
    \new_[57092]_ , \new_[57093]_ , \new_[57097]_ , \new_[57098]_ ,
    \new_[57099]_ , \new_[57103]_ , \new_[57104]_ , \new_[57107]_ ,
    \new_[57110]_ , \new_[57111]_ , \new_[57112]_ , \new_[57116]_ ,
    \new_[57117]_ , \new_[57121]_ , \new_[57122]_ , \new_[57123]_ ,
    \new_[57127]_ , \new_[57128]_ , \new_[57131]_ , \new_[57134]_ ,
    \new_[57135]_ , \new_[57136]_ , \new_[57140]_ , \new_[57141]_ ,
    \new_[57145]_ , \new_[57146]_ , \new_[57147]_ , \new_[57151]_ ,
    \new_[57152]_ , \new_[57155]_ , \new_[57158]_ , \new_[57159]_ ,
    \new_[57160]_ , \new_[57164]_ , \new_[57165]_ , \new_[57169]_ ,
    \new_[57170]_ , \new_[57171]_ , \new_[57175]_ , \new_[57176]_ ,
    \new_[57179]_ , \new_[57182]_ , \new_[57183]_ , \new_[57184]_ ,
    \new_[57188]_ , \new_[57189]_ , \new_[57193]_ , \new_[57194]_ ,
    \new_[57195]_ , \new_[57199]_ , \new_[57200]_ , \new_[57203]_ ,
    \new_[57206]_ , \new_[57207]_ , \new_[57208]_ , \new_[57212]_ ,
    \new_[57213]_ , \new_[57217]_ , \new_[57218]_ , \new_[57219]_ ,
    \new_[57223]_ , \new_[57224]_ , \new_[57227]_ , \new_[57230]_ ,
    \new_[57231]_ , \new_[57232]_ , \new_[57236]_ , \new_[57237]_ ,
    \new_[57241]_ , \new_[57242]_ , \new_[57243]_ , \new_[57247]_ ,
    \new_[57248]_ , \new_[57251]_ , \new_[57254]_ , \new_[57255]_ ,
    \new_[57256]_ , \new_[57260]_ , \new_[57261]_ , \new_[57265]_ ,
    \new_[57266]_ , \new_[57267]_ , \new_[57271]_ , \new_[57272]_ ,
    \new_[57275]_ , \new_[57278]_ , \new_[57279]_ , \new_[57280]_ ,
    \new_[57284]_ , \new_[57285]_ , \new_[57289]_ , \new_[57290]_ ,
    \new_[57291]_ , \new_[57295]_ , \new_[57296]_ , \new_[57299]_ ,
    \new_[57302]_ , \new_[57303]_ , \new_[57304]_ , \new_[57308]_ ,
    \new_[57309]_ , \new_[57313]_ , \new_[57314]_ , \new_[57315]_ ,
    \new_[57319]_ , \new_[57320]_ , \new_[57323]_ , \new_[57326]_ ,
    \new_[57327]_ , \new_[57328]_ , \new_[57332]_ , \new_[57333]_ ,
    \new_[57337]_ , \new_[57338]_ , \new_[57339]_ , \new_[57343]_ ,
    \new_[57344]_ , \new_[57347]_ , \new_[57350]_ , \new_[57351]_ ,
    \new_[57352]_ , \new_[57356]_ , \new_[57357]_ , \new_[57361]_ ,
    \new_[57362]_ , \new_[57363]_ , \new_[57367]_ , \new_[57368]_ ,
    \new_[57371]_ , \new_[57374]_ , \new_[57375]_ , \new_[57376]_ ,
    \new_[57380]_ , \new_[57381]_ , \new_[57385]_ , \new_[57386]_ ,
    \new_[57387]_ , \new_[57391]_ , \new_[57392]_ , \new_[57395]_ ,
    \new_[57398]_ , \new_[57399]_ , \new_[57400]_ , \new_[57404]_ ,
    \new_[57405]_ , \new_[57409]_ , \new_[57410]_ , \new_[57411]_ ,
    \new_[57415]_ , \new_[57416]_ , \new_[57419]_ , \new_[57422]_ ,
    \new_[57423]_ , \new_[57424]_ , \new_[57428]_ , \new_[57429]_ ,
    \new_[57433]_ , \new_[57434]_ , \new_[57435]_ , \new_[57439]_ ,
    \new_[57440]_ , \new_[57443]_ , \new_[57446]_ , \new_[57447]_ ,
    \new_[57448]_ , \new_[57452]_ , \new_[57453]_ , \new_[57457]_ ,
    \new_[57458]_ , \new_[57459]_ , \new_[57463]_ , \new_[57464]_ ,
    \new_[57467]_ , \new_[57470]_ , \new_[57471]_ , \new_[57472]_ ,
    \new_[57476]_ , \new_[57477]_ , \new_[57481]_ , \new_[57482]_ ,
    \new_[57483]_ , \new_[57487]_ , \new_[57488]_ , \new_[57491]_ ,
    \new_[57494]_ , \new_[57495]_ , \new_[57496]_ , \new_[57500]_ ,
    \new_[57501]_ , \new_[57505]_ , \new_[57506]_ , \new_[57507]_ ,
    \new_[57511]_ , \new_[57512]_ , \new_[57515]_ , \new_[57518]_ ,
    \new_[57519]_ , \new_[57520]_ , \new_[57524]_ , \new_[57525]_ ,
    \new_[57529]_ , \new_[57530]_ , \new_[57531]_ , \new_[57535]_ ,
    \new_[57536]_ , \new_[57539]_ , \new_[57542]_ , \new_[57543]_ ,
    \new_[57544]_ , \new_[57548]_ , \new_[57549]_ , \new_[57553]_ ,
    \new_[57554]_ , \new_[57555]_ , \new_[57559]_ , \new_[57560]_ ,
    \new_[57563]_ , \new_[57566]_ , \new_[57567]_ , \new_[57568]_ ,
    \new_[57572]_ , \new_[57573]_ , \new_[57577]_ , \new_[57578]_ ,
    \new_[57579]_ , \new_[57583]_ , \new_[57584]_ , \new_[57587]_ ,
    \new_[57590]_ , \new_[57591]_ , \new_[57592]_ , \new_[57596]_ ,
    \new_[57597]_ , \new_[57601]_ , \new_[57602]_ , \new_[57603]_ ,
    \new_[57607]_ , \new_[57608]_ , \new_[57611]_ , \new_[57614]_ ,
    \new_[57615]_ , \new_[57616]_ , \new_[57620]_ , \new_[57621]_ ,
    \new_[57625]_ , \new_[57626]_ , \new_[57627]_ , \new_[57631]_ ,
    \new_[57632]_ , \new_[57635]_ , \new_[57638]_ , \new_[57639]_ ,
    \new_[57640]_ , \new_[57644]_ , \new_[57645]_ , \new_[57649]_ ,
    \new_[57650]_ , \new_[57651]_ , \new_[57655]_ , \new_[57656]_ ,
    \new_[57659]_ , \new_[57662]_ , \new_[57663]_ , \new_[57664]_ ,
    \new_[57668]_ , \new_[57669]_ , \new_[57673]_ , \new_[57674]_ ,
    \new_[57675]_ , \new_[57679]_ , \new_[57680]_ , \new_[57683]_ ,
    \new_[57686]_ , \new_[57687]_ , \new_[57688]_ , \new_[57692]_ ,
    \new_[57693]_ , \new_[57697]_ , \new_[57698]_ , \new_[57699]_ ,
    \new_[57703]_ , \new_[57704]_ , \new_[57707]_ , \new_[57710]_ ,
    \new_[57711]_ , \new_[57712]_ , \new_[57716]_ , \new_[57717]_ ,
    \new_[57721]_ , \new_[57722]_ , \new_[57723]_ , \new_[57727]_ ,
    \new_[57728]_ , \new_[57731]_ , \new_[57734]_ , \new_[57735]_ ,
    \new_[57736]_ , \new_[57740]_ , \new_[57741]_ , \new_[57745]_ ,
    \new_[57746]_ , \new_[57747]_ , \new_[57751]_ , \new_[57752]_ ,
    \new_[57755]_ , \new_[57758]_ , \new_[57759]_ , \new_[57760]_ ,
    \new_[57764]_ , \new_[57765]_ , \new_[57769]_ , \new_[57770]_ ,
    \new_[57771]_ , \new_[57775]_ , \new_[57776]_ , \new_[57779]_ ,
    \new_[57782]_ , \new_[57783]_ , \new_[57784]_ , \new_[57788]_ ,
    \new_[57789]_ , \new_[57793]_ , \new_[57794]_ , \new_[57795]_ ,
    \new_[57799]_ , \new_[57800]_ , \new_[57803]_ , \new_[57806]_ ,
    \new_[57807]_ , \new_[57808]_ , \new_[57812]_ , \new_[57813]_ ,
    \new_[57817]_ , \new_[57818]_ , \new_[57819]_ , \new_[57823]_ ,
    \new_[57824]_ , \new_[57827]_ , \new_[57830]_ , \new_[57831]_ ,
    \new_[57832]_ , \new_[57836]_ , \new_[57837]_ , \new_[57841]_ ,
    \new_[57842]_ , \new_[57843]_ , \new_[57847]_ , \new_[57848]_ ,
    \new_[57851]_ , \new_[57854]_ , \new_[57855]_ , \new_[57856]_ ,
    \new_[57860]_ , \new_[57861]_ , \new_[57865]_ , \new_[57866]_ ,
    \new_[57867]_ , \new_[57871]_ , \new_[57872]_ , \new_[57875]_ ,
    \new_[57878]_ , \new_[57879]_ , \new_[57880]_ , \new_[57884]_ ,
    \new_[57885]_ , \new_[57889]_ , \new_[57890]_ , \new_[57891]_ ,
    \new_[57895]_ , \new_[57896]_ , \new_[57899]_ , \new_[57902]_ ,
    \new_[57903]_ , \new_[57904]_ , \new_[57908]_ , \new_[57909]_ ,
    \new_[57913]_ , \new_[57914]_ , \new_[57915]_ , \new_[57919]_ ,
    \new_[57920]_ , \new_[57923]_ , \new_[57926]_ , \new_[57927]_ ,
    \new_[57928]_ , \new_[57932]_ , \new_[57933]_ , \new_[57937]_ ,
    \new_[57938]_ , \new_[57939]_ , \new_[57943]_ , \new_[57944]_ ,
    \new_[57947]_ , \new_[57950]_ , \new_[57951]_ , \new_[57952]_ ,
    \new_[57956]_ , \new_[57957]_ , \new_[57961]_ , \new_[57962]_ ,
    \new_[57963]_ , \new_[57967]_ , \new_[57968]_ , \new_[57971]_ ,
    \new_[57974]_ , \new_[57975]_ , \new_[57976]_ , \new_[57980]_ ,
    \new_[57981]_ , \new_[57985]_ , \new_[57986]_ , \new_[57987]_ ,
    \new_[57991]_ , \new_[57992]_ , \new_[57995]_ , \new_[57998]_ ,
    \new_[57999]_ , \new_[58000]_ , \new_[58004]_ , \new_[58005]_ ,
    \new_[58009]_ , \new_[58010]_ , \new_[58011]_ , \new_[58015]_ ,
    \new_[58016]_ , \new_[58019]_ , \new_[58022]_ , \new_[58023]_ ,
    \new_[58024]_ , \new_[58028]_ , \new_[58029]_ , \new_[58033]_ ,
    \new_[58034]_ , \new_[58035]_ , \new_[58039]_ , \new_[58040]_ ,
    \new_[58043]_ , \new_[58046]_ , \new_[58047]_ , \new_[58048]_ ,
    \new_[58052]_ , \new_[58053]_ , \new_[58057]_ , \new_[58058]_ ,
    \new_[58059]_ , \new_[58063]_ , \new_[58064]_ , \new_[58067]_ ,
    \new_[58070]_ , \new_[58071]_ , \new_[58072]_ , \new_[58076]_ ,
    \new_[58077]_ , \new_[58081]_ , \new_[58082]_ , \new_[58083]_ ,
    \new_[58087]_ , \new_[58088]_ , \new_[58091]_ , \new_[58094]_ ,
    \new_[58095]_ , \new_[58096]_ , \new_[58100]_ , \new_[58101]_ ,
    \new_[58105]_ , \new_[58106]_ , \new_[58107]_ , \new_[58111]_ ,
    \new_[58112]_ , \new_[58115]_ , \new_[58118]_ , \new_[58119]_ ,
    \new_[58120]_ , \new_[58124]_ , \new_[58125]_ , \new_[58129]_ ,
    \new_[58130]_ , \new_[58131]_ , \new_[58135]_ , \new_[58136]_ ,
    \new_[58139]_ , \new_[58142]_ , \new_[58143]_ , \new_[58144]_ ,
    \new_[58148]_ , \new_[58149]_ , \new_[58153]_ , \new_[58154]_ ,
    \new_[58155]_ , \new_[58159]_ , \new_[58160]_ , \new_[58163]_ ,
    \new_[58166]_ , \new_[58167]_ , \new_[58168]_ , \new_[58172]_ ,
    \new_[58173]_ , \new_[58177]_ , \new_[58178]_ , \new_[58179]_ ,
    \new_[58183]_ , \new_[58184]_ , \new_[58187]_ , \new_[58190]_ ,
    \new_[58191]_ , \new_[58192]_ , \new_[58196]_ , \new_[58197]_ ,
    \new_[58201]_ , \new_[58202]_ , \new_[58203]_ , \new_[58207]_ ,
    \new_[58208]_ , \new_[58211]_ , \new_[58214]_ , \new_[58215]_ ,
    \new_[58216]_ , \new_[58220]_ , \new_[58221]_ , \new_[58225]_ ,
    \new_[58226]_ , \new_[58227]_ , \new_[58231]_ , \new_[58232]_ ,
    \new_[58235]_ , \new_[58238]_ , \new_[58239]_ , \new_[58240]_ ,
    \new_[58244]_ , \new_[58245]_ , \new_[58249]_ , \new_[58250]_ ,
    \new_[58251]_ , \new_[58255]_ , \new_[58256]_ , \new_[58259]_ ,
    \new_[58262]_ , \new_[58263]_ , \new_[58264]_ , \new_[58268]_ ,
    \new_[58269]_ , \new_[58273]_ , \new_[58274]_ , \new_[58275]_ ,
    \new_[58279]_ , \new_[58280]_ , \new_[58283]_ , \new_[58286]_ ,
    \new_[58287]_ , \new_[58288]_ , \new_[58292]_ , \new_[58293]_ ,
    \new_[58297]_ , \new_[58298]_ , \new_[58299]_ , \new_[58303]_ ,
    \new_[58304]_ , \new_[58307]_ , \new_[58310]_ , \new_[58311]_ ,
    \new_[58312]_ , \new_[58316]_ , \new_[58317]_ , \new_[58321]_ ,
    \new_[58322]_ , \new_[58323]_ , \new_[58327]_ , \new_[58328]_ ,
    \new_[58331]_ , \new_[58334]_ , \new_[58335]_ , \new_[58336]_ ,
    \new_[58340]_ , \new_[58341]_ , \new_[58345]_ , \new_[58346]_ ,
    \new_[58347]_ , \new_[58351]_ , \new_[58352]_ , \new_[58355]_ ,
    \new_[58358]_ , \new_[58359]_ , \new_[58360]_ , \new_[58364]_ ,
    \new_[58365]_ , \new_[58369]_ , \new_[58370]_ , \new_[58371]_ ,
    \new_[58375]_ , \new_[58376]_ , \new_[58379]_ , \new_[58382]_ ,
    \new_[58383]_ , \new_[58384]_ , \new_[58388]_ , \new_[58389]_ ,
    \new_[58393]_ , \new_[58394]_ , \new_[58395]_ , \new_[58399]_ ,
    \new_[58400]_ , \new_[58403]_ , \new_[58406]_ , \new_[58407]_ ,
    \new_[58408]_ , \new_[58412]_ , \new_[58413]_ , \new_[58417]_ ,
    \new_[58418]_ , \new_[58419]_ , \new_[58423]_ , \new_[58424]_ ,
    \new_[58427]_ , \new_[58430]_ , \new_[58431]_ , \new_[58432]_ ,
    \new_[58436]_ , \new_[58437]_ , \new_[58441]_ , \new_[58442]_ ,
    \new_[58443]_ , \new_[58447]_ , \new_[58448]_ , \new_[58451]_ ,
    \new_[58454]_ , \new_[58455]_ , \new_[58456]_ , \new_[58460]_ ,
    \new_[58461]_ , \new_[58465]_ , \new_[58466]_ , \new_[58467]_ ,
    \new_[58471]_ , \new_[58472]_ , \new_[58475]_ , \new_[58478]_ ,
    \new_[58479]_ , \new_[58480]_ , \new_[58484]_ , \new_[58485]_ ,
    \new_[58489]_ , \new_[58490]_ , \new_[58491]_ , \new_[58495]_ ,
    \new_[58496]_ , \new_[58499]_ , \new_[58502]_ , \new_[58503]_ ,
    \new_[58504]_ , \new_[58508]_ , \new_[58509]_ , \new_[58513]_ ,
    \new_[58514]_ , \new_[58515]_ , \new_[58519]_ , \new_[58520]_ ,
    \new_[58523]_ , \new_[58526]_ , \new_[58527]_ , \new_[58528]_ ,
    \new_[58532]_ , \new_[58533]_ , \new_[58537]_ , \new_[58538]_ ,
    \new_[58539]_ , \new_[58543]_ , \new_[58544]_ , \new_[58547]_ ,
    \new_[58550]_ , \new_[58551]_ , \new_[58552]_ , \new_[58556]_ ,
    \new_[58557]_ , \new_[58561]_ , \new_[58562]_ , \new_[58563]_ ,
    \new_[58567]_ , \new_[58568]_ , \new_[58571]_ , \new_[58574]_ ,
    \new_[58575]_ , \new_[58576]_ , \new_[58580]_ , \new_[58581]_ ,
    \new_[58585]_ , \new_[58586]_ , \new_[58587]_ , \new_[58591]_ ,
    \new_[58592]_ , \new_[58595]_ , \new_[58598]_ , \new_[58599]_ ,
    \new_[58600]_ , \new_[58604]_ , \new_[58605]_ , \new_[58609]_ ,
    \new_[58610]_ , \new_[58611]_ , \new_[58615]_ , \new_[58616]_ ,
    \new_[58619]_ , \new_[58622]_ , \new_[58623]_ , \new_[58624]_ ,
    \new_[58628]_ , \new_[58629]_ , \new_[58633]_ , \new_[58634]_ ,
    \new_[58635]_ , \new_[58639]_ , \new_[58640]_ , \new_[58643]_ ,
    \new_[58646]_ , \new_[58647]_ , \new_[58648]_ , \new_[58652]_ ,
    \new_[58653]_ , \new_[58657]_ , \new_[58658]_ , \new_[58659]_ ,
    \new_[58663]_ , \new_[58664]_ , \new_[58667]_ , \new_[58670]_ ,
    \new_[58671]_ , \new_[58672]_ , \new_[58676]_ , \new_[58677]_ ,
    \new_[58681]_ , \new_[58682]_ , \new_[58683]_ , \new_[58687]_ ,
    \new_[58688]_ , \new_[58691]_ , \new_[58694]_ , \new_[58695]_ ,
    \new_[58696]_ , \new_[58700]_ , \new_[58701]_ , \new_[58705]_ ,
    \new_[58706]_ , \new_[58707]_ , \new_[58711]_ , \new_[58712]_ ,
    \new_[58715]_ , \new_[58718]_ , \new_[58719]_ , \new_[58720]_ ,
    \new_[58724]_ , \new_[58725]_ , \new_[58729]_ , \new_[58730]_ ,
    \new_[58731]_ , \new_[58735]_ , \new_[58736]_ , \new_[58739]_ ,
    \new_[58742]_ , \new_[58743]_ , \new_[58744]_ , \new_[58748]_ ,
    \new_[58749]_ , \new_[58753]_ , \new_[58754]_ , \new_[58755]_ ,
    \new_[58759]_ , \new_[58760]_ , \new_[58763]_ , \new_[58766]_ ,
    \new_[58767]_ , \new_[58768]_ , \new_[58772]_ , \new_[58773]_ ,
    \new_[58777]_ , \new_[58778]_ , \new_[58779]_ , \new_[58783]_ ,
    \new_[58784]_ , \new_[58787]_ , \new_[58790]_ , \new_[58791]_ ,
    \new_[58792]_ , \new_[58796]_ , \new_[58797]_ , \new_[58801]_ ,
    \new_[58802]_ , \new_[58803]_ , \new_[58807]_ , \new_[58808]_ ,
    \new_[58811]_ , \new_[58814]_ , \new_[58815]_ , \new_[58816]_ ,
    \new_[58820]_ , \new_[58821]_ , \new_[58825]_ , \new_[58826]_ ,
    \new_[58827]_ , \new_[58831]_ , \new_[58832]_ , \new_[58835]_ ,
    \new_[58838]_ , \new_[58839]_ , \new_[58840]_ , \new_[58844]_ ,
    \new_[58845]_ , \new_[58849]_ , \new_[58850]_ , \new_[58851]_ ,
    \new_[58855]_ , \new_[58856]_ , \new_[58859]_ , \new_[58862]_ ,
    \new_[58863]_ , \new_[58864]_ , \new_[58868]_ , \new_[58869]_ ,
    \new_[58873]_ , \new_[58874]_ , \new_[58875]_ , \new_[58879]_ ,
    \new_[58880]_ , \new_[58883]_ , \new_[58886]_ , \new_[58887]_ ,
    \new_[58888]_ , \new_[58892]_ , \new_[58893]_ , \new_[58897]_ ,
    \new_[58898]_ , \new_[58899]_ , \new_[58903]_ , \new_[58904]_ ,
    \new_[58907]_ , \new_[58910]_ , \new_[58911]_ , \new_[58912]_ ,
    \new_[58916]_ , \new_[58917]_ , \new_[58921]_ , \new_[58922]_ ,
    \new_[58923]_ , \new_[58927]_ , \new_[58928]_ , \new_[58931]_ ,
    \new_[58934]_ , \new_[58935]_ , \new_[58936]_ , \new_[58940]_ ,
    \new_[58941]_ , \new_[58945]_ , \new_[58946]_ , \new_[58947]_ ,
    \new_[58951]_ , \new_[58952]_ , \new_[58955]_ , \new_[58958]_ ,
    \new_[58959]_ , \new_[58960]_ , \new_[58964]_ , \new_[58965]_ ,
    \new_[58969]_ , \new_[58970]_ , \new_[58971]_ , \new_[58975]_ ,
    \new_[58976]_ , \new_[58979]_ , \new_[58982]_ , \new_[58983]_ ,
    \new_[58984]_ , \new_[58988]_ , \new_[58989]_ , \new_[58993]_ ,
    \new_[58994]_ , \new_[58995]_ , \new_[58999]_ , \new_[59000]_ ,
    \new_[59003]_ , \new_[59006]_ , \new_[59007]_ , \new_[59008]_ ,
    \new_[59012]_ , \new_[59013]_ , \new_[59017]_ , \new_[59018]_ ,
    \new_[59019]_ , \new_[59023]_ , \new_[59024]_ , \new_[59027]_ ,
    \new_[59030]_ , \new_[59031]_ , \new_[59032]_ , \new_[59036]_ ,
    \new_[59037]_ , \new_[59041]_ , \new_[59042]_ , \new_[59043]_ ,
    \new_[59047]_ , \new_[59048]_ , \new_[59051]_ , \new_[59054]_ ,
    \new_[59055]_ , \new_[59056]_ , \new_[59060]_ , \new_[59061]_ ,
    \new_[59065]_ , \new_[59066]_ , \new_[59067]_ , \new_[59071]_ ,
    \new_[59072]_ , \new_[59075]_ , \new_[59078]_ , \new_[59079]_ ,
    \new_[59080]_ , \new_[59084]_ , \new_[59085]_ , \new_[59089]_ ,
    \new_[59090]_ , \new_[59091]_ , \new_[59095]_ , \new_[59096]_ ,
    \new_[59099]_ , \new_[59102]_ , \new_[59103]_ , \new_[59104]_ ,
    \new_[59108]_ , \new_[59109]_ , \new_[59113]_ , \new_[59114]_ ,
    \new_[59115]_ , \new_[59119]_ , \new_[59120]_ , \new_[59123]_ ,
    \new_[59126]_ , \new_[59127]_ , \new_[59128]_ , \new_[59132]_ ,
    \new_[59133]_ , \new_[59137]_ , \new_[59138]_ , \new_[59139]_ ,
    \new_[59143]_ , \new_[59144]_ , \new_[59147]_ , \new_[59150]_ ,
    \new_[59151]_ , \new_[59152]_ , \new_[59156]_ , \new_[59157]_ ,
    \new_[59161]_ , \new_[59162]_ , \new_[59163]_ , \new_[59167]_ ,
    \new_[59168]_ , \new_[59171]_ , \new_[59174]_ , \new_[59175]_ ,
    \new_[59176]_ , \new_[59180]_ , \new_[59181]_ , \new_[59185]_ ,
    \new_[59186]_ , \new_[59187]_ , \new_[59191]_ , \new_[59192]_ ,
    \new_[59195]_ , \new_[59198]_ , \new_[59199]_ , \new_[59200]_ ,
    \new_[59204]_ , \new_[59205]_ , \new_[59209]_ , \new_[59210]_ ,
    \new_[59211]_ , \new_[59215]_ , \new_[59216]_ , \new_[59219]_ ,
    \new_[59222]_ , \new_[59223]_ , \new_[59224]_ , \new_[59228]_ ,
    \new_[59229]_ , \new_[59233]_ , \new_[59234]_ , \new_[59235]_ ,
    \new_[59239]_ , \new_[59240]_ , \new_[59243]_ , \new_[59246]_ ,
    \new_[59247]_ , \new_[59248]_ , \new_[59252]_ , \new_[59253]_ ,
    \new_[59257]_ , \new_[59258]_ , \new_[59259]_ , \new_[59263]_ ,
    \new_[59264]_ , \new_[59267]_ , \new_[59270]_ , \new_[59271]_ ,
    \new_[59272]_ , \new_[59276]_ , \new_[59277]_ , \new_[59281]_ ,
    \new_[59282]_ , \new_[59283]_ , \new_[59287]_ , \new_[59288]_ ,
    \new_[59291]_ , \new_[59294]_ , \new_[59295]_ , \new_[59296]_ ,
    \new_[59300]_ , \new_[59301]_ , \new_[59305]_ , \new_[59306]_ ,
    \new_[59307]_ , \new_[59311]_ , \new_[59312]_ , \new_[59315]_ ,
    \new_[59318]_ , \new_[59319]_ , \new_[59320]_ , \new_[59324]_ ,
    \new_[59325]_ , \new_[59329]_ , \new_[59330]_ , \new_[59331]_ ,
    \new_[59335]_ , \new_[59336]_ , \new_[59339]_ , \new_[59342]_ ,
    \new_[59343]_ , \new_[59344]_ , \new_[59348]_ , \new_[59349]_ ,
    \new_[59353]_ , \new_[59354]_ , \new_[59355]_ , \new_[59359]_ ,
    \new_[59360]_ , \new_[59363]_ , \new_[59366]_ , \new_[59367]_ ,
    \new_[59368]_ , \new_[59372]_ , \new_[59373]_ , \new_[59377]_ ,
    \new_[59378]_ , \new_[59379]_ , \new_[59383]_ , \new_[59384]_ ,
    \new_[59387]_ , \new_[59390]_ , \new_[59391]_ , \new_[59392]_ ,
    \new_[59396]_ , \new_[59397]_ , \new_[59401]_ , \new_[59402]_ ,
    \new_[59403]_ , \new_[59407]_ , \new_[59408]_ , \new_[59411]_ ,
    \new_[59414]_ , \new_[59415]_ , \new_[59416]_ , \new_[59420]_ ,
    \new_[59421]_ , \new_[59425]_ , \new_[59426]_ , \new_[59427]_ ,
    \new_[59431]_ , \new_[59432]_ , \new_[59435]_ , \new_[59438]_ ,
    \new_[59439]_ , \new_[59440]_ , \new_[59444]_ , \new_[59445]_ ,
    \new_[59449]_ , \new_[59450]_ , \new_[59451]_ , \new_[59455]_ ,
    \new_[59456]_ , \new_[59459]_ , \new_[59462]_ , \new_[59463]_ ,
    \new_[59464]_ , \new_[59468]_ , \new_[59469]_ , \new_[59473]_ ,
    \new_[59474]_ , \new_[59475]_ , \new_[59479]_ , \new_[59480]_ ,
    \new_[59483]_ , \new_[59486]_ , \new_[59487]_ , \new_[59488]_ ,
    \new_[59492]_ , \new_[59493]_ , \new_[59497]_ , \new_[59498]_ ,
    \new_[59499]_ , \new_[59503]_ , \new_[59504]_ , \new_[59507]_ ,
    \new_[59510]_ , \new_[59511]_ , \new_[59512]_ , \new_[59516]_ ,
    \new_[59517]_ , \new_[59521]_ , \new_[59522]_ , \new_[59523]_ ,
    \new_[59527]_ , \new_[59528]_ , \new_[59531]_ , \new_[59534]_ ,
    \new_[59535]_ , \new_[59536]_ , \new_[59540]_ , \new_[59541]_ ,
    \new_[59545]_ , \new_[59546]_ , \new_[59547]_ , \new_[59551]_ ,
    \new_[59552]_ , \new_[59555]_ , \new_[59558]_ , \new_[59559]_ ,
    \new_[59560]_ , \new_[59564]_ , \new_[59565]_ , \new_[59569]_ ,
    \new_[59570]_ , \new_[59571]_ , \new_[59575]_ , \new_[59576]_ ,
    \new_[59579]_ , \new_[59582]_ , \new_[59583]_ , \new_[59584]_ ,
    \new_[59588]_ , \new_[59589]_ , \new_[59593]_ , \new_[59594]_ ,
    \new_[59595]_ , \new_[59599]_ , \new_[59600]_ , \new_[59603]_ ,
    \new_[59606]_ , \new_[59607]_ , \new_[59608]_ , \new_[59612]_ ,
    \new_[59613]_ , \new_[59617]_ , \new_[59618]_ , \new_[59619]_ ,
    \new_[59623]_ , \new_[59624]_ , \new_[59627]_ , \new_[59630]_ ,
    \new_[59631]_ , \new_[59632]_ , \new_[59636]_ , \new_[59637]_ ,
    \new_[59641]_ , \new_[59642]_ , \new_[59643]_ , \new_[59647]_ ,
    \new_[59648]_ , \new_[59651]_ , \new_[59654]_ , \new_[59655]_ ,
    \new_[59656]_ , \new_[59660]_ , \new_[59661]_ , \new_[59665]_ ,
    \new_[59666]_ , \new_[59667]_ , \new_[59671]_ , \new_[59672]_ ,
    \new_[59675]_ , \new_[59678]_ , \new_[59679]_ , \new_[59680]_ ,
    \new_[59684]_ , \new_[59685]_ , \new_[59689]_ , \new_[59690]_ ,
    \new_[59691]_ , \new_[59695]_ , \new_[59696]_ , \new_[59699]_ ,
    \new_[59702]_ , \new_[59703]_ , \new_[59704]_ , \new_[59708]_ ,
    \new_[59709]_ , \new_[59713]_ , \new_[59714]_ , \new_[59715]_ ,
    \new_[59719]_ , \new_[59720]_ , \new_[59723]_ , \new_[59726]_ ,
    \new_[59727]_ , \new_[59728]_ , \new_[59732]_ , \new_[59733]_ ,
    \new_[59737]_ , \new_[59738]_ , \new_[59739]_ , \new_[59743]_ ,
    \new_[59744]_ , \new_[59747]_ , \new_[59750]_ , \new_[59751]_ ,
    \new_[59752]_ , \new_[59756]_ , \new_[59757]_ , \new_[59761]_ ,
    \new_[59762]_ , \new_[59763]_ , \new_[59767]_ , \new_[59768]_ ,
    \new_[59771]_ , \new_[59774]_ , \new_[59775]_ , \new_[59776]_ ,
    \new_[59780]_ , \new_[59781]_ , \new_[59785]_ , \new_[59786]_ ,
    \new_[59787]_ , \new_[59791]_ , \new_[59792]_ , \new_[59795]_ ,
    \new_[59798]_ , \new_[59799]_ , \new_[59800]_ , \new_[59804]_ ,
    \new_[59805]_ , \new_[59809]_ , \new_[59810]_ , \new_[59811]_ ,
    \new_[59815]_ , \new_[59816]_ , \new_[59819]_ , \new_[59822]_ ,
    \new_[59823]_ , \new_[59824]_ , \new_[59828]_ , \new_[59829]_ ,
    \new_[59833]_ , \new_[59834]_ , \new_[59835]_ , \new_[59839]_ ,
    \new_[59840]_ , \new_[59843]_ , \new_[59846]_ , \new_[59847]_ ,
    \new_[59848]_ , \new_[59852]_ , \new_[59853]_ , \new_[59857]_ ,
    \new_[59858]_ , \new_[59859]_ , \new_[59863]_ , \new_[59864]_ ,
    \new_[59867]_ , \new_[59870]_ , \new_[59871]_ , \new_[59872]_ ,
    \new_[59876]_ , \new_[59877]_ , \new_[59881]_ , \new_[59882]_ ,
    \new_[59883]_ , \new_[59887]_ , \new_[59888]_ , \new_[59891]_ ,
    \new_[59894]_ , \new_[59895]_ , \new_[59896]_ , \new_[59900]_ ,
    \new_[59901]_ , \new_[59905]_ , \new_[59906]_ , \new_[59907]_ ,
    \new_[59911]_ , \new_[59912]_ , \new_[59915]_ , \new_[59918]_ ,
    \new_[59919]_ , \new_[59920]_ , \new_[59924]_ , \new_[59925]_ ,
    \new_[59929]_ , \new_[59930]_ , \new_[59931]_ , \new_[59935]_ ,
    \new_[59936]_ , \new_[59939]_ , \new_[59942]_ , \new_[59943]_ ,
    \new_[59944]_ , \new_[59948]_ , \new_[59949]_ , \new_[59953]_ ,
    \new_[59954]_ , \new_[59955]_ , \new_[59959]_ , \new_[59960]_ ,
    \new_[59963]_ , \new_[59966]_ , \new_[59967]_ , \new_[59968]_ ,
    \new_[59972]_ , \new_[59973]_ , \new_[59977]_ , \new_[59978]_ ,
    \new_[59979]_ , \new_[59983]_ , \new_[59984]_ , \new_[59987]_ ,
    \new_[59990]_ , \new_[59991]_ , \new_[59992]_ , \new_[59996]_ ,
    \new_[59997]_ , \new_[60001]_ , \new_[60002]_ , \new_[60003]_ ,
    \new_[60007]_ , \new_[60008]_ , \new_[60011]_ , \new_[60014]_ ,
    \new_[60015]_ , \new_[60016]_ , \new_[60020]_ , \new_[60021]_ ,
    \new_[60025]_ , \new_[60026]_ , \new_[60027]_ , \new_[60031]_ ,
    \new_[60032]_ , \new_[60035]_ , \new_[60038]_ , \new_[60039]_ ,
    \new_[60040]_ , \new_[60044]_ , \new_[60045]_ , \new_[60049]_ ,
    \new_[60050]_ , \new_[60051]_ , \new_[60055]_ , \new_[60056]_ ,
    \new_[60059]_ , \new_[60062]_ , \new_[60063]_ , \new_[60064]_ ,
    \new_[60068]_ , \new_[60069]_ , \new_[60073]_ , \new_[60074]_ ,
    \new_[60075]_ , \new_[60079]_ , \new_[60080]_ , \new_[60083]_ ,
    \new_[60086]_ , \new_[60087]_ , \new_[60088]_ , \new_[60092]_ ,
    \new_[60093]_ , \new_[60097]_ , \new_[60098]_ , \new_[60099]_ ,
    \new_[60103]_ , \new_[60104]_ , \new_[60107]_ , \new_[60110]_ ,
    \new_[60111]_ , \new_[60112]_ , \new_[60116]_ , \new_[60117]_ ,
    \new_[60120]_ , \new_[60123]_ , \new_[60124]_ , \new_[60125]_ ,
    \new_[60129]_ , \new_[60130]_ , \new_[60133]_ , \new_[60136]_ ,
    \new_[60137]_ , \new_[60138]_ , \new_[60142]_ , \new_[60143]_ ,
    \new_[60146]_ , \new_[60149]_ , \new_[60150]_ , \new_[60151]_ ,
    \new_[60155]_ , \new_[60156]_ , \new_[60159]_ , \new_[60162]_ ,
    \new_[60163]_ , \new_[60164]_ , \new_[60168]_ , \new_[60169]_ ,
    \new_[60172]_ , \new_[60175]_ , \new_[60176]_ , \new_[60177]_ ,
    \new_[60181]_ , \new_[60182]_ , \new_[60185]_ , \new_[60188]_ ,
    \new_[60189]_ , \new_[60190]_ , \new_[60194]_ , \new_[60195]_ ,
    \new_[60198]_ , \new_[60201]_ , \new_[60202]_ , \new_[60203]_ ,
    \new_[60207]_ , \new_[60208]_ , \new_[60211]_ , \new_[60214]_ ,
    \new_[60215]_ , \new_[60216]_ , \new_[60220]_ , \new_[60221]_ ,
    \new_[60224]_ , \new_[60227]_ , \new_[60228]_ , \new_[60229]_ ,
    \new_[60233]_ , \new_[60234]_ , \new_[60237]_ , \new_[60240]_ ,
    \new_[60241]_ , \new_[60242]_ , \new_[60246]_ , \new_[60247]_ ,
    \new_[60250]_ , \new_[60253]_ , \new_[60254]_ , \new_[60255]_ ,
    \new_[60259]_ , \new_[60260]_ , \new_[60263]_ , \new_[60266]_ ,
    \new_[60267]_ , \new_[60268]_ , \new_[60272]_ , \new_[60273]_ ,
    \new_[60276]_ , \new_[60279]_ , \new_[60280]_ , \new_[60281]_ ,
    \new_[60285]_ , \new_[60286]_ , \new_[60289]_ , \new_[60292]_ ,
    \new_[60293]_ , \new_[60294]_ , \new_[60298]_ , \new_[60299]_ ,
    \new_[60302]_ , \new_[60305]_ , \new_[60306]_ , \new_[60307]_ ,
    \new_[60311]_ , \new_[60312]_ , \new_[60315]_ , \new_[60318]_ ,
    \new_[60319]_ , \new_[60320]_ , \new_[60324]_ , \new_[60325]_ ,
    \new_[60328]_ , \new_[60331]_ , \new_[60332]_ , \new_[60333]_ ,
    \new_[60337]_ , \new_[60338]_ , \new_[60341]_ , \new_[60344]_ ,
    \new_[60345]_ , \new_[60346]_ , \new_[60350]_ , \new_[60351]_ ,
    \new_[60354]_ , \new_[60357]_ , \new_[60358]_ , \new_[60359]_ ,
    \new_[60363]_ , \new_[60364]_ , \new_[60367]_ , \new_[60370]_ ,
    \new_[60371]_ , \new_[60372]_ , \new_[60376]_ , \new_[60377]_ ,
    \new_[60380]_ , \new_[60383]_ , \new_[60384]_ , \new_[60385]_ ,
    \new_[60389]_ , \new_[60390]_ , \new_[60393]_ , \new_[60396]_ ,
    \new_[60397]_ , \new_[60398]_ , \new_[60402]_ , \new_[60403]_ ,
    \new_[60406]_ , \new_[60409]_ , \new_[60410]_ , \new_[60411]_ ,
    \new_[60415]_ , \new_[60416]_ , \new_[60419]_ , \new_[60422]_ ,
    \new_[60423]_ , \new_[60424]_ , \new_[60428]_ , \new_[60429]_ ,
    \new_[60432]_ , \new_[60435]_ , \new_[60436]_ , \new_[60437]_ ,
    \new_[60441]_ , \new_[60442]_ , \new_[60445]_ , \new_[60448]_ ,
    \new_[60449]_ , \new_[60450]_ , \new_[60454]_ , \new_[60455]_ ,
    \new_[60458]_ , \new_[60461]_ , \new_[60462]_ , \new_[60463]_ ,
    \new_[60467]_ , \new_[60468]_ , \new_[60471]_ , \new_[60474]_ ,
    \new_[60475]_ , \new_[60476]_ , \new_[60480]_ , \new_[60481]_ ,
    \new_[60484]_ , \new_[60487]_ , \new_[60488]_ , \new_[60489]_ ,
    \new_[60493]_ , \new_[60494]_ , \new_[60497]_ , \new_[60500]_ ,
    \new_[60501]_ , \new_[60502]_ , \new_[60506]_ , \new_[60507]_ ,
    \new_[60510]_ , \new_[60513]_ , \new_[60514]_ , \new_[60515]_ ,
    \new_[60519]_ , \new_[60520]_ , \new_[60523]_ , \new_[60526]_ ,
    \new_[60527]_ , \new_[60528]_ , \new_[60532]_ , \new_[60533]_ ,
    \new_[60536]_ , \new_[60539]_ , \new_[60540]_ , \new_[60541]_ ,
    \new_[60545]_ , \new_[60546]_ , \new_[60549]_ , \new_[60552]_ ,
    \new_[60553]_ , \new_[60554]_ , \new_[60558]_ , \new_[60559]_ ,
    \new_[60562]_ , \new_[60565]_ , \new_[60566]_ , \new_[60567]_ ,
    \new_[60571]_ , \new_[60572]_ , \new_[60575]_ , \new_[60578]_ ,
    \new_[60579]_ , \new_[60580]_ , \new_[60584]_ , \new_[60585]_ ,
    \new_[60588]_ , \new_[60591]_ , \new_[60592]_ , \new_[60593]_ ,
    \new_[60597]_ , \new_[60598]_ , \new_[60601]_ , \new_[60604]_ ,
    \new_[60605]_ , \new_[60606]_ , \new_[60610]_ , \new_[60611]_ ,
    \new_[60614]_ , \new_[60617]_ , \new_[60618]_ , \new_[60619]_ ,
    \new_[60623]_ , \new_[60624]_ , \new_[60627]_ , \new_[60630]_ ,
    \new_[60631]_ , \new_[60632]_ , \new_[60636]_ , \new_[60637]_ ,
    \new_[60640]_ , \new_[60643]_ , \new_[60644]_ , \new_[60645]_ ,
    \new_[60649]_ , \new_[60650]_ , \new_[60653]_ , \new_[60656]_ ,
    \new_[60657]_ , \new_[60658]_ , \new_[60662]_ , \new_[60663]_ ,
    \new_[60666]_ , \new_[60669]_ , \new_[60670]_ , \new_[60671]_ ,
    \new_[60675]_ , \new_[60676]_ , \new_[60679]_ , \new_[60682]_ ,
    \new_[60683]_ , \new_[60684]_ , \new_[60688]_ , \new_[60689]_ ,
    \new_[60692]_ , \new_[60695]_ , \new_[60696]_ , \new_[60697]_ ,
    \new_[60701]_ , \new_[60702]_ , \new_[60705]_ , \new_[60708]_ ,
    \new_[60709]_ , \new_[60710]_ , \new_[60714]_ , \new_[60715]_ ,
    \new_[60718]_ , \new_[60721]_ , \new_[60722]_ , \new_[60723]_ ,
    \new_[60727]_ , \new_[60728]_ , \new_[60731]_ , \new_[60734]_ ,
    \new_[60735]_ , \new_[60736]_ , \new_[60740]_ , \new_[60741]_ ,
    \new_[60744]_ , \new_[60747]_ , \new_[60748]_ , \new_[60749]_ ,
    \new_[60753]_ , \new_[60754]_ , \new_[60757]_ , \new_[60760]_ ,
    \new_[60761]_ , \new_[60762]_ , \new_[60766]_ , \new_[60767]_ ,
    \new_[60770]_ , \new_[60773]_ , \new_[60774]_ , \new_[60775]_ ,
    \new_[60779]_ , \new_[60780]_ , \new_[60783]_ , \new_[60786]_ ,
    \new_[60787]_ , \new_[60788]_ , \new_[60792]_ , \new_[60793]_ ,
    \new_[60796]_ , \new_[60799]_ , \new_[60800]_ , \new_[60801]_ ,
    \new_[60805]_ , \new_[60806]_ , \new_[60809]_ , \new_[60812]_ ,
    \new_[60813]_ , \new_[60814]_ , \new_[60818]_ , \new_[60819]_ ,
    \new_[60822]_ , \new_[60825]_ , \new_[60826]_ , \new_[60827]_ ,
    \new_[60831]_ , \new_[60832]_ , \new_[60835]_ , \new_[60838]_ ,
    \new_[60839]_ , \new_[60840]_ , \new_[60844]_ , \new_[60845]_ ,
    \new_[60848]_ , \new_[60851]_ , \new_[60852]_ , \new_[60853]_ ,
    \new_[60857]_ , \new_[60858]_ , \new_[60861]_ , \new_[60864]_ ,
    \new_[60865]_ , \new_[60866]_ , \new_[60870]_ , \new_[60871]_ ,
    \new_[60874]_ , \new_[60877]_ , \new_[60878]_ , \new_[60879]_ ,
    \new_[60883]_ , \new_[60884]_ , \new_[60887]_ , \new_[60890]_ ,
    \new_[60891]_ , \new_[60892]_ , \new_[60896]_ , \new_[60897]_ ,
    \new_[60900]_ , \new_[60903]_ , \new_[60904]_ , \new_[60905]_ ,
    \new_[60909]_ , \new_[60910]_ , \new_[60913]_ , \new_[60916]_ ,
    \new_[60917]_ , \new_[60918]_ , \new_[60922]_ , \new_[60923]_ ,
    \new_[60926]_ , \new_[60929]_ , \new_[60930]_ , \new_[60931]_ ,
    \new_[60935]_ , \new_[60936]_ , \new_[60939]_ , \new_[60942]_ ,
    \new_[60943]_ , \new_[60944]_ , \new_[60948]_ , \new_[60949]_ ,
    \new_[60952]_ , \new_[60955]_ , \new_[60956]_ , \new_[60957]_ ,
    \new_[60961]_ , \new_[60962]_ , \new_[60965]_ , \new_[60968]_ ,
    \new_[60969]_ , \new_[60970]_ , \new_[60974]_ , \new_[60975]_ ,
    \new_[60978]_ , \new_[60981]_ , \new_[60982]_ , \new_[60983]_ ,
    \new_[60987]_ , \new_[60988]_ , \new_[60991]_ , \new_[60994]_ ,
    \new_[60995]_ , \new_[60996]_ , \new_[61000]_ , \new_[61001]_ ,
    \new_[61004]_ , \new_[61007]_ , \new_[61008]_ , \new_[61009]_ ,
    \new_[61013]_ , \new_[61014]_ , \new_[61017]_ , \new_[61020]_ ,
    \new_[61021]_ , \new_[61022]_ , \new_[61026]_ , \new_[61027]_ ,
    \new_[61030]_ , \new_[61033]_ , \new_[61034]_ , \new_[61035]_ ,
    \new_[61039]_ , \new_[61040]_ , \new_[61043]_ , \new_[61046]_ ,
    \new_[61047]_ , \new_[61048]_ , \new_[61052]_ , \new_[61053]_ ,
    \new_[61056]_ , \new_[61059]_ , \new_[61060]_ , \new_[61061]_ ,
    \new_[61065]_ , \new_[61066]_ , \new_[61069]_ , \new_[61072]_ ,
    \new_[61073]_ , \new_[61074]_ , \new_[61078]_ , \new_[61079]_ ,
    \new_[61082]_ , \new_[61085]_ , \new_[61086]_ , \new_[61087]_ ,
    \new_[61091]_ , \new_[61092]_ , \new_[61095]_ , \new_[61098]_ ,
    \new_[61099]_ , \new_[61100]_ , \new_[61104]_ , \new_[61105]_ ,
    \new_[61108]_ , \new_[61111]_ , \new_[61112]_ , \new_[61113]_ ,
    \new_[61117]_ , \new_[61118]_ , \new_[61121]_ , \new_[61124]_ ,
    \new_[61125]_ , \new_[61126]_ , \new_[61130]_ , \new_[61131]_ ,
    \new_[61134]_ , \new_[61137]_ , \new_[61138]_ , \new_[61139]_ ,
    \new_[61143]_ , \new_[61144]_ , \new_[61147]_ , \new_[61150]_ ,
    \new_[61151]_ , \new_[61152]_ , \new_[61156]_ , \new_[61157]_ ,
    \new_[61160]_ , \new_[61163]_ , \new_[61164]_ , \new_[61165]_ ,
    \new_[61169]_ , \new_[61170]_ , \new_[61173]_ , \new_[61176]_ ,
    \new_[61177]_ , \new_[61178]_ , \new_[61182]_ , \new_[61183]_ ,
    \new_[61186]_ , \new_[61189]_ , \new_[61190]_ , \new_[61191]_ ,
    \new_[61195]_ , \new_[61196]_ , \new_[61199]_ , \new_[61202]_ ,
    \new_[61203]_ , \new_[61204]_ , \new_[61208]_ , \new_[61209]_ ,
    \new_[61212]_ , \new_[61215]_ , \new_[61216]_ , \new_[61217]_ ,
    \new_[61221]_ , \new_[61222]_ , \new_[61225]_ , \new_[61228]_ ,
    \new_[61229]_ , \new_[61230]_ , \new_[61234]_ , \new_[61235]_ ,
    \new_[61238]_ , \new_[61241]_ , \new_[61242]_ , \new_[61243]_ ,
    \new_[61247]_ , \new_[61248]_ , \new_[61251]_ , \new_[61254]_ ,
    \new_[61255]_ , \new_[61256]_ , \new_[61260]_ , \new_[61261]_ ,
    \new_[61264]_ , \new_[61267]_ , \new_[61268]_ , \new_[61269]_ ,
    \new_[61273]_ , \new_[61274]_ , \new_[61277]_ , \new_[61280]_ ,
    \new_[61281]_ , \new_[61282]_ , \new_[61286]_ , \new_[61287]_ ,
    \new_[61290]_ , \new_[61293]_ , \new_[61294]_ , \new_[61295]_ ,
    \new_[61299]_ , \new_[61300]_ , \new_[61303]_ , \new_[61306]_ ,
    \new_[61307]_ , \new_[61308]_ , \new_[61312]_ , \new_[61313]_ ,
    \new_[61316]_ , \new_[61319]_ , \new_[61320]_ , \new_[61321]_ ,
    \new_[61325]_ , \new_[61326]_ , \new_[61329]_ , \new_[61332]_ ,
    \new_[61333]_ , \new_[61334]_ , \new_[61338]_ , \new_[61339]_ ,
    \new_[61342]_ , \new_[61345]_ , \new_[61346]_ , \new_[61347]_ ,
    \new_[61351]_ , \new_[61352]_ , \new_[61355]_ , \new_[61358]_ ,
    \new_[61359]_ , \new_[61360]_ , \new_[61364]_ , \new_[61365]_ ,
    \new_[61368]_ , \new_[61371]_ , \new_[61372]_ , \new_[61373]_ ,
    \new_[61377]_ , \new_[61378]_ , \new_[61381]_ , \new_[61384]_ ,
    \new_[61385]_ , \new_[61386]_ , \new_[61390]_ , \new_[61391]_ ,
    \new_[61394]_ , \new_[61397]_ , \new_[61398]_ , \new_[61399]_ ,
    \new_[61403]_ , \new_[61404]_ , \new_[61407]_ , \new_[61410]_ ,
    \new_[61411]_ , \new_[61412]_ , \new_[61416]_ , \new_[61417]_ ,
    \new_[61420]_ , \new_[61423]_ , \new_[61424]_ , \new_[61425]_ ,
    \new_[61429]_ , \new_[61430]_ , \new_[61433]_ , \new_[61436]_ ,
    \new_[61437]_ , \new_[61438]_ , \new_[61442]_ , \new_[61443]_ ,
    \new_[61446]_ , \new_[61449]_ , \new_[61450]_ , \new_[61451]_ ,
    \new_[61455]_ , \new_[61456]_ , \new_[61459]_ , \new_[61462]_ ,
    \new_[61463]_ , \new_[61464]_ , \new_[61468]_ , \new_[61469]_ ,
    \new_[61472]_ , \new_[61475]_ , \new_[61476]_ , \new_[61477]_ ,
    \new_[61481]_ , \new_[61482]_ , \new_[61485]_ , \new_[61488]_ ,
    \new_[61489]_ , \new_[61490]_ , \new_[61494]_ , \new_[61495]_ ,
    \new_[61498]_ , \new_[61501]_ , \new_[61502]_ , \new_[61503]_ ,
    \new_[61507]_ , \new_[61508]_ , \new_[61511]_ , \new_[61514]_ ,
    \new_[61515]_ , \new_[61516]_ , \new_[61520]_ , \new_[61521]_ ,
    \new_[61524]_ , \new_[61527]_ , \new_[61528]_ , \new_[61529]_ ,
    \new_[61533]_ , \new_[61534]_ , \new_[61537]_ , \new_[61540]_ ,
    \new_[61541]_ , \new_[61542]_ , \new_[61546]_ , \new_[61547]_ ,
    \new_[61550]_ , \new_[61553]_ , \new_[61554]_ , \new_[61555]_ ,
    \new_[61559]_ , \new_[61560]_ , \new_[61563]_ , \new_[61566]_ ,
    \new_[61567]_ , \new_[61568]_ , \new_[61572]_ , \new_[61573]_ ,
    \new_[61576]_ , \new_[61579]_ , \new_[61580]_ , \new_[61581]_ ,
    \new_[61585]_ , \new_[61586]_ , \new_[61589]_ , \new_[61592]_ ,
    \new_[61593]_ , \new_[61594]_ , \new_[61598]_ , \new_[61599]_ ,
    \new_[61602]_ , \new_[61605]_ , \new_[61606]_ , \new_[61607]_ ,
    \new_[61611]_ , \new_[61612]_ , \new_[61615]_ , \new_[61618]_ ,
    \new_[61619]_ , \new_[61620]_ , \new_[61624]_ , \new_[61625]_ ,
    \new_[61628]_ , \new_[61631]_ , \new_[61632]_ , \new_[61633]_ ,
    \new_[61637]_ , \new_[61638]_ , \new_[61641]_ , \new_[61644]_ ,
    \new_[61645]_ , \new_[61646]_ , \new_[61650]_ , \new_[61651]_ ,
    \new_[61654]_ , \new_[61657]_ , \new_[61658]_ , \new_[61659]_ ,
    \new_[61663]_ , \new_[61664]_ , \new_[61667]_ , \new_[61670]_ ,
    \new_[61671]_ , \new_[61672]_ , \new_[61676]_ , \new_[61677]_ ,
    \new_[61680]_ , \new_[61683]_ , \new_[61684]_ , \new_[61685]_ ,
    \new_[61689]_ , \new_[61690]_ , \new_[61693]_ , \new_[61696]_ ,
    \new_[61697]_ , \new_[61698]_ , \new_[61702]_ , \new_[61703]_ ,
    \new_[61706]_ , \new_[61709]_ , \new_[61710]_ , \new_[61711]_ ,
    \new_[61715]_ , \new_[61716]_ , \new_[61719]_ , \new_[61722]_ ,
    \new_[61723]_ , \new_[61724]_ , \new_[61728]_ , \new_[61729]_ ,
    \new_[61732]_ , \new_[61735]_ , \new_[61736]_ , \new_[61737]_ ,
    \new_[61741]_ , \new_[61742]_ , \new_[61745]_ , \new_[61748]_ ,
    \new_[61749]_ , \new_[61750]_ , \new_[61754]_ , \new_[61755]_ ,
    \new_[61758]_ , \new_[61761]_ , \new_[61762]_ , \new_[61763]_ ,
    \new_[61767]_ , \new_[61768]_ , \new_[61771]_ , \new_[61774]_ ,
    \new_[61775]_ , \new_[61776]_ , \new_[61780]_ , \new_[61781]_ ,
    \new_[61784]_ , \new_[61787]_ , \new_[61788]_ , \new_[61789]_ ,
    \new_[61793]_ , \new_[61794]_ , \new_[61797]_ , \new_[61800]_ ,
    \new_[61801]_ , \new_[61802]_ , \new_[61806]_ , \new_[61807]_ ,
    \new_[61810]_ , \new_[61813]_ , \new_[61814]_ , \new_[61815]_ ,
    \new_[61819]_ , \new_[61820]_ , \new_[61823]_ , \new_[61826]_ ,
    \new_[61827]_ , \new_[61828]_ , \new_[61832]_ , \new_[61833]_ ,
    \new_[61836]_ , \new_[61839]_ , \new_[61840]_ , \new_[61841]_ ,
    \new_[61845]_ , \new_[61846]_ , \new_[61849]_ , \new_[61852]_ ,
    \new_[61853]_ , \new_[61854]_ , \new_[61858]_ , \new_[61859]_ ,
    \new_[61862]_ , \new_[61865]_ , \new_[61866]_ , \new_[61867]_ ,
    \new_[61871]_ , \new_[61872]_ , \new_[61875]_ , \new_[61878]_ ,
    \new_[61879]_ , \new_[61880]_ , \new_[61884]_ , \new_[61885]_ ,
    \new_[61888]_ , \new_[61891]_ , \new_[61892]_ , \new_[61893]_ ,
    \new_[61897]_ , \new_[61898]_ , \new_[61901]_ , \new_[61904]_ ,
    \new_[61905]_ , \new_[61906]_ , \new_[61910]_ , \new_[61911]_ ,
    \new_[61914]_ , \new_[61917]_ , \new_[61918]_ , \new_[61919]_ ,
    \new_[61923]_ , \new_[61924]_ , \new_[61927]_ , \new_[61930]_ ,
    \new_[61931]_ , \new_[61932]_ , \new_[61936]_ , \new_[61937]_ ,
    \new_[61940]_ , \new_[61943]_ , \new_[61944]_ , \new_[61945]_ ,
    \new_[61949]_ , \new_[61950]_ , \new_[61953]_ , \new_[61956]_ ,
    \new_[61957]_ , \new_[61958]_ , \new_[61962]_ , \new_[61963]_ ,
    \new_[61966]_ , \new_[61969]_ , \new_[61970]_ , \new_[61971]_ ,
    \new_[61975]_ , \new_[61976]_ , \new_[61979]_ , \new_[61982]_ ,
    \new_[61983]_ , \new_[61984]_ , \new_[61988]_ , \new_[61989]_ ,
    \new_[61992]_ , \new_[61995]_ , \new_[61996]_ , \new_[61997]_ ,
    \new_[62001]_ , \new_[62002]_ , \new_[62005]_ , \new_[62008]_ ,
    \new_[62009]_ , \new_[62010]_ , \new_[62014]_ , \new_[62015]_ ,
    \new_[62018]_ , \new_[62021]_ , \new_[62022]_ , \new_[62023]_ ,
    \new_[62027]_ , \new_[62028]_ , \new_[62031]_ , \new_[62034]_ ,
    \new_[62035]_ , \new_[62036]_ , \new_[62040]_ , \new_[62041]_ ,
    \new_[62044]_ , \new_[62047]_ , \new_[62048]_ , \new_[62049]_ ,
    \new_[62053]_ , \new_[62054]_ , \new_[62057]_ , \new_[62060]_ ,
    \new_[62061]_ , \new_[62062]_ , \new_[62066]_ , \new_[62067]_ ,
    \new_[62070]_ , \new_[62073]_ , \new_[62074]_ , \new_[62075]_ ,
    \new_[62079]_ , \new_[62080]_ , \new_[62083]_ , \new_[62086]_ ,
    \new_[62087]_ , \new_[62088]_ , \new_[62092]_ , \new_[62093]_ ,
    \new_[62096]_ , \new_[62099]_ , \new_[62100]_ , \new_[62101]_ ,
    \new_[62105]_ , \new_[62106]_ , \new_[62109]_ , \new_[62112]_ ,
    \new_[62113]_ , \new_[62114]_ , \new_[62118]_ , \new_[62119]_ ,
    \new_[62122]_ , \new_[62125]_ , \new_[62126]_ , \new_[62127]_ ,
    \new_[62131]_ , \new_[62132]_ , \new_[62135]_ , \new_[62138]_ ,
    \new_[62139]_ , \new_[62140]_ , \new_[62144]_ , \new_[62145]_ ,
    \new_[62148]_ , \new_[62151]_ , \new_[62152]_ , \new_[62153]_ ,
    \new_[62157]_ , \new_[62158]_ , \new_[62161]_ , \new_[62164]_ ,
    \new_[62165]_ , \new_[62166]_ , \new_[62170]_ , \new_[62171]_ ,
    \new_[62174]_ , \new_[62177]_ , \new_[62178]_ , \new_[62179]_ ,
    \new_[62183]_ , \new_[62184]_ , \new_[62187]_ , \new_[62190]_ ,
    \new_[62191]_ , \new_[62192]_ , \new_[62196]_ , \new_[62197]_ ,
    \new_[62200]_ , \new_[62203]_ , \new_[62204]_ , \new_[62205]_ ,
    \new_[62209]_ , \new_[62210]_ , \new_[62213]_ , \new_[62216]_ ,
    \new_[62217]_ , \new_[62218]_ , \new_[62222]_ , \new_[62223]_ ,
    \new_[62226]_ , \new_[62229]_ , \new_[62230]_ , \new_[62231]_ ,
    \new_[62235]_ , \new_[62236]_ , \new_[62239]_ , \new_[62242]_ ,
    \new_[62243]_ , \new_[62244]_ , \new_[62248]_ , \new_[62249]_ ,
    \new_[62252]_ , \new_[62255]_ , \new_[62256]_ , \new_[62257]_ ,
    \new_[62261]_ , \new_[62262]_ , \new_[62265]_ , \new_[62268]_ ,
    \new_[62269]_ , \new_[62270]_ , \new_[62274]_ , \new_[62275]_ ,
    \new_[62278]_ , \new_[62281]_ , \new_[62282]_ , \new_[62283]_ ,
    \new_[62287]_ , \new_[62288]_ , \new_[62291]_ , \new_[62294]_ ,
    \new_[62295]_ , \new_[62296]_ , \new_[62300]_ , \new_[62301]_ ,
    \new_[62304]_ , \new_[62307]_ , \new_[62308]_ , \new_[62309]_ ,
    \new_[62313]_ , \new_[62314]_ , \new_[62317]_ , \new_[62320]_ ,
    \new_[62321]_ , \new_[62322]_ , \new_[62326]_ , \new_[62327]_ ,
    \new_[62330]_ , \new_[62333]_ , \new_[62334]_ , \new_[62335]_ ,
    \new_[62339]_ , \new_[62340]_ , \new_[62343]_ , \new_[62346]_ ,
    \new_[62347]_ , \new_[62348]_ , \new_[62352]_ , \new_[62353]_ ,
    \new_[62356]_ , \new_[62359]_ , \new_[62360]_ , \new_[62361]_ ,
    \new_[62365]_ , \new_[62366]_ , \new_[62369]_ , \new_[62372]_ ,
    \new_[62373]_ , \new_[62374]_ , \new_[62378]_ , \new_[62379]_ ,
    \new_[62382]_ , \new_[62385]_ , \new_[62386]_ , \new_[62387]_ ,
    \new_[62391]_ , \new_[62392]_ , \new_[62395]_ , \new_[62398]_ ,
    \new_[62399]_ , \new_[62400]_ , \new_[62404]_ , \new_[62405]_ ,
    \new_[62408]_ , \new_[62411]_ , \new_[62412]_ , \new_[62413]_ ,
    \new_[62417]_ , \new_[62418]_ , \new_[62421]_ , \new_[62424]_ ,
    \new_[62425]_ , \new_[62426]_ , \new_[62430]_ , \new_[62431]_ ,
    \new_[62434]_ , \new_[62437]_ , \new_[62438]_ , \new_[62439]_ ,
    \new_[62443]_ , \new_[62444]_ , \new_[62447]_ , \new_[62450]_ ,
    \new_[62451]_ , \new_[62452]_ , \new_[62456]_ , \new_[62457]_ ,
    \new_[62460]_ , \new_[62463]_ , \new_[62464]_ , \new_[62465]_ ,
    \new_[62469]_ , \new_[62470]_ , \new_[62473]_ , \new_[62476]_ ,
    \new_[62477]_ , \new_[62478]_ , \new_[62482]_ , \new_[62483]_ ,
    \new_[62486]_ , \new_[62489]_ , \new_[62490]_ , \new_[62491]_ ,
    \new_[62495]_ , \new_[62496]_ , \new_[62499]_ , \new_[62502]_ ,
    \new_[62503]_ , \new_[62504]_ , \new_[62508]_ , \new_[62509]_ ,
    \new_[62512]_ , \new_[62515]_ , \new_[62516]_ , \new_[62517]_ ,
    \new_[62521]_ , \new_[62522]_ , \new_[62525]_ , \new_[62528]_ ,
    \new_[62529]_ , \new_[62530]_ , \new_[62534]_ , \new_[62535]_ ,
    \new_[62538]_ , \new_[62541]_ , \new_[62542]_ , \new_[62543]_ ,
    \new_[62547]_ , \new_[62548]_ , \new_[62551]_ , \new_[62554]_ ,
    \new_[62555]_ , \new_[62556]_ , \new_[62560]_ , \new_[62561]_ ,
    \new_[62564]_ , \new_[62567]_ , \new_[62568]_ , \new_[62569]_ ,
    \new_[62573]_ , \new_[62574]_ , \new_[62577]_ , \new_[62580]_ ,
    \new_[62581]_ , \new_[62582]_ , \new_[62586]_ , \new_[62587]_ ,
    \new_[62590]_ , \new_[62593]_ , \new_[62594]_ , \new_[62595]_ ,
    \new_[62599]_ , \new_[62600]_ , \new_[62603]_ , \new_[62606]_ ,
    \new_[62607]_ , \new_[62608]_ , \new_[62612]_ , \new_[62613]_ ,
    \new_[62616]_ , \new_[62619]_ , \new_[62620]_ , \new_[62621]_ ,
    \new_[62625]_ , \new_[62626]_ , \new_[62629]_ , \new_[62632]_ ,
    \new_[62633]_ , \new_[62634]_ , \new_[62638]_ , \new_[62639]_ ,
    \new_[62642]_ , \new_[62645]_ , \new_[62646]_ , \new_[62647]_ ,
    \new_[62651]_ , \new_[62652]_ , \new_[62655]_ , \new_[62658]_ ,
    \new_[62659]_ , \new_[62660]_ , \new_[62664]_ , \new_[62665]_ ,
    \new_[62668]_ , \new_[62671]_ , \new_[62672]_ , \new_[62673]_ ,
    \new_[62677]_ , \new_[62678]_ , \new_[62681]_ , \new_[62684]_ ,
    \new_[62685]_ , \new_[62686]_ , \new_[62690]_ , \new_[62691]_ ,
    \new_[62694]_ , \new_[62697]_ , \new_[62698]_ , \new_[62699]_ ,
    \new_[62703]_ , \new_[62704]_ , \new_[62707]_ , \new_[62710]_ ,
    \new_[62711]_ , \new_[62712]_ , \new_[62716]_ , \new_[62717]_ ,
    \new_[62720]_ , \new_[62723]_ , \new_[62724]_ , \new_[62725]_ ,
    \new_[62729]_ , \new_[62730]_ , \new_[62733]_ , \new_[62736]_ ,
    \new_[62737]_ , \new_[62738]_ , \new_[62742]_ , \new_[62743]_ ,
    \new_[62746]_ , \new_[62749]_ , \new_[62750]_ , \new_[62751]_ ,
    \new_[62755]_ , \new_[62756]_ , \new_[62759]_ , \new_[62762]_ ,
    \new_[62763]_ , \new_[62764]_ , \new_[62768]_ , \new_[62769]_ ,
    \new_[62772]_ , \new_[62775]_ , \new_[62776]_ , \new_[62777]_ ,
    \new_[62781]_ , \new_[62782]_ , \new_[62785]_ , \new_[62788]_ ,
    \new_[62789]_ , \new_[62790]_ , \new_[62794]_ , \new_[62795]_ ,
    \new_[62798]_ , \new_[62801]_ , \new_[62802]_ , \new_[62803]_ ,
    \new_[62807]_ , \new_[62808]_ , \new_[62811]_ , \new_[62814]_ ,
    \new_[62815]_ , \new_[62816]_ , \new_[62820]_ , \new_[62821]_ ,
    \new_[62824]_ , \new_[62827]_ , \new_[62828]_ , \new_[62829]_ ,
    \new_[62833]_ , \new_[62834]_ , \new_[62837]_ , \new_[62840]_ ,
    \new_[62841]_ , \new_[62842]_ , \new_[62846]_ , \new_[62847]_ ,
    \new_[62850]_ , \new_[62853]_ , \new_[62854]_ , \new_[62855]_ ,
    \new_[62859]_ , \new_[62860]_ , \new_[62863]_ , \new_[62866]_ ,
    \new_[62867]_ , \new_[62868]_ , \new_[62872]_ , \new_[62873]_ ,
    \new_[62876]_ , \new_[62879]_ , \new_[62880]_ , \new_[62881]_ ,
    \new_[62885]_ , \new_[62886]_ , \new_[62889]_ , \new_[62892]_ ,
    \new_[62893]_ , \new_[62894]_ , \new_[62898]_ , \new_[62899]_ ,
    \new_[62902]_ , \new_[62905]_ , \new_[62906]_ , \new_[62907]_ ,
    \new_[62911]_ , \new_[62912]_ , \new_[62915]_ , \new_[62918]_ ,
    \new_[62919]_ , \new_[62920]_ , \new_[62924]_ , \new_[62925]_ ,
    \new_[62928]_ , \new_[62931]_ , \new_[62932]_ , \new_[62933]_ ,
    \new_[62937]_ , \new_[62938]_ , \new_[62941]_ , \new_[62944]_ ,
    \new_[62945]_ , \new_[62946]_ , \new_[62950]_ , \new_[62951]_ ,
    \new_[62954]_ , \new_[62957]_ , \new_[62958]_ , \new_[62959]_ ,
    \new_[62963]_ , \new_[62964]_ , \new_[62967]_ , \new_[62970]_ ,
    \new_[62971]_ , \new_[62972]_ , \new_[62976]_ , \new_[62977]_ ,
    \new_[62980]_ , \new_[62983]_ , \new_[62984]_ , \new_[62985]_ ,
    \new_[62989]_ , \new_[62990]_ , \new_[62993]_ , \new_[62996]_ ,
    \new_[62997]_ , \new_[62998]_ , \new_[63002]_ , \new_[63003]_ ,
    \new_[63006]_ , \new_[63009]_ , \new_[63010]_ , \new_[63011]_ ,
    \new_[63015]_ , \new_[63016]_ , \new_[63019]_ , \new_[63022]_ ,
    \new_[63023]_ , \new_[63024]_ , \new_[63028]_ , \new_[63029]_ ,
    \new_[63032]_ , \new_[63035]_ , \new_[63036]_ , \new_[63037]_ ,
    \new_[63041]_ , \new_[63042]_ , \new_[63045]_ , \new_[63048]_ ,
    \new_[63049]_ , \new_[63050]_ , \new_[63054]_ , \new_[63055]_ ,
    \new_[63058]_ , \new_[63061]_ , \new_[63062]_ , \new_[63063]_ ,
    \new_[63067]_ , \new_[63068]_ , \new_[63071]_ , \new_[63074]_ ,
    \new_[63075]_ , \new_[63076]_ , \new_[63080]_ , \new_[63081]_ ,
    \new_[63084]_ , \new_[63087]_ , \new_[63088]_ , \new_[63089]_ ,
    \new_[63093]_ , \new_[63094]_ , \new_[63097]_ , \new_[63100]_ ,
    \new_[63101]_ , \new_[63102]_ , \new_[63106]_ , \new_[63107]_ ,
    \new_[63110]_ , \new_[63113]_ , \new_[63114]_ , \new_[63115]_ ,
    \new_[63119]_ , \new_[63120]_ , \new_[63123]_ , \new_[63126]_ ,
    \new_[63127]_ , \new_[63128]_ , \new_[63132]_ , \new_[63133]_ ,
    \new_[63136]_ , \new_[63139]_ , \new_[63140]_ , \new_[63141]_ ,
    \new_[63145]_ , \new_[63146]_ , \new_[63149]_ , \new_[63152]_ ,
    \new_[63153]_ , \new_[63154]_ , \new_[63158]_ , \new_[63159]_ ,
    \new_[63162]_ , \new_[63165]_ , \new_[63166]_ , \new_[63167]_ ,
    \new_[63171]_ , \new_[63172]_ , \new_[63175]_ , \new_[63178]_ ,
    \new_[63179]_ , \new_[63180]_ , \new_[63184]_ , \new_[63185]_ ,
    \new_[63188]_ , \new_[63191]_ , \new_[63192]_ , \new_[63193]_ ,
    \new_[63197]_ , \new_[63198]_ , \new_[63201]_ , \new_[63204]_ ,
    \new_[63205]_ , \new_[63206]_ , \new_[63210]_ , \new_[63211]_ ,
    \new_[63214]_ , \new_[63217]_ , \new_[63218]_ , \new_[63219]_ ,
    \new_[63223]_ , \new_[63224]_ , \new_[63227]_ , \new_[63230]_ ,
    \new_[63231]_ , \new_[63232]_ , \new_[63236]_ , \new_[63237]_ ,
    \new_[63240]_ , \new_[63243]_ , \new_[63244]_ , \new_[63245]_ ,
    \new_[63249]_ , \new_[63250]_ , \new_[63253]_ , \new_[63256]_ ,
    \new_[63257]_ , \new_[63258]_ , \new_[63262]_ , \new_[63263]_ ,
    \new_[63266]_ , \new_[63269]_ , \new_[63270]_ , \new_[63271]_ ,
    \new_[63275]_ , \new_[63276]_ , \new_[63279]_ , \new_[63282]_ ,
    \new_[63283]_ , \new_[63284]_ , \new_[63288]_ , \new_[63289]_ ,
    \new_[63292]_ , \new_[63295]_ , \new_[63296]_ , \new_[63297]_ ,
    \new_[63301]_ , \new_[63302]_ , \new_[63305]_ , \new_[63308]_ ,
    \new_[63309]_ , \new_[63310]_ , \new_[63314]_ , \new_[63315]_ ,
    \new_[63318]_ , \new_[63321]_ , \new_[63322]_ , \new_[63323]_ ,
    \new_[63327]_ , \new_[63328]_ , \new_[63331]_ , \new_[63334]_ ,
    \new_[63335]_ , \new_[63336]_ , \new_[63340]_ , \new_[63341]_ ,
    \new_[63344]_ , \new_[63347]_ , \new_[63348]_ , \new_[63349]_ ,
    \new_[63353]_ , \new_[63354]_ , \new_[63357]_ , \new_[63360]_ ,
    \new_[63361]_ , \new_[63362]_ , \new_[63366]_ , \new_[63367]_ ,
    \new_[63370]_ , \new_[63373]_ , \new_[63374]_ , \new_[63375]_ ,
    \new_[63379]_ , \new_[63380]_ , \new_[63383]_ , \new_[63386]_ ,
    \new_[63387]_ , \new_[63388]_ , \new_[63392]_ , \new_[63393]_ ,
    \new_[63396]_ , \new_[63399]_ , \new_[63400]_ , \new_[63401]_ ,
    \new_[63405]_ , \new_[63406]_ , \new_[63409]_ , \new_[63412]_ ,
    \new_[63413]_ , \new_[63414]_ , \new_[63418]_ , \new_[63419]_ ,
    \new_[63422]_ , \new_[63425]_ , \new_[63426]_ , \new_[63427]_ ,
    \new_[63431]_ , \new_[63432]_ , \new_[63435]_ , \new_[63438]_ ,
    \new_[63439]_ , \new_[63440]_ , \new_[63444]_ , \new_[63445]_ ,
    \new_[63448]_ , \new_[63451]_ , \new_[63452]_ , \new_[63453]_ ,
    \new_[63457]_ , \new_[63458]_ , \new_[63461]_ , \new_[63464]_ ,
    \new_[63465]_ , \new_[63466]_ , \new_[63470]_ , \new_[63471]_ ,
    \new_[63474]_ , \new_[63477]_ , \new_[63478]_ , \new_[63479]_ ,
    \new_[63483]_ , \new_[63484]_ , \new_[63487]_ , \new_[63490]_ ,
    \new_[63491]_ , \new_[63492]_ , \new_[63496]_ , \new_[63497]_ ,
    \new_[63500]_ , \new_[63503]_ , \new_[63504]_ , \new_[63505]_ ,
    \new_[63509]_ , \new_[63510]_ , \new_[63513]_ , \new_[63516]_ ,
    \new_[63517]_ , \new_[63518]_ , \new_[63522]_ , \new_[63523]_ ,
    \new_[63526]_ , \new_[63529]_ , \new_[63530]_ , \new_[63531]_ ,
    \new_[63535]_ , \new_[63536]_ , \new_[63539]_ , \new_[63542]_ ,
    \new_[63543]_ , \new_[63544]_ , \new_[63548]_ , \new_[63549]_ ,
    \new_[63552]_ , \new_[63555]_ , \new_[63556]_ , \new_[63557]_ ,
    \new_[63561]_ , \new_[63562]_ , \new_[63565]_ , \new_[63568]_ ,
    \new_[63569]_ , \new_[63570]_ , \new_[63574]_ , \new_[63575]_ ,
    \new_[63578]_ , \new_[63581]_ , \new_[63582]_ , \new_[63583]_ ,
    \new_[63587]_ , \new_[63588]_ , \new_[63591]_ , \new_[63594]_ ,
    \new_[63595]_ , \new_[63596]_ , \new_[63600]_ , \new_[63601]_ ,
    \new_[63604]_ , \new_[63607]_ , \new_[63608]_ , \new_[63609]_ ,
    \new_[63613]_ , \new_[63614]_ , \new_[63617]_ , \new_[63620]_ ,
    \new_[63621]_ , \new_[63622]_ , \new_[63626]_ , \new_[63627]_ ,
    \new_[63630]_ , \new_[63633]_ , \new_[63634]_ , \new_[63635]_ ,
    \new_[63639]_ , \new_[63640]_ , \new_[63643]_ , \new_[63646]_ ,
    \new_[63647]_ , \new_[63648]_ , \new_[63652]_ , \new_[63653]_ ,
    \new_[63656]_ , \new_[63659]_ , \new_[63660]_ , \new_[63661]_ ,
    \new_[63665]_ , \new_[63666]_ , \new_[63669]_ , \new_[63672]_ ,
    \new_[63673]_ , \new_[63674]_ , \new_[63678]_ , \new_[63679]_ ,
    \new_[63682]_ , \new_[63685]_ , \new_[63686]_ , \new_[63687]_ ,
    \new_[63691]_ , \new_[63692]_ , \new_[63695]_ , \new_[63698]_ ,
    \new_[63699]_ , \new_[63700]_ , \new_[63704]_ , \new_[63705]_ ,
    \new_[63708]_ , \new_[63711]_ , \new_[63712]_ , \new_[63713]_ ,
    \new_[63717]_ , \new_[63718]_ , \new_[63721]_ , \new_[63724]_ ,
    \new_[63725]_ , \new_[63726]_ , \new_[63730]_ , \new_[63731]_ ,
    \new_[63734]_ , \new_[63737]_ , \new_[63738]_ , \new_[63739]_ ,
    \new_[63743]_ , \new_[63744]_ , \new_[63747]_ , \new_[63750]_ ,
    \new_[63751]_ , \new_[63752]_ , \new_[63756]_ , \new_[63757]_ ,
    \new_[63760]_ , \new_[63763]_ , \new_[63764]_ , \new_[63765]_ ,
    \new_[63769]_ , \new_[63770]_ , \new_[63773]_ , \new_[63776]_ ,
    \new_[63777]_ , \new_[63778]_ , \new_[63782]_ , \new_[63783]_ ,
    \new_[63786]_ , \new_[63789]_ , \new_[63790]_ , \new_[63791]_ ,
    \new_[63795]_ , \new_[63796]_ , \new_[63799]_ , \new_[63802]_ ,
    \new_[63803]_ , \new_[63804]_ , \new_[63808]_ , \new_[63809]_ ,
    \new_[63812]_ , \new_[63815]_ , \new_[63816]_ , \new_[63817]_ ,
    \new_[63821]_ , \new_[63822]_ , \new_[63825]_ , \new_[63828]_ ,
    \new_[63829]_ , \new_[63830]_ , \new_[63834]_ , \new_[63835]_ ,
    \new_[63838]_ , \new_[63841]_ , \new_[63842]_ , \new_[63843]_ ,
    \new_[63847]_ , \new_[63848]_ , \new_[63851]_ , \new_[63854]_ ,
    \new_[63855]_ , \new_[63856]_ , \new_[63860]_ , \new_[63861]_ ,
    \new_[63864]_ , \new_[63867]_ , \new_[63868]_ , \new_[63869]_ ,
    \new_[63873]_ , \new_[63874]_ , \new_[63877]_ , \new_[63880]_ ,
    \new_[63881]_ , \new_[63882]_ , \new_[63886]_ , \new_[63887]_ ,
    \new_[63890]_ , \new_[63893]_ , \new_[63894]_ , \new_[63895]_ ,
    \new_[63899]_ , \new_[63900]_ , \new_[63903]_ , \new_[63906]_ ,
    \new_[63907]_ , \new_[63908]_ , \new_[63912]_ , \new_[63913]_ ,
    \new_[63916]_ , \new_[63919]_ , \new_[63920]_ , \new_[63921]_ ,
    \new_[63925]_ , \new_[63926]_ , \new_[63929]_ , \new_[63932]_ ,
    \new_[63933]_ , \new_[63934]_ , \new_[63938]_ , \new_[63939]_ ,
    \new_[63942]_ , \new_[63945]_ , \new_[63946]_ , \new_[63947]_ ,
    \new_[63951]_ , \new_[63952]_ , \new_[63955]_ , \new_[63958]_ ,
    \new_[63959]_ , \new_[63960]_ , \new_[63964]_ , \new_[63965]_ ,
    \new_[63968]_ , \new_[63971]_ , \new_[63972]_ , \new_[63973]_ ,
    \new_[63977]_ , \new_[63978]_ , \new_[63981]_ , \new_[63984]_ ,
    \new_[63985]_ , \new_[63986]_ , \new_[63990]_ , \new_[63991]_ ,
    \new_[63994]_ , \new_[63997]_ , \new_[63998]_ , \new_[63999]_ ,
    \new_[64003]_ , \new_[64004]_ , \new_[64007]_ , \new_[64010]_ ,
    \new_[64011]_ , \new_[64012]_ , \new_[64016]_ , \new_[64017]_ ,
    \new_[64020]_ , \new_[64023]_ , \new_[64024]_ , \new_[64025]_ ,
    \new_[64029]_ , \new_[64030]_ , \new_[64033]_ , \new_[64036]_ ,
    \new_[64037]_ , \new_[64038]_ , \new_[64042]_ , \new_[64043]_ ,
    \new_[64046]_ , \new_[64049]_ , \new_[64050]_ , \new_[64051]_ ,
    \new_[64055]_ , \new_[64056]_ , \new_[64059]_ , \new_[64062]_ ,
    \new_[64063]_ , \new_[64064]_ , \new_[64068]_ , \new_[64069]_ ,
    \new_[64072]_ , \new_[64075]_ , \new_[64076]_ , \new_[64077]_ ,
    \new_[64081]_ , \new_[64082]_ , \new_[64085]_ , \new_[64088]_ ,
    \new_[64089]_ , \new_[64090]_ , \new_[64094]_ , \new_[64095]_ ,
    \new_[64098]_ , \new_[64101]_ , \new_[64102]_ , \new_[64103]_ ,
    \new_[64107]_ , \new_[64108]_ , \new_[64111]_ , \new_[64114]_ ,
    \new_[64115]_ , \new_[64116]_ , \new_[64120]_ , \new_[64121]_ ,
    \new_[64124]_ , \new_[64127]_ , \new_[64128]_ , \new_[64129]_ ,
    \new_[64133]_ , \new_[64134]_ , \new_[64137]_ , \new_[64140]_ ,
    \new_[64141]_ , \new_[64142]_ , \new_[64146]_ , \new_[64147]_ ,
    \new_[64150]_ , \new_[64153]_ , \new_[64154]_ , \new_[64155]_ ,
    \new_[64159]_ , \new_[64160]_ , \new_[64163]_ , \new_[64166]_ ,
    \new_[64167]_ , \new_[64168]_ , \new_[64172]_ , \new_[64173]_ ,
    \new_[64176]_ , \new_[64179]_ , \new_[64180]_ , \new_[64181]_ ,
    \new_[64185]_ , \new_[64186]_ , \new_[64189]_ , \new_[64192]_ ,
    \new_[64193]_ , \new_[64194]_ , \new_[64198]_ , \new_[64199]_ ,
    \new_[64202]_ , \new_[64205]_ , \new_[64206]_ , \new_[64207]_ ,
    \new_[64211]_ , \new_[64212]_ , \new_[64215]_ , \new_[64218]_ ,
    \new_[64219]_ , \new_[64220]_ , \new_[64224]_ , \new_[64225]_ ,
    \new_[64228]_ , \new_[64231]_ , \new_[64232]_ , \new_[64233]_ ,
    \new_[64237]_ , \new_[64238]_ , \new_[64241]_ , \new_[64244]_ ,
    \new_[64245]_ , \new_[64246]_ , \new_[64250]_ , \new_[64251]_ ,
    \new_[64254]_ , \new_[64257]_ , \new_[64258]_ , \new_[64259]_ ,
    \new_[64263]_ , \new_[64264]_ , \new_[64267]_ , \new_[64270]_ ,
    \new_[64271]_ , \new_[64272]_ , \new_[64276]_ , \new_[64277]_ ,
    \new_[64280]_ , \new_[64283]_ , \new_[64284]_ , \new_[64285]_ ,
    \new_[64289]_ , \new_[64290]_ , \new_[64293]_ , \new_[64296]_ ,
    \new_[64297]_ , \new_[64298]_ , \new_[64302]_ , \new_[64303]_ ,
    \new_[64306]_ , \new_[64309]_ , \new_[64310]_ , \new_[64311]_ ,
    \new_[64315]_ , \new_[64316]_ , \new_[64319]_ , \new_[64322]_ ,
    \new_[64323]_ , \new_[64324]_ , \new_[64328]_ , \new_[64329]_ ,
    \new_[64332]_ , \new_[64335]_ , \new_[64336]_ , \new_[64337]_ ,
    \new_[64341]_ , \new_[64342]_ , \new_[64345]_ , \new_[64348]_ ,
    \new_[64349]_ , \new_[64350]_ , \new_[64354]_ , \new_[64355]_ ,
    \new_[64358]_ , \new_[64361]_ , \new_[64362]_ , \new_[64363]_ ,
    \new_[64367]_ , \new_[64368]_ , \new_[64371]_ , \new_[64374]_ ,
    \new_[64375]_ , \new_[64376]_ , \new_[64380]_ , \new_[64381]_ ,
    \new_[64384]_ , \new_[64387]_ , \new_[64388]_ , \new_[64389]_ ,
    \new_[64393]_ , \new_[64394]_ , \new_[64397]_ , \new_[64400]_ ,
    \new_[64401]_ , \new_[64402]_ , \new_[64406]_ , \new_[64407]_ ,
    \new_[64410]_ , \new_[64413]_ , \new_[64414]_ , \new_[64415]_ ,
    \new_[64419]_ , \new_[64420]_ , \new_[64423]_ , \new_[64426]_ ,
    \new_[64427]_ , \new_[64428]_ , \new_[64432]_ , \new_[64433]_ ,
    \new_[64436]_ , \new_[64439]_ , \new_[64440]_ , \new_[64441]_ ,
    \new_[64445]_ , \new_[64446]_ , \new_[64449]_ , \new_[64452]_ ,
    \new_[64453]_ , \new_[64454]_ , \new_[64458]_ , \new_[64459]_ ,
    \new_[64462]_ , \new_[64465]_ , \new_[64466]_ , \new_[64467]_ ,
    \new_[64471]_ , \new_[64472]_ , \new_[64475]_ , \new_[64478]_ ,
    \new_[64479]_ , \new_[64480]_ , \new_[64484]_ , \new_[64485]_ ,
    \new_[64488]_ , \new_[64491]_ , \new_[64492]_ , \new_[64493]_ ,
    \new_[64497]_ , \new_[64498]_ , \new_[64501]_ , \new_[64504]_ ,
    \new_[64505]_ , \new_[64506]_ , \new_[64510]_ , \new_[64511]_ ,
    \new_[64514]_ , \new_[64517]_ , \new_[64518]_ , \new_[64519]_ ,
    \new_[64523]_ , \new_[64524]_ , \new_[64527]_ , \new_[64530]_ ,
    \new_[64531]_ , \new_[64532]_ , \new_[64536]_ , \new_[64537]_ ,
    \new_[64540]_ , \new_[64543]_ , \new_[64544]_ , \new_[64545]_ ,
    \new_[64549]_ , \new_[64550]_ , \new_[64553]_ , \new_[64556]_ ,
    \new_[64557]_ , \new_[64558]_ , \new_[64562]_ , \new_[64563]_ ,
    \new_[64566]_ , \new_[64569]_ , \new_[64570]_ , \new_[64571]_ ,
    \new_[64575]_ , \new_[64576]_ , \new_[64579]_ , \new_[64582]_ ,
    \new_[64583]_ , \new_[64584]_ , \new_[64588]_ , \new_[64589]_ ,
    \new_[64592]_ , \new_[64595]_ , \new_[64596]_ , \new_[64597]_ ,
    \new_[64601]_ , \new_[64602]_ , \new_[64605]_ , \new_[64608]_ ,
    \new_[64609]_ , \new_[64610]_ , \new_[64614]_ , \new_[64615]_ ,
    \new_[64618]_ , \new_[64621]_ , \new_[64622]_ , \new_[64623]_ ,
    \new_[64627]_ , \new_[64628]_ , \new_[64631]_ , \new_[64634]_ ,
    \new_[64635]_ , \new_[64636]_ , \new_[64640]_ , \new_[64641]_ ,
    \new_[64644]_ , \new_[64647]_ , \new_[64648]_ , \new_[64649]_ ,
    \new_[64653]_ , \new_[64654]_ , \new_[64657]_ , \new_[64660]_ ,
    \new_[64661]_ , \new_[64662]_ , \new_[64666]_ , \new_[64667]_ ,
    \new_[64670]_ , \new_[64673]_ , \new_[64674]_ , \new_[64675]_ ,
    \new_[64679]_ , \new_[64680]_ , \new_[64683]_ , \new_[64686]_ ,
    \new_[64687]_ , \new_[64688]_ , \new_[64692]_ , \new_[64693]_ ,
    \new_[64696]_ , \new_[64699]_ , \new_[64700]_ , \new_[64701]_ ,
    \new_[64705]_ , \new_[64706]_ , \new_[64709]_ , \new_[64712]_ ,
    \new_[64713]_ , \new_[64714]_ , \new_[64718]_ , \new_[64719]_ ,
    \new_[64722]_ , \new_[64725]_ , \new_[64726]_ , \new_[64727]_ ,
    \new_[64731]_ , \new_[64732]_ , \new_[64735]_ , \new_[64738]_ ,
    \new_[64739]_ , \new_[64740]_ , \new_[64744]_ , \new_[64745]_ ,
    \new_[64748]_ , \new_[64751]_ , \new_[64752]_ , \new_[64753]_ ,
    \new_[64757]_ , \new_[64758]_ , \new_[64761]_ , \new_[64764]_ ,
    \new_[64765]_ , \new_[64766]_ , \new_[64770]_ , \new_[64771]_ ,
    \new_[64774]_ , \new_[64777]_ , \new_[64778]_ , \new_[64779]_ ,
    \new_[64783]_ , \new_[64784]_ , \new_[64787]_ , \new_[64790]_ ,
    \new_[64791]_ , \new_[64792]_ , \new_[64796]_ , \new_[64797]_ ,
    \new_[64800]_ , \new_[64803]_ , \new_[64804]_ , \new_[64805]_ ,
    \new_[64809]_ , \new_[64810]_ , \new_[64813]_ , \new_[64816]_ ,
    \new_[64817]_ , \new_[64818]_ , \new_[64822]_ , \new_[64823]_ ,
    \new_[64826]_ , \new_[64829]_ , \new_[64830]_ , \new_[64831]_ ,
    \new_[64835]_ , \new_[64836]_ , \new_[64839]_ , \new_[64842]_ ,
    \new_[64843]_ , \new_[64844]_ , \new_[64848]_ , \new_[64849]_ ,
    \new_[64852]_ , \new_[64855]_ , \new_[64856]_ , \new_[64857]_ ,
    \new_[64861]_ , \new_[64862]_ , \new_[64865]_ , \new_[64868]_ ,
    \new_[64869]_ , \new_[64870]_ , \new_[64874]_ , \new_[64875]_ ,
    \new_[64878]_ , \new_[64881]_ , \new_[64882]_ , \new_[64883]_ ,
    \new_[64887]_ , \new_[64888]_ , \new_[64891]_ , \new_[64894]_ ,
    \new_[64895]_ , \new_[64896]_ , \new_[64900]_ , \new_[64901]_ ,
    \new_[64904]_ , \new_[64907]_ , \new_[64908]_ , \new_[64909]_ ,
    \new_[64913]_ , \new_[64914]_ , \new_[64917]_ , \new_[64920]_ ,
    \new_[64921]_ , \new_[64922]_ , \new_[64926]_ , \new_[64927]_ ,
    \new_[64930]_ , \new_[64933]_ , \new_[64934]_ , \new_[64935]_ ,
    \new_[64939]_ , \new_[64940]_ , \new_[64943]_ , \new_[64946]_ ,
    \new_[64947]_ , \new_[64948]_ , \new_[64952]_ , \new_[64953]_ ,
    \new_[64956]_ , \new_[64959]_ , \new_[64960]_ , \new_[64961]_ ,
    \new_[64965]_ , \new_[64966]_ , \new_[64969]_ , \new_[64972]_ ,
    \new_[64973]_ , \new_[64974]_ , \new_[64978]_ , \new_[64979]_ ,
    \new_[64982]_ , \new_[64985]_ , \new_[64986]_ , \new_[64987]_ ,
    \new_[64991]_ , \new_[64992]_ , \new_[64995]_ , \new_[64998]_ ,
    \new_[64999]_ , \new_[65000]_ , \new_[65004]_ , \new_[65005]_ ,
    \new_[65008]_ , \new_[65011]_ , \new_[65012]_ , \new_[65013]_ ,
    \new_[65017]_ , \new_[65018]_ , \new_[65021]_ , \new_[65024]_ ,
    \new_[65025]_ , \new_[65026]_ , \new_[65030]_ , \new_[65031]_ ,
    \new_[65034]_ , \new_[65037]_ , \new_[65038]_ , \new_[65039]_ ,
    \new_[65043]_ , \new_[65044]_ , \new_[65047]_ , \new_[65050]_ ,
    \new_[65051]_ , \new_[65052]_ , \new_[65056]_ , \new_[65057]_ ,
    \new_[65060]_ , \new_[65063]_ , \new_[65064]_ , \new_[65065]_ ,
    \new_[65069]_ , \new_[65070]_ , \new_[65073]_ , \new_[65076]_ ,
    \new_[65077]_ , \new_[65078]_ , \new_[65082]_ , \new_[65083]_ ,
    \new_[65086]_ , \new_[65089]_ , \new_[65090]_ , \new_[65091]_ ,
    \new_[65095]_ , \new_[65096]_ , \new_[65099]_ , \new_[65102]_ ,
    \new_[65103]_ , \new_[65104]_ , \new_[65108]_ , \new_[65109]_ ,
    \new_[65112]_ , \new_[65115]_ , \new_[65116]_ , \new_[65117]_ ,
    \new_[65121]_ , \new_[65122]_ , \new_[65125]_ , \new_[65128]_ ,
    \new_[65129]_ , \new_[65130]_ , \new_[65134]_ , \new_[65135]_ ,
    \new_[65138]_ , \new_[65141]_ , \new_[65142]_ , \new_[65143]_ ,
    \new_[65147]_ , \new_[65148]_ , \new_[65151]_ , \new_[65154]_ ,
    \new_[65155]_ , \new_[65156]_ , \new_[65160]_ , \new_[65161]_ ,
    \new_[65164]_ , \new_[65167]_ , \new_[65168]_ , \new_[65169]_ ,
    \new_[65173]_ , \new_[65174]_ , \new_[65177]_ , \new_[65180]_ ,
    \new_[65181]_ , \new_[65182]_ , \new_[65186]_ , \new_[65187]_ ,
    \new_[65190]_ , \new_[65193]_ , \new_[65194]_ , \new_[65195]_ ,
    \new_[65199]_ , \new_[65200]_ , \new_[65203]_ , \new_[65206]_ ,
    \new_[65207]_ , \new_[65208]_ , \new_[65212]_ , \new_[65213]_ ,
    \new_[65216]_ , \new_[65219]_ , \new_[65220]_ , \new_[65221]_ ,
    \new_[65225]_ , \new_[65226]_ , \new_[65229]_ , \new_[65232]_ ,
    \new_[65233]_ , \new_[65234]_ , \new_[65238]_ , \new_[65239]_ ,
    \new_[65242]_ , \new_[65245]_ , \new_[65246]_ , \new_[65247]_ ,
    \new_[65251]_ , \new_[65252]_ , \new_[65255]_ , \new_[65258]_ ,
    \new_[65259]_ , \new_[65260]_ , \new_[65264]_ , \new_[65265]_ ,
    \new_[65268]_ , \new_[65271]_ , \new_[65272]_ , \new_[65273]_ ,
    \new_[65277]_ , \new_[65278]_ , \new_[65281]_ , \new_[65284]_ ,
    \new_[65285]_ , \new_[65286]_ , \new_[65290]_ , \new_[65291]_ ,
    \new_[65294]_ , \new_[65297]_ , \new_[65298]_ , \new_[65299]_ ,
    \new_[65303]_ , \new_[65304]_ , \new_[65307]_ , \new_[65310]_ ,
    \new_[65311]_ , \new_[65312]_ , \new_[65316]_ , \new_[65317]_ ,
    \new_[65320]_ , \new_[65323]_ , \new_[65324]_ , \new_[65325]_ ,
    \new_[65329]_ , \new_[65330]_ , \new_[65333]_ , \new_[65336]_ ,
    \new_[65337]_ , \new_[65338]_ , \new_[65342]_ , \new_[65343]_ ,
    \new_[65346]_ , \new_[65349]_ , \new_[65350]_ , \new_[65351]_ ,
    \new_[65355]_ , \new_[65356]_ , \new_[65359]_ , \new_[65362]_ ,
    \new_[65363]_ , \new_[65364]_ , \new_[65368]_ , \new_[65369]_ ,
    \new_[65372]_ , \new_[65375]_ , \new_[65376]_ , \new_[65377]_ ,
    \new_[65381]_ , \new_[65382]_ , \new_[65385]_ , \new_[65388]_ ,
    \new_[65389]_ , \new_[65390]_ , \new_[65394]_ , \new_[65395]_ ,
    \new_[65398]_ , \new_[65401]_ , \new_[65402]_ , \new_[65403]_ ,
    \new_[65407]_ , \new_[65408]_ , \new_[65411]_ , \new_[65414]_ ,
    \new_[65415]_ , \new_[65416]_ , \new_[65420]_ , \new_[65421]_ ,
    \new_[65424]_ , \new_[65427]_ , \new_[65428]_ , \new_[65429]_ ,
    \new_[65433]_ , \new_[65434]_ , \new_[65437]_ , \new_[65440]_ ,
    \new_[65441]_ , \new_[65442]_ , \new_[65446]_ , \new_[65447]_ ,
    \new_[65450]_ , \new_[65453]_ , \new_[65454]_ , \new_[65455]_ ,
    \new_[65459]_ , \new_[65460]_ , \new_[65463]_ , \new_[65466]_ ,
    \new_[65467]_ , \new_[65468]_ , \new_[65472]_ , \new_[65473]_ ,
    \new_[65476]_ , \new_[65479]_ , \new_[65480]_ , \new_[65481]_ ,
    \new_[65485]_ , \new_[65486]_ , \new_[65489]_ , \new_[65492]_ ,
    \new_[65493]_ , \new_[65494]_ , \new_[65498]_ , \new_[65499]_ ,
    \new_[65502]_ , \new_[65505]_ , \new_[65506]_ , \new_[65507]_ ,
    \new_[65511]_ , \new_[65512]_ , \new_[65515]_ , \new_[65518]_ ,
    \new_[65519]_ , \new_[65520]_ , \new_[65524]_ , \new_[65525]_ ,
    \new_[65528]_ , \new_[65531]_ , \new_[65532]_ , \new_[65533]_ ,
    \new_[65537]_ , \new_[65538]_ , \new_[65541]_ , \new_[65544]_ ,
    \new_[65545]_ , \new_[65546]_ , \new_[65550]_ , \new_[65551]_ ,
    \new_[65554]_ , \new_[65557]_ , \new_[65558]_ , \new_[65559]_ ,
    \new_[65563]_ , \new_[65564]_ , \new_[65567]_ , \new_[65570]_ ,
    \new_[65571]_ , \new_[65572]_ , \new_[65576]_ , \new_[65577]_ ,
    \new_[65580]_ , \new_[65583]_ , \new_[65584]_ , \new_[65585]_ ,
    \new_[65589]_ , \new_[65590]_ , \new_[65593]_ , \new_[65596]_ ,
    \new_[65597]_ , \new_[65598]_ , \new_[65602]_ , \new_[65603]_ ,
    \new_[65606]_ , \new_[65609]_ , \new_[65610]_ , \new_[65611]_ ,
    \new_[65615]_ , \new_[65616]_ , \new_[65619]_ , \new_[65622]_ ,
    \new_[65623]_ , \new_[65624]_ , \new_[65628]_ , \new_[65629]_ ,
    \new_[65632]_ , \new_[65635]_ , \new_[65636]_ , \new_[65637]_ ,
    \new_[65641]_ , \new_[65642]_ , \new_[65645]_ , \new_[65648]_ ,
    \new_[65649]_ , \new_[65650]_ , \new_[65654]_ , \new_[65655]_ ,
    \new_[65658]_ , \new_[65661]_ , \new_[65662]_ , \new_[65663]_ ,
    \new_[65667]_ , \new_[65668]_ , \new_[65671]_ , \new_[65674]_ ,
    \new_[65675]_ , \new_[65676]_ , \new_[65680]_ , \new_[65681]_ ,
    \new_[65684]_ , \new_[65687]_ , \new_[65688]_ , \new_[65689]_ ,
    \new_[65693]_ , \new_[65694]_ , \new_[65697]_ , \new_[65700]_ ,
    \new_[65701]_ , \new_[65702]_ , \new_[65706]_ , \new_[65707]_ ,
    \new_[65710]_ , \new_[65713]_ , \new_[65714]_ , \new_[65715]_ ,
    \new_[65719]_ , \new_[65720]_ , \new_[65723]_ , \new_[65726]_ ,
    \new_[65727]_ , \new_[65728]_ , \new_[65732]_ , \new_[65733]_ ,
    \new_[65736]_ , \new_[65739]_ , \new_[65740]_ , \new_[65741]_ ,
    \new_[65745]_ , \new_[65746]_ , \new_[65749]_ , \new_[65752]_ ,
    \new_[65753]_ , \new_[65754]_ , \new_[65758]_ , \new_[65759]_ ,
    \new_[65762]_ , \new_[65765]_ , \new_[65766]_ , \new_[65767]_ ,
    \new_[65771]_ , \new_[65772]_ , \new_[65775]_ , \new_[65778]_ ,
    \new_[65779]_ , \new_[65780]_ , \new_[65784]_ , \new_[65785]_ ,
    \new_[65788]_ , \new_[65791]_ , \new_[65792]_ , \new_[65793]_ ,
    \new_[65797]_ , \new_[65798]_ , \new_[65801]_ , \new_[65804]_ ,
    \new_[65805]_ , \new_[65806]_ , \new_[65810]_ , \new_[65811]_ ,
    \new_[65814]_ , \new_[65817]_ , \new_[65818]_ , \new_[65819]_ ,
    \new_[65823]_ , \new_[65824]_ , \new_[65827]_ , \new_[65830]_ ,
    \new_[65831]_ , \new_[65832]_ , \new_[65836]_ , \new_[65837]_ ,
    \new_[65840]_ , \new_[65843]_ , \new_[65844]_ , \new_[65845]_ ,
    \new_[65849]_ , \new_[65850]_ , \new_[65853]_ , \new_[65856]_ ,
    \new_[65857]_ , \new_[65858]_ , \new_[65862]_ , \new_[65863]_ ,
    \new_[65866]_ , \new_[65869]_ , \new_[65870]_ , \new_[65871]_ ,
    \new_[65875]_ , \new_[65876]_ , \new_[65879]_ , \new_[65882]_ ,
    \new_[65883]_ , \new_[65884]_ , \new_[65888]_ , \new_[65889]_ ,
    \new_[65892]_ , \new_[65895]_ , \new_[65896]_ , \new_[65897]_ ,
    \new_[65901]_ , \new_[65902]_ , \new_[65905]_ , \new_[65908]_ ,
    \new_[65909]_ , \new_[65910]_ , \new_[65914]_ , \new_[65915]_ ,
    \new_[65918]_ , \new_[65921]_ , \new_[65922]_ , \new_[65923]_ ,
    \new_[65927]_ , \new_[65928]_ , \new_[65931]_ , \new_[65934]_ ,
    \new_[65935]_ , \new_[65936]_ , \new_[65940]_ , \new_[65941]_ ,
    \new_[65944]_ , \new_[65947]_ , \new_[65948]_ , \new_[65949]_ ,
    \new_[65953]_ , \new_[65954]_ , \new_[65957]_ , \new_[65960]_ ,
    \new_[65961]_ , \new_[65962]_ , \new_[65966]_ , \new_[65967]_ ,
    \new_[65970]_ , \new_[65973]_ , \new_[65974]_ , \new_[65975]_ ,
    \new_[65979]_ , \new_[65980]_ , \new_[65983]_ , \new_[65986]_ ,
    \new_[65987]_ , \new_[65988]_ , \new_[65992]_ , \new_[65993]_ ,
    \new_[65996]_ , \new_[65999]_ , \new_[66000]_ , \new_[66001]_ ,
    \new_[66005]_ , \new_[66006]_ , \new_[66009]_ , \new_[66012]_ ,
    \new_[66013]_ , \new_[66014]_ , \new_[66018]_ , \new_[66019]_ ,
    \new_[66022]_ , \new_[66025]_ , \new_[66026]_ , \new_[66027]_ ,
    \new_[66031]_ , \new_[66032]_ , \new_[66035]_ , \new_[66038]_ ,
    \new_[66039]_ , \new_[66040]_ , \new_[66044]_ , \new_[66045]_ ,
    \new_[66048]_ , \new_[66051]_ , \new_[66052]_ , \new_[66053]_ ,
    \new_[66057]_ , \new_[66058]_ , \new_[66061]_ , \new_[66064]_ ,
    \new_[66065]_ , \new_[66066]_ , \new_[66070]_ , \new_[66071]_ ,
    \new_[66074]_ , \new_[66077]_ , \new_[66078]_ , \new_[66079]_ ,
    \new_[66083]_ , \new_[66084]_ , \new_[66087]_ , \new_[66090]_ ,
    \new_[66091]_ , \new_[66092]_ , \new_[66096]_ , \new_[66097]_ ,
    \new_[66100]_ , \new_[66103]_ , \new_[66104]_ , \new_[66105]_ ,
    \new_[66109]_ , \new_[66110]_ , \new_[66113]_ , \new_[66116]_ ,
    \new_[66117]_ , \new_[66118]_ , \new_[66122]_ , \new_[66123]_ ,
    \new_[66126]_ , \new_[66129]_ , \new_[66130]_ , \new_[66131]_ ,
    \new_[66135]_ , \new_[66136]_ , \new_[66139]_ , \new_[66142]_ ,
    \new_[66143]_ , \new_[66144]_ , \new_[66148]_ , \new_[66149]_ ,
    \new_[66152]_ , \new_[66155]_ , \new_[66156]_ , \new_[66157]_ ,
    \new_[66161]_ , \new_[66162]_ , \new_[66165]_ , \new_[66168]_ ,
    \new_[66169]_ , \new_[66170]_ , \new_[66174]_ , \new_[66175]_ ,
    \new_[66178]_ , \new_[66181]_ , \new_[66182]_ , \new_[66183]_ ,
    \new_[66187]_ , \new_[66188]_ , \new_[66191]_ , \new_[66194]_ ,
    \new_[66195]_ , \new_[66196]_ , \new_[66200]_ , \new_[66201]_ ,
    \new_[66204]_ , \new_[66207]_ , \new_[66208]_ , \new_[66209]_ ,
    \new_[66213]_ , \new_[66214]_ , \new_[66217]_ , \new_[66220]_ ,
    \new_[66221]_ , \new_[66222]_ , \new_[66226]_ , \new_[66227]_ ,
    \new_[66230]_ , \new_[66233]_ , \new_[66234]_ , \new_[66235]_ ,
    \new_[66239]_ , \new_[66240]_ , \new_[66243]_ , \new_[66246]_ ,
    \new_[66247]_ , \new_[66248]_ , \new_[66252]_ , \new_[66253]_ ,
    \new_[66256]_ , \new_[66259]_ , \new_[66260]_ , \new_[66261]_ ,
    \new_[66265]_ , \new_[66266]_ , \new_[66269]_ , \new_[66272]_ ,
    \new_[66273]_ , \new_[66274]_ , \new_[66278]_ , \new_[66279]_ ,
    \new_[66282]_ , \new_[66285]_ , \new_[66286]_ , \new_[66287]_ ,
    \new_[66291]_ , \new_[66292]_ , \new_[66295]_ , \new_[66298]_ ,
    \new_[66299]_ , \new_[66300]_ , \new_[66304]_ , \new_[66305]_ ,
    \new_[66308]_ , \new_[66311]_ , \new_[66312]_ , \new_[66313]_ ,
    \new_[66317]_ , \new_[66318]_ , \new_[66321]_ , \new_[66324]_ ,
    \new_[66325]_ , \new_[66326]_ , \new_[66330]_ , \new_[66331]_ ,
    \new_[66334]_ , \new_[66337]_ , \new_[66338]_ , \new_[66339]_ ,
    \new_[66343]_ , \new_[66344]_ , \new_[66347]_ , \new_[66350]_ ,
    \new_[66351]_ , \new_[66352]_ , \new_[66356]_ , \new_[66357]_ ,
    \new_[66360]_ , \new_[66363]_ , \new_[66364]_ , \new_[66365]_ ,
    \new_[66369]_ , \new_[66370]_ , \new_[66373]_ , \new_[66376]_ ,
    \new_[66377]_ , \new_[66378]_ , \new_[66382]_ , \new_[66383]_ ,
    \new_[66386]_ , \new_[66389]_ , \new_[66390]_ , \new_[66391]_ ,
    \new_[66395]_ , \new_[66396]_ , \new_[66399]_ , \new_[66402]_ ,
    \new_[66403]_ , \new_[66404]_ , \new_[66408]_ , \new_[66409]_ ,
    \new_[66412]_ , \new_[66415]_ , \new_[66416]_ , \new_[66417]_ ,
    \new_[66421]_ , \new_[66422]_ , \new_[66425]_ , \new_[66428]_ ,
    \new_[66429]_ , \new_[66430]_ , \new_[66434]_ , \new_[66435]_ ,
    \new_[66438]_ , \new_[66441]_ , \new_[66442]_ , \new_[66443]_ ,
    \new_[66447]_ , \new_[66448]_ , \new_[66451]_ , \new_[66454]_ ,
    \new_[66455]_ , \new_[66456]_ , \new_[66460]_ , \new_[66461]_ ,
    \new_[66464]_ , \new_[66467]_ , \new_[66468]_ , \new_[66469]_ ,
    \new_[66473]_ , \new_[66474]_ , \new_[66477]_ , \new_[66480]_ ,
    \new_[66481]_ , \new_[66482]_ , \new_[66486]_ , \new_[66487]_ ,
    \new_[66490]_ , \new_[66493]_ , \new_[66494]_ , \new_[66495]_ ,
    \new_[66499]_ , \new_[66500]_ , \new_[66503]_ , \new_[66506]_ ,
    \new_[66507]_ , \new_[66508]_ , \new_[66512]_ , \new_[66513]_ ,
    \new_[66516]_ , \new_[66519]_ , \new_[66520]_ , \new_[66521]_ ,
    \new_[66525]_ , \new_[66526]_ , \new_[66529]_ , \new_[66532]_ ,
    \new_[66533]_ , \new_[66534]_ , \new_[66538]_ , \new_[66539]_ ,
    \new_[66542]_ , \new_[66545]_ , \new_[66546]_ , \new_[66547]_ ,
    \new_[66551]_ , \new_[66552]_ , \new_[66555]_ , \new_[66558]_ ,
    \new_[66559]_ , \new_[66560]_ , \new_[66564]_ , \new_[66565]_ ,
    \new_[66568]_ , \new_[66571]_ , \new_[66572]_ , \new_[66573]_ ,
    \new_[66577]_ , \new_[66578]_ , \new_[66581]_ , \new_[66584]_ ,
    \new_[66585]_ , \new_[66586]_ , \new_[66590]_ , \new_[66591]_ ,
    \new_[66594]_ , \new_[66597]_ , \new_[66598]_ , \new_[66599]_ ,
    \new_[66603]_ , \new_[66604]_ , \new_[66607]_ , \new_[66610]_ ,
    \new_[66611]_ , \new_[66612]_ , \new_[66616]_ , \new_[66617]_ ,
    \new_[66620]_ , \new_[66623]_ , \new_[66624]_ , \new_[66625]_ ,
    \new_[66629]_ , \new_[66630]_ , \new_[66633]_ , \new_[66636]_ ,
    \new_[66637]_ , \new_[66638]_ , \new_[66642]_ , \new_[66643]_ ,
    \new_[66646]_ , \new_[66649]_ , \new_[66650]_ , \new_[66651]_ ,
    \new_[66655]_ , \new_[66656]_ , \new_[66659]_ , \new_[66662]_ ,
    \new_[66663]_ , \new_[66664]_ , \new_[66668]_ , \new_[66669]_ ,
    \new_[66672]_ , \new_[66675]_ , \new_[66676]_ , \new_[66677]_ ,
    \new_[66681]_ , \new_[66682]_ , \new_[66685]_ , \new_[66688]_ ,
    \new_[66689]_ , \new_[66690]_ , \new_[66694]_ , \new_[66695]_ ,
    \new_[66698]_ , \new_[66701]_ , \new_[66702]_ , \new_[66703]_ ,
    \new_[66707]_ , \new_[66708]_ , \new_[66711]_ , \new_[66714]_ ,
    \new_[66715]_ , \new_[66716]_ , \new_[66720]_ , \new_[66721]_ ,
    \new_[66724]_ , \new_[66727]_ , \new_[66728]_ , \new_[66729]_ ,
    \new_[66733]_ , \new_[66734]_ , \new_[66737]_ , \new_[66740]_ ,
    \new_[66741]_ , \new_[66742]_ , \new_[66746]_ , \new_[66747]_ ,
    \new_[66750]_ , \new_[66753]_ , \new_[66754]_ , \new_[66755]_ ,
    \new_[66759]_ , \new_[66760]_ , \new_[66763]_ , \new_[66766]_ ,
    \new_[66767]_ , \new_[66768]_ , \new_[66772]_ , \new_[66773]_ ,
    \new_[66776]_ , \new_[66779]_ , \new_[66780]_ , \new_[66781]_ ,
    \new_[66785]_ , \new_[66786]_ , \new_[66789]_ , \new_[66792]_ ,
    \new_[66793]_ , \new_[66794]_ , \new_[66798]_ , \new_[66799]_ ,
    \new_[66802]_ , \new_[66805]_ , \new_[66806]_ , \new_[66807]_ ,
    \new_[66811]_ , \new_[66812]_ , \new_[66815]_ , \new_[66818]_ ,
    \new_[66819]_ , \new_[66820]_ , \new_[66824]_ , \new_[66825]_ ,
    \new_[66828]_ , \new_[66831]_ , \new_[66832]_ , \new_[66833]_ ,
    \new_[66837]_ , \new_[66838]_ , \new_[66841]_ , \new_[66844]_ ,
    \new_[66845]_ , \new_[66846]_ , \new_[66850]_ , \new_[66851]_ ,
    \new_[66854]_ , \new_[66857]_ , \new_[66858]_ , \new_[66859]_ ,
    \new_[66863]_ , \new_[66864]_ , \new_[66867]_ , \new_[66870]_ ,
    \new_[66871]_ , \new_[66872]_ , \new_[66876]_ , \new_[66877]_ ,
    \new_[66880]_ , \new_[66883]_ , \new_[66884]_ , \new_[66885]_ ,
    \new_[66889]_ , \new_[66890]_ , \new_[66893]_ , \new_[66896]_ ,
    \new_[66897]_ , \new_[66898]_ , \new_[66902]_ , \new_[66903]_ ,
    \new_[66906]_ , \new_[66909]_ , \new_[66910]_ , \new_[66911]_ ,
    \new_[66915]_ , \new_[66916]_ , \new_[66919]_ , \new_[66922]_ ,
    \new_[66923]_ , \new_[66924]_ , \new_[66928]_ , \new_[66929]_ ,
    \new_[66932]_ , \new_[66935]_ , \new_[66936]_ , \new_[66937]_ ,
    \new_[66941]_ , \new_[66942]_ , \new_[66945]_ , \new_[66948]_ ,
    \new_[66949]_ , \new_[66950]_ , \new_[66954]_ , \new_[66955]_ ,
    \new_[66958]_ , \new_[66961]_ , \new_[66962]_ , \new_[66963]_ ,
    \new_[66967]_ , \new_[66968]_ , \new_[66971]_ , \new_[66974]_ ,
    \new_[66975]_ , \new_[66976]_ , \new_[66980]_ , \new_[66981]_ ,
    \new_[66984]_ , \new_[66987]_ , \new_[66988]_ , \new_[66989]_ ,
    \new_[66993]_ , \new_[66994]_ , \new_[66997]_ , \new_[67000]_ ,
    \new_[67001]_ , \new_[67002]_ , \new_[67006]_ , \new_[67007]_ ,
    \new_[67010]_ , \new_[67013]_ , \new_[67014]_ , \new_[67015]_ ,
    \new_[67019]_ , \new_[67020]_ , \new_[67023]_ , \new_[67026]_ ,
    \new_[67027]_ , \new_[67028]_ , \new_[67032]_ , \new_[67033]_ ,
    \new_[67036]_ , \new_[67039]_ , \new_[67040]_ , \new_[67041]_ ,
    \new_[67045]_ , \new_[67046]_ , \new_[67049]_ , \new_[67052]_ ,
    \new_[67053]_ , \new_[67054]_ , \new_[67058]_ , \new_[67059]_ ,
    \new_[67062]_ , \new_[67065]_ , \new_[67066]_ , \new_[67067]_ ,
    \new_[67071]_ , \new_[67072]_ , \new_[67075]_ , \new_[67078]_ ,
    \new_[67079]_ , \new_[67080]_ , \new_[67084]_ , \new_[67085]_ ,
    \new_[67088]_ , \new_[67091]_ , \new_[67092]_ , \new_[67093]_ ,
    \new_[67097]_ , \new_[67098]_ , \new_[67101]_ , \new_[67104]_ ,
    \new_[67105]_ , \new_[67106]_ , \new_[67110]_ , \new_[67111]_ ,
    \new_[67114]_ , \new_[67117]_ , \new_[67118]_ , \new_[67119]_ ,
    \new_[67123]_ , \new_[67124]_ , \new_[67127]_ , \new_[67130]_ ,
    \new_[67131]_ , \new_[67132]_ , \new_[67136]_ , \new_[67137]_ ,
    \new_[67140]_ , \new_[67143]_ , \new_[67144]_ , \new_[67145]_ ,
    \new_[67149]_ , \new_[67150]_ , \new_[67153]_ , \new_[67156]_ ,
    \new_[67157]_ , \new_[67158]_ , \new_[67162]_ , \new_[67163]_ ,
    \new_[67166]_ , \new_[67169]_ , \new_[67170]_ , \new_[67171]_ ,
    \new_[67175]_ , \new_[67176]_ , \new_[67179]_ , \new_[67182]_ ,
    \new_[67183]_ , \new_[67184]_ , \new_[67188]_ , \new_[67189]_ ,
    \new_[67192]_ , \new_[67195]_ , \new_[67196]_ , \new_[67197]_ ,
    \new_[67201]_ , \new_[67202]_ , \new_[67205]_ , \new_[67208]_ ,
    \new_[67209]_ , \new_[67210]_ , \new_[67214]_ , \new_[67215]_ ,
    \new_[67218]_ , \new_[67221]_ , \new_[67222]_ , \new_[67223]_ ,
    \new_[67227]_ , \new_[67228]_ , \new_[67231]_ , \new_[67234]_ ,
    \new_[67235]_ , \new_[67236]_ , \new_[67240]_ , \new_[67241]_ ,
    \new_[67244]_ , \new_[67247]_ , \new_[67248]_ , \new_[67249]_ ,
    \new_[67253]_ , \new_[67254]_ , \new_[67257]_ , \new_[67260]_ ,
    \new_[67261]_ , \new_[67262]_ , \new_[67266]_ , \new_[67267]_ ,
    \new_[67270]_ , \new_[67273]_ , \new_[67274]_ , \new_[67275]_ ,
    \new_[67279]_ , \new_[67280]_ , \new_[67283]_ , \new_[67286]_ ,
    \new_[67287]_ , \new_[67288]_ , \new_[67292]_ , \new_[67293]_ ,
    \new_[67296]_ , \new_[67299]_ , \new_[67300]_ , \new_[67301]_ ,
    \new_[67305]_ , \new_[67306]_ , \new_[67309]_ , \new_[67312]_ ,
    \new_[67313]_ , \new_[67314]_ , \new_[67318]_ , \new_[67319]_ ,
    \new_[67322]_ , \new_[67325]_ , \new_[67326]_ , \new_[67327]_ ,
    \new_[67331]_ , \new_[67332]_ , \new_[67335]_ , \new_[67338]_ ,
    \new_[67339]_ , \new_[67340]_ , \new_[67344]_ , \new_[67345]_ ,
    \new_[67348]_ , \new_[67351]_ , \new_[67352]_ , \new_[67353]_ ,
    \new_[67357]_ , \new_[67358]_ , \new_[67361]_ , \new_[67364]_ ,
    \new_[67365]_ , \new_[67366]_ , \new_[67370]_ , \new_[67371]_ ,
    \new_[67374]_ , \new_[67377]_ , \new_[67378]_ , \new_[67379]_ ,
    \new_[67383]_ , \new_[67384]_ , \new_[67387]_ , \new_[67390]_ ,
    \new_[67391]_ , \new_[67392]_ , \new_[67396]_ , \new_[67397]_ ,
    \new_[67400]_ , \new_[67403]_ , \new_[67404]_ , \new_[67405]_ ,
    \new_[67409]_ , \new_[67410]_ , \new_[67413]_ , \new_[67416]_ ,
    \new_[67417]_ , \new_[67418]_ , \new_[67422]_ , \new_[67423]_ ,
    \new_[67426]_ , \new_[67429]_ , \new_[67430]_ , \new_[67431]_ ,
    \new_[67435]_ , \new_[67436]_ , \new_[67439]_ , \new_[67442]_ ,
    \new_[67443]_ , \new_[67444]_ , \new_[67448]_ , \new_[67449]_ ,
    \new_[67452]_ , \new_[67455]_ , \new_[67456]_ , \new_[67457]_ ,
    \new_[67461]_ , \new_[67462]_ , \new_[67465]_ , \new_[67468]_ ,
    \new_[67469]_ , \new_[67470]_ , \new_[67474]_ , \new_[67475]_ ,
    \new_[67478]_ , \new_[67481]_ , \new_[67482]_ , \new_[67483]_ ,
    \new_[67487]_ , \new_[67488]_ , \new_[67491]_ , \new_[67494]_ ,
    \new_[67495]_ , \new_[67496]_ , \new_[67500]_ , \new_[67501]_ ,
    \new_[67504]_ , \new_[67507]_ , \new_[67508]_ , \new_[67509]_ ,
    \new_[67513]_ , \new_[67514]_ , \new_[67517]_ , \new_[67520]_ ,
    \new_[67521]_ , \new_[67522]_ , \new_[67526]_ , \new_[67527]_ ,
    \new_[67530]_ , \new_[67533]_ , \new_[67534]_ , \new_[67535]_ ,
    \new_[67539]_ , \new_[67540]_ , \new_[67543]_ , \new_[67546]_ ,
    \new_[67547]_ , \new_[67548]_ , \new_[67552]_ , \new_[67553]_ ,
    \new_[67556]_ , \new_[67559]_ , \new_[67560]_ , \new_[67561]_ ,
    \new_[67565]_ , \new_[67566]_ , \new_[67569]_ , \new_[67572]_ ,
    \new_[67573]_ , \new_[67574]_ , \new_[67578]_ , \new_[67579]_ ,
    \new_[67582]_ , \new_[67585]_ , \new_[67586]_ , \new_[67587]_ ,
    \new_[67591]_ , \new_[67592]_ , \new_[67595]_ , \new_[67598]_ ,
    \new_[67599]_ , \new_[67600]_ , \new_[67604]_ , \new_[67605]_ ,
    \new_[67608]_ , \new_[67611]_ , \new_[67612]_ , \new_[67613]_ ,
    \new_[67617]_ , \new_[67618]_ , \new_[67621]_ , \new_[67624]_ ,
    \new_[67625]_ , \new_[67626]_ , \new_[67630]_ , \new_[67631]_ ,
    \new_[67634]_ , \new_[67637]_ , \new_[67638]_ , \new_[67639]_ ,
    \new_[67643]_ , \new_[67644]_ , \new_[67647]_ , \new_[67650]_ ,
    \new_[67651]_ , \new_[67652]_ , \new_[67656]_ , \new_[67657]_ ,
    \new_[67660]_ , \new_[67663]_ , \new_[67664]_ , \new_[67665]_ ,
    \new_[67669]_ , \new_[67670]_ , \new_[67673]_ , \new_[67676]_ ,
    \new_[67677]_ , \new_[67678]_ , \new_[67682]_ , \new_[67683]_ ,
    \new_[67686]_ , \new_[67689]_ , \new_[67690]_ , \new_[67691]_ ,
    \new_[67695]_ , \new_[67696]_ , \new_[67699]_ , \new_[67702]_ ,
    \new_[67703]_ , \new_[67704]_ , \new_[67708]_ , \new_[67709]_ ,
    \new_[67712]_ , \new_[67715]_ , \new_[67716]_ , \new_[67717]_ ,
    \new_[67721]_ , \new_[67722]_ , \new_[67725]_ , \new_[67728]_ ,
    \new_[67729]_ , \new_[67730]_ , \new_[67734]_ , \new_[67735]_ ,
    \new_[67738]_ , \new_[67741]_ , \new_[67742]_ , \new_[67743]_ ,
    \new_[67747]_ , \new_[67748]_ , \new_[67751]_ , \new_[67754]_ ,
    \new_[67755]_ , \new_[67756]_ , \new_[67760]_ , \new_[67761]_ ,
    \new_[67764]_ , \new_[67767]_ , \new_[67768]_ , \new_[67769]_ ,
    \new_[67773]_ , \new_[67774]_ , \new_[67777]_ , \new_[67780]_ ,
    \new_[67781]_ , \new_[67782]_ , \new_[67786]_ , \new_[67787]_ ,
    \new_[67790]_ , \new_[67793]_ , \new_[67794]_ , \new_[67795]_ ,
    \new_[67799]_ , \new_[67800]_ , \new_[67803]_ , \new_[67806]_ ,
    \new_[67807]_ , \new_[67808]_ , \new_[67812]_ , \new_[67813]_ ,
    \new_[67816]_ , \new_[67819]_ , \new_[67820]_ , \new_[67821]_ ,
    \new_[67825]_ , \new_[67826]_ , \new_[67829]_ , \new_[67832]_ ,
    \new_[67833]_ , \new_[67834]_ , \new_[67838]_ , \new_[67839]_ ,
    \new_[67842]_ , \new_[67845]_ , \new_[67846]_ , \new_[67847]_ ,
    \new_[67851]_ , \new_[67852]_ , \new_[67855]_ , \new_[67858]_ ,
    \new_[67859]_ , \new_[67860]_ , \new_[67864]_ , \new_[67865]_ ,
    \new_[67868]_ , \new_[67871]_ , \new_[67872]_ , \new_[67873]_ ,
    \new_[67877]_ , \new_[67878]_ , \new_[67881]_ , \new_[67884]_ ,
    \new_[67885]_ , \new_[67886]_ , \new_[67890]_ , \new_[67891]_ ,
    \new_[67894]_ , \new_[67897]_ , \new_[67898]_ , \new_[67899]_ ,
    \new_[67903]_ , \new_[67904]_ , \new_[67907]_ , \new_[67910]_ ,
    \new_[67911]_ , \new_[67912]_ , \new_[67916]_ , \new_[67917]_ ,
    \new_[67920]_ , \new_[67923]_ , \new_[67924]_ , \new_[67925]_ ,
    \new_[67929]_ , \new_[67930]_ , \new_[67933]_ , \new_[67936]_ ,
    \new_[67937]_ , \new_[67938]_ , \new_[67942]_ , \new_[67943]_ ,
    \new_[67946]_ , \new_[67949]_ , \new_[67950]_ , \new_[67951]_ ,
    \new_[67955]_ , \new_[67956]_ , \new_[67959]_ , \new_[67962]_ ,
    \new_[67963]_ , \new_[67964]_ , \new_[67968]_ , \new_[67969]_ ,
    \new_[67972]_ , \new_[67975]_ , \new_[67976]_ , \new_[67977]_ ,
    \new_[67981]_ , \new_[67982]_ , \new_[67985]_ , \new_[67988]_ ,
    \new_[67989]_ , \new_[67990]_ , \new_[67994]_ , \new_[67995]_ ,
    \new_[67998]_ , \new_[68001]_ , \new_[68002]_ , \new_[68003]_ ,
    \new_[68007]_ , \new_[68008]_ , \new_[68011]_ , \new_[68014]_ ,
    \new_[68015]_ , \new_[68016]_ , \new_[68020]_ , \new_[68021]_ ,
    \new_[68024]_ , \new_[68027]_ , \new_[68028]_ , \new_[68029]_ ,
    \new_[68033]_ , \new_[68034]_ , \new_[68037]_ , \new_[68040]_ ,
    \new_[68041]_ , \new_[68042]_ , \new_[68046]_ , \new_[68047]_ ,
    \new_[68050]_ , \new_[68053]_ , \new_[68054]_ , \new_[68055]_ ,
    \new_[68059]_ , \new_[68060]_ , \new_[68063]_ , \new_[68066]_ ,
    \new_[68067]_ , \new_[68068]_ , \new_[68072]_ , \new_[68073]_ ,
    \new_[68076]_ , \new_[68079]_ , \new_[68080]_ , \new_[68081]_ ,
    \new_[68085]_ , \new_[68086]_ , \new_[68089]_ , \new_[68092]_ ,
    \new_[68093]_ , \new_[68094]_ , \new_[68098]_ , \new_[68099]_ ,
    \new_[68102]_ , \new_[68105]_ , \new_[68106]_ , \new_[68107]_ ,
    \new_[68111]_ , \new_[68112]_ , \new_[68115]_ , \new_[68118]_ ,
    \new_[68119]_ , \new_[68120]_ , \new_[68124]_ , \new_[68125]_ ,
    \new_[68128]_ , \new_[68131]_ , \new_[68132]_ , \new_[68133]_ ,
    \new_[68137]_ , \new_[68138]_ , \new_[68141]_ , \new_[68144]_ ,
    \new_[68145]_ , \new_[68146]_ , \new_[68150]_ , \new_[68151]_ ,
    \new_[68154]_ , \new_[68157]_ , \new_[68158]_ , \new_[68159]_ ,
    \new_[68163]_ , \new_[68164]_ , \new_[68167]_ , \new_[68170]_ ,
    \new_[68171]_ , \new_[68172]_ , \new_[68176]_ , \new_[68177]_ ,
    \new_[68180]_ , \new_[68183]_ , \new_[68184]_ , \new_[68185]_ ,
    \new_[68189]_ , \new_[68190]_ , \new_[68193]_ , \new_[68196]_ ,
    \new_[68197]_ , \new_[68198]_ , \new_[68202]_ , \new_[68203]_ ,
    \new_[68206]_ , \new_[68209]_ , \new_[68210]_ , \new_[68211]_ ,
    \new_[68215]_ , \new_[68216]_ , \new_[68219]_ , \new_[68222]_ ,
    \new_[68223]_ , \new_[68224]_ , \new_[68228]_ , \new_[68229]_ ,
    \new_[68232]_ , \new_[68235]_ , \new_[68236]_ , \new_[68237]_ ,
    \new_[68241]_ , \new_[68242]_ , \new_[68245]_ , \new_[68248]_ ,
    \new_[68249]_ , \new_[68250]_ , \new_[68254]_ , \new_[68255]_ ,
    \new_[68258]_ , \new_[68261]_ , \new_[68262]_ , \new_[68263]_ ,
    \new_[68267]_ , \new_[68268]_ , \new_[68271]_ , \new_[68274]_ ,
    \new_[68275]_ , \new_[68276]_ , \new_[68280]_ , \new_[68281]_ ,
    \new_[68284]_ , \new_[68287]_ , \new_[68288]_ , \new_[68289]_ ,
    \new_[68293]_ , \new_[68294]_ , \new_[68297]_ , \new_[68300]_ ,
    \new_[68301]_ , \new_[68302]_ , \new_[68306]_ , \new_[68307]_ ,
    \new_[68310]_ , \new_[68313]_ , \new_[68314]_ , \new_[68315]_ ,
    \new_[68319]_ , \new_[68320]_ , \new_[68323]_ , \new_[68326]_ ,
    \new_[68327]_ , \new_[68328]_ , \new_[68332]_ , \new_[68333]_ ,
    \new_[68336]_ , \new_[68339]_ , \new_[68340]_ , \new_[68341]_ ,
    \new_[68345]_ , \new_[68346]_ , \new_[68349]_ , \new_[68352]_ ,
    \new_[68353]_ , \new_[68354]_ , \new_[68358]_ , \new_[68359]_ ,
    \new_[68362]_ , \new_[68365]_ , \new_[68366]_ , \new_[68367]_ ,
    \new_[68371]_ , \new_[68372]_ , \new_[68375]_ , \new_[68378]_ ,
    \new_[68379]_ , \new_[68380]_ , \new_[68384]_ , \new_[68385]_ ,
    \new_[68388]_ , \new_[68391]_ , \new_[68392]_ , \new_[68393]_ ,
    \new_[68397]_ , \new_[68398]_ , \new_[68401]_ , \new_[68404]_ ,
    \new_[68405]_ , \new_[68406]_ , \new_[68410]_ , \new_[68411]_ ,
    \new_[68414]_ , \new_[68417]_ , \new_[68418]_ , \new_[68419]_ ,
    \new_[68423]_ , \new_[68424]_ , \new_[68427]_ , \new_[68430]_ ,
    \new_[68431]_ , \new_[68432]_ , \new_[68436]_ , \new_[68437]_ ,
    \new_[68440]_ , \new_[68443]_ , \new_[68444]_ , \new_[68445]_ ,
    \new_[68449]_ , \new_[68450]_ , \new_[68453]_ , \new_[68456]_ ,
    \new_[68457]_ , \new_[68458]_ , \new_[68462]_ , \new_[68463]_ ,
    \new_[68466]_ , \new_[68469]_ , \new_[68470]_ , \new_[68471]_ ,
    \new_[68475]_ , \new_[68476]_ , \new_[68479]_ , \new_[68482]_ ,
    \new_[68483]_ , \new_[68484]_ , \new_[68488]_ , \new_[68489]_ ,
    \new_[68492]_ , \new_[68495]_ , \new_[68496]_ , \new_[68497]_ ,
    \new_[68501]_ , \new_[68502]_ , \new_[68505]_ , \new_[68508]_ ,
    \new_[68509]_ , \new_[68510]_ , \new_[68514]_ , \new_[68515]_ ,
    \new_[68518]_ , \new_[68521]_ , \new_[68522]_ , \new_[68523]_ ,
    \new_[68527]_ , \new_[68528]_ , \new_[68531]_ , \new_[68534]_ ,
    \new_[68535]_ , \new_[68536]_ , \new_[68540]_ , \new_[68541]_ ,
    \new_[68544]_ , \new_[68547]_ , \new_[68548]_ , \new_[68549]_ ,
    \new_[68553]_ , \new_[68554]_ , \new_[68557]_ , \new_[68560]_ ,
    \new_[68561]_ , \new_[68562]_ , \new_[68566]_ , \new_[68567]_ ,
    \new_[68570]_ , \new_[68573]_ , \new_[68574]_ , \new_[68575]_ ,
    \new_[68579]_ , \new_[68580]_ , \new_[68583]_ , \new_[68586]_ ,
    \new_[68587]_ , \new_[68588]_ , \new_[68592]_ , \new_[68593]_ ,
    \new_[68596]_ , \new_[68599]_ , \new_[68600]_ , \new_[68601]_ ,
    \new_[68605]_ , \new_[68606]_ , \new_[68609]_ , \new_[68612]_ ,
    \new_[68613]_ , \new_[68614]_ , \new_[68618]_ , \new_[68619]_ ,
    \new_[68622]_ , \new_[68625]_ , \new_[68626]_ , \new_[68627]_ ,
    \new_[68631]_ , \new_[68632]_ , \new_[68635]_ , \new_[68638]_ ,
    \new_[68639]_ , \new_[68640]_ , \new_[68644]_ , \new_[68645]_ ,
    \new_[68648]_ , \new_[68651]_ , \new_[68652]_ , \new_[68653]_ ,
    \new_[68657]_ , \new_[68658]_ , \new_[68661]_ , \new_[68664]_ ,
    \new_[68665]_ , \new_[68666]_ , \new_[68670]_ , \new_[68671]_ ,
    \new_[68674]_ , \new_[68677]_ , \new_[68678]_ , \new_[68679]_ ,
    \new_[68683]_ , \new_[68684]_ , \new_[68687]_ , \new_[68690]_ ,
    \new_[68691]_ , \new_[68692]_ , \new_[68696]_ , \new_[68697]_ ,
    \new_[68700]_ , \new_[68703]_ , \new_[68704]_ , \new_[68705]_ ,
    \new_[68709]_ , \new_[68710]_ , \new_[68713]_ , \new_[68716]_ ,
    \new_[68717]_ , \new_[68718]_ , \new_[68722]_ , \new_[68723]_ ,
    \new_[68726]_ , \new_[68729]_ , \new_[68730]_ , \new_[68731]_ ,
    \new_[68735]_ , \new_[68736]_ , \new_[68739]_ , \new_[68742]_ ,
    \new_[68743]_ , \new_[68744]_ , \new_[68748]_ , \new_[68749]_ ,
    \new_[68752]_ , \new_[68755]_ , \new_[68756]_ , \new_[68757]_ ,
    \new_[68761]_ , \new_[68762]_ , \new_[68765]_ , \new_[68768]_ ,
    \new_[68769]_ , \new_[68770]_ , \new_[68774]_ , \new_[68775]_ ,
    \new_[68778]_ , \new_[68781]_ , \new_[68782]_ , \new_[68783]_ ,
    \new_[68787]_ , \new_[68788]_ , \new_[68791]_ , \new_[68794]_ ,
    \new_[68795]_ , \new_[68796]_ , \new_[68800]_ , \new_[68801]_ ,
    \new_[68804]_ , \new_[68807]_ , \new_[68808]_ , \new_[68809]_ ,
    \new_[68813]_ , \new_[68814]_ , \new_[68817]_ , \new_[68820]_ ,
    \new_[68821]_ , \new_[68822]_ , \new_[68826]_ , \new_[68827]_ ,
    \new_[68830]_ , \new_[68833]_ , \new_[68834]_ , \new_[68835]_ ,
    \new_[68839]_ , \new_[68840]_ , \new_[68843]_ , \new_[68846]_ ,
    \new_[68847]_ , \new_[68848]_ , \new_[68852]_ , \new_[68853]_ ,
    \new_[68856]_ , \new_[68859]_ , \new_[68860]_ , \new_[68861]_ ,
    \new_[68865]_ , \new_[68866]_ , \new_[68869]_ , \new_[68872]_ ,
    \new_[68873]_ , \new_[68874]_ , \new_[68878]_ , \new_[68879]_ ,
    \new_[68882]_ , \new_[68885]_ , \new_[68886]_ , \new_[68887]_ ,
    \new_[68891]_ , \new_[68892]_ , \new_[68895]_ , \new_[68898]_ ,
    \new_[68899]_ , \new_[68900]_ , \new_[68904]_ , \new_[68905]_ ,
    \new_[68908]_ , \new_[68911]_ , \new_[68912]_ , \new_[68913]_ ,
    \new_[68917]_ , \new_[68918]_ , \new_[68921]_ , \new_[68924]_ ,
    \new_[68925]_ , \new_[68926]_ , \new_[68930]_ , \new_[68931]_ ,
    \new_[68934]_ , \new_[68937]_ , \new_[68938]_ , \new_[68939]_ ,
    \new_[68943]_ , \new_[68944]_ , \new_[68947]_ , \new_[68950]_ ,
    \new_[68951]_ , \new_[68952]_ , \new_[68956]_ , \new_[68957]_ ,
    \new_[68960]_ , \new_[68963]_ , \new_[68964]_ , \new_[68965]_ ,
    \new_[68969]_ , \new_[68970]_ , \new_[68973]_ , \new_[68976]_ ,
    \new_[68977]_ , \new_[68978]_ , \new_[68982]_ , \new_[68983]_ ,
    \new_[68986]_ , \new_[68989]_ , \new_[68990]_ , \new_[68991]_ ,
    \new_[68995]_ , \new_[68996]_ , \new_[68999]_ , \new_[69002]_ ,
    \new_[69003]_ , \new_[69004]_ , \new_[69008]_ , \new_[69009]_ ,
    \new_[69012]_ , \new_[69015]_ , \new_[69016]_ , \new_[69017]_ ,
    \new_[69021]_ , \new_[69022]_ , \new_[69025]_ , \new_[69028]_ ,
    \new_[69029]_ , \new_[69030]_ , \new_[69034]_ , \new_[69035]_ ,
    \new_[69038]_ , \new_[69041]_ , \new_[69042]_ , \new_[69043]_ ,
    \new_[69047]_ , \new_[69048]_ , \new_[69051]_ , \new_[69054]_ ,
    \new_[69055]_ , \new_[69056]_ , \new_[69060]_ , \new_[69061]_ ,
    \new_[69064]_ , \new_[69067]_ , \new_[69068]_ , \new_[69069]_ ,
    \new_[69073]_ , \new_[69074]_ , \new_[69077]_ , \new_[69080]_ ,
    \new_[69081]_ , \new_[69082]_ , \new_[69086]_ , \new_[69087]_ ,
    \new_[69090]_ , \new_[69093]_ , \new_[69094]_ , \new_[69095]_ ,
    \new_[69099]_ , \new_[69100]_ , \new_[69103]_ , \new_[69106]_ ,
    \new_[69107]_ , \new_[69108]_ , \new_[69112]_ , \new_[69113]_ ,
    \new_[69116]_ , \new_[69119]_ , \new_[69120]_ , \new_[69121]_ ,
    \new_[69125]_ , \new_[69126]_ , \new_[69129]_ , \new_[69132]_ ,
    \new_[69133]_ , \new_[69134]_ , \new_[69138]_ , \new_[69139]_ ,
    \new_[69142]_ , \new_[69145]_ , \new_[69146]_ , \new_[69147]_ ,
    \new_[69151]_ , \new_[69152]_ , \new_[69155]_ , \new_[69158]_ ,
    \new_[69159]_ , \new_[69160]_ , \new_[69164]_ , \new_[69165]_ ,
    \new_[69168]_ , \new_[69171]_ , \new_[69172]_ , \new_[69173]_ ,
    \new_[69177]_ , \new_[69178]_ , \new_[69181]_ , \new_[69184]_ ,
    \new_[69185]_ , \new_[69186]_ , \new_[69190]_ , \new_[69191]_ ,
    \new_[69194]_ , \new_[69197]_ , \new_[69198]_ , \new_[69199]_ ,
    \new_[69203]_ , \new_[69204]_ , \new_[69207]_ , \new_[69210]_ ,
    \new_[69211]_ , \new_[69212]_ , \new_[69216]_ , \new_[69217]_ ,
    \new_[69220]_ , \new_[69223]_ , \new_[69224]_ , \new_[69225]_ ,
    \new_[69229]_ , \new_[69230]_ , \new_[69233]_ , \new_[69236]_ ,
    \new_[69237]_ , \new_[69238]_ , \new_[69242]_ , \new_[69243]_ ,
    \new_[69246]_ , \new_[69249]_ , \new_[69250]_ , \new_[69251]_ ,
    \new_[69255]_ , \new_[69256]_ , \new_[69259]_ , \new_[69262]_ ,
    \new_[69263]_ , \new_[69264]_ , \new_[69268]_ , \new_[69269]_ ,
    \new_[69272]_ , \new_[69275]_ , \new_[69276]_ , \new_[69277]_ ,
    \new_[69281]_ , \new_[69282]_ , \new_[69285]_ , \new_[69288]_ ,
    \new_[69289]_ , \new_[69290]_ , \new_[69294]_ , \new_[69295]_ ,
    \new_[69298]_ , \new_[69301]_ , \new_[69302]_ , \new_[69303]_ ,
    \new_[69307]_ , \new_[69308]_ , \new_[69311]_ , \new_[69314]_ ,
    \new_[69315]_ , \new_[69316]_ , \new_[69320]_ , \new_[69321]_ ,
    \new_[69324]_ , \new_[69327]_ , \new_[69328]_ , \new_[69329]_ ,
    \new_[69333]_ , \new_[69334]_ , \new_[69337]_ , \new_[69340]_ ,
    \new_[69341]_ , \new_[69342]_ , \new_[69346]_ , \new_[69347]_ ,
    \new_[69350]_ , \new_[69353]_ , \new_[69354]_ , \new_[69355]_ ,
    \new_[69359]_ , \new_[69360]_ , \new_[69363]_ , \new_[69366]_ ,
    \new_[69367]_ , \new_[69368]_ , \new_[69372]_ , \new_[69373]_ ,
    \new_[69376]_ , \new_[69379]_ , \new_[69380]_ , \new_[69381]_ ,
    \new_[69385]_ , \new_[69386]_ , \new_[69389]_ , \new_[69392]_ ,
    \new_[69393]_ , \new_[69394]_ , \new_[69398]_ , \new_[69399]_ ,
    \new_[69402]_ , \new_[69405]_ , \new_[69406]_ , \new_[69407]_ ,
    \new_[69411]_ , \new_[69412]_ , \new_[69415]_ , \new_[69418]_ ,
    \new_[69419]_ , \new_[69420]_ , \new_[69424]_ , \new_[69425]_ ,
    \new_[69428]_ , \new_[69431]_ , \new_[69432]_ , \new_[69433]_ ,
    \new_[69437]_ , \new_[69438]_ , \new_[69441]_ , \new_[69444]_ ,
    \new_[69445]_ , \new_[69446]_ , \new_[69450]_ , \new_[69451]_ ,
    \new_[69454]_ , \new_[69457]_ , \new_[69458]_ , \new_[69459]_ ,
    \new_[69463]_ , \new_[69464]_ , \new_[69467]_ , \new_[69470]_ ,
    \new_[69471]_ , \new_[69472]_ , \new_[69476]_ , \new_[69477]_ ,
    \new_[69480]_ , \new_[69483]_ , \new_[69484]_ , \new_[69485]_ ,
    \new_[69489]_ , \new_[69490]_ , \new_[69493]_ , \new_[69496]_ ,
    \new_[69497]_ , \new_[69498]_ , \new_[69502]_ , \new_[69503]_ ,
    \new_[69506]_ , \new_[69509]_ , \new_[69510]_ , \new_[69511]_ ,
    \new_[69515]_ , \new_[69516]_ , \new_[69519]_ , \new_[69522]_ ,
    \new_[69523]_ , \new_[69524]_ , \new_[69528]_ , \new_[69529]_ ,
    \new_[69532]_ , \new_[69535]_ , \new_[69536]_ , \new_[69537]_ ,
    \new_[69541]_ , \new_[69542]_ , \new_[69545]_ , \new_[69548]_ ,
    \new_[69549]_ , \new_[69550]_ , \new_[69554]_ , \new_[69555]_ ,
    \new_[69558]_ , \new_[69561]_ , \new_[69562]_ , \new_[69563]_ ,
    \new_[69567]_ , \new_[69568]_ , \new_[69571]_ , \new_[69574]_ ,
    \new_[69575]_ , \new_[69576]_ , \new_[69580]_ , \new_[69581]_ ,
    \new_[69584]_ , \new_[69587]_ , \new_[69588]_ , \new_[69589]_ ,
    \new_[69593]_ , \new_[69594]_ , \new_[69597]_ , \new_[69600]_ ,
    \new_[69601]_ , \new_[69602]_ , \new_[69606]_ , \new_[69607]_ ,
    \new_[69610]_ , \new_[69613]_ , \new_[69614]_ , \new_[69615]_ ,
    \new_[69619]_ , \new_[69620]_ , \new_[69623]_ , \new_[69626]_ ,
    \new_[69627]_ , \new_[69628]_ , \new_[69632]_ , \new_[69633]_ ,
    \new_[69636]_ , \new_[69639]_ , \new_[69640]_ , \new_[69641]_ ,
    \new_[69645]_ , \new_[69646]_ , \new_[69649]_ , \new_[69652]_ ,
    \new_[69653]_ , \new_[69654]_ , \new_[69658]_ , \new_[69659]_ ,
    \new_[69662]_ , \new_[69665]_ , \new_[69666]_ , \new_[69667]_ ,
    \new_[69671]_ , \new_[69672]_ , \new_[69675]_ , \new_[69678]_ ,
    \new_[69679]_ , \new_[69680]_ , \new_[69684]_ , \new_[69685]_ ,
    \new_[69688]_ , \new_[69691]_ , \new_[69692]_ , \new_[69693]_ ,
    \new_[69697]_ , \new_[69698]_ , \new_[69701]_ , \new_[69704]_ ,
    \new_[69705]_ , \new_[69706]_ , \new_[69710]_ , \new_[69711]_ ,
    \new_[69714]_ , \new_[69717]_ , \new_[69718]_ , \new_[69719]_ ,
    \new_[69723]_ , \new_[69724]_ , \new_[69727]_ , \new_[69730]_ ,
    \new_[69731]_ , \new_[69732]_ , \new_[69736]_ , \new_[69737]_ ,
    \new_[69740]_ , \new_[69743]_ , \new_[69744]_ , \new_[69745]_ ,
    \new_[69749]_ , \new_[69750]_ , \new_[69753]_ , \new_[69756]_ ,
    \new_[69757]_ , \new_[69758]_ , \new_[69762]_ , \new_[69763]_ ,
    \new_[69766]_ , \new_[69769]_ , \new_[69770]_ , \new_[69771]_ ,
    \new_[69775]_ , \new_[69776]_ , \new_[69779]_ , \new_[69782]_ ,
    \new_[69783]_ , \new_[69784]_ , \new_[69788]_ , \new_[69789]_ ,
    \new_[69792]_ , \new_[69795]_ , \new_[69796]_ , \new_[69797]_ ,
    \new_[69801]_ , \new_[69802]_ , \new_[69805]_ , \new_[69808]_ ,
    \new_[69809]_ , \new_[69810]_ , \new_[69814]_ , \new_[69815]_ ,
    \new_[69818]_ , \new_[69821]_ , \new_[69822]_ , \new_[69823]_ ,
    \new_[69827]_ , \new_[69828]_ , \new_[69831]_ , \new_[69834]_ ,
    \new_[69835]_ , \new_[69836]_ , \new_[69840]_ , \new_[69841]_ ,
    \new_[69844]_ , \new_[69847]_ , \new_[69848]_ , \new_[69849]_ ,
    \new_[69853]_ , \new_[69854]_ , \new_[69857]_ , \new_[69860]_ ,
    \new_[69861]_ , \new_[69862]_ , \new_[69866]_ , \new_[69867]_ ,
    \new_[69870]_ , \new_[69873]_ , \new_[69874]_ , \new_[69875]_ ,
    \new_[69879]_ , \new_[69880]_ , \new_[69883]_ , \new_[69886]_ ,
    \new_[69887]_ , \new_[69888]_ , \new_[69892]_ , \new_[69893]_ ,
    \new_[69896]_ , \new_[69899]_ , \new_[69900]_ , \new_[69901]_ ,
    \new_[69905]_ , \new_[69906]_ , \new_[69909]_ , \new_[69912]_ ,
    \new_[69913]_ , \new_[69914]_ , \new_[69918]_ , \new_[69919]_ ,
    \new_[69922]_ , \new_[69925]_ , \new_[69926]_ , \new_[69927]_ ,
    \new_[69931]_ , \new_[69932]_ , \new_[69935]_ , \new_[69938]_ ,
    \new_[69939]_ , \new_[69940]_ , \new_[69944]_ , \new_[69945]_ ,
    \new_[69948]_ , \new_[69951]_ , \new_[69952]_ , \new_[69953]_ ,
    \new_[69957]_ , \new_[69958]_ , \new_[69961]_ , \new_[69964]_ ,
    \new_[69965]_ , \new_[69966]_ , \new_[69970]_ , \new_[69971]_ ,
    \new_[69974]_ , \new_[69977]_ , \new_[69978]_ , \new_[69979]_ ,
    \new_[69983]_ , \new_[69984]_ , \new_[69987]_ , \new_[69990]_ ,
    \new_[69991]_ , \new_[69992]_ , \new_[69996]_ , \new_[69997]_ ,
    \new_[70000]_ , \new_[70003]_ , \new_[70004]_ , \new_[70005]_ ,
    \new_[70009]_ , \new_[70010]_ , \new_[70013]_ , \new_[70016]_ ,
    \new_[70017]_ , \new_[70018]_ , \new_[70022]_ , \new_[70023]_ ,
    \new_[70026]_ , \new_[70029]_ , \new_[70030]_ , \new_[70031]_ ,
    \new_[70035]_ , \new_[70036]_ , \new_[70039]_ , \new_[70042]_ ,
    \new_[70043]_ , \new_[70044]_ , \new_[70048]_ , \new_[70049]_ ,
    \new_[70052]_ , \new_[70055]_ , \new_[70056]_ , \new_[70057]_ ,
    \new_[70061]_ , \new_[70062]_ , \new_[70065]_ , \new_[70068]_ ,
    \new_[70069]_ , \new_[70070]_ , \new_[70074]_ , \new_[70075]_ ,
    \new_[70078]_ , \new_[70081]_ , \new_[70082]_ , \new_[70083]_ ,
    \new_[70087]_ , \new_[70088]_ , \new_[70091]_ , \new_[70094]_ ,
    \new_[70095]_ , \new_[70096]_ , \new_[70100]_ , \new_[70101]_ ,
    \new_[70104]_ , \new_[70107]_ , \new_[70108]_ , \new_[70109]_ ,
    \new_[70113]_ , \new_[70114]_ , \new_[70117]_ , \new_[70120]_ ,
    \new_[70121]_ , \new_[70122]_ , \new_[70126]_ , \new_[70127]_ ,
    \new_[70130]_ , \new_[70133]_ , \new_[70134]_ , \new_[70135]_ ,
    \new_[70139]_ , \new_[70140]_ , \new_[70143]_ , \new_[70146]_ ,
    \new_[70147]_ , \new_[70148]_ , \new_[70152]_ , \new_[70153]_ ,
    \new_[70156]_ , \new_[70159]_ , \new_[70160]_ , \new_[70161]_ ,
    \new_[70165]_ , \new_[70166]_ , \new_[70169]_ , \new_[70172]_ ,
    \new_[70173]_ , \new_[70174]_ , \new_[70178]_ , \new_[70179]_ ,
    \new_[70182]_ , \new_[70185]_ , \new_[70186]_ , \new_[70187]_ ,
    \new_[70191]_ , \new_[70192]_ , \new_[70195]_ , \new_[70198]_ ,
    \new_[70199]_ , \new_[70200]_ , \new_[70204]_ , \new_[70205]_ ,
    \new_[70208]_ , \new_[70211]_ , \new_[70212]_ , \new_[70213]_ ,
    \new_[70217]_ , \new_[70218]_ , \new_[70221]_ , \new_[70224]_ ,
    \new_[70225]_ , \new_[70226]_ , \new_[70230]_ , \new_[70231]_ ,
    \new_[70234]_ , \new_[70237]_ , \new_[70238]_ , \new_[70239]_ ,
    \new_[70243]_ , \new_[70244]_ , \new_[70247]_ , \new_[70250]_ ,
    \new_[70251]_ , \new_[70252]_ , \new_[70256]_ , \new_[70257]_ ,
    \new_[70260]_ , \new_[70263]_ , \new_[70264]_ , \new_[70265]_ ,
    \new_[70269]_ , \new_[70270]_ , \new_[70273]_ , \new_[70276]_ ,
    \new_[70277]_ , \new_[70278]_ , \new_[70282]_ , \new_[70283]_ ,
    \new_[70286]_ , \new_[70289]_ , \new_[70290]_ , \new_[70291]_ ,
    \new_[70295]_ , \new_[70296]_ , \new_[70299]_ , \new_[70302]_ ,
    \new_[70303]_ , \new_[70304]_ , \new_[70308]_ , \new_[70309]_ ,
    \new_[70312]_ , \new_[70315]_ , \new_[70316]_ , \new_[70317]_ ,
    \new_[70321]_ , \new_[70322]_ , \new_[70325]_ , \new_[70328]_ ,
    \new_[70329]_ , \new_[70330]_ , \new_[70334]_ , \new_[70335]_ ,
    \new_[70338]_ , \new_[70341]_ , \new_[70342]_ , \new_[70343]_ ,
    \new_[70347]_ , \new_[70348]_ , \new_[70351]_ , \new_[70354]_ ,
    \new_[70355]_ , \new_[70356]_ , \new_[70360]_ , \new_[70361]_ ,
    \new_[70364]_ , \new_[70367]_ , \new_[70368]_ , \new_[70369]_ ,
    \new_[70373]_ , \new_[70374]_ , \new_[70377]_ , \new_[70380]_ ,
    \new_[70381]_ , \new_[70382]_ , \new_[70386]_ , \new_[70387]_ ,
    \new_[70390]_ , \new_[70393]_ , \new_[70394]_ , \new_[70395]_ ,
    \new_[70399]_ , \new_[70400]_ , \new_[70403]_ , \new_[70406]_ ,
    \new_[70407]_ , \new_[70408]_ , \new_[70412]_ , \new_[70413]_ ,
    \new_[70416]_ , \new_[70419]_ , \new_[70420]_ , \new_[70421]_ ,
    \new_[70425]_ , \new_[70426]_ , \new_[70429]_ , \new_[70432]_ ,
    \new_[70433]_ , \new_[70434]_ , \new_[70438]_ , \new_[70439]_ ,
    \new_[70442]_ , \new_[70445]_ , \new_[70446]_ , \new_[70447]_ ,
    \new_[70451]_ , \new_[70452]_ , \new_[70455]_ , \new_[70458]_ ,
    \new_[70459]_ , \new_[70460]_ , \new_[70464]_ , \new_[70465]_ ,
    \new_[70468]_ , \new_[70471]_ , \new_[70472]_ , \new_[70473]_ ,
    \new_[70477]_ , \new_[70478]_ , \new_[70481]_ , \new_[70484]_ ,
    \new_[70485]_ , \new_[70486]_ , \new_[70490]_ , \new_[70491]_ ,
    \new_[70494]_ , \new_[70497]_ , \new_[70498]_ , \new_[70499]_ ,
    \new_[70503]_ , \new_[70504]_ , \new_[70507]_ , \new_[70510]_ ,
    \new_[70511]_ , \new_[70512]_ , \new_[70516]_ , \new_[70517]_ ,
    \new_[70520]_ , \new_[70523]_ , \new_[70524]_ , \new_[70525]_ ,
    \new_[70529]_ , \new_[70530]_ , \new_[70533]_ , \new_[70536]_ ,
    \new_[70537]_ , \new_[70538]_ , \new_[70542]_ , \new_[70543]_ ,
    \new_[70546]_ , \new_[70549]_ , \new_[70550]_ , \new_[70551]_ ,
    \new_[70555]_ , \new_[70556]_ , \new_[70559]_ , \new_[70562]_ ,
    \new_[70563]_ , \new_[70564]_ , \new_[70568]_ , \new_[70569]_ ,
    \new_[70572]_ , \new_[70575]_ , \new_[70576]_ , \new_[70577]_ ,
    \new_[70581]_ , \new_[70582]_ , \new_[70585]_ , \new_[70588]_ ,
    \new_[70589]_ , \new_[70590]_ , \new_[70594]_ , \new_[70595]_ ,
    \new_[70598]_ , \new_[70601]_ , \new_[70602]_ , \new_[70603]_ ,
    \new_[70607]_ , \new_[70608]_ , \new_[70611]_ , \new_[70614]_ ,
    \new_[70615]_ , \new_[70616]_ , \new_[70620]_ , \new_[70621]_ ,
    \new_[70624]_ , \new_[70627]_ , \new_[70628]_ , \new_[70629]_ ,
    \new_[70633]_ , \new_[70634]_ , \new_[70637]_ , \new_[70640]_ ,
    \new_[70641]_ , \new_[70642]_ , \new_[70646]_ , \new_[70647]_ ,
    \new_[70650]_ , \new_[70653]_ , \new_[70654]_ , \new_[70655]_ ,
    \new_[70659]_ , \new_[70660]_ , \new_[70663]_ , \new_[70666]_ ,
    \new_[70667]_ , \new_[70668]_ , \new_[70672]_ , \new_[70673]_ ,
    \new_[70676]_ , \new_[70679]_ , \new_[70680]_ , \new_[70681]_ ,
    \new_[70685]_ , \new_[70686]_ , \new_[70689]_ , \new_[70692]_ ,
    \new_[70693]_ , \new_[70694]_ , \new_[70698]_ , \new_[70699]_ ,
    \new_[70702]_ , \new_[70705]_ , \new_[70706]_ , \new_[70707]_ ,
    \new_[70711]_ , \new_[70712]_ , \new_[70715]_ , \new_[70718]_ ,
    \new_[70719]_ , \new_[70720]_ , \new_[70724]_ , \new_[70725]_ ,
    \new_[70728]_ , \new_[70731]_ , \new_[70732]_ , \new_[70733]_ ,
    \new_[70737]_ , \new_[70738]_ , \new_[70741]_ , \new_[70744]_ ,
    \new_[70745]_ , \new_[70746]_ , \new_[70750]_ , \new_[70751]_ ,
    \new_[70754]_ , \new_[70757]_ , \new_[70758]_ , \new_[70759]_ ,
    \new_[70763]_ , \new_[70764]_ , \new_[70767]_ , \new_[70770]_ ,
    \new_[70771]_ , \new_[70772]_ , \new_[70776]_ , \new_[70777]_ ,
    \new_[70780]_ , \new_[70783]_ , \new_[70784]_ , \new_[70785]_ ,
    \new_[70789]_ , \new_[70790]_ , \new_[70793]_ , \new_[70796]_ ,
    \new_[70797]_ , \new_[70798]_ , \new_[70802]_ , \new_[70803]_ ,
    \new_[70806]_ , \new_[70809]_ , \new_[70810]_ , \new_[70811]_ ,
    \new_[70815]_ , \new_[70816]_ , \new_[70819]_ , \new_[70822]_ ,
    \new_[70823]_ , \new_[70824]_ , \new_[70828]_ , \new_[70829]_ ,
    \new_[70832]_ , \new_[70835]_ , \new_[70836]_ , \new_[70837]_ ,
    \new_[70841]_ , \new_[70842]_ , \new_[70845]_ , \new_[70848]_ ,
    \new_[70849]_ , \new_[70850]_ , \new_[70854]_ , \new_[70855]_ ,
    \new_[70858]_ , \new_[70861]_ , \new_[70862]_ , \new_[70863]_ ,
    \new_[70867]_ , \new_[70868]_ , \new_[70871]_ , \new_[70874]_ ,
    \new_[70875]_ , \new_[70876]_ , \new_[70880]_ , \new_[70881]_ ,
    \new_[70884]_ , \new_[70887]_ , \new_[70888]_ , \new_[70889]_ ,
    \new_[70893]_ , \new_[70894]_ , \new_[70897]_ , \new_[70900]_ ,
    \new_[70901]_ , \new_[70902]_ , \new_[70906]_ , \new_[70907]_ ,
    \new_[70910]_ , \new_[70913]_ , \new_[70914]_ , \new_[70915]_ ,
    \new_[70919]_ , \new_[70920]_ , \new_[70923]_ , \new_[70926]_ ,
    \new_[70927]_ , \new_[70928]_ , \new_[70932]_ , \new_[70933]_ ,
    \new_[70936]_ , \new_[70939]_ , \new_[70940]_ , \new_[70941]_ ,
    \new_[70945]_ , \new_[70946]_ , \new_[70949]_ , \new_[70952]_ ,
    \new_[70953]_ , \new_[70954]_ , \new_[70958]_ , \new_[70959]_ ,
    \new_[70962]_ , \new_[70965]_ , \new_[70966]_ , \new_[70967]_ ,
    \new_[70971]_ , \new_[70972]_ , \new_[70975]_ , \new_[70978]_ ,
    \new_[70979]_ , \new_[70980]_ , \new_[70984]_ , \new_[70985]_ ,
    \new_[70988]_ , \new_[70991]_ , \new_[70992]_ , \new_[70993]_ ,
    \new_[70997]_ , \new_[70998]_ , \new_[71001]_ , \new_[71004]_ ,
    \new_[71005]_ , \new_[71006]_ , \new_[71010]_ , \new_[71011]_ ,
    \new_[71014]_ , \new_[71017]_ , \new_[71018]_ , \new_[71019]_ ,
    \new_[71023]_ , \new_[71024]_ , \new_[71027]_ , \new_[71030]_ ,
    \new_[71031]_ , \new_[71032]_ , \new_[71036]_ , \new_[71037]_ ,
    \new_[71040]_ , \new_[71043]_ , \new_[71044]_ , \new_[71045]_ ,
    \new_[71049]_ , \new_[71050]_ , \new_[71053]_ , \new_[71056]_ ,
    \new_[71057]_ , \new_[71058]_ , \new_[71062]_ , \new_[71063]_ ,
    \new_[71066]_ , \new_[71069]_ , \new_[71070]_ , \new_[71071]_ ,
    \new_[71075]_ , \new_[71076]_ , \new_[71079]_ , \new_[71082]_ ,
    \new_[71083]_ , \new_[71084]_ , \new_[71088]_ , \new_[71089]_ ,
    \new_[71092]_ , \new_[71095]_ , \new_[71096]_ , \new_[71097]_ ,
    \new_[71101]_ , \new_[71102]_ , \new_[71105]_ , \new_[71108]_ ,
    \new_[71109]_ , \new_[71110]_ , \new_[71114]_ , \new_[71115]_ ,
    \new_[71118]_ , \new_[71121]_ , \new_[71122]_ , \new_[71123]_ ,
    \new_[71127]_ , \new_[71128]_ , \new_[71131]_ , \new_[71134]_ ,
    \new_[71135]_ , \new_[71136]_ , \new_[71140]_ , \new_[71141]_ ,
    \new_[71144]_ , \new_[71147]_ , \new_[71148]_ , \new_[71149]_ ,
    \new_[71153]_ , \new_[71154]_ , \new_[71157]_ , \new_[71160]_ ,
    \new_[71161]_ , \new_[71162]_ , \new_[71166]_ , \new_[71167]_ ,
    \new_[71170]_ , \new_[71173]_ , \new_[71174]_ , \new_[71175]_ ,
    \new_[71179]_ , \new_[71180]_ , \new_[71183]_ , \new_[71186]_ ,
    \new_[71187]_ , \new_[71188]_ , \new_[71192]_ , \new_[71193]_ ,
    \new_[71196]_ , \new_[71199]_ , \new_[71200]_ , \new_[71201]_ ,
    \new_[71205]_ , \new_[71206]_ , \new_[71209]_ , \new_[71212]_ ,
    \new_[71213]_ , \new_[71214]_ , \new_[71218]_ , \new_[71219]_ ,
    \new_[71222]_ , \new_[71225]_ , \new_[71226]_ , \new_[71227]_ ,
    \new_[71231]_ , \new_[71232]_ , \new_[71235]_ , \new_[71238]_ ,
    \new_[71239]_ , \new_[71240]_ , \new_[71244]_ , \new_[71245]_ ,
    \new_[71248]_ , \new_[71251]_ , \new_[71252]_ , \new_[71253]_ ,
    \new_[71257]_ , \new_[71258]_ , \new_[71261]_ , \new_[71264]_ ,
    \new_[71265]_ , \new_[71266]_ , \new_[71270]_ , \new_[71271]_ ,
    \new_[71274]_ , \new_[71277]_ , \new_[71278]_ , \new_[71279]_ ,
    \new_[71283]_ , \new_[71284]_ , \new_[71287]_ , \new_[71290]_ ,
    \new_[71291]_ , \new_[71292]_ , \new_[71296]_ , \new_[71297]_ ,
    \new_[71300]_ , \new_[71303]_ , \new_[71304]_ , \new_[71305]_ ,
    \new_[71309]_ , \new_[71310]_ , \new_[71313]_ , \new_[71316]_ ,
    \new_[71317]_ , \new_[71318]_ , \new_[71322]_ , \new_[71323]_ ,
    \new_[71326]_ , \new_[71329]_ , \new_[71330]_ , \new_[71331]_ ,
    \new_[71335]_ , \new_[71336]_ , \new_[71339]_ , \new_[71342]_ ,
    \new_[71343]_ , \new_[71344]_ , \new_[71348]_ , \new_[71349]_ ,
    \new_[71352]_ , \new_[71355]_ , \new_[71356]_ , \new_[71357]_ ,
    \new_[71361]_ , \new_[71362]_ , \new_[71365]_ , \new_[71368]_ ,
    \new_[71369]_ , \new_[71370]_ , \new_[71374]_ , \new_[71375]_ ,
    \new_[71378]_ , \new_[71381]_ , \new_[71382]_ , \new_[71383]_ ,
    \new_[71387]_ , \new_[71388]_ , \new_[71391]_ , \new_[71394]_ ,
    \new_[71395]_ , \new_[71396]_ , \new_[71400]_ , \new_[71401]_ ,
    \new_[71404]_ , \new_[71407]_ , \new_[71408]_ , \new_[71409]_ ,
    \new_[71413]_ , \new_[71414]_ , \new_[71417]_ , \new_[71420]_ ,
    \new_[71421]_ , \new_[71422]_ , \new_[71426]_ , \new_[71427]_ ,
    \new_[71430]_ , \new_[71433]_ , \new_[71434]_ , \new_[71435]_ ,
    \new_[71439]_ , \new_[71440]_ , \new_[71443]_ , \new_[71446]_ ,
    \new_[71447]_ , \new_[71448]_ , \new_[71452]_ , \new_[71453]_ ,
    \new_[71456]_ , \new_[71459]_ , \new_[71460]_ , \new_[71461]_ ,
    \new_[71465]_ , \new_[71466]_ , \new_[71469]_ , \new_[71472]_ ,
    \new_[71473]_ , \new_[71474]_ , \new_[71478]_ , \new_[71479]_ ,
    \new_[71482]_ , \new_[71485]_ , \new_[71486]_ , \new_[71487]_ ,
    \new_[71491]_ , \new_[71492]_ , \new_[71495]_ , \new_[71498]_ ,
    \new_[71499]_ , \new_[71500]_ , \new_[71504]_ , \new_[71505]_ ,
    \new_[71508]_ , \new_[71511]_ , \new_[71512]_ , \new_[71513]_ ,
    \new_[71517]_ , \new_[71518]_ , \new_[71521]_ , \new_[71524]_ ,
    \new_[71525]_ , \new_[71526]_ , \new_[71530]_ , \new_[71531]_ ,
    \new_[71534]_ , \new_[71537]_ , \new_[71538]_ , \new_[71539]_ ,
    \new_[71543]_ , \new_[71544]_ , \new_[71547]_ , \new_[71550]_ ,
    \new_[71551]_ , \new_[71552]_ , \new_[71556]_ , \new_[71557]_ ,
    \new_[71560]_ , \new_[71563]_ , \new_[71564]_ , \new_[71565]_ ,
    \new_[71569]_ , \new_[71570]_ , \new_[71573]_ , \new_[71576]_ ,
    \new_[71577]_ , \new_[71578]_ , \new_[71582]_ , \new_[71583]_ ,
    \new_[71586]_ , \new_[71589]_ , \new_[71590]_ , \new_[71591]_ ,
    \new_[71595]_ , \new_[71596]_ , \new_[71599]_ , \new_[71602]_ ,
    \new_[71603]_ , \new_[71604]_ , \new_[71608]_ , \new_[71609]_ ,
    \new_[71612]_ , \new_[71615]_ , \new_[71616]_ , \new_[71617]_ ,
    \new_[71621]_ , \new_[71622]_ , \new_[71625]_ , \new_[71628]_ ,
    \new_[71629]_ , \new_[71630]_ , \new_[71634]_ , \new_[71635]_ ,
    \new_[71638]_ , \new_[71641]_ , \new_[71642]_ , \new_[71643]_ ,
    \new_[71647]_ , \new_[71648]_ , \new_[71651]_ , \new_[71654]_ ,
    \new_[71655]_ , \new_[71656]_ , \new_[71660]_ , \new_[71661]_ ,
    \new_[71664]_ , \new_[71667]_ , \new_[71668]_ , \new_[71669]_ ,
    \new_[71673]_ , \new_[71674]_ , \new_[71677]_ , \new_[71680]_ ,
    \new_[71681]_ , \new_[71682]_ , \new_[71686]_ , \new_[71687]_ ,
    \new_[71690]_ , \new_[71693]_ , \new_[71694]_ , \new_[71695]_ ,
    \new_[71699]_ , \new_[71700]_ , \new_[71703]_ , \new_[71706]_ ,
    \new_[71707]_ , \new_[71708]_ , \new_[71712]_ , \new_[71713]_ ,
    \new_[71716]_ , \new_[71719]_ , \new_[71720]_ , \new_[71721]_ ,
    \new_[71725]_ , \new_[71726]_ , \new_[71729]_ , \new_[71732]_ ,
    \new_[71733]_ , \new_[71734]_ , \new_[71738]_ , \new_[71739]_ ,
    \new_[71742]_ , \new_[71745]_ , \new_[71746]_ , \new_[71747]_ ,
    \new_[71751]_ , \new_[71752]_ , \new_[71755]_ , \new_[71758]_ ,
    \new_[71759]_ , \new_[71760]_ , \new_[71764]_ , \new_[71765]_ ,
    \new_[71768]_ , \new_[71771]_ , \new_[71772]_ , \new_[71773]_ ,
    \new_[71777]_ , \new_[71778]_ , \new_[71781]_ , \new_[71784]_ ,
    \new_[71785]_ , \new_[71786]_ , \new_[71790]_ , \new_[71791]_ ,
    \new_[71794]_ , \new_[71797]_ , \new_[71798]_ , \new_[71799]_ ,
    \new_[71803]_ , \new_[71804]_ , \new_[71807]_ , \new_[71810]_ ,
    \new_[71811]_ , \new_[71812]_ , \new_[71816]_ , \new_[71817]_ ,
    \new_[71820]_ , \new_[71823]_ , \new_[71824]_ , \new_[71825]_ ,
    \new_[71829]_ , \new_[71830]_ , \new_[71833]_ , \new_[71836]_ ,
    \new_[71837]_ , \new_[71838]_ , \new_[71842]_ , \new_[71843]_ ,
    \new_[71846]_ , \new_[71849]_ , \new_[71850]_ , \new_[71851]_ ,
    \new_[71855]_ , \new_[71856]_ , \new_[71859]_ , \new_[71862]_ ,
    \new_[71863]_ , \new_[71864]_ , \new_[71868]_ , \new_[71869]_ ,
    \new_[71872]_ , \new_[71875]_ , \new_[71876]_ , \new_[71877]_ ,
    \new_[71881]_ , \new_[71882]_ , \new_[71885]_ , \new_[71888]_ ,
    \new_[71889]_ , \new_[71890]_ , \new_[71894]_ , \new_[71895]_ ,
    \new_[71898]_ , \new_[71901]_ , \new_[71902]_ , \new_[71903]_ ,
    \new_[71907]_ , \new_[71908]_ , \new_[71911]_ , \new_[71914]_ ,
    \new_[71915]_ , \new_[71916]_ , \new_[71920]_ , \new_[71921]_ ,
    \new_[71924]_ , \new_[71927]_ , \new_[71928]_ , \new_[71929]_ ,
    \new_[71933]_ , \new_[71934]_ , \new_[71937]_ , \new_[71940]_ ,
    \new_[71941]_ , \new_[71942]_ , \new_[71946]_ , \new_[71947]_ ,
    \new_[71950]_ , \new_[71953]_ , \new_[71954]_ , \new_[71955]_ ,
    \new_[71959]_ , \new_[71960]_ , \new_[71963]_ , \new_[71966]_ ,
    \new_[71967]_ , \new_[71968]_ , \new_[71972]_ , \new_[71973]_ ,
    \new_[71976]_ , \new_[71979]_ , \new_[71980]_ , \new_[71981]_ ,
    \new_[71985]_ , \new_[71986]_ , \new_[71989]_ , \new_[71992]_ ,
    \new_[71993]_ , \new_[71994]_ , \new_[71998]_ , \new_[71999]_ ,
    \new_[72002]_ , \new_[72005]_ , \new_[72006]_ , \new_[72007]_ ,
    \new_[72011]_ , \new_[72012]_ , \new_[72015]_ , \new_[72018]_ ,
    \new_[72019]_ , \new_[72020]_ , \new_[72024]_ , \new_[72025]_ ,
    \new_[72028]_ , \new_[72031]_ , \new_[72032]_ , \new_[72033]_ ,
    \new_[72037]_ , \new_[72038]_ , \new_[72041]_ , \new_[72044]_ ,
    \new_[72045]_ , \new_[72046]_ , \new_[72050]_ , \new_[72051]_ ,
    \new_[72054]_ , \new_[72057]_ , \new_[72058]_ , \new_[72059]_ ,
    \new_[72063]_ , \new_[72064]_ , \new_[72067]_ , \new_[72070]_ ,
    \new_[72071]_ , \new_[72072]_ , \new_[72076]_ , \new_[72077]_ ,
    \new_[72080]_ , \new_[72083]_ , \new_[72084]_ , \new_[72085]_ ,
    \new_[72089]_ , \new_[72090]_ , \new_[72093]_ , \new_[72096]_ ,
    \new_[72097]_ , \new_[72098]_ , \new_[72102]_ , \new_[72103]_ ,
    \new_[72106]_ , \new_[72109]_ , \new_[72110]_ , \new_[72111]_ ,
    \new_[72115]_ , \new_[72116]_ , \new_[72119]_ , \new_[72122]_ ,
    \new_[72123]_ , \new_[72124]_ , \new_[72128]_ , \new_[72129]_ ,
    \new_[72132]_ , \new_[72135]_ , \new_[72136]_ , \new_[72137]_ ,
    \new_[72141]_ , \new_[72142]_ , \new_[72145]_ , \new_[72148]_ ,
    \new_[72149]_ , \new_[72150]_ , \new_[72154]_ , \new_[72155]_ ,
    \new_[72158]_ , \new_[72161]_ , \new_[72162]_ , \new_[72163]_ ,
    \new_[72167]_ , \new_[72168]_ , \new_[72171]_ , \new_[72174]_ ,
    \new_[72175]_ , \new_[72176]_ , \new_[72180]_ , \new_[72181]_ ,
    \new_[72184]_ , \new_[72187]_ , \new_[72188]_ , \new_[72189]_ ,
    \new_[72193]_ , \new_[72194]_ , \new_[72197]_ , \new_[72200]_ ,
    \new_[72201]_ , \new_[72202]_ , \new_[72206]_ , \new_[72207]_ ,
    \new_[72210]_ , \new_[72213]_ , \new_[72214]_ , \new_[72215]_ ,
    \new_[72219]_ , \new_[72220]_ , \new_[72223]_ , \new_[72226]_ ,
    \new_[72227]_ , \new_[72228]_ , \new_[72232]_ , \new_[72233]_ ,
    \new_[72236]_ , \new_[72239]_ , \new_[72240]_ , \new_[72241]_ ,
    \new_[72245]_ , \new_[72246]_ , \new_[72249]_ , \new_[72252]_ ,
    \new_[72253]_ , \new_[72254]_ , \new_[72258]_ , \new_[72259]_ ,
    \new_[72262]_ , \new_[72265]_ , \new_[72266]_ , \new_[72267]_ ,
    \new_[72271]_ , \new_[72272]_ , \new_[72275]_ , \new_[72278]_ ,
    \new_[72279]_ , \new_[72280]_ , \new_[72284]_ , \new_[72285]_ ,
    \new_[72288]_ , \new_[72291]_ , \new_[72292]_ , \new_[72293]_ ,
    \new_[72297]_ , \new_[72298]_ , \new_[72301]_ , \new_[72304]_ ,
    \new_[72305]_ , \new_[72306]_ , \new_[72310]_ , \new_[72311]_ ,
    \new_[72314]_ , \new_[72317]_ , \new_[72318]_ , \new_[72319]_ ,
    \new_[72323]_ , \new_[72324]_ , \new_[72327]_ , \new_[72330]_ ,
    \new_[72331]_ , \new_[72332]_ , \new_[72336]_ , \new_[72337]_ ,
    \new_[72340]_ , \new_[72343]_ , \new_[72344]_ , \new_[72345]_ ,
    \new_[72349]_ , \new_[72350]_ , \new_[72353]_ , \new_[72356]_ ,
    \new_[72357]_ , \new_[72358]_ , \new_[72362]_ , \new_[72363]_ ,
    \new_[72366]_ , \new_[72369]_ , \new_[72370]_ , \new_[72371]_ ,
    \new_[72375]_ , \new_[72376]_ , \new_[72379]_ , \new_[72382]_ ,
    \new_[72383]_ , \new_[72384]_ , \new_[72388]_ , \new_[72389]_ ,
    \new_[72392]_ , \new_[72395]_ , \new_[72396]_ , \new_[72397]_ ,
    \new_[72401]_ , \new_[72402]_ , \new_[72405]_ , \new_[72408]_ ,
    \new_[72409]_ , \new_[72410]_ , \new_[72414]_ , \new_[72415]_ ,
    \new_[72418]_ , \new_[72421]_ , \new_[72422]_ , \new_[72423]_ ,
    \new_[72427]_ , \new_[72428]_ , \new_[72431]_ , \new_[72434]_ ,
    \new_[72435]_ , \new_[72436]_ , \new_[72440]_ , \new_[72441]_ ,
    \new_[72444]_ , \new_[72447]_ , \new_[72448]_ , \new_[72449]_ ,
    \new_[72453]_ , \new_[72454]_ , \new_[72457]_ , \new_[72460]_ ,
    \new_[72461]_ , \new_[72462]_ , \new_[72466]_ , \new_[72467]_ ,
    \new_[72470]_ , \new_[72473]_ , \new_[72474]_ , \new_[72475]_ ,
    \new_[72479]_ , \new_[72480]_ , \new_[72483]_ , \new_[72486]_ ,
    \new_[72487]_ , \new_[72488]_ , \new_[72492]_ , \new_[72493]_ ,
    \new_[72496]_ , \new_[72499]_ , \new_[72500]_ , \new_[72501]_ ,
    \new_[72505]_ , \new_[72506]_ , \new_[72509]_ , \new_[72512]_ ,
    \new_[72513]_ , \new_[72514]_ , \new_[72518]_ , \new_[72519]_ ,
    \new_[72522]_ , \new_[72525]_ , \new_[72526]_ , \new_[72527]_ ,
    \new_[72531]_ , \new_[72532]_ , \new_[72535]_ , \new_[72538]_ ,
    \new_[72539]_ , \new_[72540]_ , \new_[72544]_ , \new_[72545]_ ,
    \new_[72548]_ , \new_[72551]_ , \new_[72552]_ , \new_[72553]_ ,
    \new_[72557]_ , \new_[72558]_ , \new_[72561]_ , \new_[72564]_ ,
    \new_[72565]_ , \new_[72566]_ , \new_[72570]_ , \new_[72571]_ ,
    \new_[72574]_ , \new_[72577]_ , \new_[72578]_ , \new_[72579]_ ,
    \new_[72583]_ , \new_[72584]_ , \new_[72587]_ , \new_[72590]_ ,
    \new_[72591]_ , \new_[72592]_ , \new_[72596]_ , \new_[72597]_ ,
    \new_[72600]_ , \new_[72603]_ , \new_[72604]_ , \new_[72605]_ ,
    \new_[72609]_ , \new_[72610]_ , \new_[72613]_ , \new_[72616]_ ,
    \new_[72617]_ , \new_[72618]_ , \new_[72622]_ , \new_[72623]_ ,
    \new_[72626]_ , \new_[72629]_ , \new_[72630]_ , \new_[72631]_ ,
    \new_[72635]_ , \new_[72636]_ , \new_[72639]_ , \new_[72642]_ ,
    \new_[72643]_ , \new_[72644]_ , \new_[72648]_ , \new_[72649]_ ,
    \new_[72652]_ , \new_[72655]_ , \new_[72656]_ , \new_[72657]_ ,
    \new_[72661]_ , \new_[72662]_ , \new_[72665]_ , \new_[72668]_ ,
    \new_[72669]_ , \new_[72670]_ , \new_[72674]_ , \new_[72675]_ ,
    \new_[72678]_ , \new_[72681]_ , \new_[72682]_ , \new_[72683]_ ,
    \new_[72687]_ , \new_[72688]_ , \new_[72691]_ , \new_[72694]_ ,
    \new_[72695]_ , \new_[72696]_ , \new_[72700]_ , \new_[72701]_ ,
    \new_[72704]_ , \new_[72707]_ , \new_[72708]_ , \new_[72709]_ ,
    \new_[72713]_ , \new_[72714]_ , \new_[72717]_ , \new_[72720]_ ,
    \new_[72721]_ , \new_[72722]_ , \new_[72726]_ , \new_[72727]_ ,
    \new_[72730]_ , \new_[72733]_ , \new_[72734]_ , \new_[72735]_ ,
    \new_[72739]_ , \new_[72740]_ , \new_[72743]_ , \new_[72746]_ ,
    \new_[72747]_ , \new_[72748]_ , \new_[72752]_ , \new_[72753]_ ,
    \new_[72756]_ , \new_[72759]_ , \new_[72760]_ , \new_[72761]_ ,
    \new_[72765]_ , \new_[72766]_ , \new_[72769]_ , \new_[72772]_ ,
    \new_[72773]_ , \new_[72774]_ , \new_[72778]_ , \new_[72779]_ ,
    \new_[72782]_ , \new_[72785]_ , \new_[72786]_ , \new_[72787]_ ,
    \new_[72791]_ , \new_[72792]_ , \new_[72795]_ , \new_[72798]_ ,
    \new_[72799]_ , \new_[72800]_ , \new_[72804]_ , \new_[72805]_ ,
    \new_[72808]_ , \new_[72811]_ , \new_[72812]_ , \new_[72813]_ ,
    \new_[72817]_ , \new_[72818]_ , \new_[72821]_ , \new_[72824]_ ,
    \new_[72825]_ , \new_[72826]_ , \new_[72830]_ , \new_[72831]_ ,
    \new_[72834]_ , \new_[72837]_ , \new_[72838]_ , \new_[72839]_ ,
    \new_[72843]_ , \new_[72844]_ , \new_[72847]_ , \new_[72850]_ ,
    \new_[72851]_ , \new_[72852]_ , \new_[72856]_ , \new_[72857]_ ,
    \new_[72860]_ , \new_[72863]_ , \new_[72864]_ , \new_[72865]_ ,
    \new_[72869]_ , \new_[72870]_ , \new_[72873]_ , \new_[72876]_ ,
    \new_[72877]_ , \new_[72878]_ , \new_[72882]_ , \new_[72883]_ ,
    \new_[72886]_ , \new_[72889]_ , \new_[72890]_ , \new_[72891]_ ,
    \new_[72895]_ , \new_[72896]_ , \new_[72899]_ , \new_[72902]_ ,
    \new_[72903]_ , \new_[72904]_ , \new_[72908]_ , \new_[72909]_ ,
    \new_[72912]_ , \new_[72915]_ , \new_[72916]_ , \new_[72917]_ ,
    \new_[72921]_ , \new_[72922]_ , \new_[72925]_ , \new_[72928]_ ,
    \new_[72929]_ , \new_[72930]_ , \new_[72934]_ , \new_[72935]_ ,
    \new_[72938]_ , \new_[72941]_ , \new_[72942]_ , \new_[72943]_ ,
    \new_[72947]_ , \new_[72948]_ , \new_[72951]_ , \new_[72954]_ ,
    \new_[72955]_ , \new_[72956]_ , \new_[72960]_ , \new_[72961]_ ,
    \new_[72964]_ , \new_[72967]_ , \new_[72968]_ , \new_[72969]_ ,
    \new_[72973]_ , \new_[72974]_ , \new_[72977]_ , \new_[72980]_ ,
    \new_[72981]_ , \new_[72982]_ , \new_[72986]_ , \new_[72987]_ ,
    \new_[72990]_ , \new_[72993]_ , \new_[72994]_ , \new_[72995]_ ,
    \new_[72999]_ , \new_[73000]_ , \new_[73003]_ , \new_[73006]_ ,
    \new_[73007]_ , \new_[73008]_ , \new_[73012]_ , \new_[73013]_ ,
    \new_[73016]_ , \new_[73019]_ , \new_[73020]_ , \new_[73021]_ ,
    \new_[73025]_ , \new_[73026]_ , \new_[73029]_ , \new_[73032]_ ,
    \new_[73033]_ , \new_[73034]_ , \new_[73038]_ , \new_[73039]_ ,
    \new_[73042]_ , \new_[73045]_ , \new_[73046]_ , \new_[73047]_ ,
    \new_[73051]_ , \new_[73052]_ , \new_[73055]_ , \new_[73058]_ ,
    \new_[73059]_ , \new_[73060]_ , \new_[73064]_ , \new_[73065]_ ,
    \new_[73068]_ , \new_[73071]_ , \new_[73072]_ , \new_[73073]_ ,
    \new_[73077]_ , \new_[73078]_ , \new_[73081]_ , \new_[73084]_ ,
    \new_[73085]_ , \new_[73086]_ , \new_[73090]_ , \new_[73091]_ ,
    \new_[73094]_ , \new_[73097]_ , \new_[73098]_ , \new_[73099]_ ,
    \new_[73103]_ , \new_[73104]_ , \new_[73107]_ , \new_[73110]_ ,
    \new_[73111]_ , \new_[73112]_ , \new_[73116]_ , \new_[73117]_ ,
    \new_[73120]_ , \new_[73123]_ , \new_[73124]_ , \new_[73125]_ ,
    \new_[73129]_ , \new_[73130]_ , \new_[73133]_ , \new_[73136]_ ,
    \new_[73137]_ , \new_[73138]_ , \new_[73142]_ , \new_[73143]_ ,
    \new_[73146]_ , \new_[73149]_ , \new_[73150]_ , \new_[73151]_ ,
    \new_[73155]_ , \new_[73156]_ , \new_[73159]_ , \new_[73162]_ ,
    \new_[73163]_ , \new_[73164]_ , \new_[73168]_ , \new_[73169]_ ,
    \new_[73172]_ , \new_[73175]_ , \new_[73176]_ , \new_[73177]_ ,
    \new_[73181]_ , \new_[73182]_ , \new_[73185]_ , \new_[73188]_ ,
    \new_[73189]_ , \new_[73190]_ , \new_[73194]_ , \new_[73195]_ ,
    \new_[73198]_ , \new_[73201]_ , \new_[73202]_ , \new_[73203]_ ,
    \new_[73207]_ , \new_[73208]_ , \new_[73211]_ , \new_[73214]_ ,
    \new_[73215]_ , \new_[73216]_ , \new_[73220]_ , \new_[73221]_ ,
    \new_[73224]_ , \new_[73227]_ , \new_[73228]_ , \new_[73229]_ ,
    \new_[73233]_ , \new_[73234]_ , \new_[73237]_ , \new_[73240]_ ,
    \new_[73241]_ , \new_[73242]_ , \new_[73246]_ , \new_[73247]_ ,
    \new_[73250]_ , \new_[73253]_ , \new_[73254]_ , \new_[73255]_ ,
    \new_[73259]_ , \new_[73260]_ , \new_[73263]_ , \new_[73266]_ ,
    \new_[73267]_ , \new_[73268]_ , \new_[73272]_ , \new_[73273]_ ,
    \new_[73276]_ , \new_[73279]_ , \new_[73280]_ , \new_[73281]_ ,
    \new_[73285]_ , \new_[73286]_ , \new_[73289]_ , \new_[73292]_ ,
    \new_[73293]_ , \new_[73294]_ , \new_[73298]_ , \new_[73299]_ ,
    \new_[73302]_ , \new_[73305]_ , \new_[73306]_ , \new_[73307]_ ,
    \new_[73311]_ , \new_[73312]_ , \new_[73315]_ , \new_[73318]_ ,
    \new_[73319]_ , \new_[73320]_ , \new_[73324]_ , \new_[73325]_ ,
    \new_[73328]_ , \new_[73331]_ , \new_[73332]_ , \new_[73333]_ ,
    \new_[73337]_ , \new_[73338]_ , \new_[73341]_ , \new_[73344]_ ,
    \new_[73345]_ , \new_[73346]_ , \new_[73350]_ , \new_[73351]_ ,
    \new_[73354]_ , \new_[73357]_ , \new_[73358]_ , \new_[73359]_ ,
    \new_[73363]_ , \new_[73364]_ , \new_[73367]_ , \new_[73370]_ ,
    \new_[73371]_ , \new_[73372]_ , \new_[73376]_ , \new_[73377]_ ,
    \new_[73380]_ , \new_[73383]_ , \new_[73384]_ , \new_[73385]_ ,
    \new_[73389]_ , \new_[73390]_ , \new_[73393]_ , \new_[73396]_ ,
    \new_[73397]_ , \new_[73398]_ , \new_[73402]_ , \new_[73403]_ ,
    \new_[73406]_ , \new_[73409]_ , \new_[73410]_ , \new_[73411]_ ,
    \new_[73415]_ , \new_[73416]_ , \new_[73419]_ , \new_[73422]_ ,
    \new_[73423]_ , \new_[73424]_ , \new_[73428]_ , \new_[73429]_ ,
    \new_[73432]_ , \new_[73435]_ , \new_[73436]_ , \new_[73437]_ ,
    \new_[73441]_ , \new_[73442]_ , \new_[73445]_ , \new_[73448]_ ,
    \new_[73449]_ , \new_[73450]_ , \new_[73454]_ , \new_[73455]_ ,
    \new_[73458]_ , \new_[73461]_ , \new_[73462]_ , \new_[73463]_ ,
    \new_[73467]_ , \new_[73468]_ , \new_[73471]_ , \new_[73474]_ ,
    \new_[73475]_ , \new_[73476]_ , \new_[73480]_ , \new_[73481]_ ,
    \new_[73484]_ , \new_[73487]_ , \new_[73488]_ , \new_[73489]_ ,
    \new_[73493]_ , \new_[73494]_ , \new_[73497]_ , \new_[73500]_ ,
    \new_[73501]_ , \new_[73502]_ , \new_[73506]_ , \new_[73507]_ ,
    \new_[73510]_ , \new_[73513]_ , \new_[73514]_ , \new_[73515]_ ,
    \new_[73519]_ , \new_[73520]_ , \new_[73523]_ , \new_[73526]_ ,
    \new_[73527]_ , \new_[73528]_ , \new_[73532]_ , \new_[73533]_ ,
    \new_[73536]_ , \new_[73539]_ , \new_[73540]_ , \new_[73541]_ ,
    \new_[73545]_ , \new_[73546]_ , \new_[73549]_ , \new_[73552]_ ,
    \new_[73553]_ , \new_[73554]_ , \new_[73558]_ , \new_[73559]_ ,
    \new_[73562]_ , \new_[73565]_ , \new_[73566]_ , \new_[73567]_ ,
    \new_[73571]_ , \new_[73572]_ , \new_[73575]_ , \new_[73578]_ ,
    \new_[73579]_ , \new_[73580]_ , \new_[73584]_ , \new_[73585]_ ,
    \new_[73588]_ , \new_[73591]_ , \new_[73592]_ , \new_[73593]_ ,
    \new_[73597]_ , \new_[73598]_ , \new_[73601]_ , \new_[73604]_ ,
    \new_[73605]_ , \new_[73606]_ , \new_[73610]_ , \new_[73611]_ ,
    \new_[73614]_ , \new_[73617]_ , \new_[73618]_ , \new_[73619]_ ,
    \new_[73623]_ , \new_[73624]_ , \new_[73627]_ , \new_[73630]_ ,
    \new_[73631]_ , \new_[73632]_ , \new_[73636]_ , \new_[73637]_ ,
    \new_[73640]_ , \new_[73643]_ , \new_[73644]_ , \new_[73645]_ ,
    \new_[73649]_ , \new_[73650]_ , \new_[73653]_ , \new_[73656]_ ,
    \new_[73657]_ , \new_[73658]_ , \new_[73662]_ , \new_[73663]_ ,
    \new_[73666]_ , \new_[73669]_ , \new_[73670]_ , \new_[73671]_ ,
    \new_[73675]_ , \new_[73676]_ , \new_[73679]_ , \new_[73682]_ ,
    \new_[73683]_ , \new_[73684]_ , \new_[73688]_ , \new_[73689]_ ,
    \new_[73692]_ , \new_[73695]_ , \new_[73696]_ , \new_[73697]_ ,
    \new_[73701]_ , \new_[73702]_ , \new_[73705]_ , \new_[73708]_ ,
    \new_[73709]_ , \new_[73710]_ , \new_[73714]_ , \new_[73715]_ ,
    \new_[73718]_ , \new_[73721]_ , \new_[73722]_ , \new_[73723]_ ,
    \new_[73727]_ , \new_[73728]_ , \new_[73731]_ , \new_[73734]_ ,
    \new_[73735]_ , \new_[73736]_ , \new_[73740]_ , \new_[73741]_ ,
    \new_[73744]_ , \new_[73747]_ , \new_[73748]_ , \new_[73749]_ ,
    \new_[73753]_ , \new_[73754]_ , \new_[73757]_ , \new_[73760]_ ,
    \new_[73761]_ , \new_[73762]_ , \new_[73766]_ , \new_[73767]_ ,
    \new_[73770]_ , \new_[73773]_ , \new_[73774]_ , \new_[73775]_ ,
    \new_[73779]_ , \new_[73780]_ , \new_[73783]_ , \new_[73786]_ ,
    \new_[73787]_ , \new_[73788]_ , \new_[73792]_ , \new_[73793]_ ,
    \new_[73796]_ , \new_[73799]_ , \new_[73800]_ , \new_[73801]_ ,
    \new_[73805]_ , \new_[73806]_ , \new_[73809]_ , \new_[73812]_ ,
    \new_[73813]_ , \new_[73814]_ , \new_[73818]_ , \new_[73819]_ ,
    \new_[73822]_ , \new_[73825]_ , \new_[73826]_ , \new_[73827]_ ,
    \new_[73831]_ , \new_[73832]_ , \new_[73835]_ , \new_[73838]_ ,
    \new_[73839]_ , \new_[73840]_ , \new_[73844]_ , \new_[73845]_ ,
    \new_[73848]_ , \new_[73851]_ , \new_[73852]_ , \new_[73853]_ ,
    \new_[73857]_ , \new_[73858]_ , \new_[73861]_ , \new_[73864]_ ,
    \new_[73865]_ , \new_[73866]_ , \new_[73870]_ , \new_[73871]_ ,
    \new_[73874]_ , \new_[73877]_ , \new_[73878]_ , \new_[73879]_ ,
    \new_[73883]_ , \new_[73884]_ , \new_[73887]_ , \new_[73890]_ ,
    \new_[73891]_ , \new_[73892]_ , \new_[73896]_ , \new_[73897]_ ,
    \new_[73900]_ , \new_[73903]_ , \new_[73904]_ , \new_[73905]_ ,
    \new_[73909]_ , \new_[73910]_ , \new_[73913]_ , \new_[73916]_ ,
    \new_[73917]_ , \new_[73918]_ , \new_[73922]_ , \new_[73923]_ ,
    \new_[73926]_ , \new_[73929]_ , \new_[73930]_ , \new_[73931]_ ,
    \new_[73935]_ , \new_[73936]_ , \new_[73939]_ , \new_[73942]_ ,
    \new_[73943]_ , \new_[73944]_ , \new_[73948]_ , \new_[73949]_ ,
    \new_[73952]_ , \new_[73955]_ , \new_[73956]_ , \new_[73957]_ ,
    \new_[73961]_ , \new_[73962]_ , \new_[73965]_ , \new_[73968]_ ,
    \new_[73969]_ , \new_[73970]_ , \new_[73974]_ , \new_[73975]_ ,
    \new_[73978]_ , \new_[73981]_ , \new_[73982]_ , \new_[73983]_ ,
    \new_[73987]_ , \new_[73988]_ , \new_[73991]_ , \new_[73994]_ ,
    \new_[73995]_ , \new_[73996]_ , \new_[74000]_ , \new_[74001]_ ,
    \new_[74004]_ , \new_[74007]_ , \new_[74008]_ , \new_[74009]_ ,
    \new_[74013]_ , \new_[74014]_ , \new_[74017]_ , \new_[74020]_ ,
    \new_[74021]_ , \new_[74022]_ , \new_[74026]_ , \new_[74027]_ ,
    \new_[74030]_ , \new_[74033]_ , \new_[74034]_ , \new_[74035]_ ,
    \new_[74039]_ , \new_[74040]_ , \new_[74043]_ , \new_[74046]_ ,
    \new_[74047]_ , \new_[74048]_ , \new_[74052]_ , \new_[74053]_ ,
    \new_[74056]_ , \new_[74059]_ , \new_[74060]_ , \new_[74061]_ ,
    \new_[74065]_ , \new_[74066]_ , \new_[74069]_ , \new_[74072]_ ,
    \new_[74073]_ , \new_[74074]_ , \new_[74078]_ , \new_[74079]_ ,
    \new_[74082]_ , \new_[74085]_ , \new_[74086]_ , \new_[74087]_ ,
    \new_[74091]_ , \new_[74092]_ , \new_[74095]_ , \new_[74098]_ ,
    \new_[74099]_ , \new_[74100]_ , \new_[74104]_ , \new_[74105]_ ,
    \new_[74108]_ , \new_[74111]_ , \new_[74112]_ , \new_[74113]_ ,
    \new_[74117]_ , \new_[74118]_ , \new_[74121]_ , \new_[74124]_ ,
    \new_[74125]_ , \new_[74126]_ , \new_[74130]_ , \new_[74131]_ ,
    \new_[74134]_ , \new_[74137]_ , \new_[74138]_ , \new_[74139]_ ,
    \new_[74143]_ , \new_[74144]_ , \new_[74147]_ , \new_[74150]_ ,
    \new_[74151]_ , \new_[74152]_ , \new_[74156]_ , \new_[74157]_ ,
    \new_[74160]_ , \new_[74163]_ , \new_[74164]_ , \new_[74165]_ ,
    \new_[74169]_ , \new_[74170]_ , \new_[74173]_ , \new_[74176]_ ,
    \new_[74177]_ , \new_[74178]_ , \new_[74182]_ , \new_[74183]_ ,
    \new_[74186]_ , \new_[74189]_ , \new_[74190]_ , \new_[74191]_ ,
    \new_[74195]_ , \new_[74196]_ , \new_[74199]_ , \new_[74202]_ ,
    \new_[74203]_ , \new_[74204]_ , \new_[74208]_ , \new_[74209]_ ,
    \new_[74212]_ , \new_[74215]_ , \new_[74216]_ , \new_[74217]_ ,
    \new_[74221]_ , \new_[74222]_ , \new_[74225]_ , \new_[74228]_ ,
    \new_[74229]_ , \new_[74230]_ , \new_[74234]_ , \new_[74235]_ ,
    \new_[74238]_ , \new_[74241]_ , \new_[74242]_ , \new_[74243]_ ,
    \new_[74247]_ , \new_[74248]_ , \new_[74251]_ , \new_[74254]_ ,
    \new_[74255]_ , \new_[74256]_ , \new_[74260]_ , \new_[74261]_ ,
    \new_[74264]_ , \new_[74267]_ , \new_[74268]_ , \new_[74269]_ ,
    \new_[74273]_ , \new_[74274]_ , \new_[74277]_ , \new_[74280]_ ,
    \new_[74281]_ , \new_[74282]_ , \new_[74286]_ , \new_[74287]_ ,
    \new_[74290]_ , \new_[74293]_ , \new_[74294]_ , \new_[74295]_ ,
    \new_[74299]_ , \new_[74300]_ , \new_[74303]_ , \new_[74306]_ ,
    \new_[74307]_ , \new_[74308]_ , \new_[74312]_ , \new_[74313]_ ,
    \new_[74316]_ , \new_[74319]_ , \new_[74320]_ , \new_[74321]_ ,
    \new_[74325]_ , \new_[74326]_ , \new_[74329]_ , \new_[74332]_ ,
    \new_[74333]_ , \new_[74334]_ , \new_[74338]_ , \new_[74339]_ ,
    \new_[74342]_ , \new_[74345]_ , \new_[74346]_ , \new_[74347]_ ,
    \new_[74351]_ , \new_[74352]_ , \new_[74355]_ , \new_[74358]_ ,
    \new_[74359]_ , \new_[74360]_ , \new_[74364]_ , \new_[74365]_ ,
    \new_[74368]_ , \new_[74371]_ , \new_[74372]_ , \new_[74373]_ ,
    \new_[74377]_ , \new_[74378]_ , \new_[74381]_ , \new_[74384]_ ,
    \new_[74385]_ , \new_[74386]_ , \new_[74390]_ , \new_[74391]_ ,
    \new_[74394]_ , \new_[74397]_ , \new_[74398]_ , \new_[74399]_ ,
    \new_[74403]_ , \new_[74404]_ , \new_[74407]_ , \new_[74410]_ ,
    \new_[74411]_ , \new_[74412]_ , \new_[74416]_ , \new_[74417]_ ,
    \new_[74420]_ , \new_[74423]_ , \new_[74424]_ , \new_[74425]_ ,
    \new_[74429]_ , \new_[74430]_ , \new_[74433]_ , \new_[74436]_ ,
    \new_[74437]_ , \new_[74438]_ , \new_[74442]_ , \new_[74443]_ ,
    \new_[74446]_ , \new_[74449]_ , \new_[74450]_ , \new_[74451]_ ,
    \new_[74455]_ , \new_[74456]_ , \new_[74459]_ , \new_[74462]_ ,
    \new_[74463]_ , \new_[74464]_ , \new_[74468]_ , \new_[74469]_ ,
    \new_[74472]_ , \new_[74475]_ , \new_[74476]_ , \new_[74477]_ ,
    \new_[74481]_ , \new_[74482]_ , \new_[74485]_ , \new_[74488]_ ,
    \new_[74489]_ , \new_[74490]_ , \new_[74494]_ , \new_[74495]_ ,
    \new_[74498]_ , \new_[74501]_ , \new_[74502]_ , \new_[74503]_ ,
    \new_[74507]_ , \new_[74508]_ , \new_[74511]_ , \new_[74514]_ ,
    \new_[74515]_ , \new_[74516]_ , \new_[74520]_ , \new_[74521]_ ,
    \new_[74524]_ , \new_[74527]_ , \new_[74528]_ , \new_[74529]_ ,
    \new_[74533]_ , \new_[74534]_ , \new_[74537]_ , \new_[74540]_ ,
    \new_[74541]_ , \new_[74542]_ , \new_[74546]_ , \new_[74547]_ ,
    \new_[74550]_ , \new_[74553]_ , \new_[74554]_ , \new_[74555]_ ,
    \new_[74559]_ , \new_[74560]_ , \new_[74563]_ , \new_[74566]_ ,
    \new_[74567]_ , \new_[74568]_ , \new_[74572]_ , \new_[74573]_ ,
    \new_[74576]_ , \new_[74579]_ , \new_[74580]_ , \new_[74581]_ ,
    \new_[74585]_ , \new_[74586]_ , \new_[74589]_ , \new_[74592]_ ,
    \new_[74593]_ , \new_[74594]_ , \new_[74598]_ , \new_[74599]_ ,
    \new_[74602]_ , \new_[74605]_ , \new_[74606]_ , \new_[74607]_ ,
    \new_[74611]_ , \new_[74612]_ , \new_[74615]_ , \new_[74618]_ ,
    \new_[74619]_ , \new_[74620]_ , \new_[74624]_ , \new_[74625]_ ,
    \new_[74628]_ , \new_[74631]_ , \new_[74632]_ , \new_[74633]_ ,
    \new_[74637]_ , \new_[74638]_ , \new_[74641]_ , \new_[74644]_ ,
    \new_[74645]_ , \new_[74646]_ , \new_[74650]_ , \new_[74651]_ ,
    \new_[74654]_ , \new_[74657]_ , \new_[74658]_ , \new_[74659]_ ,
    \new_[74663]_ , \new_[74664]_ , \new_[74667]_ , \new_[74670]_ ,
    \new_[74671]_ , \new_[74672]_ , \new_[74676]_ , \new_[74677]_ ,
    \new_[74680]_ , \new_[74683]_ , \new_[74684]_ , \new_[74685]_ ,
    \new_[74689]_ , \new_[74690]_ , \new_[74693]_ , \new_[74696]_ ,
    \new_[74697]_ , \new_[74698]_ , \new_[74702]_ , \new_[74703]_ ,
    \new_[74706]_ , \new_[74709]_ , \new_[74710]_ , \new_[74711]_ ,
    \new_[74715]_ , \new_[74716]_ , \new_[74719]_ , \new_[74722]_ ,
    \new_[74723]_ , \new_[74724]_ , \new_[74728]_ , \new_[74729]_ ,
    \new_[74732]_ , \new_[74735]_ , \new_[74736]_ , \new_[74737]_ ,
    \new_[74741]_ , \new_[74742]_ , \new_[74745]_ , \new_[74748]_ ,
    \new_[74749]_ , \new_[74750]_ , \new_[74754]_ , \new_[74755]_ ,
    \new_[74758]_ , \new_[74761]_ , \new_[74762]_ , \new_[74763]_ ,
    \new_[74767]_ , \new_[74768]_ , \new_[74771]_ , \new_[74774]_ ,
    \new_[74775]_ , \new_[74776]_ , \new_[74780]_ , \new_[74781]_ ,
    \new_[74784]_ , \new_[74787]_ , \new_[74788]_ , \new_[74789]_ ,
    \new_[74793]_ , \new_[74794]_ , \new_[74797]_ , \new_[74800]_ ,
    \new_[74801]_ , \new_[74802]_ , \new_[74806]_ , \new_[74807]_ ,
    \new_[74810]_ , \new_[74813]_ , \new_[74814]_ , \new_[74815]_ ,
    \new_[74819]_ , \new_[74820]_ , \new_[74823]_ , \new_[74826]_ ,
    \new_[74827]_ , \new_[74828]_ , \new_[74832]_ , \new_[74833]_ ,
    \new_[74836]_ , \new_[74839]_ , \new_[74840]_ , \new_[74841]_ ,
    \new_[74845]_ , \new_[74846]_ , \new_[74849]_ , \new_[74852]_ ,
    \new_[74853]_ , \new_[74854]_ , \new_[74858]_ , \new_[74859]_ ,
    \new_[74862]_ , \new_[74865]_ , \new_[74866]_ , \new_[74867]_ ,
    \new_[74871]_ , \new_[74872]_ , \new_[74875]_ , \new_[74878]_ ,
    \new_[74879]_ , \new_[74880]_ , \new_[74884]_ , \new_[74885]_ ,
    \new_[74888]_ , \new_[74891]_ , \new_[74892]_ , \new_[74893]_ ,
    \new_[74897]_ , \new_[74898]_ , \new_[74901]_ , \new_[74904]_ ,
    \new_[74905]_ , \new_[74906]_ , \new_[74910]_ , \new_[74911]_ ,
    \new_[74914]_ , \new_[74917]_ , \new_[74918]_ , \new_[74919]_ ,
    \new_[74923]_ , \new_[74924]_ , \new_[74927]_ , \new_[74930]_ ,
    \new_[74931]_ , \new_[74932]_ , \new_[74936]_ , \new_[74937]_ ,
    \new_[74940]_ , \new_[74943]_ , \new_[74944]_ , \new_[74945]_ ,
    \new_[74949]_ , \new_[74950]_ , \new_[74953]_ , \new_[74956]_ ,
    \new_[74957]_ , \new_[74958]_ , \new_[74962]_ , \new_[74963]_ ,
    \new_[74966]_ , \new_[74969]_ , \new_[74970]_ , \new_[74971]_ ,
    \new_[74975]_ , \new_[74976]_ , \new_[74979]_ , \new_[74982]_ ,
    \new_[74983]_ , \new_[74984]_ , \new_[74988]_ , \new_[74989]_ ,
    \new_[74992]_ , \new_[74995]_ , \new_[74996]_ , \new_[74997]_ ,
    \new_[75001]_ , \new_[75002]_ , \new_[75005]_ , \new_[75008]_ ,
    \new_[75009]_ , \new_[75010]_ , \new_[75014]_ , \new_[75015]_ ,
    \new_[75018]_ , \new_[75021]_ , \new_[75022]_ , \new_[75023]_ ,
    \new_[75027]_ , \new_[75028]_ , \new_[75031]_ , \new_[75034]_ ,
    \new_[75035]_ , \new_[75036]_ , \new_[75040]_ , \new_[75041]_ ,
    \new_[75044]_ , \new_[75047]_ , \new_[75048]_ , \new_[75049]_ ,
    \new_[75053]_ , \new_[75054]_ , \new_[75057]_ , \new_[75060]_ ,
    \new_[75061]_ , \new_[75062]_ , \new_[75066]_ , \new_[75067]_ ,
    \new_[75070]_ , \new_[75073]_ , \new_[75074]_ , \new_[75075]_ ,
    \new_[75079]_ , \new_[75080]_ , \new_[75083]_ , \new_[75086]_ ,
    \new_[75087]_ , \new_[75088]_ , \new_[75092]_ , \new_[75093]_ ,
    \new_[75096]_ , \new_[75099]_ , \new_[75100]_ , \new_[75101]_ ,
    \new_[75105]_ , \new_[75106]_ , \new_[75109]_ , \new_[75112]_ ,
    \new_[75113]_ , \new_[75114]_ , \new_[75118]_ , \new_[75119]_ ,
    \new_[75122]_ , \new_[75125]_ , \new_[75126]_ , \new_[75127]_ ,
    \new_[75131]_ , \new_[75132]_ , \new_[75135]_ , \new_[75138]_ ,
    \new_[75139]_ , \new_[75140]_ , \new_[75144]_ , \new_[75145]_ ,
    \new_[75148]_ , \new_[75151]_ , \new_[75152]_ , \new_[75153]_ ,
    \new_[75157]_ , \new_[75158]_ , \new_[75161]_ , \new_[75164]_ ,
    \new_[75165]_ , \new_[75166]_ , \new_[75170]_ , \new_[75171]_ ,
    \new_[75174]_ , \new_[75177]_ , \new_[75178]_ , \new_[75179]_ ,
    \new_[75183]_ , \new_[75184]_ , \new_[75187]_ , \new_[75190]_ ,
    \new_[75191]_ , \new_[75192]_ , \new_[75196]_ , \new_[75197]_ ,
    \new_[75200]_ , \new_[75203]_ , \new_[75204]_ , \new_[75205]_ ,
    \new_[75209]_ , \new_[75210]_ , \new_[75213]_ , \new_[75216]_ ,
    \new_[75217]_ , \new_[75218]_ , \new_[75222]_ , \new_[75223]_ ,
    \new_[75226]_ , \new_[75229]_ , \new_[75230]_ , \new_[75231]_ ,
    \new_[75235]_ , \new_[75236]_ , \new_[75239]_ , \new_[75242]_ ,
    \new_[75243]_ , \new_[75244]_ , \new_[75248]_ , \new_[75249]_ ,
    \new_[75252]_ , \new_[75255]_ , \new_[75256]_ , \new_[75257]_ ,
    \new_[75261]_ , \new_[75262]_ , \new_[75265]_ , \new_[75268]_ ,
    \new_[75269]_ , \new_[75270]_ , \new_[75274]_ , \new_[75275]_ ,
    \new_[75278]_ , \new_[75281]_ , \new_[75282]_ , \new_[75283]_ ,
    \new_[75287]_ , \new_[75288]_ , \new_[75291]_ , \new_[75294]_ ,
    \new_[75295]_ , \new_[75296]_ , \new_[75300]_ , \new_[75301]_ ,
    \new_[75304]_ , \new_[75307]_ , \new_[75308]_ , \new_[75309]_ ,
    \new_[75313]_ , \new_[75314]_ , \new_[75317]_ , \new_[75320]_ ,
    \new_[75321]_ , \new_[75322]_ , \new_[75326]_ , \new_[75327]_ ,
    \new_[75330]_ , \new_[75333]_ , \new_[75334]_ , \new_[75335]_ ,
    \new_[75339]_ , \new_[75340]_ , \new_[75343]_ , \new_[75346]_ ,
    \new_[75347]_ , \new_[75348]_ , \new_[75352]_ , \new_[75353]_ ,
    \new_[75356]_ , \new_[75359]_ , \new_[75360]_ , \new_[75361]_ ,
    \new_[75365]_ , \new_[75366]_ , \new_[75369]_ , \new_[75372]_ ,
    \new_[75373]_ , \new_[75374]_ , \new_[75378]_ , \new_[75379]_ ,
    \new_[75382]_ , \new_[75385]_ , \new_[75386]_ , \new_[75387]_ ,
    \new_[75391]_ , \new_[75392]_ , \new_[75395]_ , \new_[75398]_ ,
    \new_[75399]_ , \new_[75400]_ , \new_[75404]_ , \new_[75405]_ ,
    \new_[75408]_ , \new_[75411]_ , \new_[75412]_ , \new_[75413]_ ,
    \new_[75417]_ , \new_[75418]_ , \new_[75421]_ , \new_[75424]_ ,
    \new_[75425]_ , \new_[75426]_ , \new_[75430]_ , \new_[75431]_ ,
    \new_[75434]_ , \new_[75437]_ , \new_[75438]_ , \new_[75439]_ ,
    \new_[75443]_ , \new_[75444]_ , \new_[75447]_ , \new_[75450]_ ,
    \new_[75451]_ , \new_[75452]_ , \new_[75456]_ , \new_[75457]_ ,
    \new_[75460]_ , \new_[75463]_ , \new_[75464]_ , \new_[75465]_ ,
    \new_[75469]_ , \new_[75470]_ , \new_[75473]_ , \new_[75476]_ ,
    \new_[75477]_ , \new_[75478]_ , \new_[75482]_ , \new_[75483]_ ,
    \new_[75486]_ , \new_[75489]_ , \new_[75490]_ , \new_[75491]_ ,
    \new_[75495]_ , \new_[75496]_ , \new_[75499]_ , \new_[75502]_ ,
    \new_[75503]_ , \new_[75504]_ , \new_[75508]_ , \new_[75509]_ ,
    \new_[75512]_ , \new_[75515]_ , \new_[75516]_ , \new_[75517]_ ,
    \new_[75521]_ , \new_[75522]_ , \new_[75525]_ , \new_[75528]_ ,
    \new_[75529]_ , \new_[75530]_ , \new_[75534]_ , \new_[75535]_ ,
    \new_[75538]_ , \new_[75541]_ , \new_[75542]_ , \new_[75543]_ ,
    \new_[75547]_ , \new_[75548]_ , \new_[75551]_ , \new_[75554]_ ,
    \new_[75555]_ , \new_[75556]_ , \new_[75560]_ , \new_[75561]_ ,
    \new_[75564]_ , \new_[75567]_ , \new_[75568]_ , \new_[75569]_ ,
    \new_[75573]_ , \new_[75574]_ , \new_[75577]_ , \new_[75580]_ ,
    \new_[75581]_ , \new_[75582]_ , \new_[75586]_ , \new_[75587]_ ,
    \new_[75590]_ , \new_[75593]_ , \new_[75594]_ , \new_[75595]_ ,
    \new_[75599]_ , \new_[75600]_ , \new_[75603]_ , \new_[75606]_ ,
    \new_[75607]_ , \new_[75608]_ , \new_[75612]_ , \new_[75613]_ ,
    \new_[75616]_ , \new_[75619]_ , \new_[75620]_ , \new_[75621]_ ,
    \new_[75625]_ , \new_[75626]_ , \new_[75629]_ , \new_[75632]_ ,
    \new_[75633]_ , \new_[75634]_ , \new_[75638]_ , \new_[75639]_ ,
    \new_[75642]_ , \new_[75645]_ , \new_[75646]_ , \new_[75647]_ ,
    \new_[75651]_ , \new_[75652]_ , \new_[75655]_ , \new_[75658]_ ,
    \new_[75659]_ , \new_[75660]_ , \new_[75664]_ , \new_[75665]_ ,
    \new_[75668]_ , \new_[75671]_ , \new_[75672]_ , \new_[75673]_ ,
    \new_[75677]_ , \new_[75678]_ , \new_[75681]_ , \new_[75684]_ ,
    \new_[75685]_ , \new_[75686]_ , \new_[75690]_ , \new_[75691]_ ,
    \new_[75694]_ , \new_[75697]_ , \new_[75698]_ , \new_[75699]_ ,
    \new_[75703]_ , \new_[75704]_ , \new_[75707]_ , \new_[75710]_ ,
    \new_[75711]_ , \new_[75712]_ , \new_[75716]_ , \new_[75717]_ ,
    \new_[75720]_ , \new_[75723]_ , \new_[75724]_ , \new_[75725]_ ,
    \new_[75729]_ , \new_[75730]_ , \new_[75733]_ , \new_[75736]_ ,
    \new_[75737]_ , \new_[75738]_ , \new_[75742]_ , \new_[75743]_ ,
    \new_[75746]_ , \new_[75749]_ , \new_[75750]_ , \new_[75751]_ ,
    \new_[75755]_ , \new_[75756]_ , \new_[75759]_ , \new_[75762]_ ,
    \new_[75763]_ , \new_[75764]_ , \new_[75768]_ , \new_[75769]_ ,
    \new_[75772]_ , \new_[75775]_ , \new_[75776]_ , \new_[75777]_ ,
    \new_[75781]_ , \new_[75782]_ , \new_[75785]_ , \new_[75788]_ ,
    \new_[75789]_ , \new_[75790]_ , \new_[75794]_ , \new_[75795]_ ,
    \new_[75798]_ , \new_[75801]_ , \new_[75802]_ , \new_[75803]_ ,
    \new_[75807]_ , \new_[75808]_ , \new_[75811]_ , \new_[75814]_ ,
    \new_[75815]_ , \new_[75816]_ , \new_[75820]_ , \new_[75821]_ ,
    \new_[75824]_ , \new_[75827]_ , \new_[75828]_ , \new_[75829]_ ,
    \new_[75833]_ , \new_[75834]_ , \new_[75837]_ , \new_[75840]_ ,
    \new_[75841]_ , \new_[75842]_ , \new_[75846]_ , \new_[75847]_ ,
    \new_[75850]_ , \new_[75853]_ , \new_[75854]_ , \new_[75855]_ ,
    \new_[75859]_ , \new_[75860]_ , \new_[75863]_ , \new_[75866]_ ,
    \new_[75867]_ , \new_[75868]_ , \new_[75872]_ , \new_[75873]_ ,
    \new_[75876]_ , \new_[75879]_ , \new_[75880]_ , \new_[75881]_ ,
    \new_[75885]_ , \new_[75886]_ , \new_[75889]_ , \new_[75892]_ ,
    \new_[75893]_ , \new_[75894]_ , \new_[75898]_ , \new_[75899]_ ,
    \new_[75902]_ , \new_[75905]_ , \new_[75906]_ , \new_[75907]_ ,
    \new_[75911]_ , \new_[75912]_ , \new_[75915]_ , \new_[75918]_ ,
    \new_[75919]_ , \new_[75920]_ , \new_[75924]_ , \new_[75925]_ ,
    \new_[75928]_ , \new_[75931]_ , \new_[75932]_ , \new_[75933]_ ,
    \new_[75937]_ , \new_[75938]_ , \new_[75941]_ , \new_[75944]_ ,
    \new_[75945]_ , \new_[75946]_ , \new_[75950]_ , \new_[75951]_ ,
    \new_[75954]_ , \new_[75957]_ , \new_[75958]_ , \new_[75959]_ ,
    \new_[75963]_ , \new_[75964]_ , \new_[75967]_ , \new_[75970]_ ,
    \new_[75971]_ , \new_[75972]_ , \new_[75976]_ , \new_[75977]_ ,
    \new_[75980]_ , \new_[75983]_ , \new_[75984]_ , \new_[75985]_ ,
    \new_[75989]_ , \new_[75990]_ , \new_[75993]_ , \new_[75996]_ ,
    \new_[75997]_ , \new_[75998]_ , \new_[76002]_ , \new_[76003]_ ,
    \new_[76006]_ , \new_[76009]_ , \new_[76010]_ , \new_[76011]_ ,
    \new_[76015]_ , \new_[76016]_ , \new_[76019]_ , \new_[76022]_ ,
    \new_[76023]_ , \new_[76024]_ , \new_[76028]_ , \new_[76029]_ ,
    \new_[76032]_ , \new_[76035]_ , \new_[76036]_ , \new_[76037]_ ,
    \new_[76041]_ , \new_[76042]_ , \new_[76045]_ , \new_[76048]_ ,
    \new_[76049]_ , \new_[76050]_ , \new_[76054]_ , \new_[76055]_ ,
    \new_[76058]_ , \new_[76061]_ , \new_[76062]_ , \new_[76063]_ ,
    \new_[76067]_ , \new_[76068]_ , \new_[76071]_ , \new_[76074]_ ,
    \new_[76075]_ , \new_[76076]_ , \new_[76080]_ , \new_[76081]_ ,
    \new_[76084]_ , \new_[76087]_ , \new_[76088]_ , \new_[76089]_ ,
    \new_[76093]_ , \new_[76094]_ , \new_[76097]_ , \new_[76100]_ ,
    \new_[76101]_ , \new_[76102]_ , \new_[76106]_ , \new_[76107]_ ,
    \new_[76110]_ , \new_[76113]_ , \new_[76114]_ , \new_[76115]_ ,
    \new_[76119]_ , \new_[76120]_ , \new_[76123]_ , \new_[76126]_ ,
    \new_[76127]_ , \new_[76128]_ , \new_[76132]_ , \new_[76133]_ ,
    \new_[76136]_ , \new_[76139]_ , \new_[76140]_ , \new_[76141]_ ,
    \new_[76145]_ , \new_[76146]_ , \new_[76149]_ , \new_[76152]_ ,
    \new_[76153]_ , \new_[76154]_ , \new_[76158]_ , \new_[76159]_ ,
    \new_[76162]_ , \new_[76165]_ , \new_[76166]_ , \new_[76167]_ ,
    \new_[76171]_ , \new_[76172]_ , \new_[76175]_ , \new_[76178]_ ,
    \new_[76179]_ , \new_[76180]_ , \new_[76184]_ , \new_[76185]_ ,
    \new_[76188]_ , \new_[76191]_ , \new_[76192]_ , \new_[76193]_ ,
    \new_[76197]_ , \new_[76198]_ , \new_[76201]_ , \new_[76204]_ ,
    \new_[76205]_ , \new_[76206]_ , \new_[76210]_ , \new_[76211]_ ,
    \new_[76214]_ , \new_[76217]_ , \new_[76218]_ , \new_[76219]_ ,
    \new_[76223]_ , \new_[76224]_ , \new_[76227]_ , \new_[76230]_ ,
    \new_[76231]_ , \new_[76232]_ , \new_[76236]_ , \new_[76237]_ ,
    \new_[76240]_ , \new_[76243]_ , \new_[76244]_ , \new_[76245]_ ,
    \new_[76249]_ , \new_[76250]_ , \new_[76253]_ , \new_[76256]_ ,
    \new_[76257]_ , \new_[76258]_ , \new_[76262]_ , \new_[76263]_ ,
    \new_[76266]_ , \new_[76269]_ , \new_[76270]_ , \new_[76271]_ ,
    \new_[76275]_ , \new_[76276]_ , \new_[76279]_ , \new_[76282]_ ,
    \new_[76283]_ , \new_[76284]_ , \new_[76288]_ , \new_[76289]_ ,
    \new_[76292]_ , \new_[76295]_ , \new_[76296]_ , \new_[76297]_ ,
    \new_[76301]_ , \new_[76302]_ , \new_[76305]_ , \new_[76308]_ ,
    \new_[76309]_ , \new_[76310]_ , \new_[76314]_ , \new_[76315]_ ,
    \new_[76318]_ , \new_[76321]_ , \new_[76322]_ , \new_[76323]_ ,
    \new_[76327]_ , \new_[76328]_ , \new_[76331]_ , \new_[76334]_ ,
    \new_[76335]_ , \new_[76336]_ , \new_[76340]_ , \new_[76341]_ ,
    \new_[76344]_ , \new_[76347]_ , \new_[76348]_ , \new_[76349]_ ,
    \new_[76353]_ , \new_[76354]_ , \new_[76357]_ , \new_[76360]_ ,
    \new_[76361]_ , \new_[76362]_ , \new_[76366]_ , \new_[76367]_ ,
    \new_[76370]_ , \new_[76373]_ , \new_[76374]_ , \new_[76375]_ ,
    \new_[76379]_ , \new_[76380]_ , \new_[76383]_ , \new_[76386]_ ,
    \new_[76387]_ , \new_[76388]_ , \new_[76392]_ , \new_[76393]_ ,
    \new_[76396]_ , \new_[76399]_ , \new_[76400]_ , \new_[76401]_ ,
    \new_[76405]_ , \new_[76406]_ , \new_[76409]_ , \new_[76412]_ ,
    \new_[76413]_ , \new_[76414]_ , \new_[76418]_ , \new_[76419]_ ,
    \new_[76422]_ , \new_[76425]_ , \new_[76426]_ , \new_[76427]_ ,
    \new_[76431]_ , \new_[76432]_ , \new_[76435]_ , \new_[76438]_ ,
    \new_[76439]_ , \new_[76440]_ , \new_[76444]_ , \new_[76445]_ ,
    \new_[76448]_ , \new_[76451]_ , \new_[76452]_ , \new_[76453]_ ,
    \new_[76457]_ , \new_[76458]_ , \new_[76461]_ , \new_[76464]_ ,
    \new_[76465]_ , \new_[76466]_ , \new_[76470]_ , \new_[76471]_ ,
    \new_[76474]_ , \new_[76477]_ , \new_[76478]_ , \new_[76479]_ ,
    \new_[76483]_ , \new_[76484]_ , \new_[76487]_ , \new_[76490]_ ,
    \new_[76491]_ , \new_[76492]_ , \new_[76496]_ , \new_[76497]_ ,
    \new_[76500]_ , \new_[76503]_ , \new_[76504]_ , \new_[76505]_ ,
    \new_[76509]_ , \new_[76510]_ , \new_[76513]_ , \new_[76516]_ ,
    \new_[76517]_ , \new_[76518]_ , \new_[76522]_ , \new_[76523]_ ,
    \new_[76526]_ , \new_[76529]_ , \new_[76530]_ , \new_[76531]_ ,
    \new_[76535]_ , \new_[76536]_ , \new_[76539]_ , \new_[76542]_ ,
    \new_[76543]_ , \new_[76544]_ , \new_[76548]_ , \new_[76549]_ ,
    \new_[76552]_ , \new_[76555]_ , \new_[76556]_ , \new_[76557]_ ,
    \new_[76561]_ , \new_[76562]_ , \new_[76565]_ , \new_[76568]_ ,
    \new_[76569]_ , \new_[76570]_ , \new_[76574]_ , \new_[76575]_ ,
    \new_[76578]_ , \new_[76581]_ , \new_[76582]_ , \new_[76583]_ ,
    \new_[76587]_ , \new_[76588]_ , \new_[76591]_ , \new_[76594]_ ,
    \new_[76595]_ , \new_[76596]_ , \new_[76600]_ , \new_[76601]_ ,
    \new_[76604]_ , \new_[76607]_ , \new_[76608]_ , \new_[76609]_ ,
    \new_[76613]_ , \new_[76614]_ , \new_[76617]_ , \new_[76620]_ ,
    \new_[76621]_ , \new_[76622]_ , \new_[76626]_ , \new_[76627]_ ,
    \new_[76630]_ , \new_[76633]_ , \new_[76634]_ , \new_[76635]_ ,
    \new_[76639]_ , \new_[76640]_ , \new_[76643]_ , \new_[76646]_ ,
    \new_[76647]_ , \new_[76648]_ , \new_[76652]_ , \new_[76653]_ ,
    \new_[76656]_ , \new_[76659]_ , \new_[76660]_ , \new_[76661]_ ,
    \new_[76665]_ , \new_[76666]_ , \new_[76669]_ , \new_[76672]_ ,
    \new_[76673]_ , \new_[76674]_ , \new_[76678]_ , \new_[76679]_ ,
    \new_[76682]_ , \new_[76685]_ , \new_[76686]_ , \new_[76687]_ ,
    \new_[76691]_ , \new_[76692]_ , \new_[76695]_ , \new_[76698]_ ,
    \new_[76699]_ , \new_[76700]_ , \new_[76704]_ , \new_[76705]_ ,
    \new_[76708]_ , \new_[76711]_ , \new_[76712]_ , \new_[76713]_ ,
    \new_[76717]_ , \new_[76718]_ , \new_[76721]_ , \new_[76724]_ ,
    \new_[76725]_ , \new_[76726]_ , \new_[76730]_ , \new_[76731]_ ,
    \new_[76734]_ , \new_[76737]_ , \new_[76738]_ , \new_[76739]_ ,
    \new_[76743]_ , \new_[76744]_ , \new_[76747]_ , \new_[76750]_ ,
    \new_[76751]_ , \new_[76752]_ , \new_[76756]_ , \new_[76757]_ ,
    \new_[76760]_ , \new_[76763]_ , \new_[76764]_ , \new_[76765]_ ,
    \new_[76769]_ , \new_[76770]_ , \new_[76773]_ , \new_[76776]_ ,
    \new_[76777]_ , \new_[76778]_ , \new_[76782]_ , \new_[76783]_ ,
    \new_[76786]_ , \new_[76789]_ , \new_[76790]_ , \new_[76791]_ ,
    \new_[76795]_ , \new_[76796]_ , \new_[76799]_ , \new_[76802]_ ,
    \new_[76803]_ , \new_[76804]_ , \new_[76808]_ , \new_[76809]_ ,
    \new_[76812]_ , \new_[76815]_ , \new_[76816]_ , \new_[76817]_ ,
    \new_[76821]_ , \new_[76822]_ , \new_[76825]_ , \new_[76828]_ ,
    \new_[76829]_ , \new_[76830]_ , \new_[76834]_ , \new_[76835]_ ,
    \new_[76838]_ , \new_[76841]_ , \new_[76842]_ , \new_[76843]_ ,
    \new_[76847]_ , \new_[76848]_ , \new_[76851]_ , \new_[76854]_ ,
    \new_[76855]_ , \new_[76856]_ , \new_[76860]_ , \new_[76861]_ ,
    \new_[76864]_ , \new_[76867]_ , \new_[76868]_ , \new_[76869]_ ,
    \new_[76873]_ , \new_[76874]_ , \new_[76877]_ , \new_[76880]_ ,
    \new_[76881]_ , \new_[76882]_ , \new_[76886]_ , \new_[76887]_ ,
    \new_[76890]_ , \new_[76893]_ , \new_[76894]_ , \new_[76895]_ ,
    \new_[76899]_ , \new_[76900]_ , \new_[76903]_ , \new_[76906]_ ,
    \new_[76907]_ , \new_[76908]_ , \new_[76912]_ , \new_[76913]_ ,
    \new_[76916]_ , \new_[76919]_ , \new_[76920]_ , \new_[76921]_ ,
    \new_[76925]_ , \new_[76926]_ , \new_[76929]_ , \new_[76932]_ ,
    \new_[76933]_ , \new_[76934]_ , \new_[76938]_ , \new_[76939]_ ,
    \new_[76942]_ , \new_[76945]_ , \new_[76946]_ , \new_[76947]_ ,
    \new_[76951]_ , \new_[76952]_ , \new_[76955]_ , \new_[76958]_ ,
    \new_[76959]_ , \new_[76960]_ , \new_[76964]_ , \new_[76965]_ ,
    \new_[76968]_ , \new_[76971]_ , \new_[76972]_ , \new_[76973]_ ,
    \new_[76977]_ , \new_[76978]_ , \new_[76981]_ , \new_[76984]_ ,
    \new_[76985]_ , \new_[76986]_ , \new_[76990]_ , \new_[76991]_ ,
    \new_[76994]_ , \new_[76997]_ , \new_[76998]_ , \new_[76999]_ ,
    \new_[77003]_ , \new_[77004]_ , \new_[77007]_ , \new_[77010]_ ,
    \new_[77011]_ , \new_[77012]_ , \new_[77016]_ , \new_[77017]_ ,
    \new_[77020]_ , \new_[77023]_ , \new_[77024]_ , \new_[77025]_ ,
    \new_[77029]_ , \new_[77030]_ , \new_[77033]_ , \new_[77036]_ ,
    \new_[77037]_ , \new_[77038]_ , \new_[77042]_ , \new_[77043]_ ,
    \new_[77046]_ , \new_[77049]_ , \new_[77050]_ , \new_[77051]_ ,
    \new_[77055]_ , \new_[77056]_ , \new_[77059]_ , \new_[77062]_ ,
    \new_[77063]_ , \new_[77064]_ , \new_[77068]_ , \new_[77069]_ ,
    \new_[77072]_ , \new_[77075]_ , \new_[77076]_ , \new_[77077]_ ,
    \new_[77081]_ , \new_[77082]_ , \new_[77085]_ , \new_[77088]_ ,
    \new_[77089]_ , \new_[77090]_ , \new_[77094]_ , \new_[77095]_ ,
    \new_[77098]_ , \new_[77101]_ , \new_[77102]_ , \new_[77103]_ ,
    \new_[77107]_ , \new_[77108]_ , \new_[77111]_ , \new_[77114]_ ,
    \new_[77115]_ , \new_[77116]_ , \new_[77120]_ , \new_[77121]_ ,
    \new_[77124]_ , \new_[77127]_ , \new_[77128]_ , \new_[77129]_ ,
    \new_[77133]_ , \new_[77134]_ , \new_[77137]_ , \new_[77140]_ ,
    \new_[77141]_ , \new_[77142]_ , \new_[77146]_ , \new_[77147]_ ,
    \new_[77150]_ , \new_[77153]_ , \new_[77154]_ , \new_[77155]_ ,
    \new_[77159]_ , \new_[77160]_ , \new_[77163]_ , \new_[77166]_ ,
    \new_[77167]_ , \new_[77168]_ , \new_[77172]_ , \new_[77173]_ ,
    \new_[77176]_ , \new_[77179]_ , \new_[77180]_ , \new_[77181]_ ,
    \new_[77185]_ , \new_[77186]_ , \new_[77189]_ , \new_[77192]_ ,
    \new_[77193]_ , \new_[77194]_ , \new_[77198]_ , \new_[77199]_ ,
    \new_[77202]_ , \new_[77205]_ , \new_[77206]_ , \new_[77207]_ ,
    \new_[77211]_ , \new_[77212]_ , \new_[77215]_ , \new_[77218]_ ,
    \new_[77219]_ , \new_[77220]_ , \new_[77224]_ , \new_[77225]_ ,
    \new_[77228]_ , \new_[77231]_ , \new_[77232]_ , \new_[77233]_ ,
    \new_[77237]_ , \new_[77238]_ , \new_[77241]_ , \new_[77244]_ ,
    \new_[77245]_ , \new_[77246]_ , \new_[77250]_ , \new_[77251]_ ,
    \new_[77254]_ , \new_[77257]_ , \new_[77258]_ , \new_[77259]_ ,
    \new_[77263]_ , \new_[77264]_ , \new_[77267]_ , \new_[77270]_ ,
    \new_[77271]_ , \new_[77272]_ , \new_[77276]_ , \new_[77277]_ ,
    \new_[77280]_ , \new_[77283]_ , \new_[77284]_ , \new_[77285]_ ,
    \new_[77289]_ , \new_[77290]_ , \new_[77293]_ , \new_[77296]_ ,
    \new_[77297]_ , \new_[77298]_ , \new_[77302]_ , \new_[77303]_ ,
    \new_[77306]_ , \new_[77309]_ , \new_[77310]_ , \new_[77311]_ ,
    \new_[77315]_ , \new_[77316]_ , \new_[77319]_ , \new_[77322]_ ,
    \new_[77323]_ , \new_[77324]_ , \new_[77328]_ , \new_[77329]_ ,
    \new_[77332]_ , \new_[77335]_ , \new_[77336]_ , \new_[77337]_ ,
    \new_[77341]_ , \new_[77342]_ , \new_[77345]_ , \new_[77348]_ ,
    \new_[77349]_ , \new_[77350]_ , \new_[77354]_ , \new_[77355]_ ,
    \new_[77358]_ , \new_[77361]_ , \new_[77362]_ , \new_[77363]_ ,
    \new_[77367]_ , \new_[77368]_ , \new_[77371]_ , \new_[77374]_ ,
    \new_[77375]_ , \new_[77376]_ , \new_[77380]_ , \new_[77381]_ ,
    \new_[77384]_ , \new_[77387]_ , \new_[77388]_ , \new_[77389]_ ,
    \new_[77393]_ , \new_[77394]_ , \new_[77397]_ , \new_[77400]_ ,
    \new_[77401]_ , \new_[77402]_ , \new_[77406]_ , \new_[77407]_ ,
    \new_[77410]_ , \new_[77413]_ , \new_[77414]_ , \new_[77415]_ ,
    \new_[77419]_ , \new_[77420]_ , \new_[77423]_ , \new_[77426]_ ,
    \new_[77427]_ , \new_[77428]_ , \new_[77432]_ , \new_[77433]_ ,
    \new_[77436]_ , \new_[77439]_ , \new_[77440]_ , \new_[77441]_ ,
    \new_[77445]_ , \new_[77446]_ , \new_[77449]_ , \new_[77452]_ ,
    \new_[77453]_ , \new_[77454]_ , \new_[77458]_ , \new_[77459]_ ,
    \new_[77462]_ , \new_[77465]_ , \new_[77466]_ , \new_[77467]_ ,
    \new_[77471]_ , \new_[77472]_ , \new_[77475]_ , \new_[77478]_ ,
    \new_[77479]_ , \new_[77480]_ , \new_[77484]_ , \new_[77485]_ ,
    \new_[77488]_ , \new_[77491]_ , \new_[77492]_ , \new_[77493]_ ,
    \new_[77497]_ , \new_[77498]_ , \new_[77501]_ , \new_[77504]_ ,
    \new_[77505]_ , \new_[77506]_ , \new_[77510]_ , \new_[77511]_ ,
    \new_[77514]_ , \new_[77517]_ , \new_[77518]_ , \new_[77519]_ ,
    \new_[77523]_ , \new_[77524]_ , \new_[77527]_ , \new_[77530]_ ,
    \new_[77531]_ , \new_[77532]_ , \new_[77536]_ , \new_[77537]_ ,
    \new_[77540]_ , \new_[77543]_ , \new_[77544]_ , \new_[77545]_ ,
    \new_[77549]_ , \new_[77550]_ , \new_[77553]_ , \new_[77556]_ ,
    \new_[77557]_ , \new_[77558]_ , \new_[77562]_ , \new_[77563]_ ,
    \new_[77566]_ , \new_[77569]_ , \new_[77570]_ , \new_[77571]_ ,
    \new_[77575]_ , \new_[77576]_ , \new_[77579]_ , \new_[77582]_ ,
    \new_[77583]_ , \new_[77584]_ , \new_[77588]_ , \new_[77589]_ ,
    \new_[77592]_ , \new_[77595]_ , \new_[77596]_ , \new_[77597]_ ,
    \new_[77601]_ , \new_[77602]_ , \new_[77605]_ , \new_[77608]_ ,
    \new_[77609]_ , \new_[77610]_ , \new_[77614]_ , \new_[77615]_ ,
    \new_[77618]_ , \new_[77621]_ , \new_[77622]_ , \new_[77623]_ ,
    \new_[77627]_ , \new_[77628]_ , \new_[77631]_ , \new_[77634]_ ,
    \new_[77635]_ , \new_[77636]_ , \new_[77640]_ , \new_[77641]_ ,
    \new_[77644]_ , \new_[77647]_ , \new_[77648]_ , \new_[77649]_ ,
    \new_[77652]_ , \new_[77655]_ , \new_[77656]_ , \new_[77659]_ ,
    \new_[77662]_ , \new_[77663]_ , \new_[77664]_ , \new_[77668]_ ,
    \new_[77669]_ , \new_[77672]_ , \new_[77675]_ , \new_[77676]_ ,
    \new_[77677]_ , \new_[77680]_ , \new_[77683]_ , \new_[77684]_ ,
    \new_[77687]_ , \new_[77690]_ , \new_[77691]_ , \new_[77692]_ ,
    \new_[77696]_ , \new_[77697]_ , \new_[77700]_ , \new_[77703]_ ,
    \new_[77704]_ , \new_[77705]_ , \new_[77708]_ , \new_[77711]_ ,
    \new_[77712]_ , \new_[77715]_ , \new_[77718]_ , \new_[77719]_ ,
    \new_[77720]_ , \new_[77724]_ , \new_[77725]_ , \new_[77728]_ ,
    \new_[77731]_ , \new_[77732]_ , \new_[77733]_ , \new_[77736]_ ,
    \new_[77739]_ , \new_[77740]_ , \new_[77743]_ , \new_[77746]_ ,
    \new_[77747]_ , \new_[77748]_ , \new_[77752]_ , \new_[77753]_ ,
    \new_[77756]_ , \new_[77759]_ , \new_[77760]_ , \new_[77761]_ ,
    \new_[77764]_ , \new_[77767]_ , \new_[77768]_ , \new_[77771]_ ,
    \new_[77774]_ , \new_[77775]_ , \new_[77776]_ , \new_[77780]_ ,
    \new_[77781]_ , \new_[77784]_ , \new_[77787]_ , \new_[77788]_ ,
    \new_[77789]_ , \new_[77792]_ , \new_[77795]_ , \new_[77796]_ ,
    \new_[77799]_ , \new_[77802]_ , \new_[77803]_ , \new_[77804]_ ,
    \new_[77808]_ , \new_[77809]_ , \new_[77812]_ , \new_[77815]_ ,
    \new_[77816]_ , \new_[77817]_ , \new_[77820]_ , \new_[77823]_ ,
    \new_[77824]_ , \new_[77827]_ , \new_[77830]_ , \new_[77831]_ ,
    \new_[77832]_ , \new_[77836]_ , \new_[77837]_ , \new_[77840]_ ,
    \new_[77843]_ , \new_[77844]_ , \new_[77845]_ , \new_[77848]_ ,
    \new_[77851]_ , \new_[77852]_ , \new_[77855]_ , \new_[77858]_ ,
    \new_[77859]_ , \new_[77860]_ , \new_[77864]_ , \new_[77865]_ ,
    \new_[77868]_ , \new_[77871]_ , \new_[77872]_ , \new_[77873]_ ,
    \new_[77876]_ , \new_[77879]_ , \new_[77880]_ , \new_[77883]_ ,
    \new_[77886]_ , \new_[77887]_ , \new_[77888]_ , \new_[77892]_ ,
    \new_[77893]_ , \new_[77896]_ , \new_[77899]_ , \new_[77900]_ ,
    \new_[77901]_ , \new_[77904]_ , \new_[77907]_ , \new_[77908]_ ,
    \new_[77911]_ , \new_[77914]_ , \new_[77915]_ , \new_[77916]_ ,
    \new_[77920]_ , \new_[77921]_ , \new_[77924]_ , \new_[77927]_ ,
    \new_[77928]_ , \new_[77929]_ , \new_[77932]_ , \new_[77935]_ ,
    \new_[77936]_ , \new_[77939]_ , \new_[77942]_ , \new_[77943]_ ,
    \new_[77944]_ , \new_[77948]_ , \new_[77949]_ , \new_[77952]_ ,
    \new_[77955]_ , \new_[77956]_ , \new_[77957]_ , \new_[77960]_ ,
    \new_[77963]_ , \new_[77964]_ , \new_[77967]_ , \new_[77970]_ ,
    \new_[77971]_ , \new_[77972]_ , \new_[77976]_ , \new_[77977]_ ,
    \new_[77980]_ , \new_[77983]_ , \new_[77984]_ , \new_[77985]_ ,
    \new_[77988]_ , \new_[77991]_ , \new_[77992]_ , \new_[77995]_ ,
    \new_[77998]_ , \new_[77999]_ , \new_[78000]_ , \new_[78004]_ ,
    \new_[78005]_ , \new_[78008]_ , \new_[78011]_ , \new_[78012]_ ,
    \new_[78013]_ , \new_[78016]_ , \new_[78019]_ , \new_[78020]_ ,
    \new_[78023]_ , \new_[78026]_ , \new_[78027]_ , \new_[78028]_ ,
    \new_[78032]_ , \new_[78033]_ , \new_[78036]_ , \new_[78039]_ ,
    \new_[78040]_ , \new_[78041]_ , \new_[78044]_ , \new_[78047]_ ,
    \new_[78048]_ , \new_[78051]_ , \new_[78054]_ , \new_[78055]_ ,
    \new_[78056]_ , \new_[78060]_ , \new_[78061]_ , \new_[78064]_ ,
    \new_[78067]_ , \new_[78068]_ , \new_[78069]_ , \new_[78072]_ ,
    \new_[78075]_ , \new_[78076]_ , \new_[78079]_ , \new_[78082]_ ,
    \new_[78083]_ , \new_[78084]_ , \new_[78088]_ , \new_[78089]_ ,
    \new_[78092]_ , \new_[78095]_ , \new_[78096]_ , \new_[78097]_ ,
    \new_[78100]_ , \new_[78103]_ , \new_[78104]_ , \new_[78107]_ ,
    \new_[78110]_ , \new_[78111]_ , \new_[78112]_ , \new_[78116]_ ,
    \new_[78117]_ , \new_[78120]_ , \new_[78123]_ , \new_[78124]_ ,
    \new_[78125]_ , \new_[78128]_ , \new_[78131]_ , \new_[78132]_ ,
    \new_[78135]_ , \new_[78138]_ , \new_[78139]_ , \new_[78140]_ ,
    \new_[78144]_ , \new_[78145]_ , \new_[78148]_ , \new_[78151]_ ,
    \new_[78152]_ , \new_[78153]_ , \new_[78156]_ , \new_[78159]_ ,
    \new_[78160]_ , \new_[78163]_ , \new_[78166]_ , \new_[78167]_ ,
    \new_[78168]_ , \new_[78172]_ , \new_[78173]_ , \new_[78176]_ ,
    \new_[78179]_ , \new_[78180]_ , \new_[78181]_ , \new_[78184]_ ,
    \new_[78187]_ , \new_[78188]_ , \new_[78191]_ , \new_[78194]_ ,
    \new_[78195]_ , \new_[78196]_ , \new_[78200]_ , \new_[78201]_ ,
    \new_[78204]_ , \new_[78207]_ , \new_[78208]_ , \new_[78209]_ ,
    \new_[78212]_ , \new_[78215]_ , \new_[78216]_ , \new_[78219]_ ,
    \new_[78222]_ , \new_[78223]_ , \new_[78224]_ , \new_[78228]_ ,
    \new_[78229]_ , \new_[78232]_ , \new_[78235]_ , \new_[78236]_ ,
    \new_[78237]_ , \new_[78240]_ , \new_[78243]_ , \new_[78244]_ ,
    \new_[78247]_ , \new_[78250]_ , \new_[78251]_ , \new_[78252]_ ,
    \new_[78256]_ , \new_[78257]_ , \new_[78260]_ , \new_[78263]_ ,
    \new_[78264]_ , \new_[78265]_ , \new_[78268]_ , \new_[78271]_ ,
    \new_[78272]_ , \new_[78275]_ , \new_[78278]_ , \new_[78279]_ ,
    \new_[78280]_ , \new_[78284]_ , \new_[78285]_ , \new_[78288]_ ,
    \new_[78291]_ , \new_[78292]_ , \new_[78293]_ , \new_[78296]_ ,
    \new_[78299]_ , \new_[78300]_ , \new_[78303]_ , \new_[78306]_ ,
    \new_[78307]_ , \new_[78308]_ , \new_[78312]_ , \new_[78313]_ ,
    \new_[78316]_ , \new_[78319]_ , \new_[78320]_ , \new_[78321]_ ,
    \new_[78324]_ , \new_[78327]_ , \new_[78328]_ , \new_[78331]_ ,
    \new_[78334]_ , \new_[78335]_ , \new_[78336]_ , \new_[78340]_ ,
    \new_[78341]_ , \new_[78344]_ , \new_[78347]_ , \new_[78348]_ ,
    \new_[78349]_ , \new_[78352]_ , \new_[78355]_ , \new_[78356]_ ,
    \new_[78359]_ , \new_[78362]_ , \new_[78363]_ , \new_[78364]_ ,
    \new_[78368]_ , \new_[78369]_ , \new_[78372]_ , \new_[78375]_ ,
    \new_[78376]_ , \new_[78377]_ , \new_[78380]_ , \new_[78383]_ ,
    \new_[78384]_ , \new_[78387]_ , \new_[78390]_ , \new_[78391]_ ,
    \new_[78392]_ , \new_[78396]_ , \new_[78397]_ , \new_[78400]_ ,
    \new_[78403]_ , \new_[78404]_ , \new_[78405]_ , \new_[78408]_ ,
    \new_[78411]_ , \new_[78412]_ , \new_[78415]_ , \new_[78418]_ ,
    \new_[78419]_ , \new_[78420]_ , \new_[78424]_ , \new_[78425]_ ,
    \new_[78428]_ , \new_[78431]_ , \new_[78432]_ , \new_[78433]_ ,
    \new_[78436]_ , \new_[78439]_ , \new_[78440]_ , \new_[78443]_ ,
    \new_[78446]_ , \new_[78447]_ , \new_[78448]_ , \new_[78452]_ ,
    \new_[78453]_ , \new_[78456]_ , \new_[78459]_ , \new_[78460]_ ,
    \new_[78461]_ , \new_[78464]_ , \new_[78467]_ , \new_[78468]_ ,
    \new_[78471]_ , \new_[78474]_ , \new_[78475]_ , \new_[78476]_ ,
    \new_[78480]_ , \new_[78481]_ , \new_[78484]_ , \new_[78487]_ ,
    \new_[78488]_ , \new_[78489]_ , \new_[78492]_ , \new_[78495]_ ,
    \new_[78496]_ , \new_[78499]_ , \new_[78502]_ , \new_[78503]_ ,
    \new_[78504]_ , \new_[78508]_ , \new_[78509]_ , \new_[78512]_ ,
    \new_[78515]_ , \new_[78516]_ , \new_[78517]_ , \new_[78520]_ ,
    \new_[78523]_ , \new_[78524]_ , \new_[78527]_ , \new_[78530]_ ,
    \new_[78531]_ , \new_[78532]_ , \new_[78536]_ , \new_[78537]_ ,
    \new_[78540]_ , \new_[78543]_ , \new_[78544]_ , \new_[78545]_ ,
    \new_[78548]_ , \new_[78551]_ , \new_[78552]_ , \new_[78555]_ ,
    \new_[78558]_ , \new_[78559]_ , \new_[78560]_ , \new_[78564]_ ,
    \new_[78565]_ , \new_[78568]_ , \new_[78571]_ , \new_[78572]_ ,
    \new_[78573]_ , \new_[78576]_ , \new_[78579]_ , \new_[78580]_ ,
    \new_[78583]_ , \new_[78586]_ , \new_[78587]_ , \new_[78588]_ ,
    \new_[78592]_ , \new_[78593]_ , \new_[78596]_ , \new_[78599]_ ,
    \new_[78600]_ , \new_[78601]_ , \new_[78604]_ , \new_[78607]_ ,
    \new_[78608]_ , \new_[78611]_ , \new_[78614]_ , \new_[78615]_ ,
    \new_[78616]_ , \new_[78620]_ , \new_[78621]_ , \new_[78624]_ ,
    \new_[78627]_ , \new_[78628]_ , \new_[78629]_ , \new_[78632]_ ,
    \new_[78635]_ , \new_[78636]_ , \new_[78639]_ , \new_[78642]_ ,
    \new_[78643]_ , \new_[78644]_ , \new_[78648]_ , \new_[78649]_ ,
    \new_[78652]_ , \new_[78655]_ , \new_[78656]_ , \new_[78657]_ ,
    \new_[78660]_ , \new_[78663]_ , \new_[78664]_ , \new_[78667]_ ,
    \new_[78670]_ , \new_[78671]_ , \new_[78672]_ , \new_[78676]_ ,
    \new_[78677]_ , \new_[78680]_ , \new_[78683]_ , \new_[78684]_ ,
    \new_[78685]_ , \new_[78688]_ , \new_[78691]_ , \new_[78692]_ ,
    \new_[78695]_ , \new_[78698]_ , \new_[78699]_ , \new_[78700]_ ,
    \new_[78704]_ , \new_[78705]_ , \new_[78708]_ , \new_[78711]_ ,
    \new_[78712]_ , \new_[78713]_ , \new_[78716]_ , \new_[78719]_ ,
    \new_[78720]_ , \new_[78723]_ , \new_[78726]_ , \new_[78727]_ ,
    \new_[78728]_ , \new_[78732]_ , \new_[78733]_ , \new_[78736]_ ,
    \new_[78739]_ , \new_[78740]_ , \new_[78741]_ , \new_[78744]_ ,
    \new_[78747]_ , \new_[78748]_ , \new_[78751]_ , \new_[78754]_ ,
    \new_[78755]_ , \new_[78756]_ , \new_[78760]_ , \new_[78761]_ ,
    \new_[78764]_ , \new_[78767]_ , \new_[78768]_ , \new_[78769]_ ,
    \new_[78772]_ , \new_[78775]_ , \new_[78776]_ , \new_[78779]_ ,
    \new_[78782]_ , \new_[78783]_ , \new_[78784]_ , \new_[78788]_ ,
    \new_[78789]_ , \new_[78792]_ , \new_[78795]_ , \new_[78796]_ ,
    \new_[78797]_ , \new_[78800]_ , \new_[78803]_ , \new_[78804]_ ,
    \new_[78807]_ , \new_[78810]_ , \new_[78811]_ , \new_[78812]_ ,
    \new_[78816]_ , \new_[78817]_ , \new_[78820]_ , \new_[78823]_ ,
    \new_[78824]_ , \new_[78825]_ , \new_[78828]_ , \new_[78831]_ ,
    \new_[78832]_ , \new_[78835]_ , \new_[78838]_ , \new_[78839]_ ,
    \new_[78840]_ , \new_[78844]_ , \new_[78845]_ , \new_[78848]_ ,
    \new_[78851]_ , \new_[78852]_ , \new_[78853]_ , \new_[78856]_ ,
    \new_[78859]_ , \new_[78860]_ , \new_[78863]_ , \new_[78866]_ ,
    \new_[78867]_ , \new_[78868]_ , \new_[78872]_ , \new_[78873]_ ,
    \new_[78876]_ , \new_[78879]_ , \new_[78880]_ , \new_[78881]_ ,
    \new_[78884]_ , \new_[78887]_ , \new_[78888]_ , \new_[78891]_ ,
    \new_[78894]_ , \new_[78895]_ , \new_[78896]_ , \new_[78900]_ ,
    \new_[78901]_ , \new_[78904]_ , \new_[78907]_ , \new_[78908]_ ,
    \new_[78909]_ , \new_[78912]_ , \new_[78915]_ , \new_[78916]_ ,
    \new_[78919]_ , \new_[78922]_ , \new_[78923]_ , \new_[78924]_ ,
    \new_[78928]_ , \new_[78929]_ , \new_[78932]_ , \new_[78935]_ ,
    \new_[78936]_ , \new_[78937]_ , \new_[78940]_ , \new_[78943]_ ,
    \new_[78944]_ , \new_[78947]_ , \new_[78950]_ , \new_[78951]_ ,
    \new_[78952]_ , \new_[78956]_ , \new_[78957]_ , \new_[78960]_ ,
    \new_[78963]_ , \new_[78964]_ , \new_[78965]_ , \new_[78968]_ ,
    \new_[78971]_ , \new_[78972]_ , \new_[78975]_ , \new_[78978]_ ,
    \new_[78979]_ , \new_[78980]_ , \new_[78984]_ , \new_[78985]_ ,
    \new_[78988]_ , \new_[78991]_ , \new_[78992]_ , \new_[78993]_ ,
    \new_[78996]_ , \new_[78999]_ , \new_[79000]_ , \new_[79003]_ ,
    \new_[79006]_ , \new_[79007]_ , \new_[79008]_ , \new_[79012]_ ,
    \new_[79013]_ , \new_[79016]_ , \new_[79019]_ , \new_[79020]_ ,
    \new_[79021]_ , \new_[79024]_ , \new_[79027]_ , \new_[79028]_ ,
    \new_[79031]_ , \new_[79034]_ , \new_[79035]_ , \new_[79036]_ ,
    \new_[79040]_ , \new_[79041]_ , \new_[79044]_ , \new_[79047]_ ,
    \new_[79048]_ , \new_[79049]_ , \new_[79052]_ , \new_[79055]_ ,
    \new_[79056]_ , \new_[79059]_ , \new_[79062]_ , \new_[79063]_ ,
    \new_[79064]_ , \new_[79068]_ , \new_[79069]_ , \new_[79072]_ ,
    \new_[79075]_ , \new_[79076]_ , \new_[79077]_ , \new_[79080]_ ,
    \new_[79083]_ , \new_[79084]_ , \new_[79087]_ , \new_[79090]_ ,
    \new_[79091]_ , \new_[79092]_ , \new_[79096]_ , \new_[79097]_ ,
    \new_[79100]_ , \new_[79103]_ , \new_[79104]_ , \new_[79105]_ ,
    \new_[79108]_ , \new_[79111]_ , \new_[79112]_ , \new_[79115]_ ,
    \new_[79118]_ , \new_[79119]_ , \new_[79120]_ , \new_[79124]_ ,
    \new_[79125]_ , \new_[79128]_ , \new_[79131]_ , \new_[79132]_ ,
    \new_[79133]_ , \new_[79136]_ , \new_[79139]_ , \new_[79140]_ ,
    \new_[79143]_ , \new_[79146]_ , \new_[79147]_ , \new_[79148]_ ,
    \new_[79152]_ , \new_[79153]_ , \new_[79156]_ , \new_[79159]_ ,
    \new_[79160]_ , \new_[79161]_ , \new_[79164]_ , \new_[79167]_ ,
    \new_[79168]_ , \new_[79171]_ , \new_[79174]_ , \new_[79175]_ ,
    \new_[79176]_ , \new_[79180]_ , \new_[79181]_ , \new_[79184]_ ,
    \new_[79187]_ , \new_[79188]_ , \new_[79189]_ , \new_[79192]_ ,
    \new_[79195]_ , \new_[79196]_ , \new_[79199]_ , \new_[79202]_ ,
    \new_[79203]_ , \new_[79204]_ , \new_[79208]_ , \new_[79209]_ ,
    \new_[79212]_ , \new_[79215]_ , \new_[79216]_ , \new_[79217]_ ,
    \new_[79220]_ , \new_[79223]_ , \new_[79224]_ , \new_[79227]_ ,
    \new_[79230]_ , \new_[79231]_ , \new_[79232]_ , \new_[79236]_ ,
    \new_[79237]_ , \new_[79240]_ , \new_[79243]_ , \new_[79244]_ ,
    \new_[79245]_ , \new_[79248]_ , \new_[79251]_ , \new_[79252]_ ,
    \new_[79255]_ , \new_[79258]_ , \new_[79259]_ , \new_[79260]_ ,
    \new_[79264]_ , \new_[79265]_ , \new_[79268]_ , \new_[79271]_ ,
    \new_[79272]_ , \new_[79273]_ , \new_[79276]_ , \new_[79279]_ ,
    \new_[79280]_ , \new_[79283]_ , \new_[79286]_ , \new_[79287]_ ,
    \new_[79288]_ , \new_[79292]_ , \new_[79293]_ , \new_[79296]_ ,
    \new_[79299]_ , \new_[79300]_ , \new_[79301]_ , \new_[79304]_ ,
    \new_[79307]_ , \new_[79308]_ , \new_[79311]_ , \new_[79314]_ ,
    \new_[79315]_ , \new_[79316]_ , \new_[79320]_ , \new_[79321]_ ,
    \new_[79324]_ , \new_[79327]_ , \new_[79328]_ , \new_[79329]_ ,
    \new_[79332]_ , \new_[79335]_ , \new_[79336]_ , \new_[79339]_ ,
    \new_[79342]_ , \new_[79343]_ , \new_[79344]_ , \new_[79348]_ ,
    \new_[79349]_ , \new_[79352]_ , \new_[79355]_ , \new_[79356]_ ,
    \new_[79357]_ , \new_[79360]_ , \new_[79363]_ , \new_[79364]_ ,
    \new_[79367]_ , \new_[79370]_ , \new_[79371]_ , \new_[79372]_ ,
    \new_[79376]_ , \new_[79377]_ , \new_[79380]_ , \new_[79383]_ ,
    \new_[79384]_ , \new_[79385]_ , \new_[79388]_ , \new_[79391]_ ,
    \new_[79392]_ , \new_[79395]_ , \new_[79398]_ , \new_[79399]_ ,
    \new_[79400]_ , \new_[79404]_ , \new_[79405]_ , \new_[79408]_ ,
    \new_[79411]_ , \new_[79412]_ , \new_[79413]_ , \new_[79416]_ ,
    \new_[79419]_ , \new_[79420]_ , \new_[79423]_ , \new_[79426]_ ,
    \new_[79427]_ , \new_[79428]_ , \new_[79432]_ , \new_[79433]_ ,
    \new_[79436]_ , \new_[79439]_ , \new_[79440]_ , \new_[79441]_ ,
    \new_[79444]_ , \new_[79447]_ , \new_[79448]_ , \new_[79451]_ ,
    \new_[79454]_ , \new_[79455]_ , \new_[79456]_ , \new_[79460]_ ,
    \new_[79461]_ , \new_[79464]_ , \new_[79467]_ , \new_[79468]_ ,
    \new_[79469]_ , \new_[79472]_ , \new_[79475]_ , \new_[79476]_ ,
    \new_[79479]_ , \new_[79482]_ , \new_[79483]_ , \new_[79484]_ ,
    \new_[79488]_ , \new_[79489]_ , \new_[79492]_ , \new_[79495]_ ,
    \new_[79496]_ , \new_[79497]_ , \new_[79500]_ , \new_[79503]_ ,
    \new_[79504]_ , \new_[79507]_ , \new_[79510]_ , \new_[79511]_ ,
    \new_[79512]_ , \new_[79516]_ , \new_[79517]_ , \new_[79520]_ ,
    \new_[79523]_ , \new_[79524]_ , \new_[79525]_ , \new_[79528]_ ,
    \new_[79531]_ , \new_[79532]_ , \new_[79535]_ , \new_[79538]_ ,
    \new_[79539]_ , \new_[79540]_ , \new_[79544]_ , \new_[79545]_ ,
    \new_[79548]_ , \new_[79551]_ , \new_[79552]_ , \new_[79553]_ ,
    \new_[79556]_ , \new_[79559]_ , \new_[79560]_ , \new_[79563]_ ,
    \new_[79566]_ , \new_[79567]_ , \new_[79568]_ , \new_[79572]_ ,
    \new_[79573]_ , \new_[79576]_ , \new_[79579]_ , \new_[79580]_ ,
    \new_[79581]_ , \new_[79584]_ , \new_[79587]_ , \new_[79588]_ ,
    \new_[79591]_ , \new_[79594]_ , \new_[79595]_ , \new_[79596]_ ,
    \new_[79600]_ , \new_[79601]_ , \new_[79604]_ , \new_[79607]_ ,
    \new_[79608]_ , \new_[79609]_ , \new_[79612]_ , \new_[79615]_ ,
    \new_[79616]_ , \new_[79619]_ , \new_[79622]_ , \new_[79623]_ ,
    \new_[79624]_ , \new_[79628]_ , \new_[79629]_ , \new_[79632]_ ,
    \new_[79635]_ , \new_[79636]_ , \new_[79637]_ , \new_[79640]_ ,
    \new_[79643]_ , \new_[79644]_ , \new_[79647]_ , \new_[79650]_ ,
    \new_[79651]_ , \new_[79652]_ , \new_[79656]_ , \new_[79657]_ ,
    \new_[79660]_ , \new_[79663]_ , \new_[79664]_ , \new_[79665]_ ,
    \new_[79668]_ , \new_[79671]_ , \new_[79672]_ , \new_[79675]_ ,
    \new_[79678]_ , \new_[79679]_ , \new_[79680]_ , \new_[79684]_ ,
    \new_[79685]_ , \new_[79688]_ , \new_[79691]_ , \new_[79692]_ ,
    \new_[79693]_ , \new_[79696]_ , \new_[79699]_ , \new_[79700]_ ,
    \new_[79703]_ , \new_[79706]_ , \new_[79707]_ , \new_[79708]_ ,
    \new_[79712]_ , \new_[79713]_ , \new_[79716]_ , \new_[79719]_ ,
    \new_[79720]_ , \new_[79721]_ , \new_[79724]_ , \new_[79727]_ ,
    \new_[79728]_ , \new_[79731]_ , \new_[79734]_ , \new_[79735]_ ,
    \new_[79736]_ , \new_[79740]_ , \new_[79741]_ , \new_[79744]_ ,
    \new_[79747]_ , \new_[79748]_ , \new_[79749]_ , \new_[79752]_ ,
    \new_[79755]_ , \new_[79756]_ , \new_[79759]_ , \new_[79762]_ ,
    \new_[79763]_ , \new_[79764]_ , \new_[79768]_ , \new_[79769]_ ,
    \new_[79772]_ , \new_[79775]_ , \new_[79776]_ , \new_[79777]_ ,
    \new_[79780]_ , \new_[79783]_ , \new_[79784]_ , \new_[79787]_ ,
    \new_[79790]_ , \new_[79791]_ , \new_[79792]_ , \new_[79796]_ ,
    \new_[79797]_ , \new_[79800]_ , \new_[79803]_ , \new_[79804]_ ,
    \new_[79805]_ , \new_[79808]_ , \new_[79811]_ , \new_[79812]_ ,
    \new_[79815]_ , \new_[79818]_ , \new_[79819]_ , \new_[79820]_ ,
    \new_[79824]_ , \new_[79825]_ , \new_[79828]_ , \new_[79831]_ ,
    \new_[79832]_ , \new_[79833]_ , \new_[79836]_ , \new_[79839]_ ,
    \new_[79840]_ , \new_[79843]_ , \new_[79846]_ , \new_[79847]_ ,
    \new_[79848]_ , \new_[79852]_ , \new_[79853]_ , \new_[79856]_ ,
    \new_[79859]_ , \new_[79860]_ , \new_[79861]_ , \new_[79864]_ ,
    \new_[79867]_ , \new_[79868]_ , \new_[79871]_ , \new_[79874]_ ,
    \new_[79875]_ , \new_[79876]_ , \new_[79880]_ , \new_[79881]_ ,
    \new_[79884]_ , \new_[79887]_ , \new_[79888]_ , \new_[79889]_ ,
    \new_[79892]_ , \new_[79895]_ , \new_[79896]_ , \new_[79899]_ ,
    \new_[79902]_ , \new_[79903]_ , \new_[79904]_ , \new_[79908]_ ,
    \new_[79909]_ , \new_[79912]_ , \new_[79915]_ , \new_[79916]_ ,
    \new_[79917]_ , \new_[79920]_ , \new_[79923]_ , \new_[79924]_ ,
    \new_[79927]_ , \new_[79930]_ , \new_[79931]_ , \new_[79932]_ ,
    \new_[79936]_ , \new_[79937]_ , \new_[79940]_ , \new_[79943]_ ,
    \new_[79944]_ , \new_[79945]_ , \new_[79948]_ , \new_[79951]_ ,
    \new_[79952]_ , \new_[79955]_ , \new_[79958]_ , \new_[79959]_ ,
    \new_[79960]_ , \new_[79964]_ , \new_[79965]_ , \new_[79968]_ ,
    \new_[79971]_ , \new_[79972]_ , \new_[79973]_ , \new_[79976]_ ,
    \new_[79979]_ , \new_[79980]_ , \new_[79983]_ , \new_[79986]_ ,
    \new_[79987]_ , \new_[79988]_ , \new_[79992]_ , \new_[79993]_ ,
    \new_[79996]_ , \new_[79999]_ , \new_[80000]_ , \new_[80001]_ ,
    \new_[80004]_ , \new_[80007]_ , \new_[80008]_ , \new_[80011]_ ,
    \new_[80014]_ , \new_[80015]_ , \new_[80016]_ , \new_[80020]_ ,
    \new_[80021]_ , \new_[80024]_ , \new_[80027]_ , \new_[80028]_ ,
    \new_[80029]_ , \new_[80032]_ , \new_[80035]_ , \new_[80036]_ ,
    \new_[80039]_ , \new_[80042]_ , \new_[80043]_ , \new_[80044]_ ,
    \new_[80048]_ , \new_[80049]_ , \new_[80052]_ , \new_[80055]_ ,
    \new_[80056]_ , \new_[80057]_ , \new_[80060]_ , \new_[80063]_ ,
    \new_[80064]_ , \new_[80067]_ , \new_[80070]_ , \new_[80071]_ ,
    \new_[80072]_ , \new_[80076]_ , \new_[80077]_ , \new_[80080]_ ,
    \new_[80083]_ , \new_[80084]_ , \new_[80085]_ , \new_[80088]_ ,
    \new_[80091]_ , \new_[80092]_ , \new_[80095]_ , \new_[80098]_ ,
    \new_[80099]_ , \new_[80100]_ , \new_[80104]_ , \new_[80105]_ ,
    \new_[80108]_ , \new_[80111]_ , \new_[80112]_ , \new_[80113]_ ,
    \new_[80116]_ , \new_[80119]_ , \new_[80120]_ , \new_[80123]_ ,
    \new_[80126]_ , \new_[80127]_ , \new_[80128]_ , \new_[80132]_ ,
    \new_[80133]_ , \new_[80136]_ , \new_[80139]_ , \new_[80140]_ ,
    \new_[80141]_ , \new_[80144]_ , \new_[80147]_ , \new_[80148]_ ,
    \new_[80151]_ , \new_[80154]_ , \new_[80155]_ , \new_[80156]_ ,
    \new_[80160]_ , \new_[80161]_ , \new_[80164]_ , \new_[80167]_ ,
    \new_[80168]_ , \new_[80169]_ , \new_[80172]_ , \new_[80175]_ ,
    \new_[80176]_ , \new_[80179]_ , \new_[80182]_ , \new_[80183]_ ,
    \new_[80184]_ , \new_[80188]_ , \new_[80189]_ , \new_[80192]_ ,
    \new_[80195]_ , \new_[80196]_ , \new_[80197]_ , \new_[80200]_ ,
    \new_[80203]_ , \new_[80204]_ , \new_[80207]_ , \new_[80210]_ ,
    \new_[80211]_ , \new_[80212]_ , \new_[80216]_ , \new_[80217]_ ,
    \new_[80220]_ , \new_[80223]_ , \new_[80224]_ , \new_[80225]_ ,
    \new_[80228]_ , \new_[80231]_ , \new_[80232]_ , \new_[80235]_ ,
    \new_[80238]_ , \new_[80239]_ , \new_[80240]_ , \new_[80244]_ ,
    \new_[80245]_ , \new_[80248]_ , \new_[80251]_ , \new_[80252]_ ,
    \new_[80253]_ , \new_[80256]_ , \new_[80259]_ , \new_[80260]_ ,
    \new_[80263]_ , \new_[80266]_ , \new_[80267]_ , \new_[80268]_ ,
    \new_[80272]_ , \new_[80273]_ , \new_[80276]_ , \new_[80279]_ ,
    \new_[80280]_ , \new_[80281]_ , \new_[80284]_ , \new_[80287]_ ,
    \new_[80288]_ , \new_[80291]_ , \new_[80294]_ , \new_[80295]_ ,
    \new_[80296]_ , \new_[80300]_ , \new_[80301]_ , \new_[80304]_ ,
    \new_[80307]_ , \new_[80308]_ , \new_[80309]_ , \new_[80312]_ ,
    \new_[80315]_ , \new_[80316]_ , \new_[80319]_ , \new_[80322]_ ,
    \new_[80323]_ , \new_[80324]_ , \new_[80328]_ , \new_[80329]_ ,
    \new_[80332]_ , \new_[80335]_ , \new_[80336]_ , \new_[80337]_ ,
    \new_[80340]_ , \new_[80343]_ , \new_[80344]_ , \new_[80347]_ ,
    \new_[80350]_ , \new_[80351]_ , \new_[80352]_ , \new_[80356]_ ,
    \new_[80357]_ , \new_[80360]_ , \new_[80363]_ , \new_[80364]_ ,
    \new_[80365]_ , \new_[80368]_ , \new_[80371]_ , \new_[80372]_ ,
    \new_[80375]_ , \new_[80378]_ , \new_[80379]_ , \new_[80380]_ ,
    \new_[80384]_ , \new_[80385]_ , \new_[80388]_ , \new_[80391]_ ,
    \new_[80392]_ , \new_[80393]_ , \new_[80396]_ , \new_[80399]_ ,
    \new_[80400]_ , \new_[80403]_ , \new_[80406]_ , \new_[80407]_ ,
    \new_[80408]_ , \new_[80412]_ , \new_[80413]_ , \new_[80416]_ ,
    \new_[80419]_ , \new_[80420]_ , \new_[80421]_ , \new_[80424]_ ,
    \new_[80427]_ , \new_[80428]_ , \new_[80431]_ , \new_[80434]_ ,
    \new_[80435]_ , \new_[80436]_ , \new_[80440]_ , \new_[80441]_ ,
    \new_[80444]_ , \new_[80447]_ , \new_[80448]_ , \new_[80449]_ ,
    \new_[80452]_ , \new_[80455]_ , \new_[80456]_ , \new_[80459]_ ,
    \new_[80462]_ , \new_[80463]_ , \new_[80464]_ , \new_[80468]_ ,
    \new_[80469]_ , \new_[80472]_ , \new_[80475]_ , \new_[80476]_ ,
    \new_[80477]_ , \new_[80480]_ , \new_[80483]_ , \new_[80484]_ ,
    \new_[80487]_ , \new_[80490]_ , \new_[80491]_ , \new_[80492]_ ,
    \new_[80496]_ , \new_[80497]_ , \new_[80500]_ , \new_[80503]_ ,
    \new_[80504]_ , \new_[80505]_ , \new_[80508]_ , \new_[80511]_ ,
    \new_[80512]_ , \new_[80515]_ , \new_[80518]_ , \new_[80519]_ ,
    \new_[80520]_ , \new_[80524]_ , \new_[80525]_ , \new_[80528]_ ,
    \new_[80531]_ , \new_[80532]_ , \new_[80533]_ , \new_[80536]_ ,
    \new_[80539]_ , \new_[80540]_ , \new_[80543]_ , \new_[80546]_ ,
    \new_[80547]_ , \new_[80548]_ , \new_[80552]_ , \new_[80553]_ ,
    \new_[80556]_ , \new_[80559]_ , \new_[80560]_ , \new_[80561]_ ,
    \new_[80564]_ , \new_[80567]_ , \new_[80568]_ , \new_[80571]_ ,
    \new_[80574]_ , \new_[80575]_ , \new_[80576]_ , \new_[80580]_ ,
    \new_[80581]_ , \new_[80584]_ , \new_[80587]_ , \new_[80588]_ ,
    \new_[80589]_ , \new_[80592]_ , \new_[80595]_ , \new_[80596]_ ,
    \new_[80599]_ , \new_[80602]_ , \new_[80603]_ , \new_[80604]_ ,
    \new_[80608]_ , \new_[80609]_ , \new_[80612]_ , \new_[80615]_ ,
    \new_[80616]_ , \new_[80617]_ , \new_[80620]_ , \new_[80623]_ ,
    \new_[80624]_ , \new_[80627]_ , \new_[80630]_ , \new_[80631]_ ,
    \new_[80632]_ , \new_[80636]_ , \new_[80637]_ , \new_[80640]_ ,
    \new_[80643]_ , \new_[80644]_ , \new_[80645]_ , \new_[80648]_ ,
    \new_[80651]_ , \new_[80652]_ , \new_[80655]_ , \new_[80658]_ ,
    \new_[80659]_ , \new_[80660]_ , \new_[80664]_ , \new_[80665]_ ,
    \new_[80668]_ , \new_[80671]_ , \new_[80672]_ , \new_[80673]_ ,
    \new_[80676]_ , \new_[80679]_ , \new_[80680]_ , \new_[80683]_ ,
    \new_[80686]_ , \new_[80687]_ , \new_[80688]_ , \new_[80692]_ ,
    \new_[80693]_ , \new_[80696]_ , \new_[80699]_ , \new_[80700]_ ,
    \new_[80701]_ , \new_[80704]_ , \new_[80707]_ , \new_[80708]_ ,
    \new_[80711]_ , \new_[80714]_ , \new_[80715]_ , \new_[80716]_ ,
    \new_[80720]_ , \new_[80721]_ , \new_[80724]_ , \new_[80727]_ ,
    \new_[80728]_ , \new_[80729]_ , \new_[80732]_ , \new_[80735]_ ,
    \new_[80736]_ , \new_[80739]_ , \new_[80742]_ , \new_[80743]_ ,
    \new_[80744]_ , \new_[80748]_ , \new_[80749]_ , \new_[80752]_ ,
    \new_[80755]_ , \new_[80756]_ , \new_[80757]_ , \new_[80760]_ ,
    \new_[80763]_ , \new_[80764]_ , \new_[80767]_ , \new_[80770]_ ,
    \new_[80771]_ , \new_[80772]_ , \new_[80776]_ , \new_[80777]_ ,
    \new_[80780]_ , \new_[80783]_ , \new_[80784]_ , \new_[80785]_ ,
    \new_[80788]_ , \new_[80791]_ , \new_[80792]_ , \new_[80795]_ ,
    \new_[80798]_ , \new_[80799]_ , \new_[80800]_ , \new_[80804]_ ,
    \new_[80805]_ , \new_[80808]_ , \new_[80811]_ , \new_[80812]_ ,
    \new_[80813]_ , \new_[80816]_ , \new_[80819]_ , \new_[80820]_ ,
    \new_[80823]_ , \new_[80826]_ , \new_[80827]_ , \new_[80828]_ ,
    \new_[80832]_ , \new_[80833]_ , \new_[80836]_ , \new_[80839]_ ,
    \new_[80840]_ , \new_[80841]_ , \new_[80844]_ , \new_[80847]_ ,
    \new_[80848]_ , \new_[80851]_ , \new_[80854]_ , \new_[80855]_ ,
    \new_[80856]_ , \new_[80860]_ , \new_[80861]_ , \new_[80864]_ ,
    \new_[80867]_ , \new_[80868]_ , \new_[80869]_ , \new_[80872]_ ,
    \new_[80875]_ , \new_[80876]_ , \new_[80879]_ , \new_[80882]_ ,
    \new_[80883]_ , \new_[80884]_ , \new_[80888]_ , \new_[80889]_ ,
    \new_[80892]_ , \new_[80895]_ , \new_[80896]_ , \new_[80897]_ ,
    \new_[80900]_ , \new_[80903]_ , \new_[80904]_ , \new_[80907]_ ,
    \new_[80910]_ , \new_[80911]_ , \new_[80912]_ , \new_[80916]_ ,
    \new_[80917]_ , \new_[80920]_ , \new_[80923]_ , \new_[80924]_ ,
    \new_[80925]_ , \new_[80928]_ , \new_[80931]_ , \new_[80932]_ ,
    \new_[80935]_ , \new_[80938]_ , \new_[80939]_ , \new_[80940]_ ,
    \new_[80944]_ , \new_[80945]_ , \new_[80948]_ , \new_[80951]_ ,
    \new_[80952]_ , \new_[80953]_ , \new_[80956]_ , \new_[80959]_ ,
    \new_[80960]_ , \new_[80963]_ , \new_[80966]_ , \new_[80967]_ ,
    \new_[80968]_ , \new_[80972]_ , \new_[80973]_ , \new_[80976]_ ,
    \new_[80979]_ , \new_[80980]_ , \new_[80981]_ , \new_[80984]_ ,
    \new_[80987]_ , \new_[80988]_ , \new_[80991]_ , \new_[80994]_ ,
    \new_[80995]_ , \new_[80996]_ , \new_[81000]_ , \new_[81001]_ ,
    \new_[81004]_ , \new_[81007]_ , \new_[81008]_ , \new_[81009]_ ,
    \new_[81012]_ , \new_[81015]_ , \new_[81016]_ , \new_[81019]_ ,
    \new_[81022]_ , \new_[81023]_ , \new_[81024]_ , \new_[81028]_ ,
    \new_[81029]_ , \new_[81032]_ , \new_[81035]_ , \new_[81036]_ ,
    \new_[81037]_ , \new_[81040]_ , \new_[81043]_ , \new_[81044]_ ,
    \new_[81047]_ , \new_[81050]_ , \new_[81051]_ , \new_[81052]_ ,
    \new_[81056]_ , \new_[81057]_ , \new_[81060]_ , \new_[81063]_ ,
    \new_[81064]_ , \new_[81065]_ , \new_[81068]_ , \new_[81071]_ ,
    \new_[81072]_ , \new_[81075]_ , \new_[81078]_ , \new_[81079]_ ,
    \new_[81080]_ , \new_[81084]_ , \new_[81085]_ , \new_[81088]_ ,
    \new_[81091]_ , \new_[81092]_ , \new_[81093]_ , \new_[81096]_ ,
    \new_[81099]_ , \new_[81100]_ , \new_[81103]_ , \new_[81106]_ ,
    \new_[81107]_ , \new_[81108]_ , \new_[81112]_ , \new_[81113]_ ,
    \new_[81116]_ , \new_[81119]_ , \new_[81120]_ , \new_[81121]_ ,
    \new_[81124]_ , \new_[81127]_ , \new_[81128]_ , \new_[81131]_ ,
    \new_[81134]_ , \new_[81135]_ , \new_[81136]_ , \new_[81140]_ ,
    \new_[81141]_ , \new_[81144]_ , \new_[81147]_ , \new_[81148]_ ,
    \new_[81149]_ , \new_[81152]_ , \new_[81155]_ , \new_[81156]_ ,
    \new_[81159]_ , \new_[81162]_ , \new_[81163]_ , \new_[81164]_ ,
    \new_[81168]_ , \new_[81169]_ , \new_[81172]_ , \new_[81175]_ ,
    \new_[81176]_ , \new_[81177]_ , \new_[81180]_ , \new_[81183]_ ,
    \new_[81184]_ , \new_[81187]_ , \new_[81190]_ , \new_[81191]_ ,
    \new_[81192]_ , \new_[81196]_ , \new_[81197]_ , \new_[81200]_ ,
    \new_[81203]_ , \new_[81204]_ , \new_[81205]_ , \new_[81208]_ ,
    \new_[81211]_ , \new_[81212]_ , \new_[81215]_ , \new_[81218]_ ,
    \new_[81219]_ , \new_[81220]_ , \new_[81224]_ , \new_[81225]_ ,
    \new_[81228]_ , \new_[81231]_ , \new_[81232]_ , \new_[81233]_ ,
    \new_[81236]_ , \new_[81239]_ , \new_[81240]_ , \new_[81243]_ ,
    \new_[81246]_ , \new_[81247]_ , \new_[81248]_ , \new_[81252]_ ,
    \new_[81253]_ , \new_[81256]_ , \new_[81259]_ , \new_[81260]_ ,
    \new_[81261]_ , \new_[81264]_ , \new_[81267]_ , \new_[81268]_ ,
    \new_[81271]_ , \new_[81274]_ , \new_[81275]_ , \new_[81276]_ ,
    \new_[81280]_ , \new_[81281]_ , \new_[81284]_ , \new_[81287]_ ,
    \new_[81288]_ , \new_[81289]_ , \new_[81292]_ , \new_[81295]_ ,
    \new_[81296]_ , \new_[81299]_ , \new_[81302]_ , \new_[81303]_ ,
    \new_[81304]_ , \new_[81308]_ , \new_[81309]_ , \new_[81312]_ ,
    \new_[81315]_ , \new_[81316]_ , \new_[81317]_ , \new_[81320]_ ,
    \new_[81323]_ , \new_[81324]_ , \new_[81327]_ , \new_[81330]_ ,
    \new_[81331]_ , \new_[81332]_ , \new_[81336]_ , \new_[81337]_ ,
    \new_[81340]_ , \new_[81343]_ , \new_[81344]_ , \new_[81345]_ ,
    \new_[81348]_ , \new_[81351]_ , \new_[81352]_ , \new_[81355]_ ,
    \new_[81358]_ , \new_[81359]_ , \new_[81360]_ , \new_[81364]_ ,
    \new_[81365]_ , \new_[81368]_ , \new_[81371]_ , \new_[81372]_ ,
    \new_[81373]_ , \new_[81376]_ , \new_[81379]_ , \new_[81380]_ ,
    \new_[81383]_ , \new_[81386]_ , \new_[81387]_ , \new_[81388]_ ,
    \new_[81392]_ , \new_[81393]_ , \new_[81396]_ , \new_[81399]_ ,
    \new_[81400]_ , \new_[81401]_ , \new_[81404]_ , \new_[81407]_ ,
    \new_[81408]_ , \new_[81411]_ , \new_[81414]_ , \new_[81415]_ ,
    \new_[81416]_ , \new_[81420]_ , \new_[81421]_ , \new_[81424]_ ,
    \new_[81427]_ , \new_[81428]_ , \new_[81429]_ , \new_[81432]_ ,
    \new_[81435]_ , \new_[81436]_ , \new_[81439]_ , \new_[81442]_ ,
    \new_[81443]_ , \new_[81444]_ , \new_[81448]_ , \new_[81449]_ ,
    \new_[81452]_ , \new_[81455]_ , \new_[81456]_ , \new_[81457]_ ,
    \new_[81460]_ , \new_[81463]_ , \new_[81464]_ , \new_[81467]_ ,
    \new_[81470]_ , \new_[81471]_ , \new_[81472]_ , \new_[81476]_ ,
    \new_[81477]_ , \new_[81480]_ , \new_[81483]_ , \new_[81484]_ ,
    \new_[81485]_ , \new_[81488]_ , \new_[81491]_ , \new_[81492]_ ,
    \new_[81495]_ , \new_[81498]_ , \new_[81499]_ , \new_[81500]_ ,
    \new_[81504]_ , \new_[81505]_ , \new_[81508]_ , \new_[81511]_ ,
    \new_[81512]_ , \new_[81513]_ , \new_[81516]_ , \new_[81519]_ ,
    \new_[81520]_ , \new_[81523]_ , \new_[81526]_ , \new_[81527]_ ,
    \new_[81528]_ , \new_[81532]_ , \new_[81533]_ , \new_[81536]_ ,
    \new_[81539]_ , \new_[81540]_ , \new_[81541]_ , \new_[81544]_ ,
    \new_[81547]_ , \new_[81548]_ , \new_[81551]_ , \new_[81554]_ ,
    \new_[81555]_ , \new_[81556]_ , \new_[81560]_ , \new_[81561]_ ,
    \new_[81564]_ , \new_[81567]_ , \new_[81568]_ , \new_[81569]_ ,
    \new_[81572]_ , \new_[81575]_ , \new_[81576]_ , \new_[81579]_ ,
    \new_[81582]_ , \new_[81583]_ , \new_[81584]_ , \new_[81588]_ ,
    \new_[81589]_ , \new_[81592]_ , \new_[81595]_ , \new_[81596]_ ,
    \new_[81597]_ , \new_[81600]_ , \new_[81603]_ , \new_[81604]_ ,
    \new_[81607]_ , \new_[81610]_ , \new_[81611]_ , \new_[81612]_ ,
    \new_[81616]_ , \new_[81617]_ , \new_[81620]_ , \new_[81623]_ ,
    \new_[81624]_ , \new_[81625]_ , \new_[81628]_ , \new_[81631]_ ,
    \new_[81632]_ , \new_[81635]_ , \new_[81638]_ , \new_[81639]_ ,
    \new_[81640]_ , \new_[81644]_ , \new_[81645]_ , \new_[81648]_ ,
    \new_[81651]_ , \new_[81652]_ , \new_[81653]_ , \new_[81656]_ ,
    \new_[81659]_ , \new_[81660]_ , \new_[81663]_ , \new_[81666]_ ,
    \new_[81667]_ , \new_[81668]_ , \new_[81672]_ , \new_[81673]_ ,
    \new_[81676]_ , \new_[81679]_ , \new_[81680]_ , \new_[81681]_ ,
    \new_[81684]_ , \new_[81687]_ , \new_[81688]_ , \new_[81691]_ ,
    \new_[81694]_ , \new_[81695]_ , \new_[81696]_ , \new_[81700]_ ,
    \new_[81701]_ , \new_[81704]_ , \new_[81707]_ , \new_[81708]_ ,
    \new_[81709]_ , \new_[81712]_ , \new_[81715]_ , \new_[81716]_ ,
    \new_[81719]_ , \new_[81722]_ , \new_[81723]_ , \new_[81724]_ ,
    \new_[81728]_ , \new_[81729]_ , \new_[81732]_ , \new_[81735]_ ,
    \new_[81736]_ , \new_[81737]_ , \new_[81740]_ , \new_[81743]_ ,
    \new_[81744]_ , \new_[81747]_ , \new_[81750]_ , \new_[81751]_ ,
    \new_[81752]_ , \new_[81756]_ , \new_[81757]_ , \new_[81760]_ ,
    \new_[81763]_ , \new_[81764]_ , \new_[81765]_ , \new_[81768]_ ,
    \new_[81771]_ , \new_[81772]_ , \new_[81775]_ , \new_[81778]_ ,
    \new_[81779]_ , \new_[81780]_ , \new_[81784]_ , \new_[81785]_ ,
    \new_[81788]_ , \new_[81791]_ , \new_[81792]_ , \new_[81793]_ ,
    \new_[81796]_ , \new_[81799]_ , \new_[81800]_ , \new_[81803]_ ,
    \new_[81806]_ , \new_[81807]_ , \new_[81808]_ , \new_[81812]_ ,
    \new_[81813]_ , \new_[81816]_ , \new_[81819]_ , \new_[81820]_ ,
    \new_[81821]_ , \new_[81824]_ , \new_[81827]_ , \new_[81828]_ ,
    \new_[81831]_ , \new_[81834]_ , \new_[81835]_ , \new_[81836]_ ,
    \new_[81840]_ , \new_[81841]_ , \new_[81844]_ , \new_[81847]_ ,
    \new_[81848]_ , \new_[81849]_ , \new_[81852]_ , \new_[81855]_ ,
    \new_[81856]_ , \new_[81859]_ , \new_[81862]_ , \new_[81863]_ ,
    \new_[81864]_ , \new_[81868]_ , \new_[81869]_ , \new_[81872]_ ,
    \new_[81875]_ , \new_[81876]_ , \new_[81877]_ , \new_[81880]_ ,
    \new_[81883]_ , \new_[81884]_ , \new_[81887]_ , \new_[81890]_ ,
    \new_[81891]_ , \new_[81892]_ , \new_[81896]_ , \new_[81897]_ ,
    \new_[81900]_ , \new_[81903]_ , \new_[81904]_ , \new_[81905]_ ,
    \new_[81908]_ , \new_[81911]_ , \new_[81912]_ , \new_[81915]_ ,
    \new_[81918]_ , \new_[81919]_ , \new_[81920]_ , \new_[81924]_ ,
    \new_[81925]_ , \new_[81928]_ , \new_[81931]_ , \new_[81932]_ ,
    \new_[81933]_ , \new_[81936]_ , \new_[81939]_ , \new_[81940]_ ,
    \new_[81943]_ , \new_[81946]_ , \new_[81947]_ , \new_[81948]_ ,
    \new_[81952]_ , \new_[81953]_ , \new_[81956]_ , \new_[81959]_ ,
    \new_[81960]_ , \new_[81961]_ , \new_[81964]_ , \new_[81967]_ ,
    \new_[81968]_ , \new_[81971]_ , \new_[81974]_ , \new_[81975]_ ,
    \new_[81976]_ , \new_[81980]_ , \new_[81981]_ , \new_[81984]_ ,
    \new_[81987]_ , \new_[81988]_ , \new_[81989]_ , \new_[81992]_ ,
    \new_[81995]_ , \new_[81996]_ , \new_[81999]_ , \new_[82002]_ ,
    \new_[82003]_ , \new_[82004]_ , \new_[82008]_ , \new_[82009]_ ,
    \new_[82012]_ , \new_[82015]_ , \new_[82016]_ , \new_[82017]_ ,
    \new_[82020]_ , \new_[82023]_ , \new_[82024]_ , \new_[82027]_ ,
    \new_[82030]_ , \new_[82031]_ , \new_[82032]_ , \new_[82036]_ ,
    \new_[82037]_ , \new_[82040]_ , \new_[82043]_ , \new_[82044]_ ,
    \new_[82045]_ , \new_[82048]_ , \new_[82051]_ , \new_[82052]_ ,
    \new_[82055]_ , \new_[82058]_ , \new_[82059]_ , \new_[82060]_ ,
    \new_[82064]_ , \new_[82065]_ , \new_[82068]_ , \new_[82071]_ ,
    \new_[82072]_ , \new_[82073]_ , \new_[82076]_ , \new_[82079]_ ,
    \new_[82080]_ , \new_[82083]_ , \new_[82086]_ , \new_[82087]_ ,
    \new_[82088]_ , \new_[82092]_ , \new_[82093]_ , \new_[82096]_ ,
    \new_[82099]_ , \new_[82100]_ , \new_[82101]_ , \new_[82104]_ ,
    \new_[82107]_ , \new_[82108]_ , \new_[82111]_ , \new_[82114]_ ,
    \new_[82115]_ , \new_[82116]_ , \new_[82120]_ , \new_[82121]_ ,
    \new_[82124]_ , \new_[82127]_ , \new_[82128]_ , \new_[82129]_ ,
    \new_[82132]_ , \new_[82135]_ , \new_[82136]_ , \new_[82139]_ ,
    \new_[82142]_ , \new_[82143]_ , \new_[82144]_ , \new_[82148]_ ,
    \new_[82149]_ , \new_[82152]_ , \new_[82155]_ , \new_[82156]_ ,
    \new_[82157]_ , \new_[82160]_ , \new_[82163]_ , \new_[82164]_ ,
    \new_[82167]_ , \new_[82170]_ , \new_[82171]_ , \new_[82172]_ ,
    \new_[82176]_ , \new_[82177]_ , \new_[82180]_ , \new_[82183]_ ,
    \new_[82184]_ , \new_[82185]_ , \new_[82188]_ , \new_[82191]_ ,
    \new_[82192]_ , \new_[82195]_ , \new_[82198]_ , \new_[82199]_ ,
    \new_[82200]_ , \new_[82204]_ , \new_[82205]_ , \new_[82208]_ ,
    \new_[82211]_ , \new_[82212]_ , \new_[82213]_ , \new_[82216]_ ,
    \new_[82219]_ , \new_[82220]_ , \new_[82223]_ , \new_[82226]_ ,
    \new_[82227]_ , \new_[82228]_ , \new_[82232]_ , \new_[82233]_ ,
    \new_[82236]_ , \new_[82239]_ , \new_[82240]_ , \new_[82241]_ ,
    \new_[82244]_ , \new_[82247]_ , \new_[82248]_ , \new_[82251]_ ,
    \new_[82254]_ , \new_[82255]_ , \new_[82256]_ , \new_[82260]_ ,
    \new_[82261]_ , \new_[82264]_ , \new_[82267]_ , \new_[82268]_ ,
    \new_[82269]_ , \new_[82272]_ , \new_[82275]_ , \new_[82276]_ ,
    \new_[82279]_ , \new_[82282]_ , \new_[82283]_ , \new_[82284]_ ,
    \new_[82288]_ , \new_[82289]_ , \new_[82292]_ , \new_[82295]_ ,
    \new_[82296]_ , \new_[82297]_ , \new_[82300]_ , \new_[82303]_ ,
    \new_[82304]_ , \new_[82307]_ , \new_[82310]_ , \new_[82311]_ ,
    \new_[82312]_ , \new_[82316]_ , \new_[82317]_ , \new_[82320]_ ,
    \new_[82323]_ , \new_[82324]_ , \new_[82325]_ , \new_[82328]_ ,
    \new_[82331]_ , \new_[82332]_ , \new_[82335]_ , \new_[82338]_ ,
    \new_[82339]_ , \new_[82340]_ , \new_[82344]_ , \new_[82345]_ ,
    \new_[82348]_ , \new_[82351]_ , \new_[82352]_ , \new_[82353]_ ,
    \new_[82356]_ , \new_[82359]_ , \new_[82360]_ , \new_[82363]_ ,
    \new_[82366]_ , \new_[82367]_ , \new_[82368]_ , \new_[82372]_ ,
    \new_[82373]_ , \new_[82376]_ , \new_[82379]_ , \new_[82380]_ ,
    \new_[82381]_ , \new_[82384]_ , \new_[82387]_ , \new_[82388]_ ,
    \new_[82391]_ , \new_[82394]_ , \new_[82395]_ , \new_[82396]_ ,
    \new_[82400]_ , \new_[82401]_ , \new_[82404]_ , \new_[82407]_ ,
    \new_[82408]_ , \new_[82409]_ , \new_[82412]_ , \new_[82415]_ ,
    \new_[82416]_ , \new_[82419]_ , \new_[82422]_ , \new_[82423]_ ,
    \new_[82424]_ , \new_[82428]_ , \new_[82429]_ , \new_[82432]_ ,
    \new_[82435]_ , \new_[82436]_ , \new_[82437]_ , \new_[82440]_ ,
    \new_[82443]_ , \new_[82444]_ , \new_[82447]_ , \new_[82450]_ ,
    \new_[82451]_ , \new_[82452]_ , \new_[82456]_ , \new_[82457]_ ,
    \new_[82460]_ , \new_[82463]_ , \new_[82464]_ , \new_[82465]_ ,
    \new_[82468]_ , \new_[82471]_ , \new_[82472]_ , \new_[82475]_ ,
    \new_[82478]_ , \new_[82479]_ , \new_[82480]_ , \new_[82484]_ ,
    \new_[82485]_ , \new_[82488]_ , \new_[82491]_ , \new_[82492]_ ,
    \new_[82493]_ , \new_[82496]_ , \new_[82499]_ , \new_[82500]_ ,
    \new_[82503]_ , \new_[82506]_ , \new_[82507]_ , \new_[82508]_ ,
    \new_[82512]_ , \new_[82513]_ , \new_[82516]_ , \new_[82519]_ ,
    \new_[82520]_ , \new_[82521]_ , \new_[82524]_ , \new_[82527]_ ,
    \new_[82528]_ , \new_[82531]_ , \new_[82534]_ , \new_[82535]_ ,
    \new_[82536]_ , \new_[82540]_ , \new_[82541]_ , \new_[82544]_ ,
    \new_[82547]_ , \new_[82548]_ , \new_[82549]_ , \new_[82552]_ ,
    \new_[82555]_ , \new_[82556]_ , \new_[82559]_ , \new_[82562]_ ,
    \new_[82563]_ , \new_[82564]_ , \new_[82568]_ , \new_[82569]_ ,
    \new_[82572]_ , \new_[82575]_ , \new_[82576]_ , \new_[82577]_ ,
    \new_[82580]_ , \new_[82583]_ , \new_[82584]_ , \new_[82587]_ ,
    \new_[82590]_ , \new_[82591]_ , \new_[82592]_ , \new_[82596]_ ,
    \new_[82597]_ , \new_[82600]_ , \new_[82603]_ , \new_[82604]_ ,
    \new_[82605]_ , \new_[82608]_ , \new_[82611]_ , \new_[82612]_ ,
    \new_[82615]_ , \new_[82618]_ , \new_[82619]_ , \new_[82620]_ ,
    \new_[82624]_ , \new_[82625]_ , \new_[82628]_ , \new_[82631]_ ,
    \new_[82632]_ , \new_[82633]_ , \new_[82636]_ , \new_[82639]_ ,
    \new_[82640]_ , \new_[82643]_ , \new_[82646]_ , \new_[82647]_ ,
    \new_[82648]_ , \new_[82652]_ , \new_[82653]_ , \new_[82656]_ ,
    \new_[82659]_ , \new_[82660]_ , \new_[82661]_ , \new_[82664]_ ,
    \new_[82667]_ , \new_[82668]_ , \new_[82671]_ , \new_[82674]_ ,
    \new_[82675]_ , \new_[82676]_ , \new_[82680]_ , \new_[82681]_ ,
    \new_[82684]_ , \new_[82687]_ , \new_[82688]_ , \new_[82689]_ ,
    \new_[82692]_ , \new_[82695]_ , \new_[82696]_ , \new_[82699]_ ,
    \new_[82702]_ , \new_[82703]_ , \new_[82704]_ , \new_[82708]_ ,
    \new_[82709]_ , \new_[82712]_ , \new_[82715]_ , \new_[82716]_ ,
    \new_[82717]_ , \new_[82720]_ , \new_[82723]_ , \new_[82724]_ ,
    \new_[82727]_ , \new_[82730]_ , \new_[82731]_ , \new_[82732]_ ,
    \new_[82736]_ , \new_[82737]_ , \new_[82740]_ , \new_[82743]_ ,
    \new_[82744]_ , \new_[82745]_ , \new_[82748]_ , \new_[82751]_ ,
    \new_[82752]_ , \new_[82755]_ , \new_[82758]_ , \new_[82759]_ ,
    \new_[82760]_ , \new_[82764]_ , \new_[82765]_ , \new_[82768]_ ,
    \new_[82771]_ , \new_[82772]_ , \new_[82773]_ , \new_[82776]_ ,
    \new_[82779]_ , \new_[82780]_ , \new_[82783]_ , \new_[82786]_ ,
    \new_[82787]_ , \new_[82788]_ , \new_[82792]_ , \new_[82793]_ ,
    \new_[82796]_ , \new_[82799]_ , \new_[82800]_ , \new_[82801]_ ,
    \new_[82804]_ , \new_[82807]_ , \new_[82808]_ , \new_[82811]_ ,
    \new_[82814]_ , \new_[82815]_ , \new_[82816]_ , \new_[82820]_ ,
    \new_[82821]_ , \new_[82824]_ , \new_[82827]_ , \new_[82828]_ ,
    \new_[82829]_ , \new_[82832]_ , \new_[82835]_ , \new_[82836]_ ,
    \new_[82839]_ , \new_[82842]_ , \new_[82843]_ , \new_[82844]_ ,
    \new_[82848]_ , \new_[82849]_ , \new_[82852]_ , \new_[82855]_ ,
    \new_[82856]_ , \new_[82857]_ , \new_[82860]_ , \new_[82863]_ ,
    \new_[82864]_ , \new_[82867]_ , \new_[82870]_ , \new_[82871]_ ,
    \new_[82872]_ , \new_[82876]_ , \new_[82877]_ , \new_[82880]_ ,
    \new_[82883]_ , \new_[82884]_ , \new_[82885]_ , \new_[82888]_ ,
    \new_[82891]_ , \new_[82892]_ , \new_[82895]_ , \new_[82898]_ ,
    \new_[82899]_ , \new_[82900]_ , \new_[82904]_ , \new_[82905]_ ,
    \new_[82908]_ , \new_[82911]_ , \new_[82912]_ , \new_[82913]_ ,
    \new_[82916]_ , \new_[82919]_ , \new_[82920]_ , \new_[82923]_ ,
    \new_[82926]_ , \new_[82927]_ , \new_[82928]_ , \new_[82932]_ ,
    \new_[82933]_ , \new_[82936]_ , \new_[82939]_ , \new_[82940]_ ,
    \new_[82941]_ , \new_[82944]_ , \new_[82947]_ , \new_[82948]_ ,
    \new_[82951]_ , \new_[82954]_ , \new_[82955]_ , \new_[82956]_ ,
    \new_[82960]_ , \new_[82961]_ , \new_[82964]_ , \new_[82967]_ ,
    \new_[82968]_ , \new_[82969]_ , \new_[82972]_ , \new_[82975]_ ,
    \new_[82976]_ , \new_[82979]_ , \new_[82982]_ , \new_[82983]_ ,
    \new_[82984]_ , \new_[82988]_ , \new_[82989]_ , \new_[82992]_ ,
    \new_[82995]_ , \new_[82996]_ , \new_[82997]_ , \new_[83000]_ ,
    \new_[83003]_ , \new_[83004]_ , \new_[83007]_ , \new_[83010]_ ,
    \new_[83011]_ , \new_[83012]_ , \new_[83016]_ , \new_[83017]_ ,
    \new_[83020]_ , \new_[83023]_ , \new_[83024]_ , \new_[83025]_ ,
    \new_[83028]_ , \new_[83031]_ , \new_[83032]_ , \new_[83035]_ ,
    \new_[83038]_ , \new_[83039]_ , \new_[83040]_ , \new_[83044]_ ,
    \new_[83045]_ , \new_[83048]_ , \new_[83051]_ , \new_[83052]_ ,
    \new_[83053]_ , \new_[83056]_ , \new_[83059]_ , \new_[83060]_ ,
    \new_[83063]_ , \new_[83066]_ , \new_[83067]_ , \new_[83068]_ ,
    \new_[83072]_ , \new_[83073]_ , \new_[83076]_ , \new_[83079]_ ,
    \new_[83080]_ , \new_[83081]_ , \new_[83084]_ , \new_[83087]_ ,
    \new_[83088]_ , \new_[83091]_ , \new_[83094]_ , \new_[83095]_ ,
    \new_[83096]_ , \new_[83100]_ , \new_[83101]_ , \new_[83104]_ ,
    \new_[83107]_ , \new_[83108]_ , \new_[83109]_ , \new_[83112]_ ,
    \new_[83115]_ , \new_[83116]_ , \new_[83119]_ , \new_[83122]_ ,
    \new_[83123]_ , \new_[83124]_ , \new_[83128]_ , \new_[83129]_ ,
    \new_[83132]_ , \new_[83135]_ , \new_[83136]_ , \new_[83137]_ ,
    \new_[83140]_ , \new_[83143]_ , \new_[83144]_ , \new_[83147]_ ,
    \new_[83150]_ , \new_[83151]_ , \new_[83152]_ , \new_[83156]_ ,
    \new_[83157]_ , \new_[83160]_ , \new_[83163]_ , \new_[83164]_ ,
    \new_[83165]_ , \new_[83168]_ , \new_[83171]_ , \new_[83172]_ ,
    \new_[83175]_ , \new_[83178]_ , \new_[83179]_ , \new_[83180]_ ,
    \new_[83184]_ , \new_[83185]_ , \new_[83188]_ , \new_[83191]_ ,
    \new_[83192]_ , \new_[83193]_ , \new_[83196]_ , \new_[83199]_ ,
    \new_[83200]_ , \new_[83203]_ , \new_[83206]_ , \new_[83207]_ ,
    \new_[83208]_ , \new_[83212]_ , \new_[83213]_ , \new_[83216]_ ,
    \new_[83219]_ , \new_[83220]_ , \new_[83221]_ , \new_[83224]_ ,
    \new_[83227]_ , \new_[83228]_ , \new_[83231]_ , \new_[83234]_ ,
    \new_[83235]_ , \new_[83236]_ , \new_[83240]_ , \new_[83241]_ ,
    \new_[83244]_ , \new_[83247]_ , \new_[83248]_ , \new_[83249]_ ,
    \new_[83252]_ , \new_[83255]_ , \new_[83256]_ , \new_[83259]_ ,
    \new_[83262]_ , \new_[83263]_ , \new_[83264]_ , \new_[83268]_ ,
    \new_[83269]_ , \new_[83272]_ , \new_[83275]_ , \new_[83276]_ ,
    \new_[83277]_ , \new_[83280]_ , \new_[83283]_ , \new_[83284]_ ,
    \new_[83287]_ , \new_[83290]_ , \new_[83291]_ , \new_[83292]_ ,
    \new_[83296]_ , \new_[83297]_ , \new_[83300]_ , \new_[83303]_ ,
    \new_[83304]_ , \new_[83305]_ , \new_[83308]_ , \new_[83311]_ ,
    \new_[83312]_ , \new_[83315]_ , \new_[83318]_ , \new_[83319]_ ,
    \new_[83320]_ , \new_[83324]_ , \new_[83325]_ , \new_[83328]_ ,
    \new_[83331]_ , \new_[83332]_ , \new_[83333]_ , \new_[83336]_ ,
    \new_[83339]_ , \new_[83340]_ , \new_[83343]_ , \new_[83346]_ ,
    \new_[83347]_ , \new_[83348]_ , \new_[83352]_ , \new_[83353]_ ,
    \new_[83356]_ , \new_[83359]_ , \new_[83360]_ , \new_[83361]_ ,
    \new_[83364]_ , \new_[83367]_ , \new_[83368]_ , \new_[83371]_ ,
    \new_[83374]_ , \new_[83375]_ , \new_[83376]_ , \new_[83380]_ ,
    \new_[83381]_ , \new_[83384]_ , \new_[83387]_ , \new_[83388]_ ,
    \new_[83389]_ , \new_[83392]_ , \new_[83395]_ , \new_[83396]_ ,
    \new_[83399]_ , \new_[83402]_ , \new_[83403]_ , \new_[83404]_ ,
    \new_[83408]_ , \new_[83409]_ , \new_[83412]_ , \new_[83415]_ ,
    \new_[83416]_ , \new_[83417]_ , \new_[83420]_ , \new_[83423]_ ,
    \new_[83424]_ , \new_[83427]_ , \new_[83430]_ , \new_[83431]_ ,
    \new_[83432]_ , \new_[83436]_ , \new_[83437]_ , \new_[83440]_ ,
    \new_[83443]_ , \new_[83444]_ , \new_[83445]_ , \new_[83448]_ ,
    \new_[83451]_ , \new_[83452]_ , \new_[83455]_ , \new_[83458]_ ,
    \new_[83459]_ , \new_[83460]_ , \new_[83464]_ , \new_[83465]_ ,
    \new_[83468]_ , \new_[83471]_ , \new_[83472]_ , \new_[83473]_ ,
    \new_[83476]_ , \new_[83479]_ , \new_[83480]_ , \new_[83483]_ ,
    \new_[83486]_ , \new_[83487]_ , \new_[83488]_ , \new_[83492]_ ,
    \new_[83493]_ , \new_[83496]_ , \new_[83499]_ , \new_[83500]_ ,
    \new_[83501]_ , \new_[83504]_ , \new_[83507]_ , \new_[83508]_ ,
    \new_[83511]_ , \new_[83514]_ , \new_[83515]_ , \new_[83516]_ ,
    \new_[83520]_ , \new_[83521]_ , \new_[83524]_ , \new_[83527]_ ,
    \new_[83528]_ , \new_[83529]_ , \new_[83532]_ , \new_[83535]_ ,
    \new_[83536]_ , \new_[83539]_ , \new_[83542]_ , \new_[83543]_ ,
    \new_[83544]_ , \new_[83548]_ , \new_[83549]_ , \new_[83552]_ ,
    \new_[83555]_ , \new_[83556]_ , \new_[83557]_ , \new_[83560]_ ,
    \new_[83563]_ , \new_[83564]_ , \new_[83567]_ , \new_[83570]_ ,
    \new_[83571]_ , \new_[83572]_ , \new_[83576]_ , \new_[83577]_ ,
    \new_[83580]_ , \new_[83583]_ , \new_[83584]_ , \new_[83585]_ ,
    \new_[83588]_ , \new_[83591]_ , \new_[83592]_ , \new_[83595]_ ,
    \new_[83598]_ , \new_[83599]_ , \new_[83600]_ , \new_[83604]_ ,
    \new_[83605]_ , \new_[83608]_ , \new_[83611]_ , \new_[83612]_ ,
    \new_[83613]_ , \new_[83616]_ , \new_[83619]_ , \new_[83620]_ ,
    \new_[83623]_ , \new_[83626]_ , \new_[83627]_ , \new_[83628]_ ,
    \new_[83632]_ , \new_[83633]_ , \new_[83636]_ , \new_[83639]_ ,
    \new_[83640]_ , \new_[83641]_ , \new_[83644]_ , \new_[83647]_ ,
    \new_[83648]_ , \new_[83651]_ , \new_[83654]_ , \new_[83655]_ ,
    \new_[83656]_ , \new_[83660]_ , \new_[83661]_ , \new_[83664]_ ,
    \new_[83667]_ , \new_[83668]_ , \new_[83669]_ , \new_[83672]_ ,
    \new_[83675]_ , \new_[83676]_ , \new_[83679]_ , \new_[83682]_ ,
    \new_[83683]_ , \new_[83684]_ , \new_[83688]_ , \new_[83689]_ ,
    \new_[83692]_ , \new_[83695]_ , \new_[83696]_ , \new_[83697]_ ,
    \new_[83700]_ , \new_[83703]_ , \new_[83704]_ , \new_[83707]_ ,
    \new_[83710]_ , \new_[83711]_ , \new_[83712]_ , \new_[83716]_ ,
    \new_[83717]_ , \new_[83720]_ , \new_[83723]_ , \new_[83724]_ ,
    \new_[83725]_ , \new_[83728]_ , \new_[83731]_ , \new_[83732]_ ,
    \new_[83735]_ , \new_[83738]_ , \new_[83739]_ , \new_[83740]_ ,
    \new_[83744]_ , \new_[83745]_ , \new_[83748]_ , \new_[83751]_ ,
    \new_[83752]_ , \new_[83753]_ , \new_[83756]_ , \new_[83759]_ ,
    \new_[83760]_ , \new_[83763]_ , \new_[83766]_ , \new_[83767]_ ,
    \new_[83768]_ , \new_[83772]_ , \new_[83773]_ , \new_[83776]_ ,
    \new_[83779]_ , \new_[83780]_ , \new_[83781]_ , \new_[83784]_ ,
    \new_[83787]_ , \new_[83788]_ , \new_[83791]_ , \new_[83794]_ ,
    \new_[83795]_ , \new_[83796]_ , \new_[83800]_ , \new_[83801]_ ,
    \new_[83804]_ , \new_[83807]_ , \new_[83808]_ , \new_[83809]_ ,
    \new_[83812]_ , \new_[83815]_ , \new_[83816]_ , \new_[83819]_ ,
    \new_[83822]_ , \new_[83823]_ , \new_[83824]_ , \new_[83828]_ ,
    \new_[83829]_ , \new_[83832]_ , \new_[83835]_ , \new_[83836]_ ,
    \new_[83837]_ , \new_[83840]_ , \new_[83843]_ , \new_[83844]_ ,
    \new_[83847]_ , \new_[83850]_ , \new_[83851]_ , \new_[83852]_ ,
    \new_[83856]_ , \new_[83857]_ , \new_[83860]_ , \new_[83863]_ ,
    \new_[83864]_ , \new_[83865]_ , \new_[83868]_ , \new_[83871]_ ,
    \new_[83872]_ , \new_[83875]_ , \new_[83878]_ , \new_[83879]_ ,
    \new_[83880]_ , \new_[83884]_ , \new_[83885]_ , \new_[83888]_ ,
    \new_[83891]_ , \new_[83892]_ , \new_[83893]_ , \new_[83896]_ ,
    \new_[83899]_ , \new_[83900]_ , \new_[83903]_ , \new_[83906]_ ,
    \new_[83907]_ , \new_[83908]_ , \new_[83912]_ , \new_[83913]_ ,
    \new_[83916]_ , \new_[83919]_ , \new_[83920]_ , \new_[83921]_ ,
    \new_[83924]_ , \new_[83927]_ , \new_[83928]_ , \new_[83931]_ ,
    \new_[83934]_ , \new_[83935]_ , \new_[83936]_ , \new_[83940]_ ,
    \new_[83941]_ , \new_[83944]_ , \new_[83947]_ , \new_[83948]_ ,
    \new_[83949]_ , \new_[83952]_ , \new_[83955]_ , \new_[83956]_ ,
    \new_[83959]_ , \new_[83962]_ , \new_[83963]_ , \new_[83964]_ ,
    \new_[83968]_ , \new_[83969]_ , \new_[83972]_ , \new_[83975]_ ,
    \new_[83976]_ , \new_[83977]_ , \new_[83980]_ , \new_[83983]_ ,
    \new_[83984]_ , \new_[83987]_ , \new_[83990]_ , \new_[83991]_ ,
    \new_[83992]_ , \new_[83996]_ , \new_[83997]_ , \new_[84000]_ ,
    \new_[84003]_ , \new_[84004]_ , \new_[84005]_ , \new_[84008]_ ,
    \new_[84011]_ , \new_[84012]_ , \new_[84015]_ , \new_[84018]_ ,
    \new_[84019]_ , \new_[84020]_ , \new_[84024]_ , \new_[84025]_ ,
    \new_[84028]_ , \new_[84031]_ , \new_[84032]_ , \new_[84033]_ ,
    \new_[84036]_ , \new_[84039]_ , \new_[84040]_ , \new_[84043]_ ,
    \new_[84046]_ , \new_[84047]_ , \new_[84048]_ , \new_[84052]_ ,
    \new_[84053]_ , \new_[84056]_ , \new_[84059]_ , \new_[84060]_ ,
    \new_[84061]_ , \new_[84064]_ , \new_[84067]_ , \new_[84068]_ ,
    \new_[84071]_ , \new_[84074]_ , \new_[84075]_ , \new_[84076]_ ,
    \new_[84080]_ , \new_[84081]_ , \new_[84084]_ , \new_[84087]_ ,
    \new_[84088]_ , \new_[84089]_ , \new_[84092]_ , \new_[84095]_ ,
    \new_[84096]_ , \new_[84099]_ , \new_[84102]_ , \new_[84103]_ ,
    \new_[84104]_ , \new_[84108]_ , \new_[84109]_ , \new_[84112]_ ,
    \new_[84115]_ , \new_[84116]_ , \new_[84117]_ , \new_[84120]_ ,
    \new_[84123]_ , \new_[84124]_ , \new_[84127]_ , \new_[84130]_ ,
    \new_[84131]_ , \new_[84132]_ , \new_[84136]_ , \new_[84137]_ ,
    \new_[84140]_ , \new_[84143]_ , \new_[84144]_ , \new_[84145]_ ,
    \new_[84148]_ , \new_[84151]_ , \new_[84152]_ , \new_[84155]_ ,
    \new_[84158]_ , \new_[84159]_ , \new_[84160]_ , \new_[84164]_ ,
    \new_[84165]_ , \new_[84168]_ , \new_[84171]_ , \new_[84172]_ ,
    \new_[84173]_ , \new_[84176]_ , \new_[84179]_ , \new_[84180]_ ,
    \new_[84183]_ , \new_[84186]_ , \new_[84187]_ , \new_[84188]_ ,
    \new_[84192]_ , \new_[84193]_ , \new_[84196]_ , \new_[84199]_ ,
    \new_[84200]_ , \new_[84201]_ , \new_[84204]_ , \new_[84207]_ ,
    \new_[84208]_ , \new_[84211]_ , \new_[84214]_ , \new_[84215]_ ,
    \new_[84216]_ , \new_[84220]_ , \new_[84221]_ , \new_[84224]_ ,
    \new_[84227]_ , \new_[84228]_ , \new_[84229]_ , \new_[84232]_ ,
    \new_[84235]_ , \new_[84236]_ , \new_[84239]_ , \new_[84242]_ ,
    \new_[84243]_ , \new_[84244]_ , \new_[84248]_ , \new_[84249]_ ,
    \new_[84252]_ , \new_[84255]_ , \new_[84256]_ , \new_[84257]_ ,
    \new_[84260]_ , \new_[84263]_ , \new_[84264]_ , \new_[84267]_ ,
    \new_[84270]_ , \new_[84271]_ , \new_[84272]_ , \new_[84276]_ ,
    \new_[84277]_ , \new_[84280]_ , \new_[84283]_ , \new_[84284]_ ,
    \new_[84285]_ , \new_[84288]_ , \new_[84291]_ , \new_[84292]_ ,
    \new_[84295]_ , \new_[84298]_ , \new_[84299]_ , \new_[84300]_ ,
    \new_[84304]_ , \new_[84305]_ , \new_[84308]_ , \new_[84311]_ ,
    \new_[84312]_ , \new_[84313]_ , \new_[84316]_ , \new_[84319]_ ,
    \new_[84320]_ , \new_[84323]_ , \new_[84326]_ , \new_[84327]_ ,
    \new_[84328]_ , \new_[84332]_ , \new_[84333]_ , \new_[84336]_ ,
    \new_[84339]_ , \new_[84340]_ , \new_[84341]_ , \new_[84344]_ ,
    \new_[84347]_ , \new_[84348]_ , \new_[84351]_ , \new_[84354]_ ,
    \new_[84355]_ , \new_[84356]_ , \new_[84360]_ , \new_[84361]_ ,
    \new_[84364]_ , \new_[84367]_ , \new_[84368]_ , \new_[84369]_ ,
    \new_[84372]_ , \new_[84375]_ , \new_[84376]_ , \new_[84379]_ ,
    \new_[84382]_ , \new_[84383]_ , \new_[84384]_ , \new_[84388]_ ,
    \new_[84389]_ , \new_[84392]_ , \new_[84395]_ , \new_[84396]_ ,
    \new_[84397]_ , \new_[84400]_ , \new_[84403]_ , \new_[84404]_ ,
    \new_[84407]_ , \new_[84410]_ , \new_[84411]_ , \new_[84412]_ ,
    \new_[84416]_ , \new_[84417]_ , \new_[84420]_ , \new_[84423]_ ,
    \new_[84424]_ , \new_[84425]_ , \new_[84428]_ , \new_[84431]_ ,
    \new_[84432]_ , \new_[84435]_ , \new_[84438]_ , \new_[84439]_ ,
    \new_[84440]_ , \new_[84444]_ , \new_[84445]_ , \new_[84448]_ ,
    \new_[84451]_ , \new_[84452]_ , \new_[84453]_ , \new_[84456]_ ,
    \new_[84459]_ , \new_[84460]_ , \new_[84463]_ , \new_[84466]_ ,
    \new_[84467]_ , \new_[84468]_ , \new_[84472]_ , \new_[84473]_ ,
    \new_[84476]_ , \new_[84479]_ , \new_[84480]_ , \new_[84481]_ ,
    \new_[84484]_ , \new_[84487]_ , \new_[84488]_ , \new_[84491]_ ,
    \new_[84494]_ , \new_[84495]_ , \new_[84496]_ , \new_[84500]_ ,
    \new_[84501]_ , \new_[84504]_ , \new_[84507]_ , \new_[84508]_ ,
    \new_[84509]_ , \new_[84512]_ , \new_[84515]_ , \new_[84516]_ ,
    \new_[84519]_ , \new_[84522]_ , \new_[84523]_ , \new_[84524]_ ,
    \new_[84528]_ , \new_[84529]_ , \new_[84532]_ , \new_[84535]_ ,
    \new_[84536]_ , \new_[84537]_ , \new_[84540]_ , \new_[84543]_ ,
    \new_[84544]_ , \new_[84547]_ , \new_[84550]_ , \new_[84551]_ ,
    \new_[84552]_ , \new_[84556]_ , \new_[84557]_ , \new_[84560]_ ,
    \new_[84563]_ , \new_[84564]_ , \new_[84565]_ , \new_[84568]_ ,
    \new_[84571]_ , \new_[84572]_ , \new_[84575]_ , \new_[84578]_ ,
    \new_[84579]_ , \new_[84580]_ , \new_[84584]_ , \new_[84585]_ ,
    \new_[84588]_ , \new_[84591]_ , \new_[84592]_ , \new_[84593]_ ,
    \new_[84596]_ , \new_[84599]_ , \new_[84600]_ , \new_[84603]_ ,
    \new_[84606]_ , \new_[84607]_ , \new_[84608]_ , \new_[84612]_ ,
    \new_[84613]_ , \new_[84616]_ , \new_[84619]_ , \new_[84620]_ ,
    \new_[84621]_ , \new_[84624]_ , \new_[84627]_ , \new_[84628]_ ,
    \new_[84631]_ , \new_[84634]_ , \new_[84635]_ , \new_[84636]_ ,
    \new_[84640]_ , \new_[84641]_ , \new_[84644]_ , \new_[84647]_ ,
    \new_[84648]_ , \new_[84649]_ , \new_[84652]_ , \new_[84655]_ ,
    \new_[84656]_ , \new_[84659]_ , \new_[84662]_ , \new_[84663]_ ,
    \new_[84664]_ , \new_[84668]_ , \new_[84669]_ , \new_[84672]_ ,
    \new_[84675]_ , \new_[84676]_ , \new_[84677]_ , \new_[84680]_ ,
    \new_[84683]_ , \new_[84684]_ , \new_[84687]_ , \new_[84690]_ ,
    \new_[84691]_ , \new_[84692]_ , \new_[84696]_ , \new_[84697]_ ,
    \new_[84700]_ , \new_[84703]_ , \new_[84704]_ , \new_[84705]_ ,
    \new_[84708]_ , \new_[84711]_ , \new_[84712]_ , \new_[84715]_ ,
    \new_[84718]_ , \new_[84719]_ , \new_[84720]_ , \new_[84724]_ ,
    \new_[84725]_ , \new_[84728]_ , \new_[84731]_ , \new_[84732]_ ,
    \new_[84733]_ , \new_[84736]_ , \new_[84739]_ , \new_[84740]_ ,
    \new_[84743]_ , \new_[84746]_ , \new_[84747]_ , \new_[84748]_ ,
    \new_[84752]_ , \new_[84753]_ , \new_[84756]_ , \new_[84759]_ ,
    \new_[84760]_ , \new_[84761]_ , \new_[84764]_ , \new_[84767]_ ,
    \new_[84768]_ , \new_[84771]_ , \new_[84774]_ , \new_[84775]_ ,
    \new_[84776]_ , \new_[84780]_ , \new_[84781]_ , \new_[84784]_ ,
    \new_[84787]_ , \new_[84788]_ , \new_[84789]_ , \new_[84792]_ ,
    \new_[84795]_ , \new_[84796]_ , \new_[84799]_ , \new_[84802]_ ,
    \new_[84803]_ , \new_[84804]_ , \new_[84808]_ , \new_[84809]_ ,
    \new_[84812]_ , \new_[84815]_ , \new_[84816]_ , \new_[84817]_ ,
    \new_[84820]_ , \new_[84823]_ , \new_[84824]_ , \new_[84827]_ ,
    \new_[84830]_ , \new_[84831]_ , \new_[84832]_ , \new_[84836]_ ,
    \new_[84837]_ , \new_[84840]_ , \new_[84843]_ , \new_[84844]_ ,
    \new_[84845]_ , \new_[84848]_ , \new_[84851]_ , \new_[84852]_ ,
    \new_[84855]_ , \new_[84858]_ , \new_[84859]_ , \new_[84860]_ ,
    \new_[84864]_ , \new_[84865]_ , \new_[84868]_ , \new_[84871]_ ,
    \new_[84872]_ , \new_[84873]_ , \new_[84876]_ , \new_[84879]_ ,
    \new_[84880]_ , \new_[84883]_ , \new_[84886]_ , \new_[84887]_ ,
    \new_[84888]_ , \new_[84892]_ , \new_[84893]_ , \new_[84896]_ ,
    \new_[84899]_ , \new_[84900]_ , \new_[84901]_ , \new_[84904]_ ,
    \new_[84907]_ , \new_[84908]_ , \new_[84911]_ , \new_[84914]_ ,
    \new_[84915]_ , \new_[84916]_ , \new_[84920]_ , \new_[84921]_ ,
    \new_[84924]_ , \new_[84927]_ , \new_[84928]_ , \new_[84929]_ ,
    \new_[84932]_ , \new_[84935]_ , \new_[84936]_ , \new_[84939]_ ,
    \new_[84942]_ , \new_[84943]_ , \new_[84944]_ , \new_[84948]_ ,
    \new_[84949]_ , \new_[84952]_ , \new_[84955]_ , \new_[84956]_ ,
    \new_[84957]_ , \new_[84960]_ , \new_[84963]_ , \new_[84964]_ ,
    \new_[84967]_ , \new_[84970]_ , \new_[84971]_ , \new_[84972]_ ,
    \new_[84976]_ , \new_[84977]_ , \new_[84980]_ , \new_[84983]_ ,
    \new_[84984]_ , \new_[84985]_ , \new_[84988]_ , \new_[84991]_ ,
    \new_[84992]_ , \new_[84995]_ , \new_[84998]_ , \new_[84999]_ ,
    \new_[85000]_ , \new_[85004]_ , \new_[85005]_ , \new_[85008]_ ,
    \new_[85011]_ , \new_[85012]_ , \new_[85013]_ , \new_[85016]_ ,
    \new_[85019]_ , \new_[85020]_ , \new_[85023]_ , \new_[85026]_ ,
    \new_[85027]_ , \new_[85028]_ , \new_[85032]_ , \new_[85033]_ ,
    \new_[85036]_ , \new_[85039]_ , \new_[85040]_ , \new_[85041]_ ,
    \new_[85044]_ , \new_[85047]_ , \new_[85048]_ , \new_[85051]_ ,
    \new_[85054]_ , \new_[85055]_ , \new_[85056]_ , \new_[85060]_ ,
    \new_[85061]_ , \new_[85064]_ , \new_[85067]_ , \new_[85068]_ ,
    \new_[85069]_ , \new_[85072]_ , \new_[85075]_ , \new_[85076]_ ,
    \new_[85079]_ , \new_[85082]_ , \new_[85083]_ , \new_[85084]_ ,
    \new_[85088]_ , \new_[85089]_ , \new_[85092]_ , \new_[85095]_ ,
    \new_[85096]_ , \new_[85097]_ , \new_[85100]_ , \new_[85103]_ ,
    \new_[85104]_ , \new_[85107]_ , \new_[85110]_ , \new_[85111]_ ,
    \new_[85112]_ , \new_[85116]_ , \new_[85117]_ , \new_[85120]_ ,
    \new_[85123]_ , \new_[85124]_ , \new_[85125]_ , \new_[85128]_ ,
    \new_[85131]_ , \new_[85132]_ , \new_[85135]_ , \new_[85138]_ ,
    \new_[85139]_ , \new_[85140]_ , \new_[85144]_ , \new_[85145]_ ,
    \new_[85148]_ , \new_[85151]_ , \new_[85152]_ , \new_[85153]_ ,
    \new_[85156]_ , \new_[85159]_ , \new_[85160]_ , \new_[85163]_ ,
    \new_[85166]_ , \new_[85167]_ , \new_[85168]_ , \new_[85172]_ ,
    \new_[85173]_ , \new_[85176]_ , \new_[85179]_ , \new_[85180]_ ,
    \new_[85181]_ , \new_[85184]_ , \new_[85187]_ , \new_[85188]_ ,
    \new_[85191]_ , \new_[85194]_ , \new_[85195]_ , \new_[85196]_ ,
    \new_[85200]_ , \new_[85201]_ , \new_[85204]_ , \new_[85207]_ ,
    \new_[85208]_ , \new_[85209]_ , \new_[85212]_ , \new_[85215]_ ,
    \new_[85216]_ , \new_[85219]_ , \new_[85222]_ , \new_[85223]_ ,
    \new_[85224]_ , \new_[85228]_ , \new_[85229]_ , \new_[85232]_ ,
    \new_[85235]_ , \new_[85236]_ , \new_[85237]_ , \new_[85240]_ ,
    \new_[85243]_ , \new_[85244]_ , \new_[85247]_ , \new_[85250]_ ,
    \new_[85251]_ , \new_[85252]_ , \new_[85256]_ , \new_[85257]_ ,
    \new_[85260]_ , \new_[85263]_ , \new_[85264]_ , \new_[85265]_ ,
    \new_[85268]_ , \new_[85271]_ , \new_[85272]_ , \new_[85275]_ ,
    \new_[85278]_ , \new_[85279]_ , \new_[85280]_ , \new_[85284]_ ,
    \new_[85285]_ , \new_[85288]_ , \new_[85291]_ , \new_[85292]_ ,
    \new_[85293]_ , \new_[85296]_ , \new_[85299]_ , \new_[85300]_ ,
    \new_[85303]_ , \new_[85306]_ , \new_[85307]_ , \new_[85308]_ ,
    \new_[85312]_ , \new_[85313]_ , \new_[85316]_ , \new_[85319]_ ,
    \new_[85320]_ , \new_[85321]_ , \new_[85324]_ , \new_[85327]_ ,
    \new_[85328]_ , \new_[85331]_ , \new_[85334]_ , \new_[85335]_ ,
    \new_[85336]_ , \new_[85340]_ , \new_[85341]_ , \new_[85344]_ ,
    \new_[85347]_ , \new_[85348]_ , \new_[85349]_ , \new_[85352]_ ,
    \new_[85355]_ , \new_[85356]_ , \new_[85359]_ , \new_[85362]_ ,
    \new_[85363]_ , \new_[85364]_ , \new_[85368]_ , \new_[85369]_ ,
    \new_[85372]_ , \new_[85375]_ , \new_[85376]_ , \new_[85377]_ ,
    \new_[85380]_ , \new_[85383]_ , \new_[85384]_ , \new_[85387]_ ,
    \new_[85390]_ , \new_[85391]_ , \new_[85392]_ , \new_[85396]_ ,
    \new_[85397]_ , \new_[85400]_ , \new_[85403]_ , \new_[85404]_ ,
    \new_[85405]_ , \new_[85408]_ , \new_[85411]_ , \new_[85412]_ ,
    \new_[85415]_ , \new_[85418]_ , \new_[85419]_ , \new_[85420]_ ,
    \new_[85424]_ , \new_[85425]_ , \new_[85428]_ , \new_[85431]_ ,
    \new_[85432]_ , \new_[85433]_ , \new_[85436]_ , \new_[85439]_ ,
    \new_[85440]_ , \new_[85443]_ , \new_[85446]_ , \new_[85447]_ ,
    \new_[85448]_ , \new_[85452]_ , \new_[85453]_ , \new_[85456]_ ,
    \new_[85459]_ , \new_[85460]_ , \new_[85461]_ , \new_[85464]_ ,
    \new_[85467]_ , \new_[85468]_ , \new_[85471]_ , \new_[85474]_ ,
    \new_[85475]_ , \new_[85476]_ , \new_[85480]_ , \new_[85481]_ ,
    \new_[85484]_ , \new_[85487]_ , \new_[85488]_ , \new_[85489]_ ,
    \new_[85492]_ , \new_[85495]_ , \new_[85496]_ , \new_[85499]_ ,
    \new_[85502]_ , \new_[85503]_ , \new_[85504]_ , \new_[85508]_ ,
    \new_[85509]_ , \new_[85512]_ , \new_[85515]_ , \new_[85516]_ ,
    \new_[85517]_ , \new_[85520]_ , \new_[85523]_ , \new_[85524]_ ,
    \new_[85527]_ , \new_[85530]_ , \new_[85531]_ , \new_[85532]_ ,
    \new_[85536]_ , \new_[85537]_ , \new_[85540]_ , \new_[85543]_ ,
    \new_[85544]_ , \new_[85545]_ , \new_[85548]_ , \new_[85551]_ ,
    \new_[85552]_ , \new_[85555]_ , \new_[85558]_ , \new_[85559]_ ,
    \new_[85560]_ , \new_[85564]_ , \new_[85565]_ , \new_[85568]_ ,
    \new_[85571]_ , \new_[85572]_ , \new_[85573]_ , \new_[85576]_ ,
    \new_[85579]_ , \new_[85580]_ , \new_[85583]_ , \new_[85586]_ ,
    \new_[85587]_ , \new_[85588]_ , \new_[85592]_ , \new_[85593]_ ,
    \new_[85596]_ , \new_[85599]_ , \new_[85600]_ , \new_[85601]_ ,
    \new_[85604]_ , \new_[85607]_ , \new_[85608]_ , \new_[85611]_ ,
    \new_[85614]_ , \new_[85615]_ , \new_[85616]_ , \new_[85620]_ ,
    \new_[85621]_ , \new_[85624]_ , \new_[85627]_ , \new_[85628]_ ,
    \new_[85629]_ , \new_[85632]_ , \new_[85635]_ , \new_[85636]_ ,
    \new_[85639]_ , \new_[85642]_ , \new_[85643]_ , \new_[85644]_ ,
    \new_[85648]_ , \new_[85649]_ , \new_[85652]_ , \new_[85655]_ ,
    \new_[85656]_ , \new_[85657]_ , \new_[85660]_ , \new_[85663]_ ,
    \new_[85664]_ , \new_[85667]_ , \new_[85670]_ , \new_[85671]_ ,
    \new_[85672]_ , \new_[85676]_ , \new_[85677]_ , \new_[85680]_ ,
    \new_[85683]_ , \new_[85684]_ , \new_[85685]_ , \new_[85688]_ ,
    \new_[85691]_ , \new_[85692]_ , \new_[85695]_ , \new_[85698]_ ,
    \new_[85699]_ , \new_[85700]_ , \new_[85704]_ , \new_[85705]_ ,
    \new_[85708]_ , \new_[85711]_ , \new_[85712]_ , \new_[85713]_ ,
    \new_[85716]_ , \new_[85719]_ , \new_[85720]_ , \new_[85723]_ ,
    \new_[85726]_ , \new_[85727]_ , \new_[85728]_ , \new_[85732]_ ,
    \new_[85733]_ , \new_[85736]_ , \new_[85739]_ , \new_[85740]_ ,
    \new_[85741]_ , \new_[85744]_ , \new_[85747]_ , \new_[85748]_ ,
    \new_[85751]_ , \new_[85754]_ , \new_[85755]_ , \new_[85756]_ ,
    \new_[85760]_ , \new_[85761]_ , \new_[85764]_ , \new_[85767]_ ,
    \new_[85768]_ , \new_[85769]_ , \new_[85772]_ , \new_[85775]_ ,
    \new_[85776]_ , \new_[85779]_ , \new_[85782]_ , \new_[85783]_ ,
    \new_[85784]_ , \new_[85788]_ , \new_[85789]_ , \new_[85792]_ ,
    \new_[85795]_ , \new_[85796]_ , \new_[85797]_ , \new_[85800]_ ,
    \new_[85803]_ , \new_[85804]_ , \new_[85807]_ , \new_[85810]_ ,
    \new_[85811]_ , \new_[85812]_ , \new_[85816]_ , \new_[85817]_ ,
    \new_[85820]_ , \new_[85823]_ , \new_[85824]_ , \new_[85825]_ ,
    \new_[85828]_ , \new_[85831]_ , \new_[85832]_ , \new_[85835]_ ,
    \new_[85838]_ , \new_[85839]_ , \new_[85840]_ , \new_[85844]_ ,
    \new_[85845]_ , \new_[85848]_ , \new_[85851]_ , \new_[85852]_ ,
    \new_[85853]_ , \new_[85856]_ , \new_[85859]_ , \new_[85860]_ ,
    \new_[85863]_ , \new_[85866]_ , \new_[85867]_ , \new_[85868]_ ,
    \new_[85872]_ , \new_[85873]_ , \new_[85876]_ , \new_[85879]_ ,
    \new_[85880]_ , \new_[85881]_ , \new_[85884]_ , \new_[85887]_ ,
    \new_[85888]_ , \new_[85891]_ , \new_[85894]_ , \new_[85895]_ ,
    \new_[85896]_ , \new_[85900]_ , \new_[85901]_ , \new_[85904]_ ,
    \new_[85907]_ , \new_[85908]_ , \new_[85909]_ , \new_[85912]_ ,
    \new_[85915]_ , \new_[85916]_ , \new_[85919]_ , \new_[85922]_ ,
    \new_[85923]_ , \new_[85924]_ , \new_[85928]_ , \new_[85929]_ ,
    \new_[85932]_ , \new_[85935]_ , \new_[85936]_ , \new_[85937]_ ,
    \new_[85940]_ , \new_[85943]_ , \new_[85944]_ , \new_[85947]_ ,
    \new_[85950]_ , \new_[85951]_ , \new_[85952]_ , \new_[85956]_ ,
    \new_[85957]_ , \new_[85960]_ , \new_[85963]_ , \new_[85964]_ ,
    \new_[85965]_ , \new_[85968]_ , \new_[85971]_ , \new_[85972]_ ,
    \new_[85975]_ , \new_[85978]_ , \new_[85979]_ , \new_[85980]_ ,
    \new_[85984]_ , \new_[85985]_ , \new_[85988]_ , \new_[85991]_ ,
    \new_[85992]_ , \new_[85993]_ , \new_[85996]_ , \new_[85999]_ ,
    \new_[86000]_ , \new_[86003]_ , \new_[86006]_ , \new_[86007]_ ,
    \new_[86008]_ , \new_[86012]_ , \new_[86013]_ , \new_[86016]_ ,
    \new_[86019]_ , \new_[86020]_ , \new_[86021]_ , \new_[86024]_ ,
    \new_[86027]_ , \new_[86028]_ , \new_[86031]_ , \new_[86034]_ ,
    \new_[86035]_ , \new_[86036]_ , \new_[86040]_ , \new_[86041]_ ,
    \new_[86044]_ , \new_[86047]_ , \new_[86048]_ , \new_[86049]_ ,
    \new_[86052]_ , \new_[86055]_ , \new_[86056]_ , \new_[86059]_ ,
    \new_[86062]_ , \new_[86063]_ , \new_[86064]_ , \new_[86068]_ ,
    \new_[86069]_ , \new_[86072]_ , \new_[86075]_ , \new_[86076]_ ,
    \new_[86077]_ , \new_[86080]_ , \new_[86083]_ , \new_[86084]_ ,
    \new_[86087]_ , \new_[86090]_ , \new_[86091]_ , \new_[86092]_ ,
    \new_[86096]_ , \new_[86097]_ , \new_[86100]_ , \new_[86103]_ ,
    \new_[86104]_ , \new_[86105]_ , \new_[86108]_ , \new_[86111]_ ,
    \new_[86112]_ , \new_[86115]_ , \new_[86118]_ , \new_[86119]_ ,
    \new_[86120]_ , \new_[86124]_ , \new_[86125]_ , \new_[86128]_ ,
    \new_[86131]_ , \new_[86132]_ , \new_[86133]_ , \new_[86136]_ ,
    \new_[86139]_ , \new_[86140]_ , \new_[86143]_ , \new_[86146]_ ,
    \new_[86147]_ , \new_[86148]_ , \new_[86152]_ , \new_[86153]_ ,
    \new_[86156]_ , \new_[86159]_ , \new_[86160]_ , \new_[86161]_ ,
    \new_[86164]_ , \new_[86167]_ , \new_[86168]_ , \new_[86171]_ ,
    \new_[86174]_ , \new_[86175]_ , \new_[86176]_ , \new_[86180]_ ,
    \new_[86181]_ , \new_[86184]_ , \new_[86187]_ , \new_[86188]_ ,
    \new_[86189]_ , \new_[86192]_ , \new_[86195]_ , \new_[86196]_ ,
    \new_[86199]_ , \new_[86202]_ , \new_[86203]_ , \new_[86204]_ ,
    \new_[86208]_ , \new_[86209]_ , \new_[86212]_ , \new_[86215]_ ,
    \new_[86216]_ , \new_[86217]_ , \new_[86220]_ , \new_[86223]_ ,
    \new_[86224]_ , \new_[86227]_ , \new_[86230]_ , \new_[86231]_ ,
    \new_[86232]_ , \new_[86236]_ , \new_[86237]_ , \new_[86240]_ ,
    \new_[86243]_ , \new_[86244]_ , \new_[86245]_ , \new_[86248]_ ,
    \new_[86251]_ , \new_[86252]_ , \new_[86255]_ , \new_[86258]_ ,
    \new_[86259]_ , \new_[86260]_ , \new_[86264]_ , \new_[86265]_ ,
    \new_[86268]_ , \new_[86271]_ , \new_[86272]_ , \new_[86273]_ ,
    \new_[86276]_ , \new_[86279]_ , \new_[86280]_ , \new_[86283]_ ,
    \new_[86286]_ , \new_[86287]_ , \new_[86288]_ , \new_[86292]_ ,
    \new_[86293]_ , \new_[86296]_ , \new_[86299]_ , \new_[86300]_ ,
    \new_[86301]_ , \new_[86304]_ , \new_[86307]_ , \new_[86308]_ ,
    \new_[86311]_ , \new_[86314]_ , \new_[86315]_ , \new_[86316]_ ,
    \new_[86320]_ , \new_[86321]_ , \new_[86324]_ , \new_[86327]_ ,
    \new_[86328]_ , \new_[86329]_ , \new_[86332]_ , \new_[86335]_ ,
    \new_[86336]_ , \new_[86339]_ , \new_[86342]_ , \new_[86343]_ ,
    \new_[86344]_ , \new_[86348]_ , \new_[86349]_ , \new_[86352]_ ,
    \new_[86355]_ , \new_[86356]_ , \new_[86357]_ , \new_[86360]_ ,
    \new_[86363]_ , \new_[86364]_ , \new_[86367]_ , \new_[86370]_ ,
    \new_[86371]_ , \new_[86372]_ , \new_[86376]_ , \new_[86377]_ ,
    \new_[86380]_ , \new_[86383]_ , \new_[86384]_ , \new_[86385]_ ,
    \new_[86388]_ , \new_[86391]_ , \new_[86392]_ , \new_[86395]_ ,
    \new_[86398]_ , \new_[86399]_ , \new_[86400]_ , \new_[86404]_ ,
    \new_[86405]_ , \new_[86408]_ , \new_[86411]_ , \new_[86412]_ ,
    \new_[86413]_ , \new_[86416]_ , \new_[86419]_ , \new_[86420]_ ,
    \new_[86423]_ , \new_[86426]_ , \new_[86427]_ , \new_[86428]_ ,
    \new_[86432]_ , \new_[86433]_ , \new_[86436]_ , \new_[86439]_ ,
    \new_[86440]_ , \new_[86441]_ , \new_[86444]_ , \new_[86447]_ ,
    \new_[86448]_ , \new_[86451]_ , \new_[86454]_ , \new_[86455]_ ,
    \new_[86456]_ , \new_[86460]_ , \new_[86461]_ , \new_[86464]_ ,
    \new_[86467]_ , \new_[86468]_ , \new_[86469]_ , \new_[86472]_ ,
    \new_[86475]_ , \new_[86476]_ , \new_[86479]_ , \new_[86482]_ ,
    \new_[86483]_ , \new_[86484]_ , \new_[86488]_ , \new_[86489]_ ,
    \new_[86492]_ , \new_[86495]_ , \new_[86496]_ , \new_[86497]_ ,
    \new_[86500]_ , \new_[86503]_ , \new_[86504]_ , \new_[86507]_ ,
    \new_[86510]_ , \new_[86511]_ , \new_[86512]_ , \new_[86516]_ ,
    \new_[86517]_ , \new_[86520]_ , \new_[86523]_ , \new_[86524]_ ,
    \new_[86525]_ , \new_[86528]_ , \new_[86531]_ , \new_[86532]_ ,
    \new_[86535]_ , \new_[86538]_ , \new_[86539]_ , \new_[86540]_ ,
    \new_[86544]_ , \new_[86545]_ , \new_[86548]_ , \new_[86551]_ ,
    \new_[86552]_ , \new_[86553]_ , \new_[86556]_ , \new_[86559]_ ,
    \new_[86560]_ , \new_[86563]_ , \new_[86566]_ , \new_[86567]_ ,
    \new_[86568]_ , \new_[86572]_ , \new_[86573]_ , \new_[86576]_ ,
    \new_[86579]_ , \new_[86580]_ , \new_[86581]_ , \new_[86584]_ ,
    \new_[86587]_ , \new_[86588]_ , \new_[86591]_ , \new_[86594]_ ,
    \new_[86595]_ , \new_[86596]_ , \new_[86600]_ , \new_[86601]_ ,
    \new_[86604]_ , \new_[86607]_ , \new_[86608]_ , \new_[86609]_ ,
    \new_[86612]_ , \new_[86615]_ , \new_[86616]_ , \new_[86619]_ ,
    \new_[86622]_ , \new_[86623]_ , \new_[86624]_ , \new_[86628]_ ,
    \new_[86629]_ , \new_[86632]_ , \new_[86635]_ , \new_[86636]_ ,
    \new_[86637]_ , \new_[86640]_ , \new_[86643]_ , \new_[86644]_ ,
    \new_[86647]_ , \new_[86650]_ , \new_[86651]_ , \new_[86652]_ ,
    \new_[86656]_ , \new_[86657]_ , \new_[86660]_ , \new_[86663]_ ,
    \new_[86664]_ , \new_[86665]_ , \new_[86668]_ , \new_[86671]_ ,
    \new_[86672]_ , \new_[86675]_ , \new_[86678]_ , \new_[86679]_ ,
    \new_[86680]_ , \new_[86684]_ , \new_[86685]_ , \new_[86688]_ ,
    \new_[86691]_ , \new_[86692]_ , \new_[86693]_ , \new_[86696]_ ,
    \new_[86699]_ , \new_[86700]_ , \new_[86703]_ , \new_[86706]_ ,
    \new_[86707]_ , \new_[86708]_ , \new_[86712]_ , \new_[86713]_ ,
    \new_[86716]_ , \new_[86719]_ , \new_[86720]_ , \new_[86721]_ ,
    \new_[86724]_ , \new_[86727]_ , \new_[86728]_ , \new_[86731]_ ,
    \new_[86734]_ , \new_[86735]_ , \new_[86736]_ , \new_[86740]_ ,
    \new_[86741]_ , \new_[86744]_ , \new_[86747]_ , \new_[86748]_ ,
    \new_[86749]_ , \new_[86752]_ , \new_[86755]_ , \new_[86756]_ ,
    \new_[86759]_ , \new_[86762]_ , \new_[86763]_ , \new_[86764]_ ,
    \new_[86768]_ , \new_[86769]_ , \new_[86772]_ , \new_[86775]_ ,
    \new_[86776]_ , \new_[86777]_ , \new_[86780]_ , \new_[86783]_ ,
    \new_[86784]_ , \new_[86787]_ , \new_[86790]_ , \new_[86791]_ ,
    \new_[86792]_ , \new_[86796]_ , \new_[86797]_ , \new_[86800]_ ,
    \new_[86803]_ , \new_[86804]_ , \new_[86805]_ , \new_[86808]_ ,
    \new_[86811]_ , \new_[86812]_ , \new_[86815]_ , \new_[86818]_ ,
    \new_[86819]_ , \new_[86820]_ , \new_[86824]_ , \new_[86825]_ ,
    \new_[86828]_ , \new_[86831]_ , \new_[86832]_ , \new_[86833]_ ,
    \new_[86836]_ , \new_[86839]_ , \new_[86840]_ , \new_[86843]_ ,
    \new_[86846]_ , \new_[86847]_ , \new_[86848]_ , \new_[86852]_ ,
    \new_[86853]_ , \new_[86856]_ , \new_[86859]_ , \new_[86860]_ ,
    \new_[86861]_ , \new_[86864]_ , \new_[86867]_ , \new_[86868]_ ,
    \new_[86871]_ , \new_[86874]_ , \new_[86875]_ , \new_[86876]_ ,
    \new_[86880]_ , \new_[86881]_ , \new_[86884]_ , \new_[86887]_ ,
    \new_[86888]_ , \new_[86889]_ , \new_[86892]_ , \new_[86895]_ ,
    \new_[86896]_ , \new_[86899]_ , \new_[86902]_ , \new_[86903]_ ,
    \new_[86904]_ , \new_[86908]_ , \new_[86909]_ , \new_[86912]_ ,
    \new_[86915]_ , \new_[86916]_ , \new_[86917]_ , \new_[86920]_ ,
    \new_[86923]_ , \new_[86924]_ , \new_[86927]_ , \new_[86930]_ ,
    \new_[86931]_ , \new_[86932]_ , \new_[86936]_ , \new_[86937]_ ,
    \new_[86940]_ , \new_[86943]_ , \new_[86944]_ , \new_[86945]_ ,
    \new_[86948]_ , \new_[86951]_ , \new_[86952]_ , \new_[86955]_ ,
    \new_[86958]_ , \new_[86959]_ , \new_[86960]_ , \new_[86964]_ ,
    \new_[86965]_ , \new_[86968]_ , \new_[86971]_ , \new_[86972]_ ,
    \new_[86973]_ , \new_[86976]_ , \new_[86979]_ , \new_[86980]_ ,
    \new_[86983]_ , \new_[86986]_ , \new_[86987]_ , \new_[86988]_ ,
    \new_[86992]_ , \new_[86993]_ , \new_[86996]_ , \new_[86999]_ ,
    \new_[87000]_ , \new_[87001]_ , \new_[87004]_ , \new_[87007]_ ,
    \new_[87008]_ , \new_[87011]_ , \new_[87014]_ , \new_[87015]_ ,
    \new_[87016]_ , \new_[87020]_ , \new_[87021]_ , \new_[87024]_ ,
    \new_[87027]_ , \new_[87028]_ , \new_[87029]_ , \new_[87032]_ ,
    \new_[87035]_ , \new_[87036]_ , \new_[87039]_ , \new_[87042]_ ,
    \new_[87043]_ , \new_[87044]_ , \new_[87048]_ , \new_[87049]_ ,
    \new_[87052]_ , \new_[87055]_ , \new_[87056]_ , \new_[87057]_ ,
    \new_[87060]_ , \new_[87063]_ , \new_[87064]_ , \new_[87067]_ ,
    \new_[87070]_ , \new_[87071]_ , \new_[87072]_ , \new_[87076]_ ,
    \new_[87077]_ , \new_[87080]_ , \new_[87083]_ , \new_[87084]_ ,
    \new_[87085]_ , \new_[87088]_ , \new_[87091]_ , \new_[87092]_ ,
    \new_[87095]_ , \new_[87098]_ , \new_[87099]_ , \new_[87100]_ ,
    \new_[87104]_ , \new_[87105]_ , \new_[87108]_ , \new_[87111]_ ,
    \new_[87112]_ , \new_[87113]_ , \new_[87116]_ , \new_[87119]_ ,
    \new_[87120]_ , \new_[87123]_ , \new_[87126]_ , \new_[87127]_ ,
    \new_[87128]_ , \new_[87132]_ , \new_[87133]_ , \new_[87136]_ ,
    \new_[87139]_ , \new_[87140]_ , \new_[87141]_ , \new_[87144]_ ,
    \new_[87147]_ , \new_[87148]_ , \new_[87151]_ , \new_[87154]_ ,
    \new_[87155]_ , \new_[87156]_ , \new_[87160]_ , \new_[87161]_ ,
    \new_[87164]_ , \new_[87167]_ , \new_[87168]_ , \new_[87169]_ ,
    \new_[87172]_ , \new_[87175]_ , \new_[87176]_ , \new_[87179]_ ,
    \new_[87182]_ , \new_[87183]_ , \new_[87184]_ , \new_[87188]_ ,
    \new_[87189]_ , \new_[87192]_ , \new_[87195]_ , \new_[87196]_ ,
    \new_[87197]_ , \new_[87200]_ , \new_[87203]_ , \new_[87204]_ ,
    \new_[87207]_ , \new_[87210]_ , \new_[87211]_ , \new_[87212]_ ,
    \new_[87216]_ , \new_[87217]_ , \new_[87220]_ , \new_[87223]_ ,
    \new_[87224]_ , \new_[87225]_ , \new_[87228]_ , \new_[87231]_ ,
    \new_[87232]_ , \new_[87235]_ , \new_[87238]_ , \new_[87239]_ ,
    \new_[87240]_ , \new_[87244]_ , \new_[87245]_ , \new_[87248]_ ,
    \new_[87251]_ , \new_[87252]_ , \new_[87253]_ , \new_[87256]_ ,
    \new_[87259]_ , \new_[87260]_ , \new_[87263]_ , \new_[87266]_ ,
    \new_[87267]_ , \new_[87268]_ , \new_[87272]_ , \new_[87273]_ ,
    \new_[87276]_ , \new_[87279]_ , \new_[87280]_ , \new_[87281]_ ,
    \new_[87284]_ , \new_[87287]_ , \new_[87288]_ , \new_[87291]_ ,
    \new_[87294]_ , \new_[87295]_ , \new_[87296]_ , \new_[87300]_ ,
    \new_[87301]_ , \new_[87304]_ , \new_[87307]_ , \new_[87308]_ ,
    \new_[87309]_ , \new_[87312]_ , \new_[87315]_ , \new_[87316]_ ,
    \new_[87319]_ , \new_[87322]_ , \new_[87323]_ , \new_[87324]_ ,
    \new_[87328]_ , \new_[87329]_ , \new_[87332]_ , \new_[87335]_ ,
    \new_[87336]_ , \new_[87337]_ , \new_[87340]_ , \new_[87343]_ ,
    \new_[87344]_ , \new_[87347]_ , \new_[87350]_ , \new_[87351]_ ,
    \new_[87352]_ , \new_[87356]_ , \new_[87357]_ , \new_[87360]_ ,
    \new_[87363]_ , \new_[87364]_ , \new_[87365]_ , \new_[87368]_ ,
    \new_[87371]_ , \new_[87372]_ , \new_[87375]_ , \new_[87378]_ ,
    \new_[87379]_ , \new_[87380]_ , \new_[87384]_ , \new_[87385]_ ,
    \new_[87388]_ , \new_[87391]_ , \new_[87392]_ , \new_[87393]_ ,
    \new_[87396]_ , \new_[87399]_ , \new_[87400]_ , \new_[87403]_ ,
    \new_[87406]_ , \new_[87407]_ , \new_[87408]_ , \new_[87412]_ ,
    \new_[87413]_ , \new_[87416]_ , \new_[87419]_ , \new_[87420]_ ,
    \new_[87421]_ , \new_[87424]_ , \new_[87427]_ , \new_[87428]_ ,
    \new_[87431]_ , \new_[87434]_ , \new_[87435]_ , \new_[87436]_ ,
    \new_[87440]_ , \new_[87441]_ , \new_[87444]_ , \new_[87447]_ ,
    \new_[87448]_ , \new_[87449]_ , \new_[87452]_ , \new_[87455]_ ,
    \new_[87456]_ , \new_[87459]_ , \new_[87462]_ , \new_[87463]_ ,
    \new_[87464]_ , \new_[87468]_ , \new_[87469]_ , \new_[87472]_ ,
    \new_[87475]_ , \new_[87476]_ , \new_[87477]_ , \new_[87480]_ ,
    \new_[87483]_ , \new_[87484]_ , \new_[87487]_ , \new_[87490]_ ,
    \new_[87491]_ , \new_[87492]_ , \new_[87496]_ , \new_[87497]_ ,
    \new_[87500]_ , \new_[87503]_ , \new_[87504]_ , \new_[87505]_ ,
    \new_[87508]_ , \new_[87511]_ , \new_[87512]_ , \new_[87515]_ ,
    \new_[87518]_ , \new_[87519]_ , \new_[87520]_ , \new_[87524]_ ,
    \new_[87525]_ , \new_[87528]_ , \new_[87531]_ , \new_[87532]_ ,
    \new_[87533]_ , \new_[87536]_ , \new_[87539]_ , \new_[87540]_ ,
    \new_[87543]_ , \new_[87546]_ , \new_[87547]_ , \new_[87548]_ ,
    \new_[87552]_ , \new_[87553]_ , \new_[87556]_ , \new_[87559]_ ,
    \new_[87560]_ , \new_[87561]_ , \new_[87564]_ , \new_[87567]_ ,
    \new_[87568]_ , \new_[87571]_ , \new_[87574]_ , \new_[87575]_ ,
    \new_[87576]_ , \new_[87580]_ , \new_[87581]_ , \new_[87584]_ ,
    \new_[87587]_ , \new_[87588]_ , \new_[87589]_ , \new_[87592]_ ,
    \new_[87595]_ , \new_[87596]_ , \new_[87599]_ , \new_[87602]_ ,
    \new_[87603]_ , \new_[87604]_ , \new_[87608]_ , \new_[87609]_ ,
    \new_[87612]_ , \new_[87615]_ , \new_[87616]_ , \new_[87617]_ ,
    \new_[87620]_ , \new_[87623]_ , \new_[87624]_ , \new_[87627]_ ,
    \new_[87630]_ , \new_[87631]_ , \new_[87632]_ , \new_[87636]_ ,
    \new_[87637]_ , \new_[87640]_ , \new_[87643]_ , \new_[87644]_ ,
    \new_[87645]_ , \new_[87648]_ , \new_[87651]_ , \new_[87652]_ ,
    \new_[87655]_ , \new_[87658]_ , \new_[87659]_ , \new_[87660]_ ,
    \new_[87664]_ , \new_[87665]_ , \new_[87668]_ , \new_[87671]_ ,
    \new_[87672]_ , \new_[87673]_ , \new_[87676]_ , \new_[87679]_ ,
    \new_[87680]_ , \new_[87683]_ , \new_[87686]_ , \new_[87687]_ ,
    \new_[87688]_ , \new_[87692]_ , \new_[87693]_ , \new_[87696]_ ,
    \new_[87699]_ , \new_[87700]_ , \new_[87701]_ , \new_[87704]_ ,
    \new_[87707]_ , \new_[87708]_ , \new_[87711]_ , \new_[87714]_ ,
    \new_[87715]_ , \new_[87716]_ , \new_[87720]_ , \new_[87721]_ ,
    \new_[87724]_ , \new_[87727]_ , \new_[87728]_ , \new_[87729]_ ,
    \new_[87732]_ , \new_[87735]_ , \new_[87736]_ , \new_[87739]_ ,
    \new_[87742]_ , \new_[87743]_ , \new_[87744]_ , \new_[87748]_ ,
    \new_[87749]_ , \new_[87752]_ , \new_[87755]_ , \new_[87756]_ ,
    \new_[87757]_ , \new_[87760]_ , \new_[87763]_ , \new_[87764]_ ,
    \new_[87767]_ , \new_[87770]_ , \new_[87771]_ , \new_[87772]_ ,
    \new_[87776]_ , \new_[87777]_ , \new_[87780]_ , \new_[87783]_ ,
    \new_[87784]_ , \new_[87785]_ , \new_[87788]_ , \new_[87791]_ ,
    \new_[87792]_ , \new_[87795]_ , \new_[87798]_ , \new_[87799]_ ,
    \new_[87800]_ , \new_[87804]_ , \new_[87805]_ , \new_[87808]_ ,
    \new_[87811]_ , \new_[87812]_ , \new_[87813]_ , \new_[87816]_ ,
    \new_[87819]_ , \new_[87820]_ , \new_[87823]_ , \new_[87826]_ ,
    \new_[87827]_ , \new_[87828]_ , \new_[87832]_ , \new_[87833]_ ,
    \new_[87836]_ , \new_[87839]_ , \new_[87840]_ , \new_[87841]_ ,
    \new_[87844]_ , \new_[87847]_ , \new_[87848]_ , \new_[87851]_ ,
    \new_[87854]_ , \new_[87855]_ , \new_[87856]_ , \new_[87860]_ ,
    \new_[87861]_ , \new_[87864]_ , \new_[87867]_ , \new_[87868]_ ,
    \new_[87869]_ , \new_[87872]_ , \new_[87875]_ , \new_[87876]_ ,
    \new_[87879]_ , \new_[87882]_ , \new_[87883]_ , \new_[87884]_ ,
    \new_[87888]_ , \new_[87889]_ , \new_[87892]_ , \new_[87895]_ ,
    \new_[87896]_ , \new_[87897]_ , \new_[87900]_ , \new_[87903]_ ,
    \new_[87904]_ , \new_[87907]_ , \new_[87910]_ , \new_[87911]_ ,
    \new_[87912]_ , \new_[87916]_ , \new_[87917]_ , \new_[87920]_ ,
    \new_[87923]_ , \new_[87924]_ , \new_[87925]_ , \new_[87928]_ ,
    \new_[87931]_ , \new_[87932]_ , \new_[87935]_ , \new_[87938]_ ,
    \new_[87939]_ , \new_[87940]_ , \new_[87944]_ , \new_[87945]_ ,
    \new_[87948]_ , \new_[87951]_ , \new_[87952]_ , \new_[87953]_ ,
    \new_[87956]_ , \new_[87959]_ , \new_[87960]_ , \new_[87963]_ ,
    \new_[87966]_ , \new_[87967]_ , \new_[87968]_ , \new_[87972]_ ,
    \new_[87973]_ , \new_[87976]_ , \new_[87979]_ , \new_[87980]_ ,
    \new_[87981]_ , \new_[87984]_ , \new_[87987]_ , \new_[87988]_ ,
    \new_[87991]_ , \new_[87994]_ , \new_[87995]_ , \new_[87996]_ ,
    \new_[88000]_ , \new_[88001]_ , \new_[88004]_ , \new_[88007]_ ,
    \new_[88008]_ , \new_[88009]_ , \new_[88012]_ , \new_[88015]_ ,
    \new_[88016]_ , \new_[88019]_ , \new_[88022]_ , \new_[88023]_ ,
    \new_[88024]_ , \new_[88028]_ , \new_[88029]_ , \new_[88032]_ ,
    \new_[88035]_ , \new_[88036]_ , \new_[88037]_ , \new_[88040]_ ,
    \new_[88043]_ , \new_[88044]_ , \new_[88047]_ , \new_[88050]_ ,
    \new_[88051]_ , \new_[88052]_ , \new_[88056]_ , \new_[88057]_ ,
    \new_[88060]_ , \new_[88063]_ , \new_[88064]_ , \new_[88065]_ ,
    \new_[88068]_ , \new_[88071]_ , \new_[88072]_ , \new_[88075]_ ,
    \new_[88078]_ , \new_[88079]_ , \new_[88080]_ , \new_[88084]_ ,
    \new_[88085]_ , \new_[88088]_ , \new_[88091]_ , \new_[88092]_ ,
    \new_[88093]_ , \new_[88096]_ , \new_[88099]_ , \new_[88100]_ ,
    \new_[88103]_ , \new_[88106]_ , \new_[88107]_ , \new_[88108]_ ,
    \new_[88112]_ , \new_[88113]_ , \new_[88116]_ , \new_[88119]_ ,
    \new_[88120]_ , \new_[88121]_ , \new_[88124]_ , \new_[88127]_ ,
    \new_[88128]_ , \new_[88131]_ , \new_[88134]_ , \new_[88135]_ ,
    \new_[88136]_ , \new_[88140]_ , \new_[88141]_ , \new_[88144]_ ,
    \new_[88147]_ , \new_[88148]_ , \new_[88149]_ , \new_[88152]_ ,
    \new_[88155]_ , \new_[88156]_ , \new_[88159]_ , \new_[88162]_ ,
    \new_[88163]_ , \new_[88164]_ , \new_[88168]_ , \new_[88169]_ ,
    \new_[88172]_ , \new_[88175]_ , \new_[88176]_ , \new_[88177]_ ,
    \new_[88180]_ , \new_[88183]_ , \new_[88184]_ , \new_[88187]_ ,
    \new_[88190]_ , \new_[88191]_ , \new_[88192]_ , \new_[88196]_ ,
    \new_[88197]_ , \new_[88200]_ , \new_[88203]_ , \new_[88204]_ ,
    \new_[88205]_ , \new_[88208]_ , \new_[88211]_ , \new_[88212]_ ,
    \new_[88215]_ , \new_[88218]_ , \new_[88219]_ , \new_[88220]_ ,
    \new_[88224]_ , \new_[88225]_ , \new_[88228]_ , \new_[88231]_ ,
    \new_[88232]_ , \new_[88233]_ , \new_[88236]_ , \new_[88239]_ ,
    \new_[88240]_ , \new_[88243]_ , \new_[88246]_ , \new_[88247]_ ,
    \new_[88248]_ , \new_[88252]_ , \new_[88253]_ , \new_[88256]_ ,
    \new_[88259]_ , \new_[88260]_ , \new_[88261]_ , \new_[88264]_ ,
    \new_[88267]_ , \new_[88268]_ , \new_[88271]_ , \new_[88274]_ ,
    \new_[88275]_ , \new_[88276]_ , \new_[88280]_ , \new_[88281]_ ,
    \new_[88284]_ , \new_[88287]_ , \new_[88288]_ , \new_[88289]_ ,
    \new_[88292]_ , \new_[88295]_ , \new_[88296]_ , \new_[88299]_ ,
    \new_[88302]_ , \new_[88303]_ , \new_[88304]_ , \new_[88308]_ ,
    \new_[88309]_ , \new_[88312]_ , \new_[88315]_ , \new_[88316]_ ,
    \new_[88317]_ , \new_[88320]_ , \new_[88323]_ , \new_[88324]_ ,
    \new_[88327]_ , \new_[88330]_ , \new_[88331]_ , \new_[88332]_ ,
    \new_[88336]_ , \new_[88337]_ , \new_[88340]_ , \new_[88343]_ ,
    \new_[88344]_ , \new_[88345]_ , \new_[88348]_ , \new_[88351]_ ,
    \new_[88352]_ , \new_[88355]_ , \new_[88358]_ , \new_[88359]_ ,
    \new_[88360]_ , \new_[88364]_ , \new_[88365]_ , \new_[88368]_ ,
    \new_[88371]_ , \new_[88372]_ , \new_[88373]_ , \new_[88376]_ ,
    \new_[88379]_ , \new_[88380]_ , \new_[88383]_ , \new_[88386]_ ,
    \new_[88387]_ , \new_[88388]_ , \new_[88392]_ , \new_[88393]_ ,
    \new_[88396]_ , \new_[88399]_ , \new_[88400]_ , \new_[88401]_ ,
    \new_[88404]_ , \new_[88407]_ , \new_[88408]_ , \new_[88411]_ ,
    \new_[88414]_ , \new_[88415]_ , \new_[88416]_ , \new_[88420]_ ,
    \new_[88421]_ , \new_[88424]_ , \new_[88427]_ , \new_[88428]_ ,
    \new_[88429]_ , \new_[88432]_ , \new_[88435]_ , \new_[88436]_ ,
    \new_[88439]_ , \new_[88442]_ , \new_[88443]_ , \new_[88444]_ ,
    \new_[88448]_ , \new_[88449]_ , \new_[88452]_ , \new_[88455]_ ,
    \new_[88456]_ , \new_[88457]_ , \new_[88460]_ , \new_[88463]_ ,
    \new_[88464]_ , \new_[88467]_ , \new_[88470]_ , \new_[88471]_ ,
    \new_[88472]_ , \new_[88476]_ , \new_[88477]_ , \new_[88480]_ ,
    \new_[88483]_ , \new_[88484]_ , \new_[88485]_ , \new_[88488]_ ,
    \new_[88491]_ , \new_[88492]_ , \new_[88495]_ , \new_[88498]_ ,
    \new_[88499]_ , \new_[88500]_ , \new_[88504]_ , \new_[88505]_ ,
    \new_[88508]_ , \new_[88511]_ , \new_[88512]_ , \new_[88513]_ ,
    \new_[88516]_ , \new_[88519]_ , \new_[88520]_ , \new_[88523]_ ,
    \new_[88526]_ , \new_[88527]_ , \new_[88528]_ , \new_[88532]_ ,
    \new_[88533]_ , \new_[88536]_ , \new_[88539]_ , \new_[88540]_ ,
    \new_[88541]_ , \new_[88544]_ , \new_[88547]_ , \new_[88548]_ ,
    \new_[88551]_ , \new_[88554]_ , \new_[88555]_ , \new_[88556]_ ,
    \new_[88560]_ , \new_[88561]_ , \new_[88564]_ , \new_[88567]_ ,
    \new_[88568]_ , \new_[88569]_ , \new_[88572]_ , \new_[88575]_ ,
    \new_[88576]_ , \new_[88579]_ , \new_[88582]_ , \new_[88583]_ ,
    \new_[88584]_ , \new_[88588]_ , \new_[88589]_ , \new_[88592]_ ,
    \new_[88595]_ , \new_[88596]_ , \new_[88597]_ , \new_[88600]_ ,
    \new_[88603]_ , \new_[88604]_ , \new_[88607]_ , \new_[88610]_ ,
    \new_[88611]_ , \new_[88612]_ , \new_[88616]_ , \new_[88617]_ ,
    \new_[88620]_ , \new_[88623]_ , \new_[88624]_ , \new_[88625]_ ,
    \new_[88628]_ , \new_[88631]_ , \new_[88632]_ , \new_[88635]_ ,
    \new_[88638]_ , \new_[88639]_ , \new_[88640]_ , \new_[88644]_ ,
    \new_[88645]_ , \new_[88648]_ , \new_[88651]_ , \new_[88652]_ ,
    \new_[88653]_ , \new_[88656]_ , \new_[88659]_ , \new_[88660]_ ,
    \new_[88663]_ , \new_[88666]_ , \new_[88667]_ , \new_[88668]_ ,
    \new_[88672]_ , \new_[88673]_ , \new_[88676]_ , \new_[88679]_ ,
    \new_[88680]_ , \new_[88681]_ , \new_[88684]_ , \new_[88687]_ ,
    \new_[88688]_ , \new_[88691]_ , \new_[88694]_ , \new_[88695]_ ,
    \new_[88696]_ , \new_[88700]_ , \new_[88701]_ , \new_[88704]_ ,
    \new_[88707]_ , \new_[88708]_ , \new_[88709]_ , \new_[88712]_ ,
    \new_[88715]_ , \new_[88716]_ , \new_[88719]_ , \new_[88722]_ ,
    \new_[88723]_ , \new_[88724]_ , \new_[88728]_ , \new_[88729]_ ,
    \new_[88732]_ , \new_[88735]_ , \new_[88736]_ , \new_[88737]_ ,
    \new_[88740]_ , \new_[88743]_ , \new_[88744]_ , \new_[88747]_ ,
    \new_[88750]_ , \new_[88751]_ , \new_[88752]_ , \new_[88756]_ ,
    \new_[88757]_ , \new_[88760]_ , \new_[88763]_ , \new_[88764]_ ,
    \new_[88765]_ , \new_[88768]_ , \new_[88771]_ , \new_[88772]_ ,
    \new_[88775]_ , \new_[88778]_ , \new_[88779]_ , \new_[88780]_ ,
    \new_[88784]_ , \new_[88785]_ , \new_[88788]_ , \new_[88791]_ ,
    \new_[88792]_ , \new_[88793]_ , \new_[88796]_ , \new_[88799]_ ,
    \new_[88800]_ , \new_[88803]_ , \new_[88806]_ , \new_[88807]_ ,
    \new_[88808]_ , \new_[88812]_ , \new_[88813]_ , \new_[88816]_ ,
    \new_[88819]_ , \new_[88820]_ , \new_[88821]_ , \new_[88824]_ ,
    \new_[88827]_ , \new_[88828]_ , \new_[88831]_ , \new_[88834]_ ,
    \new_[88835]_ , \new_[88836]_ , \new_[88840]_ , \new_[88841]_ ,
    \new_[88844]_ , \new_[88847]_ , \new_[88848]_ , \new_[88849]_ ,
    \new_[88852]_ , \new_[88855]_ , \new_[88856]_ , \new_[88859]_ ,
    \new_[88862]_ , \new_[88863]_ , \new_[88864]_ , \new_[88868]_ ,
    \new_[88869]_ , \new_[88872]_ , \new_[88875]_ , \new_[88876]_ ,
    \new_[88877]_ , \new_[88880]_ , \new_[88883]_ , \new_[88884]_ ,
    \new_[88887]_ , \new_[88890]_ , \new_[88891]_ , \new_[88892]_ ,
    \new_[88896]_ , \new_[88897]_ , \new_[88900]_ , \new_[88903]_ ,
    \new_[88904]_ , \new_[88905]_ , \new_[88908]_ , \new_[88911]_ ,
    \new_[88912]_ , \new_[88915]_ , \new_[88918]_ , \new_[88919]_ ,
    \new_[88920]_ , \new_[88924]_ , \new_[88925]_ , \new_[88928]_ ,
    \new_[88931]_ , \new_[88932]_ , \new_[88933]_ , \new_[88936]_ ,
    \new_[88939]_ , \new_[88940]_ , \new_[88943]_ , \new_[88946]_ ,
    \new_[88947]_ , \new_[88948]_ , \new_[88952]_ , \new_[88953]_ ,
    \new_[88956]_ , \new_[88959]_ , \new_[88960]_ , \new_[88961]_ ,
    \new_[88964]_ , \new_[88967]_ , \new_[88968]_ , \new_[88971]_ ,
    \new_[88974]_ , \new_[88975]_ , \new_[88976]_ , \new_[88980]_ ,
    \new_[88981]_ , \new_[88984]_ , \new_[88987]_ , \new_[88988]_ ,
    \new_[88989]_ , \new_[88992]_ , \new_[88995]_ , \new_[88996]_ ,
    \new_[88999]_ , \new_[89002]_ , \new_[89003]_ , \new_[89004]_ ,
    \new_[89008]_ , \new_[89009]_ , \new_[89012]_ , \new_[89015]_ ,
    \new_[89016]_ , \new_[89017]_ , \new_[89020]_ , \new_[89023]_ ,
    \new_[89024]_ , \new_[89027]_ , \new_[89030]_ , \new_[89031]_ ,
    \new_[89032]_ , \new_[89036]_ , \new_[89037]_ , \new_[89040]_ ,
    \new_[89043]_ , \new_[89044]_ , \new_[89045]_ , \new_[89048]_ ,
    \new_[89051]_ , \new_[89052]_ , \new_[89055]_ , \new_[89058]_ ,
    \new_[89059]_ , \new_[89060]_ , \new_[89064]_ , \new_[89065]_ ,
    \new_[89068]_ , \new_[89071]_ , \new_[89072]_ , \new_[89073]_ ,
    \new_[89076]_ , \new_[89079]_ , \new_[89080]_ , \new_[89083]_ ,
    \new_[89086]_ , \new_[89087]_ , \new_[89088]_ , \new_[89092]_ ,
    \new_[89093]_ , \new_[89096]_ , \new_[89099]_ , \new_[89100]_ ,
    \new_[89101]_ , \new_[89104]_ , \new_[89107]_ , \new_[89108]_ ,
    \new_[89111]_ , \new_[89114]_ , \new_[89115]_ , \new_[89116]_ ,
    \new_[89120]_ , \new_[89121]_ , \new_[89124]_ , \new_[89127]_ ,
    \new_[89128]_ , \new_[89129]_ , \new_[89132]_ , \new_[89135]_ ,
    \new_[89136]_ , \new_[89139]_ , \new_[89142]_ , \new_[89143]_ ,
    \new_[89144]_ , \new_[89148]_ , \new_[89149]_ , \new_[89152]_ ,
    \new_[89155]_ , \new_[89156]_ , \new_[89157]_ , \new_[89160]_ ,
    \new_[89163]_ , \new_[89164]_ , \new_[89167]_ , \new_[89170]_ ,
    \new_[89171]_ , \new_[89172]_ , \new_[89176]_ , \new_[89177]_ ,
    \new_[89180]_ , \new_[89183]_ , \new_[89184]_ , \new_[89185]_ ,
    \new_[89188]_ , \new_[89191]_ , \new_[89192]_ , \new_[89195]_ ,
    \new_[89198]_ , \new_[89199]_ , \new_[89200]_ , \new_[89204]_ ,
    \new_[89205]_ , \new_[89208]_ , \new_[89211]_ , \new_[89212]_ ,
    \new_[89213]_ , \new_[89216]_ , \new_[89219]_ , \new_[89220]_ ,
    \new_[89223]_ , \new_[89226]_ , \new_[89227]_ , \new_[89228]_ ,
    \new_[89232]_ , \new_[89233]_ , \new_[89236]_ , \new_[89239]_ ,
    \new_[89240]_ , \new_[89241]_ , \new_[89244]_ , \new_[89247]_ ,
    \new_[89248]_ , \new_[89251]_ , \new_[89254]_ , \new_[89255]_ ,
    \new_[89256]_ , \new_[89260]_ , \new_[89261]_ , \new_[89264]_ ,
    \new_[89267]_ , \new_[89268]_ , \new_[89269]_ , \new_[89272]_ ,
    \new_[89275]_ , \new_[89276]_ , \new_[89279]_ , \new_[89282]_ ,
    \new_[89283]_ , \new_[89284]_ , \new_[89288]_ , \new_[89289]_ ,
    \new_[89292]_ , \new_[89295]_ , \new_[89296]_ , \new_[89297]_ ,
    \new_[89300]_ , \new_[89303]_ , \new_[89304]_ , \new_[89307]_ ,
    \new_[89310]_ , \new_[89311]_ , \new_[89312]_ , \new_[89316]_ ,
    \new_[89317]_ , \new_[89320]_ , \new_[89323]_ , \new_[89324]_ ,
    \new_[89325]_ , \new_[89328]_ , \new_[89331]_ , \new_[89332]_ ,
    \new_[89335]_ , \new_[89338]_ , \new_[89339]_ , \new_[89340]_ ,
    \new_[89344]_ , \new_[89345]_ , \new_[89348]_ , \new_[89351]_ ,
    \new_[89352]_ , \new_[89353]_ , \new_[89356]_ , \new_[89359]_ ,
    \new_[89360]_ , \new_[89363]_ , \new_[89366]_ , \new_[89367]_ ,
    \new_[89368]_ , \new_[89372]_ , \new_[89373]_ , \new_[89376]_ ,
    \new_[89379]_ , \new_[89380]_ , \new_[89381]_ , \new_[89384]_ ,
    \new_[89387]_ , \new_[89388]_ , \new_[89391]_ , \new_[89394]_ ,
    \new_[89395]_ , \new_[89396]_ , \new_[89400]_ , \new_[89401]_ ,
    \new_[89404]_ , \new_[89407]_ , \new_[89408]_ , \new_[89409]_ ,
    \new_[89412]_ , \new_[89415]_ , \new_[89416]_ , \new_[89419]_ ,
    \new_[89422]_ , \new_[89423]_ , \new_[89424]_ , \new_[89428]_ ,
    \new_[89429]_ , \new_[89432]_ , \new_[89435]_ , \new_[89436]_ ,
    \new_[89437]_ , \new_[89440]_ , \new_[89443]_ , \new_[89444]_ ,
    \new_[89447]_ , \new_[89450]_ , \new_[89451]_ , \new_[89452]_ ,
    \new_[89456]_ , \new_[89457]_ , \new_[89460]_ , \new_[89463]_ ,
    \new_[89464]_ , \new_[89465]_ , \new_[89468]_ , \new_[89471]_ ,
    \new_[89472]_ , \new_[89475]_ , \new_[89478]_ , \new_[89479]_ ,
    \new_[89480]_ , \new_[89484]_ , \new_[89485]_ , \new_[89488]_ ,
    \new_[89491]_ , \new_[89492]_ , \new_[89493]_ , \new_[89496]_ ,
    \new_[89499]_ , \new_[89500]_ , \new_[89503]_ , \new_[89506]_ ,
    \new_[89507]_ , \new_[89508]_ , \new_[89512]_ , \new_[89513]_ ,
    \new_[89516]_ , \new_[89519]_ , \new_[89520]_ , \new_[89521]_ ,
    \new_[89524]_ , \new_[89527]_ , \new_[89528]_ , \new_[89531]_ ,
    \new_[89534]_ , \new_[89535]_ , \new_[89536]_ , \new_[89540]_ ,
    \new_[89541]_ , \new_[89544]_ , \new_[89547]_ , \new_[89548]_ ,
    \new_[89549]_ , \new_[89552]_ , \new_[89555]_ , \new_[89556]_ ,
    \new_[89559]_ , \new_[89562]_ , \new_[89563]_ , \new_[89564]_ ,
    \new_[89568]_ , \new_[89569]_ , \new_[89572]_ , \new_[89575]_ ,
    \new_[89576]_ , \new_[89577]_ , \new_[89580]_ , \new_[89583]_ ,
    \new_[89584]_ , \new_[89587]_ , \new_[89590]_ , \new_[89591]_ ,
    \new_[89592]_ , \new_[89596]_ , \new_[89597]_ , \new_[89600]_ ,
    \new_[89603]_ , \new_[89604]_ , \new_[89605]_ , \new_[89608]_ ,
    \new_[89611]_ , \new_[89612]_ , \new_[89615]_ , \new_[89618]_ ,
    \new_[89619]_ , \new_[89620]_ , \new_[89624]_ , \new_[89625]_ ,
    \new_[89628]_ , \new_[89631]_ , \new_[89632]_ , \new_[89633]_ ,
    \new_[89636]_ , \new_[89639]_ , \new_[89640]_ , \new_[89643]_ ,
    \new_[89646]_ , \new_[89647]_ , \new_[89648]_ , \new_[89652]_ ,
    \new_[89653]_ , \new_[89656]_ , \new_[89659]_ , \new_[89660]_ ,
    \new_[89661]_ , \new_[89664]_ , \new_[89667]_ , \new_[89668]_ ,
    \new_[89671]_ , \new_[89674]_ , \new_[89675]_ , \new_[89676]_ ,
    \new_[89680]_ , \new_[89681]_ , \new_[89684]_ , \new_[89687]_ ,
    \new_[89688]_ , \new_[89689]_ , \new_[89692]_ , \new_[89695]_ ,
    \new_[89696]_ , \new_[89699]_ , \new_[89702]_ , \new_[89703]_ ,
    \new_[89704]_ , \new_[89708]_ , \new_[89709]_ , \new_[89712]_ ,
    \new_[89715]_ , \new_[89716]_ , \new_[89717]_ , \new_[89720]_ ,
    \new_[89723]_ , \new_[89724]_ , \new_[89727]_ , \new_[89730]_ ,
    \new_[89731]_ , \new_[89732]_ , \new_[89736]_ , \new_[89737]_ ,
    \new_[89740]_ , \new_[89743]_ , \new_[89744]_ , \new_[89745]_ ,
    \new_[89748]_ , \new_[89751]_ , \new_[89752]_ , \new_[89755]_ ,
    \new_[89758]_ , \new_[89759]_ , \new_[89760]_ , \new_[89764]_ ,
    \new_[89765]_ , \new_[89768]_ , \new_[89771]_ , \new_[89772]_ ,
    \new_[89773]_ , \new_[89776]_ , \new_[89779]_ , \new_[89780]_ ,
    \new_[89783]_ , \new_[89786]_ , \new_[89787]_ , \new_[89788]_ ,
    \new_[89792]_ , \new_[89793]_ , \new_[89796]_ , \new_[89799]_ ,
    \new_[89800]_ , \new_[89801]_ , \new_[89804]_ , \new_[89807]_ ,
    \new_[89808]_ , \new_[89811]_ , \new_[89814]_ , \new_[89815]_ ,
    \new_[89816]_ , \new_[89820]_ , \new_[89821]_ , \new_[89824]_ ,
    \new_[89827]_ , \new_[89828]_ , \new_[89829]_ , \new_[89832]_ ,
    \new_[89835]_ , \new_[89836]_ , \new_[89839]_ , \new_[89842]_ ,
    \new_[89843]_ , \new_[89844]_ , \new_[89848]_ , \new_[89849]_ ,
    \new_[89852]_ , \new_[89855]_ , \new_[89856]_ , \new_[89857]_ ,
    \new_[89860]_ , \new_[89863]_ , \new_[89864]_ , \new_[89867]_ ,
    \new_[89870]_ , \new_[89871]_ , \new_[89872]_ , \new_[89876]_ ,
    \new_[89877]_ , \new_[89880]_ , \new_[89883]_ , \new_[89884]_ ,
    \new_[89885]_ , \new_[89888]_ , \new_[89891]_ , \new_[89892]_ ,
    \new_[89895]_ , \new_[89898]_ , \new_[89899]_ , \new_[89900]_ ,
    \new_[89904]_ , \new_[89905]_ , \new_[89908]_ , \new_[89911]_ ,
    \new_[89912]_ , \new_[89913]_ , \new_[89916]_ , \new_[89919]_ ,
    \new_[89920]_ , \new_[89923]_ , \new_[89926]_ , \new_[89927]_ ,
    \new_[89928]_ , \new_[89932]_ , \new_[89933]_ , \new_[89936]_ ,
    \new_[89939]_ , \new_[89940]_ , \new_[89941]_ , \new_[89944]_ ,
    \new_[89947]_ , \new_[89948]_ , \new_[89951]_ , \new_[89954]_ ,
    \new_[89955]_ , \new_[89956]_ , \new_[89960]_ , \new_[89961]_ ,
    \new_[89964]_ , \new_[89967]_ , \new_[89968]_ , \new_[89969]_ ,
    \new_[89972]_ , \new_[89975]_ , \new_[89976]_ , \new_[89979]_ ,
    \new_[89982]_ , \new_[89983]_ , \new_[89984]_ , \new_[89988]_ ,
    \new_[89989]_ , \new_[89992]_ , \new_[89995]_ , \new_[89996]_ ,
    \new_[89997]_ , \new_[90000]_ , \new_[90003]_ , \new_[90004]_ ,
    \new_[90007]_ , \new_[90010]_ , \new_[90011]_ , \new_[90012]_ ,
    \new_[90016]_ , \new_[90017]_ , \new_[90020]_ , \new_[90023]_ ,
    \new_[90024]_ , \new_[90025]_ , \new_[90028]_ , \new_[90031]_ ,
    \new_[90032]_ , \new_[90035]_ , \new_[90038]_ , \new_[90039]_ ,
    \new_[90040]_ , \new_[90044]_ , \new_[90045]_ , \new_[90048]_ ,
    \new_[90051]_ , \new_[90052]_ , \new_[90053]_ , \new_[90056]_ ,
    \new_[90059]_ , \new_[90060]_ , \new_[90063]_ , \new_[90066]_ ,
    \new_[90067]_ , \new_[90068]_ , \new_[90072]_ , \new_[90073]_ ,
    \new_[90076]_ , \new_[90079]_ , \new_[90080]_ , \new_[90081]_ ,
    \new_[90084]_ , \new_[90087]_ , \new_[90088]_ , \new_[90091]_ ,
    \new_[90094]_ , \new_[90095]_ , \new_[90096]_ , \new_[90100]_ ,
    \new_[90101]_ , \new_[90104]_ , \new_[90107]_ , \new_[90108]_ ,
    \new_[90109]_ , \new_[90112]_ , \new_[90115]_ , \new_[90116]_ ,
    \new_[90119]_ , \new_[90122]_ , \new_[90123]_ , \new_[90124]_ ,
    \new_[90128]_ , \new_[90129]_ , \new_[90132]_ , \new_[90135]_ ,
    \new_[90136]_ , \new_[90137]_ , \new_[90140]_ , \new_[90143]_ ,
    \new_[90144]_ , \new_[90147]_ , \new_[90150]_ , \new_[90151]_ ,
    \new_[90152]_ , \new_[90156]_ , \new_[90157]_ , \new_[90160]_ ,
    \new_[90163]_ , \new_[90164]_ , \new_[90165]_ , \new_[90168]_ ,
    \new_[90171]_ , \new_[90172]_ , \new_[90175]_ , \new_[90178]_ ,
    \new_[90179]_ , \new_[90180]_ , \new_[90184]_ , \new_[90185]_ ,
    \new_[90188]_ , \new_[90191]_ , \new_[90192]_ , \new_[90193]_ ,
    \new_[90196]_ , \new_[90199]_ , \new_[90200]_ , \new_[90203]_ ,
    \new_[90206]_ , \new_[90207]_ , \new_[90208]_ , \new_[90212]_ ,
    \new_[90213]_ , \new_[90216]_ , \new_[90219]_ , \new_[90220]_ ,
    \new_[90221]_ , \new_[90224]_ , \new_[90227]_ , \new_[90228]_ ,
    \new_[90231]_ , \new_[90234]_ , \new_[90235]_ , \new_[90236]_ ,
    \new_[90240]_ , \new_[90241]_ , \new_[90244]_ , \new_[90247]_ ,
    \new_[90248]_ , \new_[90249]_ , \new_[90252]_ , \new_[90255]_ ,
    \new_[90256]_ , \new_[90259]_ , \new_[90262]_ , \new_[90263]_ ,
    \new_[90264]_ , \new_[90268]_ , \new_[90269]_ , \new_[90272]_ ,
    \new_[90275]_ , \new_[90276]_ , \new_[90277]_ , \new_[90280]_ ,
    \new_[90283]_ , \new_[90284]_ , \new_[90287]_ , \new_[90290]_ ,
    \new_[90291]_ , \new_[90292]_ , \new_[90296]_ , \new_[90297]_ ,
    \new_[90300]_ , \new_[90303]_ , \new_[90304]_ , \new_[90305]_ ,
    \new_[90308]_ , \new_[90311]_ , \new_[90312]_ , \new_[90315]_ ,
    \new_[90318]_ , \new_[90319]_ , \new_[90320]_ , \new_[90324]_ ,
    \new_[90325]_ , \new_[90328]_ , \new_[90331]_ , \new_[90332]_ ,
    \new_[90333]_ , \new_[90336]_ , \new_[90339]_ , \new_[90340]_ ,
    \new_[90343]_ , \new_[90346]_ , \new_[90347]_ , \new_[90348]_ ,
    \new_[90352]_ , \new_[90353]_ , \new_[90356]_ , \new_[90359]_ ,
    \new_[90360]_ , \new_[90361]_ , \new_[90364]_ , \new_[90367]_ ,
    \new_[90368]_ , \new_[90371]_ , \new_[90374]_ , \new_[90375]_ ,
    \new_[90376]_ , \new_[90380]_ , \new_[90381]_ , \new_[90384]_ ,
    \new_[90387]_ , \new_[90388]_ , \new_[90389]_ , \new_[90392]_ ,
    \new_[90395]_ , \new_[90396]_ , \new_[90399]_ , \new_[90402]_ ,
    \new_[90403]_ , \new_[90404]_ , \new_[90408]_ , \new_[90409]_ ,
    \new_[90412]_ , \new_[90415]_ , \new_[90416]_ , \new_[90417]_ ,
    \new_[90420]_ , \new_[90423]_ , \new_[90424]_ , \new_[90427]_ ,
    \new_[90430]_ , \new_[90431]_ , \new_[90432]_ , \new_[90436]_ ,
    \new_[90437]_ , \new_[90440]_ , \new_[90443]_ , \new_[90444]_ ,
    \new_[90445]_ , \new_[90448]_ , \new_[90451]_ , \new_[90452]_ ,
    \new_[90455]_ , \new_[90458]_ , \new_[90459]_ , \new_[90460]_ ,
    \new_[90464]_ , \new_[90465]_ , \new_[90468]_ , \new_[90471]_ ,
    \new_[90472]_ , \new_[90473]_ , \new_[90476]_ , \new_[90479]_ ,
    \new_[90480]_ , \new_[90483]_ , \new_[90486]_ , \new_[90487]_ ,
    \new_[90488]_ , \new_[90492]_ , \new_[90493]_ , \new_[90496]_ ,
    \new_[90499]_ , \new_[90500]_ , \new_[90501]_ , \new_[90504]_ ,
    \new_[90507]_ , \new_[90508]_ , \new_[90511]_ , \new_[90514]_ ,
    \new_[90515]_ , \new_[90516]_ , \new_[90520]_ , \new_[90521]_ ,
    \new_[90524]_ , \new_[90527]_ , \new_[90528]_ , \new_[90529]_ ,
    \new_[90532]_ , \new_[90535]_ , \new_[90536]_ , \new_[90539]_ ,
    \new_[90542]_ , \new_[90543]_ , \new_[90544]_ , \new_[90548]_ ,
    \new_[90549]_ , \new_[90552]_ , \new_[90555]_ , \new_[90556]_ ,
    \new_[90557]_ , \new_[90560]_ , \new_[90563]_ , \new_[90564]_ ,
    \new_[90567]_ , \new_[90570]_ , \new_[90571]_ , \new_[90572]_ ,
    \new_[90576]_ , \new_[90577]_ , \new_[90580]_ , \new_[90583]_ ,
    \new_[90584]_ , \new_[90585]_ , \new_[90588]_ , \new_[90591]_ ,
    \new_[90592]_ , \new_[90595]_ , \new_[90598]_ , \new_[90599]_ ,
    \new_[90600]_ , \new_[90604]_ , \new_[90605]_ , \new_[90608]_ ,
    \new_[90611]_ , \new_[90612]_ , \new_[90613]_ , \new_[90616]_ ,
    \new_[90619]_ , \new_[90620]_ , \new_[90623]_ , \new_[90626]_ ,
    \new_[90627]_ , \new_[90628]_ , \new_[90632]_ , \new_[90633]_ ,
    \new_[90636]_ , \new_[90639]_ , \new_[90640]_ , \new_[90641]_ ,
    \new_[90644]_ , \new_[90647]_ , \new_[90648]_ , \new_[90651]_ ,
    \new_[90654]_ , \new_[90655]_ , \new_[90656]_ , \new_[90660]_ ,
    \new_[90661]_ , \new_[90664]_ , \new_[90667]_ , \new_[90668]_ ,
    \new_[90669]_ , \new_[90672]_ , \new_[90675]_ , \new_[90676]_ ,
    \new_[90679]_ , \new_[90682]_ , \new_[90683]_ , \new_[90684]_ ,
    \new_[90688]_ , \new_[90689]_ , \new_[90692]_ , \new_[90695]_ ,
    \new_[90696]_ , \new_[90697]_ , \new_[90700]_ , \new_[90703]_ ,
    \new_[90704]_ , \new_[90707]_ , \new_[90710]_ , \new_[90711]_ ,
    \new_[90712]_ , \new_[90716]_ , \new_[90717]_ , \new_[90720]_ ,
    \new_[90723]_ , \new_[90724]_ , \new_[90725]_ , \new_[90728]_ ,
    \new_[90731]_ , \new_[90732]_ , \new_[90735]_ , \new_[90738]_ ,
    \new_[90739]_ , \new_[90740]_ , \new_[90744]_ , \new_[90745]_ ,
    \new_[90748]_ , \new_[90751]_ , \new_[90752]_ , \new_[90753]_ ,
    \new_[90756]_ , \new_[90759]_ , \new_[90760]_ , \new_[90763]_ ,
    \new_[90766]_ , \new_[90767]_ , \new_[90768]_ , \new_[90772]_ ,
    \new_[90773]_ , \new_[90776]_ , \new_[90779]_ , \new_[90780]_ ,
    \new_[90781]_ , \new_[90784]_ , \new_[90787]_ , \new_[90788]_ ,
    \new_[90791]_ , \new_[90794]_ , \new_[90795]_ , \new_[90796]_ ,
    \new_[90800]_ , \new_[90801]_ , \new_[90804]_ , \new_[90807]_ ,
    \new_[90808]_ , \new_[90809]_ , \new_[90812]_ , \new_[90815]_ ,
    \new_[90816]_ , \new_[90819]_ , \new_[90822]_ , \new_[90823]_ ,
    \new_[90824]_ , \new_[90828]_ , \new_[90829]_ , \new_[90832]_ ,
    \new_[90835]_ , \new_[90836]_ , \new_[90837]_ , \new_[90840]_ ,
    \new_[90843]_ , \new_[90844]_ , \new_[90847]_ , \new_[90850]_ ,
    \new_[90851]_ , \new_[90852]_ , \new_[90856]_ , \new_[90857]_ ,
    \new_[90860]_ , \new_[90863]_ , \new_[90864]_ , \new_[90865]_ ,
    \new_[90868]_ , \new_[90871]_ , \new_[90872]_ , \new_[90875]_ ,
    \new_[90878]_ , \new_[90879]_ , \new_[90880]_ , \new_[90884]_ ,
    \new_[90885]_ , \new_[90888]_ , \new_[90891]_ , \new_[90892]_ ,
    \new_[90893]_ , \new_[90896]_ , \new_[90899]_ , \new_[90900]_ ,
    \new_[90903]_ , \new_[90906]_ , \new_[90907]_ , \new_[90908]_ ,
    \new_[90912]_ , \new_[90913]_ , \new_[90916]_ , \new_[90919]_ ,
    \new_[90920]_ , \new_[90921]_ , \new_[90924]_ , \new_[90927]_ ,
    \new_[90928]_ , \new_[90931]_ , \new_[90934]_ , \new_[90935]_ ,
    \new_[90936]_ , \new_[90940]_ , \new_[90941]_ , \new_[90944]_ ,
    \new_[90947]_ , \new_[90948]_ , \new_[90949]_ , \new_[90952]_ ,
    \new_[90955]_ , \new_[90956]_ , \new_[90959]_ , \new_[90962]_ ,
    \new_[90963]_ , \new_[90964]_ , \new_[90968]_ , \new_[90969]_ ,
    \new_[90972]_ , \new_[90975]_ , \new_[90976]_ , \new_[90977]_ ,
    \new_[90980]_ , \new_[90983]_ , \new_[90984]_ , \new_[90987]_ ,
    \new_[90990]_ , \new_[90991]_ , \new_[90992]_ , \new_[90996]_ ,
    \new_[90997]_ , \new_[91000]_ , \new_[91003]_ , \new_[91004]_ ,
    \new_[91005]_ , \new_[91008]_ , \new_[91011]_ , \new_[91012]_ ,
    \new_[91015]_ , \new_[91018]_ , \new_[91019]_ , \new_[91020]_ ,
    \new_[91024]_ , \new_[91025]_ , \new_[91028]_ , \new_[91031]_ ,
    \new_[91032]_ , \new_[91033]_ , \new_[91036]_ , \new_[91039]_ ,
    \new_[91040]_ , \new_[91043]_ , \new_[91046]_ , \new_[91047]_ ,
    \new_[91048]_ , \new_[91052]_ , \new_[91053]_ , \new_[91056]_ ,
    \new_[91059]_ , \new_[91060]_ , \new_[91061]_ , \new_[91064]_ ,
    \new_[91067]_ , \new_[91068]_ , \new_[91071]_ , \new_[91074]_ ,
    \new_[91075]_ , \new_[91076]_ , \new_[91080]_ , \new_[91081]_ ,
    \new_[91084]_ , \new_[91087]_ , \new_[91088]_ , \new_[91089]_ ,
    \new_[91092]_ , \new_[91095]_ , \new_[91096]_ , \new_[91099]_ ,
    \new_[91102]_ , \new_[91103]_ , \new_[91104]_ , \new_[91108]_ ,
    \new_[91109]_ , \new_[91112]_ , \new_[91115]_ , \new_[91116]_ ,
    \new_[91117]_ , \new_[91120]_ , \new_[91123]_ , \new_[91124]_ ,
    \new_[91127]_ , \new_[91130]_ , \new_[91131]_ , \new_[91132]_ ,
    \new_[91136]_ , \new_[91137]_ , \new_[91140]_ , \new_[91143]_ ,
    \new_[91144]_ , \new_[91145]_ , \new_[91148]_ , \new_[91151]_ ,
    \new_[91152]_ , \new_[91155]_ , \new_[91158]_ , \new_[91159]_ ,
    \new_[91160]_ , \new_[91164]_ , \new_[91165]_ , \new_[91168]_ ,
    \new_[91171]_ , \new_[91172]_ , \new_[91173]_ , \new_[91176]_ ,
    \new_[91179]_ , \new_[91180]_ , \new_[91183]_ , \new_[91186]_ ,
    \new_[91187]_ , \new_[91188]_ , \new_[91192]_ , \new_[91193]_ ,
    \new_[91196]_ , \new_[91199]_ , \new_[91200]_ , \new_[91201]_ ,
    \new_[91204]_ , \new_[91207]_ , \new_[91208]_ , \new_[91211]_ ,
    \new_[91214]_ , \new_[91215]_ , \new_[91216]_ , \new_[91220]_ ,
    \new_[91221]_ , \new_[91224]_ , \new_[91227]_ , \new_[91228]_ ,
    \new_[91229]_ , \new_[91232]_ , \new_[91235]_ , \new_[91236]_ ,
    \new_[91239]_ , \new_[91242]_ , \new_[91243]_ , \new_[91244]_ ,
    \new_[91248]_ , \new_[91249]_ , \new_[91252]_ , \new_[91255]_ ,
    \new_[91256]_ , \new_[91257]_ , \new_[91260]_ , \new_[91263]_ ,
    \new_[91264]_ , \new_[91267]_ , \new_[91270]_ , \new_[91271]_ ,
    \new_[91272]_ , \new_[91276]_ , \new_[91277]_ , \new_[91280]_ ,
    \new_[91283]_ , \new_[91284]_ , \new_[91285]_ , \new_[91288]_ ,
    \new_[91291]_ , \new_[91292]_ , \new_[91295]_ , \new_[91298]_ ,
    \new_[91299]_ , \new_[91300]_ , \new_[91304]_ , \new_[91305]_ ,
    \new_[91308]_ , \new_[91311]_ , \new_[91312]_ , \new_[91313]_ ,
    \new_[91316]_ , \new_[91319]_ , \new_[91320]_ , \new_[91323]_ ,
    \new_[91326]_ , \new_[91327]_ , \new_[91328]_ , \new_[91332]_ ,
    \new_[91333]_ , \new_[91336]_ , \new_[91339]_ , \new_[91340]_ ,
    \new_[91341]_ , \new_[91344]_ , \new_[91347]_ , \new_[91348]_ ,
    \new_[91351]_ , \new_[91354]_ , \new_[91355]_ , \new_[91356]_ ,
    \new_[91360]_ , \new_[91361]_ , \new_[91364]_ , \new_[91367]_ ,
    \new_[91368]_ , \new_[91369]_ , \new_[91372]_ , \new_[91375]_ ,
    \new_[91376]_ , \new_[91379]_ , \new_[91382]_ , \new_[91383]_ ,
    \new_[91384]_ , \new_[91388]_ , \new_[91389]_ , \new_[91392]_ ,
    \new_[91395]_ , \new_[91396]_ , \new_[91397]_ , \new_[91400]_ ,
    \new_[91403]_ , \new_[91404]_ , \new_[91407]_ , \new_[91410]_ ,
    \new_[91411]_ , \new_[91412]_ , \new_[91416]_ , \new_[91417]_ ,
    \new_[91420]_ , \new_[91423]_ , \new_[91424]_ , \new_[91425]_ ,
    \new_[91428]_ , \new_[91431]_ , \new_[91432]_ , \new_[91435]_ ,
    \new_[91438]_ , \new_[91439]_ , \new_[91440]_ , \new_[91444]_ ,
    \new_[91445]_ , \new_[91448]_ , \new_[91451]_ , \new_[91452]_ ,
    \new_[91453]_ , \new_[91456]_ , \new_[91459]_ , \new_[91460]_ ,
    \new_[91463]_ , \new_[91466]_ , \new_[91467]_ , \new_[91468]_ ,
    \new_[91472]_ , \new_[91473]_ , \new_[91476]_ , \new_[91479]_ ,
    \new_[91480]_ , \new_[91481]_ , \new_[91484]_ , \new_[91487]_ ,
    \new_[91488]_ , \new_[91491]_ , \new_[91494]_ , \new_[91495]_ ,
    \new_[91496]_ , \new_[91500]_ , \new_[91501]_ , \new_[91504]_ ,
    \new_[91507]_ , \new_[91508]_ , \new_[91509]_ , \new_[91512]_ ,
    \new_[91515]_ , \new_[91516]_ , \new_[91519]_ , \new_[91522]_ ,
    \new_[91523]_ , \new_[91524]_ , \new_[91528]_ , \new_[91529]_ ,
    \new_[91532]_ , \new_[91535]_ , \new_[91536]_ , \new_[91537]_ ,
    \new_[91540]_ , \new_[91543]_ , \new_[91544]_ , \new_[91547]_ ,
    \new_[91550]_ , \new_[91551]_ , \new_[91552]_ , \new_[91556]_ ,
    \new_[91557]_ , \new_[91560]_ , \new_[91563]_ , \new_[91564]_ ,
    \new_[91565]_ , \new_[91568]_ , \new_[91571]_ , \new_[91572]_ ,
    \new_[91575]_ , \new_[91578]_ , \new_[91579]_ , \new_[91580]_ ,
    \new_[91584]_ , \new_[91585]_ , \new_[91588]_ , \new_[91591]_ ,
    \new_[91592]_ , \new_[91593]_ , \new_[91596]_ , \new_[91599]_ ,
    \new_[91600]_ , \new_[91603]_ , \new_[91606]_ , \new_[91607]_ ,
    \new_[91608]_ , \new_[91612]_ , \new_[91613]_ , \new_[91616]_ ,
    \new_[91619]_ , \new_[91620]_ , \new_[91621]_ , \new_[91624]_ ,
    \new_[91627]_ , \new_[91628]_ , \new_[91631]_ , \new_[91634]_ ,
    \new_[91635]_ , \new_[91636]_ , \new_[91640]_ , \new_[91641]_ ,
    \new_[91644]_ , \new_[91647]_ , \new_[91648]_ , \new_[91649]_ ,
    \new_[91652]_ , \new_[91655]_ , \new_[91656]_ , \new_[91659]_ ,
    \new_[91662]_ , \new_[91663]_ , \new_[91664]_ , \new_[91668]_ ,
    \new_[91669]_ , \new_[91672]_ , \new_[91675]_ , \new_[91676]_ ,
    \new_[91677]_ , \new_[91680]_ , \new_[91683]_ , \new_[91684]_ ,
    \new_[91687]_ , \new_[91690]_ , \new_[91691]_ , \new_[91692]_ ,
    \new_[91696]_ , \new_[91697]_ , \new_[91700]_ , \new_[91703]_ ,
    \new_[91704]_ , \new_[91705]_ , \new_[91708]_ , \new_[91711]_ ,
    \new_[91712]_ , \new_[91715]_ , \new_[91718]_ , \new_[91719]_ ,
    \new_[91720]_ , \new_[91724]_ , \new_[91725]_ , \new_[91728]_ ,
    \new_[91731]_ , \new_[91732]_ , \new_[91733]_ , \new_[91736]_ ,
    \new_[91739]_ , \new_[91740]_ , \new_[91743]_ , \new_[91746]_ ,
    \new_[91747]_ , \new_[91748]_ , \new_[91752]_ , \new_[91753]_ ,
    \new_[91756]_ , \new_[91759]_ , \new_[91760]_ , \new_[91761]_ ,
    \new_[91764]_ , \new_[91767]_ , \new_[91768]_ , \new_[91771]_ ,
    \new_[91774]_ , \new_[91775]_ , \new_[91776]_ , \new_[91780]_ ,
    \new_[91781]_ , \new_[91784]_ , \new_[91787]_ , \new_[91788]_ ,
    \new_[91789]_ , \new_[91792]_ , \new_[91795]_ , \new_[91796]_ ,
    \new_[91799]_ , \new_[91802]_ , \new_[91803]_ , \new_[91804]_ ,
    \new_[91808]_ , \new_[91809]_ , \new_[91812]_ , \new_[91815]_ ,
    \new_[91816]_ , \new_[91817]_ , \new_[91820]_ , \new_[91823]_ ,
    \new_[91824]_ , \new_[91827]_ , \new_[91830]_ , \new_[91831]_ ,
    \new_[91832]_ , \new_[91836]_ , \new_[91837]_ , \new_[91840]_ ,
    \new_[91843]_ , \new_[91844]_ , \new_[91845]_ , \new_[91848]_ ,
    \new_[91851]_ , \new_[91852]_ , \new_[91855]_ , \new_[91858]_ ,
    \new_[91859]_ , \new_[91860]_ , \new_[91864]_ , \new_[91865]_ ,
    \new_[91868]_ , \new_[91871]_ , \new_[91872]_ , \new_[91873]_ ,
    \new_[91876]_ , \new_[91879]_ , \new_[91880]_ , \new_[91883]_ ,
    \new_[91886]_ , \new_[91887]_ , \new_[91888]_ , \new_[91892]_ ,
    \new_[91893]_ , \new_[91896]_ , \new_[91899]_ , \new_[91900]_ ,
    \new_[91901]_ , \new_[91904]_ , \new_[91907]_ , \new_[91908]_ ,
    \new_[91911]_ , \new_[91914]_ , \new_[91915]_ , \new_[91916]_ ,
    \new_[91920]_ , \new_[91921]_ , \new_[91924]_ , \new_[91927]_ ,
    \new_[91928]_ , \new_[91929]_ , \new_[91932]_ , \new_[91935]_ ,
    \new_[91936]_ , \new_[91939]_ , \new_[91942]_ , \new_[91943]_ ,
    \new_[91944]_ , \new_[91948]_ , \new_[91949]_ , \new_[91952]_ ,
    \new_[91955]_ , \new_[91956]_ , \new_[91957]_ , \new_[91960]_ ,
    \new_[91963]_ , \new_[91964]_ , \new_[91967]_ , \new_[91970]_ ,
    \new_[91971]_ , \new_[91972]_ , \new_[91976]_ , \new_[91977]_ ,
    \new_[91980]_ , \new_[91983]_ , \new_[91984]_ , \new_[91985]_ ,
    \new_[91988]_ , \new_[91991]_ , \new_[91992]_ , \new_[91995]_ ,
    \new_[91998]_ , \new_[91999]_ , \new_[92000]_ , \new_[92004]_ ,
    \new_[92005]_ , \new_[92008]_ , \new_[92011]_ , \new_[92012]_ ,
    \new_[92013]_ , \new_[92016]_ , \new_[92019]_ , \new_[92020]_ ,
    \new_[92023]_ , \new_[92026]_ , \new_[92027]_ , \new_[92028]_ ,
    \new_[92032]_ , \new_[92033]_ , \new_[92036]_ , \new_[92039]_ ,
    \new_[92040]_ , \new_[92041]_ , \new_[92044]_ , \new_[92047]_ ,
    \new_[92048]_ , \new_[92051]_ , \new_[92054]_ , \new_[92055]_ ,
    \new_[92056]_ , \new_[92060]_ , \new_[92061]_ , \new_[92064]_ ,
    \new_[92067]_ , \new_[92068]_ , \new_[92069]_ , \new_[92072]_ ,
    \new_[92075]_ , \new_[92076]_ , \new_[92079]_ , \new_[92082]_ ,
    \new_[92083]_ , \new_[92084]_ , \new_[92088]_ , \new_[92089]_ ,
    \new_[92092]_ , \new_[92095]_ , \new_[92096]_ , \new_[92097]_ ,
    \new_[92100]_ , \new_[92103]_ , \new_[92104]_ , \new_[92107]_ ,
    \new_[92110]_ , \new_[92111]_ , \new_[92112]_ , \new_[92116]_ ,
    \new_[92117]_ , \new_[92120]_ , \new_[92123]_ , \new_[92124]_ ,
    \new_[92125]_ , \new_[92128]_ , \new_[92131]_ , \new_[92132]_ ,
    \new_[92135]_ , \new_[92138]_ , \new_[92139]_ , \new_[92140]_ ,
    \new_[92144]_ , \new_[92145]_ , \new_[92148]_ , \new_[92151]_ ,
    \new_[92152]_ , \new_[92153]_ , \new_[92156]_ , \new_[92159]_ ,
    \new_[92160]_ , \new_[92163]_ , \new_[92166]_ , \new_[92167]_ ,
    \new_[92168]_ , \new_[92172]_ , \new_[92173]_ , \new_[92176]_ ,
    \new_[92179]_ , \new_[92180]_ , \new_[92181]_ , \new_[92184]_ ,
    \new_[92187]_ , \new_[92188]_ , \new_[92191]_ , \new_[92194]_ ,
    \new_[92195]_ , \new_[92196]_ , \new_[92200]_ , \new_[92201]_ ,
    \new_[92204]_ , \new_[92207]_ , \new_[92208]_ , \new_[92209]_ ,
    \new_[92212]_ , \new_[92215]_ , \new_[92216]_ , \new_[92219]_ ,
    \new_[92222]_ , \new_[92223]_ , \new_[92224]_ , \new_[92228]_ ,
    \new_[92229]_ , \new_[92232]_ , \new_[92235]_ , \new_[92236]_ ,
    \new_[92237]_ , \new_[92240]_ , \new_[92243]_ , \new_[92244]_ ,
    \new_[92247]_ , \new_[92250]_ , \new_[92251]_ , \new_[92252]_ ,
    \new_[92256]_ , \new_[92257]_ , \new_[92260]_ , \new_[92263]_ ,
    \new_[92264]_ , \new_[92265]_ , \new_[92268]_ , \new_[92271]_ ,
    \new_[92272]_ , \new_[92275]_ , \new_[92278]_ , \new_[92279]_ ,
    \new_[92280]_ , \new_[92284]_ , \new_[92285]_ , \new_[92288]_ ,
    \new_[92291]_ , \new_[92292]_ , \new_[92293]_ , \new_[92296]_ ,
    \new_[92299]_ , \new_[92300]_ , \new_[92303]_ , \new_[92306]_ ,
    \new_[92307]_ , \new_[92308]_ , \new_[92312]_ , \new_[92313]_ ,
    \new_[92316]_ , \new_[92319]_ , \new_[92320]_ , \new_[92321]_ ,
    \new_[92324]_ , \new_[92327]_ , \new_[92328]_ , \new_[92331]_ ,
    \new_[92334]_ , \new_[92335]_ , \new_[92336]_ , \new_[92340]_ ,
    \new_[92341]_ , \new_[92344]_ , \new_[92347]_ , \new_[92348]_ ,
    \new_[92349]_ , \new_[92352]_ , \new_[92355]_ , \new_[92356]_ ,
    \new_[92359]_ , \new_[92362]_ , \new_[92363]_ , \new_[92364]_ ,
    \new_[92368]_ , \new_[92369]_ , \new_[92372]_ , \new_[92375]_ ,
    \new_[92376]_ , \new_[92377]_ , \new_[92380]_ , \new_[92383]_ ,
    \new_[92384]_ , \new_[92387]_ , \new_[92390]_ , \new_[92391]_ ,
    \new_[92392]_ , \new_[92396]_ , \new_[92397]_ , \new_[92400]_ ,
    \new_[92403]_ , \new_[92404]_ , \new_[92405]_ , \new_[92408]_ ,
    \new_[92411]_ , \new_[92412]_ , \new_[92415]_ , \new_[92418]_ ,
    \new_[92419]_ , \new_[92420]_ , \new_[92424]_ , \new_[92425]_ ,
    \new_[92428]_ , \new_[92431]_ , \new_[92432]_ , \new_[92433]_ ,
    \new_[92436]_ , \new_[92439]_ , \new_[92440]_ , \new_[92443]_ ,
    \new_[92446]_ , \new_[92447]_ , \new_[92448]_ , \new_[92452]_ ,
    \new_[92453]_ , \new_[92456]_ , \new_[92459]_ , \new_[92460]_ ,
    \new_[92461]_ , \new_[92464]_ , \new_[92467]_ , \new_[92468]_ ,
    \new_[92471]_ , \new_[92474]_ , \new_[92475]_ , \new_[92476]_ ,
    \new_[92480]_ , \new_[92481]_ , \new_[92484]_ , \new_[92487]_ ,
    \new_[92488]_ , \new_[92489]_ , \new_[92492]_ , \new_[92495]_ ,
    \new_[92496]_ , \new_[92499]_ , \new_[92502]_ , \new_[92503]_ ,
    \new_[92504]_ , \new_[92508]_ , \new_[92509]_ , \new_[92512]_ ,
    \new_[92515]_ , \new_[92516]_ , \new_[92517]_ , \new_[92520]_ ,
    \new_[92523]_ , \new_[92524]_ , \new_[92527]_ , \new_[92530]_ ,
    \new_[92531]_ , \new_[92532]_ , \new_[92536]_ , \new_[92537]_ ,
    \new_[92540]_ , \new_[92543]_ , \new_[92544]_ , \new_[92545]_ ,
    \new_[92548]_ , \new_[92551]_ , \new_[92552]_ , \new_[92555]_ ,
    \new_[92558]_ , \new_[92559]_ , \new_[92560]_ , \new_[92564]_ ,
    \new_[92565]_ , \new_[92568]_ , \new_[92571]_ , \new_[92572]_ ,
    \new_[92573]_ , \new_[92576]_ , \new_[92579]_ , \new_[92580]_ ,
    \new_[92583]_ , \new_[92586]_ , \new_[92587]_ , \new_[92588]_ ,
    \new_[92592]_ , \new_[92593]_ , \new_[92596]_ , \new_[92599]_ ,
    \new_[92600]_ , \new_[92601]_ , \new_[92604]_ , \new_[92607]_ ,
    \new_[92608]_ , \new_[92611]_ , \new_[92614]_ , \new_[92615]_ ,
    \new_[92616]_ , \new_[92620]_ , \new_[92621]_ , \new_[92624]_ ,
    \new_[92627]_ , \new_[92628]_ , \new_[92629]_ , \new_[92632]_ ,
    \new_[92635]_ , \new_[92636]_ , \new_[92639]_ , \new_[92642]_ ,
    \new_[92643]_ , \new_[92644]_ , \new_[92648]_ , \new_[92649]_ ,
    \new_[92652]_ , \new_[92655]_ , \new_[92656]_ , \new_[92657]_ ,
    \new_[92660]_ , \new_[92663]_ , \new_[92664]_ , \new_[92667]_ ,
    \new_[92670]_ , \new_[92671]_ , \new_[92672]_ , \new_[92676]_ ,
    \new_[92677]_ , \new_[92680]_ , \new_[92683]_ , \new_[92684]_ ,
    \new_[92685]_ , \new_[92688]_ , \new_[92691]_ , \new_[92692]_ ,
    \new_[92695]_ , \new_[92698]_ , \new_[92699]_ , \new_[92700]_ ,
    \new_[92704]_ , \new_[92705]_ , \new_[92708]_ , \new_[92711]_ ,
    \new_[92712]_ , \new_[92713]_ , \new_[92716]_ , \new_[92719]_ ,
    \new_[92720]_ , \new_[92723]_ , \new_[92726]_ , \new_[92727]_ ,
    \new_[92728]_ , \new_[92732]_ , \new_[92733]_ , \new_[92736]_ ,
    \new_[92739]_ , \new_[92740]_ , \new_[92741]_ , \new_[92744]_ ,
    \new_[92747]_ , \new_[92748]_ , \new_[92751]_ , \new_[92754]_ ,
    \new_[92755]_ , \new_[92756]_ , \new_[92760]_ , \new_[92761]_ ,
    \new_[92764]_ , \new_[92767]_ , \new_[92768]_ , \new_[92769]_ ,
    \new_[92772]_ , \new_[92775]_ , \new_[92776]_ , \new_[92779]_ ,
    \new_[92782]_ , \new_[92783]_ , \new_[92784]_ , \new_[92788]_ ,
    \new_[92789]_ , \new_[92792]_ , \new_[92795]_ , \new_[92796]_ ,
    \new_[92797]_ , \new_[92800]_ , \new_[92803]_ , \new_[92804]_ ,
    \new_[92807]_ , \new_[92810]_ , \new_[92811]_ , \new_[92812]_ ,
    \new_[92816]_ , \new_[92817]_ , \new_[92820]_ , \new_[92823]_ ,
    \new_[92824]_ , \new_[92825]_ , \new_[92828]_ , \new_[92831]_ ,
    \new_[92832]_ , \new_[92835]_ , \new_[92838]_ , \new_[92839]_ ,
    \new_[92840]_ , \new_[92844]_ , \new_[92845]_ , \new_[92848]_ ,
    \new_[92851]_ , \new_[92852]_ , \new_[92853]_ , \new_[92856]_ ,
    \new_[92859]_ , \new_[92860]_ , \new_[92863]_ , \new_[92866]_ ,
    \new_[92867]_ , \new_[92868]_ , \new_[92871]_ , \new_[92874]_ ,
    \new_[92875]_ , \new_[92878]_ , \new_[92881]_ , \new_[92882]_ ,
    \new_[92883]_ , \new_[92886]_ , \new_[92889]_ , \new_[92890]_ ,
    \new_[92893]_ , \new_[92896]_ , \new_[92897]_ , \new_[92898]_ ,
    \new_[92901]_ , \new_[92904]_ , \new_[92905]_ , \new_[92908]_ ,
    \new_[92911]_ , \new_[92912]_ , \new_[92913]_ , \new_[92916]_ ,
    \new_[92919]_ , \new_[92920]_ , \new_[92923]_ , \new_[92926]_ ,
    \new_[92927]_ , \new_[92928]_ , \new_[92931]_ , \new_[92934]_ ,
    \new_[92935]_ , \new_[92938]_ , \new_[92941]_ , \new_[92942]_ ,
    \new_[92943]_ , \new_[92946]_ , \new_[92949]_ , \new_[92950]_ ,
    \new_[92953]_ , \new_[92956]_ , \new_[92957]_ , \new_[92958]_ ,
    \new_[92961]_ , \new_[92964]_ , \new_[92965]_ , \new_[92968]_ ,
    \new_[92971]_ , \new_[92972]_ , \new_[92973]_ , \new_[92976]_ ,
    \new_[92979]_ , \new_[92980]_ , \new_[92983]_ , \new_[92986]_ ,
    \new_[92987]_ , \new_[92988]_ , \new_[92991]_ , \new_[92994]_ ,
    \new_[92995]_ , \new_[92998]_ , \new_[93001]_ , \new_[93002]_ ,
    \new_[93003]_ , \new_[93006]_ , \new_[93009]_ , \new_[93010]_ ,
    \new_[93013]_ , \new_[93016]_ , \new_[93017]_ , \new_[93018]_ ,
    \new_[93021]_ , \new_[93024]_ , \new_[93025]_ , \new_[93028]_ ,
    \new_[93031]_ , \new_[93032]_ , \new_[93033]_ , \new_[93036]_ ,
    \new_[93039]_ , \new_[93040]_ , \new_[93043]_ , \new_[93046]_ ,
    \new_[93047]_ , \new_[93048]_ , \new_[93051]_ , \new_[93054]_ ,
    \new_[93055]_ , \new_[93058]_ , \new_[93061]_ , \new_[93062]_ ,
    \new_[93063]_ , \new_[93066]_ , \new_[93069]_ , \new_[93070]_ ,
    \new_[93073]_ , \new_[93076]_ , \new_[93077]_ , \new_[93078]_ ,
    \new_[93081]_ , \new_[93084]_ , \new_[93085]_ , \new_[93088]_ ,
    \new_[93091]_ , \new_[93092]_ , \new_[93093]_ , \new_[93096]_ ,
    \new_[93099]_ , \new_[93100]_ , \new_[93103]_ , \new_[93106]_ ,
    \new_[93107]_ , \new_[93108]_ , \new_[93111]_ , \new_[93114]_ ,
    \new_[93115]_ , \new_[93118]_ , \new_[93121]_ , \new_[93122]_ ,
    \new_[93123]_ , \new_[93126]_ , \new_[93129]_ , \new_[93130]_ ,
    \new_[93133]_ , \new_[93136]_ , \new_[93137]_ , \new_[93138]_ ,
    \new_[93141]_ , \new_[93144]_ , \new_[93145]_ , \new_[93148]_ ,
    \new_[93151]_ , \new_[93152]_ , \new_[93153]_ , \new_[93156]_ ,
    \new_[93159]_ , \new_[93160]_ , \new_[93163]_ , \new_[93166]_ ,
    \new_[93167]_ , \new_[93168]_ , \new_[93171]_ , \new_[93174]_ ,
    \new_[93175]_ , \new_[93178]_ , \new_[93181]_ , \new_[93182]_ ,
    \new_[93183]_ , \new_[93186]_ , \new_[93189]_ , \new_[93190]_ ,
    \new_[93193]_ , \new_[93196]_ , \new_[93197]_ , \new_[93198]_ ,
    \new_[93201]_ , \new_[93204]_ , \new_[93205]_ , \new_[93208]_ ,
    \new_[93211]_ , \new_[93212]_ , \new_[93213]_ , \new_[93216]_ ,
    \new_[93219]_ , \new_[93220]_ , \new_[93223]_ , \new_[93226]_ ,
    \new_[93227]_ , \new_[93228]_ , \new_[93231]_ , \new_[93234]_ ,
    \new_[93235]_ , \new_[93238]_ , \new_[93241]_ , \new_[93242]_ ,
    \new_[93243]_ , \new_[93246]_ , \new_[93249]_ , \new_[93250]_ ,
    \new_[93253]_ , \new_[93256]_ , \new_[93257]_ , \new_[93258]_ ,
    \new_[93261]_ , \new_[93264]_ , \new_[93265]_ , \new_[93268]_ ,
    \new_[93271]_ , \new_[93272]_ , \new_[93273]_ , \new_[93276]_ ,
    \new_[93279]_ , \new_[93280]_ , \new_[93283]_ , \new_[93286]_ ,
    \new_[93287]_ , \new_[93288]_ , \new_[93291]_ , \new_[93294]_ ,
    \new_[93295]_ , \new_[93298]_ , \new_[93301]_ , \new_[93302]_ ,
    \new_[93303]_ , \new_[93306]_ , \new_[93309]_ , \new_[93310]_ ,
    \new_[93313]_ , \new_[93316]_ , \new_[93317]_ , \new_[93318]_ ,
    \new_[93321]_ , \new_[93324]_ , \new_[93325]_ , \new_[93328]_ ,
    \new_[93331]_ , \new_[93332]_ , \new_[93333]_ , \new_[93336]_ ,
    \new_[93339]_ , \new_[93340]_ , \new_[93343]_ , \new_[93346]_ ,
    \new_[93347]_ , \new_[93348]_ , \new_[93351]_ , \new_[93354]_ ,
    \new_[93355]_ , \new_[93358]_ , \new_[93361]_ , \new_[93362]_ ,
    \new_[93363]_ , \new_[93366]_ , \new_[93369]_ , \new_[93370]_ ,
    \new_[93373]_ , \new_[93376]_ , \new_[93377]_ , \new_[93378]_ ,
    \new_[93381]_ , \new_[93384]_ , \new_[93385]_ , \new_[93388]_ ,
    \new_[93391]_ , \new_[93392]_ , \new_[93393]_ , \new_[93396]_ ,
    \new_[93399]_ , \new_[93400]_ , \new_[93403]_ , \new_[93406]_ ,
    \new_[93407]_ , \new_[93408]_ , \new_[93411]_ , \new_[93414]_ ,
    \new_[93415]_ , \new_[93418]_ , \new_[93421]_ , \new_[93422]_ ,
    \new_[93423]_ , \new_[93426]_ , \new_[93429]_ , \new_[93430]_ ,
    \new_[93433]_ , \new_[93436]_ , \new_[93437]_ , \new_[93438]_ ,
    \new_[93441]_ , \new_[93444]_ , \new_[93445]_ , \new_[93448]_ ,
    \new_[93451]_ , \new_[93452]_ , \new_[93453]_ , \new_[93456]_ ,
    \new_[93459]_ , \new_[93460]_ , \new_[93463]_ , \new_[93466]_ ,
    \new_[93467]_ , \new_[93468]_ , \new_[93471]_ , \new_[93474]_ ,
    \new_[93475]_ , \new_[93478]_ , \new_[93481]_ , \new_[93482]_ ,
    \new_[93483]_ , \new_[93486]_ , \new_[93489]_ , \new_[93490]_ ,
    \new_[93493]_ , \new_[93496]_ , \new_[93497]_ , \new_[93498]_ ,
    \new_[93501]_ , \new_[93504]_ , \new_[93505]_ , \new_[93508]_ ,
    \new_[93511]_ , \new_[93512]_ , \new_[93513]_ , \new_[93516]_ ,
    \new_[93519]_ , \new_[93520]_ , \new_[93523]_ , \new_[93526]_ ,
    \new_[93527]_ , \new_[93528]_ , \new_[93531]_ , \new_[93534]_ ,
    \new_[93535]_ , \new_[93538]_ , \new_[93541]_ , \new_[93542]_ ,
    \new_[93543]_ , \new_[93546]_ , \new_[93549]_ , \new_[93550]_ ,
    \new_[93553]_ , \new_[93556]_ , \new_[93557]_ , \new_[93558]_ ,
    \new_[93561]_ , \new_[93564]_ , \new_[93565]_ , \new_[93568]_ ,
    \new_[93571]_ , \new_[93572]_ , \new_[93573]_ , \new_[93576]_ ,
    \new_[93579]_ , \new_[93580]_ , \new_[93583]_ , \new_[93586]_ ,
    \new_[93587]_ , \new_[93588]_ , \new_[93591]_ , \new_[93594]_ ,
    \new_[93595]_ , \new_[93598]_ , \new_[93601]_ , \new_[93602]_ ,
    \new_[93603]_ , \new_[93606]_ , \new_[93609]_ , \new_[93610]_ ,
    \new_[93613]_ , \new_[93616]_ , \new_[93617]_ , \new_[93618]_ ,
    \new_[93621]_ , \new_[93624]_ , \new_[93625]_ , \new_[93628]_ ,
    \new_[93631]_ , \new_[93632]_ , \new_[93633]_ , \new_[93636]_ ,
    \new_[93639]_ , \new_[93640]_ , \new_[93643]_ , \new_[93646]_ ,
    \new_[93647]_ , \new_[93648]_ , \new_[93651]_ , \new_[93654]_ ,
    \new_[93655]_ , \new_[93658]_ , \new_[93661]_ , \new_[93662]_ ,
    \new_[93663]_ , \new_[93666]_ , \new_[93669]_ , \new_[93670]_ ,
    \new_[93673]_ , \new_[93676]_ , \new_[93677]_ , \new_[93678]_ ,
    \new_[93681]_ , \new_[93684]_ , \new_[93685]_ , \new_[93688]_ ,
    \new_[93691]_ , \new_[93692]_ , \new_[93693]_ , \new_[93696]_ ,
    \new_[93699]_ , \new_[93700]_ , \new_[93703]_ , \new_[93706]_ ,
    \new_[93707]_ , \new_[93708]_ , \new_[93711]_ , \new_[93714]_ ,
    \new_[93715]_ , \new_[93718]_ , \new_[93721]_ , \new_[93722]_ ,
    \new_[93723]_ , \new_[93726]_ , \new_[93729]_ , \new_[93730]_ ,
    \new_[93733]_ , \new_[93736]_ , \new_[93737]_ , \new_[93738]_ ,
    \new_[93741]_ , \new_[93744]_ , \new_[93745]_ , \new_[93748]_ ,
    \new_[93751]_ , \new_[93752]_ , \new_[93753]_ , \new_[93756]_ ,
    \new_[93759]_ , \new_[93760]_ , \new_[93763]_ , \new_[93766]_ ,
    \new_[93767]_ , \new_[93768]_ , \new_[93771]_ , \new_[93774]_ ,
    \new_[93775]_ , \new_[93778]_ , \new_[93781]_ , \new_[93782]_ ,
    \new_[93783]_ , \new_[93786]_ , \new_[93789]_ , \new_[93790]_ ,
    \new_[93793]_ , \new_[93796]_ , \new_[93797]_ , \new_[93798]_ ,
    \new_[93801]_ , \new_[93804]_ , \new_[93805]_ , \new_[93808]_ ,
    \new_[93811]_ , \new_[93812]_ , \new_[93813]_ , \new_[93816]_ ,
    \new_[93819]_ , \new_[93820]_ , \new_[93823]_ , \new_[93826]_ ,
    \new_[93827]_ , \new_[93828]_ , \new_[93831]_ , \new_[93834]_ ,
    \new_[93835]_ , \new_[93838]_ , \new_[93841]_ , \new_[93842]_ ,
    \new_[93843]_ , \new_[93846]_ , \new_[93849]_ , \new_[93850]_ ,
    \new_[93853]_ , \new_[93856]_ , \new_[93857]_ , \new_[93858]_ ,
    \new_[93861]_ , \new_[93864]_ , \new_[93865]_ , \new_[93868]_ ,
    \new_[93871]_ , \new_[93872]_ , \new_[93873]_ , \new_[93876]_ ,
    \new_[93879]_ , \new_[93880]_ , \new_[93883]_ , \new_[93886]_ ,
    \new_[93887]_ , \new_[93888]_ , \new_[93891]_ , \new_[93894]_ ,
    \new_[93895]_ , \new_[93898]_ , \new_[93901]_ , \new_[93902]_ ,
    \new_[93903]_ , \new_[93906]_ , \new_[93909]_ , \new_[93910]_ ,
    \new_[93913]_ , \new_[93916]_ , \new_[93917]_ , \new_[93918]_ ,
    \new_[93921]_ , \new_[93924]_ , \new_[93925]_ , \new_[93928]_ ,
    \new_[93931]_ , \new_[93932]_ , \new_[93933]_ , \new_[93936]_ ,
    \new_[93939]_ , \new_[93940]_ , \new_[93943]_ , \new_[93946]_ ,
    \new_[93947]_ , \new_[93948]_ , \new_[93951]_ , \new_[93954]_ ,
    \new_[93955]_ , \new_[93958]_ , \new_[93961]_ , \new_[93962]_ ,
    \new_[93963]_ , \new_[93966]_ , \new_[93969]_ , \new_[93970]_ ,
    \new_[93973]_ , \new_[93976]_ , \new_[93977]_ , \new_[93978]_ ,
    \new_[93981]_ , \new_[93984]_ , \new_[93985]_ , \new_[93988]_ ,
    \new_[93991]_ , \new_[93992]_ , \new_[93993]_ , \new_[93996]_ ,
    \new_[93999]_ , \new_[94000]_ , \new_[94003]_ , \new_[94006]_ ,
    \new_[94007]_ , \new_[94008]_ , \new_[94011]_ , \new_[94014]_ ,
    \new_[94015]_ , \new_[94018]_ , \new_[94021]_ , \new_[94022]_ ,
    \new_[94023]_ , \new_[94026]_ , \new_[94029]_ , \new_[94030]_ ,
    \new_[94033]_ , \new_[94036]_ , \new_[94037]_ , \new_[94038]_ ,
    \new_[94041]_ , \new_[94044]_ , \new_[94045]_ , \new_[94048]_ ,
    \new_[94051]_ , \new_[94052]_ , \new_[94053]_ , \new_[94056]_ ,
    \new_[94059]_ , \new_[94060]_ , \new_[94063]_ , \new_[94066]_ ,
    \new_[94067]_ , \new_[94068]_ , \new_[94071]_ , \new_[94074]_ ,
    \new_[94075]_ , \new_[94078]_ , \new_[94081]_ , \new_[94082]_ ,
    \new_[94083]_ , \new_[94086]_ , \new_[94089]_ , \new_[94090]_ ,
    \new_[94093]_ , \new_[94096]_ , \new_[94097]_ , \new_[94098]_ ,
    \new_[94101]_ , \new_[94104]_ , \new_[94105]_ , \new_[94108]_ ,
    \new_[94111]_ , \new_[94112]_ , \new_[94113]_ , \new_[94116]_ ,
    \new_[94119]_ , \new_[94120]_ , \new_[94123]_ , \new_[94126]_ ,
    \new_[94127]_ , \new_[94128]_ , \new_[94131]_ , \new_[94134]_ ,
    \new_[94135]_ , \new_[94138]_ , \new_[94141]_ , \new_[94142]_ ,
    \new_[94143]_ , \new_[94146]_ , \new_[94149]_ , \new_[94150]_ ,
    \new_[94153]_ , \new_[94156]_ , \new_[94157]_ , \new_[94158]_ ,
    \new_[94161]_ , \new_[94164]_ , \new_[94165]_ , \new_[94168]_ ,
    \new_[94171]_ , \new_[94172]_ , \new_[94173]_ , \new_[94176]_ ,
    \new_[94179]_ , \new_[94180]_ , \new_[94183]_ , \new_[94186]_ ,
    \new_[94187]_ , \new_[94188]_ , \new_[94191]_ , \new_[94194]_ ,
    \new_[94195]_ , \new_[94198]_ , \new_[94201]_ , \new_[94202]_ ,
    \new_[94203]_ , \new_[94206]_ , \new_[94209]_ , \new_[94210]_ ,
    \new_[94213]_ , \new_[94216]_ , \new_[94217]_ , \new_[94218]_ ,
    \new_[94221]_ , \new_[94224]_ , \new_[94225]_ , \new_[94228]_ ,
    \new_[94231]_ , \new_[94232]_ , \new_[94233]_ , \new_[94236]_ ,
    \new_[94239]_ , \new_[94240]_ , \new_[94243]_ , \new_[94246]_ ,
    \new_[94247]_ , \new_[94248]_ , \new_[94251]_ , \new_[94254]_ ,
    \new_[94255]_ , \new_[94258]_ , \new_[94261]_ , \new_[94262]_ ,
    \new_[94263]_ , \new_[94266]_ , \new_[94269]_ , \new_[94270]_ ,
    \new_[94273]_ , \new_[94276]_ , \new_[94277]_ , \new_[94278]_ ,
    \new_[94281]_ , \new_[94284]_ , \new_[94285]_ , \new_[94288]_ ,
    \new_[94291]_ , \new_[94292]_ , \new_[94293]_ , \new_[94296]_ ,
    \new_[94299]_ , \new_[94300]_ , \new_[94303]_ , \new_[94306]_ ,
    \new_[94307]_ , \new_[94308]_ , \new_[94311]_ , \new_[94314]_ ,
    \new_[94315]_ , \new_[94318]_ , \new_[94321]_ , \new_[94322]_ ,
    \new_[94323]_ , \new_[94326]_ , \new_[94329]_ , \new_[94330]_ ,
    \new_[94333]_ , \new_[94336]_ , \new_[94337]_ , \new_[94338]_ ,
    \new_[94341]_ , \new_[94344]_ , \new_[94345]_ , \new_[94348]_ ,
    \new_[94351]_ , \new_[94352]_ , \new_[94353]_ , \new_[94356]_ ,
    \new_[94359]_ , \new_[94360]_ , \new_[94363]_ , \new_[94366]_ ,
    \new_[94367]_ , \new_[94368]_ , \new_[94371]_ , \new_[94374]_ ,
    \new_[94375]_ , \new_[94378]_ , \new_[94381]_ , \new_[94382]_ ,
    \new_[94383]_ , \new_[94386]_ , \new_[94389]_ , \new_[94390]_ ,
    \new_[94393]_ , \new_[94396]_ , \new_[94397]_ , \new_[94398]_ ,
    \new_[94401]_ , \new_[94404]_ , \new_[94405]_ , \new_[94408]_ ,
    \new_[94411]_ , \new_[94412]_ , \new_[94413]_ , \new_[94416]_ ,
    \new_[94419]_ , \new_[94420]_ , \new_[94423]_ , \new_[94426]_ ,
    \new_[94427]_ , \new_[94428]_ , \new_[94431]_ , \new_[94434]_ ,
    \new_[94435]_ , \new_[94438]_ , \new_[94441]_ , \new_[94442]_ ,
    \new_[94443]_ , \new_[94446]_ , \new_[94449]_ , \new_[94450]_ ,
    \new_[94453]_ , \new_[94456]_ , \new_[94457]_ , \new_[94458]_ ,
    \new_[94461]_ , \new_[94464]_ , \new_[94465]_ , \new_[94468]_ ,
    \new_[94471]_ , \new_[94472]_ , \new_[94473]_ , \new_[94476]_ ,
    \new_[94479]_ , \new_[94480]_ , \new_[94483]_ , \new_[94486]_ ,
    \new_[94487]_ , \new_[94488]_ , \new_[94491]_ , \new_[94494]_ ,
    \new_[94495]_ , \new_[94498]_ , \new_[94501]_ , \new_[94502]_ ,
    \new_[94503]_ , \new_[94506]_ , \new_[94509]_ , \new_[94510]_ ,
    \new_[94513]_ , \new_[94516]_ , \new_[94517]_ , \new_[94518]_ ,
    \new_[94521]_ , \new_[94524]_ , \new_[94525]_ , \new_[94528]_ ,
    \new_[94531]_ , \new_[94532]_ , \new_[94533]_ , \new_[94536]_ ,
    \new_[94539]_ , \new_[94540]_ , \new_[94543]_ , \new_[94546]_ ,
    \new_[94547]_ , \new_[94548]_ , \new_[94551]_ , \new_[94554]_ ,
    \new_[94555]_ , \new_[94558]_ , \new_[94561]_ , \new_[94562]_ ,
    \new_[94563]_ , \new_[94566]_ , \new_[94569]_ , \new_[94570]_ ,
    \new_[94573]_ , \new_[94576]_ , \new_[94577]_ , \new_[94578]_ ,
    \new_[94581]_ , \new_[94584]_ , \new_[94585]_ , \new_[94588]_ ,
    \new_[94591]_ , \new_[94592]_ , \new_[94593]_ , \new_[94596]_ ,
    \new_[94599]_ , \new_[94600]_ , \new_[94603]_ , \new_[94606]_ ,
    \new_[94607]_ , \new_[94608]_ , \new_[94611]_ , \new_[94614]_ ,
    \new_[94615]_ , \new_[94618]_ , \new_[94621]_ , \new_[94622]_ ,
    \new_[94623]_ , \new_[94626]_ , \new_[94629]_ , \new_[94630]_ ,
    \new_[94633]_ , \new_[94636]_ , \new_[94637]_ , \new_[94638]_ ,
    \new_[94641]_ , \new_[94644]_ , \new_[94645]_ , \new_[94648]_ ,
    \new_[94651]_ , \new_[94652]_ , \new_[94653]_ , \new_[94656]_ ,
    \new_[94659]_ , \new_[94660]_ , \new_[94663]_ , \new_[94666]_ ,
    \new_[94667]_ , \new_[94668]_ , \new_[94671]_ , \new_[94674]_ ,
    \new_[94675]_ , \new_[94678]_ , \new_[94681]_ , \new_[94682]_ ,
    \new_[94683]_ , \new_[94686]_ , \new_[94689]_ , \new_[94690]_ ,
    \new_[94693]_ , \new_[94696]_ , \new_[94697]_ , \new_[94698]_ ,
    \new_[94701]_ , \new_[94704]_ , \new_[94705]_ , \new_[94708]_ ,
    \new_[94711]_ , \new_[94712]_ , \new_[94713]_ , \new_[94716]_ ,
    \new_[94719]_ , \new_[94720]_ , \new_[94723]_ , \new_[94726]_ ,
    \new_[94727]_ , \new_[94728]_ , \new_[94731]_ , \new_[94734]_ ,
    \new_[94735]_ , \new_[94738]_ , \new_[94741]_ , \new_[94742]_ ,
    \new_[94743]_ , \new_[94746]_ , \new_[94749]_ , \new_[94750]_ ,
    \new_[94753]_ , \new_[94756]_ , \new_[94757]_ , \new_[94758]_ ,
    \new_[94761]_ , \new_[94764]_ , \new_[94765]_ , \new_[94768]_ ,
    \new_[94771]_ , \new_[94772]_ , \new_[94773]_ , \new_[94776]_ ,
    \new_[94779]_ , \new_[94780]_ , \new_[94783]_ , \new_[94786]_ ,
    \new_[94787]_ , \new_[94788]_ , \new_[94791]_ , \new_[94794]_ ,
    \new_[94795]_ , \new_[94798]_ , \new_[94801]_ , \new_[94802]_ ,
    \new_[94803]_ , \new_[94806]_ , \new_[94809]_ , \new_[94810]_ ,
    \new_[94813]_ , \new_[94816]_ , \new_[94817]_ , \new_[94818]_ ,
    \new_[94821]_ , \new_[94824]_ , \new_[94825]_ , \new_[94828]_ ,
    \new_[94831]_ , \new_[94832]_ , \new_[94833]_ , \new_[94836]_ ,
    \new_[94839]_ , \new_[94840]_ , \new_[94843]_ , \new_[94846]_ ,
    \new_[94847]_ , \new_[94848]_ , \new_[94851]_ , \new_[94854]_ ,
    \new_[94855]_ , \new_[94858]_ , \new_[94861]_ , \new_[94862]_ ,
    \new_[94863]_ , \new_[94866]_ , \new_[94869]_ , \new_[94870]_ ,
    \new_[94873]_ , \new_[94876]_ , \new_[94877]_ , \new_[94878]_ ,
    \new_[94881]_ , \new_[94884]_ , \new_[94885]_ , \new_[94888]_ ,
    \new_[94891]_ , \new_[94892]_ , \new_[94893]_ , \new_[94896]_ ,
    \new_[94899]_ , \new_[94900]_ , \new_[94903]_ , \new_[94906]_ ,
    \new_[94907]_ , \new_[94908]_ , \new_[94911]_ , \new_[94914]_ ,
    \new_[94915]_ , \new_[94918]_ , \new_[94921]_ , \new_[94922]_ ,
    \new_[94923]_ , \new_[94926]_ , \new_[94929]_ , \new_[94930]_ ,
    \new_[94933]_ , \new_[94936]_ , \new_[94937]_ , \new_[94938]_ ,
    \new_[94941]_ , \new_[94944]_ , \new_[94945]_ , \new_[94948]_ ,
    \new_[94951]_ , \new_[94952]_ , \new_[94953]_ , \new_[94956]_ ,
    \new_[94959]_ , \new_[94960]_ , \new_[94963]_ , \new_[94966]_ ,
    \new_[94967]_ , \new_[94968]_ , \new_[94971]_ , \new_[94974]_ ,
    \new_[94975]_ , \new_[94978]_ , \new_[94981]_ , \new_[94982]_ ,
    \new_[94983]_ , \new_[94986]_ , \new_[94989]_ , \new_[94990]_ ,
    \new_[94993]_ , \new_[94996]_ , \new_[94997]_ , \new_[94998]_ ,
    \new_[95001]_ , \new_[95004]_ , \new_[95005]_ , \new_[95008]_ ,
    \new_[95011]_ , \new_[95012]_ , \new_[95013]_ , \new_[95016]_ ,
    \new_[95019]_ , \new_[95020]_ , \new_[95023]_ , \new_[95026]_ ,
    \new_[95027]_ , \new_[95028]_ , \new_[95031]_ , \new_[95034]_ ,
    \new_[95035]_ , \new_[95038]_ , \new_[95041]_ , \new_[95042]_ ,
    \new_[95043]_ , \new_[95046]_ , \new_[95049]_ , \new_[95050]_ ,
    \new_[95053]_ , \new_[95056]_ , \new_[95057]_ , \new_[95058]_ ,
    \new_[95061]_ , \new_[95064]_ , \new_[95065]_ , \new_[95068]_ ,
    \new_[95071]_ , \new_[95072]_ , \new_[95073]_ , \new_[95076]_ ,
    \new_[95079]_ , \new_[95080]_ , \new_[95083]_ , \new_[95086]_ ,
    \new_[95087]_ , \new_[95088]_ , \new_[95091]_ , \new_[95094]_ ,
    \new_[95095]_ , \new_[95098]_ , \new_[95101]_ , \new_[95102]_ ,
    \new_[95103]_ , \new_[95106]_ , \new_[95109]_ , \new_[95110]_ ,
    \new_[95113]_ , \new_[95116]_ , \new_[95117]_ , \new_[95118]_ ,
    \new_[95121]_ , \new_[95124]_ , \new_[95125]_ , \new_[95128]_ ,
    \new_[95131]_ , \new_[95132]_ , \new_[95133]_ , \new_[95136]_ ,
    \new_[95139]_ , \new_[95140]_ , \new_[95143]_ , \new_[95146]_ ,
    \new_[95147]_ , \new_[95148]_ , \new_[95151]_ , \new_[95154]_ ,
    \new_[95155]_ , \new_[95158]_ , \new_[95161]_ , \new_[95162]_ ,
    \new_[95163]_ , \new_[95166]_ , \new_[95169]_ , \new_[95170]_ ,
    \new_[95173]_ , \new_[95176]_ , \new_[95177]_ , \new_[95178]_ ,
    \new_[95181]_ , \new_[95184]_ , \new_[95185]_ , \new_[95188]_ ,
    \new_[95191]_ , \new_[95192]_ , \new_[95193]_ , \new_[95196]_ ,
    \new_[95199]_ , \new_[95200]_ , \new_[95203]_ , \new_[95206]_ ,
    \new_[95207]_ , \new_[95208]_ , \new_[95211]_ , \new_[95214]_ ,
    \new_[95215]_ , \new_[95218]_ , \new_[95221]_ , \new_[95222]_ ,
    \new_[95223]_ , \new_[95226]_ , \new_[95229]_ , \new_[95230]_ ,
    \new_[95233]_ , \new_[95236]_ , \new_[95237]_ , \new_[95238]_ ,
    \new_[95241]_ , \new_[95244]_ , \new_[95245]_ , \new_[95248]_ ,
    \new_[95251]_ , \new_[95252]_ , \new_[95253]_ , \new_[95256]_ ,
    \new_[95259]_ , \new_[95260]_ , \new_[95263]_ , \new_[95266]_ ,
    \new_[95267]_ , \new_[95268]_ , \new_[95271]_ , \new_[95274]_ ,
    \new_[95275]_ , \new_[95278]_ , \new_[95281]_ , \new_[95282]_ ,
    \new_[95283]_ , \new_[95286]_ , \new_[95289]_ , \new_[95290]_ ,
    \new_[95293]_ , \new_[95296]_ , \new_[95297]_ , \new_[95298]_ ,
    \new_[95301]_ , \new_[95304]_ , \new_[95305]_ , \new_[95308]_ ,
    \new_[95311]_ , \new_[95312]_ , \new_[95313]_ , \new_[95316]_ ,
    \new_[95319]_ , \new_[95320]_ , \new_[95323]_ , \new_[95326]_ ,
    \new_[95327]_ , \new_[95328]_ , \new_[95331]_ , \new_[95334]_ ,
    \new_[95335]_ , \new_[95338]_ , \new_[95341]_ , \new_[95342]_ ,
    \new_[95343]_ , \new_[95346]_ , \new_[95349]_ , \new_[95350]_ ,
    \new_[95353]_ , \new_[95356]_ , \new_[95357]_ , \new_[95358]_ ,
    \new_[95361]_ , \new_[95364]_ , \new_[95365]_ , \new_[95368]_ ,
    \new_[95371]_ , \new_[95372]_ , \new_[95373]_ , \new_[95376]_ ,
    \new_[95379]_ , \new_[95380]_ , \new_[95383]_ , \new_[95386]_ ,
    \new_[95387]_ , \new_[95388]_ , \new_[95391]_ , \new_[95394]_ ,
    \new_[95395]_ , \new_[95398]_ , \new_[95401]_ , \new_[95402]_ ,
    \new_[95403]_ , \new_[95406]_ , \new_[95409]_ , \new_[95410]_ ,
    \new_[95413]_ , \new_[95416]_ , \new_[95417]_ , \new_[95418]_ ,
    \new_[95421]_ , \new_[95424]_ , \new_[95425]_ , \new_[95428]_ ,
    \new_[95431]_ , \new_[95432]_ , \new_[95433]_ , \new_[95436]_ ,
    \new_[95439]_ , \new_[95440]_ , \new_[95443]_ , \new_[95446]_ ,
    \new_[95447]_ , \new_[95448]_ , \new_[95451]_ , \new_[95454]_ ,
    \new_[95455]_ , \new_[95458]_ , \new_[95461]_ , \new_[95462]_ ,
    \new_[95463]_ , \new_[95466]_ , \new_[95469]_ , \new_[95470]_ ,
    \new_[95473]_ , \new_[95476]_ , \new_[95477]_ , \new_[95478]_ ,
    \new_[95481]_ , \new_[95484]_ , \new_[95485]_ , \new_[95488]_ ,
    \new_[95491]_ , \new_[95492]_ , \new_[95493]_ , \new_[95496]_ ,
    \new_[95499]_ , \new_[95500]_ , \new_[95503]_ , \new_[95506]_ ,
    \new_[95507]_ , \new_[95508]_ , \new_[95511]_ , \new_[95514]_ ,
    \new_[95515]_ , \new_[95518]_ , \new_[95521]_ , \new_[95522]_ ,
    \new_[95523]_ , \new_[95526]_ , \new_[95529]_ , \new_[95530]_ ,
    \new_[95533]_ , \new_[95536]_ , \new_[95537]_ , \new_[95538]_ ,
    \new_[95541]_ , \new_[95544]_ , \new_[95545]_ , \new_[95548]_ ,
    \new_[95551]_ , \new_[95552]_ , \new_[95553]_ , \new_[95556]_ ,
    \new_[95559]_ , \new_[95560]_ , \new_[95563]_ , \new_[95566]_ ,
    \new_[95567]_ , \new_[95568]_ , \new_[95571]_ , \new_[95574]_ ,
    \new_[95575]_ , \new_[95578]_ , \new_[95581]_ , \new_[95582]_ ,
    \new_[95583]_ , \new_[95586]_ , \new_[95589]_ , \new_[95590]_ ,
    \new_[95593]_ , \new_[95596]_ , \new_[95597]_ , \new_[95598]_ ,
    \new_[95601]_ , \new_[95604]_ , \new_[95605]_ , \new_[95608]_ ,
    \new_[95611]_ , \new_[95612]_ , \new_[95613]_ , \new_[95616]_ ,
    \new_[95619]_ , \new_[95620]_ , \new_[95623]_ , \new_[95626]_ ,
    \new_[95627]_ , \new_[95628]_ , \new_[95631]_ , \new_[95634]_ ,
    \new_[95635]_ , \new_[95638]_ , \new_[95641]_ , \new_[95642]_ ,
    \new_[95643]_ , \new_[95646]_ , \new_[95649]_ , \new_[95650]_ ,
    \new_[95653]_ , \new_[95656]_ , \new_[95657]_ , \new_[95658]_ ,
    \new_[95661]_ , \new_[95664]_ , \new_[95665]_ , \new_[95668]_ ,
    \new_[95671]_ , \new_[95672]_ , \new_[95673]_ , \new_[95676]_ ,
    \new_[95679]_ , \new_[95680]_ , \new_[95683]_ , \new_[95686]_ ,
    \new_[95687]_ , \new_[95688]_ , \new_[95691]_ , \new_[95694]_ ,
    \new_[95695]_ , \new_[95698]_ , \new_[95701]_ , \new_[95702]_ ,
    \new_[95703]_ , \new_[95706]_ , \new_[95709]_ , \new_[95710]_ ,
    \new_[95713]_ , \new_[95716]_ , \new_[95717]_ , \new_[95718]_ ,
    \new_[95721]_ , \new_[95724]_ , \new_[95725]_ , \new_[95728]_ ,
    \new_[95731]_ , \new_[95732]_ , \new_[95733]_ , \new_[95736]_ ,
    \new_[95739]_ , \new_[95740]_ , \new_[95743]_ , \new_[95746]_ ,
    \new_[95747]_ , \new_[95748]_ , \new_[95751]_ , \new_[95754]_ ,
    \new_[95755]_ , \new_[95758]_ , \new_[95761]_ , \new_[95762]_ ,
    \new_[95763]_ , \new_[95766]_ , \new_[95769]_ , \new_[95770]_ ,
    \new_[95773]_ , \new_[95776]_ , \new_[95777]_ , \new_[95778]_ ,
    \new_[95781]_ , \new_[95784]_ , \new_[95785]_ , \new_[95788]_ ,
    \new_[95791]_ , \new_[95792]_ , \new_[95793]_ , \new_[95796]_ ,
    \new_[95799]_ , \new_[95800]_ , \new_[95803]_ , \new_[95806]_ ,
    \new_[95807]_ , \new_[95808]_ , \new_[95811]_ , \new_[95814]_ ,
    \new_[95815]_ , \new_[95818]_ , \new_[95821]_ , \new_[95822]_ ,
    \new_[95823]_ , \new_[95826]_ , \new_[95829]_ , \new_[95830]_ ,
    \new_[95833]_ , \new_[95836]_ , \new_[95837]_ , \new_[95838]_ ,
    \new_[95841]_ , \new_[95844]_ , \new_[95845]_ , \new_[95848]_ ,
    \new_[95851]_ , \new_[95852]_ , \new_[95853]_ , \new_[95856]_ ,
    \new_[95859]_ , \new_[95860]_ , \new_[95863]_ , \new_[95866]_ ,
    \new_[95867]_ , \new_[95868]_ , \new_[95871]_ , \new_[95874]_ ,
    \new_[95875]_ , \new_[95878]_ , \new_[95881]_ , \new_[95882]_ ,
    \new_[95883]_ , \new_[95886]_ , \new_[95889]_ , \new_[95890]_ ,
    \new_[95893]_ , \new_[95896]_ , \new_[95897]_ , \new_[95898]_ ,
    \new_[95901]_ , \new_[95904]_ , \new_[95905]_ , \new_[95908]_ ,
    \new_[95911]_ , \new_[95912]_ , \new_[95913]_ , \new_[95916]_ ,
    \new_[95919]_ , \new_[95920]_ , \new_[95923]_ , \new_[95926]_ ,
    \new_[95927]_ , \new_[95928]_ , \new_[95931]_ , \new_[95934]_ ,
    \new_[95935]_ , \new_[95938]_ , \new_[95941]_ , \new_[95942]_ ,
    \new_[95943]_ , \new_[95946]_ , \new_[95949]_ , \new_[95950]_ ,
    \new_[95953]_ , \new_[95956]_ , \new_[95957]_ , \new_[95958]_ ,
    \new_[95961]_ , \new_[95964]_ , \new_[95965]_ , \new_[95968]_ ,
    \new_[95971]_ , \new_[95972]_ , \new_[95973]_ , \new_[95976]_ ,
    \new_[95979]_ , \new_[95980]_ , \new_[95983]_ , \new_[95986]_ ,
    \new_[95987]_ , \new_[95988]_ , \new_[95991]_ , \new_[95994]_ ,
    \new_[95995]_ , \new_[95998]_ , \new_[96001]_ , \new_[96002]_ ,
    \new_[96003]_ , \new_[96006]_ , \new_[96009]_ , \new_[96010]_ ,
    \new_[96013]_ , \new_[96016]_ , \new_[96017]_ , \new_[96018]_ ,
    \new_[96021]_ , \new_[96024]_ , \new_[96025]_ , \new_[96028]_ ,
    \new_[96031]_ , \new_[96032]_ , \new_[96033]_ , \new_[96036]_ ,
    \new_[96039]_ , \new_[96040]_ , \new_[96043]_ , \new_[96046]_ ,
    \new_[96047]_ , \new_[96048]_ , \new_[96051]_ , \new_[96054]_ ,
    \new_[96055]_ , \new_[96058]_ , \new_[96061]_ , \new_[96062]_ ,
    \new_[96063]_ , \new_[96066]_ , \new_[96069]_ , \new_[96070]_ ,
    \new_[96073]_ , \new_[96076]_ , \new_[96077]_ , \new_[96078]_ ,
    \new_[96081]_ , \new_[96084]_ , \new_[96085]_ , \new_[96088]_ ,
    \new_[96091]_ , \new_[96092]_ , \new_[96093]_ , \new_[96096]_ ,
    \new_[96099]_ , \new_[96100]_ , \new_[96103]_ , \new_[96106]_ ,
    \new_[96107]_ , \new_[96108]_ , \new_[96111]_ , \new_[96114]_ ,
    \new_[96115]_ , \new_[96118]_ , \new_[96121]_ , \new_[96122]_ ,
    \new_[96123]_ , \new_[96126]_ , \new_[96129]_ , \new_[96130]_ ,
    \new_[96133]_ , \new_[96136]_ , \new_[96137]_ , \new_[96138]_ ,
    \new_[96141]_ , \new_[96144]_ , \new_[96145]_ , \new_[96148]_ ,
    \new_[96151]_ , \new_[96152]_ , \new_[96153]_ , \new_[96156]_ ,
    \new_[96159]_ , \new_[96160]_ , \new_[96163]_ , \new_[96166]_ ,
    \new_[96167]_ , \new_[96168]_ , \new_[96171]_ , \new_[96174]_ ,
    \new_[96175]_ , \new_[96178]_ , \new_[96181]_ , \new_[96182]_ ,
    \new_[96183]_ , \new_[96186]_ , \new_[96189]_ , \new_[96190]_ ,
    \new_[96193]_ , \new_[96196]_ , \new_[96197]_ , \new_[96198]_ ,
    \new_[96201]_ , \new_[96204]_ , \new_[96205]_ , \new_[96208]_ ,
    \new_[96211]_ , \new_[96212]_ , \new_[96213]_ , \new_[96216]_ ,
    \new_[96219]_ , \new_[96220]_ , \new_[96223]_ , \new_[96226]_ ,
    \new_[96227]_ , \new_[96228]_ , \new_[96231]_ , \new_[96234]_ ,
    \new_[96235]_ , \new_[96238]_ , \new_[96241]_ , \new_[96242]_ ,
    \new_[96243]_ , \new_[96246]_ , \new_[96249]_ , \new_[96250]_ ,
    \new_[96253]_ , \new_[96256]_ , \new_[96257]_ , \new_[96258]_ ,
    \new_[96261]_ , \new_[96264]_ , \new_[96265]_ , \new_[96268]_ ,
    \new_[96271]_ , \new_[96272]_ , \new_[96273]_ , \new_[96276]_ ,
    \new_[96279]_ , \new_[96280]_ , \new_[96283]_ , \new_[96286]_ ,
    \new_[96287]_ , \new_[96288]_ , \new_[96291]_ , \new_[96294]_ ,
    \new_[96295]_ , \new_[96298]_ , \new_[96301]_ , \new_[96302]_ ,
    \new_[96303]_ , \new_[96306]_ , \new_[96309]_ , \new_[96310]_ ,
    \new_[96313]_ , \new_[96316]_ , \new_[96317]_ , \new_[96318]_ ,
    \new_[96321]_ , \new_[96324]_ , \new_[96325]_ , \new_[96328]_ ,
    \new_[96331]_ , \new_[96332]_ , \new_[96333]_ , \new_[96336]_ ,
    \new_[96339]_ , \new_[96340]_ , \new_[96343]_ , \new_[96346]_ ,
    \new_[96347]_ , \new_[96348]_ , \new_[96351]_ , \new_[96354]_ ,
    \new_[96355]_ , \new_[96358]_ , \new_[96361]_ , \new_[96362]_ ,
    \new_[96363]_ , \new_[96366]_ , \new_[96369]_ , \new_[96370]_ ,
    \new_[96373]_ , \new_[96376]_ , \new_[96377]_ , \new_[96378]_ ,
    \new_[96381]_ , \new_[96384]_ , \new_[96385]_ , \new_[96388]_ ,
    \new_[96391]_ , \new_[96392]_ , \new_[96393]_ , \new_[96396]_ ,
    \new_[96399]_ , \new_[96400]_ , \new_[96403]_ , \new_[96406]_ ,
    \new_[96407]_ , \new_[96408]_ , \new_[96411]_ , \new_[96414]_ ,
    \new_[96415]_ , \new_[96418]_ , \new_[96421]_ , \new_[96422]_ ,
    \new_[96423]_ , \new_[96426]_ , \new_[96429]_ , \new_[96430]_ ,
    \new_[96433]_ , \new_[96436]_ , \new_[96437]_ , \new_[96438]_ ,
    \new_[96441]_ , \new_[96444]_ , \new_[96445]_ , \new_[96448]_ ,
    \new_[96451]_ , \new_[96452]_ , \new_[96453]_ , \new_[96456]_ ,
    \new_[96459]_ , \new_[96460]_ , \new_[96463]_ , \new_[96466]_ ,
    \new_[96467]_ , \new_[96468]_ , \new_[96471]_ , \new_[96474]_ ,
    \new_[96475]_ , \new_[96478]_ , \new_[96481]_ , \new_[96482]_ ,
    \new_[96483]_ , \new_[96486]_ , \new_[96489]_ , \new_[96490]_ ,
    \new_[96493]_ , \new_[96496]_ , \new_[96497]_ , \new_[96498]_ ,
    \new_[96501]_ , \new_[96504]_ , \new_[96505]_ , \new_[96508]_ ,
    \new_[96511]_ , \new_[96512]_ , \new_[96513]_ , \new_[96516]_ ,
    \new_[96519]_ , \new_[96520]_ , \new_[96523]_ , \new_[96526]_ ,
    \new_[96527]_ , \new_[96528]_ , \new_[96531]_ , \new_[96534]_ ,
    \new_[96535]_ , \new_[96538]_ , \new_[96541]_ , \new_[96542]_ ,
    \new_[96543]_ , \new_[96546]_ , \new_[96549]_ , \new_[96550]_ ,
    \new_[96553]_ , \new_[96556]_ , \new_[96557]_ , \new_[96558]_ ,
    \new_[96561]_ , \new_[96564]_ , \new_[96565]_ , \new_[96568]_ ,
    \new_[96571]_ , \new_[96572]_ , \new_[96573]_ , \new_[96576]_ ,
    \new_[96579]_ , \new_[96580]_ , \new_[96583]_ , \new_[96586]_ ,
    \new_[96587]_ , \new_[96588]_ , \new_[96591]_ , \new_[96594]_ ,
    \new_[96595]_ , \new_[96598]_ , \new_[96601]_ , \new_[96602]_ ,
    \new_[96603]_ , \new_[96606]_ , \new_[96609]_ , \new_[96610]_ ,
    \new_[96613]_ , \new_[96616]_ , \new_[96617]_ , \new_[96618]_ ,
    \new_[96621]_ , \new_[96624]_ , \new_[96625]_ , \new_[96628]_ ,
    \new_[96631]_ , \new_[96632]_ , \new_[96633]_ , \new_[96636]_ ,
    \new_[96639]_ , \new_[96640]_ , \new_[96643]_ , \new_[96646]_ ,
    \new_[96647]_ , \new_[96648]_ , \new_[96651]_ , \new_[96654]_ ,
    \new_[96655]_ , \new_[96658]_ , \new_[96661]_ , \new_[96662]_ ,
    \new_[96663]_ , \new_[96666]_ , \new_[96669]_ , \new_[96670]_ ,
    \new_[96673]_ , \new_[96676]_ , \new_[96677]_ , \new_[96678]_ ,
    \new_[96681]_ , \new_[96684]_ , \new_[96685]_ , \new_[96688]_ ,
    \new_[96691]_ , \new_[96692]_ , \new_[96693]_ , \new_[96696]_ ,
    \new_[96699]_ , \new_[96700]_ , \new_[96703]_ , \new_[96706]_ ,
    \new_[96707]_ , \new_[96708]_ , \new_[96711]_ , \new_[96714]_ ,
    \new_[96715]_ , \new_[96718]_ , \new_[96721]_ , \new_[96722]_ ,
    \new_[96723]_ , \new_[96726]_ , \new_[96729]_ , \new_[96730]_ ,
    \new_[96733]_ , \new_[96736]_ , \new_[96737]_ , \new_[96738]_ ,
    \new_[96741]_ , \new_[96744]_ , \new_[96745]_ , \new_[96748]_ ,
    \new_[96751]_ , \new_[96752]_ , \new_[96753]_ , \new_[96756]_ ,
    \new_[96759]_ , \new_[96760]_ , \new_[96763]_ , \new_[96766]_ ,
    \new_[96767]_ , \new_[96768]_ , \new_[96771]_ , \new_[96774]_ ,
    \new_[96775]_ , \new_[96778]_ , \new_[96781]_ , \new_[96782]_ ,
    \new_[96783]_ , \new_[96786]_ , \new_[96789]_ , \new_[96790]_ ,
    \new_[96793]_ , \new_[96796]_ , \new_[96797]_ , \new_[96798]_ ,
    \new_[96801]_ , \new_[96804]_ , \new_[96805]_ , \new_[96808]_ ,
    \new_[96811]_ , \new_[96812]_ , \new_[96813]_ , \new_[96816]_ ,
    \new_[96819]_ , \new_[96820]_ , \new_[96823]_ , \new_[96826]_ ,
    \new_[96827]_ , \new_[96828]_ , \new_[96831]_ , \new_[96834]_ ,
    \new_[96835]_ , \new_[96838]_ , \new_[96841]_ , \new_[96842]_ ,
    \new_[96843]_ , \new_[96846]_ , \new_[96849]_ , \new_[96850]_ ,
    \new_[96853]_ , \new_[96856]_ , \new_[96857]_ , \new_[96858]_ ,
    \new_[96861]_ , \new_[96864]_ , \new_[96865]_ , \new_[96868]_ ,
    \new_[96871]_ , \new_[96872]_ , \new_[96873]_ , \new_[96876]_ ,
    \new_[96879]_ , \new_[96880]_ , \new_[96883]_ , \new_[96886]_ ,
    \new_[96887]_ , \new_[96888]_ , \new_[96891]_ , \new_[96894]_ ,
    \new_[96895]_ , \new_[96898]_ , \new_[96901]_ , \new_[96902]_ ,
    \new_[96903]_ , \new_[96906]_ , \new_[96909]_ , \new_[96910]_ ,
    \new_[96913]_ , \new_[96916]_ , \new_[96917]_ , \new_[96918]_ ,
    \new_[96921]_ , \new_[96924]_ , \new_[96925]_ , \new_[96928]_ ,
    \new_[96931]_ , \new_[96932]_ , \new_[96933]_ , \new_[96936]_ ,
    \new_[96939]_ , \new_[96940]_ , \new_[96943]_ , \new_[96946]_ ,
    \new_[96947]_ , \new_[96948]_ , \new_[96951]_ , \new_[96954]_ ,
    \new_[96955]_ , \new_[96958]_ , \new_[96961]_ , \new_[96962]_ ,
    \new_[96963]_ , \new_[96966]_ , \new_[96969]_ , \new_[96970]_ ,
    \new_[96973]_ , \new_[96976]_ , \new_[96977]_ , \new_[96978]_ ,
    \new_[96981]_ , \new_[96984]_ , \new_[96985]_ , \new_[96988]_ ,
    \new_[96991]_ , \new_[96992]_ , \new_[96993]_ , \new_[96996]_ ,
    \new_[96999]_ , \new_[97000]_ , \new_[97003]_ , \new_[97006]_ ,
    \new_[97007]_ , \new_[97008]_ , \new_[97011]_ , \new_[97014]_ ,
    \new_[97015]_ , \new_[97018]_ , \new_[97021]_ , \new_[97022]_ ,
    \new_[97023]_ , \new_[97026]_ , \new_[97029]_ , \new_[97030]_ ,
    \new_[97033]_ , \new_[97036]_ , \new_[97037]_ , \new_[97038]_ ,
    \new_[97041]_ , \new_[97044]_ , \new_[97045]_ , \new_[97048]_ ,
    \new_[97051]_ , \new_[97052]_ , \new_[97053]_ , \new_[97056]_ ,
    \new_[97059]_ , \new_[97060]_ , \new_[97063]_ , \new_[97066]_ ,
    \new_[97067]_ , \new_[97068]_ , \new_[97071]_ , \new_[97074]_ ,
    \new_[97075]_ , \new_[97078]_ , \new_[97081]_ , \new_[97082]_ ,
    \new_[97083]_ , \new_[97086]_ , \new_[97089]_ , \new_[97090]_ ,
    \new_[97093]_ , \new_[97096]_ , \new_[97097]_ , \new_[97098]_ ,
    \new_[97101]_ , \new_[97104]_ , \new_[97105]_ , \new_[97108]_ ,
    \new_[97111]_ , \new_[97112]_ , \new_[97113]_ , \new_[97116]_ ,
    \new_[97119]_ , \new_[97120]_ , \new_[97123]_ , \new_[97126]_ ,
    \new_[97127]_ , \new_[97128]_ , \new_[97131]_ , \new_[97134]_ ,
    \new_[97135]_ , \new_[97138]_ , \new_[97141]_ , \new_[97142]_ ,
    \new_[97143]_ , \new_[97146]_ , \new_[97149]_ , \new_[97150]_ ,
    \new_[97153]_ , \new_[97156]_ , \new_[97157]_ , \new_[97158]_ ,
    \new_[97161]_ , \new_[97164]_ , \new_[97165]_ , \new_[97168]_ ,
    \new_[97171]_ , \new_[97172]_ , \new_[97173]_ , \new_[97176]_ ,
    \new_[97179]_ , \new_[97180]_ , \new_[97183]_ , \new_[97186]_ ,
    \new_[97187]_ , \new_[97188]_ , \new_[97191]_ , \new_[97194]_ ,
    \new_[97195]_ , \new_[97198]_ , \new_[97201]_ , \new_[97202]_ ,
    \new_[97203]_ , \new_[97206]_ , \new_[97209]_ , \new_[97210]_ ,
    \new_[97213]_ , \new_[97216]_ , \new_[97217]_ , \new_[97218]_ ,
    \new_[97221]_ , \new_[97224]_ , \new_[97225]_ , \new_[97228]_ ,
    \new_[97231]_ , \new_[97232]_ , \new_[97233]_ , \new_[97236]_ ,
    \new_[97239]_ , \new_[97240]_ , \new_[97243]_ , \new_[97246]_ ,
    \new_[97247]_ , \new_[97248]_ , \new_[97251]_ , \new_[97254]_ ,
    \new_[97255]_ , \new_[97258]_ , \new_[97261]_ , \new_[97262]_ ,
    \new_[97263]_ , \new_[97266]_ , \new_[97269]_ , \new_[97270]_ ,
    \new_[97273]_ , \new_[97276]_ , \new_[97277]_ , \new_[97278]_ ,
    \new_[97281]_ , \new_[97284]_ , \new_[97285]_ , \new_[97288]_ ,
    \new_[97291]_ , \new_[97292]_ , \new_[97293]_ , \new_[97296]_ ,
    \new_[97299]_ , \new_[97300]_ , \new_[97303]_ , \new_[97306]_ ,
    \new_[97307]_ , \new_[97308]_ , \new_[97311]_ , \new_[97314]_ ,
    \new_[97315]_ , \new_[97318]_ , \new_[97321]_ , \new_[97322]_ ,
    \new_[97323]_ , \new_[97326]_ , \new_[97329]_ , \new_[97330]_ ,
    \new_[97333]_ , \new_[97336]_ , \new_[97337]_ , \new_[97338]_ ,
    \new_[97341]_ , \new_[97344]_ , \new_[97345]_ , \new_[97348]_ ,
    \new_[97351]_ , \new_[97352]_ , \new_[97353]_ , \new_[97356]_ ,
    \new_[97359]_ , \new_[97360]_ , \new_[97363]_ , \new_[97366]_ ,
    \new_[97367]_ , \new_[97368]_ , \new_[97371]_ , \new_[97374]_ ,
    \new_[97375]_ , \new_[97378]_ , \new_[97381]_ , \new_[97382]_ ,
    \new_[97383]_ , \new_[97386]_ , \new_[97389]_ , \new_[97390]_ ,
    \new_[97393]_ , \new_[97396]_ , \new_[97397]_ , \new_[97398]_ ,
    \new_[97401]_ , \new_[97404]_ , \new_[97405]_ , \new_[97408]_ ,
    \new_[97411]_ , \new_[97412]_ , \new_[97413]_ , \new_[97416]_ ,
    \new_[97419]_ , \new_[97420]_ , \new_[97423]_ , \new_[97426]_ ,
    \new_[97427]_ , \new_[97428]_ , \new_[97431]_ , \new_[97434]_ ,
    \new_[97435]_ , \new_[97438]_ , \new_[97441]_ , \new_[97442]_ ,
    \new_[97443]_ , \new_[97446]_ , \new_[97449]_ , \new_[97450]_ ,
    \new_[97453]_ , \new_[97456]_ , \new_[97457]_ , \new_[97458]_ ,
    \new_[97461]_ , \new_[97464]_ , \new_[97465]_ , \new_[97468]_ ,
    \new_[97471]_ , \new_[97472]_ , \new_[97473]_ , \new_[97476]_ ,
    \new_[97479]_ , \new_[97480]_ , \new_[97483]_ , \new_[97486]_ ,
    \new_[97487]_ , \new_[97488]_ , \new_[97491]_ , \new_[97494]_ ,
    \new_[97495]_ , \new_[97498]_ , \new_[97501]_ , \new_[97502]_ ,
    \new_[97503]_ , \new_[97506]_ , \new_[97509]_ , \new_[97510]_ ,
    \new_[97513]_ , \new_[97516]_ , \new_[97517]_ , \new_[97518]_ ,
    \new_[97521]_ , \new_[97524]_ , \new_[97525]_ , \new_[97528]_ ,
    \new_[97531]_ , \new_[97532]_ , \new_[97533]_ , \new_[97536]_ ,
    \new_[97539]_ , \new_[97540]_ , \new_[97543]_ , \new_[97546]_ ,
    \new_[97547]_ , \new_[97548]_ , \new_[97551]_ , \new_[97554]_ ,
    \new_[97555]_ , \new_[97558]_ , \new_[97561]_ , \new_[97562]_ ,
    \new_[97563]_ , \new_[97566]_ , \new_[97569]_ , \new_[97570]_ ,
    \new_[97573]_ , \new_[97576]_ , \new_[97577]_ , \new_[97578]_ ,
    \new_[97581]_ , \new_[97584]_ , \new_[97585]_ , \new_[97588]_ ,
    \new_[97591]_ , \new_[97592]_ , \new_[97593]_ , \new_[97596]_ ,
    \new_[97599]_ , \new_[97600]_ , \new_[97603]_ , \new_[97606]_ ,
    \new_[97607]_ , \new_[97608]_ , \new_[97611]_ , \new_[97614]_ ,
    \new_[97615]_ , \new_[97618]_ , \new_[97621]_ , \new_[97622]_ ,
    \new_[97623]_ , \new_[97626]_ , \new_[97629]_ , \new_[97630]_ ,
    \new_[97633]_ , \new_[97636]_ , \new_[97637]_ , \new_[97638]_ ,
    \new_[97641]_ , \new_[97644]_ , \new_[97645]_ , \new_[97648]_ ,
    \new_[97651]_ , \new_[97652]_ , \new_[97653]_ , \new_[97656]_ ,
    \new_[97659]_ , \new_[97660]_ , \new_[97663]_ , \new_[97666]_ ,
    \new_[97667]_ , \new_[97668]_ , \new_[97671]_ , \new_[97674]_ ,
    \new_[97675]_ , \new_[97678]_ , \new_[97681]_ , \new_[97682]_ ,
    \new_[97683]_ , \new_[97686]_ , \new_[97689]_ , \new_[97690]_ ,
    \new_[97693]_ , \new_[97696]_ , \new_[97697]_ , \new_[97698]_ ,
    \new_[97701]_ , \new_[97704]_ , \new_[97705]_ , \new_[97708]_ ,
    \new_[97711]_ , \new_[97712]_ , \new_[97713]_ , \new_[97716]_ ,
    \new_[97719]_ , \new_[97720]_ , \new_[97723]_ , \new_[97726]_ ,
    \new_[97727]_ , \new_[97728]_ , \new_[97731]_ , \new_[97734]_ ,
    \new_[97735]_ , \new_[97738]_ , \new_[97741]_ , \new_[97742]_ ,
    \new_[97743]_ , \new_[97746]_ , \new_[97749]_ , \new_[97750]_ ,
    \new_[97753]_ , \new_[97756]_ , \new_[97757]_ , \new_[97758]_ ,
    \new_[97761]_ , \new_[97764]_ , \new_[97765]_ , \new_[97768]_ ,
    \new_[97771]_ , \new_[97772]_ , \new_[97773]_ , \new_[97776]_ ,
    \new_[97779]_ , \new_[97780]_ , \new_[97783]_ , \new_[97786]_ ,
    \new_[97787]_ , \new_[97788]_ , \new_[97791]_ , \new_[97794]_ ,
    \new_[97795]_ , \new_[97798]_ , \new_[97801]_ , \new_[97802]_ ,
    \new_[97803]_ , \new_[97806]_ , \new_[97809]_ , \new_[97810]_ ,
    \new_[97813]_ , \new_[97816]_ , \new_[97817]_ , \new_[97818]_ ,
    \new_[97821]_ , \new_[97824]_ , \new_[97825]_ , \new_[97828]_ ,
    \new_[97831]_ , \new_[97832]_ , \new_[97833]_ , \new_[97836]_ ,
    \new_[97839]_ , \new_[97840]_ , \new_[97843]_ , \new_[97846]_ ,
    \new_[97847]_ , \new_[97848]_ , \new_[97851]_ , \new_[97854]_ ,
    \new_[97855]_ , \new_[97858]_ , \new_[97861]_ , \new_[97862]_ ,
    \new_[97863]_ , \new_[97866]_ , \new_[97869]_ , \new_[97870]_ ,
    \new_[97873]_ , \new_[97876]_ , \new_[97877]_ , \new_[97878]_ ,
    \new_[97881]_ , \new_[97884]_ , \new_[97885]_ , \new_[97888]_ ,
    \new_[97891]_ , \new_[97892]_ , \new_[97893]_ , \new_[97896]_ ,
    \new_[97899]_ , \new_[97900]_ , \new_[97903]_ , \new_[97906]_ ,
    \new_[97907]_ , \new_[97908]_ , \new_[97911]_ , \new_[97914]_ ,
    \new_[97915]_ , \new_[97918]_ , \new_[97921]_ , \new_[97922]_ ,
    \new_[97923]_ , \new_[97926]_ , \new_[97929]_ , \new_[97930]_ ,
    \new_[97933]_ , \new_[97936]_ , \new_[97937]_ , \new_[97938]_ ,
    \new_[97941]_ , \new_[97944]_ , \new_[97945]_ , \new_[97948]_ ,
    \new_[97951]_ , \new_[97952]_ , \new_[97953]_ , \new_[97956]_ ,
    \new_[97959]_ , \new_[97960]_ , \new_[97963]_ , \new_[97966]_ ,
    \new_[97967]_ , \new_[97968]_ , \new_[97971]_ , \new_[97974]_ ,
    \new_[97975]_ , \new_[97978]_ , \new_[97981]_ , \new_[97982]_ ,
    \new_[97983]_ , \new_[97986]_ , \new_[97989]_ , \new_[97990]_ ,
    \new_[97993]_ , \new_[97996]_ , \new_[97997]_ , \new_[97998]_ ,
    \new_[98001]_ , \new_[98004]_ , \new_[98005]_ , \new_[98008]_ ,
    \new_[98011]_ , \new_[98012]_ , \new_[98013]_ , \new_[98016]_ ,
    \new_[98019]_ , \new_[98020]_ , \new_[98023]_ , \new_[98026]_ ,
    \new_[98027]_ , \new_[98028]_ , \new_[98031]_ , \new_[98034]_ ,
    \new_[98035]_ , \new_[98038]_ , \new_[98041]_ , \new_[98042]_ ,
    \new_[98043]_ , \new_[98046]_ , \new_[98049]_ , \new_[98050]_ ,
    \new_[98053]_ , \new_[98056]_ , \new_[98057]_ , \new_[98058]_ ,
    \new_[98061]_ , \new_[98064]_ , \new_[98065]_ , \new_[98068]_ ,
    \new_[98071]_ , \new_[98072]_ , \new_[98073]_ , \new_[98076]_ ,
    \new_[98079]_ , \new_[98080]_ , \new_[98083]_ , \new_[98086]_ ,
    \new_[98087]_ , \new_[98088]_ , \new_[98091]_ , \new_[98094]_ ,
    \new_[98095]_ , \new_[98098]_ , \new_[98101]_ , \new_[98102]_ ,
    \new_[98103]_ , \new_[98106]_ , \new_[98109]_ , \new_[98110]_ ,
    \new_[98113]_ , \new_[98116]_ , \new_[98117]_ , \new_[98118]_ ,
    \new_[98121]_ , \new_[98124]_ , \new_[98125]_ , \new_[98128]_ ,
    \new_[98131]_ , \new_[98132]_ , \new_[98133]_ , \new_[98136]_ ,
    \new_[98139]_ , \new_[98140]_ , \new_[98143]_ , \new_[98146]_ ,
    \new_[98147]_ , \new_[98148]_ , \new_[98151]_ , \new_[98154]_ ,
    \new_[98155]_ , \new_[98158]_ , \new_[98161]_ , \new_[98162]_ ,
    \new_[98163]_ , \new_[98166]_ , \new_[98169]_ , \new_[98170]_ ,
    \new_[98173]_ , \new_[98176]_ , \new_[98177]_ , \new_[98178]_ ,
    \new_[98181]_ , \new_[98184]_ , \new_[98185]_ , \new_[98188]_ ,
    \new_[98191]_ , \new_[98192]_ , \new_[98193]_ , \new_[98196]_ ,
    \new_[98199]_ , \new_[98200]_ , \new_[98203]_ , \new_[98206]_ ,
    \new_[98207]_ , \new_[98208]_ , \new_[98211]_ , \new_[98214]_ ,
    \new_[98215]_ , \new_[98218]_ , \new_[98221]_ , \new_[98222]_ ,
    \new_[98223]_ , \new_[98226]_ , \new_[98229]_ , \new_[98230]_ ,
    \new_[98233]_ , \new_[98236]_ , \new_[98237]_ , \new_[98238]_ ,
    \new_[98241]_ , \new_[98244]_ , \new_[98245]_ , \new_[98248]_ ,
    \new_[98251]_ , \new_[98252]_ , \new_[98253]_ , \new_[98256]_ ,
    \new_[98259]_ , \new_[98260]_ , \new_[98263]_ , \new_[98266]_ ,
    \new_[98267]_ , \new_[98268]_ , \new_[98271]_ , \new_[98274]_ ,
    \new_[98275]_ , \new_[98278]_ , \new_[98281]_ , \new_[98282]_ ,
    \new_[98283]_ , \new_[98286]_ , \new_[98289]_ , \new_[98290]_ ,
    \new_[98293]_ , \new_[98296]_ , \new_[98297]_ , \new_[98298]_ ,
    \new_[98301]_ , \new_[98304]_ , \new_[98305]_ , \new_[98308]_ ,
    \new_[98311]_ , \new_[98312]_ , \new_[98313]_ , \new_[98316]_ ,
    \new_[98319]_ , \new_[98320]_ , \new_[98323]_ , \new_[98326]_ ,
    \new_[98327]_ , \new_[98328]_ , \new_[98331]_ , \new_[98334]_ ,
    \new_[98335]_ , \new_[98338]_ , \new_[98341]_ , \new_[98342]_ ,
    \new_[98343]_ , \new_[98346]_ , \new_[98349]_ , \new_[98350]_ ,
    \new_[98353]_ , \new_[98356]_ , \new_[98357]_ , \new_[98358]_ ,
    \new_[98361]_ , \new_[98364]_ , \new_[98365]_ , \new_[98368]_ ,
    \new_[98371]_ , \new_[98372]_ , \new_[98373]_ , \new_[98376]_ ,
    \new_[98379]_ , \new_[98380]_ , \new_[98383]_ , \new_[98386]_ ,
    \new_[98387]_ , \new_[98388]_ , \new_[98391]_ , \new_[98394]_ ,
    \new_[98395]_ , \new_[98398]_ , \new_[98401]_ , \new_[98402]_ ,
    \new_[98403]_ , \new_[98406]_ , \new_[98409]_ , \new_[98410]_ ,
    \new_[98413]_ , \new_[98416]_ , \new_[98417]_ , \new_[98418]_ ,
    \new_[98421]_ , \new_[98424]_ , \new_[98425]_ , \new_[98428]_ ,
    \new_[98431]_ , \new_[98432]_ , \new_[98433]_ , \new_[98436]_ ,
    \new_[98439]_ , \new_[98440]_ , \new_[98443]_ , \new_[98446]_ ,
    \new_[98447]_ , \new_[98448]_ , \new_[98451]_ , \new_[98454]_ ,
    \new_[98455]_ , \new_[98458]_ , \new_[98461]_ , \new_[98462]_ ,
    \new_[98463]_ , \new_[98466]_ , \new_[98469]_ , \new_[98470]_ ,
    \new_[98473]_ , \new_[98476]_ , \new_[98477]_ , \new_[98478]_ ,
    \new_[98481]_ , \new_[98484]_ , \new_[98485]_ , \new_[98488]_ ,
    \new_[98491]_ , \new_[98492]_ , \new_[98493]_ , \new_[98496]_ ,
    \new_[98499]_ , \new_[98500]_ , \new_[98503]_ , \new_[98506]_ ,
    \new_[98507]_ , \new_[98508]_ , \new_[98511]_ , \new_[98514]_ ,
    \new_[98515]_ , \new_[98518]_ , \new_[98521]_ , \new_[98522]_ ,
    \new_[98523]_ , \new_[98526]_ , \new_[98529]_ , \new_[98530]_ ,
    \new_[98533]_ , \new_[98536]_ , \new_[98537]_ , \new_[98538]_ ,
    \new_[98541]_ , \new_[98544]_ , \new_[98545]_ , \new_[98548]_ ,
    \new_[98551]_ , \new_[98552]_ , \new_[98553]_ , \new_[98556]_ ,
    \new_[98559]_ , \new_[98560]_ , \new_[98563]_ , \new_[98566]_ ,
    \new_[98567]_ , \new_[98568]_ , \new_[98571]_ , \new_[98574]_ ,
    \new_[98575]_ , \new_[98578]_ , \new_[98581]_ , \new_[98582]_ ,
    \new_[98583]_ , \new_[98586]_ , \new_[98589]_ , \new_[98590]_ ,
    \new_[98593]_ , \new_[98596]_ , \new_[98597]_ , \new_[98598]_ ,
    \new_[98601]_ , \new_[98604]_ , \new_[98605]_ , \new_[98608]_ ,
    \new_[98611]_ , \new_[98612]_ , \new_[98613]_ , \new_[98616]_ ,
    \new_[98619]_ , \new_[98620]_ , \new_[98623]_ , \new_[98626]_ ,
    \new_[98627]_ , \new_[98628]_ , \new_[98631]_ , \new_[98634]_ ,
    \new_[98635]_ , \new_[98638]_ , \new_[98641]_ , \new_[98642]_ ,
    \new_[98643]_ , \new_[98646]_ , \new_[98649]_ , \new_[98650]_ ,
    \new_[98653]_ , \new_[98656]_ , \new_[98657]_ , \new_[98658]_ ,
    \new_[98661]_ , \new_[98664]_ , \new_[98665]_ , \new_[98668]_ ,
    \new_[98671]_ , \new_[98672]_ , \new_[98673]_ , \new_[98676]_ ,
    \new_[98679]_ , \new_[98680]_ , \new_[98683]_ , \new_[98686]_ ,
    \new_[98687]_ , \new_[98688]_ , \new_[98691]_ , \new_[98694]_ ,
    \new_[98695]_ , \new_[98698]_ , \new_[98701]_ , \new_[98702]_ ,
    \new_[98703]_ , \new_[98706]_ , \new_[98709]_ , \new_[98710]_ ,
    \new_[98713]_ , \new_[98716]_ , \new_[98717]_ , \new_[98718]_ ,
    \new_[98721]_ , \new_[98724]_ , \new_[98725]_ , \new_[98728]_ ,
    \new_[98731]_ , \new_[98732]_ , \new_[98733]_ , \new_[98736]_ ,
    \new_[98739]_ , \new_[98740]_ , \new_[98743]_ , \new_[98746]_ ,
    \new_[98747]_ , \new_[98748]_ , \new_[98751]_ , \new_[98754]_ ,
    \new_[98755]_ , \new_[98758]_ , \new_[98761]_ , \new_[98762]_ ,
    \new_[98763]_ , \new_[98766]_ , \new_[98769]_ , \new_[98770]_ ,
    \new_[98773]_ , \new_[98776]_ , \new_[98777]_ , \new_[98778]_ ,
    \new_[98781]_ , \new_[98784]_ , \new_[98785]_ , \new_[98788]_ ,
    \new_[98791]_ , \new_[98792]_ , \new_[98793]_ , \new_[98796]_ ,
    \new_[98799]_ , \new_[98800]_ , \new_[98803]_ , \new_[98806]_ ,
    \new_[98807]_ , \new_[98808]_ , \new_[98811]_ , \new_[98814]_ ,
    \new_[98815]_ , \new_[98818]_ , \new_[98821]_ , \new_[98822]_ ,
    \new_[98823]_ , \new_[98826]_ , \new_[98829]_ , \new_[98830]_ ,
    \new_[98833]_ , \new_[98836]_ , \new_[98837]_ , \new_[98838]_ ,
    \new_[98841]_ , \new_[98844]_ , \new_[98845]_ , \new_[98848]_ ,
    \new_[98851]_ , \new_[98852]_ , \new_[98853]_ , \new_[98856]_ ,
    \new_[98859]_ , \new_[98860]_ , \new_[98863]_ , \new_[98866]_ ,
    \new_[98867]_ , \new_[98868]_ , \new_[98871]_ , \new_[98874]_ ,
    \new_[98875]_ , \new_[98878]_ , \new_[98881]_ , \new_[98882]_ ,
    \new_[98883]_ , \new_[98886]_ , \new_[98889]_ , \new_[98890]_ ,
    \new_[98893]_ , \new_[98896]_ , \new_[98897]_ , \new_[98898]_ ,
    \new_[98901]_ , \new_[98904]_ , \new_[98905]_ , \new_[98908]_ ,
    \new_[98911]_ , \new_[98912]_ , \new_[98913]_ , \new_[98916]_ ,
    \new_[98919]_ , \new_[98920]_ , \new_[98923]_ , \new_[98926]_ ,
    \new_[98927]_ , \new_[98928]_ , \new_[98931]_ , \new_[98934]_ ,
    \new_[98935]_ , \new_[98938]_ , \new_[98941]_ , \new_[98942]_ ,
    \new_[98943]_ , \new_[98946]_ , \new_[98949]_ , \new_[98950]_ ,
    \new_[98953]_ , \new_[98956]_ , \new_[98957]_ , \new_[98958]_ ,
    \new_[98961]_ , \new_[98964]_ , \new_[98965]_ , \new_[98968]_ ,
    \new_[98971]_ , \new_[98972]_ , \new_[98973]_ , \new_[98976]_ ,
    \new_[98979]_ , \new_[98980]_ , \new_[98983]_ , \new_[98986]_ ,
    \new_[98987]_ , \new_[98988]_ , \new_[98991]_ , \new_[98994]_ ,
    \new_[98995]_ , \new_[98998]_ , \new_[99001]_ , \new_[99002]_ ,
    \new_[99003]_ , \new_[99006]_ , \new_[99009]_ , \new_[99010]_ ,
    \new_[99013]_ , \new_[99016]_ , \new_[99017]_ , \new_[99018]_ ,
    \new_[99021]_ , \new_[99024]_ , \new_[99025]_ , \new_[99028]_ ,
    \new_[99031]_ , \new_[99032]_ , \new_[99033]_ , \new_[99036]_ ,
    \new_[99039]_ , \new_[99040]_ , \new_[99043]_ , \new_[99046]_ ,
    \new_[99047]_ , \new_[99048]_ , \new_[99051]_ , \new_[99054]_ ,
    \new_[99055]_ , \new_[99058]_ , \new_[99061]_ , \new_[99062]_ ,
    \new_[99063]_ , \new_[99066]_ , \new_[99069]_ , \new_[99070]_ ,
    \new_[99073]_ , \new_[99076]_ , \new_[99077]_ , \new_[99078]_ ,
    \new_[99081]_ , \new_[99084]_ , \new_[99085]_ , \new_[99088]_ ,
    \new_[99091]_ , \new_[99092]_ , \new_[99093]_ , \new_[99096]_ ,
    \new_[99099]_ , \new_[99100]_ , \new_[99103]_ , \new_[99106]_ ,
    \new_[99107]_ , \new_[99108]_ , \new_[99111]_ , \new_[99114]_ ,
    \new_[99115]_ , \new_[99118]_ , \new_[99121]_ , \new_[99122]_ ,
    \new_[99123]_ , \new_[99126]_ , \new_[99129]_ , \new_[99130]_ ,
    \new_[99133]_ , \new_[99136]_ , \new_[99137]_ , \new_[99138]_ ,
    \new_[99141]_ , \new_[99144]_ , \new_[99145]_ , \new_[99148]_ ,
    \new_[99151]_ , \new_[99152]_ , \new_[99153]_ , \new_[99156]_ ,
    \new_[99159]_ , \new_[99160]_ , \new_[99163]_ , \new_[99166]_ ,
    \new_[99167]_ , \new_[99168]_ , \new_[99171]_ , \new_[99174]_ ,
    \new_[99175]_ , \new_[99178]_ , \new_[99181]_ , \new_[99182]_ ,
    \new_[99183]_ , \new_[99186]_ , \new_[99189]_ , \new_[99190]_ ,
    \new_[99193]_ , \new_[99196]_ , \new_[99197]_ , \new_[99198]_ ,
    \new_[99201]_ , \new_[99204]_ , \new_[99205]_ , \new_[99208]_ ,
    \new_[99211]_ , \new_[99212]_ , \new_[99213]_ , \new_[99216]_ ,
    \new_[99219]_ , \new_[99220]_ , \new_[99223]_ , \new_[99226]_ ,
    \new_[99227]_ , \new_[99228]_ , \new_[99231]_ , \new_[99234]_ ,
    \new_[99235]_ , \new_[99238]_ , \new_[99241]_ , \new_[99242]_ ,
    \new_[99243]_ , \new_[99246]_ , \new_[99249]_ , \new_[99250]_ ,
    \new_[99253]_ , \new_[99256]_ , \new_[99257]_ , \new_[99258]_ ,
    \new_[99261]_ , \new_[99264]_ , \new_[99265]_ , \new_[99268]_ ,
    \new_[99271]_ , \new_[99272]_ , \new_[99273]_ , \new_[99276]_ ,
    \new_[99279]_ , \new_[99280]_ , \new_[99283]_ , \new_[99286]_ ,
    \new_[99287]_ , \new_[99288]_ , \new_[99291]_ , \new_[99294]_ ,
    \new_[99295]_ , \new_[99298]_ , \new_[99301]_ , \new_[99302]_ ,
    \new_[99303]_ , \new_[99306]_ , \new_[99309]_ , \new_[99310]_ ,
    \new_[99313]_ , \new_[99316]_ , \new_[99317]_ , \new_[99318]_ ,
    \new_[99321]_ , \new_[99324]_ , \new_[99325]_ , \new_[99328]_ ,
    \new_[99331]_ , \new_[99332]_ , \new_[99333]_ , \new_[99336]_ ,
    \new_[99339]_ , \new_[99340]_ , \new_[99343]_ , \new_[99346]_ ,
    \new_[99347]_ , \new_[99348]_ , \new_[99351]_ , \new_[99354]_ ,
    \new_[99355]_ , \new_[99358]_ , \new_[99361]_ , \new_[99362]_ ,
    \new_[99363]_ , \new_[99366]_ , \new_[99369]_ , \new_[99370]_ ,
    \new_[99373]_ , \new_[99376]_ , \new_[99377]_ , \new_[99378]_ ,
    \new_[99381]_ , \new_[99384]_ , \new_[99385]_ , \new_[99388]_ ,
    \new_[99391]_ , \new_[99392]_ , \new_[99393]_ , \new_[99396]_ ,
    \new_[99399]_ , \new_[99400]_ , \new_[99403]_ , \new_[99406]_ ,
    \new_[99407]_ , \new_[99408]_ , \new_[99411]_ , \new_[99414]_ ,
    \new_[99415]_ , \new_[99418]_ , \new_[99421]_ , \new_[99422]_ ,
    \new_[99423]_ , \new_[99426]_ , \new_[99429]_ , \new_[99430]_ ,
    \new_[99433]_ , \new_[99436]_ , \new_[99437]_ , \new_[99438]_ ,
    \new_[99441]_ , \new_[99444]_ , \new_[99445]_ , \new_[99448]_ ,
    \new_[99451]_ , \new_[99452]_ , \new_[99453]_ , \new_[99456]_ ,
    \new_[99459]_ , \new_[99460]_ , \new_[99463]_ , \new_[99466]_ ,
    \new_[99467]_ , \new_[99468]_ , \new_[99471]_ , \new_[99474]_ ,
    \new_[99475]_ , \new_[99478]_ , \new_[99481]_ , \new_[99482]_ ,
    \new_[99483]_ , \new_[99486]_ , \new_[99489]_ , \new_[99490]_ ,
    \new_[99493]_ , \new_[99496]_ , \new_[99497]_ , \new_[99498]_ ,
    \new_[99501]_ , \new_[99504]_ , \new_[99505]_ , \new_[99508]_ ,
    \new_[99511]_ , \new_[99512]_ , \new_[99513]_ , \new_[99516]_ ,
    \new_[99519]_ , \new_[99520]_ , \new_[99523]_ , \new_[99526]_ ,
    \new_[99527]_ , \new_[99528]_ , \new_[99531]_ , \new_[99534]_ ,
    \new_[99535]_ , \new_[99538]_ , \new_[99541]_ , \new_[99542]_ ,
    \new_[99543]_ , \new_[99546]_ , \new_[99549]_ , \new_[99550]_ ,
    \new_[99553]_ , \new_[99556]_ , \new_[99557]_ , \new_[99558]_ ,
    \new_[99561]_ , \new_[99564]_ , \new_[99565]_ , \new_[99568]_ ,
    \new_[99571]_ , \new_[99572]_ , \new_[99573]_ , \new_[99576]_ ,
    \new_[99579]_ , \new_[99580]_ , \new_[99583]_ , \new_[99586]_ ,
    \new_[99587]_ , \new_[99588]_ , \new_[99591]_ , \new_[99594]_ ,
    \new_[99595]_ , \new_[99598]_ , \new_[99601]_ , \new_[99602]_ ,
    \new_[99603]_ , \new_[99606]_ , \new_[99609]_ , \new_[99610]_ ,
    \new_[99613]_ , \new_[99616]_ , \new_[99617]_ , \new_[99618]_ ,
    \new_[99621]_ , \new_[99624]_ , \new_[99625]_ , \new_[99628]_ ,
    \new_[99631]_ , \new_[99632]_ , \new_[99633]_ , \new_[99636]_ ,
    \new_[99639]_ , \new_[99640]_ , \new_[99643]_ , \new_[99646]_ ,
    \new_[99647]_ , \new_[99648]_ , \new_[99651]_ , \new_[99654]_ ,
    \new_[99655]_ , \new_[99658]_ , \new_[99661]_ , \new_[99662]_ ,
    \new_[99663]_ , \new_[99666]_ , \new_[99669]_ , \new_[99670]_ ,
    \new_[99673]_ , \new_[99676]_ , \new_[99677]_ , \new_[99678]_ ,
    \new_[99681]_ , \new_[99684]_ , \new_[99685]_ , \new_[99688]_ ,
    \new_[99691]_ , \new_[99692]_ , \new_[99693]_ , \new_[99696]_ ,
    \new_[99699]_ , \new_[99700]_ , \new_[99703]_ , \new_[99706]_ ,
    \new_[99707]_ , \new_[99708]_ , \new_[99711]_ , \new_[99714]_ ,
    \new_[99715]_ , \new_[99718]_ , \new_[99721]_ , \new_[99722]_ ,
    \new_[99723]_ , \new_[99726]_ , \new_[99729]_ , \new_[99730]_ ,
    \new_[99733]_ , \new_[99736]_ , \new_[99737]_ , \new_[99738]_ ,
    \new_[99741]_ , \new_[99744]_ , \new_[99745]_ , \new_[99748]_ ,
    \new_[99751]_ , \new_[99752]_ , \new_[99753]_ , \new_[99756]_ ,
    \new_[99759]_ , \new_[99760]_ , \new_[99763]_ , \new_[99766]_ ,
    \new_[99767]_ , \new_[99768]_ , \new_[99771]_ , \new_[99774]_ ,
    \new_[99775]_ , \new_[99778]_ , \new_[99781]_ , \new_[99782]_ ,
    \new_[99783]_ , \new_[99786]_ , \new_[99789]_ , \new_[99790]_ ,
    \new_[99793]_ , \new_[99796]_ , \new_[99797]_ , \new_[99798]_ ,
    \new_[99801]_ , \new_[99804]_ , \new_[99805]_ , \new_[99808]_ ,
    \new_[99811]_ , \new_[99812]_ , \new_[99813]_ , \new_[99816]_ ,
    \new_[99819]_ , \new_[99820]_ , \new_[99823]_ , \new_[99826]_ ,
    \new_[99827]_ , \new_[99828]_ , \new_[99831]_ , \new_[99834]_ ,
    \new_[99835]_ , \new_[99838]_ , \new_[99841]_ , \new_[99842]_ ,
    \new_[99843]_ , \new_[99846]_ , \new_[99849]_ , \new_[99850]_ ,
    \new_[99853]_ , \new_[99856]_ , \new_[99857]_ , \new_[99858]_ ,
    \new_[99861]_ , \new_[99864]_ , \new_[99865]_ , \new_[99868]_ ,
    \new_[99871]_ , \new_[99872]_ , \new_[99873]_ , \new_[99876]_ ,
    \new_[99879]_ , \new_[99880]_ , \new_[99883]_ , \new_[99886]_ ,
    \new_[99887]_ , \new_[99888]_ , \new_[99891]_ , \new_[99894]_ ,
    \new_[99895]_ , \new_[99898]_ , \new_[99901]_ , \new_[99902]_ ,
    \new_[99903]_ , \new_[99906]_ , \new_[99909]_ , \new_[99910]_ ,
    \new_[99913]_ , \new_[99916]_ , \new_[99917]_ , \new_[99918]_ ,
    \new_[99921]_ , \new_[99924]_ , \new_[99925]_ , \new_[99928]_ ,
    \new_[99931]_ , \new_[99932]_ , \new_[99933]_ , \new_[99936]_ ,
    \new_[99939]_ , \new_[99940]_ , \new_[99943]_ , \new_[99946]_ ,
    \new_[99947]_ , \new_[99948]_ , \new_[99951]_ , \new_[99954]_ ,
    \new_[99955]_ , \new_[99958]_ , \new_[99961]_ , \new_[99962]_ ,
    \new_[99963]_ , \new_[99966]_ , \new_[99969]_ , \new_[99970]_ ,
    \new_[99973]_ , \new_[99976]_ , \new_[99977]_ , \new_[99978]_ ,
    \new_[99981]_ , \new_[99984]_ , \new_[99985]_ , \new_[99988]_ ,
    \new_[99991]_ , \new_[99992]_ , \new_[99993]_ , \new_[99996]_ ,
    \new_[99999]_ , \new_[100000]_ , \new_[100003]_ , \new_[100006]_ ,
    \new_[100007]_ , \new_[100008]_ , \new_[100011]_ , \new_[100014]_ ,
    \new_[100015]_ , \new_[100018]_ , \new_[100021]_ , \new_[100022]_ ,
    \new_[100023]_ , \new_[100026]_ , \new_[100029]_ , \new_[100030]_ ,
    \new_[100033]_ , \new_[100036]_ , \new_[100037]_ , \new_[100038]_ ,
    \new_[100041]_ , \new_[100044]_ , \new_[100045]_ , \new_[100048]_ ,
    \new_[100051]_ , \new_[100052]_ , \new_[100053]_ , \new_[100056]_ ,
    \new_[100059]_ , \new_[100060]_ , \new_[100063]_ , \new_[100066]_ ,
    \new_[100067]_ , \new_[100068]_ , \new_[100071]_ , \new_[100074]_ ,
    \new_[100075]_ , \new_[100078]_ , \new_[100081]_ , \new_[100082]_ ,
    \new_[100083]_ , \new_[100086]_ , \new_[100089]_ , \new_[100090]_ ,
    \new_[100093]_ , \new_[100096]_ , \new_[100097]_ , \new_[100098]_ ,
    \new_[100101]_ , \new_[100104]_ , \new_[100105]_ , \new_[100108]_ ,
    \new_[100111]_ , \new_[100112]_ , \new_[100113]_ , \new_[100116]_ ,
    \new_[100119]_ , \new_[100120]_ , \new_[100123]_ , \new_[100126]_ ,
    \new_[100127]_ , \new_[100128]_ , \new_[100131]_ , \new_[100134]_ ,
    \new_[100135]_ , \new_[100138]_ , \new_[100141]_ , \new_[100142]_ ,
    \new_[100143]_ , \new_[100146]_ , \new_[100149]_ , \new_[100150]_ ,
    \new_[100153]_ , \new_[100156]_ , \new_[100157]_ , \new_[100158]_ ,
    \new_[100161]_ , \new_[100164]_ , \new_[100165]_ , \new_[100168]_ ,
    \new_[100171]_ , \new_[100172]_ , \new_[100173]_ , \new_[100176]_ ,
    \new_[100179]_ , \new_[100180]_ , \new_[100183]_ , \new_[100186]_ ,
    \new_[100187]_ , \new_[100188]_ , \new_[100191]_ , \new_[100194]_ ,
    \new_[100195]_ , \new_[100198]_ , \new_[100201]_ , \new_[100202]_ ,
    \new_[100203]_ , \new_[100206]_ , \new_[100209]_ , \new_[100210]_ ,
    \new_[100213]_ , \new_[100216]_ , \new_[100217]_ , \new_[100218]_ ,
    \new_[100221]_ , \new_[100224]_ , \new_[100225]_ , \new_[100228]_ ,
    \new_[100231]_ , \new_[100232]_ , \new_[100233]_ , \new_[100236]_ ,
    \new_[100239]_ , \new_[100240]_ , \new_[100243]_ , \new_[100246]_ ,
    \new_[100247]_ , \new_[100248]_ , \new_[100251]_ , \new_[100254]_ ,
    \new_[100255]_ , \new_[100258]_ , \new_[100261]_ , \new_[100262]_ ,
    \new_[100263]_ , \new_[100266]_ , \new_[100269]_ , \new_[100270]_ ,
    \new_[100273]_ , \new_[100276]_ , \new_[100277]_ , \new_[100278]_ ,
    \new_[100281]_ , \new_[100284]_ , \new_[100285]_ , \new_[100288]_ ,
    \new_[100291]_ , \new_[100292]_ , \new_[100293]_ , \new_[100296]_ ,
    \new_[100299]_ , \new_[100300]_ , \new_[100303]_ , \new_[100306]_ ,
    \new_[100307]_ , \new_[100308]_ , \new_[100311]_ , \new_[100314]_ ,
    \new_[100315]_ , \new_[100318]_ , \new_[100321]_ , \new_[100322]_ ,
    \new_[100323]_ , \new_[100326]_ , \new_[100329]_ , \new_[100330]_ ,
    \new_[100333]_ , \new_[100336]_ , \new_[100337]_ , \new_[100338]_ ,
    \new_[100341]_ , \new_[100344]_ , \new_[100345]_ , \new_[100348]_ ,
    \new_[100351]_ , \new_[100352]_ , \new_[100353]_ , \new_[100356]_ ,
    \new_[100359]_ , \new_[100360]_ , \new_[100363]_ , \new_[100366]_ ,
    \new_[100367]_ , \new_[100368]_ , \new_[100371]_ , \new_[100374]_ ,
    \new_[100375]_ , \new_[100378]_ , \new_[100381]_ , \new_[100382]_ ,
    \new_[100383]_ , \new_[100386]_ , \new_[100389]_ , \new_[100390]_ ,
    \new_[100393]_ , \new_[100396]_ , \new_[100397]_ , \new_[100398]_ ,
    \new_[100401]_ , \new_[100404]_ , \new_[100405]_ , \new_[100408]_ ,
    \new_[100411]_ , \new_[100412]_ , \new_[100413]_ , \new_[100416]_ ,
    \new_[100419]_ , \new_[100420]_ , \new_[100423]_ , \new_[100426]_ ,
    \new_[100427]_ , \new_[100428]_ , \new_[100431]_ , \new_[100434]_ ,
    \new_[100435]_ , \new_[100438]_ , \new_[100441]_ , \new_[100442]_ ,
    \new_[100443]_ , \new_[100446]_ , \new_[100449]_ , \new_[100450]_ ,
    \new_[100453]_ , \new_[100456]_ , \new_[100457]_ , \new_[100458]_ ,
    \new_[100461]_ , \new_[100464]_ , \new_[100465]_ , \new_[100468]_ ,
    \new_[100471]_ , \new_[100472]_ , \new_[100473]_ , \new_[100476]_ ,
    \new_[100479]_ , \new_[100480]_ , \new_[100483]_ , \new_[100486]_ ,
    \new_[100487]_ , \new_[100488]_ , \new_[100491]_ , \new_[100494]_ ,
    \new_[100495]_ , \new_[100498]_ , \new_[100501]_ , \new_[100502]_ ,
    \new_[100503]_ , \new_[100506]_ , \new_[100509]_ , \new_[100510]_ ,
    \new_[100513]_ , \new_[100516]_ , \new_[100517]_ , \new_[100518]_ ,
    \new_[100521]_ , \new_[100524]_ , \new_[100525]_ , \new_[100528]_ ,
    \new_[100531]_ , \new_[100532]_ , \new_[100533]_ , \new_[100536]_ ,
    \new_[100539]_ , \new_[100540]_ , \new_[100543]_ , \new_[100546]_ ,
    \new_[100547]_ , \new_[100548]_ , \new_[100551]_ , \new_[100554]_ ,
    \new_[100555]_ , \new_[100558]_ , \new_[100561]_ , \new_[100562]_ ,
    \new_[100563]_ , \new_[100566]_ , \new_[100569]_ , \new_[100570]_ ,
    \new_[100573]_ , \new_[100576]_ , \new_[100577]_ , \new_[100578]_ ,
    \new_[100581]_ , \new_[100584]_ , \new_[100585]_ , \new_[100588]_ ,
    \new_[100591]_ , \new_[100592]_ , \new_[100593]_ , \new_[100596]_ ,
    \new_[100599]_ , \new_[100600]_ , \new_[100603]_ , \new_[100606]_ ,
    \new_[100607]_ , \new_[100608]_ , \new_[100611]_ , \new_[100614]_ ,
    \new_[100615]_ , \new_[100618]_ , \new_[100621]_ , \new_[100622]_ ,
    \new_[100623]_ , \new_[100626]_ , \new_[100629]_ , \new_[100630]_ ,
    \new_[100633]_ , \new_[100636]_ , \new_[100637]_ , \new_[100638]_ ,
    \new_[100641]_ , \new_[100644]_ , \new_[100645]_ , \new_[100648]_ ,
    \new_[100651]_ , \new_[100652]_ , \new_[100653]_ , \new_[100656]_ ,
    \new_[100659]_ , \new_[100660]_ , \new_[100663]_ , \new_[100666]_ ,
    \new_[100667]_ , \new_[100668]_ , \new_[100671]_ , \new_[100674]_ ,
    \new_[100675]_ , \new_[100678]_ , \new_[100681]_ , \new_[100682]_ ,
    \new_[100683]_ , \new_[100686]_ , \new_[100689]_ , \new_[100690]_ ,
    \new_[100693]_ , \new_[100696]_ , \new_[100697]_ , \new_[100698]_ ,
    \new_[100701]_ , \new_[100704]_ , \new_[100705]_ , \new_[100708]_ ,
    \new_[100711]_ , \new_[100712]_ , \new_[100713]_ , \new_[100716]_ ,
    \new_[100719]_ , \new_[100720]_ , \new_[100723]_ , \new_[100726]_ ,
    \new_[100727]_ , \new_[100728]_ , \new_[100731]_ , \new_[100734]_ ,
    \new_[100735]_ , \new_[100738]_ , \new_[100741]_ , \new_[100742]_ ,
    \new_[100743]_ , \new_[100746]_ , \new_[100749]_ , \new_[100750]_ ,
    \new_[100753]_ , \new_[100756]_ , \new_[100757]_ , \new_[100758]_ ,
    \new_[100761]_ , \new_[100764]_ , \new_[100765]_ , \new_[100768]_ ,
    \new_[100771]_ , \new_[100772]_ , \new_[100773]_ , \new_[100776]_ ,
    \new_[100779]_ , \new_[100780]_ , \new_[100783]_ , \new_[100786]_ ,
    \new_[100787]_ , \new_[100788]_ , \new_[100791]_ , \new_[100794]_ ,
    \new_[100795]_ , \new_[100798]_ , \new_[100801]_ , \new_[100802]_ ,
    \new_[100803]_ , \new_[100806]_ , \new_[100809]_ , \new_[100810]_ ,
    \new_[100813]_ , \new_[100816]_ , \new_[100817]_ , \new_[100818]_ ,
    \new_[100821]_ , \new_[100824]_ , \new_[100825]_ , \new_[100828]_ ,
    \new_[100831]_ , \new_[100832]_ , \new_[100833]_ , \new_[100836]_ ,
    \new_[100839]_ , \new_[100840]_ , \new_[100843]_ , \new_[100846]_ ,
    \new_[100847]_ , \new_[100848]_ , \new_[100851]_ , \new_[100854]_ ,
    \new_[100855]_ , \new_[100858]_ , \new_[100861]_ , \new_[100862]_ ,
    \new_[100863]_ , \new_[100866]_ , \new_[100869]_ , \new_[100870]_ ,
    \new_[100873]_ , \new_[100876]_ , \new_[100877]_ , \new_[100878]_ ,
    \new_[100881]_ , \new_[100884]_ , \new_[100885]_ , \new_[100888]_ ,
    \new_[100891]_ , \new_[100892]_ , \new_[100893]_ , \new_[100896]_ ,
    \new_[100899]_ , \new_[100900]_ , \new_[100903]_ , \new_[100906]_ ,
    \new_[100907]_ , \new_[100908]_ , \new_[100911]_ , \new_[100914]_ ,
    \new_[100915]_ , \new_[100918]_ , \new_[100921]_ , \new_[100922]_ ,
    \new_[100923]_ , \new_[100926]_ , \new_[100929]_ , \new_[100930]_ ,
    \new_[100933]_ , \new_[100936]_ , \new_[100937]_ , \new_[100938]_ ,
    \new_[100941]_ , \new_[100944]_ , \new_[100945]_ , \new_[100948]_ ,
    \new_[100951]_ , \new_[100952]_ , \new_[100953]_ , \new_[100956]_ ,
    \new_[100959]_ , \new_[100960]_ , \new_[100963]_ , \new_[100966]_ ,
    \new_[100967]_ , \new_[100968]_ , \new_[100971]_ , \new_[100974]_ ,
    \new_[100975]_ , \new_[100978]_ , \new_[100981]_ , \new_[100982]_ ,
    \new_[100983]_ , \new_[100986]_ , \new_[100989]_ , \new_[100990]_ ,
    \new_[100993]_ , \new_[100996]_ , \new_[100997]_ , \new_[100998]_ ,
    \new_[101001]_ , \new_[101004]_ , \new_[101005]_ , \new_[101008]_ ,
    \new_[101011]_ , \new_[101012]_ , \new_[101013]_ , \new_[101016]_ ,
    \new_[101019]_ , \new_[101020]_ , \new_[101023]_ , \new_[101026]_ ,
    \new_[101027]_ , \new_[101028]_ , \new_[101031]_ , \new_[101034]_ ,
    \new_[101035]_ , \new_[101038]_ , \new_[101041]_ , \new_[101042]_ ,
    \new_[101043]_ , \new_[101046]_ , \new_[101049]_ , \new_[101050]_ ,
    \new_[101053]_ , \new_[101056]_ , \new_[101057]_ , \new_[101058]_ ,
    \new_[101061]_ , \new_[101064]_ , \new_[101065]_ , \new_[101068]_ ,
    \new_[101071]_ , \new_[101072]_ , \new_[101073]_ , \new_[101076]_ ,
    \new_[101079]_ , \new_[101080]_ , \new_[101083]_ , \new_[101086]_ ,
    \new_[101087]_ , \new_[101088]_ , \new_[101091]_ , \new_[101094]_ ,
    \new_[101095]_ , \new_[101098]_ , \new_[101101]_ , \new_[101102]_ ,
    \new_[101103]_ , \new_[101106]_ , \new_[101109]_ , \new_[101110]_ ,
    \new_[101113]_ , \new_[101116]_ , \new_[101117]_ , \new_[101118]_ ,
    \new_[101121]_ , \new_[101124]_ , \new_[101125]_ , \new_[101128]_ ,
    \new_[101131]_ , \new_[101132]_ , \new_[101133]_ , \new_[101136]_ ,
    \new_[101139]_ , \new_[101140]_ , \new_[101143]_ , \new_[101146]_ ,
    \new_[101147]_ , \new_[101148]_ , \new_[101151]_ , \new_[101154]_ ,
    \new_[101155]_ , \new_[101158]_ , \new_[101161]_ , \new_[101162]_ ,
    \new_[101163]_ , \new_[101166]_ , \new_[101169]_ , \new_[101170]_ ,
    \new_[101173]_ , \new_[101176]_ , \new_[101177]_ , \new_[101178]_ ,
    \new_[101181]_ , \new_[101184]_ , \new_[101185]_ , \new_[101188]_ ,
    \new_[101191]_ , \new_[101192]_ , \new_[101193]_ , \new_[101196]_ ,
    \new_[101199]_ , \new_[101200]_ , \new_[101203]_ , \new_[101206]_ ,
    \new_[101207]_ , \new_[101208]_ , \new_[101211]_ , \new_[101214]_ ,
    \new_[101215]_ , \new_[101218]_ , \new_[101221]_ , \new_[101222]_ ,
    \new_[101223]_ , \new_[101226]_ , \new_[101229]_ , \new_[101230]_ ,
    \new_[101233]_ , \new_[101236]_ , \new_[101237]_ , \new_[101238]_ ,
    \new_[101241]_ , \new_[101244]_ , \new_[101245]_ , \new_[101248]_ ,
    \new_[101251]_ , \new_[101252]_ , \new_[101253]_ , \new_[101256]_ ,
    \new_[101259]_ , \new_[101260]_ , \new_[101263]_ , \new_[101266]_ ,
    \new_[101267]_ , \new_[101268]_ , \new_[101271]_ , \new_[101274]_ ,
    \new_[101275]_ , \new_[101278]_ , \new_[101281]_ , \new_[101282]_ ,
    \new_[101283]_ , \new_[101286]_ , \new_[101289]_ , \new_[101290]_ ,
    \new_[101293]_ , \new_[101296]_ , \new_[101297]_ , \new_[101298]_ ,
    \new_[101301]_ , \new_[101304]_ , \new_[101305]_ , \new_[101308]_ ,
    \new_[101311]_ , \new_[101312]_ , \new_[101313]_ , \new_[101316]_ ,
    \new_[101319]_ , \new_[101320]_ , \new_[101323]_ , \new_[101326]_ ,
    \new_[101327]_ , \new_[101328]_ , \new_[101331]_ , \new_[101334]_ ,
    \new_[101335]_ , \new_[101338]_ , \new_[101341]_ , \new_[101342]_ ,
    \new_[101343]_ , \new_[101346]_ , \new_[101349]_ , \new_[101350]_ ,
    \new_[101353]_ , \new_[101356]_ , \new_[101357]_ , \new_[101358]_ ,
    \new_[101361]_ , \new_[101364]_ , \new_[101365]_ , \new_[101368]_ ,
    \new_[101371]_ , \new_[101372]_ , \new_[101373]_ , \new_[101376]_ ,
    \new_[101379]_ , \new_[101380]_ , \new_[101383]_ , \new_[101386]_ ,
    \new_[101387]_ , \new_[101388]_ , \new_[101391]_ , \new_[101394]_ ,
    \new_[101395]_ , \new_[101398]_ , \new_[101401]_ , \new_[101402]_ ,
    \new_[101403]_ , \new_[101406]_ , \new_[101409]_ , \new_[101410]_ ,
    \new_[101413]_ , \new_[101416]_ , \new_[101417]_ , \new_[101418]_ ,
    \new_[101421]_ , \new_[101424]_ , \new_[101425]_ , \new_[101428]_ ,
    \new_[101431]_ , \new_[101432]_ , \new_[101433]_ , \new_[101436]_ ,
    \new_[101439]_ , \new_[101440]_ , \new_[101443]_ , \new_[101446]_ ,
    \new_[101447]_ , \new_[101448]_ , \new_[101451]_ , \new_[101454]_ ,
    \new_[101455]_ , \new_[101458]_ , \new_[101461]_ , \new_[101462]_ ,
    \new_[101463]_ , \new_[101466]_ , \new_[101469]_ , \new_[101470]_ ,
    \new_[101473]_ , \new_[101476]_ , \new_[101477]_ , \new_[101478]_ ,
    \new_[101481]_ , \new_[101484]_ , \new_[101485]_ , \new_[101488]_ ,
    \new_[101491]_ , \new_[101492]_ , \new_[101493]_ , \new_[101496]_ ,
    \new_[101499]_ , \new_[101500]_ , \new_[101503]_ , \new_[101506]_ ,
    \new_[101507]_ , \new_[101508]_ , \new_[101511]_ , \new_[101514]_ ,
    \new_[101515]_ , \new_[101518]_ , \new_[101521]_ , \new_[101522]_ ,
    \new_[101523]_ , \new_[101526]_ , \new_[101529]_ , \new_[101530]_ ,
    \new_[101533]_ , \new_[101536]_ , \new_[101537]_ , \new_[101538]_ ,
    \new_[101541]_ , \new_[101544]_ , \new_[101545]_ , \new_[101548]_ ,
    \new_[101551]_ , \new_[101552]_ , \new_[101553]_ , \new_[101556]_ ,
    \new_[101559]_ , \new_[101560]_ , \new_[101563]_ , \new_[101566]_ ,
    \new_[101567]_ , \new_[101568]_ , \new_[101571]_ , \new_[101574]_ ,
    \new_[101575]_ , \new_[101578]_ , \new_[101581]_ , \new_[101582]_ ,
    \new_[101583]_ , \new_[101586]_ , \new_[101589]_ , \new_[101590]_ ,
    \new_[101593]_ , \new_[101596]_ , \new_[101597]_ , \new_[101598]_ ,
    \new_[101601]_ , \new_[101604]_ , \new_[101605]_ , \new_[101608]_ ,
    \new_[101611]_ , \new_[101612]_ , \new_[101613]_ , \new_[101616]_ ,
    \new_[101619]_ , \new_[101620]_ , \new_[101623]_ , \new_[101626]_ ,
    \new_[101627]_ , \new_[101628]_ , \new_[101631]_ , \new_[101634]_ ,
    \new_[101635]_ , \new_[101638]_ , \new_[101641]_ , \new_[101642]_ ,
    \new_[101643]_ , \new_[101646]_ , \new_[101649]_ , \new_[101650]_ ,
    \new_[101653]_ , \new_[101656]_ , \new_[101657]_ , \new_[101658]_ ,
    \new_[101661]_ , \new_[101664]_ , \new_[101665]_ , \new_[101668]_ ,
    \new_[101671]_ , \new_[101672]_ , \new_[101673]_ , \new_[101676]_ ,
    \new_[101679]_ , \new_[101680]_ , \new_[101683]_ , \new_[101686]_ ,
    \new_[101687]_ , \new_[101688]_ , \new_[101691]_ , \new_[101694]_ ,
    \new_[101695]_ , \new_[101698]_ , \new_[101701]_ , \new_[101702]_ ,
    \new_[101703]_ , \new_[101706]_ , \new_[101709]_ , \new_[101710]_ ,
    \new_[101713]_ , \new_[101716]_ , \new_[101717]_ , \new_[101718]_ ,
    \new_[101721]_ , \new_[101724]_ , \new_[101725]_ , \new_[101728]_ ,
    \new_[101731]_ , \new_[101732]_ , \new_[101733]_ , \new_[101736]_ ,
    \new_[101739]_ , \new_[101740]_ , \new_[101743]_ , \new_[101746]_ ,
    \new_[101747]_ , \new_[101748]_ , \new_[101751]_ , \new_[101754]_ ,
    \new_[101755]_ , \new_[101758]_ , \new_[101761]_ , \new_[101762]_ ,
    \new_[101763]_ , \new_[101766]_ , \new_[101769]_ , \new_[101770]_ ,
    \new_[101773]_ , \new_[101777]_ , \new_[101778]_ , \new_[101779]_ ,
    \new_[101780]_ , \new_[101783]_ , \new_[101786]_ , \new_[101787]_ ,
    \new_[101790]_ , \new_[101793]_ , \new_[101794]_ , \new_[101795]_ ,
    \new_[101798]_ , \new_[101801]_ , \new_[101802]_ , \new_[101805]_ ,
    \new_[101809]_ , \new_[101810]_ , \new_[101811]_ , \new_[101812]_ ,
    \new_[101815]_ , \new_[101818]_ , \new_[101819]_ , \new_[101822]_ ,
    \new_[101825]_ , \new_[101826]_ , \new_[101827]_ , \new_[101830]_ ,
    \new_[101833]_ , \new_[101834]_ , \new_[101837]_ , \new_[101841]_ ,
    \new_[101842]_ , \new_[101843]_ , \new_[101844]_ , \new_[101847]_ ,
    \new_[101850]_ , \new_[101851]_ , \new_[101854]_ , \new_[101857]_ ,
    \new_[101858]_ , \new_[101859]_ , \new_[101862]_ , \new_[101865]_ ,
    \new_[101866]_ , \new_[101869]_ , \new_[101873]_ , \new_[101874]_ ,
    \new_[101875]_ , \new_[101876]_ , \new_[101879]_ , \new_[101882]_ ,
    \new_[101883]_ , \new_[101886]_ , \new_[101889]_ , \new_[101890]_ ,
    \new_[101891]_ , \new_[101894]_ , \new_[101897]_ , \new_[101898]_ ,
    \new_[101901]_ , \new_[101905]_ , \new_[101906]_ , \new_[101907]_ ,
    \new_[101908]_ , \new_[101911]_ , \new_[101914]_ , \new_[101915]_ ,
    \new_[101918]_ , \new_[101921]_ , \new_[101922]_ , \new_[101923]_ ,
    \new_[101926]_ , \new_[101929]_ , \new_[101930]_ , \new_[101933]_ ,
    \new_[101937]_ , \new_[101938]_ , \new_[101939]_ , \new_[101940]_ ,
    \new_[101943]_ , \new_[101946]_ , \new_[101947]_ , \new_[101950]_ ,
    \new_[101953]_ , \new_[101954]_ , \new_[101955]_ , \new_[101958]_ ,
    \new_[101961]_ , \new_[101962]_ , \new_[101965]_ , \new_[101969]_ ,
    \new_[101970]_ , \new_[101971]_ , \new_[101972]_ , \new_[101975]_ ,
    \new_[101978]_ , \new_[101979]_ , \new_[101982]_ , \new_[101985]_ ,
    \new_[101986]_ , \new_[101987]_ , \new_[101990]_ , \new_[101993]_ ,
    \new_[101994]_ , \new_[101997]_ , \new_[102001]_ , \new_[102002]_ ,
    \new_[102003]_ , \new_[102004]_ , \new_[102007]_ , \new_[102010]_ ,
    \new_[102011]_ , \new_[102014]_ , \new_[102017]_ , \new_[102018]_ ,
    \new_[102019]_ , \new_[102022]_ , \new_[102025]_ , \new_[102026]_ ,
    \new_[102029]_ , \new_[102033]_ , \new_[102034]_ , \new_[102035]_ ,
    \new_[102036]_ , \new_[102039]_ , \new_[102042]_ , \new_[102043]_ ,
    \new_[102046]_ , \new_[102049]_ , \new_[102050]_ , \new_[102051]_ ,
    \new_[102054]_ , \new_[102057]_ , \new_[102058]_ , \new_[102061]_ ,
    \new_[102065]_ , \new_[102066]_ , \new_[102067]_ , \new_[102068]_ ,
    \new_[102071]_ , \new_[102074]_ , \new_[102075]_ , \new_[102078]_ ,
    \new_[102081]_ , \new_[102082]_ , \new_[102083]_ , \new_[102086]_ ,
    \new_[102089]_ , \new_[102090]_ , \new_[102093]_ , \new_[102097]_ ,
    \new_[102098]_ , \new_[102099]_ , \new_[102100]_ , \new_[102103]_ ,
    \new_[102106]_ , \new_[102107]_ , \new_[102110]_ , \new_[102113]_ ,
    \new_[102114]_ , \new_[102115]_ , \new_[102118]_ , \new_[102121]_ ,
    \new_[102122]_ , \new_[102125]_ , \new_[102129]_ , \new_[102130]_ ,
    \new_[102131]_ , \new_[102132]_ , \new_[102135]_ , \new_[102138]_ ,
    \new_[102139]_ , \new_[102142]_ , \new_[102145]_ , \new_[102146]_ ,
    \new_[102147]_ , \new_[102150]_ , \new_[102153]_ , \new_[102154]_ ,
    \new_[102157]_ , \new_[102161]_ , \new_[102162]_ , \new_[102163]_ ,
    \new_[102164]_ , \new_[102167]_ , \new_[102170]_ , \new_[102171]_ ,
    \new_[102174]_ , \new_[102177]_ , \new_[102178]_ , \new_[102179]_ ,
    \new_[102182]_ , \new_[102185]_ , \new_[102186]_ , \new_[102189]_ ,
    \new_[102193]_ , \new_[102194]_ , \new_[102195]_ , \new_[102196]_ ,
    \new_[102199]_ , \new_[102202]_ , \new_[102203]_ , \new_[102206]_ ,
    \new_[102209]_ , \new_[102210]_ , \new_[102211]_ , \new_[102214]_ ,
    \new_[102217]_ , \new_[102218]_ , \new_[102221]_ , \new_[102225]_ ,
    \new_[102226]_ , \new_[102227]_ , \new_[102228]_ , \new_[102231]_ ,
    \new_[102234]_ , \new_[102235]_ , \new_[102238]_ , \new_[102241]_ ,
    \new_[102242]_ , \new_[102243]_ , \new_[102246]_ , \new_[102249]_ ,
    \new_[102250]_ , \new_[102253]_ , \new_[102257]_ , \new_[102258]_ ,
    \new_[102259]_ , \new_[102260]_ , \new_[102263]_ , \new_[102266]_ ,
    \new_[102267]_ , \new_[102270]_ , \new_[102273]_ , \new_[102274]_ ,
    \new_[102275]_ , \new_[102278]_ , \new_[102281]_ , \new_[102282]_ ,
    \new_[102285]_ , \new_[102289]_ , \new_[102290]_ , \new_[102291]_ ,
    \new_[102292]_ , \new_[102295]_ , \new_[102298]_ , \new_[102299]_ ,
    \new_[102302]_ , \new_[102305]_ , \new_[102306]_ , \new_[102307]_ ,
    \new_[102310]_ , \new_[102313]_ , \new_[102314]_ , \new_[102317]_ ,
    \new_[102321]_ , \new_[102322]_ , \new_[102323]_ , \new_[102324]_ ,
    \new_[102327]_ , \new_[102330]_ , \new_[102331]_ , \new_[102334]_ ,
    \new_[102337]_ , \new_[102338]_ , \new_[102339]_ , \new_[102342]_ ,
    \new_[102345]_ , \new_[102346]_ , \new_[102349]_ , \new_[102353]_ ,
    \new_[102354]_ , \new_[102355]_ , \new_[102356]_ , \new_[102359]_ ,
    \new_[102362]_ , \new_[102363]_ , \new_[102366]_ , \new_[102369]_ ,
    \new_[102370]_ , \new_[102371]_ , \new_[102374]_ , \new_[102377]_ ,
    \new_[102378]_ , \new_[102381]_ , \new_[102385]_ , \new_[102386]_ ,
    \new_[102387]_ , \new_[102388]_ , \new_[102391]_ , \new_[102394]_ ,
    \new_[102395]_ , \new_[102398]_ , \new_[102401]_ , \new_[102402]_ ,
    \new_[102403]_ , \new_[102406]_ , \new_[102409]_ , \new_[102410]_ ,
    \new_[102413]_ , \new_[102417]_ , \new_[102418]_ , \new_[102419]_ ,
    \new_[102420]_ , \new_[102423]_ , \new_[102426]_ , \new_[102427]_ ,
    \new_[102430]_ , \new_[102433]_ , \new_[102434]_ , \new_[102435]_ ,
    \new_[102438]_ , \new_[102441]_ , \new_[102442]_ , \new_[102445]_ ,
    \new_[102449]_ , \new_[102450]_ , \new_[102451]_ , \new_[102452]_ ,
    \new_[102455]_ , \new_[102458]_ , \new_[102459]_ , \new_[102462]_ ,
    \new_[102465]_ , \new_[102466]_ , \new_[102467]_ , \new_[102470]_ ,
    \new_[102473]_ , \new_[102474]_ , \new_[102477]_ , \new_[102481]_ ,
    \new_[102482]_ , \new_[102483]_ , \new_[102484]_ , \new_[102487]_ ,
    \new_[102490]_ , \new_[102491]_ , \new_[102494]_ , \new_[102497]_ ,
    \new_[102498]_ , \new_[102499]_ , \new_[102502]_ , \new_[102505]_ ,
    \new_[102506]_ , \new_[102509]_ , \new_[102513]_ , \new_[102514]_ ,
    \new_[102515]_ , \new_[102516]_ , \new_[102519]_ , \new_[102522]_ ,
    \new_[102523]_ , \new_[102526]_ , \new_[102529]_ , \new_[102530]_ ,
    \new_[102531]_ , \new_[102534]_ , \new_[102537]_ , \new_[102538]_ ,
    \new_[102541]_ , \new_[102545]_ , \new_[102546]_ , \new_[102547]_ ,
    \new_[102548]_ , \new_[102551]_ , \new_[102554]_ , \new_[102555]_ ,
    \new_[102558]_ , \new_[102561]_ , \new_[102562]_ , \new_[102563]_ ,
    \new_[102566]_ , \new_[102569]_ , \new_[102570]_ , \new_[102573]_ ,
    \new_[102577]_ , \new_[102578]_ , \new_[102579]_ , \new_[102580]_ ,
    \new_[102583]_ , \new_[102586]_ , \new_[102587]_ , \new_[102590]_ ,
    \new_[102593]_ , \new_[102594]_ , \new_[102595]_ , \new_[102598]_ ,
    \new_[102601]_ , \new_[102602]_ , \new_[102605]_ , \new_[102609]_ ,
    \new_[102610]_ , \new_[102611]_ , \new_[102612]_ , \new_[102615]_ ,
    \new_[102618]_ , \new_[102619]_ , \new_[102622]_ , \new_[102625]_ ,
    \new_[102626]_ , \new_[102627]_ , \new_[102630]_ , \new_[102633]_ ,
    \new_[102634]_ , \new_[102637]_ , \new_[102641]_ , \new_[102642]_ ,
    \new_[102643]_ , \new_[102644]_ , \new_[102647]_ , \new_[102650]_ ,
    \new_[102651]_ , \new_[102654]_ , \new_[102657]_ , \new_[102658]_ ,
    \new_[102659]_ , \new_[102662]_ , \new_[102665]_ , \new_[102666]_ ,
    \new_[102669]_ , \new_[102673]_ , \new_[102674]_ , \new_[102675]_ ,
    \new_[102676]_ , \new_[102679]_ , \new_[102682]_ , \new_[102683]_ ,
    \new_[102686]_ , \new_[102689]_ , \new_[102690]_ , \new_[102691]_ ,
    \new_[102694]_ , \new_[102697]_ , \new_[102698]_ , \new_[102701]_ ,
    \new_[102705]_ , \new_[102706]_ , \new_[102707]_ , \new_[102708]_ ,
    \new_[102711]_ , \new_[102714]_ , \new_[102715]_ , \new_[102718]_ ,
    \new_[102721]_ , \new_[102722]_ , \new_[102723]_ , \new_[102726]_ ,
    \new_[102729]_ , \new_[102730]_ , \new_[102733]_ , \new_[102737]_ ,
    \new_[102738]_ , \new_[102739]_ , \new_[102740]_ , \new_[102743]_ ,
    \new_[102746]_ , \new_[102747]_ , \new_[102750]_ , \new_[102753]_ ,
    \new_[102754]_ , \new_[102755]_ , \new_[102758]_ , \new_[102761]_ ,
    \new_[102762]_ , \new_[102765]_ , \new_[102769]_ , \new_[102770]_ ,
    \new_[102771]_ , \new_[102772]_ , \new_[102775]_ , \new_[102778]_ ,
    \new_[102779]_ , \new_[102782]_ , \new_[102785]_ , \new_[102786]_ ,
    \new_[102787]_ , \new_[102790]_ , \new_[102793]_ , \new_[102794]_ ,
    \new_[102797]_ , \new_[102801]_ , \new_[102802]_ , \new_[102803]_ ,
    \new_[102804]_ , \new_[102807]_ , \new_[102810]_ , \new_[102811]_ ,
    \new_[102814]_ , \new_[102817]_ , \new_[102818]_ , \new_[102819]_ ,
    \new_[102822]_ , \new_[102825]_ , \new_[102826]_ , \new_[102829]_ ,
    \new_[102833]_ , \new_[102834]_ , \new_[102835]_ , \new_[102836]_ ,
    \new_[102839]_ , \new_[102842]_ , \new_[102843]_ , \new_[102846]_ ,
    \new_[102849]_ , \new_[102850]_ , \new_[102851]_ , \new_[102854]_ ,
    \new_[102857]_ , \new_[102858]_ , \new_[102861]_ , \new_[102865]_ ,
    \new_[102866]_ , \new_[102867]_ , \new_[102868]_ , \new_[102871]_ ,
    \new_[102874]_ , \new_[102875]_ , \new_[102878]_ , \new_[102881]_ ,
    \new_[102882]_ , \new_[102883]_ , \new_[102886]_ , \new_[102889]_ ,
    \new_[102890]_ , \new_[102893]_ , \new_[102897]_ , \new_[102898]_ ,
    \new_[102899]_ , \new_[102900]_ , \new_[102903]_ , \new_[102906]_ ,
    \new_[102907]_ , \new_[102910]_ , \new_[102913]_ , \new_[102914]_ ,
    \new_[102915]_ , \new_[102918]_ , \new_[102921]_ , \new_[102922]_ ,
    \new_[102925]_ , \new_[102929]_ , \new_[102930]_ , \new_[102931]_ ,
    \new_[102932]_ , \new_[102935]_ , \new_[102938]_ , \new_[102939]_ ,
    \new_[102942]_ , \new_[102945]_ , \new_[102946]_ , \new_[102947]_ ,
    \new_[102950]_ , \new_[102953]_ , \new_[102954]_ , \new_[102957]_ ,
    \new_[102961]_ , \new_[102962]_ , \new_[102963]_ , \new_[102964]_ ,
    \new_[102967]_ , \new_[102970]_ , \new_[102971]_ , \new_[102974]_ ,
    \new_[102977]_ , \new_[102978]_ , \new_[102979]_ , \new_[102982]_ ,
    \new_[102985]_ , \new_[102986]_ , \new_[102989]_ , \new_[102993]_ ,
    \new_[102994]_ , \new_[102995]_ , \new_[102996]_ , \new_[102999]_ ,
    \new_[103002]_ , \new_[103003]_ , \new_[103006]_ , \new_[103009]_ ,
    \new_[103010]_ , \new_[103011]_ , \new_[103014]_ , \new_[103017]_ ,
    \new_[103018]_ , \new_[103021]_ , \new_[103025]_ , \new_[103026]_ ,
    \new_[103027]_ , \new_[103028]_ , \new_[103031]_ , \new_[103034]_ ,
    \new_[103035]_ , \new_[103038]_ , \new_[103041]_ , \new_[103042]_ ,
    \new_[103043]_ , \new_[103046]_ , \new_[103049]_ , \new_[103050]_ ,
    \new_[103053]_ , \new_[103057]_ , \new_[103058]_ , \new_[103059]_ ,
    \new_[103060]_ , \new_[103063]_ , \new_[103066]_ , \new_[103067]_ ,
    \new_[103070]_ , \new_[103073]_ , \new_[103074]_ , \new_[103075]_ ,
    \new_[103078]_ , \new_[103081]_ , \new_[103082]_ , \new_[103085]_ ,
    \new_[103089]_ , \new_[103090]_ , \new_[103091]_ , \new_[103092]_ ,
    \new_[103095]_ , \new_[103098]_ , \new_[103099]_ , \new_[103102]_ ,
    \new_[103105]_ , \new_[103106]_ , \new_[103107]_ , \new_[103110]_ ,
    \new_[103113]_ , \new_[103114]_ , \new_[103117]_ , \new_[103121]_ ,
    \new_[103122]_ , \new_[103123]_ , \new_[103124]_ , \new_[103127]_ ,
    \new_[103130]_ , \new_[103131]_ , \new_[103134]_ , \new_[103137]_ ,
    \new_[103138]_ , \new_[103139]_ , \new_[103142]_ , \new_[103145]_ ,
    \new_[103146]_ , \new_[103149]_ , \new_[103153]_ , \new_[103154]_ ,
    \new_[103155]_ , \new_[103156]_ , \new_[103159]_ , \new_[103162]_ ,
    \new_[103163]_ , \new_[103166]_ , \new_[103169]_ , \new_[103170]_ ,
    \new_[103171]_ , \new_[103174]_ , \new_[103177]_ , \new_[103178]_ ,
    \new_[103181]_ , \new_[103185]_ , \new_[103186]_ , \new_[103187]_ ,
    \new_[103188]_ , \new_[103191]_ , \new_[103194]_ , \new_[103195]_ ,
    \new_[103198]_ , \new_[103201]_ , \new_[103202]_ , \new_[103203]_ ,
    \new_[103206]_ , \new_[103209]_ , \new_[103210]_ , \new_[103213]_ ,
    \new_[103217]_ , \new_[103218]_ , \new_[103219]_ , \new_[103220]_ ,
    \new_[103223]_ , \new_[103226]_ , \new_[103227]_ , \new_[103230]_ ,
    \new_[103233]_ , \new_[103234]_ , \new_[103235]_ , \new_[103238]_ ,
    \new_[103241]_ , \new_[103242]_ , \new_[103245]_ , \new_[103249]_ ,
    \new_[103250]_ , \new_[103251]_ , \new_[103252]_ , \new_[103255]_ ,
    \new_[103258]_ , \new_[103259]_ , \new_[103262]_ , \new_[103265]_ ,
    \new_[103266]_ , \new_[103267]_ , \new_[103270]_ , \new_[103273]_ ,
    \new_[103274]_ , \new_[103277]_ , \new_[103281]_ , \new_[103282]_ ,
    \new_[103283]_ , \new_[103284]_ , \new_[103287]_ , \new_[103290]_ ,
    \new_[103291]_ , \new_[103294]_ , \new_[103297]_ , \new_[103298]_ ,
    \new_[103299]_ , \new_[103302]_ , \new_[103305]_ , \new_[103306]_ ,
    \new_[103309]_ , \new_[103313]_ , \new_[103314]_ , \new_[103315]_ ,
    \new_[103316]_ , \new_[103319]_ , \new_[103322]_ , \new_[103323]_ ,
    \new_[103326]_ , \new_[103329]_ , \new_[103330]_ , \new_[103331]_ ,
    \new_[103334]_ , \new_[103337]_ , \new_[103338]_ , \new_[103341]_ ,
    \new_[103345]_ , \new_[103346]_ , \new_[103347]_ , \new_[103348]_ ,
    \new_[103351]_ , \new_[103354]_ , \new_[103355]_ , \new_[103358]_ ,
    \new_[103361]_ , \new_[103362]_ , \new_[103363]_ , \new_[103366]_ ,
    \new_[103369]_ , \new_[103370]_ , \new_[103373]_ , \new_[103377]_ ,
    \new_[103378]_ , \new_[103379]_ , \new_[103380]_ , \new_[103383]_ ,
    \new_[103386]_ , \new_[103387]_ , \new_[103390]_ , \new_[103393]_ ,
    \new_[103394]_ , \new_[103395]_ , \new_[103398]_ , \new_[103401]_ ,
    \new_[103402]_ , \new_[103405]_ , \new_[103409]_ , \new_[103410]_ ,
    \new_[103411]_ , \new_[103412]_ , \new_[103415]_ , \new_[103418]_ ,
    \new_[103419]_ , \new_[103422]_ , \new_[103425]_ , \new_[103426]_ ,
    \new_[103427]_ , \new_[103430]_ , \new_[103433]_ , \new_[103434]_ ,
    \new_[103437]_ , \new_[103441]_ , \new_[103442]_ , \new_[103443]_ ,
    \new_[103444]_ , \new_[103447]_ , \new_[103450]_ , \new_[103451]_ ,
    \new_[103454]_ , \new_[103457]_ , \new_[103458]_ , \new_[103459]_ ,
    \new_[103462]_ , \new_[103465]_ , \new_[103466]_ , \new_[103469]_ ,
    \new_[103473]_ , \new_[103474]_ , \new_[103475]_ , \new_[103476]_ ,
    \new_[103479]_ , \new_[103482]_ , \new_[103483]_ , \new_[103486]_ ,
    \new_[103489]_ , \new_[103490]_ , \new_[103491]_ , \new_[103494]_ ,
    \new_[103497]_ , \new_[103498]_ , \new_[103501]_ , \new_[103505]_ ,
    \new_[103506]_ , \new_[103507]_ , \new_[103508]_ , \new_[103511]_ ,
    \new_[103514]_ , \new_[103515]_ , \new_[103518]_ , \new_[103521]_ ,
    \new_[103522]_ , \new_[103523]_ , \new_[103526]_ , \new_[103529]_ ,
    \new_[103530]_ , \new_[103533]_ , \new_[103537]_ , \new_[103538]_ ,
    \new_[103539]_ , \new_[103540]_ , \new_[103543]_ , \new_[103546]_ ,
    \new_[103547]_ , \new_[103550]_ , \new_[103553]_ , \new_[103554]_ ,
    \new_[103555]_ , \new_[103558]_ , \new_[103561]_ , \new_[103562]_ ,
    \new_[103565]_ , \new_[103569]_ , \new_[103570]_ , \new_[103571]_ ,
    \new_[103572]_ , \new_[103575]_ , \new_[103578]_ , \new_[103579]_ ,
    \new_[103582]_ , \new_[103585]_ , \new_[103586]_ , \new_[103587]_ ,
    \new_[103590]_ , \new_[103593]_ , \new_[103594]_ , \new_[103597]_ ,
    \new_[103601]_ , \new_[103602]_ , \new_[103603]_ , \new_[103604]_ ,
    \new_[103607]_ , \new_[103610]_ , \new_[103611]_ , \new_[103614]_ ,
    \new_[103617]_ , \new_[103618]_ , \new_[103619]_ , \new_[103622]_ ,
    \new_[103625]_ , \new_[103626]_ , \new_[103629]_ , \new_[103633]_ ,
    \new_[103634]_ , \new_[103635]_ , \new_[103636]_ , \new_[103639]_ ,
    \new_[103642]_ , \new_[103643]_ , \new_[103646]_ , \new_[103649]_ ,
    \new_[103650]_ , \new_[103651]_ , \new_[103654]_ , \new_[103657]_ ,
    \new_[103658]_ , \new_[103661]_ , \new_[103665]_ , \new_[103666]_ ,
    \new_[103667]_ , \new_[103668]_ , \new_[103671]_ , \new_[103674]_ ,
    \new_[103675]_ , \new_[103678]_ , \new_[103681]_ , \new_[103682]_ ,
    \new_[103683]_ , \new_[103686]_ , \new_[103689]_ , \new_[103690]_ ,
    \new_[103693]_ , \new_[103697]_ , \new_[103698]_ , \new_[103699]_ ,
    \new_[103700]_ , \new_[103703]_ , \new_[103706]_ , \new_[103707]_ ,
    \new_[103710]_ , \new_[103713]_ , \new_[103714]_ , \new_[103715]_ ,
    \new_[103718]_ , \new_[103721]_ , \new_[103722]_ , \new_[103725]_ ,
    \new_[103729]_ , \new_[103730]_ , \new_[103731]_ , \new_[103732]_ ,
    \new_[103735]_ , \new_[103738]_ , \new_[103739]_ , \new_[103742]_ ,
    \new_[103745]_ , \new_[103746]_ , \new_[103747]_ , \new_[103750]_ ,
    \new_[103753]_ , \new_[103754]_ , \new_[103757]_ , \new_[103761]_ ,
    \new_[103762]_ , \new_[103763]_ , \new_[103764]_ , \new_[103767]_ ,
    \new_[103770]_ , \new_[103771]_ , \new_[103774]_ , \new_[103777]_ ,
    \new_[103778]_ , \new_[103779]_ , \new_[103782]_ , \new_[103785]_ ,
    \new_[103786]_ , \new_[103789]_ , \new_[103793]_ , \new_[103794]_ ,
    \new_[103795]_ , \new_[103796]_ , \new_[103799]_ , \new_[103802]_ ,
    \new_[103803]_ , \new_[103806]_ , \new_[103809]_ , \new_[103810]_ ,
    \new_[103811]_ , \new_[103814]_ , \new_[103817]_ , \new_[103818]_ ,
    \new_[103821]_ , \new_[103825]_ , \new_[103826]_ , \new_[103827]_ ,
    \new_[103828]_ , \new_[103831]_ , \new_[103834]_ , \new_[103835]_ ,
    \new_[103838]_ , \new_[103841]_ , \new_[103842]_ , \new_[103843]_ ,
    \new_[103846]_ , \new_[103849]_ , \new_[103850]_ , \new_[103853]_ ,
    \new_[103857]_ , \new_[103858]_ , \new_[103859]_ , \new_[103860]_ ,
    \new_[103863]_ , \new_[103866]_ , \new_[103867]_ , \new_[103870]_ ,
    \new_[103873]_ , \new_[103874]_ , \new_[103875]_ , \new_[103878]_ ,
    \new_[103881]_ , \new_[103882]_ , \new_[103885]_ , \new_[103889]_ ,
    \new_[103890]_ , \new_[103891]_ , \new_[103892]_ , \new_[103895]_ ,
    \new_[103898]_ , \new_[103899]_ , \new_[103902]_ , \new_[103905]_ ,
    \new_[103906]_ , \new_[103907]_ , \new_[103910]_ , \new_[103913]_ ,
    \new_[103914]_ , \new_[103917]_ , \new_[103921]_ , \new_[103922]_ ,
    \new_[103923]_ , \new_[103924]_ , \new_[103927]_ , \new_[103930]_ ,
    \new_[103931]_ , \new_[103934]_ , \new_[103937]_ , \new_[103938]_ ,
    \new_[103939]_ , \new_[103942]_ , \new_[103945]_ , \new_[103946]_ ,
    \new_[103949]_ , \new_[103953]_ , \new_[103954]_ , \new_[103955]_ ,
    \new_[103956]_ , \new_[103959]_ , \new_[103962]_ , \new_[103963]_ ,
    \new_[103966]_ , \new_[103969]_ , \new_[103970]_ , \new_[103971]_ ,
    \new_[103974]_ , \new_[103977]_ , \new_[103978]_ , \new_[103981]_ ,
    \new_[103985]_ , \new_[103986]_ , \new_[103987]_ , \new_[103988]_ ,
    \new_[103991]_ , \new_[103994]_ , \new_[103995]_ , \new_[103998]_ ,
    \new_[104001]_ , \new_[104002]_ , \new_[104003]_ , \new_[104006]_ ,
    \new_[104009]_ , \new_[104010]_ , \new_[104013]_ , \new_[104017]_ ,
    \new_[104018]_ , \new_[104019]_ , \new_[104020]_ , \new_[104023]_ ,
    \new_[104026]_ , \new_[104027]_ , \new_[104030]_ , \new_[104033]_ ,
    \new_[104034]_ , \new_[104035]_ , \new_[104038]_ , \new_[104041]_ ,
    \new_[104042]_ , \new_[104045]_ , \new_[104049]_ , \new_[104050]_ ,
    \new_[104051]_ , \new_[104052]_ , \new_[104055]_ , \new_[104058]_ ,
    \new_[104059]_ , \new_[104062]_ , \new_[104065]_ , \new_[104066]_ ,
    \new_[104067]_ , \new_[104070]_ , \new_[104073]_ , \new_[104074]_ ,
    \new_[104077]_ , \new_[104081]_ , \new_[104082]_ , \new_[104083]_ ,
    \new_[104084]_ , \new_[104087]_ , \new_[104090]_ , \new_[104091]_ ,
    \new_[104094]_ , \new_[104097]_ , \new_[104098]_ , \new_[104099]_ ,
    \new_[104102]_ , \new_[104105]_ , \new_[104106]_ , \new_[104109]_ ,
    \new_[104113]_ , \new_[104114]_ , \new_[104115]_ , \new_[104116]_ ,
    \new_[104119]_ , \new_[104122]_ , \new_[104123]_ , \new_[104126]_ ,
    \new_[104129]_ , \new_[104130]_ , \new_[104131]_ , \new_[104134]_ ,
    \new_[104137]_ , \new_[104138]_ , \new_[104141]_ , \new_[104145]_ ,
    \new_[104146]_ , \new_[104147]_ , \new_[104148]_ , \new_[104151]_ ,
    \new_[104154]_ , \new_[104155]_ , \new_[104158]_ , \new_[104161]_ ,
    \new_[104162]_ , \new_[104163]_ , \new_[104166]_ , \new_[104169]_ ,
    \new_[104170]_ , \new_[104173]_ , \new_[104177]_ , \new_[104178]_ ,
    \new_[104179]_ , \new_[104180]_ , \new_[104183]_ , \new_[104186]_ ,
    \new_[104187]_ , \new_[104190]_ , \new_[104193]_ , \new_[104194]_ ,
    \new_[104195]_ , \new_[104198]_ , \new_[104201]_ , \new_[104202]_ ,
    \new_[104205]_ , \new_[104209]_ , \new_[104210]_ , \new_[104211]_ ,
    \new_[104212]_ , \new_[104215]_ , \new_[104218]_ , \new_[104219]_ ,
    \new_[104222]_ , \new_[104225]_ , \new_[104226]_ , \new_[104227]_ ,
    \new_[104230]_ , \new_[104233]_ , \new_[104234]_ , \new_[104237]_ ,
    \new_[104241]_ , \new_[104242]_ , \new_[104243]_ , \new_[104244]_ ,
    \new_[104247]_ , \new_[104250]_ , \new_[104251]_ , \new_[104254]_ ,
    \new_[104257]_ , \new_[104258]_ , \new_[104259]_ , \new_[104262]_ ,
    \new_[104265]_ , \new_[104266]_ , \new_[104269]_ , \new_[104273]_ ,
    \new_[104274]_ , \new_[104275]_ , \new_[104276]_ , \new_[104279]_ ,
    \new_[104282]_ , \new_[104283]_ , \new_[104286]_ , \new_[104289]_ ,
    \new_[104290]_ , \new_[104291]_ , \new_[104294]_ , \new_[104297]_ ,
    \new_[104298]_ , \new_[104301]_ , \new_[104305]_ , \new_[104306]_ ,
    \new_[104307]_ , \new_[104308]_ , \new_[104311]_ , \new_[104314]_ ,
    \new_[104315]_ , \new_[104318]_ , \new_[104322]_ , \new_[104323]_ ,
    \new_[104324]_ , \new_[104325]_ , \new_[104328]_ , \new_[104331]_ ,
    \new_[104332]_ , \new_[104335]_ , \new_[104339]_ , \new_[104340]_ ,
    \new_[104341]_ , \new_[104342]_ , \new_[104345]_ , \new_[104348]_ ,
    \new_[104349]_ , \new_[104352]_ , \new_[104356]_ , \new_[104357]_ ,
    \new_[104358]_ , \new_[104359]_ , \new_[104362]_ , \new_[104365]_ ,
    \new_[104366]_ , \new_[104369]_ , \new_[104373]_ , \new_[104374]_ ,
    \new_[104375]_ , \new_[104376]_ , \new_[104379]_ , \new_[104382]_ ,
    \new_[104383]_ , \new_[104386]_ , \new_[104390]_ , \new_[104391]_ ,
    \new_[104392]_ , \new_[104393]_ , \new_[104396]_ , \new_[104399]_ ,
    \new_[104400]_ , \new_[104403]_ , \new_[104407]_ , \new_[104408]_ ,
    \new_[104409]_ , \new_[104410]_ , \new_[104413]_ , \new_[104416]_ ,
    \new_[104417]_ , \new_[104420]_ , \new_[104424]_ , \new_[104425]_ ,
    \new_[104426]_ , \new_[104427]_ , \new_[104430]_ , \new_[104433]_ ,
    \new_[104434]_ , \new_[104437]_ , \new_[104441]_ , \new_[104442]_ ,
    \new_[104443]_ , \new_[104444]_ , \new_[104447]_ , \new_[104450]_ ,
    \new_[104451]_ , \new_[104454]_ , \new_[104458]_ , \new_[104459]_ ,
    \new_[104460]_ , \new_[104461]_ , \new_[104464]_ , \new_[104467]_ ,
    \new_[104468]_ , \new_[104471]_ , \new_[104475]_ , \new_[104476]_ ,
    \new_[104477]_ , \new_[104478]_ , \new_[104481]_ , \new_[104484]_ ,
    \new_[104485]_ , \new_[104488]_ , \new_[104492]_ , \new_[104493]_ ,
    \new_[104494]_ , \new_[104495]_ , \new_[104498]_ , \new_[104501]_ ,
    \new_[104502]_ , \new_[104505]_ , \new_[104509]_ , \new_[104510]_ ,
    \new_[104511]_ , \new_[104512]_ , \new_[104515]_ , \new_[104518]_ ,
    \new_[104519]_ , \new_[104522]_ , \new_[104526]_ , \new_[104527]_ ,
    \new_[104528]_ , \new_[104529]_ , \new_[104532]_ , \new_[104535]_ ,
    \new_[104536]_ , \new_[104539]_ , \new_[104543]_ , \new_[104544]_ ,
    \new_[104545]_ , \new_[104546]_ , \new_[104549]_ , \new_[104552]_ ,
    \new_[104553]_ , \new_[104556]_ , \new_[104560]_ , \new_[104561]_ ,
    \new_[104562]_ , \new_[104563]_ , \new_[104566]_ , \new_[104569]_ ,
    \new_[104570]_ , \new_[104573]_ , \new_[104577]_ , \new_[104578]_ ,
    \new_[104579]_ , \new_[104580]_ ;
  assign A7 = \new_[11512]_  | \new_[7675]_ ;
  assign \new_[1]_  = \new_[104580]_  & \new_[104563]_ ;
  assign \new_[2]_  = \new_[104546]_  & \new_[104529]_ ;
  assign \new_[3]_  = \new_[104512]_  & \new_[104495]_ ;
  assign \new_[4]_  = \new_[104478]_  & \new_[104461]_ ;
  assign \new_[5]_  = \new_[104444]_  & \new_[104427]_ ;
  assign \new_[6]_  = \new_[104410]_  & \new_[104393]_ ;
  assign \new_[7]_  = \new_[104376]_  & \new_[104359]_ ;
  assign \new_[8]_  = \new_[104342]_  & \new_[104325]_ ;
  assign \new_[9]_  = \new_[104308]_  & \new_[104291]_ ;
  assign \new_[10]_  = \new_[104276]_  & \new_[104259]_ ;
  assign \new_[11]_  = \new_[104244]_  & \new_[104227]_ ;
  assign \new_[12]_  = \new_[104212]_  & \new_[104195]_ ;
  assign \new_[13]_  = \new_[104180]_  & \new_[104163]_ ;
  assign \new_[14]_  = \new_[104148]_  & \new_[104131]_ ;
  assign \new_[15]_  = \new_[104116]_  & \new_[104099]_ ;
  assign \new_[16]_  = \new_[104084]_  & \new_[104067]_ ;
  assign \new_[17]_  = \new_[104052]_  & \new_[104035]_ ;
  assign \new_[18]_  = \new_[104020]_  & \new_[104003]_ ;
  assign \new_[19]_  = \new_[103988]_  & \new_[103971]_ ;
  assign \new_[20]_  = \new_[103956]_  & \new_[103939]_ ;
  assign \new_[21]_  = \new_[103924]_  & \new_[103907]_ ;
  assign \new_[22]_  = \new_[103892]_  & \new_[103875]_ ;
  assign \new_[23]_  = \new_[103860]_  & \new_[103843]_ ;
  assign \new_[24]_  = \new_[103828]_  & \new_[103811]_ ;
  assign \new_[25]_  = \new_[103796]_  & \new_[103779]_ ;
  assign \new_[26]_  = \new_[103764]_  & \new_[103747]_ ;
  assign \new_[27]_  = \new_[103732]_  & \new_[103715]_ ;
  assign \new_[28]_  = \new_[103700]_  & \new_[103683]_ ;
  assign \new_[29]_  = \new_[103668]_  & \new_[103651]_ ;
  assign \new_[30]_  = \new_[103636]_  & \new_[103619]_ ;
  assign \new_[31]_  = \new_[103604]_  & \new_[103587]_ ;
  assign \new_[32]_  = \new_[103572]_  & \new_[103555]_ ;
  assign \new_[33]_  = \new_[103540]_  & \new_[103523]_ ;
  assign \new_[34]_  = \new_[103508]_  & \new_[103491]_ ;
  assign \new_[35]_  = \new_[103476]_  & \new_[103459]_ ;
  assign \new_[36]_  = \new_[103444]_  & \new_[103427]_ ;
  assign \new_[37]_  = \new_[103412]_  & \new_[103395]_ ;
  assign \new_[38]_  = \new_[103380]_  & \new_[103363]_ ;
  assign \new_[39]_  = \new_[103348]_  & \new_[103331]_ ;
  assign \new_[40]_  = \new_[103316]_  & \new_[103299]_ ;
  assign \new_[41]_  = \new_[103284]_  & \new_[103267]_ ;
  assign \new_[42]_  = \new_[103252]_  & \new_[103235]_ ;
  assign \new_[43]_  = \new_[103220]_  & \new_[103203]_ ;
  assign \new_[44]_  = \new_[103188]_  & \new_[103171]_ ;
  assign \new_[45]_  = \new_[103156]_  & \new_[103139]_ ;
  assign \new_[46]_  = \new_[103124]_  & \new_[103107]_ ;
  assign \new_[47]_  = \new_[103092]_  & \new_[103075]_ ;
  assign \new_[48]_  = \new_[103060]_  & \new_[103043]_ ;
  assign \new_[49]_  = \new_[103028]_  & \new_[103011]_ ;
  assign \new_[50]_  = \new_[102996]_  & \new_[102979]_ ;
  assign \new_[51]_  = \new_[102964]_  & \new_[102947]_ ;
  assign \new_[52]_  = \new_[102932]_  & \new_[102915]_ ;
  assign \new_[53]_  = \new_[102900]_  & \new_[102883]_ ;
  assign \new_[54]_  = \new_[102868]_  & \new_[102851]_ ;
  assign \new_[55]_  = \new_[102836]_  & \new_[102819]_ ;
  assign \new_[56]_  = \new_[102804]_  & \new_[102787]_ ;
  assign \new_[57]_  = \new_[102772]_  & \new_[102755]_ ;
  assign \new_[58]_  = \new_[102740]_  & \new_[102723]_ ;
  assign \new_[59]_  = \new_[102708]_  & \new_[102691]_ ;
  assign \new_[60]_  = \new_[102676]_  & \new_[102659]_ ;
  assign \new_[61]_  = \new_[102644]_  & \new_[102627]_ ;
  assign \new_[62]_  = \new_[102612]_  & \new_[102595]_ ;
  assign \new_[63]_  = \new_[102580]_  & \new_[102563]_ ;
  assign \new_[64]_  = \new_[102548]_  & \new_[102531]_ ;
  assign \new_[65]_  = \new_[102516]_  & \new_[102499]_ ;
  assign \new_[66]_  = \new_[102484]_  & \new_[102467]_ ;
  assign \new_[67]_  = \new_[102452]_  & \new_[102435]_ ;
  assign \new_[68]_  = \new_[102420]_  & \new_[102403]_ ;
  assign \new_[69]_  = \new_[102388]_  & \new_[102371]_ ;
  assign \new_[70]_  = \new_[102356]_  & \new_[102339]_ ;
  assign \new_[71]_  = \new_[102324]_  & \new_[102307]_ ;
  assign \new_[72]_  = \new_[102292]_  & \new_[102275]_ ;
  assign \new_[73]_  = \new_[102260]_  & \new_[102243]_ ;
  assign \new_[74]_  = \new_[102228]_  & \new_[102211]_ ;
  assign \new_[75]_  = \new_[102196]_  & \new_[102179]_ ;
  assign \new_[76]_  = \new_[102164]_  & \new_[102147]_ ;
  assign \new_[77]_  = \new_[102132]_  & \new_[102115]_ ;
  assign \new_[78]_  = \new_[102100]_  & \new_[102083]_ ;
  assign \new_[79]_  = \new_[102068]_  & \new_[102051]_ ;
  assign \new_[80]_  = \new_[102036]_  & \new_[102019]_ ;
  assign \new_[81]_  = \new_[102004]_  & \new_[101987]_ ;
  assign \new_[82]_  = \new_[101972]_  & \new_[101955]_ ;
  assign \new_[83]_  = \new_[101940]_  & \new_[101923]_ ;
  assign \new_[84]_  = \new_[101908]_  & \new_[101891]_ ;
  assign \new_[85]_  = \new_[101876]_  & \new_[101859]_ ;
  assign \new_[86]_  = \new_[101844]_  & \new_[101827]_ ;
  assign \new_[87]_  = \new_[101812]_  & \new_[101795]_ ;
  assign \new_[88]_  = \new_[101780]_  & \new_[101763]_ ;
  assign \new_[89]_  = \new_[101748]_  & \new_[101733]_ ;
  assign \new_[90]_  = \new_[101718]_  & \new_[101703]_ ;
  assign \new_[91]_  = \new_[101688]_  & \new_[101673]_ ;
  assign \new_[92]_  = \new_[101658]_  & \new_[101643]_ ;
  assign \new_[93]_  = \new_[101628]_  & \new_[101613]_ ;
  assign \new_[94]_  = \new_[101598]_  & \new_[101583]_ ;
  assign \new_[95]_  = \new_[101568]_  & \new_[101553]_ ;
  assign \new_[96]_  = \new_[101538]_  & \new_[101523]_ ;
  assign \new_[97]_  = \new_[101508]_  & \new_[101493]_ ;
  assign \new_[98]_  = \new_[101478]_  & \new_[101463]_ ;
  assign \new_[99]_  = \new_[101448]_  & \new_[101433]_ ;
  assign \new_[100]_  = \new_[101418]_  & \new_[101403]_ ;
  assign \new_[101]_  = \new_[101388]_  & \new_[101373]_ ;
  assign \new_[102]_  = \new_[101358]_  & \new_[101343]_ ;
  assign \new_[103]_  = \new_[101328]_  & \new_[101313]_ ;
  assign \new_[104]_  = \new_[101298]_  & \new_[101283]_ ;
  assign \new_[105]_  = \new_[101268]_  & \new_[101253]_ ;
  assign \new_[106]_  = \new_[101238]_  & \new_[101223]_ ;
  assign \new_[107]_  = \new_[101208]_  & \new_[101193]_ ;
  assign \new_[108]_  = \new_[101178]_  & \new_[101163]_ ;
  assign \new_[109]_  = \new_[101148]_  & \new_[101133]_ ;
  assign \new_[110]_  = \new_[101118]_  & \new_[101103]_ ;
  assign \new_[111]_  = \new_[101088]_  & \new_[101073]_ ;
  assign \new_[112]_  = \new_[101058]_  & \new_[101043]_ ;
  assign \new_[113]_  = \new_[101028]_  & \new_[101013]_ ;
  assign \new_[114]_  = \new_[100998]_  & \new_[100983]_ ;
  assign \new_[115]_  = \new_[100968]_  & \new_[100953]_ ;
  assign \new_[116]_  = \new_[100938]_  & \new_[100923]_ ;
  assign \new_[117]_  = \new_[100908]_  & \new_[100893]_ ;
  assign \new_[118]_  = \new_[100878]_  & \new_[100863]_ ;
  assign \new_[119]_  = \new_[100848]_  & \new_[100833]_ ;
  assign \new_[120]_  = \new_[100818]_  & \new_[100803]_ ;
  assign \new_[121]_  = \new_[100788]_  & \new_[100773]_ ;
  assign \new_[122]_  = \new_[100758]_  & \new_[100743]_ ;
  assign \new_[123]_  = \new_[100728]_  & \new_[100713]_ ;
  assign \new_[124]_  = \new_[100698]_  & \new_[100683]_ ;
  assign \new_[125]_  = \new_[100668]_  & \new_[100653]_ ;
  assign \new_[126]_  = \new_[100638]_  & \new_[100623]_ ;
  assign \new_[127]_  = \new_[100608]_  & \new_[100593]_ ;
  assign \new_[128]_  = \new_[100578]_  & \new_[100563]_ ;
  assign \new_[129]_  = \new_[100548]_  & \new_[100533]_ ;
  assign \new_[130]_  = \new_[100518]_  & \new_[100503]_ ;
  assign \new_[131]_  = \new_[100488]_  & \new_[100473]_ ;
  assign \new_[132]_  = \new_[100458]_  & \new_[100443]_ ;
  assign \new_[133]_  = \new_[100428]_  & \new_[100413]_ ;
  assign \new_[134]_  = \new_[100398]_  & \new_[100383]_ ;
  assign \new_[135]_  = \new_[100368]_  & \new_[100353]_ ;
  assign \new_[136]_  = \new_[100338]_  & \new_[100323]_ ;
  assign \new_[137]_  = \new_[100308]_  & \new_[100293]_ ;
  assign \new_[138]_  = \new_[100278]_  & \new_[100263]_ ;
  assign \new_[139]_  = \new_[100248]_  & \new_[100233]_ ;
  assign \new_[140]_  = \new_[100218]_  & \new_[100203]_ ;
  assign \new_[141]_  = \new_[100188]_  & \new_[100173]_ ;
  assign \new_[142]_  = \new_[100158]_  & \new_[100143]_ ;
  assign \new_[143]_  = \new_[100128]_  & \new_[100113]_ ;
  assign \new_[144]_  = \new_[100098]_  & \new_[100083]_ ;
  assign \new_[145]_  = \new_[100068]_  & \new_[100053]_ ;
  assign \new_[146]_  = \new_[100038]_  & \new_[100023]_ ;
  assign \new_[147]_  = \new_[100008]_  & \new_[99993]_ ;
  assign \new_[148]_  = \new_[99978]_  & \new_[99963]_ ;
  assign \new_[149]_  = \new_[99948]_  & \new_[99933]_ ;
  assign \new_[150]_  = \new_[99918]_  & \new_[99903]_ ;
  assign \new_[151]_  = \new_[99888]_  & \new_[99873]_ ;
  assign \new_[152]_  = \new_[99858]_  & \new_[99843]_ ;
  assign \new_[153]_  = \new_[99828]_  & \new_[99813]_ ;
  assign \new_[154]_  = \new_[99798]_  & \new_[99783]_ ;
  assign \new_[155]_  = \new_[99768]_  & \new_[99753]_ ;
  assign \new_[156]_  = \new_[99738]_  & \new_[99723]_ ;
  assign \new_[157]_  = \new_[99708]_  & \new_[99693]_ ;
  assign \new_[158]_  = \new_[99678]_  & \new_[99663]_ ;
  assign \new_[159]_  = \new_[99648]_  & \new_[99633]_ ;
  assign \new_[160]_  = \new_[99618]_  & \new_[99603]_ ;
  assign \new_[161]_  = \new_[99588]_  & \new_[99573]_ ;
  assign \new_[162]_  = \new_[99558]_  & \new_[99543]_ ;
  assign \new_[163]_  = \new_[99528]_  & \new_[99513]_ ;
  assign \new_[164]_  = \new_[99498]_  & \new_[99483]_ ;
  assign \new_[165]_  = \new_[99468]_  & \new_[99453]_ ;
  assign \new_[166]_  = \new_[99438]_  & \new_[99423]_ ;
  assign \new_[167]_  = \new_[99408]_  & \new_[99393]_ ;
  assign \new_[168]_  = \new_[99378]_  & \new_[99363]_ ;
  assign \new_[169]_  = \new_[99348]_  & \new_[99333]_ ;
  assign \new_[170]_  = \new_[99318]_  & \new_[99303]_ ;
  assign \new_[171]_  = \new_[99288]_  & \new_[99273]_ ;
  assign \new_[172]_  = \new_[99258]_  & \new_[99243]_ ;
  assign \new_[173]_  = \new_[99228]_  & \new_[99213]_ ;
  assign \new_[174]_  = \new_[99198]_  & \new_[99183]_ ;
  assign \new_[175]_  = \new_[99168]_  & \new_[99153]_ ;
  assign \new_[176]_  = \new_[99138]_  & \new_[99123]_ ;
  assign \new_[177]_  = \new_[99108]_  & \new_[99093]_ ;
  assign \new_[178]_  = \new_[99078]_  & \new_[99063]_ ;
  assign \new_[179]_  = \new_[99048]_  & \new_[99033]_ ;
  assign \new_[180]_  = \new_[99018]_  & \new_[99003]_ ;
  assign \new_[181]_  = \new_[98988]_  & \new_[98973]_ ;
  assign \new_[182]_  = \new_[98958]_  & \new_[98943]_ ;
  assign \new_[183]_  = \new_[98928]_  & \new_[98913]_ ;
  assign \new_[184]_  = \new_[98898]_  & \new_[98883]_ ;
  assign \new_[185]_  = \new_[98868]_  & \new_[98853]_ ;
  assign \new_[186]_  = \new_[98838]_  & \new_[98823]_ ;
  assign \new_[187]_  = \new_[98808]_  & \new_[98793]_ ;
  assign \new_[188]_  = \new_[98778]_  & \new_[98763]_ ;
  assign \new_[189]_  = \new_[98748]_  & \new_[98733]_ ;
  assign \new_[190]_  = \new_[98718]_  & \new_[98703]_ ;
  assign \new_[191]_  = \new_[98688]_  & \new_[98673]_ ;
  assign \new_[192]_  = \new_[98658]_  & \new_[98643]_ ;
  assign \new_[193]_  = \new_[98628]_  & \new_[98613]_ ;
  assign \new_[194]_  = \new_[98598]_  & \new_[98583]_ ;
  assign \new_[195]_  = \new_[98568]_  & \new_[98553]_ ;
  assign \new_[196]_  = \new_[98538]_  & \new_[98523]_ ;
  assign \new_[197]_  = \new_[98508]_  & \new_[98493]_ ;
  assign \new_[198]_  = \new_[98478]_  & \new_[98463]_ ;
  assign \new_[199]_  = \new_[98448]_  & \new_[98433]_ ;
  assign \new_[200]_  = \new_[98418]_  & \new_[98403]_ ;
  assign \new_[201]_  = \new_[98388]_  & \new_[98373]_ ;
  assign \new_[202]_  = \new_[98358]_  & \new_[98343]_ ;
  assign \new_[203]_  = \new_[98328]_  & \new_[98313]_ ;
  assign \new_[204]_  = \new_[98298]_  & \new_[98283]_ ;
  assign \new_[205]_  = \new_[98268]_  & \new_[98253]_ ;
  assign \new_[206]_  = \new_[98238]_  & \new_[98223]_ ;
  assign \new_[207]_  = \new_[98208]_  & \new_[98193]_ ;
  assign \new_[208]_  = \new_[98178]_  & \new_[98163]_ ;
  assign \new_[209]_  = \new_[98148]_  & \new_[98133]_ ;
  assign \new_[210]_  = \new_[98118]_  & \new_[98103]_ ;
  assign \new_[211]_  = \new_[98088]_  & \new_[98073]_ ;
  assign \new_[212]_  = \new_[98058]_  & \new_[98043]_ ;
  assign \new_[213]_  = \new_[98028]_  & \new_[98013]_ ;
  assign \new_[214]_  = \new_[97998]_  & \new_[97983]_ ;
  assign \new_[215]_  = \new_[97968]_  & \new_[97953]_ ;
  assign \new_[216]_  = \new_[97938]_  & \new_[97923]_ ;
  assign \new_[217]_  = \new_[97908]_  & \new_[97893]_ ;
  assign \new_[218]_  = \new_[97878]_  & \new_[97863]_ ;
  assign \new_[219]_  = \new_[97848]_  & \new_[97833]_ ;
  assign \new_[220]_  = \new_[97818]_  & \new_[97803]_ ;
  assign \new_[221]_  = \new_[97788]_  & \new_[97773]_ ;
  assign \new_[222]_  = \new_[97758]_  & \new_[97743]_ ;
  assign \new_[223]_  = \new_[97728]_  & \new_[97713]_ ;
  assign \new_[224]_  = \new_[97698]_  & \new_[97683]_ ;
  assign \new_[225]_  = \new_[97668]_  & \new_[97653]_ ;
  assign \new_[226]_  = \new_[97638]_  & \new_[97623]_ ;
  assign \new_[227]_  = \new_[97608]_  & \new_[97593]_ ;
  assign \new_[228]_  = \new_[97578]_  & \new_[97563]_ ;
  assign \new_[229]_  = \new_[97548]_  & \new_[97533]_ ;
  assign \new_[230]_  = \new_[97518]_  & \new_[97503]_ ;
  assign \new_[231]_  = \new_[97488]_  & \new_[97473]_ ;
  assign \new_[232]_  = \new_[97458]_  & \new_[97443]_ ;
  assign \new_[233]_  = \new_[97428]_  & \new_[97413]_ ;
  assign \new_[234]_  = \new_[97398]_  & \new_[97383]_ ;
  assign \new_[235]_  = \new_[97368]_  & \new_[97353]_ ;
  assign \new_[236]_  = \new_[97338]_  & \new_[97323]_ ;
  assign \new_[237]_  = \new_[97308]_  & \new_[97293]_ ;
  assign \new_[238]_  = \new_[97278]_  & \new_[97263]_ ;
  assign \new_[239]_  = \new_[97248]_  & \new_[97233]_ ;
  assign \new_[240]_  = \new_[97218]_  & \new_[97203]_ ;
  assign \new_[241]_  = \new_[97188]_  & \new_[97173]_ ;
  assign \new_[242]_  = \new_[97158]_  & \new_[97143]_ ;
  assign \new_[243]_  = \new_[97128]_  & \new_[97113]_ ;
  assign \new_[244]_  = \new_[97098]_  & \new_[97083]_ ;
  assign \new_[245]_  = \new_[97068]_  & \new_[97053]_ ;
  assign \new_[246]_  = \new_[97038]_  & \new_[97023]_ ;
  assign \new_[247]_  = \new_[97008]_  & \new_[96993]_ ;
  assign \new_[248]_  = \new_[96978]_  & \new_[96963]_ ;
  assign \new_[249]_  = \new_[96948]_  & \new_[96933]_ ;
  assign \new_[250]_  = \new_[96918]_  & \new_[96903]_ ;
  assign \new_[251]_  = \new_[96888]_  & \new_[96873]_ ;
  assign \new_[252]_  = \new_[96858]_  & \new_[96843]_ ;
  assign \new_[253]_  = \new_[96828]_  & \new_[96813]_ ;
  assign \new_[254]_  = \new_[96798]_  & \new_[96783]_ ;
  assign \new_[255]_  = \new_[96768]_  & \new_[96753]_ ;
  assign \new_[256]_  = \new_[96738]_  & \new_[96723]_ ;
  assign \new_[257]_  = \new_[96708]_  & \new_[96693]_ ;
  assign \new_[258]_  = \new_[96678]_  & \new_[96663]_ ;
  assign \new_[259]_  = \new_[96648]_  & \new_[96633]_ ;
  assign \new_[260]_  = \new_[96618]_  & \new_[96603]_ ;
  assign \new_[261]_  = \new_[96588]_  & \new_[96573]_ ;
  assign \new_[262]_  = \new_[96558]_  & \new_[96543]_ ;
  assign \new_[263]_  = \new_[96528]_  & \new_[96513]_ ;
  assign \new_[264]_  = \new_[96498]_  & \new_[96483]_ ;
  assign \new_[265]_  = \new_[96468]_  & \new_[96453]_ ;
  assign \new_[266]_  = \new_[96438]_  & \new_[96423]_ ;
  assign \new_[267]_  = \new_[96408]_  & \new_[96393]_ ;
  assign \new_[268]_  = \new_[96378]_  & \new_[96363]_ ;
  assign \new_[269]_  = \new_[96348]_  & \new_[96333]_ ;
  assign \new_[270]_  = \new_[96318]_  & \new_[96303]_ ;
  assign \new_[271]_  = \new_[96288]_  & \new_[96273]_ ;
  assign \new_[272]_  = \new_[96258]_  & \new_[96243]_ ;
  assign \new_[273]_  = \new_[96228]_  & \new_[96213]_ ;
  assign \new_[274]_  = \new_[96198]_  & \new_[96183]_ ;
  assign \new_[275]_  = \new_[96168]_  & \new_[96153]_ ;
  assign \new_[276]_  = \new_[96138]_  & \new_[96123]_ ;
  assign \new_[277]_  = \new_[96108]_  & \new_[96093]_ ;
  assign \new_[278]_  = \new_[96078]_  & \new_[96063]_ ;
  assign \new_[279]_  = \new_[96048]_  & \new_[96033]_ ;
  assign \new_[280]_  = \new_[96018]_  & \new_[96003]_ ;
  assign \new_[281]_  = \new_[95988]_  & \new_[95973]_ ;
  assign \new_[282]_  = \new_[95958]_  & \new_[95943]_ ;
  assign \new_[283]_  = \new_[95928]_  & \new_[95913]_ ;
  assign \new_[284]_  = \new_[95898]_  & \new_[95883]_ ;
  assign \new_[285]_  = \new_[95868]_  & \new_[95853]_ ;
  assign \new_[286]_  = \new_[95838]_  & \new_[95823]_ ;
  assign \new_[287]_  = \new_[95808]_  & \new_[95793]_ ;
  assign \new_[288]_  = \new_[95778]_  & \new_[95763]_ ;
  assign \new_[289]_  = \new_[95748]_  & \new_[95733]_ ;
  assign \new_[290]_  = \new_[95718]_  & \new_[95703]_ ;
  assign \new_[291]_  = \new_[95688]_  & \new_[95673]_ ;
  assign \new_[292]_  = \new_[95658]_  & \new_[95643]_ ;
  assign \new_[293]_  = \new_[95628]_  & \new_[95613]_ ;
  assign \new_[294]_  = \new_[95598]_  & \new_[95583]_ ;
  assign \new_[295]_  = \new_[95568]_  & \new_[95553]_ ;
  assign \new_[296]_  = \new_[95538]_  & \new_[95523]_ ;
  assign \new_[297]_  = \new_[95508]_  & \new_[95493]_ ;
  assign \new_[298]_  = \new_[95478]_  & \new_[95463]_ ;
  assign \new_[299]_  = \new_[95448]_  & \new_[95433]_ ;
  assign \new_[300]_  = \new_[95418]_  & \new_[95403]_ ;
  assign \new_[301]_  = \new_[95388]_  & \new_[95373]_ ;
  assign \new_[302]_  = \new_[95358]_  & \new_[95343]_ ;
  assign \new_[303]_  = \new_[95328]_  & \new_[95313]_ ;
  assign \new_[304]_  = \new_[95298]_  & \new_[95283]_ ;
  assign \new_[305]_  = \new_[95268]_  & \new_[95253]_ ;
  assign \new_[306]_  = \new_[95238]_  & \new_[95223]_ ;
  assign \new_[307]_  = \new_[95208]_  & \new_[95193]_ ;
  assign \new_[308]_  = \new_[95178]_  & \new_[95163]_ ;
  assign \new_[309]_  = \new_[95148]_  & \new_[95133]_ ;
  assign \new_[310]_  = \new_[95118]_  & \new_[95103]_ ;
  assign \new_[311]_  = \new_[95088]_  & \new_[95073]_ ;
  assign \new_[312]_  = \new_[95058]_  & \new_[95043]_ ;
  assign \new_[313]_  = \new_[95028]_  & \new_[95013]_ ;
  assign \new_[314]_  = \new_[94998]_  & \new_[94983]_ ;
  assign \new_[315]_  = \new_[94968]_  & \new_[94953]_ ;
  assign \new_[316]_  = \new_[94938]_  & \new_[94923]_ ;
  assign \new_[317]_  = \new_[94908]_  & \new_[94893]_ ;
  assign \new_[318]_  = \new_[94878]_  & \new_[94863]_ ;
  assign \new_[319]_  = \new_[94848]_  & \new_[94833]_ ;
  assign \new_[320]_  = \new_[94818]_  & \new_[94803]_ ;
  assign \new_[321]_  = \new_[94788]_  & \new_[94773]_ ;
  assign \new_[322]_  = \new_[94758]_  & \new_[94743]_ ;
  assign \new_[323]_  = \new_[94728]_  & \new_[94713]_ ;
  assign \new_[324]_  = \new_[94698]_  & \new_[94683]_ ;
  assign \new_[325]_  = \new_[94668]_  & \new_[94653]_ ;
  assign \new_[326]_  = \new_[94638]_  & \new_[94623]_ ;
  assign \new_[327]_  = \new_[94608]_  & \new_[94593]_ ;
  assign \new_[328]_  = \new_[94578]_  & \new_[94563]_ ;
  assign \new_[329]_  = \new_[94548]_  & \new_[94533]_ ;
  assign \new_[330]_  = \new_[94518]_  & \new_[94503]_ ;
  assign \new_[331]_  = \new_[94488]_  & \new_[94473]_ ;
  assign \new_[332]_  = \new_[94458]_  & \new_[94443]_ ;
  assign \new_[333]_  = \new_[94428]_  & \new_[94413]_ ;
  assign \new_[334]_  = \new_[94398]_  & \new_[94383]_ ;
  assign \new_[335]_  = \new_[94368]_  & \new_[94353]_ ;
  assign \new_[336]_  = \new_[94338]_  & \new_[94323]_ ;
  assign \new_[337]_  = \new_[94308]_  & \new_[94293]_ ;
  assign \new_[338]_  = \new_[94278]_  & \new_[94263]_ ;
  assign \new_[339]_  = \new_[94248]_  & \new_[94233]_ ;
  assign \new_[340]_  = \new_[94218]_  & \new_[94203]_ ;
  assign \new_[341]_  = \new_[94188]_  & \new_[94173]_ ;
  assign \new_[342]_  = \new_[94158]_  & \new_[94143]_ ;
  assign \new_[343]_  = \new_[94128]_  & \new_[94113]_ ;
  assign \new_[344]_  = \new_[94098]_  & \new_[94083]_ ;
  assign \new_[345]_  = \new_[94068]_  & \new_[94053]_ ;
  assign \new_[346]_  = \new_[94038]_  & \new_[94023]_ ;
  assign \new_[347]_  = \new_[94008]_  & \new_[93993]_ ;
  assign \new_[348]_  = \new_[93978]_  & \new_[93963]_ ;
  assign \new_[349]_  = \new_[93948]_  & \new_[93933]_ ;
  assign \new_[350]_  = \new_[93918]_  & \new_[93903]_ ;
  assign \new_[351]_  = \new_[93888]_  & \new_[93873]_ ;
  assign \new_[352]_  = \new_[93858]_  & \new_[93843]_ ;
  assign \new_[353]_  = \new_[93828]_  & \new_[93813]_ ;
  assign \new_[354]_  = \new_[93798]_  & \new_[93783]_ ;
  assign \new_[355]_  = \new_[93768]_  & \new_[93753]_ ;
  assign \new_[356]_  = \new_[93738]_  & \new_[93723]_ ;
  assign \new_[357]_  = \new_[93708]_  & \new_[93693]_ ;
  assign \new_[358]_  = \new_[93678]_  & \new_[93663]_ ;
  assign \new_[359]_  = \new_[93648]_  & \new_[93633]_ ;
  assign \new_[360]_  = \new_[93618]_  & \new_[93603]_ ;
  assign \new_[361]_  = \new_[93588]_  & \new_[93573]_ ;
  assign \new_[362]_  = \new_[93558]_  & \new_[93543]_ ;
  assign \new_[363]_  = \new_[93528]_  & \new_[93513]_ ;
  assign \new_[364]_  = \new_[93498]_  & \new_[93483]_ ;
  assign \new_[365]_  = \new_[93468]_  & \new_[93453]_ ;
  assign \new_[366]_  = \new_[93438]_  & \new_[93423]_ ;
  assign \new_[367]_  = \new_[93408]_  & \new_[93393]_ ;
  assign \new_[368]_  = \new_[93378]_  & \new_[93363]_ ;
  assign \new_[369]_  = \new_[93348]_  & \new_[93333]_ ;
  assign \new_[370]_  = \new_[93318]_  & \new_[93303]_ ;
  assign \new_[371]_  = \new_[93288]_  & \new_[93273]_ ;
  assign \new_[372]_  = \new_[93258]_  & \new_[93243]_ ;
  assign \new_[373]_  = \new_[93228]_  & \new_[93213]_ ;
  assign \new_[374]_  = \new_[93198]_  & \new_[93183]_ ;
  assign \new_[375]_  = \new_[93168]_  & \new_[93153]_ ;
  assign \new_[376]_  = \new_[93138]_  & \new_[93123]_ ;
  assign \new_[377]_  = \new_[93108]_  & \new_[93093]_ ;
  assign \new_[378]_  = \new_[93078]_  & \new_[93063]_ ;
  assign \new_[379]_  = \new_[93048]_  & \new_[93033]_ ;
  assign \new_[380]_  = \new_[93018]_  & \new_[93003]_ ;
  assign \new_[381]_  = \new_[92988]_  & \new_[92973]_ ;
  assign \new_[382]_  = \new_[92958]_  & \new_[92943]_ ;
  assign \new_[383]_  = \new_[92928]_  & \new_[92913]_ ;
  assign \new_[384]_  = \new_[92898]_  & \new_[92883]_ ;
  assign \new_[385]_  = \new_[92868]_  & \new_[92853]_ ;
  assign \new_[386]_  = \new_[92840]_  & \new_[92825]_ ;
  assign \new_[387]_  = \new_[92812]_  & \new_[92797]_ ;
  assign \new_[388]_  = \new_[92784]_  & \new_[92769]_ ;
  assign \new_[389]_  = \new_[92756]_  & \new_[92741]_ ;
  assign \new_[390]_  = \new_[92728]_  & \new_[92713]_ ;
  assign \new_[391]_  = \new_[92700]_  & \new_[92685]_ ;
  assign \new_[392]_  = \new_[92672]_  & \new_[92657]_ ;
  assign \new_[393]_  = \new_[92644]_  & \new_[92629]_ ;
  assign \new_[394]_  = \new_[92616]_  & \new_[92601]_ ;
  assign \new_[395]_  = \new_[92588]_  & \new_[92573]_ ;
  assign \new_[396]_  = \new_[92560]_  & \new_[92545]_ ;
  assign \new_[397]_  = \new_[92532]_  & \new_[92517]_ ;
  assign \new_[398]_  = \new_[92504]_  & \new_[92489]_ ;
  assign \new_[399]_  = \new_[92476]_  & \new_[92461]_ ;
  assign \new_[400]_  = \new_[92448]_  & \new_[92433]_ ;
  assign \new_[401]_  = \new_[92420]_  & \new_[92405]_ ;
  assign \new_[402]_  = \new_[92392]_  & \new_[92377]_ ;
  assign \new_[403]_  = \new_[92364]_  & \new_[92349]_ ;
  assign \new_[404]_  = \new_[92336]_  & \new_[92321]_ ;
  assign \new_[405]_  = \new_[92308]_  & \new_[92293]_ ;
  assign \new_[406]_  = \new_[92280]_  & \new_[92265]_ ;
  assign \new_[407]_  = \new_[92252]_  & \new_[92237]_ ;
  assign \new_[408]_  = \new_[92224]_  & \new_[92209]_ ;
  assign \new_[409]_  = \new_[92196]_  & \new_[92181]_ ;
  assign \new_[410]_  = \new_[92168]_  & \new_[92153]_ ;
  assign \new_[411]_  = \new_[92140]_  & \new_[92125]_ ;
  assign \new_[412]_  = \new_[92112]_  & \new_[92097]_ ;
  assign \new_[413]_  = \new_[92084]_  & \new_[92069]_ ;
  assign \new_[414]_  = \new_[92056]_  & \new_[92041]_ ;
  assign \new_[415]_  = \new_[92028]_  & \new_[92013]_ ;
  assign \new_[416]_  = \new_[92000]_  & \new_[91985]_ ;
  assign \new_[417]_  = \new_[91972]_  & \new_[91957]_ ;
  assign \new_[418]_  = \new_[91944]_  & \new_[91929]_ ;
  assign \new_[419]_  = \new_[91916]_  & \new_[91901]_ ;
  assign \new_[420]_  = \new_[91888]_  & \new_[91873]_ ;
  assign \new_[421]_  = \new_[91860]_  & \new_[91845]_ ;
  assign \new_[422]_  = \new_[91832]_  & \new_[91817]_ ;
  assign \new_[423]_  = \new_[91804]_  & \new_[91789]_ ;
  assign \new_[424]_  = \new_[91776]_  & \new_[91761]_ ;
  assign \new_[425]_  = \new_[91748]_  & \new_[91733]_ ;
  assign \new_[426]_  = \new_[91720]_  & \new_[91705]_ ;
  assign \new_[427]_  = \new_[91692]_  & \new_[91677]_ ;
  assign \new_[428]_  = \new_[91664]_  & \new_[91649]_ ;
  assign \new_[429]_  = \new_[91636]_  & \new_[91621]_ ;
  assign \new_[430]_  = \new_[91608]_  & \new_[91593]_ ;
  assign \new_[431]_  = \new_[91580]_  & \new_[91565]_ ;
  assign \new_[432]_  = \new_[91552]_  & \new_[91537]_ ;
  assign \new_[433]_  = \new_[91524]_  & \new_[91509]_ ;
  assign \new_[434]_  = \new_[91496]_  & \new_[91481]_ ;
  assign \new_[435]_  = \new_[91468]_  & \new_[91453]_ ;
  assign \new_[436]_  = \new_[91440]_  & \new_[91425]_ ;
  assign \new_[437]_  = \new_[91412]_  & \new_[91397]_ ;
  assign \new_[438]_  = \new_[91384]_  & \new_[91369]_ ;
  assign \new_[439]_  = \new_[91356]_  & \new_[91341]_ ;
  assign \new_[440]_  = \new_[91328]_  & \new_[91313]_ ;
  assign \new_[441]_  = \new_[91300]_  & \new_[91285]_ ;
  assign \new_[442]_  = \new_[91272]_  & \new_[91257]_ ;
  assign \new_[443]_  = \new_[91244]_  & \new_[91229]_ ;
  assign \new_[444]_  = \new_[91216]_  & \new_[91201]_ ;
  assign \new_[445]_  = \new_[91188]_  & \new_[91173]_ ;
  assign \new_[446]_  = \new_[91160]_  & \new_[91145]_ ;
  assign \new_[447]_  = \new_[91132]_  & \new_[91117]_ ;
  assign \new_[448]_  = \new_[91104]_  & \new_[91089]_ ;
  assign \new_[449]_  = \new_[91076]_  & \new_[91061]_ ;
  assign \new_[450]_  = \new_[91048]_  & \new_[91033]_ ;
  assign \new_[451]_  = \new_[91020]_  & \new_[91005]_ ;
  assign \new_[452]_  = \new_[90992]_  & \new_[90977]_ ;
  assign \new_[453]_  = \new_[90964]_  & \new_[90949]_ ;
  assign \new_[454]_  = \new_[90936]_  & \new_[90921]_ ;
  assign \new_[455]_  = \new_[90908]_  & \new_[90893]_ ;
  assign \new_[456]_  = \new_[90880]_  & \new_[90865]_ ;
  assign \new_[457]_  = \new_[90852]_  & \new_[90837]_ ;
  assign \new_[458]_  = \new_[90824]_  & \new_[90809]_ ;
  assign \new_[459]_  = \new_[90796]_  & \new_[90781]_ ;
  assign \new_[460]_  = \new_[90768]_  & \new_[90753]_ ;
  assign \new_[461]_  = \new_[90740]_  & \new_[90725]_ ;
  assign \new_[462]_  = \new_[90712]_  & \new_[90697]_ ;
  assign \new_[463]_  = \new_[90684]_  & \new_[90669]_ ;
  assign \new_[464]_  = \new_[90656]_  & \new_[90641]_ ;
  assign \new_[465]_  = \new_[90628]_  & \new_[90613]_ ;
  assign \new_[466]_  = \new_[90600]_  & \new_[90585]_ ;
  assign \new_[467]_  = \new_[90572]_  & \new_[90557]_ ;
  assign \new_[468]_  = \new_[90544]_  & \new_[90529]_ ;
  assign \new_[469]_  = \new_[90516]_  & \new_[90501]_ ;
  assign \new_[470]_  = \new_[90488]_  & \new_[90473]_ ;
  assign \new_[471]_  = \new_[90460]_  & \new_[90445]_ ;
  assign \new_[472]_  = \new_[90432]_  & \new_[90417]_ ;
  assign \new_[473]_  = \new_[90404]_  & \new_[90389]_ ;
  assign \new_[474]_  = \new_[90376]_  & \new_[90361]_ ;
  assign \new_[475]_  = \new_[90348]_  & \new_[90333]_ ;
  assign \new_[476]_  = \new_[90320]_  & \new_[90305]_ ;
  assign \new_[477]_  = \new_[90292]_  & \new_[90277]_ ;
  assign \new_[478]_  = \new_[90264]_  & \new_[90249]_ ;
  assign \new_[479]_  = \new_[90236]_  & \new_[90221]_ ;
  assign \new_[480]_  = \new_[90208]_  & \new_[90193]_ ;
  assign \new_[481]_  = \new_[90180]_  & \new_[90165]_ ;
  assign \new_[482]_  = \new_[90152]_  & \new_[90137]_ ;
  assign \new_[483]_  = \new_[90124]_  & \new_[90109]_ ;
  assign \new_[484]_  = \new_[90096]_  & \new_[90081]_ ;
  assign \new_[485]_  = \new_[90068]_  & \new_[90053]_ ;
  assign \new_[486]_  = \new_[90040]_  & \new_[90025]_ ;
  assign \new_[487]_  = \new_[90012]_  & \new_[89997]_ ;
  assign \new_[488]_  = \new_[89984]_  & \new_[89969]_ ;
  assign \new_[489]_  = \new_[89956]_  & \new_[89941]_ ;
  assign \new_[490]_  = \new_[89928]_  & \new_[89913]_ ;
  assign \new_[491]_  = \new_[89900]_  & \new_[89885]_ ;
  assign \new_[492]_  = \new_[89872]_  & \new_[89857]_ ;
  assign \new_[493]_  = \new_[89844]_  & \new_[89829]_ ;
  assign \new_[494]_  = \new_[89816]_  & \new_[89801]_ ;
  assign \new_[495]_  = \new_[89788]_  & \new_[89773]_ ;
  assign \new_[496]_  = \new_[89760]_  & \new_[89745]_ ;
  assign \new_[497]_  = \new_[89732]_  & \new_[89717]_ ;
  assign \new_[498]_  = \new_[89704]_  & \new_[89689]_ ;
  assign \new_[499]_  = \new_[89676]_  & \new_[89661]_ ;
  assign \new_[500]_  = \new_[89648]_  & \new_[89633]_ ;
  assign \new_[501]_  = \new_[89620]_  & \new_[89605]_ ;
  assign \new_[502]_  = \new_[89592]_  & \new_[89577]_ ;
  assign \new_[503]_  = \new_[89564]_  & \new_[89549]_ ;
  assign \new_[504]_  = \new_[89536]_  & \new_[89521]_ ;
  assign \new_[505]_  = \new_[89508]_  & \new_[89493]_ ;
  assign \new_[506]_  = \new_[89480]_  & \new_[89465]_ ;
  assign \new_[507]_  = \new_[89452]_  & \new_[89437]_ ;
  assign \new_[508]_  = \new_[89424]_  & \new_[89409]_ ;
  assign \new_[509]_  = \new_[89396]_  & \new_[89381]_ ;
  assign \new_[510]_  = \new_[89368]_  & \new_[89353]_ ;
  assign \new_[511]_  = \new_[89340]_  & \new_[89325]_ ;
  assign \new_[512]_  = \new_[89312]_  & \new_[89297]_ ;
  assign \new_[513]_  = \new_[89284]_  & \new_[89269]_ ;
  assign \new_[514]_  = \new_[89256]_  & \new_[89241]_ ;
  assign \new_[515]_  = \new_[89228]_  & \new_[89213]_ ;
  assign \new_[516]_  = \new_[89200]_  & \new_[89185]_ ;
  assign \new_[517]_  = \new_[89172]_  & \new_[89157]_ ;
  assign \new_[518]_  = \new_[89144]_  & \new_[89129]_ ;
  assign \new_[519]_  = \new_[89116]_  & \new_[89101]_ ;
  assign \new_[520]_  = \new_[89088]_  & \new_[89073]_ ;
  assign \new_[521]_  = \new_[89060]_  & \new_[89045]_ ;
  assign \new_[522]_  = \new_[89032]_  & \new_[89017]_ ;
  assign \new_[523]_  = \new_[89004]_  & \new_[88989]_ ;
  assign \new_[524]_  = \new_[88976]_  & \new_[88961]_ ;
  assign \new_[525]_  = \new_[88948]_  & \new_[88933]_ ;
  assign \new_[526]_  = \new_[88920]_  & \new_[88905]_ ;
  assign \new_[527]_  = \new_[88892]_  & \new_[88877]_ ;
  assign \new_[528]_  = \new_[88864]_  & \new_[88849]_ ;
  assign \new_[529]_  = \new_[88836]_  & \new_[88821]_ ;
  assign \new_[530]_  = \new_[88808]_  & \new_[88793]_ ;
  assign \new_[531]_  = \new_[88780]_  & \new_[88765]_ ;
  assign \new_[532]_  = \new_[88752]_  & \new_[88737]_ ;
  assign \new_[533]_  = \new_[88724]_  & \new_[88709]_ ;
  assign \new_[534]_  = \new_[88696]_  & \new_[88681]_ ;
  assign \new_[535]_  = \new_[88668]_  & \new_[88653]_ ;
  assign \new_[536]_  = \new_[88640]_  & \new_[88625]_ ;
  assign \new_[537]_  = \new_[88612]_  & \new_[88597]_ ;
  assign \new_[538]_  = \new_[88584]_  & \new_[88569]_ ;
  assign \new_[539]_  = \new_[88556]_  & \new_[88541]_ ;
  assign \new_[540]_  = \new_[88528]_  & \new_[88513]_ ;
  assign \new_[541]_  = \new_[88500]_  & \new_[88485]_ ;
  assign \new_[542]_  = \new_[88472]_  & \new_[88457]_ ;
  assign \new_[543]_  = \new_[88444]_  & \new_[88429]_ ;
  assign \new_[544]_  = \new_[88416]_  & \new_[88401]_ ;
  assign \new_[545]_  = \new_[88388]_  & \new_[88373]_ ;
  assign \new_[546]_  = \new_[88360]_  & \new_[88345]_ ;
  assign \new_[547]_  = \new_[88332]_  & \new_[88317]_ ;
  assign \new_[548]_  = \new_[88304]_  & \new_[88289]_ ;
  assign \new_[549]_  = \new_[88276]_  & \new_[88261]_ ;
  assign \new_[550]_  = \new_[88248]_  & \new_[88233]_ ;
  assign \new_[551]_  = \new_[88220]_  & \new_[88205]_ ;
  assign \new_[552]_  = \new_[88192]_  & \new_[88177]_ ;
  assign \new_[553]_  = \new_[88164]_  & \new_[88149]_ ;
  assign \new_[554]_  = \new_[88136]_  & \new_[88121]_ ;
  assign \new_[555]_  = \new_[88108]_  & \new_[88093]_ ;
  assign \new_[556]_  = \new_[88080]_  & \new_[88065]_ ;
  assign \new_[557]_  = \new_[88052]_  & \new_[88037]_ ;
  assign \new_[558]_  = \new_[88024]_  & \new_[88009]_ ;
  assign \new_[559]_  = \new_[87996]_  & \new_[87981]_ ;
  assign \new_[560]_  = \new_[87968]_  & \new_[87953]_ ;
  assign \new_[561]_  = \new_[87940]_  & \new_[87925]_ ;
  assign \new_[562]_  = \new_[87912]_  & \new_[87897]_ ;
  assign \new_[563]_  = \new_[87884]_  & \new_[87869]_ ;
  assign \new_[564]_  = \new_[87856]_  & \new_[87841]_ ;
  assign \new_[565]_  = \new_[87828]_  & \new_[87813]_ ;
  assign \new_[566]_  = \new_[87800]_  & \new_[87785]_ ;
  assign \new_[567]_  = \new_[87772]_  & \new_[87757]_ ;
  assign \new_[568]_  = \new_[87744]_  & \new_[87729]_ ;
  assign \new_[569]_  = \new_[87716]_  & \new_[87701]_ ;
  assign \new_[570]_  = \new_[87688]_  & \new_[87673]_ ;
  assign \new_[571]_  = \new_[87660]_  & \new_[87645]_ ;
  assign \new_[572]_  = \new_[87632]_  & \new_[87617]_ ;
  assign \new_[573]_  = \new_[87604]_  & \new_[87589]_ ;
  assign \new_[574]_  = \new_[87576]_  & \new_[87561]_ ;
  assign \new_[575]_  = \new_[87548]_  & \new_[87533]_ ;
  assign \new_[576]_  = \new_[87520]_  & \new_[87505]_ ;
  assign \new_[577]_  = \new_[87492]_  & \new_[87477]_ ;
  assign \new_[578]_  = \new_[87464]_  & \new_[87449]_ ;
  assign \new_[579]_  = \new_[87436]_  & \new_[87421]_ ;
  assign \new_[580]_  = \new_[87408]_  & \new_[87393]_ ;
  assign \new_[581]_  = \new_[87380]_  & \new_[87365]_ ;
  assign \new_[582]_  = \new_[87352]_  & \new_[87337]_ ;
  assign \new_[583]_  = \new_[87324]_  & \new_[87309]_ ;
  assign \new_[584]_  = \new_[87296]_  & \new_[87281]_ ;
  assign \new_[585]_  = \new_[87268]_  & \new_[87253]_ ;
  assign \new_[586]_  = \new_[87240]_  & \new_[87225]_ ;
  assign \new_[587]_  = \new_[87212]_  & \new_[87197]_ ;
  assign \new_[588]_  = \new_[87184]_  & \new_[87169]_ ;
  assign \new_[589]_  = \new_[87156]_  & \new_[87141]_ ;
  assign \new_[590]_  = \new_[87128]_  & \new_[87113]_ ;
  assign \new_[591]_  = \new_[87100]_  & \new_[87085]_ ;
  assign \new_[592]_  = \new_[87072]_  & \new_[87057]_ ;
  assign \new_[593]_  = \new_[87044]_  & \new_[87029]_ ;
  assign \new_[594]_  = \new_[87016]_  & \new_[87001]_ ;
  assign \new_[595]_  = \new_[86988]_  & \new_[86973]_ ;
  assign \new_[596]_  = \new_[86960]_  & \new_[86945]_ ;
  assign \new_[597]_  = \new_[86932]_  & \new_[86917]_ ;
  assign \new_[598]_  = \new_[86904]_  & \new_[86889]_ ;
  assign \new_[599]_  = \new_[86876]_  & \new_[86861]_ ;
  assign \new_[600]_  = \new_[86848]_  & \new_[86833]_ ;
  assign \new_[601]_  = \new_[86820]_  & \new_[86805]_ ;
  assign \new_[602]_  = \new_[86792]_  & \new_[86777]_ ;
  assign \new_[603]_  = \new_[86764]_  & \new_[86749]_ ;
  assign \new_[604]_  = \new_[86736]_  & \new_[86721]_ ;
  assign \new_[605]_  = \new_[86708]_  & \new_[86693]_ ;
  assign \new_[606]_  = \new_[86680]_  & \new_[86665]_ ;
  assign \new_[607]_  = \new_[86652]_  & \new_[86637]_ ;
  assign \new_[608]_  = \new_[86624]_  & \new_[86609]_ ;
  assign \new_[609]_  = \new_[86596]_  & \new_[86581]_ ;
  assign \new_[610]_  = \new_[86568]_  & \new_[86553]_ ;
  assign \new_[611]_  = \new_[86540]_  & \new_[86525]_ ;
  assign \new_[612]_  = \new_[86512]_  & \new_[86497]_ ;
  assign \new_[613]_  = \new_[86484]_  & \new_[86469]_ ;
  assign \new_[614]_  = \new_[86456]_  & \new_[86441]_ ;
  assign \new_[615]_  = \new_[86428]_  & \new_[86413]_ ;
  assign \new_[616]_  = \new_[86400]_  & \new_[86385]_ ;
  assign \new_[617]_  = \new_[86372]_  & \new_[86357]_ ;
  assign \new_[618]_  = \new_[86344]_  & \new_[86329]_ ;
  assign \new_[619]_  = \new_[86316]_  & \new_[86301]_ ;
  assign \new_[620]_  = \new_[86288]_  & \new_[86273]_ ;
  assign \new_[621]_  = \new_[86260]_  & \new_[86245]_ ;
  assign \new_[622]_  = \new_[86232]_  & \new_[86217]_ ;
  assign \new_[623]_  = \new_[86204]_  & \new_[86189]_ ;
  assign \new_[624]_  = \new_[86176]_  & \new_[86161]_ ;
  assign \new_[625]_  = \new_[86148]_  & \new_[86133]_ ;
  assign \new_[626]_  = \new_[86120]_  & \new_[86105]_ ;
  assign \new_[627]_  = \new_[86092]_  & \new_[86077]_ ;
  assign \new_[628]_  = \new_[86064]_  & \new_[86049]_ ;
  assign \new_[629]_  = \new_[86036]_  & \new_[86021]_ ;
  assign \new_[630]_  = \new_[86008]_  & \new_[85993]_ ;
  assign \new_[631]_  = \new_[85980]_  & \new_[85965]_ ;
  assign \new_[632]_  = \new_[85952]_  & \new_[85937]_ ;
  assign \new_[633]_  = \new_[85924]_  & \new_[85909]_ ;
  assign \new_[634]_  = \new_[85896]_  & \new_[85881]_ ;
  assign \new_[635]_  = \new_[85868]_  & \new_[85853]_ ;
  assign \new_[636]_  = \new_[85840]_  & \new_[85825]_ ;
  assign \new_[637]_  = \new_[85812]_  & \new_[85797]_ ;
  assign \new_[638]_  = \new_[85784]_  & \new_[85769]_ ;
  assign \new_[639]_  = \new_[85756]_  & \new_[85741]_ ;
  assign \new_[640]_  = \new_[85728]_  & \new_[85713]_ ;
  assign \new_[641]_  = \new_[85700]_  & \new_[85685]_ ;
  assign \new_[642]_  = \new_[85672]_  & \new_[85657]_ ;
  assign \new_[643]_  = \new_[85644]_  & \new_[85629]_ ;
  assign \new_[644]_  = \new_[85616]_  & \new_[85601]_ ;
  assign \new_[645]_  = \new_[85588]_  & \new_[85573]_ ;
  assign \new_[646]_  = \new_[85560]_  & \new_[85545]_ ;
  assign \new_[647]_  = \new_[85532]_  & \new_[85517]_ ;
  assign \new_[648]_  = \new_[85504]_  & \new_[85489]_ ;
  assign \new_[649]_  = \new_[85476]_  & \new_[85461]_ ;
  assign \new_[650]_  = \new_[85448]_  & \new_[85433]_ ;
  assign \new_[651]_  = \new_[85420]_  & \new_[85405]_ ;
  assign \new_[652]_  = \new_[85392]_  & \new_[85377]_ ;
  assign \new_[653]_  = \new_[85364]_  & \new_[85349]_ ;
  assign \new_[654]_  = \new_[85336]_  & \new_[85321]_ ;
  assign \new_[655]_  = \new_[85308]_  & \new_[85293]_ ;
  assign \new_[656]_  = \new_[85280]_  & \new_[85265]_ ;
  assign \new_[657]_  = \new_[85252]_  & \new_[85237]_ ;
  assign \new_[658]_  = \new_[85224]_  & \new_[85209]_ ;
  assign \new_[659]_  = \new_[85196]_  & \new_[85181]_ ;
  assign \new_[660]_  = \new_[85168]_  & \new_[85153]_ ;
  assign \new_[661]_  = \new_[85140]_  & \new_[85125]_ ;
  assign \new_[662]_  = \new_[85112]_  & \new_[85097]_ ;
  assign \new_[663]_  = \new_[85084]_  & \new_[85069]_ ;
  assign \new_[664]_  = \new_[85056]_  & \new_[85041]_ ;
  assign \new_[665]_  = \new_[85028]_  & \new_[85013]_ ;
  assign \new_[666]_  = \new_[85000]_  & \new_[84985]_ ;
  assign \new_[667]_  = \new_[84972]_  & \new_[84957]_ ;
  assign \new_[668]_  = \new_[84944]_  & \new_[84929]_ ;
  assign \new_[669]_  = \new_[84916]_  & \new_[84901]_ ;
  assign \new_[670]_  = \new_[84888]_  & \new_[84873]_ ;
  assign \new_[671]_  = \new_[84860]_  & \new_[84845]_ ;
  assign \new_[672]_  = \new_[84832]_  & \new_[84817]_ ;
  assign \new_[673]_  = \new_[84804]_  & \new_[84789]_ ;
  assign \new_[674]_  = \new_[84776]_  & \new_[84761]_ ;
  assign \new_[675]_  = \new_[84748]_  & \new_[84733]_ ;
  assign \new_[676]_  = \new_[84720]_  & \new_[84705]_ ;
  assign \new_[677]_  = \new_[84692]_  & \new_[84677]_ ;
  assign \new_[678]_  = \new_[84664]_  & \new_[84649]_ ;
  assign \new_[679]_  = \new_[84636]_  & \new_[84621]_ ;
  assign \new_[680]_  = \new_[84608]_  & \new_[84593]_ ;
  assign \new_[681]_  = \new_[84580]_  & \new_[84565]_ ;
  assign \new_[682]_  = \new_[84552]_  & \new_[84537]_ ;
  assign \new_[683]_  = \new_[84524]_  & \new_[84509]_ ;
  assign \new_[684]_  = \new_[84496]_  & \new_[84481]_ ;
  assign \new_[685]_  = \new_[84468]_  & \new_[84453]_ ;
  assign \new_[686]_  = \new_[84440]_  & \new_[84425]_ ;
  assign \new_[687]_  = \new_[84412]_  & \new_[84397]_ ;
  assign \new_[688]_  = \new_[84384]_  & \new_[84369]_ ;
  assign \new_[689]_  = \new_[84356]_  & \new_[84341]_ ;
  assign \new_[690]_  = \new_[84328]_  & \new_[84313]_ ;
  assign \new_[691]_  = \new_[84300]_  & \new_[84285]_ ;
  assign \new_[692]_  = \new_[84272]_  & \new_[84257]_ ;
  assign \new_[693]_  = \new_[84244]_  & \new_[84229]_ ;
  assign \new_[694]_  = \new_[84216]_  & \new_[84201]_ ;
  assign \new_[695]_  = \new_[84188]_  & \new_[84173]_ ;
  assign \new_[696]_  = \new_[84160]_  & \new_[84145]_ ;
  assign \new_[697]_  = \new_[84132]_  & \new_[84117]_ ;
  assign \new_[698]_  = \new_[84104]_  & \new_[84089]_ ;
  assign \new_[699]_  = \new_[84076]_  & \new_[84061]_ ;
  assign \new_[700]_  = \new_[84048]_  & \new_[84033]_ ;
  assign \new_[701]_  = \new_[84020]_  & \new_[84005]_ ;
  assign \new_[702]_  = \new_[83992]_  & \new_[83977]_ ;
  assign \new_[703]_  = \new_[83964]_  & \new_[83949]_ ;
  assign \new_[704]_  = \new_[83936]_  & \new_[83921]_ ;
  assign \new_[705]_  = \new_[83908]_  & \new_[83893]_ ;
  assign \new_[706]_  = \new_[83880]_  & \new_[83865]_ ;
  assign \new_[707]_  = \new_[83852]_  & \new_[83837]_ ;
  assign \new_[708]_  = \new_[83824]_  & \new_[83809]_ ;
  assign \new_[709]_  = \new_[83796]_  & \new_[83781]_ ;
  assign \new_[710]_  = \new_[83768]_  & \new_[83753]_ ;
  assign \new_[711]_  = \new_[83740]_  & \new_[83725]_ ;
  assign \new_[712]_  = \new_[83712]_  & \new_[83697]_ ;
  assign \new_[713]_  = \new_[83684]_  & \new_[83669]_ ;
  assign \new_[714]_  = \new_[83656]_  & \new_[83641]_ ;
  assign \new_[715]_  = \new_[83628]_  & \new_[83613]_ ;
  assign \new_[716]_  = \new_[83600]_  & \new_[83585]_ ;
  assign \new_[717]_  = \new_[83572]_  & \new_[83557]_ ;
  assign \new_[718]_  = \new_[83544]_  & \new_[83529]_ ;
  assign \new_[719]_  = \new_[83516]_  & \new_[83501]_ ;
  assign \new_[720]_  = \new_[83488]_  & \new_[83473]_ ;
  assign \new_[721]_  = \new_[83460]_  & \new_[83445]_ ;
  assign \new_[722]_  = \new_[83432]_  & \new_[83417]_ ;
  assign \new_[723]_  = \new_[83404]_  & \new_[83389]_ ;
  assign \new_[724]_  = \new_[83376]_  & \new_[83361]_ ;
  assign \new_[725]_  = \new_[83348]_  & \new_[83333]_ ;
  assign \new_[726]_  = \new_[83320]_  & \new_[83305]_ ;
  assign \new_[727]_  = \new_[83292]_  & \new_[83277]_ ;
  assign \new_[728]_  = \new_[83264]_  & \new_[83249]_ ;
  assign \new_[729]_  = \new_[83236]_  & \new_[83221]_ ;
  assign \new_[730]_  = \new_[83208]_  & \new_[83193]_ ;
  assign \new_[731]_  = \new_[83180]_  & \new_[83165]_ ;
  assign \new_[732]_  = \new_[83152]_  & \new_[83137]_ ;
  assign \new_[733]_  = \new_[83124]_  & \new_[83109]_ ;
  assign \new_[734]_  = \new_[83096]_  & \new_[83081]_ ;
  assign \new_[735]_  = \new_[83068]_  & \new_[83053]_ ;
  assign \new_[736]_  = \new_[83040]_  & \new_[83025]_ ;
  assign \new_[737]_  = \new_[83012]_  & \new_[82997]_ ;
  assign \new_[738]_  = \new_[82984]_  & \new_[82969]_ ;
  assign \new_[739]_  = \new_[82956]_  & \new_[82941]_ ;
  assign \new_[740]_  = \new_[82928]_  & \new_[82913]_ ;
  assign \new_[741]_  = \new_[82900]_  & \new_[82885]_ ;
  assign \new_[742]_  = \new_[82872]_  & \new_[82857]_ ;
  assign \new_[743]_  = \new_[82844]_  & \new_[82829]_ ;
  assign \new_[744]_  = \new_[82816]_  & \new_[82801]_ ;
  assign \new_[745]_  = \new_[82788]_  & \new_[82773]_ ;
  assign \new_[746]_  = \new_[82760]_  & \new_[82745]_ ;
  assign \new_[747]_  = \new_[82732]_  & \new_[82717]_ ;
  assign \new_[748]_  = \new_[82704]_  & \new_[82689]_ ;
  assign \new_[749]_  = \new_[82676]_  & \new_[82661]_ ;
  assign \new_[750]_  = \new_[82648]_  & \new_[82633]_ ;
  assign \new_[751]_  = \new_[82620]_  & \new_[82605]_ ;
  assign \new_[752]_  = \new_[82592]_  & \new_[82577]_ ;
  assign \new_[753]_  = \new_[82564]_  & \new_[82549]_ ;
  assign \new_[754]_  = \new_[82536]_  & \new_[82521]_ ;
  assign \new_[755]_  = \new_[82508]_  & \new_[82493]_ ;
  assign \new_[756]_  = \new_[82480]_  & \new_[82465]_ ;
  assign \new_[757]_  = \new_[82452]_  & \new_[82437]_ ;
  assign \new_[758]_  = \new_[82424]_  & \new_[82409]_ ;
  assign \new_[759]_  = \new_[82396]_  & \new_[82381]_ ;
  assign \new_[760]_  = \new_[82368]_  & \new_[82353]_ ;
  assign \new_[761]_  = \new_[82340]_  & \new_[82325]_ ;
  assign \new_[762]_  = \new_[82312]_  & \new_[82297]_ ;
  assign \new_[763]_  = \new_[82284]_  & \new_[82269]_ ;
  assign \new_[764]_  = \new_[82256]_  & \new_[82241]_ ;
  assign \new_[765]_  = \new_[82228]_  & \new_[82213]_ ;
  assign \new_[766]_  = \new_[82200]_  & \new_[82185]_ ;
  assign \new_[767]_  = \new_[82172]_  & \new_[82157]_ ;
  assign \new_[768]_  = \new_[82144]_  & \new_[82129]_ ;
  assign \new_[769]_  = \new_[82116]_  & \new_[82101]_ ;
  assign \new_[770]_  = \new_[82088]_  & \new_[82073]_ ;
  assign \new_[771]_  = \new_[82060]_  & \new_[82045]_ ;
  assign \new_[772]_  = \new_[82032]_  & \new_[82017]_ ;
  assign \new_[773]_  = \new_[82004]_  & \new_[81989]_ ;
  assign \new_[774]_  = \new_[81976]_  & \new_[81961]_ ;
  assign \new_[775]_  = \new_[81948]_  & \new_[81933]_ ;
  assign \new_[776]_  = \new_[81920]_  & \new_[81905]_ ;
  assign \new_[777]_  = \new_[81892]_  & \new_[81877]_ ;
  assign \new_[778]_  = \new_[81864]_  & \new_[81849]_ ;
  assign \new_[779]_  = \new_[81836]_  & \new_[81821]_ ;
  assign \new_[780]_  = \new_[81808]_  & \new_[81793]_ ;
  assign \new_[781]_  = \new_[81780]_  & \new_[81765]_ ;
  assign \new_[782]_  = \new_[81752]_  & \new_[81737]_ ;
  assign \new_[783]_  = \new_[81724]_  & \new_[81709]_ ;
  assign \new_[784]_  = \new_[81696]_  & \new_[81681]_ ;
  assign \new_[785]_  = \new_[81668]_  & \new_[81653]_ ;
  assign \new_[786]_  = \new_[81640]_  & \new_[81625]_ ;
  assign \new_[787]_  = \new_[81612]_  & \new_[81597]_ ;
  assign \new_[788]_  = \new_[81584]_  & \new_[81569]_ ;
  assign \new_[789]_  = \new_[81556]_  & \new_[81541]_ ;
  assign \new_[790]_  = \new_[81528]_  & \new_[81513]_ ;
  assign \new_[791]_  = \new_[81500]_  & \new_[81485]_ ;
  assign \new_[792]_  = \new_[81472]_  & \new_[81457]_ ;
  assign \new_[793]_  = \new_[81444]_  & \new_[81429]_ ;
  assign \new_[794]_  = \new_[81416]_  & \new_[81401]_ ;
  assign \new_[795]_  = \new_[81388]_  & \new_[81373]_ ;
  assign \new_[796]_  = \new_[81360]_  & \new_[81345]_ ;
  assign \new_[797]_  = \new_[81332]_  & \new_[81317]_ ;
  assign \new_[798]_  = \new_[81304]_  & \new_[81289]_ ;
  assign \new_[799]_  = \new_[81276]_  & \new_[81261]_ ;
  assign \new_[800]_  = \new_[81248]_  & \new_[81233]_ ;
  assign \new_[801]_  = \new_[81220]_  & \new_[81205]_ ;
  assign \new_[802]_  = \new_[81192]_  & \new_[81177]_ ;
  assign \new_[803]_  = \new_[81164]_  & \new_[81149]_ ;
  assign \new_[804]_  = \new_[81136]_  & \new_[81121]_ ;
  assign \new_[805]_  = \new_[81108]_  & \new_[81093]_ ;
  assign \new_[806]_  = \new_[81080]_  & \new_[81065]_ ;
  assign \new_[807]_  = \new_[81052]_  & \new_[81037]_ ;
  assign \new_[808]_  = \new_[81024]_  & \new_[81009]_ ;
  assign \new_[809]_  = \new_[80996]_  & \new_[80981]_ ;
  assign \new_[810]_  = \new_[80968]_  & \new_[80953]_ ;
  assign \new_[811]_  = \new_[80940]_  & \new_[80925]_ ;
  assign \new_[812]_  = \new_[80912]_  & \new_[80897]_ ;
  assign \new_[813]_  = \new_[80884]_  & \new_[80869]_ ;
  assign \new_[814]_  = \new_[80856]_  & \new_[80841]_ ;
  assign \new_[815]_  = \new_[80828]_  & \new_[80813]_ ;
  assign \new_[816]_  = \new_[80800]_  & \new_[80785]_ ;
  assign \new_[817]_  = \new_[80772]_  & \new_[80757]_ ;
  assign \new_[818]_  = \new_[80744]_  & \new_[80729]_ ;
  assign \new_[819]_  = \new_[80716]_  & \new_[80701]_ ;
  assign \new_[820]_  = \new_[80688]_  & \new_[80673]_ ;
  assign \new_[821]_  = \new_[80660]_  & \new_[80645]_ ;
  assign \new_[822]_  = \new_[80632]_  & \new_[80617]_ ;
  assign \new_[823]_  = \new_[80604]_  & \new_[80589]_ ;
  assign \new_[824]_  = \new_[80576]_  & \new_[80561]_ ;
  assign \new_[825]_  = \new_[80548]_  & \new_[80533]_ ;
  assign \new_[826]_  = \new_[80520]_  & \new_[80505]_ ;
  assign \new_[827]_  = \new_[80492]_  & \new_[80477]_ ;
  assign \new_[828]_  = \new_[80464]_  & \new_[80449]_ ;
  assign \new_[829]_  = \new_[80436]_  & \new_[80421]_ ;
  assign \new_[830]_  = \new_[80408]_  & \new_[80393]_ ;
  assign \new_[831]_  = \new_[80380]_  & \new_[80365]_ ;
  assign \new_[832]_  = \new_[80352]_  & \new_[80337]_ ;
  assign \new_[833]_  = \new_[80324]_  & \new_[80309]_ ;
  assign \new_[834]_  = \new_[80296]_  & \new_[80281]_ ;
  assign \new_[835]_  = \new_[80268]_  & \new_[80253]_ ;
  assign \new_[836]_  = \new_[80240]_  & \new_[80225]_ ;
  assign \new_[837]_  = \new_[80212]_  & \new_[80197]_ ;
  assign \new_[838]_  = \new_[80184]_  & \new_[80169]_ ;
  assign \new_[839]_  = \new_[80156]_  & \new_[80141]_ ;
  assign \new_[840]_  = \new_[80128]_  & \new_[80113]_ ;
  assign \new_[841]_  = \new_[80100]_  & \new_[80085]_ ;
  assign \new_[842]_  = \new_[80072]_  & \new_[80057]_ ;
  assign \new_[843]_  = \new_[80044]_  & \new_[80029]_ ;
  assign \new_[844]_  = \new_[80016]_  & \new_[80001]_ ;
  assign \new_[845]_  = \new_[79988]_  & \new_[79973]_ ;
  assign \new_[846]_  = \new_[79960]_  & \new_[79945]_ ;
  assign \new_[847]_  = \new_[79932]_  & \new_[79917]_ ;
  assign \new_[848]_  = \new_[79904]_  & \new_[79889]_ ;
  assign \new_[849]_  = \new_[79876]_  & \new_[79861]_ ;
  assign \new_[850]_  = \new_[79848]_  & \new_[79833]_ ;
  assign \new_[851]_  = \new_[79820]_  & \new_[79805]_ ;
  assign \new_[852]_  = \new_[79792]_  & \new_[79777]_ ;
  assign \new_[853]_  = \new_[79764]_  & \new_[79749]_ ;
  assign \new_[854]_  = \new_[79736]_  & \new_[79721]_ ;
  assign \new_[855]_  = \new_[79708]_  & \new_[79693]_ ;
  assign \new_[856]_  = \new_[79680]_  & \new_[79665]_ ;
  assign \new_[857]_  = \new_[79652]_  & \new_[79637]_ ;
  assign \new_[858]_  = \new_[79624]_  & \new_[79609]_ ;
  assign \new_[859]_  = \new_[79596]_  & \new_[79581]_ ;
  assign \new_[860]_  = \new_[79568]_  & \new_[79553]_ ;
  assign \new_[861]_  = \new_[79540]_  & \new_[79525]_ ;
  assign \new_[862]_  = \new_[79512]_  & \new_[79497]_ ;
  assign \new_[863]_  = \new_[79484]_  & \new_[79469]_ ;
  assign \new_[864]_  = \new_[79456]_  & \new_[79441]_ ;
  assign \new_[865]_  = \new_[79428]_  & \new_[79413]_ ;
  assign \new_[866]_  = \new_[79400]_  & \new_[79385]_ ;
  assign \new_[867]_  = \new_[79372]_  & \new_[79357]_ ;
  assign \new_[868]_  = \new_[79344]_  & \new_[79329]_ ;
  assign \new_[869]_  = \new_[79316]_  & \new_[79301]_ ;
  assign \new_[870]_  = \new_[79288]_  & \new_[79273]_ ;
  assign \new_[871]_  = \new_[79260]_  & \new_[79245]_ ;
  assign \new_[872]_  = \new_[79232]_  & \new_[79217]_ ;
  assign \new_[873]_  = \new_[79204]_  & \new_[79189]_ ;
  assign \new_[874]_  = \new_[79176]_  & \new_[79161]_ ;
  assign \new_[875]_  = \new_[79148]_  & \new_[79133]_ ;
  assign \new_[876]_  = \new_[79120]_  & \new_[79105]_ ;
  assign \new_[877]_  = \new_[79092]_  & \new_[79077]_ ;
  assign \new_[878]_  = \new_[79064]_  & \new_[79049]_ ;
  assign \new_[879]_  = \new_[79036]_  & \new_[79021]_ ;
  assign \new_[880]_  = \new_[79008]_  & \new_[78993]_ ;
  assign \new_[881]_  = \new_[78980]_  & \new_[78965]_ ;
  assign \new_[882]_  = \new_[78952]_  & \new_[78937]_ ;
  assign \new_[883]_  = \new_[78924]_  & \new_[78909]_ ;
  assign \new_[884]_  = \new_[78896]_  & \new_[78881]_ ;
  assign \new_[885]_  = \new_[78868]_  & \new_[78853]_ ;
  assign \new_[886]_  = \new_[78840]_  & \new_[78825]_ ;
  assign \new_[887]_  = \new_[78812]_  & \new_[78797]_ ;
  assign \new_[888]_  = \new_[78784]_  & \new_[78769]_ ;
  assign \new_[889]_  = \new_[78756]_  & \new_[78741]_ ;
  assign \new_[890]_  = \new_[78728]_  & \new_[78713]_ ;
  assign \new_[891]_  = \new_[78700]_  & \new_[78685]_ ;
  assign \new_[892]_  = \new_[78672]_  & \new_[78657]_ ;
  assign \new_[893]_  = \new_[78644]_  & \new_[78629]_ ;
  assign \new_[894]_  = \new_[78616]_  & \new_[78601]_ ;
  assign \new_[895]_  = \new_[78588]_  & \new_[78573]_ ;
  assign \new_[896]_  = \new_[78560]_  & \new_[78545]_ ;
  assign \new_[897]_  = \new_[78532]_  & \new_[78517]_ ;
  assign \new_[898]_  = \new_[78504]_  & \new_[78489]_ ;
  assign \new_[899]_  = \new_[78476]_  & \new_[78461]_ ;
  assign \new_[900]_  = \new_[78448]_  & \new_[78433]_ ;
  assign \new_[901]_  = \new_[78420]_  & \new_[78405]_ ;
  assign \new_[902]_  = \new_[78392]_  & \new_[78377]_ ;
  assign \new_[903]_  = \new_[78364]_  & \new_[78349]_ ;
  assign \new_[904]_  = \new_[78336]_  & \new_[78321]_ ;
  assign \new_[905]_  = \new_[78308]_  & \new_[78293]_ ;
  assign \new_[906]_  = \new_[78280]_  & \new_[78265]_ ;
  assign \new_[907]_  = \new_[78252]_  & \new_[78237]_ ;
  assign \new_[908]_  = \new_[78224]_  & \new_[78209]_ ;
  assign \new_[909]_  = \new_[78196]_  & \new_[78181]_ ;
  assign \new_[910]_  = \new_[78168]_  & \new_[78153]_ ;
  assign \new_[911]_  = \new_[78140]_  & \new_[78125]_ ;
  assign \new_[912]_  = \new_[78112]_  & \new_[78097]_ ;
  assign \new_[913]_  = \new_[78084]_  & \new_[78069]_ ;
  assign \new_[914]_  = \new_[78056]_  & \new_[78041]_ ;
  assign \new_[915]_  = \new_[78028]_  & \new_[78013]_ ;
  assign \new_[916]_  = \new_[78000]_  & \new_[77985]_ ;
  assign \new_[917]_  = \new_[77972]_  & \new_[77957]_ ;
  assign \new_[918]_  = \new_[77944]_  & \new_[77929]_ ;
  assign \new_[919]_  = \new_[77916]_  & \new_[77901]_ ;
  assign \new_[920]_  = \new_[77888]_  & \new_[77873]_ ;
  assign \new_[921]_  = \new_[77860]_  & \new_[77845]_ ;
  assign \new_[922]_  = \new_[77832]_  & \new_[77817]_ ;
  assign \new_[923]_  = \new_[77804]_  & \new_[77789]_ ;
  assign \new_[924]_  = \new_[77776]_  & \new_[77761]_ ;
  assign \new_[925]_  = \new_[77748]_  & \new_[77733]_ ;
  assign \new_[926]_  = \new_[77720]_  & \new_[77705]_ ;
  assign \new_[927]_  = \new_[77692]_  & \new_[77677]_ ;
  assign \new_[928]_  = \new_[77664]_  & \new_[77649]_ ;
  assign \new_[929]_  = \new_[77636]_  & \new_[77623]_ ;
  assign \new_[930]_  = \new_[77610]_  & \new_[77597]_ ;
  assign \new_[931]_  = \new_[77584]_  & \new_[77571]_ ;
  assign \new_[932]_  = \new_[77558]_  & \new_[77545]_ ;
  assign \new_[933]_  = \new_[77532]_  & \new_[77519]_ ;
  assign \new_[934]_  = \new_[77506]_  & \new_[77493]_ ;
  assign \new_[935]_  = \new_[77480]_  & \new_[77467]_ ;
  assign \new_[936]_  = \new_[77454]_  & \new_[77441]_ ;
  assign \new_[937]_  = \new_[77428]_  & \new_[77415]_ ;
  assign \new_[938]_  = \new_[77402]_  & \new_[77389]_ ;
  assign \new_[939]_  = \new_[77376]_  & \new_[77363]_ ;
  assign \new_[940]_  = \new_[77350]_  & \new_[77337]_ ;
  assign \new_[941]_  = \new_[77324]_  & \new_[77311]_ ;
  assign \new_[942]_  = \new_[77298]_  & \new_[77285]_ ;
  assign \new_[943]_  = \new_[77272]_  & \new_[77259]_ ;
  assign \new_[944]_  = \new_[77246]_  & \new_[77233]_ ;
  assign \new_[945]_  = \new_[77220]_  & \new_[77207]_ ;
  assign \new_[946]_  = \new_[77194]_  & \new_[77181]_ ;
  assign \new_[947]_  = \new_[77168]_  & \new_[77155]_ ;
  assign \new_[948]_  = \new_[77142]_  & \new_[77129]_ ;
  assign \new_[949]_  = \new_[77116]_  & \new_[77103]_ ;
  assign \new_[950]_  = \new_[77090]_  & \new_[77077]_ ;
  assign \new_[951]_  = \new_[77064]_  & \new_[77051]_ ;
  assign \new_[952]_  = \new_[77038]_  & \new_[77025]_ ;
  assign \new_[953]_  = \new_[77012]_  & \new_[76999]_ ;
  assign \new_[954]_  = \new_[76986]_  & \new_[76973]_ ;
  assign \new_[955]_  = \new_[76960]_  & \new_[76947]_ ;
  assign \new_[956]_  = \new_[76934]_  & \new_[76921]_ ;
  assign \new_[957]_  = \new_[76908]_  & \new_[76895]_ ;
  assign \new_[958]_  = \new_[76882]_  & \new_[76869]_ ;
  assign \new_[959]_  = \new_[76856]_  & \new_[76843]_ ;
  assign \new_[960]_  = \new_[76830]_  & \new_[76817]_ ;
  assign \new_[961]_  = \new_[76804]_  & \new_[76791]_ ;
  assign \new_[962]_  = \new_[76778]_  & \new_[76765]_ ;
  assign \new_[963]_  = \new_[76752]_  & \new_[76739]_ ;
  assign \new_[964]_  = \new_[76726]_  & \new_[76713]_ ;
  assign \new_[965]_  = \new_[76700]_  & \new_[76687]_ ;
  assign \new_[966]_  = \new_[76674]_  & \new_[76661]_ ;
  assign \new_[967]_  = \new_[76648]_  & \new_[76635]_ ;
  assign \new_[968]_  = \new_[76622]_  & \new_[76609]_ ;
  assign \new_[969]_  = \new_[76596]_  & \new_[76583]_ ;
  assign \new_[970]_  = \new_[76570]_  & \new_[76557]_ ;
  assign \new_[971]_  = \new_[76544]_  & \new_[76531]_ ;
  assign \new_[972]_  = \new_[76518]_  & \new_[76505]_ ;
  assign \new_[973]_  = \new_[76492]_  & \new_[76479]_ ;
  assign \new_[974]_  = \new_[76466]_  & \new_[76453]_ ;
  assign \new_[975]_  = \new_[76440]_  & \new_[76427]_ ;
  assign \new_[976]_  = \new_[76414]_  & \new_[76401]_ ;
  assign \new_[977]_  = \new_[76388]_  & \new_[76375]_ ;
  assign \new_[978]_  = \new_[76362]_  & \new_[76349]_ ;
  assign \new_[979]_  = \new_[76336]_  & \new_[76323]_ ;
  assign \new_[980]_  = \new_[76310]_  & \new_[76297]_ ;
  assign \new_[981]_  = \new_[76284]_  & \new_[76271]_ ;
  assign \new_[982]_  = \new_[76258]_  & \new_[76245]_ ;
  assign \new_[983]_  = \new_[76232]_  & \new_[76219]_ ;
  assign \new_[984]_  = \new_[76206]_  & \new_[76193]_ ;
  assign \new_[985]_  = \new_[76180]_  & \new_[76167]_ ;
  assign \new_[986]_  = \new_[76154]_  & \new_[76141]_ ;
  assign \new_[987]_  = \new_[76128]_  & \new_[76115]_ ;
  assign \new_[988]_  = \new_[76102]_  & \new_[76089]_ ;
  assign \new_[989]_  = \new_[76076]_  & \new_[76063]_ ;
  assign \new_[990]_  = \new_[76050]_  & \new_[76037]_ ;
  assign \new_[991]_  = \new_[76024]_  & \new_[76011]_ ;
  assign \new_[992]_  = \new_[75998]_  & \new_[75985]_ ;
  assign \new_[993]_  = \new_[75972]_  & \new_[75959]_ ;
  assign \new_[994]_  = \new_[75946]_  & \new_[75933]_ ;
  assign \new_[995]_  = \new_[75920]_  & \new_[75907]_ ;
  assign \new_[996]_  = \new_[75894]_  & \new_[75881]_ ;
  assign \new_[997]_  = \new_[75868]_  & \new_[75855]_ ;
  assign \new_[998]_  = \new_[75842]_  & \new_[75829]_ ;
  assign \new_[999]_  = \new_[75816]_  & \new_[75803]_ ;
  assign \new_[1000]_  = \new_[75790]_  & \new_[75777]_ ;
  assign \new_[1001]_  = \new_[75764]_  & \new_[75751]_ ;
  assign \new_[1002]_  = \new_[75738]_  & \new_[75725]_ ;
  assign \new_[1003]_  = \new_[75712]_  & \new_[75699]_ ;
  assign \new_[1004]_  = \new_[75686]_  & \new_[75673]_ ;
  assign \new_[1005]_  = \new_[75660]_  & \new_[75647]_ ;
  assign \new_[1006]_  = \new_[75634]_  & \new_[75621]_ ;
  assign \new_[1007]_  = \new_[75608]_  & \new_[75595]_ ;
  assign \new_[1008]_  = \new_[75582]_  & \new_[75569]_ ;
  assign \new_[1009]_  = \new_[75556]_  & \new_[75543]_ ;
  assign \new_[1010]_  = \new_[75530]_  & \new_[75517]_ ;
  assign \new_[1011]_  = \new_[75504]_  & \new_[75491]_ ;
  assign \new_[1012]_  = \new_[75478]_  & \new_[75465]_ ;
  assign \new_[1013]_  = \new_[75452]_  & \new_[75439]_ ;
  assign \new_[1014]_  = \new_[75426]_  & \new_[75413]_ ;
  assign \new_[1015]_  = \new_[75400]_  & \new_[75387]_ ;
  assign \new_[1016]_  = \new_[75374]_  & \new_[75361]_ ;
  assign \new_[1017]_  = \new_[75348]_  & \new_[75335]_ ;
  assign \new_[1018]_  = \new_[75322]_  & \new_[75309]_ ;
  assign \new_[1019]_  = \new_[75296]_  & \new_[75283]_ ;
  assign \new_[1020]_  = \new_[75270]_  & \new_[75257]_ ;
  assign \new_[1021]_  = \new_[75244]_  & \new_[75231]_ ;
  assign \new_[1022]_  = \new_[75218]_  & \new_[75205]_ ;
  assign \new_[1023]_  = \new_[75192]_  & \new_[75179]_ ;
  assign \new_[1024]_  = \new_[75166]_  & \new_[75153]_ ;
  assign \new_[1025]_  = \new_[75140]_  & \new_[75127]_ ;
  assign \new_[1026]_  = \new_[75114]_  & \new_[75101]_ ;
  assign \new_[1027]_  = \new_[75088]_  & \new_[75075]_ ;
  assign \new_[1028]_  = \new_[75062]_  & \new_[75049]_ ;
  assign \new_[1029]_  = \new_[75036]_  & \new_[75023]_ ;
  assign \new_[1030]_  = \new_[75010]_  & \new_[74997]_ ;
  assign \new_[1031]_  = \new_[74984]_  & \new_[74971]_ ;
  assign \new_[1032]_  = \new_[74958]_  & \new_[74945]_ ;
  assign \new_[1033]_  = \new_[74932]_  & \new_[74919]_ ;
  assign \new_[1034]_  = \new_[74906]_  & \new_[74893]_ ;
  assign \new_[1035]_  = \new_[74880]_  & \new_[74867]_ ;
  assign \new_[1036]_  = \new_[74854]_  & \new_[74841]_ ;
  assign \new_[1037]_  = \new_[74828]_  & \new_[74815]_ ;
  assign \new_[1038]_  = \new_[74802]_  & \new_[74789]_ ;
  assign \new_[1039]_  = \new_[74776]_  & \new_[74763]_ ;
  assign \new_[1040]_  = \new_[74750]_  & \new_[74737]_ ;
  assign \new_[1041]_  = \new_[74724]_  & \new_[74711]_ ;
  assign \new_[1042]_  = \new_[74698]_  & \new_[74685]_ ;
  assign \new_[1043]_  = \new_[74672]_  & \new_[74659]_ ;
  assign \new_[1044]_  = \new_[74646]_  & \new_[74633]_ ;
  assign \new_[1045]_  = \new_[74620]_  & \new_[74607]_ ;
  assign \new_[1046]_  = \new_[74594]_  & \new_[74581]_ ;
  assign \new_[1047]_  = \new_[74568]_  & \new_[74555]_ ;
  assign \new_[1048]_  = \new_[74542]_  & \new_[74529]_ ;
  assign \new_[1049]_  = \new_[74516]_  & \new_[74503]_ ;
  assign \new_[1050]_  = \new_[74490]_  & \new_[74477]_ ;
  assign \new_[1051]_  = \new_[74464]_  & \new_[74451]_ ;
  assign \new_[1052]_  = \new_[74438]_  & \new_[74425]_ ;
  assign \new_[1053]_  = \new_[74412]_  & \new_[74399]_ ;
  assign \new_[1054]_  = \new_[74386]_  & \new_[74373]_ ;
  assign \new_[1055]_  = \new_[74360]_  & \new_[74347]_ ;
  assign \new_[1056]_  = \new_[74334]_  & \new_[74321]_ ;
  assign \new_[1057]_  = \new_[74308]_  & \new_[74295]_ ;
  assign \new_[1058]_  = \new_[74282]_  & \new_[74269]_ ;
  assign \new_[1059]_  = \new_[74256]_  & \new_[74243]_ ;
  assign \new_[1060]_  = \new_[74230]_  & \new_[74217]_ ;
  assign \new_[1061]_  = \new_[74204]_  & \new_[74191]_ ;
  assign \new_[1062]_  = \new_[74178]_  & \new_[74165]_ ;
  assign \new_[1063]_  = \new_[74152]_  & \new_[74139]_ ;
  assign \new_[1064]_  = \new_[74126]_  & \new_[74113]_ ;
  assign \new_[1065]_  = \new_[74100]_  & \new_[74087]_ ;
  assign \new_[1066]_  = \new_[74074]_  & \new_[74061]_ ;
  assign \new_[1067]_  = \new_[74048]_  & \new_[74035]_ ;
  assign \new_[1068]_  = \new_[74022]_  & \new_[74009]_ ;
  assign \new_[1069]_  = \new_[73996]_  & \new_[73983]_ ;
  assign \new_[1070]_  = \new_[73970]_  & \new_[73957]_ ;
  assign \new_[1071]_  = \new_[73944]_  & \new_[73931]_ ;
  assign \new_[1072]_  = \new_[73918]_  & \new_[73905]_ ;
  assign \new_[1073]_  = \new_[73892]_  & \new_[73879]_ ;
  assign \new_[1074]_  = \new_[73866]_  & \new_[73853]_ ;
  assign \new_[1075]_  = \new_[73840]_  & \new_[73827]_ ;
  assign \new_[1076]_  = \new_[73814]_  & \new_[73801]_ ;
  assign \new_[1077]_  = \new_[73788]_  & \new_[73775]_ ;
  assign \new_[1078]_  = \new_[73762]_  & \new_[73749]_ ;
  assign \new_[1079]_  = \new_[73736]_  & \new_[73723]_ ;
  assign \new_[1080]_  = \new_[73710]_  & \new_[73697]_ ;
  assign \new_[1081]_  = \new_[73684]_  & \new_[73671]_ ;
  assign \new_[1082]_  = \new_[73658]_  & \new_[73645]_ ;
  assign \new_[1083]_  = \new_[73632]_  & \new_[73619]_ ;
  assign \new_[1084]_  = \new_[73606]_  & \new_[73593]_ ;
  assign \new_[1085]_  = \new_[73580]_  & \new_[73567]_ ;
  assign \new_[1086]_  = \new_[73554]_  & \new_[73541]_ ;
  assign \new_[1087]_  = \new_[73528]_  & \new_[73515]_ ;
  assign \new_[1088]_  = \new_[73502]_  & \new_[73489]_ ;
  assign \new_[1089]_  = \new_[73476]_  & \new_[73463]_ ;
  assign \new_[1090]_  = \new_[73450]_  & \new_[73437]_ ;
  assign \new_[1091]_  = \new_[73424]_  & \new_[73411]_ ;
  assign \new_[1092]_  = \new_[73398]_  & \new_[73385]_ ;
  assign \new_[1093]_  = \new_[73372]_  & \new_[73359]_ ;
  assign \new_[1094]_  = \new_[73346]_  & \new_[73333]_ ;
  assign \new_[1095]_  = \new_[73320]_  & \new_[73307]_ ;
  assign \new_[1096]_  = \new_[73294]_  & \new_[73281]_ ;
  assign \new_[1097]_  = \new_[73268]_  & \new_[73255]_ ;
  assign \new_[1098]_  = \new_[73242]_  & \new_[73229]_ ;
  assign \new_[1099]_  = \new_[73216]_  & \new_[73203]_ ;
  assign \new_[1100]_  = \new_[73190]_  & \new_[73177]_ ;
  assign \new_[1101]_  = \new_[73164]_  & \new_[73151]_ ;
  assign \new_[1102]_  = \new_[73138]_  & \new_[73125]_ ;
  assign \new_[1103]_  = \new_[73112]_  & \new_[73099]_ ;
  assign \new_[1104]_  = \new_[73086]_  & \new_[73073]_ ;
  assign \new_[1105]_  = \new_[73060]_  & \new_[73047]_ ;
  assign \new_[1106]_  = \new_[73034]_  & \new_[73021]_ ;
  assign \new_[1107]_  = \new_[73008]_  & \new_[72995]_ ;
  assign \new_[1108]_  = \new_[72982]_  & \new_[72969]_ ;
  assign \new_[1109]_  = \new_[72956]_  & \new_[72943]_ ;
  assign \new_[1110]_  = \new_[72930]_  & \new_[72917]_ ;
  assign \new_[1111]_  = \new_[72904]_  & \new_[72891]_ ;
  assign \new_[1112]_  = \new_[72878]_  & \new_[72865]_ ;
  assign \new_[1113]_  = \new_[72852]_  & \new_[72839]_ ;
  assign \new_[1114]_  = \new_[72826]_  & \new_[72813]_ ;
  assign \new_[1115]_  = \new_[72800]_  & \new_[72787]_ ;
  assign \new_[1116]_  = \new_[72774]_  & \new_[72761]_ ;
  assign \new_[1117]_  = \new_[72748]_  & \new_[72735]_ ;
  assign \new_[1118]_  = \new_[72722]_  & \new_[72709]_ ;
  assign \new_[1119]_  = \new_[72696]_  & \new_[72683]_ ;
  assign \new_[1120]_  = \new_[72670]_  & \new_[72657]_ ;
  assign \new_[1121]_  = \new_[72644]_  & \new_[72631]_ ;
  assign \new_[1122]_  = \new_[72618]_  & \new_[72605]_ ;
  assign \new_[1123]_  = \new_[72592]_  & \new_[72579]_ ;
  assign \new_[1124]_  = \new_[72566]_  & \new_[72553]_ ;
  assign \new_[1125]_  = \new_[72540]_  & \new_[72527]_ ;
  assign \new_[1126]_  = \new_[72514]_  & \new_[72501]_ ;
  assign \new_[1127]_  = \new_[72488]_  & \new_[72475]_ ;
  assign \new_[1128]_  = \new_[72462]_  & \new_[72449]_ ;
  assign \new_[1129]_  = \new_[72436]_  & \new_[72423]_ ;
  assign \new_[1130]_  = \new_[72410]_  & \new_[72397]_ ;
  assign \new_[1131]_  = \new_[72384]_  & \new_[72371]_ ;
  assign \new_[1132]_  = \new_[72358]_  & \new_[72345]_ ;
  assign \new_[1133]_  = \new_[72332]_  & \new_[72319]_ ;
  assign \new_[1134]_  = \new_[72306]_  & \new_[72293]_ ;
  assign \new_[1135]_  = \new_[72280]_  & \new_[72267]_ ;
  assign \new_[1136]_  = \new_[72254]_  & \new_[72241]_ ;
  assign \new_[1137]_  = \new_[72228]_  & \new_[72215]_ ;
  assign \new_[1138]_  = \new_[72202]_  & \new_[72189]_ ;
  assign \new_[1139]_  = \new_[72176]_  & \new_[72163]_ ;
  assign \new_[1140]_  = \new_[72150]_  & \new_[72137]_ ;
  assign \new_[1141]_  = \new_[72124]_  & \new_[72111]_ ;
  assign \new_[1142]_  = \new_[72098]_  & \new_[72085]_ ;
  assign \new_[1143]_  = \new_[72072]_  & \new_[72059]_ ;
  assign \new_[1144]_  = \new_[72046]_  & \new_[72033]_ ;
  assign \new_[1145]_  = \new_[72020]_  & \new_[72007]_ ;
  assign \new_[1146]_  = \new_[71994]_  & \new_[71981]_ ;
  assign \new_[1147]_  = \new_[71968]_  & \new_[71955]_ ;
  assign \new_[1148]_  = \new_[71942]_  & \new_[71929]_ ;
  assign \new_[1149]_  = \new_[71916]_  & \new_[71903]_ ;
  assign \new_[1150]_  = \new_[71890]_  & \new_[71877]_ ;
  assign \new_[1151]_  = \new_[71864]_  & \new_[71851]_ ;
  assign \new_[1152]_  = \new_[71838]_  & \new_[71825]_ ;
  assign \new_[1153]_  = \new_[71812]_  & \new_[71799]_ ;
  assign \new_[1154]_  = \new_[71786]_  & \new_[71773]_ ;
  assign \new_[1155]_  = \new_[71760]_  & \new_[71747]_ ;
  assign \new_[1156]_  = \new_[71734]_  & \new_[71721]_ ;
  assign \new_[1157]_  = \new_[71708]_  & \new_[71695]_ ;
  assign \new_[1158]_  = \new_[71682]_  & \new_[71669]_ ;
  assign \new_[1159]_  = \new_[71656]_  & \new_[71643]_ ;
  assign \new_[1160]_  = \new_[71630]_  & \new_[71617]_ ;
  assign \new_[1161]_  = \new_[71604]_  & \new_[71591]_ ;
  assign \new_[1162]_  = \new_[71578]_  & \new_[71565]_ ;
  assign \new_[1163]_  = \new_[71552]_  & \new_[71539]_ ;
  assign \new_[1164]_  = \new_[71526]_  & \new_[71513]_ ;
  assign \new_[1165]_  = \new_[71500]_  & \new_[71487]_ ;
  assign \new_[1166]_  = \new_[71474]_  & \new_[71461]_ ;
  assign \new_[1167]_  = \new_[71448]_  & \new_[71435]_ ;
  assign \new_[1168]_  = \new_[71422]_  & \new_[71409]_ ;
  assign \new_[1169]_  = \new_[71396]_  & \new_[71383]_ ;
  assign \new_[1170]_  = \new_[71370]_  & \new_[71357]_ ;
  assign \new_[1171]_  = \new_[71344]_  & \new_[71331]_ ;
  assign \new_[1172]_  = \new_[71318]_  & \new_[71305]_ ;
  assign \new_[1173]_  = \new_[71292]_  & \new_[71279]_ ;
  assign \new_[1174]_  = \new_[71266]_  & \new_[71253]_ ;
  assign \new_[1175]_  = \new_[71240]_  & \new_[71227]_ ;
  assign \new_[1176]_  = \new_[71214]_  & \new_[71201]_ ;
  assign \new_[1177]_  = \new_[71188]_  & \new_[71175]_ ;
  assign \new_[1178]_  = \new_[71162]_  & \new_[71149]_ ;
  assign \new_[1179]_  = \new_[71136]_  & \new_[71123]_ ;
  assign \new_[1180]_  = \new_[71110]_  & \new_[71097]_ ;
  assign \new_[1181]_  = \new_[71084]_  & \new_[71071]_ ;
  assign \new_[1182]_  = \new_[71058]_  & \new_[71045]_ ;
  assign \new_[1183]_  = \new_[71032]_  & \new_[71019]_ ;
  assign \new_[1184]_  = \new_[71006]_  & \new_[70993]_ ;
  assign \new_[1185]_  = \new_[70980]_  & \new_[70967]_ ;
  assign \new_[1186]_  = \new_[70954]_  & \new_[70941]_ ;
  assign \new_[1187]_  = \new_[70928]_  & \new_[70915]_ ;
  assign \new_[1188]_  = \new_[70902]_  & \new_[70889]_ ;
  assign \new_[1189]_  = \new_[70876]_  & \new_[70863]_ ;
  assign \new_[1190]_  = \new_[70850]_  & \new_[70837]_ ;
  assign \new_[1191]_  = \new_[70824]_  & \new_[70811]_ ;
  assign \new_[1192]_  = \new_[70798]_  & \new_[70785]_ ;
  assign \new_[1193]_  = \new_[70772]_  & \new_[70759]_ ;
  assign \new_[1194]_  = \new_[70746]_  & \new_[70733]_ ;
  assign \new_[1195]_  = \new_[70720]_  & \new_[70707]_ ;
  assign \new_[1196]_  = \new_[70694]_  & \new_[70681]_ ;
  assign \new_[1197]_  = \new_[70668]_  & \new_[70655]_ ;
  assign \new_[1198]_  = \new_[70642]_  & \new_[70629]_ ;
  assign \new_[1199]_  = \new_[70616]_  & \new_[70603]_ ;
  assign \new_[1200]_  = \new_[70590]_  & \new_[70577]_ ;
  assign \new_[1201]_  = \new_[70564]_  & \new_[70551]_ ;
  assign \new_[1202]_  = \new_[70538]_  & \new_[70525]_ ;
  assign \new_[1203]_  = \new_[70512]_  & \new_[70499]_ ;
  assign \new_[1204]_  = \new_[70486]_  & \new_[70473]_ ;
  assign \new_[1205]_  = \new_[70460]_  & \new_[70447]_ ;
  assign \new_[1206]_  = \new_[70434]_  & \new_[70421]_ ;
  assign \new_[1207]_  = \new_[70408]_  & \new_[70395]_ ;
  assign \new_[1208]_  = \new_[70382]_  & \new_[70369]_ ;
  assign \new_[1209]_  = \new_[70356]_  & \new_[70343]_ ;
  assign \new_[1210]_  = \new_[70330]_  & \new_[70317]_ ;
  assign \new_[1211]_  = \new_[70304]_  & \new_[70291]_ ;
  assign \new_[1212]_  = \new_[70278]_  & \new_[70265]_ ;
  assign \new_[1213]_  = \new_[70252]_  & \new_[70239]_ ;
  assign \new_[1214]_  = \new_[70226]_  & \new_[70213]_ ;
  assign \new_[1215]_  = \new_[70200]_  & \new_[70187]_ ;
  assign \new_[1216]_  = \new_[70174]_  & \new_[70161]_ ;
  assign \new_[1217]_  = \new_[70148]_  & \new_[70135]_ ;
  assign \new_[1218]_  = \new_[70122]_  & \new_[70109]_ ;
  assign \new_[1219]_  = \new_[70096]_  & \new_[70083]_ ;
  assign \new_[1220]_  = \new_[70070]_  & \new_[70057]_ ;
  assign \new_[1221]_  = \new_[70044]_  & \new_[70031]_ ;
  assign \new_[1222]_  = \new_[70018]_  & \new_[70005]_ ;
  assign \new_[1223]_  = \new_[69992]_  & \new_[69979]_ ;
  assign \new_[1224]_  = \new_[69966]_  & \new_[69953]_ ;
  assign \new_[1225]_  = \new_[69940]_  & \new_[69927]_ ;
  assign \new_[1226]_  = \new_[69914]_  & \new_[69901]_ ;
  assign \new_[1227]_  = \new_[69888]_  & \new_[69875]_ ;
  assign \new_[1228]_  = \new_[69862]_  & \new_[69849]_ ;
  assign \new_[1229]_  = \new_[69836]_  & \new_[69823]_ ;
  assign \new_[1230]_  = \new_[69810]_  & \new_[69797]_ ;
  assign \new_[1231]_  = \new_[69784]_  & \new_[69771]_ ;
  assign \new_[1232]_  = \new_[69758]_  & \new_[69745]_ ;
  assign \new_[1233]_  = \new_[69732]_  & \new_[69719]_ ;
  assign \new_[1234]_  = \new_[69706]_  & \new_[69693]_ ;
  assign \new_[1235]_  = \new_[69680]_  & \new_[69667]_ ;
  assign \new_[1236]_  = \new_[69654]_  & \new_[69641]_ ;
  assign \new_[1237]_  = \new_[69628]_  & \new_[69615]_ ;
  assign \new_[1238]_  = \new_[69602]_  & \new_[69589]_ ;
  assign \new_[1239]_  = \new_[69576]_  & \new_[69563]_ ;
  assign \new_[1240]_  = \new_[69550]_  & \new_[69537]_ ;
  assign \new_[1241]_  = \new_[69524]_  & \new_[69511]_ ;
  assign \new_[1242]_  = \new_[69498]_  & \new_[69485]_ ;
  assign \new_[1243]_  = \new_[69472]_  & \new_[69459]_ ;
  assign \new_[1244]_  = \new_[69446]_  & \new_[69433]_ ;
  assign \new_[1245]_  = \new_[69420]_  & \new_[69407]_ ;
  assign \new_[1246]_  = \new_[69394]_  & \new_[69381]_ ;
  assign \new_[1247]_  = \new_[69368]_  & \new_[69355]_ ;
  assign \new_[1248]_  = \new_[69342]_  & \new_[69329]_ ;
  assign \new_[1249]_  = \new_[69316]_  & \new_[69303]_ ;
  assign \new_[1250]_  = \new_[69290]_  & \new_[69277]_ ;
  assign \new_[1251]_  = \new_[69264]_  & \new_[69251]_ ;
  assign \new_[1252]_  = \new_[69238]_  & \new_[69225]_ ;
  assign \new_[1253]_  = \new_[69212]_  & \new_[69199]_ ;
  assign \new_[1254]_  = \new_[69186]_  & \new_[69173]_ ;
  assign \new_[1255]_  = \new_[69160]_  & \new_[69147]_ ;
  assign \new_[1256]_  = \new_[69134]_  & \new_[69121]_ ;
  assign \new_[1257]_  = \new_[69108]_  & \new_[69095]_ ;
  assign \new_[1258]_  = \new_[69082]_  & \new_[69069]_ ;
  assign \new_[1259]_  = \new_[69056]_  & \new_[69043]_ ;
  assign \new_[1260]_  = \new_[69030]_  & \new_[69017]_ ;
  assign \new_[1261]_  = \new_[69004]_  & \new_[68991]_ ;
  assign \new_[1262]_  = \new_[68978]_  & \new_[68965]_ ;
  assign \new_[1263]_  = \new_[68952]_  & \new_[68939]_ ;
  assign \new_[1264]_  = \new_[68926]_  & \new_[68913]_ ;
  assign \new_[1265]_  = \new_[68900]_  & \new_[68887]_ ;
  assign \new_[1266]_  = \new_[68874]_  & \new_[68861]_ ;
  assign \new_[1267]_  = \new_[68848]_  & \new_[68835]_ ;
  assign \new_[1268]_  = \new_[68822]_  & \new_[68809]_ ;
  assign \new_[1269]_  = \new_[68796]_  & \new_[68783]_ ;
  assign \new_[1270]_  = \new_[68770]_  & \new_[68757]_ ;
  assign \new_[1271]_  = \new_[68744]_  & \new_[68731]_ ;
  assign \new_[1272]_  = \new_[68718]_  & \new_[68705]_ ;
  assign \new_[1273]_  = \new_[68692]_  & \new_[68679]_ ;
  assign \new_[1274]_  = \new_[68666]_  & \new_[68653]_ ;
  assign \new_[1275]_  = \new_[68640]_  & \new_[68627]_ ;
  assign \new_[1276]_  = \new_[68614]_  & \new_[68601]_ ;
  assign \new_[1277]_  = \new_[68588]_  & \new_[68575]_ ;
  assign \new_[1278]_  = \new_[68562]_  & \new_[68549]_ ;
  assign \new_[1279]_  = \new_[68536]_  & \new_[68523]_ ;
  assign \new_[1280]_  = \new_[68510]_  & \new_[68497]_ ;
  assign \new_[1281]_  = \new_[68484]_  & \new_[68471]_ ;
  assign \new_[1282]_  = \new_[68458]_  & \new_[68445]_ ;
  assign \new_[1283]_  = \new_[68432]_  & \new_[68419]_ ;
  assign \new_[1284]_  = \new_[68406]_  & \new_[68393]_ ;
  assign \new_[1285]_  = \new_[68380]_  & \new_[68367]_ ;
  assign \new_[1286]_  = \new_[68354]_  & \new_[68341]_ ;
  assign \new_[1287]_  = \new_[68328]_  & \new_[68315]_ ;
  assign \new_[1288]_  = \new_[68302]_  & \new_[68289]_ ;
  assign \new_[1289]_  = \new_[68276]_  & \new_[68263]_ ;
  assign \new_[1290]_  = \new_[68250]_  & \new_[68237]_ ;
  assign \new_[1291]_  = \new_[68224]_  & \new_[68211]_ ;
  assign \new_[1292]_  = \new_[68198]_  & \new_[68185]_ ;
  assign \new_[1293]_  = \new_[68172]_  & \new_[68159]_ ;
  assign \new_[1294]_  = \new_[68146]_  & \new_[68133]_ ;
  assign \new_[1295]_  = \new_[68120]_  & \new_[68107]_ ;
  assign \new_[1296]_  = \new_[68094]_  & \new_[68081]_ ;
  assign \new_[1297]_  = \new_[68068]_  & \new_[68055]_ ;
  assign \new_[1298]_  = \new_[68042]_  & \new_[68029]_ ;
  assign \new_[1299]_  = \new_[68016]_  & \new_[68003]_ ;
  assign \new_[1300]_  = \new_[67990]_  & \new_[67977]_ ;
  assign \new_[1301]_  = \new_[67964]_  & \new_[67951]_ ;
  assign \new_[1302]_  = \new_[67938]_  & \new_[67925]_ ;
  assign \new_[1303]_  = \new_[67912]_  & \new_[67899]_ ;
  assign \new_[1304]_  = \new_[67886]_  & \new_[67873]_ ;
  assign \new_[1305]_  = \new_[67860]_  & \new_[67847]_ ;
  assign \new_[1306]_  = \new_[67834]_  & \new_[67821]_ ;
  assign \new_[1307]_  = \new_[67808]_  & \new_[67795]_ ;
  assign \new_[1308]_  = \new_[67782]_  & \new_[67769]_ ;
  assign \new_[1309]_  = \new_[67756]_  & \new_[67743]_ ;
  assign \new_[1310]_  = \new_[67730]_  & \new_[67717]_ ;
  assign \new_[1311]_  = \new_[67704]_  & \new_[67691]_ ;
  assign \new_[1312]_  = \new_[67678]_  & \new_[67665]_ ;
  assign \new_[1313]_  = \new_[67652]_  & \new_[67639]_ ;
  assign \new_[1314]_  = \new_[67626]_  & \new_[67613]_ ;
  assign \new_[1315]_  = \new_[67600]_  & \new_[67587]_ ;
  assign \new_[1316]_  = \new_[67574]_  & \new_[67561]_ ;
  assign \new_[1317]_  = \new_[67548]_  & \new_[67535]_ ;
  assign \new_[1318]_  = \new_[67522]_  & \new_[67509]_ ;
  assign \new_[1319]_  = \new_[67496]_  & \new_[67483]_ ;
  assign \new_[1320]_  = \new_[67470]_  & \new_[67457]_ ;
  assign \new_[1321]_  = \new_[67444]_  & \new_[67431]_ ;
  assign \new_[1322]_  = \new_[67418]_  & \new_[67405]_ ;
  assign \new_[1323]_  = \new_[67392]_  & \new_[67379]_ ;
  assign \new_[1324]_  = \new_[67366]_  & \new_[67353]_ ;
  assign \new_[1325]_  = \new_[67340]_  & \new_[67327]_ ;
  assign \new_[1326]_  = \new_[67314]_  & \new_[67301]_ ;
  assign \new_[1327]_  = \new_[67288]_  & \new_[67275]_ ;
  assign \new_[1328]_  = \new_[67262]_  & \new_[67249]_ ;
  assign \new_[1329]_  = \new_[67236]_  & \new_[67223]_ ;
  assign \new_[1330]_  = \new_[67210]_  & \new_[67197]_ ;
  assign \new_[1331]_  = \new_[67184]_  & \new_[67171]_ ;
  assign \new_[1332]_  = \new_[67158]_  & \new_[67145]_ ;
  assign \new_[1333]_  = \new_[67132]_  & \new_[67119]_ ;
  assign \new_[1334]_  = \new_[67106]_  & \new_[67093]_ ;
  assign \new_[1335]_  = \new_[67080]_  & \new_[67067]_ ;
  assign \new_[1336]_  = \new_[67054]_  & \new_[67041]_ ;
  assign \new_[1337]_  = \new_[67028]_  & \new_[67015]_ ;
  assign \new_[1338]_  = \new_[67002]_  & \new_[66989]_ ;
  assign \new_[1339]_  = \new_[66976]_  & \new_[66963]_ ;
  assign \new_[1340]_  = \new_[66950]_  & \new_[66937]_ ;
  assign \new_[1341]_  = \new_[66924]_  & \new_[66911]_ ;
  assign \new_[1342]_  = \new_[66898]_  & \new_[66885]_ ;
  assign \new_[1343]_  = \new_[66872]_  & \new_[66859]_ ;
  assign \new_[1344]_  = \new_[66846]_  & \new_[66833]_ ;
  assign \new_[1345]_  = \new_[66820]_  & \new_[66807]_ ;
  assign \new_[1346]_  = \new_[66794]_  & \new_[66781]_ ;
  assign \new_[1347]_  = \new_[66768]_  & \new_[66755]_ ;
  assign \new_[1348]_  = \new_[66742]_  & \new_[66729]_ ;
  assign \new_[1349]_  = \new_[66716]_  & \new_[66703]_ ;
  assign \new_[1350]_  = \new_[66690]_  & \new_[66677]_ ;
  assign \new_[1351]_  = \new_[66664]_  & \new_[66651]_ ;
  assign \new_[1352]_  = \new_[66638]_  & \new_[66625]_ ;
  assign \new_[1353]_  = \new_[66612]_  & \new_[66599]_ ;
  assign \new_[1354]_  = \new_[66586]_  & \new_[66573]_ ;
  assign \new_[1355]_  = \new_[66560]_  & \new_[66547]_ ;
  assign \new_[1356]_  = \new_[66534]_  & \new_[66521]_ ;
  assign \new_[1357]_  = \new_[66508]_  & \new_[66495]_ ;
  assign \new_[1358]_  = \new_[66482]_  & \new_[66469]_ ;
  assign \new_[1359]_  = \new_[66456]_  & \new_[66443]_ ;
  assign \new_[1360]_  = \new_[66430]_  & \new_[66417]_ ;
  assign \new_[1361]_  = \new_[66404]_  & \new_[66391]_ ;
  assign \new_[1362]_  = \new_[66378]_  & \new_[66365]_ ;
  assign \new_[1363]_  = \new_[66352]_  & \new_[66339]_ ;
  assign \new_[1364]_  = \new_[66326]_  & \new_[66313]_ ;
  assign \new_[1365]_  = \new_[66300]_  & \new_[66287]_ ;
  assign \new_[1366]_  = \new_[66274]_  & \new_[66261]_ ;
  assign \new_[1367]_  = \new_[66248]_  & \new_[66235]_ ;
  assign \new_[1368]_  = \new_[66222]_  & \new_[66209]_ ;
  assign \new_[1369]_  = \new_[66196]_  & \new_[66183]_ ;
  assign \new_[1370]_  = \new_[66170]_  & \new_[66157]_ ;
  assign \new_[1371]_  = \new_[66144]_  & \new_[66131]_ ;
  assign \new_[1372]_  = \new_[66118]_  & \new_[66105]_ ;
  assign \new_[1373]_  = \new_[66092]_  & \new_[66079]_ ;
  assign \new_[1374]_  = \new_[66066]_  & \new_[66053]_ ;
  assign \new_[1375]_  = \new_[66040]_  & \new_[66027]_ ;
  assign \new_[1376]_  = \new_[66014]_  & \new_[66001]_ ;
  assign \new_[1377]_  = \new_[65988]_  & \new_[65975]_ ;
  assign \new_[1378]_  = \new_[65962]_  & \new_[65949]_ ;
  assign \new_[1379]_  = \new_[65936]_  & \new_[65923]_ ;
  assign \new_[1380]_  = \new_[65910]_  & \new_[65897]_ ;
  assign \new_[1381]_  = \new_[65884]_  & \new_[65871]_ ;
  assign \new_[1382]_  = \new_[65858]_  & \new_[65845]_ ;
  assign \new_[1383]_  = \new_[65832]_  & \new_[65819]_ ;
  assign \new_[1384]_  = \new_[65806]_  & \new_[65793]_ ;
  assign \new_[1385]_  = \new_[65780]_  & \new_[65767]_ ;
  assign \new_[1386]_  = \new_[65754]_  & \new_[65741]_ ;
  assign \new_[1387]_  = \new_[65728]_  & \new_[65715]_ ;
  assign \new_[1388]_  = \new_[65702]_  & \new_[65689]_ ;
  assign \new_[1389]_  = \new_[65676]_  & \new_[65663]_ ;
  assign \new_[1390]_  = \new_[65650]_  & \new_[65637]_ ;
  assign \new_[1391]_  = \new_[65624]_  & \new_[65611]_ ;
  assign \new_[1392]_  = \new_[65598]_  & \new_[65585]_ ;
  assign \new_[1393]_  = \new_[65572]_  & \new_[65559]_ ;
  assign \new_[1394]_  = \new_[65546]_  & \new_[65533]_ ;
  assign \new_[1395]_  = \new_[65520]_  & \new_[65507]_ ;
  assign \new_[1396]_  = \new_[65494]_  & \new_[65481]_ ;
  assign \new_[1397]_  = \new_[65468]_  & \new_[65455]_ ;
  assign \new_[1398]_  = \new_[65442]_  & \new_[65429]_ ;
  assign \new_[1399]_  = \new_[65416]_  & \new_[65403]_ ;
  assign \new_[1400]_  = \new_[65390]_  & \new_[65377]_ ;
  assign \new_[1401]_  = \new_[65364]_  & \new_[65351]_ ;
  assign \new_[1402]_  = \new_[65338]_  & \new_[65325]_ ;
  assign \new_[1403]_  = \new_[65312]_  & \new_[65299]_ ;
  assign \new_[1404]_  = \new_[65286]_  & \new_[65273]_ ;
  assign \new_[1405]_  = \new_[65260]_  & \new_[65247]_ ;
  assign \new_[1406]_  = \new_[65234]_  & \new_[65221]_ ;
  assign \new_[1407]_  = \new_[65208]_  & \new_[65195]_ ;
  assign \new_[1408]_  = \new_[65182]_  & \new_[65169]_ ;
  assign \new_[1409]_  = \new_[65156]_  & \new_[65143]_ ;
  assign \new_[1410]_  = \new_[65130]_  & \new_[65117]_ ;
  assign \new_[1411]_  = \new_[65104]_  & \new_[65091]_ ;
  assign \new_[1412]_  = \new_[65078]_  & \new_[65065]_ ;
  assign \new_[1413]_  = \new_[65052]_  & \new_[65039]_ ;
  assign \new_[1414]_  = \new_[65026]_  & \new_[65013]_ ;
  assign \new_[1415]_  = \new_[65000]_  & \new_[64987]_ ;
  assign \new_[1416]_  = \new_[64974]_  & \new_[64961]_ ;
  assign \new_[1417]_  = \new_[64948]_  & \new_[64935]_ ;
  assign \new_[1418]_  = \new_[64922]_  & \new_[64909]_ ;
  assign \new_[1419]_  = \new_[64896]_  & \new_[64883]_ ;
  assign \new_[1420]_  = \new_[64870]_  & \new_[64857]_ ;
  assign \new_[1421]_  = \new_[64844]_  & \new_[64831]_ ;
  assign \new_[1422]_  = \new_[64818]_  & \new_[64805]_ ;
  assign \new_[1423]_  = \new_[64792]_  & \new_[64779]_ ;
  assign \new_[1424]_  = \new_[64766]_  & \new_[64753]_ ;
  assign \new_[1425]_  = \new_[64740]_  & \new_[64727]_ ;
  assign \new_[1426]_  = \new_[64714]_  & \new_[64701]_ ;
  assign \new_[1427]_  = \new_[64688]_  & \new_[64675]_ ;
  assign \new_[1428]_  = \new_[64662]_  & \new_[64649]_ ;
  assign \new_[1429]_  = \new_[64636]_  & \new_[64623]_ ;
  assign \new_[1430]_  = \new_[64610]_  & \new_[64597]_ ;
  assign \new_[1431]_  = \new_[64584]_  & \new_[64571]_ ;
  assign \new_[1432]_  = \new_[64558]_  & \new_[64545]_ ;
  assign \new_[1433]_  = \new_[64532]_  & \new_[64519]_ ;
  assign \new_[1434]_  = \new_[64506]_  & \new_[64493]_ ;
  assign \new_[1435]_  = \new_[64480]_  & \new_[64467]_ ;
  assign \new_[1436]_  = \new_[64454]_  & \new_[64441]_ ;
  assign \new_[1437]_  = \new_[64428]_  & \new_[64415]_ ;
  assign \new_[1438]_  = \new_[64402]_  & \new_[64389]_ ;
  assign \new_[1439]_  = \new_[64376]_  & \new_[64363]_ ;
  assign \new_[1440]_  = \new_[64350]_  & \new_[64337]_ ;
  assign \new_[1441]_  = \new_[64324]_  & \new_[64311]_ ;
  assign \new_[1442]_  = \new_[64298]_  & \new_[64285]_ ;
  assign \new_[1443]_  = \new_[64272]_  & \new_[64259]_ ;
  assign \new_[1444]_  = \new_[64246]_  & \new_[64233]_ ;
  assign \new_[1445]_  = \new_[64220]_  & \new_[64207]_ ;
  assign \new_[1446]_  = \new_[64194]_  & \new_[64181]_ ;
  assign \new_[1447]_  = \new_[64168]_  & \new_[64155]_ ;
  assign \new_[1448]_  = \new_[64142]_  & \new_[64129]_ ;
  assign \new_[1449]_  = \new_[64116]_  & \new_[64103]_ ;
  assign \new_[1450]_  = \new_[64090]_  & \new_[64077]_ ;
  assign \new_[1451]_  = \new_[64064]_  & \new_[64051]_ ;
  assign \new_[1452]_  = \new_[64038]_  & \new_[64025]_ ;
  assign \new_[1453]_  = \new_[64012]_  & \new_[63999]_ ;
  assign \new_[1454]_  = \new_[63986]_  & \new_[63973]_ ;
  assign \new_[1455]_  = \new_[63960]_  & \new_[63947]_ ;
  assign \new_[1456]_  = \new_[63934]_  & \new_[63921]_ ;
  assign \new_[1457]_  = \new_[63908]_  & \new_[63895]_ ;
  assign \new_[1458]_  = \new_[63882]_  & \new_[63869]_ ;
  assign \new_[1459]_  = \new_[63856]_  & \new_[63843]_ ;
  assign \new_[1460]_  = \new_[63830]_  & \new_[63817]_ ;
  assign \new_[1461]_  = \new_[63804]_  & \new_[63791]_ ;
  assign \new_[1462]_  = \new_[63778]_  & \new_[63765]_ ;
  assign \new_[1463]_  = \new_[63752]_  & \new_[63739]_ ;
  assign \new_[1464]_  = \new_[63726]_  & \new_[63713]_ ;
  assign \new_[1465]_  = \new_[63700]_  & \new_[63687]_ ;
  assign \new_[1466]_  = \new_[63674]_  & \new_[63661]_ ;
  assign \new_[1467]_  = \new_[63648]_  & \new_[63635]_ ;
  assign \new_[1468]_  = \new_[63622]_  & \new_[63609]_ ;
  assign \new_[1469]_  = \new_[63596]_  & \new_[63583]_ ;
  assign \new_[1470]_  = \new_[63570]_  & \new_[63557]_ ;
  assign \new_[1471]_  = \new_[63544]_  & \new_[63531]_ ;
  assign \new_[1472]_  = \new_[63518]_  & \new_[63505]_ ;
  assign \new_[1473]_  = \new_[63492]_  & \new_[63479]_ ;
  assign \new_[1474]_  = \new_[63466]_  & \new_[63453]_ ;
  assign \new_[1475]_  = \new_[63440]_  & \new_[63427]_ ;
  assign \new_[1476]_  = \new_[63414]_  & \new_[63401]_ ;
  assign \new_[1477]_  = \new_[63388]_  & \new_[63375]_ ;
  assign \new_[1478]_  = \new_[63362]_  & \new_[63349]_ ;
  assign \new_[1479]_  = \new_[63336]_  & \new_[63323]_ ;
  assign \new_[1480]_  = \new_[63310]_  & \new_[63297]_ ;
  assign \new_[1481]_  = \new_[63284]_  & \new_[63271]_ ;
  assign \new_[1482]_  = \new_[63258]_  & \new_[63245]_ ;
  assign \new_[1483]_  = \new_[63232]_  & \new_[63219]_ ;
  assign \new_[1484]_  = \new_[63206]_  & \new_[63193]_ ;
  assign \new_[1485]_  = \new_[63180]_  & \new_[63167]_ ;
  assign \new_[1486]_  = \new_[63154]_  & \new_[63141]_ ;
  assign \new_[1487]_  = \new_[63128]_  & \new_[63115]_ ;
  assign \new_[1488]_  = \new_[63102]_  & \new_[63089]_ ;
  assign \new_[1489]_  = \new_[63076]_  & \new_[63063]_ ;
  assign \new_[1490]_  = \new_[63050]_  & \new_[63037]_ ;
  assign \new_[1491]_  = \new_[63024]_  & \new_[63011]_ ;
  assign \new_[1492]_  = \new_[62998]_  & \new_[62985]_ ;
  assign \new_[1493]_  = \new_[62972]_  & \new_[62959]_ ;
  assign \new_[1494]_  = \new_[62946]_  & \new_[62933]_ ;
  assign \new_[1495]_  = \new_[62920]_  & \new_[62907]_ ;
  assign \new_[1496]_  = \new_[62894]_  & \new_[62881]_ ;
  assign \new_[1497]_  = \new_[62868]_  & \new_[62855]_ ;
  assign \new_[1498]_  = \new_[62842]_  & \new_[62829]_ ;
  assign \new_[1499]_  = \new_[62816]_  & \new_[62803]_ ;
  assign \new_[1500]_  = \new_[62790]_  & \new_[62777]_ ;
  assign \new_[1501]_  = \new_[62764]_  & \new_[62751]_ ;
  assign \new_[1502]_  = \new_[62738]_  & \new_[62725]_ ;
  assign \new_[1503]_  = \new_[62712]_  & \new_[62699]_ ;
  assign \new_[1504]_  = \new_[62686]_  & \new_[62673]_ ;
  assign \new_[1505]_  = \new_[62660]_  & \new_[62647]_ ;
  assign \new_[1506]_  = \new_[62634]_  & \new_[62621]_ ;
  assign \new_[1507]_  = \new_[62608]_  & \new_[62595]_ ;
  assign \new_[1508]_  = \new_[62582]_  & \new_[62569]_ ;
  assign \new_[1509]_  = \new_[62556]_  & \new_[62543]_ ;
  assign \new_[1510]_  = \new_[62530]_  & \new_[62517]_ ;
  assign \new_[1511]_  = \new_[62504]_  & \new_[62491]_ ;
  assign \new_[1512]_  = \new_[62478]_  & \new_[62465]_ ;
  assign \new_[1513]_  = \new_[62452]_  & \new_[62439]_ ;
  assign \new_[1514]_  = \new_[62426]_  & \new_[62413]_ ;
  assign \new_[1515]_  = \new_[62400]_  & \new_[62387]_ ;
  assign \new_[1516]_  = \new_[62374]_  & \new_[62361]_ ;
  assign \new_[1517]_  = \new_[62348]_  & \new_[62335]_ ;
  assign \new_[1518]_  = \new_[62322]_  & \new_[62309]_ ;
  assign \new_[1519]_  = \new_[62296]_  & \new_[62283]_ ;
  assign \new_[1520]_  = \new_[62270]_  & \new_[62257]_ ;
  assign \new_[1521]_  = \new_[62244]_  & \new_[62231]_ ;
  assign \new_[1522]_  = \new_[62218]_  & \new_[62205]_ ;
  assign \new_[1523]_  = \new_[62192]_  & \new_[62179]_ ;
  assign \new_[1524]_  = \new_[62166]_  & \new_[62153]_ ;
  assign \new_[1525]_  = \new_[62140]_  & \new_[62127]_ ;
  assign \new_[1526]_  = \new_[62114]_  & \new_[62101]_ ;
  assign \new_[1527]_  = \new_[62088]_  & \new_[62075]_ ;
  assign \new_[1528]_  = \new_[62062]_  & \new_[62049]_ ;
  assign \new_[1529]_  = \new_[62036]_  & \new_[62023]_ ;
  assign \new_[1530]_  = \new_[62010]_  & \new_[61997]_ ;
  assign \new_[1531]_  = \new_[61984]_  & \new_[61971]_ ;
  assign \new_[1532]_  = \new_[61958]_  & \new_[61945]_ ;
  assign \new_[1533]_  = \new_[61932]_  & \new_[61919]_ ;
  assign \new_[1534]_  = \new_[61906]_  & \new_[61893]_ ;
  assign \new_[1535]_  = \new_[61880]_  & \new_[61867]_ ;
  assign \new_[1536]_  = \new_[61854]_  & \new_[61841]_ ;
  assign \new_[1537]_  = \new_[61828]_  & \new_[61815]_ ;
  assign \new_[1538]_  = \new_[61802]_  & \new_[61789]_ ;
  assign \new_[1539]_  = \new_[61776]_  & \new_[61763]_ ;
  assign \new_[1540]_  = \new_[61750]_  & \new_[61737]_ ;
  assign \new_[1541]_  = \new_[61724]_  & \new_[61711]_ ;
  assign \new_[1542]_  = \new_[61698]_  & \new_[61685]_ ;
  assign \new_[1543]_  = \new_[61672]_  & \new_[61659]_ ;
  assign \new_[1544]_  = \new_[61646]_  & \new_[61633]_ ;
  assign \new_[1545]_  = \new_[61620]_  & \new_[61607]_ ;
  assign \new_[1546]_  = \new_[61594]_  & \new_[61581]_ ;
  assign \new_[1547]_  = \new_[61568]_  & \new_[61555]_ ;
  assign \new_[1548]_  = \new_[61542]_  & \new_[61529]_ ;
  assign \new_[1549]_  = \new_[61516]_  & \new_[61503]_ ;
  assign \new_[1550]_  = \new_[61490]_  & \new_[61477]_ ;
  assign \new_[1551]_  = \new_[61464]_  & \new_[61451]_ ;
  assign \new_[1552]_  = \new_[61438]_  & \new_[61425]_ ;
  assign \new_[1553]_  = \new_[61412]_  & \new_[61399]_ ;
  assign \new_[1554]_  = \new_[61386]_  & \new_[61373]_ ;
  assign \new_[1555]_  = \new_[61360]_  & \new_[61347]_ ;
  assign \new_[1556]_  = \new_[61334]_  & \new_[61321]_ ;
  assign \new_[1557]_  = \new_[61308]_  & \new_[61295]_ ;
  assign \new_[1558]_  = \new_[61282]_  & \new_[61269]_ ;
  assign \new_[1559]_  = \new_[61256]_  & \new_[61243]_ ;
  assign \new_[1560]_  = \new_[61230]_  & \new_[61217]_ ;
  assign \new_[1561]_  = \new_[61204]_  & \new_[61191]_ ;
  assign \new_[1562]_  = \new_[61178]_  & \new_[61165]_ ;
  assign \new_[1563]_  = \new_[61152]_  & \new_[61139]_ ;
  assign \new_[1564]_  = \new_[61126]_  & \new_[61113]_ ;
  assign \new_[1565]_  = \new_[61100]_  & \new_[61087]_ ;
  assign \new_[1566]_  = \new_[61074]_  & \new_[61061]_ ;
  assign \new_[1567]_  = \new_[61048]_  & \new_[61035]_ ;
  assign \new_[1568]_  = \new_[61022]_  & \new_[61009]_ ;
  assign \new_[1569]_  = \new_[60996]_  & \new_[60983]_ ;
  assign \new_[1570]_  = \new_[60970]_  & \new_[60957]_ ;
  assign \new_[1571]_  = \new_[60944]_  & \new_[60931]_ ;
  assign \new_[1572]_  = \new_[60918]_  & \new_[60905]_ ;
  assign \new_[1573]_  = \new_[60892]_  & \new_[60879]_ ;
  assign \new_[1574]_  = \new_[60866]_  & \new_[60853]_ ;
  assign \new_[1575]_  = \new_[60840]_  & \new_[60827]_ ;
  assign \new_[1576]_  = \new_[60814]_  & \new_[60801]_ ;
  assign \new_[1577]_  = \new_[60788]_  & \new_[60775]_ ;
  assign \new_[1578]_  = \new_[60762]_  & \new_[60749]_ ;
  assign \new_[1579]_  = \new_[60736]_  & \new_[60723]_ ;
  assign \new_[1580]_  = \new_[60710]_  & \new_[60697]_ ;
  assign \new_[1581]_  = \new_[60684]_  & \new_[60671]_ ;
  assign \new_[1582]_  = \new_[60658]_  & \new_[60645]_ ;
  assign \new_[1583]_  = \new_[60632]_  & \new_[60619]_ ;
  assign \new_[1584]_  = \new_[60606]_  & \new_[60593]_ ;
  assign \new_[1585]_  = \new_[60580]_  & \new_[60567]_ ;
  assign \new_[1586]_  = \new_[60554]_  & \new_[60541]_ ;
  assign \new_[1587]_  = \new_[60528]_  & \new_[60515]_ ;
  assign \new_[1588]_  = \new_[60502]_  & \new_[60489]_ ;
  assign \new_[1589]_  = \new_[60476]_  & \new_[60463]_ ;
  assign \new_[1590]_  = \new_[60450]_  & \new_[60437]_ ;
  assign \new_[1591]_  = \new_[60424]_  & \new_[60411]_ ;
  assign \new_[1592]_  = \new_[60398]_  & \new_[60385]_ ;
  assign \new_[1593]_  = \new_[60372]_  & \new_[60359]_ ;
  assign \new_[1594]_  = \new_[60346]_  & \new_[60333]_ ;
  assign \new_[1595]_  = \new_[60320]_  & \new_[60307]_ ;
  assign \new_[1596]_  = \new_[60294]_  & \new_[60281]_ ;
  assign \new_[1597]_  = \new_[60268]_  & \new_[60255]_ ;
  assign \new_[1598]_  = \new_[60242]_  & \new_[60229]_ ;
  assign \new_[1599]_  = \new_[60216]_  & \new_[60203]_ ;
  assign \new_[1600]_  = \new_[60190]_  & \new_[60177]_ ;
  assign \new_[1601]_  = \new_[60164]_  & \new_[60151]_ ;
  assign \new_[1602]_  = \new_[60138]_  & \new_[60125]_ ;
  assign \new_[1603]_  = \new_[60112]_  & \new_[60099]_ ;
  assign \new_[1604]_  = \new_[60088]_  & \new_[60075]_ ;
  assign \new_[1605]_  = \new_[60064]_  & \new_[60051]_ ;
  assign \new_[1606]_  = \new_[60040]_  & \new_[60027]_ ;
  assign \new_[1607]_  = \new_[60016]_  & \new_[60003]_ ;
  assign \new_[1608]_  = \new_[59992]_  & \new_[59979]_ ;
  assign \new_[1609]_  = \new_[59968]_  & \new_[59955]_ ;
  assign \new_[1610]_  = \new_[59944]_  & \new_[59931]_ ;
  assign \new_[1611]_  = \new_[59920]_  & \new_[59907]_ ;
  assign \new_[1612]_  = \new_[59896]_  & \new_[59883]_ ;
  assign \new_[1613]_  = \new_[59872]_  & \new_[59859]_ ;
  assign \new_[1614]_  = \new_[59848]_  & \new_[59835]_ ;
  assign \new_[1615]_  = \new_[59824]_  & \new_[59811]_ ;
  assign \new_[1616]_  = \new_[59800]_  & \new_[59787]_ ;
  assign \new_[1617]_  = \new_[59776]_  & \new_[59763]_ ;
  assign \new_[1618]_  = \new_[59752]_  & \new_[59739]_ ;
  assign \new_[1619]_  = \new_[59728]_  & \new_[59715]_ ;
  assign \new_[1620]_  = \new_[59704]_  & \new_[59691]_ ;
  assign \new_[1621]_  = \new_[59680]_  & \new_[59667]_ ;
  assign \new_[1622]_  = \new_[59656]_  & \new_[59643]_ ;
  assign \new_[1623]_  = \new_[59632]_  & \new_[59619]_ ;
  assign \new_[1624]_  = \new_[59608]_  & \new_[59595]_ ;
  assign \new_[1625]_  = \new_[59584]_  & \new_[59571]_ ;
  assign \new_[1626]_  = \new_[59560]_  & \new_[59547]_ ;
  assign \new_[1627]_  = \new_[59536]_  & \new_[59523]_ ;
  assign \new_[1628]_  = \new_[59512]_  & \new_[59499]_ ;
  assign \new_[1629]_  = \new_[59488]_  & \new_[59475]_ ;
  assign \new_[1630]_  = \new_[59464]_  & \new_[59451]_ ;
  assign \new_[1631]_  = \new_[59440]_  & \new_[59427]_ ;
  assign \new_[1632]_  = \new_[59416]_  & \new_[59403]_ ;
  assign \new_[1633]_  = \new_[59392]_  & \new_[59379]_ ;
  assign \new_[1634]_  = \new_[59368]_  & \new_[59355]_ ;
  assign \new_[1635]_  = \new_[59344]_  & \new_[59331]_ ;
  assign \new_[1636]_  = \new_[59320]_  & \new_[59307]_ ;
  assign \new_[1637]_  = \new_[59296]_  & \new_[59283]_ ;
  assign \new_[1638]_  = \new_[59272]_  & \new_[59259]_ ;
  assign \new_[1639]_  = \new_[59248]_  & \new_[59235]_ ;
  assign \new_[1640]_  = \new_[59224]_  & \new_[59211]_ ;
  assign \new_[1641]_  = \new_[59200]_  & \new_[59187]_ ;
  assign \new_[1642]_  = \new_[59176]_  & \new_[59163]_ ;
  assign \new_[1643]_  = \new_[59152]_  & \new_[59139]_ ;
  assign \new_[1644]_  = \new_[59128]_  & \new_[59115]_ ;
  assign \new_[1645]_  = \new_[59104]_  & \new_[59091]_ ;
  assign \new_[1646]_  = \new_[59080]_  & \new_[59067]_ ;
  assign \new_[1647]_  = \new_[59056]_  & \new_[59043]_ ;
  assign \new_[1648]_  = \new_[59032]_  & \new_[59019]_ ;
  assign \new_[1649]_  = \new_[59008]_  & \new_[58995]_ ;
  assign \new_[1650]_  = \new_[58984]_  & \new_[58971]_ ;
  assign \new_[1651]_  = \new_[58960]_  & \new_[58947]_ ;
  assign \new_[1652]_  = \new_[58936]_  & \new_[58923]_ ;
  assign \new_[1653]_  = \new_[58912]_  & \new_[58899]_ ;
  assign \new_[1654]_  = \new_[58888]_  & \new_[58875]_ ;
  assign \new_[1655]_  = \new_[58864]_  & \new_[58851]_ ;
  assign \new_[1656]_  = \new_[58840]_  & \new_[58827]_ ;
  assign \new_[1657]_  = \new_[58816]_  & \new_[58803]_ ;
  assign \new_[1658]_  = \new_[58792]_  & \new_[58779]_ ;
  assign \new_[1659]_  = \new_[58768]_  & \new_[58755]_ ;
  assign \new_[1660]_  = \new_[58744]_  & \new_[58731]_ ;
  assign \new_[1661]_  = \new_[58720]_  & \new_[58707]_ ;
  assign \new_[1662]_  = \new_[58696]_  & \new_[58683]_ ;
  assign \new_[1663]_  = \new_[58672]_  & \new_[58659]_ ;
  assign \new_[1664]_  = \new_[58648]_  & \new_[58635]_ ;
  assign \new_[1665]_  = \new_[58624]_  & \new_[58611]_ ;
  assign \new_[1666]_  = \new_[58600]_  & \new_[58587]_ ;
  assign \new_[1667]_  = \new_[58576]_  & \new_[58563]_ ;
  assign \new_[1668]_  = \new_[58552]_  & \new_[58539]_ ;
  assign \new_[1669]_  = \new_[58528]_  & \new_[58515]_ ;
  assign \new_[1670]_  = \new_[58504]_  & \new_[58491]_ ;
  assign \new_[1671]_  = \new_[58480]_  & \new_[58467]_ ;
  assign \new_[1672]_  = \new_[58456]_  & \new_[58443]_ ;
  assign \new_[1673]_  = \new_[58432]_  & \new_[58419]_ ;
  assign \new_[1674]_  = \new_[58408]_  & \new_[58395]_ ;
  assign \new_[1675]_  = \new_[58384]_  & \new_[58371]_ ;
  assign \new_[1676]_  = \new_[58360]_  & \new_[58347]_ ;
  assign \new_[1677]_  = \new_[58336]_  & \new_[58323]_ ;
  assign \new_[1678]_  = \new_[58312]_  & \new_[58299]_ ;
  assign \new_[1679]_  = \new_[58288]_  & \new_[58275]_ ;
  assign \new_[1680]_  = \new_[58264]_  & \new_[58251]_ ;
  assign \new_[1681]_  = \new_[58240]_  & \new_[58227]_ ;
  assign \new_[1682]_  = \new_[58216]_  & \new_[58203]_ ;
  assign \new_[1683]_  = \new_[58192]_  & \new_[58179]_ ;
  assign \new_[1684]_  = \new_[58168]_  & \new_[58155]_ ;
  assign \new_[1685]_  = \new_[58144]_  & \new_[58131]_ ;
  assign \new_[1686]_  = \new_[58120]_  & \new_[58107]_ ;
  assign \new_[1687]_  = \new_[58096]_  & \new_[58083]_ ;
  assign \new_[1688]_  = \new_[58072]_  & \new_[58059]_ ;
  assign \new_[1689]_  = \new_[58048]_  & \new_[58035]_ ;
  assign \new_[1690]_  = \new_[58024]_  & \new_[58011]_ ;
  assign \new_[1691]_  = \new_[58000]_  & \new_[57987]_ ;
  assign \new_[1692]_  = \new_[57976]_  & \new_[57963]_ ;
  assign \new_[1693]_  = \new_[57952]_  & \new_[57939]_ ;
  assign \new_[1694]_  = \new_[57928]_  & \new_[57915]_ ;
  assign \new_[1695]_  = \new_[57904]_  & \new_[57891]_ ;
  assign \new_[1696]_  = \new_[57880]_  & \new_[57867]_ ;
  assign \new_[1697]_  = \new_[57856]_  & \new_[57843]_ ;
  assign \new_[1698]_  = \new_[57832]_  & \new_[57819]_ ;
  assign \new_[1699]_  = \new_[57808]_  & \new_[57795]_ ;
  assign \new_[1700]_  = \new_[57784]_  & \new_[57771]_ ;
  assign \new_[1701]_  = \new_[57760]_  & \new_[57747]_ ;
  assign \new_[1702]_  = \new_[57736]_  & \new_[57723]_ ;
  assign \new_[1703]_  = \new_[57712]_  & \new_[57699]_ ;
  assign \new_[1704]_  = \new_[57688]_  & \new_[57675]_ ;
  assign \new_[1705]_  = \new_[57664]_  & \new_[57651]_ ;
  assign \new_[1706]_  = \new_[57640]_  & \new_[57627]_ ;
  assign \new_[1707]_  = \new_[57616]_  & \new_[57603]_ ;
  assign \new_[1708]_  = \new_[57592]_  & \new_[57579]_ ;
  assign \new_[1709]_  = \new_[57568]_  & \new_[57555]_ ;
  assign \new_[1710]_  = \new_[57544]_  & \new_[57531]_ ;
  assign \new_[1711]_  = \new_[57520]_  & \new_[57507]_ ;
  assign \new_[1712]_  = \new_[57496]_  & \new_[57483]_ ;
  assign \new_[1713]_  = \new_[57472]_  & \new_[57459]_ ;
  assign \new_[1714]_  = \new_[57448]_  & \new_[57435]_ ;
  assign \new_[1715]_  = \new_[57424]_  & \new_[57411]_ ;
  assign \new_[1716]_  = \new_[57400]_  & \new_[57387]_ ;
  assign \new_[1717]_  = \new_[57376]_  & \new_[57363]_ ;
  assign \new_[1718]_  = \new_[57352]_  & \new_[57339]_ ;
  assign \new_[1719]_  = \new_[57328]_  & \new_[57315]_ ;
  assign \new_[1720]_  = \new_[57304]_  & \new_[57291]_ ;
  assign \new_[1721]_  = \new_[57280]_  & \new_[57267]_ ;
  assign \new_[1722]_  = \new_[57256]_  & \new_[57243]_ ;
  assign \new_[1723]_  = \new_[57232]_  & \new_[57219]_ ;
  assign \new_[1724]_  = \new_[57208]_  & \new_[57195]_ ;
  assign \new_[1725]_  = \new_[57184]_  & \new_[57171]_ ;
  assign \new_[1726]_  = \new_[57160]_  & \new_[57147]_ ;
  assign \new_[1727]_  = \new_[57136]_  & \new_[57123]_ ;
  assign \new_[1728]_  = \new_[57112]_  & \new_[57099]_ ;
  assign \new_[1729]_  = \new_[57088]_  & \new_[57075]_ ;
  assign \new_[1730]_  = \new_[57064]_  & \new_[57051]_ ;
  assign \new_[1731]_  = \new_[57040]_  & \new_[57027]_ ;
  assign \new_[1732]_  = \new_[57016]_  & \new_[57003]_ ;
  assign \new_[1733]_  = \new_[56992]_  & \new_[56979]_ ;
  assign \new_[1734]_  = \new_[56968]_  & \new_[56955]_ ;
  assign \new_[1735]_  = \new_[56944]_  & \new_[56931]_ ;
  assign \new_[1736]_  = \new_[56920]_  & \new_[56907]_ ;
  assign \new_[1737]_  = \new_[56896]_  & \new_[56883]_ ;
  assign \new_[1738]_  = \new_[56872]_  & \new_[56859]_ ;
  assign \new_[1739]_  = \new_[56848]_  & \new_[56835]_ ;
  assign \new_[1740]_  = \new_[56824]_  & \new_[56811]_ ;
  assign \new_[1741]_  = \new_[56800]_  & \new_[56787]_ ;
  assign \new_[1742]_  = \new_[56776]_  & \new_[56763]_ ;
  assign \new_[1743]_  = \new_[56752]_  & \new_[56739]_ ;
  assign \new_[1744]_  = \new_[56728]_  & \new_[56715]_ ;
  assign \new_[1745]_  = \new_[56704]_  & \new_[56691]_ ;
  assign \new_[1746]_  = \new_[56680]_  & \new_[56667]_ ;
  assign \new_[1747]_  = \new_[56656]_  & \new_[56643]_ ;
  assign \new_[1748]_  = \new_[56632]_  & \new_[56619]_ ;
  assign \new_[1749]_  = \new_[56608]_  & \new_[56595]_ ;
  assign \new_[1750]_  = \new_[56584]_  & \new_[56571]_ ;
  assign \new_[1751]_  = \new_[56560]_  & \new_[56547]_ ;
  assign \new_[1752]_  = \new_[56536]_  & \new_[56523]_ ;
  assign \new_[1753]_  = \new_[56512]_  & \new_[56499]_ ;
  assign \new_[1754]_  = \new_[56488]_  & \new_[56475]_ ;
  assign \new_[1755]_  = \new_[56464]_  & \new_[56451]_ ;
  assign \new_[1756]_  = \new_[56440]_  & \new_[56427]_ ;
  assign \new_[1757]_  = \new_[56416]_  & \new_[56403]_ ;
  assign \new_[1758]_  = \new_[56392]_  & \new_[56379]_ ;
  assign \new_[1759]_  = \new_[56368]_  & \new_[56355]_ ;
  assign \new_[1760]_  = \new_[56344]_  & \new_[56331]_ ;
  assign \new_[1761]_  = \new_[56320]_  & \new_[56307]_ ;
  assign \new_[1762]_  = \new_[56296]_  & \new_[56283]_ ;
  assign \new_[1763]_  = \new_[56272]_  & \new_[56259]_ ;
  assign \new_[1764]_  = \new_[56248]_  & \new_[56235]_ ;
  assign \new_[1765]_  = \new_[56224]_  & \new_[56211]_ ;
  assign \new_[1766]_  = \new_[56200]_  & \new_[56187]_ ;
  assign \new_[1767]_  = \new_[56176]_  & \new_[56163]_ ;
  assign \new_[1768]_  = \new_[56152]_  & \new_[56139]_ ;
  assign \new_[1769]_  = \new_[56128]_  & \new_[56115]_ ;
  assign \new_[1770]_  = \new_[56104]_  & \new_[56091]_ ;
  assign \new_[1771]_  = \new_[56080]_  & \new_[56067]_ ;
  assign \new_[1772]_  = \new_[56056]_  & \new_[56043]_ ;
  assign \new_[1773]_  = \new_[56032]_  & \new_[56019]_ ;
  assign \new_[1774]_  = \new_[56008]_  & \new_[55995]_ ;
  assign \new_[1775]_  = \new_[55984]_  & \new_[55971]_ ;
  assign \new_[1776]_  = \new_[55960]_  & \new_[55947]_ ;
  assign \new_[1777]_  = \new_[55936]_  & \new_[55923]_ ;
  assign \new_[1778]_  = \new_[55912]_  & \new_[55899]_ ;
  assign \new_[1779]_  = \new_[55888]_  & \new_[55875]_ ;
  assign \new_[1780]_  = \new_[55864]_  & \new_[55851]_ ;
  assign \new_[1781]_  = \new_[55840]_  & \new_[55827]_ ;
  assign \new_[1782]_  = \new_[55816]_  & \new_[55803]_ ;
  assign \new_[1783]_  = \new_[55792]_  & \new_[55779]_ ;
  assign \new_[1784]_  = \new_[55768]_  & \new_[55755]_ ;
  assign \new_[1785]_  = \new_[55744]_  & \new_[55731]_ ;
  assign \new_[1786]_  = \new_[55720]_  & \new_[55707]_ ;
  assign \new_[1787]_  = \new_[55696]_  & \new_[55683]_ ;
  assign \new_[1788]_  = \new_[55672]_  & \new_[55659]_ ;
  assign \new_[1789]_  = \new_[55648]_  & \new_[55635]_ ;
  assign \new_[1790]_  = \new_[55624]_  & \new_[55611]_ ;
  assign \new_[1791]_  = \new_[55600]_  & \new_[55587]_ ;
  assign \new_[1792]_  = \new_[55576]_  & \new_[55563]_ ;
  assign \new_[1793]_  = \new_[55552]_  & \new_[55539]_ ;
  assign \new_[1794]_  = \new_[55528]_  & \new_[55515]_ ;
  assign \new_[1795]_  = \new_[55504]_  & \new_[55491]_ ;
  assign \new_[1796]_  = \new_[55480]_  & \new_[55467]_ ;
  assign \new_[1797]_  = \new_[55456]_  & \new_[55443]_ ;
  assign \new_[1798]_  = \new_[55432]_  & \new_[55419]_ ;
  assign \new_[1799]_  = \new_[55408]_  & \new_[55395]_ ;
  assign \new_[1800]_  = \new_[55384]_  & \new_[55371]_ ;
  assign \new_[1801]_  = \new_[55360]_  & \new_[55347]_ ;
  assign \new_[1802]_  = \new_[55336]_  & \new_[55323]_ ;
  assign \new_[1803]_  = \new_[55312]_  & \new_[55299]_ ;
  assign \new_[1804]_  = \new_[55288]_  & \new_[55275]_ ;
  assign \new_[1805]_  = \new_[55264]_  & \new_[55251]_ ;
  assign \new_[1806]_  = \new_[55240]_  & \new_[55227]_ ;
  assign \new_[1807]_  = \new_[55216]_  & \new_[55203]_ ;
  assign \new_[1808]_  = \new_[55192]_  & \new_[55179]_ ;
  assign \new_[1809]_  = \new_[55168]_  & \new_[55155]_ ;
  assign \new_[1810]_  = \new_[55144]_  & \new_[55131]_ ;
  assign \new_[1811]_  = \new_[55120]_  & \new_[55107]_ ;
  assign \new_[1812]_  = \new_[55096]_  & \new_[55083]_ ;
  assign \new_[1813]_  = \new_[55072]_  & \new_[55059]_ ;
  assign \new_[1814]_  = \new_[55048]_  & \new_[55035]_ ;
  assign \new_[1815]_  = \new_[55024]_  & \new_[55011]_ ;
  assign \new_[1816]_  = \new_[55000]_  & \new_[54987]_ ;
  assign \new_[1817]_  = \new_[54976]_  & \new_[54963]_ ;
  assign \new_[1818]_  = \new_[54952]_  & \new_[54939]_ ;
  assign \new_[1819]_  = \new_[54928]_  & \new_[54915]_ ;
  assign \new_[1820]_  = \new_[54904]_  & \new_[54891]_ ;
  assign \new_[1821]_  = \new_[54880]_  & \new_[54867]_ ;
  assign \new_[1822]_  = \new_[54856]_  & \new_[54843]_ ;
  assign \new_[1823]_  = \new_[54832]_  & \new_[54819]_ ;
  assign \new_[1824]_  = \new_[54808]_  & \new_[54795]_ ;
  assign \new_[1825]_  = \new_[54784]_  & \new_[54771]_ ;
  assign \new_[1826]_  = \new_[54760]_  & \new_[54747]_ ;
  assign \new_[1827]_  = \new_[54736]_  & \new_[54723]_ ;
  assign \new_[1828]_  = \new_[54712]_  & \new_[54699]_ ;
  assign \new_[1829]_  = \new_[54688]_  & \new_[54675]_ ;
  assign \new_[1830]_  = \new_[54664]_  & \new_[54651]_ ;
  assign \new_[1831]_  = \new_[54640]_  & \new_[54627]_ ;
  assign \new_[1832]_  = \new_[54616]_  & \new_[54603]_ ;
  assign \new_[1833]_  = \new_[54592]_  & \new_[54579]_ ;
  assign \new_[1834]_  = \new_[54568]_  & \new_[54555]_ ;
  assign \new_[1835]_  = \new_[54544]_  & \new_[54531]_ ;
  assign \new_[1836]_  = \new_[54520]_  & \new_[54507]_ ;
  assign \new_[1837]_  = \new_[54496]_  & \new_[54483]_ ;
  assign \new_[1838]_  = \new_[54472]_  & \new_[54459]_ ;
  assign \new_[1839]_  = \new_[54448]_  & \new_[54435]_ ;
  assign \new_[1840]_  = \new_[54424]_  & \new_[54411]_ ;
  assign \new_[1841]_  = \new_[54400]_  & \new_[54387]_ ;
  assign \new_[1842]_  = \new_[54376]_  & \new_[54363]_ ;
  assign \new_[1843]_  = \new_[54352]_  & \new_[54339]_ ;
  assign \new_[1844]_  = \new_[54328]_  & \new_[54315]_ ;
  assign \new_[1845]_  = \new_[54304]_  & \new_[54291]_ ;
  assign \new_[1846]_  = \new_[54280]_  & \new_[54267]_ ;
  assign \new_[1847]_  = \new_[54256]_  & \new_[54243]_ ;
  assign \new_[1848]_  = \new_[54232]_  & \new_[54219]_ ;
  assign \new_[1849]_  = \new_[54208]_  & \new_[54195]_ ;
  assign \new_[1850]_  = \new_[54184]_  & \new_[54171]_ ;
  assign \new_[1851]_  = \new_[54160]_  & \new_[54147]_ ;
  assign \new_[1852]_  = \new_[54136]_  & \new_[54123]_ ;
  assign \new_[1853]_  = \new_[54112]_  & \new_[54099]_ ;
  assign \new_[1854]_  = \new_[54088]_  & \new_[54075]_ ;
  assign \new_[1855]_  = \new_[54064]_  & \new_[54051]_ ;
  assign \new_[1856]_  = \new_[54040]_  & \new_[54027]_ ;
  assign \new_[1857]_  = \new_[54016]_  & \new_[54003]_ ;
  assign \new_[1858]_  = \new_[53992]_  & \new_[53979]_ ;
  assign \new_[1859]_  = \new_[53968]_  & \new_[53955]_ ;
  assign \new_[1860]_  = \new_[53944]_  & \new_[53931]_ ;
  assign \new_[1861]_  = \new_[53920]_  & \new_[53907]_ ;
  assign \new_[1862]_  = \new_[53896]_  & \new_[53883]_ ;
  assign \new_[1863]_  = \new_[53872]_  & \new_[53859]_ ;
  assign \new_[1864]_  = \new_[53848]_  & \new_[53835]_ ;
  assign \new_[1865]_  = \new_[53824]_  & \new_[53811]_ ;
  assign \new_[1866]_  = \new_[53800]_  & \new_[53787]_ ;
  assign \new_[1867]_  = \new_[53776]_  & \new_[53763]_ ;
  assign \new_[1868]_  = \new_[53752]_  & \new_[53739]_ ;
  assign \new_[1869]_  = \new_[53728]_  & \new_[53715]_ ;
  assign \new_[1870]_  = \new_[53704]_  & \new_[53691]_ ;
  assign \new_[1871]_  = \new_[53680]_  & \new_[53667]_ ;
  assign \new_[1872]_  = \new_[53656]_  & \new_[53643]_ ;
  assign \new_[1873]_  = \new_[53632]_  & \new_[53619]_ ;
  assign \new_[1874]_  = \new_[53608]_  & \new_[53595]_ ;
  assign \new_[1875]_  = \new_[53584]_  & \new_[53571]_ ;
  assign \new_[1876]_  = \new_[53560]_  & \new_[53547]_ ;
  assign \new_[1877]_  = \new_[53536]_  & \new_[53523]_ ;
  assign \new_[1878]_  = \new_[53512]_  & \new_[53499]_ ;
  assign \new_[1879]_  = \new_[53488]_  & \new_[53475]_ ;
  assign \new_[1880]_  = \new_[53464]_  & \new_[53451]_ ;
  assign \new_[1881]_  = \new_[53440]_  & \new_[53427]_ ;
  assign \new_[1882]_  = \new_[53416]_  & \new_[53403]_ ;
  assign \new_[1883]_  = \new_[53392]_  & \new_[53379]_ ;
  assign \new_[1884]_  = \new_[53368]_  & \new_[53355]_ ;
  assign \new_[1885]_  = \new_[53344]_  & \new_[53331]_ ;
  assign \new_[1886]_  = \new_[53320]_  & \new_[53307]_ ;
  assign \new_[1887]_  = \new_[53296]_  & \new_[53283]_ ;
  assign \new_[1888]_  = \new_[53272]_  & \new_[53259]_ ;
  assign \new_[1889]_  = \new_[53248]_  & \new_[53235]_ ;
  assign \new_[1890]_  = \new_[53224]_  & \new_[53211]_ ;
  assign \new_[1891]_  = \new_[53200]_  & \new_[53187]_ ;
  assign \new_[1892]_  = \new_[53176]_  & \new_[53163]_ ;
  assign \new_[1893]_  = \new_[53152]_  & \new_[53139]_ ;
  assign \new_[1894]_  = \new_[53128]_  & \new_[53115]_ ;
  assign \new_[1895]_  = \new_[53104]_  & \new_[53091]_ ;
  assign \new_[1896]_  = \new_[53080]_  & \new_[53067]_ ;
  assign \new_[1897]_  = \new_[53056]_  & \new_[53043]_ ;
  assign \new_[1898]_  = \new_[53032]_  & \new_[53019]_ ;
  assign \new_[1899]_  = \new_[53008]_  & \new_[52995]_ ;
  assign \new_[1900]_  = \new_[52984]_  & \new_[52971]_ ;
  assign \new_[1901]_  = \new_[52960]_  & \new_[52947]_ ;
  assign \new_[1902]_  = \new_[52936]_  & \new_[52923]_ ;
  assign \new_[1903]_  = \new_[52912]_  & \new_[52899]_ ;
  assign \new_[1904]_  = \new_[52888]_  & \new_[52875]_ ;
  assign \new_[1905]_  = \new_[52864]_  & \new_[52851]_ ;
  assign \new_[1906]_  = \new_[52840]_  & \new_[52827]_ ;
  assign \new_[1907]_  = \new_[52816]_  & \new_[52803]_ ;
  assign \new_[1908]_  = \new_[52792]_  & \new_[52779]_ ;
  assign \new_[1909]_  = \new_[52768]_  & \new_[52755]_ ;
  assign \new_[1910]_  = \new_[52744]_  & \new_[52731]_ ;
  assign \new_[1911]_  = \new_[52720]_  & \new_[52707]_ ;
  assign \new_[1912]_  = \new_[52696]_  & \new_[52683]_ ;
  assign \new_[1913]_  = \new_[52672]_  & \new_[52659]_ ;
  assign \new_[1914]_  = \new_[52648]_  & \new_[52635]_ ;
  assign \new_[1915]_  = \new_[52624]_  & \new_[52611]_ ;
  assign \new_[1916]_  = \new_[52600]_  & \new_[52587]_ ;
  assign \new_[1917]_  = \new_[52576]_  & \new_[52563]_ ;
  assign \new_[1918]_  = \new_[52552]_  & \new_[52539]_ ;
  assign \new_[1919]_  = \new_[52528]_  & \new_[52515]_ ;
  assign \new_[1920]_  = \new_[52504]_  & \new_[52491]_ ;
  assign \new_[1921]_  = \new_[52480]_  & \new_[52467]_ ;
  assign \new_[1922]_  = \new_[52456]_  & \new_[52443]_ ;
  assign \new_[1923]_  = \new_[52432]_  & \new_[52419]_ ;
  assign \new_[1924]_  = \new_[52408]_  & \new_[52395]_ ;
  assign \new_[1925]_  = \new_[52384]_  & \new_[52371]_ ;
  assign \new_[1926]_  = \new_[52360]_  & \new_[52347]_ ;
  assign \new_[1927]_  = \new_[52336]_  & \new_[52323]_ ;
  assign \new_[1928]_  = \new_[52312]_  & \new_[52299]_ ;
  assign \new_[1929]_  = \new_[52288]_  & \new_[52275]_ ;
  assign \new_[1930]_  = \new_[52264]_  & \new_[52251]_ ;
  assign \new_[1931]_  = \new_[52240]_  & \new_[52227]_ ;
  assign \new_[1932]_  = \new_[52216]_  & \new_[52203]_ ;
  assign \new_[1933]_  = \new_[52192]_  & \new_[52179]_ ;
  assign \new_[1934]_  = \new_[52168]_  & \new_[52155]_ ;
  assign \new_[1935]_  = \new_[52144]_  & \new_[52131]_ ;
  assign \new_[1936]_  = \new_[52120]_  & \new_[52107]_ ;
  assign \new_[1937]_  = \new_[52096]_  & \new_[52083]_ ;
  assign \new_[1938]_  = \new_[52072]_  & \new_[52059]_ ;
  assign \new_[1939]_  = \new_[52048]_  & \new_[52035]_ ;
  assign \new_[1940]_  = \new_[52024]_  & \new_[52011]_ ;
  assign \new_[1941]_  = \new_[52000]_  & \new_[51987]_ ;
  assign \new_[1942]_  = \new_[51976]_  & \new_[51963]_ ;
  assign \new_[1943]_  = \new_[51952]_  & \new_[51939]_ ;
  assign \new_[1944]_  = \new_[51928]_  & \new_[51915]_ ;
  assign \new_[1945]_  = \new_[51904]_  & \new_[51891]_ ;
  assign \new_[1946]_  = \new_[51880]_  & \new_[51867]_ ;
  assign \new_[1947]_  = \new_[51856]_  & \new_[51843]_ ;
  assign \new_[1948]_  = \new_[51832]_  & \new_[51819]_ ;
  assign \new_[1949]_  = \new_[51808]_  & \new_[51795]_ ;
  assign \new_[1950]_  = \new_[51784]_  & \new_[51771]_ ;
  assign \new_[1951]_  = \new_[51760]_  & \new_[51747]_ ;
  assign \new_[1952]_  = \new_[51736]_  & \new_[51723]_ ;
  assign \new_[1953]_  = \new_[51712]_  & \new_[51699]_ ;
  assign \new_[1954]_  = \new_[51688]_  & \new_[51675]_ ;
  assign \new_[1955]_  = \new_[51664]_  & \new_[51651]_ ;
  assign \new_[1956]_  = \new_[51640]_  & \new_[51627]_ ;
  assign \new_[1957]_  = \new_[51616]_  & \new_[51603]_ ;
  assign \new_[1958]_  = \new_[51592]_  & \new_[51579]_ ;
  assign \new_[1959]_  = \new_[51568]_  & \new_[51555]_ ;
  assign \new_[1960]_  = \new_[51544]_  & \new_[51531]_ ;
  assign \new_[1961]_  = \new_[51520]_  & \new_[51507]_ ;
  assign \new_[1962]_  = \new_[51496]_  & \new_[51483]_ ;
  assign \new_[1963]_  = \new_[51472]_  & \new_[51459]_ ;
  assign \new_[1964]_  = \new_[51448]_  & \new_[51435]_ ;
  assign \new_[1965]_  = \new_[51424]_  & \new_[51411]_ ;
  assign \new_[1966]_  = \new_[51400]_  & \new_[51387]_ ;
  assign \new_[1967]_  = \new_[51376]_  & \new_[51363]_ ;
  assign \new_[1968]_  = \new_[51352]_  & \new_[51339]_ ;
  assign \new_[1969]_  = \new_[51328]_  & \new_[51315]_ ;
  assign \new_[1970]_  = \new_[51304]_  & \new_[51291]_ ;
  assign \new_[1971]_  = \new_[51280]_  & \new_[51267]_ ;
  assign \new_[1972]_  = \new_[51256]_  & \new_[51243]_ ;
  assign \new_[1973]_  = \new_[51232]_  & \new_[51219]_ ;
  assign \new_[1974]_  = \new_[51208]_  & \new_[51195]_ ;
  assign \new_[1975]_  = \new_[51184]_  & \new_[51171]_ ;
  assign \new_[1976]_  = \new_[51160]_  & \new_[51147]_ ;
  assign \new_[1977]_  = \new_[51136]_  & \new_[51123]_ ;
  assign \new_[1978]_  = \new_[51112]_  & \new_[51099]_ ;
  assign \new_[1979]_  = \new_[51088]_  & \new_[51075]_ ;
  assign \new_[1980]_  = \new_[51064]_  & \new_[51051]_ ;
  assign \new_[1981]_  = \new_[51040]_  & \new_[51027]_ ;
  assign \new_[1982]_  = \new_[51016]_  & \new_[51003]_ ;
  assign \new_[1983]_  = \new_[50992]_  & \new_[50979]_ ;
  assign \new_[1984]_  = \new_[50968]_  & \new_[50955]_ ;
  assign \new_[1985]_  = \new_[50944]_  & \new_[50931]_ ;
  assign \new_[1986]_  = \new_[50920]_  & \new_[50907]_ ;
  assign \new_[1987]_  = \new_[50896]_  & \new_[50883]_ ;
  assign \new_[1988]_  = \new_[50872]_  & \new_[50859]_ ;
  assign \new_[1989]_  = \new_[50848]_  & \new_[50835]_ ;
  assign \new_[1990]_  = \new_[50824]_  & \new_[50811]_ ;
  assign \new_[1991]_  = \new_[50800]_  & \new_[50787]_ ;
  assign \new_[1992]_  = \new_[50776]_  & \new_[50763]_ ;
  assign \new_[1993]_  = \new_[50752]_  & \new_[50739]_ ;
  assign \new_[1994]_  = \new_[50728]_  & \new_[50715]_ ;
  assign \new_[1995]_  = \new_[50704]_  & \new_[50691]_ ;
  assign \new_[1996]_  = \new_[50680]_  & \new_[50667]_ ;
  assign \new_[1997]_  = \new_[50656]_  & \new_[50643]_ ;
  assign \new_[1998]_  = \new_[50632]_  & \new_[50619]_ ;
  assign \new_[1999]_  = \new_[50608]_  & \new_[50595]_ ;
  assign \new_[2000]_  = \new_[50584]_  & \new_[50571]_ ;
  assign \new_[2001]_  = \new_[50560]_  & \new_[50547]_ ;
  assign \new_[2002]_  = \new_[50536]_  & \new_[50523]_ ;
  assign \new_[2003]_  = \new_[50512]_  & \new_[50499]_ ;
  assign \new_[2004]_  = \new_[50488]_  & \new_[50475]_ ;
  assign \new_[2005]_  = \new_[50464]_  & \new_[50451]_ ;
  assign \new_[2006]_  = \new_[50440]_  & \new_[50427]_ ;
  assign \new_[2007]_  = \new_[50416]_  & \new_[50403]_ ;
  assign \new_[2008]_  = \new_[50392]_  & \new_[50379]_ ;
  assign \new_[2009]_  = \new_[50368]_  & \new_[50355]_ ;
  assign \new_[2010]_  = \new_[50344]_  & \new_[50331]_ ;
  assign \new_[2011]_  = \new_[50320]_  & \new_[50307]_ ;
  assign \new_[2012]_  = \new_[50296]_  & \new_[50283]_ ;
  assign \new_[2013]_  = \new_[50272]_  & \new_[50259]_ ;
  assign \new_[2014]_  = \new_[50248]_  & \new_[50235]_ ;
  assign \new_[2015]_  = \new_[50224]_  & \new_[50211]_ ;
  assign \new_[2016]_  = \new_[50200]_  & \new_[50187]_ ;
  assign \new_[2017]_  = \new_[50176]_  & \new_[50163]_ ;
  assign \new_[2018]_  = \new_[50152]_  & \new_[50139]_ ;
  assign \new_[2019]_  = \new_[50128]_  & \new_[50115]_ ;
  assign \new_[2020]_  = \new_[50104]_  & \new_[50091]_ ;
  assign \new_[2021]_  = \new_[50080]_  & \new_[50067]_ ;
  assign \new_[2022]_  = \new_[50056]_  & \new_[50043]_ ;
  assign \new_[2023]_  = \new_[50032]_  & \new_[50019]_ ;
  assign \new_[2024]_  = \new_[50008]_  & \new_[49995]_ ;
  assign \new_[2025]_  = \new_[49984]_  & \new_[49971]_ ;
  assign \new_[2026]_  = \new_[49960]_  & \new_[49947]_ ;
  assign \new_[2027]_  = \new_[49936]_  & \new_[49923]_ ;
  assign \new_[2028]_  = \new_[49912]_  & \new_[49899]_ ;
  assign \new_[2029]_  = \new_[49888]_  & \new_[49875]_ ;
  assign \new_[2030]_  = \new_[49864]_  & \new_[49851]_ ;
  assign \new_[2031]_  = \new_[49840]_  & \new_[49827]_ ;
  assign \new_[2032]_  = \new_[49816]_  & \new_[49803]_ ;
  assign \new_[2033]_  = \new_[49792]_  & \new_[49779]_ ;
  assign \new_[2034]_  = \new_[49768]_  & \new_[49755]_ ;
  assign \new_[2035]_  = \new_[49744]_  & \new_[49731]_ ;
  assign \new_[2036]_  = \new_[49720]_  & \new_[49707]_ ;
  assign \new_[2037]_  = \new_[49696]_  & \new_[49683]_ ;
  assign \new_[2038]_  = \new_[49672]_  & \new_[49659]_ ;
  assign \new_[2039]_  = \new_[49648]_  & \new_[49635]_ ;
  assign \new_[2040]_  = \new_[49624]_  & \new_[49611]_ ;
  assign \new_[2041]_  = \new_[49600]_  & \new_[49587]_ ;
  assign \new_[2042]_  = \new_[49576]_  & \new_[49563]_ ;
  assign \new_[2043]_  = \new_[49552]_  & \new_[49539]_ ;
  assign \new_[2044]_  = \new_[49528]_  & \new_[49515]_ ;
  assign \new_[2045]_  = \new_[49504]_  & \new_[49491]_ ;
  assign \new_[2046]_  = \new_[49480]_  & \new_[49467]_ ;
  assign \new_[2047]_  = \new_[49456]_  & \new_[49443]_ ;
  assign \new_[2048]_  = \new_[49432]_  & \new_[49419]_ ;
  assign \new_[2049]_  = \new_[49408]_  & \new_[49395]_ ;
  assign \new_[2050]_  = \new_[49384]_  & \new_[49371]_ ;
  assign \new_[2051]_  = \new_[49360]_  & \new_[49347]_ ;
  assign \new_[2052]_  = \new_[49336]_  & \new_[49323]_ ;
  assign \new_[2053]_  = \new_[49312]_  & \new_[49299]_ ;
  assign \new_[2054]_  = \new_[49288]_  & \new_[49275]_ ;
  assign \new_[2055]_  = \new_[49264]_  & \new_[49251]_ ;
  assign \new_[2056]_  = \new_[49240]_  & \new_[49227]_ ;
  assign \new_[2057]_  = \new_[49216]_  & \new_[49203]_ ;
  assign \new_[2058]_  = \new_[49192]_  & \new_[49179]_ ;
  assign \new_[2059]_  = \new_[49168]_  & \new_[49155]_ ;
  assign \new_[2060]_  = \new_[49144]_  & \new_[49131]_ ;
  assign \new_[2061]_  = \new_[49120]_  & \new_[49107]_ ;
  assign \new_[2062]_  = \new_[49096]_  & \new_[49083]_ ;
  assign \new_[2063]_  = \new_[49072]_  & \new_[49059]_ ;
  assign \new_[2064]_  = \new_[49048]_  & \new_[49035]_ ;
  assign \new_[2065]_  = \new_[49024]_  & \new_[49011]_ ;
  assign \new_[2066]_  = \new_[49000]_  & \new_[48987]_ ;
  assign \new_[2067]_  = \new_[48976]_  & \new_[48963]_ ;
  assign \new_[2068]_  = \new_[48952]_  & \new_[48939]_ ;
  assign \new_[2069]_  = \new_[48928]_  & \new_[48915]_ ;
  assign \new_[2070]_  = \new_[48904]_  & \new_[48891]_ ;
  assign \new_[2071]_  = \new_[48880]_  & \new_[48867]_ ;
  assign \new_[2072]_  = \new_[48856]_  & \new_[48843]_ ;
  assign \new_[2073]_  = \new_[48832]_  & \new_[48819]_ ;
  assign \new_[2074]_  = \new_[48808]_  & \new_[48795]_ ;
  assign \new_[2075]_  = \new_[48784]_  & \new_[48771]_ ;
  assign \new_[2076]_  = \new_[48760]_  & \new_[48747]_ ;
  assign \new_[2077]_  = \new_[48736]_  & \new_[48723]_ ;
  assign \new_[2078]_  = \new_[48712]_  & \new_[48699]_ ;
  assign \new_[2079]_  = \new_[48688]_  & \new_[48675]_ ;
  assign \new_[2080]_  = \new_[48664]_  & \new_[48651]_ ;
  assign \new_[2081]_  = \new_[48640]_  & \new_[48627]_ ;
  assign \new_[2082]_  = \new_[48616]_  & \new_[48603]_ ;
  assign \new_[2083]_  = \new_[48592]_  & \new_[48579]_ ;
  assign \new_[2084]_  = \new_[48568]_  & \new_[48555]_ ;
  assign \new_[2085]_  = \new_[48544]_  & \new_[48531]_ ;
  assign \new_[2086]_  = \new_[48520]_  & \new_[48507]_ ;
  assign \new_[2087]_  = \new_[48496]_  & \new_[48483]_ ;
  assign \new_[2088]_  = \new_[48472]_  & \new_[48459]_ ;
  assign \new_[2089]_  = \new_[48448]_  & \new_[48435]_ ;
  assign \new_[2090]_  = \new_[48424]_  & \new_[48411]_ ;
  assign \new_[2091]_  = \new_[48400]_  & \new_[48387]_ ;
  assign \new_[2092]_  = \new_[48376]_  & \new_[48363]_ ;
  assign \new_[2093]_  = \new_[48352]_  & \new_[48339]_ ;
  assign \new_[2094]_  = \new_[48328]_  & \new_[48315]_ ;
  assign \new_[2095]_  = \new_[48304]_  & \new_[48291]_ ;
  assign \new_[2096]_  = \new_[48280]_  & \new_[48267]_ ;
  assign \new_[2097]_  = \new_[48256]_  & \new_[48243]_ ;
  assign \new_[2098]_  = \new_[48232]_  & \new_[48219]_ ;
  assign \new_[2099]_  = \new_[48208]_  & \new_[48195]_ ;
  assign \new_[2100]_  = \new_[48184]_  & \new_[48171]_ ;
  assign \new_[2101]_  = \new_[48160]_  & \new_[48147]_ ;
  assign \new_[2102]_  = \new_[48136]_  & \new_[48123]_ ;
  assign \new_[2103]_  = \new_[48112]_  & \new_[48099]_ ;
  assign \new_[2104]_  = \new_[48088]_  & \new_[48075]_ ;
  assign \new_[2105]_  = \new_[48064]_  & \new_[48051]_ ;
  assign \new_[2106]_  = \new_[48040]_  & \new_[48027]_ ;
  assign \new_[2107]_  = \new_[48016]_  & \new_[48003]_ ;
  assign \new_[2108]_  = \new_[47992]_  & \new_[47979]_ ;
  assign \new_[2109]_  = \new_[47968]_  & \new_[47955]_ ;
  assign \new_[2110]_  = \new_[47944]_  & \new_[47931]_ ;
  assign \new_[2111]_  = \new_[47920]_  & \new_[47907]_ ;
  assign \new_[2112]_  = \new_[47896]_  & \new_[47883]_ ;
  assign \new_[2113]_  = \new_[47872]_  & \new_[47859]_ ;
  assign \new_[2114]_  = \new_[47848]_  & \new_[47835]_ ;
  assign \new_[2115]_  = \new_[47824]_  & \new_[47811]_ ;
  assign \new_[2116]_  = \new_[47800]_  & \new_[47787]_ ;
  assign \new_[2117]_  = \new_[47776]_  & \new_[47763]_ ;
  assign \new_[2118]_  = \new_[47752]_  & \new_[47739]_ ;
  assign \new_[2119]_  = \new_[47728]_  & \new_[47715]_ ;
  assign \new_[2120]_  = \new_[47704]_  & \new_[47691]_ ;
  assign \new_[2121]_  = \new_[47680]_  & \new_[47667]_ ;
  assign \new_[2122]_  = \new_[47656]_  & \new_[47643]_ ;
  assign \new_[2123]_  = \new_[47632]_  & \new_[47619]_ ;
  assign \new_[2124]_  = \new_[47608]_  & \new_[47595]_ ;
  assign \new_[2125]_  = \new_[47584]_  & \new_[47571]_ ;
  assign \new_[2126]_  = \new_[47560]_  & \new_[47547]_ ;
  assign \new_[2127]_  = \new_[47536]_  & \new_[47523]_ ;
  assign \new_[2128]_  = \new_[47512]_  & \new_[47499]_ ;
  assign \new_[2129]_  = \new_[47488]_  & \new_[47475]_ ;
  assign \new_[2130]_  = \new_[47464]_  & \new_[47451]_ ;
  assign \new_[2131]_  = \new_[47440]_  & \new_[47427]_ ;
  assign \new_[2132]_  = \new_[47416]_  & \new_[47403]_ ;
  assign \new_[2133]_  = \new_[47392]_  & \new_[47379]_ ;
  assign \new_[2134]_  = \new_[47368]_  & \new_[47355]_ ;
  assign \new_[2135]_  = \new_[47344]_  & \new_[47331]_ ;
  assign \new_[2136]_  = \new_[47320]_  & \new_[47307]_ ;
  assign \new_[2137]_  = \new_[47296]_  & \new_[47283]_ ;
  assign \new_[2138]_  = \new_[47272]_  & \new_[47259]_ ;
  assign \new_[2139]_  = \new_[47248]_  & \new_[47235]_ ;
  assign \new_[2140]_  = \new_[47224]_  & \new_[47211]_ ;
  assign \new_[2141]_  = \new_[47200]_  & \new_[47187]_ ;
  assign \new_[2142]_  = \new_[47176]_  & \new_[47163]_ ;
  assign \new_[2143]_  = \new_[47152]_  & \new_[47139]_ ;
  assign \new_[2144]_  = \new_[47128]_  & \new_[47115]_ ;
  assign \new_[2145]_  = \new_[47104]_  & \new_[47091]_ ;
  assign \new_[2146]_  = \new_[47080]_  & \new_[47067]_ ;
  assign \new_[2147]_  = \new_[47056]_  & \new_[47043]_ ;
  assign \new_[2148]_  = \new_[47032]_  & \new_[47019]_ ;
  assign \new_[2149]_  = \new_[47008]_  & \new_[46995]_ ;
  assign \new_[2150]_  = \new_[46984]_  & \new_[46971]_ ;
  assign \new_[2151]_  = \new_[46960]_  & \new_[46947]_ ;
  assign \new_[2152]_  = \new_[46936]_  & \new_[46923]_ ;
  assign \new_[2153]_  = \new_[46912]_  & \new_[46899]_ ;
  assign \new_[2154]_  = \new_[46888]_  & \new_[46875]_ ;
  assign \new_[2155]_  = \new_[46864]_  & \new_[46851]_ ;
  assign \new_[2156]_  = \new_[46840]_  & \new_[46827]_ ;
  assign \new_[2157]_  = \new_[46816]_  & \new_[46803]_ ;
  assign \new_[2158]_  = \new_[46792]_  & \new_[46779]_ ;
  assign \new_[2159]_  = \new_[46768]_  & \new_[46755]_ ;
  assign \new_[2160]_  = \new_[46744]_  & \new_[46731]_ ;
  assign \new_[2161]_  = \new_[46720]_  & \new_[46707]_ ;
  assign \new_[2162]_  = \new_[46696]_  & \new_[46683]_ ;
  assign \new_[2163]_  = \new_[46672]_  & \new_[46659]_ ;
  assign \new_[2164]_  = \new_[46648]_  & \new_[46635]_ ;
  assign \new_[2165]_  = \new_[46624]_  & \new_[46611]_ ;
  assign \new_[2166]_  = \new_[46600]_  & \new_[46587]_ ;
  assign \new_[2167]_  = \new_[46576]_  & \new_[46563]_ ;
  assign \new_[2168]_  = \new_[46552]_  & \new_[46539]_ ;
  assign \new_[2169]_  = \new_[46528]_  & \new_[46515]_ ;
  assign \new_[2170]_  = \new_[46504]_  & \new_[46491]_ ;
  assign \new_[2171]_  = \new_[46480]_  & \new_[46467]_ ;
  assign \new_[2172]_  = \new_[46456]_  & \new_[46443]_ ;
  assign \new_[2173]_  = \new_[46432]_  & \new_[46419]_ ;
  assign \new_[2174]_  = \new_[46408]_  & \new_[46395]_ ;
  assign \new_[2175]_  = \new_[46384]_  & \new_[46371]_ ;
  assign \new_[2176]_  = \new_[46360]_  & \new_[46347]_ ;
  assign \new_[2177]_  = \new_[46336]_  & \new_[46323]_ ;
  assign \new_[2178]_  = \new_[46312]_  & \new_[46299]_ ;
  assign \new_[2179]_  = \new_[46288]_  & \new_[46275]_ ;
  assign \new_[2180]_  = \new_[46264]_  & \new_[46251]_ ;
  assign \new_[2181]_  = \new_[46240]_  & \new_[46227]_ ;
  assign \new_[2182]_  = \new_[46216]_  & \new_[46203]_ ;
  assign \new_[2183]_  = \new_[46192]_  & \new_[46179]_ ;
  assign \new_[2184]_  = \new_[46168]_  & \new_[46155]_ ;
  assign \new_[2185]_  = \new_[46144]_  & \new_[46131]_ ;
  assign \new_[2186]_  = \new_[46120]_  & \new_[46107]_ ;
  assign \new_[2187]_  = \new_[46096]_  & \new_[46083]_ ;
  assign \new_[2188]_  = \new_[46072]_  & \new_[46059]_ ;
  assign \new_[2189]_  = \new_[46048]_  & \new_[46035]_ ;
  assign \new_[2190]_  = \new_[46024]_  & \new_[46011]_ ;
  assign \new_[2191]_  = \new_[46000]_  & \new_[45987]_ ;
  assign \new_[2192]_  = \new_[45976]_  & \new_[45963]_ ;
  assign \new_[2193]_  = \new_[45952]_  & \new_[45939]_ ;
  assign \new_[2194]_  = \new_[45928]_  & \new_[45915]_ ;
  assign \new_[2195]_  = \new_[45904]_  & \new_[45891]_ ;
  assign \new_[2196]_  = \new_[45880]_  & \new_[45867]_ ;
  assign \new_[2197]_  = \new_[45856]_  & \new_[45843]_ ;
  assign \new_[2198]_  = \new_[45832]_  & \new_[45819]_ ;
  assign \new_[2199]_  = \new_[45808]_  & \new_[45795]_ ;
  assign \new_[2200]_  = \new_[45784]_  & \new_[45771]_ ;
  assign \new_[2201]_  = \new_[45760]_  & \new_[45747]_ ;
  assign \new_[2202]_  = \new_[45736]_  & \new_[45723]_ ;
  assign \new_[2203]_  = \new_[45712]_  & \new_[45699]_ ;
  assign \new_[2204]_  = \new_[45688]_  & \new_[45675]_ ;
  assign \new_[2205]_  = \new_[45664]_  & \new_[45651]_ ;
  assign \new_[2206]_  = \new_[45640]_  & \new_[45627]_ ;
  assign \new_[2207]_  = \new_[45616]_  & \new_[45603]_ ;
  assign \new_[2208]_  = \new_[45592]_  & \new_[45579]_ ;
  assign \new_[2209]_  = \new_[45568]_  & \new_[45555]_ ;
  assign \new_[2210]_  = \new_[45544]_  & \new_[45531]_ ;
  assign \new_[2211]_  = \new_[45520]_  & \new_[45507]_ ;
  assign \new_[2212]_  = \new_[45496]_  & \new_[45483]_ ;
  assign \new_[2213]_  = \new_[45472]_  & \new_[45459]_ ;
  assign \new_[2214]_  = \new_[45448]_  & \new_[45435]_ ;
  assign \new_[2215]_  = \new_[45424]_  & \new_[45411]_ ;
  assign \new_[2216]_  = \new_[45400]_  & \new_[45387]_ ;
  assign \new_[2217]_  = \new_[45376]_  & \new_[45363]_ ;
  assign \new_[2218]_  = \new_[45352]_  & \new_[45339]_ ;
  assign \new_[2219]_  = \new_[45328]_  & \new_[45315]_ ;
  assign \new_[2220]_  = \new_[45304]_  & \new_[45291]_ ;
  assign \new_[2221]_  = \new_[45280]_  & \new_[45267]_ ;
  assign \new_[2222]_  = \new_[45256]_  & \new_[45243]_ ;
  assign \new_[2223]_  = \new_[45232]_  & \new_[45219]_ ;
  assign \new_[2224]_  = \new_[45208]_  & \new_[45195]_ ;
  assign \new_[2225]_  = \new_[45184]_  & \new_[45171]_ ;
  assign \new_[2226]_  = \new_[45160]_  & \new_[45147]_ ;
  assign \new_[2227]_  = \new_[45136]_  & \new_[45123]_ ;
  assign \new_[2228]_  = \new_[45112]_  & \new_[45099]_ ;
  assign \new_[2229]_  = \new_[45088]_  & \new_[45075]_ ;
  assign \new_[2230]_  = \new_[45064]_  & \new_[45051]_ ;
  assign \new_[2231]_  = \new_[45040]_  & \new_[45027]_ ;
  assign \new_[2232]_  = \new_[45016]_  & \new_[45003]_ ;
  assign \new_[2233]_  = \new_[44992]_  & \new_[44979]_ ;
  assign \new_[2234]_  = \new_[44968]_  & \new_[44955]_ ;
  assign \new_[2235]_  = \new_[44944]_  & \new_[44931]_ ;
  assign \new_[2236]_  = \new_[44920]_  & \new_[44907]_ ;
  assign \new_[2237]_  = \new_[44896]_  & \new_[44883]_ ;
  assign \new_[2238]_  = \new_[44872]_  & \new_[44859]_ ;
  assign \new_[2239]_  = \new_[44848]_  & \new_[44835]_ ;
  assign \new_[2240]_  = \new_[44824]_  & \new_[44811]_ ;
  assign \new_[2241]_  = \new_[44800]_  & \new_[44787]_ ;
  assign \new_[2242]_  = \new_[44776]_  & \new_[44763]_ ;
  assign \new_[2243]_  = \new_[44752]_  & \new_[44739]_ ;
  assign \new_[2244]_  = \new_[44728]_  & \new_[44715]_ ;
  assign \new_[2245]_  = \new_[44704]_  & \new_[44691]_ ;
  assign \new_[2246]_  = \new_[44680]_  & \new_[44667]_ ;
  assign \new_[2247]_  = \new_[44656]_  & \new_[44643]_ ;
  assign \new_[2248]_  = \new_[44632]_  & \new_[44619]_ ;
  assign \new_[2249]_  = \new_[44608]_  & \new_[44595]_ ;
  assign \new_[2250]_  = \new_[44584]_  & \new_[44571]_ ;
  assign \new_[2251]_  = \new_[44560]_  & \new_[44547]_ ;
  assign \new_[2252]_  = \new_[44536]_  & \new_[44523]_ ;
  assign \new_[2253]_  = \new_[44512]_  & \new_[44499]_ ;
  assign \new_[2254]_  = \new_[44488]_  & \new_[44475]_ ;
  assign \new_[2255]_  = \new_[44464]_  & \new_[44451]_ ;
  assign \new_[2256]_  = \new_[44440]_  & \new_[44427]_ ;
  assign \new_[2257]_  = \new_[44416]_  & \new_[44403]_ ;
  assign \new_[2258]_  = \new_[44392]_  & \new_[44379]_ ;
  assign \new_[2259]_  = \new_[44368]_  & \new_[44355]_ ;
  assign \new_[2260]_  = \new_[44344]_  & \new_[44331]_ ;
  assign \new_[2261]_  = \new_[44320]_  & \new_[44307]_ ;
  assign \new_[2262]_  = \new_[44296]_  & \new_[44283]_ ;
  assign \new_[2263]_  = \new_[44272]_  & \new_[44259]_ ;
  assign \new_[2264]_  = \new_[44248]_  & \new_[44235]_ ;
  assign \new_[2265]_  = \new_[44224]_  & \new_[44211]_ ;
  assign \new_[2266]_  = \new_[44200]_  & \new_[44187]_ ;
  assign \new_[2267]_  = \new_[44176]_  & \new_[44163]_ ;
  assign \new_[2268]_  = \new_[44152]_  & \new_[44139]_ ;
  assign \new_[2269]_  = \new_[44128]_  & \new_[44115]_ ;
  assign \new_[2270]_  = \new_[44104]_  & \new_[44091]_ ;
  assign \new_[2271]_  = \new_[44080]_  & \new_[44067]_ ;
  assign \new_[2272]_  = \new_[44056]_  & \new_[44043]_ ;
  assign \new_[2273]_  = \new_[44032]_  & \new_[44019]_ ;
  assign \new_[2274]_  = \new_[44008]_  & \new_[43995]_ ;
  assign \new_[2275]_  = \new_[43984]_  & \new_[43971]_ ;
  assign \new_[2276]_  = \new_[43960]_  & \new_[43947]_ ;
  assign \new_[2277]_  = \new_[43936]_  & \new_[43923]_ ;
  assign \new_[2278]_  = \new_[43912]_  & \new_[43899]_ ;
  assign \new_[2279]_  = \new_[43888]_  & \new_[43875]_ ;
  assign \new_[2280]_  = \new_[43864]_  & \new_[43851]_ ;
  assign \new_[2281]_  = \new_[43840]_  & \new_[43827]_ ;
  assign \new_[2282]_  = \new_[43816]_  & \new_[43803]_ ;
  assign \new_[2283]_  = \new_[43792]_  & \new_[43779]_ ;
  assign \new_[2284]_  = \new_[43768]_  & \new_[43755]_ ;
  assign \new_[2285]_  = \new_[43744]_  & \new_[43731]_ ;
  assign \new_[2286]_  = \new_[43720]_  & \new_[43707]_ ;
  assign \new_[2287]_  = \new_[43696]_  & \new_[43683]_ ;
  assign \new_[2288]_  = \new_[43672]_  & \new_[43659]_ ;
  assign \new_[2289]_  = \new_[43648]_  & \new_[43635]_ ;
  assign \new_[2290]_  = \new_[43624]_  & \new_[43611]_ ;
  assign \new_[2291]_  = \new_[43600]_  & \new_[43587]_ ;
  assign \new_[2292]_  = \new_[43576]_  & \new_[43563]_ ;
  assign \new_[2293]_  = \new_[43552]_  & \new_[43539]_ ;
  assign \new_[2294]_  = \new_[43528]_  & \new_[43515]_ ;
  assign \new_[2295]_  = \new_[43504]_  & \new_[43491]_ ;
  assign \new_[2296]_  = \new_[43480]_  & \new_[43467]_ ;
  assign \new_[2297]_  = \new_[43456]_  & \new_[43443]_ ;
  assign \new_[2298]_  = \new_[43432]_  & \new_[43419]_ ;
  assign \new_[2299]_  = \new_[43408]_  & \new_[43395]_ ;
  assign \new_[2300]_  = \new_[43384]_  & \new_[43371]_ ;
  assign \new_[2301]_  = \new_[43360]_  & \new_[43347]_ ;
  assign \new_[2302]_  = \new_[43336]_  & \new_[43323]_ ;
  assign \new_[2303]_  = \new_[43312]_  & \new_[43299]_ ;
  assign \new_[2304]_  = \new_[43288]_  & \new_[43275]_ ;
  assign \new_[2305]_  = \new_[43264]_  & \new_[43251]_ ;
  assign \new_[2306]_  = \new_[43240]_  & \new_[43227]_ ;
  assign \new_[2307]_  = \new_[43216]_  & \new_[43203]_ ;
  assign \new_[2308]_  = \new_[43192]_  & \new_[43179]_ ;
  assign \new_[2309]_  = \new_[43168]_  & \new_[43155]_ ;
  assign \new_[2310]_  = \new_[43144]_  & \new_[43131]_ ;
  assign \new_[2311]_  = \new_[43120]_  & \new_[43107]_ ;
  assign \new_[2312]_  = \new_[43096]_  & \new_[43083]_ ;
  assign \new_[2313]_  = \new_[43072]_  & \new_[43059]_ ;
  assign \new_[2314]_  = \new_[43048]_  & \new_[43035]_ ;
  assign \new_[2315]_  = \new_[43024]_  & \new_[43011]_ ;
  assign \new_[2316]_  = \new_[43000]_  & \new_[42987]_ ;
  assign \new_[2317]_  = \new_[42976]_  & \new_[42963]_ ;
  assign \new_[2318]_  = \new_[42952]_  & \new_[42939]_ ;
  assign \new_[2319]_  = \new_[42928]_  & \new_[42915]_ ;
  assign \new_[2320]_  = \new_[42904]_  & \new_[42891]_ ;
  assign \new_[2321]_  = \new_[42880]_  & \new_[42867]_ ;
  assign \new_[2322]_  = \new_[42856]_  & \new_[42843]_ ;
  assign \new_[2323]_  = \new_[42832]_  & \new_[42819]_ ;
  assign \new_[2324]_  = \new_[42808]_  & \new_[42795]_ ;
  assign \new_[2325]_  = \new_[42784]_  & \new_[42771]_ ;
  assign \new_[2326]_  = \new_[42760]_  & \new_[42747]_ ;
  assign \new_[2327]_  = \new_[42736]_  & \new_[42723]_ ;
  assign \new_[2328]_  = \new_[42712]_  & \new_[42699]_ ;
  assign \new_[2329]_  = \new_[42688]_  & \new_[42675]_ ;
  assign \new_[2330]_  = \new_[42664]_  & \new_[42651]_ ;
  assign \new_[2331]_  = \new_[42640]_  & \new_[42627]_ ;
  assign \new_[2332]_  = \new_[42616]_  & \new_[42603]_ ;
  assign \new_[2333]_  = \new_[42592]_  & \new_[42579]_ ;
  assign \new_[2334]_  = \new_[42568]_  & \new_[42555]_ ;
  assign \new_[2335]_  = \new_[42544]_  & \new_[42531]_ ;
  assign \new_[2336]_  = \new_[42520]_  & \new_[42507]_ ;
  assign \new_[2337]_  = \new_[42496]_  & \new_[42483]_ ;
  assign \new_[2338]_  = \new_[42472]_  & \new_[42459]_ ;
  assign \new_[2339]_  = \new_[42448]_  & \new_[42435]_ ;
  assign \new_[2340]_  = \new_[42424]_  & \new_[42411]_ ;
  assign \new_[2341]_  = \new_[42400]_  & \new_[42387]_ ;
  assign \new_[2342]_  = \new_[42376]_  & \new_[42363]_ ;
  assign \new_[2343]_  = \new_[42352]_  & \new_[42339]_ ;
  assign \new_[2344]_  = \new_[42328]_  & \new_[42315]_ ;
  assign \new_[2345]_  = \new_[42304]_  & \new_[42291]_ ;
  assign \new_[2346]_  = \new_[42280]_  & \new_[42267]_ ;
  assign \new_[2347]_  = \new_[42256]_  & \new_[42243]_ ;
  assign \new_[2348]_  = \new_[42232]_  & \new_[42219]_ ;
  assign \new_[2349]_  = \new_[42208]_  & \new_[42195]_ ;
  assign \new_[2350]_  = \new_[42184]_  & \new_[42171]_ ;
  assign \new_[2351]_  = \new_[42160]_  & \new_[42147]_ ;
  assign \new_[2352]_  = \new_[42136]_  & \new_[42123]_ ;
  assign \new_[2353]_  = \new_[42112]_  & \new_[42099]_ ;
  assign \new_[2354]_  = \new_[42088]_  & \new_[42075]_ ;
  assign \new_[2355]_  = \new_[42064]_  & \new_[42051]_ ;
  assign \new_[2356]_  = \new_[42040]_  & \new_[42027]_ ;
  assign \new_[2357]_  = \new_[42016]_  & \new_[42003]_ ;
  assign \new_[2358]_  = \new_[41992]_  & \new_[41979]_ ;
  assign \new_[2359]_  = \new_[41968]_  & \new_[41955]_ ;
  assign \new_[2360]_  = \new_[41944]_  & \new_[41931]_ ;
  assign \new_[2361]_  = \new_[41920]_  & \new_[41907]_ ;
  assign \new_[2362]_  = \new_[41896]_  & \new_[41883]_ ;
  assign \new_[2363]_  = \new_[41872]_  & \new_[41859]_ ;
  assign \new_[2364]_  = \new_[41848]_  & \new_[41835]_ ;
  assign \new_[2365]_  = \new_[41824]_  & \new_[41811]_ ;
  assign \new_[2366]_  = \new_[41800]_  & \new_[41787]_ ;
  assign \new_[2367]_  = \new_[41776]_  & \new_[41763]_ ;
  assign \new_[2368]_  = \new_[41752]_  & \new_[41739]_ ;
  assign \new_[2369]_  = \new_[41728]_  & \new_[41715]_ ;
  assign \new_[2370]_  = \new_[41704]_  & \new_[41691]_ ;
  assign \new_[2371]_  = \new_[41680]_  & \new_[41667]_ ;
  assign \new_[2372]_  = \new_[41656]_  & \new_[41643]_ ;
  assign \new_[2373]_  = \new_[41632]_  & \new_[41619]_ ;
  assign \new_[2374]_  = \new_[41608]_  & \new_[41595]_ ;
  assign \new_[2375]_  = \new_[41584]_  & \new_[41571]_ ;
  assign \new_[2376]_  = \new_[41560]_  & \new_[41547]_ ;
  assign \new_[2377]_  = \new_[41536]_  & \new_[41523]_ ;
  assign \new_[2378]_  = \new_[41512]_  & \new_[41499]_ ;
  assign \new_[2379]_  = \new_[41488]_  & \new_[41475]_ ;
  assign \new_[2380]_  = \new_[41464]_  & \new_[41451]_ ;
  assign \new_[2381]_  = \new_[41440]_  & \new_[41427]_ ;
  assign \new_[2382]_  = \new_[41416]_  & \new_[41403]_ ;
  assign \new_[2383]_  = \new_[41392]_  & \new_[41379]_ ;
  assign \new_[2384]_  = \new_[41368]_  & \new_[41355]_ ;
  assign \new_[2385]_  = \new_[41344]_  & \new_[41331]_ ;
  assign \new_[2386]_  = \new_[41320]_  & \new_[41307]_ ;
  assign \new_[2387]_  = \new_[41296]_  & \new_[41283]_ ;
  assign \new_[2388]_  = \new_[41272]_  & \new_[41259]_ ;
  assign \new_[2389]_  = \new_[41248]_  & \new_[41235]_ ;
  assign \new_[2390]_  = \new_[41224]_  & \new_[41211]_ ;
  assign \new_[2391]_  = \new_[41200]_  & \new_[41187]_ ;
  assign \new_[2392]_  = \new_[41176]_  & \new_[41163]_ ;
  assign \new_[2393]_  = \new_[41152]_  & \new_[41139]_ ;
  assign \new_[2394]_  = \new_[41128]_  & \new_[41115]_ ;
  assign \new_[2395]_  = \new_[41104]_  & \new_[41091]_ ;
  assign \new_[2396]_  = \new_[41080]_  & \new_[41067]_ ;
  assign \new_[2397]_  = \new_[41056]_  & \new_[41043]_ ;
  assign \new_[2398]_  = \new_[41032]_  & \new_[41019]_ ;
  assign \new_[2399]_  = \new_[41008]_  & \new_[40995]_ ;
  assign \new_[2400]_  = \new_[40984]_  & \new_[40971]_ ;
  assign \new_[2401]_  = \new_[40960]_  & \new_[40947]_ ;
  assign \new_[2402]_  = \new_[40936]_  & \new_[40923]_ ;
  assign \new_[2403]_  = \new_[40912]_  & \new_[40899]_ ;
  assign \new_[2404]_  = \new_[40888]_  & \new_[40875]_ ;
  assign \new_[2405]_  = \new_[40864]_  & \new_[40851]_ ;
  assign \new_[2406]_  = \new_[40840]_  & \new_[40827]_ ;
  assign \new_[2407]_  = \new_[40816]_  & \new_[40803]_ ;
  assign \new_[2408]_  = \new_[40792]_  & \new_[40779]_ ;
  assign \new_[2409]_  = \new_[40768]_  & \new_[40755]_ ;
  assign \new_[2410]_  = \new_[40744]_  & \new_[40731]_ ;
  assign \new_[2411]_  = \new_[40720]_  & \new_[40707]_ ;
  assign \new_[2412]_  = \new_[40696]_  & \new_[40683]_ ;
  assign \new_[2413]_  = \new_[40672]_  & \new_[40659]_ ;
  assign \new_[2414]_  = \new_[40648]_  & \new_[40635]_ ;
  assign \new_[2415]_  = \new_[40624]_  & \new_[40611]_ ;
  assign \new_[2416]_  = \new_[40600]_  & \new_[40587]_ ;
  assign \new_[2417]_  = \new_[40576]_  & \new_[40563]_ ;
  assign \new_[2418]_  = \new_[40552]_  & \new_[40539]_ ;
  assign \new_[2419]_  = \new_[40528]_  & \new_[40515]_ ;
  assign \new_[2420]_  = \new_[40504]_  & \new_[40491]_ ;
  assign \new_[2421]_  = \new_[40480]_  & \new_[40467]_ ;
  assign \new_[2422]_  = \new_[40456]_  & \new_[40443]_ ;
  assign \new_[2423]_  = \new_[40432]_  & \new_[40419]_ ;
  assign \new_[2424]_  = \new_[40408]_  & \new_[40395]_ ;
  assign \new_[2425]_  = \new_[40384]_  & \new_[40371]_ ;
  assign \new_[2426]_  = \new_[40360]_  & \new_[40347]_ ;
  assign \new_[2427]_  = \new_[40336]_  & \new_[40325]_ ;
  assign \new_[2428]_  = \new_[40314]_  & \new_[40303]_ ;
  assign \new_[2429]_  = \new_[40292]_  & \new_[40281]_ ;
  assign \new_[2430]_  = \new_[40270]_  & \new_[40259]_ ;
  assign \new_[2431]_  = \new_[40248]_  & \new_[40237]_ ;
  assign \new_[2432]_  = \new_[40226]_  & \new_[40215]_ ;
  assign \new_[2433]_  = \new_[40204]_  & \new_[40193]_ ;
  assign \new_[2434]_  = \new_[40182]_  & \new_[40171]_ ;
  assign \new_[2435]_  = \new_[40160]_  & \new_[40149]_ ;
  assign \new_[2436]_  = \new_[40138]_  & \new_[40127]_ ;
  assign \new_[2437]_  = \new_[40116]_  & \new_[40105]_ ;
  assign \new_[2438]_  = \new_[40094]_  & \new_[40083]_ ;
  assign \new_[2439]_  = \new_[40072]_  & \new_[40061]_ ;
  assign \new_[2440]_  = \new_[40050]_  & \new_[40039]_ ;
  assign \new_[2441]_  = \new_[40028]_  & \new_[40017]_ ;
  assign \new_[2442]_  = \new_[40006]_  & \new_[39995]_ ;
  assign \new_[2443]_  = \new_[39984]_  & \new_[39973]_ ;
  assign \new_[2444]_  = \new_[39962]_  & \new_[39951]_ ;
  assign \new_[2445]_  = \new_[39940]_  & \new_[39929]_ ;
  assign \new_[2446]_  = \new_[39918]_  & \new_[39907]_ ;
  assign \new_[2447]_  = \new_[39896]_  & \new_[39885]_ ;
  assign \new_[2448]_  = \new_[39874]_  & \new_[39863]_ ;
  assign \new_[2449]_  = \new_[39852]_  & \new_[39841]_ ;
  assign \new_[2450]_  = \new_[39830]_  & \new_[39819]_ ;
  assign \new_[2451]_  = \new_[39808]_  & \new_[39797]_ ;
  assign \new_[2452]_  = \new_[39786]_  & \new_[39775]_ ;
  assign \new_[2453]_  = \new_[39764]_  & \new_[39753]_ ;
  assign \new_[2454]_  = \new_[39742]_  & \new_[39731]_ ;
  assign \new_[2455]_  = \new_[39720]_  & \new_[39709]_ ;
  assign \new_[2456]_  = \new_[39698]_  & \new_[39687]_ ;
  assign \new_[2457]_  = \new_[39676]_  & \new_[39665]_ ;
  assign \new_[2458]_  = \new_[39654]_  & \new_[39643]_ ;
  assign \new_[2459]_  = \new_[39632]_  & \new_[39621]_ ;
  assign \new_[2460]_  = \new_[39610]_  & \new_[39599]_ ;
  assign \new_[2461]_  = \new_[39588]_  & \new_[39577]_ ;
  assign \new_[2462]_  = \new_[39566]_  & \new_[39555]_ ;
  assign \new_[2463]_  = \new_[39544]_  & \new_[39533]_ ;
  assign \new_[2464]_  = \new_[39522]_  & \new_[39511]_ ;
  assign \new_[2465]_  = \new_[39500]_  & \new_[39489]_ ;
  assign \new_[2466]_  = \new_[39478]_  & \new_[39467]_ ;
  assign \new_[2467]_  = \new_[39456]_  & \new_[39445]_ ;
  assign \new_[2468]_  = \new_[39434]_  & \new_[39423]_ ;
  assign \new_[2469]_  = \new_[39412]_  & \new_[39401]_ ;
  assign \new_[2470]_  = \new_[39390]_  & \new_[39379]_ ;
  assign \new_[2471]_  = \new_[39368]_  & \new_[39357]_ ;
  assign \new_[2472]_  = \new_[39346]_  & \new_[39335]_ ;
  assign \new_[2473]_  = \new_[39324]_  & \new_[39313]_ ;
  assign \new_[2474]_  = \new_[39302]_  & \new_[39291]_ ;
  assign \new_[2475]_  = \new_[39280]_  & \new_[39269]_ ;
  assign \new_[2476]_  = \new_[39258]_  & \new_[39247]_ ;
  assign \new_[2477]_  = \new_[39236]_  & \new_[39225]_ ;
  assign \new_[2478]_  = \new_[39214]_  & \new_[39203]_ ;
  assign \new_[2479]_  = \new_[39192]_  & \new_[39181]_ ;
  assign \new_[2480]_  = \new_[39170]_  & \new_[39159]_ ;
  assign \new_[2481]_  = \new_[39148]_  & \new_[39137]_ ;
  assign \new_[2482]_  = \new_[39126]_  & \new_[39115]_ ;
  assign \new_[2483]_  = \new_[39104]_  & \new_[39093]_ ;
  assign \new_[2484]_  = \new_[39082]_  & \new_[39071]_ ;
  assign \new_[2485]_  = \new_[39060]_  & \new_[39049]_ ;
  assign \new_[2486]_  = \new_[39038]_  & \new_[39027]_ ;
  assign \new_[2487]_  = \new_[39016]_  & \new_[39005]_ ;
  assign \new_[2488]_  = \new_[38994]_  & \new_[38983]_ ;
  assign \new_[2489]_  = \new_[38972]_  & \new_[38961]_ ;
  assign \new_[2490]_  = \new_[38950]_  & \new_[38939]_ ;
  assign \new_[2491]_  = \new_[38928]_  & \new_[38917]_ ;
  assign \new_[2492]_  = \new_[38906]_  & \new_[38895]_ ;
  assign \new_[2493]_  = \new_[38884]_  & \new_[38873]_ ;
  assign \new_[2494]_  = \new_[38862]_  & \new_[38851]_ ;
  assign \new_[2495]_  = \new_[38840]_  & \new_[38829]_ ;
  assign \new_[2496]_  = \new_[38818]_  & \new_[38807]_ ;
  assign \new_[2497]_  = \new_[38796]_  & \new_[38785]_ ;
  assign \new_[2498]_  = \new_[38774]_  & \new_[38763]_ ;
  assign \new_[2499]_  = \new_[38752]_  & \new_[38741]_ ;
  assign \new_[2500]_  = \new_[38730]_  & \new_[38719]_ ;
  assign \new_[2501]_  = \new_[38708]_  & \new_[38697]_ ;
  assign \new_[2502]_  = \new_[38686]_  & \new_[38675]_ ;
  assign \new_[2503]_  = \new_[38664]_  & \new_[38653]_ ;
  assign \new_[2504]_  = \new_[38642]_  & \new_[38631]_ ;
  assign \new_[2505]_  = \new_[38620]_  & \new_[38609]_ ;
  assign \new_[2506]_  = \new_[38598]_  & \new_[38587]_ ;
  assign \new_[2507]_  = \new_[38576]_  & \new_[38565]_ ;
  assign \new_[2508]_  = \new_[38554]_  & \new_[38543]_ ;
  assign \new_[2509]_  = \new_[38532]_  & \new_[38521]_ ;
  assign \new_[2510]_  = \new_[38510]_  & \new_[38499]_ ;
  assign \new_[2511]_  = \new_[38488]_  & \new_[38477]_ ;
  assign \new_[2512]_  = \new_[38466]_  & \new_[38455]_ ;
  assign \new_[2513]_  = \new_[38444]_  & \new_[38433]_ ;
  assign \new_[2514]_  = \new_[38422]_  & \new_[38411]_ ;
  assign \new_[2515]_  = \new_[38400]_  & \new_[38389]_ ;
  assign \new_[2516]_  = \new_[38378]_  & \new_[38367]_ ;
  assign \new_[2517]_  = \new_[38356]_  & \new_[38345]_ ;
  assign \new_[2518]_  = \new_[38334]_  & \new_[38323]_ ;
  assign \new_[2519]_  = \new_[38312]_  & \new_[38301]_ ;
  assign \new_[2520]_  = \new_[38290]_  & \new_[38279]_ ;
  assign \new_[2521]_  = \new_[38268]_  & \new_[38257]_ ;
  assign \new_[2522]_  = \new_[38246]_  & \new_[38235]_ ;
  assign \new_[2523]_  = \new_[38224]_  & \new_[38213]_ ;
  assign \new_[2524]_  = \new_[38202]_  & \new_[38191]_ ;
  assign \new_[2525]_  = \new_[38180]_  & \new_[38169]_ ;
  assign \new_[2526]_  = \new_[38158]_  & \new_[38147]_ ;
  assign \new_[2527]_  = \new_[38136]_  & \new_[38125]_ ;
  assign \new_[2528]_  = \new_[38114]_  & \new_[38103]_ ;
  assign \new_[2529]_  = \new_[38092]_  & \new_[38081]_ ;
  assign \new_[2530]_  = \new_[38070]_  & \new_[38059]_ ;
  assign \new_[2531]_  = \new_[38048]_  & \new_[38037]_ ;
  assign \new_[2532]_  = \new_[38026]_  & \new_[38015]_ ;
  assign \new_[2533]_  = \new_[38004]_  & \new_[37993]_ ;
  assign \new_[2534]_  = \new_[37982]_  & \new_[37971]_ ;
  assign \new_[2535]_  = \new_[37960]_  & \new_[37949]_ ;
  assign \new_[2536]_  = \new_[37938]_  & \new_[37927]_ ;
  assign \new_[2537]_  = \new_[37916]_  & \new_[37905]_ ;
  assign \new_[2538]_  = \new_[37894]_  & \new_[37883]_ ;
  assign \new_[2539]_  = \new_[37872]_  & \new_[37861]_ ;
  assign \new_[2540]_  = \new_[37850]_  & \new_[37839]_ ;
  assign \new_[2541]_  = \new_[37828]_  & \new_[37817]_ ;
  assign \new_[2542]_  = \new_[37806]_  & \new_[37795]_ ;
  assign \new_[2543]_  = \new_[37784]_  & \new_[37773]_ ;
  assign \new_[2544]_  = \new_[37762]_  & \new_[37751]_ ;
  assign \new_[2545]_  = \new_[37740]_  & \new_[37729]_ ;
  assign \new_[2546]_  = \new_[37718]_  & \new_[37707]_ ;
  assign \new_[2547]_  = \new_[37696]_  & \new_[37685]_ ;
  assign \new_[2548]_  = \new_[37674]_  & \new_[37663]_ ;
  assign \new_[2549]_  = \new_[37652]_  & \new_[37641]_ ;
  assign \new_[2550]_  = \new_[37630]_  & \new_[37619]_ ;
  assign \new_[2551]_  = \new_[37608]_  & \new_[37597]_ ;
  assign \new_[2552]_  = \new_[37586]_  & \new_[37575]_ ;
  assign \new_[2553]_  = \new_[37564]_  & \new_[37553]_ ;
  assign \new_[2554]_  = \new_[37542]_  & \new_[37531]_ ;
  assign \new_[2555]_  = \new_[37520]_  & \new_[37509]_ ;
  assign \new_[2556]_  = \new_[37498]_  & \new_[37487]_ ;
  assign \new_[2557]_  = \new_[37476]_  & \new_[37465]_ ;
  assign \new_[2558]_  = \new_[37454]_  & \new_[37443]_ ;
  assign \new_[2559]_  = \new_[37432]_  & \new_[37421]_ ;
  assign \new_[2560]_  = \new_[37410]_  & \new_[37399]_ ;
  assign \new_[2561]_  = \new_[37388]_  & \new_[37377]_ ;
  assign \new_[2562]_  = \new_[37366]_  & \new_[37355]_ ;
  assign \new_[2563]_  = \new_[37344]_  & \new_[37333]_ ;
  assign \new_[2564]_  = \new_[37322]_  & \new_[37311]_ ;
  assign \new_[2565]_  = \new_[37300]_  & \new_[37289]_ ;
  assign \new_[2566]_  = \new_[37278]_  & \new_[37267]_ ;
  assign \new_[2567]_  = \new_[37256]_  & \new_[37245]_ ;
  assign \new_[2568]_  = \new_[37234]_  & \new_[37223]_ ;
  assign \new_[2569]_  = \new_[37212]_  & \new_[37201]_ ;
  assign \new_[2570]_  = \new_[37190]_  & \new_[37179]_ ;
  assign \new_[2571]_  = \new_[37168]_  & \new_[37157]_ ;
  assign \new_[2572]_  = \new_[37146]_  & \new_[37135]_ ;
  assign \new_[2573]_  = \new_[37124]_  & \new_[37113]_ ;
  assign \new_[2574]_  = \new_[37102]_  & \new_[37091]_ ;
  assign \new_[2575]_  = \new_[37080]_  & \new_[37069]_ ;
  assign \new_[2576]_  = \new_[37058]_  & \new_[37047]_ ;
  assign \new_[2577]_  = \new_[37036]_  & \new_[37025]_ ;
  assign \new_[2578]_  = \new_[37014]_  & \new_[37003]_ ;
  assign \new_[2579]_  = \new_[36992]_  & \new_[36981]_ ;
  assign \new_[2580]_  = \new_[36970]_  & \new_[36959]_ ;
  assign \new_[2581]_  = \new_[36948]_  & \new_[36937]_ ;
  assign \new_[2582]_  = \new_[36926]_  & \new_[36915]_ ;
  assign \new_[2583]_  = \new_[36904]_  & \new_[36893]_ ;
  assign \new_[2584]_  = \new_[36882]_  & \new_[36871]_ ;
  assign \new_[2585]_  = \new_[36860]_  & \new_[36849]_ ;
  assign \new_[2586]_  = \new_[36838]_  & \new_[36827]_ ;
  assign \new_[2587]_  = \new_[36816]_  & \new_[36805]_ ;
  assign \new_[2588]_  = \new_[36794]_  & \new_[36783]_ ;
  assign \new_[2589]_  = \new_[36772]_  & \new_[36761]_ ;
  assign \new_[2590]_  = \new_[36750]_  & \new_[36739]_ ;
  assign \new_[2591]_  = \new_[36728]_  & \new_[36717]_ ;
  assign \new_[2592]_  = \new_[36706]_  & \new_[36695]_ ;
  assign \new_[2593]_  = \new_[36684]_  & \new_[36673]_ ;
  assign \new_[2594]_  = \new_[36662]_  & \new_[36651]_ ;
  assign \new_[2595]_  = \new_[36640]_  & \new_[36629]_ ;
  assign \new_[2596]_  = \new_[36618]_  & \new_[36607]_ ;
  assign \new_[2597]_  = \new_[36596]_  & \new_[36585]_ ;
  assign \new_[2598]_  = \new_[36574]_  & \new_[36563]_ ;
  assign \new_[2599]_  = \new_[36552]_  & \new_[36541]_ ;
  assign \new_[2600]_  = \new_[36530]_  & \new_[36519]_ ;
  assign \new_[2601]_  = \new_[36508]_  & \new_[36497]_ ;
  assign \new_[2602]_  = \new_[36486]_  & \new_[36475]_ ;
  assign \new_[2603]_  = \new_[36464]_  & \new_[36453]_ ;
  assign \new_[2604]_  = \new_[36442]_  & \new_[36431]_ ;
  assign \new_[2605]_  = \new_[36420]_  & \new_[36409]_ ;
  assign \new_[2606]_  = \new_[36398]_  & \new_[36387]_ ;
  assign \new_[2607]_  = \new_[36376]_  & \new_[36365]_ ;
  assign \new_[2608]_  = \new_[36354]_  & \new_[36343]_ ;
  assign \new_[2609]_  = \new_[36332]_  & \new_[36321]_ ;
  assign \new_[2610]_  = \new_[36310]_  & \new_[36299]_ ;
  assign \new_[2611]_  = \new_[36288]_  & \new_[36277]_ ;
  assign \new_[2612]_  = \new_[36266]_  & \new_[36255]_ ;
  assign \new_[2613]_  = \new_[36244]_  & \new_[36233]_ ;
  assign \new_[2614]_  = \new_[36222]_  & \new_[36211]_ ;
  assign \new_[2615]_  = \new_[36200]_  & \new_[36189]_ ;
  assign \new_[2616]_  = \new_[36178]_  & \new_[36167]_ ;
  assign \new_[2617]_  = \new_[36156]_  & \new_[36145]_ ;
  assign \new_[2618]_  = \new_[36134]_  & \new_[36123]_ ;
  assign \new_[2619]_  = \new_[36112]_  & \new_[36101]_ ;
  assign \new_[2620]_  = \new_[36090]_  & \new_[36079]_ ;
  assign \new_[2621]_  = \new_[36068]_  & \new_[36057]_ ;
  assign \new_[2622]_  = \new_[36046]_  & \new_[36035]_ ;
  assign \new_[2623]_  = \new_[36024]_  & \new_[36013]_ ;
  assign \new_[2624]_  = \new_[36002]_  & \new_[35991]_ ;
  assign \new_[2625]_  = \new_[35980]_  & \new_[35969]_ ;
  assign \new_[2626]_  = \new_[35958]_  & \new_[35947]_ ;
  assign \new_[2627]_  = \new_[35936]_  & \new_[35925]_ ;
  assign \new_[2628]_  = \new_[35914]_  & \new_[35903]_ ;
  assign \new_[2629]_  = \new_[35892]_  & \new_[35881]_ ;
  assign \new_[2630]_  = \new_[35870]_  & \new_[35859]_ ;
  assign \new_[2631]_  = \new_[35848]_  & \new_[35837]_ ;
  assign \new_[2632]_  = \new_[35826]_  & \new_[35815]_ ;
  assign \new_[2633]_  = \new_[35804]_  & \new_[35793]_ ;
  assign \new_[2634]_  = \new_[35782]_  & \new_[35771]_ ;
  assign \new_[2635]_  = \new_[35760]_  & \new_[35749]_ ;
  assign \new_[2636]_  = \new_[35738]_  & \new_[35727]_ ;
  assign \new_[2637]_  = \new_[35716]_  & \new_[35705]_ ;
  assign \new_[2638]_  = \new_[35694]_  & \new_[35683]_ ;
  assign \new_[2639]_  = \new_[35672]_  & \new_[35661]_ ;
  assign \new_[2640]_  = \new_[35650]_  & \new_[35639]_ ;
  assign \new_[2641]_  = \new_[35628]_  & \new_[35617]_ ;
  assign \new_[2642]_  = \new_[35606]_  & \new_[35595]_ ;
  assign \new_[2643]_  = \new_[35584]_  & \new_[35573]_ ;
  assign \new_[2644]_  = \new_[35562]_  & \new_[35551]_ ;
  assign \new_[2645]_  = \new_[35540]_  & \new_[35529]_ ;
  assign \new_[2646]_  = \new_[35518]_  & \new_[35507]_ ;
  assign \new_[2647]_  = \new_[35496]_  & \new_[35485]_ ;
  assign \new_[2648]_  = \new_[35474]_  & \new_[35463]_ ;
  assign \new_[2649]_  = \new_[35452]_  & \new_[35441]_ ;
  assign \new_[2650]_  = \new_[35430]_  & \new_[35419]_ ;
  assign \new_[2651]_  = \new_[35408]_  & \new_[35397]_ ;
  assign \new_[2652]_  = \new_[35386]_  & \new_[35375]_ ;
  assign \new_[2653]_  = \new_[35364]_  & \new_[35353]_ ;
  assign \new_[2654]_  = \new_[35342]_  & \new_[35331]_ ;
  assign \new_[2655]_  = \new_[35320]_  & \new_[35309]_ ;
  assign \new_[2656]_  = \new_[35298]_  & \new_[35287]_ ;
  assign \new_[2657]_  = \new_[35276]_  & \new_[35265]_ ;
  assign \new_[2658]_  = \new_[35254]_  & \new_[35243]_ ;
  assign \new_[2659]_  = \new_[35232]_  & \new_[35221]_ ;
  assign \new_[2660]_  = \new_[35210]_  & \new_[35199]_ ;
  assign \new_[2661]_  = \new_[35188]_  & \new_[35177]_ ;
  assign \new_[2662]_  = \new_[35166]_  & \new_[35155]_ ;
  assign \new_[2663]_  = \new_[35144]_  & \new_[35133]_ ;
  assign \new_[2664]_  = \new_[35122]_  & \new_[35111]_ ;
  assign \new_[2665]_  = \new_[35100]_  & \new_[35089]_ ;
  assign \new_[2666]_  = \new_[35078]_  & \new_[35067]_ ;
  assign \new_[2667]_  = \new_[35056]_  & \new_[35045]_ ;
  assign \new_[2668]_  = \new_[35034]_  & \new_[35023]_ ;
  assign \new_[2669]_  = \new_[35012]_  & \new_[35001]_ ;
  assign \new_[2670]_  = \new_[34990]_  & \new_[34979]_ ;
  assign \new_[2671]_  = \new_[34968]_  & \new_[34957]_ ;
  assign \new_[2672]_  = \new_[34946]_  & \new_[34935]_ ;
  assign \new_[2673]_  = \new_[34924]_  & \new_[34913]_ ;
  assign \new_[2674]_  = \new_[34902]_  & \new_[34891]_ ;
  assign \new_[2675]_  = \new_[34880]_  & \new_[34869]_ ;
  assign \new_[2676]_  = \new_[34858]_  & \new_[34847]_ ;
  assign \new_[2677]_  = \new_[34836]_  & \new_[34825]_ ;
  assign \new_[2678]_  = \new_[34814]_  & \new_[34803]_ ;
  assign \new_[2679]_  = \new_[34792]_  & \new_[34781]_ ;
  assign \new_[2680]_  = \new_[34770]_  & \new_[34759]_ ;
  assign \new_[2681]_  = \new_[34748]_  & \new_[34737]_ ;
  assign \new_[2682]_  = \new_[34726]_  & \new_[34715]_ ;
  assign \new_[2683]_  = \new_[34704]_  & \new_[34693]_ ;
  assign \new_[2684]_  = \new_[34682]_  & \new_[34671]_ ;
  assign \new_[2685]_  = \new_[34660]_  & \new_[34649]_ ;
  assign \new_[2686]_  = \new_[34638]_  & \new_[34627]_ ;
  assign \new_[2687]_  = \new_[34616]_  & \new_[34605]_ ;
  assign \new_[2688]_  = \new_[34594]_  & \new_[34583]_ ;
  assign \new_[2689]_  = \new_[34572]_  & \new_[34561]_ ;
  assign \new_[2690]_  = \new_[34550]_  & \new_[34539]_ ;
  assign \new_[2691]_  = \new_[34528]_  & \new_[34517]_ ;
  assign \new_[2692]_  = \new_[34506]_  & \new_[34495]_ ;
  assign \new_[2693]_  = \new_[34484]_  & \new_[34473]_ ;
  assign \new_[2694]_  = \new_[34462]_  & \new_[34451]_ ;
  assign \new_[2695]_  = \new_[34440]_  & \new_[34429]_ ;
  assign \new_[2696]_  = \new_[34418]_  & \new_[34407]_ ;
  assign \new_[2697]_  = \new_[34396]_  & \new_[34385]_ ;
  assign \new_[2698]_  = \new_[34374]_  & \new_[34363]_ ;
  assign \new_[2699]_  = \new_[34352]_  & \new_[34341]_ ;
  assign \new_[2700]_  = \new_[34330]_  & \new_[34319]_ ;
  assign \new_[2701]_  = \new_[34308]_  & \new_[34297]_ ;
  assign \new_[2702]_  = \new_[34286]_  & \new_[34275]_ ;
  assign \new_[2703]_  = \new_[34264]_  & \new_[34253]_ ;
  assign \new_[2704]_  = \new_[34242]_  & \new_[34231]_ ;
  assign \new_[2705]_  = \new_[34220]_  & \new_[34209]_ ;
  assign \new_[2706]_  = \new_[34198]_  & \new_[34187]_ ;
  assign \new_[2707]_  = \new_[34176]_  & \new_[34165]_ ;
  assign \new_[2708]_  = \new_[34154]_  & \new_[34143]_ ;
  assign \new_[2709]_  = \new_[34132]_  & \new_[34121]_ ;
  assign \new_[2710]_  = \new_[34110]_  & \new_[34099]_ ;
  assign \new_[2711]_  = \new_[34088]_  & \new_[34077]_ ;
  assign \new_[2712]_  = \new_[34066]_  & \new_[34055]_ ;
  assign \new_[2713]_  = \new_[34044]_  & \new_[34033]_ ;
  assign \new_[2714]_  = \new_[34022]_  & \new_[34011]_ ;
  assign \new_[2715]_  = \new_[34000]_  & \new_[33989]_ ;
  assign \new_[2716]_  = \new_[33978]_  & \new_[33967]_ ;
  assign \new_[2717]_  = \new_[33956]_  & \new_[33945]_ ;
  assign \new_[2718]_  = \new_[33934]_  & \new_[33923]_ ;
  assign \new_[2719]_  = \new_[33912]_  & \new_[33901]_ ;
  assign \new_[2720]_  = \new_[33890]_  & \new_[33879]_ ;
  assign \new_[2721]_  = \new_[33868]_  & \new_[33857]_ ;
  assign \new_[2722]_  = \new_[33846]_  & \new_[33835]_ ;
  assign \new_[2723]_  = \new_[33824]_  & \new_[33813]_ ;
  assign \new_[2724]_  = \new_[33802]_  & \new_[33791]_ ;
  assign \new_[2725]_  = \new_[33780]_  & \new_[33769]_ ;
  assign \new_[2726]_  = \new_[33758]_  & \new_[33747]_ ;
  assign \new_[2727]_  = \new_[33736]_  & \new_[33725]_ ;
  assign \new_[2728]_  = \new_[33714]_  & \new_[33703]_ ;
  assign \new_[2729]_  = \new_[33692]_  & \new_[33681]_ ;
  assign \new_[2730]_  = \new_[33670]_  & \new_[33659]_ ;
  assign \new_[2731]_  = \new_[33648]_  & \new_[33637]_ ;
  assign \new_[2732]_  = \new_[33626]_  & \new_[33615]_ ;
  assign \new_[2733]_  = \new_[33604]_  & \new_[33593]_ ;
  assign \new_[2734]_  = \new_[33582]_  & \new_[33571]_ ;
  assign \new_[2735]_  = \new_[33560]_  & \new_[33549]_ ;
  assign \new_[2736]_  = \new_[33538]_  & \new_[33527]_ ;
  assign \new_[2737]_  = \new_[33516]_  & \new_[33505]_ ;
  assign \new_[2738]_  = \new_[33494]_  & \new_[33483]_ ;
  assign \new_[2739]_  = \new_[33472]_  & \new_[33461]_ ;
  assign \new_[2740]_  = \new_[33450]_  & \new_[33439]_ ;
  assign \new_[2741]_  = \new_[33428]_  & \new_[33417]_ ;
  assign \new_[2742]_  = \new_[33406]_  & \new_[33395]_ ;
  assign \new_[2743]_  = \new_[33384]_  & \new_[33373]_ ;
  assign \new_[2744]_  = \new_[33362]_  & \new_[33351]_ ;
  assign \new_[2745]_  = \new_[33340]_  & \new_[33329]_ ;
  assign \new_[2746]_  = \new_[33318]_  & \new_[33307]_ ;
  assign \new_[2747]_  = \new_[33296]_  & \new_[33285]_ ;
  assign \new_[2748]_  = \new_[33274]_  & \new_[33263]_ ;
  assign \new_[2749]_  = \new_[33252]_  & \new_[33241]_ ;
  assign \new_[2750]_  = \new_[33230]_  & \new_[33219]_ ;
  assign \new_[2751]_  = \new_[33208]_  & \new_[33197]_ ;
  assign \new_[2752]_  = \new_[33186]_  & \new_[33175]_ ;
  assign \new_[2753]_  = \new_[33164]_  & \new_[33153]_ ;
  assign \new_[2754]_  = \new_[33142]_  & \new_[33131]_ ;
  assign \new_[2755]_  = \new_[33120]_  & \new_[33109]_ ;
  assign \new_[2756]_  = \new_[33098]_  & \new_[33087]_ ;
  assign \new_[2757]_  = \new_[33076]_  & \new_[33065]_ ;
  assign \new_[2758]_  = \new_[33054]_  & \new_[33043]_ ;
  assign \new_[2759]_  = \new_[33032]_  & \new_[33021]_ ;
  assign \new_[2760]_  = \new_[33010]_  & \new_[32999]_ ;
  assign \new_[2761]_  = \new_[32988]_  & \new_[32977]_ ;
  assign \new_[2762]_  = \new_[32966]_  & \new_[32955]_ ;
  assign \new_[2763]_  = \new_[32944]_  & \new_[32933]_ ;
  assign \new_[2764]_  = \new_[32922]_  & \new_[32911]_ ;
  assign \new_[2765]_  = \new_[32900]_  & \new_[32889]_ ;
  assign \new_[2766]_  = \new_[32878]_  & \new_[32867]_ ;
  assign \new_[2767]_  = \new_[32856]_  & \new_[32845]_ ;
  assign \new_[2768]_  = \new_[32834]_  & \new_[32823]_ ;
  assign \new_[2769]_  = \new_[32812]_  & \new_[32801]_ ;
  assign \new_[2770]_  = \new_[32790]_  & \new_[32779]_ ;
  assign \new_[2771]_  = \new_[32768]_  & \new_[32757]_ ;
  assign \new_[2772]_  = \new_[32746]_  & \new_[32735]_ ;
  assign \new_[2773]_  = \new_[32724]_  & \new_[32713]_ ;
  assign \new_[2774]_  = \new_[32702]_  & \new_[32691]_ ;
  assign \new_[2775]_  = \new_[32680]_  & \new_[32669]_ ;
  assign \new_[2776]_  = \new_[32658]_  & \new_[32647]_ ;
  assign \new_[2777]_  = \new_[32636]_  & \new_[32625]_ ;
  assign \new_[2778]_  = \new_[32614]_  & \new_[32603]_ ;
  assign \new_[2779]_  = \new_[32592]_  & \new_[32581]_ ;
  assign \new_[2780]_  = \new_[32570]_  & \new_[32559]_ ;
  assign \new_[2781]_  = \new_[32548]_  & \new_[32537]_ ;
  assign \new_[2782]_  = \new_[32526]_  & \new_[32515]_ ;
  assign \new_[2783]_  = \new_[32504]_  & \new_[32493]_ ;
  assign \new_[2784]_  = \new_[32482]_  & \new_[32471]_ ;
  assign \new_[2785]_  = \new_[32460]_  & \new_[32449]_ ;
  assign \new_[2786]_  = \new_[32438]_  & \new_[32427]_ ;
  assign \new_[2787]_  = \new_[32416]_  & \new_[32405]_ ;
  assign \new_[2788]_  = \new_[32394]_  & \new_[32383]_ ;
  assign \new_[2789]_  = \new_[32372]_  & \new_[32361]_ ;
  assign \new_[2790]_  = \new_[32350]_  & \new_[32339]_ ;
  assign \new_[2791]_  = \new_[32328]_  & \new_[32317]_ ;
  assign \new_[2792]_  = \new_[32306]_  & \new_[32295]_ ;
  assign \new_[2793]_  = \new_[32284]_  & \new_[32273]_ ;
  assign \new_[2794]_  = \new_[32262]_  & \new_[32251]_ ;
  assign \new_[2795]_  = \new_[32240]_  & \new_[32229]_ ;
  assign \new_[2796]_  = \new_[32218]_  & \new_[32207]_ ;
  assign \new_[2797]_  = \new_[32196]_  & \new_[32185]_ ;
  assign \new_[2798]_  = \new_[32174]_  & \new_[32163]_ ;
  assign \new_[2799]_  = \new_[32152]_  & \new_[32141]_ ;
  assign \new_[2800]_  = \new_[32130]_  & \new_[32119]_ ;
  assign \new_[2801]_  = \new_[32108]_  & \new_[32097]_ ;
  assign \new_[2802]_  = \new_[32086]_  & \new_[32075]_ ;
  assign \new_[2803]_  = \new_[32064]_  & \new_[32053]_ ;
  assign \new_[2804]_  = \new_[32042]_  & \new_[32031]_ ;
  assign \new_[2805]_  = \new_[32020]_  & \new_[32009]_ ;
  assign \new_[2806]_  = \new_[31998]_  & \new_[31987]_ ;
  assign \new_[2807]_  = \new_[31976]_  & \new_[31965]_ ;
  assign \new_[2808]_  = \new_[31954]_  & \new_[31943]_ ;
  assign \new_[2809]_  = \new_[31932]_  & \new_[31921]_ ;
  assign \new_[2810]_  = \new_[31910]_  & \new_[31899]_ ;
  assign \new_[2811]_  = \new_[31888]_  & \new_[31877]_ ;
  assign \new_[2812]_  = \new_[31866]_  & \new_[31855]_ ;
  assign \new_[2813]_  = \new_[31844]_  & \new_[31833]_ ;
  assign \new_[2814]_  = \new_[31822]_  & \new_[31811]_ ;
  assign \new_[2815]_  = \new_[31800]_  & \new_[31789]_ ;
  assign \new_[2816]_  = \new_[31778]_  & \new_[31767]_ ;
  assign \new_[2817]_  = \new_[31756]_  & \new_[31745]_ ;
  assign \new_[2818]_  = \new_[31734]_  & \new_[31723]_ ;
  assign \new_[2819]_  = \new_[31712]_  & \new_[31701]_ ;
  assign \new_[2820]_  = \new_[31690]_  & \new_[31679]_ ;
  assign \new_[2821]_  = \new_[31668]_  & \new_[31657]_ ;
  assign \new_[2822]_  = \new_[31646]_  & \new_[31635]_ ;
  assign \new_[2823]_  = \new_[31624]_  & \new_[31613]_ ;
  assign \new_[2824]_  = \new_[31602]_  & \new_[31591]_ ;
  assign \new_[2825]_  = \new_[31580]_  & \new_[31569]_ ;
  assign \new_[2826]_  = \new_[31558]_  & \new_[31547]_ ;
  assign \new_[2827]_  = \new_[31536]_  & \new_[31525]_ ;
  assign \new_[2828]_  = \new_[31514]_  & \new_[31503]_ ;
  assign \new_[2829]_  = \new_[31492]_  & \new_[31481]_ ;
  assign \new_[2830]_  = \new_[31470]_  & \new_[31459]_ ;
  assign \new_[2831]_  = \new_[31448]_  & \new_[31437]_ ;
  assign \new_[2832]_  = \new_[31426]_  & \new_[31415]_ ;
  assign \new_[2833]_  = \new_[31404]_  & \new_[31393]_ ;
  assign \new_[2834]_  = \new_[31382]_  & \new_[31371]_ ;
  assign \new_[2835]_  = \new_[31360]_  & \new_[31349]_ ;
  assign \new_[2836]_  = \new_[31338]_  & \new_[31327]_ ;
  assign \new_[2837]_  = \new_[31316]_  & \new_[31305]_ ;
  assign \new_[2838]_  = \new_[31294]_  & \new_[31283]_ ;
  assign \new_[2839]_  = \new_[31272]_  & \new_[31261]_ ;
  assign \new_[2840]_  = \new_[31250]_  & \new_[31239]_ ;
  assign \new_[2841]_  = \new_[31228]_  & \new_[31217]_ ;
  assign \new_[2842]_  = \new_[31206]_  & \new_[31195]_ ;
  assign \new_[2843]_  = \new_[31184]_  & \new_[31173]_ ;
  assign \new_[2844]_  = \new_[31162]_  & \new_[31151]_ ;
  assign \new_[2845]_  = \new_[31140]_  & \new_[31129]_ ;
  assign \new_[2846]_  = \new_[31118]_  & \new_[31107]_ ;
  assign \new_[2847]_  = \new_[31096]_  & \new_[31085]_ ;
  assign \new_[2848]_  = \new_[31074]_  & \new_[31063]_ ;
  assign \new_[2849]_  = \new_[31052]_  & \new_[31041]_ ;
  assign \new_[2850]_  = \new_[31030]_  & \new_[31019]_ ;
  assign \new_[2851]_  = \new_[31008]_  & \new_[30997]_ ;
  assign \new_[2852]_  = \new_[30986]_  & \new_[30975]_ ;
  assign \new_[2853]_  = \new_[30964]_  & \new_[30953]_ ;
  assign \new_[2854]_  = \new_[30942]_  & \new_[30931]_ ;
  assign \new_[2855]_  = \new_[30920]_  & \new_[30909]_ ;
  assign \new_[2856]_  = \new_[30898]_  & \new_[30887]_ ;
  assign \new_[2857]_  = \new_[30876]_  & \new_[30865]_ ;
  assign \new_[2858]_  = \new_[30854]_  & \new_[30843]_ ;
  assign \new_[2859]_  = \new_[30832]_  & \new_[30821]_ ;
  assign \new_[2860]_  = \new_[30810]_  & \new_[30799]_ ;
  assign \new_[2861]_  = \new_[30788]_  & \new_[30777]_ ;
  assign \new_[2862]_  = \new_[30766]_  & \new_[30755]_ ;
  assign \new_[2863]_  = \new_[30744]_  & \new_[30733]_ ;
  assign \new_[2864]_  = \new_[30722]_  & \new_[30711]_ ;
  assign \new_[2865]_  = \new_[30700]_  & \new_[30689]_ ;
  assign \new_[2866]_  = \new_[30678]_  & \new_[30667]_ ;
  assign \new_[2867]_  = \new_[30656]_  & \new_[30645]_ ;
  assign \new_[2868]_  = \new_[30634]_  & \new_[30623]_ ;
  assign \new_[2869]_  = \new_[30612]_  & \new_[30601]_ ;
  assign \new_[2870]_  = \new_[30590]_  & \new_[30579]_ ;
  assign \new_[2871]_  = \new_[30568]_  & \new_[30557]_ ;
  assign \new_[2872]_  = \new_[30546]_  & \new_[30535]_ ;
  assign \new_[2873]_  = \new_[30524]_  & \new_[30513]_ ;
  assign \new_[2874]_  = \new_[30502]_  & \new_[30491]_ ;
  assign \new_[2875]_  = \new_[30480]_  & \new_[30469]_ ;
  assign \new_[2876]_  = \new_[30458]_  & \new_[30447]_ ;
  assign \new_[2877]_  = \new_[30436]_  & \new_[30425]_ ;
  assign \new_[2878]_  = \new_[30414]_  & \new_[30403]_ ;
  assign \new_[2879]_  = \new_[30392]_  & \new_[30381]_ ;
  assign \new_[2880]_  = \new_[30370]_  & \new_[30359]_ ;
  assign \new_[2881]_  = \new_[30348]_  & \new_[30337]_ ;
  assign \new_[2882]_  = \new_[30326]_  & \new_[30315]_ ;
  assign \new_[2883]_  = \new_[30304]_  & \new_[30293]_ ;
  assign \new_[2884]_  = \new_[30282]_  & \new_[30271]_ ;
  assign \new_[2885]_  = \new_[30260]_  & \new_[30249]_ ;
  assign \new_[2886]_  = \new_[30238]_  & \new_[30227]_ ;
  assign \new_[2887]_  = \new_[30216]_  & \new_[30205]_ ;
  assign \new_[2888]_  = \new_[30194]_  & \new_[30183]_ ;
  assign \new_[2889]_  = \new_[30172]_  & \new_[30161]_ ;
  assign \new_[2890]_  = \new_[30150]_  & \new_[30139]_ ;
  assign \new_[2891]_  = \new_[30128]_  & \new_[30117]_ ;
  assign \new_[2892]_  = \new_[30106]_  & \new_[30095]_ ;
  assign \new_[2893]_  = \new_[30084]_  & \new_[30073]_ ;
  assign \new_[2894]_  = \new_[30062]_  & \new_[30051]_ ;
  assign \new_[2895]_  = \new_[30040]_  & \new_[30029]_ ;
  assign \new_[2896]_  = \new_[30018]_  & \new_[30007]_ ;
  assign \new_[2897]_  = \new_[29996]_  & \new_[29985]_ ;
  assign \new_[2898]_  = \new_[29974]_  & \new_[29963]_ ;
  assign \new_[2899]_  = \new_[29952]_  & \new_[29941]_ ;
  assign \new_[2900]_  = \new_[29930]_  & \new_[29919]_ ;
  assign \new_[2901]_  = \new_[29908]_  & \new_[29897]_ ;
  assign \new_[2902]_  = \new_[29886]_  & \new_[29875]_ ;
  assign \new_[2903]_  = \new_[29864]_  & \new_[29853]_ ;
  assign \new_[2904]_  = \new_[29842]_  & \new_[29831]_ ;
  assign \new_[2905]_  = \new_[29820]_  & \new_[29809]_ ;
  assign \new_[2906]_  = \new_[29798]_  & \new_[29787]_ ;
  assign \new_[2907]_  = \new_[29776]_  & \new_[29765]_ ;
  assign \new_[2908]_  = \new_[29754]_  & \new_[29743]_ ;
  assign \new_[2909]_  = \new_[29732]_  & \new_[29721]_ ;
  assign \new_[2910]_  = \new_[29710]_  & \new_[29699]_ ;
  assign \new_[2911]_  = \new_[29688]_  & \new_[29677]_ ;
  assign \new_[2912]_  = \new_[29666]_  & \new_[29655]_ ;
  assign \new_[2913]_  = \new_[29644]_  & \new_[29633]_ ;
  assign \new_[2914]_  = \new_[29622]_  & \new_[29611]_ ;
  assign \new_[2915]_  = \new_[29600]_  & \new_[29589]_ ;
  assign \new_[2916]_  = \new_[29578]_  & \new_[29567]_ ;
  assign \new_[2917]_  = \new_[29556]_  & \new_[29545]_ ;
  assign \new_[2918]_  = \new_[29534]_  & \new_[29523]_ ;
  assign \new_[2919]_  = \new_[29512]_  & \new_[29501]_ ;
  assign \new_[2920]_  = \new_[29490]_  & \new_[29479]_ ;
  assign \new_[2921]_  = \new_[29468]_  & \new_[29457]_ ;
  assign \new_[2922]_  = \new_[29446]_  & \new_[29435]_ ;
  assign \new_[2923]_  = \new_[29424]_  & \new_[29413]_ ;
  assign \new_[2924]_  = \new_[29402]_  & \new_[29391]_ ;
  assign \new_[2925]_  = \new_[29380]_  & \new_[29369]_ ;
  assign \new_[2926]_  = \new_[29358]_  & \new_[29347]_ ;
  assign \new_[2927]_  = \new_[29336]_  & \new_[29325]_ ;
  assign \new_[2928]_  = \new_[29314]_  & \new_[29303]_ ;
  assign \new_[2929]_  = \new_[29292]_  & \new_[29281]_ ;
  assign \new_[2930]_  = \new_[29270]_  & \new_[29259]_ ;
  assign \new_[2931]_  = \new_[29248]_  & \new_[29237]_ ;
  assign \new_[2932]_  = \new_[29226]_  & \new_[29215]_ ;
  assign \new_[2933]_  = \new_[29204]_  & \new_[29193]_ ;
  assign \new_[2934]_  = \new_[29182]_  & \new_[29171]_ ;
  assign \new_[2935]_  = \new_[29160]_  & \new_[29149]_ ;
  assign \new_[2936]_  = \new_[29138]_  & \new_[29127]_ ;
  assign \new_[2937]_  = \new_[29116]_  & \new_[29105]_ ;
  assign \new_[2938]_  = \new_[29094]_  & \new_[29083]_ ;
  assign \new_[2939]_  = \new_[29072]_  & \new_[29061]_ ;
  assign \new_[2940]_  = \new_[29050]_  & \new_[29039]_ ;
  assign \new_[2941]_  = \new_[29028]_  & \new_[29017]_ ;
  assign \new_[2942]_  = \new_[29006]_  & \new_[28995]_ ;
  assign \new_[2943]_  = \new_[28984]_  & \new_[28973]_ ;
  assign \new_[2944]_  = \new_[28962]_  & \new_[28951]_ ;
  assign \new_[2945]_  = \new_[28940]_  & \new_[28929]_ ;
  assign \new_[2946]_  = \new_[28918]_  & \new_[28907]_ ;
  assign \new_[2947]_  = \new_[28896]_  & \new_[28885]_ ;
  assign \new_[2948]_  = \new_[28874]_  & \new_[28863]_ ;
  assign \new_[2949]_  = \new_[28852]_  & \new_[28841]_ ;
  assign \new_[2950]_  = \new_[28830]_  & \new_[28819]_ ;
  assign \new_[2951]_  = \new_[28808]_  & \new_[28797]_ ;
  assign \new_[2952]_  = \new_[28786]_  & \new_[28775]_ ;
  assign \new_[2953]_  = \new_[28764]_  & \new_[28753]_ ;
  assign \new_[2954]_  = \new_[28742]_  & \new_[28731]_ ;
  assign \new_[2955]_  = \new_[28720]_  & \new_[28709]_ ;
  assign \new_[2956]_  = \new_[28698]_  & \new_[28687]_ ;
  assign \new_[2957]_  = \new_[28676]_  & \new_[28665]_ ;
  assign \new_[2958]_  = \new_[28654]_  & \new_[28643]_ ;
  assign \new_[2959]_  = \new_[28632]_  & \new_[28621]_ ;
  assign \new_[2960]_  = \new_[28610]_  & \new_[28599]_ ;
  assign \new_[2961]_  = \new_[28588]_  & \new_[28577]_ ;
  assign \new_[2962]_  = \new_[28566]_  & \new_[28555]_ ;
  assign \new_[2963]_  = \new_[28544]_  & \new_[28533]_ ;
  assign \new_[2964]_  = \new_[28522]_  & \new_[28511]_ ;
  assign \new_[2965]_  = \new_[28500]_  & \new_[28489]_ ;
  assign \new_[2966]_  = \new_[28478]_  & \new_[28467]_ ;
  assign \new_[2967]_  = \new_[28456]_  & \new_[28445]_ ;
  assign \new_[2968]_  = \new_[28434]_  & \new_[28423]_ ;
  assign \new_[2969]_  = \new_[28412]_  & \new_[28401]_ ;
  assign \new_[2970]_  = \new_[28390]_  & \new_[28379]_ ;
  assign \new_[2971]_  = \new_[28368]_  & \new_[28357]_ ;
  assign \new_[2972]_  = \new_[28346]_  & \new_[28335]_ ;
  assign \new_[2973]_  = \new_[28324]_  & \new_[28313]_ ;
  assign \new_[2974]_  = \new_[28302]_  & \new_[28291]_ ;
  assign \new_[2975]_  = \new_[28280]_  & \new_[28269]_ ;
  assign \new_[2976]_  = \new_[28258]_  & \new_[28247]_ ;
  assign \new_[2977]_  = \new_[28236]_  & \new_[28225]_ ;
  assign \new_[2978]_  = \new_[28214]_  & \new_[28203]_ ;
  assign \new_[2979]_  = \new_[28192]_  & \new_[28181]_ ;
  assign \new_[2980]_  = \new_[28170]_  & \new_[28159]_ ;
  assign \new_[2981]_  = \new_[28148]_  & \new_[28137]_ ;
  assign \new_[2982]_  = \new_[28126]_  & \new_[28115]_ ;
  assign \new_[2983]_  = \new_[28104]_  & \new_[28093]_ ;
  assign \new_[2984]_  = \new_[28082]_  & \new_[28071]_ ;
  assign \new_[2985]_  = \new_[28060]_  & \new_[28049]_ ;
  assign \new_[2986]_  = \new_[28038]_  & \new_[28027]_ ;
  assign \new_[2987]_  = \new_[28016]_  & \new_[28005]_ ;
  assign \new_[2988]_  = \new_[27994]_  & \new_[27983]_ ;
  assign \new_[2989]_  = \new_[27972]_  & \new_[27961]_ ;
  assign \new_[2990]_  = \new_[27950]_  & \new_[27939]_ ;
  assign \new_[2991]_  = \new_[27928]_  & \new_[27917]_ ;
  assign \new_[2992]_  = \new_[27906]_  & \new_[27895]_ ;
  assign \new_[2993]_  = \new_[27884]_  & \new_[27873]_ ;
  assign \new_[2994]_  = \new_[27862]_  & \new_[27851]_ ;
  assign \new_[2995]_  = \new_[27840]_  & \new_[27829]_ ;
  assign \new_[2996]_  = \new_[27818]_  & \new_[27807]_ ;
  assign \new_[2997]_  = \new_[27796]_  & \new_[27785]_ ;
  assign \new_[2998]_  = \new_[27774]_  & \new_[27763]_ ;
  assign \new_[2999]_  = \new_[27752]_  & \new_[27741]_ ;
  assign \new_[3000]_  = \new_[27730]_  & \new_[27719]_ ;
  assign \new_[3001]_  = \new_[27708]_  & \new_[27697]_ ;
  assign \new_[3002]_  = \new_[27686]_  & \new_[27675]_ ;
  assign \new_[3003]_  = \new_[27664]_  & \new_[27653]_ ;
  assign \new_[3004]_  = \new_[27642]_  & \new_[27631]_ ;
  assign \new_[3005]_  = \new_[27620]_  & \new_[27609]_ ;
  assign \new_[3006]_  = \new_[27598]_  & \new_[27587]_ ;
  assign \new_[3007]_  = \new_[27576]_  & \new_[27565]_ ;
  assign \new_[3008]_  = \new_[27554]_  & \new_[27543]_ ;
  assign \new_[3009]_  = \new_[27532]_  & \new_[27521]_ ;
  assign \new_[3010]_  = \new_[27510]_  & \new_[27499]_ ;
  assign \new_[3011]_  = \new_[27488]_  & \new_[27477]_ ;
  assign \new_[3012]_  = \new_[27466]_  & \new_[27455]_ ;
  assign \new_[3013]_  = \new_[27444]_  & \new_[27433]_ ;
  assign \new_[3014]_  = \new_[27422]_  & \new_[27411]_ ;
  assign \new_[3015]_  = \new_[27400]_  & \new_[27389]_ ;
  assign \new_[3016]_  = \new_[27378]_  & \new_[27367]_ ;
  assign \new_[3017]_  = \new_[27356]_  & \new_[27345]_ ;
  assign \new_[3018]_  = \new_[27334]_  & \new_[27323]_ ;
  assign \new_[3019]_  = \new_[27312]_  & \new_[27301]_ ;
  assign \new_[3020]_  = \new_[27290]_  & \new_[27279]_ ;
  assign \new_[3021]_  = \new_[27268]_  & \new_[27257]_ ;
  assign \new_[3022]_  = \new_[27246]_  & \new_[27235]_ ;
  assign \new_[3023]_  = \new_[27224]_  & \new_[27213]_ ;
  assign \new_[3024]_  = \new_[27202]_  & \new_[27191]_ ;
  assign \new_[3025]_  = \new_[27180]_  & \new_[27169]_ ;
  assign \new_[3026]_  = \new_[27158]_  & \new_[27147]_ ;
  assign \new_[3027]_  = \new_[27136]_  & \new_[27125]_ ;
  assign \new_[3028]_  = \new_[27114]_  & \new_[27103]_ ;
  assign \new_[3029]_  = \new_[27092]_  & \new_[27081]_ ;
  assign \new_[3030]_  = \new_[27070]_  & \new_[27059]_ ;
  assign \new_[3031]_  = \new_[27048]_  & \new_[27037]_ ;
  assign \new_[3032]_  = \new_[27026]_  & \new_[27015]_ ;
  assign \new_[3033]_  = \new_[27004]_  & \new_[26993]_ ;
  assign \new_[3034]_  = \new_[26982]_  & \new_[26971]_ ;
  assign \new_[3035]_  = \new_[26960]_  & \new_[26949]_ ;
  assign \new_[3036]_  = \new_[26938]_  & \new_[26927]_ ;
  assign \new_[3037]_  = \new_[26916]_  & \new_[26905]_ ;
  assign \new_[3038]_  = \new_[26894]_  & \new_[26883]_ ;
  assign \new_[3039]_  = \new_[26872]_  & \new_[26861]_ ;
  assign \new_[3040]_  = \new_[26850]_  & \new_[26839]_ ;
  assign \new_[3041]_  = \new_[26828]_  & \new_[26817]_ ;
  assign \new_[3042]_  = \new_[26806]_  & \new_[26795]_ ;
  assign \new_[3043]_  = \new_[26784]_  & \new_[26773]_ ;
  assign \new_[3044]_  = \new_[26762]_  & \new_[26751]_ ;
  assign \new_[3045]_  = \new_[26740]_  & \new_[26729]_ ;
  assign \new_[3046]_  = \new_[26718]_  & \new_[26707]_ ;
  assign \new_[3047]_  = \new_[26696]_  & \new_[26685]_ ;
  assign \new_[3048]_  = \new_[26674]_  & \new_[26663]_ ;
  assign \new_[3049]_  = \new_[26652]_  & \new_[26641]_ ;
  assign \new_[3050]_  = \new_[26630]_  & \new_[26619]_ ;
  assign \new_[3051]_  = \new_[26608]_  & \new_[26597]_ ;
  assign \new_[3052]_  = \new_[26586]_  & \new_[26575]_ ;
  assign \new_[3053]_  = \new_[26564]_  & \new_[26553]_ ;
  assign \new_[3054]_  = \new_[26542]_  & \new_[26531]_ ;
  assign \new_[3055]_  = \new_[26520]_  & \new_[26509]_ ;
  assign \new_[3056]_  = \new_[26498]_  & \new_[26487]_ ;
  assign \new_[3057]_  = \new_[26476]_  & \new_[26465]_ ;
  assign \new_[3058]_  = \new_[26454]_  & \new_[26443]_ ;
  assign \new_[3059]_  = \new_[26432]_  & \new_[26421]_ ;
  assign \new_[3060]_  = \new_[26410]_  & \new_[26399]_ ;
  assign \new_[3061]_  = \new_[26388]_  & \new_[26377]_ ;
  assign \new_[3062]_  = \new_[26366]_  & \new_[26355]_ ;
  assign \new_[3063]_  = \new_[26344]_  & \new_[26333]_ ;
  assign \new_[3064]_  = \new_[26322]_  & \new_[26311]_ ;
  assign \new_[3065]_  = \new_[26300]_  & \new_[26289]_ ;
  assign \new_[3066]_  = \new_[26278]_  & \new_[26267]_ ;
  assign \new_[3067]_  = \new_[26256]_  & \new_[26245]_ ;
  assign \new_[3068]_  = \new_[26234]_  & \new_[26223]_ ;
  assign \new_[3069]_  = \new_[26212]_  & \new_[26201]_ ;
  assign \new_[3070]_  = \new_[26190]_  & \new_[26179]_ ;
  assign \new_[3071]_  = \new_[26168]_  & \new_[26157]_ ;
  assign \new_[3072]_  = \new_[26146]_  & \new_[26135]_ ;
  assign \new_[3073]_  = \new_[26124]_  & \new_[26113]_ ;
  assign \new_[3074]_  = \new_[26102]_  & \new_[26091]_ ;
  assign \new_[3075]_  = \new_[26080]_  & \new_[26069]_ ;
  assign \new_[3076]_  = \new_[26058]_  & \new_[26047]_ ;
  assign \new_[3077]_  = \new_[26036]_  & \new_[26025]_ ;
  assign \new_[3078]_  = \new_[26014]_  & \new_[26003]_ ;
  assign \new_[3079]_  = \new_[25992]_  & \new_[25981]_ ;
  assign \new_[3080]_  = \new_[25970]_  & \new_[25959]_ ;
  assign \new_[3081]_  = \new_[25948]_  & \new_[25937]_ ;
  assign \new_[3082]_  = \new_[25926]_  & \new_[25915]_ ;
  assign \new_[3083]_  = \new_[25904]_  & \new_[25893]_ ;
  assign \new_[3084]_  = \new_[25882]_  & \new_[25871]_ ;
  assign \new_[3085]_  = \new_[25860]_  & \new_[25849]_ ;
  assign \new_[3086]_  = \new_[25838]_  & \new_[25827]_ ;
  assign \new_[3087]_  = \new_[25816]_  & \new_[25805]_ ;
  assign \new_[3088]_  = \new_[25794]_  & \new_[25783]_ ;
  assign \new_[3089]_  = \new_[25772]_  & \new_[25761]_ ;
  assign \new_[3090]_  = \new_[25750]_  & \new_[25739]_ ;
  assign \new_[3091]_  = \new_[25728]_  & \new_[25717]_ ;
  assign \new_[3092]_  = \new_[25706]_  & \new_[25695]_ ;
  assign \new_[3093]_  = \new_[25684]_  & \new_[25673]_ ;
  assign \new_[3094]_  = \new_[25662]_  & \new_[25651]_ ;
  assign \new_[3095]_  = \new_[25640]_  & \new_[25629]_ ;
  assign \new_[3096]_  = \new_[25618]_  & \new_[25607]_ ;
  assign \new_[3097]_  = \new_[25596]_  & \new_[25585]_ ;
  assign \new_[3098]_  = \new_[25574]_  & \new_[25563]_ ;
  assign \new_[3099]_  = \new_[25552]_  & \new_[25541]_ ;
  assign \new_[3100]_  = \new_[25530]_  & \new_[25519]_ ;
  assign \new_[3101]_  = \new_[25508]_  & \new_[25497]_ ;
  assign \new_[3102]_  = \new_[25486]_  & \new_[25475]_ ;
  assign \new_[3103]_  = \new_[25464]_  & \new_[25453]_ ;
  assign \new_[3104]_  = \new_[25442]_  & \new_[25431]_ ;
  assign \new_[3105]_  = \new_[25420]_  & \new_[25409]_ ;
  assign \new_[3106]_  = \new_[25398]_  & \new_[25387]_ ;
  assign \new_[3107]_  = \new_[25376]_  & \new_[25365]_ ;
  assign \new_[3108]_  = \new_[25354]_  & \new_[25343]_ ;
  assign \new_[3109]_  = \new_[25332]_  & \new_[25321]_ ;
  assign \new_[3110]_  = \new_[25310]_  & \new_[25299]_ ;
  assign \new_[3111]_  = \new_[25288]_  & \new_[25277]_ ;
  assign \new_[3112]_  = \new_[25266]_  & \new_[25255]_ ;
  assign \new_[3113]_  = \new_[25244]_  & \new_[25233]_ ;
  assign \new_[3114]_  = \new_[25222]_  & \new_[25211]_ ;
  assign \new_[3115]_  = \new_[25200]_  & \new_[25189]_ ;
  assign \new_[3116]_  = \new_[25178]_  & \new_[25167]_ ;
  assign \new_[3117]_  = \new_[25156]_  & \new_[25145]_ ;
  assign \new_[3118]_  = \new_[25134]_  & \new_[25123]_ ;
  assign \new_[3119]_  = \new_[25112]_  & \new_[25101]_ ;
  assign \new_[3120]_  = \new_[25090]_  & \new_[25079]_ ;
  assign \new_[3121]_  = \new_[25068]_  & \new_[25057]_ ;
  assign \new_[3122]_  = \new_[25046]_  & \new_[25035]_ ;
  assign \new_[3123]_  = \new_[25024]_  & \new_[25013]_ ;
  assign \new_[3124]_  = \new_[25002]_  & \new_[24991]_ ;
  assign \new_[3125]_  = \new_[24980]_  & \new_[24969]_ ;
  assign \new_[3126]_  = \new_[24958]_  & \new_[24947]_ ;
  assign \new_[3127]_  = \new_[24936]_  & \new_[24925]_ ;
  assign \new_[3128]_  = \new_[24914]_  & \new_[24903]_ ;
  assign \new_[3129]_  = \new_[24892]_  & \new_[24881]_ ;
  assign \new_[3130]_  = \new_[24870]_  & \new_[24859]_ ;
  assign \new_[3131]_  = \new_[24848]_  & \new_[24837]_ ;
  assign \new_[3132]_  = \new_[24826]_  & \new_[24815]_ ;
  assign \new_[3133]_  = \new_[24804]_  & \new_[24793]_ ;
  assign \new_[3134]_  = \new_[24782]_  & \new_[24771]_ ;
  assign \new_[3135]_  = \new_[24760]_  & \new_[24749]_ ;
  assign \new_[3136]_  = \new_[24738]_  & \new_[24727]_ ;
  assign \new_[3137]_  = \new_[24716]_  & \new_[24705]_ ;
  assign \new_[3138]_  = \new_[24694]_  & \new_[24683]_ ;
  assign \new_[3139]_  = \new_[24672]_  & \new_[24661]_ ;
  assign \new_[3140]_  = \new_[24650]_  & \new_[24639]_ ;
  assign \new_[3141]_  = \new_[24628]_  & \new_[24617]_ ;
  assign \new_[3142]_  = \new_[24606]_  & \new_[24595]_ ;
  assign \new_[3143]_  = \new_[24584]_  & \new_[24573]_ ;
  assign \new_[3144]_  = \new_[24562]_  & \new_[24551]_ ;
  assign \new_[3145]_  = \new_[24540]_  & \new_[24529]_ ;
  assign \new_[3146]_  = \new_[24518]_  & \new_[24507]_ ;
  assign \new_[3147]_  = \new_[24496]_  & \new_[24485]_ ;
  assign \new_[3148]_  = \new_[24476]_  & \new_[24465]_ ;
  assign \new_[3149]_  = \new_[24456]_  & \new_[24445]_ ;
  assign \new_[3150]_  = \new_[24436]_  & \new_[24425]_ ;
  assign \new_[3151]_  = \new_[24416]_  & \new_[24405]_ ;
  assign \new_[3152]_  = \new_[24396]_  & \new_[24385]_ ;
  assign \new_[3153]_  = \new_[24376]_  & \new_[24365]_ ;
  assign \new_[3154]_  = \new_[24356]_  & \new_[24345]_ ;
  assign \new_[3155]_  = \new_[24336]_  & \new_[24325]_ ;
  assign \new_[3156]_  = \new_[24316]_  & \new_[24305]_ ;
  assign \new_[3157]_  = \new_[24296]_  & \new_[24285]_ ;
  assign \new_[3158]_  = \new_[24276]_  & \new_[24265]_ ;
  assign \new_[3159]_  = \new_[24256]_  & \new_[24245]_ ;
  assign \new_[3160]_  = \new_[24236]_  & \new_[24225]_ ;
  assign \new_[3161]_  = \new_[24216]_  & \new_[24205]_ ;
  assign \new_[3162]_  = \new_[24196]_  & \new_[24185]_ ;
  assign \new_[3163]_  = \new_[24176]_  & \new_[24165]_ ;
  assign \new_[3164]_  = \new_[24156]_  & \new_[24145]_ ;
  assign \new_[3165]_  = \new_[24136]_  & \new_[24125]_ ;
  assign \new_[3166]_  = \new_[24116]_  & \new_[24105]_ ;
  assign \new_[3167]_  = \new_[24096]_  & \new_[24085]_ ;
  assign \new_[3168]_  = \new_[24076]_  & \new_[24065]_ ;
  assign \new_[3169]_  = \new_[24056]_  & \new_[24045]_ ;
  assign \new_[3170]_  = \new_[24036]_  & \new_[24025]_ ;
  assign \new_[3171]_  = \new_[24016]_  & \new_[24005]_ ;
  assign \new_[3172]_  = \new_[23996]_  & \new_[23985]_ ;
  assign \new_[3173]_  = \new_[23976]_  & \new_[23965]_ ;
  assign \new_[3174]_  = \new_[23956]_  & \new_[23945]_ ;
  assign \new_[3175]_  = \new_[23936]_  & \new_[23925]_ ;
  assign \new_[3176]_  = \new_[23916]_  & \new_[23905]_ ;
  assign \new_[3177]_  = \new_[23896]_  & \new_[23885]_ ;
  assign \new_[3178]_  = \new_[23876]_  & \new_[23865]_ ;
  assign \new_[3179]_  = \new_[23856]_  & \new_[23845]_ ;
  assign \new_[3180]_  = \new_[23836]_  & \new_[23825]_ ;
  assign \new_[3181]_  = \new_[23816]_  & \new_[23805]_ ;
  assign \new_[3182]_  = \new_[23796]_  & \new_[23785]_ ;
  assign \new_[3183]_  = \new_[23776]_  & \new_[23765]_ ;
  assign \new_[3184]_  = \new_[23756]_  & \new_[23745]_ ;
  assign \new_[3185]_  = \new_[23736]_  & \new_[23725]_ ;
  assign \new_[3186]_  = \new_[23716]_  & \new_[23705]_ ;
  assign \new_[3187]_  = \new_[23696]_  & \new_[23685]_ ;
  assign \new_[3188]_  = \new_[23676]_  & \new_[23665]_ ;
  assign \new_[3189]_  = \new_[23656]_  & \new_[23645]_ ;
  assign \new_[3190]_  = \new_[23636]_  & \new_[23625]_ ;
  assign \new_[3191]_  = \new_[23616]_  & \new_[23605]_ ;
  assign \new_[3192]_  = \new_[23596]_  & \new_[23585]_ ;
  assign \new_[3193]_  = \new_[23576]_  & \new_[23565]_ ;
  assign \new_[3194]_  = \new_[23556]_  & \new_[23545]_ ;
  assign \new_[3195]_  = \new_[23536]_  & \new_[23525]_ ;
  assign \new_[3196]_  = \new_[23516]_  & \new_[23505]_ ;
  assign \new_[3197]_  = \new_[23496]_  & \new_[23485]_ ;
  assign \new_[3198]_  = \new_[23476]_  & \new_[23465]_ ;
  assign \new_[3199]_  = \new_[23456]_  & \new_[23445]_ ;
  assign \new_[3200]_  = \new_[23436]_  & \new_[23425]_ ;
  assign \new_[3201]_  = \new_[23416]_  & \new_[23405]_ ;
  assign \new_[3202]_  = \new_[23396]_  & \new_[23385]_ ;
  assign \new_[3203]_  = \new_[23376]_  & \new_[23365]_ ;
  assign \new_[3204]_  = \new_[23356]_  & \new_[23345]_ ;
  assign \new_[3205]_  = \new_[23336]_  & \new_[23325]_ ;
  assign \new_[3206]_  = \new_[23316]_  & \new_[23305]_ ;
  assign \new_[3207]_  = \new_[23296]_  & \new_[23285]_ ;
  assign \new_[3208]_  = \new_[23276]_  & \new_[23265]_ ;
  assign \new_[3209]_  = \new_[23256]_  & \new_[23245]_ ;
  assign \new_[3210]_  = \new_[23236]_  & \new_[23225]_ ;
  assign \new_[3211]_  = \new_[23216]_  & \new_[23205]_ ;
  assign \new_[3212]_  = \new_[23196]_  & \new_[23185]_ ;
  assign \new_[3213]_  = \new_[23176]_  & \new_[23165]_ ;
  assign \new_[3214]_  = \new_[23156]_  & \new_[23145]_ ;
  assign \new_[3215]_  = \new_[23136]_  & \new_[23125]_ ;
  assign \new_[3216]_  = \new_[23116]_  & \new_[23105]_ ;
  assign \new_[3217]_  = \new_[23096]_  & \new_[23085]_ ;
  assign \new_[3218]_  = \new_[23076]_  & \new_[23065]_ ;
  assign \new_[3219]_  = \new_[23056]_  & \new_[23045]_ ;
  assign \new_[3220]_  = \new_[23036]_  & \new_[23025]_ ;
  assign \new_[3221]_  = \new_[23016]_  & \new_[23005]_ ;
  assign \new_[3222]_  = \new_[22996]_  & \new_[22985]_ ;
  assign \new_[3223]_  = \new_[22976]_  & \new_[22965]_ ;
  assign \new_[3224]_  = \new_[22956]_  & \new_[22945]_ ;
  assign \new_[3225]_  = \new_[22936]_  & \new_[22925]_ ;
  assign \new_[3226]_  = \new_[22916]_  & \new_[22905]_ ;
  assign \new_[3227]_  = \new_[22896]_  & \new_[22885]_ ;
  assign \new_[3228]_  = \new_[22876]_  & \new_[22865]_ ;
  assign \new_[3229]_  = \new_[22856]_  & \new_[22845]_ ;
  assign \new_[3230]_  = \new_[22836]_  & \new_[22825]_ ;
  assign \new_[3231]_  = \new_[22816]_  & \new_[22805]_ ;
  assign \new_[3232]_  = \new_[22796]_  & \new_[22785]_ ;
  assign \new_[3233]_  = \new_[22776]_  & \new_[22765]_ ;
  assign \new_[3234]_  = \new_[22756]_  & \new_[22745]_ ;
  assign \new_[3235]_  = \new_[22736]_  & \new_[22725]_ ;
  assign \new_[3236]_  = \new_[22716]_  & \new_[22705]_ ;
  assign \new_[3237]_  = \new_[22696]_  & \new_[22685]_ ;
  assign \new_[3238]_  = \new_[22676]_  & \new_[22665]_ ;
  assign \new_[3239]_  = \new_[22656]_  & \new_[22645]_ ;
  assign \new_[3240]_  = \new_[22636]_  & \new_[22625]_ ;
  assign \new_[3241]_  = \new_[22616]_  & \new_[22605]_ ;
  assign \new_[3242]_  = \new_[22596]_  & \new_[22585]_ ;
  assign \new_[3243]_  = \new_[22576]_  & \new_[22565]_ ;
  assign \new_[3244]_  = \new_[22556]_  & \new_[22545]_ ;
  assign \new_[3245]_  = \new_[22536]_  & \new_[22525]_ ;
  assign \new_[3246]_  = \new_[22516]_  & \new_[22505]_ ;
  assign \new_[3247]_  = \new_[22496]_  & \new_[22485]_ ;
  assign \new_[3248]_  = \new_[22476]_  & \new_[22465]_ ;
  assign \new_[3249]_  = \new_[22456]_  & \new_[22445]_ ;
  assign \new_[3250]_  = \new_[22436]_  & \new_[22425]_ ;
  assign \new_[3251]_  = \new_[22416]_  & \new_[22405]_ ;
  assign \new_[3252]_  = \new_[22396]_  & \new_[22385]_ ;
  assign \new_[3253]_  = \new_[22376]_  & \new_[22365]_ ;
  assign \new_[3254]_  = \new_[22356]_  & \new_[22345]_ ;
  assign \new_[3255]_  = \new_[22336]_  & \new_[22325]_ ;
  assign \new_[3256]_  = \new_[22316]_  & \new_[22305]_ ;
  assign \new_[3257]_  = \new_[22296]_  & \new_[22285]_ ;
  assign \new_[3258]_  = \new_[22276]_  & \new_[22265]_ ;
  assign \new_[3259]_  = \new_[22256]_  & \new_[22245]_ ;
  assign \new_[3260]_  = \new_[22236]_  & \new_[22225]_ ;
  assign \new_[3261]_  = \new_[22216]_  & \new_[22205]_ ;
  assign \new_[3262]_  = \new_[22196]_  & \new_[22185]_ ;
  assign \new_[3263]_  = \new_[22176]_  & \new_[22165]_ ;
  assign \new_[3264]_  = \new_[22156]_  & \new_[22145]_ ;
  assign \new_[3265]_  = \new_[22136]_  & \new_[22125]_ ;
  assign \new_[3266]_  = \new_[22116]_  & \new_[22105]_ ;
  assign \new_[3267]_  = \new_[22096]_  & \new_[22085]_ ;
  assign \new_[3268]_  = \new_[22076]_  & \new_[22065]_ ;
  assign \new_[3269]_  = \new_[22056]_  & \new_[22045]_ ;
  assign \new_[3270]_  = \new_[22036]_  & \new_[22025]_ ;
  assign \new_[3271]_  = \new_[22016]_  & \new_[22005]_ ;
  assign \new_[3272]_  = \new_[21996]_  & \new_[21985]_ ;
  assign \new_[3273]_  = \new_[21976]_  & \new_[21965]_ ;
  assign \new_[3274]_  = \new_[21956]_  & \new_[21945]_ ;
  assign \new_[3275]_  = \new_[21936]_  & \new_[21925]_ ;
  assign \new_[3276]_  = \new_[21916]_  & \new_[21905]_ ;
  assign \new_[3277]_  = \new_[21896]_  & \new_[21885]_ ;
  assign \new_[3278]_  = \new_[21876]_  & \new_[21865]_ ;
  assign \new_[3279]_  = \new_[21856]_  & \new_[21845]_ ;
  assign \new_[3280]_  = \new_[21836]_  & \new_[21825]_ ;
  assign \new_[3281]_  = \new_[21816]_  & \new_[21805]_ ;
  assign \new_[3282]_  = \new_[21796]_  & \new_[21785]_ ;
  assign \new_[3283]_  = \new_[21776]_  & \new_[21765]_ ;
  assign \new_[3284]_  = \new_[21756]_  & \new_[21745]_ ;
  assign \new_[3285]_  = \new_[21736]_  & \new_[21725]_ ;
  assign \new_[3286]_  = \new_[21716]_  & \new_[21705]_ ;
  assign \new_[3287]_  = \new_[21696]_  & \new_[21685]_ ;
  assign \new_[3288]_  = \new_[21676]_  & \new_[21665]_ ;
  assign \new_[3289]_  = \new_[21656]_  & \new_[21645]_ ;
  assign \new_[3290]_  = \new_[21636]_  & \new_[21625]_ ;
  assign \new_[3291]_  = \new_[21616]_  & \new_[21605]_ ;
  assign \new_[3292]_  = \new_[21596]_  & \new_[21585]_ ;
  assign \new_[3293]_  = \new_[21576]_  & \new_[21565]_ ;
  assign \new_[3294]_  = \new_[21556]_  & \new_[21545]_ ;
  assign \new_[3295]_  = \new_[21536]_  & \new_[21525]_ ;
  assign \new_[3296]_  = \new_[21516]_  & \new_[21505]_ ;
  assign \new_[3297]_  = \new_[21496]_  & \new_[21485]_ ;
  assign \new_[3298]_  = \new_[21476]_  & \new_[21465]_ ;
  assign \new_[3299]_  = \new_[21456]_  & \new_[21445]_ ;
  assign \new_[3300]_  = \new_[21436]_  & \new_[21425]_ ;
  assign \new_[3301]_  = \new_[21416]_  & \new_[21405]_ ;
  assign \new_[3302]_  = \new_[21396]_  & \new_[21385]_ ;
  assign \new_[3303]_  = \new_[21376]_  & \new_[21365]_ ;
  assign \new_[3304]_  = \new_[21356]_  & \new_[21345]_ ;
  assign \new_[3305]_  = \new_[21336]_  & \new_[21325]_ ;
  assign \new_[3306]_  = \new_[21316]_  & \new_[21305]_ ;
  assign \new_[3307]_  = \new_[21296]_  & \new_[21285]_ ;
  assign \new_[3308]_  = \new_[21276]_  & \new_[21265]_ ;
  assign \new_[3309]_  = \new_[21256]_  & \new_[21245]_ ;
  assign \new_[3310]_  = \new_[21236]_  & \new_[21225]_ ;
  assign \new_[3311]_  = \new_[21216]_  & \new_[21205]_ ;
  assign \new_[3312]_  = \new_[21196]_  & \new_[21185]_ ;
  assign \new_[3313]_  = \new_[21176]_  & \new_[21165]_ ;
  assign \new_[3314]_  = \new_[21156]_  & \new_[21145]_ ;
  assign \new_[3315]_  = \new_[21136]_  & \new_[21125]_ ;
  assign \new_[3316]_  = \new_[21116]_  & \new_[21105]_ ;
  assign \new_[3317]_  = \new_[21096]_  & \new_[21085]_ ;
  assign \new_[3318]_  = \new_[21076]_  & \new_[21065]_ ;
  assign \new_[3319]_  = \new_[21056]_  & \new_[21045]_ ;
  assign \new_[3320]_  = \new_[21036]_  & \new_[21025]_ ;
  assign \new_[3321]_  = \new_[21016]_  & \new_[21005]_ ;
  assign \new_[3322]_  = \new_[20996]_  & \new_[20985]_ ;
  assign \new_[3323]_  = \new_[20976]_  & \new_[20965]_ ;
  assign \new_[3324]_  = \new_[20956]_  & \new_[20945]_ ;
  assign \new_[3325]_  = \new_[20936]_  & \new_[20925]_ ;
  assign \new_[3326]_  = \new_[20916]_  & \new_[20905]_ ;
  assign \new_[3327]_  = \new_[20896]_  & \new_[20885]_ ;
  assign \new_[3328]_  = \new_[20876]_  & \new_[20865]_ ;
  assign \new_[3329]_  = \new_[20856]_  & \new_[20845]_ ;
  assign \new_[3330]_  = \new_[20836]_  & \new_[20825]_ ;
  assign \new_[3331]_  = \new_[20816]_  & \new_[20805]_ ;
  assign \new_[3332]_  = \new_[20796]_  & \new_[20785]_ ;
  assign \new_[3333]_  = \new_[20776]_  & \new_[20765]_ ;
  assign \new_[3334]_  = \new_[20756]_  & \new_[20745]_ ;
  assign \new_[3335]_  = \new_[20736]_  & \new_[20725]_ ;
  assign \new_[3336]_  = \new_[20716]_  & \new_[20705]_ ;
  assign \new_[3337]_  = \new_[20696]_  & \new_[20685]_ ;
  assign \new_[3338]_  = \new_[20676]_  & \new_[20665]_ ;
  assign \new_[3339]_  = \new_[20656]_  & \new_[20645]_ ;
  assign \new_[3340]_  = \new_[20636]_  & \new_[20625]_ ;
  assign \new_[3341]_  = \new_[20616]_  & \new_[20605]_ ;
  assign \new_[3342]_  = \new_[20596]_  & \new_[20585]_ ;
  assign \new_[3343]_  = \new_[20576]_  & \new_[20565]_ ;
  assign \new_[3344]_  = \new_[20556]_  & \new_[20545]_ ;
  assign \new_[3345]_  = \new_[20536]_  & \new_[20525]_ ;
  assign \new_[3346]_  = \new_[20516]_  & \new_[20505]_ ;
  assign \new_[3347]_  = \new_[20496]_  & \new_[20485]_ ;
  assign \new_[3348]_  = \new_[20476]_  & \new_[20465]_ ;
  assign \new_[3349]_  = \new_[20456]_  & \new_[20445]_ ;
  assign \new_[3350]_  = \new_[20436]_  & \new_[20425]_ ;
  assign \new_[3351]_  = \new_[20416]_  & \new_[20405]_ ;
  assign \new_[3352]_  = \new_[20396]_  & \new_[20385]_ ;
  assign \new_[3353]_  = \new_[20376]_  & \new_[20365]_ ;
  assign \new_[3354]_  = \new_[20356]_  & \new_[20345]_ ;
  assign \new_[3355]_  = \new_[20336]_  & \new_[20325]_ ;
  assign \new_[3356]_  = \new_[20316]_  & \new_[20305]_ ;
  assign \new_[3357]_  = \new_[20296]_  & \new_[20285]_ ;
  assign \new_[3358]_  = \new_[20276]_  & \new_[20265]_ ;
  assign \new_[3359]_  = \new_[20256]_  & \new_[20245]_ ;
  assign \new_[3360]_  = \new_[20236]_  & \new_[20225]_ ;
  assign \new_[3361]_  = \new_[20216]_  & \new_[20205]_ ;
  assign \new_[3362]_  = \new_[20196]_  & \new_[20185]_ ;
  assign \new_[3363]_  = \new_[20176]_  & \new_[20165]_ ;
  assign \new_[3364]_  = \new_[20156]_  & \new_[20145]_ ;
  assign \new_[3365]_  = \new_[20136]_  & \new_[20125]_ ;
  assign \new_[3366]_  = \new_[20116]_  & \new_[20105]_ ;
  assign \new_[3367]_  = \new_[20096]_  & \new_[20085]_ ;
  assign \new_[3368]_  = \new_[20076]_  & \new_[20065]_ ;
  assign \new_[3369]_  = \new_[20056]_  & \new_[20045]_ ;
  assign \new_[3370]_  = \new_[20036]_  & \new_[20025]_ ;
  assign \new_[3371]_  = \new_[20016]_  & \new_[20005]_ ;
  assign \new_[3372]_  = \new_[19996]_  & \new_[19985]_ ;
  assign \new_[3373]_  = \new_[19976]_  & \new_[19965]_ ;
  assign \new_[3374]_  = \new_[19956]_  & \new_[19945]_ ;
  assign \new_[3375]_  = \new_[19936]_  & \new_[19925]_ ;
  assign \new_[3376]_  = \new_[19916]_  & \new_[19905]_ ;
  assign \new_[3377]_  = \new_[19896]_  & \new_[19885]_ ;
  assign \new_[3378]_  = \new_[19876]_  & \new_[19865]_ ;
  assign \new_[3379]_  = \new_[19856]_  & \new_[19845]_ ;
  assign \new_[3380]_  = \new_[19836]_  & \new_[19825]_ ;
  assign \new_[3381]_  = \new_[19816]_  & \new_[19805]_ ;
  assign \new_[3382]_  = \new_[19796]_  & \new_[19785]_ ;
  assign \new_[3383]_  = \new_[19776]_  & \new_[19765]_ ;
  assign \new_[3384]_  = \new_[19756]_  & \new_[19745]_ ;
  assign \new_[3385]_  = \new_[19736]_  & \new_[19725]_ ;
  assign \new_[3386]_  = \new_[19716]_  & \new_[19705]_ ;
  assign \new_[3387]_  = \new_[19696]_  & \new_[19685]_ ;
  assign \new_[3388]_  = \new_[19676]_  & \new_[19665]_ ;
  assign \new_[3389]_  = \new_[19656]_  & \new_[19645]_ ;
  assign \new_[3390]_  = \new_[19636]_  & \new_[19625]_ ;
  assign \new_[3391]_  = \new_[19616]_  & \new_[19605]_ ;
  assign \new_[3392]_  = \new_[19596]_  & \new_[19585]_ ;
  assign \new_[3393]_  = \new_[19576]_  & \new_[19565]_ ;
  assign \new_[3394]_  = \new_[19556]_  & \new_[19545]_ ;
  assign \new_[3395]_  = \new_[19536]_  & \new_[19525]_ ;
  assign \new_[3396]_  = \new_[19516]_  & \new_[19505]_ ;
  assign \new_[3397]_  = \new_[19496]_  & \new_[19485]_ ;
  assign \new_[3398]_  = \new_[19476]_  & \new_[19465]_ ;
  assign \new_[3399]_  = \new_[19456]_  & \new_[19445]_ ;
  assign \new_[3400]_  = \new_[19436]_  & \new_[19425]_ ;
  assign \new_[3401]_  = \new_[19416]_  & \new_[19405]_ ;
  assign \new_[3402]_  = \new_[19396]_  & \new_[19385]_ ;
  assign \new_[3403]_  = \new_[19376]_  & \new_[19365]_ ;
  assign \new_[3404]_  = \new_[19356]_  & \new_[19345]_ ;
  assign \new_[3405]_  = \new_[19336]_  & \new_[19325]_ ;
  assign \new_[3406]_  = \new_[19316]_  & \new_[19305]_ ;
  assign \new_[3407]_  = \new_[19296]_  & \new_[19285]_ ;
  assign \new_[3408]_  = \new_[19276]_  & \new_[19265]_ ;
  assign \new_[3409]_  = \new_[19256]_  & \new_[19245]_ ;
  assign \new_[3410]_  = \new_[19236]_  & \new_[19225]_ ;
  assign \new_[3411]_  = \new_[19216]_  & \new_[19205]_ ;
  assign \new_[3412]_  = \new_[19196]_  & \new_[19185]_ ;
  assign \new_[3413]_  = \new_[19176]_  & \new_[19165]_ ;
  assign \new_[3414]_  = \new_[19156]_  & \new_[19145]_ ;
  assign \new_[3415]_  = \new_[19136]_  & \new_[19125]_ ;
  assign \new_[3416]_  = \new_[19116]_  & \new_[19105]_ ;
  assign \new_[3417]_  = \new_[19096]_  & \new_[19085]_ ;
  assign \new_[3418]_  = \new_[19076]_  & \new_[19065]_ ;
  assign \new_[3419]_  = \new_[19056]_  & \new_[19045]_ ;
  assign \new_[3420]_  = \new_[19036]_  & \new_[19025]_ ;
  assign \new_[3421]_  = \new_[19016]_  & \new_[19005]_ ;
  assign \new_[3422]_  = \new_[18996]_  & \new_[18985]_ ;
  assign \new_[3423]_  = \new_[18976]_  & \new_[18965]_ ;
  assign \new_[3424]_  = \new_[18956]_  & \new_[18945]_ ;
  assign \new_[3425]_  = \new_[18936]_  & \new_[18925]_ ;
  assign \new_[3426]_  = \new_[18916]_  & \new_[18905]_ ;
  assign \new_[3427]_  = \new_[18896]_  & \new_[18885]_ ;
  assign \new_[3428]_  = \new_[18876]_  & \new_[18865]_ ;
  assign \new_[3429]_  = \new_[18856]_  & \new_[18845]_ ;
  assign \new_[3430]_  = \new_[18836]_  & \new_[18825]_ ;
  assign \new_[3431]_  = \new_[18816]_  & \new_[18805]_ ;
  assign \new_[3432]_  = \new_[18796]_  & \new_[18785]_ ;
  assign \new_[3433]_  = \new_[18776]_  & \new_[18765]_ ;
  assign \new_[3434]_  = \new_[18756]_  & \new_[18745]_ ;
  assign \new_[3435]_  = \new_[18736]_  & \new_[18725]_ ;
  assign \new_[3436]_  = \new_[18716]_  & \new_[18705]_ ;
  assign \new_[3437]_  = \new_[18696]_  & \new_[18685]_ ;
  assign \new_[3438]_  = \new_[18676]_  & \new_[18665]_ ;
  assign \new_[3439]_  = \new_[18656]_  & \new_[18645]_ ;
  assign \new_[3440]_  = \new_[18636]_  & \new_[18625]_ ;
  assign \new_[3441]_  = \new_[18616]_  & \new_[18605]_ ;
  assign \new_[3442]_  = \new_[18596]_  & \new_[18585]_ ;
  assign \new_[3443]_  = \new_[18576]_  & \new_[18565]_ ;
  assign \new_[3444]_  = \new_[18556]_  & \new_[18545]_ ;
  assign \new_[3445]_  = \new_[18536]_  & \new_[18525]_ ;
  assign \new_[3446]_  = \new_[18516]_  & \new_[18505]_ ;
  assign \new_[3447]_  = \new_[18496]_  & \new_[18485]_ ;
  assign \new_[3448]_  = \new_[18476]_  & \new_[18465]_ ;
  assign \new_[3449]_  = \new_[18456]_  & \new_[18445]_ ;
  assign \new_[3450]_  = \new_[18436]_  & \new_[18425]_ ;
  assign \new_[3451]_  = \new_[18416]_  & \new_[18405]_ ;
  assign \new_[3452]_  = \new_[18396]_  & \new_[18385]_ ;
  assign \new_[3453]_  = \new_[18376]_  & \new_[18365]_ ;
  assign \new_[3454]_  = \new_[18356]_  & \new_[18345]_ ;
  assign \new_[3455]_  = \new_[18336]_  & \new_[18325]_ ;
  assign \new_[3456]_  = \new_[18316]_  & \new_[18305]_ ;
  assign \new_[3457]_  = \new_[18296]_  & \new_[18285]_ ;
  assign \new_[3458]_  = \new_[18276]_  & \new_[18265]_ ;
  assign \new_[3459]_  = \new_[18256]_  & \new_[18245]_ ;
  assign \new_[3460]_  = \new_[18236]_  & \new_[18225]_ ;
  assign \new_[3461]_  = \new_[18216]_  & \new_[18205]_ ;
  assign \new_[3462]_  = \new_[18196]_  & \new_[18185]_ ;
  assign \new_[3463]_  = \new_[18176]_  & \new_[18165]_ ;
  assign \new_[3464]_  = \new_[18156]_  & \new_[18145]_ ;
  assign \new_[3465]_  = \new_[18136]_  & \new_[18125]_ ;
  assign \new_[3466]_  = \new_[18116]_  & \new_[18105]_ ;
  assign \new_[3467]_  = \new_[18096]_  & \new_[18085]_ ;
  assign \new_[3468]_  = \new_[18076]_  & \new_[18065]_ ;
  assign \new_[3469]_  = \new_[18056]_  & \new_[18045]_ ;
  assign \new_[3470]_  = \new_[18036]_  & \new_[18025]_ ;
  assign \new_[3471]_  = \new_[18016]_  & \new_[18005]_ ;
  assign \new_[3472]_  = \new_[17996]_  & \new_[17985]_ ;
  assign \new_[3473]_  = \new_[17976]_  & \new_[17965]_ ;
  assign \new_[3474]_  = \new_[17956]_  & \new_[17945]_ ;
  assign \new_[3475]_  = \new_[17936]_  & \new_[17925]_ ;
  assign \new_[3476]_  = \new_[17916]_  & \new_[17905]_ ;
  assign \new_[3477]_  = \new_[17896]_  & \new_[17885]_ ;
  assign \new_[3478]_  = \new_[17876]_  & \new_[17865]_ ;
  assign \new_[3479]_  = \new_[17856]_  & \new_[17845]_ ;
  assign \new_[3480]_  = \new_[17836]_  & \new_[17825]_ ;
  assign \new_[3481]_  = \new_[17816]_  & \new_[17805]_ ;
  assign \new_[3482]_  = \new_[17796]_  & \new_[17785]_ ;
  assign \new_[3483]_  = \new_[17776]_  & \new_[17765]_ ;
  assign \new_[3484]_  = \new_[17756]_  & \new_[17745]_ ;
  assign \new_[3485]_  = \new_[17736]_  & \new_[17725]_ ;
  assign \new_[3486]_  = \new_[17716]_  & \new_[17705]_ ;
  assign \new_[3487]_  = \new_[17696]_  & \new_[17685]_ ;
  assign \new_[3488]_  = \new_[17676]_  & \new_[17665]_ ;
  assign \new_[3489]_  = \new_[17656]_  & \new_[17645]_ ;
  assign \new_[3490]_  = \new_[17636]_  & \new_[17625]_ ;
  assign \new_[3491]_  = \new_[17616]_  & \new_[17605]_ ;
  assign \new_[3492]_  = \new_[17596]_  & \new_[17585]_ ;
  assign \new_[3493]_  = \new_[17576]_  & \new_[17565]_ ;
  assign \new_[3494]_  = \new_[17556]_  & \new_[17545]_ ;
  assign \new_[3495]_  = \new_[17536]_  & \new_[17525]_ ;
  assign \new_[3496]_  = \new_[17516]_  & \new_[17505]_ ;
  assign \new_[3497]_  = \new_[17496]_  & \new_[17485]_ ;
  assign \new_[3498]_  = \new_[17476]_  & \new_[17465]_ ;
  assign \new_[3499]_  = \new_[17456]_  & \new_[17447]_ ;
  assign \new_[3500]_  = \new_[17438]_  & \new_[17429]_ ;
  assign \new_[3501]_  = \new_[17420]_  & \new_[17411]_ ;
  assign \new_[3502]_  = \new_[17402]_  & \new_[17393]_ ;
  assign \new_[3503]_  = \new_[17384]_  & \new_[17375]_ ;
  assign \new_[3504]_  = \new_[17366]_  & \new_[17357]_ ;
  assign \new_[3505]_  = \new_[17348]_  & \new_[17339]_ ;
  assign \new_[3506]_  = \new_[17330]_  & \new_[17321]_ ;
  assign \new_[3507]_  = \new_[17312]_  & \new_[17303]_ ;
  assign \new_[3508]_  = \new_[17294]_  & \new_[17285]_ ;
  assign \new_[3509]_  = \new_[17276]_  & \new_[17267]_ ;
  assign \new_[3510]_  = \new_[17258]_  & \new_[17249]_ ;
  assign \new_[3511]_  = \new_[17240]_  & \new_[17231]_ ;
  assign \new_[3512]_  = \new_[17222]_  & \new_[17213]_ ;
  assign \new_[3513]_  = \new_[17204]_  & \new_[17195]_ ;
  assign \new_[3514]_  = \new_[17186]_  & \new_[17177]_ ;
  assign \new_[3515]_  = \new_[17168]_  & \new_[17159]_ ;
  assign \new_[3516]_  = \new_[17150]_  & \new_[17141]_ ;
  assign \new_[3517]_  = \new_[17132]_  & \new_[17123]_ ;
  assign \new_[3518]_  = \new_[17114]_  & \new_[17105]_ ;
  assign \new_[3519]_  = \new_[17096]_  & \new_[17087]_ ;
  assign \new_[3520]_  = \new_[17078]_  & \new_[17069]_ ;
  assign \new_[3521]_  = \new_[17060]_  & \new_[17051]_ ;
  assign \new_[3522]_  = \new_[17042]_  & \new_[17033]_ ;
  assign \new_[3523]_  = \new_[17024]_  & \new_[17015]_ ;
  assign \new_[3524]_  = \new_[17006]_  & \new_[16997]_ ;
  assign \new_[3525]_  = \new_[16988]_  & \new_[16979]_ ;
  assign \new_[3526]_  = \new_[16970]_  & \new_[16961]_ ;
  assign \new_[3527]_  = \new_[16952]_  & \new_[16943]_ ;
  assign \new_[3528]_  = \new_[16934]_  & \new_[16925]_ ;
  assign \new_[3529]_  = \new_[16916]_  & \new_[16907]_ ;
  assign \new_[3530]_  = \new_[16898]_  & \new_[16889]_ ;
  assign \new_[3531]_  = \new_[16880]_  & \new_[16871]_ ;
  assign \new_[3532]_  = \new_[16862]_  & \new_[16853]_ ;
  assign \new_[3533]_  = \new_[16844]_  & \new_[16835]_ ;
  assign \new_[3534]_  = \new_[16826]_  & \new_[16817]_ ;
  assign \new_[3535]_  = \new_[16808]_  & \new_[16799]_ ;
  assign \new_[3536]_  = \new_[16790]_  & \new_[16781]_ ;
  assign \new_[3537]_  = \new_[16772]_  & \new_[16763]_ ;
  assign \new_[3538]_  = \new_[16754]_  & \new_[16745]_ ;
  assign \new_[3539]_  = \new_[16736]_  & \new_[16727]_ ;
  assign \new_[3540]_  = \new_[16718]_  & \new_[16709]_ ;
  assign \new_[3541]_  = \new_[16700]_  & \new_[16691]_ ;
  assign \new_[3542]_  = \new_[16682]_  & \new_[16673]_ ;
  assign \new_[3543]_  = \new_[16664]_  & \new_[16655]_ ;
  assign \new_[3544]_  = \new_[16646]_  & \new_[16637]_ ;
  assign \new_[3545]_  = \new_[16628]_  & \new_[16619]_ ;
  assign \new_[3546]_  = \new_[16610]_  & \new_[16601]_ ;
  assign \new_[3547]_  = \new_[16592]_  & \new_[16583]_ ;
  assign \new_[3548]_  = \new_[16574]_  & \new_[16565]_ ;
  assign \new_[3549]_  = \new_[16556]_  & \new_[16547]_ ;
  assign \new_[3550]_  = \new_[16538]_  & \new_[16529]_ ;
  assign \new_[3551]_  = \new_[16520]_  & \new_[16511]_ ;
  assign \new_[3552]_  = \new_[16502]_  & \new_[16493]_ ;
  assign \new_[3553]_  = \new_[16484]_  & \new_[16475]_ ;
  assign \new_[3554]_  = \new_[16466]_  & \new_[16457]_ ;
  assign \new_[3555]_  = \new_[16448]_  & \new_[16439]_ ;
  assign \new_[3556]_  = \new_[16430]_  & \new_[16421]_ ;
  assign \new_[3557]_  = \new_[16412]_  & \new_[16403]_ ;
  assign \new_[3558]_  = \new_[16394]_  & \new_[16385]_ ;
  assign \new_[3559]_  = \new_[16376]_  & \new_[16367]_ ;
  assign \new_[3560]_  = \new_[16358]_  & \new_[16349]_ ;
  assign \new_[3561]_  = \new_[16340]_  & \new_[16331]_ ;
  assign \new_[3562]_  = \new_[16322]_  & \new_[16313]_ ;
  assign \new_[3563]_  = \new_[16304]_  & \new_[16295]_ ;
  assign \new_[3564]_  = \new_[16286]_  & \new_[16277]_ ;
  assign \new_[3565]_  = \new_[16268]_  & \new_[16259]_ ;
  assign \new_[3566]_  = \new_[16250]_  & \new_[16241]_ ;
  assign \new_[3567]_  = \new_[16232]_  & \new_[16223]_ ;
  assign \new_[3568]_  = \new_[16214]_  & \new_[16205]_ ;
  assign \new_[3569]_  = \new_[16196]_  & \new_[16187]_ ;
  assign \new_[3570]_  = \new_[16178]_  & \new_[16169]_ ;
  assign \new_[3571]_  = \new_[16160]_  & \new_[16151]_ ;
  assign \new_[3572]_  = \new_[16142]_  & \new_[16133]_ ;
  assign \new_[3573]_  = \new_[16124]_  & \new_[16115]_ ;
  assign \new_[3574]_  = \new_[16106]_  & \new_[16097]_ ;
  assign \new_[3575]_  = \new_[16088]_  & \new_[16079]_ ;
  assign \new_[3576]_  = \new_[16070]_  & \new_[16061]_ ;
  assign \new_[3577]_  = \new_[16052]_  & \new_[16043]_ ;
  assign \new_[3578]_  = \new_[16034]_  & \new_[16025]_ ;
  assign \new_[3579]_  = \new_[16016]_  & \new_[16007]_ ;
  assign \new_[3580]_  = \new_[15998]_  & \new_[15989]_ ;
  assign \new_[3581]_  = \new_[15980]_  & \new_[15971]_ ;
  assign \new_[3582]_  = \new_[15962]_  & \new_[15953]_ ;
  assign \new_[3583]_  = \new_[15944]_  & \new_[15935]_ ;
  assign \new_[3584]_  = \new_[15926]_  & \new_[15917]_ ;
  assign \new_[3585]_  = \new_[15908]_  & \new_[15899]_ ;
  assign \new_[3586]_  = \new_[15890]_  & \new_[15881]_ ;
  assign \new_[3587]_  = \new_[15872]_  & \new_[15863]_ ;
  assign \new_[3588]_  = \new_[15854]_  & \new_[15845]_ ;
  assign \new_[3589]_  = \new_[15836]_  & \new_[15827]_ ;
  assign \new_[3590]_  = \new_[15818]_  & \new_[15809]_ ;
  assign \new_[3591]_  = \new_[15800]_  & \new_[15791]_ ;
  assign \new_[3592]_  = \new_[15782]_  & \new_[15773]_ ;
  assign \new_[3593]_  = \new_[15764]_  & \new_[15755]_ ;
  assign \new_[3594]_  = \new_[15746]_  & \new_[15737]_ ;
  assign \new_[3595]_  = \new_[15728]_  & \new_[15719]_ ;
  assign \new_[3596]_  = \new_[15710]_  & \new_[15701]_ ;
  assign \new_[3597]_  = \new_[15692]_  & \new_[15683]_ ;
  assign \new_[3598]_  = \new_[15674]_  & \new_[15665]_ ;
  assign \new_[3599]_  = \new_[15656]_  & \new_[15647]_ ;
  assign \new_[3600]_  = \new_[15638]_  & \new_[15629]_ ;
  assign \new_[3601]_  = \new_[15620]_  & \new_[15611]_ ;
  assign \new_[3602]_  = \new_[15602]_  & \new_[15593]_ ;
  assign \new_[3603]_  = \new_[15584]_  & \new_[15575]_ ;
  assign \new_[3604]_  = \new_[15566]_  & \new_[15557]_ ;
  assign \new_[3605]_  = \new_[15548]_  & \new_[15539]_ ;
  assign \new_[3606]_  = \new_[15530]_  & \new_[15521]_ ;
  assign \new_[3607]_  = \new_[15512]_  & \new_[15503]_ ;
  assign \new_[3608]_  = \new_[15494]_  & \new_[15485]_ ;
  assign \new_[3609]_  = \new_[15476]_  & \new_[15467]_ ;
  assign \new_[3610]_  = \new_[15458]_  & \new_[15449]_ ;
  assign \new_[3611]_  = \new_[15440]_  & \new_[15431]_ ;
  assign \new_[3612]_  = \new_[15422]_  & \new_[15413]_ ;
  assign \new_[3613]_  = \new_[15404]_  & \new_[15395]_ ;
  assign \new_[3614]_  = \new_[15386]_  & \new_[15377]_ ;
  assign \new_[3615]_  = \new_[15368]_  & \new_[15359]_ ;
  assign \new_[3616]_  = \new_[15350]_  & \new_[15341]_ ;
  assign \new_[3617]_  = \new_[15332]_  & \new_[15323]_ ;
  assign \new_[3618]_  = \new_[15314]_  & \new_[15305]_ ;
  assign \new_[3619]_  = \new_[15296]_  & \new_[15287]_ ;
  assign \new_[3620]_  = \new_[15278]_  & \new_[15269]_ ;
  assign \new_[3621]_  = \new_[15260]_  & \new_[15251]_ ;
  assign \new_[3622]_  = \new_[15242]_  & \new_[15233]_ ;
  assign \new_[3623]_  = \new_[15224]_  & \new_[15215]_ ;
  assign \new_[3624]_  = \new_[15206]_  & \new_[15197]_ ;
  assign \new_[3625]_  = \new_[15188]_  & \new_[15179]_ ;
  assign \new_[3626]_  = \new_[15170]_  & \new_[15161]_ ;
  assign \new_[3627]_  = \new_[15152]_  & \new_[15143]_ ;
  assign \new_[3628]_  = \new_[15134]_  & \new_[15125]_ ;
  assign \new_[3629]_  = \new_[15116]_  & \new_[15107]_ ;
  assign \new_[3630]_  = \new_[15098]_  & \new_[15089]_ ;
  assign \new_[3631]_  = \new_[15080]_  & \new_[15071]_ ;
  assign \new_[3632]_  = \new_[15062]_  & \new_[15053]_ ;
  assign \new_[3633]_  = \new_[15044]_  & \new_[15035]_ ;
  assign \new_[3634]_  = \new_[15026]_  & \new_[15017]_ ;
  assign \new_[3635]_  = \new_[15008]_  & \new_[14999]_ ;
  assign \new_[3636]_  = \new_[14990]_  & \new_[14981]_ ;
  assign \new_[3637]_  = \new_[14972]_  & \new_[14963]_ ;
  assign \new_[3638]_  = \new_[14954]_  & \new_[14945]_ ;
  assign \new_[3639]_  = \new_[14936]_  & \new_[14927]_ ;
  assign \new_[3640]_  = \new_[14918]_  & \new_[14909]_ ;
  assign \new_[3641]_  = \new_[14900]_  & \new_[14891]_ ;
  assign \new_[3642]_  = \new_[14882]_  & \new_[14873]_ ;
  assign \new_[3643]_  = \new_[14864]_  & \new_[14855]_ ;
  assign \new_[3644]_  = \new_[14846]_  & \new_[14837]_ ;
  assign \new_[3645]_  = \new_[14828]_  & \new_[14819]_ ;
  assign \new_[3646]_  = \new_[14810]_  & \new_[14801]_ ;
  assign \new_[3647]_  = \new_[14792]_  & \new_[14783]_ ;
  assign \new_[3648]_  = \new_[14774]_  & \new_[14765]_ ;
  assign \new_[3649]_  = \new_[14756]_  & \new_[14747]_ ;
  assign \new_[3650]_  = \new_[14738]_  & \new_[14729]_ ;
  assign \new_[3651]_  = \new_[14720]_  & \new_[14711]_ ;
  assign \new_[3652]_  = \new_[14702]_  & \new_[14693]_ ;
  assign \new_[3653]_  = \new_[14684]_  & \new_[14675]_ ;
  assign \new_[3654]_  = \new_[14666]_  & \new_[14657]_ ;
  assign \new_[3655]_  = \new_[14648]_  & \new_[14639]_ ;
  assign \new_[3656]_  = \new_[14630]_  & \new_[14621]_ ;
  assign \new_[3657]_  = \new_[14612]_  & \new_[14603]_ ;
  assign \new_[3658]_  = \new_[14594]_  & \new_[14585]_ ;
  assign \new_[3659]_  = \new_[14576]_  & \new_[14567]_ ;
  assign \new_[3660]_  = \new_[14558]_  & \new_[14549]_ ;
  assign \new_[3661]_  = \new_[14540]_  & \new_[14531]_ ;
  assign \new_[3662]_  = \new_[14522]_  & \new_[14513]_ ;
  assign \new_[3663]_  = \new_[14504]_  & \new_[14495]_ ;
  assign \new_[3664]_  = \new_[14486]_  & \new_[14477]_ ;
  assign \new_[3665]_  = \new_[14468]_  & \new_[14459]_ ;
  assign \new_[3666]_  = \new_[14450]_  & \new_[14441]_ ;
  assign \new_[3667]_  = \new_[14432]_  & \new_[14423]_ ;
  assign \new_[3668]_  = \new_[14414]_  & \new_[14405]_ ;
  assign \new_[3669]_  = \new_[14396]_  & \new_[14387]_ ;
  assign \new_[3670]_  = \new_[14378]_  & \new_[14369]_ ;
  assign \new_[3671]_  = \new_[14360]_  & \new_[14351]_ ;
  assign \new_[3672]_  = \new_[14342]_  & \new_[14333]_ ;
  assign \new_[3673]_  = \new_[14324]_  & \new_[14315]_ ;
  assign \new_[3674]_  = \new_[14306]_  & \new_[14297]_ ;
  assign \new_[3675]_  = \new_[14288]_  & \new_[14279]_ ;
  assign \new_[3676]_  = \new_[14270]_  & \new_[14261]_ ;
  assign \new_[3677]_  = \new_[14252]_  & \new_[14243]_ ;
  assign \new_[3678]_  = \new_[14234]_  & \new_[14225]_ ;
  assign \new_[3679]_  = \new_[14216]_  & \new_[14207]_ ;
  assign \new_[3680]_  = \new_[14198]_  & \new_[14189]_ ;
  assign \new_[3681]_  = \new_[14180]_  & \new_[14171]_ ;
  assign \new_[3682]_  = \new_[14162]_  & \new_[14153]_ ;
  assign \new_[3683]_  = \new_[14144]_  & \new_[14135]_ ;
  assign \new_[3684]_  = \new_[14126]_  & \new_[14117]_ ;
  assign \new_[3685]_  = \new_[14108]_  & \new_[14099]_ ;
  assign \new_[3686]_  = \new_[14090]_  & \new_[14081]_ ;
  assign \new_[3687]_  = \new_[14072]_  & \new_[14063]_ ;
  assign \new_[3688]_  = \new_[14054]_  & \new_[14045]_ ;
  assign \new_[3689]_  = \new_[14036]_  & \new_[14027]_ ;
  assign \new_[3690]_  = \new_[14018]_  & \new_[14009]_ ;
  assign \new_[3691]_  = \new_[14000]_  & \new_[13991]_ ;
  assign \new_[3692]_  = \new_[13982]_  & \new_[13973]_ ;
  assign \new_[3693]_  = \new_[13964]_  & \new_[13955]_ ;
  assign \new_[3694]_  = \new_[13946]_  & \new_[13937]_ ;
  assign \new_[3695]_  = \new_[13928]_  & \new_[13919]_ ;
  assign \new_[3696]_  = \new_[13910]_  & \new_[13901]_ ;
  assign \new_[3697]_  = \new_[13892]_  & \new_[13883]_ ;
  assign \new_[3698]_  = \new_[13874]_  & \new_[13865]_ ;
  assign \new_[3699]_  = \new_[13856]_  & \new_[13847]_ ;
  assign \new_[3700]_  = \new_[13838]_  & \new_[13829]_ ;
  assign \new_[3701]_  = \new_[13820]_  & \new_[13811]_ ;
  assign \new_[3702]_  = \new_[13802]_  & \new_[13793]_ ;
  assign \new_[3703]_  = \new_[13784]_  & \new_[13775]_ ;
  assign \new_[3704]_  = \new_[13766]_  & \new_[13757]_ ;
  assign \new_[3705]_  = \new_[13748]_  & \new_[13739]_ ;
  assign \new_[3706]_  = \new_[13730]_  & \new_[13721]_ ;
  assign \new_[3707]_  = \new_[13712]_  & \new_[13703]_ ;
  assign \new_[3708]_  = \new_[13694]_  & \new_[13685]_ ;
  assign \new_[3709]_  = \new_[13676]_  & \new_[13667]_ ;
  assign \new_[3710]_  = \new_[13658]_  & \new_[13649]_ ;
  assign \new_[3711]_  = \new_[13640]_  & \new_[13631]_ ;
  assign \new_[3712]_  = \new_[13622]_  & \new_[13613]_ ;
  assign \new_[3713]_  = \new_[13604]_  & \new_[13595]_ ;
  assign \new_[3714]_  = \new_[13586]_  & \new_[13577]_ ;
  assign \new_[3715]_  = \new_[13568]_  & \new_[13559]_ ;
  assign \new_[3716]_  = \new_[13550]_  & \new_[13541]_ ;
  assign \new_[3717]_  = \new_[13532]_  & \new_[13523]_ ;
  assign \new_[3718]_  = \new_[13514]_  & \new_[13505]_ ;
  assign \new_[3719]_  = \new_[13496]_  & \new_[13487]_ ;
  assign \new_[3720]_  = \new_[13478]_  & \new_[13469]_ ;
  assign \new_[3721]_  = \new_[13460]_  & \new_[13451]_ ;
  assign \new_[3722]_  = \new_[13442]_  & \new_[13433]_ ;
  assign \new_[3723]_  = \new_[13424]_  & \new_[13415]_ ;
  assign \new_[3724]_  = \new_[13406]_  & \new_[13397]_ ;
  assign \new_[3725]_  = \new_[13388]_  & \new_[13379]_ ;
  assign \new_[3726]_  = \new_[13370]_  & \new_[13361]_ ;
  assign \new_[3727]_  = \new_[13352]_  & \new_[13343]_ ;
  assign \new_[3728]_  = \new_[13334]_  & \new_[13325]_ ;
  assign \new_[3729]_  = \new_[13316]_  & \new_[13307]_ ;
  assign \new_[3730]_  = \new_[13298]_  & \new_[13289]_ ;
  assign \new_[3731]_  = \new_[13280]_  & \new_[13271]_ ;
  assign \new_[3732]_  = \new_[13262]_  & \new_[13253]_ ;
  assign \new_[3733]_  = \new_[13244]_  & \new_[13235]_ ;
  assign \new_[3734]_  = \new_[13226]_  & \new_[13217]_ ;
  assign \new_[3735]_  = \new_[13208]_  & \new_[13199]_ ;
  assign \new_[3736]_  = \new_[13190]_  & \new_[13181]_ ;
  assign \new_[3737]_  = \new_[13172]_  & \new_[13163]_ ;
  assign \new_[3738]_  = \new_[13154]_  & \new_[13145]_ ;
  assign \new_[3739]_  = \new_[13136]_  & \new_[13127]_ ;
  assign \new_[3740]_  = \new_[13118]_  & \new_[13109]_ ;
  assign \new_[3741]_  = \new_[13100]_  & \new_[13091]_ ;
  assign \new_[3742]_  = \new_[13082]_  & \new_[13073]_ ;
  assign \new_[3743]_  = \new_[13064]_  & \new_[13055]_ ;
  assign \new_[3744]_  = \new_[13046]_  & \new_[13037]_ ;
  assign \new_[3745]_  = \new_[13028]_  & \new_[13019]_ ;
  assign \new_[3746]_  = \new_[13010]_  & \new_[13001]_ ;
  assign \new_[3747]_  = \new_[12992]_  & \new_[12983]_ ;
  assign \new_[3748]_  = \new_[12974]_  & \new_[12965]_ ;
  assign \new_[3749]_  = \new_[12956]_  & \new_[12947]_ ;
  assign \new_[3750]_  = \new_[12938]_  & \new_[12929]_ ;
  assign \new_[3751]_  = \new_[12920]_  & \new_[12911]_ ;
  assign \new_[3752]_  = \new_[12902]_  & \new_[12893]_ ;
  assign \new_[3753]_  = \new_[12884]_  & \new_[12875]_ ;
  assign \new_[3754]_  = \new_[12866]_  & \new_[12857]_ ;
  assign \new_[3755]_  = \new_[12848]_  & \new_[12839]_ ;
  assign \new_[3756]_  = \new_[12830]_  & \new_[12821]_ ;
  assign \new_[3757]_  = \new_[12812]_  & \new_[12803]_ ;
  assign \new_[3758]_  = \new_[12794]_  & \new_[12785]_ ;
  assign \new_[3759]_  = \new_[12776]_  & \new_[12767]_ ;
  assign \new_[3760]_  = \new_[12758]_  & \new_[12749]_ ;
  assign \new_[3761]_  = \new_[12740]_  & \new_[12731]_ ;
  assign \new_[3762]_  = \new_[12722]_  & \new_[12713]_ ;
  assign \new_[3763]_  = \new_[12704]_  & \new_[12695]_ ;
  assign \new_[3764]_  = \new_[12686]_  & \new_[12677]_ ;
  assign \new_[3765]_  = \new_[12668]_  & \new_[12659]_ ;
  assign \new_[3766]_  = \new_[12650]_  & \new_[12641]_ ;
  assign \new_[3767]_  = \new_[12632]_  & \new_[12623]_ ;
  assign \new_[3768]_  = \new_[12614]_  & \new_[12605]_ ;
  assign \new_[3769]_  = \new_[12596]_  & \new_[12587]_ ;
  assign \new_[3770]_  = \new_[12578]_  & \new_[12569]_ ;
  assign \new_[3771]_  = \new_[12560]_  & \new_[12551]_ ;
  assign \new_[3772]_  = \new_[12542]_  & \new_[12533]_ ;
  assign \new_[3773]_  = \new_[12524]_  & \new_[12515]_ ;
  assign \new_[3774]_  = \new_[12506]_  & \new_[12497]_ ;
  assign \new_[3775]_  = \new_[12488]_  & \new_[12479]_ ;
  assign \new_[3776]_  = \new_[12470]_  & \new_[12461]_ ;
  assign \new_[3777]_  = \new_[12452]_  & \new_[12443]_ ;
  assign \new_[3778]_  = \new_[12434]_  & \new_[12425]_ ;
  assign \new_[3779]_  = \new_[12416]_  & \new_[12407]_ ;
  assign \new_[3780]_  = \new_[12398]_  & \new_[12389]_ ;
  assign \new_[3781]_  = \new_[12380]_  & \new_[12371]_ ;
  assign \new_[3782]_  = \new_[12362]_  & \new_[12353]_ ;
  assign \new_[3783]_  = \new_[12344]_  & \new_[12335]_ ;
  assign \new_[3784]_  = \new_[12328]_  & \new_[12319]_ ;
  assign \new_[3785]_  = \new_[12312]_  & \new_[12303]_ ;
  assign \new_[3786]_  = \new_[12296]_  & \new_[12287]_ ;
  assign \new_[3787]_  = \new_[12280]_  & \new_[12271]_ ;
  assign \new_[3788]_  = \new_[12264]_  & \new_[12255]_ ;
  assign \new_[3789]_  = \new_[12248]_  & \new_[12239]_ ;
  assign \new_[3790]_  = \new_[12232]_  & \new_[12223]_ ;
  assign \new_[3791]_  = \new_[12216]_  & \new_[12207]_ ;
  assign \new_[3792]_  = \new_[12200]_  & \new_[12191]_ ;
  assign \new_[3793]_  = \new_[12184]_  & \new_[12175]_ ;
  assign \new_[3794]_  = \new_[12168]_  & \new_[12159]_ ;
  assign \new_[3795]_  = \new_[12152]_  & \new_[12143]_ ;
  assign \new_[3796]_  = \new_[12136]_  & \new_[12127]_ ;
  assign \new_[3797]_  = \new_[12120]_  & \new_[12111]_ ;
  assign \new_[3798]_  = \new_[12104]_  & \new_[12095]_ ;
  assign \new_[3799]_  = \new_[12088]_  & \new_[12079]_ ;
  assign \new_[3800]_  = \new_[12072]_  & \new_[12063]_ ;
  assign \new_[3801]_  = \new_[12056]_  & \new_[12047]_ ;
  assign \new_[3802]_  = \new_[12040]_  & \new_[12031]_ ;
  assign \new_[3803]_  = \new_[12024]_  & \new_[12015]_ ;
  assign \new_[3804]_  = \new_[12008]_  & \new_[11999]_ ;
  assign \new_[3805]_  = \new_[11992]_  & \new_[11983]_ ;
  assign \new_[3806]_  = \new_[11976]_  & \new_[11967]_ ;
  assign \new_[3807]_  = \new_[11960]_  & \new_[11953]_ ;
  assign \new_[3808]_  = \new_[11946]_  & \new_[11939]_ ;
  assign \new_[3809]_  = \new_[11932]_  & \new_[11925]_ ;
  assign \new_[3810]_  = \new_[11918]_  & \new_[11911]_ ;
  assign \new_[3811]_  = \new_[11904]_  & \new_[11897]_ ;
  assign \new_[3812]_  = \new_[11890]_  & \new_[11883]_ ;
  assign \new_[3813]_  = \new_[11876]_  & \new_[11869]_ ;
  assign \new_[3814]_  = \new_[11862]_  & \new_[11855]_ ;
  assign \new_[3815]_  = \new_[11848]_  & \new_[11841]_ ;
  assign \new_[3816]_  = \new_[11834]_  & \new_[11827]_ ;
  assign \new_[3817]_  = \new_[11820]_  & \new_[11813]_ ;
  assign \new_[3818]_  = \new_[11806]_  & \new_[11799]_ ;
  assign \new_[3819]_  = \new_[11792]_  & \new_[11785]_ ;
  assign \new_[3820]_  = \new_[11778]_  & \new_[11771]_ ;
  assign \new_[3821]_  = \new_[11764]_  & \new_[11757]_ ;
  assign \new_[3822]_  = \new_[11750]_  & \new_[11743]_ ;
  assign \new_[3823]_  = \new_[11736]_  & \new_[11729]_ ;
  assign \new_[3824]_  = \new_[11722]_  & \new_[11715]_ ;
  assign \new_[3825]_  = \new_[11708]_  & \new_[11701]_ ;
  assign \new_[3826]_  = \new_[11694]_  & \new_[11687]_ ;
  assign \new_[3827]_  = \new_[11680]_  & \new_[11673]_ ;
  assign \new_[3828]_  = \new_[11666]_  & \new_[11659]_ ;
  assign \new_[3829]_  = \new_[11652]_  & \new_[11645]_ ;
  assign \new_[3830]_  = \new_[11638]_  & \new_[11631]_ ;
  assign \new_[3831]_  = \new_[11624]_  & \new_[11617]_ ;
  assign \new_[3832]_  = \new_[11610]_  & \new_[11603]_ ;
  assign \new_[3833]_  = \new_[11596]_  & \new_[11589]_ ;
  assign \new_[3834]_  = \new_[11582]_  & \new_[11575]_ ;
  assign \new_[3835]_  = \new_[11568]_  & \new_[11561]_ ;
  assign \new_[3836]_  = \new_[11554]_  & \new_[11547]_ ;
  assign \new_[3837]_  = \new_[11540]_  & \new_[11533]_ ;
  assign \new_[3838]_  = \new_[11526]_  & \new_[11519]_ ;
  assign \new_[3842]_  = \new_[3836]_  | \new_[3837]_ ;
  assign \new_[3843]_  = \new_[3838]_  | \new_[3842]_ ;
  assign \new_[3846]_  = \new_[3834]_  | \new_[3835]_ ;
  assign \new_[3849]_  = \new_[3832]_  | \new_[3833]_ ;
  assign \new_[3850]_  = \new_[3849]_  | \new_[3846]_ ;
  assign \new_[3851]_  = \new_[3850]_  | \new_[3843]_ ;
  assign \new_[3855]_  = \new_[3829]_  | \new_[3830]_ ;
  assign \new_[3856]_  = \new_[3831]_  | \new_[3855]_ ;
  assign \new_[3859]_  = \new_[3827]_  | \new_[3828]_ ;
  assign \new_[3862]_  = \new_[3825]_  | \new_[3826]_ ;
  assign \new_[3863]_  = \new_[3862]_  | \new_[3859]_ ;
  assign \new_[3864]_  = \new_[3863]_  | \new_[3856]_ ;
  assign \new_[3865]_  = \new_[3864]_  | \new_[3851]_ ;
  assign \new_[3869]_  = \new_[3822]_  | \new_[3823]_ ;
  assign \new_[3870]_  = \new_[3824]_  | \new_[3869]_ ;
  assign \new_[3873]_  = \new_[3820]_  | \new_[3821]_ ;
  assign \new_[3876]_  = \new_[3818]_  | \new_[3819]_ ;
  assign \new_[3877]_  = \new_[3876]_  | \new_[3873]_ ;
  assign \new_[3878]_  = \new_[3877]_  | \new_[3870]_ ;
  assign \new_[3881]_  = \new_[3816]_  | \new_[3817]_ ;
  assign \new_[3884]_  = \new_[3814]_  | \new_[3815]_ ;
  assign \new_[3885]_  = \new_[3884]_  | \new_[3881]_ ;
  assign \new_[3888]_  = \new_[3812]_  | \new_[3813]_ ;
  assign \new_[3891]_  = \new_[3810]_  | \new_[3811]_ ;
  assign \new_[3892]_  = \new_[3891]_  | \new_[3888]_ ;
  assign \new_[3893]_  = \new_[3892]_  | \new_[3885]_ ;
  assign \new_[3894]_  = \new_[3893]_  | \new_[3878]_ ;
  assign \new_[3895]_  = \new_[3894]_  | \new_[3865]_ ;
  assign \new_[3899]_  = \new_[3807]_  | \new_[3808]_ ;
  assign \new_[3900]_  = \new_[3809]_  | \new_[3899]_ ;
  assign \new_[3903]_  = \new_[3805]_  | \new_[3806]_ ;
  assign \new_[3906]_  = \new_[3803]_  | \new_[3804]_ ;
  assign \new_[3907]_  = \new_[3906]_  | \new_[3903]_ ;
  assign \new_[3908]_  = \new_[3907]_  | \new_[3900]_ ;
  assign \new_[3911]_  = \new_[3801]_  | \new_[3802]_ ;
  assign \new_[3914]_  = \new_[3799]_  | \new_[3800]_ ;
  assign \new_[3915]_  = \new_[3914]_  | \new_[3911]_ ;
  assign \new_[3918]_  = \new_[3797]_  | \new_[3798]_ ;
  assign \new_[3921]_  = \new_[3795]_  | \new_[3796]_ ;
  assign \new_[3922]_  = \new_[3921]_  | \new_[3918]_ ;
  assign \new_[3923]_  = \new_[3922]_  | \new_[3915]_ ;
  assign \new_[3924]_  = \new_[3923]_  | \new_[3908]_ ;
  assign \new_[3928]_  = \new_[3792]_  | \new_[3793]_ ;
  assign \new_[3929]_  = \new_[3794]_  | \new_[3928]_ ;
  assign \new_[3932]_  = \new_[3790]_  | \new_[3791]_ ;
  assign \new_[3935]_  = \new_[3788]_  | \new_[3789]_ ;
  assign \new_[3936]_  = \new_[3935]_  | \new_[3932]_ ;
  assign \new_[3937]_  = \new_[3936]_  | \new_[3929]_ ;
  assign \new_[3940]_  = \new_[3786]_  | \new_[3787]_ ;
  assign \new_[3943]_  = \new_[3784]_  | \new_[3785]_ ;
  assign \new_[3944]_  = \new_[3943]_  | \new_[3940]_ ;
  assign \new_[3947]_  = \new_[3782]_  | \new_[3783]_ ;
  assign \new_[3950]_  = \new_[3780]_  | \new_[3781]_ ;
  assign \new_[3951]_  = \new_[3950]_  | \new_[3947]_ ;
  assign \new_[3952]_  = \new_[3951]_  | \new_[3944]_ ;
  assign \new_[3953]_  = \new_[3952]_  | \new_[3937]_ ;
  assign \new_[3954]_  = \new_[3953]_  | \new_[3924]_ ;
  assign \new_[3955]_  = \new_[3954]_  | \new_[3895]_ ;
  assign \new_[3959]_  = \new_[3777]_  | \new_[3778]_ ;
  assign \new_[3960]_  = \new_[3779]_  | \new_[3959]_ ;
  assign \new_[3963]_  = \new_[3775]_  | \new_[3776]_ ;
  assign \new_[3966]_  = \new_[3773]_  | \new_[3774]_ ;
  assign \new_[3967]_  = \new_[3966]_  | \new_[3963]_ ;
  assign \new_[3968]_  = \new_[3967]_  | \new_[3960]_ ;
  assign \new_[3971]_  = \new_[3771]_  | \new_[3772]_ ;
  assign \new_[3974]_  = \new_[3769]_  | \new_[3770]_ ;
  assign \new_[3975]_  = \new_[3974]_  | \new_[3971]_ ;
  assign \new_[3978]_  = \new_[3767]_  | \new_[3768]_ ;
  assign \new_[3981]_  = \new_[3765]_  | \new_[3766]_ ;
  assign \new_[3982]_  = \new_[3981]_  | \new_[3978]_ ;
  assign \new_[3983]_  = \new_[3982]_  | \new_[3975]_ ;
  assign \new_[3984]_  = \new_[3983]_  | \new_[3968]_ ;
  assign \new_[3988]_  = \new_[3762]_  | \new_[3763]_ ;
  assign \new_[3989]_  = \new_[3764]_  | \new_[3988]_ ;
  assign \new_[3992]_  = \new_[3760]_  | \new_[3761]_ ;
  assign \new_[3995]_  = \new_[3758]_  | \new_[3759]_ ;
  assign \new_[3996]_  = \new_[3995]_  | \new_[3992]_ ;
  assign \new_[3997]_  = \new_[3996]_  | \new_[3989]_ ;
  assign \new_[4000]_  = \new_[3756]_  | \new_[3757]_ ;
  assign \new_[4003]_  = \new_[3754]_  | \new_[3755]_ ;
  assign \new_[4004]_  = \new_[4003]_  | \new_[4000]_ ;
  assign \new_[4007]_  = \new_[3752]_  | \new_[3753]_ ;
  assign \new_[4010]_  = \new_[3750]_  | \new_[3751]_ ;
  assign \new_[4011]_  = \new_[4010]_  | \new_[4007]_ ;
  assign \new_[4012]_  = \new_[4011]_  | \new_[4004]_ ;
  assign \new_[4013]_  = \new_[4012]_  | \new_[3997]_ ;
  assign \new_[4014]_  = \new_[4013]_  | \new_[3984]_ ;
  assign \new_[4018]_  = \new_[3747]_  | \new_[3748]_ ;
  assign \new_[4019]_  = \new_[3749]_  | \new_[4018]_ ;
  assign \new_[4022]_  = \new_[3745]_  | \new_[3746]_ ;
  assign \new_[4025]_  = \new_[3743]_  | \new_[3744]_ ;
  assign \new_[4026]_  = \new_[4025]_  | \new_[4022]_ ;
  assign \new_[4027]_  = \new_[4026]_  | \new_[4019]_ ;
  assign \new_[4030]_  = \new_[3741]_  | \new_[3742]_ ;
  assign \new_[4033]_  = \new_[3739]_  | \new_[3740]_ ;
  assign \new_[4034]_  = \new_[4033]_  | \new_[4030]_ ;
  assign \new_[4037]_  = \new_[3737]_  | \new_[3738]_ ;
  assign \new_[4040]_  = \new_[3735]_  | \new_[3736]_ ;
  assign \new_[4041]_  = \new_[4040]_  | \new_[4037]_ ;
  assign \new_[4042]_  = \new_[4041]_  | \new_[4034]_ ;
  assign \new_[4043]_  = \new_[4042]_  | \new_[4027]_ ;
  assign \new_[4047]_  = \new_[3732]_  | \new_[3733]_ ;
  assign \new_[4048]_  = \new_[3734]_  | \new_[4047]_ ;
  assign \new_[4051]_  = \new_[3730]_  | \new_[3731]_ ;
  assign \new_[4054]_  = \new_[3728]_  | \new_[3729]_ ;
  assign \new_[4055]_  = \new_[4054]_  | \new_[4051]_ ;
  assign \new_[4056]_  = \new_[4055]_  | \new_[4048]_ ;
  assign \new_[4059]_  = \new_[3726]_  | \new_[3727]_ ;
  assign \new_[4062]_  = \new_[3724]_  | \new_[3725]_ ;
  assign \new_[4063]_  = \new_[4062]_  | \new_[4059]_ ;
  assign \new_[4066]_  = \new_[3722]_  | \new_[3723]_ ;
  assign \new_[4069]_  = \new_[3720]_  | \new_[3721]_ ;
  assign \new_[4070]_  = \new_[4069]_  | \new_[4066]_ ;
  assign \new_[4071]_  = \new_[4070]_  | \new_[4063]_ ;
  assign \new_[4072]_  = \new_[4071]_  | \new_[4056]_ ;
  assign \new_[4073]_  = \new_[4072]_  | \new_[4043]_ ;
  assign \new_[4074]_  = \new_[4073]_  | \new_[4014]_ ;
  assign \new_[4075]_  = \new_[4074]_  | \new_[3955]_ ;
  assign \new_[4079]_  = \new_[3717]_  | \new_[3718]_ ;
  assign \new_[4080]_  = \new_[3719]_  | \new_[4079]_ ;
  assign \new_[4083]_  = \new_[3715]_  | \new_[3716]_ ;
  assign \new_[4086]_  = \new_[3713]_  | \new_[3714]_ ;
  assign \new_[4087]_  = \new_[4086]_  | \new_[4083]_ ;
  assign \new_[4088]_  = \new_[4087]_  | \new_[4080]_ ;
  assign \new_[4091]_  = \new_[3711]_  | \new_[3712]_ ;
  assign \new_[4094]_  = \new_[3709]_  | \new_[3710]_ ;
  assign \new_[4095]_  = \new_[4094]_  | \new_[4091]_ ;
  assign \new_[4098]_  = \new_[3707]_  | \new_[3708]_ ;
  assign \new_[4101]_  = \new_[3705]_  | \new_[3706]_ ;
  assign \new_[4102]_  = \new_[4101]_  | \new_[4098]_ ;
  assign \new_[4103]_  = \new_[4102]_  | \new_[4095]_ ;
  assign \new_[4104]_  = \new_[4103]_  | \new_[4088]_ ;
  assign \new_[4108]_  = \new_[3702]_  | \new_[3703]_ ;
  assign \new_[4109]_  = \new_[3704]_  | \new_[4108]_ ;
  assign \new_[4112]_  = \new_[3700]_  | \new_[3701]_ ;
  assign \new_[4115]_  = \new_[3698]_  | \new_[3699]_ ;
  assign \new_[4116]_  = \new_[4115]_  | \new_[4112]_ ;
  assign \new_[4117]_  = \new_[4116]_  | \new_[4109]_ ;
  assign \new_[4120]_  = \new_[3696]_  | \new_[3697]_ ;
  assign \new_[4123]_  = \new_[3694]_  | \new_[3695]_ ;
  assign \new_[4124]_  = \new_[4123]_  | \new_[4120]_ ;
  assign \new_[4127]_  = \new_[3692]_  | \new_[3693]_ ;
  assign \new_[4130]_  = \new_[3690]_  | \new_[3691]_ ;
  assign \new_[4131]_  = \new_[4130]_  | \new_[4127]_ ;
  assign \new_[4132]_  = \new_[4131]_  | \new_[4124]_ ;
  assign \new_[4133]_  = \new_[4132]_  | \new_[4117]_ ;
  assign \new_[4134]_  = \new_[4133]_  | \new_[4104]_ ;
  assign \new_[4138]_  = \new_[3687]_  | \new_[3688]_ ;
  assign \new_[4139]_  = \new_[3689]_  | \new_[4138]_ ;
  assign \new_[4142]_  = \new_[3685]_  | \new_[3686]_ ;
  assign \new_[4145]_  = \new_[3683]_  | \new_[3684]_ ;
  assign \new_[4146]_  = \new_[4145]_  | \new_[4142]_ ;
  assign \new_[4147]_  = \new_[4146]_  | \new_[4139]_ ;
  assign \new_[4150]_  = \new_[3681]_  | \new_[3682]_ ;
  assign \new_[4153]_  = \new_[3679]_  | \new_[3680]_ ;
  assign \new_[4154]_  = \new_[4153]_  | \new_[4150]_ ;
  assign \new_[4157]_  = \new_[3677]_  | \new_[3678]_ ;
  assign \new_[4160]_  = \new_[3675]_  | \new_[3676]_ ;
  assign \new_[4161]_  = \new_[4160]_  | \new_[4157]_ ;
  assign \new_[4162]_  = \new_[4161]_  | \new_[4154]_ ;
  assign \new_[4163]_  = \new_[4162]_  | \new_[4147]_ ;
  assign \new_[4167]_  = \new_[3672]_  | \new_[3673]_ ;
  assign \new_[4168]_  = \new_[3674]_  | \new_[4167]_ ;
  assign \new_[4171]_  = \new_[3670]_  | \new_[3671]_ ;
  assign \new_[4174]_  = \new_[3668]_  | \new_[3669]_ ;
  assign \new_[4175]_  = \new_[4174]_  | \new_[4171]_ ;
  assign \new_[4176]_  = \new_[4175]_  | \new_[4168]_ ;
  assign \new_[4179]_  = \new_[3666]_  | \new_[3667]_ ;
  assign \new_[4182]_  = \new_[3664]_  | \new_[3665]_ ;
  assign \new_[4183]_  = \new_[4182]_  | \new_[4179]_ ;
  assign \new_[4186]_  = \new_[3662]_  | \new_[3663]_ ;
  assign \new_[4189]_  = \new_[3660]_  | \new_[3661]_ ;
  assign \new_[4190]_  = \new_[4189]_  | \new_[4186]_ ;
  assign \new_[4191]_  = \new_[4190]_  | \new_[4183]_ ;
  assign \new_[4192]_  = \new_[4191]_  | \new_[4176]_ ;
  assign \new_[4193]_  = \new_[4192]_  | \new_[4163]_ ;
  assign \new_[4194]_  = \new_[4193]_  | \new_[4134]_ ;
  assign \new_[4198]_  = \new_[3657]_  | \new_[3658]_ ;
  assign \new_[4199]_  = \new_[3659]_  | \new_[4198]_ ;
  assign \new_[4202]_  = \new_[3655]_  | \new_[3656]_ ;
  assign \new_[4205]_  = \new_[3653]_  | \new_[3654]_ ;
  assign \new_[4206]_  = \new_[4205]_  | \new_[4202]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4199]_ ;
  assign \new_[4210]_  = \new_[3651]_  | \new_[3652]_ ;
  assign \new_[4213]_  = \new_[3649]_  | \new_[3650]_ ;
  assign \new_[4214]_  = \new_[4213]_  | \new_[4210]_ ;
  assign \new_[4217]_  = \new_[3647]_  | \new_[3648]_ ;
  assign \new_[4220]_  = \new_[3645]_  | \new_[3646]_ ;
  assign \new_[4221]_  = \new_[4220]_  | \new_[4217]_ ;
  assign \new_[4222]_  = \new_[4221]_  | \new_[4214]_ ;
  assign \new_[4223]_  = \new_[4222]_  | \new_[4207]_ ;
  assign \new_[4227]_  = \new_[3642]_  | \new_[3643]_ ;
  assign \new_[4228]_  = \new_[3644]_  | \new_[4227]_ ;
  assign \new_[4231]_  = \new_[3640]_  | \new_[3641]_ ;
  assign \new_[4234]_  = \new_[3638]_  | \new_[3639]_ ;
  assign \new_[4235]_  = \new_[4234]_  | \new_[4231]_ ;
  assign \new_[4236]_  = \new_[4235]_  | \new_[4228]_ ;
  assign \new_[4239]_  = \new_[3636]_  | \new_[3637]_ ;
  assign \new_[4242]_  = \new_[3634]_  | \new_[3635]_ ;
  assign \new_[4243]_  = \new_[4242]_  | \new_[4239]_ ;
  assign \new_[4246]_  = \new_[3632]_  | \new_[3633]_ ;
  assign \new_[4249]_  = \new_[3630]_  | \new_[3631]_ ;
  assign \new_[4250]_  = \new_[4249]_  | \new_[4246]_ ;
  assign \new_[4251]_  = \new_[4250]_  | \new_[4243]_ ;
  assign \new_[4252]_  = \new_[4251]_  | \new_[4236]_ ;
  assign \new_[4253]_  = \new_[4252]_  | \new_[4223]_ ;
  assign \new_[4257]_  = \new_[3627]_  | \new_[3628]_ ;
  assign \new_[4258]_  = \new_[3629]_  | \new_[4257]_ ;
  assign \new_[4261]_  = \new_[3625]_  | \new_[3626]_ ;
  assign \new_[4264]_  = \new_[3623]_  | \new_[3624]_ ;
  assign \new_[4265]_  = \new_[4264]_  | \new_[4261]_ ;
  assign \new_[4266]_  = \new_[4265]_  | \new_[4258]_ ;
  assign \new_[4269]_  = \new_[3621]_  | \new_[3622]_ ;
  assign \new_[4272]_  = \new_[3619]_  | \new_[3620]_ ;
  assign \new_[4273]_  = \new_[4272]_  | \new_[4269]_ ;
  assign \new_[4276]_  = \new_[3617]_  | \new_[3618]_ ;
  assign \new_[4279]_  = \new_[3615]_  | \new_[3616]_ ;
  assign \new_[4280]_  = \new_[4279]_  | \new_[4276]_ ;
  assign \new_[4281]_  = \new_[4280]_  | \new_[4273]_ ;
  assign \new_[4282]_  = \new_[4281]_  | \new_[4266]_ ;
  assign \new_[4286]_  = \new_[3612]_  | \new_[3613]_ ;
  assign \new_[4287]_  = \new_[3614]_  | \new_[4286]_ ;
  assign \new_[4290]_  = \new_[3610]_  | \new_[3611]_ ;
  assign \new_[4293]_  = \new_[3608]_  | \new_[3609]_ ;
  assign \new_[4294]_  = \new_[4293]_  | \new_[4290]_ ;
  assign \new_[4295]_  = \new_[4294]_  | \new_[4287]_ ;
  assign \new_[4298]_  = \new_[3606]_  | \new_[3607]_ ;
  assign \new_[4301]_  = \new_[3604]_  | \new_[3605]_ ;
  assign \new_[4302]_  = \new_[4301]_  | \new_[4298]_ ;
  assign \new_[4305]_  = \new_[3602]_  | \new_[3603]_ ;
  assign \new_[4308]_  = \new_[3600]_  | \new_[3601]_ ;
  assign \new_[4309]_  = \new_[4308]_  | \new_[4305]_ ;
  assign \new_[4310]_  = \new_[4309]_  | \new_[4302]_ ;
  assign \new_[4311]_  = \new_[4310]_  | \new_[4295]_ ;
  assign \new_[4312]_  = \new_[4311]_  | \new_[4282]_ ;
  assign \new_[4313]_  = \new_[4312]_  | \new_[4253]_ ;
  assign \new_[4314]_  = \new_[4313]_  | \new_[4194]_ ;
  assign \new_[4315]_  = \new_[4314]_  | \new_[4075]_ ;
  assign \new_[4319]_  = \new_[3597]_  | \new_[3598]_ ;
  assign \new_[4320]_  = \new_[3599]_  | \new_[4319]_ ;
  assign \new_[4323]_  = \new_[3595]_  | \new_[3596]_ ;
  assign \new_[4326]_  = \new_[3593]_  | \new_[3594]_ ;
  assign \new_[4327]_  = \new_[4326]_  | \new_[4323]_ ;
  assign \new_[4328]_  = \new_[4327]_  | \new_[4320]_ ;
  assign \new_[4331]_  = \new_[3591]_  | \new_[3592]_ ;
  assign \new_[4334]_  = \new_[3589]_  | \new_[3590]_ ;
  assign \new_[4335]_  = \new_[4334]_  | \new_[4331]_ ;
  assign \new_[4338]_  = \new_[3587]_  | \new_[3588]_ ;
  assign \new_[4341]_  = \new_[3585]_  | \new_[3586]_ ;
  assign \new_[4342]_  = \new_[4341]_  | \new_[4338]_ ;
  assign \new_[4343]_  = \new_[4342]_  | \new_[4335]_ ;
  assign \new_[4344]_  = \new_[4343]_  | \new_[4328]_ ;
  assign \new_[4348]_  = \new_[3582]_  | \new_[3583]_ ;
  assign \new_[4349]_  = \new_[3584]_  | \new_[4348]_ ;
  assign \new_[4352]_  = \new_[3580]_  | \new_[3581]_ ;
  assign \new_[4355]_  = \new_[3578]_  | \new_[3579]_ ;
  assign \new_[4356]_  = \new_[4355]_  | \new_[4352]_ ;
  assign \new_[4357]_  = \new_[4356]_  | \new_[4349]_ ;
  assign \new_[4360]_  = \new_[3576]_  | \new_[3577]_ ;
  assign \new_[4363]_  = \new_[3574]_  | \new_[3575]_ ;
  assign \new_[4364]_  = \new_[4363]_  | \new_[4360]_ ;
  assign \new_[4367]_  = \new_[3572]_  | \new_[3573]_ ;
  assign \new_[4370]_  = \new_[3570]_  | \new_[3571]_ ;
  assign \new_[4371]_  = \new_[4370]_  | \new_[4367]_ ;
  assign \new_[4372]_  = \new_[4371]_  | \new_[4364]_ ;
  assign \new_[4373]_  = \new_[4372]_  | \new_[4357]_ ;
  assign \new_[4374]_  = \new_[4373]_  | \new_[4344]_ ;
  assign \new_[4378]_  = \new_[3567]_  | \new_[3568]_ ;
  assign \new_[4379]_  = \new_[3569]_  | \new_[4378]_ ;
  assign \new_[4382]_  = \new_[3565]_  | \new_[3566]_ ;
  assign \new_[4385]_  = \new_[3563]_  | \new_[3564]_ ;
  assign \new_[4386]_  = \new_[4385]_  | \new_[4382]_ ;
  assign \new_[4387]_  = \new_[4386]_  | \new_[4379]_ ;
  assign \new_[4390]_  = \new_[3561]_  | \new_[3562]_ ;
  assign \new_[4393]_  = \new_[3559]_  | \new_[3560]_ ;
  assign \new_[4394]_  = \new_[4393]_  | \new_[4390]_ ;
  assign \new_[4397]_  = \new_[3557]_  | \new_[3558]_ ;
  assign \new_[4400]_  = \new_[3555]_  | \new_[3556]_ ;
  assign \new_[4401]_  = \new_[4400]_  | \new_[4397]_ ;
  assign \new_[4402]_  = \new_[4401]_  | \new_[4394]_ ;
  assign \new_[4403]_  = \new_[4402]_  | \new_[4387]_ ;
  assign \new_[4407]_  = \new_[3552]_  | \new_[3553]_ ;
  assign \new_[4408]_  = \new_[3554]_  | \new_[4407]_ ;
  assign \new_[4411]_  = \new_[3550]_  | \new_[3551]_ ;
  assign \new_[4414]_  = \new_[3548]_  | \new_[3549]_ ;
  assign \new_[4415]_  = \new_[4414]_  | \new_[4411]_ ;
  assign \new_[4416]_  = \new_[4415]_  | \new_[4408]_ ;
  assign \new_[4419]_  = \new_[3546]_  | \new_[3547]_ ;
  assign \new_[4422]_  = \new_[3544]_  | \new_[3545]_ ;
  assign \new_[4423]_  = \new_[4422]_  | \new_[4419]_ ;
  assign \new_[4426]_  = \new_[3542]_  | \new_[3543]_ ;
  assign \new_[4429]_  = \new_[3540]_  | \new_[3541]_ ;
  assign \new_[4430]_  = \new_[4429]_  | \new_[4426]_ ;
  assign \new_[4431]_  = \new_[4430]_  | \new_[4423]_ ;
  assign \new_[4432]_  = \new_[4431]_  | \new_[4416]_ ;
  assign \new_[4433]_  = \new_[4432]_  | \new_[4403]_ ;
  assign \new_[4434]_  = \new_[4433]_  | \new_[4374]_ ;
  assign \new_[4438]_  = \new_[3537]_  | \new_[3538]_ ;
  assign \new_[4439]_  = \new_[3539]_  | \new_[4438]_ ;
  assign \new_[4442]_  = \new_[3535]_  | \new_[3536]_ ;
  assign \new_[4445]_  = \new_[3533]_  | \new_[3534]_ ;
  assign \new_[4446]_  = \new_[4445]_  | \new_[4442]_ ;
  assign \new_[4447]_  = \new_[4446]_  | \new_[4439]_ ;
  assign \new_[4450]_  = \new_[3531]_  | \new_[3532]_ ;
  assign \new_[4453]_  = \new_[3529]_  | \new_[3530]_ ;
  assign \new_[4454]_  = \new_[4453]_  | \new_[4450]_ ;
  assign \new_[4457]_  = \new_[3527]_  | \new_[3528]_ ;
  assign \new_[4460]_  = \new_[3525]_  | \new_[3526]_ ;
  assign \new_[4461]_  = \new_[4460]_  | \new_[4457]_ ;
  assign \new_[4462]_  = \new_[4461]_  | \new_[4454]_ ;
  assign \new_[4463]_  = \new_[4462]_  | \new_[4447]_ ;
  assign \new_[4467]_  = \new_[3522]_  | \new_[3523]_ ;
  assign \new_[4468]_  = \new_[3524]_  | \new_[4467]_ ;
  assign \new_[4471]_  = \new_[3520]_  | \new_[3521]_ ;
  assign \new_[4474]_  = \new_[3518]_  | \new_[3519]_ ;
  assign \new_[4475]_  = \new_[4474]_  | \new_[4471]_ ;
  assign \new_[4476]_  = \new_[4475]_  | \new_[4468]_ ;
  assign \new_[4479]_  = \new_[3516]_  | \new_[3517]_ ;
  assign \new_[4482]_  = \new_[3514]_  | \new_[3515]_ ;
  assign \new_[4483]_  = \new_[4482]_  | \new_[4479]_ ;
  assign \new_[4486]_  = \new_[3512]_  | \new_[3513]_ ;
  assign \new_[4489]_  = \new_[3510]_  | \new_[3511]_ ;
  assign \new_[4490]_  = \new_[4489]_  | \new_[4486]_ ;
  assign \new_[4491]_  = \new_[4490]_  | \new_[4483]_ ;
  assign \new_[4492]_  = \new_[4491]_  | \new_[4476]_ ;
  assign \new_[4493]_  = \new_[4492]_  | \new_[4463]_ ;
  assign \new_[4497]_  = \new_[3507]_  | \new_[3508]_ ;
  assign \new_[4498]_  = \new_[3509]_  | \new_[4497]_ ;
  assign \new_[4501]_  = \new_[3505]_  | \new_[3506]_ ;
  assign \new_[4504]_  = \new_[3503]_  | \new_[3504]_ ;
  assign \new_[4505]_  = \new_[4504]_  | \new_[4501]_ ;
  assign \new_[4506]_  = \new_[4505]_  | \new_[4498]_ ;
  assign \new_[4509]_  = \new_[3501]_  | \new_[3502]_ ;
  assign \new_[4512]_  = \new_[3499]_  | \new_[3500]_ ;
  assign \new_[4513]_  = \new_[4512]_  | \new_[4509]_ ;
  assign \new_[4516]_  = \new_[3497]_  | \new_[3498]_ ;
  assign \new_[4519]_  = \new_[3495]_  | \new_[3496]_ ;
  assign \new_[4520]_  = \new_[4519]_  | \new_[4516]_ ;
  assign \new_[4521]_  = \new_[4520]_  | \new_[4513]_ ;
  assign \new_[4522]_  = \new_[4521]_  | \new_[4506]_ ;
  assign \new_[4526]_  = \new_[3492]_  | \new_[3493]_ ;
  assign \new_[4527]_  = \new_[3494]_  | \new_[4526]_ ;
  assign \new_[4530]_  = \new_[3490]_  | \new_[3491]_ ;
  assign \new_[4533]_  = \new_[3488]_  | \new_[3489]_ ;
  assign \new_[4534]_  = \new_[4533]_  | \new_[4530]_ ;
  assign \new_[4535]_  = \new_[4534]_  | \new_[4527]_ ;
  assign \new_[4538]_  = \new_[3486]_  | \new_[3487]_ ;
  assign \new_[4541]_  = \new_[3484]_  | \new_[3485]_ ;
  assign \new_[4542]_  = \new_[4541]_  | \new_[4538]_ ;
  assign \new_[4545]_  = \new_[3482]_  | \new_[3483]_ ;
  assign \new_[4548]_  = \new_[3480]_  | \new_[3481]_ ;
  assign \new_[4549]_  = \new_[4548]_  | \new_[4545]_ ;
  assign \new_[4550]_  = \new_[4549]_  | \new_[4542]_ ;
  assign \new_[4551]_  = \new_[4550]_  | \new_[4535]_ ;
  assign \new_[4552]_  = \new_[4551]_  | \new_[4522]_ ;
  assign \new_[4553]_  = \new_[4552]_  | \new_[4493]_ ;
  assign \new_[4554]_  = \new_[4553]_  | \new_[4434]_ ;
  assign \new_[4558]_  = \new_[3477]_  | \new_[3478]_ ;
  assign \new_[4559]_  = \new_[3479]_  | \new_[4558]_ ;
  assign \new_[4562]_  = \new_[3475]_  | \new_[3476]_ ;
  assign \new_[4565]_  = \new_[3473]_  | \new_[3474]_ ;
  assign \new_[4566]_  = \new_[4565]_  | \new_[4562]_ ;
  assign \new_[4567]_  = \new_[4566]_  | \new_[4559]_ ;
  assign \new_[4570]_  = \new_[3471]_  | \new_[3472]_ ;
  assign \new_[4573]_  = \new_[3469]_  | \new_[3470]_ ;
  assign \new_[4574]_  = \new_[4573]_  | \new_[4570]_ ;
  assign \new_[4577]_  = \new_[3467]_  | \new_[3468]_ ;
  assign \new_[4580]_  = \new_[3465]_  | \new_[3466]_ ;
  assign \new_[4581]_  = \new_[4580]_  | \new_[4577]_ ;
  assign \new_[4582]_  = \new_[4581]_  | \new_[4574]_ ;
  assign \new_[4583]_  = \new_[4582]_  | \new_[4567]_ ;
  assign \new_[4587]_  = \new_[3462]_  | \new_[3463]_ ;
  assign \new_[4588]_  = \new_[3464]_  | \new_[4587]_ ;
  assign \new_[4591]_  = \new_[3460]_  | \new_[3461]_ ;
  assign \new_[4594]_  = \new_[3458]_  | \new_[3459]_ ;
  assign \new_[4595]_  = \new_[4594]_  | \new_[4591]_ ;
  assign \new_[4596]_  = \new_[4595]_  | \new_[4588]_ ;
  assign \new_[4599]_  = \new_[3456]_  | \new_[3457]_ ;
  assign \new_[4602]_  = \new_[3454]_  | \new_[3455]_ ;
  assign \new_[4603]_  = \new_[4602]_  | \new_[4599]_ ;
  assign \new_[4606]_  = \new_[3452]_  | \new_[3453]_ ;
  assign \new_[4609]_  = \new_[3450]_  | \new_[3451]_ ;
  assign \new_[4610]_  = \new_[4609]_  | \new_[4606]_ ;
  assign \new_[4611]_  = \new_[4610]_  | \new_[4603]_ ;
  assign \new_[4612]_  = \new_[4611]_  | \new_[4596]_ ;
  assign \new_[4613]_  = \new_[4612]_  | \new_[4583]_ ;
  assign \new_[4617]_  = \new_[3447]_  | \new_[3448]_ ;
  assign \new_[4618]_  = \new_[3449]_  | \new_[4617]_ ;
  assign \new_[4621]_  = \new_[3445]_  | \new_[3446]_ ;
  assign \new_[4624]_  = \new_[3443]_  | \new_[3444]_ ;
  assign \new_[4625]_  = \new_[4624]_  | \new_[4621]_ ;
  assign \new_[4626]_  = \new_[4625]_  | \new_[4618]_ ;
  assign \new_[4629]_  = \new_[3441]_  | \new_[3442]_ ;
  assign \new_[4632]_  = \new_[3439]_  | \new_[3440]_ ;
  assign \new_[4633]_  = \new_[4632]_  | \new_[4629]_ ;
  assign \new_[4636]_  = \new_[3437]_  | \new_[3438]_ ;
  assign \new_[4639]_  = \new_[3435]_  | \new_[3436]_ ;
  assign \new_[4640]_  = \new_[4639]_  | \new_[4636]_ ;
  assign \new_[4641]_  = \new_[4640]_  | \new_[4633]_ ;
  assign \new_[4642]_  = \new_[4641]_  | \new_[4626]_ ;
  assign \new_[4646]_  = \new_[3432]_  | \new_[3433]_ ;
  assign \new_[4647]_  = \new_[3434]_  | \new_[4646]_ ;
  assign \new_[4650]_  = \new_[3430]_  | \new_[3431]_ ;
  assign \new_[4653]_  = \new_[3428]_  | \new_[3429]_ ;
  assign \new_[4654]_  = \new_[4653]_  | \new_[4650]_ ;
  assign \new_[4655]_  = \new_[4654]_  | \new_[4647]_ ;
  assign \new_[4658]_  = \new_[3426]_  | \new_[3427]_ ;
  assign \new_[4661]_  = \new_[3424]_  | \new_[3425]_ ;
  assign \new_[4662]_  = \new_[4661]_  | \new_[4658]_ ;
  assign \new_[4665]_  = \new_[3422]_  | \new_[3423]_ ;
  assign \new_[4668]_  = \new_[3420]_  | \new_[3421]_ ;
  assign \new_[4669]_  = \new_[4668]_  | \new_[4665]_ ;
  assign \new_[4670]_  = \new_[4669]_  | \new_[4662]_ ;
  assign \new_[4671]_  = \new_[4670]_  | \new_[4655]_ ;
  assign \new_[4672]_  = \new_[4671]_  | \new_[4642]_ ;
  assign \new_[4673]_  = \new_[4672]_  | \new_[4613]_ ;
  assign \new_[4677]_  = \new_[3417]_  | \new_[3418]_ ;
  assign \new_[4678]_  = \new_[3419]_  | \new_[4677]_ ;
  assign \new_[4681]_  = \new_[3415]_  | \new_[3416]_ ;
  assign \new_[4684]_  = \new_[3413]_  | \new_[3414]_ ;
  assign \new_[4685]_  = \new_[4684]_  | \new_[4681]_ ;
  assign \new_[4686]_  = \new_[4685]_  | \new_[4678]_ ;
  assign \new_[4689]_  = \new_[3411]_  | \new_[3412]_ ;
  assign \new_[4692]_  = \new_[3409]_  | \new_[3410]_ ;
  assign \new_[4693]_  = \new_[4692]_  | \new_[4689]_ ;
  assign \new_[4696]_  = \new_[3407]_  | \new_[3408]_ ;
  assign \new_[4699]_  = \new_[3405]_  | \new_[3406]_ ;
  assign \new_[4700]_  = \new_[4699]_  | \new_[4696]_ ;
  assign \new_[4701]_  = \new_[4700]_  | \new_[4693]_ ;
  assign \new_[4702]_  = \new_[4701]_  | \new_[4686]_ ;
  assign \new_[4706]_  = \new_[3402]_  | \new_[3403]_ ;
  assign \new_[4707]_  = \new_[3404]_  | \new_[4706]_ ;
  assign \new_[4710]_  = \new_[3400]_  | \new_[3401]_ ;
  assign \new_[4713]_  = \new_[3398]_  | \new_[3399]_ ;
  assign \new_[4714]_  = \new_[4713]_  | \new_[4710]_ ;
  assign \new_[4715]_  = \new_[4714]_  | \new_[4707]_ ;
  assign \new_[4718]_  = \new_[3396]_  | \new_[3397]_ ;
  assign \new_[4721]_  = \new_[3394]_  | \new_[3395]_ ;
  assign \new_[4722]_  = \new_[4721]_  | \new_[4718]_ ;
  assign \new_[4725]_  = \new_[3392]_  | \new_[3393]_ ;
  assign \new_[4728]_  = \new_[3390]_  | \new_[3391]_ ;
  assign \new_[4729]_  = \new_[4728]_  | \new_[4725]_ ;
  assign \new_[4730]_  = \new_[4729]_  | \new_[4722]_ ;
  assign \new_[4731]_  = \new_[4730]_  | \new_[4715]_ ;
  assign \new_[4732]_  = \new_[4731]_  | \new_[4702]_ ;
  assign \new_[4736]_  = \new_[3387]_  | \new_[3388]_ ;
  assign \new_[4737]_  = \new_[3389]_  | \new_[4736]_ ;
  assign \new_[4740]_  = \new_[3385]_  | \new_[3386]_ ;
  assign \new_[4743]_  = \new_[3383]_  | \new_[3384]_ ;
  assign \new_[4744]_  = \new_[4743]_  | \new_[4740]_ ;
  assign \new_[4745]_  = \new_[4744]_  | \new_[4737]_ ;
  assign \new_[4748]_  = \new_[3381]_  | \new_[3382]_ ;
  assign \new_[4751]_  = \new_[3379]_  | \new_[3380]_ ;
  assign \new_[4752]_  = \new_[4751]_  | \new_[4748]_ ;
  assign \new_[4755]_  = \new_[3377]_  | \new_[3378]_ ;
  assign \new_[4758]_  = \new_[3375]_  | \new_[3376]_ ;
  assign \new_[4759]_  = \new_[4758]_  | \new_[4755]_ ;
  assign \new_[4760]_  = \new_[4759]_  | \new_[4752]_ ;
  assign \new_[4761]_  = \new_[4760]_  | \new_[4745]_ ;
  assign \new_[4765]_  = \new_[3372]_  | \new_[3373]_ ;
  assign \new_[4766]_  = \new_[3374]_  | \new_[4765]_ ;
  assign \new_[4769]_  = \new_[3370]_  | \new_[3371]_ ;
  assign \new_[4772]_  = \new_[3368]_  | \new_[3369]_ ;
  assign \new_[4773]_  = \new_[4772]_  | \new_[4769]_ ;
  assign \new_[4774]_  = \new_[4773]_  | \new_[4766]_ ;
  assign \new_[4777]_  = \new_[3366]_  | \new_[3367]_ ;
  assign \new_[4780]_  = \new_[3364]_  | \new_[3365]_ ;
  assign \new_[4781]_  = \new_[4780]_  | \new_[4777]_ ;
  assign \new_[4784]_  = \new_[3362]_  | \new_[3363]_ ;
  assign \new_[4787]_  = \new_[3360]_  | \new_[3361]_ ;
  assign \new_[4788]_  = \new_[4787]_  | \new_[4784]_ ;
  assign \new_[4789]_  = \new_[4788]_  | \new_[4781]_ ;
  assign \new_[4790]_  = \new_[4789]_  | \new_[4774]_ ;
  assign \new_[4791]_  = \new_[4790]_  | \new_[4761]_ ;
  assign \new_[4792]_  = \new_[4791]_  | \new_[4732]_ ;
  assign \new_[4793]_  = \new_[4792]_  | \new_[4673]_ ;
  assign \new_[4794]_  = \new_[4793]_  | \new_[4554]_ ;
  assign \new_[4795]_  = \new_[4794]_  | \new_[4315]_ ;
  assign \new_[4799]_  = \new_[3357]_  | \new_[3358]_ ;
  assign \new_[4800]_  = \new_[3359]_  | \new_[4799]_ ;
  assign \new_[4803]_  = \new_[3355]_  | \new_[3356]_ ;
  assign \new_[4806]_  = \new_[3353]_  | \new_[3354]_ ;
  assign \new_[4807]_  = \new_[4806]_  | \new_[4803]_ ;
  assign \new_[4808]_  = \new_[4807]_  | \new_[4800]_ ;
  assign \new_[4811]_  = \new_[3351]_  | \new_[3352]_ ;
  assign \new_[4814]_  = \new_[3349]_  | \new_[3350]_ ;
  assign \new_[4815]_  = \new_[4814]_  | \new_[4811]_ ;
  assign \new_[4818]_  = \new_[3347]_  | \new_[3348]_ ;
  assign \new_[4821]_  = \new_[3345]_  | \new_[3346]_ ;
  assign \new_[4822]_  = \new_[4821]_  | \new_[4818]_ ;
  assign \new_[4823]_  = \new_[4822]_  | \new_[4815]_ ;
  assign \new_[4824]_  = \new_[4823]_  | \new_[4808]_ ;
  assign \new_[4828]_  = \new_[3342]_  | \new_[3343]_ ;
  assign \new_[4829]_  = \new_[3344]_  | \new_[4828]_ ;
  assign \new_[4832]_  = \new_[3340]_  | \new_[3341]_ ;
  assign \new_[4835]_  = \new_[3338]_  | \new_[3339]_ ;
  assign \new_[4836]_  = \new_[4835]_  | \new_[4832]_ ;
  assign \new_[4837]_  = \new_[4836]_  | \new_[4829]_ ;
  assign \new_[4840]_  = \new_[3336]_  | \new_[3337]_ ;
  assign \new_[4843]_  = \new_[3334]_  | \new_[3335]_ ;
  assign \new_[4844]_  = \new_[4843]_  | \new_[4840]_ ;
  assign \new_[4847]_  = \new_[3332]_  | \new_[3333]_ ;
  assign \new_[4850]_  = \new_[3330]_  | \new_[3331]_ ;
  assign \new_[4851]_  = \new_[4850]_  | \new_[4847]_ ;
  assign \new_[4852]_  = \new_[4851]_  | \new_[4844]_ ;
  assign \new_[4853]_  = \new_[4852]_  | \new_[4837]_ ;
  assign \new_[4854]_  = \new_[4853]_  | \new_[4824]_ ;
  assign \new_[4858]_  = \new_[3327]_  | \new_[3328]_ ;
  assign \new_[4859]_  = \new_[3329]_  | \new_[4858]_ ;
  assign \new_[4862]_  = \new_[3325]_  | \new_[3326]_ ;
  assign \new_[4865]_  = \new_[3323]_  | \new_[3324]_ ;
  assign \new_[4866]_  = \new_[4865]_  | \new_[4862]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4859]_ ;
  assign \new_[4870]_  = \new_[3321]_  | \new_[3322]_ ;
  assign \new_[4873]_  = \new_[3319]_  | \new_[3320]_ ;
  assign \new_[4874]_  = \new_[4873]_  | \new_[4870]_ ;
  assign \new_[4877]_  = \new_[3317]_  | \new_[3318]_ ;
  assign \new_[4880]_  = \new_[3315]_  | \new_[3316]_ ;
  assign \new_[4881]_  = \new_[4880]_  | \new_[4877]_ ;
  assign \new_[4882]_  = \new_[4881]_  | \new_[4874]_ ;
  assign \new_[4883]_  = \new_[4882]_  | \new_[4867]_ ;
  assign \new_[4887]_  = \new_[3312]_  | \new_[3313]_ ;
  assign \new_[4888]_  = \new_[3314]_  | \new_[4887]_ ;
  assign \new_[4891]_  = \new_[3310]_  | \new_[3311]_ ;
  assign \new_[4894]_  = \new_[3308]_  | \new_[3309]_ ;
  assign \new_[4895]_  = \new_[4894]_  | \new_[4891]_ ;
  assign \new_[4896]_  = \new_[4895]_  | \new_[4888]_ ;
  assign \new_[4899]_  = \new_[3306]_  | \new_[3307]_ ;
  assign \new_[4902]_  = \new_[3304]_  | \new_[3305]_ ;
  assign \new_[4903]_  = \new_[4902]_  | \new_[4899]_ ;
  assign \new_[4906]_  = \new_[3302]_  | \new_[3303]_ ;
  assign \new_[4909]_  = \new_[3300]_  | \new_[3301]_ ;
  assign \new_[4910]_  = \new_[4909]_  | \new_[4906]_ ;
  assign \new_[4911]_  = \new_[4910]_  | \new_[4903]_ ;
  assign \new_[4912]_  = \new_[4911]_  | \new_[4896]_ ;
  assign \new_[4913]_  = \new_[4912]_  | \new_[4883]_ ;
  assign \new_[4914]_  = \new_[4913]_  | \new_[4854]_ ;
  assign \new_[4918]_  = \new_[3297]_  | \new_[3298]_ ;
  assign \new_[4919]_  = \new_[3299]_  | \new_[4918]_ ;
  assign \new_[4922]_  = \new_[3295]_  | \new_[3296]_ ;
  assign \new_[4925]_  = \new_[3293]_  | \new_[3294]_ ;
  assign \new_[4926]_  = \new_[4925]_  | \new_[4922]_ ;
  assign \new_[4927]_  = \new_[4926]_  | \new_[4919]_ ;
  assign \new_[4930]_  = \new_[3291]_  | \new_[3292]_ ;
  assign \new_[4933]_  = \new_[3289]_  | \new_[3290]_ ;
  assign \new_[4934]_  = \new_[4933]_  | \new_[4930]_ ;
  assign \new_[4937]_  = \new_[3287]_  | \new_[3288]_ ;
  assign \new_[4940]_  = \new_[3285]_  | \new_[3286]_ ;
  assign \new_[4941]_  = \new_[4940]_  | \new_[4937]_ ;
  assign \new_[4942]_  = \new_[4941]_  | \new_[4934]_ ;
  assign \new_[4943]_  = \new_[4942]_  | \new_[4927]_ ;
  assign \new_[4947]_  = \new_[3282]_  | \new_[3283]_ ;
  assign \new_[4948]_  = \new_[3284]_  | \new_[4947]_ ;
  assign \new_[4951]_  = \new_[3280]_  | \new_[3281]_ ;
  assign \new_[4954]_  = \new_[3278]_  | \new_[3279]_ ;
  assign \new_[4955]_  = \new_[4954]_  | \new_[4951]_ ;
  assign \new_[4956]_  = \new_[4955]_  | \new_[4948]_ ;
  assign \new_[4959]_  = \new_[3276]_  | \new_[3277]_ ;
  assign \new_[4962]_  = \new_[3274]_  | \new_[3275]_ ;
  assign \new_[4963]_  = \new_[4962]_  | \new_[4959]_ ;
  assign \new_[4966]_  = \new_[3272]_  | \new_[3273]_ ;
  assign \new_[4969]_  = \new_[3270]_  | \new_[3271]_ ;
  assign \new_[4970]_  = \new_[4969]_  | \new_[4966]_ ;
  assign \new_[4971]_  = \new_[4970]_  | \new_[4963]_ ;
  assign \new_[4972]_  = \new_[4971]_  | \new_[4956]_ ;
  assign \new_[4973]_  = \new_[4972]_  | \new_[4943]_ ;
  assign \new_[4977]_  = \new_[3267]_  | \new_[3268]_ ;
  assign \new_[4978]_  = \new_[3269]_  | \new_[4977]_ ;
  assign \new_[4981]_  = \new_[3265]_  | \new_[3266]_ ;
  assign \new_[4984]_  = \new_[3263]_  | \new_[3264]_ ;
  assign \new_[4985]_  = \new_[4984]_  | \new_[4981]_ ;
  assign \new_[4986]_  = \new_[4985]_  | \new_[4978]_ ;
  assign \new_[4989]_  = \new_[3261]_  | \new_[3262]_ ;
  assign \new_[4992]_  = \new_[3259]_  | \new_[3260]_ ;
  assign \new_[4993]_  = \new_[4992]_  | \new_[4989]_ ;
  assign \new_[4996]_  = \new_[3257]_  | \new_[3258]_ ;
  assign \new_[4999]_  = \new_[3255]_  | \new_[3256]_ ;
  assign \new_[5000]_  = \new_[4999]_  | \new_[4996]_ ;
  assign \new_[5001]_  = \new_[5000]_  | \new_[4993]_ ;
  assign \new_[5002]_  = \new_[5001]_  | \new_[4986]_ ;
  assign \new_[5006]_  = \new_[3252]_  | \new_[3253]_ ;
  assign \new_[5007]_  = \new_[3254]_  | \new_[5006]_ ;
  assign \new_[5010]_  = \new_[3250]_  | \new_[3251]_ ;
  assign \new_[5013]_  = \new_[3248]_  | \new_[3249]_ ;
  assign \new_[5014]_  = \new_[5013]_  | \new_[5010]_ ;
  assign \new_[5015]_  = \new_[5014]_  | \new_[5007]_ ;
  assign \new_[5018]_  = \new_[3246]_  | \new_[3247]_ ;
  assign \new_[5021]_  = \new_[3244]_  | \new_[3245]_ ;
  assign \new_[5022]_  = \new_[5021]_  | \new_[5018]_ ;
  assign \new_[5025]_  = \new_[3242]_  | \new_[3243]_ ;
  assign \new_[5028]_  = \new_[3240]_  | \new_[3241]_ ;
  assign \new_[5029]_  = \new_[5028]_  | \new_[5025]_ ;
  assign \new_[5030]_  = \new_[5029]_  | \new_[5022]_ ;
  assign \new_[5031]_  = \new_[5030]_  | \new_[5015]_ ;
  assign \new_[5032]_  = \new_[5031]_  | \new_[5002]_ ;
  assign \new_[5033]_  = \new_[5032]_  | \new_[4973]_ ;
  assign \new_[5034]_  = \new_[5033]_  | \new_[4914]_ ;
  assign \new_[5038]_  = \new_[3237]_  | \new_[3238]_ ;
  assign \new_[5039]_  = \new_[3239]_  | \new_[5038]_ ;
  assign \new_[5042]_  = \new_[3235]_  | \new_[3236]_ ;
  assign \new_[5045]_  = \new_[3233]_  | \new_[3234]_ ;
  assign \new_[5046]_  = \new_[5045]_  | \new_[5042]_ ;
  assign \new_[5047]_  = \new_[5046]_  | \new_[5039]_ ;
  assign \new_[5050]_  = \new_[3231]_  | \new_[3232]_ ;
  assign \new_[5053]_  = \new_[3229]_  | \new_[3230]_ ;
  assign \new_[5054]_  = \new_[5053]_  | \new_[5050]_ ;
  assign \new_[5057]_  = \new_[3227]_  | \new_[3228]_ ;
  assign \new_[5060]_  = \new_[3225]_  | \new_[3226]_ ;
  assign \new_[5061]_  = \new_[5060]_  | \new_[5057]_ ;
  assign \new_[5062]_  = \new_[5061]_  | \new_[5054]_ ;
  assign \new_[5063]_  = \new_[5062]_  | \new_[5047]_ ;
  assign \new_[5067]_  = \new_[3222]_  | \new_[3223]_ ;
  assign \new_[5068]_  = \new_[3224]_  | \new_[5067]_ ;
  assign \new_[5071]_  = \new_[3220]_  | \new_[3221]_ ;
  assign \new_[5074]_  = \new_[3218]_  | \new_[3219]_ ;
  assign \new_[5075]_  = \new_[5074]_  | \new_[5071]_ ;
  assign \new_[5076]_  = \new_[5075]_  | \new_[5068]_ ;
  assign \new_[5079]_  = \new_[3216]_  | \new_[3217]_ ;
  assign \new_[5082]_  = \new_[3214]_  | \new_[3215]_ ;
  assign \new_[5083]_  = \new_[5082]_  | \new_[5079]_ ;
  assign \new_[5086]_  = \new_[3212]_  | \new_[3213]_ ;
  assign \new_[5089]_  = \new_[3210]_  | \new_[3211]_ ;
  assign \new_[5090]_  = \new_[5089]_  | \new_[5086]_ ;
  assign \new_[5091]_  = \new_[5090]_  | \new_[5083]_ ;
  assign \new_[5092]_  = \new_[5091]_  | \new_[5076]_ ;
  assign \new_[5093]_  = \new_[5092]_  | \new_[5063]_ ;
  assign \new_[5097]_  = \new_[3207]_  | \new_[3208]_ ;
  assign \new_[5098]_  = \new_[3209]_  | \new_[5097]_ ;
  assign \new_[5101]_  = \new_[3205]_  | \new_[3206]_ ;
  assign \new_[5104]_  = \new_[3203]_  | \new_[3204]_ ;
  assign \new_[5105]_  = \new_[5104]_  | \new_[5101]_ ;
  assign \new_[5106]_  = \new_[5105]_  | \new_[5098]_ ;
  assign \new_[5109]_  = \new_[3201]_  | \new_[3202]_ ;
  assign \new_[5112]_  = \new_[3199]_  | \new_[3200]_ ;
  assign \new_[5113]_  = \new_[5112]_  | \new_[5109]_ ;
  assign \new_[5116]_  = \new_[3197]_  | \new_[3198]_ ;
  assign \new_[5119]_  = \new_[3195]_  | \new_[3196]_ ;
  assign \new_[5120]_  = \new_[5119]_  | \new_[5116]_ ;
  assign \new_[5121]_  = \new_[5120]_  | \new_[5113]_ ;
  assign \new_[5122]_  = \new_[5121]_  | \new_[5106]_ ;
  assign \new_[5126]_  = \new_[3192]_  | \new_[3193]_ ;
  assign \new_[5127]_  = \new_[3194]_  | \new_[5126]_ ;
  assign \new_[5130]_  = \new_[3190]_  | \new_[3191]_ ;
  assign \new_[5133]_  = \new_[3188]_  | \new_[3189]_ ;
  assign \new_[5134]_  = \new_[5133]_  | \new_[5130]_ ;
  assign \new_[5135]_  = \new_[5134]_  | \new_[5127]_ ;
  assign \new_[5138]_  = \new_[3186]_  | \new_[3187]_ ;
  assign \new_[5141]_  = \new_[3184]_  | \new_[3185]_ ;
  assign \new_[5142]_  = \new_[5141]_  | \new_[5138]_ ;
  assign \new_[5145]_  = \new_[3182]_  | \new_[3183]_ ;
  assign \new_[5148]_  = \new_[3180]_  | \new_[3181]_ ;
  assign \new_[5149]_  = \new_[5148]_  | \new_[5145]_ ;
  assign \new_[5150]_  = \new_[5149]_  | \new_[5142]_ ;
  assign \new_[5151]_  = \new_[5150]_  | \new_[5135]_ ;
  assign \new_[5152]_  = \new_[5151]_  | \new_[5122]_ ;
  assign \new_[5153]_  = \new_[5152]_  | \new_[5093]_ ;
  assign \new_[5157]_  = \new_[3177]_  | \new_[3178]_ ;
  assign \new_[5158]_  = \new_[3179]_  | \new_[5157]_ ;
  assign \new_[5161]_  = \new_[3175]_  | \new_[3176]_ ;
  assign \new_[5164]_  = \new_[3173]_  | \new_[3174]_ ;
  assign \new_[5165]_  = \new_[5164]_  | \new_[5161]_ ;
  assign \new_[5166]_  = \new_[5165]_  | \new_[5158]_ ;
  assign \new_[5169]_  = \new_[3171]_  | \new_[3172]_ ;
  assign \new_[5172]_  = \new_[3169]_  | \new_[3170]_ ;
  assign \new_[5173]_  = \new_[5172]_  | \new_[5169]_ ;
  assign \new_[5176]_  = \new_[3167]_  | \new_[3168]_ ;
  assign \new_[5179]_  = \new_[3165]_  | \new_[3166]_ ;
  assign \new_[5180]_  = \new_[5179]_  | \new_[5176]_ ;
  assign \new_[5181]_  = \new_[5180]_  | \new_[5173]_ ;
  assign \new_[5182]_  = \new_[5181]_  | \new_[5166]_ ;
  assign \new_[5186]_  = \new_[3162]_  | \new_[3163]_ ;
  assign \new_[5187]_  = \new_[3164]_  | \new_[5186]_ ;
  assign \new_[5190]_  = \new_[3160]_  | \new_[3161]_ ;
  assign \new_[5193]_  = \new_[3158]_  | \new_[3159]_ ;
  assign \new_[5194]_  = \new_[5193]_  | \new_[5190]_ ;
  assign \new_[5195]_  = \new_[5194]_  | \new_[5187]_ ;
  assign \new_[5198]_  = \new_[3156]_  | \new_[3157]_ ;
  assign \new_[5201]_  = \new_[3154]_  | \new_[3155]_ ;
  assign \new_[5202]_  = \new_[5201]_  | \new_[5198]_ ;
  assign \new_[5205]_  = \new_[3152]_  | \new_[3153]_ ;
  assign \new_[5208]_  = \new_[3150]_  | \new_[3151]_ ;
  assign \new_[5209]_  = \new_[5208]_  | \new_[5205]_ ;
  assign \new_[5210]_  = \new_[5209]_  | \new_[5202]_ ;
  assign \new_[5211]_  = \new_[5210]_  | \new_[5195]_ ;
  assign \new_[5212]_  = \new_[5211]_  | \new_[5182]_ ;
  assign \new_[5216]_  = \new_[3147]_  | \new_[3148]_ ;
  assign \new_[5217]_  = \new_[3149]_  | \new_[5216]_ ;
  assign \new_[5220]_  = \new_[3145]_  | \new_[3146]_ ;
  assign \new_[5223]_  = \new_[3143]_  | \new_[3144]_ ;
  assign \new_[5224]_  = \new_[5223]_  | \new_[5220]_ ;
  assign \new_[5225]_  = \new_[5224]_  | \new_[5217]_ ;
  assign \new_[5228]_  = \new_[3141]_  | \new_[3142]_ ;
  assign \new_[5231]_  = \new_[3139]_  | \new_[3140]_ ;
  assign \new_[5232]_  = \new_[5231]_  | \new_[5228]_ ;
  assign \new_[5235]_  = \new_[3137]_  | \new_[3138]_ ;
  assign \new_[5238]_  = \new_[3135]_  | \new_[3136]_ ;
  assign \new_[5239]_  = \new_[5238]_  | \new_[5235]_ ;
  assign \new_[5240]_  = \new_[5239]_  | \new_[5232]_ ;
  assign \new_[5241]_  = \new_[5240]_  | \new_[5225]_ ;
  assign \new_[5245]_  = \new_[3132]_  | \new_[3133]_ ;
  assign \new_[5246]_  = \new_[3134]_  | \new_[5245]_ ;
  assign \new_[5249]_  = \new_[3130]_  | \new_[3131]_ ;
  assign \new_[5252]_  = \new_[3128]_  | \new_[3129]_ ;
  assign \new_[5253]_  = \new_[5252]_  | \new_[5249]_ ;
  assign \new_[5254]_  = \new_[5253]_  | \new_[5246]_ ;
  assign \new_[5257]_  = \new_[3126]_  | \new_[3127]_ ;
  assign \new_[5260]_  = \new_[3124]_  | \new_[3125]_ ;
  assign \new_[5261]_  = \new_[5260]_  | \new_[5257]_ ;
  assign \new_[5264]_  = \new_[3122]_  | \new_[3123]_ ;
  assign \new_[5267]_  = \new_[3120]_  | \new_[3121]_ ;
  assign \new_[5268]_  = \new_[5267]_  | \new_[5264]_ ;
  assign \new_[5269]_  = \new_[5268]_  | \new_[5261]_ ;
  assign \new_[5270]_  = \new_[5269]_  | \new_[5254]_ ;
  assign \new_[5271]_  = \new_[5270]_  | \new_[5241]_ ;
  assign \new_[5272]_  = \new_[5271]_  | \new_[5212]_ ;
  assign \new_[5273]_  = \new_[5272]_  | \new_[5153]_ ;
  assign \new_[5274]_  = \new_[5273]_  | \new_[5034]_ ;
  assign \new_[5278]_  = \new_[3117]_  | \new_[3118]_ ;
  assign \new_[5279]_  = \new_[3119]_  | \new_[5278]_ ;
  assign \new_[5282]_  = \new_[3115]_  | \new_[3116]_ ;
  assign \new_[5285]_  = \new_[3113]_  | \new_[3114]_ ;
  assign \new_[5286]_  = \new_[5285]_  | \new_[5282]_ ;
  assign \new_[5287]_  = \new_[5286]_  | \new_[5279]_ ;
  assign \new_[5290]_  = \new_[3111]_  | \new_[3112]_ ;
  assign \new_[5293]_  = \new_[3109]_  | \new_[3110]_ ;
  assign \new_[5294]_  = \new_[5293]_  | \new_[5290]_ ;
  assign \new_[5297]_  = \new_[3107]_  | \new_[3108]_ ;
  assign \new_[5300]_  = \new_[3105]_  | \new_[3106]_ ;
  assign \new_[5301]_  = \new_[5300]_  | \new_[5297]_ ;
  assign \new_[5302]_  = \new_[5301]_  | \new_[5294]_ ;
  assign \new_[5303]_  = \new_[5302]_  | \new_[5287]_ ;
  assign \new_[5307]_  = \new_[3102]_  | \new_[3103]_ ;
  assign \new_[5308]_  = \new_[3104]_  | \new_[5307]_ ;
  assign \new_[5311]_  = \new_[3100]_  | \new_[3101]_ ;
  assign \new_[5314]_  = \new_[3098]_  | \new_[3099]_ ;
  assign \new_[5315]_  = \new_[5314]_  | \new_[5311]_ ;
  assign \new_[5316]_  = \new_[5315]_  | \new_[5308]_ ;
  assign \new_[5319]_  = \new_[3096]_  | \new_[3097]_ ;
  assign \new_[5322]_  = \new_[3094]_  | \new_[3095]_ ;
  assign \new_[5323]_  = \new_[5322]_  | \new_[5319]_ ;
  assign \new_[5326]_  = \new_[3092]_  | \new_[3093]_ ;
  assign \new_[5329]_  = \new_[3090]_  | \new_[3091]_ ;
  assign \new_[5330]_  = \new_[5329]_  | \new_[5326]_ ;
  assign \new_[5331]_  = \new_[5330]_  | \new_[5323]_ ;
  assign \new_[5332]_  = \new_[5331]_  | \new_[5316]_ ;
  assign \new_[5333]_  = \new_[5332]_  | \new_[5303]_ ;
  assign \new_[5337]_  = \new_[3087]_  | \new_[3088]_ ;
  assign \new_[5338]_  = \new_[3089]_  | \new_[5337]_ ;
  assign \new_[5341]_  = \new_[3085]_  | \new_[3086]_ ;
  assign \new_[5344]_  = \new_[3083]_  | \new_[3084]_ ;
  assign \new_[5345]_  = \new_[5344]_  | \new_[5341]_ ;
  assign \new_[5346]_  = \new_[5345]_  | \new_[5338]_ ;
  assign \new_[5349]_  = \new_[3081]_  | \new_[3082]_ ;
  assign \new_[5352]_  = \new_[3079]_  | \new_[3080]_ ;
  assign \new_[5353]_  = \new_[5352]_  | \new_[5349]_ ;
  assign \new_[5356]_  = \new_[3077]_  | \new_[3078]_ ;
  assign \new_[5359]_  = \new_[3075]_  | \new_[3076]_ ;
  assign \new_[5360]_  = \new_[5359]_  | \new_[5356]_ ;
  assign \new_[5361]_  = \new_[5360]_  | \new_[5353]_ ;
  assign \new_[5362]_  = \new_[5361]_  | \new_[5346]_ ;
  assign \new_[5366]_  = \new_[3072]_  | \new_[3073]_ ;
  assign \new_[5367]_  = \new_[3074]_  | \new_[5366]_ ;
  assign \new_[5370]_  = \new_[3070]_  | \new_[3071]_ ;
  assign \new_[5373]_  = \new_[3068]_  | \new_[3069]_ ;
  assign \new_[5374]_  = \new_[5373]_  | \new_[5370]_ ;
  assign \new_[5375]_  = \new_[5374]_  | \new_[5367]_ ;
  assign \new_[5378]_  = \new_[3066]_  | \new_[3067]_ ;
  assign \new_[5381]_  = \new_[3064]_  | \new_[3065]_ ;
  assign \new_[5382]_  = \new_[5381]_  | \new_[5378]_ ;
  assign \new_[5385]_  = \new_[3062]_  | \new_[3063]_ ;
  assign \new_[5388]_  = \new_[3060]_  | \new_[3061]_ ;
  assign \new_[5389]_  = \new_[5388]_  | \new_[5385]_ ;
  assign \new_[5390]_  = \new_[5389]_  | \new_[5382]_ ;
  assign \new_[5391]_  = \new_[5390]_  | \new_[5375]_ ;
  assign \new_[5392]_  = \new_[5391]_  | \new_[5362]_ ;
  assign \new_[5393]_  = \new_[5392]_  | \new_[5333]_ ;
  assign \new_[5397]_  = \new_[3057]_  | \new_[3058]_ ;
  assign \new_[5398]_  = \new_[3059]_  | \new_[5397]_ ;
  assign \new_[5401]_  = \new_[3055]_  | \new_[3056]_ ;
  assign \new_[5404]_  = \new_[3053]_  | \new_[3054]_ ;
  assign \new_[5405]_  = \new_[5404]_  | \new_[5401]_ ;
  assign \new_[5406]_  = \new_[5405]_  | \new_[5398]_ ;
  assign \new_[5409]_  = \new_[3051]_  | \new_[3052]_ ;
  assign \new_[5412]_  = \new_[3049]_  | \new_[3050]_ ;
  assign \new_[5413]_  = \new_[5412]_  | \new_[5409]_ ;
  assign \new_[5416]_  = \new_[3047]_  | \new_[3048]_ ;
  assign \new_[5419]_  = \new_[3045]_  | \new_[3046]_ ;
  assign \new_[5420]_  = \new_[5419]_  | \new_[5416]_ ;
  assign \new_[5421]_  = \new_[5420]_  | \new_[5413]_ ;
  assign \new_[5422]_  = \new_[5421]_  | \new_[5406]_ ;
  assign \new_[5426]_  = \new_[3042]_  | \new_[3043]_ ;
  assign \new_[5427]_  = \new_[3044]_  | \new_[5426]_ ;
  assign \new_[5430]_  = \new_[3040]_  | \new_[3041]_ ;
  assign \new_[5433]_  = \new_[3038]_  | \new_[3039]_ ;
  assign \new_[5434]_  = \new_[5433]_  | \new_[5430]_ ;
  assign \new_[5435]_  = \new_[5434]_  | \new_[5427]_ ;
  assign \new_[5438]_  = \new_[3036]_  | \new_[3037]_ ;
  assign \new_[5441]_  = \new_[3034]_  | \new_[3035]_ ;
  assign \new_[5442]_  = \new_[5441]_  | \new_[5438]_ ;
  assign \new_[5445]_  = \new_[3032]_  | \new_[3033]_ ;
  assign \new_[5448]_  = \new_[3030]_  | \new_[3031]_ ;
  assign \new_[5449]_  = \new_[5448]_  | \new_[5445]_ ;
  assign \new_[5450]_  = \new_[5449]_  | \new_[5442]_ ;
  assign \new_[5451]_  = \new_[5450]_  | \new_[5435]_ ;
  assign \new_[5452]_  = \new_[5451]_  | \new_[5422]_ ;
  assign \new_[5456]_  = \new_[3027]_  | \new_[3028]_ ;
  assign \new_[5457]_  = \new_[3029]_  | \new_[5456]_ ;
  assign \new_[5460]_  = \new_[3025]_  | \new_[3026]_ ;
  assign \new_[5463]_  = \new_[3023]_  | \new_[3024]_ ;
  assign \new_[5464]_  = \new_[5463]_  | \new_[5460]_ ;
  assign \new_[5465]_  = \new_[5464]_  | \new_[5457]_ ;
  assign \new_[5468]_  = \new_[3021]_  | \new_[3022]_ ;
  assign \new_[5471]_  = \new_[3019]_  | \new_[3020]_ ;
  assign \new_[5472]_  = \new_[5471]_  | \new_[5468]_ ;
  assign \new_[5475]_  = \new_[3017]_  | \new_[3018]_ ;
  assign \new_[5478]_  = \new_[3015]_  | \new_[3016]_ ;
  assign \new_[5479]_  = \new_[5478]_  | \new_[5475]_ ;
  assign \new_[5480]_  = \new_[5479]_  | \new_[5472]_ ;
  assign \new_[5481]_  = \new_[5480]_  | \new_[5465]_ ;
  assign \new_[5485]_  = \new_[3012]_  | \new_[3013]_ ;
  assign \new_[5486]_  = \new_[3014]_  | \new_[5485]_ ;
  assign \new_[5489]_  = \new_[3010]_  | \new_[3011]_ ;
  assign \new_[5492]_  = \new_[3008]_  | \new_[3009]_ ;
  assign \new_[5493]_  = \new_[5492]_  | \new_[5489]_ ;
  assign \new_[5494]_  = \new_[5493]_  | \new_[5486]_ ;
  assign \new_[5497]_  = \new_[3006]_  | \new_[3007]_ ;
  assign \new_[5500]_  = \new_[3004]_  | \new_[3005]_ ;
  assign \new_[5501]_  = \new_[5500]_  | \new_[5497]_ ;
  assign \new_[5504]_  = \new_[3002]_  | \new_[3003]_ ;
  assign \new_[5507]_  = \new_[3000]_  | \new_[3001]_ ;
  assign \new_[5508]_  = \new_[5507]_  | \new_[5504]_ ;
  assign \new_[5509]_  = \new_[5508]_  | \new_[5501]_ ;
  assign \new_[5510]_  = \new_[5509]_  | \new_[5494]_ ;
  assign \new_[5511]_  = \new_[5510]_  | \new_[5481]_ ;
  assign \new_[5512]_  = \new_[5511]_  | \new_[5452]_ ;
  assign \new_[5513]_  = \new_[5512]_  | \new_[5393]_ ;
  assign \new_[5517]_  = \new_[2997]_  | \new_[2998]_ ;
  assign \new_[5518]_  = \new_[2999]_  | \new_[5517]_ ;
  assign \new_[5521]_  = \new_[2995]_  | \new_[2996]_ ;
  assign \new_[5524]_  = \new_[2993]_  | \new_[2994]_ ;
  assign \new_[5525]_  = \new_[5524]_  | \new_[5521]_ ;
  assign \new_[5526]_  = \new_[5525]_  | \new_[5518]_ ;
  assign \new_[5529]_  = \new_[2991]_  | \new_[2992]_ ;
  assign \new_[5532]_  = \new_[2989]_  | \new_[2990]_ ;
  assign \new_[5533]_  = \new_[5532]_  | \new_[5529]_ ;
  assign \new_[5536]_  = \new_[2987]_  | \new_[2988]_ ;
  assign \new_[5539]_  = \new_[2985]_  | \new_[2986]_ ;
  assign \new_[5540]_  = \new_[5539]_  | \new_[5536]_ ;
  assign \new_[5541]_  = \new_[5540]_  | \new_[5533]_ ;
  assign \new_[5542]_  = \new_[5541]_  | \new_[5526]_ ;
  assign \new_[5546]_  = \new_[2982]_  | \new_[2983]_ ;
  assign \new_[5547]_  = \new_[2984]_  | \new_[5546]_ ;
  assign \new_[5550]_  = \new_[2980]_  | \new_[2981]_ ;
  assign \new_[5553]_  = \new_[2978]_  | \new_[2979]_ ;
  assign \new_[5554]_  = \new_[5553]_  | \new_[5550]_ ;
  assign \new_[5555]_  = \new_[5554]_  | \new_[5547]_ ;
  assign \new_[5558]_  = \new_[2976]_  | \new_[2977]_ ;
  assign \new_[5561]_  = \new_[2974]_  | \new_[2975]_ ;
  assign \new_[5562]_  = \new_[5561]_  | \new_[5558]_ ;
  assign \new_[5565]_  = \new_[2972]_  | \new_[2973]_ ;
  assign \new_[5568]_  = \new_[2970]_  | \new_[2971]_ ;
  assign \new_[5569]_  = \new_[5568]_  | \new_[5565]_ ;
  assign \new_[5570]_  = \new_[5569]_  | \new_[5562]_ ;
  assign \new_[5571]_  = \new_[5570]_  | \new_[5555]_ ;
  assign \new_[5572]_  = \new_[5571]_  | \new_[5542]_ ;
  assign \new_[5576]_  = \new_[2967]_  | \new_[2968]_ ;
  assign \new_[5577]_  = \new_[2969]_  | \new_[5576]_ ;
  assign \new_[5580]_  = \new_[2965]_  | \new_[2966]_ ;
  assign \new_[5583]_  = \new_[2963]_  | \new_[2964]_ ;
  assign \new_[5584]_  = \new_[5583]_  | \new_[5580]_ ;
  assign \new_[5585]_  = \new_[5584]_  | \new_[5577]_ ;
  assign \new_[5588]_  = \new_[2961]_  | \new_[2962]_ ;
  assign \new_[5591]_  = \new_[2959]_  | \new_[2960]_ ;
  assign \new_[5592]_  = \new_[5591]_  | \new_[5588]_ ;
  assign \new_[5595]_  = \new_[2957]_  | \new_[2958]_ ;
  assign \new_[5598]_  = \new_[2955]_  | \new_[2956]_ ;
  assign \new_[5599]_  = \new_[5598]_  | \new_[5595]_ ;
  assign \new_[5600]_  = \new_[5599]_  | \new_[5592]_ ;
  assign \new_[5601]_  = \new_[5600]_  | \new_[5585]_ ;
  assign \new_[5605]_  = \new_[2952]_  | \new_[2953]_ ;
  assign \new_[5606]_  = \new_[2954]_  | \new_[5605]_ ;
  assign \new_[5609]_  = \new_[2950]_  | \new_[2951]_ ;
  assign \new_[5612]_  = \new_[2948]_  | \new_[2949]_ ;
  assign \new_[5613]_  = \new_[5612]_  | \new_[5609]_ ;
  assign \new_[5614]_  = \new_[5613]_  | \new_[5606]_ ;
  assign \new_[5617]_  = \new_[2946]_  | \new_[2947]_ ;
  assign \new_[5620]_  = \new_[2944]_  | \new_[2945]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5617]_ ;
  assign \new_[5624]_  = \new_[2942]_  | \new_[2943]_ ;
  assign \new_[5627]_  = \new_[2940]_  | \new_[2941]_ ;
  assign \new_[5628]_  = \new_[5627]_  | \new_[5624]_ ;
  assign \new_[5629]_  = \new_[5628]_  | \new_[5621]_ ;
  assign \new_[5630]_  = \new_[5629]_  | \new_[5614]_ ;
  assign \new_[5631]_  = \new_[5630]_  | \new_[5601]_ ;
  assign \new_[5632]_  = \new_[5631]_  | \new_[5572]_ ;
  assign \new_[5636]_  = \new_[2937]_  | \new_[2938]_ ;
  assign \new_[5637]_  = \new_[2939]_  | \new_[5636]_ ;
  assign \new_[5640]_  = \new_[2935]_  | \new_[2936]_ ;
  assign \new_[5643]_  = \new_[2933]_  | \new_[2934]_ ;
  assign \new_[5644]_  = \new_[5643]_  | \new_[5640]_ ;
  assign \new_[5645]_  = \new_[5644]_  | \new_[5637]_ ;
  assign \new_[5648]_  = \new_[2931]_  | \new_[2932]_ ;
  assign \new_[5651]_  = \new_[2929]_  | \new_[2930]_ ;
  assign \new_[5652]_  = \new_[5651]_  | \new_[5648]_ ;
  assign \new_[5655]_  = \new_[2927]_  | \new_[2928]_ ;
  assign \new_[5658]_  = \new_[2925]_  | \new_[2926]_ ;
  assign \new_[5659]_  = \new_[5658]_  | \new_[5655]_ ;
  assign \new_[5660]_  = \new_[5659]_  | \new_[5652]_ ;
  assign \new_[5661]_  = \new_[5660]_  | \new_[5645]_ ;
  assign \new_[5665]_  = \new_[2922]_  | \new_[2923]_ ;
  assign \new_[5666]_  = \new_[2924]_  | \new_[5665]_ ;
  assign \new_[5669]_  = \new_[2920]_  | \new_[2921]_ ;
  assign \new_[5672]_  = \new_[2918]_  | \new_[2919]_ ;
  assign \new_[5673]_  = \new_[5672]_  | \new_[5669]_ ;
  assign \new_[5674]_  = \new_[5673]_  | \new_[5666]_ ;
  assign \new_[5677]_  = \new_[2916]_  | \new_[2917]_ ;
  assign \new_[5680]_  = \new_[2914]_  | \new_[2915]_ ;
  assign \new_[5681]_  = \new_[5680]_  | \new_[5677]_ ;
  assign \new_[5684]_  = \new_[2912]_  | \new_[2913]_ ;
  assign \new_[5687]_  = \new_[2910]_  | \new_[2911]_ ;
  assign \new_[5688]_  = \new_[5687]_  | \new_[5684]_ ;
  assign \new_[5689]_  = \new_[5688]_  | \new_[5681]_ ;
  assign \new_[5690]_  = \new_[5689]_  | \new_[5674]_ ;
  assign \new_[5691]_  = \new_[5690]_  | \new_[5661]_ ;
  assign \new_[5695]_  = \new_[2907]_  | \new_[2908]_ ;
  assign \new_[5696]_  = \new_[2909]_  | \new_[5695]_ ;
  assign \new_[5699]_  = \new_[2905]_  | \new_[2906]_ ;
  assign \new_[5702]_  = \new_[2903]_  | \new_[2904]_ ;
  assign \new_[5703]_  = \new_[5702]_  | \new_[5699]_ ;
  assign \new_[5704]_  = \new_[5703]_  | \new_[5696]_ ;
  assign \new_[5707]_  = \new_[2901]_  | \new_[2902]_ ;
  assign \new_[5710]_  = \new_[2899]_  | \new_[2900]_ ;
  assign \new_[5711]_  = \new_[5710]_  | \new_[5707]_ ;
  assign \new_[5714]_  = \new_[2897]_  | \new_[2898]_ ;
  assign \new_[5717]_  = \new_[2895]_  | \new_[2896]_ ;
  assign \new_[5718]_  = \new_[5717]_  | \new_[5714]_ ;
  assign \new_[5719]_  = \new_[5718]_  | \new_[5711]_ ;
  assign \new_[5720]_  = \new_[5719]_  | \new_[5704]_ ;
  assign \new_[5724]_  = \new_[2892]_  | \new_[2893]_ ;
  assign \new_[5725]_  = \new_[2894]_  | \new_[5724]_ ;
  assign \new_[5728]_  = \new_[2890]_  | \new_[2891]_ ;
  assign \new_[5731]_  = \new_[2888]_  | \new_[2889]_ ;
  assign \new_[5732]_  = \new_[5731]_  | \new_[5728]_ ;
  assign \new_[5733]_  = \new_[5732]_  | \new_[5725]_ ;
  assign \new_[5736]_  = \new_[2886]_  | \new_[2887]_ ;
  assign \new_[5739]_  = \new_[2884]_  | \new_[2885]_ ;
  assign \new_[5740]_  = \new_[5739]_  | \new_[5736]_ ;
  assign \new_[5743]_  = \new_[2882]_  | \new_[2883]_ ;
  assign \new_[5746]_  = \new_[2880]_  | \new_[2881]_ ;
  assign \new_[5747]_  = \new_[5746]_  | \new_[5743]_ ;
  assign \new_[5748]_  = \new_[5747]_  | \new_[5740]_ ;
  assign \new_[5749]_  = \new_[5748]_  | \new_[5733]_ ;
  assign \new_[5750]_  = \new_[5749]_  | \new_[5720]_ ;
  assign \new_[5751]_  = \new_[5750]_  | \new_[5691]_ ;
  assign \new_[5752]_  = \new_[5751]_  | \new_[5632]_ ;
  assign \new_[5753]_  = \new_[5752]_  | \new_[5513]_ ;
  assign \new_[5754]_  = \new_[5753]_  | \new_[5274]_ ;
  assign \new_[5755]_  = \new_[5754]_  | \new_[4795]_ ;
  assign \new_[5759]_  = \new_[2877]_  | \new_[2878]_ ;
  assign \new_[5760]_  = \new_[2879]_  | \new_[5759]_ ;
  assign \new_[5763]_  = \new_[2875]_  | \new_[2876]_ ;
  assign \new_[5766]_  = \new_[2873]_  | \new_[2874]_ ;
  assign \new_[5767]_  = \new_[5766]_  | \new_[5763]_ ;
  assign \new_[5768]_  = \new_[5767]_  | \new_[5760]_ ;
  assign \new_[5771]_  = \new_[2871]_  | \new_[2872]_ ;
  assign \new_[5774]_  = \new_[2869]_  | \new_[2870]_ ;
  assign \new_[5775]_  = \new_[5774]_  | \new_[5771]_ ;
  assign \new_[5778]_  = \new_[2867]_  | \new_[2868]_ ;
  assign \new_[5781]_  = \new_[2865]_  | \new_[2866]_ ;
  assign \new_[5782]_  = \new_[5781]_  | \new_[5778]_ ;
  assign \new_[5783]_  = \new_[5782]_  | \new_[5775]_ ;
  assign \new_[5784]_  = \new_[5783]_  | \new_[5768]_ ;
  assign \new_[5788]_  = \new_[2862]_  | \new_[2863]_ ;
  assign \new_[5789]_  = \new_[2864]_  | \new_[5788]_ ;
  assign \new_[5792]_  = \new_[2860]_  | \new_[2861]_ ;
  assign \new_[5795]_  = \new_[2858]_  | \new_[2859]_ ;
  assign \new_[5796]_  = \new_[5795]_  | \new_[5792]_ ;
  assign \new_[5797]_  = \new_[5796]_  | \new_[5789]_ ;
  assign \new_[5800]_  = \new_[2856]_  | \new_[2857]_ ;
  assign \new_[5803]_  = \new_[2854]_  | \new_[2855]_ ;
  assign \new_[5804]_  = \new_[5803]_  | \new_[5800]_ ;
  assign \new_[5807]_  = \new_[2852]_  | \new_[2853]_ ;
  assign \new_[5810]_  = \new_[2850]_  | \new_[2851]_ ;
  assign \new_[5811]_  = \new_[5810]_  | \new_[5807]_ ;
  assign \new_[5812]_  = \new_[5811]_  | \new_[5804]_ ;
  assign \new_[5813]_  = \new_[5812]_  | \new_[5797]_ ;
  assign \new_[5814]_  = \new_[5813]_  | \new_[5784]_ ;
  assign \new_[5818]_  = \new_[2847]_  | \new_[2848]_ ;
  assign \new_[5819]_  = \new_[2849]_  | \new_[5818]_ ;
  assign \new_[5822]_  = \new_[2845]_  | \new_[2846]_ ;
  assign \new_[5825]_  = \new_[2843]_  | \new_[2844]_ ;
  assign \new_[5826]_  = \new_[5825]_  | \new_[5822]_ ;
  assign \new_[5827]_  = \new_[5826]_  | \new_[5819]_ ;
  assign \new_[5830]_  = \new_[2841]_  | \new_[2842]_ ;
  assign \new_[5833]_  = \new_[2839]_  | \new_[2840]_ ;
  assign \new_[5834]_  = \new_[5833]_  | \new_[5830]_ ;
  assign \new_[5837]_  = \new_[2837]_  | \new_[2838]_ ;
  assign \new_[5840]_  = \new_[2835]_  | \new_[2836]_ ;
  assign \new_[5841]_  = \new_[5840]_  | \new_[5837]_ ;
  assign \new_[5842]_  = \new_[5841]_  | \new_[5834]_ ;
  assign \new_[5843]_  = \new_[5842]_  | \new_[5827]_ ;
  assign \new_[5847]_  = \new_[2832]_  | \new_[2833]_ ;
  assign \new_[5848]_  = \new_[2834]_  | \new_[5847]_ ;
  assign \new_[5851]_  = \new_[2830]_  | \new_[2831]_ ;
  assign \new_[5854]_  = \new_[2828]_  | \new_[2829]_ ;
  assign \new_[5855]_  = \new_[5854]_  | \new_[5851]_ ;
  assign \new_[5856]_  = \new_[5855]_  | \new_[5848]_ ;
  assign \new_[5859]_  = \new_[2826]_  | \new_[2827]_ ;
  assign \new_[5862]_  = \new_[2824]_  | \new_[2825]_ ;
  assign \new_[5863]_  = \new_[5862]_  | \new_[5859]_ ;
  assign \new_[5866]_  = \new_[2822]_  | \new_[2823]_ ;
  assign \new_[5869]_  = \new_[2820]_  | \new_[2821]_ ;
  assign \new_[5870]_  = \new_[5869]_  | \new_[5866]_ ;
  assign \new_[5871]_  = \new_[5870]_  | \new_[5863]_ ;
  assign \new_[5872]_  = \new_[5871]_  | \new_[5856]_ ;
  assign \new_[5873]_  = \new_[5872]_  | \new_[5843]_ ;
  assign \new_[5874]_  = \new_[5873]_  | \new_[5814]_ ;
  assign \new_[5878]_  = \new_[2817]_  | \new_[2818]_ ;
  assign \new_[5879]_  = \new_[2819]_  | \new_[5878]_ ;
  assign \new_[5882]_  = \new_[2815]_  | \new_[2816]_ ;
  assign \new_[5885]_  = \new_[2813]_  | \new_[2814]_ ;
  assign \new_[5886]_  = \new_[5885]_  | \new_[5882]_ ;
  assign \new_[5887]_  = \new_[5886]_  | \new_[5879]_ ;
  assign \new_[5890]_  = \new_[2811]_  | \new_[2812]_ ;
  assign \new_[5893]_  = \new_[2809]_  | \new_[2810]_ ;
  assign \new_[5894]_  = \new_[5893]_  | \new_[5890]_ ;
  assign \new_[5897]_  = \new_[2807]_  | \new_[2808]_ ;
  assign \new_[5900]_  = \new_[2805]_  | \new_[2806]_ ;
  assign \new_[5901]_  = \new_[5900]_  | \new_[5897]_ ;
  assign \new_[5902]_  = \new_[5901]_  | \new_[5894]_ ;
  assign \new_[5903]_  = \new_[5902]_  | \new_[5887]_ ;
  assign \new_[5907]_  = \new_[2802]_  | \new_[2803]_ ;
  assign \new_[5908]_  = \new_[2804]_  | \new_[5907]_ ;
  assign \new_[5911]_  = \new_[2800]_  | \new_[2801]_ ;
  assign \new_[5914]_  = \new_[2798]_  | \new_[2799]_ ;
  assign \new_[5915]_  = \new_[5914]_  | \new_[5911]_ ;
  assign \new_[5916]_  = \new_[5915]_  | \new_[5908]_ ;
  assign \new_[5919]_  = \new_[2796]_  | \new_[2797]_ ;
  assign \new_[5922]_  = \new_[2794]_  | \new_[2795]_ ;
  assign \new_[5923]_  = \new_[5922]_  | \new_[5919]_ ;
  assign \new_[5926]_  = \new_[2792]_  | \new_[2793]_ ;
  assign \new_[5929]_  = \new_[2790]_  | \new_[2791]_ ;
  assign \new_[5930]_  = \new_[5929]_  | \new_[5926]_ ;
  assign \new_[5931]_  = \new_[5930]_  | \new_[5923]_ ;
  assign \new_[5932]_  = \new_[5931]_  | \new_[5916]_ ;
  assign \new_[5933]_  = \new_[5932]_  | \new_[5903]_ ;
  assign \new_[5937]_  = \new_[2787]_  | \new_[2788]_ ;
  assign \new_[5938]_  = \new_[2789]_  | \new_[5937]_ ;
  assign \new_[5941]_  = \new_[2785]_  | \new_[2786]_ ;
  assign \new_[5944]_  = \new_[2783]_  | \new_[2784]_ ;
  assign \new_[5945]_  = \new_[5944]_  | \new_[5941]_ ;
  assign \new_[5946]_  = \new_[5945]_  | \new_[5938]_ ;
  assign \new_[5949]_  = \new_[2781]_  | \new_[2782]_ ;
  assign \new_[5952]_  = \new_[2779]_  | \new_[2780]_ ;
  assign \new_[5953]_  = \new_[5952]_  | \new_[5949]_ ;
  assign \new_[5956]_  = \new_[2777]_  | \new_[2778]_ ;
  assign \new_[5959]_  = \new_[2775]_  | \new_[2776]_ ;
  assign \new_[5960]_  = \new_[5959]_  | \new_[5956]_ ;
  assign \new_[5961]_  = \new_[5960]_  | \new_[5953]_ ;
  assign \new_[5962]_  = \new_[5961]_  | \new_[5946]_ ;
  assign \new_[5966]_  = \new_[2772]_  | \new_[2773]_ ;
  assign \new_[5967]_  = \new_[2774]_  | \new_[5966]_ ;
  assign \new_[5970]_  = \new_[2770]_  | \new_[2771]_ ;
  assign \new_[5973]_  = \new_[2768]_  | \new_[2769]_ ;
  assign \new_[5974]_  = \new_[5973]_  | \new_[5970]_ ;
  assign \new_[5975]_  = \new_[5974]_  | \new_[5967]_ ;
  assign \new_[5978]_  = \new_[2766]_  | \new_[2767]_ ;
  assign \new_[5981]_  = \new_[2764]_  | \new_[2765]_ ;
  assign \new_[5982]_  = \new_[5981]_  | \new_[5978]_ ;
  assign \new_[5985]_  = \new_[2762]_  | \new_[2763]_ ;
  assign \new_[5988]_  = \new_[2760]_  | \new_[2761]_ ;
  assign \new_[5989]_  = \new_[5988]_  | \new_[5985]_ ;
  assign \new_[5990]_  = \new_[5989]_  | \new_[5982]_ ;
  assign \new_[5991]_  = \new_[5990]_  | \new_[5975]_ ;
  assign \new_[5992]_  = \new_[5991]_  | \new_[5962]_ ;
  assign \new_[5993]_  = \new_[5992]_  | \new_[5933]_ ;
  assign \new_[5994]_  = \new_[5993]_  | \new_[5874]_ ;
  assign \new_[5998]_  = \new_[2757]_  | \new_[2758]_ ;
  assign \new_[5999]_  = \new_[2759]_  | \new_[5998]_ ;
  assign \new_[6002]_  = \new_[2755]_  | \new_[2756]_ ;
  assign \new_[6005]_  = \new_[2753]_  | \new_[2754]_ ;
  assign \new_[6006]_  = \new_[6005]_  | \new_[6002]_ ;
  assign \new_[6007]_  = \new_[6006]_  | \new_[5999]_ ;
  assign \new_[6010]_  = \new_[2751]_  | \new_[2752]_ ;
  assign \new_[6013]_  = \new_[2749]_  | \new_[2750]_ ;
  assign \new_[6014]_  = \new_[6013]_  | \new_[6010]_ ;
  assign \new_[6017]_  = \new_[2747]_  | \new_[2748]_ ;
  assign \new_[6020]_  = \new_[2745]_  | \new_[2746]_ ;
  assign \new_[6021]_  = \new_[6020]_  | \new_[6017]_ ;
  assign \new_[6022]_  = \new_[6021]_  | \new_[6014]_ ;
  assign \new_[6023]_  = \new_[6022]_  | \new_[6007]_ ;
  assign \new_[6027]_  = \new_[2742]_  | \new_[2743]_ ;
  assign \new_[6028]_  = \new_[2744]_  | \new_[6027]_ ;
  assign \new_[6031]_  = \new_[2740]_  | \new_[2741]_ ;
  assign \new_[6034]_  = \new_[2738]_  | \new_[2739]_ ;
  assign \new_[6035]_  = \new_[6034]_  | \new_[6031]_ ;
  assign \new_[6036]_  = \new_[6035]_  | \new_[6028]_ ;
  assign \new_[6039]_  = \new_[2736]_  | \new_[2737]_ ;
  assign \new_[6042]_  = \new_[2734]_  | \new_[2735]_ ;
  assign \new_[6043]_  = \new_[6042]_  | \new_[6039]_ ;
  assign \new_[6046]_  = \new_[2732]_  | \new_[2733]_ ;
  assign \new_[6049]_  = \new_[2730]_  | \new_[2731]_ ;
  assign \new_[6050]_  = \new_[6049]_  | \new_[6046]_ ;
  assign \new_[6051]_  = \new_[6050]_  | \new_[6043]_ ;
  assign \new_[6052]_  = \new_[6051]_  | \new_[6036]_ ;
  assign \new_[6053]_  = \new_[6052]_  | \new_[6023]_ ;
  assign \new_[6057]_  = \new_[2727]_  | \new_[2728]_ ;
  assign \new_[6058]_  = \new_[2729]_  | \new_[6057]_ ;
  assign \new_[6061]_  = \new_[2725]_  | \new_[2726]_ ;
  assign \new_[6064]_  = \new_[2723]_  | \new_[2724]_ ;
  assign \new_[6065]_  = \new_[6064]_  | \new_[6061]_ ;
  assign \new_[6066]_  = \new_[6065]_  | \new_[6058]_ ;
  assign \new_[6069]_  = \new_[2721]_  | \new_[2722]_ ;
  assign \new_[6072]_  = \new_[2719]_  | \new_[2720]_ ;
  assign \new_[6073]_  = \new_[6072]_  | \new_[6069]_ ;
  assign \new_[6076]_  = \new_[2717]_  | \new_[2718]_ ;
  assign \new_[6079]_  = \new_[2715]_  | \new_[2716]_ ;
  assign \new_[6080]_  = \new_[6079]_  | \new_[6076]_ ;
  assign \new_[6081]_  = \new_[6080]_  | \new_[6073]_ ;
  assign \new_[6082]_  = \new_[6081]_  | \new_[6066]_ ;
  assign \new_[6086]_  = \new_[2712]_  | \new_[2713]_ ;
  assign \new_[6087]_  = \new_[2714]_  | \new_[6086]_ ;
  assign \new_[6090]_  = \new_[2710]_  | \new_[2711]_ ;
  assign \new_[6093]_  = \new_[2708]_  | \new_[2709]_ ;
  assign \new_[6094]_  = \new_[6093]_  | \new_[6090]_ ;
  assign \new_[6095]_  = \new_[6094]_  | \new_[6087]_ ;
  assign \new_[6098]_  = \new_[2706]_  | \new_[2707]_ ;
  assign \new_[6101]_  = \new_[2704]_  | \new_[2705]_ ;
  assign \new_[6102]_  = \new_[6101]_  | \new_[6098]_ ;
  assign \new_[6105]_  = \new_[2702]_  | \new_[2703]_ ;
  assign \new_[6108]_  = \new_[2700]_  | \new_[2701]_ ;
  assign \new_[6109]_  = \new_[6108]_  | \new_[6105]_ ;
  assign \new_[6110]_  = \new_[6109]_  | \new_[6102]_ ;
  assign \new_[6111]_  = \new_[6110]_  | \new_[6095]_ ;
  assign \new_[6112]_  = \new_[6111]_  | \new_[6082]_ ;
  assign \new_[6113]_  = \new_[6112]_  | \new_[6053]_ ;
  assign \new_[6117]_  = \new_[2697]_  | \new_[2698]_ ;
  assign \new_[6118]_  = \new_[2699]_  | \new_[6117]_ ;
  assign \new_[6121]_  = \new_[2695]_  | \new_[2696]_ ;
  assign \new_[6124]_  = \new_[2693]_  | \new_[2694]_ ;
  assign \new_[6125]_  = \new_[6124]_  | \new_[6121]_ ;
  assign \new_[6126]_  = \new_[6125]_  | \new_[6118]_ ;
  assign \new_[6129]_  = \new_[2691]_  | \new_[2692]_ ;
  assign \new_[6132]_  = \new_[2689]_  | \new_[2690]_ ;
  assign \new_[6133]_  = \new_[6132]_  | \new_[6129]_ ;
  assign \new_[6136]_  = \new_[2687]_  | \new_[2688]_ ;
  assign \new_[6139]_  = \new_[2685]_  | \new_[2686]_ ;
  assign \new_[6140]_  = \new_[6139]_  | \new_[6136]_ ;
  assign \new_[6141]_  = \new_[6140]_  | \new_[6133]_ ;
  assign \new_[6142]_  = \new_[6141]_  | \new_[6126]_ ;
  assign \new_[6146]_  = \new_[2682]_  | \new_[2683]_ ;
  assign \new_[6147]_  = \new_[2684]_  | \new_[6146]_ ;
  assign \new_[6150]_  = \new_[2680]_  | \new_[2681]_ ;
  assign \new_[6153]_  = \new_[2678]_  | \new_[2679]_ ;
  assign \new_[6154]_  = \new_[6153]_  | \new_[6150]_ ;
  assign \new_[6155]_  = \new_[6154]_  | \new_[6147]_ ;
  assign \new_[6158]_  = \new_[2676]_  | \new_[2677]_ ;
  assign \new_[6161]_  = \new_[2674]_  | \new_[2675]_ ;
  assign \new_[6162]_  = \new_[6161]_  | \new_[6158]_ ;
  assign \new_[6165]_  = \new_[2672]_  | \new_[2673]_ ;
  assign \new_[6168]_  = \new_[2670]_  | \new_[2671]_ ;
  assign \new_[6169]_  = \new_[6168]_  | \new_[6165]_ ;
  assign \new_[6170]_  = \new_[6169]_  | \new_[6162]_ ;
  assign \new_[6171]_  = \new_[6170]_  | \new_[6155]_ ;
  assign \new_[6172]_  = \new_[6171]_  | \new_[6142]_ ;
  assign \new_[6176]_  = \new_[2667]_  | \new_[2668]_ ;
  assign \new_[6177]_  = \new_[2669]_  | \new_[6176]_ ;
  assign \new_[6180]_  = \new_[2665]_  | \new_[2666]_ ;
  assign \new_[6183]_  = \new_[2663]_  | \new_[2664]_ ;
  assign \new_[6184]_  = \new_[6183]_  | \new_[6180]_ ;
  assign \new_[6185]_  = \new_[6184]_  | \new_[6177]_ ;
  assign \new_[6188]_  = \new_[2661]_  | \new_[2662]_ ;
  assign \new_[6191]_  = \new_[2659]_  | \new_[2660]_ ;
  assign \new_[6192]_  = \new_[6191]_  | \new_[6188]_ ;
  assign \new_[6195]_  = \new_[2657]_  | \new_[2658]_ ;
  assign \new_[6198]_  = \new_[2655]_  | \new_[2656]_ ;
  assign \new_[6199]_  = \new_[6198]_  | \new_[6195]_ ;
  assign \new_[6200]_  = \new_[6199]_  | \new_[6192]_ ;
  assign \new_[6201]_  = \new_[6200]_  | \new_[6185]_ ;
  assign \new_[6205]_  = \new_[2652]_  | \new_[2653]_ ;
  assign \new_[6206]_  = \new_[2654]_  | \new_[6205]_ ;
  assign \new_[6209]_  = \new_[2650]_  | \new_[2651]_ ;
  assign \new_[6212]_  = \new_[2648]_  | \new_[2649]_ ;
  assign \new_[6213]_  = \new_[6212]_  | \new_[6209]_ ;
  assign \new_[6214]_  = \new_[6213]_  | \new_[6206]_ ;
  assign \new_[6217]_  = \new_[2646]_  | \new_[2647]_ ;
  assign \new_[6220]_  = \new_[2644]_  | \new_[2645]_ ;
  assign \new_[6221]_  = \new_[6220]_  | \new_[6217]_ ;
  assign \new_[6224]_  = \new_[2642]_  | \new_[2643]_ ;
  assign \new_[6227]_  = \new_[2640]_  | \new_[2641]_ ;
  assign \new_[6228]_  = \new_[6227]_  | \new_[6224]_ ;
  assign \new_[6229]_  = \new_[6228]_  | \new_[6221]_ ;
  assign \new_[6230]_  = \new_[6229]_  | \new_[6214]_ ;
  assign \new_[6231]_  = \new_[6230]_  | \new_[6201]_ ;
  assign \new_[6232]_  = \new_[6231]_  | \new_[6172]_ ;
  assign \new_[6233]_  = \new_[6232]_  | \new_[6113]_ ;
  assign \new_[6234]_  = \new_[6233]_  | \new_[5994]_ ;
  assign \new_[6238]_  = \new_[2637]_  | \new_[2638]_ ;
  assign \new_[6239]_  = \new_[2639]_  | \new_[6238]_ ;
  assign \new_[6242]_  = \new_[2635]_  | \new_[2636]_ ;
  assign \new_[6245]_  = \new_[2633]_  | \new_[2634]_ ;
  assign \new_[6246]_  = \new_[6245]_  | \new_[6242]_ ;
  assign \new_[6247]_  = \new_[6246]_  | \new_[6239]_ ;
  assign \new_[6250]_  = \new_[2631]_  | \new_[2632]_ ;
  assign \new_[6253]_  = \new_[2629]_  | \new_[2630]_ ;
  assign \new_[6254]_  = \new_[6253]_  | \new_[6250]_ ;
  assign \new_[6257]_  = \new_[2627]_  | \new_[2628]_ ;
  assign \new_[6260]_  = \new_[2625]_  | \new_[2626]_ ;
  assign \new_[6261]_  = \new_[6260]_  | \new_[6257]_ ;
  assign \new_[6262]_  = \new_[6261]_  | \new_[6254]_ ;
  assign \new_[6263]_  = \new_[6262]_  | \new_[6247]_ ;
  assign \new_[6267]_  = \new_[2622]_  | \new_[2623]_ ;
  assign \new_[6268]_  = \new_[2624]_  | \new_[6267]_ ;
  assign \new_[6271]_  = \new_[2620]_  | \new_[2621]_ ;
  assign \new_[6274]_  = \new_[2618]_  | \new_[2619]_ ;
  assign \new_[6275]_  = \new_[6274]_  | \new_[6271]_ ;
  assign \new_[6276]_  = \new_[6275]_  | \new_[6268]_ ;
  assign \new_[6279]_  = \new_[2616]_  | \new_[2617]_ ;
  assign \new_[6282]_  = \new_[2614]_  | \new_[2615]_ ;
  assign \new_[6283]_  = \new_[6282]_  | \new_[6279]_ ;
  assign \new_[6286]_  = \new_[2612]_  | \new_[2613]_ ;
  assign \new_[6289]_  = \new_[2610]_  | \new_[2611]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6286]_ ;
  assign \new_[6291]_  = \new_[6290]_  | \new_[6283]_ ;
  assign \new_[6292]_  = \new_[6291]_  | \new_[6276]_ ;
  assign \new_[6293]_  = \new_[6292]_  | \new_[6263]_ ;
  assign \new_[6297]_  = \new_[2607]_  | \new_[2608]_ ;
  assign \new_[6298]_  = \new_[2609]_  | \new_[6297]_ ;
  assign \new_[6301]_  = \new_[2605]_  | \new_[2606]_ ;
  assign \new_[6304]_  = \new_[2603]_  | \new_[2604]_ ;
  assign \new_[6305]_  = \new_[6304]_  | \new_[6301]_ ;
  assign \new_[6306]_  = \new_[6305]_  | \new_[6298]_ ;
  assign \new_[6309]_  = \new_[2601]_  | \new_[2602]_ ;
  assign \new_[6312]_  = \new_[2599]_  | \new_[2600]_ ;
  assign \new_[6313]_  = \new_[6312]_  | \new_[6309]_ ;
  assign \new_[6316]_  = \new_[2597]_  | \new_[2598]_ ;
  assign \new_[6319]_  = \new_[2595]_  | \new_[2596]_ ;
  assign \new_[6320]_  = \new_[6319]_  | \new_[6316]_ ;
  assign \new_[6321]_  = \new_[6320]_  | \new_[6313]_ ;
  assign \new_[6322]_  = \new_[6321]_  | \new_[6306]_ ;
  assign \new_[6326]_  = \new_[2592]_  | \new_[2593]_ ;
  assign \new_[6327]_  = \new_[2594]_  | \new_[6326]_ ;
  assign \new_[6330]_  = \new_[2590]_  | \new_[2591]_ ;
  assign \new_[6333]_  = \new_[2588]_  | \new_[2589]_ ;
  assign \new_[6334]_  = \new_[6333]_  | \new_[6330]_ ;
  assign \new_[6335]_  = \new_[6334]_  | \new_[6327]_ ;
  assign \new_[6338]_  = \new_[2586]_  | \new_[2587]_ ;
  assign \new_[6341]_  = \new_[2584]_  | \new_[2585]_ ;
  assign \new_[6342]_  = \new_[6341]_  | \new_[6338]_ ;
  assign \new_[6345]_  = \new_[2582]_  | \new_[2583]_ ;
  assign \new_[6348]_  = \new_[2580]_  | \new_[2581]_ ;
  assign \new_[6349]_  = \new_[6348]_  | \new_[6345]_ ;
  assign \new_[6350]_  = \new_[6349]_  | \new_[6342]_ ;
  assign \new_[6351]_  = \new_[6350]_  | \new_[6335]_ ;
  assign \new_[6352]_  = \new_[6351]_  | \new_[6322]_ ;
  assign \new_[6353]_  = \new_[6352]_  | \new_[6293]_ ;
  assign \new_[6357]_  = \new_[2577]_  | \new_[2578]_ ;
  assign \new_[6358]_  = \new_[2579]_  | \new_[6357]_ ;
  assign \new_[6361]_  = \new_[2575]_  | \new_[2576]_ ;
  assign \new_[6364]_  = \new_[2573]_  | \new_[2574]_ ;
  assign \new_[6365]_  = \new_[6364]_  | \new_[6361]_ ;
  assign \new_[6366]_  = \new_[6365]_  | \new_[6358]_ ;
  assign \new_[6369]_  = \new_[2571]_  | \new_[2572]_ ;
  assign \new_[6372]_  = \new_[2569]_  | \new_[2570]_ ;
  assign \new_[6373]_  = \new_[6372]_  | \new_[6369]_ ;
  assign \new_[6376]_  = \new_[2567]_  | \new_[2568]_ ;
  assign \new_[6379]_  = \new_[2565]_  | \new_[2566]_ ;
  assign \new_[6380]_  = \new_[6379]_  | \new_[6376]_ ;
  assign \new_[6381]_  = \new_[6380]_  | \new_[6373]_ ;
  assign \new_[6382]_  = \new_[6381]_  | \new_[6366]_ ;
  assign \new_[6386]_  = \new_[2562]_  | \new_[2563]_ ;
  assign \new_[6387]_  = \new_[2564]_  | \new_[6386]_ ;
  assign \new_[6390]_  = \new_[2560]_  | \new_[2561]_ ;
  assign \new_[6393]_  = \new_[2558]_  | \new_[2559]_ ;
  assign \new_[6394]_  = \new_[6393]_  | \new_[6390]_ ;
  assign \new_[6395]_  = \new_[6394]_  | \new_[6387]_ ;
  assign \new_[6398]_  = \new_[2556]_  | \new_[2557]_ ;
  assign \new_[6401]_  = \new_[2554]_  | \new_[2555]_ ;
  assign \new_[6402]_  = \new_[6401]_  | \new_[6398]_ ;
  assign \new_[6405]_  = \new_[2552]_  | \new_[2553]_ ;
  assign \new_[6408]_  = \new_[2550]_  | \new_[2551]_ ;
  assign \new_[6409]_  = \new_[6408]_  | \new_[6405]_ ;
  assign \new_[6410]_  = \new_[6409]_  | \new_[6402]_ ;
  assign \new_[6411]_  = \new_[6410]_  | \new_[6395]_ ;
  assign \new_[6412]_  = \new_[6411]_  | \new_[6382]_ ;
  assign \new_[6416]_  = \new_[2547]_  | \new_[2548]_ ;
  assign \new_[6417]_  = \new_[2549]_  | \new_[6416]_ ;
  assign \new_[6420]_  = \new_[2545]_  | \new_[2546]_ ;
  assign \new_[6423]_  = \new_[2543]_  | \new_[2544]_ ;
  assign \new_[6424]_  = \new_[6423]_  | \new_[6420]_ ;
  assign \new_[6425]_  = \new_[6424]_  | \new_[6417]_ ;
  assign \new_[6428]_  = \new_[2541]_  | \new_[2542]_ ;
  assign \new_[6431]_  = \new_[2539]_  | \new_[2540]_ ;
  assign \new_[6432]_  = \new_[6431]_  | \new_[6428]_ ;
  assign \new_[6435]_  = \new_[2537]_  | \new_[2538]_ ;
  assign \new_[6438]_  = \new_[2535]_  | \new_[2536]_ ;
  assign \new_[6439]_  = \new_[6438]_  | \new_[6435]_ ;
  assign \new_[6440]_  = \new_[6439]_  | \new_[6432]_ ;
  assign \new_[6441]_  = \new_[6440]_  | \new_[6425]_ ;
  assign \new_[6445]_  = \new_[2532]_  | \new_[2533]_ ;
  assign \new_[6446]_  = \new_[2534]_  | \new_[6445]_ ;
  assign \new_[6449]_  = \new_[2530]_  | \new_[2531]_ ;
  assign \new_[6452]_  = \new_[2528]_  | \new_[2529]_ ;
  assign \new_[6453]_  = \new_[6452]_  | \new_[6449]_ ;
  assign \new_[6454]_  = \new_[6453]_  | \new_[6446]_ ;
  assign \new_[6457]_  = \new_[2526]_  | \new_[2527]_ ;
  assign \new_[6460]_  = \new_[2524]_  | \new_[2525]_ ;
  assign \new_[6461]_  = \new_[6460]_  | \new_[6457]_ ;
  assign \new_[6464]_  = \new_[2522]_  | \new_[2523]_ ;
  assign \new_[6467]_  = \new_[2520]_  | \new_[2521]_ ;
  assign \new_[6468]_  = \new_[6467]_  | \new_[6464]_ ;
  assign \new_[6469]_  = \new_[6468]_  | \new_[6461]_ ;
  assign \new_[6470]_  = \new_[6469]_  | \new_[6454]_ ;
  assign \new_[6471]_  = \new_[6470]_  | \new_[6441]_ ;
  assign \new_[6472]_  = \new_[6471]_  | \new_[6412]_ ;
  assign \new_[6473]_  = \new_[6472]_  | \new_[6353]_ ;
  assign \new_[6477]_  = \new_[2517]_  | \new_[2518]_ ;
  assign \new_[6478]_  = \new_[2519]_  | \new_[6477]_ ;
  assign \new_[6481]_  = \new_[2515]_  | \new_[2516]_ ;
  assign \new_[6484]_  = \new_[2513]_  | \new_[2514]_ ;
  assign \new_[6485]_  = \new_[6484]_  | \new_[6481]_ ;
  assign \new_[6486]_  = \new_[6485]_  | \new_[6478]_ ;
  assign \new_[6489]_  = \new_[2511]_  | \new_[2512]_ ;
  assign \new_[6492]_  = \new_[2509]_  | \new_[2510]_ ;
  assign \new_[6493]_  = \new_[6492]_  | \new_[6489]_ ;
  assign \new_[6496]_  = \new_[2507]_  | \new_[2508]_ ;
  assign \new_[6499]_  = \new_[2505]_  | \new_[2506]_ ;
  assign \new_[6500]_  = \new_[6499]_  | \new_[6496]_ ;
  assign \new_[6501]_  = \new_[6500]_  | \new_[6493]_ ;
  assign \new_[6502]_  = \new_[6501]_  | \new_[6486]_ ;
  assign \new_[6506]_  = \new_[2502]_  | \new_[2503]_ ;
  assign \new_[6507]_  = \new_[2504]_  | \new_[6506]_ ;
  assign \new_[6510]_  = \new_[2500]_  | \new_[2501]_ ;
  assign \new_[6513]_  = \new_[2498]_  | \new_[2499]_ ;
  assign \new_[6514]_  = \new_[6513]_  | \new_[6510]_ ;
  assign \new_[6515]_  = \new_[6514]_  | \new_[6507]_ ;
  assign \new_[6518]_  = \new_[2496]_  | \new_[2497]_ ;
  assign \new_[6521]_  = \new_[2494]_  | \new_[2495]_ ;
  assign \new_[6522]_  = \new_[6521]_  | \new_[6518]_ ;
  assign \new_[6525]_  = \new_[2492]_  | \new_[2493]_ ;
  assign \new_[6528]_  = \new_[2490]_  | \new_[2491]_ ;
  assign \new_[6529]_  = \new_[6528]_  | \new_[6525]_ ;
  assign \new_[6530]_  = \new_[6529]_  | \new_[6522]_ ;
  assign \new_[6531]_  = \new_[6530]_  | \new_[6515]_ ;
  assign \new_[6532]_  = \new_[6531]_  | \new_[6502]_ ;
  assign \new_[6536]_  = \new_[2487]_  | \new_[2488]_ ;
  assign \new_[6537]_  = \new_[2489]_  | \new_[6536]_ ;
  assign \new_[6540]_  = \new_[2485]_  | \new_[2486]_ ;
  assign \new_[6543]_  = \new_[2483]_  | \new_[2484]_ ;
  assign \new_[6544]_  = \new_[6543]_  | \new_[6540]_ ;
  assign \new_[6545]_  = \new_[6544]_  | \new_[6537]_ ;
  assign \new_[6548]_  = \new_[2481]_  | \new_[2482]_ ;
  assign \new_[6551]_  = \new_[2479]_  | \new_[2480]_ ;
  assign \new_[6552]_  = \new_[6551]_  | \new_[6548]_ ;
  assign \new_[6555]_  = \new_[2477]_  | \new_[2478]_ ;
  assign \new_[6558]_  = \new_[2475]_  | \new_[2476]_ ;
  assign \new_[6559]_  = \new_[6558]_  | \new_[6555]_ ;
  assign \new_[6560]_  = \new_[6559]_  | \new_[6552]_ ;
  assign \new_[6561]_  = \new_[6560]_  | \new_[6545]_ ;
  assign \new_[6565]_  = \new_[2472]_  | \new_[2473]_ ;
  assign \new_[6566]_  = \new_[2474]_  | \new_[6565]_ ;
  assign \new_[6569]_  = \new_[2470]_  | \new_[2471]_ ;
  assign \new_[6572]_  = \new_[2468]_  | \new_[2469]_ ;
  assign \new_[6573]_  = \new_[6572]_  | \new_[6569]_ ;
  assign \new_[6574]_  = \new_[6573]_  | \new_[6566]_ ;
  assign \new_[6577]_  = \new_[2466]_  | \new_[2467]_ ;
  assign \new_[6580]_  = \new_[2464]_  | \new_[2465]_ ;
  assign \new_[6581]_  = \new_[6580]_  | \new_[6577]_ ;
  assign \new_[6584]_  = \new_[2462]_  | \new_[2463]_ ;
  assign \new_[6587]_  = \new_[2460]_  | \new_[2461]_ ;
  assign \new_[6588]_  = \new_[6587]_  | \new_[6584]_ ;
  assign \new_[6589]_  = \new_[6588]_  | \new_[6581]_ ;
  assign \new_[6590]_  = \new_[6589]_  | \new_[6574]_ ;
  assign \new_[6591]_  = \new_[6590]_  | \new_[6561]_ ;
  assign \new_[6592]_  = \new_[6591]_  | \new_[6532]_ ;
  assign \new_[6596]_  = \new_[2457]_  | \new_[2458]_ ;
  assign \new_[6597]_  = \new_[2459]_  | \new_[6596]_ ;
  assign \new_[6600]_  = \new_[2455]_  | \new_[2456]_ ;
  assign \new_[6603]_  = \new_[2453]_  | \new_[2454]_ ;
  assign \new_[6604]_  = \new_[6603]_  | \new_[6600]_ ;
  assign \new_[6605]_  = \new_[6604]_  | \new_[6597]_ ;
  assign \new_[6608]_  = \new_[2451]_  | \new_[2452]_ ;
  assign \new_[6611]_  = \new_[2449]_  | \new_[2450]_ ;
  assign \new_[6612]_  = \new_[6611]_  | \new_[6608]_ ;
  assign \new_[6615]_  = \new_[2447]_  | \new_[2448]_ ;
  assign \new_[6618]_  = \new_[2445]_  | \new_[2446]_ ;
  assign \new_[6619]_  = \new_[6618]_  | \new_[6615]_ ;
  assign \new_[6620]_  = \new_[6619]_  | \new_[6612]_ ;
  assign \new_[6621]_  = \new_[6620]_  | \new_[6605]_ ;
  assign \new_[6625]_  = \new_[2442]_  | \new_[2443]_ ;
  assign \new_[6626]_  = \new_[2444]_  | \new_[6625]_ ;
  assign \new_[6629]_  = \new_[2440]_  | \new_[2441]_ ;
  assign \new_[6632]_  = \new_[2438]_  | \new_[2439]_ ;
  assign \new_[6633]_  = \new_[6632]_  | \new_[6629]_ ;
  assign \new_[6634]_  = \new_[6633]_  | \new_[6626]_ ;
  assign \new_[6637]_  = \new_[2436]_  | \new_[2437]_ ;
  assign \new_[6640]_  = \new_[2434]_  | \new_[2435]_ ;
  assign \new_[6641]_  = \new_[6640]_  | \new_[6637]_ ;
  assign \new_[6644]_  = \new_[2432]_  | \new_[2433]_ ;
  assign \new_[6647]_  = \new_[2430]_  | \new_[2431]_ ;
  assign \new_[6648]_  = \new_[6647]_  | \new_[6644]_ ;
  assign \new_[6649]_  = \new_[6648]_  | \new_[6641]_ ;
  assign \new_[6650]_  = \new_[6649]_  | \new_[6634]_ ;
  assign \new_[6651]_  = \new_[6650]_  | \new_[6621]_ ;
  assign \new_[6655]_  = \new_[2427]_  | \new_[2428]_ ;
  assign \new_[6656]_  = \new_[2429]_  | \new_[6655]_ ;
  assign \new_[6659]_  = \new_[2425]_  | \new_[2426]_ ;
  assign \new_[6662]_  = \new_[2423]_  | \new_[2424]_ ;
  assign \new_[6663]_  = \new_[6662]_  | \new_[6659]_ ;
  assign \new_[6664]_  = \new_[6663]_  | \new_[6656]_ ;
  assign \new_[6667]_  = \new_[2421]_  | \new_[2422]_ ;
  assign \new_[6670]_  = \new_[2419]_  | \new_[2420]_ ;
  assign \new_[6671]_  = \new_[6670]_  | \new_[6667]_ ;
  assign \new_[6674]_  = \new_[2417]_  | \new_[2418]_ ;
  assign \new_[6677]_  = \new_[2415]_  | \new_[2416]_ ;
  assign \new_[6678]_  = \new_[6677]_  | \new_[6674]_ ;
  assign \new_[6679]_  = \new_[6678]_  | \new_[6671]_ ;
  assign \new_[6680]_  = \new_[6679]_  | \new_[6664]_ ;
  assign \new_[6684]_  = \new_[2412]_  | \new_[2413]_ ;
  assign \new_[6685]_  = \new_[2414]_  | \new_[6684]_ ;
  assign \new_[6688]_  = \new_[2410]_  | \new_[2411]_ ;
  assign \new_[6691]_  = \new_[2408]_  | \new_[2409]_ ;
  assign \new_[6692]_  = \new_[6691]_  | \new_[6688]_ ;
  assign \new_[6693]_  = \new_[6692]_  | \new_[6685]_ ;
  assign \new_[6696]_  = \new_[2406]_  | \new_[2407]_ ;
  assign \new_[6699]_  = \new_[2404]_  | \new_[2405]_ ;
  assign \new_[6700]_  = \new_[6699]_  | \new_[6696]_ ;
  assign \new_[6703]_  = \new_[2402]_  | \new_[2403]_ ;
  assign \new_[6706]_  = \new_[2400]_  | \new_[2401]_ ;
  assign \new_[6707]_  = \new_[6706]_  | \new_[6703]_ ;
  assign \new_[6708]_  = \new_[6707]_  | \new_[6700]_ ;
  assign \new_[6709]_  = \new_[6708]_  | \new_[6693]_ ;
  assign \new_[6710]_  = \new_[6709]_  | \new_[6680]_ ;
  assign \new_[6711]_  = \new_[6710]_  | \new_[6651]_ ;
  assign \new_[6712]_  = \new_[6711]_  | \new_[6592]_ ;
  assign \new_[6713]_  = \new_[6712]_  | \new_[6473]_ ;
  assign \new_[6714]_  = \new_[6713]_  | \new_[6234]_ ;
  assign \new_[6718]_  = \new_[2397]_  | \new_[2398]_ ;
  assign \new_[6719]_  = \new_[2399]_  | \new_[6718]_ ;
  assign \new_[6722]_  = \new_[2395]_  | \new_[2396]_ ;
  assign \new_[6725]_  = \new_[2393]_  | \new_[2394]_ ;
  assign \new_[6726]_  = \new_[6725]_  | \new_[6722]_ ;
  assign \new_[6727]_  = \new_[6726]_  | \new_[6719]_ ;
  assign \new_[6730]_  = \new_[2391]_  | \new_[2392]_ ;
  assign \new_[6733]_  = \new_[2389]_  | \new_[2390]_ ;
  assign \new_[6734]_  = \new_[6733]_  | \new_[6730]_ ;
  assign \new_[6737]_  = \new_[2387]_  | \new_[2388]_ ;
  assign \new_[6740]_  = \new_[2385]_  | \new_[2386]_ ;
  assign \new_[6741]_  = \new_[6740]_  | \new_[6737]_ ;
  assign \new_[6742]_  = \new_[6741]_  | \new_[6734]_ ;
  assign \new_[6743]_  = \new_[6742]_  | \new_[6727]_ ;
  assign \new_[6747]_  = \new_[2382]_  | \new_[2383]_ ;
  assign \new_[6748]_  = \new_[2384]_  | \new_[6747]_ ;
  assign \new_[6751]_  = \new_[2380]_  | \new_[2381]_ ;
  assign \new_[6754]_  = \new_[2378]_  | \new_[2379]_ ;
  assign \new_[6755]_  = \new_[6754]_  | \new_[6751]_ ;
  assign \new_[6756]_  = \new_[6755]_  | \new_[6748]_ ;
  assign \new_[6759]_  = \new_[2376]_  | \new_[2377]_ ;
  assign \new_[6762]_  = \new_[2374]_  | \new_[2375]_ ;
  assign \new_[6763]_  = \new_[6762]_  | \new_[6759]_ ;
  assign \new_[6766]_  = \new_[2372]_  | \new_[2373]_ ;
  assign \new_[6769]_  = \new_[2370]_  | \new_[2371]_ ;
  assign \new_[6770]_  = \new_[6769]_  | \new_[6766]_ ;
  assign \new_[6771]_  = \new_[6770]_  | \new_[6763]_ ;
  assign \new_[6772]_  = \new_[6771]_  | \new_[6756]_ ;
  assign \new_[6773]_  = \new_[6772]_  | \new_[6743]_ ;
  assign \new_[6777]_  = \new_[2367]_  | \new_[2368]_ ;
  assign \new_[6778]_  = \new_[2369]_  | \new_[6777]_ ;
  assign \new_[6781]_  = \new_[2365]_  | \new_[2366]_ ;
  assign \new_[6784]_  = \new_[2363]_  | \new_[2364]_ ;
  assign \new_[6785]_  = \new_[6784]_  | \new_[6781]_ ;
  assign \new_[6786]_  = \new_[6785]_  | \new_[6778]_ ;
  assign \new_[6789]_  = \new_[2361]_  | \new_[2362]_ ;
  assign \new_[6792]_  = \new_[2359]_  | \new_[2360]_ ;
  assign \new_[6793]_  = \new_[6792]_  | \new_[6789]_ ;
  assign \new_[6796]_  = \new_[2357]_  | \new_[2358]_ ;
  assign \new_[6799]_  = \new_[2355]_  | \new_[2356]_ ;
  assign \new_[6800]_  = \new_[6799]_  | \new_[6796]_ ;
  assign \new_[6801]_  = \new_[6800]_  | \new_[6793]_ ;
  assign \new_[6802]_  = \new_[6801]_  | \new_[6786]_ ;
  assign \new_[6806]_  = \new_[2352]_  | \new_[2353]_ ;
  assign \new_[6807]_  = \new_[2354]_  | \new_[6806]_ ;
  assign \new_[6810]_  = \new_[2350]_  | \new_[2351]_ ;
  assign \new_[6813]_  = \new_[2348]_  | \new_[2349]_ ;
  assign \new_[6814]_  = \new_[6813]_  | \new_[6810]_ ;
  assign \new_[6815]_  = \new_[6814]_  | \new_[6807]_ ;
  assign \new_[6818]_  = \new_[2346]_  | \new_[2347]_ ;
  assign \new_[6821]_  = \new_[2344]_  | \new_[2345]_ ;
  assign \new_[6822]_  = \new_[6821]_  | \new_[6818]_ ;
  assign \new_[6825]_  = \new_[2342]_  | \new_[2343]_ ;
  assign \new_[6828]_  = \new_[2340]_  | \new_[2341]_ ;
  assign \new_[6829]_  = \new_[6828]_  | \new_[6825]_ ;
  assign \new_[6830]_  = \new_[6829]_  | \new_[6822]_ ;
  assign \new_[6831]_  = \new_[6830]_  | \new_[6815]_ ;
  assign \new_[6832]_  = \new_[6831]_  | \new_[6802]_ ;
  assign \new_[6833]_  = \new_[6832]_  | \new_[6773]_ ;
  assign \new_[6837]_  = \new_[2337]_  | \new_[2338]_ ;
  assign \new_[6838]_  = \new_[2339]_  | \new_[6837]_ ;
  assign \new_[6841]_  = \new_[2335]_  | \new_[2336]_ ;
  assign \new_[6844]_  = \new_[2333]_  | \new_[2334]_ ;
  assign \new_[6845]_  = \new_[6844]_  | \new_[6841]_ ;
  assign \new_[6846]_  = \new_[6845]_  | \new_[6838]_ ;
  assign \new_[6849]_  = \new_[2331]_  | \new_[2332]_ ;
  assign \new_[6852]_  = \new_[2329]_  | \new_[2330]_ ;
  assign \new_[6853]_  = \new_[6852]_  | \new_[6849]_ ;
  assign \new_[6856]_  = \new_[2327]_  | \new_[2328]_ ;
  assign \new_[6859]_  = \new_[2325]_  | \new_[2326]_ ;
  assign \new_[6860]_  = \new_[6859]_  | \new_[6856]_ ;
  assign \new_[6861]_  = \new_[6860]_  | \new_[6853]_ ;
  assign \new_[6862]_  = \new_[6861]_  | \new_[6846]_ ;
  assign \new_[6866]_  = \new_[2322]_  | \new_[2323]_ ;
  assign \new_[6867]_  = \new_[2324]_  | \new_[6866]_ ;
  assign \new_[6870]_  = \new_[2320]_  | \new_[2321]_ ;
  assign \new_[6873]_  = \new_[2318]_  | \new_[2319]_ ;
  assign \new_[6874]_  = \new_[6873]_  | \new_[6870]_ ;
  assign \new_[6875]_  = \new_[6874]_  | \new_[6867]_ ;
  assign \new_[6878]_  = \new_[2316]_  | \new_[2317]_ ;
  assign \new_[6881]_  = \new_[2314]_  | \new_[2315]_ ;
  assign \new_[6882]_  = \new_[6881]_  | \new_[6878]_ ;
  assign \new_[6885]_  = \new_[2312]_  | \new_[2313]_ ;
  assign \new_[6888]_  = \new_[2310]_  | \new_[2311]_ ;
  assign \new_[6889]_  = \new_[6888]_  | \new_[6885]_ ;
  assign \new_[6890]_  = \new_[6889]_  | \new_[6882]_ ;
  assign \new_[6891]_  = \new_[6890]_  | \new_[6875]_ ;
  assign \new_[6892]_  = \new_[6891]_  | \new_[6862]_ ;
  assign \new_[6896]_  = \new_[2307]_  | \new_[2308]_ ;
  assign \new_[6897]_  = \new_[2309]_  | \new_[6896]_ ;
  assign \new_[6900]_  = \new_[2305]_  | \new_[2306]_ ;
  assign \new_[6903]_  = \new_[2303]_  | \new_[2304]_ ;
  assign \new_[6904]_  = \new_[6903]_  | \new_[6900]_ ;
  assign \new_[6905]_  = \new_[6904]_  | \new_[6897]_ ;
  assign \new_[6908]_  = \new_[2301]_  | \new_[2302]_ ;
  assign \new_[6911]_  = \new_[2299]_  | \new_[2300]_ ;
  assign \new_[6912]_  = \new_[6911]_  | \new_[6908]_ ;
  assign \new_[6915]_  = \new_[2297]_  | \new_[2298]_ ;
  assign \new_[6918]_  = \new_[2295]_  | \new_[2296]_ ;
  assign \new_[6919]_  = \new_[6918]_  | \new_[6915]_ ;
  assign \new_[6920]_  = \new_[6919]_  | \new_[6912]_ ;
  assign \new_[6921]_  = \new_[6920]_  | \new_[6905]_ ;
  assign \new_[6925]_  = \new_[2292]_  | \new_[2293]_ ;
  assign \new_[6926]_  = \new_[2294]_  | \new_[6925]_ ;
  assign \new_[6929]_  = \new_[2290]_  | \new_[2291]_ ;
  assign \new_[6932]_  = \new_[2288]_  | \new_[2289]_ ;
  assign \new_[6933]_  = \new_[6932]_  | \new_[6929]_ ;
  assign \new_[6934]_  = \new_[6933]_  | \new_[6926]_ ;
  assign \new_[6937]_  = \new_[2286]_  | \new_[2287]_ ;
  assign \new_[6940]_  = \new_[2284]_  | \new_[2285]_ ;
  assign \new_[6941]_  = \new_[6940]_  | \new_[6937]_ ;
  assign \new_[6944]_  = \new_[2282]_  | \new_[2283]_ ;
  assign \new_[6947]_  = \new_[2280]_  | \new_[2281]_ ;
  assign \new_[6948]_  = \new_[6947]_  | \new_[6944]_ ;
  assign \new_[6949]_  = \new_[6948]_  | \new_[6941]_ ;
  assign \new_[6950]_  = \new_[6949]_  | \new_[6934]_ ;
  assign \new_[6951]_  = \new_[6950]_  | \new_[6921]_ ;
  assign \new_[6952]_  = \new_[6951]_  | \new_[6892]_ ;
  assign \new_[6953]_  = \new_[6952]_  | \new_[6833]_ ;
  assign \new_[6957]_  = \new_[2277]_  | \new_[2278]_ ;
  assign \new_[6958]_  = \new_[2279]_  | \new_[6957]_ ;
  assign \new_[6961]_  = \new_[2275]_  | \new_[2276]_ ;
  assign \new_[6964]_  = \new_[2273]_  | \new_[2274]_ ;
  assign \new_[6965]_  = \new_[6964]_  | \new_[6961]_ ;
  assign \new_[6966]_  = \new_[6965]_  | \new_[6958]_ ;
  assign \new_[6969]_  = \new_[2271]_  | \new_[2272]_ ;
  assign \new_[6972]_  = \new_[2269]_  | \new_[2270]_ ;
  assign \new_[6973]_  = \new_[6972]_  | \new_[6969]_ ;
  assign \new_[6976]_  = \new_[2267]_  | \new_[2268]_ ;
  assign \new_[6979]_  = \new_[2265]_  | \new_[2266]_ ;
  assign \new_[6980]_  = \new_[6979]_  | \new_[6976]_ ;
  assign \new_[6981]_  = \new_[6980]_  | \new_[6973]_ ;
  assign \new_[6982]_  = \new_[6981]_  | \new_[6966]_ ;
  assign \new_[6986]_  = \new_[2262]_  | \new_[2263]_ ;
  assign \new_[6987]_  = \new_[2264]_  | \new_[6986]_ ;
  assign \new_[6990]_  = \new_[2260]_  | \new_[2261]_ ;
  assign \new_[6993]_  = \new_[2258]_  | \new_[2259]_ ;
  assign \new_[6994]_  = \new_[6993]_  | \new_[6990]_ ;
  assign \new_[6995]_  = \new_[6994]_  | \new_[6987]_ ;
  assign \new_[6998]_  = \new_[2256]_  | \new_[2257]_ ;
  assign \new_[7001]_  = \new_[2254]_  | \new_[2255]_ ;
  assign \new_[7002]_  = \new_[7001]_  | \new_[6998]_ ;
  assign \new_[7005]_  = \new_[2252]_  | \new_[2253]_ ;
  assign \new_[7008]_  = \new_[2250]_  | \new_[2251]_ ;
  assign \new_[7009]_  = \new_[7008]_  | \new_[7005]_ ;
  assign \new_[7010]_  = \new_[7009]_  | \new_[7002]_ ;
  assign \new_[7011]_  = \new_[7010]_  | \new_[6995]_ ;
  assign \new_[7012]_  = \new_[7011]_  | \new_[6982]_ ;
  assign \new_[7016]_  = \new_[2247]_  | \new_[2248]_ ;
  assign \new_[7017]_  = \new_[2249]_  | \new_[7016]_ ;
  assign \new_[7020]_  = \new_[2245]_  | \new_[2246]_ ;
  assign \new_[7023]_  = \new_[2243]_  | \new_[2244]_ ;
  assign \new_[7024]_  = \new_[7023]_  | \new_[7020]_ ;
  assign \new_[7025]_  = \new_[7024]_  | \new_[7017]_ ;
  assign \new_[7028]_  = \new_[2241]_  | \new_[2242]_ ;
  assign \new_[7031]_  = \new_[2239]_  | \new_[2240]_ ;
  assign \new_[7032]_  = \new_[7031]_  | \new_[7028]_ ;
  assign \new_[7035]_  = \new_[2237]_  | \new_[2238]_ ;
  assign \new_[7038]_  = \new_[2235]_  | \new_[2236]_ ;
  assign \new_[7039]_  = \new_[7038]_  | \new_[7035]_ ;
  assign \new_[7040]_  = \new_[7039]_  | \new_[7032]_ ;
  assign \new_[7041]_  = \new_[7040]_  | \new_[7025]_ ;
  assign \new_[7045]_  = \new_[2232]_  | \new_[2233]_ ;
  assign \new_[7046]_  = \new_[2234]_  | \new_[7045]_ ;
  assign \new_[7049]_  = \new_[2230]_  | \new_[2231]_ ;
  assign \new_[7052]_  = \new_[2228]_  | \new_[2229]_ ;
  assign \new_[7053]_  = \new_[7052]_  | \new_[7049]_ ;
  assign \new_[7054]_  = \new_[7053]_  | \new_[7046]_ ;
  assign \new_[7057]_  = \new_[2226]_  | \new_[2227]_ ;
  assign \new_[7060]_  = \new_[2224]_  | \new_[2225]_ ;
  assign \new_[7061]_  = \new_[7060]_  | \new_[7057]_ ;
  assign \new_[7064]_  = \new_[2222]_  | \new_[2223]_ ;
  assign \new_[7067]_  = \new_[2220]_  | \new_[2221]_ ;
  assign \new_[7068]_  = \new_[7067]_  | \new_[7064]_ ;
  assign \new_[7069]_  = \new_[7068]_  | \new_[7061]_ ;
  assign \new_[7070]_  = \new_[7069]_  | \new_[7054]_ ;
  assign \new_[7071]_  = \new_[7070]_  | \new_[7041]_ ;
  assign \new_[7072]_  = \new_[7071]_  | \new_[7012]_ ;
  assign \new_[7076]_  = \new_[2217]_  | \new_[2218]_ ;
  assign \new_[7077]_  = \new_[2219]_  | \new_[7076]_ ;
  assign \new_[7080]_  = \new_[2215]_  | \new_[2216]_ ;
  assign \new_[7083]_  = \new_[2213]_  | \new_[2214]_ ;
  assign \new_[7084]_  = \new_[7083]_  | \new_[7080]_ ;
  assign \new_[7085]_  = \new_[7084]_  | \new_[7077]_ ;
  assign \new_[7088]_  = \new_[2211]_  | \new_[2212]_ ;
  assign \new_[7091]_  = \new_[2209]_  | \new_[2210]_ ;
  assign \new_[7092]_  = \new_[7091]_  | \new_[7088]_ ;
  assign \new_[7095]_  = \new_[2207]_  | \new_[2208]_ ;
  assign \new_[7098]_  = \new_[2205]_  | \new_[2206]_ ;
  assign \new_[7099]_  = \new_[7098]_  | \new_[7095]_ ;
  assign \new_[7100]_  = \new_[7099]_  | \new_[7092]_ ;
  assign \new_[7101]_  = \new_[7100]_  | \new_[7085]_ ;
  assign \new_[7105]_  = \new_[2202]_  | \new_[2203]_ ;
  assign \new_[7106]_  = \new_[2204]_  | \new_[7105]_ ;
  assign \new_[7109]_  = \new_[2200]_  | \new_[2201]_ ;
  assign \new_[7112]_  = \new_[2198]_  | \new_[2199]_ ;
  assign \new_[7113]_  = \new_[7112]_  | \new_[7109]_ ;
  assign \new_[7114]_  = \new_[7113]_  | \new_[7106]_ ;
  assign \new_[7117]_  = \new_[2196]_  | \new_[2197]_ ;
  assign \new_[7120]_  = \new_[2194]_  | \new_[2195]_ ;
  assign \new_[7121]_  = \new_[7120]_  | \new_[7117]_ ;
  assign \new_[7124]_  = \new_[2192]_  | \new_[2193]_ ;
  assign \new_[7127]_  = \new_[2190]_  | \new_[2191]_ ;
  assign \new_[7128]_  = \new_[7127]_  | \new_[7124]_ ;
  assign \new_[7129]_  = \new_[7128]_  | \new_[7121]_ ;
  assign \new_[7130]_  = \new_[7129]_  | \new_[7114]_ ;
  assign \new_[7131]_  = \new_[7130]_  | \new_[7101]_ ;
  assign \new_[7135]_  = \new_[2187]_  | \new_[2188]_ ;
  assign \new_[7136]_  = \new_[2189]_  | \new_[7135]_ ;
  assign \new_[7139]_  = \new_[2185]_  | \new_[2186]_ ;
  assign \new_[7142]_  = \new_[2183]_  | \new_[2184]_ ;
  assign \new_[7143]_  = \new_[7142]_  | \new_[7139]_ ;
  assign \new_[7144]_  = \new_[7143]_  | \new_[7136]_ ;
  assign \new_[7147]_  = \new_[2181]_  | \new_[2182]_ ;
  assign \new_[7150]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[7151]_  = \new_[7150]_  | \new_[7147]_ ;
  assign \new_[7154]_  = \new_[2177]_  | \new_[2178]_ ;
  assign \new_[7157]_  = \new_[2175]_  | \new_[2176]_ ;
  assign \new_[7158]_  = \new_[7157]_  | \new_[7154]_ ;
  assign \new_[7159]_  = \new_[7158]_  | \new_[7151]_ ;
  assign \new_[7160]_  = \new_[7159]_  | \new_[7144]_ ;
  assign \new_[7164]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[7165]_  = \new_[2174]_  | \new_[7164]_ ;
  assign \new_[7168]_  = \new_[2170]_  | \new_[2171]_ ;
  assign \new_[7171]_  = \new_[2168]_  | \new_[2169]_ ;
  assign \new_[7172]_  = \new_[7171]_  | \new_[7168]_ ;
  assign \new_[7173]_  = \new_[7172]_  | \new_[7165]_ ;
  assign \new_[7176]_  = \new_[2166]_  | \new_[2167]_ ;
  assign \new_[7179]_  = \new_[2164]_  | \new_[2165]_ ;
  assign \new_[7180]_  = \new_[7179]_  | \new_[7176]_ ;
  assign \new_[7183]_  = \new_[2162]_  | \new_[2163]_ ;
  assign \new_[7186]_  = \new_[2160]_  | \new_[2161]_ ;
  assign \new_[7187]_  = \new_[7186]_  | \new_[7183]_ ;
  assign \new_[7188]_  = \new_[7187]_  | \new_[7180]_ ;
  assign \new_[7189]_  = \new_[7188]_  | \new_[7173]_ ;
  assign \new_[7190]_  = \new_[7189]_  | \new_[7160]_ ;
  assign \new_[7191]_  = \new_[7190]_  | \new_[7131]_ ;
  assign \new_[7192]_  = \new_[7191]_  | \new_[7072]_ ;
  assign \new_[7193]_  = \new_[7192]_  | \new_[6953]_ ;
  assign \new_[7197]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[7198]_  = \new_[2159]_  | \new_[7197]_ ;
  assign \new_[7201]_  = \new_[2155]_  | \new_[2156]_ ;
  assign \new_[7204]_  = \new_[2153]_  | \new_[2154]_ ;
  assign \new_[7205]_  = \new_[7204]_  | \new_[7201]_ ;
  assign \new_[7206]_  = \new_[7205]_  | \new_[7198]_ ;
  assign \new_[7209]_  = \new_[2151]_  | \new_[2152]_ ;
  assign \new_[7212]_  = \new_[2149]_  | \new_[2150]_ ;
  assign \new_[7213]_  = \new_[7212]_  | \new_[7209]_ ;
  assign \new_[7216]_  = \new_[2147]_  | \new_[2148]_ ;
  assign \new_[7219]_  = \new_[2145]_  | \new_[2146]_ ;
  assign \new_[7220]_  = \new_[7219]_  | \new_[7216]_ ;
  assign \new_[7221]_  = \new_[7220]_  | \new_[7213]_ ;
  assign \new_[7222]_  = \new_[7221]_  | \new_[7206]_ ;
  assign \new_[7226]_  = \new_[2142]_  | \new_[2143]_ ;
  assign \new_[7227]_  = \new_[2144]_  | \new_[7226]_ ;
  assign \new_[7230]_  = \new_[2140]_  | \new_[2141]_ ;
  assign \new_[7233]_  = \new_[2138]_  | \new_[2139]_ ;
  assign \new_[7234]_  = \new_[7233]_  | \new_[7230]_ ;
  assign \new_[7235]_  = \new_[7234]_  | \new_[7227]_ ;
  assign \new_[7238]_  = \new_[2136]_  | \new_[2137]_ ;
  assign \new_[7241]_  = \new_[2134]_  | \new_[2135]_ ;
  assign \new_[7242]_  = \new_[7241]_  | \new_[7238]_ ;
  assign \new_[7245]_  = \new_[2132]_  | \new_[2133]_ ;
  assign \new_[7248]_  = \new_[2130]_  | \new_[2131]_ ;
  assign \new_[7249]_  = \new_[7248]_  | \new_[7245]_ ;
  assign \new_[7250]_  = \new_[7249]_  | \new_[7242]_ ;
  assign \new_[7251]_  = \new_[7250]_  | \new_[7235]_ ;
  assign \new_[7252]_  = \new_[7251]_  | \new_[7222]_ ;
  assign \new_[7256]_  = \new_[2127]_  | \new_[2128]_ ;
  assign \new_[7257]_  = \new_[2129]_  | \new_[7256]_ ;
  assign \new_[7260]_  = \new_[2125]_  | \new_[2126]_ ;
  assign \new_[7263]_  = \new_[2123]_  | \new_[2124]_ ;
  assign \new_[7264]_  = \new_[7263]_  | \new_[7260]_ ;
  assign \new_[7265]_  = \new_[7264]_  | \new_[7257]_ ;
  assign \new_[7268]_  = \new_[2121]_  | \new_[2122]_ ;
  assign \new_[7271]_  = \new_[2119]_  | \new_[2120]_ ;
  assign \new_[7272]_  = \new_[7271]_  | \new_[7268]_ ;
  assign \new_[7275]_  = \new_[2117]_  | \new_[2118]_ ;
  assign \new_[7278]_  = \new_[2115]_  | \new_[2116]_ ;
  assign \new_[7279]_  = \new_[7278]_  | \new_[7275]_ ;
  assign \new_[7280]_  = \new_[7279]_  | \new_[7272]_ ;
  assign \new_[7281]_  = \new_[7280]_  | \new_[7265]_ ;
  assign \new_[7285]_  = \new_[2112]_  | \new_[2113]_ ;
  assign \new_[7286]_  = \new_[2114]_  | \new_[7285]_ ;
  assign \new_[7289]_  = \new_[2110]_  | \new_[2111]_ ;
  assign \new_[7292]_  = \new_[2108]_  | \new_[2109]_ ;
  assign \new_[7293]_  = \new_[7292]_  | \new_[7289]_ ;
  assign \new_[7294]_  = \new_[7293]_  | \new_[7286]_ ;
  assign \new_[7297]_  = \new_[2106]_  | \new_[2107]_ ;
  assign \new_[7300]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[7301]_  = \new_[7300]_  | \new_[7297]_ ;
  assign \new_[7304]_  = \new_[2102]_  | \new_[2103]_ ;
  assign \new_[7307]_  = \new_[2100]_  | \new_[2101]_ ;
  assign \new_[7308]_  = \new_[7307]_  | \new_[7304]_ ;
  assign \new_[7309]_  = \new_[7308]_  | \new_[7301]_ ;
  assign \new_[7310]_  = \new_[7309]_  | \new_[7294]_ ;
  assign \new_[7311]_  = \new_[7310]_  | \new_[7281]_ ;
  assign \new_[7312]_  = \new_[7311]_  | \new_[7252]_ ;
  assign \new_[7316]_  = \new_[2097]_  | \new_[2098]_ ;
  assign \new_[7317]_  = \new_[2099]_  | \new_[7316]_ ;
  assign \new_[7320]_  = \new_[2095]_  | \new_[2096]_ ;
  assign \new_[7323]_  = \new_[2093]_  | \new_[2094]_ ;
  assign \new_[7324]_  = \new_[7323]_  | \new_[7320]_ ;
  assign \new_[7325]_  = \new_[7324]_  | \new_[7317]_ ;
  assign \new_[7328]_  = \new_[2091]_  | \new_[2092]_ ;
  assign \new_[7331]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[7332]_  = \new_[7331]_  | \new_[7328]_ ;
  assign \new_[7335]_  = \new_[2087]_  | \new_[2088]_ ;
  assign \new_[7338]_  = \new_[2085]_  | \new_[2086]_ ;
  assign \new_[7339]_  = \new_[7338]_  | \new_[7335]_ ;
  assign \new_[7340]_  = \new_[7339]_  | \new_[7332]_ ;
  assign \new_[7341]_  = \new_[7340]_  | \new_[7325]_ ;
  assign \new_[7345]_  = \new_[2082]_  | \new_[2083]_ ;
  assign \new_[7346]_  = \new_[2084]_  | \new_[7345]_ ;
  assign \new_[7349]_  = \new_[2080]_  | \new_[2081]_ ;
  assign \new_[7352]_  = \new_[2078]_  | \new_[2079]_ ;
  assign \new_[7353]_  = \new_[7352]_  | \new_[7349]_ ;
  assign \new_[7354]_  = \new_[7353]_  | \new_[7346]_ ;
  assign \new_[7357]_  = \new_[2076]_  | \new_[2077]_ ;
  assign \new_[7360]_  = \new_[2074]_  | \new_[2075]_ ;
  assign \new_[7361]_  = \new_[7360]_  | \new_[7357]_ ;
  assign \new_[7364]_  = \new_[2072]_  | \new_[2073]_ ;
  assign \new_[7367]_  = \new_[2070]_  | \new_[2071]_ ;
  assign \new_[7368]_  = \new_[7367]_  | \new_[7364]_ ;
  assign \new_[7369]_  = \new_[7368]_  | \new_[7361]_ ;
  assign \new_[7370]_  = \new_[7369]_  | \new_[7354]_ ;
  assign \new_[7371]_  = \new_[7370]_  | \new_[7341]_ ;
  assign \new_[7375]_  = \new_[2067]_  | \new_[2068]_ ;
  assign \new_[7376]_  = \new_[2069]_  | \new_[7375]_ ;
  assign \new_[7379]_  = \new_[2065]_  | \new_[2066]_ ;
  assign \new_[7382]_  = \new_[2063]_  | \new_[2064]_ ;
  assign \new_[7383]_  = \new_[7382]_  | \new_[7379]_ ;
  assign \new_[7384]_  = \new_[7383]_  | \new_[7376]_ ;
  assign \new_[7387]_  = \new_[2061]_  | \new_[2062]_ ;
  assign \new_[7390]_  = \new_[2059]_  | \new_[2060]_ ;
  assign \new_[7391]_  = \new_[7390]_  | \new_[7387]_ ;
  assign \new_[7394]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[7397]_  = \new_[2055]_  | \new_[2056]_ ;
  assign \new_[7398]_  = \new_[7397]_  | \new_[7394]_ ;
  assign \new_[7399]_  = \new_[7398]_  | \new_[7391]_ ;
  assign \new_[7400]_  = \new_[7399]_  | \new_[7384]_ ;
  assign \new_[7404]_  = \new_[2052]_  | \new_[2053]_ ;
  assign \new_[7405]_  = \new_[2054]_  | \new_[7404]_ ;
  assign \new_[7408]_  = \new_[2050]_  | \new_[2051]_ ;
  assign \new_[7411]_  = \new_[2048]_  | \new_[2049]_ ;
  assign \new_[7412]_  = \new_[7411]_  | \new_[7408]_ ;
  assign \new_[7413]_  = \new_[7412]_  | \new_[7405]_ ;
  assign \new_[7416]_  = \new_[2046]_  | \new_[2047]_ ;
  assign \new_[7419]_  = \new_[2044]_  | \new_[2045]_ ;
  assign \new_[7420]_  = \new_[7419]_  | \new_[7416]_ ;
  assign \new_[7423]_  = \new_[2042]_  | \new_[2043]_ ;
  assign \new_[7426]_  = \new_[2040]_  | \new_[2041]_ ;
  assign \new_[7427]_  = \new_[7426]_  | \new_[7423]_ ;
  assign \new_[7428]_  = \new_[7427]_  | \new_[7420]_ ;
  assign \new_[7429]_  = \new_[7428]_  | \new_[7413]_ ;
  assign \new_[7430]_  = \new_[7429]_  | \new_[7400]_ ;
  assign \new_[7431]_  = \new_[7430]_  | \new_[7371]_ ;
  assign \new_[7432]_  = \new_[7431]_  | \new_[7312]_ ;
  assign \new_[7436]_  = \new_[2037]_  | \new_[2038]_ ;
  assign \new_[7437]_  = \new_[2039]_  | \new_[7436]_ ;
  assign \new_[7440]_  = \new_[2035]_  | \new_[2036]_ ;
  assign \new_[7443]_  = \new_[2033]_  | \new_[2034]_ ;
  assign \new_[7444]_  = \new_[7443]_  | \new_[7440]_ ;
  assign \new_[7445]_  = \new_[7444]_  | \new_[7437]_ ;
  assign \new_[7448]_  = \new_[2031]_  | \new_[2032]_ ;
  assign \new_[7451]_  = \new_[2029]_  | \new_[2030]_ ;
  assign \new_[7452]_  = \new_[7451]_  | \new_[7448]_ ;
  assign \new_[7455]_  = \new_[2027]_  | \new_[2028]_ ;
  assign \new_[7458]_  = \new_[2025]_  | \new_[2026]_ ;
  assign \new_[7459]_  = \new_[7458]_  | \new_[7455]_ ;
  assign \new_[7460]_  = \new_[7459]_  | \new_[7452]_ ;
  assign \new_[7461]_  = \new_[7460]_  | \new_[7445]_ ;
  assign \new_[7465]_  = \new_[2022]_  | \new_[2023]_ ;
  assign \new_[7466]_  = \new_[2024]_  | \new_[7465]_ ;
  assign \new_[7469]_  = \new_[2020]_  | \new_[2021]_ ;
  assign \new_[7472]_  = \new_[2018]_  | \new_[2019]_ ;
  assign \new_[7473]_  = \new_[7472]_  | \new_[7469]_ ;
  assign \new_[7474]_  = \new_[7473]_  | \new_[7466]_ ;
  assign \new_[7477]_  = \new_[2016]_  | \new_[2017]_ ;
  assign \new_[7480]_  = \new_[2014]_  | \new_[2015]_ ;
  assign \new_[7481]_  = \new_[7480]_  | \new_[7477]_ ;
  assign \new_[7484]_  = \new_[2012]_  | \new_[2013]_ ;
  assign \new_[7487]_  = \new_[2010]_  | \new_[2011]_ ;
  assign \new_[7488]_  = \new_[7487]_  | \new_[7484]_ ;
  assign \new_[7489]_  = \new_[7488]_  | \new_[7481]_ ;
  assign \new_[7490]_  = \new_[7489]_  | \new_[7474]_ ;
  assign \new_[7491]_  = \new_[7490]_  | \new_[7461]_ ;
  assign \new_[7495]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[7496]_  = \new_[2009]_  | \new_[7495]_ ;
  assign \new_[7499]_  = \new_[2005]_  | \new_[2006]_ ;
  assign \new_[7502]_  = \new_[2003]_  | \new_[2004]_ ;
  assign \new_[7503]_  = \new_[7502]_  | \new_[7499]_ ;
  assign \new_[7504]_  = \new_[7503]_  | \new_[7496]_ ;
  assign \new_[7507]_  = \new_[2001]_  | \new_[2002]_ ;
  assign \new_[7510]_  = \new_[1999]_  | \new_[2000]_ ;
  assign \new_[7511]_  = \new_[7510]_  | \new_[7507]_ ;
  assign \new_[7514]_  = \new_[1997]_  | \new_[1998]_ ;
  assign \new_[7517]_  = \new_[1995]_  | \new_[1996]_ ;
  assign \new_[7518]_  = \new_[7517]_  | \new_[7514]_ ;
  assign \new_[7519]_  = \new_[7518]_  | \new_[7511]_ ;
  assign \new_[7520]_  = \new_[7519]_  | \new_[7504]_ ;
  assign \new_[7524]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[7525]_  = \new_[1994]_  | \new_[7524]_ ;
  assign \new_[7528]_  = \new_[1990]_  | \new_[1991]_ ;
  assign \new_[7531]_  = \new_[1988]_  | \new_[1989]_ ;
  assign \new_[7532]_  = \new_[7531]_  | \new_[7528]_ ;
  assign \new_[7533]_  = \new_[7532]_  | \new_[7525]_ ;
  assign \new_[7536]_  = \new_[1986]_  | \new_[1987]_ ;
  assign \new_[7539]_  = \new_[1984]_  | \new_[1985]_ ;
  assign \new_[7540]_  = \new_[7539]_  | \new_[7536]_ ;
  assign \new_[7543]_  = \new_[1982]_  | \new_[1983]_ ;
  assign \new_[7546]_  = \new_[1980]_  | \new_[1981]_ ;
  assign \new_[7547]_  = \new_[7546]_  | \new_[7543]_ ;
  assign \new_[7548]_  = \new_[7547]_  | \new_[7540]_ ;
  assign \new_[7549]_  = \new_[7548]_  | \new_[7533]_ ;
  assign \new_[7550]_  = \new_[7549]_  | \new_[7520]_ ;
  assign \new_[7551]_  = \new_[7550]_  | \new_[7491]_ ;
  assign \new_[7555]_  = \new_[1977]_  | \new_[1978]_ ;
  assign \new_[7556]_  = \new_[1979]_  | \new_[7555]_ ;
  assign \new_[7559]_  = \new_[1975]_  | \new_[1976]_ ;
  assign \new_[7562]_  = \new_[1973]_  | \new_[1974]_ ;
  assign \new_[7563]_  = \new_[7562]_  | \new_[7559]_ ;
  assign \new_[7564]_  = \new_[7563]_  | \new_[7556]_ ;
  assign \new_[7567]_  = \new_[1971]_  | \new_[1972]_ ;
  assign \new_[7570]_  = \new_[1969]_  | \new_[1970]_ ;
  assign \new_[7571]_  = \new_[7570]_  | \new_[7567]_ ;
  assign \new_[7574]_  = \new_[1967]_  | \new_[1968]_ ;
  assign \new_[7577]_  = \new_[1965]_  | \new_[1966]_ ;
  assign \new_[7578]_  = \new_[7577]_  | \new_[7574]_ ;
  assign \new_[7579]_  = \new_[7578]_  | \new_[7571]_ ;
  assign \new_[7580]_  = \new_[7579]_  | \new_[7564]_ ;
  assign \new_[7584]_  = \new_[1962]_  | \new_[1963]_ ;
  assign \new_[7585]_  = \new_[1964]_  | \new_[7584]_ ;
  assign \new_[7588]_  = \new_[1960]_  | \new_[1961]_ ;
  assign \new_[7591]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[7592]_  = \new_[7591]_  | \new_[7588]_ ;
  assign \new_[7593]_  = \new_[7592]_  | \new_[7585]_ ;
  assign \new_[7596]_  = \new_[1956]_  | \new_[1957]_ ;
  assign \new_[7599]_  = \new_[1954]_  | \new_[1955]_ ;
  assign \new_[7600]_  = \new_[7599]_  | \new_[7596]_ ;
  assign \new_[7603]_  = \new_[1952]_  | \new_[1953]_ ;
  assign \new_[7606]_  = \new_[1950]_  | \new_[1951]_ ;
  assign \new_[7607]_  = \new_[7606]_  | \new_[7603]_ ;
  assign \new_[7608]_  = \new_[7607]_  | \new_[7600]_ ;
  assign \new_[7609]_  = \new_[7608]_  | \new_[7593]_ ;
  assign \new_[7610]_  = \new_[7609]_  | \new_[7580]_ ;
  assign \new_[7614]_  = \new_[1947]_  | \new_[1948]_ ;
  assign \new_[7615]_  = \new_[1949]_  | \new_[7614]_ ;
  assign \new_[7618]_  = \new_[1945]_  | \new_[1946]_ ;
  assign \new_[7621]_  = \new_[1943]_  | \new_[1944]_ ;
  assign \new_[7622]_  = \new_[7621]_  | \new_[7618]_ ;
  assign \new_[7623]_  = \new_[7622]_  | \new_[7615]_ ;
  assign \new_[7626]_  = \new_[1941]_  | \new_[1942]_ ;
  assign \new_[7629]_  = \new_[1939]_  | \new_[1940]_ ;
  assign \new_[7630]_  = \new_[7629]_  | \new_[7626]_ ;
  assign \new_[7633]_  = \new_[1937]_  | \new_[1938]_ ;
  assign \new_[7636]_  = \new_[1935]_  | \new_[1936]_ ;
  assign \new_[7637]_  = \new_[7636]_  | \new_[7633]_ ;
  assign \new_[7638]_  = \new_[7637]_  | \new_[7630]_ ;
  assign \new_[7639]_  = \new_[7638]_  | \new_[7623]_ ;
  assign \new_[7643]_  = \new_[1932]_  | \new_[1933]_ ;
  assign \new_[7644]_  = \new_[1934]_  | \new_[7643]_ ;
  assign \new_[7647]_  = \new_[1930]_  | \new_[1931]_ ;
  assign \new_[7650]_  = \new_[1928]_  | \new_[1929]_ ;
  assign \new_[7651]_  = \new_[7650]_  | \new_[7647]_ ;
  assign \new_[7652]_  = \new_[7651]_  | \new_[7644]_ ;
  assign \new_[7655]_  = \new_[1926]_  | \new_[1927]_ ;
  assign \new_[7658]_  = \new_[1924]_  | \new_[1925]_ ;
  assign \new_[7659]_  = \new_[7658]_  | \new_[7655]_ ;
  assign \new_[7662]_  = \new_[1922]_  | \new_[1923]_ ;
  assign \new_[7665]_  = \new_[1920]_  | \new_[1921]_ ;
  assign \new_[7666]_  = \new_[7665]_  | \new_[7662]_ ;
  assign \new_[7667]_  = \new_[7666]_  | \new_[7659]_ ;
  assign \new_[7668]_  = \new_[7667]_  | \new_[7652]_ ;
  assign \new_[7669]_  = \new_[7668]_  | \new_[7639]_ ;
  assign \new_[7670]_  = \new_[7669]_  | \new_[7610]_ ;
  assign \new_[7671]_  = \new_[7670]_  | \new_[7551]_ ;
  assign \new_[7672]_  = \new_[7671]_  | \new_[7432]_ ;
  assign \new_[7673]_  = \new_[7672]_  | \new_[7193]_ ;
  assign \new_[7674]_  = \new_[7673]_  | \new_[6714]_ ;
  assign \new_[7675]_  = \new_[7674]_  | \new_[5755]_ ;
  assign \new_[7679]_  = \new_[1917]_  | \new_[1918]_ ;
  assign \new_[7680]_  = \new_[1919]_  | \new_[7679]_ ;
  assign \new_[7683]_  = \new_[1915]_  | \new_[1916]_ ;
  assign \new_[7686]_  = \new_[1913]_  | \new_[1914]_ ;
  assign \new_[7687]_  = \new_[7686]_  | \new_[7683]_ ;
  assign \new_[7688]_  = \new_[7687]_  | \new_[7680]_ ;
  assign \new_[7692]_  = \new_[1910]_  | \new_[1911]_ ;
  assign \new_[7693]_  = \new_[1912]_  | \new_[7692]_ ;
  assign \new_[7696]_  = \new_[1908]_  | \new_[1909]_ ;
  assign \new_[7699]_  = \new_[1906]_  | \new_[1907]_ ;
  assign \new_[7700]_  = \new_[7699]_  | \new_[7696]_ ;
  assign \new_[7701]_  = \new_[7700]_  | \new_[7693]_ ;
  assign \new_[7702]_  = \new_[7701]_  | \new_[7688]_ ;
  assign \new_[7706]_  = \new_[1903]_  | \new_[1904]_ ;
  assign \new_[7707]_  = \new_[1905]_  | \new_[7706]_ ;
  assign \new_[7710]_  = \new_[1901]_  | \new_[1902]_ ;
  assign \new_[7713]_  = \new_[1899]_  | \new_[1900]_ ;
  assign \new_[7714]_  = \new_[7713]_  | \new_[7710]_ ;
  assign \new_[7715]_  = \new_[7714]_  | \new_[7707]_ ;
  assign \new_[7718]_  = \new_[1897]_  | \new_[1898]_ ;
  assign \new_[7721]_  = \new_[1895]_  | \new_[1896]_ ;
  assign \new_[7722]_  = \new_[7721]_  | \new_[7718]_ ;
  assign \new_[7725]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[7728]_  = \new_[1891]_  | \new_[1892]_ ;
  assign \new_[7729]_  = \new_[7728]_  | \new_[7725]_ ;
  assign \new_[7730]_  = \new_[7729]_  | \new_[7722]_ ;
  assign \new_[7731]_  = \new_[7730]_  | \new_[7715]_ ;
  assign \new_[7732]_  = \new_[7731]_  | \new_[7702]_ ;
  assign \new_[7736]_  = \new_[1888]_  | \new_[1889]_ ;
  assign \new_[7737]_  = \new_[1890]_  | \new_[7736]_ ;
  assign \new_[7740]_  = \new_[1886]_  | \new_[1887]_ ;
  assign \new_[7743]_  = \new_[1884]_  | \new_[1885]_ ;
  assign \new_[7744]_  = \new_[7743]_  | \new_[7740]_ ;
  assign \new_[7745]_  = \new_[7744]_  | \new_[7737]_ ;
  assign \new_[7748]_  = \new_[1882]_  | \new_[1883]_ ;
  assign \new_[7751]_  = \new_[1880]_  | \new_[1881]_ ;
  assign \new_[7752]_  = \new_[7751]_  | \new_[7748]_ ;
  assign \new_[7755]_  = \new_[1878]_  | \new_[1879]_ ;
  assign \new_[7758]_  = \new_[1876]_  | \new_[1877]_ ;
  assign \new_[7759]_  = \new_[7758]_  | \new_[7755]_ ;
  assign \new_[7760]_  = \new_[7759]_  | \new_[7752]_ ;
  assign \new_[7761]_  = \new_[7760]_  | \new_[7745]_ ;
  assign \new_[7765]_  = \new_[1873]_  | \new_[1874]_ ;
  assign \new_[7766]_  = \new_[1875]_  | \new_[7765]_ ;
  assign \new_[7769]_  = \new_[1871]_  | \new_[1872]_ ;
  assign \new_[7772]_  = \new_[1869]_  | \new_[1870]_ ;
  assign \new_[7773]_  = \new_[7772]_  | \new_[7769]_ ;
  assign \new_[7774]_  = \new_[7773]_  | \new_[7766]_ ;
  assign \new_[7777]_  = \new_[1867]_  | \new_[1868]_ ;
  assign \new_[7780]_  = \new_[1865]_  | \new_[1866]_ ;
  assign \new_[7781]_  = \new_[7780]_  | \new_[7777]_ ;
  assign \new_[7784]_  = \new_[1863]_  | \new_[1864]_ ;
  assign \new_[7787]_  = \new_[1861]_  | \new_[1862]_ ;
  assign \new_[7788]_  = \new_[7787]_  | \new_[7784]_ ;
  assign \new_[7789]_  = \new_[7788]_  | \new_[7781]_ ;
  assign \new_[7790]_  = \new_[7789]_  | \new_[7774]_ ;
  assign \new_[7791]_  = \new_[7790]_  | \new_[7761]_ ;
  assign \new_[7792]_  = \new_[7791]_  | \new_[7732]_ ;
  assign \new_[7796]_  = \new_[1858]_  | \new_[1859]_ ;
  assign \new_[7797]_  = \new_[1860]_  | \new_[7796]_ ;
  assign \new_[7800]_  = \new_[1856]_  | \new_[1857]_ ;
  assign \new_[7803]_  = \new_[1854]_  | \new_[1855]_ ;
  assign \new_[7804]_  = \new_[7803]_  | \new_[7800]_ ;
  assign \new_[7805]_  = \new_[7804]_  | \new_[7797]_ ;
  assign \new_[7808]_  = \new_[1852]_  | \new_[1853]_ ;
  assign \new_[7811]_  = \new_[1850]_  | \new_[1851]_ ;
  assign \new_[7812]_  = \new_[7811]_  | \new_[7808]_ ;
  assign \new_[7815]_  = \new_[1848]_  | \new_[1849]_ ;
  assign \new_[7818]_  = \new_[1846]_  | \new_[1847]_ ;
  assign \new_[7819]_  = \new_[7818]_  | \new_[7815]_ ;
  assign \new_[7820]_  = \new_[7819]_  | \new_[7812]_ ;
  assign \new_[7821]_  = \new_[7820]_  | \new_[7805]_ ;
  assign \new_[7825]_  = \new_[1843]_  | \new_[1844]_ ;
  assign \new_[7826]_  = \new_[1845]_  | \new_[7825]_ ;
  assign \new_[7829]_  = \new_[1841]_  | \new_[1842]_ ;
  assign \new_[7832]_  = \new_[1839]_  | \new_[1840]_ ;
  assign \new_[7833]_  = \new_[7832]_  | \new_[7829]_ ;
  assign \new_[7834]_  = \new_[7833]_  | \new_[7826]_ ;
  assign \new_[7837]_  = \new_[1837]_  | \new_[1838]_ ;
  assign \new_[7840]_  = \new_[1835]_  | \new_[1836]_ ;
  assign \new_[7841]_  = \new_[7840]_  | \new_[7837]_ ;
  assign \new_[7844]_  = \new_[1833]_  | \new_[1834]_ ;
  assign \new_[7847]_  = \new_[1831]_  | \new_[1832]_ ;
  assign \new_[7848]_  = \new_[7847]_  | \new_[7844]_ ;
  assign \new_[7849]_  = \new_[7848]_  | \new_[7841]_ ;
  assign \new_[7850]_  = \new_[7849]_  | \new_[7834]_ ;
  assign \new_[7851]_  = \new_[7850]_  | \new_[7821]_ ;
  assign \new_[7855]_  = \new_[1828]_  | \new_[1829]_ ;
  assign \new_[7856]_  = \new_[1830]_  | \new_[7855]_ ;
  assign \new_[7859]_  = \new_[1826]_  | \new_[1827]_ ;
  assign \new_[7862]_  = \new_[1824]_  | \new_[1825]_ ;
  assign \new_[7863]_  = \new_[7862]_  | \new_[7859]_ ;
  assign \new_[7864]_  = \new_[7863]_  | \new_[7856]_ ;
  assign \new_[7867]_  = \new_[1822]_  | \new_[1823]_ ;
  assign \new_[7870]_  = \new_[1820]_  | \new_[1821]_ ;
  assign \new_[7871]_  = \new_[7870]_  | \new_[7867]_ ;
  assign \new_[7874]_  = \new_[1818]_  | \new_[1819]_ ;
  assign \new_[7877]_  = \new_[1816]_  | \new_[1817]_ ;
  assign \new_[7878]_  = \new_[7877]_  | \new_[7874]_ ;
  assign \new_[7879]_  = \new_[7878]_  | \new_[7871]_ ;
  assign \new_[7880]_  = \new_[7879]_  | \new_[7864]_ ;
  assign \new_[7884]_  = \new_[1813]_  | \new_[1814]_ ;
  assign \new_[7885]_  = \new_[1815]_  | \new_[7884]_ ;
  assign \new_[7888]_  = \new_[1811]_  | \new_[1812]_ ;
  assign \new_[7891]_  = \new_[1809]_  | \new_[1810]_ ;
  assign \new_[7892]_  = \new_[7891]_  | \new_[7888]_ ;
  assign \new_[7893]_  = \new_[7892]_  | \new_[7885]_ ;
  assign \new_[7896]_  = \new_[1807]_  | \new_[1808]_ ;
  assign \new_[7899]_  = \new_[1805]_  | \new_[1806]_ ;
  assign \new_[7900]_  = \new_[7899]_  | \new_[7896]_ ;
  assign \new_[7903]_  = \new_[1803]_  | \new_[1804]_ ;
  assign \new_[7906]_  = \new_[1801]_  | \new_[1802]_ ;
  assign \new_[7907]_  = \new_[7906]_  | \new_[7903]_ ;
  assign \new_[7908]_  = \new_[7907]_  | \new_[7900]_ ;
  assign \new_[7909]_  = \new_[7908]_  | \new_[7893]_ ;
  assign \new_[7910]_  = \new_[7909]_  | \new_[7880]_ ;
  assign \new_[7911]_  = \new_[7910]_  | \new_[7851]_ ;
  assign \new_[7912]_  = \new_[7911]_  | \new_[7792]_ ;
  assign \new_[7916]_  = \new_[1798]_  | \new_[1799]_ ;
  assign \new_[7917]_  = \new_[1800]_  | \new_[7916]_ ;
  assign \new_[7920]_  = \new_[1796]_  | \new_[1797]_ ;
  assign \new_[7923]_  = \new_[1794]_  | \new_[1795]_ ;
  assign \new_[7924]_  = \new_[7923]_  | \new_[7920]_ ;
  assign \new_[7925]_  = \new_[7924]_  | \new_[7917]_ ;
  assign \new_[7928]_  = \new_[1792]_  | \new_[1793]_ ;
  assign \new_[7931]_  = \new_[1790]_  | \new_[1791]_ ;
  assign \new_[7932]_  = \new_[7931]_  | \new_[7928]_ ;
  assign \new_[7935]_  = \new_[1788]_  | \new_[1789]_ ;
  assign \new_[7938]_  = \new_[1786]_  | \new_[1787]_ ;
  assign \new_[7939]_  = \new_[7938]_  | \new_[7935]_ ;
  assign \new_[7940]_  = \new_[7939]_  | \new_[7932]_ ;
  assign \new_[7941]_  = \new_[7940]_  | \new_[7925]_ ;
  assign \new_[7945]_  = \new_[1783]_  | \new_[1784]_ ;
  assign \new_[7946]_  = \new_[1785]_  | \new_[7945]_ ;
  assign \new_[7949]_  = \new_[1781]_  | \new_[1782]_ ;
  assign \new_[7952]_  = \new_[1779]_  | \new_[1780]_ ;
  assign \new_[7953]_  = \new_[7952]_  | \new_[7949]_ ;
  assign \new_[7954]_  = \new_[7953]_  | \new_[7946]_ ;
  assign \new_[7957]_  = \new_[1777]_  | \new_[1778]_ ;
  assign \new_[7960]_  = \new_[1775]_  | \new_[1776]_ ;
  assign \new_[7961]_  = \new_[7960]_  | \new_[7957]_ ;
  assign \new_[7964]_  = \new_[1773]_  | \new_[1774]_ ;
  assign \new_[7967]_  = \new_[1771]_  | \new_[1772]_ ;
  assign \new_[7968]_  = \new_[7967]_  | \new_[7964]_ ;
  assign \new_[7969]_  = \new_[7968]_  | \new_[7961]_ ;
  assign \new_[7970]_  = \new_[7969]_  | \new_[7954]_ ;
  assign \new_[7971]_  = \new_[7970]_  | \new_[7941]_ ;
  assign \new_[7975]_  = \new_[1768]_  | \new_[1769]_ ;
  assign \new_[7976]_  = \new_[1770]_  | \new_[7975]_ ;
  assign \new_[7979]_  = \new_[1766]_  | \new_[1767]_ ;
  assign \new_[7982]_  = \new_[1764]_  | \new_[1765]_ ;
  assign \new_[7983]_  = \new_[7982]_  | \new_[7979]_ ;
  assign \new_[7984]_  = \new_[7983]_  | \new_[7976]_ ;
  assign \new_[7987]_  = \new_[1762]_  | \new_[1763]_ ;
  assign \new_[7990]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[7991]_  = \new_[7990]_  | \new_[7987]_ ;
  assign \new_[7994]_  = \new_[1758]_  | \new_[1759]_ ;
  assign \new_[7997]_  = \new_[1756]_  | \new_[1757]_ ;
  assign \new_[7998]_  = \new_[7997]_  | \new_[7994]_ ;
  assign \new_[7999]_  = \new_[7998]_  | \new_[7991]_ ;
  assign \new_[8000]_  = \new_[7999]_  | \new_[7984]_ ;
  assign \new_[8004]_  = \new_[1753]_  | \new_[1754]_ ;
  assign \new_[8005]_  = \new_[1755]_  | \new_[8004]_ ;
  assign \new_[8008]_  = \new_[1751]_  | \new_[1752]_ ;
  assign \new_[8011]_  = \new_[1749]_  | \new_[1750]_ ;
  assign \new_[8012]_  = \new_[8011]_  | \new_[8008]_ ;
  assign \new_[8013]_  = \new_[8012]_  | \new_[8005]_ ;
  assign \new_[8016]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[8019]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[8020]_  = \new_[8019]_  | \new_[8016]_ ;
  assign \new_[8023]_  = \new_[1743]_  | \new_[1744]_ ;
  assign \new_[8026]_  = \new_[1741]_  | \new_[1742]_ ;
  assign \new_[8027]_  = \new_[8026]_  | \new_[8023]_ ;
  assign \new_[8028]_  = \new_[8027]_  | \new_[8020]_ ;
  assign \new_[8029]_  = \new_[8028]_  | \new_[8013]_ ;
  assign \new_[8030]_  = \new_[8029]_  | \new_[8000]_ ;
  assign \new_[8031]_  = \new_[8030]_  | \new_[7971]_ ;
  assign \new_[8035]_  = \new_[1738]_  | \new_[1739]_ ;
  assign \new_[8036]_  = \new_[1740]_  | \new_[8035]_ ;
  assign \new_[8039]_  = \new_[1736]_  | \new_[1737]_ ;
  assign \new_[8042]_  = \new_[1734]_  | \new_[1735]_ ;
  assign \new_[8043]_  = \new_[8042]_  | \new_[8039]_ ;
  assign \new_[8044]_  = \new_[8043]_  | \new_[8036]_ ;
  assign \new_[8047]_  = \new_[1732]_  | \new_[1733]_ ;
  assign \new_[8050]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[8051]_  = \new_[8050]_  | \new_[8047]_ ;
  assign \new_[8054]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[8057]_  = \new_[1726]_  | \new_[1727]_ ;
  assign \new_[8058]_  = \new_[8057]_  | \new_[8054]_ ;
  assign \new_[8059]_  = \new_[8058]_  | \new_[8051]_ ;
  assign \new_[8060]_  = \new_[8059]_  | \new_[8044]_ ;
  assign \new_[8064]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[8065]_  = \new_[1725]_  | \new_[8064]_ ;
  assign \new_[8068]_  = \new_[1721]_  | \new_[1722]_ ;
  assign \new_[8071]_  = \new_[1719]_  | \new_[1720]_ ;
  assign \new_[8072]_  = \new_[8071]_  | \new_[8068]_ ;
  assign \new_[8073]_  = \new_[8072]_  | \new_[8065]_ ;
  assign \new_[8076]_  = \new_[1717]_  | \new_[1718]_ ;
  assign \new_[8079]_  = \new_[1715]_  | \new_[1716]_ ;
  assign \new_[8080]_  = \new_[8079]_  | \new_[8076]_ ;
  assign \new_[8083]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[8086]_  = \new_[1711]_  | \new_[1712]_ ;
  assign \new_[8087]_  = \new_[8086]_  | \new_[8083]_ ;
  assign \new_[8088]_  = \new_[8087]_  | \new_[8080]_ ;
  assign \new_[8089]_  = \new_[8088]_  | \new_[8073]_ ;
  assign \new_[8090]_  = \new_[8089]_  | \new_[8060]_ ;
  assign \new_[8094]_  = \new_[1708]_  | \new_[1709]_ ;
  assign \new_[8095]_  = \new_[1710]_  | \new_[8094]_ ;
  assign \new_[8098]_  = \new_[1706]_  | \new_[1707]_ ;
  assign \new_[8101]_  = \new_[1704]_  | \new_[1705]_ ;
  assign \new_[8102]_  = \new_[8101]_  | \new_[8098]_ ;
  assign \new_[8103]_  = \new_[8102]_  | \new_[8095]_ ;
  assign \new_[8106]_  = \new_[1702]_  | \new_[1703]_ ;
  assign \new_[8109]_  = \new_[1700]_  | \new_[1701]_ ;
  assign \new_[8110]_  = \new_[8109]_  | \new_[8106]_ ;
  assign \new_[8113]_  = \new_[1698]_  | \new_[1699]_ ;
  assign \new_[8116]_  = \new_[1696]_  | \new_[1697]_ ;
  assign \new_[8117]_  = \new_[8116]_  | \new_[8113]_ ;
  assign \new_[8118]_  = \new_[8117]_  | \new_[8110]_ ;
  assign \new_[8119]_  = \new_[8118]_  | \new_[8103]_ ;
  assign \new_[8123]_  = \new_[1693]_  | \new_[1694]_ ;
  assign \new_[8124]_  = \new_[1695]_  | \new_[8123]_ ;
  assign \new_[8127]_  = \new_[1691]_  | \new_[1692]_ ;
  assign \new_[8130]_  = \new_[1689]_  | \new_[1690]_ ;
  assign \new_[8131]_  = \new_[8130]_  | \new_[8127]_ ;
  assign \new_[8132]_  = \new_[8131]_  | \new_[8124]_ ;
  assign \new_[8135]_  = \new_[1687]_  | \new_[1688]_ ;
  assign \new_[8138]_  = \new_[1685]_  | \new_[1686]_ ;
  assign \new_[8139]_  = \new_[8138]_  | \new_[8135]_ ;
  assign \new_[8142]_  = \new_[1683]_  | \new_[1684]_ ;
  assign \new_[8145]_  = \new_[1681]_  | \new_[1682]_ ;
  assign \new_[8146]_  = \new_[8145]_  | \new_[8142]_ ;
  assign \new_[8147]_  = \new_[8146]_  | \new_[8139]_ ;
  assign \new_[8148]_  = \new_[8147]_  | \new_[8132]_ ;
  assign \new_[8149]_  = \new_[8148]_  | \new_[8119]_ ;
  assign \new_[8150]_  = \new_[8149]_  | \new_[8090]_ ;
  assign \new_[8151]_  = \new_[8150]_  | \new_[8031]_ ;
  assign \new_[8152]_  = \new_[8151]_  | \new_[7912]_ ;
  assign \new_[8156]_  = \new_[1678]_  | \new_[1679]_ ;
  assign \new_[8157]_  = \new_[1680]_  | \new_[8156]_ ;
  assign \new_[8160]_  = \new_[1676]_  | \new_[1677]_ ;
  assign \new_[8163]_  = \new_[1674]_  | \new_[1675]_ ;
  assign \new_[8164]_  = \new_[8163]_  | \new_[8160]_ ;
  assign \new_[8165]_  = \new_[8164]_  | \new_[8157]_ ;
  assign \new_[8168]_  = \new_[1672]_  | \new_[1673]_ ;
  assign \new_[8171]_  = \new_[1670]_  | \new_[1671]_ ;
  assign \new_[8172]_  = \new_[8171]_  | \new_[8168]_ ;
  assign \new_[8175]_  = \new_[1668]_  | \new_[1669]_ ;
  assign \new_[8178]_  = \new_[1666]_  | \new_[1667]_ ;
  assign \new_[8179]_  = \new_[8178]_  | \new_[8175]_ ;
  assign \new_[8180]_  = \new_[8179]_  | \new_[8172]_ ;
  assign \new_[8181]_  = \new_[8180]_  | \new_[8165]_ ;
  assign \new_[8185]_  = \new_[1663]_  | \new_[1664]_ ;
  assign \new_[8186]_  = \new_[1665]_  | \new_[8185]_ ;
  assign \new_[8189]_  = \new_[1661]_  | \new_[1662]_ ;
  assign \new_[8192]_  = \new_[1659]_  | \new_[1660]_ ;
  assign \new_[8193]_  = \new_[8192]_  | \new_[8189]_ ;
  assign \new_[8194]_  = \new_[8193]_  | \new_[8186]_ ;
  assign \new_[8197]_  = \new_[1657]_  | \new_[1658]_ ;
  assign \new_[8200]_  = \new_[1655]_  | \new_[1656]_ ;
  assign \new_[8201]_  = \new_[8200]_  | \new_[8197]_ ;
  assign \new_[8204]_  = \new_[1653]_  | \new_[1654]_ ;
  assign \new_[8207]_  = \new_[1651]_  | \new_[1652]_ ;
  assign \new_[8208]_  = \new_[8207]_  | \new_[8204]_ ;
  assign \new_[8209]_  = \new_[8208]_  | \new_[8201]_ ;
  assign \new_[8210]_  = \new_[8209]_  | \new_[8194]_ ;
  assign \new_[8211]_  = \new_[8210]_  | \new_[8181]_ ;
  assign \new_[8215]_  = \new_[1648]_  | \new_[1649]_ ;
  assign \new_[8216]_  = \new_[1650]_  | \new_[8215]_ ;
  assign \new_[8219]_  = \new_[1646]_  | \new_[1647]_ ;
  assign \new_[8222]_  = \new_[1644]_  | \new_[1645]_ ;
  assign \new_[8223]_  = \new_[8222]_  | \new_[8219]_ ;
  assign \new_[8224]_  = \new_[8223]_  | \new_[8216]_ ;
  assign \new_[8227]_  = \new_[1642]_  | \new_[1643]_ ;
  assign \new_[8230]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[8231]_  = \new_[8230]_  | \new_[8227]_ ;
  assign \new_[8234]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[8237]_  = \new_[1636]_  | \new_[1637]_ ;
  assign \new_[8238]_  = \new_[8237]_  | \new_[8234]_ ;
  assign \new_[8239]_  = \new_[8238]_  | \new_[8231]_ ;
  assign \new_[8240]_  = \new_[8239]_  | \new_[8224]_ ;
  assign \new_[8244]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[8245]_  = \new_[1635]_  | \new_[8244]_ ;
  assign \new_[8248]_  = \new_[1631]_  | \new_[1632]_ ;
  assign \new_[8251]_  = \new_[1629]_  | \new_[1630]_ ;
  assign \new_[8252]_  = \new_[8251]_  | \new_[8248]_ ;
  assign \new_[8253]_  = \new_[8252]_  | \new_[8245]_ ;
  assign \new_[8256]_  = \new_[1627]_  | \new_[1628]_ ;
  assign \new_[8259]_  = \new_[1625]_  | \new_[1626]_ ;
  assign \new_[8260]_  = \new_[8259]_  | \new_[8256]_ ;
  assign \new_[8263]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[8266]_  = \new_[1621]_  | \new_[1622]_ ;
  assign \new_[8267]_  = \new_[8266]_  | \new_[8263]_ ;
  assign \new_[8268]_  = \new_[8267]_  | \new_[8260]_ ;
  assign \new_[8269]_  = \new_[8268]_  | \new_[8253]_ ;
  assign \new_[8270]_  = \new_[8269]_  | \new_[8240]_ ;
  assign \new_[8271]_  = \new_[8270]_  | \new_[8211]_ ;
  assign \new_[8275]_  = \new_[1618]_  | \new_[1619]_ ;
  assign \new_[8276]_  = \new_[1620]_  | \new_[8275]_ ;
  assign \new_[8279]_  = \new_[1616]_  | \new_[1617]_ ;
  assign \new_[8282]_  = \new_[1614]_  | \new_[1615]_ ;
  assign \new_[8283]_  = \new_[8282]_  | \new_[8279]_ ;
  assign \new_[8284]_  = \new_[8283]_  | \new_[8276]_ ;
  assign \new_[8287]_  = \new_[1612]_  | \new_[1613]_ ;
  assign \new_[8290]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[8291]_  = \new_[8290]_  | \new_[8287]_ ;
  assign \new_[8294]_  = \new_[1608]_  | \new_[1609]_ ;
  assign \new_[8297]_  = \new_[1606]_  | \new_[1607]_ ;
  assign \new_[8298]_  = \new_[8297]_  | \new_[8294]_ ;
  assign \new_[8299]_  = \new_[8298]_  | \new_[8291]_ ;
  assign \new_[8300]_  = \new_[8299]_  | \new_[8284]_ ;
  assign \new_[8304]_  = \new_[1603]_  | \new_[1604]_ ;
  assign \new_[8305]_  = \new_[1605]_  | \new_[8304]_ ;
  assign \new_[8308]_  = \new_[1601]_  | \new_[1602]_ ;
  assign \new_[8311]_  = \new_[1599]_  | \new_[1600]_ ;
  assign \new_[8312]_  = \new_[8311]_  | \new_[8308]_ ;
  assign \new_[8313]_  = \new_[8312]_  | \new_[8305]_ ;
  assign \new_[8316]_  = \new_[1597]_  | \new_[1598]_ ;
  assign \new_[8319]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[8320]_  = \new_[8319]_  | \new_[8316]_ ;
  assign \new_[8323]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[8326]_  = \new_[1591]_  | \new_[1592]_ ;
  assign \new_[8327]_  = \new_[8326]_  | \new_[8323]_ ;
  assign \new_[8328]_  = \new_[8327]_  | \new_[8320]_ ;
  assign \new_[8329]_  = \new_[8328]_  | \new_[8313]_ ;
  assign \new_[8330]_  = \new_[8329]_  | \new_[8300]_ ;
  assign \new_[8334]_  = \new_[1588]_  | \new_[1589]_ ;
  assign \new_[8335]_  = \new_[1590]_  | \new_[8334]_ ;
  assign \new_[8338]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[8341]_  = \new_[1584]_  | \new_[1585]_ ;
  assign \new_[8342]_  = \new_[8341]_  | \new_[8338]_ ;
  assign \new_[8343]_  = \new_[8342]_  | \new_[8335]_ ;
  assign \new_[8346]_  = \new_[1582]_  | \new_[1583]_ ;
  assign \new_[8349]_  = \new_[1580]_  | \new_[1581]_ ;
  assign \new_[8350]_  = \new_[8349]_  | \new_[8346]_ ;
  assign \new_[8353]_  = \new_[1578]_  | \new_[1579]_ ;
  assign \new_[8356]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[8357]_  = \new_[8356]_  | \new_[8353]_ ;
  assign \new_[8358]_  = \new_[8357]_  | \new_[8350]_ ;
  assign \new_[8359]_  = \new_[8358]_  | \new_[8343]_ ;
  assign \new_[8363]_  = \new_[1573]_  | \new_[1574]_ ;
  assign \new_[8364]_  = \new_[1575]_  | \new_[8363]_ ;
  assign \new_[8367]_  = \new_[1571]_  | \new_[1572]_ ;
  assign \new_[8370]_  = \new_[1569]_  | \new_[1570]_ ;
  assign \new_[8371]_  = \new_[8370]_  | \new_[8367]_ ;
  assign \new_[8372]_  = \new_[8371]_  | \new_[8364]_ ;
  assign \new_[8375]_  = \new_[1567]_  | \new_[1568]_ ;
  assign \new_[8378]_  = \new_[1565]_  | \new_[1566]_ ;
  assign \new_[8379]_  = \new_[8378]_  | \new_[8375]_ ;
  assign \new_[8382]_  = \new_[1563]_  | \new_[1564]_ ;
  assign \new_[8385]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[8386]_  = \new_[8385]_  | \new_[8382]_ ;
  assign \new_[8387]_  = \new_[8386]_  | \new_[8379]_ ;
  assign \new_[8388]_  = \new_[8387]_  | \new_[8372]_ ;
  assign \new_[8389]_  = \new_[8388]_  | \new_[8359]_ ;
  assign \new_[8390]_  = \new_[8389]_  | \new_[8330]_ ;
  assign \new_[8391]_  = \new_[8390]_  | \new_[8271]_ ;
  assign \new_[8395]_  = \new_[1558]_  | \new_[1559]_ ;
  assign \new_[8396]_  = \new_[1560]_  | \new_[8395]_ ;
  assign \new_[8399]_  = \new_[1556]_  | \new_[1557]_ ;
  assign \new_[8402]_  = \new_[1554]_  | \new_[1555]_ ;
  assign \new_[8403]_  = \new_[8402]_  | \new_[8399]_ ;
  assign \new_[8404]_  = \new_[8403]_  | \new_[8396]_ ;
  assign \new_[8407]_  = \new_[1552]_  | \new_[1553]_ ;
  assign \new_[8410]_  = \new_[1550]_  | \new_[1551]_ ;
  assign \new_[8411]_  = \new_[8410]_  | \new_[8407]_ ;
  assign \new_[8414]_  = \new_[1548]_  | \new_[1549]_ ;
  assign \new_[8417]_  = \new_[1546]_  | \new_[1547]_ ;
  assign \new_[8418]_  = \new_[8417]_  | \new_[8414]_ ;
  assign \new_[8419]_  = \new_[8418]_  | \new_[8411]_ ;
  assign \new_[8420]_  = \new_[8419]_  | \new_[8404]_ ;
  assign \new_[8424]_  = \new_[1543]_  | \new_[1544]_ ;
  assign \new_[8425]_  = \new_[1545]_  | \new_[8424]_ ;
  assign \new_[8428]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[8431]_  = \new_[1539]_  | \new_[1540]_ ;
  assign \new_[8432]_  = \new_[8431]_  | \new_[8428]_ ;
  assign \new_[8433]_  = \new_[8432]_  | \new_[8425]_ ;
  assign \new_[8436]_  = \new_[1537]_  | \new_[1538]_ ;
  assign \new_[8439]_  = \new_[1535]_  | \new_[1536]_ ;
  assign \new_[8440]_  = \new_[8439]_  | \new_[8436]_ ;
  assign \new_[8443]_  = \new_[1533]_  | \new_[1534]_ ;
  assign \new_[8446]_  = \new_[1531]_  | \new_[1532]_ ;
  assign \new_[8447]_  = \new_[8446]_  | \new_[8443]_ ;
  assign \new_[8448]_  = \new_[8447]_  | \new_[8440]_ ;
  assign \new_[8449]_  = \new_[8448]_  | \new_[8433]_ ;
  assign \new_[8450]_  = \new_[8449]_  | \new_[8420]_ ;
  assign \new_[8454]_  = \new_[1528]_  | \new_[1529]_ ;
  assign \new_[8455]_  = \new_[1530]_  | \new_[8454]_ ;
  assign \new_[8458]_  = \new_[1526]_  | \new_[1527]_ ;
  assign \new_[8461]_  = \new_[1524]_  | \new_[1525]_ ;
  assign \new_[8462]_  = \new_[8461]_  | \new_[8458]_ ;
  assign \new_[8463]_  = \new_[8462]_  | \new_[8455]_ ;
  assign \new_[8466]_  = \new_[1522]_  | \new_[1523]_ ;
  assign \new_[8469]_  = \new_[1520]_  | \new_[1521]_ ;
  assign \new_[8470]_  = \new_[8469]_  | \new_[8466]_ ;
  assign \new_[8473]_  = \new_[1518]_  | \new_[1519]_ ;
  assign \new_[8476]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[8477]_  = \new_[8476]_  | \new_[8473]_ ;
  assign \new_[8478]_  = \new_[8477]_  | \new_[8470]_ ;
  assign \new_[8479]_  = \new_[8478]_  | \new_[8463]_ ;
  assign \new_[8483]_  = \new_[1513]_  | \new_[1514]_ ;
  assign \new_[8484]_  = \new_[1515]_  | \new_[8483]_ ;
  assign \new_[8487]_  = \new_[1511]_  | \new_[1512]_ ;
  assign \new_[8490]_  = \new_[1509]_  | \new_[1510]_ ;
  assign \new_[8491]_  = \new_[8490]_  | \new_[8487]_ ;
  assign \new_[8492]_  = \new_[8491]_  | \new_[8484]_ ;
  assign \new_[8495]_  = \new_[1507]_  | \new_[1508]_ ;
  assign \new_[8498]_  = \new_[1505]_  | \new_[1506]_ ;
  assign \new_[8499]_  = \new_[8498]_  | \new_[8495]_ ;
  assign \new_[8502]_  = \new_[1503]_  | \new_[1504]_ ;
  assign \new_[8505]_  = \new_[1501]_  | \new_[1502]_ ;
  assign \new_[8506]_  = \new_[8505]_  | \new_[8502]_ ;
  assign \new_[8507]_  = \new_[8506]_  | \new_[8499]_ ;
  assign \new_[8508]_  = \new_[8507]_  | \new_[8492]_ ;
  assign \new_[8509]_  = \new_[8508]_  | \new_[8479]_ ;
  assign \new_[8510]_  = \new_[8509]_  | \new_[8450]_ ;
  assign \new_[8514]_  = \new_[1498]_  | \new_[1499]_ ;
  assign \new_[8515]_  = \new_[1500]_  | \new_[8514]_ ;
  assign \new_[8518]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[8521]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[8522]_  = \new_[8521]_  | \new_[8518]_ ;
  assign \new_[8523]_  = \new_[8522]_  | \new_[8515]_ ;
  assign \new_[8526]_  = \new_[1492]_  | \new_[1493]_ ;
  assign \new_[8529]_  = \new_[1490]_  | \new_[1491]_ ;
  assign \new_[8530]_  = \new_[8529]_  | \new_[8526]_ ;
  assign \new_[8533]_  = \new_[1488]_  | \new_[1489]_ ;
  assign \new_[8536]_  = \new_[1486]_  | \new_[1487]_ ;
  assign \new_[8537]_  = \new_[8536]_  | \new_[8533]_ ;
  assign \new_[8538]_  = \new_[8537]_  | \new_[8530]_ ;
  assign \new_[8539]_  = \new_[8538]_  | \new_[8523]_ ;
  assign \new_[8543]_  = \new_[1483]_  | \new_[1484]_ ;
  assign \new_[8544]_  = \new_[1485]_  | \new_[8543]_ ;
  assign \new_[8547]_  = \new_[1481]_  | \new_[1482]_ ;
  assign \new_[8550]_  = \new_[1479]_  | \new_[1480]_ ;
  assign \new_[8551]_  = \new_[8550]_  | \new_[8547]_ ;
  assign \new_[8552]_  = \new_[8551]_  | \new_[8544]_ ;
  assign \new_[8555]_  = \new_[1477]_  | \new_[1478]_ ;
  assign \new_[8558]_  = \new_[1475]_  | \new_[1476]_ ;
  assign \new_[8559]_  = \new_[8558]_  | \new_[8555]_ ;
  assign \new_[8562]_  = \new_[1473]_  | \new_[1474]_ ;
  assign \new_[8565]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[8566]_  = \new_[8565]_  | \new_[8562]_ ;
  assign \new_[8567]_  = \new_[8566]_  | \new_[8559]_ ;
  assign \new_[8568]_  = \new_[8567]_  | \new_[8552]_ ;
  assign \new_[8569]_  = \new_[8568]_  | \new_[8539]_ ;
  assign \new_[8573]_  = \new_[1468]_  | \new_[1469]_ ;
  assign \new_[8574]_  = \new_[1470]_  | \new_[8573]_ ;
  assign \new_[8577]_  = \new_[1466]_  | \new_[1467]_ ;
  assign \new_[8580]_  = \new_[1464]_  | \new_[1465]_ ;
  assign \new_[8581]_  = \new_[8580]_  | \new_[8577]_ ;
  assign \new_[8582]_  = \new_[8581]_  | \new_[8574]_ ;
  assign \new_[8585]_  = \new_[1462]_  | \new_[1463]_ ;
  assign \new_[8588]_  = \new_[1460]_  | \new_[1461]_ ;
  assign \new_[8589]_  = \new_[8588]_  | \new_[8585]_ ;
  assign \new_[8592]_  = \new_[1458]_  | \new_[1459]_ ;
  assign \new_[8595]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[8596]_  = \new_[8595]_  | \new_[8592]_ ;
  assign \new_[8597]_  = \new_[8596]_  | \new_[8589]_ ;
  assign \new_[8598]_  = \new_[8597]_  | \new_[8582]_ ;
  assign \new_[8602]_  = \new_[1453]_  | \new_[1454]_ ;
  assign \new_[8603]_  = \new_[1455]_  | \new_[8602]_ ;
  assign \new_[8606]_  = \new_[1451]_  | \new_[1452]_ ;
  assign \new_[8609]_  = \new_[1449]_  | \new_[1450]_ ;
  assign \new_[8610]_  = \new_[8609]_  | \new_[8606]_ ;
  assign \new_[8611]_  = \new_[8610]_  | \new_[8603]_ ;
  assign \new_[8614]_  = \new_[1447]_  | \new_[1448]_ ;
  assign \new_[8617]_  = \new_[1445]_  | \new_[1446]_ ;
  assign \new_[8618]_  = \new_[8617]_  | \new_[8614]_ ;
  assign \new_[8621]_  = \new_[1443]_  | \new_[1444]_ ;
  assign \new_[8624]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[8625]_  = \new_[8624]_  | \new_[8621]_ ;
  assign \new_[8626]_  = \new_[8625]_  | \new_[8618]_ ;
  assign \new_[8627]_  = \new_[8626]_  | \new_[8611]_ ;
  assign \new_[8628]_  = \new_[8627]_  | \new_[8598]_ ;
  assign \new_[8629]_  = \new_[8628]_  | \new_[8569]_ ;
  assign \new_[8630]_  = \new_[8629]_  | \new_[8510]_ ;
  assign \new_[8631]_  = \new_[8630]_  | \new_[8391]_ ;
  assign \new_[8632]_  = \new_[8631]_  | \new_[8152]_ ;
  assign \new_[8636]_  = \new_[1438]_  | \new_[1439]_ ;
  assign \new_[8637]_  = \new_[1440]_  | \new_[8636]_ ;
  assign \new_[8640]_  = \new_[1436]_  | \new_[1437]_ ;
  assign \new_[8643]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[8644]_  = \new_[8643]_  | \new_[8640]_ ;
  assign \new_[8645]_  = \new_[8644]_  | \new_[8637]_ ;
  assign \new_[8648]_  = \new_[1432]_  | \new_[1433]_ ;
  assign \new_[8651]_  = \new_[1430]_  | \new_[1431]_ ;
  assign \new_[8652]_  = \new_[8651]_  | \new_[8648]_ ;
  assign \new_[8655]_  = \new_[1428]_  | \new_[1429]_ ;
  assign \new_[8658]_  = \new_[1426]_  | \new_[1427]_ ;
  assign \new_[8659]_  = \new_[8658]_  | \new_[8655]_ ;
  assign \new_[8660]_  = \new_[8659]_  | \new_[8652]_ ;
  assign \new_[8661]_  = \new_[8660]_  | \new_[8645]_ ;
  assign \new_[8665]_  = \new_[1423]_  | \new_[1424]_ ;
  assign \new_[8666]_  = \new_[1425]_  | \new_[8665]_ ;
  assign \new_[8669]_  = \new_[1421]_  | \new_[1422]_ ;
  assign \new_[8672]_  = \new_[1419]_  | \new_[1420]_ ;
  assign \new_[8673]_  = \new_[8672]_  | \new_[8669]_ ;
  assign \new_[8674]_  = \new_[8673]_  | \new_[8666]_ ;
  assign \new_[8677]_  = \new_[1417]_  | \new_[1418]_ ;
  assign \new_[8680]_  = \new_[1415]_  | \new_[1416]_ ;
  assign \new_[8681]_  = \new_[8680]_  | \new_[8677]_ ;
  assign \new_[8684]_  = \new_[1413]_  | \new_[1414]_ ;
  assign \new_[8687]_  = \new_[1411]_  | \new_[1412]_ ;
  assign \new_[8688]_  = \new_[8687]_  | \new_[8684]_ ;
  assign \new_[8689]_  = \new_[8688]_  | \new_[8681]_ ;
  assign \new_[8690]_  = \new_[8689]_  | \new_[8674]_ ;
  assign \new_[8691]_  = \new_[8690]_  | \new_[8661]_ ;
  assign \new_[8695]_  = \new_[1408]_  | \new_[1409]_ ;
  assign \new_[8696]_  = \new_[1410]_  | \new_[8695]_ ;
  assign \new_[8699]_  = \new_[1406]_  | \new_[1407]_ ;
  assign \new_[8702]_  = \new_[1404]_  | \new_[1405]_ ;
  assign \new_[8703]_  = \new_[8702]_  | \new_[8699]_ ;
  assign \new_[8704]_  = \new_[8703]_  | \new_[8696]_ ;
  assign \new_[8707]_  = \new_[1402]_  | \new_[1403]_ ;
  assign \new_[8710]_  = \new_[1400]_  | \new_[1401]_ ;
  assign \new_[8711]_  = \new_[8710]_  | \new_[8707]_ ;
  assign \new_[8714]_  = \new_[1398]_  | \new_[1399]_ ;
  assign \new_[8717]_  = \new_[1396]_  | \new_[1397]_ ;
  assign \new_[8718]_  = \new_[8717]_  | \new_[8714]_ ;
  assign \new_[8719]_  = \new_[8718]_  | \new_[8711]_ ;
  assign \new_[8720]_  = \new_[8719]_  | \new_[8704]_ ;
  assign \new_[8724]_  = \new_[1393]_  | \new_[1394]_ ;
  assign \new_[8725]_  = \new_[1395]_  | \new_[8724]_ ;
  assign \new_[8728]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[8731]_  = \new_[1389]_  | \new_[1390]_ ;
  assign \new_[8732]_  = \new_[8731]_  | \new_[8728]_ ;
  assign \new_[8733]_  = \new_[8732]_  | \new_[8725]_ ;
  assign \new_[8736]_  = \new_[1387]_  | \new_[1388]_ ;
  assign \new_[8739]_  = \new_[1385]_  | \new_[1386]_ ;
  assign \new_[8740]_  = \new_[8739]_  | \new_[8736]_ ;
  assign \new_[8743]_  = \new_[1383]_  | \new_[1384]_ ;
  assign \new_[8746]_  = \new_[1381]_  | \new_[1382]_ ;
  assign \new_[8747]_  = \new_[8746]_  | \new_[8743]_ ;
  assign \new_[8748]_  = \new_[8747]_  | \new_[8740]_ ;
  assign \new_[8749]_  = \new_[8748]_  | \new_[8733]_ ;
  assign \new_[8750]_  = \new_[8749]_  | \new_[8720]_ ;
  assign \new_[8751]_  = \new_[8750]_  | \new_[8691]_ ;
  assign \new_[8755]_  = \new_[1378]_  | \new_[1379]_ ;
  assign \new_[8756]_  = \new_[1380]_  | \new_[8755]_ ;
  assign \new_[8759]_  = \new_[1376]_  | \new_[1377]_ ;
  assign \new_[8762]_  = \new_[1374]_  | \new_[1375]_ ;
  assign \new_[8763]_  = \new_[8762]_  | \new_[8759]_ ;
  assign \new_[8764]_  = \new_[8763]_  | \new_[8756]_ ;
  assign \new_[8767]_  = \new_[1372]_  | \new_[1373]_ ;
  assign \new_[8770]_  = \new_[1370]_  | \new_[1371]_ ;
  assign \new_[8771]_  = \new_[8770]_  | \new_[8767]_ ;
  assign \new_[8774]_  = \new_[1368]_  | \new_[1369]_ ;
  assign \new_[8777]_  = \new_[1366]_  | \new_[1367]_ ;
  assign \new_[8778]_  = \new_[8777]_  | \new_[8774]_ ;
  assign \new_[8779]_  = \new_[8778]_  | \new_[8771]_ ;
  assign \new_[8780]_  = \new_[8779]_  | \new_[8764]_ ;
  assign \new_[8784]_  = \new_[1363]_  | \new_[1364]_ ;
  assign \new_[8785]_  = \new_[1365]_  | \new_[8784]_ ;
  assign \new_[8788]_  = \new_[1361]_  | \new_[1362]_ ;
  assign \new_[8791]_  = \new_[1359]_  | \new_[1360]_ ;
  assign \new_[8792]_  = \new_[8791]_  | \new_[8788]_ ;
  assign \new_[8793]_  = \new_[8792]_  | \new_[8785]_ ;
  assign \new_[8796]_  = \new_[1357]_  | \new_[1358]_ ;
  assign \new_[8799]_  = \new_[1355]_  | \new_[1356]_ ;
  assign \new_[8800]_  = \new_[8799]_  | \new_[8796]_ ;
  assign \new_[8803]_  = \new_[1353]_  | \new_[1354]_ ;
  assign \new_[8806]_  = \new_[1351]_  | \new_[1352]_ ;
  assign \new_[8807]_  = \new_[8806]_  | \new_[8803]_ ;
  assign \new_[8808]_  = \new_[8807]_  | \new_[8800]_ ;
  assign \new_[8809]_  = \new_[8808]_  | \new_[8793]_ ;
  assign \new_[8810]_  = \new_[8809]_  | \new_[8780]_ ;
  assign \new_[8814]_  = \new_[1348]_  | \new_[1349]_ ;
  assign \new_[8815]_  = \new_[1350]_  | \new_[8814]_ ;
  assign \new_[8818]_  = \new_[1346]_  | \new_[1347]_ ;
  assign \new_[8821]_  = \new_[1344]_  | \new_[1345]_ ;
  assign \new_[8822]_  = \new_[8821]_  | \new_[8818]_ ;
  assign \new_[8823]_  = \new_[8822]_  | \new_[8815]_ ;
  assign \new_[8826]_  = \new_[1342]_  | \new_[1343]_ ;
  assign \new_[8829]_  = \new_[1340]_  | \new_[1341]_ ;
  assign \new_[8830]_  = \new_[8829]_  | \new_[8826]_ ;
  assign \new_[8833]_  = \new_[1338]_  | \new_[1339]_ ;
  assign \new_[8836]_  = \new_[1336]_  | \new_[1337]_ ;
  assign \new_[8837]_  = \new_[8836]_  | \new_[8833]_ ;
  assign \new_[8838]_  = \new_[8837]_  | \new_[8830]_ ;
  assign \new_[8839]_  = \new_[8838]_  | \new_[8823]_ ;
  assign \new_[8843]_  = \new_[1333]_  | \new_[1334]_ ;
  assign \new_[8844]_  = \new_[1335]_  | \new_[8843]_ ;
  assign \new_[8847]_  = \new_[1331]_  | \new_[1332]_ ;
  assign \new_[8850]_  = \new_[1329]_  | \new_[1330]_ ;
  assign \new_[8851]_  = \new_[8850]_  | \new_[8847]_ ;
  assign \new_[8852]_  = \new_[8851]_  | \new_[8844]_ ;
  assign \new_[8855]_  = \new_[1327]_  | \new_[1328]_ ;
  assign \new_[8858]_  = \new_[1325]_  | \new_[1326]_ ;
  assign \new_[8859]_  = \new_[8858]_  | \new_[8855]_ ;
  assign \new_[8862]_  = \new_[1323]_  | \new_[1324]_ ;
  assign \new_[8865]_  = \new_[1321]_  | \new_[1322]_ ;
  assign \new_[8866]_  = \new_[8865]_  | \new_[8862]_ ;
  assign \new_[8867]_  = \new_[8866]_  | \new_[8859]_ ;
  assign \new_[8868]_  = \new_[8867]_  | \new_[8852]_ ;
  assign \new_[8869]_  = \new_[8868]_  | \new_[8839]_ ;
  assign \new_[8870]_  = \new_[8869]_  | \new_[8810]_ ;
  assign \new_[8871]_  = \new_[8870]_  | \new_[8751]_ ;
  assign \new_[8875]_  = \new_[1318]_  | \new_[1319]_ ;
  assign \new_[8876]_  = \new_[1320]_  | \new_[8875]_ ;
  assign \new_[8879]_  = \new_[1316]_  | \new_[1317]_ ;
  assign \new_[8882]_  = \new_[1314]_  | \new_[1315]_ ;
  assign \new_[8883]_  = \new_[8882]_  | \new_[8879]_ ;
  assign \new_[8884]_  = \new_[8883]_  | \new_[8876]_ ;
  assign \new_[8887]_  = \new_[1312]_  | \new_[1313]_ ;
  assign \new_[8890]_  = \new_[1310]_  | \new_[1311]_ ;
  assign \new_[8891]_  = \new_[8890]_  | \new_[8887]_ ;
  assign \new_[8894]_  = \new_[1308]_  | \new_[1309]_ ;
  assign \new_[8897]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[8898]_  = \new_[8897]_  | \new_[8894]_ ;
  assign \new_[8899]_  = \new_[8898]_  | \new_[8891]_ ;
  assign \new_[8900]_  = \new_[8899]_  | \new_[8884]_ ;
  assign \new_[8904]_  = \new_[1303]_  | \new_[1304]_ ;
  assign \new_[8905]_  = \new_[1305]_  | \new_[8904]_ ;
  assign \new_[8908]_  = \new_[1301]_  | \new_[1302]_ ;
  assign \new_[8911]_  = \new_[1299]_  | \new_[1300]_ ;
  assign \new_[8912]_  = \new_[8911]_  | \new_[8908]_ ;
  assign \new_[8913]_  = \new_[8912]_  | \new_[8905]_ ;
  assign \new_[8916]_  = \new_[1297]_  | \new_[1298]_ ;
  assign \new_[8919]_  = \new_[1295]_  | \new_[1296]_ ;
  assign \new_[8920]_  = \new_[8919]_  | \new_[8916]_ ;
  assign \new_[8923]_  = \new_[1293]_  | \new_[1294]_ ;
  assign \new_[8926]_  = \new_[1291]_  | \new_[1292]_ ;
  assign \new_[8927]_  = \new_[8926]_  | \new_[8923]_ ;
  assign \new_[8928]_  = \new_[8927]_  | \new_[8920]_ ;
  assign \new_[8929]_  = \new_[8928]_  | \new_[8913]_ ;
  assign \new_[8930]_  = \new_[8929]_  | \new_[8900]_ ;
  assign \new_[8934]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[8935]_  = \new_[1290]_  | \new_[8934]_ ;
  assign \new_[8938]_  = \new_[1286]_  | \new_[1287]_ ;
  assign \new_[8941]_  = \new_[1284]_  | \new_[1285]_ ;
  assign \new_[8942]_  = \new_[8941]_  | \new_[8938]_ ;
  assign \new_[8943]_  = \new_[8942]_  | \new_[8935]_ ;
  assign \new_[8946]_  = \new_[1282]_  | \new_[1283]_ ;
  assign \new_[8949]_  = \new_[1280]_  | \new_[1281]_ ;
  assign \new_[8950]_  = \new_[8949]_  | \new_[8946]_ ;
  assign \new_[8953]_  = \new_[1278]_  | \new_[1279]_ ;
  assign \new_[8956]_  = \new_[1276]_  | \new_[1277]_ ;
  assign \new_[8957]_  = \new_[8956]_  | \new_[8953]_ ;
  assign \new_[8958]_  = \new_[8957]_  | \new_[8950]_ ;
  assign \new_[8959]_  = \new_[8958]_  | \new_[8943]_ ;
  assign \new_[8963]_  = \new_[1273]_  | \new_[1274]_ ;
  assign \new_[8964]_  = \new_[1275]_  | \new_[8963]_ ;
  assign \new_[8967]_  = \new_[1271]_  | \new_[1272]_ ;
  assign \new_[8970]_  = \new_[1269]_  | \new_[1270]_ ;
  assign \new_[8971]_  = \new_[8970]_  | \new_[8967]_ ;
  assign \new_[8972]_  = \new_[8971]_  | \new_[8964]_ ;
  assign \new_[8975]_  = \new_[1267]_  | \new_[1268]_ ;
  assign \new_[8978]_  = \new_[1265]_  | \new_[1266]_ ;
  assign \new_[8979]_  = \new_[8978]_  | \new_[8975]_ ;
  assign \new_[8982]_  = \new_[1263]_  | \new_[1264]_ ;
  assign \new_[8985]_  = \new_[1261]_  | \new_[1262]_ ;
  assign \new_[8986]_  = \new_[8985]_  | \new_[8982]_ ;
  assign \new_[8987]_  = \new_[8986]_  | \new_[8979]_ ;
  assign \new_[8988]_  = \new_[8987]_  | \new_[8972]_ ;
  assign \new_[8989]_  = \new_[8988]_  | \new_[8959]_ ;
  assign \new_[8990]_  = \new_[8989]_  | \new_[8930]_ ;
  assign \new_[8994]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[8995]_  = \new_[1260]_  | \new_[8994]_ ;
  assign \new_[8998]_  = \new_[1256]_  | \new_[1257]_ ;
  assign \new_[9001]_  = \new_[1254]_  | \new_[1255]_ ;
  assign \new_[9002]_  = \new_[9001]_  | \new_[8998]_ ;
  assign \new_[9003]_  = \new_[9002]_  | \new_[8995]_ ;
  assign \new_[9006]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[9009]_  = \new_[1250]_  | \new_[1251]_ ;
  assign \new_[9010]_  = \new_[9009]_  | \new_[9006]_ ;
  assign \new_[9013]_  = \new_[1248]_  | \new_[1249]_ ;
  assign \new_[9016]_  = \new_[1246]_  | \new_[1247]_ ;
  assign \new_[9017]_  = \new_[9016]_  | \new_[9013]_ ;
  assign \new_[9018]_  = \new_[9017]_  | \new_[9010]_ ;
  assign \new_[9019]_  = \new_[9018]_  | \new_[9003]_ ;
  assign \new_[9023]_  = \new_[1243]_  | \new_[1244]_ ;
  assign \new_[9024]_  = \new_[1245]_  | \new_[9023]_ ;
  assign \new_[9027]_  = \new_[1241]_  | \new_[1242]_ ;
  assign \new_[9030]_  = \new_[1239]_  | \new_[1240]_ ;
  assign \new_[9031]_  = \new_[9030]_  | \new_[9027]_ ;
  assign \new_[9032]_  = \new_[9031]_  | \new_[9024]_ ;
  assign \new_[9035]_  = \new_[1237]_  | \new_[1238]_ ;
  assign \new_[9038]_  = \new_[1235]_  | \new_[1236]_ ;
  assign \new_[9039]_  = \new_[9038]_  | \new_[9035]_ ;
  assign \new_[9042]_  = \new_[1233]_  | \new_[1234]_ ;
  assign \new_[9045]_  = \new_[1231]_  | \new_[1232]_ ;
  assign \new_[9046]_  = \new_[9045]_  | \new_[9042]_ ;
  assign \new_[9047]_  = \new_[9046]_  | \new_[9039]_ ;
  assign \new_[9048]_  = \new_[9047]_  | \new_[9032]_ ;
  assign \new_[9049]_  = \new_[9048]_  | \new_[9019]_ ;
  assign \new_[9053]_  = \new_[1228]_  | \new_[1229]_ ;
  assign \new_[9054]_  = \new_[1230]_  | \new_[9053]_ ;
  assign \new_[9057]_  = \new_[1226]_  | \new_[1227]_ ;
  assign \new_[9060]_  = \new_[1224]_  | \new_[1225]_ ;
  assign \new_[9061]_  = \new_[9060]_  | \new_[9057]_ ;
  assign \new_[9062]_  = \new_[9061]_  | \new_[9054]_ ;
  assign \new_[9065]_  = \new_[1222]_  | \new_[1223]_ ;
  assign \new_[9068]_  = \new_[1220]_  | \new_[1221]_ ;
  assign \new_[9069]_  = \new_[9068]_  | \new_[9065]_ ;
  assign \new_[9072]_  = \new_[1218]_  | \new_[1219]_ ;
  assign \new_[9075]_  = \new_[1216]_  | \new_[1217]_ ;
  assign \new_[9076]_  = \new_[9075]_  | \new_[9072]_ ;
  assign \new_[9077]_  = \new_[9076]_  | \new_[9069]_ ;
  assign \new_[9078]_  = \new_[9077]_  | \new_[9062]_ ;
  assign \new_[9082]_  = \new_[1213]_  | \new_[1214]_ ;
  assign \new_[9083]_  = \new_[1215]_  | \new_[9082]_ ;
  assign \new_[9086]_  = \new_[1211]_  | \new_[1212]_ ;
  assign \new_[9089]_  = \new_[1209]_  | \new_[1210]_ ;
  assign \new_[9090]_  = \new_[9089]_  | \new_[9086]_ ;
  assign \new_[9091]_  = \new_[9090]_  | \new_[9083]_ ;
  assign \new_[9094]_  = \new_[1207]_  | \new_[1208]_ ;
  assign \new_[9097]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[9098]_  = \new_[9097]_  | \new_[9094]_ ;
  assign \new_[9101]_  = \new_[1203]_  | \new_[1204]_ ;
  assign \new_[9104]_  = \new_[1201]_  | \new_[1202]_ ;
  assign \new_[9105]_  = \new_[9104]_  | \new_[9101]_ ;
  assign \new_[9106]_  = \new_[9105]_  | \new_[9098]_ ;
  assign \new_[9107]_  = \new_[9106]_  | \new_[9091]_ ;
  assign \new_[9108]_  = \new_[9107]_  | \new_[9078]_ ;
  assign \new_[9109]_  = \new_[9108]_  | \new_[9049]_ ;
  assign \new_[9110]_  = \new_[9109]_  | \new_[8990]_ ;
  assign \new_[9111]_  = \new_[9110]_  | \new_[8871]_ ;
  assign \new_[9115]_  = \new_[1198]_  | \new_[1199]_ ;
  assign \new_[9116]_  = \new_[1200]_  | \new_[9115]_ ;
  assign \new_[9119]_  = \new_[1196]_  | \new_[1197]_ ;
  assign \new_[9122]_  = \new_[1194]_  | \new_[1195]_ ;
  assign \new_[9123]_  = \new_[9122]_  | \new_[9119]_ ;
  assign \new_[9124]_  = \new_[9123]_  | \new_[9116]_ ;
  assign \new_[9127]_  = \new_[1192]_  | \new_[1193]_ ;
  assign \new_[9130]_  = \new_[1190]_  | \new_[1191]_ ;
  assign \new_[9131]_  = \new_[9130]_  | \new_[9127]_ ;
  assign \new_[9134]_  = \new_[1188]_  | \new_[1189]_ ;
  assign \new_[9137]_  = \new_[1186]_  | \new_[1187]_ ;
  assign \new_[9138]_  = \new_[9137]_  | \new_[9134]_ ;
  assign \new_[9139]_  = \new_[9138]_  | \new_[9131]_ ;
  assign \new_[9140]_  = \new_[9139]_  | \new_[9124]_ ;
  assign \new_[9144]_  = \new_[1183]_  | \new_[1184]_ ;
  assign \new_[9145]_  = \new_[1185]_  | \new_[9144]_ ;
  assign \new_[9148]_  = \new_[1181]_  | \new_[1182]_ ;
  assign \new_[9151]_  = \new_[1179]_  | \new_[1180]_ ;
  assign \new_[9152]_  = \new_[9151]_  | \new_[9148]_ ;
  assign \new_[9153]_  = \new_[9152]_  | \new_[9145]_ ;
  assign \new_[9156]_  = \new_[1177]_  | \new_[1178]_ ;
  assign \new_[9159]_  = \new_[1175]_  | \new_[1176]_ ;
  assign \new_[9160]_  = \new_[9159]_  | \new_[9156]_ ;
  assign \new_[9163]_  = \new_[1173]_  | \new_[1174]_ ;
  assign \new_[9166]_  = \new_[1171]_  | \new_[1172]_ ;
  assign \new_[9167]_  = \new_[9166]_  | \new_[9163]_ ;
  assign \new_[9168]_  = \new_[9167]_  | \new_[9160]_ ;
  assign \new_[9169]_  = \new_[9168]_  | \new_[9153]_ ;
  assign \new_[9170]_  = \new_[9169]_  | \new_[9140]_ ;
  assign \new_[9174]_  = \new_[1168]_  | \new_[1169]_ ;
  assign \new_[9175]_  = \new_[1170]_  | \new_[9174]_ ;
  assign \new_[9178]_  = \new_[1166]_  | \new_[1167]_ ;
  assign \new_[9181]_  = \new_[1164]_  | \new_[1165]_ ;
  assign \new_[9182]_  = \new_[9181]_  | \new_[9178]_ ;
  assign \new_[9183]_  = \new_[9182]_  | \new_[9175]_ ;
  assign \new_[9186]_  = \new_[1162]_  | \new_[1163]_ ;
  assign \new_[9189]_  = \new_[1160]_  | \new_[1161]_ ;
  assign \new_[9190]_  = \new_[9189]_  | \new_[9186]_ ;
  assign \new_[9193]_  = \new_[1158]_  | \new_[1159]_ ;
  assign \new_[9196]_  = \new_[1156]_  | \new_[1157]_ ;
  assign \new_[9197]_  = \new_[9196]_  | \new_[9193]_ ;
  assign \new_[9198]_  = \new_[9197]_  | \new_[9190]_ ;
  assign \new_[9199]_  = \new_[9198]_  | \new_[9183]_ ;
  assign \new_[9203]_  = \new_[1153]_  | \new_[1154]_ ;
  assign \new_[9204]_  = \new_[1155]_  | \new_[9203]_ ;
  assign \new_[9207]_  = \new_[1151]_  | \new_[1152]_ ;
  assign \new_[9210]_  = \new_[1149]_  | \new_[1150]_ ;
  assign \new_[9211]_  = \new_[9210]_  | \new_[9207]_ ;
  assign \new_[9212]_  = \new_[9211]_  | \new_[9204]_ ;
  assign \new_[9215]_  = \new_[1147]_  | \new_[1148]_ ;
  assign \new_[9218]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[9219]_  = \new_[9218]_  | \new_[9215]_ ;
  assign \new_[9222]_  = \new_[1143]_  | \new_[1144]_ ;
  assign \new_[9225]_  = \new_[1141]_  | \new_[1142]_ ;
  assign \new_[9226]_  = \new_[9225]_  | \new_[9222]_ ;
  assign \new_[9227]_  = \new_[9226]_  | \new_[9219]_ ;
  assign \new_[9228]_  = \new_[9227]_  | \new_[9212]_ ;
  assign \new_[9229]_  = \new_[9228]_  | \new_[9199]_ ;
  assign \new_[9230]_  = \new_[9229]_  | \new_[9170]_ ;
  assign \new_[9234]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[9235]_  = \new_[1140]_  | \new_[9234]_ ;
  assign \new_[9238]_  = \new_[1136]_  | \new_[1137]_ ;
  assign \new_[9241]_  = \new_[1134]_  | \new_[1135]_ ;
  assign \new_[9242]_  = \new_[9241]_  | \new_[9238]_ ;
  assign \new_[9243]_  = \new_[9242]_  | \new_[9235]_ ;
  assign \new_[9246]_  = \new_[1132]_  | \new_[1133]_ ;
  assign \new_[9249]_  = \new_[1130]_  | \new_[1131]_ ;
  assign \new_[9250]_  = \new_[9249]_  | \new_[9246]_ ;
  assign \new_[9253]_  = \new_[1128]_  | \new_[1129]_ ;
  assign \new_[9256]_  = \new_[1126]_  | \new_[1127]_ ;
  assign \new_[9257]_  = \new_[9256]_  | \new_[9253]_ ;
  assign \new_[9258]_  = \new_[9257]_  | \new_[9250]_ ;
  assign \new_[9259]_  = \new_[9258]_  | \new_[9243]_ ;
  assign \new_[9263]_  = \new_[1123]_  | \new_[1124]_ ;
  assign \new_[9264]_  = \new_[1125]_  | \new_[9263]_ ;
  assign \new_[9267]_  = \new_[1121]_  | \new_[1122]_ ;
  assign \new_[9270]_  = \new_[1119]_  | \new_[1120]_ ;
  assign \new_[9271]_  = \new_[9270]_  | \new_[9267]_ ;
  assign \new_[9272]_  = \new_[9271]_  | \new_[9264]_ ;
  assign \new_[9275]_  = \new_[1117]_  | \new_[1118]_ ;
  assign \new_[9278]_  = \new_[1115]_  | \new_[1116]_ ;
  assign \new_[9279]_  = \new_[9278]_  | \new_[9275]_ ;
  assign \new_[9282]_  = \new_[1113]_  | \new_[1114]_ ;
  assign \new_[9285]_  = \new_[1111]_  | \new_[1112]_ ;
  assign \new_[9286]_  = \new_[9285]_  | \new_[9282]_ ;
  assign \new_[9287]_  = \new_[9286]_  | \new_[9279]_ ;
  assign \new_[9288]_  = \new_[9287]_  | \new_[9272]_ ;
  assign \new_[9289]_  = \new_[9288]_  | \new_[9259]_ ;
  assign \new_[9293]_  = \new_[1108]_  | \new_[1109]_ ;
  assign \new_[9294]_  = \new_[1110]_  | \new_[9293]_ ;
  assign \new_[9297]_  = \new_[1106]_  | \new_[1107]_ ;
  assign \new_[9300]_  = \new_[1104]_  | \new_[1105]_ ;
  assign \new_[9301]_  = \new_[9300]_  | \new_[9297]_ ;
  assign \new_[9302]_  = \new_[9301]_  | \new_[9294]_ ;
  assign \new_[9305]_  = \new_[1102]_  | \new_[1103]_ ;
  assign \new_[9308]_  = \new_[1100]_  | \new_[1101]_ ;
  assign \new_[9309]_  = \new_[9308]_  | \new_[9305]_ ;
  assign \new_[9312]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[9315]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[9316]_  = \new_[9315]_  | \new_[9312]_ ;
  assign \new_[9317]_  = \new_[9316]_  | \new_[9309]_ ;
  assign \new_[9318]_  = \new_[9317]_  | \new_[9302]_ ;
  assign \new_[9322]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[9323]_  = \new_[1095]_  | \new_[9322]_ ;
  assign \new_[9326]_  = \new_[1091]_  | \new_[1092]_ ;
  assign \new_[9329]_  = \new_[1089]_  | \new_[1090]_ ;
  assign \new_[9330]_  = \new_[9329]_  | \new_[9326]_ ;
  assign \new_[9331]_  = \new_[9330]_  | \new_[9323]_ ;
  assign \new_[9334]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[9337]_  = \new_[1085]_  | \new_[1086]_ ;
  assign \new_[9338]_  = \new_[9337]_  | \new_[9334]_ ;
  assign \new_[9341]_  = \new_[1083]_  | \new_[1084]_ ;
  assign \new_[9344]_  = \new_[1081]_  | \new_[1082]_ ;
  assign \new_[9345]_  = \new_[9344]_  | \new_[9341]_ ;
  assign \new_[9346]_  = \new_[9345]_  | \new_[9338]_ ;
  assign \new_[9347]_  = \new_[9346]_  | \new_[9331]_ ;
  assign \new_[9348]_  = \new_[9347]_  | \new_[9318]_ ;
  assign \new_[9349]_  = \new_[9348]_  | \new_[9289]_ ;
  assign \new_[9350]_  = \new_[9349]_  | \new_[9230]_ ;
  assign \new_[9354]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[9355]_  = \new_[1080]_  | \new_[9354]_ ;
  assign \new_[9358]_  = \new_[1076]_  | \new_[1077]_ ;
  assign \new_[9361]_  = \new_[1074]_  | \new_[1075]_ ;
  assign \new_[9362]_  = \new_[9361]_  | \new_[9358]_ ;
  assign \new_[9363]_  = \new_[9362]_  | \new_[9355]_ ;
  assign \new_[9366]_  = \new_[1072]_  | \new_[1073]_ ;
  assign \new_[9369]_  = \new_[1070]_  | \new_[1071]_ ;
  assign \new_[9370]_  = \new_[9369]_  | \new_[9366]_ ;
  assign \new_[9373]_  = \new_[1068]_  | \new_[1069]_ ;
  assign \new_[9376]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[9377]_  = \new_[9376]_  | \new_[9373]_ ;
  assign \new_[9378]_  = \new_[9377]_  | \new_[9370]_ ;
  assign \new_[9379]_  = \new_[9378]_  | \new_[9363]_ ;
  assign \new_[9383]_  = \new_[1063]_  | \new_[1064]_ ;
  assign \new_[9384]_  = \new_[1065]_  | \new_[9383]_ ;
  assign \new_[9387]_  = \new_[1061]_  | \new_[1062]_ ;
  assign \new_[9390]_  = \new_[1059]_  | \new_[1060]_ ;
  assign \new_[9391]_  = \new_[9390]_  | \new_[9387]_ ;
  assign \new_[9392]_  = \new_[9391]_  | \new_[9384]_ ;
  assign \new_[9395]_  = \new_[1057]_  | \new_[1058]_ ;
  assign \new_[9398]_  = \new_[1055]_  | \new_[1056]_ ;
  assign \new_[9399]_  = \new_[9398]_  | \new_[9395]_ ;
  assign \new_[9402]_  = \new_[1053]_  | \new_[1054]_ ;
  assign \new_[9405]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[9406]_  = \new_[9405]_  | \new_[9402]_ ;
  assign \new_[9407]_  = \new_[9406]_  | \new_[9399]_ ;
  assign \new_[9408]_  = \new_[9407]_  | \new_[9392]_ ;
  assign \new_[9409]_  = \new_[9408]_  | \new_[9379]_ ;
  assign \new_[9413]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[9414]_  = \new_[1050]_  | \new_[9413]_ ;
  assign \new_[9417]_  = \new_[1046]_  | \new_[1047]_ ;
  assign \new_[9420]_  = \new_[1044]_  | \new_[1045]_ ;
  assign \new_[9421]_  = \new_[9420]_  | \new_[9417]_ ;
  assign \new_[9422]_  = \new_[9421]_  | \new_[9414]_ ;
  assign \new_[9425]_  = \new_[1042]_  | \new_[1043]_ ;
  assign \new_[9428]_  = \new_[1040]_  | \new_[1041]_ ;
  assign \new_[9429]_  = \new_[9428]_  | \new_[9425]_ ;
  assign \new_[9432]_  = \new_[1038]_  | \new_[1039]_ ;
  assign \new_[9435]_  = \new_[1036]_  | \new_[1037]_ ;
  assign \new_[9436]_  = \new_[9435]_  | \new_[9432]_ ;
  assign \new_[9437]_  = \new_[9436]_  | \new_[9429]_ ;
  assign \new_[9438]_  = \new_[9437]_  | \new_[9422]_ ;
  assign \new_[9442]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[9443]_  = \new_[1035]_  | \new_[9442]_ ;
  assign \new_[9446]_  = \new_[1031]_  | \new_[1032]_ ;
  assign \new_[9449]_  = \new_[1029]_  | \new_[1030]_ ;
  assign \new_[9450]_  = \new_[9449]_  | \new_[9446]_ ;
  assign \new_[9451]_  = \new_[9450]_  | \new_[9443]_ ;
  assign \new_[9454]_  = \new_[1027]_  | \new_[1028]_ ;
  assign \new_[9457]_  = \new_[1025]_  | \new_[1026]_ ;
  assign \new_[9458]_  = \new_[9457]_  | \new_[9454]_ ;
  assign \new_[9461]_  = \new_[1023]_  | \new_[1024]_ ;
  assign \new_[9464]_  = \new_[1021]_  | \new_[1022]_ ;
  assign \new_[9465]_  = \new_[9464]_  | \new_[9461]_ ;
  assign \new_[9466]_  = \new_[9465]_  | \new_[9458]_ ;
  assign \new_[9467]_  = \new_[9466]_  | \new_[9451]_ ;
  assign \new_[9468]_  = \new_[9467]_  | \new_[9438]_ ;
  assign \new_[9469]_  = \new_[9468]_  | \new_[9409]_ ;
  assign \new_[9473]_  = \new_[1018]_  | \new_[1019]_ ;
  assign \new_[9474]_  = \new_[1020]_  | \new_[9473]_ ;
  assign \new_[9477]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[9480]_  = \new_[1014]_  | \new_[1015]_ ;
  assign \new_[9481]_  = \new_[9480]_  | \new_[9477]_ ;
  assign \new_[9482]_  = \new_[9481]_  | \new_[9474]_ ;
  assign \new_[9485]_  = \new_[1012]_  | \new_[1013]_ ;
  assign \new_[9488]_  = \new_[1010]_  | \new_[1011]_ ;
  assign \new_[9489]_  = \new_[9488]_  | \new_[9485]_ ;
  assign \new_[9492]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[9495]_  = \new_[1006]_  | \new_[1007]_ ;
  assign \new_[9496]_  = \new_[9495]_  | \new_[9492]_ ;
  assign \new_[9497]_  = \new_[9496]_  | \new_[9489]_ ;
  assign \new_[9498]_  = \new_[9497]_  | \new_[9482]_ ;
  assign \new_[9502]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[9503]_  = \new_[1005]_  | \new_[9502]_ ;
  assign \new_[9506]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[9509]_  = \new_[999]_  | \new_[1000]_ ;
  assign \new_[9510]_  = \new_[9509]_  | \new_[9506]_ ;
  assign \new_[9511]_  = \new_[9510]_  | \new_[9503]_ ;
  assign \new_[9514]_  = \new_[997]_  | \new_[998]_ ;
  assign \new_[9517]_  = \new_[995]_  | \new_[996]_ ;
  assign \new_[9518]_  = \new_[9517]_  | \new_[9514]_ ;
  assign \new_[9521]_  = \new_[993]_  | \new_[994]_ ;
  assign \new_[9524]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[9525]_  = \new_[9524]_  | \new_[9521]_ ;
  assign \new_[9526]_  = \new_[9525]_  | \new_[9518]_ ;
  assign \new_[9527]_  = \new_[9526]_  | \new_[9511]_ ;
  assign \new_[9528]_  = \new_[9527]_  | \new_[9498]_ ;
  assign \new_[9532]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[9533]_  = \new_[990]_  | \new_[9532]_ ;
  assign \new_[9536]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[9539]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[9540]_  = \new_[9539]_  | \new_[9536]_ ;
  assign \new_[9541]_  = \new_[9540]_  | \new_[9533]_ ;
  assign \new_[9544]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[9547]_  = \new_[980]_  | \new_[981]_ ;
  assign \new_[9548]_  = \new_[9547]_  | \new_[9544]_ ;
  assign \new_[9551]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[9554]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[9555]_  = \new_[9554]_  | \new_[9551]_ ;
  assign \new_[9556]_  = \new_[9555]_  | \new_[9548]_ ;
  assign \new_[9557]_  = \new_[9556]_  | \new_[9541]_ ;
  assign \new_[9561]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[9562]_  = \new_[975]_  | \new_[9561]_ ;
  assign \new_[9565]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[9568]_  = \new_[969]_  | \new_[970]_ ;
  assign \new_[9569]_  = \new_[9568]_  | \new_[9565]_ ;
  assign \new_[9570]_  = \new_[9569]_  | \new_[9562]_ ;
  assign \new_[9573]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[9576]_  = \new_[965]_  | \new_[966]_ ;
  assign \new_[9577]_  = \new_[9576]_  | \new_[9573]_ ;
  assign \new_[9580]_  = \new_[963]_  | \new_[964]_ ;
  assign \new_[9583]_  = \new_[961]_  | \new_[962]_ ;
  assign \new_[9584]_  = \new_[9583]_  | \new_[9580]_ ;
  assign \new_[9585]_  = \new_[9584]_  | \new_[9577]_ ;
  assign \new_[9586]_  = \new_[9585]_  | \new_[9570]_ ;
  assign \new_[9587]_  = \new_[9586]_  | \new_[9557]_ ;
  assign \new_[9588]_  = \new_[9587]_  | \new_[9528]_ ;
  assign \new_[9589]_  = \new_[9588]_  | \new_[9469]_ ;
  assign \new_[9590]_  = \new_[9589]_  | \new_[9350]_ ;
  assign \new_[9591]_  = \new_[9590]_  | \new_[9111]_ ;
  assign \new_[9592]_  = \new_[9591]_  | \new_[8632]_ ;
  assign \new_[9596]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[9597]_  = \new_[960]_  | \new_[9596]_ ;
  assign \new_[9600]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[9603]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[9604]_  = \new_[9603]_  | \new_[9600]_ ;
  assign \new_[9605]_  = \new_[9604]_  | \new_[9597]_ ;
  assign \new_[9608]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[9611]_  = \new_[950]_  | \new_[951]_ ;
  assign \new_[9612]_  = \new_[9611]_  | \new_[9608]_ ;
  assign \new_[9615]_  = \new_[948]_  | \new_[949]_ ;
  assign \new_[9618]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[9619]_  = \new_[9618]_  | \new_[9615]_ ;
  assign \new_[9620]_  = \new_[9619]_  | \new_[9612]_ ;
  assign \new_[9621]_  = \new_[9620]_  | \new_[9605]_ ;
  assign \new_[9625]_  = \new_[943]_  | \new_[944]_ ;
  assign \new_[9626]_  = \new_[945]_  | \new_[9625]_ ;
  assign \new_[9629]_  = \new_[941]_  | \new_[942]_ ;
  assign \new_[9632]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[9633]_  = \new_[9632]_  | \new_[9629]_ ;
  assign \new_[9634]_  = \new_[9633]_  | \new_[9626]_ ;
  assign \new_[9637]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[9640]_  = \new_[935]_  | \new_[936]_ ;
  assign \new_[9641]_  = \new_[9640]_  | \new_[9637]_ ;
  assign \new_[9644]_  = \new_[933]_  | \new_[934]_ ;
  assign \new_[9647]_  = \new_[931]_  | \new_[932]_ ;
  assign \new_[9648]_  = \new_[9647]_  | \new_[9644]_ ;
  assign \new_[9649]_  = \new_[9648]_  | \new_[9641]_ ;
  assign \new_[9650]_  = \new_[9649]_  | \new_[9634]_ ;
  assign \new_[9651]_  = \new_[9650]_  | \new_[9621]_ ;
  assign \new_[9655]_  = \new_[928]_  | \new_[929]_ ;
  assign \new_[9656]_  = \new_[930]_  | \new_[9655]_ ;
  assign \new_[9659]_  = \new_[926]_  | \new_[927]_ ;
  assign \new_[9662]_  = \new_[924]_  | \new_[925]_ ;
  assign \new_[9663]_  = \new_[9662]_  | \new_[9659]_ ;
  assign \new_[9664]_  = \new_[9663]_  | \new_[9656]_ ;
  assign \new_[9667]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[9670]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[9671]_  = \new_[9670]_  | \new_[9667]_ ;
  assign \new_[9674]_  = \new_[918]_  | \new_[919]_ ;
  assign \new_[9677]_  = \new_[916]_  | \new_[917]_ ;
  assign \new_[9678]_  = \new_[9677]_  | \new_[9674]_ ;
  assign \new_[9679]_  = \new_[9678]_  | \new_[9671]_ ;
  assign \new_[9680]_  = \new_[9679]_  | \new_[9664]_ ;
  assign \new_[9684]_  = \new_[913]_  | \new_[914]_ ;
  assign \new_[9685]_  = \new_[915]_  | \new_[9684]_ ;
  assign \new_[9688]_  = \new_[911]_  | \new_[912]_ ;
  assign \new_[9691]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[9692]_  = \new_[9691]_  | \new_[9688]_ ;
  assign \new_[9693]_  = \new_[9692]_  | \new_[9685]_ ;
  assign \new_[9696]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[9699]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[9700]_  = \new_[9699]_  | \new_[9696]_ ;
  assign \new_[9703]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[9706]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[9707]_  = \new_[9706]_  | \new_[9703]_ ;
  assign \new_[9708]_  = \new_[9707]_  | \new_[9700]_ ;
  assign \new_[9709]_  = \new_[9708]_  | \new_[9693]_ ;
  assign \new_[9710]_  = \new_[9709]_  | \new_[9680]_ ;
  assign \new_[9711]_  = \new_[9710]_  | \new_[9651]_ ;
  assign \new_[9715]_  = \new_[898]_  | \new_[899]_ ;
  assign \new_[9716]_  = \new_[900]_  | \new_[9715]_ ;
  assign \new_[9719]_  = \new_[896]_  | \new_[897]_ ;
  assign \new_[9722]_  = \new_[894]_  | \new_[895]_ ;
  assign \new_[9723]_  = \new_[9722]_  | \new_[9719]_ ;
  assign \new_[9724]_  = \new_[9723]_  | \new_[9716]_ ;
  assign \new_[9727]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[9730]_  = \new_[890]_  | \new_[891]_ ;
  assign \new_[9731]_  = \new_[9730]_  | \new_[9727]_ ;
  assign \new_[9734]_  = \new_[888]_  | \new_[889]_ ;
  assign \new_[9737]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[9738]_  = \new_[9737]_  | \new_[9734]_ ;
  assign \new_[9739]_  = \new_[9738]_  | \new_[9731]_ ;
  assign \new_[9740]_  = \new_[9739]_  | \new_[9724]_ ;
  assign \new_[9744]_  = \new_[883]_  | \new_[884]_ ;
  assign \new_[9745]_  = \new_[885]_  | \new_[9744]_ ;
  assign \new_[9748]_  = \new_[881]_  | \new_[882]_ ;
  assign \new_[9751]_  = \new_[879]_  | \new_[880]_ ;
  assign \new_[9752]_  = \new_[9751]_  | \new_[9748]_ ;
  assign \new_[9753]_  = \new_[9752]_  | \new_[9745]_ ;
  assign \new_[9756]_  = \new_[877]_  | \new_[878]_ ;
  assign \new_[9759]_  = \new_[875]_  | \new_[876]_ ;
  assign \new_[9760]_  = \new_[9759]_  | \new_[9756]_ ;
  assign \new_[9763]_  = \new_[873]_  | \new_[874]_ ;
  assign \new_[9766]_  = \new_[871]_  | \new_[872]_ ;
  assign \new_[9767]_  = \new_[9766]_  | \new_[9763]_ ;
  assign \new_[9768]_  = \new_[9767]_  | \new_[9760]_ ;
  assign \new_[9769]_  = \new_[9768]_  | \new_[9753]_ ;
  assign \new_[9770]_  = \new_[9769]_  | \new_[9740]_ ;
  assign \new_[9774]_  = \new_[868]_  | \new_[869]_ ;
  assign \new_[9775]_  = \new_[870]_  | \new_[9774]_ ;
  assign \new_[9778]_  = \new_[866]_  | \new_[867]_ ;
  assign \new_[9781]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[9782]_  = \new_[9781]_  | \new_[9778]_ ;
  assign \new_[9783]_  = \new_[9782]_  | \new_[9775]_ ;
  assign \new_[9786]_  = \new_[862]_  | \new_[863]_ ;
  assign \new_[9789]_  = \new_[860]_  | \new_[861]_ ;
  assign \new_[9790]_  = \new_[9789]_  | \new_[9786]_ ;
  assign \new_[9793]_  = \new_[858]_  | \new_[859]_ ;
  assign \new_[9796]_  = \new_[856]_  | \new_[857]_ ;
  assign \new_[9797]_  = \new_[9796]_  | \new_[9793]_ ;
  assign \new_[9798]_  = \new_[9797]_  | \new_[9790]_ ;
  assign \new_[9799]_  = \new_[9798]_  | \new_[9783]_ ;
  assign \new_[9803]_  = \new_[853]_  | \new_[854]_ ;
  assign \new_[9804]_  = \new_[855]_  | \new_[9803]_ ;
  assign \new_[9807]_  = \new_[851]_  | \new_[852]_ ;
  assign \new_[9810]_  = \new_[849]_  | \new_[850]_ ;
  assign \new_[9811]_  = \new_[9810]_  | \new_[9807]_ ;
  assign \new_[9812]_  = \new_[9811]_  | \new_[9804]_ ;
  assign \new_[9815]_  = \new_[847]_  | \new_[848]_ ;
  assign \new_[9818]_  = \new_[845]_  | \new_[846]_ ;
  assign \new_[9819]_  = \new_[9818]_  | \new_[9815]_ ;
  assign \new_[9822]_  = \new_[843]_  | \new_[844]_ ;
  assign \new_[9825]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[9826]_  = \new_[9825]_  | \new_[9822]_ ;
  assign \new_[9827]_  = \new_[9826]_  | \new_[9819]_ ;
  assign \new_[9828]_  = \new_[9827]_  | \new_[9812]_ ;
  assign \new_[9829]_  = \new_[9828]_  | \new_[9799]_ ;
  assign \new_[9830]_  = \new_[9829]_  | \new_[9770]_ ;
  assign \new_[9831]_  = \new_[9830]_  | \new_[9711]_ ;
  assign \new_[9835]_  = \new_[838]_  | \new_[839]_ ;
  assign \new_[9836]_  = \new_[840]_  | \new_[9835]_ ;
  assign \new_[9839]_  = \new_[836]_  | \new_[837]_ ;
  assign \new_[9842]_  = \new_[834]_  | \new_[835]_ ;
  assign \new_[9843]_  = \new_[9842]_  | \new_[9839]_ ;
  assign \new_[9844]_  = \new_[9843]_  | \new_[9836]_ ;
  assign \new_[9847]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[9850]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[9851]_  = \new_[9850]_  | \new_[9847]_ ;
  assign \new_[9854]_  = \new_[828]_  | \new_[829]_ ;
  assign \new_[9857]_  = \new_[826]_  | \new_[827]_ ;
  assign \new_[9858]_  = \new_[9857]_  | \new_[9854]_ ;
  assign \new_[9859]_  = \new_[9858]_  | \new_[9851]_ ;
  assign \new_[9860]_  = \new_[9859]_  | \new_[9844]_ ;
  assign \new_[9864]_  = \new_[823]_  | \new_[824]_ ;
  assign \new_[9865]_  = \new_[825]_  | \new_[9864]_ ;
  assign \new_[9868]_  = \new_[821]_  | \new_[822]_ ;
  assign \new_[9871]_  = \new_[819]_  | \new_[820]_ ;
  assign \new_[9872]_  = \new_[9871]_  | \new_[9868]_ ;
  assign \new_[9873]_  = \new_[9872]_  | \new_[9865]_ ;
  assign \new_[9876]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[9879]_  = \new_[815]_  | \new_[816]_ ;
  assign \new_[9880]_  = \new_[9879]_  | \new_[9876]_ ;
  assign \new_[9883]_  = \new_[813]_  | \new_[814]_ ;
  assign \new_[9886]_  = \new_[811]_  | \new_[812]_ ;
  assign \new_[9887]_  = \new_[9886]_  | \new_[9883]_ ;
  assign \new_[9888]_  = \new_[9887]_  | \new_[9880]_ ;
  assign \new_[9889]_  = \new_[9888]_  | \new_[9873]_ ;
  assign \new_[9890]_  = \new_[9889]_  | \new_[9860]_ ;
  assign \new_[9894]_  = \new_[808]_  | \new_[809]_ ;
  assign \new_[9895]_  = \new_[810]_  | \new_[9894]_ ;
  assign \new_[9898]_  = \new_[806]_  | \new_[807]_ ;
  assign \new_[9901]_  = \new_[804]_  | \new_[805]_ ;
  assign \new_[9902]_  = \new_[9901]_  | \new_[9898]_ ;
  assign \new_[9903]_  = \new_[9902]_  | \new_[9895]_ ;
  assign \new_[9906]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[9909]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[9910]_  = \new_[9909]_  | \new_[9906]_ ;
  assign \new_[9913]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[9916]_  = \new_[796]_  | \new_[797]_ ;
  assign \new_[9917]_  = \new_[9916]_  | \new_[9913]_ ;
  assign \new_[9918]_  = \new_[9917]_  | \new_[9910]_ ;
  assign \new_[9919]_  = \new_[9918]_  | \new_[9903]_ ;
  assign \new_[9923]_  = \new_[793]_  | \new_[794]_ ;
  assign \new_[9924]_  = \new_[795]_  | \new_[9923]_ ;
  assign \new_[9927]_  = \new_[791]_  | \new_[792]_ ;
  assign \new_[9930]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[9931]_  = \new_[9930]_  | \new_[9927]_ ;
  assign \new_[9932]_  = \new_[9931]_  | \new_[9924]_ ;
  assign \new_[9935]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[9938]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[9939]_  = \new_[9938]_  | \new_[9935]_ ;
  assign \new_[9942]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[9945]_  = \new_[781]_  | \new_[782]_ ;
  assign \new_[9946]_  = \new_[9945]_  | \new_[9942]_ ;
  assign \new_[9947]_  = \new_[9946]_  | \new_[9939]_ ;
  assign \new_[9948]_  = \new_[9947]_  | \new_[9932]_ ;
  assign \new_[9949]_  = \new_[9948]_  | \new_[9919]_ ;
  assign \new_[9950]_  = \new_[9949]_  | \new_[9890]_ ;
  assign \new_[9954]_  = \new_[778]_  | \new_[779]_ ;
  assign \new_[9955]_  = \new_[780]_  | \new_[9954]_ ;
  assign \new_[9958]_  = \new_[776]_  | \new_[777]_ ;
  assign \new_[9961]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[9962]_  = \new_[9961]_  | \new_[9958]_ ;
  assign \new_[9963]_  = \new_[9962]_  | \new_[9955]_ ;
  assign \new_[9966]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[9969]_  = \new_[770]_  | \new_[771]_ ;
  assign \new_[9970]_  = \new_[9969]_  | \new_[9966]_ ;
  assign \new_[9973]_  = \new_[768]_  | \new_[769]_ ;
  assign \new_[9976]_  = \new_[766]_  | \new_[767]_ ;
  assign \new_[9977]_  = \new_[9976]_  | \new_[9973]_ ;
  assign \new_[9978]_  = \new_[9977]_  | \new_[9970]_ ;
  assign \new_[9979]_  = \new_[9978]_  | \new_[9963]_ ;
  assign \new_[9983]_  = \new_[763]_  | \new_[764]_ ;
  assign \new_[9984]_  = \new_[765]_  | \new_[9983]_ ;
  assign \new_[9987]_  = \new_[761]_  | \new_[762]_ ;
  assign \new_[9990]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[9991]_  = \new_[9990]_  | \new_[9987]_ ;
  assign \new_[9992]_  = \new_[9991]_  | \new_[9984]_ ;
  assign \new_[9995]_  = \new_[757]_  | \new_[758]_ ;
  assign \new_[9998]_  = \new_[755]_  | \new_[756]_ ;
  assign \new_[9999]_  = \new_[9998]_  | \new_[9995]_ ;
  assign \new_[10002]_  = \new_[753]_  | \new_[754]_ ;
  assign \new_[10005]_  = \new_[751]_  | \new_[752]_ ;
  assign \new_[10006]_  = \new_[10005]_  | \new_[10002]_ ;
  assign \new_[10007]_  = \new_[10006]_  | \new_[9999]_ ;
  assign \new_[10008]_  = \new_[10007]_  | \new_[9992]_ ;
  assign \new_[10009]_  = \new_[10008]_  | \new_[9979]_ ;
  assign \new_[10013]_  = \new_[748]_  | \new_[749]_ ;
  assign \new_[10014]_  = \new_[750]_  | \new_[10013]_ ;
  assign \new_[10017]_  = \new_[746]_  | \new_[747]_ ;
  assign \new_[10020]_  = \new_[744]_  | \new_[745]_ ;
  assign \new_[10021]_  = \new_[10020]_  | \new_[10017]_ ;
  assign \new_[10022]_  = \new_[10021]_  | \new_[10014]_ ;
  assign \new_[10025]_  = \new_[742]_  | \new_[743]_ ;
  assign \new_[10028]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[10029]_  = \new_[10028]_  | \new_[10025]_ ;
  assign \new_[10032]_  = \new_[738]_  | \new_[739]_ ;
  assign \new_[10035]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[10036]_  = \new_[10035]_  | \new_[10032]_ ;
  assign \new_[10037]_  = \new_[10036]_  | \new_[10029]_ ;
  assign \new_[10038]_  = \new_[10037]_  | \new_[10022]_ ;
  assign \new_[10042]_  = \new_[733]_  | \new_[734]_ ;
  assign \new_[10043]_  = \new_[735]_  | \new_[10042]_ ;
  assign \new_[10046]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[10049]_  = \new_[729]_  | \new_[730]_ ;
  assign \new_[10050]_  = \new_[10049]_  | \new_[10046]_ ;
  assign \new_[10051]_  = \new_[10050]_  | \new_[10043]_ ;
  assign \new_[10054]_  = \new_[727]_  | \new_[728]_ ;
  assign \new_[10057]_  = \new_[725]_  | \new_[726]_ ;
  assign \new_[10058]_  = \new_[10057]_  | \new_[10054]_ ;
  assign \new_[10061]_  = \new_[723]_  | \new_[724]_ ;
  assign \new_[10064]_  = \new_[721]_  | \new_[722]_ ;
  assign \new_[10065]_  = \new_[10064]_  | \new_[10061]_ ;
  assign \new_[10066]_  = \new_[10065]_  | \new_[10058]_ ;
  assign \new_[10067]_  = \new_[10066]_  | \new_[10051]_ ;
  assign \new_[10068]_  = \new_[10067]_  | \new_[10038]_ ;
  assign \new_[10069]_  = \new_[10068]_  | \new_[10009]_ ;
  assign \new_[10070]_  = \new_[10069]_  | \new_[9950]_ ;
  assign \new_[10071]_  = \new_[10070]_  | \new_[9831]_ ;
  assign \new_[10075]_  = \new_[718]_  | \new_[719]_ ;
  assign \new_[10076]_  = \new_[720]_  | \new_[10075]_ ;
  assign \new_[10079]_  = \new_[716]_  | \new_[717]_ ;
  assign \new_[10082]_  = \new_[714]_  | \new_[715]_ ;
  assign \new_[10083]_  = \new_[10082]_  | \new_[10079]_ ;
  assign \new_[10084]_  = \new_[10083]_  | \new_[10076]_ ;
  assign \new_[10087]_  = \new_[712]_  | \new_[713]_ ;
  assign \new_[10090]_  = \new_[710]_  | \new_[711]_ ;
  assign \new_[10091]_  = \new_[10090]_  | \new_[10087]_ ;
  assign \new_[10094]_  = \new_[708]_  | \new_[709]_ ;
  assign \new_[10097]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[10098]_  = \new_[10097]_  | \new_[10094]_ ;
  assign \new_[10099]_  = \new_[10098]_  | \new_[10091]_ ;
  assign \new_[10100]_  = \new_[10099]_  | \new_[10084]_ ;
  assign \new_[10104]_  = \new_[703]_  | \new_[704]_ ;
  assign \new_[10105]_  = \new_[705]_  | \new_[10104]_ ;
  assign \new_[10108]_  = \new_[701]_  | \new_[702]_ ;
  assign \new_[10111]_  = \new_[699]_  | \new_[700]_ ;
  assign \new_[10112]_  = \new_[10111]_  | \new_[10108]_ ;
  assign \new_[10113]_  = \new_[10112]_  | \new_[10105]_ ;
  assign \new_[10116]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[10119]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[10120]_  = \new_[10119]_  | \new_[10116]_ ;
  assign \new_[10123]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[10126]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[10127]_  = \new_[10126]_  | \new_[10123]_ ;
  assign \new_[10128]_  = \new_[10127]_  | \new_[10120]_ ;
  assign \new_[10129]_  = \new_[10128]_  | \new_[10113]_ ;
  assign \new_[10130]_  = \new_[10129]_  | \new_[10100]_ ;
  assign \new_[10134]_  = \new_[688]_  | \new_[689]_ ;
  assign \new_[10135]_  = \new_[690]_  | \new_[10134]_ ;
  assign \new_[10138]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[10141]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[10142]_  = \new_[10141]_  | \new_[10138]_ ;
  assign \new_[10143]_  = \new_[10142]_  | \new_[10135]_ ;
  assign \new_[10146]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[10149]_  = \new_[680]_  | \new_[681]_ ;
  assign \new_[10150]_  = \new_[10149]_  | \new_[10146]_ ;
  assign \new_[10153]_  = \new_[678]_  | \new_[679]_ ;
  assign \new_[10156]_  = \new_[676]_  | \new_[677]_ ;
  assign \new_[10157]_  = \new_[10156]_  | \new_[10153]_ ;
  assign \new_[10158]_  = \new_[10157]_  | \new_[10150]_ ;
  assign \new_[10159]_  = \new_[10158]_  | \new_[10143]_ ;
  assign \new_[10163]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[10164]_  = \new_[675]_  | \new_[10163]_ ;
  assign \new_[10167]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[10170]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[10171]_  = \new_[10170]_  | \new_[10167]_ ;
  assign \new_[10172]_  = \new_[10171]_  | \new_[10164]_ ;
  assign \new_[10175]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[10178]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[10179]_  = \new_[10178]_  | \new_[10175]_ ;
  assign \new_[10182]_  = \new_[663]_  | \new_[664]_ ;
  assign \new_[10185]_  = \new_[661]_  | \new_[662]_ ;
  assign \new_[10186]_  = \new_[10185]_  | \new_[10182]_ ;
  assign \new_[10187]_  = \new_[10186]_  | \new_[10179]_ ;
  assign \new_[10188]_  = \new_[10187]_  | \new_[10172]_ ;
  assign \new_[10189]_  = \new_[10188]_  | \new_[10159]_ ;
  assign \new_[10190]_  = \new_[10189]_  | \new_[10130]_ ;
  assign \new_[10194]_  = \new_[658]_  | \new_[659]_ ;
  assign \new_[10195]_  = \new_[660]_  | \new_[10194]_ ;
  assign \new_[10198]_  = \new_[656]_  | \new_[657]_ ;
  assign \new_[10201]_  = \new_[654]_  | \new_[655]_ ;
  assign \new_[10202]_  = \new_[10201]_  | \new_[10198]_ ;
  assign \new_[10203]_  = \new_[10202]_  | \new_[10195]_ ;
  assign \new_[10206]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[10209]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[10210]_  = \new_[10209]_  | \new_[10206]_ ;
  assign \new_[10213]_  = \new_[648]_  | \new_[649]_ ;
  assign \new_[10216]_  = \new_[646]_  | \new_[647]_ ;
  assign \new_[10217]_  = \new_[10216]_  | \new_[10213]_ ;
  assign \new_[10218]_  = \new_[10217]_  | \new_[10210]_ ;
  assign \new_[10219]_  = \new_[10218]_  | \new_[10203]_ ;
  assign \new_[10223]_  = \new_[643]_  | \new_[644]_ ;
  assign \new_[10224]_  = \new_[645]_  | \new_[10223]_ ;
  assign \new_[10227]_  = \new_[641]_  | \new_[642]_ ;
  assign \new_[10230]_  = \new_[639]_  | \new_[640]_ ;
  assign \new_[10231]_  = \new_[10230]_  | \new_[10227]_ ;
  assign \new_[10232]_  = \new_[10231]_  | \new_[10224]_ ;
  assign \new_[10235]_  = \new_[637]_  | \new_[638]_ ;
  assign \new_[10238]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[10239]_  = \new_[10238]_  | \new_[10235]_ ;
  assign \new_[10242]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[10245]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[10246]_  = \new_[10245]_  | \new_[10242]_ ;
  assign \new_[10247]_  = \new_[10246]_  | \new_[10239]_ ;
  assign \new_[10248]_  = \new_[10247]_  | \new_[10232]_ ;
  assign \new_[10249]_  = \new_[10248]_  | \new_[10219]_ ;
  assign \new_[10253]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[10254]_  = \new_[630]_  | \new_[10253]_ ;
  assign \new_[10257]_  = \new_[626]_  | \new_[627]_ ;
  assign \new_[10260]_  = \new_[624]_  | \new_[625]_ ;
  assign \new_[10261]_  = \new_[10260]_  | \new_[10257]_ ;
  assign \new_[10262]_  = \new_[10261]_  | \new_[10254]_ ;
  assign \new_[10265]_  = \new_[622]_  | \new_[623]_ ;
  assign \new_[10268]_  = \new_[620]_  | \new_[621]_ ;
  assign \new_[10269]_  = \new_[10268]_  | \new_[10265]_ ;
  assign \new_[10272]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[10275]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[10276]_  = \new_[10275]_  | \new_[10272]_ ;
  assign \new_[10277]_  = \new_[10276]_  | \new_[10269]_ ;
  assign \new_[10278]_  = \new_[10277]_  | \new_[10262]_ ;
  assign \new_[10282]_  = \new_[613]_  | \new_[614]_ ;
  assign \new_[10283]_  = \new_[615]_  | \new_[10282]_ ;
  assign \new_[10286]_  = \new_[611]_  | \new_[612]_ ;
  assign \new_[10289]_  = \new_[609]_  | \new_[610]_ ;
  assign \new_[10290]_  = \new_[10289]_  | \new_[10286]_ ;
  assign \new_[10291]_  = \new_[10290]_  | \new_[10283]_ ;
  assign \new_[10294]_  = \new_[607]_  | \new_[608]_ ;
  assign \new_[10297]_  = \new_[605]_  | \new_[606]_ ;
  assign \new_[10298]_  = \new_[10297]_  | \new_[10294]_ ;
  assign \new_[10301]_  = \new_[603]_  | \new_[604]_ ;
  assign \new_[10304]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[10305]_  = \new_[10304]_  | \new_[10301]_ ;
  assign \new_[10306]_  = \new_[10305]_  | \new_[10298]_ ;
  assign \new_[10307]_  = \new_[10306]_  | \new_[10291]_ ;
  assign \new_[10308]_  = \new_[10307]_  | \new_[10278]_ ;
  assign \new_[10309]_  = \new_[10308]_  | \new_[10249]_ ;
  assign \new_[10310]_  = \new_[10309]_  | \new_[10190]_ ;
  assign \new_[10314]_  = \new_[598]_  | \new_[599]_ ;
  assign \new_[10315]_  = \new_[600]_  | \new_[10314]_ ;
  assign \new_[10318]_  = \new_[596]_  | \new_[597]_ ;
  assign \new_[10321]_  = \new_[594]_  | \new_[595]_ ;
  assign \new_[10322]_  = \new_[10321]_  | \new_[10318]_ ;
  assign \new_[10323]_  = \new_[10322]_  | \new_[10315]_ ;
  assign \new_[10326]_  = \new_[592]_  | \new_[593]_ ;
  assign \new_[10329]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[10330]_  = \new_[10329]_  | \new_[10326]_ ;
  assign \new_[10333]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[10336]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[10337]_  = \new_[10336]_  | \new_[10333]_ ;
  assign \new_[10338]_  = \new_[10337]_  | \new_[10330]_ ;
  assign \new_[10339]_  = \new_[10338]_  | \new_[10323]_ ;
  assign \new_[10343]_  = \new_[583]_  | \new_[584]_ ;
  assign \new_[10344]_  = \new_[585]_  | \new_[10343]_ ;
  assign \new_[10347]_  = \new_[581]_  | \new_[582]_ ;
  assign \new_[10350]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[10351]_  = \new_[10350]_  | \new_[10347]_ ;
  assign \new_[10352]_  = \new_[10351]_  | \new_[10344]_ ;
  assign \new_[10355]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[10358]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[10359]_  = \new_[10358]_  | \new_[10355]_ ;
  assign \new_[10362]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[10365]_  = \new_[571]_  | \new_[572]_ ;
  assign \new_[10366]_  = \new_[10365]_  | \new_[10362]_ ;
  assign \new_[10367]_  = \new_[10366]_  | \new_[10359]_ ;
  assign \new_[10368]_  = \new_[10367]_  | \new_[10352]_ ;
  assign \new_[10369]_  = \new_[10368]_  | \new_[10339]_ ;
  assign \new_[10373]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[10374]_  = \new_[570]_  | \new_[10373]_ ;
  assign \new_[10377]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[10380]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[10381]_  = \new_[10380]_  | \new_[10377]_ ;
  assign \new_[10382]_  = \new_[10381]_  | \new_[10374]_ ;
  assign \new_[10385]_  = \new_[562]_  | \new_[563]_ ;
  assign \new_[10388]_  = \new_[560]_  | \new_[561]_ ;
  assign \new_[10389]_  = \new_[10388]_  | \new_[10385]_ ;
  assign \new_[10392]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[10395]_  = \new_[556]_  | \new_[557]_ ;
  assign \new_[10396]_  = \new_[10395]_  | \new_[10392]_ ;
  assign \new_[10397]_  = \new_[10396]_  | \new_[10389]_ ;
  assign \new_[10398]_  = \new_[10397]_  | \new_[10382]_ ;
  assign \new_[10402]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[10403]_  = \new_[555]_  | \new_[10402]_ ;
  assign \new_[10406]_  = \new_[551]_  | \new_[552]_ ;
  assign \new_[10409]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[10410]_  = \new_[10409]_  | \new_[10406]_ ;
  assign \new_[10411]_  = \new_[10410]_  | \new_[10403]_ ;
  assign \new_[10414]_  = \new_[547]_  | \new_[548]_ ;
  assign \new_[10417]_  = \new_[545]_  | \new_[546]_ ;
  assign \new_[10418]_  = \new_[10417]_  | \new_[10414]_ ;
  assign \new_[10421]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[10424]_  = \new_[541]_  | \new_[542]_ ;
  assign \new_[10425]_  = \new_[10424]_  | \new_[10421]_ ;
  assign \new_[10426]_  = \new_[10425]_  | \new_[10418]_ ;
  assign \new_[10427]_  = \new_[10426]_  | \new_[10411]_ ;
  assign \new_[10428]_  = \new_[10427]_  | \new_[10398]_ ;
  assign \new_[10429]_  = \new_[10428]_  | \new_[10369]_ ;
  assign \new_[10433]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[10434]_  = \new_[540]_  | \new_[10433]_ ;
  assign \new_[10437]_  = \new_[536]_  | \new_[537]_ ;
  assign \new_[10440]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[10441]_  = \new_[10440]_  | \new_[10437]_ ;
  assign \new_[10442]_  = \new_[10441]_  | \new_[10434]_ ;
  assign \new_[10445]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[10448]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[10449]_  = \new_[10448]_  | \new_[10445]_ ;
  assign \new_[10452]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[10455]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[10456]_  = \new_[10455]_  | \new_[10452]_ ;
  assign \new_[10457]_  = \new_[10456]_  | \new_[10449]_ ;
  assign \new_[10458]_  = \new_[10457]_  | \new_[10442]_ ;
  assign \new_[10462]_  = \new_[523]_  | \new_[524]_ ;
  assign \new_[10463]_  = \new_[525]_  | \new_[10462]_ ;
  assign \new_[10466]_  = \new_[521]_  | \new_[522]_ ;
  assign \new_[10469]_  = \new_[519]_  | \new_[520]_ ;
  assign \new_[10470]_  = \new_[10469]_  | \new_[10466]_ ;
  assign \new_[10471]_  = \new_[10470]_  | \new_[10463]_ ;
  assign \new_[10474]_  = \new_[517]_  | \new_[518]_ ;
  assign \new_[10477]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[10478]_  = \new_[10477]_  | \new_[10474]_ ;
  assign \new_[10481]_  = \new_[513]_  | \new_[514]_ ;
  assign \new_[10484]_  = \new_[511]_  | \new_[512]_ ;
  assign \new_[10485]_  = \new_[10484]_  | \new_[10481]_ ;
  assign \new_[10486]_  = \new_[10485]_  | \new_[10478]_ ;
  assign \new_[10487]_  = \new_[10486]_  | \new_[10471]_ ;
  assign \new_[10488]_  = \new_[10487]_  | \new_[10458]_ ;
  assign \new_[10492]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[10493]_  = \new_[510]_  | \new_[10492]_ ;
  assign \new_[10496]_  = \new_[506]_  | \new_[507]_ ;
  assign \new_[10499]_  = \new_[504]_  | \new_[505]_ ;
  assign \new_[10500]_  = \new_[10499]_  | \new_[10496]_ ;
  assign \new_[10501]_  = \new_[10500]_  | \new_[10493]_ ;
  assign \new_[10504]_  = \new_[502]_  | \new_[503]_ ;
  assign \new_[10507]_  = \new_[500]_  | \new_[501]_ ;
  assign \new_[10508]_  = \new_[10507]_  | \new_[10504]_ ;
  assign \new_[10511]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[10514]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[10515]_  = \new_[10514]_  | \new_[10511]_ ;
  assign \new_[10516]_  = \new_[10515]_  | \new_[10508]_ ;
  assign \new_[10517]_  = \new_[10516]_  | \new_[10501]_ ;
  assign \new_[10521]_  = \new_[493]_  | \new_[494]_ ;
  assign \new_[10522]_  = \new_[495]_  | \new_[10521]_ ;
  assign \new_[10525]_  = \new_[491]_  | \new_[492]_ ;
  assign \new_[10528]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[10529]_  = \new_[10528]_  | \new_[10525]_ ;
  assign \new_[10530]_  = \new_[10529]_  | \new_[10522]_ ;
  assign \new_[10533]_  = \new_[487]_  | \new_[488]_ ;
  assign \new_[10536]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[10537]_  = \new_[10536]_  | \new_[10533]_ ;
  assign \new_[10540]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[10543]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[10544]_  = \new_[10543]_  | \new_[10540]_ ;
  assign \new_[10545]_  = \new_[10544]_  | \new_[10537]_ ;
  assign \new_[10546]_  = \new_[10545]_  | \new_[10530]_ ;
  assign \new_[10547]_  = \new_[10546]_  | \new_[10517]_ ;
  assign \new_[10548]_  = \new_[10547]_  | \new_[10488]_ ;
  assign \new_[10549]_  = \new_[10548]_  | \new_[10429]_ ;
  assign \new_[10550]_  = \new_[10549]_  | \new_[10310]_ ;
  assign \new_[10551]_  = \new_[10550]_  | \new_[10071]_ ;
  assign \new_[10555]_  = \new_[478]_  | \new_[479]_ ;
  assign \new_[10556]_  = \new_[480]_  | \new_[10555]_ ;
  assign \new_[10559]_  = \new_[476]_  | \new_[477]_ ;
  assign \new_[10562]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[10563]_  = \new_[10562]_  | \new_[10559]_ ;
  assign \new_[10564]_  = \new_[10563]_  | \new_[10556]_ ;
  assign \new_[10567]_  = \new_[472]_  | \new_[473]_ ;
  assign \new_[10570]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[10571]_  = \new_[10570]_  | \new_[10567]_ ;
  assign \new_[10574]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[10577]_  = \new_[466]_  | \new_[467]_ ;
  assign \new_[10578]_  = \new_[10577]_  | \new_[10574]_ ;
  assign \new_[10579]_  = \new_[10578]_  | \new_[10571]_ ;
  assign \new_[10580]_  = \new_[10579]_  | \new_[10564]_ ;
  assign \new_[10584]_  = \new_[463]_  | \new_[464]_ ;
  assign \new_[10585]_  = \new_[465]_  | \new_[10584]_ ;
  assign \new_[10588]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[10591]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[10592]_  = \new_[10591]_  | \new_[10588]_ ;
  assign \new_[10593]_  = \new_[10592]_  | \new_[10585]_ ;
  assign \new_[10596]_  = \new_[457]_  | \new_[458]_ ;
  assign \new_[10599]_  = \new_[455]_  | \new_[456]_ ;
  assign \new_[10600]_  = \new_[10599]_  | \new_[10596]_ ;
  assign \new_[10603]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[10606]_  = \new_[451]_  | \new_[452]_ ;
  assign \new_[10607]_  = \new_[10606]_  | \new_[10603]_ ;
  assign \new_[10608]_  = \new_[10607]_  | \new_[10600]_ ;
  assign \new_[10609]_  = \new_[10608]_  | \new_[10593]_ ;
  assign \new_[10610]_  = \new_[10609]_  | \new_[10580]_ ;
  assign \new_[10614]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[10615]_  = \new_[450]_  | \new_[10614]_ ;
  assign \new_[10618]_  = \new_[446]_  | \new_[447]_ ;
  assign \new_[10621]_  = \new_[444]_  | \new_[445]_ ;
  assign \new_[10622]_  = \new_[10621]_  | \new_[10618]_ ;
  assign \new_[10623]_  = \new_[10622]_  | \new_[10615]_ ;
  assign \new_[10626]_  = \new_[442]_  | \new_[443]_ ;
  assign \new_[10629]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[10630]_  = \new_[10629]_  | \new_[10626]_ ;
  assign \new_[10633]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[10636]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[10637]_  = \new_[10636]_  | \new_[10633]_ ;
  assign \new_[10638]_  = \new_[10637]_  | \new_[10630]_ ;
  assign \new_[10639]_  = \new_[10638]_  | \new_[10623]_ ;
  assign \new_[10643]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[10644]_  = \new_[435]_  | \new_[10643]_ ;
  assign \new_[10647]_  = \new_[431]_  | \new_[432]_ ;
  assign \new_[10650]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[10651]_  = \new_[10650]_  | \new_[10647]_ ;
  assign \new_[10652]_  = \new_[10651]_  | \new_[10644]_ ;
  assign \new_[10655]_  = \new_[427]_  | \new_[428]_ ;
  assign \new_[10658]_  = \new_[425]_  | \new_[426]_ ;
  assign \new_[10659]_  = \new_[10658]_  | \new_[10655]_ ;
  assign \new_[10662]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[10665]_  = \new_[421]_  | \new_[422]_ ;
  assign \new_[10666]_  = \new_[10665]_  | \new_[10662]_ ;
  assign \new_[10667]_  = \new_[10666]_  | \new_[10659]_ ;
  assign \new_[10668]_  = \new_[10667]_  | \new_[10652]_ ;
  assign \new_[10669]_  = \new_[10668]_  | \new_[10639]_ ;
  assign \new_[10670]_  = \new_[10669]_  | \new_[10610]_ ;
  assign \new_[10674]_  = \new_[418]_  | \new_[419]_ ;
  assign \new_[10675]_  = \new_[420]_  | \new_[10674]_ ;
  assign \new_[10678]_  = \new_[416]_  | \new_[417]_ ;
  assign \new_[10681]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[10682]_  = \new_[10681]_  | \new_[10678]_ ;
  assign \new_[10683]_  = \new_[10682]_  | \new_[10675]_ ;
  assign \new_[10686]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[10689]_  = \new_[410]_  | \new_[411]_ ;
  assign \new_[10690]_  = \new_[10689]_  | \new_[10686]_ ;
  assign \new_[10693]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[10696]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[10697]_  = \new_[10696]_  | \new_[10693]_ ;
  assign \new_[10698]_  = \new_[10697]_  | \new_[10690]_ ;
  assign \new_[10699]_  = \new_[10698]_  | \new_[10683]_ ;
  assign \new_[10703]_  = \new_[403]_  | \new_[404]_ ;
  assign \new_[10704]_  = \new_[405]_  | \new_[10703]_ ;
  assign \new_[10707]_  = \new_[401]_  | \new_[402]_ ;
  assign \new_[10710]_  = \new_[399]_  | \new_[400]_ ;
  assign \new_[10711]_  = \new_[10710]_  | \new_[10707]_ ;
  assign \new_[10712]_  = \new_[10711]_  | \new_[10704]_ ;
  assign \new_[10715]_  = \new_[397]_  | \new_[398]_ ;
  assign \new_[10718]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[10719]_  = \new_[10718]_  | \new_[10715]_ ;
  assign \new_[10722]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[10725]_  = \new_[391]_  | \new_[392]_ ;
  assign \new_[10726]_  = \new_[10725]_  | \new_[10722]_ ;
  assign \new_[10727]_  = \new_[10726]_  | \new_[10719]_ ;
  assign \new_[10728]_  = \new_[10727]_  | \new_[10712]_ ;
  assign \new_[10729]_  = \new_[10728]_  | \new_[10699]_ ;
  assign \new_[10733]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[10734]_  = \new_[390]_  | \new_[10733]_ ;
  assign \new_[10737]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[10740]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[10741]_  = \new_[10740]_  | \new_[10737]_ ;
  assign \new_[10742]_  = \new_[10741]_  | \new_[10734]_ ;
  assign \new_[10745]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[10748]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[10749]_  = \new_[10748]_  | \new_[10745]_ ;
  assign \new_[10752]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[10755]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[10756]_  = \new_[10755]_  | \new_[10752]_ ;
  assign \new_[10757]_  = \new_[10756]_  | \new_[10749]_ ;
  assign \new_[10758]_  = \new_[10757]_  | \new_[10742]_ ;
  assign \new_[10762]_  = \new_[373]_  | \new_[374]_ ;
  assign \new_[10763]_  = \new_[375]_  | \new_[10762]_ ;
  assign \new_[10766]_  = \new_[371]_  | \new_[372]_ ;
  assign \new_[10769]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[10770]_  = \new_[10769]_  | \new_[10766]_ ;
  assign \new_[10771]_  = \new_[10770]_  | \new_[10763]_ ;
  assign \new_[10774]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[10777]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[10778]_  = \new_[10777]_  | \new_[10774]_ ;
  assign \new_[10781]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[10784]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[10785]_  = \new_[10784]_  | \new_[10781]_ ;
  assign \new_[10786]_  = \new_[10785]_  | \new_[10778]_ ;
  assign \new_[10787]_  = \new_[10786]_  | \new_[10771]_ ;
  assign \new_[10788]_  = \new_[10787]_  | \new_[10758]_ ;
  assign \new_[10789]_  = \new_[10788]_  | \new_[10729]_ ;
  assign \new_[10790]_  = \new_[10789]_  | \new_[10670]_ ;
  assign \new_[10794]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[10795]_  = \new_[360]_  | \new_[10794]_ ;
  assign \new_[10798]_  = \new_[356]_  | \new_[357]_ ;
  assign \new_[10801]_  = \new_[354]_  | \new_[355]_ ;
  assign \new_[10802]_  = \new_[10801]_  | \new_[10798]_ ;
  assign \new_[10803]_  = \new_[10802]_  | \new_[10795]_ ;
  assign \new_[10806]_  = \new_[352]_  | \new_[353]_ ;
  assign \new_[10809]_  = \new_[350]_  | \new_[351]_ ;
  assign \new_[10810]_  = \new_[10809]_  | \new_[10806]_ ;
  assign \new_[10813]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[10816]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[10817]_  = \new_[10816]_  | \new_[10813]_ ;
  assign \new_[10818]_  = \new_[10817]_  | \new_[10810]_ ;
  assign \new_[10819]_  = \new_[10818]_  | \new_[10803]_ ;
  assign \new_[10823]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[10824]_  = \new_[345]_  | \new_[10823]_ ;
  assign \new_[10827]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[10830]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[10831]_  = \new_[10830]_  | \new_[10827]_ ;
  assign \new_[10832]_  = \new_[10831]_  | \new_[10824]_ ;
  assign \new_[10835]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[10838]_  = \new_[335]_  | \new_[336]_ ;
  assign \new_[10839]_  = \new_[10838]_  | \new_[10835]_ ;
  assign \new_[10842]_  = \new_[333]_  | \new_[334]_ ;
  assign \new_[10845]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[10846]_  = \new_[10845]_  | \new_[10842]_ ;
  assign \new_[10847]_  = \new_[10846]_  | \new_[10839]_ ;
  assign \new_[10848]_  = \new_[10847]_  | \new_[10832]_ ;
  assign \new_[10849]_  = \new_[10848]_  | \new_[10819]_ ;
  assign \new_[10853]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[10854]_  = \new_[330]_  | \new_[10853]_ ;
  assign \new_[10857]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[10860]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[10861]_  = \new_[10860]_  | \new_[10857]_ ;
  assign \new_[10862]_  = \new_[10861]_  | \new_[10854]_ ;
  assign \new_[10865]_  = \new_[322]_  | \new_[323]_ ;
  assign \new_[10868]_  = \new_[320]_  | \new_[321]_ ;
  assign \new_[10869]_  = \new_[10868]_  | \new_[10865]_ ;
  assign \new_[10872]_  = \new_[318]_  | \new_[319]_ ;
  assign \new_[10875]_  = \new_[316]_  | \new_[317]_ ;
  assign \new_[10876]_  = \new_[10875]_  | \new_[10872]_ ;
  assign \new_[10877]_  = \new_[10876]_  | \new_[10869]_ ;
  assign \new_[10878]_  = \new_[10877]_  | \new_[10862]_ ;
  assign \new_[10882]_  = \new_[313]_  | \new_[314]_ ;
  assign \new_[10883]_  = \new_[315]_  | \new_[10882]_ ;
  assign \new_[10886]_  = \new_[311]_  | \new_[312]_ ;
  assign \new_[10889]_  = \new_[309]_  | \new_[310]_ ;
  assign \new_[10890]_  = \new_[10889]_  | \new_[10886]_ ;
  assign \new_[10891]_  = \new_[10890]_  | \new_[10883]_ ;
  assign \new_[10894]_  = \new_[307]_  | \new_[308]_ ;
  assign \new_[10897]_  = \new_[305]_  | \new_[306]_ ;
  assign \new_[10898]_  = \new_[10897]_  | \new_[10894]_ ;
  assign \new_[10901]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[10904]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[10905]_  = \new_[10904]_  | \new_[10901]_ ;
  assign \new_[10906]_  = \new_[10905]_  | \new_[10898]_ ;
  assign \new_[10907]_  = \new_[10906]_  | \new_[10891]_ ;
  assign \new_[10908]_  = \new_[10907]_  | \new_[10878]_ ;
  assign \new_[10909]_  = \new_[10908]_  | \new_[10849]_ ;
  assign \new_[10913]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[10914]_  = \new_[300]_  | \new_[10913]_ ;
  assign \new_[10917]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[10920]_  = \new_[294]_  | \new_[295]_ ;
  assign \new_[10921]_  = \new_[10920]_  | \new_[10917]_ ;
  assign \new_[10922]_  = \new_[10921]_  | \new_[10914]_ ;
  assign \new_[10925]_  = \new_[292]_  | \new_[293]_ ;
  assign \new_[10928]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[10929]_  = \new_[10928]_  | \new_[10925]_ ;
  assign \new_[10932]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[10935]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[10936]_  = \new_[10935]_  | \new_[10932]_ ;
  assign \new_[10937]_  = \new_[10936]_  | \new_[10929]_ ;
  assign \new_[10938]_  = \new_[10937]_  | \new_[10922]_ ;
  assign \new_[10942]_  = \new_[283]_  | \new_[284]_ ;
  assign \new_[10943]_  = \new_[285]_  | \new_[10942]_ ;
  assign \new_[10946]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[10949]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[10950]_  = \new_[10949]_  | \new_[10946]_ ;
  assign \new_[10951]_  = \new_[10950]_  | \new_[10943]_ ;
  assign \new_[10954]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[10957]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[10958]_  = \new_[10957]_  | \new_[10954]_ ;
  assign \new_[10961]_  = \new_[273]_  | \new_[274]_ ;
  assign \new_[10964]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[10965]_  = \new_[10964]_  | \new_[10961]_ ;
  assign \new_[10966]_  = \new_[10965]_  | \new_[10958]_ ;
  assign \new_[10967]_  = \new_[10966]_  | \new_[10951]_ ;
  assign \new_[10968]_  = \new_[10967]_  | \new_[10938]_ ;
  assign \new_[10972]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[10973]_  = \new_[270]_  | \new_[10972]_ ;
  assign \new_[10976]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[10979]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[10980]_  = \new_[10979]_  | \new_[10976]_ ;
  assign \new_[10981]_  = \new_[10980]_  | \new_[10973]_ ;
  assign \new_[10984]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[10987]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[10988]_  = \new_[10987]_  | \new_[10984]_ ;
  assign \new_[10991]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[10994]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[10995]_  = \new_[10994]_  | \new_[10991]_ ;
  assign \new_[10996]_  = \new_[10995]_  | \new_[10988]_ ;
  assign \new_[10997]_  = \new_[10996]_  | \new_[10981]_ ;
  assign \new_[11001]_  = \new_[253]_  | \new_[254]_ ;
  assign \new_[11002]_  = \new_[255]_  | \new_[11001]_ ;
  assign \new_[11005]_  = \new_[251]_  | \new_[252]_ ;
  assign \new_[11008]_  = \new_[249]_  | \new_[250]_ ;
  assign \new_[11009]_  = \new_[11008]_  | \new_[11005]_ ;
  assign \new_[11010]_  = \new_[11009]_  | \new_[11002]_ ;
  assign \new_[11013]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[11016]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[11017]_  = \new_[11016]_  | \new_[11013]_ ;
  assign \new_[11020]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[11023]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[11024]_  = \new_[11023]_  | \new_[11020]_ ;
  assign \new_[11025]_  = \new_[11024]_  | \new_[11017]_ ;
  assign \new_[11026]_  = \new_[11025]_  | \new_[11010]_ ;
  assign \new_[11027]_  = \new_[11026]_  | \new_[10997]_ ;
  assign \new_[11028]_  = \new_[11027]_  | \new_[10968]_ ;
  assign \new_[11029]_  = \new_[11028]_  | \new_[10909]_ ;
  assign \new_[11030]_  = \new_[11029]_  | \new_[10790]_ ;
  assign \new_[11034]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[11035]_  = \new_[240]_  | \new_[11034]_ ;
  assign \new_[11038]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[11041]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[11042]_  = \new_[11041]_  | \new_[11038]_ ;
  assign \new_[11043]_  = \new_[11042]_  | \new_[11035]_ ;
  assign \new_[11046]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[11049]_  = \new_[230]_  | \new_[231]_ ;
  assign \new_[11050]_  = \new_[11049]_  | \new_[11046]_ ;
  assign \new_[11053]_  = \new_[228]_  | \new_[229]_ ;
  assign \new_[11056]_  = \new_[226]_  | \new_[227]_ ;
  assign \new_[11057]_  = \new_[11056]_  | \new_[11053]_ ;
  assign \new_[11058]_  = \new_[11057]_  | \new_[11050]_ ;
  assign \new_[11059]_  = \new_[11058]_  | \new_[11043]_ ;
  assign \new_[11063]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[11064]_  = \new_[225]_  | \new_[11063]_ ;
  assign \new_[11067]_  = \new_[221]_  | \new_[222]_ ;
  assign \new_[11070]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[11071]_  = \new_[11070]_  | \new_[11067]_ ;
  assign \new_[11072]_  = \new_[11071]_  | \new_[11064]_ ;
  assign \new_[11075]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[11078]_  = \new_[215]_  | \new_[216]_ ;
  assign \new_[11079]_  = \new_[11078]_  | \new_[11075]_ ;
  assign \new_[11082]_  = \new_[213]_  | \new_[214]_ ;
  assign \new_[11085]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[11086]_  = \new_[11085]_  | \new_[11082]_ ;
  assign \new_[11087]_  = \new_[11086]_  | \new_[11079]_ ;
  assign \new_[11088]_  = \new_[11087]_  | \new_[11072]_ ;
  assign \new_[11089]_  = \new_[11088]_  | \new_[11059]_ ;
  assign \new_[11093]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[11094]_  = \new_[210]_  | \new_[11093]_ ;
  assign \new_[11097]_  = \new_[206]_  | \new_[207]_ ;
  assign \new_[11100]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[11101]_  = \new_[11100]_  | \new_[11097]_ ;
  assign \new_[11102]_  = \new_[11101]_  | \new_[11094]_ ;
  assign \new_[11105]_  = \new_[202]_  | \new_[203]_ ;
  assign \new_[11108]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[11109]_  = \new_[11108]_  | \new_[11105]_ ;
  assign \new_[11112]_  = \new_[198]_  | \new_[199]_ ;
  assign \new_[11115]_  = \new_[196]_  | \new_[197]_ ;
  assign \new_[11116]_  = \new_[11115]_  | \new_[11112]_ ;
  assign \new_[11117]_  = \new_[11116]_  | \new_[11109]_ ;
  assign \new_[11118]_  = \new_[11117]_  | \new_[11102]_ ;
  assign \new_[11122]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[11123]_  = \new_[195]_  | \new_[11122]_ ;
  assign \new_[11126]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[11129]_  = \new_[189]_  | \new_[190]_ ;
  assign \new_[11130]_  = \new_[11129]_  | \new_[11126]_ ;
  assign \new_[11131]_  = \new_[11130]_  | \new_[11123]_ ;
  assign \new_[11134]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[11137]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[11138]_  = \new_[11137]_  | \new_[11134]_ ;
  assign \new_[11141]_  = \new_[183]_  | \new_[184]_ ;
  assign \new_[11144]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[11145]_  = \new_[11144]_  | \new_[11141]_ ;
  assign \new_[11146]_  = \new_[11145]_  | \new_[11138]_ ;
  assign \new_[11147]_  = \new_[11146]_  | \new_[11131]_ ;
  assign \new_[11148]_  = \new_[11147]_  | \new_[11118]_ ;
  assign \new_[11149]_  = \new_[11148]_  | \new_[11089]_ ;
  assign \new_[11153]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[11154]_  = \new_[180]_  | \new_[11153]_ ;
  assign \new_[11157]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[11160]_  = \new_[174]_  | \new_[175]_ ;
  assign \new_[11161]_  = \new_[11160]_  | \new_[11157]_ ;
  assign \new_[11162]_  = \new_[11161]_  | \new_[11154]_ ;
  assign \new_[11165]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[11168]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[11169]_  = \new_[11168]_  | \new_[11165]_ ;
  assign \new_[11172]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[11175]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[11176]_  = \new_[11175]_  | \new_[11172]_ ;
  assign \new_[11177]_  = \new_[11176]_  | \new_[11169]_ ;
  assign \new_[11178]_  = \new_[11177]_  | \new_[11162]_ ;
  assign \new_[11182]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[11183]_  = \new_[165]_  | \new_[11182]_ ;
  assign \new_[11186]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[11189]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[11190]_  = \new_[11189]_  | \new_[11186]_ ;
  assign \new_[11191]_  = \new_[11190]_  | \new_[11183]_ ;
  assign \new_[11194]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[11197]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[11198]_  = \new_[11197]_  | \new_[11194]_ ;
  assign \new_[11201]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[11204]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[11205]_  = \new_[11204]_  | \new_[11201]_ ;
  assign \new_[11206]_  = \new_[11205]_  | \new_[11198]_ ;
  assign \new_[11207]_  = \new_[11206]_  | \new_[11191]_ ;
  assign \new_[11208]_  = \new_[11207]_  | \new_[11178]_ ;
  assign \new_[11212]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[11213]_  = \new_[150]_  | \new_[11212]_ ;
  assign \new_[11216]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[11219]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[11220]_  = \new_[11219]_  | \new_[11216]_ ;
  assign \new_[11221]_  = \new_[11220]_  | \new_[11213]_ ;
  assign \new_[11224]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[11227]_  = \new_[140]_  | \new_[141]_ ;
  assign \new_[11228]_  = \new_[11227]_  | \new_[11224]_ ;
  assign \new_[11231]_  = \new_[138]_  | \new_[139]_ ;
  assign \new_[11234]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[11235]_  = \new_[11234]_  | \new_[11231]_ ;
  assign \new_[11236]_  = \new_[11235]_  | \new_[11228]_ ;
  assign \new_[11237]_  = \new_[11236]_  | \new_[11221]_ ;
  assign \new_[11241]_  = \new_[133]_  | \new_[134]_ ;
  assign \new_[11242]_  = \new_[135]_  | \new_[11241]_ ;
  assign \new_[11245]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[11248]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[11249]_  = \new_[11248]_  | \new_[11245]_ ;
  assign \new_[11250]_  = \new_[11249]_  | \new_[11242]_ ;
  assign \new_[11253]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[11256]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[11257]_  = \new_[11256]_  | \new_[11253]_ ;
  assign \new_[11260]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[11263]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[11264]_  = \new_[11263]_  | \new_[11260]_ ;
  assign \new_[11265]_  = \new_[11264]_  | \new_[11257]_ ;
  assign \new_[11266]_  = \new_[11265]_  | \new_[11250]_ ;
  assign \new_[11267]_  = \new_[11266]_  | \new_[11237]_ ;
  assign \new_[11268]_  = \new_[11267]_  | \new_[11208]_ ;
  assign \new_[11269]_  = \new_[11268]_  | \new_[11149]_ ;
  assign \new_[11273]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[11274]_  = \new_[120]_  | \new_[11273]_ ;
  assign \new_[11277]_  = \new_[116]_  | \new_[117]_ ;
  assign \new_[11280]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[11281]_  = \new_[11280]_  | \new_[11277]_ ;
  assign \new_[11282]_  = \new_[11281]_  | \new_[11274]_ ;
  assign \new_[11285]_  = \new_[112]_  | \new_[113]_ ;
  assign \new_[11288]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[11289]_  = \new_[11288]_  | \new_[11285]_ ;
  assign \new_[11292]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[11295]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[11296]_  = \new_[11295]_  | \new_[11292]_ ;
  assign \new_[11297]_  = \new_[11296]_  | \new_[11289]_ ;
  assign \new_[11298]_  = \new_[11297]_  | \new_[11282]_ ;
  assign \new_[11302]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[11303]_  = \new_[105]_  | \new_[11302]_ ;
  assign \new_[11306]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[11309]_  = \new_[99]_  | \new_[100]_ ;
  assign \new_[11310]_  = \new_[11309]_  | \new_[11306]_ ;
  assign \new_[11311]_  = \new_[11310]_  | \new_[11303]_ ;
  assign \new_[11314]_  = \new_[97]_  | \new_[98]_ ;
  assign \new_[11317]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[11318]_  = \new_[11317]_  | \new_[11314]_ ;
  assign \new_[11321]_  = \new_[93]_  | \new_[94]_ ;
  assign \new_[11324]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[11325]_  = \new_[11324]_  | \new_[11321]_ ;
  assign \new_[11326]_  = \new_[11325]_  | \new_[11318]_ ;
  assign \new_[11327]_  = \new_[11326]_  | \new_[11311]_ ;
  assign \new_[11328]_  = \new_[11327]_  | \new_[11298]_ ;
  assign \new_[11332]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[11333]_  = \new_[90]_  | \new_[11332]_ ;
  assign \new_[11336]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[11339]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[11340]_  = \new_[11339]_  | \new_[11336]_ ;
  assign \new_[11341]_  = \new_[11340]_  | \new_[11333]_ ;
  assign \new_[11344]_  = \new_[82]_  | \new_[83]_ ;
  assign \new_[11347]_  = \new_[80]_  | \new_[81]_ ;
  assign \new_[11348]_  = \new_[11347]_  | \new_[11344]_ ;
  assign \new_[11351]_  = \new_[78]_  | \new_[79]_ ;
  assign \new_[11354]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[11355]_  = \new_[11354]_  | \new_[11351]_ ;
  assign \new_[11356]_  = \new_[11355]_  | \new_[11348]_ ;
  assign \new_[11357]_  = \new_[11356]_  | \new_[11341]_ ;
  assign \new_[11361]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[11362]_  = \new_[75]_  | \new_[11361]_ ;
  assign \new_[11365]_  = \new_[71]_  | \new_[72]_ ;
  assign \new_[11368]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[11369]_  = \new_[11368]_  | \new_[11365]_ ;
  assign \new_[11370]_  = \new_[11369]_  | \new_[11362]_ ;
  assign \new_[11373]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[11376]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[11377]_  = \new_[11376]_  | \new_[11373]_ ;
  assign \new_[11380]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[11383]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[11384]_  = \new_[11383]_  | \new_[11380]_ ;
  assign \new_[11385]_  = \new_[11384]_  | \new_[11377]_ ;
  assign \new_[11386]_  = \new_[11385]_  | \new_[11370]_ ;
  assign \new_[11387]_  = \new_[11386]_  | \new_[11357]_ ;
  assign \new_[11388]_  = \new_[11387]_  | \new_[11328]_ ;
  assign \new_[11392]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[11393]_  = \new_[60]_  | \new_[11392]_ ;
  assign \new_[11396]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[11399]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[11400]_  = \new_[11399]_  | \new_[11396]_ ;
  assign \new_[11401]_  = \new_[11400]_  | \new_[11393]_ ;
  assign \new_[11404]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[11407]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[11408]_  = \new_[11407]_  | \new_[11404]_ ;
  assign \new_[11411]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[11414]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[11415]_  = \new_[11414]_  | \new_[11411]_ ;
  assign \new_[11416]_  = \new_[11415]_  | \new_[11408]_ ;
  assign \new_[11417]_  = \new_[11416]_  | \new_[11401]_ ;
  assign \new_[11421]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[11422]_  = \new_[45]_  | \new_[11421]_ ;
  assign \new_[11425]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[11428]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[11429]_  = \new_[11428]_  | \new_[11425]_ ;
  assign \new_[11430]_  = \new_[11429]_  | \new_[11422]_ ;
  assign \new_[11433]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[11436]_  = \new_[35]_  | \new_[36]_ ;
  assign \new_[11437]_  = \new_[11436]_  | \new_[11433]_ ;
  assign \new_[11440]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[11443]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[11444]_  = \new_[11443]_  | \new_[11440]_ ;
  assign \new_[11445]_  = \new_[11444]_  | \new_[11437]_ ;
  assign \new_[11446]_  = \new_[11445]_  | \new_[11430]_ ;
  assign \new_[11447]_  = \new_[11446]_  | \new_[11417]_ ;
  assign \new_[11451]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[11452]_  = \new_[30]_  | \new_[11451]_ ;
  assign \new_[11455]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[11458]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[11459]_  = \new_[11458]_  | \new_[11455]_ ;
  assign \new_[11460]_  = \new_[11459]_  | \new_[11452]_ ;
  assign \new_[11463]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[11466]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[11467]_  = \new_[11466]_  | \new_[11463]_ ;
  assign \new_[11470]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[11473]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[11474]_  = \new_[11473]_  | \new_[11470]_ ;
  assign \new_[11475]_  = \new_[11474]_  | \new_[11467]_ ;
  assign \new_[11476]_  = \new_[11475]_  | \new_[11460]_ ;
  assign \new_[11480]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[11481]_  = \new_[15]_  | \new_[11480]_ ;
  assign \new_[11484]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[11487]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[11488]_  = \new_[11487]_  | \new_[11484]_ ;
  assign \new_[11489]_  = \new_[11488]_  | \new_[11481]_ ;
  assign \new_[11492]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[11495]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[11496]_  = \new_[11495]_  | \new_[11492]_ ;
  assign \new_[11499]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[11502]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[11503]_  = \new_[11502]_  | \new_[11499]_ ;
  assign \new_[11504]_  = \new_[11503]_  | \new_[11496]_ ;
  assign \new_[11505]_  = \new_[11504]_  | \new_[11489]_ ;
  assign \new_[11506]_  = \new_[11505]_  | \new_[11476]_ ;
  assign \new_[11507]_  = \new_[11506]_  | \new_[11447]_ ;
  assign \new_[11508]_  = \new_[11507]_  | \new_[11388]_ ;
  assign \new_[11509]_  = \new_[11508]_  | \new_[11269]_ ;
  assign \new_[11510]_  = \new_[11509]_  | \new_[11030]_ ;
  assign \new_[11511]_  = \new_[11510]_  | \new_[10551]_ ;
  assign \new_[11512]_  = \new_[11511]_  | \new_[9592]_ ;
  assign \new_[11515]_  = A233 & ~A232;
  assign \new_[11518]_  = A235 & A234;
  assign \new_[11519]_  = \new_[11518]_  & \new_[11515]_ ;
  assign \new_[11522]_  = ~A299 & A298;
  assign \new_[11525]_  = A301 & A300;
  assign \new_[11526]_  = \new_[11525]_  & \new_[11522]_ ;
  assign \new_[11529]_  = A233 & ~A232;
  assign \new_[11532]_  = A235 & A234;
  assign \new_[11533]_  = \new_[11532]_  & \new_[11529]_ ;
  assign \new_[11536]_  = ~A299 & A298;
  assign \new_[11539]_  = ~A302 & A300;
  assign \new_[11540]_  = \new_[11539]_  & \new_[11536]_ ;
  assign \new_[11543]_  = A233 & ~A232;
  assign \new_[11546]_  = A235 & A234;
  assign \new_[11547]_  = \new_[11546]_  & \new_[11543]_ ;
  assign \new_[11550]_  = A299 & ~A298;
  assign \new_[11553]_  = A301 & A300;
  assign \new_[11554]_  = \new_[11553]_  & \new_[11550]_ ;
  assign \new_[11557]_  = A233 & ~A232;
  assign \new_[11560]_  = A235 & A234;
  assign \new_[11561]_  = \new_[11560]_  & \new_[11557]_ ;
  assign \new_[11564]_  = A299 & ~A298;
  assign \new_[11567]_  = ~A302 & A300;
  assign \new_[11568]_  = \new_[11567]_  & \new_[11564]_ ;
  assign \new_[11571]_  = A233 & ~A232;
  assign \new_[11574]_  = A235 & A234;
  assign \new_[11575]_  = \new_[11574]_  & \new_[11571]_ ;
  assign \new_[11578]_  = A266 & ~A265;
  assign \new_[11581]_  = A268 & A267;
  assign \new_[11582]_  = \new_[11581]_  & \new_[11578]_ ;
  assign \new_[11585]_  = A233 & ~A232;
  assign \new_[11588]_  = A235 & A234;
  assign \new_[11589]_  = \new_[11588]_  & \new_[11585]_ ;
  assign \new_[11592]_  = A266 & ~A265;
  assign \new_[11595]_  = ~A269 & A267;
  assign \new_[11596]_  = \new_[11595]_  & \new_[11592]_ ;
  assign \new_[11599]_  = A233 & ~A232;
  assign \new_[11602]_  = A235 & A234;
  assign \new_[11603]_  = \new_[11602]_  & \new_[11599]_ ;
  assign \new_[11606]_  = ~A266 & A265;
  assign \new_[11609]_  = A268 & A267;
  assign \new_[11610]_  = \new_[11609]_  & \new_[11606]_ ;
  assign \new_[11613]_  = A233 & ~A232;
  assign \new_[11616]_  = A235 & A234;
  assign \new_[11617]_  = \new_[11616]_  & \new_[11613]_ ;
  assign \new_[11620]_  = ~A266 & A265;
  assign \new_[11623]_  = ~A269 & A267;
  assign \new_[11624]_  = \new_[11623]_  & \new_[11620]_ ;
  assign \new_[11627]_  = A233 & ~A232;
  assign \new_[11630]_  = ~A236 & A234;
  assign \new_[11631]_  = \new_[11630]_  & \new_[11627]_ ;
  assign \new_[11634]_  = ~A299 & A298;
  assign \new_[11637]_  = A301 & A300;
  assign \new_[11638]_  = \new_[11637]_  & \new_[11634]_ ;
  assign \new_[11641]_  = A233 & ~A232;
  assign \new_[11644]_  = ~A236 & A234;
  assign \new_[11645]_  = \new_[11644]_  & \new_[11641]_ ;
  assign \new_[11648]_  = ~A299 & A298;
  assign \new_[11651]_  = ~A302 & A300;
  assign \new_[11652]_  = \new_[11651]_  & \new_[11648]_ ;
  assign \new_[11655]_  = A233 & ~A232;
  assign \new_[11658]_  = ~A236 & A234;
  assign \new_[11659]_  = \new_[11658]_  & \new_[11655]_ ;
  assign \new_[11662]_  = A299 & ~A298;
  assign \new_[11665]_  = A301 & A300;
  assign \new_[11666]_  = \new_[11665]_  & \new_[11662]_ ;
  assign \new_[11669]_  = A233 & ~A232;
  assign \new_[11672]_  = ~A236 & A234;
  assign \new_[11673]_  = \new_[11672]_  & \new_[11669]_ ;
  assign \new_[11676]_  = A299 & ~A298;
  assign \new_[11679]_  = ~A302 & A300;
  assign \new_[11680]_  = \new_[11679]_  & \new_[11676]_ ;
  assign \new_[11683]_  = A233 & ~A232;
  assign \new_[11686]_  = ~A236 & A234;
  assign \new_[11687]_  = \new_[11686]_  & \new_[11683]_ ;
  assign \new_[11690]_  = A266 & ~A265;
  assign \new_[11693]_  = A268 & A267;
  assign \new_[11694]_  = \new_[11693]_  & \new_[11690]_ ;
  assign \new_[11697]_  = A233 & ~A232;
  assign \new_[11700]_  = ~A236 & A234;
  assign \new_[11701]_  = \new_[11700]_  & \new_[11697]_ ;
  assign \new_[11704]_  = A266 & ~A265;
  assign \new_[11707]_  = ~A269 & A267;
  assign \new_[11708]_  = \new_[11707]_  & \new_[11704]_ ;
  assign \new_[11711]_  = A233 & ~A232;
  assign \new_[11714]_  = ~A236 & A234;
  assign \new_[11715]_  = \new_[11714]_  & \new_[11711]_ ;
  assign \new_[11718]_  = ~A266 & A265;
  assign \new_[11721]_  = A268 & A267;
  assign \new_[11722]_  = \new_[11721]_  & \new_[11718]_ ;
  assign \new_[11725]_  = A233 & ~A232;
  assign \new_[11728]_  = ~A236 & A234;
  assign \new_[11729]_  = \new_[11728]_  & \new_[11725]_ ;
  assign \new_[11732]_  = ~A266 & A265;
  assign \new_[11735]_  = ~A269 & A267;
  assign \new_[11736]_  = \new_[11735]_  & \new_[11732]_ ;
  assign \new_[11739]_  = ~A233 & A232;
  assign \new_[11742]_  = A235 & A234;
  assign \new_[11743]_  = \new_[11742]_  & \new_[11739]_ ;
  assign \new_[11746]_  = ~A299 & A298;
  assign \new_[11749]_  = A301 & A300;
  assign \new_[11750]_  = \new_[11749]_  & \new_[11746]_ ;
  assign \new_[11753]_  = ~A233 & A232;
  assign \new_[11756]_  = A235 & A234;
  assign \new_[11757]_  = \new_[11756]_  & \new_[11753]_ ;
  assign \new_[11760]_  = ~A299 & A298;
  assign \new_[11763]_  = ~A302 & A300;
  assign \new_[11764]_  = \new_[11763]_  & \new_[11760]_ ;
  assign \new_[11767]_  = ~A233 & A232;
  assign \new_[11770]_  = A235 & A234;
  assign \new_[11771]_  = \new_[11770]_  & \new_[11767]_ ;
  assign \new_[11774]_  = A299 & ~A298;
  assign \new_[11777]_  = A301 & A300;
  assign \new_[11778]_  = \new_[11777]_  & \new_[11774]_ ;
  assign \new_[11781]_  = ~A233 & A232;
  assign \new_[11784]_  = A235 & A234;
  assign \new_[11785]_  = \new_[11784]_  & \new_[11781]_ ;
  assign \new_[11788]_  = A299 & ~A298;
  assign \new_[11791]_  = ~A302 & A300;
  assign \new_[11792]_  = \new_[11791]_  & \new_[11788]_ ;
  assign \new_[11795]_  = ~A233 & A232;
  assign \new_[11798]_  = A235 & A234;
  assign \new_[11799]_  = \new_[11798]_  & \new_[11795]_ ;
  assign \new_[11802]_  = A266 & ~A265;
  assign \new_[11805]_  = A268 & A267;
  assign \new_[11806]_  = \new_[11805]_  & \new_[11802]_ ;
  assign \new_[11809]_  = ~A233 & A232;
  assign \new_[11812]_  = A235 & A234;
  assign \new_[11813]_  = \new_[11812]_  & \new_[11809]_ ;
  assign \new_[11816]_  = A266 & ~A265;
  assign \new_[11819]_  = ~A269 & A267;
  assign \new_[11820]_  = \new_[11819]_  & \new_[11816]_ ;
  assign \new_[11823]_  = ~A233 & A232;
  assign \new_[11826]_  = A235 & A234;
  assign \new_[11827]_  = \new_[11826]_  & \new_[11823]_ ;
  assign \new_[11830]_  = ~A266 & A265;
  assign \new_[11833]_  = A268 & A267;
  assign \new_[11834]_  = \new_[11833]_  & \new_[11830]_ ;
  assign \new_[11837]_  = ~A233 & A232;
  assign \new_[11840]_  = A235 & A234;
  assign \new_[11841]_  = \new_[11840]_  & \new_[11837]_ ;
  assign \new_[11844]_  = ~A266 & A265;
  assign \new_[11847]_  = ~A269 & A267;
  assign \new_[11848]_  = \new_[11847]_  & \new_[11844]_ ;
  assign \new_[11851]_  = ~A233 & A232;
  assign \new_[11854]_  = ~A236 & A234;
  assign \new_[11855]_  = \new_[11854]_  & \new_[11851]_ ;
  assign \new_[11858]_  = ~A299 & A298;
  assign \new_[11861]_  = A301 & A300;
  assign \new_[11862]_  = \new_[11861]_  & \new_[11858]_ ;
  assign \new_[11865]_  = ~A233 & A232;
  assign \new_[11868]_  = ~A236 & A234;
  assign \new_[11869]_  = \new_[11868]_  & \new_[11865]_ ;
  assign \new_[11872]_  = ~A299 & A298;
  assign \new_[11875]_  = ~A302 & A300;
  assign \new_[11876]_  = \new_[11875]_  & \new_[11872]_ ;
  assign \new_[11879]_  = ~A233 & A232;
  assign \new_[11882]_  = ~A236 & A234;
  assign \new_[11883]_  = \new_[11882]_  & \new_[11879]_ ;
  assign \new_[11886]_  = A299 & ~A298;
  assign \new_[11889]_  = A301 & A300;
  assign \new_[11890]_  = \new_[11889]_  & \new_[11886]_ ;
  assign \new_[11893]_  = ~A233 & A232;
  assign \new_[11896]_  = ~A236 & A234;
  assign \new_[11897]_  = \new_[11896]_  & \new_[11893]_ ;
  assign \new_[11900]_  = A299 & ~A298;
  assign \new_[11903]_  = ~A302 & A300;
  assign \new_[11904]_  = \new_[11903]_  & \new_[11900]_ ;
  assign \new_[11907]_  = ~A233 & A232;
  assign \new_[11910]_  = ~A236 & A234;
  assign \new_[11911]_  = \new_[11910]_  & \new_[11907]_ ;
  assign \new_[11914]_  = A266 & ~A265;
  assign \new_[11917]_  = A268 & A267;
  assign \new_[11918]_  = \new_[11917]_  & \new_[11914]_ ;
  assign \new_[11921]_  = ~A233 & A232;
  assign \new_[11924]_  = ~A236 & A234;
  assign \new_[11925]_  = \new_[11924]_  & \new_[11921]_ ;
  assign \new_[11928]_  = A266 & ~A265;
  assign \new_[11931]_  = ~A269 & A267;
  assign \new_[11932]_  = \new_[11931]_  & \new_[11928]_ ;
  assign \new_[11935]_  = ~A233 & A232;
  assign \new_[11938]_  = ~A236 & A234;
  assign \new_[11939]_  = \new_[11938]_  & \new_[11935]_ ;
  assign \new_[11942]_  = ~A266 & A265;
  assign \new_[11945]_  = A268 & A267;
  assign \new_[11946]_  = \new_[11945]_  & \new_[11942]_ ;
  assign \new_[11949]_  = ~A233 & A232;
  assign \new_[11952]_  = ~A236 & A234;
  assign \new_[11953]_  = \new_[11952]_  & \new_[11949]_ ;
  assign \new_[11956]_  = ~A266 & A265;
  assign \new_[11959]_  = ~A269 & A267;
  assign \new_[11960]_  = \new_[11959]_  & \new_[11956]_ ;
  assign \new_[11963]_  = A233 & ~A232;
  assign \new_[11966]_  = A235 & A234;
  assign \new_[11967]_  = \new_[11966]_  & \new_[11963]_ ;
  assign \new_[11970]_  = ~A299 & A298;
  assign \new_[11974]_  = A302 & ~A301;
  assign \new_[11975]_  = ~A300 & \new_[11974]_ ;
  assign \new_[11976]_  = \new_[11975]_  & \new_[11970]_ ;
  assign \new_[11979]_  = A233 & ~A232;
  assign \new_[11982]_  = A235 & A234;
  assign \new_[11983]_  = \new_[11982]_  & \new_[11979]_ ;
  assign \new_[11986]_  = A299 & ~A298;
  assign \new_[11990]_  = A302 & ~A301;
  assign \new_[11991]_  = ~A300 & \new_[11990]_ ;
  assign \new_[11992]_  = \new_[11991]_  & \new_[11986]_ ;
  assign \new_[11995]_  = A233 & ~A232;
  assign \new_[11998]_  = ~A236 & A234;
  assign \new_[11999]_  = \new_[11998]_  & \new_[11995]_ ;
  assign \new_[12002]_  = ~A299 & A298;
  assign \new_[12006]_  = A302 & ~A301;
  assign \new_[12007]_  = ~A300 & \new_[12006]_ ;
  assign \new_[12008]_  = \new_[12007]_  & \new_[12002]_ ;
  assign \new_[12011]_  = A233 & ~A232;
  assign \new_[12014]_  = ~A236 & A234;
  assign \new_[12015]_  = \new_[12014]_  & \new_[12011]_ ;
  assign \new_[12018]_  = A299 & ~A298;
  assign \new_[12022]_  = A302 & ~A301;
  assign \new_[12023]_  = ~A300 & \new_[12022]_ ;
  assign \new_[12024]_  = \new_[12023]_  & \new_[12018]_ ;
  assign \new_[12027]_  = A233 & ~A232;
  assign \new_[12030]_  = ~A235 & ~A234;
  assign \new_[12031]_  = \new_[12030]_  & \new_[12027]_ ;
  assign \new_[12034]_  = A298 & A236;
  assign \new_[12038]_  = A301 & A300;
  assign \new_[12039]_  = ~A299 & \new_[12038]_ ;
  assign \new_[12040]_  = \new_[12039]_  & \new_[12034]_ ;
  assign \new_[12043]_  = A233 & ~A232;
  assign \new_[12046]_  = ~A235 & ~A234;
  assign \new_[12047]_  = \new_[12046]_  & \new_[12043]_ ;
  assign \new_[12050]_  = A298 & A236;
  assign \new_[12054]_  = ~A302 & A300;
  assign \new_[12055]_  = ~A299 & \new_[12054]_ ;
  assign \new_[12056]_  = \new_[12055]_  & \new_[12050]_ ;
  assign \new_[12059]_  = A233 & ~A232;
  assign \new_[12062]_  = ~A235 & ~A234;
  assign \new_[12063]_  = \new_[12062]_  & \new_[12059]_ ;
  assign \new_[12066]_  = ~A298 & A236;
  assign \new_[12070]_  = A301 & A300;
  assign \new_[12071]_  = A299 & \new_[12070]_ ;
  assign \new_[12072]_  = \new_[12071]_  & \new_[12066]_ ;
  assign \new_[12075]_  = A233 & ~A232;
  assign \new_[12078]_  = ~A235 & ~A234;
  assign \new_[12079]_  = \new_[12078]_  & \new_[12075]_ ;
  assign \new_[12082]_  = ~A298 & A236;
  assign \new_[12086]_  = ~A302 & A300;
  assign \new_[12087]_  = A299 & \new_[12086]_ ;
  assign \new_[12088]_  = \new_[12087]_  & \new_[12082]_ ;
  assign \new_[12091]_  = A233 & ~A232;
  assign \new_[12094]_  = ~A235 & ~A234;
  assign \new_[12095]_  = \new_[12094]_  & \new_[12091]_ ;
  assign \new_[12098]_  = ~A265 & A236;
  assign \new_[12102]_  = A268 & A267;
  assign \new_[12103]_  = A266 & \new_[12102]_ ;
  assign \new_[12104]_  = \new_[12103]_  & \new_[12098]_ ;
  assign \new_[12107]_  = A233 & ~A232;
  assign \new_[12110]_  = ~A235 & ~A234;
  assign \new_[12111]_  = \new_[12110]_  & \new_[12107]_ ;
  assign \new_[12114]_  = ~A265 & A236;
  assign \new_[12118]_  = ~A269 & A267;
  assign \new_[12119]_  = A266 & \new_[12118]_ ;
  assign \new_[12120]_  = \new_[12119]_  & \new_[12114]_ ;
  assign \new_[12123]_  = A233 & ~A232;
  assign \new_[12126]_  = ~A235 & ~A234;
  assign \new_[12127]_  = \new_[12126]_  & \new_[12123]_ ;
  assign \new_[12130]_  = A265 & A236;
  assign \new_[12134]_  = A268 & A267;
  assign \new_[12135]_  = ~A266 & \new_[12134]_ ;
  assign \new_[12136]_  = \new_[12135]_  & \new_[12130]_ ;
  assign \new_[12139]_  = A233 & ~A232;
  assign \new_[12142]_  = ~A235 & ~A234;
  assign \new_[12143]_  = \new_[12142]_  & \new_[12139]_ ;
  assign \new_[12146]_  = A265 & A236;
  assign \new_[12150]_  = ~A269 & A267;
  assign \new_[12151]_  = ~A266 & \new_[12150]_ ;
  assign \new_[12152]_  = \new_[12151]_  & \new_[12146]_ ;
  assign \new_[12155]_  = ~A233 & A232;
  assign \new_[12158]_  = A235 & A234;
  assign \new_[12159]_  = \new_[12158]_  & \new_[12155]_ ;
  assign \new_[12162]_  = ~A299 & A298;
  assign \new_[12166]_  = A302 & ~A301;
  assign \new_[12167]_  = ~A300 & \new_[12166]_ ;
  assign \new_[12168]_  = \new_[12167]_  & \new_[12162]_ ;
  assign \new_[12171]_  = ~A233 & A232;
  assign \new_[12174]_  = A235 & A234;
  assign \new_[12175]_  = \new_[12174]_  & \new_[12171]_ ;
  assign \new_[12178]_  = A299 & ~A298;
  assign \new_[12182]_  = A302 & ~A301;
  assign \new_[12183]_  = ~A300 & \new_[12182]_ ;
  assign \new_[12184]_  = \new_[12183]_  & \new_[12178]_ ;
  assign \new_[12187]_  = ~A233 & A232;
  assign \new_[12190]_  = ~A236 & A234;
  assign \new_[12191]_  = \new_[12190]_  & \new_[12187]_ ;
  assign \new_[12194]_  = ~A299 & A298;
  assign \new_[12198]_  = A302 & ~A301;
  assign \new_[12199]_  = ~A300 & \new_[12198]_ ;
  assign \new_[12200]_  = \new_[12199]_  & \new_[12194]_ ;
  assign \new_[12203]_  = ~A233 & A232;
  assign \new_[12206]_  = ~A236 & A234;
  assign \new_[12207]_  = \new_[12206]_  & \new_[12203]_ ;
  assign \new_[12210]_  = A299 & ~A298;
  assign \new_[12214]_  = A302 & ~A301;
  assign \new_[12215]_  = ~A300 & \new_[12214]_ ;
  assign \new_[12216]_  = \new_[12215]_  & \new_[12210]_ ;
  assign \new_[12219]_  = ~A233 & A232;
  assign \new_[12222]_  = ~A235 & ~A234;
  assign \new_[12223]_  = \new_[12222]_  & \new_[12219]_ ;
  assign \new_[12226]_  = A298 & A236;
  assign \new_[12230]_  = A301 & A300;
  assign \new_[12231]_  = ~A299 & \new_[12230]_ ;
  assign \new_[12232]_  = \new_[12231]_  & \new_[12226]_ ;
  assign \new_[12235]_  = ~A233 & A232;
  assign \new_[12238]_  = ~A235 & ~A234;
  assign \new_[12239]_  = \new_[12238]_  & \new_[12235]_ ;
  assign \new_[12242]_  = A298 & A236;
  assign \new_[12246]_  = ~A302 & A300;
  assign \new_[12247]_  = ~A299 & \new_[12246]_ ;
  assign \new_[12248]_  = \new_[12247]_  & \new_[12242]_ ;
  assign \new_[12251]_  = ~A233 & A232;
  assign \new_[12254]_  = ~A235 & ~A234;
  assign \new_[12255]_  = \new_[12254]_  & \new_[12251]_ ;
  assign \new_[12258]_  = ~A298 & A236;
  assign \new_[12262]_  = A301 & A300;
  assign \new_[12263]_  = A299 & \new_[12262]_ ;
  assign \new_[12264]_  = \new_[12263]_  & \new_[12258]_ ;
  assign \new_[12267]_  = ~A233 & A232;
  assign \new_[12270]_  = ~A235 & ~A234;
  assign \new_[12271]_  = \new_[12270]_  & \new_[12267]_ ;
  assign \new_[12274]_  = ~A298 & A236;
  assign \new_[12278]_  = ~A302 & A300;
  assign \new_[12279]_  = A299 & \new_[12278]_ ;
  assign \new_[12280]_  = \new_[12279]_  & \new_[12274]_ ;
  assign \new_[12283]_  = ~A233 & A232;
  assign \new_[12286]_  = ~A235 & ~A234;
  assign \new_[12287]_  = \new_[12286]_  & \new_[12283]_ ;
  assign \new_[12290]_  = ~A265 & A236;
  assign \new_[12294]_  = A268 & A267;
  assign \new_[12295]_  = A266 & \new_[12294]_ ;
  assign \new_[12296]_  = \new_[12295]_  & \new_[12290]_ ;
  assign \new_[12299]_  = ~A233 & A232;
  assign \new_[12302]_  = ~A235 & ~A234;
  assign \new_[12303]_  = \new_[12302]_  & \new_[12299]_ ;
  assign \new_[12306]_  = ~A265 & A236;
  assign \new_[12310]_  = ~A269 & A267;
  assign \new_[12311]_  = A266 & \new_[12310]_ ;
  assign \new_[12312]_  = \new_[12311]_  & \new_[12306]_ ;
  assign \new_[12315]_  = ~A233 & A232;
  assign \new_[12318]_  = ~A235 & ~A234;
  assign \new_[12319]_  = \new_[12318]_  & \new_[12315]_ ;
  assign \new_[12322]_  = A265 & A236;
  assign \new_[12326]_  = A268 & A267;
  assign \new_[12327]_  = ~A266 & \new_[12326]_ ;
  assign \new_[12328]_  = \new_[12327]_  & \new_[12322]_ ;
  assign \new_[12331]_  = ~A233 & A232;
  assign \new_[12334]_  = ~A235 & ~A234;
  assign \new_[12335]_  = \new_[12334]_  & \new_[12331]_ ;
  assign \new_[12338]_  = A265 & A236;
  assign \new_[12342]_  = ~A269 & A267;
  assign \new_[12343]_  = ~A266 & \new_[12342]_ ;
  assign \new_[12344]_  = \new_[12343]_  & \new_[12338]_ ;
  assign \new_[12347]_  = A233 & ~A232;
  assign \new_[12351]_  = ~A265 & A235;
  assign \new_[12352]_  = A234 & \new_[12351]_ ;
  assign \new_[12353]_  = \new_[12352]_  & \new_[12347]_ ;
  assign \new_[12356]_  = ~A267 & A266;
  assign \new_[12360]_  = A300 & A269;
  assign \new_[12361]_  = ~A268 & \new_[12360]_ ;
  assign \new_[12362]_  = \new_[12361]_  & \new_[12356]_ ;
  assign \new_[12365]_  = A233 & ~A232;
  assign \new_[12369]_  = A265 & A235;
  assign \new_[12370]_  = A234 & \new_[12369]_ ;
  assign \new_[12371]_  = \new_[12370]_  & \new_[12365]_ ;
  assign \new_[12374]_  = ~A267 & ~A266;
  assign \new_[12378]_  = A300 & A269;
  assign \new_[12379]_  = ~A268 & \new_[12378]_ ;
  assign \new_[12380]_  = \new_[12379]_  & \new_[12374]_ ;
  assign \new_[12383]_  = A233 & ~A232;
  assign \new_[12387]_  = ~A265 & ~A236;
  assign \new_[12388]_  = A234 & \new_[12387]_ ;
  assign \new_[12389]_  = \new_[12388]_  & \new_[12383]_ ;
  assign \new_[12392]_  = ~A267 & A266;
  assign \new_[12396]_  = A300 & A269;
  assign \new_[12397]_  = ~A268 & \new_[12396]_ ;
  assign \new_[12398]_  = \new_[12397]_  & \new_[12392]_ ;
  assign \new_[12401]_  = A233 & ~A232;
  assign \new_[12405]_  = A265 & ~A236;
  assign \new_[12406]_  = A234 & \new_[12405]_ ;
  assign \new_[12407]_  = \new_[12406]_  & \new_[12401]_ ;
  assign \new_[12410]_  = ~A267 & ~A266;
  assign \new_[12414]_  = A300 & A269;
  assign \new_[12415]_  = ~A268 & \new_[12414]_ ;
  assign \new_[12416]_  = \new_[12415]_  & \new_[12410]_ ;
  assign \new_[12419]_  = A233 & ~A232;
  assign \new_[12423]_  = A236 & ~A235;
  assign \new_[12424]_  = ~A234 & \new_[12423]_ ;
  assign \new_[12425]_  = \new_[12424]_  & \new_[12419]_ ;
  assign \new_[12428]_  = ~A299 & A298;
  assign \new_[12432]_  = A302 & ~A301;
  assign \new_[12433]_  = ~A300 & \new_[12432]_ ;
  assign \new_[12434]_  = \new_[12433]_  & \new_[12428]_ ;
  assign \new_[12437]_  = A233 & ~A232;
  assign \new_[12441]_  = A236 & ~A235;
  assign \new_[12442]_  = ~A234 & \new_[12441]_ ;
  assign \new_[12443]_  = \new_[12442]_  & \new_[12437]_ ;
  assign \new_[12446]_  = A299 & ~A298;
  assign \new_[12450]_  = A302 & ~A301;
  assign \new_[12451]_  = ~A300 & \new_[12450]_ ;
  assign \new_[12452]_  = \new_[12451]_  & \new_[12446]_ ;
  assign \new_[12455]_  = ~A233 & A232;
  assign \new_[12459]_  = ~A265 & A235;
  assign \new_[12460]_  = A234 & \new_[12459]_ ;
  assign \new_[12461]_  = \new_[12460]_  & \new_[12455]_ ;
  assign \new_[12464]_  = ~A267 & A266;
  assign \new_[12468]_  = A300 & A269;
  assign \new_[12469]_  = ~A268 & \new_[12468]_ ;
  assign \new_[12470]_  = \new_[12469]_  & \new_[12464]_ ;
  assign \new_[12473]_  = ~A233 & A232;
  assign \new_[12477]_  = A265 & A235;
  assign \new_[12478]_  = A234 & \new_[12477]_ ;
  assign \new_[12479]_  = \new_[12478]_  & \new_[12473]_ ;
  assign \new_[12482]_  = ~A267 & ~A266;
  assign \new_[12486]_  = A300 & A269;
  assign \new_[12487]_  = ~A268 & \new_[12486]_ ;
  assign \new_[12488]_  = \new_[12487]_  & \new_[12482]_ ;
  assign \new_[12491]_  = ~A233 & A232;
  assign \new_[12495]_  = ~A265 & ~A236;
  assign \new_[12496]_  = A234 & \new_[12495]_ ;
  assign \new_[12497]_  = \new_[12496]_  & \new_[12491]_ ;
  assign \new_[12500]_  = ~A267 & A266;
  assign \new_[12504]_  = A300 & A269;
  assign \new_[12505]_  = ~A268 & \new_[12504]_ ;
  assign \new_[12506]_  = \new_[12505]_  & \new_[12500]_ ;
  assign \new_[12509]_  = ~A233 & A232;
  assign \new_[12513]_  = A265 & ~A236;
  assign \new_[12514]_  = A234 & \new_[12513]_ ;
  assign \new_[12515]_  = \new_[12514]_  & \new_[12509]_ ;
  assign \new_[12518]_  = ~A267 & ~A266;
  assign \new_[12522]_  = A300 & A269;
  assign \new_[12523]_  = ~A268 & \new_[12522]_ ;
  assign \new_[12524]_  = \new_[12523]_  & \new_[12518]_ ;
  assign \new_[12527]_  = ~A233 & A232;
  assign \new_[12531]_  = A236 & ~A235;
  assign \new_[12532]_  = ~A234 & \new_[12531]_ ;
  assign \new_[12533]_  = \new_[12532]_  & \new_[12527]_ ;
  assign \new_[12536]_  = ~A299 & A298;
  assign \new_[12540]_  = A302 & ~A301;
  assign \new_[12541]_  = ~A300 & \new_[12540]_ ;
  assign \new_[12542]_  = \new_[12541]_  & \new_[12536]_ ;
  assign \new_[12545]_  = ~A233 & A232;
  assign \new_[12549]_  = A236 & ~A235;
  assign \new_[12550]_  = ~A234 & \new_[12549]_ ;
  assign \new_[12551]_  = \new_[12550]_  & \new_[12545]_ ;
  assign \new_[12554]_  = A299 & ~A298;
  assign \new_[12558]_  = A302 & ~A301;
  assign \new_[12559]_  = ~A300 & \new_[12558]_ ;
  assign \new_[12560]_  = \new_[12559]_  & \new_[12554]_ ;
  assign \new_[12563]_  = ~A232 & ~A201;
  assign \new_[12567]_  = A235 & A234;
  assign \new_[12568]_  = A233 & \new_[12567]_ ;
  assign \new_[12569]_  = \new_[12568]_  & \new_[12563]_ ;
  assign \new_[12572]_  = A266 & ~A265;
  assign \new_[12576]_  = A269 & ~A268;
  assign \new_[12577]_  = ~A267 & \new_[12576]_ ;
  assign \new_[12578]_  = \new_[12577]_  & \new_[12572]_ ;
  assign \new_[12581]_  = ~A232 & ~A201;
  assign \new_[12585]_  = A235 & A234;
  assign \new_[12586]_  = A233 & \new_[12585]_ ;
  assign \new_[12587]_  = \new_[12586]_  & \new_[12581]_ ;
  assign \new_[12590]_  = ~A266 & A265;
  assign \new_[12594]_  = A269 & ~A268;
  assign \new_[12595]_  = ~A267 & \new_[12594]_ ;
  assign \new_[12596]_  = \new_[12595]_  & \new_[12590]_ ;
  assign \new_[12599]_  = ~A232 & ~A201;
  assign \new_[12603]_  = ~A236 & A234;
  assign \new_[12604]_  = A233 & \new_[12603]_ ;
  assign \new_[12605]_  = \new_[12604]_  & \new_[12599]_ ;
  assign \new_[12608]_  = A266 & ~A265;
  assign \new_[12612]_  = A269 & ~A268;
  assign \new_[12613]_  = ~A267 & \new_[12612]_ ;
  assign \new_[12614]_  = \new_[12613]_  & \new_[12608]_ ;
  assign \new_[12617]_  = ~A232 & ~A201;
  assign \new_[12621]_  = ~A236 & A234;
  assign \new_[12622]_  = A233 & \new_[12621]_ ;
  assign \new_[12623]_  = \new_[12622]_  & \new_[12617]_ ;
  assign \new_[12626]_  = ~A266 & A265;
  assign \new_[12630]_  = A269 & ~A268;
  assign \new_[12631]_  = ~A267 & \new_[12630]_ ;
  assign \new_[12632]_  = \new_[12631]_  & \new_[12626]_ ;
  assign \new_[12635]_  = A232 & ~A201;
  assign \new_[12639]_  = A235 & A234;
  assign \new_[12640]_  = ~A233 & \new_[12639]_ ;
  assign \new_[12641]_  = \new_[12640]_  & \new_[12635]_ ;
  assign \new_[12644]_  = A266 & ~A265;
  assign \new_[12648]_  = A269 & ~A268;
  assign \new_[12649]_  = ~A267 & \new_[12648]_ ;
  assign \new_[12650]_  = \new_[12649]_  & \new_[12644]_ ;
  assign \new_[12653]_  = A232 & ~A201;
  assign \new_[12657]_  = A235 & A234;
  assign \new_[12658]_  = ~A233 & \new_[12657]_ ;
  assign \new_[12659]_  = \new_[12658]_  & \new_[12653]_ ;
  assign \new_[12662]_  = ~A266 & A265;
  assign \new_[12666]_  = A269 & ~A268;
  assign \new_[12667]_  = ~A267 & \new_[12666]_ ;
  assign \new_[12668]_  = \new_[12667]_  & \new_[12662]_ ;
  assign \new_[12671]_  = A232 & ~A201;
  assign \new_[12675]_  = ~A236 & A234;
  assign \new_[12676]_  = ~A233 & \new_[12675]_ ;
  assign \new_[12677]_  = \new_[12676]_  & \new_[12671]_ ;
  assign \new_[12680]_  = A266 & ~A265;
  assign \new_[12684]_  = A269 & ~A268;
  assign \new_[12685]_  = ~A267 & \new_[12684]_ ;
  assign \new_[12686]_  = \new_[12685]_  & \new_[12680]_ ;
  assign \new_[12689]_  = A232 & ~A201;
  assign \new_[12693]_  = ~A236 & A234;
  assign \new_[12694]_  = ~A233 & \new_[12693]_ ;
  assign \new_[12695]_  = \new_[12694]_  & \new_[12689]_ ;
  assign \new_[12698]_  = ~A266 & A265;
  assign \new_[12702]_  = A269 & ~A268;
  assign \new_[12703]_  = ~A267 & \new_[12702]_ ;
  assign \new_[12704]_  = \new_[12703]_  & \new_[12698]_ ;
  assign \new_[12707]_  = A166 & A167;
  assign \new_[12711]_  = A201 & A200;
  assign \new_[12712]_  = ~A199 & \new_[12711]_ ;
  assign \new_[12713]_  = \new_[12712]_  & \new_[12707]_ ;
  assign \new_[12716]_  = ~A267 & A202;
  assign \new_[12720]_  = A301 & ~A300;
  assign \new_[12721]_  = A268 & \new_[12720]_ ;
  assign \new_[12722]_  = \new_[12721]_  & \new_[12716]_ ;
  assign \new_[12725]_  = A166 & A167;
  assign \new_[12729]_  = A201 & A200;
  assign \new_[12730]_  = ~A199 & \new_[12729]_ ;
  assign \new_[12731]_  = \new_[12730]_  & \new_[12725]_ ;
  assign \new_[12734]_  = ~A267 & A202;
  assign \new_[12738]_  = ~A302 & ~A300;
  assign \new_[12739]_  = A268 & \new_[12738]_ ;
  assign \new_[12740]_  = \new_[12739]_  & \new_[12734]_ ;
  assign \new_[12743]_  = A166 & A167;
  assign \new_[12747]_  = A201 & A200;
  assign \new_[12748]_  = ~A199 & \new_[12747]_ ;
  assign \new_[12749]_  = \new_[12748]_  & \new_[12743]_ ;
  assign \new_[12752]_  = ~A267 & A202;
  assign \new_[12756]_  = A299 & A298;
  assign \new_[12757]_  = A268 & \new_[12756]_ ;
  assign \new_[12758]_  = \new_[12757]_  & \new_[12752]_ ;
  assign \new_[12761]_  = A166 & A167;
  assign \new_[12765]_  = A201 & A200;
  assign \new_[12766]_  = ~A199 & \new_[12765]_ ;
  assign \new_[12767]_  = \new_[12766]_  & \new_[12761]_ ;
  assign \new_[12770]_  = ~A267 & A202;
  assign \new_[12774]_  = ~A299 & ~A298;
  assign \new_[12775]_  = A268 & \new_[12774]_ ;
  assign \new_[12776]_  = \new_[12775]_  & \new_[12770]_ ;
  assign \new_[12779]_  = A166 & A167;
  assign \new_[12783]_  = A201 & A200;
  assign \new_[12784]_  = ~A199 & \new_[12783]_ ;
  assign \new_[12785]_  = \new_[12784]_  & \new_[12779]_ ;
  assign \new_[12788]_  = ~A267 & A202;
  assign \new_[12792]_  = A301 & ~A300;
  assign \new_[12793]_  = ~A269 & \new_[12792]_ ;
  assign \new_[12794]_  = \new_[12793]_  & \new_[12788]_ ;
  assign \new_[12797]_  = A166 & A167;
  assign \new_[12801]_  = A201 & A200;
  assign \new_[12802]_  = ~A199 & \new_[12801]_ ;
  assign \new_[12803]_  = \new_[12802]_  & \new_[12797]_ ;
  assign \new_[12806]_  = ~A267 & A202;
  assign \new_[12810]_  = ~A302 & ~A300;
  assign \new_[12811]_  = ~A269 & \new_[12810]_ ;
  assign \new_[12812]_  = \new_[12811]_  & \new_[12806]_ ;
  assign \new_[12815]_  = A166 & A167;
  assign \new_[12819]_  = A201 & A200;
  assign \new_[12820]_  = ~A199 & \new_[12819]_ ;
  assign \new_[12821]_  = \new_[12820]_  & \new_[12815]_ ;
  assign \new_[12824]_  = ~A267 & A202;
  assign \new_[12828]_  = A299 & A298;
  assign \new_[12829]_  = ~A269 & \new_[12828]_ ;
  assign \new_[12830]_  = \new_[12829]_  & \new_[12824]_ ;
  assign \new_[12833]_  = A166 & A167;
  assign \new_[12837]_  = A201 & A200;
  assign \new_[12838]_  = ~A199 & \new_[12837]_ ;
  assign \new_[12839]_  = \new_[12838]_  & \new_[12833]_ ;
  assign \new_[12842]_  = ~A267 & A202;
  assign \new_[12846]_  = ~A299 & ~A298;
  assign \new_[12847]_  = ~A269 & \new_[12846]_ ;
  assign \new_[12848]_  = \new_[12847]_  & \new_[12842]_ ;
  assign \new_[12851]_  = A166 & A167;
  assign \new_[12855]_  = A201 & A200;
  assign \new_[12856]_  = ~A199 & \new_[12855]_ ;
  assign \new_[12857]_  = \new_[12856]_  & \new_[12851]_ ;
  assign \new_[12860]_  = A265 & A202;
  assign \new_[12864]_  = A301 & ~A300;
  assign \new_[12865]_  = A266 & \new_[12864]_ ;
  assign \new_[12866]_  = \new_[12865]_  & \new_[12860]_ ;
  assign \new_[12869]_  = A166 & A167;
  assign \new_[12873]_  = A201 & A200;
  assign \new_[12874]_  = ~A199 & \new_[12873]_ ;
  assign \new_[12875]_  = \new_[12874]_  & \new_[12869]_ ;
  assign \new_[12878]_  = A265 & A202;
  assign \new_[12882]_  = ~A302 & ~A300;
  assign \new_[12883]_  = A266 & \new_[12882]_ ;
  assign \new_[12884]_  = \new_[12883]_  & \new_[12878]_ ;
  assign \new_[12887]_  = A166 & A167;
  assign \new_[12891]_  = A201 & A200;
  assign \new_[12892]_  = ~A199 & \new_[12891]_ ;
  assign \new_[12893]_  = \new_[12892]_  & \new_[12887]_ ;
  assign \new_[12896]_  = A265 & A202;
  assign \new_[12900]_  = A299 & A298;
  assign \new_[12901]_  = A266 & \new_[12900]_ ;
  assign \new_[12902]_  = \new_[12901]_  & \new_[12896]_ ;
  assign \new_[12905]_  = A166 & A167;
  assign \new_[12909]_  = A201 & A200;
  assign \new_[12910]_  = ~A199 & \new_[12909]_ ;
  assign \new_[12911]_  = \new_[12910]_  & \new_[12905]_ ;
  assign \new_[12914]_  = A265 & A202;
  assign \new_[12918]_  = ~A299 & ~A298;
  assign \new_[12919]_  = A266 & \new_[12918]_ ;
  assign \new_[12920]_  = \new_[12919]_  & \new_[12914]_ ;
  assign \new_[12923]_  = A166 & A167;
  assign \new_[12927]_  = A201 & A200;
  assign \new_[12928]_  = ~A199 & \new_[12927]_ ;
  assign \new_[12929]_  = \new_[12928]_  & \new_[12923]_ ;
  assign \new_[12932]_  = ~A265 & A202;
  assign \new_[12936]_  = A301 & ~A300;
  assign \new_[12937]_  = ~A266 & \new_[12936]_ ;
  assign \new_[12938]_  = \new_[12937]_  & \new_[12932]_ ;
  assign \new_[12941]_  = A166 & A167;
  assign \new_[12945]_  = A201 & A200;
  assign \new_[12946]_  = ~A199 & \new_[12945]_ ;
  assign \new_[12947]_  = \new_[12946]_  & \new_[12941]_ ;
  assign \new_[12950]_  = ~A265 & A202;
  assign \new_[12954]_  = ~A302 & ~A300;
  assign \new_[12955]_  = ~A266 & \new_[12954]_ ;
  assign \new_[12956]_  = \new_[12955]_  & \new_[12950]_ ;
  assign \new_[12959]_  = A166 & A167;
  assign \new_[12963]_  = A201 & A200;
  assign \new_[12964]_  = ~A199 & \new_[12963]_ ;
  assign \new_[12965]_  = \new_[12964]_  & \new_[12959]_ ;
  assign \new_[12968]_  = ~A265 & A202;
  assign \new_[12972]_  = A299 & A298;
  assign \new_[12973]_  = ~A266 & \new_[12972]_ ;
  assign \new_[12974]_  = \new_[12973]_  & \new_[12968]_ ;
  assign \new_[12977]_  = A166 & A167;
  assign \new_[12981]_  = A201 & A200;
  assign \new_[12982]_  = ~A199 & \new_[12981]_ ;
  assign \new_[12983]_  = \new_[12982]_  & \new_[12977]_ ;
  assign \new_[12986]_  = ~A265 & A202;
  assign \new_[12990]_  = ~A299 & ~A298;
  assign \new_[12991]_  = ~A266 & \new_[12990]_ ;
  assign \new_[12992]_  = \new_[12991]_  & \new_[12986]_ ;
  assign \new_[12995]_  = A166 & A167;
  assign \new_[12999]_  = A201 & A200;
  assign \new_[13000]_  = ~A199 & \new_[12999]_ ;
  assign \new_[13001]_  = \new_[13000]_  & \new_[12995]_ ;
  assign \new_[13004]_  = ~A267 & ~A203;
  assign \new_[13008]_  = A301 & ~A300;
  assign \new_[13009]_  = A268 & \new_[13008]_ ;
  assign \new_[13010]_  = \new_[13009]_  & \new_[13004]_ ;
  assign \new_[13013]_  = A166 & A167;
  assign \new_[13017]_  = A201 & A200;
  assign \new_[13018]_  = ~A199 & \new_[13017]_ ;
  assign \new_[13019]_  = \new_[13018]_  & \new_[13013]_ ;
  assign \new_[13022]_  = ~A267 & ~A203;
  assign \new_[13026]_  = ~A302 & ~A300;
  assign \new_[13027]_  = A268 & \new_[13026]_ ;
  assign \new_[13028]_  = \new_[13027]_  & \new_[13022]_ ;
  assign \new_[13031]_  = A166 & A167;
  assign \new_[13035]_  = A201 & A200;
  assign \new_[13036]_  = ~A199 & \new_[13035]_ ;
  assign \new_[13037]_  = \new_[13036]_  & \new_[13031]_ ;
  assign \new_[13040]_  = ~A267 & ~A203;
  assign \new_[13044]_  = A299 & A298;
  assign \new_[13045]_  = A268 & \new_[13044]_ ;
  assign \new_[13046]_  = \new_[13045]_  & \new_[13040]_ ;
  assign \new_[13049]_  = A166 & A167;
  assign \new_[13053]_  = A201 & A200;
  assign \new_[13054]_  = ~A199 & \new_[13053]_ ;
  assign \new_[13055]_  = \new_[13054]_  & \new_[13049]_ ;
  assign \new_[13058]_  = ~A267 & ~A203;
  assign \new_[13062]_  = ~A299 & ~A298;
  assign \new_[13063]_  = A268 & \new_[13062]_ ;
  assign \new_[13064]_  = \new_[13063]_  & \new_[13058]_ ;
  assign \new_[13067]_  = A166 & A167;
  assign \new_[13071]_  = A201 & A200;
  assign \new_[13072]_  = ~A199 & \new_[13071]_ ;
  assign \new_[13073]_  = \new_[13072]_  & \new_[13067]_ ;
  assign \new_[13076]_  = ~A267 & ~A203;
  assign \new_[13080]_  = A301 & ~A300;
  assign \new_[13081]_  = ~A269 & \new_[13080]_ ;
  assign \new_[13082]_  = \new_[13081]_  & \new_[13076]_ ;
  assign \new_[13085]_  = A166 & A167;
  assign \new_[13089]_  = A201 & A200;
  assign \new_[13090]_  = ~A199 & \new_[13089]_ ;
  assign \new_[13091]_  = \new_[13090]_  & \new_[13085]_ ;
  assign \new_[13094]_  = ~A267 & ~A203;
  assign \new_[13098]_  = ~A302 & ~A300;
  assign \new_[13099]_  = ~A269 & \new_[13098]_ ;
  assign \new_[13100]_  = \new_[13099]_  & \new_[13094]_ ;
  assign \new_[13103]_  = A166 & A167;
  assign \new_[13107]_  = A201 & A200;
  assign \new_[13108]_  = ~A199 & \new_[13107]_ ;
  assign \new_[13109]_  = \new_[13108]_  & \new_[13103]_ ;
  assign \new_[13112]_  = ~A267 & ~A203;
  assign \new_[13116]_  = A299 & A298;
  assign \new_[13117]_  = ~A269 & \new_[13116]_ ;
  assign \new_[13118]_  = \new_[13117]_  & \new_[13112]_ ;
  assign \new_[13121]_  = A166 & A167;
  assign \new_[13125]_  = A201 & A200;
  assign \new_[13126]_  = ~A199 & \new_[13125]_ ;
  assign \new_[13127]_  = \new_[13126]_  & \new_[13121]_ ;
  assign \new_[13130]_  = ~A267 & ~A203;
  assign \new_[13134]_  = ~A299 & ~A298;
  assign \new_[13135]_  = ~A269 & \new_[13134]_ ;
  assign \new_[13136]_  = \new_[13135]_  & \new_[13130]_ ;
  assign \new_[13139]_  = A166 & A167;
  assign \new_[13143]_  = A201 & A200;
  assign \new_[13144]_  = ~A199 & \new_[13143]_ ;
  assign \new_[13145]_  = \new_[13144]_  & \new_[13139]_ ;
  assign \new_[13148]_  = A265 & ~A203;
  assign \new_[13152]_  = A301 & ~A300;
  assign \new_[13153]_  = A266 & \new_[13152]_ ;
  assign \new_[13154]_  = \new_[13153]_  & \new_[13148]_ ;
  assign \new_[13157]_  = A166 & A167;
  assign \new_[13161]_  = A201 & A200;
  assign \new_[13162]_  = ~A199 & \new_[13161]_ ;
  assign \new_[13163]_  = \new_[13162]_  & \new_[13157]_ ;
  assign \new_[13166]_  = A265 & ~A203;
  assign \new_[13170]_  = ~A302 & ~A300;
  assign \new_[13171]_  = A266 & \new_[13170]_ ;
  assign \new_[13172]_  = \new_[13171]_  & \new_[13166]_ ;
  assign \new_[13175]_  = A166 & A167;
  assign \new_[13179]_  = A201 & A200;
  assign \new_[13180]_  = ~A199 & \new_[13179]_ ;
  assign \new_[13181]_  = \new_[13180]_  & \new_[13175]_ ;
  assign \new_[13184]_  = A265 & ~A203;
  assign \new_[13188]_  = A299 & A298;
  assign \new_[13189]_  = A266 & \new_[13188]_ ;
  assign \new_[13190]_  = \new_[13189]_  & \new_[13184]_ ;
  assign \new_[13193]_  = A166 & A167;
  assign \new_[13197]_  = A201 & A200;
  assign \new_[13198]_  = ~A199 & \new_[13197]_ ;
  assign \new_[13199]_  = \new_[13198]_  & \new_[13193]_ ;
  assign \new_[13202]_  = A265 & ~A203;
  assign \new_[13206]_  = ~A299 & ~A298;
  assign \new_[13207]_  = A266 & \new_[13206]_ ;
  assign \new_[13208]_  = \new_[13207]_  & \new_[13202]_ ;
  assign \new_[13211]_  = A166 & A167;
  assign \new_[13215]_  = A201 & A200;
  assign \new_[13216]_  = ~A199 & \new_[13215]_ ;
  assign \new_[13217]_  = \new_[13216]_  & \new_[13211]_ ;
  assign \new_[13220]_  = ~A265 & ~A203;
  assign \new_[13224]_  = A301 & ~A300;
  assign \new_[13225]_  = ~A266 & \new_[13224]_ ;
  assign \new_[13226]_  = \new_[13225]_  & \new_[13220]_ ;
  assign \new_[13229]_  = A166 & A167;
  assign \new_[13233]_  = A201 & A200;
  assign \new_[13234]_  = ~A199 & \new_[13233]_ ;
  assign \new_[13235]_  = \new_[13234]_  & \new_[13229]_ ;
  assign \new_[13238]_  = ~A265 & ~A203;
  assign \new_[13242]_  = ~A302 & ~A300;
  assign \new_[13243]_  = ~A266 & \new_[13242]_ ;
  assign \new_[13244]_  = \new_[13243]_  & \new_[13238]_ ;
  assign \new_[13247]_  = A166 & A167;
  assign \new_[13251]_  = A201 & A200;
  assign \new_[13252]_  = ~A199 & \new_[13251]_ ;
  assign \new_[13253]_  = \new_[13252]_  & \new_[13247]_ ;
  assign \new_[13256]_  = ~A265 & ~A203;
  assign \new_[13260]_  = A299 & A298;
  assign \new_[13261]_  = ~A266 & \new_[13260]_ ;
  assign \new_[13262]_  = \new_[13261]_  & \new_[13256]_ ;
  assign \new_[13265]_  = A166 & A167;
  assign \new_[13269]_  = A201 & A200;
  assign \new_[13270]_  = ~A199 & \new_[13269]_ ;
  assign \new_[13271]_  = \new_[13270]_  & \new_[13265]_ ;
  assign \new_[13274]_  = ~A265 & ~A203;
  assign \new_[13278]_  = ~A299 & ~A298;
  assign \new_[13279]_  = ~A266 & \new_[13278]_ ;
  assign \new_[13280]_  = \new_[13279]_  & \new_[13274]_ ;
  assign \new_[13283]_  = A166 & A167;
  assign \new_[13287]_  = A201 & ~A200;
  assign \new_[13288]_  = A199 & \new_[13287]_ ;
  assign \new_[13289]_  = \new_[13288]_  & \new_[13283]_ ;
  assign \new_[13292]_  = ~A267 & A202;
  assign \new_[13296]_  = A301 & ~A300;
  assign \new_[13297]_  = A268 & \new_[13296]_ ;
  assign \new_[13298]_  = \new_[13297]_  & \new_[13292]_ ;
  assign \new_[13301]_  = A166 & A167;
  assign \new_[13305]_  = A201 & ~A200;
  assign \new_[13306]_  = A199 & \new_[13305]_ ;
  assign \new_[13307]_  = \new_[13306]_  & \new_[13301]_ ;
  assign \new_[13310]_  = ~A267 & A202;
  assign \new_[13314]_  = ~A302 & ~A300;
  assign \new_[13315]_  = A268 & \new_[13314]_ ;
  assign \new_[13316]_  = \new_[13315]_  & \new_[13310]_ ;
  assign \new_[13319]_  = A166 & A167;
  assign \new_[13323]_  = A201 & ~A200;
  assign \new_[13324]_  = A199 & \new_[13323]_ ;
  assign \new_[13325]_  = \new_[13324]_  & \new_[13319]_ ;
  assign \new_[13328]_  = ~A267 & A202;
  assign \new_[13332]_  = A299 & A298;
  assign \new_[13333]_  = A268 & \new_[13332]_ ;
  assign \new_[13334]_  = \new_[13333]_  & \new_[13328]_ ;
  assign \new_[13337]_  = A166 & A167;
  assign \new_[13341]_  = A201 & ~A200;
  assign \new_[13342]_  = A199 & \new_[13341]_ ;
  assign \new_[13343]_  = \new_[13342]_  & \new_[13337]_ ;
  assign \new_[13346]_  = ~A267 & A202;
  assign \new_[13350]_  = ~A299 & ~A298;
  assign \new_[13351]_  = A268 & \new_[13350]_ ;
  assign \new_[13352]_  = \new_[13351]_  & \new_[13346]_ ;
  assign \new_[13355]_  = A166 & A167;
  assign \new_[13359]_  = A201 & ~A200;
  assign \new_[13360]_  = A199 & \new_[13359]_ ;
  assign \new_[13361]_  = \new_[13360]_  & \new_[13355]_ ;
  assign \new_[13364]_  = ~A267 & A202;
  assign \new_[13368]_  = A301 & ~A300;
  assign \new_[13369]_  = ~A269 & \new_[13368]_ ;
  assign \new_[13370]_  = \new_[13369]_  & \new_[13364]_ ;
  assign \new_[13373]_  = A166 & A167;
  assign \new_[13377]_  = A201 & ~A200;
  assign \new_[13378]_  = A199 & \new_[13377]_ ;
  assign \new_[13379]_  = \new_[13378]_  & \new_[13373]_ ;
  assign \new_[13382]_  = ~A267 & A202;
  assign \new_[13386]_  = ~A302 & ~A300;
  assign \new_[13387]_  = ~A269 & \new_[13386]_ ;
  assign \new_[13388]_  = \new_[13387]_  & \new_[13382]_ ;
  assign \new_[13391]_  = A166 & A167;
  assign \new_[13395]_  = A201 & ~A200;
  assign \new_[13396]_  = A199 & \new_[13395]_ ;
  assign \new_[13397]_  = \new_[13396]_  & \new_[13391]_ ;
  assign \new_[13400]_  = ~A267 & A202;
  assign \new_[13404]_  = A299 & A298;
  assign \new_[13405]_  = ~A269 & \new_[13404]_ ;
  assign \new_[13406]_  = \new_[13405]_  & \new_[13400]_ ;
  assign \new_[13409]_  = A166 & A167;
  assign \new_[13413]_  = A201 & ~A200;
  assign \new_[13414]_  = A199 & \new_[13413]_ ;
  assign \new_[13415]_  = \new_[13414]_  & \new_[13409]_ ;
  assign \new_[13418]_  = ~A267 & A202;
  assign \new_[13422]_  = ~A299 & ~A298;
  assign \new_[13423]_  = ~A269 & \new_[13422]_ ;
  assign \new_[13424]_  = \new_[13423]_  & \new_[13418]_ ;
  assign \new_[13427]_  = A166 & A167;
  assign \new_[13431]_  = A201 & ~A200;
  assign \new_[13432]_  = A199 & \new_[13431]_ ;
  assign \new_[13433]_  = \new_[13432]_  & \new_[13427]_ ;
  assign \new_[13436]_  = A265 & A202;
  assign \new_[13440]_  = A301 & ~A300;
  assign \new_[13441]_  = A266 & \new_[13440]_ ;
  assign \new_[13442]_  = \new_[13441]_  & \new_[13436]_ ;
  assign \new_[13445]_  = A166 & A167;
  assign \new_[13449]_  = A201 & ~A200;
  assign \new_[13450]_  = A199 & \new_[13449]_ ;
  assign \new_[13451]_  = \new_[13450]_  & \new_[13445]_ ;
  assign \new_[13454]_  = A265 & A202;
  assign \new_[13458]_  = ~A302 & ~A300;
  assign \new_[13459]_  = A266 & \new_[13458]_ ;
  assign \new_[13460]_  = \new_[13459]_  & \new_[13454]_ ;
  assign \new_[13463]_  = A166 & A167;
  assign \new_[13467]_  = A201 & ~A200;
  assign \new_[13468]_  = A199 & \new_[13467]_ ;
  assign \new_[13469]_  = \new_[13468]_  & \new_[13463]_ ;
  assign \new_[13472]_  = A265 & A202;
  assign \new_[13476]_  = A299 & A298;
  assign \new_[13477]_  = A266 & \new_[13476]_ ;
  assign \new_[13478]_  = \new_[13477]_  & \new_[13472]_ ;
  assign \new_[13481]_  = A166 & A167;
  assign \new_[13485]_  = A201 & ~A200;
  assign \new_[13486]_  = A199 & \new_[13485]_ ;
  assign \new_[13487]_  = \new_[13486]_  & \new_[13481]_ ;
  assign \new_[13490]_  = A265 & A202;
  assign \new_[13494]_  = ~A299 & ~A298;
  assign \new_[13495]_  = A266 & \new_[13494]_ ;
  assign \new_[13496]_  = \new_[13495]_  & \new_[13490]_ ;
  assign \new_[13499]_  = A166 & A167;
  assign \new_[13503]_  = A201 & ~A200;
  assign \new_[13504]_  = A199 & \new_[13503]_ ;
  assign \new_[13505]_  = \new_[13504]_  & \new_[13499]_ ;
  assign \new_[13508]_  = ~A265 & A202;
  assign \new_[13512]_  = A301 & ~A300;
  assign \new_[13513]_  = ~A266 & \new_[13512]_ ;
  assign \new_[13514]_  = \new_[13513]_  & \new_[13508]_ ;
  assign \new_[13517]_  = A166 & A167;
  assign \new_[13521]_  = A201 & ~A200;
  assign \new_[13522]_  = A199 & \new_[13521]_ ;
  assign \new_[13523]_  = \new_[13522]_  & \new_[13517]_ ;
  assign \new_[13526]_  = ~A265 & A202;
  assign \new_[13530]_  = ~A302 & ~A300;
  assign \new_[13531]_  = ~A266 & \new_[13530]_ ;
  assign \new_[13532]_  = \new_[13531]_  & \new_[13526]_ ;
  assign \new_[13535]_  = A166 & A167;
  assign \new_[13539]_  = A201 & ~A200;
  assign \new_[13540]_  = A199 & \new_[13539]_ ;
  assign \new_[13541]_  = \new_[13540]_  & \new_[13535]_ ;
  assign \new_[13544]_  = ~A265 & A202;
  assign \new_[13548]_  = A299 & A298;
  assign \new_[13549]_  = ~A266 & \new_[13548]_ ;
  assign \new_[13550]_  = \new_[13549]_  & \new_[13544]_ ;
  assign \new_[13553]_  = A166 & A167;
  assign \new_[13557]_  = A201 & ~A200;
  assign \new_[13558]_  = A199 & \new_[13557]_ ;
  assign \new_[13559]_  = \new_[13558]_  & \new_[13553]_ ;
  assign \new_[13562]_  = ~A265 & A202;
  assign \new_[13566]_  = ~A299 & ~A298;
  assign \new_[13567]_  = ~A266 & \new_[13566]_ ;
  assign \new_[13568]_  = \new_[13567]_  & \new_[13562]_ ;
  assign \new_[13571]_  = A166 & A167;
  assign \new_[13575]_  = A201 & ~A200;
  assign \new_[13576]_  = A199 & \new_[13575]_ ;
  assign \new_[13577]_  = \new_[13576]_  & \new_[13571]_ ;
  assign \new_[13580]_  = ~A267 & ~A203;
  assign \new_[13584]_  = A301 & ~A300;
  assign \new_[13585]_  = A268 & \new_[13584]_ ;
  assign \new_[13586]_  = \new_[13585]_  & \new_[13580]_ ;
  assign \new_[13589]_  = A166 & A167;
  assign \new_[13593]_  = A201 & ~A200;
  assign \new_[13594]_  = A199 & \new_[13593]_ ;
  assign \new_[13595]_  = \new_[13594]_  & \new_[13589]_ ;
  assign \new_[13598]_  = ~A267 & ~A203;
  assign \new_[13602]_  = ~A302 & ~A300;
  assign \new_[13603]_  = A268 & \new_[13602]_ ;
  assign \new_[13604]_  = \new_[13603]_  & \new_[13598]_ ;
  assign \new_[13607]_  = A166 & A167;
  assign \new_[13611]_  = A201 & ~A200;
  assign \new_[13612]_  = A199 & \new_[13611]_ ;
  assign \new_[13613]_  = \new_[13612]_  & \new_[13607]_ ;
  assign \new_[13616]_  = ~A267 & ~A203;
  assign \new_[13620]_  = A299 & A298;
  assign \new_[13621]_  = A268 & \new_[13620]_ ;
  assign \new_[13622]_  = \new_[13621]_  & \new_[13616]_ ;
  assign \new_[13625]_  = A166 & A167;
  assign \new_[13629]_  = A201 & ~A200;
  assign \new_[13630]_  = A199 & \new_[13629]_ ;
  assign \new_[13631]_  = \new_[13630]_  & \new_[13625]_ ;
  assign \new_[13634]_  = ~A267 & ~A203;
  assign \new_[13638]_  = ~A299 & ~A298;
  assign \new_[13639]_  = A268 & \new_[13638]_ ;
  assign \new_[13640]_  = \new_[13639]_  & \new_[13634]_ ;
  assign \new_[13643]_  = A166 & A167;
  assign \new_[13647]_  = A201 & ~A200;
  assign \new_[13648]_  = A199 & \new_[13647]_ ;
  assign \new_[13649]_  = \new_[13648]_  & \new_[13643]_ ;
  assign \new_[13652]_  = ~A267 & ~A203;
  assign \new_[13656]_  = A301 & ~A300;
  assign \new_[13657]_  = ~A269 & \new_[13656]_ ;
  assign \new_[13658]_  = \new_[13657]_  & \new_[13652]_ ;
  assign \new_[13661]_  = A166 & A167;
  assign \new_[13665]_  = A201 & ~A200;
  assign \new_[13666]_  = A199 & \new_[13665]_ ;
  assign \new_[13667]_  = \new_[13666]_  & \new_[13661]_ ;
  assign \new_[13670]_  = ~A267 & ~A203;
  assign \new_[13674]_  = ~A302 & ~A300;
  assign \new_[13675]_  = ~A269 & \new_[13674]_ ;
  assign \new_[13676]_  = \new_[13675]_  & \new_[13670]_ ;
  assign \new_[13679]_  = A166 & A167;
  assign \new_[13683]_  = A201 & ~A200;
  assign \new_[13684]_  = A199 & \new_[13683]_ ;
  assign \new_[13685]_  = \new_[13684]_  & \new_[13679]_ ;
  assign \new_[13688]_  = ~A267 & ~A203;
  assign \new_[13692]_  = A299 & A298;
  assign \new_[13693]_  = ~A269 & \new_[13692]_ ;
  assign \new_[13694]_  = \new_[13693]_  & \new_[13688]_ ;
  assign \new_[13697]_  = A166 & A167;
  assign \new_[13701]_  = A201 & ~A200;
  assign \new_[13702]_  = A199 & \new_[13701]_ ;
  assign \new_[13703]_  = \new_[13702]_  & \new_[13697]_ ;
  assign \new_[13706]_  = ~A267 & ~A203;
  assign \new_[13710]_  = ~A299 & ~A298;
  assign \new_[13711]_  = ~A269 & \new_[13710]_ ;
  assign \new_[13712]_  = \new_[13711]_  & \new_[13706]_ ;
  assign \new_[13715]_  = A166 & A167;
  assign \new_[13719]_  = A201 & ~A200;
  assign \new_[13720]_  = A199 & \new_[13719]_ ;
  assign \new_[13721]_  = \new_[13720]_  & \new_[13715]_ ;
  assign \new_[13724]_  = A265 & ~A203;
  assign \new_[13728]_  = A301 & ~A300;
  assign \new_[13729]_  = A266 & \new_[13728]_ ;
  assign \new_[13730]_  = \new_[13729]_  & \new_[13724]_ ;
  assign \new_[13733]_  = A166 & A167;
  assign \new_[13737]_  = A201 & ~A200;
  assign \new_[13738]_  = A199 & \new_[13737]_ ;
  assign \new_[13739]_  = \new_[13738]_  & \new_[13733]_ ;
  assign \new_[13742]_  = A265 & ~A203;
  assign \new_[13746]_  = ~A302 & ~A300;
  assign \new_[13747]_  = A266 & \new_[13746]_ ;
  assign \new_[13748]_  = \new_[13747]_  & \new_[13742]_ ;
  assign \new_[13751]_  = A166 & A167;
  assign \new_[13755]_  = A201 & ~A200;
  assign \new_[13756]_  = A199 & \new_[13755]_ ;
  assign \new_[13757]_  = \new_[13756]_  & \new_[13751]_ ;
  assign \new_[13760]_  = A265 & ~A203;
  assign \new_[13764]_  = A299 & A298;
  assign \new_[13765]_  = A266 & \new_[13764]_ ;
  assign \new_[13766]_  = \new_[13765]_  & \new_[13760]_ ;
  assign \new_[13769]_  = A166 & A167;
  assign \new_[13773]_  = A201 & ~A200;
  assign \new_[13774]_  = A199 & \new_[13773]_ ;
  assign \new_[13775]_  = \new_[13774]_  & \new_[13769]_ ;
  assign \new_[13778]_  = A265 & ~A203;
  assign \new_[13782]_  = ~A299 & ~A298;
  assign \new_[13783]_  = A266 & \new_[13782]_ ;
  assign \new_[13784]_  = \new_[13783]_  & \new_[13778]_ ;
  assign \new_[13787]_  = A166 & A167;
  assign \new_[13791]_  = A201 & ~A200;
  assign \new_[13792]_  = A199 & \new_[13791]_ ;
  assign \new_[13793]_  = \new_[13792]_  & \new_[13787]_ ;
  assign \new_[13796]_  = ~A265 & ~A203;
  assign \new_[13800]_  = A301 & ~A300;
  assign \new_[13801]_  = ~A266 & \new_[13800]_ ;
  assign \new_[13802]_  = \new_[13801]_  & \new_[13796]_ ;
  assign \new_[13805]_  = A166 & A167;
  assign \new_[13809]_  = A201 & ~A200;
  assign \new_[13810]_  = A199 & \new_[13809]_ ;
  assign \new_[13811]_  = \new_[13810]_  & \new_[13805]_ ;
  assign \new_[13814]_  = ~A265 & ~A203;
  assign \new_[13818]_  = ~A302 & ~A300;
  assign \new_[13819]_  = ~A266 & \new_[13818]_ ;
  assign \new_[13820]_  = \new_[13819]_  & \new_[13814]_ ;
  assign \new_[13823]_  = A166 & A167;
  assign \new_[13827]_  = A201 & ~A200;
  assign \new_[13828]_  = A199 & \new_[13827]_ ;
  assign \new_[13829]_  = \new_[13828]_  & \new_[13823]_ ;
  assign \new_[13832]_  = ~A265 & ~A203;
  assign \new_[13836]_  = A299 & A298;
  assign \new_[13837]_  = ~A266 & \new_[13836]_ ;
  assign \new_[13838]_  = \new_[13837]_  & \new_[13832]_ ;
  assign \new_[13841]_  = A166 & A167;
  assign \new_[13845]_  = A201 & ~A200;
  assign \new_[13846]_  = A199 & \new_[13845]_ ;
  assign \new_[13847]_  = \new_[13846]_  & \new_[13841]_ ;
  assign \new_[13850]_  = ~A265 & ~A203;
  assign \new_[13854]_  = ~A299 & ~A298;
  assign \new_[13855]_  = ~A266 & \new_[13854]_ ;
  assign \new_[13856]_  = \new_[13855]_  & \new_[13850]_ ;
  assign \new_[13859]_  = ~A166 & ~A167;
  assign \new_[13863]_  = A201 & A200;
  assign \new_[13864]_  = ~A199 & \new_[13863]_ ;
  assign \new_[13865]_  = \new_[13864]_  & \new_[13859]_ ;
  assign \new_[13868]_  = ~A267 & A202;
  assign \new_[13872]_  = A301 & ~A300;
  assign \new_[13873]_  = A268 & \new_[13872]_ ;
  assign \new_[13874]_  = \new_[13873]_  & \new_[13868]_ ;
  assign \new_[13877]_  = ~A166 & ~A167;
  assign \new_[13881]_  = A201 & A200;
  assign \new_[13882]_  = ~A199 & \new_[13881]_ ;
  assign \new_[13883]_  = \new_[13882]_  & \new_[13877]_ ;
  assign \new_[13886]_  = ~A267 & A202;
  assign \new_[13890]_  = ~A302 & ~A300;
  assign \new_[13891]_  = A268 & \new_[13890]_ ;
  assign \new_[13892]_  = \new_[13891]_  & \new_[13886]_ ;
  assign \new_[13895]_  = ~A166 & ~A167;
  assign \new_[13899]_  = A201 & A200;
  assign \new_[13900]_  = ~A199 & \new_[13899]_ ;
  assign \new_[13901]_  = \new_[13900]_  & \new_[13895]_ ;
  assign \new_[13904]_  = ~A267 & A202;
  assign \new_[13908]_  = A299 & A298;
  assign \new_[13909]_  = A268 & \new_[13908]_ ;
  assign \new_[13910]_  = \new_[13909]_  & \new_[13904]_ ;
  assign \new_[13913]_  = ~A166 & ~A167;
  assign \new_[13917]_  = A201 & A200;
  assign \new_[13918]_  = ~A199 & \new_[13917]_ ;
  assign \new_[13919]_  = \new_[13918]_  & \new_[13913]_ ;
  assign \new_[13922]_  = ~A267 & A202;
  assign \new_[13926]_  = ~A299 & ~A298;
  assign \new_[13927]_  = A268 & \new_[13926]_ ;
  assign \new_[13928]_  = \new_[13927]_  & \new_[13922]_ ;
  assign \new_[13931]_  = ~A166 & ~A167;
  assign \new_[13935]_  = A201 & A200;
  assign \new_[13936]_  = ~A199 & \new_[13935]_ ;
  assign \new_[13937]_  = \new_[13936]_  & \new_[13931]_ ;
  assign \new_[13940]_  = ~A267 & A202;
  assign \new_[13944]_  = A301 & ~A300;
  assign \new_[13945]_  = ~A269 & \new_[13944]_ ;
  assign \new_[13946]_  = \new_[13945]_  & \new_[13940]_ ;
  assign \new_[13949]_  = ~A166 & ~A167;
  assign \new_[13953]_  = A201 & A200;
  assign \new_[13954]_  = ~A199 & \new_[13953]_ ;
  assign \new_[13955]_  = \new_[13954]_  & \new_[13949]_ ;
  assign \new_[13958]_  = ~A267 & A202;
  assign \new_[13962]_  = ~A302 & ~A300;
  assign \new_[13963]_  = ~A269 & \new_[13962]_ ;
  assign \new_[13964]_  = \new_[13963]_  & \new_[13958]_ ;
  assign \new_[13967]_  = ~A166 & ~A167;
  assign \new_[13971]_  = A201 & A200;
  assign \new_[13972]_  = ~A199 & \new_[13971]_ ;
  assign \new_[13973]_  = \new_[13972]_  & \new_[13967]_ ;
  assign \new_[13976]_  = ~A267 & A202;
  assign \new_[13980]_  = A299 & A298;
  assign \new_[13981]_  = ~A269 & \new_[13980]_ ;
  assign \new_[13982]_  = \new_[13981]_  & \new_[13976]_ ;
  assign \new_[13985]_  = ~A166 & ~A167;
  assign \new_[13989]_  = A201 & A200;
  assign \new_[13990]_  = ~A199 & \new_[13989]_ ;
  assign \new_[13991]_  = \new_[13990]_  & \new_[13985]_ ;
  assign \new_[13994]_  = ~A267 & A202;
  assign \new_[13998]_  = ~A299 & ~A298;
  assign \new_[13999]_  = ~A269 & \new_[13998]_ ;
  assign \new_[14000]_  = \new_[13999]_  & \new_[13994]_ ;
  assign \new_[14003]_  = ~A166 & ~A167;
  assign \new_[14007]_  = A201 & A200;
  assign \new_[14008]_  = ~A199 & \new_[14007]_ ;
  assign \new_[14009]_  = \new_[14008]_  & \new_[14003]_ ;
  assign \new_[14012]_  = A265 & A202;
  assign \new_[14016]_  = A301 & ~A300;
  assign \new_[14017]_  = A266 & \new_[14016]_ ;
  assign \new_[14018]_  = \new_[14017]_  & \new_[14012]_ ;
  assign \new_[14021]_  = ~A166 & ~A167;
  assign \new_[14025]_  = A201 & A200;
  assign \new_[14026]_  = ~A199 & \new_[14025]_ ;
  assign \new_[14027]_  = \new_[14026]_  & \new_[14021]_ ;
  assign \new_[14030]_  = A265 & A202;
  assign \new_[14034]_  = ~A302 & ~A300;
  assign \new_[14035]_  = A266 & \new_[14034]_ ;
  assign \new_[14036]_  = \new_[14035]_  & \new_[14030]_ ;
  assign \new_[14039]_  = ~A166 & ~A167;
  assign \new_[14043]_  = A201 & A200;
  assign \new_[14044]_  = ~A199 & \new_[14043]_ ;
  assign \new_[14045]_  = \new_[14044]_  & \new_[14039]_ ;
  assign \new_[14048]_  = A265 & A202;
  assign \new_[14052]_  = A299 & A298;
  assign \new_[14053]_  = A266 & \new_[14052]_ ;
  assign \new_[14054]_  = \new_[14053]_  & \new_[14048]_ ;
  assign \new_[14057]_  = ~A166 & ~A167;
  assign \new_[14061]_  = A201 & A200;
  assign \new_[14062]_  = ~A199 & \new_[14061]_ ;
  assign \new_[14063]_  = \new_[14062]_  & \new_[14057]_ ;
  assign \new_[14066]_  = A265 & A202;
  assign \new_[14070]_  = ~A299 & ~A298;
  assign \new_[14071]_  = A266 & \new_[14070]_ ;
  assign \new_[14072]_  = \new_[14071]_  & \new_[14066]_ ;
  assign \new_[14075]_  = ~A166 & ~A167;
  assign \new_[14079]_  = A201 & A200;
  assign \new_[14080]_  = ~A199 & \new_[14079]_ ;
  assign \new_[14081]_  = \new_[14080]_  & \new_[14075]_ ;
  assign \new_[14084]_  = ~A265 & A202;
  assign \new_[14088]_  = A301 & ~A300;
  assign \new_[14089]_  = ~A266 & \new_[14088]_ ;
  assign \new_[14090]_  = \new_[14089]_  & \new_[14084]_ ;
  assign \new_[14093]_  = ~A166 & ~A167;
  assign \new_[14097]_  = A201 & A200;
  assign \new_[14098]_  = ~A199 & \new_[14097]_ ;
  assign \new_[14099]_  = \new_[14098]_  & \new_[14093]_ ;
  assign \new_[14102]_  = ~A265 & A202;
  assign \new_[14106]_  = ~A302 & ~A300;
  assign \new_[14107]_  = ~A266 & \new_[14106]_ ;
  assign \new_[14108]_  = \new_[14107]_  & \new_[14102]_ ;
  assign \new_[14111]_  = ~A166 & ~A167;
  assign \new_[14115]_  = A201 & A200;
  assign \new_[14116]_  = ~A199 & \new_[14115]_ ;
  assign \new_[14117]_  = \new_[14116]_  & \new_[14111]_ ;
  assign \new_[14120]_  = ~A265 & A202;
  assign \new_[14124]_  = A299 & A298;
  assign \new_[14125]_  = ~A266 & \new_[14124]_ ;
  assign \new_[14126]_  = \new_[14125]_  & \new_[14120]_ ;
  assign \new_[14129]_  = ~A166 & ~A167;
  assign \new_[14133]_  = A201 & A200;
  assign \new_[14134]_  = ~A199 & \new_[14133]_ ;
  assign \new_[14135]_  = \new_[14134]_  & \new_[14129]_ ;
  assign \new_[14138]_  = ~A265 & A202;
  assign \new_[14142]_  = ~A299 & ~A298;
  assign \new_[14143]_  = ~A266 & \new_[14142]_ ;
  assign \new_[14144]_  = \new_[14143]_  & \new_[14138]_ ;
  assign \new_[14147]_  = ~A166 & ~A167;
  assign \new_[14151]_  = A201 & A200;
  assign \new_[14152]_  = ~A199 & \new_[14151]_ ;
  assign \new_[14153]_  = \new_[14152]_  & \new_[14147]_ ;
  assign \new_[14156]_  = ~A267 & ~A203;
  assign \new_[14160]_  = A301 & ~A300;
  assign \new_[14161]_  = A268 & \new_[14160]_ ;
  assign \new_[14162]_  = \new_[14161]_  & \new_[14156]_ ;
  assign \new_[14165]_  = ~A166 & ~A167;
  assign \new_[14169]_  = A201 & A200;
  assign \new_[14170]_  = ~A199 & \new_[14169]_ ;
  assign \new_[14171]_  = \new_[14170]_  & \new_[14165]_ ;
  assign \new_[14174]_  = ~A267 & ~A203;
  assign \new_[14178]_  = ~A302 & ~A300;
  assign \new_[14179]_  = A268 & \new_[14178]_ ;
  assign \new_[14180]_  = \new_[14179]_  & \new_[14174]_ ;
  assign \new_[14183]_  = ~A166 & ~A167;
  assign \new_[14187]_  = A201 & A200;
  assign \new_[14188]_  = ~A199 & \new_[14187]_ ;
  assign \new_[14189]_  = \new_[14188]_  & \new_[14183]_ ;
  assign \new_[14192]_  = ~A267 & ~A203;
  assign \new_[14196]_  = A299 & A298;
  assign \new_[14197]_  = A268 & \new_[14196]_ ;
  assign \new_[14198]_  = \new_[14197]_  & \new_[14192]_ ;
  assign \new_[14201]_  = ~A166 & ~A167;
  assign \new_[14205]_  = A201 & A200;
  assign \new_[14206]_  = ~A199 & \new_[14205]_ ;
  assign \new_[14207]_  = \new_[14206]_  & \new_[14201]_ ;
  assign \new_[14210]_  = ~A267 & ~A203;
  assign \new_[14214]_  = ~A299 & ~A298;
  assign \new_[14215]_  = A268 & \new_[14214]_ ;
  assign \new_[14216]_  = \new_[14215]_  & \new_[14210]_ ;
  assign \new_[14219]_  = ~A166 & ~A167;
  assign \new_[14223]_  = A201 & A200;
  assign \new_[14224]_  = ~A199 & \new_[14223]_ ;
  assign \new_[14225]_  = \new_[14224]_  & \new_[14219]_ ;
  assign \new_[14228]_  = ~A267 & ~A203;
  assign \new_[14232]_  = A301 & ~A300;
  assign \new_[14233]_  = ~A269 & \new_[14232]_ ;
  assign \new_[14234]_  = \new_[14233]_  & \new_[14228]_ ;
  assign \new_[14237]_  = ~A166 & ~A167;
  assign \new_[14241]_  = A201 & A200;
  assign \new_[14242]_  = ~A199 & \new_[14241]_ ;
  assign \new_[14243]_  = \new_[14242]_  & \new_[14237]_ ;
  assign \new_[14246]_  = ~A267 & ~A203;
  assign \new_[14250]_  = ~A302 & ~A300;
  assign \new_[14251]_  = ~A269 & \new_[14250]_ ;
  assign \new_[14252]_  = \new_[14251]_  & \new_[14246]_ ;
  assign \new_[14255]_  = ~A166 & ~A167;
  assign \new_[14259]_  = A201 & A200;
  assign \new_[14260]_  = ~A199 & \new_[14259]_ ;
  assign \new_[14261]_  = \new_[14260]_  & \new_[14255]_ ;
  assign \new_[14264]_  = ~A267 & ~A203;
  assign \new_[14268]_  = A299 & A298;
  assign \new_[14269]_  = ~A269 & \new_[14268]_ ;
  assign \new_[14270]_  = \new_[14269]_  & \new_[14264]_ ;
  assign \new_[14273]_  = ~A166 & ~A167;
  assign \new_[14277]_  = A201 & A200;
  assign \new_[14278]_  = ~A199 & \new_[14277]_ ;
  assign \new_[14279]_  = \new_[14278]_  & \new_[14273]_ ;
  assign \new_[14282]_  = ~A267 & ~A203;
  assign \new_[14286]_  = ~A299 & ~A298;
  assign \new_[14287]_  = ~A269 & \new_[14286]_ ;
  assign \new_[14288]_  = \new_[14287]_  & \new_[14282]_ ;
  assign \new_[14291]_  = ~A166 & ~A167;
  assign \new_[14295]_  = A201 & A200;
  assign \new_[14296]_  = ~A199 & \new_[14295]_ ;
  assign \new_[14297]_  = \new_[14296]_  & \new_[14291]_ ;
  assign \new_[14300]_  = A265 & ~A203;
  assign \new_[14304]_  = A301 & ~A300;
  assign \new_[14305]_  = A266 & \new_[14304]_ ;
  assign \new_[14306]_  = \new_[14305]_  & \new_[14300]_ ;
  assign \new_[14309]_  = ~A166 & ~A167;
  assign \new_[14313]_  = A201 & A200;
  assign \new_[14314]_  = ~A199 & \new_[14313]_ ;
  assign \new_[14315]_  = \new_[14314]_  & \new_[14309]_ ;
  assign \new_[14318]_  = A265 & ~A203;
  assign \new_[14322]_  = ~A302 & ~A300;
  assign \new_[14323]_  = A266 & \new_[14322]_ ;
  assign \new_[14324]_  = \new_[14323]_  & \new_[14318]_ ;
  assign \new_[14327]_  = ~A166 & ~A167;
  assign \new_[14331]_  = A201 & A200;
  assign \new_[14332]_  = ~A199 & \new_[14331]_ ;
  assign \new_[14333]_  = \new_[14332]_  & \new_[14327]_ ;
  assign \new_[14336]_  = A265 & ~A203;
  assign \new_[14340]_  = A299 & A298;
  assign \new_[14341]_  = A266 & \new_[14340]_ ;
  assign \new_[14342]_  = \new_[14341]_  & \new_[14336]_ ;
  assign \new_[14345]_  = ~A166 & ~A167;
  assign \new_[14349]_  = A201 & A200;
  assign \new_[14350]_  = ~A199 & \new_[14349]_ ;
  assign \new_[14351]_  = \new_[14350]_  & \new_[14345]_ ;
  assign \new_[14354]_  = A265 & ~A203;
  assign \new_[14358]_  = ~A299 & ~A298;
  assign \new_[14359]_  = A266 & \new_[14358]_ ;
  assign \new_[14360]_  = \new_[14359]_  & \new_[14354]_ ;
  assign \new_[14363]_  = ~A166 & ~A167;
  assign \new_[14367]_  = A201 & A200;
  assign \new_[14368]_  = ~A199 & \new_[14367]_ ;
  assign \new_[14369]_  = \new_[14368]_  & \new_[14363]_ ;
  assign \new_[14372]_  = ~A265 & ~A203;
  assign \new_[14376]_  = A301 & ~A300;
  assign \new_[14377]_  = ~A266 & \new_[14376]_ ;
  assign \new_[14378]_  = \new_[14377]_  & \new_[14372]_ ;
  assign \new_[14381]_  = ~A166 & ~A167;
  assign \new_[14385]_  = A201 & A200;
  assign \new_[14386]_  = ~A199 & \new_[14385]_ ;
  assign \new_[14387]_  = \new_[14386]_  & \new_[14381]_ ;
  assign \new_[14390]_  = ~A265 & ~A203;
  assign \new_[14394]_  = ~A302 & ~A300;
  assign \new_[14395]_  = ~A266 & \new_[14394]_ ;
  assign \new_[14396]_  = \new_[14395]_  & \new_[14390]_ ;
  assign \new_[14399]_  = ~A166 & ~A167;
  assign \new_[14403]_  = A201 & A200;
  assign \new_[14404]_  = ~A199 & \new_[14403]_ ;
  assign \new_[14405]_  = \new_[14404]_  & \new_[14399]_ ;
  assign \new_[14408]_  = ~A265 & ~A203;
  assign \new_[14412]_  = A299 & A298;
  assign \new_[14413]_  = ~A266 & \new_[14412]_ ;
  assign \new_[14414]_  = \new_[14413]_  & \new_[14408]_ ;
  assign \new_[14417]_  = ~A166 & ~A167;
  assign \new_[14421]_  = A201 & A200;
  assign \new_[14422]_  = ~A199 & \new_[14421]_ ;
  assign \new_[14423]_  = \new_[14422]_  & \new_[14417]_ ;
  assign \new_[14426]_  = ~A265 & ~A203;
  assign \new_[14430]_  = ~A299 & ~A298;
  assign \new_[14431]_  = ~A266 & \new_[14430]_ ;
  assign \new_[14432]_  = \new_[14431]_  & \new_[14426]_ ;
  assign \new_[14435]_  = ~A166 & ~A167;
  assign \new_[14439]_  = A201 & ~A200;
  assign \new_[14440]_  = A199 & \new_[14439]_ ;
  assign \new_[14441]_  = \new_[14440]_  & \new_[14435]_ ;
  assign \new_[14444]_  = ~A267 & A202;
  assign \new_[14448]_  = A301 & ~A300;
  assign \new_[14449]_  = A268 & \new_[14448]_ ;
  assign \new_[14450]_  = \new_[14449]_  & \new_[14444]_ ;
  assign \new_[14453]_  = ~A166 & ~A167;
  assign \new_[14457]_  = A201 & ~A200;
  assign \new_[14458]_  = A199 & \new_[14457]_ ;
  assign \new_[14459]_  = \new_[14458]_  & \new_[14453]_ ;
  assign \new_[14462]_  = ~A267 & A202;
  assign \new_[14466]_  = ~A302 & ~A300;
  assign \new_[14467]_  = A268 & \new_[14466]_ ;
  assign \new_[14468]_  = \new_[14467]_  & \new_[14462]_ ;
  assign \new_[14471]_  = ~A166 & ~A167;
  assign \new_[14475]_  = A201 & ~A200;
  assign \new_[14476]_  = A199 & \new_[14475]_ ;
  assign \new_[14477]_  = \new_[14476]_  & \new_[14471]_ ;
  assign \new_[14480]_  = ~A267 & A202;
  assign \new_[14484]_  = A299 & A298;
  assign \new_[14485]_  = A268 & \new_[14484]_ ;
  assign \new_[14486]_  = \new_[14485]_  & \new_[14480]_ ;
  assign \new_[14489]_  = ~A166 & ~A167;
  assign \new_[14493]_  = A201 & ~A200;
  assign \new_[14494]_  = A199 & \new_[14493]_ ;
  assign \new_[14495]_  = \new_[14494]_  & \new_[14489]_ ;
  assign \new_[14498]_  = ~A267 & A202;
  assign \new_[14502]_  = ~A299 & ~A298;
  assign \new_[14503]_  = A268 & \new_[14502]_ ;
  assign \new_[14504]_  = \new_[14503]_  & \new_[14498]_ ;
  assign \new_[14507]_  = ~A166 & ~A167;
  assign \new_[14511]_  = A201 & ~A200;
  assign \new_[14512]_  = A199 & \new_[14511]_ ;
  assign \new_[14513]_  = \new_[14512]_  & \new_[14507]_ ;
  assign \new_[14516]_  = ~A267 & A202;
  assign \new_[14520]_  = A301 & ~A300;
  assign \new_[14521]_  = ~A269 & \new_[14520]_ ;
  assign \new_[14522]_  = \new_[14521]_  & \new_[14516]_ ;
  assign \new_[14525]_  = ~A166 & ~A167;
  assign \new_[14529]_  = A201 & ~A200;
  assign \new_[14530]_  = A199 & \new_[14529]_ ;
  assign \new_[14531]_  = \new_[14530]_  & \new_[14525]_ ;
  assign \new_[14534]_  = ~A267 & A202;
  assign \new_[14538]_  = ~A302 & ~A300;
  assign \new_[14539]_  = ~A269 & \new_[14538]_ ;
  assign \new_[14540]_  = \new_[14539]_  & \new_[14534]_ ;
  assign \new_[14543]_  = ~A166 & ~A167;
  assign \new_[14547]_  = A201 & ~A200;
  assign \new_[14548]_  = A199 & \new_[14547]_ ;
  assign \new_[14549]_  = \new_[14548]_  & \new_[14543]_ ;
  assign \new_[14552]_  = ~A267 & A202;
  assign \new_[14556]_  = A299 & A298;
  assign \new_[14557]_  = ~A269 & \new_[14556]_ ;
  assign \new_[14558]_  = \new_[14557]_  & \new_[14552]_ ;
  assign \new_[14561]_  = ~A166 & ~A167;
  assign \new_[14565]_  = A201 & ~A200;
  assign \new_[14566]_  = A199 & \new_[14565]_ ;
  assign \new_[14567]_  = \new_[14566]_  & \new_[14561]_ ;
  assign \new_[14570]_  = ~A267 & A202;
  assign \new_[14574]_  = ~A299 & ~A298;
  assign \new_[14575]_  = ~A269 & \new_[14574]_ ;
  assign \new_[14576]_  = \new_[14575]_  & \new_[14570]_ ;
  assign \new_[14579]_  = ~A166 & ~A167;
  assign \new_[14583]_  = A201 & ~A200;
  assign \new_[14584]_  = A199 & \new_[14583]_ ;
  assign \new_[14585]_  = \new_[14584]_  & \new_[14579]_ ;
  assign \new_[14588]_  = A265 & A202;
  assign \new_[14592]_  = A301 & ~A300;
  assign \new_[14593]_  = A266 & \new_[14592]_ ;
  assign \new_[14594]_  = \new_[14593]_  & \new_[14588]_ ;
  assign \new_[14597]_  = ~A166 & ~A167;
  assign \new_[14601]_  = A201 & ~A200;
  assign \new_[14602]_  = A199 & \new_[14601]_ ;
  assign \new_[14603]_  = \new_[14602]_  & \new_[14597]_ ;
  assign \new_[14606]_  = A265 & A202;
  assign \new_[14610]_  = ~A302 & ~A300;
  assign \new_[14611]_  = A266 & \new_[14610]_ ;
  assign \new_[14612]_  = \new_[14611]_  & \new_[14606]_ ;
  assign \new_[14615]_  = ~A166 & ~A167;
  assign \new_[14619]_  = A201 & ~A200;
  assign \new_[14620]_  = A199 & \new_[14619]_ ;
  assign \new_[14621]_  = \new_[14620]_  & \new_[14615]_ ;
  assign \new_[14624]_  = A265 & A202;
  assign \new_[14628]_  = A299 & A298;
  assign \new_[14629]_  = A266 & \new_[14628]_ ;
  assign \new_[14630]_  = \new_[14629]_  & \new_[14624]_ ;
  assign \new_[14633]_  = ~A166 & ~A167;
  assign \new_[14637]_  = A201 & ~A200;
  assign \new_[14638]_  = A199 & \new_[14637]_ ;
  assign \new_[14639]_  = \new_[14638]_  & \new_[14633]_ ;
  assign \new_[14642]_  = A265 & A202;
  assign \new_[14646]_  = ~A299 & ~A298;
  assign \new_[14647]_  = A266 & \new_[14646]_ ;
  assign \new_[14648]_  = \new_[14647]_  & \new_[14642]_ ;
  assign \new_[14651]_  = ~A166 & ~A167;
  assign \new_[14655]_  = A201 & ~A200;
  assign \new_[14656]_  = A199 & \new_[14655]_ ;
  assign \new_[14657]_  = \new_[14656]_  & \new_[14651]_ ;
  assign \new_[14660]_  = ~A265 & A202;
  assign \new_[14664]_  = A301 & ~A300;
  assign \new_[14665]_  = ~A266 & \new_[14664]_ ;
  assign \new_[14666]_  = \new_[14665]_  & \new_[14660]_ ;
  assign \new_[14669]_  = ~A166 & ~A167;
  assign \new_[14673]_  = A201 & ~A200;
  assign \new_[14674]_  = A199 & \new_[14673]_ ;
  assign \new_[14675]_  = \new_[14674]_  & \new_[14669]_ ;
  assign \new_[14678]_  = ~A265 & A202;
  assign \new_[14682]_  = ~A302 & ~A300;
  assign \new_[14683]_  = ~A266 & \new_[14682]_ ;
  assign \new_[14684]_  = \new_[14683]_  & \new_[14678]_ ;
  assign \new_[14687]_  = ~A166 & ~A167;
  assign \new_[14691]_  = A201 & ~A200;
  assign \new_[14692]_  = A199 & \new_[14691]_ ;
  assign \new_[14693]_  = \new_[14692]_  & \new_[14687]_ ;
  assign \new_[14696]_  = ~A265 & A202;
  assign \new_[14700]_  = A299 & A298;
  assign \new_[14701]_  = ~A266 & \new_[14700]_ ;
  assign \new_[14702]_  = \new_[14701]_  & \new_[14696]_ ;
  assign \new_[14705]_  = ~A166 & ~A167;
  assign \new_[14709]_  = A201 & ~A200;
  assign \new_[14710]_  = A199 & \new_[14709]_ ;
  assign \new_[14711]_  = \new_[14710]_  & \new_[14705]_ ;
  assign \new_[14714]_  = ~A265 & A202;
  assign \new_[14718]_  = ~A299 & ~A298;
  assign \new_[14719]_  = ~A266 & \new_[14718]_ ;
  assign \new_[14720]_  = \new_[14719]_  & \new_[14714]_ ;
  assign \new_[14723]_  = ~A166 & ~A167;
  assign \new_[14727]_  = A201 & ~A200;
  assign \new_[14728]_  = A199 & \new_[14727]_ ;
  assign \new_[14729]_  = \new_[14728]_  & \new_[14723]_ ;
  assign \new_[14732]_  = ~A267 & ~A203;
  assign \new_[14736]_  = A301 & ~A300;
  assign \new_[14737]_  = A268 & \new_[14736]_ ;
  assign \new_[14738]_  = \new_[14737]_  & \new_[14732]_ ;
  assign \new_[14741]_  = ~A166 & ~A167;
  assign \new_[14745]_  = A201 & ~A200;
  assign \new_[14746]_  = A199 & \new_[14745]_ ;
  assign \new_[14747]_  = \new_[14746]_  & \new_[14741]_ ;
  assign \new_[14750]_  = ~A267 & ~A203;
  assign \new_[14754]_  = ~A302 & ~A300;
  assign \new_[14755]_  = A268 & \new_[14754]_ ;
  assign \new_[14756]_  = \new_[14755]_  & \new_[14750]_ ;
  assign \new_[14759]_  = ~A166 & ~A167;
  assign \new_[14763]_  = A201 & ~A200;
  assign \new_[14764]_  = A199 & \new_[14763]_ ;
  assign \new_[14765]_  = \new_[14764]_  & \new_[14759]_ ;
  assign \new_[14768]_  = ~A267 & ~A203;
  assign \new_[14772]_  = A299 & A298;
  assign \new_[14773]_  = A268 & \new_[14772]_ ;
  assign \new_[14774]_  = \new_[14773]_  & \new_[14768]_ ;
  assign \new_[14777]_  = ~A166 & ~A167;
  assign \new_[14781]_  = A201 & ~A200;
  assign \new_[14782]_  = A199 & \new_[14781]_ ;
  assign \new_[14783]_  = \new_[14782]_  & \new_[14777]_ ;
  assign \new_[14786]_  = ~A267 & ~A203;
  assign \new_[14790]_  = ~A299 & ~A298;
  assign \new_[14791]_  = A268 & \new_[14790]_ ;
  assign \new_[14792]_  = \new_[14791]_  & \new_[14786]_ ;
  assign \new_[14795]_  = ~A166 & ~A167;
  assign \new_[14799]_  = A201 & ~A200;
  assign \new_[14800]_  = A199 & \new_[14799]_ ;
  assign \new_[14801]_  = \new_[14800]_  & \new_[14795]_ ;
  assign \new_[14804]_  = ~A267 & ~A203;
  assign \new_[14808]_  = A301 & ~A300;
  assign \new_[14809]_  = ~A269 & \new_[14808]_ ;
  assign \new_[14810]_  = \new_[14809]_  & \new_[14804]_ ;
  assign \new_[14813]_  = ~A166 & ~A167;
  assign \new_[14817]_  = A201 & ~A200;
  assign \new_[14818]_  = A199 & \new_[14817]_ ;
  assign \new_[14819]_  = \new_[14818]_  & \new_[14813]_ ;
  assign \new_[14822]_  = ~A267 & ~A203;
  assign \new_[14826]_  = ~A302 & ~A300;
  assign \new_[14827]_  = ~A269 & \new_[14826]_ ;
  assign \new_[14828]_  = \new_[14827]_  & \new_[14822]_ ;
  assign \new_[14831]_  = ~A166 & ~A167;
  assign \new_[14835]_  = A201 & ~A200;
  assign \new_[14836]_  = A199 & \new_[14835]_ ;
  assign \new_[14837]_  = \new_[14836]_  & \new_[14831]_ ;
  assign \new_[14840]_  = ~A267 & ~A203;
  assign \new_[14844]_  = A299 & A298;
  assign \new_[14845]_  = ~A269 & \new_[14844]_ ;
  assign \new_[14846]_  = \new_[14845]_  & \new_[14840]_ ;
  assign \new_[14849]_  = ~A166 & ~A167;
  assign \new_[14853]_  = A201 & ~A200;
  assign \new_[14854]_  = A199 & \new_[14853]_ ;
  assign \new_[14855]_  = \new_[14854]_  & \new_[14849]_ ;
  assign \new_[14858]_  = ~A267 & ~A203;
  assign \new_[14862]_  = ~A299 & ~A298;
  assign \new_[14863]_  = ~A269 & \new_[14862]_ ;
  assign \new_[14864]_  = \new_[14863]_  & \new_[14858]_ ;
  assign \new_[14867]_  = ~A166 & ~A167;
  assign \new_[14871]_  = A201 & ~A200;
  assign \new_[14872]_  = A199 & \new_[14871]_ ;
  assign \new_[14873]_  = \new_[14872]_  & \new_[14867]_ ;
  assign \new_[14876]_  = A265 & ~A203;
  assign \new_[14880]_  = A301 & ~A300;
  assign \new_[14881]_  = A266 & \new_[14880]_ ;
  assign \new_[14882]_  = \new_[14881]_  & \new_[14876]_ ;
  assign \new_[14885]_  = ~A166 & ~A167;
  assign \new_[14889]_  = A201 & ~A200;
  assign \new_[14890]_  = A199 & \new_[14889]_ ;
  assign \new_[14891]_  = \new_[14890]_  & \new_[14885]_ ;
  assign \new_[14894]_  = A265 & ~A203;
  assign \new_[14898]_  = ~A302 & ~A300;
  assign \new_[14899]_  = A266 & \new_[14898]_ ;
  assign \new_[14900]_  = \new_[14899]_  & \new_[14894]_ ;
  assign \new_[14903]_  = ~A166 & ~A167;
  assign \new_[14907]_  = A201 & ~A200;
  assign \new_[14908]_  = A199 & \new_[14907]_ ;
  assign \new_[14909]_  = \new_[14908]_  & \new_[14903]_ ;
  assign \new_[14912]_  = A265 & ~A203;
  assign \new_[14916]_  = A299 & A298;
  assign \new_[14917]_  = A266 & \new_[14916]_ ;
  assign \new_[14918]_  = \new_[14917]_  & \new_[14912]_ ;
  assign \new_[14921]_  = ~A166 & ~A167;
  assign \new_[14925]_  = A201 & ~A200;
  assign \new_[14926]_  = A199 & \new_[14925]_ ;
  assign \new_[14927]_  = \new_[14926]_  & \new_[14921]_ ;
  assign \new_[14930]_  = A265 & ~A203;
  assign \new_[14934]_  = ~A299 & ~A298;
  assign \new_[14935]_  = A266 & \new_[14934]_ ;
  assign \new_[14936]_  = \new_[14935]_  & \new_[14930]_ ;
  assign \new_[14939]_  = ~A166 & ~A167;
  assign \new_[14943]_  = A201 & ~A200;
  assign \new_[14944]_  = A199 & \new_[14943]_ ;
  assign \new_[14945]_  = \new_[14944]_  & \new_[14939]_ ;
  assign \new_[14948]_  = ~A265 & ~A203;
  assign \new_[14952]_  = A301 & ~A300;
  assign \new_[14953]_  = ~A266 & \new_[14952]_ ;
  assign \new_[14954]_  = \new_[14953]_  & \new_[14948]_ ;
  assign \new_[14957]_  = ~A166 & ~A167;
  assign \new_[14961]_  = A201 & ~A200;
  assign \new_[14962]_  = A199 & \new_[14961]_ ;
  assign \new_[14963]_  = \new_[14962]_  & \new_[14957]_ ;
  assign \new_[14966]_  = ~A265 & ~A203;
  assign \new_[14970]_  = ~A302 & ~A300;
  assign \new_[14971]_  = ~A266 & \new_[14970]_ ;
  assign \new_[14972]_  = \new_[14971]_  & \new_[14966]_ ;
  assign \new_[14975]_  = ~A166 & ~A167;
  assign \new_[14979]_  = A201 & ~A200;
  assign \new_[14980]_  = A199 & \new_[14979]_ ;
  assign \new_[14981]_  = \new_[14980]_  & \new_[14975]_ ;
  assign \new_[14984]_  = ~A265 & ~A203;
  assign \new_[14988]_  = A299 & A298;
  assign \new_[14989]_  = ~A266 & \new_[14988]_ ;
  assign \new_[14990]_  = \new_[14989]_  & \new_[14984]_ ;
  assign \new_[14993]_  = ~A166 & ~A167;
  assign \new_[14997]_  = A201 & ~A200;
  assign \new_[14998]_  = A199 & \new_[14997]_ ;
  assign \new_[14999]_  = \new_[14998]_  & \new_[14993]_ ;
  assign \new_[15002]_  = ~A265 & ~A203;
  assign \new_[15006]_  = ~A299 & ~A298;
  assign \new_[15007]_  = ~A266 & \new_[15006]_ ;
  assign \new_[15008]_  = \new_[15007]_  & \new_[15002]_ ;
  assign \new_[15011]_  = ~A232 & ~A168;
  assign \new_[15015]_  = A235 & A234;
  assign \new_[15016]_  = A233 & \new_[15015]_ ;
  assign \new_[15017]_  = \new_[15016]_  & \new_[15011]_ ;
  assign \new_[15020]_  = A266 & ~A265;
  assign \new_[15024]_  = A269 & ~A268;
  assign \new_[15025]_  = ~A267 & \new_[15024]_ ;
  assign \new_[15026]_  = \new_[15025]_  & \new_[15020]_ ;
  assign \new_[15029]_  = ~A232 & ~A168;
  assign \new_[15033]_  = A235 & A234;
  assign \new_[15034]_  = A233 & \new_[15033]_ ;
  assign \new_[15035]_  = \new_[15034]_  & \new_[15029]_ ;
  assign \new_[15038]_  = ~A266 & A265;
  assign \new_[15042]_  = A269 & ~A268;
  assign \new_[15043]_  = ~A267 & \new_[15042]_ ;
  assign \new_[15044]_  = \new_[15043]_  & \new_[15038]_ ;
  assign \new_[15047]_  = ~A232 & ~A168;
  assign \new_[15051]_  = ~A236 & A234;
  assign \new_[15052]_  = A233 & \new_[15051]_ ;
  assign \new_[15053]_  = \new_[15052]_  & \new_[15047]_ ;
  assign \new_[15056]_  = A266 & ~A265;
  assign \new_[15060]_  = A269 & ~A268;
  assign \new_[15061]_  = ~A267 & \new_[15060]_ ;
  assign \new_[15062]_  = \new_[15061]_  & \new_[15056]_ ;
  assign \new_[15065]_  = ~A232 & ~A168;
  assign \new_[15069]_  = ~A236 & A234;
  assign \new_[15070]_  = A233 & \new_[15069]_ ;
  assign \new_[15071]_  = \new_[15070]_  & \new_[15065]_ ;
  assign \new_[15074]_  = ~A266 & A265;
  assign \new_[15078]_  = A269 & ~A268;
  assign \new_[15079]_  = ~A267 & \new_[15078]_ ;
  assign \new_[15080]_  = \new_[15079]_  & \new_[15074]_ ;
  assign \new_[15083]_  = A232 & ~A168;
  assign \new_[15087]_  = A235 & A234;
  assign \new_[15088]_  = ~A233 & \new_[15087]_ ;
  assign \new_[15089]_  = \new_[15088]_  & \new_[15083]_ ;
  assign \new_[15092]_  = A266 & ~A265;
  assign \new_[15096]_  = A269 & ~A268;
  assign \new_[15097]_  = ~A267 & \new_[15096]_ ;
  assign \new_[15098]_  = \new_[15097]_  & \new_[15092]_ ;
  assign \new_[15101]_  = A232 & ~A168;
  assign \new_[15105]_  = A235 & A234;
  assign \new_[15106]_  = ~A233 & \new_[15105]_ ;
  assign \new_[15107]_  = \new_[15106]_  & \new_[15101]_ ;
  assign \new_[15110]_  = ~A266 & A265;
  assign \new_[15114]_  = A269 & ~A268;
  assign \new_[15115]_  = ~A267 & \new_[15114]_ ;
  assign \new_[15116]_  = \new_[15115]_  & \new_[15110]_ ;
  assign \new_[15119]_  = A232 & ~A168;
  assign \new_[15123]_  = ~A236 & A234;
  assign \new_[15124]_  = ~A233 & \new_[15123]_ ;
  assign \new_[15125]_  = \new_[15124]_  & \new_[15119]_ ;
  assign \new_[15128]_  = A266 & ~A265;
  assign \new_[15132]_  = A269 & ~A268;
  assign \new_[15133]_  = ~A267 & \new_[15132]_ ;
  assign \new_[15134]_  = \new_[15133]_  & \new_[15128]_ ;
  assign \new_[15137]_  = A232 & ~A168;
  assign \new_[15141]_  = ~A236 & A234;
  assign \new_[15142]_  = ~A233 & \new_[15141]_ ;
  assign \new_[15143]_  = \new_[15142]_  & \new_[15137]_ ;
  assign \new_[15146]_  = ~A266 & A265;
  assign \new_[15150]_  = A269 & ~A268;
  assign \new_[15151]_  = ~A267 & \new_[15150]_ ;
  assign \new_[15152]_  = \new_[15151]_  & \new_[15146]_ ;
  assign \new_[15155]_  = ~A168 & A170;
  assign \new_[15159]_  = A201 & A200;
  assign \new_[15160]_  = ~A199 & \new_[15159]_ ;
  assign \new_[15161]_  = \new_[15160]_  & \new_[15155]_ ;
  assign \new_[15164]_  = ~A267 & A202;
  assign \new_[15168]_  = A301 & ~A300;
  assign \new_[15169]_  = A268 & \new_[15168]_ ;
  assign \new_[15170]_  = \new_[15169]_  & \new_[15164]_ ;
  assign \new_[15173]_  = ~A168 & A170;
  assign \new_[15177]_  = A201 & A200;
  assign \new_[15178]_  = ~A199 & \new_[15177]_ ;
  assign \new_[15179]_  = \new_[15178]_  & \new_[15173]_ ;
  assign \new_[15182]_  = ~A267 & A202;
  assign \new_[15186]_  = ~A302 & ~A300;
  assign \new_[15187]_  = A268 & \new_[15186]_ ;
  assign \new_[15188]_  = \new_[15187]_  & \new_[15182]_ ;
  assign \new_[15191]_  = ~A168 & A170;
  assign \new_[15195]_  = A201 & A200;
  assign \new_[15196]_  = ~A199 & \new_[15195]_ ;
  assign \new_[15197]_  = \new_[15196]_  & \new_[15191]_ ;
  assign \new_[15200]_  = ~A267 & A202;
  assign \new_[15204]_  = A299 & A298;
  assign \new_[15205]_  = A268 & \new_[15204]_ ;
  assign \new_[15206]_  = \new_[15205]_  & \new_[15200]_ ;
  assign \new_[15209]_  = ~A168 & A170;
  assign \new_[15213]_  = A201 & A200;
  assign \new_[15214]_  = ~A199 & \new_[15213]_ ;
  assign \new_[15215]_  = \new_[15214]_  & \new_[15209]_ ;
  assign \new_[15218]_  = ~A267 & A202;
  assign \new_[15222]_  = ~A299 & ~A298;
  assign \new_[15223]_  = A268 & \new_[15222]_ ;
  assign \new_[15224]_  = \new_[15223]_  & \new_[15218]_ ;
  assign \new_[15227]_  = ~A168 & A170;
  assign \new_[15231]_  = A201 & A200;
  assign \new_[15232]_  = ~A199 & \new_[15231]_ ;
  assign \new_[15233]_  = \new_[15232]_  & \new_[15227]_ ;
  assign \new_[15236]_  = ~A267 & A202;
  assign \new_[15240]_  = A301 & ~A300;
  assign \new_[15241]_  = ~A269 & \new_[15240]_ ;
  assign \new_[15242]_  = \new_[15241]_  & \new_[15236]_ ;
  assign \new_[15245]_  = ~A168 & A170;
  assign \new_[15249]_  = A201 & A200;
  assign \new_[15250]_  = ~A199 & \new_[15249]_ ;
  assign \new_[15251]_  = \new_[15250]_  & \new_[15245]_ ;
  assign \new_[15254]_  = ~A267 & A202;
  assign \new_[15258]_  = ~A302 & ~A300;
  assign \new_[15259]_  = ~A269 & \new_[15258]_ ;
  assign \new_[15260]_  = \new_[15259]_  & \new_[15254]_ ;
  assign \new_[15263]_  = ~A168 & A170;
  assign \new_[15267]_  = A201 & A200;
  assign \new_[15268]_  = ~A199 & \new_[15267]_ ;
  assign \new_[15269]_  = \new_[15268]_  & \new_[15263]_ ;
  assign \new_[15272]_  = ~A267 & A202;
  assign \new_[15276]_  = A299 & A298;
  assign \new_[15277]_  = ~A269 & \new_[15276]_ ;
  assign \new_[15278]_  = \new_[15277]_  & \new_[15272]_ ;
  assign \new_[15281]_  = ~A168 & A170;
  assign \new_[15285]_  = A201 & A200;
  assign \new_[15286]_  = ~A199 & \new_[15285]_ ;
  assign \new_[15287]_  = \new_[15286]_  & \new_[15281]_ ;
  assign \new_[15290]_  = ~A267 & A202;
  assign \new_[15294]_  = ~A299 & ~A298;
  assign \new_[15295]_  = ~A269 & \new_[15294]_ ;
  assign \new_[15296]_  = \new_[15295]_  & \new_[15290]_ ;
  assign \new_[15299]_  = ~A168 & A170;
  assign \new_[15303]_  = A201 & A200;
  assign \new_[15304]_  = ~A199 & \new_[15303]_ ;
  assign \new_[15305]_  = \new_[15304]_  & \new_[15299]_ ;
  assign \new_[15308]_  = A265 & A202;
  assign \new_[15312]_  = A301 & ~A300;
  assign \new_[15313]_  = A266 & \new_[15312]_ ;
  assign \new_[15314]_  = \new_[15313]_  & \new_[15308]_ ;
  assign \new_[15317]_  = ~A168 & A170;
  assign \new_[15321]_  = A201 & A200;
  assign \new_[15322]_  = ~A199 & \new_[15321]_ ;
  assign \new_[15323]_  = \new_[15322]_  & \new_[15317]_ ;
  assign \new_[15326]_  = A265 & A202;
  assign \new_[15330]_  = ~A302 & ~A300;
  assign \new_[15331]_  = A266 & \new_[15330]_ ;
  assign \new_[15332]_  = \new_[15331]_  & \new_[15326]_ ;
  assign \new_[15335]_  = ~A168 & A170;
  assign \new_[15339]_  = A201 & A200;
  assign \new_[15340]_  = ~A199 & \new_[15339]_ ;
  assign \new_[15341]_  = \new_[15340]_  & \new_[15335]_ ;
  assign \new_[15344]_  = A265 & A202;
  assign \new_[15348]_  = A299 & A298;
  assign \new_[15349]_  = A266 & \new_[15348]_ ;
  assign \new_[15350]_  = \new_[15349]_  & \new_[15344]_ ;
  assign \new_[15353]_  = ~A168 & A170;
  assign \new_[15357]_  = A201 & A200;
  assign \new_[15358]_  = ~A199 & \new_[15357]_ ;
  assign \new_[15359]_  = \new_[15358]_  & \new_[15353]_ ;
  assign \new_[15362]_  = A265 & A202;
  assign \new_[15366]_  = ~A299 & ~A298;
  assign \new_[15367]_  = A266 & \new_[15366]_ ;
  assign \new_[15368]_  = \new_[15367]_  & \new_[15362]_ ;
  assign \new_[15371]_  = ~A168 & A170;
  assign \new_[15375]_  = A201 & A200;
  assign \new_[15376]_  = ~A199 & \new_[15375]_ ;
  assign \new_[15377]_  = \new_[15376]_  & \new_[15371]_ ;
  assign \new_[15380]_  = ~A265 & A202;
  assign \new_[15384]_  = A301 & ~A300;
  assign \new_[15385]_  = ~A266 & \new_[15384]_ ;
  assign \new_[15386]_  = \new_[15385]_  & \new_[15380]_ ;
  assign \new_[15389]_  = ~A168 & A170;
  assign \new_[15393]_  = A201 & A200;
  assign \new_[15394]_  = ~A199 & \new_[15393]_ ;
  assign \new_[15395]_  = \new_[15394]_  & \new_[15389]_ ;
  assign \new_[15398]_  = ~A265 & A202;
  assign \new_[15402]_  = ~A302 & ~A300;
  assign \new_[15403]_  = ~A266 & \new_[15402]_ ;
  assign \new_[15404]_  = \new_[15403]_  & \new_[15398]_ ;
  assign \new_[15407]_  = ~A168 & A170;
  assign \new_[15411]_  = A201 & A200;
  assign \new_[15412]_  = ~A199 & \new_[15411]_ ;
  assign \new_[15413]_  = \new_[15412]_  & \new_[15407]_ ;
  assign \new_[15416]_  = ~A265 & A202;
  assign \new_[15420]_  = A299 & A298;
  assign \new_[15421]_  = ~A266 & \new_[15420]_ ;
  assign \new_[15422]_  = \new_[15421]_  & \new_[15416]_ ;
  assign \new_[15425]_  = ~A168 & A170;
  assign \new_[15429]_  = A201 & A200;
  assign \new_[15430]_  = ~A199 & \new_[15429]_ ;
  assign \new_[15431]_  = \new_[15430]_  & \new_[15425]_ ;
  assign \new_[15434]_  = ~A265 & A202;
  assign \new_[15438]_  = ~A299 & ~A298;
  assign \new_[15439]_  = ~A266 & \new_[15438]_ ;
  assign \new_[15440]_  = \new_[15439]_  & \new_[15434]_ ;
  assign \new_[15443]_  = ~A168 & A170;
  assign \new_[15447]_  = A201 & A200;
  assign \new_[15448]_  = ~A199 & \new_[15447]_ ;
  assign \new_[15449]_  = \new_[15448]_  & \new_[15443]_ ;
  assign \new_[15452]_  = ~A267 & ~A203;
  assign \new_[15456]_  = A301 & ~A300;
  assign \new_[15457]_  = A268 & \new_[15456]_ ;
  assign \new_[15458]_  = \new_[15457]_  & \new_[15452]_ ;
  assign \new_[15461]_  = ~A168 & A170;
  assign \new_[15465]_  = A201 & A200;
  assign \new_[15466]_  = ~A199 & \new_[15465]_ ;
  assign \new_[15467]_  = \new_[15466]_  & \new_[15461]_ ;
  assign \new_[15470]_  = ~A267 & ~A203;
  assign \new_[15474]_  = ~A302 & ~A300;
  assign \new_[15475]_  = A268 & \new_[15474]_ ;
  assign \new_[15476]_  = \new_[15475]_  & \new_[15470]_ ;
  assign \new_[15479]_  = ~A168 & A170;
  assign \new_[15483]_  = A201 & A200;
  assign \new_[15484]_  = ~A199 & \new_[15483]_ ;
  assign \new_[15485]_  = \new_[15484]_  & \new_[15479]_ ;
  assign \new_[15488]_  = ~A267 & ~A203;
  assign \new_[15492]_  = A299 & A298;
  assign \new_[15493]_  = A268 & \new_[15492]_ ;
  assign \new_[15494]_  = \new_[15493]_  & \new_[15488]_ ;
  assign \new_[15497]_  = ~A168 & A170;
  assign \new_[15501]_  = A201 & A200;
  assign \new_[15502]_  = ~A199 & \new_[15501]_ ;
  assign \new_[15503]_  = \new_[15502]_  & \new_[15497]_ ;
  assign \new_[15506]_  = ~A267 & ~A203;
  assign \new_[15510]_  = ~A299 & ~A298;
  assign \new_[15511]_  = A268 & \new_[15510]_ ;
  assign \new_[15512]_  = \new_[15511]_  & \new_[15506]_ ;
  assign \new_[15515]_  = ~A168 & A170;
  assign \new_[15519]_  = A201 & A200;
  assign \new_[15520]_  = ~A199 & \new_[15519]_ ;
  assign \new_[15521]_  = \new_[15520]_  & \new_[15515]_ ;
  assign \new_[15524]_  = ~A267 & ~A203;
  assign \new_[15528]_  = A301 & ~A300;
  assign \new_[15529]_  = ~A269 & \new_[15528]_ ;
  assign \new_[15530]_  = \new_[15529]_  & \new_[15524]_ ;
  assign \new_[15533]_  = ~A168 & A170;
  assign \new_[15537]_  = A201 & A200;
  assign \new_[15538]_  = ~A199 & \new_[15537]_ ;
  assign \new_[15539]_  = \new_[15538]_  & \new_[15533]_ ;
  assign \new_[15542]_  = ~A267 & ~A203;
  assign \new_[15546]_  = ~A302 & ~A300;
  assign \new_[15547]_  = ~A269 & \new_[15546]_ ;
  assign \new_[15548]_  = \new_[15547]_  & \new_[15542]_ ;
  assign \new_[15551]_  = ~A168 & A170;
  assign \new_[15555]_  = A201 & A200;
  assign \new_[15556]_  = ~A199 & \new_[15555]_ ;
  assign \new_[15557]_  = \new_[15556]_  & \new_[15551]_ ;
  assign \new_[15560]_  = ~A267 & ~A203;
  assign \new_[15564]_  = A299 & A298;
  assign \new_[15565]_  = ~A269 & \new_[15564]_ ;
  assign \new_[15566]_  = \new_[15565]_  & \new_[15560]_ ;
  assign \new_[15569]_  = ~A168 & A170;
  assign \new_[15573]_  = A201 & A200;
  assign \new_[15574]_  = ~A199 & \new_[15573]_ ;
  assign \new_[15575]_  = \new_[15574]_  & \new_[15569]_ ;
  assign \new_[15578]_  = ~A267 & ~A203;
  assign \new_[15582]_  = ~A299 & ~A298;
  assign \new_[15583]_  = ~A269 & \new_[15582]_ ;
  assign \new_[15584]_  = \new_[15583]_  & \new_[15578]_ ;
  assign \new_[15587]_  = ~A168 & A170;
  assign \new_[15591]_  = A201 & A200;
  assign \new_[15592]_  = ~A199 & \new_[15591]_ ;
  assign \new_[15593]_  = \new_[15592]_  & \new_[15587]_ ;
  assign \new_[15596]_  = A265 & ~A203;
  assign \new_[15600]_  = A301 & ~A300;
  assign \new_[15601]_  = A266 & \new_[15600]_ ;
  assign \new_[15602]_  = \new_[15601]_  & \new_[15596]_ ;
  assign \new_[15605]_  = ~A168 & A170;
  assign \new_[15609]_  = A201 & A200;
  assign \new_[15610]_  = ~A199 & \new_[15609]_ ;
  assign \new_[15611]_  = \new_[15610]_  & \new_[15605]_ ;
  assign \new_[15614]_  = A265 & ~A203;
  assign \new_[15618]_  = ~A302 & ~A300;
  assign \new_[15619]_  = A266 & \new_[15618]_ ;
  assign \new_[15620]_  = \new_[15619]_  & \new_[15614]_ ;
  assign \new_[15623]_  = ~A168 & A170;
  assign \new_[15627]_  = A201 & A200;
  assign \new_[15628]_  = ~A199 & \new_[15627]_ ;
  assign \new_[15629]_  = \new_[15628]_  & \new_[15623]_ ;
  assign \new_[15632]_  = A265 & ~A203;
  assign \new_[15636]_  = A299 & A298;
  assign \new_[15637]_  = A266 & \new_[15636]_ ;
  assign \new_[15638]_  = \new_[15637]_  & \new_[15632]_ ;
  assign \new_[15641]_  = ~A168 & A170;
  assign \new_[15645]_  = A201 & A200;
  assign \new_[15646]_  = ~A199 & \new_[15645]_ ;
  assign \new_[15647]_  = \new_[15646]_  & \new_[15641]_ ;
  assign \new_[15650]_  = A265 & ~A203;
  assign \new_[15654]_  = ~A299 & ~A298;
  assign \new_[15655]_  = A266 & \new_[15654]_ ;
  assign \new_[15656]_  = \new_[15655]_  & \new_[15650]_ ;
  assign \new_[15659]_  = ~A168 & A170;
  assign \new_[15663]_  = A201 & A200;
  assign \new_[15664]_  = ~A199 & \new_[15663]_ ;
  assign \new_[15665]_  = \new_[15664]_  & \new_[15659]_ ;
  assign \new_[15668]_  = ~A265 & ~A203;
  assign \new_[15672]_  = A301 & ~A300;
  assign \new_[15673]_  = ~A266 & \new_[15672]_ ;
  assign \new_[15674]_  = \new_[15673]_  & \new_[15668]_ ;
  assign \new_[15677]_  = ~A168 & A170;
  assign \new_[15681]_  = A201 & A200;
  assign \new_[15682]_  = ~A199 & \new_[15681]_ ;
  assign \new_[15683]_  = \new_[15682]_  & \new_[15677]_ ;
  assign \new_[15686]_  = ~A265 & ~A203;
  assign \new_[15690]_  = ~A302 & ~A300;
  assign \new_[15691]_  = ~A266 & \new_[15690]_ ;
  assign \new_[15692]_  = \new_[15691]_  & \new_[15686]_ ;
  assign \new_[15695]_  = ~A168 & A170;
  assign \new_[15699]_  = A201 & A200;
  assign \new_[15700]_  = ~A199 & \new_[15699]_ ;
  assign \new_[15701]_  = \new_[15700]_  & \new_[15695]_ ;
  assign \new_[15704]_  = ~A265 & ~A203;
  assign \new_[15708]_  = A299 & A298;
  assign \new_[15709]_  = ~A266 & \new_[15708]_ ;
  assign \new_[15710]_  = \new_[15709]_  & \new_[15704]_ ;
  assign \new_[15713]_  = ~A168 & A170;
  assign \new_[15717]_  = A201 & A200;
  assign \new_[15718]_  = ~A199 & \new_[15717]_ ;
  assign \new_[15719]_  = \new_[15718]_  & \new_[15713]_ ;
  assign \new_[15722]_  = ~A265 & ~A203;
  assign \new_[15726]_  = ~A299 & ~A298;
  assign \new_[15727]_  = ~A266 & \new_[15726]_ ;
  assign \new_[15728]_  = \new_[15727]_  & \new_[15722]_ ;
  assign \new_[15731]_  = ~A168 & A170;
  assign \new_[15735]_  = A201 & ~A200;
  assign \new_[15736]_  = A199 & \new_[15735]_ ;
  assign \new_[15737]_  = \new_[15736]_  & \new_[15731]_ ;
  assign \new_[15740]_  = ~A267 & A202;
  assign \new_[15744]_  = A301 & ~A300;
  assign \new_[15745]_  = A268 & \new_[15744]_ ;
  assign \new_[15746]_  = \new_[15745]_  & \new_[15740]_ ;
  assign \new_[15749]_  = ~A168 & A170;
  assign \new_[15753]_  = A201 & ~A200;
  assign \new_[15754]_  = A199 & \new_[15753]_ ;
  assign \new_[15755]_  = \new_[15754]_  & \new_[15749]_ ;
  assign \new_[15758]_  = ~A267 & A202;
  assign \new_[15762]_  = ~A302 & ~A300;
  assign \new_[15763]_  = A268 & \new_[15762]_ ;
  assign \new_[15764]_  = \new_[15763]_  & \new_[15758]_ ;
  assign \new_[15767]_  = ~A168 & A170;
  assign \new_[15771]_  = A201 & ~A200;
  assign \new_[15772]_  = A199 & \new_[15771]_ ;
  assign \new_[15773]_  = \new_[15772]_  & \new_[15767]_ ;
  assign \new_[15776]_  = ~A267 & A202;
  assign \new_[15780]_  = A299 & A298;
  assign \new_[15781]_  = A268 & \new_[15780]_ ;
  assign \new_[15782]_  = \new_[15781]_  & \new_[15776]_ ;
  assign \new_[15785]_  = ~A168 & A170;
  assign \new_[15789]_  = A201 & ~A200;
  assign \new_[15790]_  = A199 & \new_[15789]_ ;
  assign \new_[15791]_  = \new_[15790]_  & \new_[15785]_ ;
  assign \new_[15794]_  = ~A267 & A202;
  assign \new_[15798]_  = ~A299 & ~A298;
  assign \new_[15799]_  = A268 & \new_[15798]_ ;
  assign \new_[15800]_  = \new_[15799]_  & \new_[15794]_ ;
  assign \new_[15803]_  = ~A168 & A170;
  assign \new_[15807]_  = A201 & ~A200;
  assign \new_[15808]_  = A199 & \new_[15807]_ ;
  assign \new_[15809]_  = \new_[15808]_  & \new_[15803]_ ;
  assign \new_[15812]_  = ~A267 & A202;
  assign \new_[15816]_  = A301 & ~A300;
  assign \new_[15817]_  = ~A269 & \new_[15816]_ ;
  assign \new_[15818]_  = \new_[15817]_  & \new_[15812]_ ;
  assign \new_[15821]_  = ~A168 & A170;
  assign \new_[15825]_  = A201 & ~A200;
  assign \new_[15826]_  = A199 & \new_[15825]_ ;
  assign \new_[15827]_  = \new_[15826]_  & \new_[15821]_ ;
  assign \new_[15830]_  = ~A267 & A202;
  assign \new_[15834]_  = ~A302 & ~A300;
  assign \new_[15835]_  = ~A269 & \new_[15834]_ ;
  assign \new_[15836]_  = \new_[15835]_  & \new_[15830]_ ;
  assign \new_[15839]_  = ~A168 & A170;
  assign \new_[15843]_  = A201 & ~A200;
  assign \new_[15844]_  = A199 & \new_[15843]_ ;
  assign \new_[15845]_  = \new_[15844]_  & \new_[15839]_ ;
  assign \new_[15848]_  = ~A267 & A202;
  assign \new_[15852]_  = A299 & A298;
  assign \new_[15853]_  = ~A269 & \new_[15852]_ ;
  assign \new_[15854]_  = \new_[15853]_  & \new_[15848]_ ;
  assign \new_[15857]_  = ~A168 & A170;
  assign \new_[15861]_  = A201 & ~A200;
  assign \new_[15862]_  = A199 & \new_[15861]_ ;
  assign \new_[15863]_  = \new_[15862]_  & \new_[15857]_ ;
  assign \new_[15866]_  = ~A267 & A202;
  assign \new_[15870]_  = ~A299 & ~A298;
  assign \new_[15871]_  = ~A269 & \new_[15870]_ ;
  assign \new_[15872]_  = \new_[15871]_  & \new_[15866]_ ;
  assign \new_[15875]_  = ~A168 & A170;
  assign \new_[15879]_  = A201 & ~A200;
  assign \new_[15880]_  = A199 & \new_[15879]_ ;
  assign \new_[15881]_  = \new_[15880]_  & \new_[15875]_ ;
  assign \new_[15884]_  = A265 & A202;
  assign \new_[15888]_  = A301 & ~A300;
  assign \new_[15889]_  = A266 & \new_[15888]_ ;
  assign \new_[15890]_  = \new_[15889]_  & \new_[15884]_ ;
  assign \new_[15893]_  = ~A168 & A170;
  assign \new_[15897]_  = A201 & ~A200;
  assign \new_[15898]_  = A199 & \new_[15897]_ ;
  assign \new_[15899]_  = \new_[15898]_  & \new_[15893]_ ;
  assign \new_[15902]_  = A265 & A202;
  assign \new_[15906]_  = ~A302 & ~A300;
  assign \new_[15907]_  = A266 & \new_[15906]_ ;
  assign \new_[15908]_  = \new_[15907]_  & \new_[15902]_ ;
  assign \new_[15911]_  = ~A168 & A170;
  assign \new_[15915]_  = A201 & ~A200;
  assign \new_[15916]_  = A199 & \new_[15915]_ ;
  assign \new_[15917]_  = \new_[15916]_  & \new_[15911]_ ;
  assign \new_[15920]_  = A265 & A202;
  assign \new_[15924]_  = A299 & A298;
  assign \new_[15925]_  = A266 & \new_[15924]_ ;
  assign \new_[15926]_  = \new_[15925]_  & \new_[15920]_ ;
  assign \new_[15929]_  = ~A168 & A170;
  assign \new_[15933]_  = A201 & ~A200;
  assign \new_[15934]_  = A199 & \new_[15933]_ ;
  assign \new_[15935]_  = \new_[15934]_  & \new_[15929]_ ;
  assign \new_[15938]_  = A265 & A202;
  assign \new_[15942]_  = ~A299 & ~A298;
  assign \new_[15943]_  = A266 & \new_[15942]_ ;
  assign \new_[15944]_  = \new_[15943]_  & \new_[15938]_ ;
  assign \new_[15947]_  = ~A168 & A170;
  assign \new_[15951]_  = A201 & ~A200;
  assign \new_[15952]_  = A199 & \new_[15951]_ ;
  assign \new_[15953]_  = \new_[15952]_  & \new_[15947]_ ;
  assign \new_[15956]_  = ~A265 & A202;
  assign \new_[15960]_  = A301 & ~A300;
  assign \new_[15961]_  = ~A266 & \new_[15960]_ ;
  assign \new_[15962]_  = \new_[15961]_  & \new_[15956]_ ;
  assign \new_[15965]_  = ~A168 & A170;
  assign \new_[15969]_  = A201 & ~A200;
  assign \new_[15970]_  = A199 & \new_[15969]_ ;
  assign \new_[15971]_  = \new_[15970]_  & \new_[15965]_ ;
  assign \new_[15974]_  = ~A265 & A202;
  assign \new_[15978]_  = ~A302 & ~A300;
  assign \new_[15979]_  = ~A266 & \new_[15978]_ ;
  assign \new_[15980]_  = \new_[15979]_  & \new_[15974]_ ;
  assign \new_[15983]_  = ~A168 & A170;
  assign \new_[15987]_  = A201 & ~A200;
  assign \new_[15988]_  = A199 & \new_[15987]_ ;
  assign \new_[15989]_  = \new_[15988]_  & \new_[15983]_ ;
  assign \new_[15992]_  = ~A265 & A202;
  assign \new_[15996]_  = A299 & A298;
  assign \new_[15997]_  = ~A266 & \new_[15996]_ ;
  assign \new_[15998]_  = \new_[15997]_  & \new_[15992]_ ;
  assign \new_[16001]_  = ~A168 & A170;
  assign \new_[16005]_  = A201 & ~A200;
  assign \new_[16006]_  = A199 & \new_[16005]_ ;
  assign \new_[16007]_  = \new_[16006]_  & \new_[16001]_ ;
  assign \new_[16010]_  = ~A265 & A202;
  assign \new_[16014]_  = ~A299 & ~A298;
  assign \new_[16015]_  = ~A266 & \new_[16014]_ ;
  assign \new_[16016]_  = \new_[16015]_  & \new_[16010]_ ;
  assign \new_[16019]_  = ~A168 & A170;
  assign \new_[16023]_  = A201 & ~A200;
  assign \new_[16024]_  = A199 & \new_[16023]_ ;
  assign \new_[16025]_  = \new_[16024]_  & \new_[16019]_ ;
  assign \new_[16028]_  = ~A267 & ~A203;
  assign \new_[16032]_  = A301 & ~A300;
  assign \new_[16033]_  = A268 & \new_[16032]_ ;
  assign \new_[16034]_  = \new_[16033]_  & \new_[16028]_ ;
  assign \new_[16037]_  = ~A168 & A170;
  assign \new_[16041]_  = A201 & ~A200;
  assign \new_[16042]_  = A199 & \new_[16041]_ ;
  assign \new_[16043]_  = \new_[16042]_  & \new_[16037]_ ;
  assign \new_[16046]_  = ~A267 & ~A203;
  assign \new_[16050]_  = ~A302 & ~A300;
  assign \new_[16051]_  = A268 & \new_[16050]_ ;
  assign \new_[16052]_  = \new_[16051]_  & \new_[16046]_ ;
  assign \new_[16055]_  = ~A168 & A170;
  assign \new_[16059]_  = A201 & ~A200;
  assign \new_[16060]_  = A199 & \new_[16059]_ ;
  assign \new_[16061]_  = \new_[16060]_  & \new_[16055]_ ;
  assign \new_[16064]_  = ~A267 & ~A203;
  assign \new_[16068]_  = A299 & A298;
  assign \new_[16069]_  = A268 & \new_[16068]_ ;
  assign \new_[16070]_  = \new_[16069]_  & \new_[16064]_ ;
  assign \new_[16073]_  = ~A168 & A170;
  assign \new_[16077]_  = A201 & ~A200;
  assign \new_[16078]_  = A199 & \new_[16077]_ ;
  assign \new_[16079]_  = \new_[16078]_  & \new_[16073]_ ;
  assign \new_[16082]_  = ~A267 & ~A203;
  assign \new_[16086]_  = ~A299 & ~A298;
  assign \new_[16087]_  = A268 & \new_[16086]_ ;
  assign \new_[16088]_  = \new_[16087]_  & \new_[16082]_ ;
  assign \new_[16091]_  = ~A168 & A170;
  assign \new_[16095]_  = A201 & ~A200;
  assign \new_[16096]_  = A199 & \new_[16095]_ ;
  assign \new_[16097]_  = \new_[16096]_  & \new_[16091]_ ;
  assign \new_[16100]_  = ~A267 & ~A203;
  assign \new_[16104]_  = A301 & ~A300;
  assign \new_[16105]_  = ~A269 & \new_[16104]_ ;
  assign \new_[16106]_  = \new_[16105]_  & \new_[16100]_ ;
  assign \new_[16109]_  = ~A168 & A170;
  assign \new_[16113]_  = A201 & ~A200;
  assign \new_[16114]_  = A199 & \new_[16113]_ ;
  assign \new_[16115]_  = \new_[16114]_  & \new_[16109]_ ;
  assign \new_[16118]_  = ~A267 & ~A203;
  assign \new_[16122]_  = ~A302 & ~A300;
  assign \new_[16123]_  = ~A269 & \new_[16122]_ ;
  assign \new_[16124]_  = \new_[16123]_  & \new_[16118]_ ;
  assign \new_[16127]_  = ~A168 & A170;
  assign \new_[16131]_  = A201 & ~A200;
  assign \new_[16132]_  = A199 & \new_[16131]_ ;
  assign \new_[16133]_  = \new_[16132]_  & \new_[16127]_ ;
  assign \new_[16136]_  = ~A267 & ~A203;
  assign \new_[16140]_  = A299 & A298;
  assign \new_[16141]_  = ~A269 & \new_[16140]_ ;
  assign \new_[16142]_  = \new_[16141]_  & \new_[16136]_ ;
  assign \new_[16145]_  = ~A168 & A170;
  assign \new_[16149]_  = A201 & ~A200;
  assign \new_[16150]_  = A199 & \new_[16149]_ ;
  assign \new_[16151]_  = \new_[16150]_  & \new_[16145]_ ;
  assign \new_[16154]_  = ~A267 & ~A203;
  assign \new_[16158]_  = ~A299 & ~A298;
  assign \new_[16159]_  = ~A269 & \new_[16158]_ ;
  assign \new_[16160]_  = \new_[16159]_  & \new_[16154]_ ;
  assign \new_[16163]_  = ~A168 & A170;
  assign \new_[16167]_  = A201 & ~A200;
  assign \new_[16168]_  = A199 & \new_[16167]_ ;
  assign \new_[16169]_  = \new_[16168]_  & \new_[16163]_ ;
  assign \new_[16172]_  = A265 & ~A203;
  assign \new_[16176]_  = A301 & ~A300;
  assign \new_[16177]_  = A266 & \new_[16176]_ ;
  assign \new_[16178]_  = \new_[16177]_  & \new_[16172]_ ;
  assign \new_[16181]_  = ~A168 & A170;
  assign \new_[16185]_  = A201 & ~A200;
  assign \new_[16186]_  = A199 & \new_[16185]_ ;
  assign \new_[16187]_  = \new_[16186]_  & \new_[16181]_ ;
  assign \new_[16190]_  = A265 & ~A203;
  assign \new_[16194]_  = ~A302 & ~A300;
  assign \new_[16195]_  = A266 & \new_[16194]_ ;
  assign \new_[16196]_  = \new_[16195]_  & \new_[16190]_ ;
  assign \new_[16199]_  = ~A168 & A170;
  assign \new_[16203]_  = A201 & ~A200;
  assign \new_[16204]_  = A199 & \new_[16203]_ ;
  assign \new_[16205]_  = \new_[16204]_  & \new_[16199]_ ;
  assign \new_[16208]_  = A265 & ~A203;
  assign \new_[16212]_  = A299 & A298;
  assign \new_[16213]_  = A266 & \new_[16212]_ ;
  assign \new_[16214]_  = \new_[16213]_  & \new_[16208]_ ;
  assign \new_[16217]_  = ~A168 & A170;
  assign \new_[16221]_  = A201 & ~A200;
  assign \new_[16222]_  = A199 & \new_[16221]_ ;
  assign \new_[16223]_  = \new_[16222]_  & \new_[16217]_ ;
  assign \new_[16226]_  = A265 & ~A203;
  assign \new_[16230]_  = ~A299 & ~A298;
  assign \new_[16231]_  = A266 & \new_[16230]_ ;
  assign \new_[16232]_  = \new_[16231]_  & \new_[16226]_ ;
  assign \new_[16235]_  = ~A168 & A170;
  assign \new_[16239]_  = A201 & ~A200;
  assign \new_[16240]_  = A199 & \new_[16239]_ ;
  assign \new_[16241]_  = \new_[16240]_  & \new_[16235]_ ;
  assign \new_[16244]_  = ~A265 & ~A203;
  assign \new_[16248]_  = A301 & ~A300;
  assign \new_[16249]_  = ~A266 & \new_[16248]_ ;
  assign \new_[16250]_  = \new_[16249]_  & \new_[16244]_ ;
  assign \new_[16253]_  = ~A168 & A170;
  assign \new_[16257]_  = A201 & ~A200;
  assign \new_[16258]_  = A199 & \new_[16257]_ ;
  assign \new_[16259]_  = \new_[16258]_  & \new_[16253]_ ;
  assign \new_[16262]_  = ~A265 & ~A203;
  assign \new_[16266]_  = ~A302 & ~A300;
  assign \new_[16267]_  = ~A266 & \new_[16266]_ ;
  assign \new_[16268]_  = \new_[16267]_  & \new_[16262]_ ;
  assign \new_[16271]_  = ~A168 & A170;
  assign \new_[16275]_  = A201 & ~A200;
  assign \new_[16276]_  = A199 & \new_[16275]_ ;
  assign \new_[16277]_  = \new_[16276]_  & \new_[16271]_ ;
  assign \new_[16280]_  = ~A265 & ~A203;
  assign \new_[16284]_  = A299 & A298;
  assign \new_[16285]_  = ~A266 & \new_[16284]_ ;
  assign \new_[16286]_  = \new_[16285]_  & \new_[16280]_ ;
  assign \new_[16289]_  = ~A168 & A170;
  assign \new_[16293]_  = A201 & ~A200;
  assign \new_[16294]_  = A199 & \new_[16293]_ ;
  assign \new_[16295]_  = \new_[16294]_  & \new_[16289]_ ;
  assign \new_[16298]_  = ~A265 & ~A203;
  assign \new_[16302]_  = ~A299 & ~A298;
  assign \new_[16303]_  = ~A266 & \new_[16302]_ ;
  assign \new_[16304]_  = \new_[16303]_  & \new_[16298]_ ;
  assign \new_[16307]_  = ~A168 & A169;
  assign \new_[16311]_  = A201 & A200;
  assign \new_[16312]_  = ~A199 & \new_[16311]_ ;
  assign \new_[16313]_  = \new_[16312]_  & \new_[16307]_ ;
  assign \new_[16316]_  = ~A267 & A202;
  assign \new_[16320]_  = A301 & ~A300;
  assign \new_[16321]_  = A268 & \new_[16320]_ ;
  assign \new_[16322]_  = \new_[16321]_  & \new_[16316]_ ;
  assign \new_[16325]_  = ~A168 & A169;
  assign \new_[16329]_  = A201 & A200;
  assign \new_[16330]_  = ~A199 & \new_[16329]_ ;
  assign \new_[16331]_  = \new_[16330]_  & \new_[16325]_ ;
  assign \new_[16334]_  = ~A267 & A202;
  assign \new_[16338]_  = ~A302 & ~A300;
  assign \new_[16339]_  = A268 & \new_[16338]_ ;
  assign \new_[16340]_  = \new_[16339]_  & \new_[16334]_ ;
  assign \new_[16343]_  = ~A168 & A169;
  assign \new_[16347]_  = A201 & A200;
  assign \new_[16348]_  = ~A199 & \new_[16347]_ ;
  assign \new_[16349]_  = \new_[16348]_  & \new_[16343]_ ;
  assign \new_[16352]_  = ~A267 & A202;
  assign \new_[16356]_  = A299 & A298;
  assign \new_[16357]_  = A268 & \new_[16356]_ ;
  assign \new_[16358]_  = \new_[16357]_  & \new_[16352]_ ;
  assign \new_[16361]_  = ~A168 & A169;
  assign \new_[16365]_  = A201 & A200;
  assign \new_[16366]_  = ~A199 & \new_[16365]_ ;
  assign \new_[16367]_  = \new_[16366]_  & \new_[16361]_ ;
  assign \new_[16370]_  = ~A267 & A202;
  assign \new_[16374]_  = ~A299 & ~A298;
  assign \new_[16375]_  = A268 & \new_[16374]_ ;
  assign \new_[16376]_  = \new_[16375]_  & \new_[16370]_ ;
  assign \new_[16379]_  = ~A168 & A169;
  assign \new_[16383]_  = A201 & A200;
  assign \new_[16384]_  = ~A199 & \new_[16383]_ ;
  assign \new_[16385]_  = \new_[16384]_  & \new_[16379]_ ;
  assign \new_[16388]_  = ~A267 & A202;
  assign \new_[16392]_  = A301 & ~A300;
  assign \new_[16393]_  = ~A269 & \new_[16392]_ ;
  assign \new_[16394]_  = \new_[16393]_  & \new_[16388]_ ;
  assign \new_[16397]_  = ~A168 & A169;
  assign \new_[16401]_  = A201 & A200;
  assign \new_[16402]_  = ~A199 & \new_[16401]_ ;
  assign \new_[16403]_  = \new_[16402]_  & \new_[16397]_ ;
  assign \new_[16406]_  = ~A267 & A202;
  assign \new_[16410]_  = ~A302 & ~A300;
  assign \new_[16411]_  = ~A269 & \new_[16410]_ ;
  assign \new_[16412]_  = \new_[16411]_  & \new_[16406]_ ;
  assign \new_[16415]_  = ~A168 & A169;
  assign \new_[16419]_  = A201 & A200;
  assign \new_[16420]_  = ~A199 & \new_[16419]_ ;
  assign \new_[16421]_  = \new_[16420]_  & \new_[16415]_ ;
  assign \new_[16424]_  = ~A267 & A202;
  assign \new_[16428]_  = A299 & A298;
  assign \new_[16429]_  = ~A269 & \new_[16428]_ ;
  assign \new_[16430]_  = \new_[16429]_  & \new_[16424]_ ;
  assign \new_[16433]_  = ~A168 & A169;
  assign \new_[16437]_  = A201 & A200;
  assign \new_[16438]_  = ~A199 & \new_[16437]_ ;
  assign \new_[16439]_  = \new_[16438]_  & \new_[16433]_ ;
  assign \new_[16442]_  = ~A267 & A202;
  assign \new_[16446]_  = ~A299 & ~A298;
  assign \new_[16447]_  = ~A269 & \new_[16446]_ ;
  assign \new_[16448]_  = \new_[16447]_  & \new_[16442]_ ;
  assign \new_[16451]_  = ~A168 & A169;
  assign \new_[16455]_  = A201 & A200;
  assign \new_[16456]_  = ~A199 & \new_[16455]_ ;
  assign \new_[16457]_  = \new_[16456]_  & \new_[16451]_ ;
  assign \new_[16460]_  = A265 & A202;
  assign \new_[16464]_  = A301 & ~A300;
  assign \new_[16465]_  = A266 & \new_[16464]_ ;
  assign \new_[16466]_  = \new_[16465]_  & \new_[16460]_ ;
  assign \new_[16469]_  = ~A168 & A169;
  assign \new_[16473]_  = A201 & A200;
  assign \new_[16474]_  = ~A199 & \new_[16473]_ ;
  assign \new_[16475]_  = \new_[16474]_  & \new_[16469]_ ;
  assign \new_[16478]_  = A265 & A202;
  assign \new_[16482]_  = ~A302 & ~A300;
  assign \new_[16483]_  = A266 & \new_[16482]_ ;
  assign \new_[16484]_  = \new_[16483]_  & \new_[16478]_ ;
  assign \new_[16487]_  = ~A168 & A169;
  assign \new_[16491]_  = A201 & A200;
  assign \new_[16492]_  = ~A199 & \new_[16491]_ ;
  assign \new_[16493]_  = \new_[16492]_  & \new_[16487]_ ;
  assign \new_[16496]_  = A265 & A202;
  assign \new_[16500]_  = A299 & A298;
  assign \new_[16501]_  = A266 & \new_[16500]_ ;
  assign \new_[16502]_  = \new_[16501]_  & \new_[16496]_ ;
  assign \new_[16505]_  = ~A168 & A169;
  assign \new_[16509]_  = A201 & A200;
  assign \new_[16510]_  = ~A199 & \new_[16509]_ ;
  assign \new_[16511]_  = \new_[16510]_  & \new_[16505]_ ;
  assign \new_[16514]_  = A265 & A202;
  assign \new_[16518]_  = ~A299 & ~A298;
  assign \new_[16519]_  = A266 & \new_[16518]_ ;
  assign \new_[16520]_  = \new_[16519]_  & \new_[16514]_ ;
  assign \new_[16523]_  = ~A168 & A169;
  assign \new_[16527]_  = A201 & A200;
  assign \new_[16528]_  = ~A199 & \new_[16527]_ ;
  assign \new_[16529]_  = \new_[16528]_  & \new_[16523]_ ;
  assign \new_[16532]_  = ~A265 & A202;
  assign \new_[16536]_  = A301 & ~A300;
  assign \new_[16537]_  = ~A266 & \new_[16536]_ ;
  assign \new_[16538]_  = \new_[16537]_  & \new_[16532]_ ;
  assign \new_[16541]_  = ~A168 & A169;
  assign \new_[16545]_  = A201 & A200;
  assign \new_[16546]_  = ~A199 & \new_[16545]_ ;
  assign \new_[16547]_  = \new_[16546]_  & \new_[16541]_ ;
  assign \new_[16550]_  = ~A265 & A202;
  assign \new_[16554]_  = ~A302 & ~A300;
  assign \new_[16555]_  = ~A266 & \new_[16554]_ ;
  assign \new_[16556]_  = \new_[16555]_  & \new_[16550]_ ;
  assign \new_[16559]_  = ~A168 & A169;
  assign \new_[16563]_  = A201 & A200;
  assign \new_[16564]_  = ~A199 & \new_[16563]_ ;
  assign \new_[16565]_  = \new_[16564]_  & \new_[16559]_ ;
  assign \new_[16568]_  = ~A265 & A202;
  assign \new_[16572]_  = A299 & A298;
  assign \new_[16573]_  = ~A266 & \new_[16572]_ ;
  assign \new_[16574]_  = \new_[16573]_  & \new_[16568]_ ;
  assign \new_[16577]_  = ~A168 & A169;
  assign \new_[16581]_  = A201 & A200;
  assign \new_[16582]_  = ~A199 & \new_[16581]_ ;
  assign \new_[16583]_  = \new_[16582]_  & \new_[16577]_ ;
  assign \new_[16586]_  = ~A265 & A202;
  assign \new_[16590]_  = ~A299 & ~A298;
  assign \new_[16591]_  = ~A266 & \new_[16590]_ ;
  assign \new_[16592]_  = \new_[16591]_  & \new_[16586]_ ;
  assign \new_[16595]_  = ~A168 & A169;
  assign \new_[16599]_  = A201 & A200;
  assign \new_[16600]_  = ~A199 & \new_[16599]_ ;
  assign \new_[16601]_  = \new_[16600]_  & \new_[16595]_ ;
  assign \new_[16604]_  = ~A267 & ~A203;
  assign \new_[16608]_  = A301 & ~A300;
  assign \new_[16609]_  = A268 & \new_[16608]_ ;
  assign \new_[16610]_  = \new_[16609]_  & \new_[16604]_ ;
  assign \new_[16613]_  = ~A168 & A169;
  assign \new_[16617]_  = A201 & A200;
  assign \new_[16618]_  = ~A199 & \new_[16617]_ ;
  assign \new_[16619]_  = \new_[16618]_  & \new_[16613]_ ;
  assign \new_[16622]_  = ~A267 & ~A203;
  assign \new_[16626]_  = ~A302 & ~A300;
  assign \new_[16627]_  = A268 & \new_[16626]_ ;
  assign \new_[16628]_  = \new_[16627]_  & \new_[16622]_ ;
  assign \new_[16631]_  = ~A168 & A169;
  assign \new_[16635]_  = A201 & A200;
  assign \new_[16636]_  = ~A199 & \new_[16635]_ ;
  assign \new_[16637]_  = \new_[16636]_  & \new_[16631]_ ;
  assign \new_[16640]_  = ~A267 & ~A203;
  assign \new_[16644]_  = A299 & A298;
  assign \new_[16645]_  = A268 & \new_[16644]_ ;
  assign \new_[16646]_  = \new_[16645]_  & \new_[16640]_ ;
  assign \new_[16649]_  = ~A168 & A169;
  assign \new_[16653]_  = A201 & A200;
  assign \new_[16654]_  = ~A199 & \new_[16653]_ ;
  assign \new_[16655]_  = \new_[16654]_  & \new_[16649]_ ;
  assign \new_[16658]_  = ~A267 & ~A203;
  assign \new_[16662]_  = ~A299 & ~A298;
  assign \new_[16663]_  = A268 & \new_[16662]_ ;
  assign \new_[16664]_  = \new_[16663]_  & \new_[16658]_ ;
  assign \new_[16667]_  = ~A168 & A169;
  assign \new_[16671]_  = A201 & A200;
  assign \new_[16672]_  = ~A199 & \new_[16671]_ ;
  assign \new_[16673]_  = \new_[16672]_  & \new_[16667]_ ;
  assign \new_[16676]_  = ~A267 & ~A203;
  assign \new_[16680]_  = A301 & ~A300;
  assign \new_[16681]_  = ~A269 & \new_[16680]_ ;
  assign \new_[16682]_  = \new_[16681]_  & \new_[16676]_ ;
  assign \new_[16685]_  = ~A168 & A169;
  assign \new_[16689]_  = A201 & A200;
  assign \new_[16690]_  = ~A199 & \new_[16689]_ ;
  assign \new_[16691]_  = \new_[16690]_  & \new_[16685]_ ;
  assign \new_[16694]_  = ~A267 & ~A203;
  assign \new_[16698]_  = ~A302 & ~A300;
  assign \new_[16699]_  = ~A269 & \new_[16698]_ ;
  assign \new_[16700]_  = \new_[16699]_  & \new_[16694]_ ;
  assign \new_[16703]_  = ~A168 & A169;
  assign \new_[16707]_  = A201 & A200;
  assign \new_[16708]_  = ~A199 & \new_[16707]_ ;
  assign \new_[16709]_  = \new_[16708]_  & \new_[16703]_ ;
  assign \new_[16712]_  = ~A267 & ~A203;
  assign \new_[16716]_  = A299 & A298;
  assign \new_[16717]_  = ~A269 & \new_[16716]_ ;
  assign \new_[16718]_  = \new_[16717]_  & \new_[16712]_ ;
  assign \new_[16721]_  = ~A168 & A169;
  assign \new_[16725]_  = A201 & A200;
  assign \new_[16726]_  = ~A199 & \new_[16725]_ ;
  assign \new_[16727]_  = \new_[16726]_  & \new_[16721]_ ;
  assign \new_[16730]_  = ~A267 & ~A203;
  assign \new_[16734]_  = ~A299 & ~A298;
  assign \new_[16735]_  = ~A269 & \new_[16734]_ ;
  assign \new_[16736]_  = \new_[16735]_  & \new_[16730]_ ;
  assign \new_[16739]_  = ~A168 & A169;
  assign \new_[16743]_  = A201 & A200;
  assign \new_[16744]_  = ~A199 & \new_[16743]_ ;
  assign \new_[16745]_  = \new_[16744]_  & \new_[16739]_ ;
  assign \new_[16748]_  = A265 & ~A203;
  assign \new_[16752]_  = A301 & ~A300;
  assign \new_[16753]_  = A266 & \new_[16752]_ ;
  assign \new_[16754]_  = \new_[16753]_  & \new_[16748]_ ;
  assign \new_[16757]_  = ~A168 & A169;
  assign \new_[16761]_  = A201 & A200;
  assign \new_[16762]_  = ~A199 & \new_[16761]_ ;
  assign \new_[16763]_  = \new_[16762]_  & \new_[16757]_ ;
  assign \new_[16766]_  = A265 & ~A203;
  assign \new_[16770]_  = ~A302 & ~A300;
  assign \new_[16771]_  = A266 & \new_[16770]_ ;
  assign \new_[16772]_  = \new_[16771]_  & \new_[16766]_ ;
  assign \new_[16775]_  = ~A168 & A169;
  assign \new_[16779]_  = A201 & A200;
  assign \new_[16780]_  = ~A199 & \new_[16779]_ ;
  assign \new_[16781]_  = \new_[16780]_  & \new_[16775]_ ;
  assign \new_[16784]_  = A265 & ~A203;
  assign \new_[16788]_  = A299 & A298;
  assign \new_[16789]_  = A266 & \new_[16788]_ ;
  assign \new_[16790]_  = \new_[16789]_  & \new_[16784]_ ;
  assign \new_[16793]_  = ~A168 & A169;
  assign \new_[16797]_  = A201 & A200;
  assign \new_[16798]_  = ~A199 & \new_[16797]_ ;
  assign \new_[16799]_  = \new_[16798]_  & \new_[16793]_ ;
  assign \new_[16802]_  = A265 & ~A203;
  assign \new_[16806]_  = ~A299 & ~A298;
  assign \new_[16807]_  = A266 & \new_[16806]_ ;
  assign \new_[16808]_  = \new_[16807]_  & \new_[16802]_ ;
  assign \new_[16811]_  = ~A168 & A169;
  assign \new_[16815]_  = A201 & A200;
  assign \new_[16816]_  = ~A199 & \new_[16815]_ ;
  assign \new_[16817]_  = \new_[16816]_  & \new_[16811]_ ;
  assign \new_[16820]_  = ~A265 & ~A203;
  assign \new_[16824]_  = A301 & ~A300;
  assign \new_[16825]_  = ~A266 & \new_[16824]_ ;
  assign \new_[16826]_  = \new_[16825]_  & \new_[16820]_ ;
  assign \new_[16829]_  = ~A168 & A169;
  assign \new_[16833]_  = A201 & A200;
  assign \new_[16834]_  = ~A199 & \new_[16833]_ ;
  assign \new_[16835]_  = \new_[16834]_  & \new_[16829]_ ;
  assign \new_[16838]_  = ~A265 & ~A203;
  assign \new_[16842]_  = ~A302 & ~A300;
  assign \new_[16843]_  = ~A266 & \new_[16842]_ ;
  assign \new_[16844]_  = \new_[16843]_  & \new_[16838]_ ;
  assign \new_[16847]_  = ~A168 & A169;
  assign \new_[16851]_  = A201 & A200;
  assign \new_[16852]_  = ~A199 & \new_[16851]_ ;
  assign \new_[16853]_  = \new_[16852]_  & \new_[16847]_ ;
  assign \new_[16856]_  = ~A265 & ~A203;
  assign \new_[16860]_  = A299 & A298;
  assign \new_[16861]_  = ~A266 & \new_[16860]_ ;
  assign \new_[16862]_  = \new_[16861]_  & \new_[16856]_ ;
  assign \new_[16865]_  = ~A168 & A169;
  assign \new_[16869]_  = A201 & A200;
  assign \new_[16870]_  = ~A199 & \new_[16869]_ ;
  assign \new_[16871]_  = \new_[16870]_  & \new_[16865]_ ;
  assign \new_[16874]_  = ~A265 & ~A203;
  assign \new_[16878]_  = ~A299 & ~A298;
  assign \new_[16879]_  = ~A266 & \new_[16878]_ ;
  assign \new_[16880]_  = \new_[16879]_  & \new_[16874]_ ;
  assign \new_[16883]_  = ~A168 & A169;
  assign \new_[16887]_  = A201 & ~A200;
  assign \new_[16888]_  = A199 & \new_[16887]_ ;
  assign \new_[16889]_  = \new_[16888]_  & \new_[16883]_ ;
  assign \new_[16892]_  = ~A267 & A202;
  assign \new_[16896]_  = A301 & ~A300;
  assign \new_[16897]_  = A268 & \new_[16896]_ ;
  assign \new_[16898]_  = \new_[16897]_  & \new_[16892]_ ;
  assign \new_[16901]_  = ~A168 & A169;
  assign \new_[16905]_  = A201 & ~A200;
  assign \new_[16906]_  = A199 & \new_[16905]_ ;
  assign \new_[16907]_  = \new_[16906]_  & \new_[16901]_ ;
  assign \new_[16910]_  = ~A267 & A202;
  assign \new_[16914]_  = ~A302 & ~A300;
  assign \new_[16915]_  = A268 & \new_[16914]_ ;
  assign \new_[16916]_  = \new_[16915]_  & \new_[16910]_ ;
  assign \new_[16919]_  = ~A168 & A169;
  assign \new_[16923]_  = A201 & ~A200;
  assign \new_[16924]_  = A199 & \new_[16923]_ ;
  assign \new_[16925]_  = \new_[16924]_  & \new_[16919]_ ;
  assign \new_[16928]_  = ~A267 & A202;
  assign \new_[16932]_  = A299 & A298;
  assign \new_[16933]_  = A268 & \new_[16932]_ ;
  assign \new_[16934]_  = \new_[16933]_  & \new_[16928]_ ;
  assign \new_[16937]_  = ~A168 & A169;
  assign \new_[16941]_  = A201 & ~A200;
  assign \new_[16942]_  = A199 & \new_[16941]_ ;
  assign \new_[16943]_  = \new_[16942]_  & \new_[16937]_ ;
  assign \new_[16946]_  = ~A267 & A202;
  assign \new_[16950]_  = ~A299 & ~A298;
  assign \new_[16951]_  = A268 & \new_[16950]_ ;
  assign \new_[16952]_  = \new_[16951]_  & \new_[16946]_ ;
  assign \new_[16955]_  = ~A168 & A169;
  assign \new_[16959]_  = A201 & ~A200;
  assign \new_[16960]_  = A199 & \new_[16959]_ ;
  assign \new_[16961]_  = \new_[16960]_  & \new_[16955]_ ;
  assign \new_[16964]_  = ~A267 & A202;
  assign \new_[16968]_  = A301 & ~A300;
  assign \new_[16969]_  = ~A269 & \new_[16968]_ ;
  assign \new_[16970]_  = \new_[16969]_  & \new_[16964]_ ;
  assign \new_[16973]_  = ~A168 & A169;
  assign \new_[16977]_  = A201 & ~A200;
  assign \new_[16978]_  = A199 & \new_[16977]_ ;
  assign \new_[16979]_  = \new_[16978]_  & \new_[16973]_ ;
  assign \new_[16982]_  = ~A267 & A202;
  assign \new_[16986]_  = ~A302 & ~A300;
  assign \new_[16987]_  = ~A269 & \new_[16986]_ ;
  assign \new_[16988]_  = \new_[16987]_  & \new_[16982]_ ;
  assign \new_[16991]_  = ~A168 & A169;
  assign \new_[16995]_  = A201 & ~A200;
  assign \new_[16996]_  = A199 & \new_[16995]_ ;
  assign \new_[16997]_  = \new_[16996]_  & \new_[16991]_ ;
  assign \new_[17000]_  = ~A267 & A202;
  assign \new_[17004]_  = A299 & A298;
  assign \new_[17005]_  = ~A269 & \new_[17004]_ ;
  assign \new_[17006]_  = \new_[17005]_  & \new_[17000]_ ;
  assign \new_[17009]_  = ~A168 & A169;
  assign \new_[17013]_  = A201 & ~A200;
  assign \new_[17014]_  = A199 & \new_[17013]_ ;
  assign \new_[17015]_  = \new_[17014]_  & \new_[17009]_ ;
  assign \new_[17018]_  = ~A267 & A202;
  assign \new_[17022]_  = ~A299 & ~A298;
  assign \new_[17023]_  = ~A269 & \new_[17022]_ ;
  assign \new_[17024]_  = \new_[17023]_  & \new_[17018]_ ;
  assign \new_[17027]_  = ~A168 & A169;
  assign \new_[17031]_  = A201 & ~A200;
  assign \new_[17032]_  = A199 & \new_[17031]_ ;
  assign \new_[17033]_  = \new_[17032]_  & \new_[17027]_ ;
  assign \new_[17036]_  = A265 & A202;
  assign \new_[17040]_  = A301 & ~A300;
  assign \new_[17041]_  = A266 & \new_[17040]_ ;
  assign \new_[17042]_  = \new_[17041]_  & \new_[17036]_ ;
  assign \new_[17045]_  = ~A168 & A169;
  assign \new_[17049]_  = A201 & ~A200;
  assign \new_[17050]_  = A199 & \new_[17049]_ ;
  assign \new_[17051]_  = \new_[17050]_  & \new_[17045]_ ;
  assign \new_[17054]_  = A265 & A202;
  assign \new_[17058]_  = ~A302 & ~A300;
  assign \new_[17059]_  = A266 & \new_[17058]_ ;
  assign \new_[17060]_  = \new_[17059]_  & \new_[17054]_ ;
  assign \new_[17063]_  = ~A168 & A169;
  assign \new_[17067]_  = A201 & ~A200;
  assign \new_[17068]_  = A199 & \new_[17067]_ ;
  assign \new_[17069]_  = \new_[17068]_  & \new_[17063]_ ;
  assign \new_[17072]_  = A265 & A202;
  assign \new_[17076]_  = A299 & A298;
  assign \new_[17077]_  = A266 & \new_[17076]_ ;
  assign \new_[17078]_  = \new_[17077]_  & \new_[17072]_ ;
  assign \new_[17081]_  = ~A168 & A169;
  assign \new_[17085]_  = A201 & ~A200;
  assign \new_[17086]_  = A199 & \new_[17085]_ ;
  assign \new_[17087]_  = \new_[17086]_  & \new_[17081]_ ;
  assign \new_[17090]_  = A265 & A202;
  assign \new_[17094]_  = ~A299 & ~A298;
  assign \new_[17095]_  = A266 & \new_[17094]_ ;
  assign \new_[17096]_  = \new_[17095]_  & \new_[17090]_ ;
  assign \new_[17099]_  = ~A168 & A169;
  assign \new_[17103]_  = A201 & ~A200;
  assign \new_[17104]_  = A199 & \new_[17103]_ ;
  assign \new_[17105]_  = \new_[17104]_  & \new_[17099]_ ;
  assign \new_[17108]_  = ~A265 & A202;
  assign \new_[17112]_  = A301 & ~A300;
  assign \new_[17113]_  = ~A266 & \new_[17112]_ ;
  assign \new_[17114]_  = \new_[17113]_  & \new_[17108]_ ;
  assign \new_[17117]_  = ~A168 & A169;
  assign \new_[17121]_  = A201 & ~A200;
  assign \new_[17122]_  = A199 & \new_[17121]_ ;
  assign \new_[17123]_  = \new_[17122]_  & \new_[17117]_ ;
  assign \new_[17126]_  = ~A265 & A202;
  assign \new_[17130]_  = ~A302 & ~A300;
  assign \new_[17131]_  = ~A266 & \new_[17130]_ ;
  assign \new_[17132]_  = \new_[17131]_  & \new_[17126]_ ;
  assign \new_[17135]_  = ~A168 & A169;
  assign \new_[17139]_  = A201 & ~A200;
  assign \new_[17140]_  = A199 & \new_[17139]_ ;
  assign \new_[17141]_  = \new_[17140]_  & \new_[17135]_ ;
  assign \new_[17144]_  = ~A265 & A202;
  assign \new_[17148]_  = A299 & A298;
  assign \new_[17149]_  = ~A266 & \new_[17148]_ ;
  assign \new_[17150]_  = \new_[17149]_  & \new_[17144]_ ;
  assign \new_[17153]_  = ~A168 & A169;
  assign \new_[17157]_  = A201 & ~A200;
  assign \new_[17158]_  = A199 & \new_[17157]_ ;
  assign \new_[17159]_  = \new_[17158]_  & \new_[17153]_ ;
  assign \new_[17162]_  = ~A265 & A202;
  assign \new_[17166]_  = ~A299 & ~A298;
  assign \new_[17167]_  = ~A266 & \new_[17166]_ ;
  assign \new_[17168]_  = \new_[17167]_  & \new_[17162]_ ;
  assign \new_[17171]_  = ~A168 & A169;
  assign \new_[17175]_  = A201 & ~A200;
  assign \new_[17176]_  = A199 & \new_[17175]_ ;
  assign \new_[17177]_  = \new_[17176]_  & \new_[17171]_ ;
  assign \new_[17180]_  = ~A267 & ~A203;
  assign \new_[17184]_  = A301 & ~A300;
  assign \new_[17185]_  = A268 & \new_[17184]_ ;
  assign \new_[17186]_  = \new_[17185]_  & \new_[17180]_ ;
  assign \new_[17189]_  = ~A168 & A169;
  assign \new_[17193]_  = A201 & ~A200;
  assign \new_[17194]_  = A199 & \new_[17193]_ ;
  assign \new_[17195]_  = \new_[17194]_  & \new_[17189]_ ;
  assign \new_[17198]_  = ~A267 & ~A203;
  assign \new_[17202]_  = ~A302 & ~A300;
  assign \new_[17203]_  = A268 & \new_[17202]_ ;
  assign \new_[17204]_  = \new_[17203]_  & \new_[17198]_ ;
  assign \new_[17207]_  = ~A168 & A169;
  assign \new_[17211]_  = A201 & ~A200;
  assign \new_[17212]_  = A199 & \new_[17211]_ ;
  assign \new_[17213]_  = \new_[17212]_  & \new_[17207]_ ;
  assign \new_[17216]_  = ~A267 & ~A203;
  assign \new_[17220]_  = A299 & A298;
  assign \new_[17221]_  = A268 & \new_[17220]_ ;
  assign \new_[17222]_  = \new_[17221]_  & \new_[17216]_ ;
  assign \new_[17225]_  = ~A168 & A169;
  assign \new_[17229]_  = A201 & ~A200;
  assign \new_[17230]_  = A199 & \new_[17229]_ ;
  assign \new_[17231]_  = \new_[17230]_  & \new_[17225]_ ;
  assign \new_[17234]_  = ~A267 & ~A203;
  assign \new_[17238]_  = ~A299 & ~A298;
  assign \new_[17239]_  = A268 & \new_[17238]_ ;
  assign \new_[17240]_  = \new_[17239]_  & \new_[17234]_ ;
  assign \new_[17243]_  = ~A168 & A169;
  assign \new_[17247]_  = A201 & ~A200;
  assign \new_[17248]_  = A199 & \new_[17247]_ ;
  assign \new_[17249]_  = \new_[17248]_  & \new_[17243]_ ;
  assign \new_[17252]_  = ~A267 & ~A203;
  assign \new_[17256]_  = A301 & ~A300;
  assign \new_[17257]_  = ~A269 & \new_[17256]_ ;
  assign \new_[17258]_  = \new_[17257]_  & \new_[17252]_ ;
  assign \new_[17261]_  = ~A168 & A169;
  assign \new_[17265]_  = A201 & ~A200;
  assign \new_[17266]_  = A199 & \new_[17265]_ ;
  assign \new_[17267]_  = \new_[17266]_  & \new_[17261]_ ;
  assign \new_[17270]_  = ~A267 & ~A203;
  assign \new_[17274]_  = ~A302 & ~A300;
  assign \new_[17275]_  = ~A269 & \new_[17274]_ ;
  assign \new_[17276]_  = \new_[17275]_  & \new_[17270]_ ;
  assign \new_[17279]_  = ~A168 & A169;
  assign \new_[17283]_  = A201 & ~A200;
  assign \new_[17284]_  = A199 & \new_[17283]_ ;
  assign \new_[17285]_  = \new_[17284]_  & \new_[17279]_ ;
  assign \new_[17288]_  = ~A267 & ~A203;
  assign \new_[17292]_  = A299 & A298;
  assign \new_[17293]_  = ~A269 & \new_[17292]_ ;
  assign \new_[17294]_  = \new_[17293]_  & \new_[17288]_ ;
  assign \new_[17297]_  = ~A168 & A169;
  assign \new_[17301]_  = A201 & ~A200;
  assign \new_[17302]_  = A199 & \new_[17301]_ ;
  assign \new_[17303]_  = \new_[17302]_  & \new_[17297]_ ;
  assign \new_[17306]_  = ~A267 & ~A203;
  assign \new_[17310]_  = ~A299 & ~A298;
  assign \new_[17311]_  = ~A269 & \new_[17310]_ ;
  assign \new_[17312]_  = \new_[17311]_  & \new_[17306]_ ;
  assign \new_[17315]_  = ~A168 & A169;
  assign \new_[17319]_  = A201 & ~A200;
  assign \new_[17320]_  = A199 & \new_[17319]_ ;
  assign \new_[17321]_  = \new_[17320]_  & \new_[17315]_ ;
  assign \new_[17324]_  = A265 & ~A203;
  assign \new_[17328]_  = A301 & ~A300;
  assign \new_[17329]_  = A266 & \new_[17328]_ ;
  assign \new_[17330]_  = \new_[17329]_  & \new_[17324]_ ;
  assign \new_[17333]_  = ~A168 & A169;
  assign \new_[17337]_  = A201 & ~A200;
  assign \new_[17338]_  = A199 & \new_[17337]_ ;
  assign \new_[17339]_  = \new_[17338]_  & \new_[17333]_ ;
  assign \new_[17342]_  = A265 & ~A203;
  assign \new_[17346]_  = ~A302 & ~A300;
  assign \new_[17347]_  = A266 & \new_[17346]_ ;
  assign \new_[17348]_  = \new_[17347]_  & \new_[17342]_ ;
  assign \new_[17351]_  = ~A168 & A169;
  assign \new_[17355]_  = A201 & ~A200;
  assign \new_[17356]_  = A199 & \new_[17355]_ ;
  assign \new_[17357]_  = \new_[17356]_  & \new_[17351]_ ;
  assign \new_[17360]_  = A265 & ~A203;
  assign \new_[17364]_  = A299 & A298;
  assign \new_[17365]_  = A266 & \new_[17364]_ ;
  assign \new_[17366]_  = \new_[17365]_  & \new_[17360]_ ;
  assign \new_[17369]_  = ~A168 & A169;
  assign \new_[17373]_  = A201 & ~A200;
  assign \new_[17374]_  = A199 & \new_[17373]_ ;
  assign \new_[17375]_  = \new_[17374]_  & \new_[17369]_ ;
  assign \new_[17378]_  = A265 & ~A203;
  assign \new_[17382]_  = ~A299 & ~A298;
  assign \new_[17383]_  = A266 & \new_[17382]_ ;
  assign \new_[17384]_  = \new_[17383]_  & \new_[17378]_ ;
  assign \new_[17387]_  = ~A168 & A169;
  assign \new_[17391]_  = A201 & ~A200;
  assign \new_[17392]_  = A199 & \new_[17391]_ ;
  assign \new_[17393]_  = \new_[17392]_  & \new_[17387]_ ;
  assign \new_[17396]_  = ~A265 & ~A203;
  assign \new_[17400]_  = A301 & ~A300;
  assign \new_[17401]_  = ~A266 & \new_[17400]_ ;
  assign \new_[17402]_  = \new_[17401]_  & \new_[17396]_ ;
  assign \new_[17405]_  = ~A168 & A169;
  assign \new_[17409]_  = A201 & ~A200;
  assign \new_[17410]_  = A199 & \new_[17409]_ ;
  assign \new_[17411]_  = \new_[17410]_  & \new_[17405]_ ;
  assign \new_[17414]_  = ~A265 & ~A203;
  assign \new_[17418]_  = ~A302 & ~A300;
  assign \new_[17419]_  = ~A266 & \new_[17418]_ ;
  assign \new_[17420]_  = \new_[17419]_  & \new_[17414]_ ;
  assign \new_[17423]_  = ~A168 & A169;
  assign \new_[17427]_  = A201 & ~A200;
  assign \new_[17428]_  = A199 & \new_[17427]_ ;
  assign \new_[17429]_  = \new_[17428]_  & \new_[17423]_ ;
  assign \new_[17432]_  = ~A265 & ~A203;
  assign \new_[17436]_  = A299 & A298;
  assign \new_[17437]_  = ~A266 & \new_[17436]_ ;
  assign \new_[17438]_  = \new_[17437]_  & \new_[17432]_ ;
  assign \new_[17441]_  = ~A168 & A169;
  assign \new_[17445]_  = A201 & ~A200;
  assign \new_[17446]_  = A199 & \new_[17445]_ ;
  assign \new_[17447]_  = \new_[17446]_  & \new_[17441]_ ;
  assign \new_[17450]_  = ~A265 & ~A203;
  assign \new_[17454]_  = ~A299 & ~A298;
  assign \new_[17455]_  = ~A266 & \new_[17454]_ ;
  assign \new_[17456]_  = \new_[17455]_  & \new_[17450]_ ;
  assign \new_[17459]_  = A233 & ~A232;
  assign \new_[17463]_  = A236 & ~A235;
  assign \new_[17464]_  = ~A234 & \new_[17463]_ ;
  assign \new_[17465]_  = \new_[17464]_  & \new_[17459]_ ;
  assign \new_[17469]_  = ~A267 & A266;
  assign \new_[17470]_  = ~A265 & \new_[17469]_ ;
  assign \new_[17474]_  = A300 & A269;
  assign \new_[17475]_  = ~A268 & \new_[17474]_ ;
  assign \new_[17476]_  = \new_[17475]_  & \new_[17470]_ ;
  assign \new_[17479]_  = A233 & ~A232;
  assign \new_[17483]_  = A236 & ~A235;
  assign \new_[17484]_  = ~A234 & \new_[17483]_ ;
  assign \new_[17485]_  = \new_[17484]_  & \new_[17479]_ ;
  assign \new_[17489]_  = ~A267 & ~A266;
  assign \new_[17490]_  = A265 & \new_[17489]_ ;
  assign \new_[17494]_  = A300 & A269;
  assign \new_[17495]_  = ~A268 & \new_[17494]_ ;
  assign \new_[17496]_  = \new_[17495]_  & \new_[17490]_ ;
  assign \new_[17499]_  = ~A233 & A232;
  assign \new_[17503]_  = A236 & ~A235;
  assign \new_[17504]_  = ~A234 & \new_[17503]_ ;
  assign \new_[17505]_  = \new_[17504]_  & \new_[17499]_ ;
  assign \new_[17509]_  = ~A267 & A266;
  assign \new_[17510]_  = ~A265 & \new_[17509]_ ;
  assign \new_[17514]_  = A300 & A269;
  assign \new_[17515]_  = ~A268 & \new_[17514]_ ;
  assign \new_[17516]_  = \new_[17515]_  & \new_[17510]_ ;
  assign \new_[17519]_  = ~A233 & A232;
  assign \new_[17523]_  = A236 & ~A235;
  assign \new_[17524]_  = ~A234 & \new_[17523]_ ;
  assign \new_[17525]_  = \new_[17524]_  & \new_[17519]_ ;
  assign \new_[17529]_  = ~A267 & ~A266;
  assign \new_[17530]_  = A265 & \new_[17529]_ ;
  assign \new_[17534]_  = A300 & A269;
  assign \new_[17535]_  = ~A268 & \new_[17534]_ ;
  assign \new_[17536]_  = \new_[17535]_  & \new_[17530]_ ;
  assign \new_[17539]_  = ~A232 & ~A201;
  assign \new_[17543]_  = ~A235 & ~A234;
  assign \new_[17544]_  = A233 & \new_[17543]_ ;
  assign \new_[17545]_  = \new_[17544]_  & \new_[17539]_ ;
  assign \new_[17549]_  = A266 & ~A265;
  assign \new_[17550]_  = A236 & \new_[17549]_ ;
  assign \new_[17554]_  = A269 & ~A268;
  assign \new_[17555]_  = ~A267 & \new_[17554]_ ;
  assign \new_[17556]_  = \new_[17555]_  & \new_[17550]_ ;
  assign \new_[17559]_  = ~A232 & ~A201;
  assign \new_[17563]_  = ~A235 & ~A234;
  assign \new_[17564]_  = A233 & \new_[17563]_ ;
  assign \new_[17565]_  = \new_[17564]_  & \new_[17559]_ ;
  assign \new_[17569]_  = ~A266 & A265;
  assign \new_[17570]_  = A236 & \new_[17569]_ ;
  assign \new_[17574]_  = A269 & ~A268;
  assign \new_[17575]_  = ~A267 & \new_[17574]_ ;
  assign \new_[17576]_  = \new_[17575]_  & \new_[17570]_ ;
  assign \new_[17579]_  = A232 & ~A201;
  assign \new_[17583]_  = ~A235 & ~A234;
  assign \new_[17584]_  = ~A233 & \new_[17583]_ ;
  assign \new_[17585]_  = \new_[17584]_  & \new_[17579]_ ;
  assign \new_[17589]_  = A266 & ~A265;
  assign \new_[17590]_  = A236 & \new_[17589]_ ;
  assign \new_[17594]_  = A269 & ~A268;
  assign \new_[17595]_  = ~A267 & \new_[17594]_ ;
  assign \new_[17596]_  = \new_[17595]_  & \new_[17590]_ ;
  assign \new_[17599]_  = A232 & ~A201;
  assign \new_[17603]_  = ~A235 & ~A234;
  assign \new_[17604]_  = ~A233 & \new_[17603]_ ;
  assign \new_[17605]_  = \new_[17604]_  & \new_[17599]_ ;
  assign \new_[17609]_  = ~A266 & A265;
  assign \new_[17610]_  = A236 & \new_[17609]_ ;
  assign \new_[17614]_  = A269 & ~A268;
  assign \new_[17615]_  = ~A267 & \new_[17614]_ ;
  assign \new_[17616]_  = \new_[17615]_  & \new_[17610]_ ;
  assign \new_[17619]_  = A166 & A167;
  assign \new_[17623]_  = A234 & A233;
  assign \new_[17624]_  = ~A232 & \new_[17623]_ ;
  assign \new_[17625]_  = \new_[17624]_  & \new_[17619]_ ;
  assign \new_[17629]_  = A266 & ~A265;
  assign \new_[17630]_  = A235 & \new_[17629]_ ;
  assign \new_[17634]_  = A269 & ~A268;
  assign \new_[17635]_  = ~A267 & \new_[17634]_ ;
  assign \new_[17636]_  = \new_[17635]_  & \new_[17630]_ ;
  assign \new_[17639]_  = A166 & A167;
  assign \new_[17643]_  = A234 & A233;
  assign \new_[17644]_  = ~A232 & \new_[17643]_ ;
  assign \new_[17645]_  = \new_[17644]_  & \new_[17639]_ ;
  assign \new_[17649]_  = ~A266 & A265;
  assign \new_[17650]_  = A235 & \new_[17649]_ ;
  assign \new_[17654]_  = A269 & ~A268;
  assign \new_[17655]_  = ~A267 & \new_[17654]_ ;
  assign \new_[17656]_  = \new_[17655]_  & \new_[17650]_ ;
  assign \new_[17659]_  = A166 & A167;
  assign \new_[17663]_  = A234 & A233;
  assign \new_[17664]_  = ~A232 & \new_[17663]_ ;
  assign \new_[17665]_  = \new_[17664]_  & \new_[17659]_ ;
  assign \new_[17669]_  = A266 & ~A265;
  assign \new_[17670]_  = ~A236 & \new_[17669]_ ;
  assign \new_[17674]_  = A269 & ~A268;
  assign \new_[17675]_  = ~A267 & \new_[17674]_ ;
  assign \new_[17676]_  = \new_[17675]_  & \new_[17670]_ ;
  assign \new_[17679]_  = A166 & A167;
  assign \new_[17683]_  = A234 & A233;
  assign \new_[17684]_  = ~A232 & \new_[17683]_ ;
  assign \new_[17685]_  = \new_[17684]_  & \new_[17679]_ ;
  assign \new_[17689]_  = ~A266 & A265;
  assign \new_[17690]_  = ~A236 & \new_[17689]_ ;
  assign \new_[17694]_  = A269 & ~A268;
  assign \new_[17695]_  = ~A267 & \new_[17694]_ ;
  assign \new_[17696]_  = \new_[17695]_  & \new_[17690]_ ;
  assign \new_[17699]_  = A166 & A167;
  assign \new_[17703]_  = A234 & ~A233;
  assign \new_[17704]_  = A232 & \new_[17703]_ ;
  assign \new_[17705]_  = \new_[17704]_  & \new_[17699]_ ;
  assign \new_[17709]_  = A266 & ~A265;
  assign \new_[17710]_  = A235 & \new_[17709]_ ;
  assign \new_[17714]_  = A269 & ~A268;
  assign \new_[17715]_  = ~A267 & \new_[17714]_ ;
  assign \new_[17716]_  = \new_[17715]_  & \new_[17710]_ ;
  assign \new_[17719]_  = A166 & A167;
  assign \new_[17723]_  = A234 & ~A233;
  assign \new_[17724]_  = A232 & \new_[17723]_ ;
  assign \new_[17725]_  = \new_[17724]_  & \new_[17719]_ ;
  assign \new_[17729]_  = ~A266 & A265;
  assign \new_[17730]_  = A235 & \new_[17729]_ ;
  assign \new_[17734]_  = A269 & ~A268;
  assign \new_[17735]_  = ~A267 & \new_[17734]_ ;
  assign \new_[17736]_  = \new_[17735]_  & \new_[17730]_ ;
  assign \new_[17739]_  = A166 & A167;
  assign \new_[17743]_  = A234 & ~A233;
  assign \new_[17744]_  = A232 & \new_[17743]_ ;
  assign \new_[17745]_  = \new_[17744]_  & \new_[17739]_ ;
  assign \new_[17749]_  = A266 & ~A265;
  assign \new_[17750]_  = ~A236 & \new_[17749]_ ;
  assign \new_[17754]_  = A269 & ~A268;
  assign \new_[17755]_  = ~A267 & \new_[17754]_ ;
  assign \new_[17756]_  = \new_[17755]_  & \new_[17750]_ ;
  assign \new_[17759]_  = A166 & A167;
  assign \new_[17763]_  = A234 & ~A233;
  assign \new_[17764]_  = A232 & \new_[17763]_ ;
  assign \new_[17765]_  = \new_[17764]_  & \new_[17759]_ ;
  assign \new_[17769]_  = ~A266 & A265;
  assign \new_[17770]_  = ~A236 & \new_[17769]_ ;
  assign \new_[17774]_  = A269 & ~A268;
  assign \new_[17775]_  = ~A267 & \new_[17774]_ ;
  assign \new_[17776]_  = \new_[17775]_  & \new_[17770]_ ;
  assign \new_[17779]_  = A166 & A167;
  assign \new_[17783]_  = A201 & A200;
  assign \new_[17784]_  = ~A199 & \new_[17783]_ ;
  assign \new_[17785]_  = \new_[17784]_  & \new_[17779]_ ;
  assign \new_[17789]_  = ~A268 & A267;
  assign \new_[17790]_  = A202 & \new_[17789]_ ;
  assign \new_[17794]_  = A301 & ~A300;
  assign \new_[17795]_  = A269 & \new_[17794]_ ;
  assign \new_[17796]_  = \new_[17795]_  & \new_[17790]_ ;
  assign \new_[17799]_  = A166 & A167;
  assign \new_[17803]_  = A201 & A200;
  assign \new_[17804]_  = ~A199 & \new_[17803]_ ;
  assign \new_[17805]_  = \new_[17804]_  & \new_[17799]_ ;
  assign \new_[17809]_  = ~A268 & A267;
  assign \new_[17810]_  = A202 & \new_[17809]_ ;
  assign \new_[17814]_  = ~A302 & ~A300;
  assign \new_[17815]_  = A269 & \new_[17814]_ ;
  assign \new_[17816]_  = \new_[17815]_  & \new_[17810]_ ;
  assign \new_[17819]_  = A166 & A167;
  assign \new_[17823]_  = A201 & A200;
  assign \new_[17824]_  = ~A199 & \new_[17823]_ ;
  assign \new_[17825]_  = \new_[17824]_  & \new_[17819]_ ;
  assign \new_[17829]_  = ~A268 & A267;
  assign \new_[17830]_  = A202 & \new_[17829]_ ;
  assign \new_[17834]_  = A299 & A298;
  assign \new_[17835]_  = A269 & \new_[17834]_ ;
  assign \new_[17836]_  = \new_[17835]_  & \new_[17830]_ ;
  assign \new_[17839]_  = A166 & A167;
  assign \new_[17843]_  = A201 & A200;
  assign \new_[17844]_  = ~A199 & \new_[17843]_ ;
  assign \new_[17845]_  = \new_[17844]_  & \new_[17839]_ ;
  assign \new_[17849]_  = ~A268 & A267;
  assign \new_[17850]_  = A202 & \new_[17849]_ ;
  assign \new_[17854]_  = ~A299 & ~A298;
  assign \new_[17855]_  = A269 & \new_[17854]_ ;
  assign \new_[17856]_  = \new_[17855]_  & \new_[17850]_ ;
  assign \new_[17859]_  = A166 & A167;
  assign \new_[17863]_  = A201 & A200;
  assign \new_[17864]_  = ~A199 & \new_[17863]_ ;
  assign \new_[17865]_  = \new_[17864]_  & \new_[17859]_ ;
  assign \new_[17869]_  = A268 & ~A267;
  assign \new_[17870]_  = A202 & \new_[17869]_ ;
  assign \new_[17874]_  = A302 & ~A301;
  assign \new_[17875]_  = A300 & \new_[17874]_ ;
  assign \new_[17876]_  = \new_[17875]_  & \new_[17870]_ ;
  assign \new_[17879]_  = A166 & A167;
  assign \new_[17883]_  = A201 & A200;
  assign \new_[17884]_  = ~A199 & \new_[17883]_ ;
  assign \new_[17885]_  = \new_[17884]_  & \new_[17879]_ ;
  assign \new_[17889]_  = ~A269 & ~A267;
  assign \new_[17890]_  = A202 & \new_[17889]_ ;
  assign \new_[17894]_  = A302 & ~A301;
  assign \new_[17895]_  = A300 & \new_[17894]_ ;
  assign \new_[17896]_  = \new_[17895]_  & \new_[17890]_ ;
  assign \new_[17899]_  = A166 & A167;
  assign \new_[17903]_  = A201 & A200;
  assign \new_[17904]_  = ~A199 & \new_[17903]_ ;
  assign \new_[17905]_  = \new_[17904]_  & \new_[17899]_ ;
  assign \new_[17909]_  = A266 & A265;
  assign \new_[17910]_  = A202 & \new_[17909]_ ;
  assign \new_[17914]_  = A302 & ~A301;
  assign \new_[17915]_  = A300 & \new_[17914]_ ;
  assign \new_[17916]_  = \new_[17915]_  & \new_[17910]_ ;
  assign \new_[17919]_  = A166 & A167;
  assign \new_[17923]_  = A201 & A200;
  assign \new_[17924]_  = ~A199 & \new_[17923]_ ;
  assign \new_[17925]_  = \new_[17924]_  & \new_[17919]_ ;
  assign \new_[17929]_  = ~A266 & ~A265;
  assign \new_[17930]_  = A202 & \new_[17929]_ ;
  assign \new_[17934]_  = A302 & ~A301;
  assign \new_[17935]_  = A300 & \new_[17934]_ ;
  assign \new_[17936]_  = \new_[17935]_  & \new_[17930]_ ;
  assign \new_[17939]_  = A166 & A167;
  assign \new_[17943]_  = A201 & A200;
  assign \new_[17944]_  = ~A199 & \new_[17943]_ ;
  assign \new_[17945]_  = \new_[17944]_  & \new_[17939]_ ;
  assign \new_[17949]_  = ~A268 & A267;
  assign \new_[17950]_  = ~A203 & \new_[17949]_ ;
  assign \new_[17954]_  = A301 & ~A300;
  assign \new_[17955]_  = A269 & \new_[17954]_ ;
  assign \new_[17956]_  = \new_[17955]_  & \new_[17950]_ ;
  assign \new_[17959]_  = A166 & A167;
  assign \new_[17963]_  = A201 & A200;
  assign \new_[17964]_  = ~A199 & \new_[17963]_ ;
  assign \new_[17965]_  = \new_[17964]_  & \new_[17959]_ ;
  assign \new_[17969]_  = ~A268 & A267;
  assign \new_[17970]_  = ~A203 & \new_[17969]_ ;
  assign \new_[17974]_  = ~A302 & ~A300;
  assign \new_[17975]_  = A269 & \new_[17974]_ ;
  assign \new_[17976]_  = \new_[17975]_  & \new_[17970]_ ;
  assign \new_[17979]_  = A166 & A167;
  assign \new_[17983]_  = A201 & A200;
  assign \new_[17984]_  = ~A199 & \new_[17983]_ ;
  assign \new_[17985]_  = \new_[17984]_  & \new_[17979]_ ;
  assign \new_[17989]_  = ~A268 & A267;
  assign \new_[17990]_  = ~A203 & \new_[17989]_ ;
  assign \new_[17994]_  = A299 & A298;
  assign \new_[17995]_  = A269 & \new_[17994]_ ;
  assign \new_[17996]_  = \new_[17995]_  & \new_[17990]_ ;
  assign \new_[17999]_  = A166 & A167;
  assign \new_[18003]_  = A201 & A200;
  assign \new_[18004]_  = ~A199 & \new_[18003]_ ;
  assign \new_[18005]_  = \new_[18004]_  & \new_[17999]_ ;
  assign \new_[18009]_  = ~A268 & A267;
  assign \new_[18010]_  = ~A203 & \new_[18009]_ ;
  assign \new_[18014]_  = ~A299 & ~A298;
  assign \new_[18015]_  = A269 & \new_[18014]_ ;
  assign \new_[18016]_  = \new_[18015]_  & \new_[18010]_ ;
  assign \new_[18019]_  = A166 & A167;
  assign \new_[18023]_  = A201 & A200;
  assign \new_[18024]_  = ~A199 & \new_[18023]_ ;
  assign \new_[18025]_  = \new_[18024]_  & \new_[18019]_ ;
  assign \new_[18029]_  = A268 & ~A267;
  assign \new_[18030]_  = ~A203 & \new_[18029]_ ;
  assign \new_[18034]_  = A302 & ~A301;
  assign \new_[18035]_  = A300 & \new_[18034]_ ;
  assign \new_[18036]_  = \new_[18035]_  & \new_[18030]_ ;
  assign \new_[18039]_  = A166 & A167;
  assign \new_[18043]_  = A201 & A200;
  assign \new_[18044]_  = ~A199 & \new_[18043]_ ;
  assign \new_[18045]_  = \new_[18044]_  & \new_[18039]_ ;
  assign \new_[18049]_  = ~A269 & ~A267;
  assign \new_[18050]_  = ~A203 & \new_[18049]_ ;
  assign \new_[18054]_  = A302 & ~A301;
  assign \new_[18055]_  = A300 & \new_[18054]_ ;
  assign \new_[18056]_  = \new_[18055]_  & \new_[18050]_ ;
  assign \new_[18059]_  = A166 & A167;
  assign \new_[18063]_  = A201 & A200;
  assign \new_[18064]_  = ~A199 & \new_[18063]_ ;
  assign \new_[18065]_  = \new_[18064]_  & \new_[18059]_ ;
  assign \new_[18069]_  = A266 & A265;
  assign \new_[18070]_  = ~A203 & \new_[18069]_ ;
  assign \new_[18074]_  = A302 & ~A301;
  assign \new_[18075]_  = A300 & \new_[18074]_ ;
  assign \new_[18076]_  = \new_[18075]_  & \new_[18070]_ ;
  assign \new_[18079]_  = A166 & A167;
  assign \new_[18083]_  = A201 & A200;
  assign \new_[18084]_  = ~A199 & \new_[18083]_ ;
  assign \new_[18085]_  = \new_[18084]_  & \new_[18079]_ ;
  assign \new_[18089]_  = ~A266 & ~A265;
  assign \new_[18090]_  = ~A203 & \new_[18089]_ ;
  assign \new_[18094]_  = A302 & ~A301;
  assign \new_[18095]_  = A300 & \new_[18094]_ ;
  assign \new_[18096]_  = \new_[18095]_  & \new_[18090]_ ;
  assign \new_[18099]_  = A166 & A167;
  assign \new_[18103]_  = ~A201 & A200;
  assign \new_[18104]_  = ~A199 & \new_[18103]_ ;
  assign \new_[18105]_  = \new_[18104]_  & \new_[18099]_ ;
  assign \new_[18109]_  = ~A267 & A203;
  assign \new_[18110]_  = ~A202 & \new_[18109]_ ;
  assign \new_[18114]_  = A301 & ~A300;
  assign \new_[18115]_  = A268 & \new_[18114]_ ;
  assign \new_[18116]_  = \new_[18115]_  & \new_[18110]_ ;
  assign \new_[18119]_  = A166 & A167;
  assign \new_[18123]_  = ~A201 & A200;
  assign \new_[18124]_  = ~A199 & \new_[18123]_ ;
  assign \new_[18125]_  = \new_[18124]_  & \new_[18119]_ ;
  assign \new_[18129]_  = ~A267 & A203;
  assign \new_[18130]_  = ~A202 & \new_[18129]_ ;
  assign \new_[18134]_  = ~A302 & ~A300;
  assign \new_[18135]_  = A268 & \new_[18134]_ ;
  assign \new_[18136]_  = \new_[18135]_  & \new_[18130]_ ;
  assign \new_[18139]_  = A166 & A167;
  assign \new_[18143]_  = ~A201 & A200;
  assign \new_[18144]_  = ~A199 & \new_[18143]_ ;
  assign \new_[18145]_  = \new_[18144]_  & \new_[18139]_ ;
  assign \new_[18149]_  = ~A267 & A203;
  assign \new_[18150]_  = ~A202 & \new_[18149]_ ;
  assign \new_[18154]_  = A299 & A298;
  assign \new_[18155]_  = A268 & \new_[18154]_ ;
  assign \new_[18156]_  = \new_[18155]_  & \new_[18150]_ ;
  assign \new_[18159]_  = A166 & A167;
  assign \new_[18163]_  = ~A201 & A200;
  assign \new_[18164]_  = ~A199 & \new_[18163]_ ;
  assign \new_[18165]_  = \new_[18164]_  & \new_[18159]_ ;
  assign \new_[18169]_  = ~A267 & A203;
  assign \new_[18170]_  = ~A202 & \new_[18169]_ ;
  assign \new_[18174]_  = ~A299 & ~A298;
  assign \new_[18175]_  = A268 & \new_[18174]_ ;
  assign \new_[18176]_  = \new_[18175]_  & \new_[18170]_ ;
  assign \new_[18179]_  = A166 & A167;
  assign \new_[18183]_  = ~A201 & A200;
  assign \new_[18184]_  = ~A199 & \new_[18183]_ ;
  assign \new_[18185]_  = \new_[18184]_  & \new_[18179]_ ;
  assign \new_[18189]_  = ~A267 & A203;
  assign \new_[18190]_  = ~A202 & \new_[18189]_ ;
  assign \new_[18194]_  = A301 & ~A300;
  assign \new_[18195]_  = ~A269 & \new_[18194]_ ;
  assign \new_[18196]_  = \new_[18195]_  & \new_[18190]_ ;
  assign \new_[18199]_  = A166 & A167;
  assign \new_[18203]_  = ~A201 & A200;
  assign \new_[18204]_  = ~A199 & \new_[18203]_ ;
  assign \new_[18205]_  = \new_[18204]_  & \new_[18199]_ ;
  assign \new_[18209]_  = ~A267 & A203;
  assign \new_[18210]_  = ~A202 & \new_[18209]_ ;
  assign \new_[18214]_  = ~A302 & ~A300;
  assign \new_[18215]_  = ~A269 & \new_[18214]_ ;
  assign \new_[18216]_  = \new_[18215]_  & \new_[18210]_ ;
  assign \new_[18219]_  = A166 & A167;
  assign \new_[18223]_  = ~A201 & A200;
  assign \new_[18224]_  = ~A199 & \new_[18223]_ ;
  assign \new_[18225]_  = \new_[18224]_  & \new_[18219]_ ;
  assign \new_[18229]_  = ~A267 & A203;
  assign \new_[18230]_  = ~A202 & \new_[18229]_ ;
  assign \new_[18234]_  = A299 & A298;
  assign \new_[18235]_  = ~A269 & \new_[18234]_ ;
  assign \new_[18236]_  = \new_[18235]_  & \new_[18230]_ ;
  assign \new_[18239]_  = A166 & A167;
  assign \new_[18243]_  = ~A201 & A200;
  assign \new_[18244]_  = ~A199 & \new_[18243]_ ;
  assign \new_[18245]_  = \new_[18244]_  & \new_[18239]_ ;
  assign \new_[18249]_  = ~A267 & A203;
  assign \new_[18250]_  = ~A202 & \new_[18249]_ ;
  assign \new_[18254]_  = ~A299 & ~A298;
  assign \new_[18255]_  = ~A269 & \new_[18254]_ ;
  assign \new_[18256]_  = \new_[18255]_  & \new_[18250]_ ;
  assign \new_[18259]_  = A166 & A167;
  assign \new_[18263]_  = ~A201 & A200;
  assign \new_[18264]_  = ~A199 & \new_[18263]_ ;
  assign \new_[18265]_  = \new_[18264]_  & \new_[18259]_ ;
  assign \new_[18269]_  = A265 & A203;
  assign \new_[18270]_  = ~A202 & \new_[18269]_ ;
  assign \new_[18274]_  = A301 & ~A300;
  assign \new_[18275]_  = A266 & \new_[18274]_ ;
  assign \new_[18276]_  = \new_[18275]_  & \new_[18270]_ ;
  assign \new_[18279]_  = A166 & A167;
  assign \new_[18283]_  = ~A201 & A200;
  assign \new_[18284]_  = ~A199 & \new_[18283]_ ;
  assign \new_[18285]_  = \new_[18284]_  & \new_[18279]_ ;
  assign \new_[18289]_  = A265 & A203;
  assign \new_[18290]_  = ~A202 & \new_[18289]_ ;
  assign \new_[18294]_  = ~A302 & ~A300;
  assign \new_[18295]_  = A266 & \new_[18294]_ ;
  assign \new_[18296]_  = \new_[18295]_  & \new_[18290]_ ;
  assign \new_[18299]_  = A166 & A167;
  assign \new_[18303]_  = ~A201 & A200;
  assign \new_[18304]_  = ~A199 & \new_[18303]_ ;
  assign \new_[18305]_  = \new_[18304]_  & \new_[18299]_ ;
  assign \new_[18309]_  = A265 & A203;
  assign \new_[18310]_  = ~A202 & \new_[18309]_ ;
  assign \new_[18314]_  = A299 & A298;
  assign \new_[18315]_  = A266 & \new_[18314]_ ;
  assign \new_[18316]_  = \new_[18315]_  & \new_[18310]_ ;
  assign \new_[18319]_  = A166 & A167;
  assign \new_[18323]_  = ~A201 & A200;
  assign \new_[18324]_  = ~A199 & \new_[18323]_ ;
  assign \new_[18325]_  = \new_[18324]_  & \new_[18319]_ ;
  assign \new_[18329]_  = A265 & A203;
  assign \new_[18330]_  = ~A202 & \new_[18329]_ ;
  assign \new_[18334]_  = ~A299 & ~A298;
  assign \new_[18335]_  = A266 & \new_[18334]_ ;
  assign \new_[18336]_  = \new_[18335]_  & \new_[18330]_ ;
  assign \new_[18339]_  = A166 & A167;
  assign \new_[18343]_  = ~A201 & A200;
  assign \new_[18344]_  = ~A199 & \new_[18343]_ ;
  assign \new_[18345]_  = \new_[18344]_  & \new_[18339]_ ;
  assign \new_[18349]_  = ~A265 & A203;
  assign \new_[18350]_  = ~A202 & \new_[18349]_ ;
  assign \new_[18354]_  = A301 & ~A300;
  assign \new_[18355]_  = ~A266 & \new_[18354]_ ;
  assign \new_[18356]_  = \new_[18355]_  & \new_[18350]_ ;
  assign \new_[18359]_  = A166 & A167;
  assign \new_[18363]_  = ~A201 & A200;
  assign \new_[18364]_  = ~A199 & \new_[18363]_ ;
  assign \new_[18365]_  = \new_[18364]_  & \new_[18359]_ ;
  assign \new_[18369]_  = ~A265 & A203;
  assign \new_[18370]_  = ~A202 & \new_[18369]_ ;
  assign \new_[18374]_  = ~A302 & ~A300;
  assign \new_[18375]_  = ~A266 & \new_[18374]_ ;
  assign \new_[18376]_  = \new_[18375]_  & \new_[18370]_ ;
  assign \new_[18379]_  = A166 & A167;
  assign \new_[18383]_  = ~A201 & A200;
  assign \new_[18384]_  = ~A199 & \new_[18383]_ ;
  assign \new_[18385]_  = \new_[18384]_  & \new_[18379]_ ;
  assign \new_[18389]_  = ~A265 & A203;
  assign \new_[18390]_  = ~A202 & \new_[18389]_ ;
  assign \new_[18394]_  = A299 & A298;
  assign \new_[18395]_  = ~A266 & \new_[18394]_ ;
  assign \new_[18396]_  = \new_[18395]_  & \new_[18390]_ ;
  assign \new_[18399]_  = A166 & A167;
  assign \new_[18403]_  = ~A201 & A200;
  assign \new_[18404]_  = ~A199 & \new_[18403]_ ;
  assign \new_[18405]_  = \new_[18404]_  & \new_[18399]_ ;
  assign \new_[18409]_  = ~A265 & A203;
  assign \new_[18410]_  = ~A202 & \new_[18409]_ ;
  assign \new_[18414]_  = ~A299 & ~A298;
  assign \new_[18415]_  = ~A266 & \new_[18414]_ ;
  assign \new_[18416]_  = \new_[18415]_  & \new_[18410]_ ;
  assign \new_[18419]_  = A166 & A167;
  assign \new_[18423]_  = A201 & ~A200;
  assign \new_[18424]_  = A199 & \new_[18423]_ ;
  assign \new_[18425]_  = \new_[18424]_  & \new_[18419]_ ;
  assign \new_[18429]_  = ~A268 & A267;
  assign \new_[18430]_  = A202 & \new_[18429]_ ;
  assign \new_[18434]_  = A301 & ~A300;
  assign \new_[18435]_  = A269 & \new_[18434]_ ;
  assign \new_[18436]_  = \new_[18435]_  & \new_[18430]_ ;
  assign \new_[18439]_  = A166 & A167;
  assign \new_[18443]_  = A201 & ~A200;
  assign \new_[18444]_  = A199 & \new_[18443]_ ;
  assign \new_[18445]_  = \new_[18444]_  & \new_[18439]_ ;
  assign \new_[18449]_  = ~A268 & A267;
  assign \new_[18450]_  = A202 & \new_[18449]_ ;
  assign \new_[18454]_  = ~A302 & ~A300;
  assign \new_[18455]_  = A269 & \new_[18454]_ ;
  assign \new_[18456]_  = \new_[18455]_  & \new_[18450]_ ;
  assign \new_[18459]_  = A166 & A167;
  assign \new_[18463]_  = A201 & ~A200;
  assign \new_[18464]_  = A199 & \new_[18463]_ ;
  assign \new_[18465]_  = \new_[18464]_  & \new_[18459]_ ;
  assign \new_[18469]_  = ~A268 & A267;
  assign \new_[18470]_  = A202 & \new_[18469]_ ;
  assign \new_[18474]_  = A299 & A298;
  assign \new_[18475]_  = A269 & \new_[18474]_ ;
  assign \new_[18476]_  = \new_[18475]_  & \new_[18470]_ ;
  assign \new_[18479]_  = A166 & A167;
  assign \new_[18483]_  = A201 & ~A200;
  assign \new_[18484]_  = A199 & \new_[18483]_ ;
  assign \new_[18485]_  = \new_[18484]_  & \new_[18479]_ ;
  assign \new_[18489]_  = ~A268 & A267;
  assign \new_[18490]_  = A202 & \new_[18489]_ ;
  assign \new_[18494]_  = ~A299 & ~A298;
  assign \new_[18495]_  = A269 & \new_[18494]_ ;
  assign \new_[18496]_  = \new_[18495]_  & \new_[18490]_ ;
  assign \new_[18499]_  = A166 & A167;
  assign \new_[18503]_  = A201 & ~A200;
  assign \new_[18504]_  = A199 & \new_[18503]_ ;
  assign \new_[18505]_  = \new_[18504]_  & \new_[18499]_ ;
  assign \new_[18509]_  = A268 & ~A267;
  assign \new_[18510]_  = A202 & \new_[18509]_ ;
  assign \new_[18514]_  = A302 & ~A301;
  assign \new_[18515]_  = A300 & \new_[18514]_ ;
  assign \new_[18516]_  = \new_[18515]_  & \new_[18510]_ ;
  assign \new_[18519]_  = A166 & A167;
  assign \new_[18523]_  = A201 & ~A200;
  assign \new_[18524]_  = A199 & \new_[18523]_ ;
  assign \new_[18525]_  = \new_[18524]_  & \new_[18519]_ ;
  assign \new_[18529]_  = ~A269 & ~A267;
  assign \new_[18530]_  = A202 & \new_[18529]_ ;
  assign \new_[18534]_  = A302 & ~A301;
  assign \new_[18535]_  = A300 & \new_[18534]_ ;
  assign \new_[18536]_  = \new_[18535]_  & \new_[18530]_ ;
  assign \new_[18539]_  = A166 & A167;
  assign \new_[18543]_  = A201 & ~A200;
  assign \new_[18544]_  = A199 & \new_[18543]_ ;
  assign \new_[18545]_  = \new_[18544]_  & \new_[18539]_ ;
  assign \new_[18549]_  = A266 & A265;
  assign \new_[18550]_  = A202 & \new_[18549]_ ;
  assign \new_[18554]_  = A302 & ~A301;
  assign \new_[18555]_  = A300 & \new_[18554]_ ;
  assign \new_[18556]_  = \new_[18555]_  & \new_[18550]_ ;
  assign \new_[18559]_  = A166 & A167;
  assign \new_[18563]_  = A201 & ~A200;
  assign \new_[18564]_  = A199 & \new_[18563]_ ;
  assign \new_[18565]_  = \new_[18564]_  & \new_[18559]_ ;
  assign \new_[18569]_  = ~A266 & ~A265;
  assign \new_[18570]_  = A202 & \new_[18569]_ ;
  assign \new_[18574]_  = A302 & ~A301;
  assign \new_[18575]_  = A300 & \new_[18574]_ ;
  assign \new_[18576]_  = \new_[18575]_  & \new_[18570]_ ;
  assign \new_[18579]_  = A166 & A167;
  assign \new_[18583]_  = A201 & ~A200;
  assign \new_[18584]_  = A199 & \new_[18583]_ ;
  assign \new_[18585]_  = \new_[18584]_  & \new_[18579]_ ;
  assign \new_[18589]_  = ~A268 & A267;
  assign \new_[18590]_  = ~A203 & \new_[18589]_ ;
  assign \new_[18594]_  = A301 & ~A300;
  assign \new_[18595]_  = A269 & \new_[18594]_ ;
  assign \new_[18596]_  = \new_[18595]_  & \new_[18590]_ ;
  assign \new_[18599]_  = A166 & A167;
  assign \new_[18603]_  = A201 & ~A200;
  assign \new_[18604]_  = A199 & \new_[18603]_ ;
  assign \new_[18605]_  = \new_[18604]_  & \new_[18599]_ ;
  assign \new_[18609]_  = ~A268 & A267;
  assign \new_[18610]_  = ~A203 & \new_[18609]_ ;
  assign \new_[18614]_  = ~A302 & ~A300;
  assign \new_[18615]_  = A269 & \new_[18614]_ ;
  assign \new_[18616]_  = \new_[18615]_  & \new_[18610]_ ;
  assign \new_[18619]_  = A166 & A167;
  assign \new_[18623]_  = A201 & ~A200;
  assign \new_[18624]_  = A199 & \new_[18623]_ ;
  assign \new_[18625]_  = \new_[18624]_  & \new_[18619]_ ;
  assign \new_[18629]_  = ~A268 & A267;
  assign \new_[18630]_  = ~A203 & \new_[18629]_ ;
  assign \new_[18634]_  = A299 & A298;
  assign \new_[18635]_  = A269 & \new_[18634]_ ;
  assign \new_[18636]_  = \new_[18635]_  & \new_[18630]_ ;
  assign \new_[18639]_  = A166 & A167;
  assign \new_[18643]_  = A201 & ~A200;
  assign \new_[18644]_  = A199 & \new_[18643]_ ;
  assign \new_[18645]_  = \new_[18644]_  & \new_[18639]_ ;
  assign \new_[18649]_  = ~A268 & A267;
  assign \new_[18650]_  = ~A203 & \new_[18649]_ ;
  assign \new_[18654]_  = ~A299 & ~A298;
  assign \new_[18655]_  = A269 & \new_[18654]_ ;
  assign \new_[18656]_  = \new_[18655]_  & \new_[18650]_ ;
  assign \new_[18659]_  = A166 & A167;
  assign \new_[18663]_  = A201 & ~A200;
  assign \new_[18664]_  = A199 & \new_[18663]_ ;
  assign \new_[18665]_  = \new_[18664]_  & \new_[18659]_ ;
  assign \new_[18669]_  = A268 & ~A267;
  assign \new_[18670]_  = ~A203 & \new_[18669]_ ;
  assign \new_[18674]_  = A302 & ~A301;
  assign \new_[18675]_  = A300 & \new_[18674]_ ;
  assign \new_[18676]_  = \new_[18675]_  & \new_[18670]_ ;
  assign \new_[18679]_  = A166 & A167;
  assign \new_[18683]_  = A201 & ~A200;
  assign \new_[18684]_  = A199 & \new_[18683]_ ;
  assign \new_[18685]_  = \new_[18684]_  & \new_[18679]_ ;
  assign \new_[18689]_  = ~A269 & ~A267;
  assign \new_[18690]_  = ~A203 & \new_[18689]_ ;
  assign \new_[18694]_  = A302 & ~A301;
  assign \new_[18695]_  = A300 & \new_[18694]_ ;
  assign \new_[18696]_  = \new_[18695]_  & \new_[18690]_ ;
  assign \new_[18699]_  = A166 & A167;
  assign \new_[18703]_  = A201 & ~A200;
  assign \new_[18704]_  = A199 & \new_[18703]_ ;
  assign \new_[18705]_  = \new_[18704]_  & \new_[18699]_ ;
  assign \new_[18709]_  = A266 & A265;
  assign \new_[18710]_  = ~A203 & \new_[18709]_ ;
  assign \new_[18714]_  = A302 & ~A301;
  assign \new_[18715]_  = A300 & \new_[18714]_ ;
  assign \new_[18716]_  = \new_[18715]_  & \new_[18710]_ ;
  assign \new_[18719]_  = A166 & A167;
  assign \new_[18723]_  = A201 & ~A200;
  assign \new_[18724]_  = A199 & \new_[18723]_ ;
  assign \new_[18725]_  = \new_[18724]_  & \new_[18719]_ ;
  assign \new_[18729]_  = ~A266 & ~A265;
  assign \new_[18730]_  = ~A203 & \new_[18729]_ ;
  assign \new_[18734]_  = A302 & ~A301;
  assign \new_[18735]_  = A300 & \new_[18734]_ ;
  assign \new_[18736]_  = \new_[18735]_  & \new_[18730]_ ;
  assign \new_[18739]_  = A166 & A167;
  assign \new_[18743]_  = ~A201 & ~A200;
  assign \new_[18744]_  = A199 & \new_[18743]_ ;
  assign \new_[18745]_  = \new_[18744]_  & \new_[18739]_ ;
  assign \new_[18749]_  = ~A267 & A203;
  assign \new_[18750]_  = ~A202 & \new_[18749]_ ;
  assign \new_[18754]_  = A301 & ~A300;
  assign \new_[18755]_  = A268 & \new_[18754]_ ;
  assign \new_[18756]_  = \new_[18755]_  & \new_[18750]_ ;
  assign \new_[18759]_  = A166 & A167;
  assign \new_[18763]_  = ~A201 & ~A200;
  assign \new_[18764]_  = A199 & \new_[18763]_ ;
  assign \new_[18765]_  = \new_[18764]_  & \new_[18759]_ ;
  assign \new_[18769]_  = ~A267 & A203;
  assign \new_[18770]_  = ~A202 & \new_[18769]_ ;
  assign \new_[18774]_  = ~A302 & ~A300;
  assign \new_[18775]_  = A268 & \new_[18774]_ ;
  assign \new_[18776]_  = \new_[18775]_  & \new_[18770]_ ;
  assign \new_[18779]_  = A166 & A167;
  assign \new_[18783]_  = ~A201 & ~A200;
  assign \new_[18784]_  = A199 & \new_[18783]_ ;
  assign \new_[18785]_  = \new_[18784]_  & \new_[18779]_ ;
  assign \new_[18789]_  = ~A267 & A203;
  assign \new_[18790]_  = ~A202 & \new_[18789]_ ;
  assign \new_[18794]_  = A299 & A298;
  assign \new_[18795]_  = A268 & \new_[18794]_ ;
  assign \new_[18796]_  = \new_[18795]_  & \new_[18790]_ ;
  assign \new_[18799]_  = A166 & A167;
  assign \new_[18803]_  = ~A201 & ~A200;
  assign \new_[18804]_  = A199 & \new_[18803]_ ;
  assign \new_[18805]_  = \new_[18804]_  & \new_[18799]_ ;
  assign \new_[18809]_  = ~A267 & A203;
  assign \new_[18810]_  = ~A202 & \new_[18809]_ ;
  assign \new_[18814]_  = ~A299 & ~A298;
  assign \new_[18815]_  = A268 & \new_[18814]_ ;
  assign \new_[18816]_  = \new_[18815]_  & \new_[18810]_ ;
  assign \new_[18819]_  = A166 & A167;
  assign \new_[18823]_  = ~A201 & ~A200;
  assign \new_[18824]_  = A199 & \new_[18823]_ ;
  assign \new_[18825]_  = \new_[18824]_  & \new_[18819]_ ;
  assign \new_[18829]_  = ~A267 & A203;
  assign \new_[18830]_  = ~A202 & \new_[18829]_ ;
  assign \new_[18834]_  = A301 & ~A300;
  assign \new_[18835]_  = ~A269 & \new_[18834]_ ;
  assign \new_[18836]_  = \new_[18835]_  & \new_[18830]_ ;
  assign \new_[18839]_  = A166 & A167;
  assign \new_[18843]_  = ~A201 & ~A200;
  assign \new_[18844]_  = A199 & \new_[18843]_ ;
  assign \new_[18845]_  = \new_[18844]_  & \new_[18839]_ ;
  assign \new_[18849]_  = ~A267 & A203;
  assign \new_[18850]_  = ~A202 & \new_[18849]_ ;
  assign \new_[18854]_  = ~A302 & ~A300;
  assign \new_[18855]_  = ~A269 & \new_[18854]_ ;
  assign \new_[18856]_  = \new_[18855]_  & \new_[18850]_ ;
  assign \new_[18859]_  = A166 & A167;
  assign \new_[18863]_  = ~A201 & ~A200;
  assign \new_[18864]_  = A199 & \new_[18863]_ ;
  assign \new_[18865]_  = \new_[18864]_  & \new_[18859]_ ;
  assign \new_[18869]_  = ~A267 & A203;
  assign \new_[18870]_  = ~A202 & \new_[18869]_ ;
  assign \new_[18874]_  = A299 & A298;
  assign \new_[18875]_  = ~A269 & \new_[18874]_ ;
  assign \new_[18876]_  = \new_[18875]_  & \new_[18870]_ ;
  assign \new_[18879]_  = A166 & A167;
  assign \new_[18883]_  = ~A201 & ~A200;
  assign \new_[18884]_  = A199 & \new_[18883]_ ;
  assign \new_[18885]_  = \new_[18884]_  & \new_[18879]_ ;
  assign \new_[18889]_  = ~A267 & A203;
  assign \new_[18890]_  = ~A202 & \new_[18889]_ ;
  assign \new_[18894]_  = ~A299 & ~A298;
  assign \new_[18895]_  = ~A269 & \new_[18894]_ ;
  assign \new_[18896]_  = \new_[18895]_  & \new_[18890]_ ;
  assign \new_[18899]_  = A166 & A167;
  assign \new_[18903]_  = ~A201 & ~A200;
  assign \new_[18904]_  = A199 & \new_[18903]_ ;
  assign \new_[18905]_  = \new_[18904]_  & \new_[18899]_ ;
  assign \new_[18909]_  = A265 & A203;
  assign \new_[18910]_  = ~A202 & \new_[18909]_ ;
  assign \new_[18914]_  = A301 & ~A300;
  assign \new_[18915]_  = A266 & \new_[18914]_ ;
  assign \new_[18916]_  = \new_[18915]_  & \new_[18910]_ ;
  assign \new_[18919]_  = A166 & A167;
  assign \new_[18923]_  = ~A201 & ~A200;
  assign \new_[18924]_  = A199 & \new_[18923]_ ;
  assign \new_[18925]_  = \new_[18924]_  & \new_[18919]_ ;
  assign \new_[18929]_  = A265 & A203;
  assign \new_[18930]_  = ~A202 & \new_[18929]_ ;
  assign \new_[18934]_  = ~A302 & ~A300;
  assign \new_[18935]_  = A266 & \new_[18934]_ ;
  assign \new_[18936]_  = \new_[18935]_  & \new_[18930]_ ;
  assign \new_[18939]_  = A166 & A167;
  assign \new_[18943]_  = ~A201 & ~A200;
  assign \new_[18944]_  = A199 & \new_[18943]_ ;
  assign \new_[18945]_  = \new_[18944]_  & \new_[18939]_ ;
  assign \new_[18949]_  = A265 & A203;
  assign \new_[18950]_  = ~A202 & \new_[18949]_ ;
  assign \new_[18954]_  = A299 & A298;
  assign \new_[18955]_  = A266 & \new_[18954]_ ;
  assign \new_[18956]_  = \new_[18955]_  & \new_[18950]_ ;
  assign \new_[18959]_  = A166 & A167;
  assign \new_[18963]_  = ~A201 & ~A200;
  assign \new_[18964]_  = A199 & \new_[18963]_ ;
  assign \new_[18965]_  = \new_[18964]_  & \new_[18959]_ ;
  assign \new_[18969]_  = A265 & A203;
  assign \new_[18970]_  = ~A202 & \new_[18969]_ ;
  assign \new_[18974]_  = ~A299 & ~A298;
  assign \new_[18975]_  = A266 & \new_[18974]_ ;
  assign \new_[18976]_  = \new_[18975]_  & \new_[18970]_ ;
  assign \new_[18979]_  = A166 & A167;
  assign \new_[18983]_  = ~A201 & ~A200;
  assign \new_[18984]_  = A199 & \new_[18983]_ ;
  assign \new_[18985]_  = \new_[18984]_  & \new_[18979]_ ;
  assign \new_[18989]_  = ~A265 & A203;
  assign \new_[18990]_  = ~A202 & \new_[18989]_ ;
  assign \new_[18994]_  = A301 & ~A300;
  assign \new_[18995]_  = ~A266 & \new_[18994]_ ;
  assign \new_[18996]_  = \new_[18995]_  & \new_[18990]_ ;
  assign \new_[18999]_  = A166 & A167;
  assign \new_[19003]_  = ~A201 & ~A200;
  assign \new_[19004]_  = A199 & \new_[19003]_ ;
  assign \new_[19005]_  = \new_[19004]_  & \new_[18999]_ ;
  assign \new_[19009]_  = ~A265 & A203;
  assign \new_[19010]_  = ~A202 & \new_[19009]_ ;
  assign \new_[19014]_  = ~A302 & ~A300;
  assign \new_[19015]_  = ~A266 & \new_[19014]_ ;
  assign \new_[19016]_  = \new_[19015]_  & \new_[19010]_ ;
  assign \new_[19019]_  = A166 & A167;
  assign \new_[19023]_  = ~A201 & ~A200;
  assign \new_[19024]_  = A199 & \new_[19023]_ ;
  assign \new_[19025]_  = \new_[19024]_  & \new_[19019]_ ;
  assign \new_[19029]_  = ~A265 & A203;
  assign \new_[19030]_  = ~A202 & \new_[19029]_ ;
  assign \new_[19034]_  = A299 & A298;
  assign \new_[19035]_  = ~A266 & \new_[19034]_ ;
  assign \new_[19036]_  = \new_[19035]_  & \new_[19030]_ ;
  assign \new_[19039]_  = A166 & A167;
  assign \new_[19043]_  = ~A201 & ~A200;
  assign \new_[19044]_  = A199 & \new_[19043]_ ;
  assign \new_[19045]_  = \new_[19044]_  & \new_[19039]_ ;
  assign \new_[19049]_  = ~A265 & A203;
  assign \new_[19050]_  = ~A202 & \new_[19049]_ ;
  assign \new_[19054]_  = ~A299 & ~A298;
  assign \new_[19055]_  = ~A266 & \new_[19054]_ ;
  assign \new_[19056]_  = \new_[19055]_  & \new_[19050]_ ;
  assign \new_[19059]_  = ~A166 & ~A167;
  assign \new_[19063]_  = A234 & A233;
  assign \new_[19064]_  = ~A232 & \new_[19063]_ ;
  assign \new_[19065]_  = \new_[19064]_  & \new_[19059]_ ;
  assign \new_[19069]_  = A266 & ~A265;
  assign \new_[19070]_  = A235 & \new_[19069]_ ;
  assign \new_[19074]_  = A269 & ~A268;
  assign \new_[19075]_  = ~A267 & \new_[19074]_ ;
  assign \new_[19076]_  = \new_[19075]_  & \new_[19070]_ ;
  assign \new_[19079]_  = ~A166 & ~A167;
  assign \new_[19083]_  = A234 & A233;
  assign \new_[19084]_  = ~A232 & \new_[19083]_ ;
  assign \new_[19085]_  = \new_[19084]_  & \new_[19079]_ ;
  assign \new_[19089]_  = ~A266 & A265;
  assign \new_[19090]_  = A235 & \new_[19089]_ ;
  assign \new_[19094]_  = A269 & ~A268;
  assign \new_[19095]_  = ~A267 & \new_[19094]_ ;
  assign \new_[19096]_  = \new_[19095]_  & \new_[19090]_ ;
  assign \new_[19099]_  = ~A166 & ~A167;
  assign \new_[19103]_  = A234 & A233;
  assign \new_[19104]_  = ~A232 & \new_[19103]_ ;
  assign \new_[19105]_  = \new_[19104]_  & \new_[19099]_ ;
  assign \new_[19109]_  = A266 & ~A265;
  assign \new_[19110]_  = ~A236 & \new_[19109]_ ;
  assign \new_[19114]_  = A269 & ~A268;
  assign \new_[19115]_  = ~A267 & \new_[19114]_ ;
  assign \new_[19116]_  = \new_[19115]_  & \new_[19110]_ ;
  assign \new_[19119]_  = ~A166 & ~A167;
  assign \new_[19123]_  = A234 & A233;
  assign \new_[19124]_  = ~A232 & \new_[19123]_ ;
  assign \new_[19125]_  = \new_[19124]_  & \new_[19119]_ ;
  assign \new_[19129]_  = ~A266 & A265;
  assign \new_[19130]_  = ~A236 & \new_[19129]_ ;
  assign \new_[19134]_  = A269 & ~A268;
  assign \new_[19135]_  = ~A267 & \new_[19134]_ ;
  assign \new_[19136]_  = \new_[19135]_  & \new_[19130]_ ;
  assign \new_[19139]_  = ~A166 & ~A167;
  assign \new_[19143]_  = A234 & ~A233;
  assign \new_[19144]_  = A232 & \new_[19143]_ ;
  assign \new_[19145]_  = \new_[19144]_  & \new_[19139]_ ;
  assign \new_[19149]_  = A266 & ~A265;
  assign \new_[19150]_  = A235 & \new_[19149]_ ;
  assign \new_[19154]_  = A269 & ~A268;
  assign \new_[19155]_  = ~A267 & \new_[19154]_ ;
  assign \new_[19156]_  = \new_[19155]_  & \new_[19150]_ ;
  assign \new_[19159]_  = ~A166 & ~A167;
  assign \new_[19163]_  = A234 & ~A233;
  assign \new_[19164]_  = A232 & \new_[19163]_ ;
  assign \new_[19165]_  = \new_[19164]_  & \new_[19159]_ ;
  assign \new_[19169]_  = ~A266 & A265;
  assign \new_[19170]_  = A235 & \new_[19169]_ ;
  assign \new_[19174]_  = A269 & ~A268;
  assign \new_[19175]_  = ~A267 & \new_[19174]_ ;
  assign \new_[19176]_  = \new_[19175]_  & \new_[19170]_ ;
  assign \new_[19179]_  = ~A166 & ~A167;
  assign \new_[19183]_  = A234 & ~A233;
  assign \new_[19184]_  = A232 & \new_[19183]_ ;
  assign \new_[19185]_  = \new_[19184]_  & \new_[19179]_ ;
  assign \new_[19189]_  = A266 & ~A265;
  assign \new_[19190]_  = ~A236 & \new_[19189]_ ;
  assign \new_[19194]_  = A269 & ~A268;
  assign \new_[19195]_  = ~A267 & \new_[19194]_ ;
  assign \new_[19196]_  = \new_[19195]_  & \new_[19190]_ ;
  assign \new_[19199]_  = ~A166 & ~A167;
  assign \new_[19203]_  = A234 & ~A233;
  assign \new_[19204]_  = A232 & \new_[19203]_ ;
  assign \new_[19205]_  = \new_[19204]_  & \new_[19199]_ ;
  assign \new_[19209]_  = ~A266 & A265;
  assign \new_[19210]_  = ~A236 & \new_[19209]_ ;
  assign \new_[19214]_  = A269 & ~A268;
  assign \new_[19215]_  = ~A267 & \new_[19214]_ ;
  assign \new_[19216]_  = \new_[19215]_  & \new_[19210]_ ;
  assign \new_[19219]_  = ~A166 & ~A167;
  assign \new_[19223]_  = A201 & A200;
  assign \new_[19224]_  = ~A199 & \new_[19223]_ ;
  assign \new_[19225]_  = \new_[19224]_  & \new_[19219]_ ;
  assign \new_[19229]_  = ~A268 & A267;
  assign \new_[19230]_  = A202 & \new_[19229]_ ;
  assign \new_[19234]_  = A301 & ~A300;
  assign \new_[19235]_  = A269 & \new_[19234]_ ;
  assign \new_[19236]_  = \new_[19235]_  & \new_[19230]_ ;
  assign \new_[19239]_  = ~A166 & ~A167;
  assign \new_[19243]_  = A201 & A200;
  assign \new_[19244]_  = ~A199 & \new_[19243]_ ;
  assign \new_[19245]_  = \new_[19244]_  & \new_[19239]_ ;
  assign \new_[19249]_  = ~A268 & A267;
  assign \new_[19250]_  = A202 & \new_[19249]_ ;
  assign \new_[19254]_  = ~A302 & ~A300;
  assign \new_[19255]_  = A269 & \new_[19254]_ ;
  assign \new_[19256]_  = \new_[19255]_  & \new_[19250]_ ;
  assign \new_[19259]_  = ~A166 & ~A167;
  assign \new_[19263]_  = A201 & A200;
  assign \new_[19264]_  = ~A199 & \new_[19263]_ ;
  assign \new_[19265]_  = \new_[19264]_  & \new_[19259]_ ;
  assign \new_[19269]_  = ~A268 & A267;
  assign \new_[19270]_  = A202 & \new_[19269]_ ;
  assign \new_[19274]_  = A299 & A298;
  assign \new_[19275]_  = A269 & \new_[19274]_ ;
  assign \new_[19276]_  = \new_[19275]_  & \new_[19270]_ ;
  assign \new_[19279]_  = ~A166 & ~A167;
  assign \new_[19283]_  = A201 & A200;
  assign \new_[19284]_  = ~A199 & \new_[19283]_ ;
  assign \new_[19285]_  = \new_[19284]_  & \new_[19279]_ ;
  assign \new_[19289]_  = ~A268 & A267;
  assign \new_[19290]_  = A202 & \new_[19289]_ ;
  assign \new_[19294]_  = ~A299 & ~A298;
  assign \new_[19295]_  = A269 & \new_[19294]_ ;
  assign \new_[19296]_  = \new_[19295]_  & \new_[19290]_ ;
  assign \new_[19299]_  = ~A166 & ~A167;
  assign \new_[19303]_  = A201 & A200;
  assign \new_[19304]_  = ~A199 & \new_[19303]_ ;
  assign \new_[19305]_  = \new_[19304]_  & \new_[19299]_ ;
  assign \new_[19309]_  = A268 & ~A267;
  assign \new_[19310]_  = A202 & \new_[19309]_ ;
  assign \new_[19314]_  = A302 & ~A301;
  assign \new_[19315]_  = A300 & \new_[19314]_ ;
  assign \new_[19316]_  = \new_[19315]_  & \new_[19310]_ ;
  assign \new_[19319]_  = ~A166 & ~A167;
  assign \new_[19323]_  = A201 & A200;
  assign \new_[19324]_  = ~A199 & \new_[19323]_ ;
  assign \new_[19325]_  = \new_[19324]_  & \new_[19319]_ ;
  assign \new_[19329]_  = ~A269 & ~A267;
  assign \new_[19330]_  = A202 & \new_[19329]_ ;
  assign \new_[19334]_  = A302 & ~A301;
  assign \new_[19335]_  = A300 & \new_[19334]_ ;
  assign \new_[19336]_  = \new_[19335]_  & \new_[19330]_ ;
  assign \new_[19339]_  = ~A166 & ~A167;
  assign \new_[19343]_  = A201 & A200;
  assign \new_[19344]_  = ~A199 & \new_[19343]_ ;
  assign \new_[19345]_  = \new_[19344]_  & \new_[19339]_ ;
  assign \new_[19349]_  = A266 & A265;
  assign \new_[19350]_  = A202 & \new_[19349]_ ;
  assign \new_[19354]_  = A302 & ~A301;
  assign \new_[19355]_  = A300 & \new_[19354]_ ;
  assign \new_[19356]_  = \new_[19355]_  & \new_[19350]_ ;
  assign \new_[19359]_  = ~A166 & ~A167;
  assign \new_[19363]_  = A201 & A200;
  assign \new_[19364]_  = ~A199 & \new_[19363]_ ;
  assign \new_[19365]_  = \new_[19364]_  & \new_[19359]_ ;
  assign \new_[19369]_  = ~A266 & ~A265;
  assign \new_[19370]_  = A202 & \new_[19369]_ ;
  assign \new_[19374]_  = A302 & ~A301;
  assign \new_[19375]_  = A300 & \new_[19374]_ ;
  assign \new_[19376]_  = \new_[19375]_  & \new_[19370]_ ;
  assign \new_[19379]_  = ~A166 & ~A167;
  assign \new_[19383]_  = A201 & A200;
  assign \new_[19384]_  = ~A199 & \new_[19383]_ ;
  assign \new_[19385]_  = \new_[19384]_  & \new_[19379]_ ;
  assign \new_[19389]_  = ~A268 & A267;
  assign \new_[19390]_  = ~A203 & \new_[19389]_ ;
  assign \new_[19394]_  = A301 & ~A300;
  assign \new_[19395]_  = A269 & \new_[19394]_ ;
  assign \new_[19396]_  = \new_[19395]_  & \new_[19390]_ ;
  assign \new_[19399]_  = ~A166 & ~A167;
  assign \new_[19403]_  = A201 & A200;
  assign \new_[19404]_  = ~A199 & \new_[19403]_ ;
  assign \new_[19405]_  = \new_[19404]_  & \new_[19399]_ ;
  assign \new_[19409]_  = ~A268 & A267;
  assign \new_[19410]_  = ~A203 & \new_[19409]_ ;
  assign \new_[19414]_  = ~A302 & ~A300;
  assign \new_[19415]_  = A269 & \new_[19414]_ ;
  assign \new_[19416]_  = \new_[19415]_  & \new_[19410]_ ;
  assign \new_[19419]_  = ~A166 & ~A167;
  assign \new_[19423]_  = A201 & A200;
  assign \new_[19424]_  = ~A199 & \new_[19423]_ ;
  assign \new_[19425]_  = \new_[19424]_  & \new_[19419]_ ;
  assign \new_[19429]_  = ~A268 & A267;
  assign \new_[19430]_  = ~A203 & \new_[19429]_ ;
  assign \new_[19434]_  = A299 & A298;
  assign \new_[19435]_  = A269 & \new_[19434]_ ;
  assign \new_[19436]_  = \new_[19435]_  & \new_[19430]_ ;
  assign \new_[19439]_  = ~A166 & ~A167;
  assign \new_[19443]_  = A201 & A200;
  assign \new_[19444]_  = ~A199 & \new_[19443]_ ;
  assign \new_[19445]_  = \new_[19444]_  & \new_[19439]_ ;
  assign \new_[19449]_  = ~A268 & A267;
  assign \new_[19450]_  = ~A203 & \new_[19449]_ ;
  assign \new_[19454]_  = ~A299 & ~A298;
  assign \new_[19455]_  = A269 & \new_[19454]_ ;
  assign \new_[19456]_  = \new_[19455]_  & \new_[19450]_ ;
  assign \new_[19459]_  = ~A166 & ~A167;
  assign \new_[19463]_  = A201 & A200;
  assign \new_[19464]_  = ~A199 & \new_[19463]_ ;
  assign \new_[19465]_  = \new_[19464]_  & \new_[19459]_ ;
  assign \new_[19469]_  = A268 & ~A267;
  assign \new_[19470]_  = ~A203 & \new_[19469]_ ;
  assign \new_[19474]_  = A302 & ~A301;
  assign \new_[19475]_  = A300 & \new_[19474]_ ;
  assign \new_[19476]_  = \new_[19475]_  & \new_[19470]_ ;
  assign \new_[19479]_  = ~A166 & ~A167;
  assign \new_[19483]_  = A201 & A200;
  assign \new_[19484]_  = ~A199 & \new_[19483]_ ;
  assign \new_[19485]_  = \new_[19484]_  & \new_[19479]_ ;
  assign \new_[19489]_  = ~A269 & ~A267;
  assign \new_[19490]_  = ~A203 & \new_[19489]_ ;
  assign \new_[19494]_  = A302 & ~A301;
  assign \new_[19495]_  = A300 & \new_[19494]_ ;
  assign \new_[19496]_  = \new_[19495]_  & \new_[19490]_ ;
  assign \new_[19499]_  = ~A166 & ~A167;
  assign \new_[19503]_  = A201 & A200;
  assign \new_[19504]_  = ~A199 & \new_[19503]_ ;
  assign \new_[19505]_  = \new_[19504]_  & \new_[19499]_ ;
  assign \new_[19509]_  = A266 & A265;
  assign \new_[19510]_  = ~A203 & \new_[19509]_ ;
  assign \new_[19514]_  = A302 & ~A301;
  assign \new_[19515]_  = A300 & \new_[19514]_ ;
  assign \new_[19516]_  = \new_[19515]_  & \new_[19510]_ ;
  assign \new_[19519]_  = ~A166 & ~A167;
  assign \new_[19523]_  = A201 & A200;
  assign \new_[19524]_  = ~A199 & \new_[19523]_ ;
  assign \new_[19525]_  = \new_[19524]_  & \new_[19519]_ ;
  assign \new_[19529]_  = ~A266 & ~A265;
  assign \new_[19530]_  = ~A203 & \new_[19529]_ ;
  assign \new_[19534]_  = A302 & ~A301;
  assign \new_[19535]_  = A300 & \new_[19534]_ ;
  assign \new_[19536]_  = \new_[19535]_  & \new_[19530]_ ;
  assign \new_[19539]_  = ~A166 & ~A167;
  assign \new_[19543]_  = ~A201 & A200;
  assign \new_[19544]_  = ~A199 & \new_[19543]_ ;
  assign \new_[19545]_  = \new_[19544]_  & \new_[19539]_ ;
  assign \new_[19549]_  = ~A267 & A203;
  assign \new_[19550]_  = ~A202 & \new_[19549]_ ;
  assign \new_[19554]_  = A301 & ~A300;
  assign \new_[19555]_  = A268 & \new_[19554]_ ;
  assign \new_[19556]_  = \new_[19555]_  & \new_[19550]_ ;
  assign \new_[19559]_  = ~A166 & ~A167;
  assign \new_[19563]_  = ~A201 & A200;
  assign \new_[19564]_  = ~A199 & \new_[19563]_ ;
  assign \new_[19565]_  = \new_[19564]_  & \new_[19559]_ ;
  assign \new_[19569]_  = ~A267 & A203;
  assign \new_[19570]_  = ~A202 & \new_[19569]_ ;
  assign \new_[19574]_  = ~A302 & ~A300;
  assign \new_[19575]_  = A268 & \new_[19574]_ ;
  assign \new_[19576]_  = \new_[19575]_  & \new_[19570]_ ;
  assign \new_[19579]_  = ~A166 & ~A167;
  assign \new_[19583]_  = ~A201 & A200;
  assign \new_[19584]_  = ~A199 & \new_[19583]_ ;
  assign \new_[19585]_  = \new_[19584]_  & \new_[19579]_ ;
  assign \new_[19589]_  = ~A267 & A203;
  assign \new_[19590]_  = ~A202 & \new_[19589]_ ;
  assign \new_[19594]_  = A299 & A298;
  assign \new_[19595]_  = A268 & \new_[19594]_ ;
  assign \new_[19596]_  = \new_[19595]_  & \new_[19590]_ ;
  assign \new_[19599]_  = ~A166 & ~A167;
  assign \new_[19603]_  = ~A201 & A200;
  assign \new_[19604]_  = ~A199 & \new_[19603]_ ;
  assign \new_[19605]_  = \new_[19604]_  & \new_[19599]_ ;
  assign \new_[19609]_  = ~A267 & A203;
  assign \new_[19610]_  = ~A202 & \new_[19609]_ ;
  assign \new_[19614]_  = ~A299 & ~A298;
  assign \new_[19615]_  = A268 & \new_[19614]_ ;
  assign \new_[19616]_  = \new_[19615]_  & \new_[19610]_ ;
  assign \new_[19619]_  = ~A166 & ~A167;
  assign \new_[19623]_  = ~A201 & A200;
  assign \new_[19624]_  = ~A199 & \new_[19623]_ ;
  assign \new_[19625]_  = \new_[19624]_  & \new_[19619]_ ;
  assign \new_[19629]_  = ~A267 & A203;
  assign \new_[19630]_  = ~A202 & \new_[19629]_ ;
  assign \new_[19634]_  = A301 & ~A300;
  assign \new_[19635]_  = ~A269 & \new_[19634]_ ;
  assign \new_[19636]_  = \new_[19635]_  & \new_[19630]_ ;
  assign \new_[19639]_  = ~A166 & ~A167;
  assign \new_[19643]_  = ~A201 & A200;
  assign \new_[19644]_  = ~A199 & \new_[19643]_ ;
  assign \new_[19645]_  = \new_[19644]_  & \new_[19639]_ ;
  assign \new_[19649]_  = ~A267 & A203;
  assign \new_[19650]_  = ~A202 & \new_[19649]_ ;
  assign \new_[19654]_  = ~A302 & ~A300;
  assign \new_[19655]_  = ~A269 & \new_[19654]_ ;
  assign \new_[19656]_  = \new_[19655]_  & \new_[19650]_ ;
  assign \new_[19659]_  = ~A166 & ~A167;
  assign \new_[19663]_  = ~A201 & A200;
  assign \new_[19664]_  = ~A199 & \new_[19663]_ ;
  assign \new_[19665]_  = \new_[19664]_  & \new_[19659]_ ;
  assign \new_[19669]_  = ~A267 & A203;
  assign \new_[19670]_  = ~A202 & \new_[19669]_ ;
  assign \new_[19674]_  = A299 & A298;
  assign \new_[19675]_  = ~A269 & \new_[19674]_ ;
  assign \new_[19676]_  = \new_[19675]_  & \new_[19670]_ ;
  assign \new_[19679]_  = ~A166 & ~A167;
  assign \new_[19683]_  = ~A201 & A200;
  assign \new_[19684]_  = ~A199 & \new_[19683]_ ;
  assign \new_[19685]_  = \new_[19684]_  & \new_[19679]_ ;
  assign \new_[19689]_  = ~A267 & A203;
  assign \new_[19690]_  = ~A202 & \new_[19689]_ ;
  assign \new_[19694]_  = ~A299 & ~A298;
  assign \new_[19695]_  = ~A269 & \new_[19694]_ ;
  assign \new_[19696]_  = \new_[19695]_  & \new_[19690]_ ;
  assign \new_[19699]_  = ~A166 & ~A167;
  assign \new_[19703]_  = ~A201 & A200;
  assign \new_[19704]_  = ~A199 & \new_[19703]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19699]_ ;
  assign \new_[19709]_  = A265 & A203;
  assign \new_[19710]_  = ~A202 & \new_[19709]_ ;
  assign \new_[19714]_  = A301 & ~A300;
  assign \new_[19715]_  = A266 & \new_[19714]_ ;
  assign \new_[19716]_  = \new_[19715]_  & \new_[19710]_ ;
  assign \new_[19719]_  = ~A166 & ~A167;
  assign \new_[19723]_  = ~A201 & A200;
  assign \new_[19724]_  = ~A199 & \new_[19723]_ ;
  assign \new_[19725]_  = \new_[19724]_  & \new_[19719]_ ;
  assign \new_[19729]_  = A265 & A203;
  assign \new_[19730]_  = ~A202 & \new_[19729]_ ;
  assign \new_[19734]_  = ~A302 & ~A300;
  assign \new_[19735]_  = A266 & \new_[19734]_ ;
  assign \new_[19736]_  = \new_[19735]_  & \new_[19730]_ ;
  assign \new_[19739]_  = ~A166 & ~A167;
  assign \new_[19743]_  = ~A201 & A200;
  assign \new_[19744]_  = ~A199 & \new_[19743]_ ;
  assign \new_[19745]_  = \new_[19744]_  & \new_[19739]_ ;
  assign \new_[19749]_  = A265 & A203;
  assign \new_[19750]_  = ~A202 & \new_[19749]_ ;
  assign \new_[19754]_  = A299 & A298;
  assign \new_[19755]_  = A266 & \new_[19754]_ ;
  assign \new_[19756]_  = \new_[19755]_  & \new_[19750]_ ;
  assign \new_[19759]_  = ~A166 & ~A167;
  assign \new_[19763]_  = ~A201 & A200;
  assign \new_[19764]_  = ~A199 & \new_[19763]_ ;
  assign \new_[19765]_  = \new_[19764]_  & \new_[19759]_ ;
  assign \new_[19769]_  = A265 & A203;
  assign \new_[19770]_  = ~A202 & \new_[19769]_ ;
  assign \new_[19774]_  = ~A299 & ~A298;
  assign \new_[19775]_  = A266 & \new_[19774]_ ;
  assign \new_[19776]_  = \new_[19775]_  & \new_[19770]_ ;
  assign \new_[19779]_  = ~A166 & ~A167;
  assign \new_[19783]_  = ~A201 & A200;
  assign \new_[19784]_  = ~A199 & \new_[19783]_ ;
  assign \new_[19785]_  = \new_[19784]_  & \new_[19779]_ ;
  assign \new_[19789]_  = ~A265 & A203;
  assign \new_[19790]_  = ~A202 & \new_[19789]_ ;
  assign \new_[19794]_  = A301 & ~A300;
  assign \new_[19795]_  = ~A266 & \new_[19794]_ ;
  assign \new_[19796]_  = \new_[19795]_  & \new_[19790]_ ;
  assign \new_[19799]_  = ~A166 & ~A167;
  assign \new_[19803]_  = ~A201 & A200;
  assign \new_[19804]_  = ~A199 & \new_[19803]_ ;
  assign \new_[19805]_  = \new_[19804]_  & \new_[19799]_ ;
  assign \new_[19809]_  = ~A265 & A203;
  assign \new_[19810]_  = ~A202 & \new_[19809]_ ;
  assign \new_[19814]_  = ~A302 & ~A300;
  assign \new_[19815]_  = ~A266 & \new_[19814]_ ;
  assign \new_[19816]_  = \new_[19815]_  & \new_[19810]_ ;
  assign \new_[19819]_  = ~A166 & ~A167;
  assign \new_[19823]_  = ~A201 & A200;
  assign \new_[19824]_  = ~A199 & \new_[19823]_ ;
  assign \new_[19825]_  = \new_[19824]_  & \new_[19819]_ ;
  assign \new_[19829]_  = ~A265 & A203;
  assign \new_[19830]_  = ~A202 & \new_[19829]_ ;
  assign \new_[19834]_  = A299 & A298;
  assign \new_[19835]_  = ~A266 & \new_[19834]_ ;
  assign \new_[19836]_  = \new_[19835]_  & \new_[19830]_ ;
  assign \new_[19839]_  = ~A166 & ~A167;
  assign \new_[19843]_  = ~A201 & A200;
  assign \new_[19844]_  = ~A199 & \new_[19843]_ ;
  assign \new_[19845]_  = \new_[19844]_  & \new_[19839]_ ;
  assign \new_[19849]_  = ~A265 & A203;
  assign \new_[19850]_  = ~A202 & \new_[19849]_ ;
  assign \new_[19854]_  = ~A299 & ~A298;
  assign \new_[19855]_  = ~A266 & \new_[19854]_ ;
  assign \new_[19856]_  = \new_[19855]_  & \new_[19850]_ ;
  assign \new_[19859]_  = ~A166 & ~A167;
  assign \new_[19863]_  = A201 & ~A200;
  assign \new_[19864]_  = A199 & \new_[19863]_ ;
  assign \new_[19865]_  = \new_[19864]_  & \new_[19859]_ ;
  assign \new_[19869]_  = ~A268 & A267;
  assign \new_[19870]_  = A202 & \new_[19869]_ ;
  assign \new_[19874]_  = A301 & ~A300;
  assign \new_[19875]_  = A269 & \new_[19874]_ ;
  assign \new_[19876]_  = \new_[19875]_  & \new_[19870]_ ;
  assign \new_[19879]_  = ~A166 & ~A167;
  assign \new_[19883]_  = A201 & ~A200;
  assign \new_[19884]_  = A199 & \new_[19883]_ ;
  assign \new_[19885]_  = \new_[19884]_  & \new_[19879]_ ;
  assign \new_[19889]_  = ~A268 & A267;
  assign \new_[19890]_  = A202 & \new_[19889]_ ;
  assign \new_[19894]_  = ~A302 & ~A300;
  assign \new_[19895]_  = A269 & \new_[19894]_ ;
  assign \new_[19896]_  = \new_[19895]_  & \new_[19890]_ ;
  assign \new_[19899]_  = ~A166 & ~A167;
  assign \new_[19903]_  = A201 & ~A200;
  assign \new_[19904]_  = A199 & \new_[19903]_ ;
  assign \new_[19905]_  = \new_[19904]_  & \new_[19899]_ ;
  assign \new_[19909]_  = ~A268 & A267;
  assign \new_[19910]_  = A202 & \new_[19909]_ ;
  assign \new_[19914]_  = A299 & A298;
  assign \new_[19915]_  = A269 & \new_[19914]_ ;
  assign \new_[19916]_  = \new_[19915]_  & \new_[19910]_ ;
  assign \new_[19919]_  = ~A166 & ~A167;
  assign \new_[19923]_  = A201 & ~A200;
  assign \new_[19924]_  = A199 & \new_[19923]_ ;
  assign \new_[19925]_  = \new_[19924]_  & \new_[19919]_ ;
  assign \new_[19929]_  = ~A268 & A267;
  assign \new_[19930]_  = A202 & \new_[19929]_ ;
  assign \new_[19934]_  = ~A299 & ~A298;
  assign \new_[19935]_  = A269 & \new_[19934]_ ;
  assign \new_[19936]_  = \new_[19935]_  & \new_[19930]_ ;
  assign \new_[19939]_  = ~A166 & ~A167;
  assign \new_[19943]_  = A201 & ~A200;
  assign \new_[19944]_  = A199 & \new_[19943]_ ;
  assign \new_[19945]_  = \new_[19944]_  & \new_[19939]_ ;
  assign \new_[19949]_  = A268 & ~A267;
  assign \new_[19950]_  = A202 & \new_[19949]_ ;
  assign \new_[19954]_  = A302 & ~A301;
  assign \new_[19955]_  = A300 & \new_[19954]_ ;
  assign \new_[19956]_  = \new_[19955]_  & \new_[19950]_ ;
  assign \new_[19959]_  = ~A166 & ~A167;
  assign \new_[19963]_  = A201 & ~A200;
  assign \new_[19964]_  = A199 & \new_[19963]_ ;
  assign \new_[19965]_  = \new_[19964]_  & \new_[19959]_ ;
  assign \new_[19969]_  = ~A269 & ~A267;
  assign \new_[19970]_  = A202 & \new_[19969]_ ;
  assign \new_[19974]_  = A302 & ~A301;
  assign \new_[19975]_  = A300 & \new_[19974]_ ;
  assign \new_[19976]_  = \new_[19975]_  & \new_[19970]_ ;
  assign \new_[19979]_  = ~A166 & ~A167;
  assign \new_[19983]_  = A201 & ~A200;
  assign \new_[19984]_  = A199 & \new_[19983]_ ;
  assign \new_[19985]_  = \new_[19984]_  & \new_[19979]_ ;
  assign \new_[19989]_  = A266 & A265;
  assign \new_[19990]_  = A202 & \new_[19989]_ ;
  assign \new_[19994]_  = A302 & ~A301;
  assign \new_[19995]_  = A300 & \new_[19994]_ ;
  assign \new_[19996]_  = \new_[19995]_  & \new_[19990]_ ;
  assign \new_[19999]_  = ~A166 & ~A167;
  assign \new_[20003]_  = A201 & ~A200;
  assign \new_[20004]_  = A199 & \new_[20003]_ ;
  assign \new_[20005]_  = \new_[20004]_  & \new_[19999]_ ;
  assign \new_[20009]_  = ~A266 & ~A265;
  assign \new_[20010]_  = A202 & \new_[20009]_ ;
  assign \new_[20014]_  = A302 & ~A301;
  assign \new_[20015]_  = A300 & \new_[20014]_ ;
  assign \new_[20016]_  = \new_[20015]_  & \new_[20010]_ ;
  assign \new_[20019]_  = ~A166 & ~A167;
  assign \new_[20023]_  = A201 & ~A200;
  assign \new_[20024]_  = A199 & \new_[20023]_ ;
  assign \new_[20025]_  = \new_[20024]_  & \new_[20019]_ ;
  assign \new_[20029]_  = ~A268 & A267;
  assign \new_[20030]_  = ~A203 & \new_[20029]_ ;
  assign \new_[20034]_  = A301 & ~A300;
  assign \new_[20035]_  = A269 & \new_[20034]_ ;
  assign \new_[20036]_  = \new_[20035]_  & \new_[20030]_ ;
  assign \new_[20039]_  = ~A166 & ~A167;
  assign \new_[20043]_  = A201 & ~A200;
  assign \new_[20044]_  = A199 & \new_[20043]_ ;
  assign \new_[20045]_  = \new_[20044]_  & \new_[20039]_ ;
  assign \new_[20049]_  = ~A268 & A267;
  assign \new_[20050]_  = ~A203 & \new_[20049]_ ;
  assign \new_[20054]_  = ~A302 & ~A300;
  assign \new_[20055]_  = A269 & \new_[20054]_ ;
  assign \new_[20056]_  = \new_[20055]_  & \new_[20050]_ ;
  assign \new_[20059]_  = ~A166 & ~A167;
  assign \new_[20063]_  = A201 & ~A200;
  assign \new_[20064]_  = A199 & \new_[20063]_ ;
  assign \new_[20065]_  = \new_[20064]_  & \new_[20059]_ ;
  assign \new_[20069]_  = ~A268 & A267;
  assign \new_[20070]_  = ~A203 & \new_[20069]_ ;
  assign \new_[20074]_  = A299 & A298;
  assign \new_[20075]_  = A269 & \new_[20074]_ ;
  assign \new_[20076]_  = \new_[20075]_  & \new_[20070]_ ;
  assign \new_[20079]_  = ~A166 & ~A167;
  assign \new_[20083]_  = A201 & ~A200;
  assign \new_[20084]_  = A199 & \new_[20083]_ ;
  assign \new_[20085]_  = \new_[20084]_  & \new_[20079]_ ;
  assign \new_[20089]_  = ~A268 & A267;
  assign \new_[20090]_  = ~A203 & \new_[20089]_ ;
  assign \new_[20094]_  = ~A299 & ~A298;
  assign \new_[20095]_  = A269 & \new_[20094]_ ;
  assign \new_[20096]_  = \new_[20095]_  & \new_[20090]_ ;
  assign \new_[20099]_  = ~A166 & ~A167;
  assign \new_[20103]_  = A201 & ~A200;
  assign \new_[20104]_  = A199 & \new_[20103]_ ;
  assign \new_[20105]_  = \new_[20104]_  & \new_[20099]_ ;
  assign \new_[20109]_  = A268 & ~A267;
  assign \new_[20110]_  = ~A203 & \new_[20109]_ ;
  assign \new_[20114]_  = A302 & ~A301;
  assign \new_[20115]_  = A300 & \new_[20114]_ ;
  assign \new_[20116]_  = \new_[20115]_  & \new_[20110]_ ;
  assign \new_[20119]_  = ~A166 & ~A167;
  assign \new_[20123]_  = A201 & ~A200;
  assign \new_[20124]_  = A199 & \new_[20123]_ ;
  assign \new_[20125]_  = \new_[20124]_  & \new_[20119]_ ;
  assign \new_[20129]_  = ~A269 & ~A267;
  assign \new_[20130]_  = ~A203 & \new_[20129]_ ;
  assign \new_[20134]_  = A302 & ~A301;
  assign \new_[20135]_  = A300 & \new_[20134]_ ;
  assign \new_[20136]_  = \new_[20135]_  & \new_[20130]_ ;
  assign \new_[20139]_  = ~A166 & ~A167;
  assign \new_[20143]_  = A201 & ~A200;
  assign \new_[20144]_  = A199 & \new_[20143]_ ;
  assign \new_[20145]_  = \new_[20144]_  & \new_[20139]_ ;
  assign \new_[20149]_  = A266 & A265;
  assign \new_[20150]_  = ~A203 & \new_[20149]_ ;
  assign \new_[20154]_  = A302 & ~A301;
  assign \new_[20155]_  = A300 & \new_[20154]_ ;
  assign \new_[20156]_  = \new_[20155]_  & \new_[20150]_ ;
  assign \new_[20159]_  = ~A166 & ~A167;
  assign \new_[20163]_  = A201 & ~A200;
  assign \new_[20164]_  = A199 & \new_[20163]_ ;
  assign \new_[20165]_  = \new_[20164]_  & \new_[20159]_ ;
  assign \new_[20169]_  = ~A266 & ~A265;
  assign \new_[20170]_  = ~A203 & \new_[20169]_ ;
  assign \new_[20174]_  = A302 & ~A301;
  assign \new_[20175]_  = A300 & \new_[20174]_ ;
  assign \new_[20176]_  = \new_[20175]_  & \new_[20170]_ ;
  assign \new_[20179]_  = ~A166 & ~A167;
  assign \new_[20183]_  = ~A201 & ~A200;
  assign \new_[20184]_  = A199 & \new_[20183]_ ;
  assign \new_[20185]_  = \new_[20184]_  & \new_[20179]_ ;
  assign \new_[20189]_  = ~A267 & A203;
  assign \new_[20190]_  = ~A202 & \new_[20189]_ ;
  assign \new_[20194]_  = A301 & ~A300;
  assign \new_[20195]_  = A268 & \new_[20194]_ ;
  assign \new_[20196]_  = \new_[20195]_  & \new_[20190]_ ;
  assign \new_[20199]_  = ~A166 & ~A167;
  assign \new_[20203]_  = ~A201 & ~A200;
  assign \new_[20204]_  = A199 & \new_[20203]_ ;
  assign \new_[20205]_  = \new_[20204]_  & \new_[20199]_ ;
  assign \new_[20209]_  = ~A267 & A203;
  assign \new_[20210]_  = ~A202 & \new_[20209]_ ;
  assign \new_[20214]_  = ~A302 & ~A300;
  assign \new_[20215]_  = A268 & \new_[20214]_ ;
  assign \new_[20216]_  = \new_[20215]_  & \new_[20210]_ ;
  assign \new_[20219]_  = ~A166 & ~A167;
  assign \new_[20223]_  = ~A201 & ~A200;
  assign \new_[20224]_  = A199 & \new_[20223]_ ;
  assign \new_[20225]_  = \new_[20224]_  & \new_[20219]_ ;
  assign \new_[20229]_  = ~A267 & A203;
  assign \new_[20230]_  = ~A202 & \new_[20229]_ ;
  assign \new_[20234]_  = A299 & A298;
  assign \new_[20235]_  = A268 & \new_[20234]_ ;
  assign \new_[20236]_  = \new_[20235]_  & \new_[20230]_ ;
  assign \new_[20239]_  = ~A166 & ~A167;
  assign \new_[20243]_  = ~A201 & ~A200;
  assign \new_[20244]_  = A199 & \new_[20243]_ ;
  assign \new_[20245]_  = \new_[20244]_  & \new_[20239]_ ;
  assign \new_[20249]_  = ~A267 & A203;
  assign \new_[20250]_  = ~A202 & \new_[20249]_ ;
  assign \new_[20254]_  = ~A299 & ~A298;
  assign \new_[20255]_  = A268 & \new_[20254]_ ;
  assign \new_[20256]_  = \new_[20255]_  & \new_[20250]_ ;
  assign \new_[20259]_  = ~A166 & ~A167;
  assign \new_[20263]_  = ~A201 & ~A200;
  assign \new_[20264]_  = A199 & \new_[20263]_ ;
  assign \new_[20265]_  = \new_[20264]_  & \new_[20259]_ ;
  assign \new_[20269]_  = ~A267 & A203;
  assign \new_[20270]_  = ~A202 & \new_[20269]_ ;
  assign \new_[20274]_  = A301 & ~A300;
  assign \new_[20275]_  = ~A269 & \new_[20274]_ ;
  assign \new_[20276]_  = \new_[20275]_  & \new_[20270]_ ;
  assign \new_[20279]_  = ~A166 & ~A167;
  assign \new_[20283]_  = ~A201 & ~A200;
  assign \new_[20284]_  = A199 & \new_[20283]_ ;
  assign \new_[20285]_  = \new_[20284]_  & \new_[20279]_ ;
  assign \new_[20289]_  = ~A267 & A203;
  assign \new_[20290]_  = ~A202 & \new_[20289]_ ;
  assign \new_[20294]_  = ~A302 & ~A300;
  assign \new_[20295]_  = ~A269 & \new_[20294]_ ;
  assign \new_[20296]_  = \new_[20295]_  & \new_[20290]_ ;
  assign \new_[20299]_  = ~A166 & ~A167;
  assign \new_[20303]_  = ~A201 & ~A200;
  assign \new_[20304]_  = A199 & \new_[20303]_ ;
  assign \new_[20305]_  = \new_[20304]_  & \new_[20299]_ ;
  assign \new_[20309]_  = ~A267 & A203;
  assign \new_[20310]_  = ~A202 & \new_[20309]_ ;
  assign \new_[20314]_  = A299 & A298;
  assign \new_[20315]_  = ~A269 & \new_[20314]_ ;
  assign \new_[20316]_  = \new_[20315]_  & \new_[20310]_ ;
  assign \new_[20319]_  = ~A166 & ~A167;
  assign \new_[20323]_  = ~A201 & ~A200;
  assign \new_[20324]_  = A199 & \new_[20323]_ ;
  assign \new_[20325]_  = \new_[20324]_  & \new_[20319]_ ;
  assign \new_[20329]_  = ~A267 & A203;
  assign \new_[20330]_  = ~A202 & \new_[20329]_ ;
  assign \new_[20334]_  = ~A299 & ~A298;
  assign \new_[20335]_  = ~A269 & \new_[20334]_ ;
  assign \new_[20336]_  = \new_[20335]_  & \new_[20330]_ ;
  assign \new_[20339]_  = ~A166 & ~A167;
  assign \new_[20343]_  = ~A201 & ~A200;
  assign \new_[20344]_  = A199 & \new_[20343]_ ;
  assign \new_[20345]_  = \new_[20344]_  & \new_[20339]_ ;
  assign \new_[20349]_  = A265 & A203;
  assign \new_[20350]_  = ~A202 & \new_[20349]_ ;
  assign \new_[20354]_  = A301 & ~A300;
  assign \new_[20355]_  = A266 & \new_[20354]_ ;
  assign \new_[20356]_  = \new_[20355]_  & \new_[20350]_ ;
  assign \new_[20359]_  = ~A166 & ~A167;
  assign \new_[20363]_  = ~A201 & ~A200;
  assign \new_[20364]_  = A199 & \new_[20363]_ ;
  assign \new_[20365]_  = \new_[20364]_  & \new_[20359]_ ;
  assign \new_[20369]_  = A265 & A203;
  assign \new_[20370]_  = ~A202 & \new_[20369]_ ;
  assign \new_[20374]_  = ~A302 & ~A300;
  assign \new_[20375]_  = A266 & \new_[20374]_ ;
  assign \new_[20376]_  = \new_[20375]_  & \new_[20370]_ ;
  assign \new_[20379]_  = ~A166 & ~A167;
  assign \new_[20383]_  = ~A201 & ~A200;
  assign \new_[20384]_  = A199 & \new_[20383]_ ;
  assign \new_[20385]_  = \new_[20384]_  & \new_[20379]_ ;
  assign \new_[20389]_  = A265 & A203;
  assign \new_[20390]_  = ~A202 & \new_[20389]_ ;
  assign \new_[20394]_  = A299 & A298;
  assign \new_[20395]_  = A266 & \new_[20394]_ ;
  assign \new_[20396]_  = \new_[20395]_  & \new_[20390]_ ;
  assign \new_[20399]_  = ~A166 & ~A167;
  assign \new_[20403]_  = ~A201 & ~A200;
  assign \new_[20404]_  = A199 & \new_[20403]_ ;
  assign \new_[20405]_  = \new_[20404]_  & \new_[20399]_ ;
  assign \new_[20409]_  = A265 & A203;
  assign \new_[20410]_  = ~A202 & \new_[20409]_ ;
  assign \new_[20414]_  = ~A299 & ~A298;
  assign \new_[20415]_  = A266 & \new_[20414]_ ;
  assign \new_[20416]_  = \new_[20415]_  & \new_[20410]_ ;
  assign \new_[20419]_  = ~A166 & ~A167;
  assign \new_[20423]_  = ~A201 & ~A200;
  assign \new_[20424]_  = A199 & \new_[20423]_ ;
  assign \new_[20425]_  = \new_[20424]_  & \new_[20419]_ ;
  assign \new_[20429]_  = ~A265 & A203;
  assign \new_[20430]_  = ~A202 & \new_[20429]_ ;
  assign \new_[20434]_  = A301 & ~A300;
  assign \new_[20435]_  = ~A266 & \new_[20434]_ ;
  assign \new_[20436]_  = \new_[20435]_  & \new_[20430]_ ;
  assign \new_[20439]_  = ~A166 & ~A167;
  assign \new_[20443]_  = ~A201 & ~A200;
  assign \new_[20444]_  = A199 & \new_[20443]_ ;
  assign \new_[20445]_  = \new_[20444]_  & \new_[20439]_ ;
  assign \new_[20449]_  = ~A265 & A203;
  assign \new_[20450]_  = ~A202 & \new_[20449]_ ;
  assign \new_[20454]_  = ~A302 & ~A300;
  assign \new_[20455]_  = ~A266 & \new_[20454]_ ;
  assign \new_[20456]_  = \new_[20455]_  & \new_[20450]_ ;
  assign \new_[20459]_  = ~A166 & ~A167;
  assign \new_[20463]_  = ~A201 & ~A200;
  assign \new_[20464]_  = A199 & \new_[20463]_ ;
  assign \new_[20465]_  = \new_[20464]_  & \new_[20459]_ ;
  assign \new_[20469]_  = ~A265 & A203;
  assign \new_[20470]_  = ~A202 & \new_[20469]_ ;
  assign \new_[20474]_  = A299 & A298;
  assign \new_[20475]_  = ~A266 & \new_[20474]_ ;
  assign \new_[20476]_  = \new_[20475]_  & \new_[20470]_ ;
  assign \new_[20479]_  = ~A166 & ~A167;
  assign \new_[20483]_  = ~A201 & ~A200;
  assign \new_[20484]_  = A199 & \new_[20483]_ ;
  assign \new_[20485]_  = \new_[20484]_  & \new_[20479]_ ;
  assign \new_[20489]_  = ~A265 & A203;
  assign \new_[20490]_  = ~A202 & \new_[20489]_ ;
  assign \new_[20494]_  = ~A299 & ~A298;
  assign \new_[20495]_  = ~A266 & \new_[20494]_ ;
  assign \new_[20496]_  = \new_[20495]_  & \new_[20490]_ ;
  assign \new_[20499]_  = ~A168 & A170;
  assign \new_[20503]_  = A201 & A200;
  assign \new_[20504]_  = ~A199 & \new_[20503]_ ;
  assign \new_[20505]_  = \new_[20504]_  & \new_[20499]_ ;
  assign \new_[20509]_  = ~A268 & A267;
  assign \new_[20510]_  = A202 & \new_[20509]_ ;
  assign \new_[20514]_  = A301 & ~A300;
  assign \new_[20515]_  = A269 & \new_[20514]_ ;
  assign \new_[20516]_  = \new_[20515]_  & \new_[20510]_ ;
  assign \new_[20519]_  = ~A168 & A170;
  assign \new_[20523]_  = A201 & A200;
  assign \new_[20524]_  = ~A199 & \new_[20523]_ ;
  assign \new_[20525]_  = \new_[20524]_  & \new_[20519]_ ;
  assign \new_[20529]_  = ~A268 & A267;
  assign \new_[20530]_  = A202 & \new_[20529]_ ;
  assign \new_[20534]_  = ~A302 & ~A300;
  assign \new_[20535]_  = A269 & \new_[20534]_ ;
  assign \new_[20536]_  = \new_[20535]_  & \new_[20530]_ ;
  assign \new_[20539]_  = ~A168 & A170;
  assign \new_[20543]_  = A201 & A200;
  assign \new_[20544]_  = ~A199 & \new_[20543]_ ;
  assign \new_[20545]_  = \new_[20544]_  & \new_[20539]_ ;
  assign \new_[20549]_  = ~A268 & A267;
  assign \new_[20550]_  = A202 & \new_[20549]_ ;
  assign \new_[20554]_  = A299 & A298;
  assign \new_[20555]_  = A269 & \new_[20554]_ ;
  assign \new_[20556]_  = \new_[20555]_  & \new_[20550]_ ;
  assign \new_[20559]_  = ~A168 & A170;
  assign \new_[20563]_  = A201 & A200;
  assign \new_[20564]_  = ~A199 & \new_[20563]_ ;
  assign \new_[20565]_  = \new_[20564]_  & \new_[20559]_ ;
  assign \new_[20569]_  = ~A268 & A267;
  assign \new_[20570]_  = A202 & \new_[20569]_ ;
  assign \new_[20574]_  = ~A299 & ~A298;
  assign \new_[20575]_  = A269 & \new_[20574]_ ;
  assign \new_[20576]_  = \new_[20575]_  & \new_[20570]_ ;
  assign \new_[20579]_  = ~A168 & A170;
  assign \new_[20583]_  = A201 & A200;
  assign \new_[20584]_  = ~A199 & \new_[20583]_ ;
  assign \new_[20585]_  = \new_[20584]_  & \new_[20579]_ ;
  assign \new_[20589]_  = A268 & ~A267;
  assign \new_[20590]_  = A202 & \new_[20589]_ ;
  assign \new_[20594]_  = A302 & ~A301;
  assign \new_[20595]_  = A300 & \new_[20594]_ ;
  assign \new_[20596]_  = \new_[20595]_  & \new_[20590]_ ;
  assign \new_[20599]_  = ~A168 & A170;
  assign \new_[20603]_  = A201 & A200;
  assign \new_[20604]_  = ~A199 & \new_[20603]_ ;
  assign \new_[20605]_  = \new_[20604]_  & \new_[20599]_ ;
  assign \new_[20609]_  = ~A269 & ~A267;
  assign \new_[20610]_  = A202 & \new_[20609]_ ;
  assign \new_[20614]_  = A302 & ~A301;
  assign \new_[20615]_  = A300 & \new_[20614]_ ;
  assign \new_[20616]_  = \new_[20615]_  & \new_[20610]_ ;
  assign \new_[20619]_  = ~A168 & A170;
  assign \new_[20623]_  = A201 & A200;
  assign \new_[20624]_  = ~A199 & \new_[20623]_ ;
  assign \new_[20625]_  = \new_[20624]_  & \new_[20619]_ ;
  assign \new_[20629]_  = A266 & A265;
  assign \new_[20630]_  = A202 & \new_[20629]_ ;
  assign \new_[20634]_  = A302 & ~A301;
  assign \new_[20635]_  = A300 & \new_[20634]_ ;
  assign \new_[20636]_  = \new_[20635]_  & \new_[20630]_ ;
  assign \new_[20639]_  = ~A168 & A170;
  assign \new_[20643]_  = A201 & A200;
  assign \new_[20644]_  = ~A199 & \new_[20643]_ ;
  assign \new_[20645]_  = \new_[20644]_  & \new_[20639]_ ;
  assign \new_[20649]_  = ~A266 & ~A265;
  assign \new_[20650]_  = A202 & \new_[20649]_ ;
  assign \new_[20654]_  = A302 & ~A301;
  assign \new_[20655]_  = A300 & \new_[20654]_ ;
  assign \new_[20656]_  = \new_[20655]_  & \new_[20650]_ ;
  assign \new_[20659]_  = ~A168 & A170;
  assign \new_[20663]_  = A201 & A200;
  assign \new_[20664]_  = ~A199 & \new_[20663]_ ;
  assign \new_[20665]_  = \new_[20664]_  & \new_[20659]_ ;
  assign \new_[20669]_  = ~A268 & A267;
  assign \new_[20670]_  = ~A203 & \new_[20669]_ ;
  assign \new_[20674]_  = A301 & ~A300;
  assign \new_[20675]_  = A269 & \new_[20674]_ ;
  assign \new_[20676]_  = \new_[20675]_  & \new_[20670]_ ;
  assign \new_[20679]_  = ~A168 & A170;
  assign \new_[20683]_  = A201 & A200;
  assign \new_[20684]_  = ~A199 & \new_[20683]_ ;
  assign \new_[20685]_  = \new_[20684]_  & \new_[20679]_ ;
  assign \new_[20689]_  = ~A268 & A267;
  assign \new_[20690]_  = ~A203 & \new_[20689]_ ;
  assign \new_[20694]_  = ~A302 & ~A300;
  assign \new_[20695]_  = A269 & \new_[20694]_ ;
  assign \new_[20696]_  = \new_[20695]_  & \new_[20690]_ ;
  assign \new_[20699]_  = ~A168 & A170;
  assign \new_[20703]_  = A201 & A200;
  assign \new_[20704]_  = ~A199 & \new_[20703]_ ;
  assign \new_[20705]_  = \new_[20704]_  & \new_[20699]_ ;
  assign \new_[20709]_  = ~A268 & A267;
  assign \new_[20710]_  = ~A203 & \new_[20709]_ ;
  assign \new_[20714]_  = A299 & A298;
  assign \new_[20715]_  = A269 & \new_[20714]_ ;
  assign \new_[20716]_  = \new_[20715]_  & \new_[20710]_ ;
  assign \new_[20719]_  = ~A168 & A170;
  assign \new_[20723]_  = A201 & A200;
  assign \new_[20724]_  = ~A199 & \new_[20723]_ ;
  assign \new_[20725]_  = \new_[20724]_  & \new_[20719]_ ;
  assign \new_[20729]_  = ~A268 & A267;
  assign \new_[20730]_  = ~A203 & \new_[20729]_ ;
  assign \new_[20734]_  = ~A299 & ~A298;
  assign \new_[20735]_  = A269 & \new_[20734]_ ;
  assign \new_[20736]_  = \new_[20735]_  & \new_[20730]_ ;
  assign \new_[20739]_  = ~A168 & A170;
  assign \new_[20743]_  = A201 & A200;
  assign \new_[20744]_  = ~A199 & \new_[20743]_ ;
  assign \new_[20745]_  = \new_[20744]_  & \new_[20739]_ ;
  assign \new_[20749]_  = A268 & ~A267;
  assign \new_[20750]_  = ~A203 & \new_[20749]_ ;
  assign \new_[20754]_  = A302 & ~A301;
  assign \new_[20755]_  = A300 & \new_[20754]_ ;
  assign \new_[20756]_  = \new_[20755]_  & \new_[20750]_ ;
  assign \new_[20759]_  = ~A168 & A170;
  assign \new_[20763]_  = A201 & A200;
  assign \new_[20764]_  = ~A199 & \new_[20763]_ ;
  assign \new_[20765]_  = \new_[20764]_  & \new_[20759]_ ;
  assign \new_[20769]_  = ~A269 & ~A267;
  assign \new_[20770]_  = ~A203 & \new_[20769]_ ;
  assign \new_[20774]_  = A302 & ~A301;
  assign \new_[20775]_  = A300 & \new_[20774]_ ;
  assign \new_[20776]_  = \new_[20775]_  & \new_[20770]_ ;
  assign \new_[20779]_  = ~A168 & A170;
  assign \new_[20783]_  = A201 & A200;
  assign \new_[20784]_  = ~A199 & \new_[20783]_ ;
  assign \new_[20785]_  = \new_[20784]_  & \new_[20779]_ ;
  assign \new_[20789]_  = A266 & A265;
  assign \new_[20790]_  = ~A203 & \new_[20789]_ ;
  assign \new_[20794]_  = A302 & ~A301;
  assign \new_[20795]_  = A300 & \new_[20794]_ ;
  assign \new_[20796]_  = \new_[20795]_  & \new_[20790]_ ;
  assign \new_[20799]_  = ~A168 & A170;
  assign \new_[20803]_  = A201 & A200;
  assign \new_[20804]_  = ~A199 & \new_[20803]_ ;
  assign \new_[20805]_  = \new_[20804]_  & \new_[20799]_ ;
  assign \new_[20809]_  = ~A266 & ~A265;
  assign \new_[20810]_  = ~A203 & \new_[20809]_ ;
  assign \new_[20814]_  = A302 & ~A301;
  assign \new_[20815]_  = A300 & \new_[20814]_ ;
  assign \new_[20816]_  = \new_[20815]_  & \new_[20810]_ ;
  assign \new_[20819]_  = ~A168 & A170;
  assign \new_[20823]_  = ~A201 & A200;
  assign \new_[20824]_  = ~A199 & \new_[20823]_ ;
  assign \new_[20825]_  = \new_[20824]_  & \new_[20819]_ ;
  assign \new_[20829]_  = ~A267 & A203;
  assign \new_[20830]_  = ~A202 & \new_[20829]_ ;
  assign \new_[20834]_  = A301 & ~A300;
  assign \new_[20835]_  = A268 & \new_[20834]_ ;
  assign \new_[20836]_  = \new_[20835]_  & \new_[20830]_ ;
  assign \new_[20839]_  = ~A168 & A170;
  assign \new_[20843]_  = ~A201 & A200;
  assign \new_[20844]_  = ~A199 & \new_[20843]_ ;
  assign \new_[20845]_  = \new_[20844]_  & \new_[20839]_ ;
  assign \new_[20849]_  = ~A267 & A203;
  assign \new_[20850]_  = ~A202 & \new_[20849]_ ;
  assign \new_[20854]_  = ~A302 & ~A300;
  assign \new_[20855]_  = A268 & \new_[20854]_ ;
  assign \new_[20856]_  = \new_[20855]_  & \new_[20850]_ ;
  assign \new_[20859]_  = ~A168 & A170;
  assign \new_[20863]_  = ~A201 & A200;
  assign \new_[20864]_  = ~A199 & \new_[20863]_ ;
  assign \new_[20865]_  = \new_[20864]_  & \new_[20859]_ ;
  assign \new_[20869]_  = ~A267 & A203;
  assign \new_[20870]_  = ~A202 & \new_[20869]_ ;
  assign \new_[20874]_  = A299 & A298;
  assign \new_[20875]_  = A268 & \new_[20874]_ ;
  assign \new_[20876]_  = \new_[20875]_  & \new_[20870]_ ;
  assign \new_[20879]_  = ~A168 & A170;
  assign \new_[20883]_  = ~A201 & A200;
  assign \new_[20884]_  = ~A199 & \new_[20883]_ ;
  assign \new_[20885]_  = \new_[20884]_  & \new_[20879]_ ;
  assign \new_[20889]_  = ~A267 & A203;
  assign \new_[20890]_  = ~A202 & \new_[20889]_ ;
  assign \new_[20894]_  = ~A299 & ~A298;
  assign \new_[20895]_  = A268 & \new_[20894]_ ;
  assign \new_[20896]_  = \new_[20895]_  & \new_[20890]_ ;
  assign \new_[20899]_  = ~A168 & A170;
  assign \new_[20903]_  = ~A201 & A200;
  assign \new_[20904]_  = ~A199 & \new_[20903]_ ;
  assign \new_[20905]_  = \new_[20904]_  & \new_[20899]_ ;
  assign \new_[20909]_  = ~A267 & A203;
  assign \new_[20910]_  = ~A202 & \new_[20909]_ ;
  assign \new_[20914]_  = A301 & ~A300;
  assign \new_[20915]_  = ~A269 & \new_[20914]_ ;
  assign \new_[20916]_  = \new_[20915]_  & \new_[20910]_ ;
  assign \new_[20919]_  = ~A168 & A170;
  assign \new_[20923]_  = ~A201 & A200;
  assign \new_[20924]_  = ~A199 & \new_[20923]_ ;
  assign \new_[20925]_  = \new_[20924]_  & \new_[20919]_ ;
  assign \new_[20929]_  = ~A267 & A203;
  assign \new_[20930]_  = ~A202 & \new_[20929]_ ;
  assign \new_[20934]_  = ~A302 & ~A300;
  assign \new_[20935]_  = ~A269 & \new_[20934]_ ;
  assign \new_[20936]_  = \new_[20935]_  & \new_[20930]_ ;
  assign \new_[20939]_  = ~A168 & A170;
  assign \new_[20943]_  = ~A201 & A200;
  assign \new_[20944]_  = ~A199 & \new_[20943]_ ;
  assign \new_[20945]_  = \new_[20944]_  & \new_[20939]_ ;
  assign \new_[20949]_  = ~A267 & A203;
  assign \new_[20950]_  = ~A202 & \new_[20949]_ ;
  assign \new_[20954]_  = A299 & A298;
  assign \new_[20955]_  = ~A269 & \new_[20954]_ ;
  assign \new_[20956]_  = \new_[20955]_  & \new_[20950]_ ;
  assign \new_[20959]_  = ~A168 & A170;
  assign \new_[20963]_  = ~A201 & A200;
  assign \new_[20964]_  = ~A199 & \new_[20963]_ ;
  assign \new_[20965]_  = \new_[20964]_  & \new_[20959]_ ;
  assign \new_[20969]_  = ~A267 & A203;
  assign \new_[20970]_  = ~A202 & \new_[20969]_ ;
  assign \new_[20974]_  = ~A299 & ~A298;
  assign \new_[20975]_  = ~A269 & \new_[20974]_ ;
  assign \new_[20976]_  = \new_[20975]_  & \new_[20970]_ ;
  assign \new_[20979]_  = ~A168 & A170;
  assign \new_[20983]_  = ~A201 & A200;
  assign \new_[20984]_  = ~A199 & \new_[20983]_ ;
  assign \new_[20985]_  = \new_[20984]_  & \new_[20979]_ ;
  assign \new_[20989]_  = A265 & A203;
  assign \new_[20990]_  = ~A202 & \new_[20989]_ ;
  assign \new_[20994]_  = A301 & ~A300;
  assign \new_[20995]_  = A266 & \new_[20994]_ ;
  assign \new_[20996]_  = \new_[20995]_  & \new_[20990]_ ;
  assign \new_[20999]_  = ~A168 & A170;
  assign \new_[21003]_  = ~A201 & A200;
  assign \new_[21004]_  = ~A199 & \new_[21003]_ ;
  assign \new_[21005]_  = \new_[21004]_  & \new_[20999]_ ;
  assign \new_[21009]_  = A265 & A203;
  assign \new_[21010]_  = ~A202 & \new_[21009]_ ;
  assign \new_[21014]_  = ~A302 & ~A300;
  assign \new_[21015]_  = A266 & \new_[21014]_ ;
  assign \new_[21016]_  = \new_[21015]_  & \new_[21010]_ ;
  assign \new_[21019]_  = ~A168 & A170;
  assign \new_[21023]_  = ~A201 & A200;
  assign \new_[21024]_  = ~A199 & \new_[21023]_ ;
  assign \new_[21025]_  = \new_[21024]_  & \new_[21019]_ ;
  assign \new_[21029]_  = A265 & A203;
  assign \new_[21030]_  = ~A202 & \new_[21029]_ ;
  assign \new_[21034]_  = A299 & A298;
  assign \new_[21035]_  = A266 & \new_[21034]_ ;
  assign \new_[21036]_  = \new_[21035]_  & \new_[21030]_ ;
  assign \new_[21039]_  = ~A168 & A170;
  assign \new_[21043]_  = ~A201 & A200;
  assign \new_[21044]_  = ~A199 & \new_[21043]_ ;
  assign \new_[21045]_  = \new_[21044]_  & \new_[21039]_ ;
  assign \new_[21049]_  = A265 & A203;
  assign \new_[21050]_  = ~A202 & \new_[21049]_ ;
  assign \new_[21054]_  = ~A299 & ~A298;
  assign \new_[21055]_  = A266 & \new_[21054]_ ;
  assign \new_[21056]_  = \new_[21055]_  & \new_[21050]_ ;
  assign \new_[21059]_  = ~A168 & A170;
  assign \new_[21063]_  = ~A201 & A200;
  assign \new_[21064]_  = ~A199 & \new_[21063]_ ;
  assign \new_[21065]_  = \new_[21064]_  & \new_[21059]_ ;
  assign \new_[21069]_  = ~A265 & A203;
  assign \new_[21070]_  = ~A202 & \new_[21069]_ ;
  assign \new_[21074]_  = A301 & ~A300;
  assign \new_[21075]_  = ~A266 & \new_[21074]_ ;
  assign \new_[21076]_  = \new_[21075]_  & \new_[21070]_ ;
  assign \new_[21079]_  = ~A168 & A170;
  assign \new_[21083]_  = ~A201 & A200;
  assign \new_[21084]_  = ~A199 & \new_[21083]_ ;
  assign \new_[21085]_  = \new_[21084]_  & \new_[21079]_ ;
  assign \new_[21089]_  = ~A265 & A203;
  assign \new_[21090]_  = ~A202 & \new_[21089]_ ;
  assign \new_[21094]_  = ~A302 & ~A300;
  assign \new_[21095]_  = ~A266 & \new_[21094]_ ;
  assign \new_[21096]_  = \new_[21095]_  & \new_[21090]_ ;
  assign \new_[21099]_  = ~A168 & A170;
  assign \new_[21103]_  = ~A201 & A200;
  assign \new_[21104]_  = ~A199 & \new_[21103]_ ;
  assign \new_[21105]_  = \new_[21104]_  & \new_[21099]_ ;
  assign \new_[21109]_  = ~A265 & A203;
  assign \new_[21110]_  = ~A202 & \new_[21109]_ ;
  assign \new_[21114]_  = A299 & A298;
  assign \new_[21115]_  = ~A266 & \new_[21114]_ ;
  assign \new_[21116]_  = \new_[21115]_  & \new_[21110]_ ;
  assign \new_[21119]_  = ~A168 & A170;
  assign \new_[21123]_  = ~A201 & A200;
  assign \new_[21124]_  = ~A199 & \new_[21123]_ ;
  assign \new_[21125]_  = \new_[21124]_  & \new_[21119]_ ;
  assign \new_[21129]_  = ~A265 & A203;
  assign \new_[21130]_  = ~A202 & \new_[21129]_ ;
  assign \new_[21134]_  = ~A299 & ~A298;
  assign \new_[21135]_  = ~A266 & \new_[21134]_ ;
  assign \new_[21136]_  = \new_[21135]_  & \new_[21130]_ ;
  assign \new_[21139]_  = ~A168 & A170;
  assign \new_[21143]_  = A201 & ~A200;
  assign \new_[21144]_  = A199 & \new_[21143]_ ;
  assign \new_[21145]_  = \new_[21144]_  & \new_[21139]_ ;
  assign \new_[21149]_  = ~A268 & A267;
  assign \new_[21150]_  = A202 & \new_[21149]_ ;
  assign \new_[21154]_  = A301 & ~A300;
  assign \new_[21155]_  = A269 & \new_[21154]_ ;
  assign \new_[21156]_  = \new_[21155]_  & \new_[21150]_ ;
  assign \new_[21159]_  = ~A168 & A170;
  assign \new_[21163]_  = A201 & ~A200;
  assign \new_[21164]_  = A199 & \new_[21163]_ ;
  assign \new_[21165]_  = \new_[21164]_  & \new_[21159]_ ;
  assign \new_[21169]_  = ~A268 & A267;
  assign \new_[21170]_  = A202 & \new_[21169]_ ;
  assign \new_[21174]_  = ~A302 & ~A300;
  assign \new_[21175]_  = A269 & \new_[21174]_ ;
  assign \new_[21176]_  = \new_[21175]_  & \new_[21170]_ ;
  assign \new_[21179]_  = ~A168 & A170;
  assign \new_[21183]_  = A201 & ~A200;
  assign \new_[21184]_  = A199 & \new_[21183]_ ;
  assign \new_[21185]_  = \new_[21184]_  & \new_[21179]_ ;
  assign \new_[21189]_  = ~A268 & A267;
  assign \new_[21190]_  = A202 & \new_[21189]_ ;
  assign \new_[21194]_  = A299 & A298;
  assign \new_[21195]_  = A269 & \new_[21194]_ ;
  assign \new_[21196]_  = \new_[21195]_  & \new_[21190]_ ;
  assign \new_[21199]_  = ~A168 & A170;
  assign \new_[21203]_  = A201 & ~A200;
  assign \new_[21204]_  = A199 & \new_[21203]_ ;
  assign \new_[21205]_  = \new_[21204]_  & \new_[21199]_ ;
  assign \new_[21209]_  = ~A268 & A267;
  assign \new_[21210]_  = A202 & \new_[21209]_ ;
  assign \new_[21214]_  = ~A299 & ~A298;
  assign \new_[21215]_  = A269 & \new_[21214]_ ;
  assign \new_[21216]_  = \new_[21215]_  & \new_[21210]_ ;
  assign \new_[21219]_  = ~A168 & A170;
  assign \new_[21223]_  = A201 & ~A200;
  assign \new_[21224]_  = A199 & \new_[21223]_ ;
  assign \new_[21225]_  = \new_[21224]_  & \new_[21219]_ ;
  assign \new_[21229]_  = A268 & ~A267;
  assign \new_[21230]_  = A202 & \new_[21229]_ ;
  assign \new_[21234]_  = A302 & ~A301;
  assign \new_[21235]_  = A300 & \new_[21234]_ ;
  assign \new_[21236]_  = \new_[21235]_  & \new_[21230]_ ;
  assign \new_[21239]_  = ~A168 & A170;
  assign \new_[21243]_  = A201 & ~A200;
  assign \new_[21244]_  = A199 & \new_[21243]_ ;
  assign \new_[21245]_  = \new_[21244]_  & \new_[21239]_ ;
  assign \new_[21249]_  = ~A269 & ~A267;
  assign \new_[21250]_  = A202 & \new_[21249]_ ;
  assign \new_[21254]_  = A302 & ~A301;
  assign \new_[21255]_  = A300 & \new_[21254]_ ;
  assign \new_[21256]_  = \new_[21255]_  & \new_[21250]_ ;
  assign \new_[21259]_  = ~A168 & A170;
  assign \new_[21263]_  = A201 & ~A200;
  assign \new_[21264]_  = A199 & \new_[21263]_ ;
  assign \new_[21265]_  = \new_[21264]_  & \new_[21259]_ ;
  assign \new_[21269]_  = A266 & A265;
  assign \new_[21270]_  = A202 & \new_[21269]_ ;
  assign \new_[21274]_  = A302 & ~A301;
  assign \new_[21275]_  = A300 & \new_[21274]_ ;
  assign \new_[21276]_  = \new_[21275]_  & \new_[21270]_ ;
  assign \new_[21279]_  = ~A168 & A170;
  assign \new_[21283]_  = A201 & ~A200;
  assign \new_[21284]_  = A199 & \new_[21283]_ ;
  assign \new_[21285]_  = \new_[21284]_  & \new_[21279]_ ;
  assign \new_[21289]_  = ~A266 & ~A265;
  assign \new_[21290]_  = A202 & \new_[21289]_ ;
  assign \new_[21294]_  = A302 & ~A301;
  assign \new_[21295]_  = A300 & \new_[21294]_ ;
  assign \new_[21296]_  = \new_[21295]_  & \new_[21290]_ ;
  assign \new_[21299]_  = ~A168 & A170;
  assign \new_[21303]_  = A201 & ~A200;
  assign \new_[21304]_  = A199 & \new_[21303]_ ;
  assign \new_[21305]_  = \new_[21304]_  & \new_[21299]_ ;
  assign \new_[21309]_  = ~A268 & A267;
  assign \new_[21310]_  = ~A203 & \new_[21309]_ ;
  assign \new_[21314]_  = A301 & ~A300;
  assign \new_[21315]_  = A269 & \new_[21314]_ ;
  assign \new_[21316]_  = \new_[21315]_  & \new_[21310]_ ;
  assign \new_[21319]_  = ~A168 & A170;
  assign \new_[21323]_  = A201 & ~A200;
  assign \new_[21324]_  = A199 & \new_[21323]_ ;
  assign \new_[21325]_  = \new_[21324]_  & \new_[21319]_ ;
  assign \new_[21329]_  = ~A268 & A267;
  assign \new_[21330]_  = ~A203 & \new_[21329]_ ;
  assign \new_[21334]_  = ~A302 & ~A300;
  assign \new_[21335]_  = A269 & \new_[21334]_ ;
  assign \new_[21336]_  = \new_[21335]_  & \new_[21330]_ ;
  assign \new_[21339]_  = ~A168 & A170;
  assign \new_[21343]_  = A201 & ~A200;
  assign \new_[21344]_  = A199 & \new_[21343]_ ;
  assign \new_[21345]_  = \new_[21344]_  & \new_[21339]_ ;
  assign \new_[21349]_  = ~A268 & A267;
  assign \new_[21350]_  = ~A203 & \new_[21349]_ ;
  assign \new_[21354]_  = A299 & A298;
  assign \new_[21355]_  = A269 & \new_[21354]_ ;
  assign \new_[21356]_  = \new_[21355]_  & \new_[21350]_ ;
  assign \new_[21359]_  = ~A168 & A170;
  assign \new_[21363]_  = A201 & ~A200;
  assign \new_[21364]_  = A199 & \new_[21363]_ ;
  assign \new_[21365]_  = \new_[21364]_  & \new_[21359]_ ;
  assign \new_[21369]_  = ~A268 & A267;
  assign \new_[21370]_  = ~A203 & \new_[21369]_ ;
  assign \new_[21374]_  = ~A299 & ~A298;
  assign \new_[21375]_  = A269 & \new_[21374]_ ;
  assign \new_[21376]_  = \new_[21375]_  & \new_[21370]_ ;
  assign \new_[21379]_  = ~A168 & A170;
  assign \new_[21383]_  = A201 & ~A200;
  assign \new_[21384]_  = A199 & \new_[21383]_ ;
  assign \new_[21385]_  = \new_[21384]_  & \new_[21379]_ ;
  assign \new_[21389]_  = A268 & ~A267;
  assign \new_[21390]_  = ~A203 & \new_[21389]_ ;
  assign \new_[21394]_  = A302 & ~A301;
  assign \new_[21395]_  = A300 & \new_[21394]_ ;
  assign \new_[21396]_  = \new_[21395]_  & \new_[21390]_ ;
  assign \new_[21399]_  = ~A168 & A170;
  assign \new_[21403]_  = A201 & ~A200;
  assign \new_[21404]_  = A199 & \new_[21403]_ ;
  assign \new_[21405]_  = \new_[21404]_  & \new_[21399]_ ;
  assign \new_[21409]_  = ~A269 & ~A267;
  assign \new_[21410]_  = ~A203 & \new_[21409]_ ;
  assign \new_[21414]_  = A302 & ~A301;
  assign \new_[21415]_  = A300 & \new_[21414]_ ;
  assign \new_[21416]_  = \new_[21415]_  & \new_[21410]_ ;
  assign \new_[21419]_  = ~A168 & A170;
  assign \new_[21423]_  = A201 & ~A200;
  assign \new_[21424]_  = A199 & \new_[21423]_ ;
  assign \new_[21425]_  = \new_[21424]_  & \new_[21419]_ ;
  assign \new_[21429]_  = A266 & A265;
  assign \new_[21430]_  = ~A203 & \new_[21429]_ ;
  assign \new_[21434]_  = A302 & ~A301;
  assign \new_[21435]_  = A300 & \new_[21434]_ ;
  assign \new_[21436]_  = \new_[21435]_  & \new_[21430]_ ;
  assign \new_[21439]_  = ~A168 & A170;
  assign \new_[21443]_  = A201 & ~A200;
  assign \new_[21444]_  = A199 & \new_[21443]_ ;
  assign \new_[21445]_  = \new_[21444]_  & \new_[21439]_ ;
  assign \new_[21449]_  = ~A266 & ~A265;
  assign \new_[21450]_  = ~A203 & \new_[21449]_ ;
  assign \new_[21454]_  = A302 & ~A301;
  assign \new_[21455]_  = A300 & \new_[21454]_ ;
  assign \new_[21456]_  = \new_[21455]_  & \new_[21450]_ ;
  assign \new_[21459]_  = ~A168 & A170;
  assign \new_[21463]_  = ~A201 & ~A200;
  assign \new_[21464]_  = A199 & \new_[21463]_ ;
  assign \new_[21465]_  = \new_[21464]_  & \new_[21459]_ ;
  assign \new_[21469]_  = ~A267 & A203;
  assign \new_[21470]_  = ~A202 & \new_[21469]_ ;
  assign \new_[21474]_  = A301 & ~A300;
  assign \new_[21475]_  = A268 & \new_[21474]_ ;
  assign \new_[21476]_  = \new_[21475]_  & \new_[21470]_ ;
  assign \new_[21479]_  = ~A168 & A170;
  assign \new_[21483]_  = ~A201 & ~A200;
  assign \new_[21484]_  = A199 & \new_[21483]_ ;
  assign \new_[21485]_  = \new_[21484]_  & \new_[21479]_ ;
  assign \new_[21489]_  = ~A267 & A203;
  assign \new_[21490]_  = ~A202 & \new_[21489]_ ;
  assign \new_[21494]_  = ~A302 & ~A300;
  assign \new_[21495]_  = A268 & \new_[21494]_ ;
  assign \new_[21496]_  = \new_[21495]_  & \new_[21490]_ ;
  assign \new_[21499]_  = ~A168 & A170;
  assign \new_[21503]_  = ~A201 & ~A200;
  assign \new_[21504]_  = A199 & \new_[21503]_ ;
  assign \new_[21505]_  = \new_[21504]_  & \new_[21499]_ ;
  assign \new_[21509]_  = ~A267 & A203;
  assign \new_[21510]_  = ~A202 & \new_[21509]_ ;
  assign \new_[21514]_  = A299 & A298;
  assign \new_[21515]_  = A268 & \new_[21514]_ ;
  assign \new_[21516]_  = \new_[21515]_  & \new_[21510]_ ;
  assign \new_[21519]_  = ~A168 & A170;
  assign \new_[21523]_  = ~A201 & ~A200;
  assign \new_[21524]_  = A199 & \new_[21523]_ ;
  assign \new_[21525]_  = \new_[21524]_  & \new_[21519]_ ;
  assign \new_[21529]_  = ~A267 & A203;
  assign \new_[21530]_  = ~A202 & \new_[21529]_ ;
  assign \new_[21534]_  = ~A299 & ~A298;
  assign \new_[21535]_  = A268 & \new_[21534]_ ;
  assign \new_[21536]_  = \new_[21535]_  & \new_[21530]_ ;
  assign \new_[21539]_  = ~A168 & A170;
  assign \new_[21543]_  = ~A201 & ~A200;
  assign \new_[21544]_  = A199 & \new_[21543]_ ;
  assign \new_[21545]_  = \new_[21544]_  & \new_[21539]_ ;
  assign \new_[21549]_  = ~A267 & A203;
  assign \new_[21550]_  = ~A202 & \new_[21549]_ ;
  assign \new_[21554]_  = A301 & ~A300;
  assign \new_[21555]_  = ~A269 & \new_[21554]_ ;
  assign \new_[21556]_  = \new_[21555]_  & \new_[21550]_ ;
  assign \new_[21559]_  = ~A168 & A170;
  assign \new_[21563]_  = ~A201 & ~A200;
  assign \new_[21564]_  = A199 & \new_[21563]_ ;
  assign \new_[21565]_  = \new_[21564]_  & \new_[21559]_ ;
  assign \new_[21569]_  = ~A267 & A203;
  assign \new_[21570]_  = ~A202 & \new_[21569]_ ;
  assign \new_[21574]_  = ~A302 & ~A300;
  assign \new_[21575]_  = ~A269 & \new_[21574]_ ;
  assign \new_[21576]_  = \new_[21575]_  & \new_[21570]_ ;
  assign \new_[21579]_  = ~A168 & A170;
  assign \new_[21583]_  = ~A201 & ~A200;
  assign \new_[21584]_  = A199 & \new_[21583]_ ;
  assign \new_[21585]_  = \new_[21584]_  & \new_[21579]_ ;
  assign \new_[21589]_  = ~A267 & A203;
  assign \new_[21590]_  = ~A202 & \new_[21589]_ ;
  assign \new_[21594]_  = A299 & A298;
  assign \new_[21595]_  = ~A269 & \new_[21594]_ ;
  assign \new_[21596]_  = \new_[21595]_  & \new_[21590]_ ;
  assign \new_[21599]_  = ~A168 & A170;
  assign \new_[21603]_  = ~A201 & ~A200;
  assign \new_[21604]_  = A199 & \new_[21603]_ ;
  assign \new_[21605]_  = \new_[21604]_  & \new_[21599]_ ;
  assign \new_[21609]_  = ~A267 & A203;
  assign \new_[21610]_  = ~A202 & \new_[21609]_ ;
  assign \new_[21614]_  = ~A299 & ~A298;
  assign \new_[21615]_  = ~A269 & \new_[21614]_ ;
  assign \new_[21616]_  = \new_[21615]_  & \new_[21610]_ ;
  assign \new_[21619]_  = ~A168 & A170;
  assign \new_[21623]_  = ~A201 & ~A200;
  assign \new_[21624]_  = A199 & \new_[21623]_ ;
  assign \new_[21625]_  = \new_[21624]_  & \new_[21619]_ ;
  assign \new_[21629]_  = A265 & A203;
  assign \new_[21630]_  = ~A202 & \new_[21629]_ ;
  assign \new_[21634]_  = A301 & ~A300;
  assign \new_[21635]_  = A266 & \new_[21634]_ ;
  assign \new_[21636]_  = \new_[21635]_  & \new_[21630]_ ;
  assign \new_[21639]_  = ~A168 & A170;
  assign \new_[21643]_  = ~A201 & ~A200;
  assign \new_[21644]_  = A199 & \new_[21643]_ ;
  assign \new_[21645]_  = \new_[21644]_  & \new_[21639]_ ;
  assign \new_[21649]_  = A265 & A203;
  assign \new_[21650]_  = ~A202 & \new_[21649]_ ;
  assign \new_[21654]_  = ~A302 & ~A300;
  assign \new_[21655]_  = A266 & \new_[21654]_ ;
  assign \new_[21656]_  = \new_[21655]_  & \new_[21650]_ ;
  assign \new_[21659]_  = ~A168 & A170;
  assign \new_[21663]_  = ~A201 & ~A200;
  assign \new_[21664]_  = A199 & \new_[21663]_ ;
  assign \new_[21665]_  = \new_[21664]_  & \new_[21659]_ ;
  assign \new_[21669]_  = A265 & A203;
  assign \new_[21670]_  = ~A202 & \new_[21669]_ ;
  assign \new_[21674]_  = A299 & A298;
  assign \new_[21675]_  = A266 & \new_[21674]_ ;
  assign \new_[21676]_  = \new_[21675]_  & \new_[21670]_ ;
  assign \new_[21679]_  = ~A168 & A170;
  assign \new_[21683]_  = ~A201 & ~A200;
  assign \new_[21684]_  = A199 & \new_[21683]_ ;
  assign \new_[21685]_  = \new_[21684]_  & \new_[21679]_ ;
  assign \new_[21689]_  = A265 & A203;
  assign \new_[21690]_  = ~A202 & \new_[21689]_ ;
  assign \new_[21694]_  = ~A299 & ~A298;
  assign \new_[21695]_  = A266 & \new_[21694]_ ;
  assign \new_[21696]_  = \new_[21695]_  & \new_[21690]_ ;
  assign \new_[21699]_  = ~A168 & A170;
  assign \new_[21703]_  = ~A201 & ~A200;
  assign \new_[21704]_  = A199 & \new_[21703]_ ;
  assign \new_[21705]_  = \new_[21704]_  & \new_[21699]_ ;
  assign \new_[21709]_  = ~A265 & A203;
  assign \new_[21710]_  = ~A202 & \new_[21709]_ ;
  assign \new_[21714]_  = A301 & ~A300;
  assign \new_[21715]_  = ~A266 & \new_[21714]_ ;
  assign \new_[21716]_  = \new_[21715]_  & \new_[21710]_ ;
  assign \new_[21719]_  = ~A168 & A170;
  assign \new_[21723]_  = ~A201 & ~A200;
  assign \new_[21724]_  = A199 & \new_[21723]_ ;
  assign \new_[21725]_  = \new_[21724]_  & \new_[21719]_ ;
  assign \new_[21729]_  = ~A265 & A203;
  assign \new_[21730]_  = ~A202 & \new_[21729]_ ;
  assign \new_[21734]_  = ~A302 & ~A300;
  assign \new_[21735]_  = ~A266 & \new_[21734]_ ;
  assign \new_[21736]_  = \new_[21735]_  & \new_[21730]_ ;
  assign \new_[21739]_  = ~A168 & A170;
  assign \new_[21743]_  = ~A201 & ~A200;
  assign \new_[21744]_  = A199 & \new_[21743]_ ;
  assign \new_[21745]_  = \new_[21744]_  & \new_[21739]_ ;
  assign \new_[21749]_  = ~A265 & A203;
  assign \new_[21750]_  = ~A202 & \new_[21749]_ ;
  assign \new_[21754]_  = A299 & A298;
  assign \new_[21755]_  = ~A266 & \new_[21754]_ ;
  assign \new_[21756]_  = \new_[21755]_  & \new_[21750]_ ;
  assign \new_[21759]_  = ~A168 & A170;
  assign \new_[21763]_  = ~A201 & ~A200;
  assign \new_[21764]_  = A199 & \new_[21763]_ ;
  assign \new_[21765]_  = \new_[21764]_  & \new_[21759]_ ;
  assign \new_[21769]_  = ~A265 & A203;
  assign \new_[21770]_  = ~A202 & \new_[21769]_ ;
  assign \new_[21774]_  = ~A299 & ~A298;
  assign \new_[21775]_  = ~A266 & \new_[21774]_ ;
  assign \new_[21776]_  = \new_[21775]_  & \new_[21770]_ ;
  assign \new_[21779]_  = ~A168 & A169;
  assign \new_[21783]_  = A201 & A200;
  assign \new_[21784]_  = ~A199 & \new_[21783]_ ;
  assign \new_[21785]_  = \new_[21784]_  & \new_[21779]_ ;
  assign \new_[21789]_  = ~A268 & A267;
  assign \new_[21790]_  = A202 & \new_[21789]_ ;
  assign \new_[21794]_  = A301 & ~A300;
  assign \new_[21795]_  = A269 & \new_[21794]_ ;
  assign \new_[21796]_  = \new_[21795]_  & \new_[21790]_ ;
  assign \new_[21799]_  = ~A168 & A169;
  assign \new_[21803]_  = A201 & A200;
  assign \new_[21804]_  = ~A199 & \new_[21803]_ ;
  assign \new_[21805]_  = \new_[21804]_  & \new_[21799]_ ;
  assign \new_[21809]_  = ~A268 & A267;
  assign \new_[21810]_  = A202 & \new_[21809]_ ;
  assign \new_[21814]_  = ~A302 & ~A300;
  assign \new_[21815]_  = A269 & \new_[21814]_ ;
  assign \new_[21816]_  = \new_[21815]_  & \new_[21810]_ ;
  assign \new_[21819]_  = ~A168 & A169;
  assign \new_[21823]_  = A201 & A200;
  assign \new_[21824]_  = ~A199 & \new_[21823]_ ;
  assign \new_[21825]_  = \new_[21824]_  & \new_[21819]_ ;
  assign \new_[21829]_  = ~A268 & A267;
  assign \new_[21830]_  = A202 & \new_[21829]_ ;
  assign \new_[21834]_  = A299 & A298;
  assign \new_[21835]_  = A269 & \new_[21834]_ ;
  assign \new_[21836]_  = \new_[21835]_  & \new_[21830]_ ;
  assign \new_[21839]_  = ~A168 & A169;
  assign \new_[21843]_  = A201 & A200;
  assign \new_[21844]_  = ~A199 & \new_[21843]_ ;
  assign \new_[21845]_  = \new_[21844]_  & \new_[21839]_ ;
  assign \new_[21849]_  = ~A268 & A267;
  assign \new_[21850]_  = A202 & \new_[21849]_ ;
  assign \new_[21854]_  = ~A299 & ~A298;
  assign \new_[21855]_  = A269 & \new_[21854]_ ;
  assign \new_[21856]_  = \new_[21855]_  & \new_[21850]_ ;
  assign \new_[21859]_  = ~A168 & A169;
  assign \new_[21863]_  = A201 & A200;
  assign \new_[21864]_  = ~A199 & \new_[21863]_ ;
  assign \new_[21865]_  = \new_[21864]_  & \new_[21859]_ ;
  assign \new_[21869]_  = A268 & ~A267;
  assign \new_[21870]_  = A202 & \new_[21869]_ ;
  assign \new_[21874]_  = A302 & ~A301;
  assign \new_[21875]_  = A300 & \new_[21874]_ ;
  assign \new_[21876]_  = \new_[21875]_  & \new_[21870]_ ;
  assign \new_[21879]_  = ~A168 & A169;
  assign \new_[21883]_  = A201 & A200;
  assign \new_[21884]_  = ~A199 & \new_[21883]_ ;
  assign \new_[21885]_  = \new_[21884]_  & \new_[21879]_ ;
  assign \new_[21889]_  = ~A269 & ~A267;
  assign \new_[21890]_  = A202 & \new_[21889]_ ;
  assign \new_[21894]_  = A302 & ~A301;
  assign \new_[21895]_  = A300 & \new_[21894]_ ;
  assign \new_[21896]_  = \new_[21895]_  & \new_[21890]_ ;
  assign \new_[21899]_  = ~A168 & A169;
  assign \new_[21903]_  = A201 & A200;
  assign \new_[21904]_  = ~A199 & \new_[21903]_ ;
  assign \new_[21905]_  = \new_[21904]_  & \new_[21899]_ ;
  assign \new_[21909]_  = A266 & A265;
  assign \new_[21910]_  = A202 & \new_[21909]_ ;
  assign \new_[21914]_  = A302 & ~A301;
  assign \new_[21915]_  = A300 & \new_[21914]_ ;
  assign \new_[21916]_  = \new_[21915]_  & \new_[21910]_ ;
  assign \new_[21919]_  = ~A168 & A169;
  assign \new_[21923]_  = A201 & A200;
  assign \new_[21924]_  = ~A199 & \new_[21923]_ ;
  assign \new_[21925]_  = \new_[21924]_  & \new_[21919]_ ;
  assign \new_[21929]_  = ~A266 & ~A265;
  assign \new_[21930]_  = A202 & \new_[21929]_ ;
  assign \new_[21934]_  = A302 & ~A301;
  assign \new_[21935]_  = A300 & \new_[21934]_ ;
  assign \new_[21936]_  = \new_[21935]_  & \new_[21930]_ ;
  assign \new_[21939]_  = ~A168 & A169;
  assign \new_[21943]_  = A201 & A200;
  assign \new_[21944]_  = ~A199 & \new_[21943]_ ;
  assign \new_[21945]_  = \new_[21944]_  & \new_[21939]_ ;
  assign \new_[21949]_  = ~A268 & A267;
  assign \new_[21950]_  = ~A203 & \new_[21949]_ ;
  assign \new_[21954]_  = A301 & ~A300;
  assign \new_[21955]_  = A269 & \new_[21954]_ ;
  assign \new_[21956]_  = \new_[21955]_  & \new_[21950]_ ;
  assign \new_[21959]_  = ~A168 & A169;
  assign \new_[21963]_  = A201 & A200;
  assign \new_[21964]_  = ~A199 & \new_[21963]_ ;
  assign \new_[21965]_  = \new_[21964]_  & \new_[21959]_ ;
  assign \new_[21969]_  = ~A268 & A267;
  assign \new_[21970]_  = ~A203 & \new_[21969]_ ;
  assign \new_[21974]_  = ~A302 & ~A300;
  assign \new_[21975]_  = A269 & \new_[21974]_ ;
  assign \new_[21976]_  = \new_[21975]_  & \new_[21970]_ ;
  assign \new_[21979]_  = ~A168 & A169;
  assign \new_[21983]_  = A201 & A200;
  assign \new_[21984]_  = ~A199 & \new_[21983]_ ;
  assign \new_[21985]_  = \new_[21984]_  & \new_[21979]_ ;
  assign \new_[21989]_  = ~A268 & A267;
  assign \new_[21990]_  = ~A203 & \new_[21989]_ ;
  assign \new_[21994]_  = A299 & A298;
  assign \new_[21995]_  = A269 & \new_[21994]_ ;
  assign \new_[21996]_  = \new_[21995]_  & \new_[21990]_ ;
  assign \new_[21999]_  = ~A168 & A169;
  assign \new_[22003]_  = A201 & A200;
  assign \new_[22004]_  = ~A199 & \new_[22003]_ ;
  assign \new_[22005]_  = \new_[22004]_  & \new_[21999]_ ;
  assign \new_[22009]_  = ~A268 & A267;
  assign \new_[22010]_  = ~A203 & \new_[22009]_ ;
  assign \new_[22014]_  = ~A299 & ~A298;
  assign \new_[22015]_  = A269 & \new_[22014]_ ;
  assign \new_[22016]_  = \new_[22015]_  & \new_[22010]_ ;
  assign \new_[22019]_  = ~A168 & A169;
  assign \new_[22023]_  = A201 & A200;
  assign \new_[22024]_  = ~A199 & \new_[22023]_ ;
  assign \new_[22025]_  = \new_[22024]_  & \new_[22019]_ ;
  assign \new_[22029]_  = A268 & ~A267;
  assign \new_[22030]_  = ~A203 & \new_[22029]_ ;
  assign \new_[22034]_  = A302 & ~A301;
  assign \new_[22035]_  = A300 & \new_[22034]_ ;
  assign \new_[22036]_  = \new_[22035]_  & \new_[22030]_ ;
  assign \new_[22039]_  = ~A168 & A169;
  assign \new_[22043]_  = A201 & A200;
  assign \new_[22044]_  = ~A199 & \new_[22043]_ ;
  assign \new_[22045]_  = \new_[22044]_  & \new_[22039]_ ;
  assign \new_[22049]_  = ~A269 & ~A267;
  assign \new_[22050]_  = ~A203 & \new_[22049]_ ;
  assign \new_[22054]_  = A302 & ~A301;
  assign \new_[22055]_  = A300 & \new_[22054]_ ;
  assign \new_[22056]_  = \new_[22055]_  & \new_[22050]_ ;
  assign \new_[22059]_  = ~A168 & A169;
  assign \new_[22063]_  = A201 & A200;
  assign \new_[22064]_  = ~A199 & \new_[22063]_ ;
  assign \new_[22065]_  = \new_[22064]_  & \new_[22059]_ ;
  assign \new_[22069]_  = A266 & A265;
  assign \new_[22070]_  = ~A203 & \new_[22069]_ ;
  assign \new_[22074]_  = A302 & ~A301;
  assign \new_[22075]_  = A300 & \new_[22074]_ ;
  assign \new_[22076]_  = \new_[22075]_  & \new_[22070]_ ;
  assign \new_[22079]_  = ~A168 & A169;
  assign \new_[22083]_  = A201 & A200;
  assign \new_[22084]_  = ~A199 & \new_[22083]_ ;
  assign \new_[22085]_  = \new_[22084]_  & \new_[22079]_ ;
  assign \new_[22089]_  = ~A266 & ~A265;
  assign \new_[22090]_  = ~A203 & \new_[22089]_ ;
  assign \new_[22094]_  = A302 & ~A301;
  assign \new_[22095]_  = A300 & \new_[22094]_ ;
  assign \new_[22096]_  = \new_[22095]_  & \new_[22090]_ ;
  assign \new_[22099]_  = ~A168 & A169;
  assign \new_[22103]_  = ~A201 & A200;
  assign \new_[22104]_  = ~A199 & \new_[22103]_ ;
  assign \new_[22105]_  = \new_[22104]_  & \new_[22099]_ ;
  assign \new_[22109]_  = ~A267 & A203;
  assign \new_[22110]_  = ~A202 & \new_[22109]_ ;
  assign \new_[22114]_  = A301 & ~A300;
  assign \new_[22115]_  = A268 & \new_[22114]_ ;
  assign \new_[22116]_  = \new_[22115]_  & \new_[22110]_ ;
  assign \new_[22119]_  = ~A168 & A169;
  assign \new_[22123]_  = ~A201 & A200;
  assign \new_[22124]_  = ~A199 & \new_[22123]_ ;
  assign \new_[22125]_  = \new_[22124]_  & \new_[22119]_ ;
  assign \new_[22129]_  = ~A267 & A203;
  assign \new_[22130]_  = ~A202 & \new_[22129]_ ;
  assign \new_[22134]_  = ~A302 & ~A300;
  assign \new_[22135]_  = A268 & \new_[22134]_ ;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22130]_ ;
  assign \new_[22139]_  = ~A168 & A169;
  assign \new_[22143]_  = ~A201 & A200;
  assign \new_[22144]_  = ~A199 & \new_[22143]_ ;
  assign \new_[22145]_  = \new_[22144]_  & \new_[22139]_ ;
  assign \new_[22149]_  = ~A267 & A203;
  assign \new_[22150]_  = ~A202 & \new_[22149]_ ;
  assign \new_[22154]_  = A299 & A298;
  assign \new_[22155]_  = A268 & \new_[22154]_ ;
  assign \new_[22156]_  = \new_[22155]_  & \new_[22150]_ ;
  assign \new_[22159]_  = ~A168 & A169;
  assign \new_[22163]_  = ~A201 & A200;
  assign \new_[22164]_  = ~A199 & \new_[22163]_ ;
  assign \new_[22165]_  = \new_[22164]_  & \new_[22159]_ ;
  assign \new_[22169]_  = ~A267 & A203;
  assign \new_[22170]_  = ~A202 & \new_[22169]_ ;
  assign \new_[22174]_  = ~A299 & ~A298;
  assign \new_[22175]_  = A268 & \new_[22174]_ ;
  assign \new_[22176]_  = \new_[22175]_  & \new_[22170]_ ;
  assign \new_[22179]_  = ~A168 & A169;
  assign \new_[22183]_  = ~A201 & A200;
  assign \new_[22184]_  = ~A199 & \new_[22183]_ ;
  assign \new_[22185]_  = \new_[22184]_  & \new_[22179]_ ;
  assign \new_[22189]_  = ~A267 & A203;
  assign \new_[22190]_  = ~A202 & \new_[22189]_ ;
  assign \new_[22194]_  = A301 & ~A300;
  assign \new_[22195]_  = ~A269 & \new_[22194]_ ;
  assign \new_[22196]_  = \new_[22195]_  & \new_[22190]_ ;
  assign \new_[22199]_  = ~A168 & A169;
  assign \new_[22203]_  = ~A201 & A200;
  assign \new_[22204]_  = ~A199 & \new_[22203]_ ;
  assign \new_[22205]_  = \new_[22204]_  & \new_[22199]_ ;
  assign \new_[22209]_  = ~A267 & A203;
  assign \new_[22210]_  = ~A202 & \new_[22209]_ ;
  assign \new_[22214]_  = ~A302 & ~A300;
  assign \new_[22215]_  = ~A269 & \new_[22214]_ ;
  assign \new_[22216]_  = \new_[22215]_  & \new_[22210]_ ;
  assign \new_[22219]_  = ~A168 & A169;
  assign \new_[22223]_  = ~A201 & A200;
  assign \new_[22224]_  = ~A199 & \new_[22223]_ ;
  assign \new_[22225]_  = \new_[22224]_  & \new_[22219]_ ;
  assign \new_[22229]_  = ~A267 & A203;
  assign \new_[22230]_  = ~A202 & \new_[22229]_ ;
  assign \new_[22234]_  = A299 & A298;
  assign \new_[22235]_  = ~A269 & \new_[22234]_ ;
  assign \new_[22236]_  = \new_[22235]_  & \new_[22230]_ ;
  assign \new_[22239]_  = ~A168 & A169;
  assign \new_[22243]_  = ~A201 & A200;
  assign \new_[22244]_  = ~A199 & \new_[22243]_ ;
  assign \new_[22245]_  = \new_[22244]_  & \new_[22239]_ ;
  assign \new_[22249]_  = ~A267 & A203;
  assign \new_[22250]_  = ~A202 & \new_[22249]_ ;
  assign \new_[22254]_  = ~A299 & ~A298;
  assign \new_[22255]_  = ~A269 & \new_[22254]_ ;
  assign \new_[22256]_  = \new_[22255]_  & \new_[22250]_ ;
  assign \new_[22259]_  = ~A168 & A169;
  assign \new_[22263]_  = ~A201 & A200;
  assign \new_[22264]_  = ~A199 & \new_[22263]_ ;
  assign \new_[22265]_  = \new_[22264]_  & \new_[22259]_ ;
  assign \new_[22269]_  = A265 & A203;
  assign \new_[22270]_  = ~A202 & \new_[22269]_ ;
  assign \new_[22274]_  = A301 & ~A300;
  assign \new_[22275]_  = A266 & \new_[22274]_ ;
  assign \new_[22276]_  = \new_[22275]_  & \new_[22270]_ ;
  assign \new_[22279]_  = ~A168 & A169;
  assign \new_[22283]_  = ~A201 & A200;
  assign \new_[22284]_  = ~A199 & \new_[22283]_ ;
  assign \new_[22285]_  = \new_[22284]_  & \new_[22279]_ ;
  assign \new_[22289]_  = A265 & A203;
  assign \new_[22290]_  = ~A202 & \new_[22289]_ ;
  assign \new_[22294]_  = ~A302 & ~A300;
  assign \new_[22295]_  = A266 & \new_[22294]_ ;
  assign \new_[22296]_  = \new_[22295]_  & \new_[22290]_ ;
  assign \new_[22299]_  = ~A168 & A169;
  assign \new_[22303]_  = ~A201 & A200;
  assign \new_[22304]_  = ~A199 & \new_[22303]_ ;
  assign \new_[22305]_  = \new_[22304]_  & \new_[22299]_ ;
  assign \new_[22309]_  = A265 & A203;
  assign \new_[22310]_  = ~A202 & \new_[22309]_ ;
  assign \new_[22314]_  = A299 & A298;
  assign \new_[22315]_  = A266 & \new_[22314]_ ;
  assign \new_[22316]_  = \new_[22315]_  & \new_[22310]_ ;
  assign \new_[22319]_  = ~A168 & A169;
  assign \new_[22323]_  = ~A201 & A200;
  assign \new_[22324]_  = ~A199 & \new_[22323]_ ;
  assign \new_[22325]_  = \new_[22324]_  & \new_[22319]_ ;
  assign \new_[22329]_  = A265 & A203;
  assign \new_[22330]_  = ~A202 & \new_[22329]_ ;
  assign \new_[22334]_  = ~A299 & ~A298;
  assign \new_[22335]_  = A266 & \new_[22334]_ ;
  assign \new_[22336]_  = \new_[22335]_  & \new_[22330]_ ;
  assign \new_[22339]_  = ~A168 & A169;
  assign \new_[22343]_  = ~A201 & A200;
  assign \new_[22344]_  = ~A199 & \new_[22343]_ ;
  assign \new_[22345]_  = \new_[22344]_  & \new_[22339]_ ;
  assign \new_[22349]_  = ~A265 & A203;
  assign \new_[22350]_  = ~A202 & \new_[22349]_ ;
  assign \new_[22354]_  = A301 & ~A300;
  assign \new_[22355]_  = ~A266 & \new_[22354]_ ;
  assign \new_[22356]_  = \new_[22355]_  & \new_[22350]_ ;
  assign \new_[22359]_  = ~A168 & A169;
  assign \new_[22363]_  = ~A201 & A200;
  assign \new_[22364]_  = ~A199 & \new_[22363]_ ;
  assign \new_[22365]_  = \new_[22364]_  & \new_[22359]_ ;
  assign \new_[22369]_  = ~A265 & A203;
  assign \new_[22370]_  = ~A202 & \new_[22369]_ ;
  assign \new_[22374]_  = ~A302 & ~A300;
  assign \new_[22375]_  = ~A266 & \new_[22374]_ ;
  assign \new_[22376]_  = \new_[22375]_  & \new_[22370]_ ;
  assign \new_[22379]_  = ~A168 & A169;
  assign \new_[22383]_  = ~A201 & A200;
  assign \new_[22384]_  = ~A199 & \new_[22383]_ ;
  assign \new_[22385]_  = \new_[22384]_  & \new_[22379]_ ;
  assign \new_[22389]_  = ~A265 & A203;
  assign \new_[22390]_  = ~A202 & \new_[22389]_ ;
  assign \new_[22394]_  = A299 & A298;
  assign \new_[22395]_  = ~A266 & \new_[22394]_ ;
  assign \new_[22396]_  = \new_[22395]_  & \new_[22390]_ ;
  assign \new_[22399]_  = ~A168 & A169;
  assign \new_[22403]_  = ~A201 & A200;
  assign \new_[22404]_  = ~A199 & \new_[22403]_ ;
  assign \new_[22405]_  = \new_[22404]_  & \new_[22399]_ ;
  assign \new_[22409]_  = ~A265 & A203;
  assign \new_[22410]_  = ~A202 & \new_[22409]_ ;
  assign \new_[22414]_  = ~A299 & ~A298;
  assign \new_[22415]_  = ~A266 & \new_[22414]_ ;
  assign \new_[22416]_  = \new_[22415]_  & \new_[22410]_ ;
  assign \new_[22419]_  = ~A168 & A169;
  assign \new_[22423]_  = A201 & ~A200;
  assign \new_[22424]_  = A199 & \new_[22423]_ ;
  assign \new_[22425]_  = \new_[22424]_  & \new_[22419]_ ;
  assign \new_[22429]_  = ~A268 & A267;
  assign \new_[22430]_  = A202 & \new_[22429]_ ;
  assign \new_[22434]_  = A301 & ~A300;
  assign \new_[22435]_  = A269 & \new_[22434]_ ;
  assign \new_[22436]_  = \new_[22435]_  & \new_[22430]_ ;
  assign \new_[22439]_  = ~A168 & A169;
  assign \new_[22443]_  = A201 & ~A200;
  assign \new_[22444]_  = A199 & \new_[22443]_ ;
  assign \new_[22445]_  = \new_[22444]_  & \new_[22439]_ ;
  assign \new_[22449]_  = ~A268 & A267;
  assign \new_[22450]_  = A202 & \new_[22449]_ ;
  assign \new_[22454]_  = ~A302 & ~A300;
  assign \new_[22455]_  = A269 & \new_[22454]_ ;
  assign \new_[22456]_  = \new_[22455]_  & \new_[22450]_ ;
  assign \new_[22459]_  = ~A168 & A169;
  assign \new_[22463]_  = A201 & ~A200;
  assign \new_[22464]_  = A199 & \new_[22463]_ ;
  assign \new_[22465]_  = \new_[22464]_  & \new_[22459]_ ;
  assign \new_[22469]_  = ~A268 & A267;
  assign \new_[22470]_  = A202 & \new_[22469]_ ;
  assign \new_[22474]_  = A299 & A298;
  assign \new_[22475]_  = A269 & \new_[22474]_ ;
  assign \new_[22476]_  = \new_[22475]_  & \new_[22470]_ ;
  assign \new_[22479]_  = ~A168 & A169;
  assign \new_[22483]_  = A201 & ~A200;
  assign \new_[22484]_  = A199 & \new_[22483]_ ;
  assign \new_[22485]_  = \new_[22484]_  & \new_[22479]_ ;
  assign \new_[22489]_  = ~A268 & A267;
  assign \new_[22490]_  = A202 & \new_[22489]_ ;
  assign \new_[22494]_  = ~A299 & ~A298;
  assign \new_[22495]_  = A269 & \new_[22494]_ ;
  assign \new_[22496]_  = \new_[22495]_  & \new_[22490]_ ;
  assign \new_[22499]_  = ~A168 & A169;
  assign \new_[22503]_  = A201 & ~A200;
  assign \new_[22504]_  = A199 & \new_[22503]_ ;
  assign \new_[22505]_  = \new_[22504]_  & \new_[22499]_ ;
  assign \new_[22509]_  = A268 & ~A267;
  assign \new_[22510]_  = A202 & \new_[22509]_ ;
  assign \new_[22514]_  = A302 & ~A301;
  assign \new_[22515]_  = A300 & \new_[22514]_ ;
  assign \new_[22516]_  = \new_[22515]_  & \new_[22510]_ ;
  assign \new_[22519]_  = ~A168 & A169;
  assign \new_[22523]_  = A201 & ~A200;
  assign \new_[22524]_  = A199 & \new_[22523]_ ;
  assign \new_[22525]_  = \new_[22524]_  & \new_[22519]_ ;
  assign \new_[22529]_  = ~A269 & ~A267;
  assign \new_[22530]_  = A202 & \new_[22529]_ ;
  assign \new_[22534]_  = A302 & ~A301;
  assign \new_[22535]_  = A300 & \new_[22534]_ ;
  assign \new_[22536]_  = \new_[22535]_  & \new_[22530]_ ;
  assign \new_[22539]_  = ~A168 & A169;
  assign \new_[22543]_  = A201 & ~A200;
  assign \new_[22544]_  = A199 & \new_[22543]_ ;
  assign \new_[22545]_  = \new_[22544]_  & \new_[22539]_ ;
  assign \new_[22549]_  = A266 & A265;
  assign \new_[22550]_  = A202 & \new_[22549]_ ;
  assign \new_[22554]_  = A302 & ~A301;
  assign \new_[22555]_  = A300 & \new_[22554]_ ;
  assign \new_[22556]_  = \new_[22555]_  & \new_[22550]_ ;
  assign \new_[22559]_  = ~A168 & A169;
  assign \new_[22563]_  = A201 & ~A200;
  assign \new_[22564]_  = A199 & \new_[22563]_ ;
  assign \new_[22565]_  = \new_[22564]_  & \new_[22559]_ ;
  assign \new_[22569]_  = ~A266 & ~A265;
  assign \new_[22570]_  = A202 & \new_[22569]_ ;
  assign \new_[22574]_  = A302 & ~A301;
  assign \new_[22575]_  = A300 & \new_[22574]_ ;
  assign \new_[22576]_  = \new_[22575]_  & \new_[22570]_ ;
  assign \new_[22579]_  = ~A168 & A169;
  assign \new_[22583]_  = A201 & ~A200;
  assign \new_[22584]_  = A199 & \new_[22583]_ ;
  assign \new_[22585]_  = \new_[22584]_  & \new_[22579]_ ;
  assign \new_[22589]_  = ~A268 & A267;
  assign \new_[22590]_  = ~A203 & \new_[22589]_ ;
  assign \new_[22594]_  = A301 & ~A300;
  assign \new_[22595]_  = A269 & \new_[22594]_ ;
  assign \new_[22596]_  = \new_[22595]_  & \new_[22590]_ ;
  assign \new_[22599]_  = ~A168 & A169;
  assign \new_[22603]_  = A201 & ~A200;
  assign \new_[22604]_  = A199 & \new_[22603]_ ;
  assign \new_[22605]_  = \new_[22604]_  & \new_[22599]_ ;
  assign \new_[22609]_  = ~A268 & A267;
  assign \new_[22610]_  = ~A203 & \new_[22609]_ ;
  assign \new_[22614]_  = ~A302 & ~A300;
  assign \new_[22615]_  = A269 & \new_[22614]_ ;
  assign \new_[22616]_  = \new_[22615]_  & \new_[22610]_ ;
  assign \new_[22619]_  = ~A168 & A169;
  assign \new_[22623]_  = A201 & ~A200;
  assign \new_[22624]_  = A199 & \new_[22623]_ ;
  assign \new_[22625]_  = \new_[22624]_  & \new_[22619]_ ;
  assign \new_[22629]_  = ~A268 & A267;
  assign \new_[22630]_  = ~A203 & \new_[22629]_ ;
  assign \new_[22634]_  = A299 & A298;
  assign \new_[22635]_  = A269 & \new_[22634]_ ;
  assign \new_[22636]_  = \new_[22635]_  & \new_[22630]_ ;
  assign \new_[22639]_  = ~A168 & A169;
  assign \new_[22643]_  = A201 & ~A200;
  assign \new_[22644]_  = A199 & \new_[22643]_ ;
  assign \new_[22645]_  = \new_[22644]_  & \new_[22639]_ ;
  assign \new_[22649]_  = ~A268 & A267;
  assign \new_[22650]_  = ~A203 & \new_[22649]_ ;
  assign \new_[22654]_  = ~A299 & ~A298;
  assign \new_[22655]_  = A269 & \new_[22654]_ ;
  assign \new_[22656]_  = \new_[22655]_  & \new_[22650]_ ;
  assign \new_[22659]_  = ~A168 & A169;
  assign \new_[22663]_  = A201 & ~A200;
  assign \new_[22664]_  = A199 & \new_[22663]_ ;
  assign \new_[22665]_  = \new_[22664]_  & \new_[22659]_ ;
  assign \new_[22669]_  = A268 & ~A267;
  assign \new_[22670]_  = ~A203 & \new_[22669]_ ;
  assign \new_[22674]_  = A302 & ~A301;
  assign \new_[22675]_  = A300 & \new_[22674]_ ;
  assign \new_[22676]_  = \new_[22675]_  & \new_[22670]_ ;
  assign \new_[22679]_  = ~A168 & A169;
  assign \new_[22683]_  = A201 & ~A200;
  assign \new_[22684]_  = A199 & \new_[22683]_ ;
  assign \new_[22685]_  = \new_[22684]_  & \new_[22679]_ ;
  assign \new_[22689]_  = ~A269 & ~A267;
  assign \new_[22690]_  = ~A203 & \new_[22689]_ ;
  assign \new_[22694]_  = A302 & ~A301;
  assign \new_[22695]_  = A300 & \new_[22694]_ ;
  assign \new_[22696]_  = \new_[22695]_  & \new_[22690]_ ;
  assign \new_[22699]_  = ~A168 & A169;
  assign \new_[22703]_  = A201 & ~A200;
  assign \new_[22704]_  = A199 & \new_[22703]_ ;
  assign \new_[22705]_  = \new_[22704]_  & \new_[22699]_ ;
  assign \new_[22709]_  = A266 & A265;
  assign \new_[22710]_  = ~A203 & \new_[22709]_ ;
  assign \new_[22714]_  = A302 & ~A301;
  assign \new_[22715]_  = A300 & \new_[22714]_ ;
  assign \new_[22716]_  = \new_[22715]_  & \new_[22710]_ ;
  assign \new_[22719]_  = ~A168 & A169;
  assign \new_[22723]_  = A201 & ~A200;
  assign \new_[22724]_  = A199 & \new_[22723]_ ;
  assign \new_[22725]_  = \new_[22724]_  & \new_[22719]_ ;
  assign \new_[22729]_  = ~A266 & ~A265;
  assign \new_[22730]_  = ~A203 & \new_[22729]_ ;
  assign \new_[22734]_  = A302 & ~A301;
  assign \new_[22735]_  = A300 & \new_[22734]_ ;
  assign \new_[22736]_  = \new_[22735]_  & \new_[22730]_ ;
  assign \new_[22739]_  = ~A168 & A169;
  assign \new_[22743]_  = ~A201 & ~A200;
  assign \new_[22744]_  = A199 & \new_[22743]_ ;
  assign \new_[22745]_  = \new_[22744]_  & \new_[22739]_ ;
  assign \new_[22749]_  = ~A267 & A203;
  assign \new_[22750]_  = ~A202 & \new_[22749]_ ;
  assign \new_[22754]_  = A301 & ~A300;
  assign \new_[22755]_  = A268 & \new_[22754]_ ;
  assign \new_[22756]_  = \new_[22755]_  & \new_[22750]_ ;
  assign \new_[22759]_  = ~A168 & A169;
  assign \new_[22763]_  = ~A201 & ~A200;
  assign \new_[22764]_  = A199 & \new_[22763]_ ;
  assign \new_[22765]_  = \new_[22764]_  & \new_[22759]_ ;
  assign \new_[22769]_  = ~A267 & A203;
  assign \new_[22770]_  = ~A202 & \new_[22769]_ ;
  assign \new_[22774]_  = ~A302 & ~A300;
  assign \new_[22775]_  = A268 & \new_[22774]_ ;
  assign \new_[22776]_  = \new_[22775]_  & \new_[22770]_ ;
  assign \new_[22779]_  = ~A168 & A169;
  assign \new_[22783]_  = ~A201 & ~A200;
  assign \new_[22784]_  = A199 & \new_[22783]_ ;
  assign \new_[22785]_  = \new_[22784]_  & \new_[22779]_ ;
  assign \new_[22789]_  = ~A267 & A203;
  assign \new_[22790]_  = ~A202 & \new_[22789]_ ;
  assign \new_[22794]_  = A299 & A298;
  assign \new_[22795]_  = A268 & \new_[22794]_ ;
  assign \new_[22796]_  = \new_[22795]_  & \new_[22790]_ ;
  assign \new_[22799]_  = ~A168 & A169;
  assign \new_[22803]_  = ~A201 & ~A200;
  assign \new_[22804]_  = A199 & \new_[22803]_ ;
  assign \new_[22805]_  = \new_[22804]_  & \new_[22799]_ ;
  assign \new_[22809]_  = ~A267 & A203;
  assign \new_[22810]_  = ~A202 & \new_[22809]_ ;
  assign \new_[22814]_  = ~A299 & ~A298;
  assign \new_[22815]_  = A268 & \new_[22814]_ ;
  assign \new_[22816]_  = \new_[22815]_  & \new_[22810]_ ;
  assign \new_[22819]_  = ~A168 & A169;
  assign \new_[22823]_  = ~A201 & ~A200;
  assign \new_[22824]_  = A199 & \new_[22823]_ ;
  assign \new_[22825]_  = \new_[22824]_  & \new_[22819]_ ;
  assign \new_[22829]_  = ~A267 & A203;
  assign \new_[22830]_  = ~A202 & \new_[22829]_ ;
  assign \new_[22834]_  = A301 & ~A300;
  assign \new_[22835]_  = ~A269 & \new_[22834]_ ;
  assign \new_[22836]_  = \new_[22835]_  & \new_[22830]_ ;
  assign \new_[22839]_  = ~A168 & A169;
  assign \new_[22843]_  = ~A201 & ~A200;
  assign \new_[22844]_  = A199 & \new_[22843]_ ;
  assign \new_[22845]_  = \new_[22844]_  & \new_[22839]_ ;
  assign \new_[22849]_  = ~A267 & A203;
  assign \new_[22850]_  = ~A202 & \new_[22849]_ ;
  assign \new_[22854]_  = ~A302 & ~A300;
  assign \new_[22855]_  = ~A269 & \new_[22854]_ ;
  assign \new_[22856]_  = \new_[22855]_  & \new_[22850]_ ;
  assign \new_[22859]_  = ~A168 & A169;
  assign \new_[22863]_  = ~A201 & ~A200;
  assign \new_[22864]_  = A199 & \new_[22863]_ ;
  assign \new_[22865]_  = \new_[22864]_  & \new_[22859]_ ;
  assign \new_[22869]_  = ~A267 & A203;
  assign \new_[22870]_  = ~A202 & \new_[22869]_ ;
  assign \new_[22874]_  = A299 & A298;
  assign \new_[22875]_  = ~A269 & \new_[22874]_ ;
  assign \new_[22876]_  = \new_[22875]_  & \new_[22870]_ ;
  assign \new_[22879]_  = ~A168 & A169;
  assign \new_[22883]_  = ~A201 & ~A200;
  assign \new_[22884]_  = A199 & \new_[22883]_ ;
  assign \new_[22885]_  = \new_[22884]_  & \new_[22879]_ ;
  assign \new_[22889]_  = ~A267 & A203;
  assign \new_[22890]_  = ~A202 & \new_[22889]_ ;
  assign \new_[22894]_  = ~A299 & ~A298;
  assign \new_[22895]_  = ~A269 & \new_[22894]_ ;
  assign \new_[22896]_  = \new_[22895]_  & \new_[22890]_ ;
  assign \new_[22899]_  = ~A168 & A169;
  assign \new_[22903]_  = ~A201 & ~A200;
  assign \new_[22904]_  = A199 & \new_[22903]_ ;
  assign \new_[22905]_  = \new_[22904]_  & \new_[22899]_ ;
  assign \new_[22909]_  = A265 & A203;
  assign \new_[22910]_  = ~A202 & \new_[22909]_ ;
  assign \new_[22914]_  = A301 & ~A300;
  assign \new_[22915]_  = A266 & \new_[22914]_ ;
  assign \new_[22916]_  = \new_[22915]_  & \new_[22910]_ ;
  assign \new_[22919]_  = ~A168 & A169;
  assign \new_[22923]_  = ~A201 & ~A200;
  assign \new_[22924]_  = A199 & \new_[22923]_ ;
  assign \new_[22925]_  = \new_[22924]_  & \new_[22919]_ ;
  assign \new_[22929]_  = A265 & A203;
  assign \new_[22930]_  = ~A202 & \new_[22929]_ ;
  assign \new_[22934]_  = ~A302 & ~A300;
  assign \new_[22935]_  = A266 & \new_[22934]_ ;
  assign \new_[22936]_  = \new_[22935]_  & \new_[22930]_ ;
  assign \new_[22939]_  = ~A168 & A169;
  assign \new_[22943]_  = ~A201 & ~A200;
  assign \new_[22944]_  = A199 & \new_[22943]_ ;
  assign \new_[22945]_  = \new_[22944]_  & \new_[22939]_ ;
  assign \new_[22949]_  = A265 & A203;
  assign \new_[22950]_  = ~A202 & \new_[22949]_ ;
  assign \new_[22954]_  = A299 & A298;
  assign \new_[22955]_  = A266 & \new_[22954]_ ;
  assign \new_[22956]_  = \new_[22955]_  & \new_[22950]_ ;
  assign \new_[22959]_  = ~A168 & A169;
  assign \new_[22963]_  = ~A201 & ~A200;
  assign \new_[22964]_  = A199 & \new_[22963]_ ;
  assign \new_[22965]_  = \new_[22964]_  & \new_[22959]_ ;
  assign \new_[22969]_  = A265 & A203;
  assign \new_[22970]_  = ~A202 & \new_[22969]_ ;
  assign \new_[22974]_  = ~A299 & ~A298;
  assign \new_[22975]_  = A266 & \new_[22974]_ ;
  assign \new_[22976]_  = \new_[22975]_  & \new_[22970]_ ;
  assign \new_[22979]_  = ~A168 & A169;
  assign \new_[22983]_  = ~A201 & ~A200;
  assign \new_[22984]_  = A199 & \new_[22983]_ ;
  assign \new_[22985]_  = \new_[22984]_  & \new_[22979]_ ;
  assign \new_[22989]_  = ~A265 & A203;
  assign \new_[22990]_  = ~A202 & \new_[22989]_ ;
  assign \new_[22994]_  = A301 & ~A300;
  assign \new_[22995]_  = ~A266 & \new_[22994]_ ;
  assign \new_[22996]_  = \new_[22995]_  & \new_[22990]_ ;
  assign \new_[22999]_  = ~A168 & A169;
  assign \new_[23003]_  = ~A201 & ~A200;
  assign \new_[23004]_  = A199 & \new_[23003]_ ;
  assign \new_[23005]_  = \new_[23004]_  & \new_[22999]_ ;
  assign \new_[23009]_  = ~A265 & A203;
  assign \new_[23010]_  = ~A202 & \new_[23009]_ ;
  assign \new_[23014]_  = ~A302 & ~A300;
  assign \new_[23015]_  = ~A266 & \new_[23014]_ ;
  assign \new_[23016]_  = \new_[23015]_  & \new_[23010]_ ;
  assign \new_[23019]_  = ~A168 & A169;
  assign \new_[23023]_  = ~A201 & ~A200;
  assign \new_[23024]_  = A199 & \new_[23023]_ ;
  assign \new_[23025]_  = \new_[23024]_  & \new_[23019]_ ;
  assign \new_[23029]_  = ~A265 & A203;
  assign \new_[23030]_  = ~A202 & \new_[23029]_ ;
  assign \new_[23034]_  = A299 & A298;
  assign \new_[23035]_  = ~A266 & \new_[23034]_ ;
  assign \new_[23036]_  = \new_[23035]_  & \new_[23030]_ ;
  assign \new_[23039]_  = ~A168 & A169;
  assign \new_[23043]_  = ~A201 & ~A200;
  assign \new_[23044]_  = A199 & \new_[23043]_ ;
  assign \new_[23045]_  = \new_[23044]_  & \new_[23039]_ ;
  assign \new_[23049]_  = ~A265 & A203;
  assign \new_[23050]_  = ~A202 & \new_[23049]_ ;
  assign \new_[23054]_  = ~A299 & ~A298;
  assign \new_[23055]_  = ~A266 & \new_[23054]_ ;
  assign \new_[23056]_  = \new_[23055]_  & \new_[23050]_ ;
  assign \new_[23059]_  = ~A169 & ~A170;
  assign \new_[23063]_  = A234 & A233;
  assign \new_[23064]_  = ~A232 & \new_[23063]_ ;
  assign \new_[23065]_  = \new_[23064]_  & \new_[23059]_ ;
  assign \new_[23069]_  = A266 & ~A265;
  assign \new_[23070]_  = A235 & \new_[23069]_ ;
  assign \new_[23074]_  = A269 & ~A268;
  assign \new_[23075]_  = ~A267 & \new_[23074]_ ;
  assign \new_[23076]_  = \new_[23075]_  & \new_[23070]_ ;
  assign \new_[23079]_  = ~A169 & ~A170;
  assign \new_[23083]_  = A234 & A233;
  assign \new_[23084]_  = ~A232 & \new_[23083]_ ;
  assign \new_[23085]_  = \new_[23084]_  & \new_[23079]_ ;
  assign \new_[23089]_  = ~A266 & A265;
  assign \new_[23090]_  = A235 & \new_[23089]_ ;
  assign \new_[23094]_  = A269 & ~A268;
  assign \new_[23095]_  = ~A267 & \new_[23094]_ ;
  assign \new_[23096]_  = \new_[23095]_  & \new_[23090]_ ;
  assign \new_[23099]_  = ~A169 & ~A170;
  assign \new_[23103]_  = A234 & A233;
  assign \new_[23104]_  = ~A232 & \new_[23103]_ ;
  assign \new_[23105]_  = \new_[23104]_  & \new_[23099]_ ;
  assign \new_[23109]_  = A266 & ~A265;
  assign \new_[23110]_  = ~A236 & \new_[23109]_ ;
  assign \new_[23114]_  = A269 & ~A268;
  assign \new_[23115]_  = ~A267 & \new_[23114]_ ;
  assign \new_[23116]_  = \new_[23115]_  & \new_[23110]_ ;
  assign \new_[23119]_  = ~A169 & ~A170;
  assign \new_[23123]_  = A234 & A233;
  assign \new_[23124]_  = ~A232 & \new_[23123]_ ;
  assign \new_[23125]_  = \new_[23124]_  & \new_[23119]_ ;
  assign \new_[23129]_  = ~A266 & A265;
  assign \new_[23130]_  = ~A236 & \new_[23129]_ ;
  assign \new_[23134]_  = A269 & ~A268;
  assign \new_[23135]_  = ~A267 & \new_[23134]_ ;
  assign \new_[23136]_  = \new_[23135]_  & \new_[23130]_ ;
  assign \new_[23139]_  = ~A169 & ~A170;
  assign \new_[23143]_  = A234 & ~A233;
  assign \new_[23144]_  = A232 & \new_[23143]_ ;
  assign \new_[23145]_  = \new_[23144]_  & \new_[23139]_ ;
  assign \new_[23149]_  = A266 & ~A265;
  assign \new_[23150]_  = A235 & \new_[23149]_ ;
  assign \new_[23154]_  = A269 & ~A268;
  assign \new_[23155]_  = ~A267 & \new_[23154]_ ;
  assign \new_[23156]_  = \new_[23155]_  & \new_[23150]_ ;
  assign \new_[23159]_  = ~A169 & ~A170;
  assign \new_[23163]_  = A234 & ~A233;
  assign \new_[23164]_  = A232 & \new_[23163]_ ;
  assign \new_[23165]_  = \new_[23164]_  & \new_[23159]_ ;
  assign \new_[23169]_  = ~A266 & A265;
  assign \new_[23170]_  = A235 & \new_[23169]_ ;
  assign \new_[23174]_  = A269 & ~A268;
  assign \new_[23175]_  = ~A267 & \new_[23174]_ ;
  assign \new_[23176]_  = \new_[23175]_  & \new_[23170]_ ;
  assign \new_[23179]_  = ~A169 & ~A170;
  assign \new_[23183]_  = A234 & ~A233;
  assign \new_[23184]_  = A232 & \new_[23183]_ ;
  assign \new_[23185]_  = \new_[23184]_  & \new_[23179]_ ;
  assign \new_[23189]_  = A266 & ~A265;
  assign \new_[23190]_  = ~A236 & \new_[23189]_ ;
  assign \new_[23194]_  = A269 & ~A268;
  assign \new_[23195]_  = ~A267 & \new_[23194]_ ;
  assign \new_[23196]_  = \new_[23195]_  & \new_[23190]_ ;
  assign \new_[23199]_  = ~A169 & ~A170;
  assign \new_[23203]_  = A234 & ~A233;
  assign \new_[23204]_  = A232 & \new_[23203]_ ;
  assign \new_[23205]_  = \new_[23204]_  & \new_[23199]_ ;
  assign \new_[23209]_  = ~A266 & A265;
  assign \new_[23210]_  = ~A236 & \new_[23209]_ ;
  assign \new_[23214]_  = A269 & ~A268;
  assign \new_[23215]_  = ~A267 & \new_[23214]_ ;
  assign \new_[23216]_  = \new_[23215]_  & \new_[23210]_ ;
  assign \new_[23219]_  = ~A169 & ~A170;
  assign \new_[23223]_  = A200 & ~A199;
  assign \new_[23224]_  = A168 & \new_[23223]_ ;
  assign \new_[23225]_  = \new_[23224]_  & \new_[23219]_ ;
  assign \new_[23229]_  = ~A267 & A202;
  assign \new_[23230]_  = A201 & \new_[23229]_ ;
  assign \new_[23234]_  = A301 & ~A300;
  assign \new_[23235]_  = A268 & \new_[23234]_ ;
  assign \new_[23236]_  = \new_[23235]_  & \new_[23230]_ ;
  assign \new_[23239]_  = ~A169 & ~A170;
  assign \new_[23243]_  = A200 & ~A199;
  assign \new_[23244]_  = A168 & \new_[23243]_ ;
  assign \new_[23245]_  = \new_[23244]_  & \new_[23239]_ ;
  assign \new_[23249]_  = ~A267 & A202;
  assign \new_[23250]_  = A201 & \new_[23249]_ ;
  assign \new_[23254]_  = ~A302 & ~A300;
  assign \new_[23255]_  = A268 & \new_[23254]_ ;
  assign \new_[23256]_  = \new_[23255]_  & \new_[23250]_ ;
  assign \new_[23259]_  = ~A169 & ~A170;
  assign \new_[23263]_  = A200 & ~A199;
  assign \new_[23264]_  = A168 & \new_[23263]_ ;
  assign \new_[23265]_  = \new_[23264]_  & \new_[23259]_ ;
  assign \new_[23269]_  = ~A267 & A202;
  assign \new_[23270]_  = A201 & \new_[23269]_ ;
  assign \new_[23274]_  = A299 & A298;
  assign \new_[23275]_  = A268 & \new_[23274]_ ;
  assign \new_[23276]_  = \new_[23275]_  & \new_[23270]_ ;
  assign \new_[23279]_  = ~A169 & ~A170;
  assign \new_[23283]_  = A200 & ~A199;
  assign \new_[23284]_  = A168 & \new_[23283]_ ;
  assign \new_[23285]_  = \new_[23284]_  & \new_[23279]_ ;
  assign \new_[23289]_  = ~A267 & A202;
  assign \new_[23290]_  = A201 & \new_[23289]_ ;
  assign \new_[23294]_  = ~A299 & ~A298;
  assign \new_[23295]_  = A268 & \new_[23294]_ ;
  assign \new_[23296]_  = \new_[23295]_  & \new_[23290]_ ;
  assign \new_[23299]_  = ~A169 & ~A170;
  assign \new_[23303]_  = A200 & ~A199;
  assign \new_[23304]_  = A168 & \new_[23303]_ ;
  assign \new_[23305]_  = \new_[23304]_  & \new_[23299]_ ;
  assign \new_[23309]_  = ~A267 & A202;
  assign \new_[23310]_  = A201 & \new_[23309]_ ;
  assign \new_[23314]_  = A301 & ~A300;
  assign \new_[23315]_  = ~A269 & \new_[23314]_ ;
  assign \new_[23316]_  = \new_[23315]_  & \new_[23310]_ ;
  assign \new_[23319]_  = ~A169 & ~A170;
  assign \new_[23323]_  = A200 & ~A199;
  assign \new_[23324]_  = A168 & \new_[23323]_ ;
  assign \new_[23325]_  = \new_[23324]_  & \new_[23319]_ ;
  assign \new_[23329]_  = ~A267 & A202;
  assign \new_[23330]_  = A201 & \new_[23329]_ ;
  assign \new_[23334]_  = ~A302 & ~A300;
  assign \new_[23335]_  = ~A269 & \new_[23334]_ ;
  assign \new_[23336]_  = \new_[23335]_  & \new_[23330]_ ;
  assign \new_[23339]_  = ~A169 & ~A170;
  assign \new_[23343]_  = A200 & ~A199;
  assign \new_[23344]_  = A168 & \new_[23343]_ ;
  assign \new_[23345]_  = \new_[23344]_  & \new_[23339]_ ;
  assign \new_[23349]_  = ~A267 & A202;
  assign \new_[23350]_  = A201 & \new_[23349]_ ;
  assign \new_[23354]_  = A299 & A298;
  assign \new_[23355]_  = ~A269 & \new_[23354]_ ;
  assign \new_[23356]_  = \new_[23355]_  & \new_[23350]_ ;
  assign \new_[23359]_  = ~A169 & ~A170;
  assign \new_[23363]_  = A200 & ~A199;
  assign \new_[23364]_  = A168 & \new_[23363]_ ;
  assign \new_[23365]_  = \new_[23364]_  & \new_[23359]_ ;
  assign \new_[23369]_  = ~A267 & A202;
  assign \new_[23370]_  = A201 & \new_[23369]_ ;
  assign \new_[23374]_  = ~A299 & ~A298;
  assign \new_[23375]_  = ~A269 & \new_[23374]_ ;
  assign \new_[23376]_  = \new_[23375]_  & \new_[23370]_ ;
  assign \new_[23379]_  = ~A169 & ~A170;
  assign \new_[23383]_  = A200 & ~A199;
  assign \new_[23384]_  = A168 & \new_[23383]_ ;
  assign \new_[23385]_  = \new_[23384]_  & \new_[23379]_ ;
  assign \new_[23389]_  = A265 & A202;
  assign \new_[23390]_  = A201 & \new_[23389]_ ;
  assign \new_[23394]_  = A301 & ~A300;
  assign \new_[23395]_  = A266 & \new_[23394]_ ;
  assign \new_[23396]_  = \new_[23395]_  & \new_[23390]_ ;
  assign \new_[23399]_  = ~A169 & ~A170;
  assign \new_[23403]_  = A200 & ~A199;
  assign \new_[23404]_  = A168 & \new_[23403]_ ;
  assign \new_[23405]_  = \new_[23404]_  & \new_[23399]_ ;
  assign \new_[23409]_  = A265 & A202;
  assign \new_[23410]_  = A201 & \new_[23409]_ ;
  assign \new_[23414]_  = ~A302 & ~A300;
  assign \new_[23415]_  = A266 & \new_[23414]_ ;
  assign \new_[23416]_  = \new_[23415]_  & \new_[23410]_ ;
  assign \new_[23419]_  = ~A169 & ~A170;
  assign \new_[23423]_  = A200 & ~A199;
  assign \new_[23424]_  = A168 & \new_[23423]_ ;
  assign \new_[23425]_  = \new_[23424]_  & \new_[23419]_ ;
  assign \new_[23429]_  = A265 & A202;
  assign \new_[23430]_  = A201 & \new_[23429]_ ;
  assign \new_[23434]_  = A299 & A298;
  assign \new_[23435]_  = A266 & \new_[23434]_ ;
  assign \new_[23436]_  = \new_[23435]_  & \new_[23430]_ ;
  assign \new_[23439]_  = ~A169 & ~A170;
  assign \new_[23443]_  = A200 & ~A199;
  assign \new_[23444]_  = A168 & \new_[23443]_ ;
  assign \new_[23445]_  = \new_[23444]_  & \new_[23439]_ ;
  assign \new_[23449]_  = A265 & A202;
  assign \new_[23450]_  = A201 & \new_[23449]_ ;
  assign \new_[23454]_  = ~A299 & ~A298;
  assign \new_[23455]_  = A266 & \new_[23454]_ ;
  assign \new_[23456]_  = \new_[23455]_  & \new_[23450]_ ;
  assign \new_[23459]_  = ~A169 & ~A170;
  assign \new_[23463]_  = A200 & ~A199;
  assign \new_[23464]_  = A168 & \new_[23463]_ ;
  assign \new_[23465]_  = \new_[23464]_  & \new_[23459]_ ;
  assign \new_[23469]_  = ~A265 & A202;
  assign \new_[23470]_  = A201 & \new_[23469]_ ;
  assign \new_[23474]_  = A301 & ~A300;
  assign \new_[23475]_  = ~A266 & \new_[23474]_ ;
  assign \new_[23476]_  = \new_[23475]_  & \new_[23470]_ ;
  assign \new_[23479]_  = ~A169 & ~A170;
  assign \new_[23483]_  = A200 & ~A199;
  assign \new_[23484]_  = A168 & \new_[23483]_ ;
  assign \new_[23485]_  = \new_[23484]_  & \new_[23479]_ ;
  assign \new_[23489]_  = ~A265 & A202;
  assign \new_[23490]_  = A201 & \new_[23489]_ ;
  assign \new_[23494]_  = ~A302 & ~A300;
  assign \new_[23495]_  = ~A266 & \new_[23494]_ ;
  assign \new_[23496]_  = \new_[23495]_  & \new_[23490]_ ;
  assign \new_[23499]_  = ~A169 & ~A170;
  assign \new_[23503]_  = A200 & ~A199;
  assign \new_[23504]_  = A168 & \new_[23503]_ ;
  assign \new_[23505]_  = \new_[23504]_  & \new_[23499]_ ;
  assign \new_[23509]_  = ~A265 & A202;
  assign \new_[23510]_  = A201 & \new_[23509]_ ;
  assign \new_[23514]_  = A299 & A298;
  assign \new_[23515]_  = ~A266 & \new_[23514]_ ;
  assign \new_[23516]_  = \new_[23515]_  & \new_[23510]_ ;
  assign \new_[23519]_  = ~A169 & ~A170;
  assign \new_[23523]_  = A200 & ~A199;
  assign \new_[23524]_  = A168 & \new_[23523]_ ;
  assign \new_[23525]_  = \new_[23524]_  & \new_[23519]_ ;
  assign \new_[23529]_  = ~A265 & A202;
  assign \new_[23530]_  = A201 & \new_[23529]_ ;
  assign \new_[23534]_  = ~A299 & ~A298;
  assign \new_[23535]_  = ~A266 & \new_[23534]_ ;
  assign \new_[23536]_  = \new_[23535]_  & \new_[23530]_ ;
  assign \new_[23539]_  = ~A169 & ~A170;
  assign \new_[23543]_  = A200 & ~A199;
  assign \new_[23544]_  = A168 & \new_[23543]_ ;
  assign \new_[23545]_  = \new_[23544]_  & \new_[23539]_ ;
  assign \new_[23549]_  = ~A267 & ~A203;
  assign \new_[23550]_  = A201 & \new_[23549]_ ;
  assign \new_[23554]_  = A301 & ~A300;
  assign \new_[23555]_  = A268 & \new_[23554]_ ;
  assign \new_[23556]_  = \new_[23555]_  & \new_[23550]_ ;
  assign \new_[23559]_  = ~A169 & ~A170;
  assign \new_[23563]_  = A200 & ~A199;
  assign \new_[23564]_  = A168 & \new_[23563]_ ;
  assign \new_[23565]_  = \new_[23564]_  & \new_[23559]_ ;
  assign \new_[23569]_  = ~A267 & ~A203;
  assign \new_[23570]_  = A201 & \new_[23569]_ ;
  assign \new_[23574]_  = ~A302 & ~A300;
  assign \new_[23575]_  = A268 & \new_[23574]_ ;
  assign \new_[23576]_  = \new_[23575]_  & \new_[23570]_ ;
  assign \new_[23579]_  = ~A169 & ~A170;
  assign \new_[23583]_  = A200 & ~A199;
  assign \new_[23584]_  = A168 & \new_[23583]_ ;
  assign \new_[23585]_  = \new_[23584]_  & \new_[23579]_ ;
  assign \new_[23589]_  = ~A267 & ~A203;
  assign \new_[23590]_  = A201 & \new_[23589]_ ;
  assign \new_[23594]_  = A299 & A298;
  assign \new_[23595]_  = A268 & \new_[23594]_ ;
  assign \new_[23596]_  = \new_[23595]_  & \new_[23590]_ ;
  assign \new_[23599]_  = ~A169 & ~A170;
  assign \new_[23603]_  = A200 & ~A199;
  assign \new_[23604]_  = A168 & \new_[23603]_ ;
  assign \new_[23605]_  = \new_[23604]_  & \new_[23599]_ ;
  assign \new_[23609]_  = ~A267 & ~A203;
  assign \new_[23610]_  = A201 & \new_[23609]_ ;
  assign \new_[23614]_  = ~A299 & ~A298;
  assign \new_[23615]_  = A268 & \new_[23614]_ ;
  assign \new_[23616]_  = \new_[23615]_  & \new_[23610]_ ;
  assign \new_[23619]_  = ~A169 & ~A170;
  assign \new_[23623]_  = A200 & ~A199;
  assign \new_[23624]_  = A168 & \new_[23623]_ ;
  assign \new_[23625]_  = \new_[23624]_  & \new_[23619]_ ;
  assign \new_[23629]_  = ~A267 & ~A203;
  assign \new_[23630]_  = A201 & \new_[23629]_ ;
  assign \new_[23634]_  = A301 & ~A300;
  assign \new_[23635]_  = ~A269 & \new_[23634]_ ;
  assign \new_[23636]_  = \new_[23635]_  & \new_[23630]_ ;
  assign \new_[23639]_  = ~A169 & ~A170;
  assign \new_[23643]_  = A200 & ~A199;
  assign \new_[23644]_  = A168 & \new_[23643]_ ;
  assign \new_[23645]_  = \new_[23644]_  & \new_[23639]_ ;
  assign \new_[23649]_  = ~A267 & ~A203;
  assign \new_[23650]_  = A201 & \new_[23649]_ ;
  assign \new_[23654]_  = ~A302 & ~A300;
  assign \new_[23655]_  = ~A269 & \new_[23654]_ ;
  assign \new_[23656]_  = \new_[23655]_  & \new_[23650]_ ;
  assign \new_[23659]_  = ~A169 & ~A170;
  assign \new_[23663]_  = A200 & ~A199;
  assign \new_[23664]_  = A168 & \new_[23663]_ ;
  assign \new_[23665]_  = \new_[23664]_  & \new_[23659]_ ;
  assign \new_[23669]_  = ~A267 & ~A203;
  assign \new_[23670]_  = A201 & \new_[23669]_ ;
  assign \new_[23674]_  = A299 & A298;
  assign \new_[23675]_  = ~A269 & \new_[23674]_ ;
  assign \new_[23676]_  = \new_[23675]_  & \new_[23670]_ ;
  assign \new_[23679]_  = ~A169 & ~A170;
  assign \new_[23683]_  = A200 & ~A199;
  assign \new_[23684]_  = A168 & \new_[23683]_ ;
  assign \new_[23685]_  = \new_[23684]_  & \new_[23679]_ ;
  assign \new_[23689]_  = ~A267 & ~A203;
  assign \new_[23690]_  = A201 & \new_[23689]_ ;
  assign \new_[23694]_  = ~A299 & ~A298;
  assign \new_[23695]_  = ~A269 & \new_[23694]_ ;
  assign \new_[23696]_  = \new_[23695]_  & \new_[23690]_ ;
  assign \new_[23699]_  = ~A169 & ~A170;
  assign \new_[23703]_  = A200 & ~A199;
  assign \new_[23704]_  = A168 & \new_[23703]_ ;
  assign \new_[23705]_  = \new_[23704]_  & \new_[23699]_ ;
  assign \new_[23709]_  = A265 & ~A203;
  assign \new_[23710]_  = A201 & \new_[23709]_ ;
  assign \new_[23714]_  = A301 & ~A300;
  assign \new_[23715]_  = A266 & \new_[23714]_ ;
  assign \new_[23716]_  = \new_[23715]_  & \new_[23710]_ ;
  assign \new_[23719]_  = ~A169 & ~A170;
  assign \new_[23723]_  = A200 & ~A199;
  assign \new_[23724]_  = A168 & \new_[23723]_ ;
  assign \new_[23725]_  = \new_[23724]_  & \new_[23719]_ ;
  assign \new_[23729]_  = A265 & ~A203;
  assign \new_[23730]_  = A201 & \new_[23729]_ ;
  assign \new_[23734]_  = ~A302 & ~A300;
  assign \new_[23735]_  = A266 & \new_[23734]_ ;
  assign \new_[23736]_  = \new_[23735]_  & \new_[23730]_ ;
  assign \new_[23739]_  = ~A169 & ~A170;
  assign \new_[23743]_  = A200 & ~A199;
  assign \new_[23744]_  = A168 & \new_[23743]_ ;
  assign \new_[23745]_  = \new_[23744]_  & \new_[23739]_ ;
  assign \new_[23749]_  = A265 & ~A203;
  assign \new_[23750]_  = A201 & \new_[23749]_ ;
  assign \new_[23754]_  = A299 & A298;
  assign \new_[23755]_  = A266 & \new_[23754]_ ;
  assign \new_[23756]_  = \new_[23755]_  & \new_[23750]_ ;
  assign \new_[23759]_  = ~A169 & ~A170;
  assign \new_[23763]_  = A200 & ~A199;
  assign \new_[23764]_  = A168 & \new_[23763]_ ;
  assign \new_[23765]_  = \new_[23764]_  & \new_[23759]_ ;
  assign \new_[23769]_  = A265 & ~A203;
  assign \new_[23770]_  = A201 & \new_[23769]_ ;
  assign \new_[23774]_  = ~A299 & ~A298;
  assign \new_[23775]_  = A266 & \new_[23774]_ ;
  assign \new_[23776]_  = \new_[23775]_  & \new_[23770]_ ;
  assign \new_[23779]_  = ~A169 & ~A170;
  assign \new_[23783]_  = A200 & ~A199;
  assign \new_[23784]_  = A168 & \new_[23783]_ ;
  assign \new_[23785]_  = \new_[23784]_  & \new_[23779]_ ;
  assign \new_[23789]_  = ~A265 & ~A203;
  assign \new_[23790]_  = A201 & \new_[23789]_ ;
  assign \new_[23794]_  = A301 & ~A300;
  assign \new_[23795]_  = ~A266 & \new_[23794]_ ;
  assign \new_[23796]_  = \new_[23795]_  & \new_[23790]_ ;
  assign \new_[23799]_  = ~A169 & ~A170;
  assign \new_[23803]_  = A200 & ~A199;
  assign \new_[23804]_  = A168 & \new_[23803]_ ;
  assign \new_[23805]_  = \new_[23804]_  & \new_[23799]_ ;
  assign \new_[23809]_  = ~A265 & ~A203;
  assign \new_[23810]_  = A201 & \new_[23809]_ ;
  assign \new_[23814]_  = ~A302 & ~A300;
  assign \new_[23815]_  = ~A266 & \new_[23814]_ ;
  assign \new_[23816]_  = \new_[23815]_  & \new_[23810]_ ;
  assign \new_[23819]_  = ~A169 & ~A170;
  assign \new_[23823]_  = A200 & ~A199;
  assign \new_[23824]_  = A168 & \new_[23823]_ ;
  assign \new_[23825]_  = \new_[23824]_  & \new_[23819]_ ;
  assign \new_[23829]_  = ~A265 & ~A203;
  assign \new_[23830]_  = A201 & \new_[23829]_ ;
  assign \new_[23834]_  = A299 & A298;
  assign \new_[23835]_  = ~A266 & \new_[23834]_ ;
  assign \new_[23836]_  = \new_[23835]_  & \new_[23830]_ ;
  assign \new_[23839]_  = ~A169 & ~A170;
  assign \new_[23843]_  = A200 & ~A199;
  assign \new_[23844]_  = A168 & \new_[23843]_ ;
  assign \new_[23845]_  = \new_[23844]_  & \new_[23839]_ ;
  assign \new_[23849]_  = ~A265 & ~A203;
  assign \new_[23850]_  = A201 & \new_[23849]_ ;
  assign \new_[23854]_  = ~A299 & ~A298;
  assign \new_[23855]_  = ~A266 & \new_[23854]_ ;
  assign \new_[23856]_  = \new_[23855]_  & \new_[23850]_ ;
  assign \new_[23859]_  = ~A169 & ~A170;
  assign \new_[23863]_  = ~A200 & A199;
  assign \new_[23864]_  = A168 & \new_[23863]_ ;
  assign \new_[23865]_  = \new_[23864]_  & \new_[23859]_ ;
  assign \new_[23869]_  = ~A267 & A202;
  assign \new_[23870]_  = A201 & \new_[23869]_ ;
  assign \new_[23874]_  = A301 & ~A300;
  assign \new_[23875]_  = A268 & \new_[23874]_ ;
  assign \new_[23876]_  = \new_[23875]_  & \new_[23870]_ ;
  assign \new_[23879]_  = ~A169 & ~A170;
  assign \new_[23883]_  = ~A200 & A199;
  assign \new_[23884]_  = A168 & \new_[23883]_ ;
  assign \new_[23885]_  = \new_[23884]_  & \new_[23879]_ ;
  assign \new_[23889]_  = ~A267 & A202;
  assign \new_[23890]_  = A201 & \new_[23889]_ ;
  assign \new_[23894]_  = ~A302 & ~A300;
  assign \new_[23895]_  = A268 & \new_[23894]_ ;
  assign \new_[23896]_  = \new_[23895]_  & \new_[23890]_ ;
  assign \new_[23899]_  = ~A169 & ~A170;
  assign \new_[23903]_  = ~A200 & A199;
  assign \new_[23904]_  = A168 & \new_[23903]_ ;
  assign \new_[23905]_  = \new_[23904]_  & \new_[23899]_ ;
  assign \new_[23909]_  = ~A267 & A202;
  assign \new_[23910]_  = A201 & \new_[23909]_ ;
  assign \new_[23914]_  = A299 & A298;
  assign \new_[23915]_  = A268 & \new_[23914]_ ;
  assign \new_[23916]_  = \new_[23915]_  & \new_[23910]_ ;
  assign \new_[23919]_  = ~A169 & ~A170;
  assign \new_[23923]_  = ~A200 & A199;
  assign \new_[23924]_  = A168 & \new_[23923]_ ;
  assign \new_[23925]_  = \new_[23924]_  & \new_[23919]_ ;
  assign \new_[23929]_  = ~A267 & A202;
  assign \new_[23930]_  = A201 & \new_[23929]_ ;
  assign \new_[23934]_  = ~A299 & ~A298;
  assign \new_[23935]_  = A268 & \new_[23934]_ ;
  assign \new_[23936]_  = \new_[23935]_  & \new_[23930]_ ;
  assign \new_[23939]_  = ~A169 & ~A170;
  assign \new_[23943]_  = ~A200 & A199;
  assign \new_[23944]_  = A168 & \new_[23943]_ ;
  assign \new_[23945]_  = \new_[23944]_  & \new_[23939]_ ;
  assign \new_[23949]_  = ~A267 & A202;
  assign \new_[23950]_  = A201 & \new_[23949]_ ;
  assign \new_[23954]_  = A301 & ~A300;
  assign \new_[23955]_  = ~A269 & \new_[23954]_ ;
  assign \new_[23956]_  = \new_[23955]_  & \new_[23950]_ ;
  assign \new_[23959]_  = ~A169 & ~A170;
  assign \new_[23963]_  = ~A200 & A199;
  assign \new_[23964]_  = A168 & \new_[23963]_ ;
  assign \new_[23965]_  = \new_[23964]_  & \new_[23959]_ ;
  assign \new_[23969]_  = ~A267 & A202;
  assign \new_[23970]_  = A201 & \new_[23969]_ ;
  assign \new_[23974]_  = ~A302 & ~A300;
  assign \new_[23975]_  = ~A269 & \new_[23974]_ ;
  assign \new_[23976]_  = \new_[23975]_  & \new_[23970]_ ;
  assign \new_[23979]_  = ~A169 & ~A170;
  assign \new_[23983]_  = ~A200 & A199;
  assign \new_[23984]_  = A168 & \new_[23983]_ ;
  assign \new_[23985]_  = \new_[23984]_  & \new_[23979]_ ;
  assign \new_[23989]_  = ~A267 & A202;
  assign \new_[23990]_  = A201 & \new_[23989]_ ;
  assign \new_[23994]_  = A299 & A298;
  assign \new_[23995]_  = ~A269 & \new_[23994]_ ;
  assign \new_[23996]_  = \new_[23995]_  & \new_[23990]_ ;
  assign \new_[23999]_  = ~A169 & ~A170;
  assign \new_[24003]_  = ~A200 & A199;
  assign \new_[24004]_  = A168 & \new_[24003]_ ;
  assign \new_[24005]_  = \new_[24004]_  & \new_[23999]_ ;
  assign \new_[24009]_  = ~A267 & A202;
  assign \new_[24010]_  = A201 & \new_[24009]_ ;
  assign \new_[24014]_  = ~A299 & ~A298;
  assign \new_[24015]_  = ~A269 & \new_[24014]_ ;
  assign \new_[24016]_  = \new_[24015]_  & \new_[24010]_ ;
  assign \new_[24019]_  = ~A169 & ~A170;
  assign \new_[24023]_  = ~A200 & A199;
  assign \new_[24024]_  = A168 & \new_[24023]_ ;
  assign \new_[24025]_  = \new_[24024]_  & \new_[24019]_ ;
  assign \new_[24029]_  = A265 & A202;
  assign \new_[24030]_  = A201 & \new_[24029]_ ;
  assign \new_[24034]_  = A301 & ~A300;
  assign \new_[24035]_  = A266 & \new_[24034]_ ;
  assign \new_[24036]_  = \new_[24035]_  & \new_[24030]_ ;
  assign \new_[24039]_  = ~A169 & ~A170;
  assign \new_[24043]_  = ~A200 & A199;
  assign \new_[24044]_  = A168 & \new_[24043]_ ;
  assign \new_[24045]_  = \new_[24044]_  & \new_[24039]_ ;
  assign \new_[24049]_  = A265 & A202;
  assign \new_[24050]_  = A201 & \new_[24049]_ ;
  assign \new_[24054]_  = ~A302 & ~A300;
  assign \new_[24055]_  = A266 & \new_[24054]_ ;
  assign \new_[24056]_  = \new_[24055]_  & \new_[24050]_ ;
  assign \new_[24059]_  = ~A169 & ~A170;
  assign \new_[24063]_  = ~A200 & A199;
  assign \new_[24064]_  = A168 & \new_[24063]_ ;
  assign \new_[24065]_  = \new_[24064]_  & \new_[24059]_ ;
  assign \new_[24069]_  = A265 & A202;
  assign \new_[24070]_  = A201 & \new_[24069]_ ;
  assign \new_[24074]_  = A299 & A298;
  assign \new_[24075]_  = A266 & \new_[24074]_ ;
  assign \new_[24076]_  = \new_[24075]_  & \new_[24070]_ ;
  assign \new_[24079]_  = ~A169 & ~A170;
  assign \new_[24083]_  = ~A200 & A199;
  assign \new_[24084]_  = A168 & \new_[24083]_ ;
  assign \new_[24085]_  = \new_[24084]_  & \new_[24079]_ ;
  assign \new_[24089]_  = A265 & A202;
  assign \new_[24090]_  = A201 & \new_[24089]_ ;
  assign \new_[24094]_  = ~A299 & ~A298;
  assign \new_[24095]_  = A266 & \new_[24094]_ ;
  assign \new_[24096]_  = \new_[24095]_  & \new_[24090]_ ;
  assign \new_[24099]_  = ~A169 & ~A170;
  assign \new_[24103]_  = ~A200 & A199;
  assign \new_[24104]_  = A168 & \new_[24103]_ ;
  assign \new_[24105]_  = \new_[24104]_  & \new_[24099]_ ;
  assign \new_[24109]_  = ~A265 & A202;
  assign \new_[24110]_  = A201 & \new_[24109]_ ;
  assign \new_[24114]_  = A301 & ~A300;
  assign \new_[24115]_  = ~A266 & \new_[24114]_ ;
  assign \new_[24116]_  = \new_[24115]_  & \new_[24110]_ ;
  assign \new_[24119]_  = ~A169 & ~A170;
  assign \new_[24123]_  = ~A200 & A199;
  assign \new_[24124]_  = A168 & \new_[24123]_ ;
  assign \new_[24125]_  = \new_[24124]_  & \new_[24119]_ ;
  assign \new_[24129]_  = ~A265 & A202;
  assign \new_[24130]_  = A201 & \new_[24129]_ ;
  assign \new_[24134]_  = ~A302 & ~A300;
  assign \new_[24135]_  = ~A266 & \new_[24134]_ ;
  assign \new_[24136]_  = \new_[24135]_  & \new_[24130]_ ;
  assign \new_[24139]_  = ~A169 & ~A170;
  assign \new_[24143]_  = ~A200 & A199;
  assign \new_[24144]_  = A168 & \new_[24143]_ ;
  assign \new_[24145]_  = \new_[24144]_  & \new_[24139]_ ;
  assign \new_[24149]_  = ~A265 & A202;
  assign \new_[24150]_  = A201 & \new_[24149]_ ;
  assign \new_[24154]_  = A299 & A298;
  assign \new_[24155]_  = ~A266 & \new_[24154]_ ;
  assign \new_[24156]_  = \new_[24155]_  & \new_[24150]_ ;
  assign \new_[24159]_  = ~A169 & ~A170;
  assign \new_[24163]_  = ~A200 & A199;
  assign \new_[24164]_  = A168 & \new_[24163]_ ;
  assign \new_[24165]_  = \new_[24164]_  & \new_[24159]_ ;
  assign \new_[24169]_  = ~A265 & A202;
  assign \new_[24170]_  = A201 & \new_[24169]_ ;
  assign \new_[24174]_  = ~A299 & ~A298;
  assign \new_[24175]_  = ~A266 & \new_[24174]_ ;
  assign \new_[24176]_  = \new_[24175]_  & \new_[24170]_ ;
  assign \new_[24179]_  = ~A169 & ~A170;
  assign \new_[24183]_  = ~A200 & A199;
  assign \new_[24184]_  = A168 & \new_[24183]_ ;
  assign \new_[24185]_  = \new_[24184]_  & \new_[24179]_ ;
  assign \new_[24189]_  = ~A267 & ~A203;
  assign \new_[24190]_  = A201 & \new_[24189]_ ;
  assign \new_[24194]_  = A301 & ~A300;
  assign \new_[24195]_  = A268 & \new_[24194]_ ;
  assign \new_[24196]_  = \new_[24195]_  & \new_[24190]_ ;
  assign \new_[24199]_  = ~A169 & ~A170;
  assign \new_[24203]_  = ~A200 & A199;
  assign \new_[24204]_  = A168 & \new_[24203]_ ;
  assign \new_[24205]_  = \new_[24204]_  & \new_[24199]_ ;
  assign \new_[24209]_  = ~A267 & ~A203;
  assign \new_[24210]_  = A201 & \new_[24209]_ ;
  assign \new_[24214]_  = ~A302 & ~A300;
  assign \new_[24215]_  = A268 & \new_[24214]_ ;
  assign \new_[24216]_  = \new_[24215]_  & \new_[24210]_ ;
  assign \new_[24219]_  = ~A169 & ~A170;
  assign \new_[24223]_  = ~A200 & A199;
  assign \new_[24224]_  = A168 & \new_[24223]_ ;
  assign \new_[24225]_  = \new_[24224]_  & \new_[24219]_ ;
  assign \new_[24229]_  = ~A267 & ~A203;
  assign \new_[24230]_  = A201 & \new_[24229]_ ;
  assign \new_[24234]_  = A299 & A298;
  assign \new_[24235]_  = A268 & \new_[24234]_ ;
  assign \new_[24236]_  = \new_[24235]_  & \new_[24230]_ ;
  assign \new_[24239]_  = ~A169 & ~A170;
  assign \new_[24243]_  = ~A200 & A199;
  assign \new_[24244]_  = A168 & \new_[24243]_ ;
  assign \new_[24245]_  = \new_[24244]_  & \new_[24239]_ ;
  assign \new_[24249]_  = ~A267 & ~A203;
  assign \new_[24250]_  = A201 & \new_[24249]_ ;
  assign \new_[24254]_  = ~A299 & ~A298;
  assign \new_[24255]_  = A268 & \new_[24254]_ ;
  assign \new_[24256]_  = \new_[24255]_  & \new_[24250]_ ;
  assign \new_[24259]_  = ~A169 & ~A170;
  assign \new_[24263]_  = ~A200 & A199;
  assign \new_[24264]_  = A168 & \new_[24263]_ ;
  assign \new_[24265]_  = \new_[24264]_  & \new_[24259]_ ;
  assign \new_[24269]_  = ~A267 & ~A203;
  assign \new_[24270]_  = A201 & \new_[24269]_ ;
  assign \new_[24274]_  = A301 & ~A300;
  assign \new_[24275]_  = ~A269 & \new_[24274]_ ;
  assign \new_[24276]_  = \new_[24275]_  & \new_[24270]_ ;
  assign \new_[24279]_  = ~A169 & ~A170;
  assign \new_[24283]_  = ~A200 & A199;
  assign \new_[24284]_  = A168 & \new_[24283]_ ;
  assign \new_[24285]_  = \new_[24284]_  & \new_[24279]_ ;
  assign \new_[24289]_  = ~A267 & ~A203;
  assign \new_[24290]_  = A201 & \new_[24289]_ ;
  assign \new_[24294]_  = ~A302 & ~A300;
  assign \new_[24295]_  = ~A269 & \new_[24294]_ ;
  assign \new_[24296]_  = \new_[24295]_  & \new_[24290]_ ;
  assign \new_[24299]_  = ~A169 & ~A170;
  assign \new_[24303]_  = ~A200 & A199;
  assign \new_[24304]_  = A168 & \new_[24303]_ ;
  assign \new_[24305]_  = \new_[24304]_  & \new_[24299]_ ;
  assign \new_[24309]_  = ~A267 & ~A203;
  assign \new_[24310]_  = A201 & \new_[24309]_ ;
  assign \new_[24314]_  = A299 & A298;
  assign \new_[24315]_  = ~A269 & \new_[24314]_ ;
  assign \new_[24316]_  = \new_[24315]_  & \new_[24310]_ ;
  assign \new_[24319]_  = ~A169 & ~A170;
  assign \new_[24323]_  = ~A200 & A199;
  assign \new_[24324]_  = A168 & \new_[24323]_ ;
  assign \new_[24325]_  = \new_[24324]_  & \new_[24319]_ ;
  assign \new_[24329]_  = ~A267 & ~A203;
  assign \new_[24330]_  = A201 & \new_[24329]_ ;
  assign \new_[24334]_  = ~A299 & ~A298;
  assign \new_[24335]_  = ~A269 & \new_[24334]_ ;
  assign \new_[24336]_  = \new_[24335]_  & \new_[24330]_ ;
  assign \new_[24339]_  = ~A169 & ~A170;
  assign \new_[24343]_  = ~A200 & A199;
  assign \new_[24344]_  = A168 & \new_[24343]_ ;
  assign \new_[24345]_  = \new_[24344]_  & \new_[24339]_ ;
  assign \new_[24349]_  = A265 & ~A203;
  assign \new_[24350]_  = A201 & \new_[24349]_ ;
  assign \new_[24354]_  = A301 & ~A300;
  assign \new_[24355]_  = A266 & \new_[24354]_ ;
  assign \new_[24356]_  = \new_[24355]_  & \new_[24350]_ ;
  assign \new_[24359]_  = ~A169 & ~A170;
  assign \new_[24363]_  = ~A200 & A199;
  assign \new_[24364]_  = A168 & \new_[24363]_ ;
  assign \new_[24365]_  = \new_[24364]_  & \new_[24359]_ ;
  assign \new_[24369]_  = A265 & ~A203;
  assign \new_[24370]_  = A201 & \new_[24369]_ ;
  assign \new_[24374]_  = ~A302 & ~A300;
  assign \new_[24375]_  = A266 & \new_[24374]_ ;
  assign \new_[24376]_  = \new_[24375]_  & \new_[24370]_ ;
  assign \new_[24379]_  = ~A169 & ~A170;
  assign \new_[24383]_  = ~A200 & A199;
  assign \new_[24384]_  = A168 & \new_[24383]_ ;
  assign \new_[24385]_  = \new_[24384]_  & \new_[24379]_ ;
  assign \new_[24389]_  = A265 & ~A203;
  assign \new_[24390]_  = A201 & \new_[24389]_ ;
  assign \new_[24394]_  = A299 & A298;
  assign \new_[24395]_  = A266 & \new_[24394]_ ;
  assign \new_[24396]_  = \new_[24395]_  & \new_[24390]_ ;
  assign \new_[24399]_  = ~A169 & ~A170;
  assign \new_[24403]_  = ~A200 & A199;
  assign \new_[24404]_  = A168 & \new_[24403]_ ;
  assign \new_[24405]_  = \new_[24404]_  & \new_[24399]_ ;
  assign \new_[24409]_  = A265 & ~A203;
  assign \new_[24410]_  = A201 & \new_[24409]_ ;
  assign \new_[24414]_  = ~A299 & ~A298;
  assign \new_[24415]_  = A266 & \new_[24414]_ ;
  assign \new_[24416]_  = \new_[24415]_  & \new_[24410]_ ;
  assign \new_[24419]_  = ~A169 & ~A170;
  assign \new_[24423]_  = ~A200 & A199;
  assign \new_[24424]_  = A168 & \new_[24423]_ ;
  assign \new_[24425]_  = \new_[24424]_  & \new_[24419]_ ;
  assign \new_[24429]_  = ~A265 & ~A203;
  assign \new_[24430]_  = A201 & \new_[24429]_ ;
  assign \new_[24434]_  = A301 & ~A300;
  assign \new_[24435]_  = ~A266 & \new_[24434]_ ;
  assign \new_[24436]_  = \new_[24435]_  & \new_[24430]_ ;
  assign \new_[24439]_  = ~A169 & ~A170;
  assign \new_[24443]_  = ~A200 & A199;
  assign \new_[24444]_  = A168 & \new_[24443]_ ;
  assign \new_[24445]_  = \new_[24444]_  & \new_[24439]_ ;
  assign \new_[24449]_  = ~A265 & ~A203;
  assign \new_[24450]_  = A201 & \new_[24449]_ ;
  assign \new_[24454]_  = ~A302 & ~A300;
  assign \new_[24455]_  = ~A266 & \new_[24454]_ ;
  assign \new_[24456]_  = \new_[24455]_  & \new_[24450]_ ;
  assign \new_[24459]_  = ~A169 & ~A170;
  assign \new_[24463]_  = ~A200 & A199;
  assign \new_[24464]_  = A168 & \new_[24463]_ ;
  assign \new_[24465]_  = \new_[24464]_  & \new_[24459]_ ;
  assign \new_[24469]_  = ~A265 & ~A203;
  assign \new_[24470]_  = A201 & \new_[24469]_ ;
  assign \new_[24474]_  = A299 & A298;
  assign \new_[24475]_  = ~A266 & \new_[24474]_ ;
  assign \new_[24476]_  = \new_[24475]_  & \new_[24470]_ ;
  assign \new_[24479]_  = ~A169 & ~A170;
  assign \new_[24483]_  = ~A200 & A199;
  assign \new_[24484]_  = A168 & \new_[24483]_ ;
  assign \new_[24485]_  = \new_[24484]_  & \new_[24479]_ ;
  assign \new_[24489]_  = ~A265 & ~A203;
  assign \new_[24490]_  = A201 & \new_[24489]_ ;
  assign \new_[24494]_  = ~A299 & ~A298;
  assign \new_[24495]_  = ~A266 & \new_[24494]_ ;
  assign \new_[24496]_  = \new_[24495]_  & \new_[24490]_ ;
  assign \new_[24500]_  = A202 & A200;
  assign \new_[24501]_  = ~A199 & \new_[24500]_ ;
  assign \new_[24505]_  = A234 & A233;
  assign \new_[24506]_  = ~A232 & \new_[24505]_ ;
  assign \new_[24507]_  = \new_[24506]_  & \new_[24501]_ ;
  assign \new_[24511]_  = A266 & ~A265;
  assign \new_[24512]_  = A235 & \new_[24511]_ ;
  assign \new_[24516]_  = A269 & ~A268;
  assign \new_[24517]_  = ~A267 & \new_[24516]_ ;
  assign \new_[24518]_  = \new_[24517]_  & \new_[24512]_ ;
  assign \new_[24522]_  = A202 & A200;
  assign \new_[24523]_  = ~A199 & \new_[24522]_ ;
  assign \new_[24527]_  = A234 & A233;
  assign \new_[24528]_  = ~A232 & \new_[24527]_ ;
  assign \new_[24529]_  = \new_[24528]_  & \new_[24523]_ ;
  assign \new_[24533]_  = ~A266 & A265;
  assign \new_[24534]_  = A235 & \new_[24533]_ ;
  assign \new_[24538]_  = A269 & ~A268;
  assign \new_[24539]_  = ~A267 & \new_[24538]_ ;
  assign \new_[24540]_  = \new_[24539]_  & \new_[24534]_ ;
  assign \new_[24544]_  = A202 & A200;
  assign \new_[24545]_  = ~A199 & \new_[24544]_ ;
  assign \new_[24549]_  = A234 & A233;
  assign \new_[24550]_  = ~A232 & \new_[24549]_ ;
  assign \new_[24551]_  = \new_[24550]_  & \new_[24545]_ ;
  assign \new_[24555]_  = A266 & ~A265;
  assign \new_[24556]_  = ~A236 & \new_[24555]_ ;
  assign \new_[24560]_  = A269 & ~A268;
  assign \new_[24561]_  = ~A267 & \new_[24560]_ ;
  assign \new_[24562]_  = \new_[24561]_  & \new_[24556]_ ;
  assign \new_[24566]_  = A202 & A200;
  assign \new_[24567]_  = ~A199 & \new_[24566]_ ;
  assign \new_[24571]_  = A234 & A233;
  assign \new_[24572]_  = ~A232 & \new_[24571]_ ;
  assign \new_[24573]_  = \new_[24572]_  & \new_[24567]_ ;
  assign \new_[24577]_  = ~A266 & A265;
  assign \new_[24578]_  = ~A236 & \new_[24577]_ ;
  assign \new_[24582]_  = A269 & ~A268;
  assign \new_[24583]_  = ~A267 & \new_[24582]_ ;
  assign \new_[24584]_  = \new_[24583]_  & \new_[24578]_ ;
  assign \new_[24588]_  = A202 & A200;
  assign \new_[24589]_  = ~A199 & \new_[24588]_ ;
  assign \new_[24593]_  = A234 & ~A233;
  assign \new_[24594]_  = A232 & \new_[24593]_ ;
  assign \new_[24595]_  = \new_[24594]_  & \new_[24589]_ ;
  assign \new_[24599]_  = A266 & ~A265;
  assign \new_[24600]_  = A235 & \new_[24599]_ ;
  assign \new_[24604]_  = A269 & ~A268;
  assign \new_[24605]_  = ~A267 & \new_[24604]_ ;
  assign \new_[24606]_  = \new_[24605]_  & \new_[24600]_ ;
  assign \new_[24610]_  = A202 & A200;
  assign \new_[24611]_  = ~A199 & \new_[24610]_ ;
  assign \new_[24615]_  = A234 & ~A233;
  assign \new_[24616]_  = A232 & \new_[24615]_ ;
  assign \new_[24617]_  = \new_[24616]_  & \new_[24611]_ ;
  assign \new_[24621]_  = ~A266 & A265;
  assign \new_[24622]_  = A235 & \new_[24621]_ ;
  assign \new_[24626]_  = A269 & ~A268;
  assign \new_[24627]_  = ~A267 & \new_[24626]_ ;
  assign \new_[24628]_  = \new_[24627]_  & \new_[24622]_ ;
  assign \new_[24632]_  = A202 & A200;
  assign \new_[24633]_  = ~A199 & \new_[24632]_ ;
  assign \new_[24637]_  = A234 & ~A233;
  assign \new_[24638]_  = A232 & \new_[24637]_ ;
  assign \new_[24639]_  = \new_[24638]_  & \new_[24633]_ ;
  assign \new_[24643]_  = A266 & ~A265;
  assign \new_[24644]_  = ~A236 & \new_[24643]_ ;
  assign \new_[24648]_  = A269 & ~A268;
  assign \new_[24649]_  = ~A267 & \new_[24648]_ ;
  assign \new_[24650]_  = \new_[24649]_  & \new_[24644]_ ;
  assign \new_[24654]_  = A202 & A200;
  assign \new_[24655]_  = ~A199 & \new_[24654]_ ;
  assign \new_[24659]_  = A234 & ~A233;
  assign \new_[24660]_  = A232 & \new_[24659]_ ;
  assign \new_[24661]_  = \new_[24660]_  & \new_[24655]_ ;
  assign \new_[24665]_  = ~A266 & A265;
  assign \new_[24666]_  = ~A236 & \new_[24665]_ ;
  assign \new_[24670]_  = A269 & ~A268;
  assign \new_[24671]_  = ~A267 & \new_[24670]_ ;
  assign \new_[24672]_  = \new_[24671]_  & \new_[24666]_ ;
  assign \new_[24676]_  = ~A203 & A200;
  assign \new_[24677]_  = ~A199 & \new_[24676]_ ;
  assign \new_[24681]_  = A234 & A233;
  assign \new_[24682]_  = ~A232 & \new_[24681]_ ;
  assign \new_[24683]_  = \new_[24682]_  & \new_[24677]_ ;
  assign \new_[24687]_  = A266 & ~A265;
  assign \new_[24688]_  = A235 & \new_[24687]_ ;
  assign \new_[24692]_  = A269 & ~A268;
  assign \new_[24693]_  = ~A267 & \new_[24692]_ ;
  assign \new_[24694]_  = \new_[24693]_  & \new_[24688]_ ;
  assign \new_[24698]_  = ~A203 & A200;
  assign \new_[24699]_  = ~A199 & \new_[24698]_ ;
  assign \new_[24703]_  = A234 & A233;
  assign \new_[24704]_  = ~A232 & \new_[24703]_ ;
  assign \new_[24705]_  = \new_[24704]_  & \new_[24699]_ ;
  assign \new_[24709]_  = ~A266 & A265;
  assign \new_[24710]_  = A235 & \new_[24709]_ ;
  assign \new_[24714]_  = A269 & ~A268;
  assign \new_[24715]_  = ~A267 & \new_[24714]_ ;
  assign \new_[24716]_  = \new_[24715]_  & \new_[24710]_ ;
  assign \new_[24720]_  = ~A203 & A200;
  assign \new_[24721]_  = ~A199 & \new_[24720]_ ;
  assign \new_[24725]_  = A234 & A233;
  assign \new_[24726]_  = ~A232 & \new_[24725]_ ;
  assign \new_[24727]_  = \new_[24726]_  & \new_[24721]_ ;
  assign \new_[24731]_  = A266 & ~A265;
  assign \new_[24732]_  = ~A236 & \new_[24731]_ ;
  assign \new_[24736]_  = A269 & ~A268;
  assign \new_[24737]_  = ~A267 & \new_[24736]_ ;
  assign \new_[24738]_  = \new_[24737]_  & \new_[24732]_ ;
  assign \new_[24742]_  = ~A203 & A200;
  assign \new_[24743]_  = ~A199 & \new_[24742]_ ;
  assign \new_[24747]_  = A234 & A233;
  assign \new_[24748]_  = ~A232 & \new_[24747]_ ;
  assign \new_[24749]_  = \new_[24748]_  & \new_[24743]_ ;
  assign \new_[24753]_  = ~A266 & A265;
  assign \new_[24754]_  = ~A236 & \new_[24753]_ ;
  assign \new_[24758]_  = A269 & ~A268;
  assign \new_[24759]_  = ~A267 & \new_[24758]_ ;
  assign \new_[24760]_  = \new_[24759]_  & \new_[24754]_ ;
  assign \new_[24764]_  = ~A203 & A200;
  assign \new_[24765]_  = ~A199 & \new_[24764]_ ;
  assign \new_[24769]_  = A234 & ~A233;
  assign \new_[24770]_  = A232 & \new_[24769]_ ;
  assign \new_[24771]_  = \new_[24770]_  & \new_[24765]_ ;
  assign \new_[24775]_  = A266 & ~A265;
  assign \new_[24776]_  = A235 & \new_[24775]_ ;
  assign \new_[24780]_  = A269 & ~A268;
  assign \new_[24781]_  = ~A267 & \new_[24780]_ ;
  assign \new_[24782]_  = \new_[24781]_  & \new_[24776]_ ;
  assign \new_[24786]_  = ~A203 & A200;
  assign \new_[24787]_  = ~A199 & \new_[24786]_ ;
  assign \new_[24791]_  = A234 & ~A233;
  assign \new_[24792]_  = A232 & \new_[24791]_ ;
  assign \new_[24793]_  = \new_[24792]_  & \new_[24787]_ ;
  assign \new_[24797]_  = ~A266 & A265;
  assign \new_[24798]_  = A235 & \new_[24797]_ ;
  assign \new_[24802]_  = A269 & ~A268;
  assign \new_[24803]_  = ~A267 & \new_[24802]_ ;
  assign \new_[24804]_  = \new_[24803]_  & \new_[24798]_ ;
  assign \new_[24808]_  = ~A203 & A200;
  assign \new_[24809]_  = ~A199 & \new_[24808]_ ;
  assign \new_[24813]_  = A234 & ~A233;
  assign \new_[24814]_  = A232 & \new_[24813]_ ;
  assign \new_[24815]_  = \new_[24814]_  & \new_[24809]_ ;
  assign \new_[24819]_  = A266 & ~A265;
  assign \new_[24820]_  = ~A236 & \new_[24819]_ ;
  assign \new_[24824]_  = A269 & ~A268;
  assign \new_[24825]_  = ~A267 & \new_[24824]_ ;
  assign \new_[24826]_  = \new_[24825]_  & \new_[24820]_ ;
  assign \new_[24830]_  = ~A203 & A200;
  assign \new_[24831]_  = ~A199 & \new_[24830]_ ;
  assign \new_[24835]_  = A234 & ~A233;
  assign \new_[24836]_  = A232 & \new_[24835]_ ;
  assign \new_[24837]_  = \new_[24836]_  & \new_[24831]_ ;
  assign \new_[24841]_  = ~A266 & A265;
  assign \new_[24842]_  = ~A236 & \new_[24841]_ ;
  assign \new_[24846]_  = A269 & ~A268;
  assign \new_[24847]_  = ~A267 & \new_[24846]_ ;
  assign \new_[24848]_  = \new_[24847]_  & \new_[24842]_ ;
  assign \new_[24852]_  = A202 & ~A200;
  assign \new_[24853]_  = A199 & \new_[24852]_ ;
  assign \new_[24857]_  = A234 & A233;
  assign \new_[24858]_  = ~A232 & \new_[24857]_ ;
  assign \new_[24859]_  = \new_[24858]_  & \new_[24853]_ ;
  assign \new_[24863]_  = A266 & ~A265;
  assign \new_[24864]_  = A235 & \new_[24863]_ ;
  assign \new_[24868]_  = A269 & ~A268;
  assign \new_[24869]_  = ~A267 & \new_[24868]_ ;
  assign \new_[24870]_  = \new_[24869]_  & \new_[24864]_ ;
  assign \new_[24874]_  = A202 & ~A200;
  assign \new_[24875]_  = A199 & \new_[24874]_ ;
  assign \new_[24879]_  = A234 & A233;
  assign \new_[24880]_  = ~A232 & \new_[24879]_ ;
  assign \new_[24881]_  = \new_[24880]_  & \new_[24875]_ ;
  assign \new_[24885]_  = ~A266 & A265;
  assign \new_[24886]_  = A235 & \new_[24885]_ ;
  assign \new_[24890]_  = A269 & ~A268;
  assign \new_[24891]_  = ~A267 & \new_[24890]_ ;
  assign \new_[24892]_  = \new_[24891]_  & \new_[24886]_ ;
  assign \new_[24896]_  = A202 & ~A200;
  assign \new_[24897]_  = A199 & \new_[24896]_ ;
  assign \new_[24901]_  = A234 & A233;
  assign \new_[24902]_  = ~A232 & \new_[24901]_ ;
  assign \new_[24903]_  = \new_[24902]_  & \new_[24897]_ ;
  assign \new_[24907]_  = A266 & ~A265;
  assign \new_[24908]_  = ~A236 & \new_[24907]_ ;
  assign \new_[24912]_  = A269 & ~A268;
  assign \new_[24913]_  = ~A267 & \new_[24912]_ ;
  assign \new_[24914]_  = \new_[24913]_  & \new_[24908]_ ;
  assign \new_[24918]_  = A202 & ~A200;
  assign \new_[24919]_  = A199 & \new_[24918]_ ;
  assign \new_[24923]_  = A234 & A233;
  assign \new_[24924]_  = ~A232 & \new_[24923]_ ;
  assign \new_[24925]_  = \new_[24924]_  & \new_[24919]_ ;
  assign \new_[24929]_  = ~A266 & A265;
  assign \new_[24930]_  = ~A236 & \new_[24929]_ ;
  assign \new_[24934]_  = A269 & ~A268;
  assign \new_[24935]_  = ~A267 & \new_[24934]_ ;
  assign \new_[24936]_  = \new_[24935]_  & \new_[24930]_ ;
  assign \new_[24940]_  = A202 & ~A200;
  assign \new_[24941]_  = A199 & \new_[24940]_ ;
  assign \new_[24945]_  = A234 & ~A233;
  assign \new_[24946]_  = A232 & \new_[24945]_ ;
  assign \new_[24947]_  = \new_[24946]_  & \new_[24941]_ ;
  assign \new_[24951]_  = A266 & ~A265;
  assign \new_[24952]_  = A235 & \new_[24951]_ ;
  assign \new_[24956]_  = A269 & ~A268;
  assign \new_[24957]_  = ~A267 & \new_[24956]_ ;
  assign \new_[24958]_  = \new_[24957]_  & \new_[24952]_ ;
  assign \new_[24962]_  = A202 & ~A200;
  assign \new_[24963]_  = A199 & \new_[24962]_ ;
  assign \new_[24967]_  = A234 & ~A233;
  assign \new_[24968]_  = A232 & \new_[24967]_ ;
  assign \new_[24969]_  = \new_[24968]_  & \new_[24963]_ ;
  assign \new_[24973]_  = ~A266 & A265;
  assign \new_[24974]_  = A235 & \new_[24973]_ ;
  assign \new_[24978]_  = A269 & ~A268;
  assign \new_[24979]_  = ~A267 & \new_[24978]_ ;
  assign \new_[24980]_  = \new_[24979]_  & \new_[24974]_ ;
  assign \new_[24984]_  = A202 & ~A200;
  assign \new_[24985]_  = A199 & \new_[24984]_ ;
  assign \new_[24989]_  = A234 & ~A233;
  assign \new_[24990]_  = A232 & \new_[24989]_ ;
  assign \new_[24991]_  = \new_[24990]_  & \new_[24985]_ ;
  assign \new_[24995]_  = A266 & ~A265;
  assign \new_[24996]_  = ~A236 & \new_[24995]_ ;
  assign \new_[25000]_  = A269 & ~A268;
  assign \new_[25001]_  = ~A267 & \new_[25000]_ ;
  assign \new_[25002]_  = \new_[25001]_  & \new_[24996]_ ;
  assign \new_[25006]_  = A202 & ~A200;
  assign \new_[25007]_  = A199 & \new_[25006]_ ;
  assign \new_[25011]_  = A234 & ~A233;
  assign \new_[25012]_  = A232 & \new_[25011]_ ;
  assign \new_[25013]_  = \new_[25012]_  & \new_[25007]_ ;
  assign \new_[25017]_  = ~A266 & A265;
  assign \new_[25018]_  = ~A236 & \new_[25017]_ ;
  assign \new_[25022]_  = A269 & ~A268;
  assign \new_[25023]_  = ~A267 & \new_[25022]_ ;
  assign \new_[25024]_  = \new_[25023]_  & \new_[25018]_ ;
  assign \new_[25028]_  = ~A203 & ~A200;
  assign \new_[25029]_  = A199 & \new_[25028]_ ;
  assign \new_[25033]_  = A234 & A233;
  assign \new_[25034]_  = ~A232 & \new_[25033]_ ;
  assign \new_[25035]_  = \new_[25034]_  & \new_[25029]_ ;
  assign \new_[25039]_  = A266 & ~A265;
  assign \new_[25040]_  = A235 & \new_[25039]_ ;
  assign \new_[25044]_  = A269 & ~A268;
  assign \new_[25045]_  = ~A267 & \new_[25044]_ ;
  assign \new_[25046]_  = \new_[25045]_  & \new_[25040]_ ;
  assign \new_[25050]_  = ~A203 & ~A200;
  assign \new_[25051]_  = A199 & \new_[25050]_ ;
  assign \new_[25055]_  = A234 & A233;
  assign \new_[25056]_  = ~A232 & \new_[25055]_ ;
  assign \new_[25057]_  = \new_[25056]_  & \new_[25051]_ ;
  assign \new_[25061]_  = ~A266 & A265;
  assign \new_[25062]_  = A235 & \new_[25061]_ ;
  assign \new_[25066]_  = A269 & ~A268;
  assign \new_[25067]_  = ~A267 & \new_[25066]_ ;
  assign \new_[25068]_  = \new_[25067]_  & \new_[25062]_ ;
  assign \new_[25072]_  = ~A203 & ~A200;
  assign \new_[25073]_  = A199 & \new_[25072]_ ;
  assign \new_[25077]_  = A234 & A233;
  assign \new_[25078]_  = ~A232 & \new_[25077]_ ;
  assign \new_[25079]_  = \new_[25078]_  & \new_[25073]_ ;
  assign \new_[25083]_  = A266 & ~A265;
  assign \new_[25084]_  = ~A236 & \new_[25083]_ ;
  assign \new_[25088]_  = A269 & ~A268;
  assign \new_[25089]_  = ~A267 & \new_[25088]_ ;
  assign \new_[25090]_  = \new_[25089]_  & \new_[25084]_ ;
  assign \new_[25094]_  = ~A203 & ~A200;
  assign \new_[25095]_  = A199 & \new_[25094]_ ;
  assign \new_[25099]_  = A234 & A233;
  assign \new_[25100]_  = ~A232 & \new_[25099]_ ;
  assign \new_[25101]_  = \new_[25100]_  & \new_[25095]_ ;
  assign \new_[25105]_  = ~A266 & A265;
  assign \new_[25106]_  = ~A236 & \new_[25105]_ ;
  assign \new_[25110]_  = A269 & ~A268;
  assign \new_[25111]_  = ~A267 & \new_[25110]_ ;
  assign \new_[25112]_  = \new_[25111]_  & \new_[25106]_ ;
  assign \new_[25116]_  = ~A203 & ~A200;
  assign \new_[25117]_  = A199 & \new_[25116]_ ;
  assign \new_[25121]_  = A234 & ~A233;
  assign \new_[25122]_  = A232 & \new_[25121]_ ;
  assign \new_[25123]_  = \new_[25122]_  & \new_[25117]_ ;
  assign \new_[25127]_  = A266 & ~A265;
  assign \new_[25128]_  = A235 & \new_[25127]_ ;
  assign \new_[25132]_  = A269 & ~A268;
  assign \new_[25133]_  = ~A267 & \new_[25132]_ ;
  assign \new_[25134]_  = \new_[25133]_  & \new_[25128]_ ;
  assign \new_[25138]_  = ~A203 & ~A200;
  assign \new_[25139]_  = A199 & \new_[25138]_ ;
  assign \new_[25143]_  = A234 & ~A233;
  assign \new_[25144]_  = A232 & \new_[25143]_ ;
  assign \new_[25145]_  = \new_[25144]_  & \new_[25139]_ ;
  assign \new_[25149]_  = ~A266 & A265;
  assign \new_[25150]_  = A235 & \new_[25149]_ ;
  assign \new_[25154]_  = A269 & ~A268;
  assign \new_[25155]_  = ~A267 & \new_[25154]_ ;
  assign \new_[25156]_  = \new_[25155]_  & \new_[25150]_ ;
  assign \new_[25160]_  = ~A203 & ~A200;
  assign \new_[25161]_  = A199 & \new_[25160]_ ;
  assign \new_[25165]_  = A234 & ~A233;
  assign \new_[25166]_  = A232 & \new_[25165]_ ;
  assign \new_[25167]_  = \new_[25166]_  & \new_[25161]_ ;
  assign \new_[25171]_  = A266 & ~A265;
  assign \new_[25172]_  = ~A236 & \new_[25171]_ ;
  assign \new_[25176]_  = A269 & ~A268;
  assign \new_[25177]_  = ~A267 & \new_[25176]_ ;
  assign \new_[25178]_  = \new_[25177]_  & \new_[25172]_ ;
  assign \new_[25182]_  = ~A203 & ~A200;
  assign \new_[25183]_  = A199 & \new_[25182]_ ;
  assign \new_[25187]_  = A234 & ~A233;
  assign \new_[25188]_  = A232 & \new_[25187]_ ;
  assign \new_[25189]_  = \new_[25188]_  & \new_[25183]_ ;
  assign \new_[25193]_  = ~A266 & A265;
  assign \new_[25194]_  = ~A236 & \new_[25193]_ ;
  assign \new_[25198]_  = A269 & ~A268;
  assign \new_[25199]_  = ~A267 & \new_[25198]_ ;
  assign \new_[25200]_  = \new_[25199]_  & \new_[25194]_ ;
  assign \new_[25204]_  = ~A232 & A166;
  assign \new_[25205]_  = A167 & \new_[25204]_ ;
  assign \new_[25209]_  = ~A235 & ~A234;
  assign \new_[25210]_  = A233 & \new_[25209]_ ;
  assign \new_[25211]_  = \new_[25210]_  & \new_[25205]_ ;
  assign \new_[25215]_  = A266 & ~A265;
  assign \new_[25216]_  = A236 & \new_[25215]_ ;
  assign \new_[25220]_  = A269 & ~A268;
  assign \new_[25221]_  = ~A267 & \new_[25220]_ ;
  assign \new_[25222]_  = \new_[25221]_  & \new_[25216]_ ;
  assign \new_[25226]_  = ~A232 & A166;
  assign \new_[25227]_  = A167 & \new_[25226]_ ;
  assign \new_[25231]_  = ~A235 & ~A234;
  assign \new_[25232]_  = A233 & \new_[25231]_ ;
  assign \new_[25233]_  = \new_[25232]_  & \new_[25227]_ ;
  assign \new_[25237]_  = ~A266 & A265;
  assign \new_[25238]_  = A236 & \new_[25237]_ ;
  assign \new_[25242]_  = A269 & ~A268;
  assign \new_[25243]_  = ~A267 & \new_[25242]_ ;
  assign \new_[25244]_  = \new_[25243]_  & \new_[25238]_ ;
  assign \new_[25248]_  = A232 & A166;
  assign \new_[25249]_  = A167 & \new_[25248]_ ;
  assign \new_[25253]_  = ~A235 & ~A234;
  assign \new_[25254]_  = ~A233 & \new_[25253]_ ;
  assign \new_[25255]_  = \new_[25254]_  & \new_[25249]_ ;
  assign \new_[25259]_  = A266 & ~A265;
  assign \new_[25260]_  = A236 & \new_[25259]_ ;
  assign \new_[25264]_  = A269 & ~A268;
  assign \new_[25265]_  = ~A267 & \new_[25264]_ ;
  assign \new_[25266]_  = \new_[25265]_  & \new_[25260]_ ;
  assign \new_[25270]_  = A232 & A166;
  assign \new_[25271]_  = A167 & \new_[25270]_ ;
  assign \new_[25275]_  = ~A235 & ~A234;
  assign \new_[25276]_  = ~A233 & \new_[25275]_ ;
  assign \new_[25277]_  = \new_[25276]_  & \new_[25271]_ ;
  assign \new_[25281]_  = ~A266 & A265;
  assign \new_[25282]_  = A236 & \new_[25281]_ ;
  assign \new_[25286]_  = A269 & ~A268;
  assign \new_[25287]_  = ~A267 & \new_[25286]_ ;
  assign \new_[25288]_  = \new_[25287]_  & \new_[25282]_ ;
  assign \new_[25292]_  = ~A199 & A166;
  assign \new_[25293]_  = A167 & \new_[25292]_ ;
  assign \new_[25297]_  = A202 & A201;
  assign \new_[25298]_  = A200 & \new_[25297]_ ;
  assign \new_[25299]_  = \new_[25298]_  & \new_[25293]_ ;
  assign \new_[25303]_  = A269 & ~A268;
  assign \new_[25304]_  = A267 & \new_[25303]_ ;
  assign \new_[25308]_  = A302 & ~A301;
  assign \new_[25309]_  = A300 & \new_[25308]_ ;
  assign \new_[25310]_  = \new_[25309]_  & \new_[25304]_ ;
  assign \new_[25314]_  = ~A199 & A166;
  assign \new_[25315]_  = A167 & \new_[25314]_ ;
  assign \new_[25319]_  = ~A203 & A201;
  assign \new_[25320]_  = A200 & \new_[25319]_ ;
  assign \new_[25321]_  = \new_[25320]_  & \new_[25315]_ ;
  assign \new_[25325]_  = A269 & ~A268;
  assign \new_[25326]_  = A267 & \new_[25325]_ ;
  assign \new_[25330]_  = A302 & ~A301;
  assign \new_[25331]_  = A300 & \new_[25330]_ ;
  assign \new_[25332]_  = \new_[25331]_  & \new_[25326]_ ;
  assign \new_[25336]_  = ~A199 & A166;
  assign \new_[25337]_  = A167 & \new_[25336]_ ;
  assign \new_[25341]_  = ~A202 & ~A201;
  assign \new_[25342]_  = A200 & \new_[25341]_ ;
  assign \new_[25343]_  = \new_[25342]_  & \new_[25337]_ ;
  assign \new_[25347]_  = ~A268 & A267;
  assign \new_[25348]_  = A203 & \new_[25347]_ ;
  assign \new_[25352]_  = A301 & ~A300;
  assign \new_[25353]_  = A269 & \new_[25352]_ ;
  assign \new_[25354]_  = \new_[25353]_  & \new_[25348]_ ;
  assign \new_[25358]_  = ~A199 & A166;
  assign \new_[25359]_  = A167 & \new_[25358]_ ;
  assign \new_[25363]_  = ~A202 & ~A201;
  assign \new_[25364]_  = A200 & \new_[25363]_ ;
  assign \new_[25365]_  = \new_[25364]_  & \new_[25359]_ ;
  assign \new_[25369]_  = ~A268 & A267;
  assign \new_[25370]_  = A203 & \new_[25369]_ ;
  assign \new_[25374]_  = ~A302 & ~A300;
  assign \new_[25375]_  = A269 & \new_[25374]_ ;
  assign \new_[25376]_  = \new_[25375]_  & \new_[25370]_ ;
  assign \new_[25380]_  = ~A199 & A166;
  assign \new_[25381]_  = A167 & \new_[25380]_ ;
  assign \new_[25385]_  = ~A202 & ~A201;
  assign \new_[25386]_  = A200 & \new_[25385]_ ;
  assign \new_[25387]_  = \new_[25386]_  & \new_[25381]_ ;
  assign \new_[25391]_  = ~A268 & A267;
  assign \new_[25392]_  = A203 & \new_[25391]_ ;
  assign \new_[25396]_  = A299 & A298;
  assign \new_[25397]_  = A269 & \new_[25396]_ ;
  assign \new_[25398]_  = \new_[25397]_  & \new_[25392]_ ;
  assign \new_[25402]_  = ~A199 & A166;
  assign \new_[25403]_  = A167 & \new_[25402]_ ;
  assign \new_[25407]_  = ~A202 & ~A201;
  assign \new_[25408]_  = A200 & \new_[25407]_ ;
  assign \new_[25409]_  = \new_[25408]_  & \new_[25403]_ ;
  assign \new_[25413]_  = ~A268 & A267;
  assign \new_[25414]_  = A203 & \new_[25413]_ ;
  assign \new_[25418]_  = ~A299 & ~A298;
  assign \new_[25419]_  = A269 & \new_[25418]_ ;
  assign \new_[25420]_  = \new_[25419]_  & \new_[25414]_ ;
  assign \new_[25424]_  = ~A199 & A166;
  assign \new_[25425]_  = A167 & \new_[25424]_ ;
  assign \new_[25429]_  = ~A202 & ~A201;
  assign \new_[25430]_  = A200 & \new_[25429]_ ;
  assign \new_[25431]_  = \new_[25430]_  & \new_[25425]_ ;
  assign \new_[25435]_  = A268 & ~A267;
  assign \new_[25436]_  = A203 & \new_[25435]_ ;
  assign \new_[25440]_  = A302 & ~A301;
  assign \new_[25441]_  = A300 & \new_[25440]_ ;
  assign \new_[25442]_  = \new_[25441]_  & \new_[25436]_ ;
  assign \new_[25446]_  = ~A199 & A166;
  assign \new_[25447]_  = A167 & \new_[25446]_ ;
  assign \new_[25451]_  = ~A202 & ~A201;
  assign \new_[25452]_  = A200 & \new_[25451]_ ;
  assign \new_[25453]_  = \new_[25452]_  & \new_[25447]_ ;
  assign \new_[25457]_  = ~A269 & ~A267;
  assign \new_[25458]_  = A203 & \new_[25457]_ ;
  assign \new_[25462]_  = A302 & ~A301;
  assign \new_[25463]_  = A300 & \new_[25462]_ ;
  assign \new_[25464]_  = \new_[25463]_  & \new_[25458]_ ;
  assign \new_[25468]_  = ~A199 & A166;
  assign \new_[25469]_  = A167 & \new_[25468]_ ;
  assign \new_[25473]_  = ~A202 & ~A201;
  assign \new_[25474]_  = A200 & \new_[25473]_ ;
  assign \new_[25475]_  = \new_[25474]_  & \new_[25469]_ ;
  assign \new_[25479]_  = A266 & A265;
  assign \new_[25480]_  = A203 & \new_[25479]_ ;
  assign \new_[25484]_  = A302 & ~A301;
  assign \new_[25485]_  = A300 & \new_[25484]_ ;
  assign \new_[25486]_  = \new_[25485]_  & \new_[25480]_ ;
  assign \new_[25490]_  = ~A199 & A166;
  assign \new_[25491]_  = A167 & \new_[25490]_ ;
  assign \new_[25495]_  = ~A202 & ~A201;
  assign \new_[25496]_  = A200 & \new_[25495]_ ;
  assign \new_[25497]_  = \new_[25496]_  & \new_[25491]_ ;
  assign \new_[25501]_  = ~A266 & ~A265;
  assign \new_[25502]_  = A203 & \new_[25501]_ ;
  assign \new_[25506]_  = A302 & ~A301;
  assign \new_[25507]_  = A300 & \new_[25506]_ ;
  assign \new_[25508]_  = \new_[25507]_  & \new_[25502]_ ;
  assign \new_[25512]_  = A199 & A166;
  assign \new_[25513]_  = A167 & \new_[25512]_ ;
  assign \new_[25517]_  = A202 & A201;
  assign \new_[25518]_  = ~A200 & \new_[25517]_ ;
  assign \new_[25519]_  = \new_[25518]_  & \new_[25513]_ ;
  assign \new_[25523]_  = A269 & ~A268;
  assign \new_[25524]_  = A267 & \new_[25523]_ ;
  assign \new_[25528]_  = A302 & ~A301;
  assign \new_[25529]_  = A300 & \new_[25528]_ ;
  assign \new_[25530]_  = \new_[25529]_  & \new_[25524]_ ;
  assign \new_[25534]_  = A199 & A166;
  assign \new_[25535]_  = A167 & \new_[25534]_ ;
  assign \new_[25539]_  = ~A203 & A201;
  assign \new_[25540]_  = ~A200 & \new_[25539]_ ;
  assign \new_[25541]_  = \new_[25540]_  & \new_[25535]_ ;
  assign \new_[25545]_  = A269 & ~A268;
  assign \new_[25546]_  = A267 & \new_[25545]_ ;
  assign \new_[25550]_  = A302 & ~A301;
  assign \new_[25551]_  = A300 & \new_[25550]_ ;
  assign \new_[25552]_  = \new_[25551]_  & \new_[25546]_ ;
  assign \new_[25556]_  = A199 & A166;
  assign \new_[25557]_  = A167 & \new_[25556]_ ;
  assign \new_[25561]_  = ~A202 & ~A201;
  assign \new_[25562]_  = ~A200 & \new_[25561]_ ;
  assign \new_[25563]_  = \new_[25562]_  & \new_[25557]_ ;
  assign \new_[25567]_  = ~A268 & A267;
  assign \new_[25568]_  = A203 & \new_[25567]_ ;
  assign \new_[25572]_  = A301 & ~A300;
  assign \new_[25573]_  = A269 & \new_[25572]_ ;
  assign \new_[25574]_  = \new_[25573]_  & \new_[25568]_ ;
  assign \new_[25578]_  = A199 & A166;
  assign \new_[25579]_  = A167 & \new_[25578]_ ;
  assign \new_[25583]_  = ~A202 & ~A201;
  assign \new_[25584]_  = ~A200 & \new_[25583]_ ;
  assign \new_[25585]_  = \new_[25584]_  & \new_[25579]_ ;
  assign \new_[25589]_  = ~A268 & A267;
  assign \new_[25590]_  = A203 & \new_[25589]_ ;
  assign \new_[25594]_  = ~A302 & ~A300;
  assign \new_[25595]_  = A269 & \new_[25594]_ ;
  assign \new_[25596]_  = \new_[25595]_  & \new_[25590]_ ;
  assign \new_[25600]_  = A199 & A166;
  assign \new_[25601]_  = A167 & \new_[25600]_ ;
  assign \new_[25605]_  = ~A202 & ~A201;
  assign \new_[25606]_  = ~A200 & \new_[25605]_ ;
  assign \new_[25607]_  = \new_[25606]_  & \new_[25601]_ ;
  assign \new_[25611]_  = ~A268 & A267;
  assign \new_[25612]_  = A203 & \new_[25611]_ ;
  assign \new_[25616]_  = A299 & A298;
  assign \new_[25617]_  = A269 & \new_[25616]_ ;
  assign \new_[25618]_  = \new_[25617]_  & \new_[25612]_ ;
  assign \new_[25622]_  = A199 & A166;
  assign \new_[25623]_  = A167 & \new_[25622]_ ;
  assign \new_[25627]_  = ~A202 & ~A201;
  assign \new_[25628]_  = ~A200 & \new_[25627]_ ;
  assign \new_[25629]_  = \new_[25628]_  & \new_[25623]_ ;
  assign \new_[25633]_  = ~A268 & A267;
  assign \new_[25634]_  = A203 & \new_[25633]_ ;
  assign \new_[25638]_  = ~A299 & ~A298;
  assign \new_[25639]_  = A269 & \new_[25638]_ ;
  assign \new_[25640]_  = \new_[25639]_  & \new_[25634]_ ;
  assign \new_[25644]_  = A199 & A166;
  assign \new_[25645]_  = A167 & \new_[25644]_ ;
  assign \new_[25649]_  = ~A202 & ~A201;
  assign \new_[25650]_  = ~A200 & \new_[25649]_ ;
  assign \new_[25651]_  = \new_[25650]_  & \new_[25645]_ ;
  assign \new_[25655]_  = A268 & ~A267;
  assign \new_[25656]_  = A203 & \new_[25655]_ ;
  assign \new_[25660]_  = A302 & ~A301;
  assign \new_[25661]_  = A300 & \new_[25660]_ ;
  assign \new_[25662]_  = \new_[25661]_  & \new_[25656]_ ;
  assign \new_[25666]_  = A199 & A166;
  assign \new_[25667]_  = A167 & \new_[25666]_ ;
  assign \new_[25671]_  = ~A202 & ~A201;
  assign \new_[25672]_  = ~A200 & \new_[25671]_ ;
  assign \new_[25673]_  = \new_[25672]_  & \new_[25667]_ ;
  assign \new_[25677]_  = ~A269 & ~A267;
  assign \new_[25678]_  = A203 & \new_[25677]_ ;
  assign \new_[25682]_  = A302 & ~A301;
  assign \new_[25683]_  = A300 & \new_[25682]_ ;
  assign \new_[25684]_  = \new_[25683]_  & \new_[25678]_ ;
  assign \new_[25688]_  = A199 & A166;
  assign \new_[25689]_  = A167 & \new_[25688]_ ;
  assign \new_[25693]_  = ~A202 & ~A201;
  assign \new_[25694]_  = ~A200 & \new_[25693]_ ;
  assign \new_[25695]_  = \new_[25694]_  & \new_[25689]_ ;
  assign \new_[25699]_  = A266 & A265;
  assign \new_[25700]_  = A203 & \new_[25699]_ ;
  assign \new_[25704]_  = A302 & ~A301;
  assign \new_[25705]_  = A300 & \new_[25704]_ ;
  assign \new_[25706]_  = \new_[25705]_  & \new_[25700]_ ;
  assign \new_[25710]_  = A199 & A166;
  assign \new_[25711]_  = A167 & \new_[25710]_ ;
  assign \new_[25715]_  = ~A202 & ~A201;
  assign \new_[25716]_  = ~A200 & \new_[25715]_ ;
  assign \new_[25717]_  = \new_[25716]_  & \new_[25711]_ ;
  assign \new_[25721]_  = ~A266 & ~A265;
  assign \new_[25722]_  = A203 & \new_[25721]_ ;
  assign \new_[25726]_  = A302 & ~A301;
  assign \new_[25727]_  = A300 & \new_[25726]_ ;
  assign \new_[25728]_  = \new_[25727]_  & \new_[25722]_ ;
  assign \new_[25732]_  = ~A232 & ~A166;
  assign \new_[25733]_  = ~A167 & \new_[25732]_ ;
  assign \new_[25737]_  = ~A235 & ~A234;
  assign \new_[25738]_  = A233 & \new_[25737]_ ;
  assign \new_[25739]_  = \new_[25738]_  & \new_[25733]_ ;
  assign \new_[25743]_  = A266 & ~A265;
  assign \new_[25744]_  = A236 & \new_[25743]_ ;
  assign \new_[25748]_  = A269 & ~A268;
  assign \new_[25749]_  = ~A267 & \new_[25748]_ ;
  assign \new_[25750]_  = \new_[25749]_  & \new_[25744]_ ;
  assign \new_[25754]_  = ~A232 & ~A166;
  assign \new_[25755]_  = ~A167 & \new_[25754]_ ;
  assign \new_[25759]_  = ~A235 & ~A234;
  assign \new_[25760]_  = A233 & \new_[25759]_ ;
  assign \new_[25761]_  = \new_[25760]_  & \new_[25755]_ ;
  assign \new_[25765]_  = ~A266 & A265;
  assign \new_[25766]_  = A236 & \new_[25765]_ ;
  assign \new_[25770]_  = A269 & ~A268;
  assign \new_[25771]_  = ~A267 & \new_[25770]_ ;
  assign \new_[25772]_  = \new_[25771]_  & \new_[25766]_ ;
  assign \new_[25776]_  = A232 & ~A166;
  assign \new_[25777]_  = ~A167 & \new_[25776]_ ;
  assign \new_[25781]_  = ~A235 & ~A234;
  assign \new_[25782]_  = ~A233 & \new_[25781]_ ;
  assign \new_[25783]_  = \new_[25782]_  & \new_[25777]_ ;
  assign \new_[25787]_  = A266 & ~A265;
  assign \new_[25788]_  = A236 & \new_[25787]_ ;
  assign \new_[25792]_  = A269 & ~A268;
  assign \new_[25793]_  = ~A267 & \new_[25792]_ ;
  assign \new_[25794]_  = \new_[25793]_  & \new_[25788]_ ;
  assign \new_[25798]_  = A232 & ~A166;
  assign \new_[25799]_  = ~A167 & \new_[25798]_ ;
  assign \new_[25803]_  = ~A235 & ~A234;
  assign \new_[25804]_  = ~A233 & \new_[25803]_ ;
  assign \new_[25805]_  = \new_[25804]_  & \new_[25799]_ ;
  assign \new_[25809]_  = ~A266 & A265;
  assign \new_[25810]_  = A236 & \new_[25809]_ ;
  assign \new_[25814]_  = A269 & ~A268;
  assign \new_[25815]_  = ~A267 & \new_[25814]_ ;
  assign \new_[25816]_  = \new_[25815]_  & \new_[25810]_ ;
  assign \new_[25820]_  = ~A199 & ~A166;
  assign \new_[25821]_  = ~A167 & \new_[25820]_ ;
  assign \new_[25825]_  = A202 & A201;
  assign \new_[25826]_  = A200 & \new_[25825]_ ;
  assign \new_[25827]_  = \new_[25826]_  & \new_[25821]_ ;
  assign \new_[25831]_  = A269 & ~A268;
  assign \new_[25832]_  = A267 & \new_[25831]_ ;
  assign \new_[25836]_  = A302 & ~A301;
  assign \new_[25837]_  = A300 & \new_[25836]_ ;
  assign \new_[25838]_  = \new_[25837]_  & \new_[25832]_ ;
  assign \new_[25842]_  = ~A199 & ~A166;
  assign \new_[25843]_  = ~A167 & \new_[25842]_ ;
  assign \new_[25847]_  = ~A203 & A201;
  assign \new_[25848]_  = A200 & \new_[25847]_ ;
  assign \new_[25849]_  = \new_[25848]_  & \new_[25843]_ ;
  assign \new_[25853]_  = A269 & ~A268;
  assign \new_[25854]_  = A267 & \new_[25853]_ ;
  assign \new_[25858]_  = A302 & ~A301;
  assign \new_[25859]_  = A300 & \new_[25858]_ ;
  assign \new_[25860]_  = \new_[25859]_  & \new_[25854]_ ;
  assign \new_[25864]_  = ~A199 & ~A166;
  assign \new_[25865]_  = ~A167 & \new_[25864]_ ;
  assign \new_[25869]_  = ~A202 & ~A201;
  assign \new_[25870]_  = A200 & \new_[25869]_ ;
  assign \new_[25871]_  = \new_[25870]_  & \new_[25865]_ ;
  assign \new_[25875]_  = ~A268 & A267;
  assign \new_[25876]_  = A203 & \new_[25875]_ ;
  assign \new_[25880]_  = A301 & ~A300;
  assign \new_[25881]_  = A269 & \new_[25880]_ ;
  assign \new_[25882]_  = \new_[25881]_  & \new_[25876]_ ;
  assign \new_[25886]_  = ~A199 & ~A166;
  assign \new_[25887]_  = ~A167 & \new_[25886]_ ;
  assign \new_[25891]_  = ~A202 & ~A201;
  assign \new_[25892]_  = A200 & \new_[25891]_ ;
  assign \new_[25893]_  = \new_[25892]_  & \new_[25887]_ ;
  assign \new_[25897]_  = ~A268 & A267;
  assign \new_[25898]_  = A203 & \new_[25897]_ ;
  assign \new_[25902]_  = ~A302 & ~A300;
  assign \new_[25903]_  = A269 & \new_[25902]_ ;
  assign \new_[25904]_  = \new_[25903]_  & \new_[25898]_ ;
  assign \new_[25908]_  = ~A199 & ~A166;
  assign \new_[25909]_  = ~A167 & \new_[25908]_ ;
  assign \new_[25913]_  = ~A202 & ~A201;
  assign \new_[25914]_  = A200 & \new_[25913]_ ;
  assign \new_[25915]_  = \new_[25914]_  & \new_[25909]_ ;
  assign \new_[25919]_  = ~A268 & A267;
  assign \new_[25920]_  = A203 & \new_[25919]_ ;
  assign \new_[25924]_  = A299 & A298;
  assign \new_[25925]_  = A269 & \new_[25924]_ ;
  assign \new_[25926]_  = \new_[25925]_  & \new_[25920]_ ;
  assign \new_[25930]_  = ~A199 & ~A166;
  assign \new_[25931]_  = ~A167 & \new_[25930]_ ;
  assign \new_[25935]_  = ~A202 & ~A201;
  assign \new_[25936]_  = A200 & \new_[25935]_ ;
  assign \new_[25937]_  = \new_[25936]_  & \new_[25931]_ ;
  assign \new_[25941]_  = ~A268 & A267;
  assign \new_[25942]_  = A203 & \new_[25941]_ ;
  assign \new_[25946]_  = ~A299 & ~A298;
  assign \new_[25947]_  = A269 & \new_[25946]_ ;
  assign \new_[25948]_  = \new_[25947]_  & \new_[25942]_ ;
  assign \new_[25952]_  = ~A199 & ~A166;
  assign \new_[25953]_  = ~A167 & \new_[25952]_ ;
  assign \new_[25957]_  = ~A202 & ~A201;
  assign \new_[25958]_  = A200 & \new_[25957]_ ;
  assign \new_[25959]_  = \new_[25958]_  & \new_[25953]_ ;
  assign \new_[25963]_  = A268 & ~A267;
  assign \new_[25964]_  = A203 & \new_[25963]_ ;
  assign \new_[25968]_  = A302 & ~A301;
  assign \new_[25969]_  = A300 & \new_[25968]_ ;
  assign \new_[25970]_  = \new_[25969]_  & \new_[25964]_ ;
  assign \new_[25974]_  = ~A199 & ~A166;
  assign \new_[25975]_  = ~A167 & \new_[25974]_ ;
  assign \new_[25979]_  = ~A202 & ~A201;
  assign \new_[25980]_  = A200 & \new_[25979]_ ;
  assign \new_[25981]_  = \new_[25980]_  & \new_[25975]_ ;
  assign \new_[25985]_  = ~A269 & ~A267;
  assign \new_[25986]_  = A203 & \new_[25985]_ ;
  assign \new_[25990]_  = A302 & ~A301;
  assign \new_[25991]_  = A300 & \new_[25990]_ ;
  assign \new_[25992]_  = \new_[25991]_  & \new_[25986]_ ;
  assign \new_[25996]_  = ~A199 & ~A166;
  assign \new_[25997]_  = ~A167 & \new_[25996]_ ;
  assign \new_[26001]_  = ~A202 & ~A201;
  assign \new_[26002]_  = A200 & \new_[26001]_ ;
  assign \new_[26003]_  = \new_[26002]_  & \new_[25997]_ ;
  assign \new_[26007]_  = A266 & A265;
  assign \new_[26008]_  = A203 & \new_[26007]_ ;
  assign \new_[26012]_  = A302 & ~A301;
  assign \new_[26013]_  = A300 & \new_[26012]_ ;
  assign \new_[26014]_  = \new_[26013]_  & \new_[26008]_ ;
  assign \new_[26018]_  = ~A199 & ~A166;
  assign \new_[26019]_  = ~A167 & \new_[26018]_ ;
  assign \new_[26023]_  = ~A202 & ~A201;
  assign \new_[26024]_  = A200 & \new_[26023]_ ;
  assign \new_[26025]_  = \new_[26024]_  & \new_[26019]_ ;
  assign \new_[26029]_  = ~A266 & ~A265;
  assign \new_[26030]_  = A203 & \new_[26029]_ ;
  assign \new_[26034]_  = A302 & ~A301;
  assign \new_[26035]_  = A300 & \new_[26034]_ ;
  assign \new_[26036]_  = \new_[26035]_  & \new_[26030]_ ;
  assign \new_[26040]_  = A199 & ~A166;
  assign \new_[26041]_  = ~A167 & \new_[26040]_ ;
  assign \new_[26045]_  = A202 & A201;
  assign \new_[26046]_  = ~A200 & \new_[26045]_ ;
  assign \new_[26047]_  = \new_[26046]_  & \new_[26041]_ ;
  assign \new_[26051]_  = A269 & ~A268;
  assign \new_[26052]_  = A267 & \new_[26051]_ ;
  assign \new_[26056]_  = A302 & ~A301;
  assign \new_[26057]_  = A300 & \new_[26056]_ ;
  assign \new_[26058]_  = \new_[26057]_  & \new_[26052]_ ;
  assign \new_[26062]_  = A199 & ~A166;
  assign \new_[26063]_  = ~A167 & \new_[26062]_ ;
  assign \new_[26067]_  = ~A203 & A201;
  assign \new_[26068]_  = ~A200 & \new_[26067]_ ;
  assign \new_[26069]_  = \new_[26068]_  & \new_[26063]_ ;
  assign \new_[26073]_  = A269 & ~A268;
  assign \new_[26074]_  = A267 & \new_[26073]_ ;
  assign \new_[26078]_  = A302 & ~A301;
  assign \new_[26079]_  = A300 & \new_[26078]_ ;
  assign \new_[26080]_  = \new_[26079]_  & \new_[26074]_ ;
  assign \new_[26084]_  = A199 & ~A166;
  assign \new_[26085]_  = ~A167 & \new_[26084]_ ;
  assign \new_[26089]_  = ~A202 & ~A201;
  assign \new_[26090]_  = ~A200 & \new_[26089]_ ;
  assign \new_[26091]_  = \new_[26090]_  & \new_[26085]_ ;
  assign \new_[26095]_  = ~A268 & A267;
  assign \new_[26096]_  = A203 & \new_[26095]_ ;
  assign \new_[26100]_  = A301 & ~A300;
  assign \new_[26101]_  = A269 & \new_[26100]_ ;
  assign \new_[26102]_  = \new_[26101]_  & \new_[26096]_ ;
  assign \new_[26106]_  = A199 & ~A166;
  assign \new_[26107]_  = ~A167 & \new_[26106]_ ;
  assign \new_[26111]_  = ~A202 & ~A201;
  assign \new_[26112]_  = ~A200 & \new_[26111]_ ;
  assign \new_[26113]_  = \new_[26112]_  & \new_[26107]_ ;
  assign \new_[26117]_  = ~A268 & A267;
  assign \new_[26118]_  = A203 & \new_[26117]_ ;
  assign \new_[26122]_  = ~A302 & ~A300;
  assign \new_[26123]_  = A269 & \new_[26122]_ ;
  assign \new_[26124]_  = \new_[26123]_  & \new_[26118]_ ;
  assign \new_[26128]_  = A199 & ~A166;
  assign \new_[26129]_  = ~A167 & \new_[26128]_ ;
  assign \new_[26133]_  = ~A202 & ~A201;
  assign \new_[26134]_  = ~A200 & \new_[26133]_ ;
  assign \new_[26135]_  = \new_[26134]_  & \new_[26129]_ ;
  assign \new_[26139]_  = ~A268 & A267;
  assign \new_[26140]_  = A203 & \new_[26139]_ ;
  assign \new_[26144]_  = A299 & A298;
  assign \new_[26145]_  = A269 & \new_[26144]_ ;
  assign \new_[26146]_  = \new_[26145]_  & \new_[26140]_ ;
  assign \new_[26150]_  = A199 & ~A166;
  assign \new_[26151]_  = ~A167 & \new_[26150]_ ;
  assign \new_[26155]_  = ~A202 & ~A201;
  assign \new_[26156]_  = ~A200 & \new_[26155]_ ;
  assign \new_[26157]_  = \new_[26156]_  & \new_[26151]_ ;
  assign \new_[26161]_  = ~A268 & A267;
  assign \new_[26162]_  = A203 & \new_[26161]_ ;
  assign \new_[26166]_  = ~A299 & ~A298;
  assign \new_[26167]_  = A269 & \new_[26166]_ ;
  assign \new_[26168]_  = \new_[26167]_  & \new_[26162]_ ;
  assign \new_[26172]_  = A199 & ~A166;
  assign \new_[26173]_  = ~A167 & \new_[26172]_ ;
  assign \new_[26177]_  = ~A202 & ~A201;
  assign \new_[26178]_  = ~A200 & \new_[26177]_ ;
  assign \new_[26179]_  = \new_[26178]_  & \new_[26173]_ ;
  assign \new_[26183]_  = A268 & ~A267;
  assign \new_[26184]_  = A203 & \new_[26183]_ ;
  assign \new_[26188]_  = A302 & ~A301;
  assign \new_[26189]_  = A300 & \new_[26188]_ ;
  assign \new_[26190]_  = \new_[26189]_  & \new_[26184]_ ;
  assign \new_[26194]_  = A199 & ~A166;
  assign \new_[26195]_  = ~A167 & \new_[26194]_ ;
  assign \new_[26199]_  = ~A202 & ~A201;
  assign \new_[26200]_  = ~A200 & \new_[26199]_ ;
  assign \new_[26201]_  = \new_[26200]_  & \new_[26195]_ ;
  assign \new_[26205]_  = ~A269 & ~A267;
  assign \new_[26206]_  = A203 & \new_[26205]_ ;
  assign \new_[26210]_  = A302 & ~A301;
  assign \new_[26211]_  = A300 & \new_[26210]_ ;
  assign \new_[26212]_  = \new_[26211]_  & \new_[26206]_ ;
  assign \new_[26216]_  = A199 & ~A166;
  assign \new_[26217]_  = ~A167 & \new_[26216]_ ;
  assign \new_[26221]_  = ~A202 & ~A201;
  assign \new_[26222]_  = ~A200 & \new_[26221]_ ;
  assign \new_[26223]_  = \new_[26222]_  & \new_[26217]_ ;
  assign \new_[26227]_  = A266 & A265;
  assign \new_[26228]_  = A203 & \new_[26227]_ ;
  assign \new_[26232]_  = A302 & ~A301;
  assign \new_[26233]_  = A300 & \new_[26232]_ ;
  assign \new_[26234]_  = \new_[26233]_  & \new_[26228]_ ;
  assign \new_[26238]_  = A199 & ~A166;
  assign \new_[26239]_  = ~A167 & \new_[26238]_ ;
  assign \new_[26243]_  = ~A202 & ~A201;
  assign \new_[26244]_  = ~A200 & \new_[26243]_ ;
  assign \new_[26245]_  = \new_[26244]_  & \new_[26239]_ ;
  assign \new_[26249]_  = ~A266 & ~A265;
  assign \new_[26250]_  = A203 & \new_[26249]_ ;
  assign \new_[26254]_  = A302 & ~A301;
  assign \new_[26255]_  = A300 & \new_[26254]_ ;
  assign \new_[26256]_  = \new_[26255]_  & \new_[26250]_ ;
  assign \new_[26260]_  = A200 & ~A199;
  assign \new_[26261]_  = A170 & \new_[26260]_ ;
  assign \new_[26265]_  = A234 & A233;
  assign \new_[26266]_  = ~A232 & \new_[26265]_ ;
  assign \new_[26267]_  = \new_[26266]_  & \new_[26261]_ ;
  assign \new_[26271]_  = A266 & ~A265;
  assign \new_[26272]_  = A235 & \new_[26271]_ ;
  assign \new_[26276]_  = A269 & ~A268;
  assign \new_[26277]_  = ~A267 & \new_[26276]_ ;
  assign \new_[26278]_  = \new_[26277]_  & \new_[26272]_ ;
  assign \new_[26282]_  = A200 & ~A199;
  assign \new_[26283]_  = A170 & \new_[26282]_ ;
  assign \new_[26287]_  = A234 & A233;
  assign \new_[26288]_  = ~A232 & \new_[26287]_ ;
  assign \new_[26289]_  = \new_[26288]_  & \new_[26283]_ ;
  assign \new_[26293]_  = ~A266 & A265;
  assign \new_[26294]_  = A235 & \new_[26293]_ ;
  assign \new_[26298]_  = A269 & ~A268;
  assign \new_[26299]_  = ~A267 & \new_[26298]_ ;
  assign \new_[26300]_  = \new_[26299]_  & \new_[26294]_ ;
  assign \new_[26304]_  = A200 & ~A199;
  assign \new_[26305]_  = A170 & \new_[26304]_ ;
  assign \new_[26309]_  = A234 & A233;
  assign \new_[26310]_  = ~A232 & \new_[26309]_ ;
  assign \new_[26311]_  = \new_[26310]_  & \new_[26305]_ ;
  assign \new_[26315]_  = A266 & ~A265;
  assign \new_[26316]_  = ~A236 & \new_[26315]_ ;
  assign \new_[26320]_  = A269 & ~A268;
  assign \new_[26321]_  = ~A267 & \new_[26320]_ ;
  assign \new_[26322]_  = \new_[26321]_  & \new_[26316]_ ;
  assign \new_[26326]_  = A200 & ~A199;
  assign \new_[26327]_  = A170 & \new_[26326]_ ;
  assign \new_[26331]_  = A234 & A233;
  assign \new_[26332]_  = ~A232 & \new_[26331]_ ;
  assign \new_[26333]_  = \new_[26332]_  & \new_[26327]_ ;
  assign \new_[26337]_  = ~A266 & A265;
  assign \new_[26338]_  = ~A236 & \new_[26337]_ ;
  assign \new_[26342]_  = A269 & ~A268;
  assign \new_[26343]_  = ~A267 & \new_[26342]_ ;
  assign \new_[26344]_  = \new_[26343]_  & \new_[26338]_ ;
  assign \new_[26348]_  = A200 & ~A199;
  assign \new_[26349]_  = A170 & \new_[26348]_ ;
  assign \new_[26353]_  = A234 & ~A233;
  assign \new_[26354]_  = A232 & \new_[26353]_ ;
  assign \new_[26355]_  = \new_[26354]_  & \new_[26349]_ ;
  assign \new_[26359]_  = A266 & ~A265;
  assign \new_[26360]_  = A235 & \new_[26359]_ ;
  assign \new_[26364]_  = A269 & ~A268;
  assign \new_[26365]_  = ~A267 & \new_[26364]_ ;
  assign \new_[26366]_  = \new_[26365]_  & \new_[26360]_ ;
  assign \new_[26370]_  = A200 & ~A199;
  assign \new_[26371]_  = A170 & \new_[26370]_ ;
  assign \new_[26375]_  = A234 & ~A233;
  assign \new_[26376]_  = A232 & \new_[26375]_ ;
  assign \new_[26377]_  = \new_[26376]_  & \new_[26371]_ ;
  assign \new_[26381]_  = ~A266 & A265;
  assign \new_[26382]_  = A235 & \new_[26381]_ ;
  assign \new_[26386]_  = A269 & ~A268;
  assign \new_[26387]_  = ~A267 & \new_[26386]_ ;
  assign \new_[26388]_  = \new_[26387]_  & \new_[26382]_ ;
  assign \new_[26392]_  = A200 & ~A199;
  assign \new_[26393]_  = A170 & \new_[26392]_ ;
  assign \new_[26397]_  = A234 & ~A233;
  assign \new_[26398]_  = A232 & \new_[26397]_ ;
  assign \new_[26399]_  = \new_[26398]_  & \new_[26393]_ ;
  assign \new_[26403]_  = A266 & ~A265;
  assign \new_[26404]_  = ~A236 & \new_[26403]_ ;
  assign \new_[26408]_  = A269 & ~A268;
  assign \new_[26409]_  = ~A267 & \new_[26408]_ ;
  assign \new_[26410]_  = \new_[26409]_  & \new_[26404]_ ;
  assign \new_[26414]_  = A200 & ~A199;
  assign \new_[26415]_  = A170 & \new_[26414]_ ;
  assign \new_[26419]_  = A234 & ~A233;
  assign \new_[26420]_  = A232 & \new_[26419]_ ;
  assign \new_[26421]_  = \new_[26420]_  & \new_[26415]_ ;
  assign \new_[26425]_  = ~A266 & A265;
  assign \new_[26426]_  = ~A236 & \new_[26425]_ ;
  assign \new_[26430]_  = A269 & ~A268;
  assign \new_[26431]_  = ~A267 & \new_[26430]_ ;
  assign \new_[26432]_  = \new_[26431]_  & \new_[26426]_ ;
  assign \new_[26436]_  = ~A200 & A199;
  assign \new_[26437]_  = A170 & \new_[26436]_ ;
  assign \new_[26441]_  = A234 & A233;
  assign \new_[26442]_  = ~A232 & \new_[26441]_ ;
  assign \new_[26443]_  = \new_[26442]_  & \new_[26437]_ ;
  assign \new_[26447]_  = A266 & ~A265;
  assign \new_[26448]_  = A235 & \new_[26447]_ ;
  assign \new_[26452]_  = A269 & ~A268;
  assign \new_[26453]_  = ~A267 & \new_[26452]_ ;
  assign \new_[26454]_  = \new_[26453]_  & \new_[26448]_ ;
  assign \new_[26458]_  = ~A200 & A199;
  assign \new_[26459]_  = A170 & \new_[26458]_ ;
  assign \new_[26463]_  = A234 & A233;
  assign \new_[26464]_  = ~A232 & \new_[26463]_ ;
  assign \new_[26465]_  = \new_[26464]_  & \new_[26459]_ ;
  assign \new_[26469]_  = ~A266 & A265;
  assign \new_[26470]_  = A235 & \new_[26469]_ ;
  assign \new_[26474]_  = A269 & ~A268;
  assign \new_[26475]_  = ~A267 & \new_[26474]_ ;
  assign \new_[26476]_  = \new_[26475]_  & \new_[26470]_ ;
  assign \new_[26480]_  = ~A200 & A199;
  assign \new_[26481]_  = A170 & \new_[26480]_ ;
  assign \new_[26485]_  = A234 & A233;
  assign \new_[26486]_  = ~A232 & \new_[26485]_ ;
  assign \new_[26487]_  = \new_[26486]_  & \new_[26481]_ ;
  assign \new_[26491]_  = A266 & ~A265;
  assign \new_[26492]_  = ~A236 & \new_[26491]_ ;
  assign \new_[26496]_  = A269 & ~A268;
  assign \new_[26497]_  = ~A267 & \new_[26496]_ ;
  assign \new_[26498]_  = \new_[26497]_  & \new_[26492]_ ;
  assign \new_[26502]_  = ~A200 & A199;
  assign \new_[26503]_  = A170 & \new_[26502]_ ;
  assign \new_[26507]_  = A234 & A233;
  assign \new_[26508]_  = ~A232 & \new_[26507]_ ;
  assign \new_[26509]_  = \new_[26508]_  & \new_[26503]_ ;
  assign \new_[26513]_  = ~A266 & A265;
  assign \new_[26514]_  = ~A236 & \new_[26513]_ ;
  assign \new_[26518]_  = A269 & ~A268;
  assign \new_[26519]_  = ~A267 & \new_[26518]_ ;
  assign \new_[26520]_  = \new_[26519]_  & \new_[26514]_ ;
  assign \new_[26524]_  = ~A200 & A199;
  assign \new_[26525]_  = A170 & \new_[26524]_ ;
  assign \new_[26529]_  = A234 & ~A233;
  assign \new_[26530]_  = A232 & \new_[26529]_ ;
  assign \new_[26531]_  = \new_[26530]_  & \new_[26525]_ ;
  assign \new_[26535]_  = A266 & ~A265;
  assign \new_[26536]_  = A235 & \new_[26535]_ ;
  assign \new_[26540]_  = A269 & ~A268;
  assign \new_[26541]_  = ~A267 & \new_[26540]_ ;
  assign \new_[26542]_  = \new_[26541]_  & \new_[26536]_ ;
  assign \new_[26546]_  = ~A200 & A199;
  assign \new_[26547]_  = A170 & \new_[26546]_ ;
  assign \new_[26551]_  = A234 & ~A233;
  assign \new_[26552]_  = A232 & \new_[26551]_ ;
  assign \new_[26553]_  = \new_[26552]_  & \new_[26547]_ ;
  assign \new_[26557]_  = ~A266 & A265;
  assign \new_[26558]_  = A235 & \new_[26557]_ ;
  assign \new_[26562]_  = A269 & ~A268;
  assign \new_[26563]_  = ~A267 & \new_[26562]_ ;
  assign \new_[26564]_  = \new_[26563]_  & \new_[26558]_ ;
  assign \new_[26568]_  = ~A200 & A199;
  assign \new_[26569]_  = A170 & \new_[26568]_ ;
  assign \new_[26573]_  = A234 & ~A233;
  assign \new_[26574]_  = A232 & \new_[26573]_ ;
  assign \new_[26575]_  = \new_[26574]_  & \new_[26569]_ ;
  assign \new_[26579]_  = A266 & ~A265;
  assign \new_[26580]_  = ~A236 & \new_[26579]_ ;
  assign \new_[26584]_  = A269 & ~A268;
  assign \new_[26585]_  = ~A267 & \new_[26584]_ ;
  assign \new_[26586]_  = \new_[26585]_  & \new_[26580]_ ;
  assign \new_[26590]_  = ~A200 & A199;
  assign \new_[26591]_  = A170 & \new_[26590]_ ;
  assign \new_[26595]_  = A234 & ~A233;
  assign \new_[26596]_  = A232 & \new_[26595]_ ;
  assign \new_[26597]_  = \new_[26596]_  & \new_[26591]_ ;
  assign \new_[26601]_  = ~A266 & A265;
  assign \new_[26602]_  = ~A236 & \new_[26601]_ ;
  assign \new_[26606]_  = A269 & ~A268;
  assign \new_[26607]_  = ~A267 & \new_[26606]_ ;
  assign \new_[26608]_  = \new_[26607]_  & \new_[26602]_ ;
  assign \new_[26612]_  = A167 & A168;
  assign \new_[26613]_  = A170 & \new_[26612]_ ;
  assign \new_[26617]_  = A202 & ~A201;
  assign \new_[26618]_  = ~A166 & \new_[26617]_ ;
  assign \new_[26619]_  = \new_[26618]_  & \new_[26613]_ ;
  assign \new_[26623]_  = A298 & A268;
  assign \new_[26624]_  = ~A267 & \new_[26623]_ ;
  assign \new_[26628]_  = A301 & A300;
  assign \new_[26629]_  = ~A299 & \new_[26628]_ ;
  assign \new_[26630]_  = \new_[26629]_  & \new_[26624]_ ;
  assign \new_[26634]_  = A167 & A168;
  assign \new_[26635]_  = A170 & \new_[26634]_ ;
  assign \new_[26639]_  = A202 & ~A201;
  assign \new_[26640]_  = ~A166 & \new_[26639]_ ;
  assign \new_[26641]_  = \new_[26640]_  & \new_[26635]_ ;
  assign \new_[26645]_  = A298 & A268;
  assign \new_[26646]_  = ~A267 & \new_[26645]_ ;
  assign \new_[26650]_  = ~A302 & A300;
  assign \new_[26651]_  = ~A299 & \new_[26650]_ ;
  assign \new_[26652]_  = \new_[26651]_  & \new_[26646]_ ;
  assign \new_[26656]_  = A167 & A168;
  assign \new_[26657]_  = A170 & \new_[26656]_ ;
  assign \new_[26661]_  = A202 & ~A201;
  assign \new_[26662]_  = ~A166 & \new_[26661]_ ;
  assign \new_[26663]_  = \new_[26662]_  & \new_[26657]_ ;
  assign \new_[26667]_  = ~A298 & A268;
  assign \new_[26668]_  = ~A267 & \new_[26667]_ ;
  assign \new_[26672]_  = A301 & A300;
  assign \new_[26673]_  = A299 & \new_[26672]_ ;
  assign \new_[26674]_  = \new_[26673]_  & \new_[26668]_ ;
  assign \new_[26678]_  = A167 & A168;
  assign \new_[26679]_  = A170 & \new_[26678]_ ;
  assign \new_[26683]_  = A202 & ~A201;
  assign \new_[26684]_  = ~A166 & \new_[26683]_ ;
  assign \new_[26685]_  = \new_[26684]_  & \new_[26679]_ ;
  assign \new_[26689]_  = ~A298 & A268;
  assign \new_[26690]_  = ~A267 & \new_[26689]_ ;
  assign \new_[26694]_  = ~A302 & A300;
  assign \new_[26695]_  = A299 & \new_[26694]_ ;
  assign \new_[26696]_  = \new_[26695]_  & \new_[26690]_ ;
  assign \new_[26700]_  = A167 & A168;
  assign \new_[26701]_  = A170 & \new_[26700]_ ;
  assign \new_[26705]_  = A202 & ~A201;
  assign \new_[26706]_  = ~A166 & \new_[26705]_ ;
  assign \new_[26707]_  = \new_[26706]_  & \new_[26701]_ ;
  assign \new_[26711]_  = A298 & ~A269;
  assign \new_[26712]_  = ~A267 & \new_[26711]_ ;
  assign \new_[26716]_  = A301 & A300;
  assign \new_[26717]_  = ~A299 & \new_[26716]_ ;
  assign \new_[26718]_  = \new_[26717]_  & \new_[26712]_ ;
  assign \new_[26722]_  = A167 & A168;
  assign \new_[26723]_  = A170 & \new_[26722]_ ;
  assign \new_[26727]_  = A202 & ~A201;
  assign \new_[26728]_  = ~A166 & \new_[26727]_ ;
  assign \new_[26729]_  = \new_[26728]_  & \new_[26723]_ ;
  assign \new_[26733]_  = A298 & ~A269;
  assign \new_[26734]_  = ~A267 & \new_[26733]_ ;
  assign \new_[26738]_  = ~A302 & A300;
  assign \new_[26739]_  = ~A299 & \new_[26738]_ ;
  assign \new_[26740]_  = \new_[26739]_  & \new_[26734]_ ;
  assign \new_[26744]_  = A167 & A168;
  assign \new_[26745]_  = A170 & \new_[26744]_ ;
  assign \new_[26749]_  = A202 & ~A201;
  assign \new_[26750]_  = ~A166 & \new_[26749]_ ;
  assign \new_[26751]_  = \new_[26750]_  & \new_[26745]_ ;
  assign \new_[26755]_  = ~A298 & ~A269;
  assign \new_[26756]_  = ~A267 & \new_[26755]_ ;
  assign \new_[26760]_  = A301 & A300;
  assign \new_[26761]_  = A299 & \new_[26760]_ ;
  assign \new_[26762]_  = \new_[26761]_  & \new_[26756]_ ;
  assign \new_[26766]_  = A167 & A168;
  assign \new_[26767]_  = A170 & \new_[26766]_ ;
  assign \new_[26771]_  = A202 & ~A201;
  assign \new_[26772]_  = ~A166 & \new_[26771]_ ;
  assign \new_[26773]_  = \new_[26772]_  & \new_[26767]_ ;
  assign \new_[26777]_  = ~A298 & ~A269;
  assign \new_[26778]_  = ~A267 & \new_[26777]_ ;
  assign \new_[26782]_  = ~A302 & A300;
  assign \new_[26783]_  = A299 & \new_[26782]_ ;
  assign \new_[26784]_  = \new_[26783]_  & \new_[26778]_ ;
  assign \new_[26788]_  = A167 & A168;
  assign \new_[26789]_  = A170 & \new_[26788]_ ;
  assign \new_[26793]_  = A202 & ~A201;
  assign \new_[26794]_  = ~A166 & \new_[26793]_ ;
  assign \new_[26795]_  = \new_[26794]_  & \new_[26789]_ ;
  assign \new_[26799]_  = A298 & A266;
  assign \new_[26800]_  = A265 & \new_[26799]_ ;
  assign \new_[26804]_  = A301 & A300;
  assign \new_[26805]_  = ~A299 & \new_[26804]_ ;
  assign \new_[26806]_  = \new_[26805]_  & \new_[26800]_ ;
  assign \new_[26810]_  = A167 & A168;
  assign \new_[26811]_  = A170 & \new_[26810]_ ;
  assign \new_[26815]_  = A202 & ~A201;
  assign \new_[26816]_  = ~A166 & \new_[26815]_ ;
  assign \new_[26817]_  = \new_[26816]_  & \new_[26811]_ ;
  assign \new_[26821]_  = A298 & A266;
  assign \new_[26822]_  = A265 & \new_[26821]_ ;
  assign \new_[26826]_  = ~A302 & A300;
  assign \new_[26827]_  = ~A299 & \new_[26826]_ ;
  assign \new_[26828]_  = \new_[26827]_  & \new_[26822]_ ;
  assign \new_[26832]_  = A167 & A168;
  assign \new_[26833]_  = A170 & \new_[26832]_ ;
  assign \new_[26837]_  = A202 & ~A201;
  assign \new_[26838]_  = ~A166 & \new_[26837]_ ;
  assign \new_[26839]_  = \new_[26838]_  & \new_[26833]_ ;
  assign \new_[26843]_  = ~A298 & A266;
  assign \new_[26844]_  = A265 & \new_[26843]_ ;
  assign \new_[26848]_  = A301 & A300;
  assign \new_[26849]_  = A299 & \new_[26848]_ ;
  assign \new_[26850]_  = \new_[26849]_  & \new_[26844]_ ;
  assign \new_[26854]_  = A167 & A168;
  assign \new_[26855]_  = A170 & \new_[26854]_ ;
  assign \new_[26859]_  = A202 & ~A201;
  assign \new_[26860]_  = ~A166 & \new_[26859]_ ;
  assign \new_[26861]_  = \new_[26860]_  & \new_[26855]_ ;
  assign \new_[26865]_  = ~A298 & A266;
  assign \new_[26866]_  = A265 & \new_[26865]_ ;
  assign \new_[26870]_  = ~A302 & A300;
  assign \new_[26871]_  = A299 & \new_[26870]_ ;
  assign \new_[26872]_  = \new_[26871]_  & \new_[26866]_ ;
  assign \new_[26876]_  = A167 & A168;
  assign \new_[26877]_  = A170 & \new_[26876]_ ;
  assign \new_[26881]_  = A202 & ~A201;
  assign \new_[26882]_  = ~A166 & \new_[26881]_ ;
  assign \new_[26883]_  = \new_[26882]_  & \new_[26877]_ ;
  assign \new_[26887]_  = A267 & A266;
  assign \new_[26888]_  = ~A265 & \new_[26887]_ ;
  assign \new_[26892]_  = A301 & ~A300;
  assign \new_[26893]_  = A268 & \new_[26892]_ ;
  assign \new_[26894]_  = \new_[26893]_  & \new_[26888]_ ;
  assign \new_[26898]_  = A167 & A168;
  assign \new_[26899]_  = A170 & \new_[26898]_ ;
  assign \new_[26903]_  = A202 & ~A201;
  assign \new_[26904]_  = ~A166 & \new_[26903]_ ;
  assign \new_[26905]_  = \new_[26904]_  & \new_[26899]_ ;
  assign \new_[26909]_  = A267 & A266;
  assign \new_[26910]_  = ~A265 & \new_[26909]_ ;
  assign \new_[26914]_  = ~A302 & ~A300;
  assign \new_[26915]_  = A268 & \new_[26914]_ ;
  assign \new_[26916]_  = \new_[26915]_  & \new_[26910]_ ;
  assign \new_[26920]_  = A167 & A168;
  assign \new_[26921]_  = A170 & \new_[26920]_ ;
  assign \new_[26925]_  = A202 & ~A201;
  assign \new_[26926]_  = ~A166 & \new_[26925]_ ;
  assign \new_[26927]_  = \new_[26926]_  & \new_[26921]_ ;
  assign \new_[26931]_  = A267 & A266;
  assign \new_[26932]_  = ~A265 & \new_[26931]_ ;
  assign \new_[26936]_  = A299 & A298;
  assign \new_[26937]_  = A268 & \new_[26936]_ ;
  assign \new_[26938]_  = \new_[26937]_  & \new_[26932]_ ;
  assign \new_[26942]_  = A167 & A168;
  assign \new_[26943]_  = A170 & \new_[26942]_ ;
  assign \new_[26947]_  = A202 & ~A201;
  assign \new_[26948]_  = ~A166 & \new_[26947]_ ;
  assign \new_[26949]_  = \new_[26948]_  & \new_[26943]_ ;
  assign \new_[26953]_  = A267 & A266;
  assign \new_[26954]_  = ~A265 & \new_[26953]_ ;
  assign \new_[26958]_  = ~A299 & ~A298;
  assign \new_[26959]_  = A268 & \new_[26958]_ ;
  assign \new_[26960]_  = \new_[26959]_  & \new_[26954]_ ;
  assign \new_[26964]_  = A167 & A168;
  assign \new_[26965]_  = A170 & \new_[26964]_ ;
  assign \new_[26969]_  = A202 & ~A201;
  assign \new_[26970]_  = ~A166 & \new_[26969]_ ;
  assign \new_[26971]_  = \new_[26970]_  & \new_[26965]_ ;
  assign \new_[26975]_  = A267 & A266;
  assign \new_[26976]_  = ~A265 & \new_[26975]_ ;
  assign \new_[26980]_  = A301 & ~A300;
  assign \new_[26981]_  = ~A269 & \new_[26980]_ ;
  assign \new_[26982]_  = \new_[26981]_  & \new_[26976]_ ;
  assign \new_[26986]_  = A167 & A168;
  assign \new_[26987]_  = A170 & \new_[26986]_ ;
  assign \new_[26991]_  = A202 & ~A201;
  assign \new_[26992]_  = ~A166 & \new_[26991]_ ;
  assign \new_[26993]_  = \new_[26992]_  & \new_[26987]_ ;
  assign \new_[26997]_  = A267 & A266;
  assign \new_[26998]_  = ~A265 & \new_[26997]_ ;
  assign \new_[27002]_  = ~A302 & ~A300;
  assign \new_[27003]_  = ~A269 & \new_[27002]_ ;
  assign \new_[27004]_  = \new_[27003]_  & \new_[26998]_ ;
  assign \new_[27008]_  = A167 & A168;
  assign \new_[27009]_  = A170 & \new_[27008]_ ;
  assign \new_[27013]_  = A202 & ~A201;
  assign \new_[27014]_  = ~A166 & \new_[27013]_ ;
  assign \new_[27015]_  = \new_[27014]_  & \new_[27009]_ ;
  assign \new_[27019]_  = A267 & A266;
  assign \new_[27020]_  = ~A265 & \new_[27019]_ ;
  assign \new_[27024]_  = A299 & A298;
  assign \new_[27025]_  = ~A269 & \new_[27024]_ ;
  assign \new_[27026]_  = \new_[27025]_  & \new_[27020]_ ;
  assign \new_[27030]_  = A167 & A168;
  assign \new_[27031]_  = A170 & \new_[27030]_ ;
  assign \new_[27035]_  = A202 & ~A201;
  assign \new_[27036]_  = ~A166 & \new_[27035]_ ;
  assign \new_[27037]_  = \new_[27036]_  & \new_[27031]_ ;
  assign \new_[27041]_  = A267 & A266;
  assign \new_[27042]_  = ~A265 & \new_[27041]_ ;
  assign \new_[27046]_  = ~A299 & ~A298;
  assign \new_[27047]_  = ~A269 & \new_[27046]_ ;
  assign \new_[27048]_  = \new_[27047]_  & \new_[27042]_ ;
  assign \new_[27052]_  = A167 & A168;
  assign \new_[27053]_  = A170 & \new_[27052]_ ;
  assign \new_[27057]_  = A202 & ~A201;
  assign \new_[27058]_  = ~A166 & \new_[27057]_ ;
  assign \new_[27059]_  = \new_[27058]_  & \new_[27053]_ ;
  assign \new_[27063]_  = A267 & ~A266;
  assign \new_[27064]_  = A265 & \new_[27063]_ ;
  assign \new_[27068]_  = A301 & ~A300;
  assign \new_[27069]_  = A268 & \new_[27068]_ ;
  assign \new_[27070]_  = \new_[27069]_  & \new_[27064]_ ;
  assign \new_[27074]_  = A167 & A168;
  assign \new_[27075]_  = A170 & \new_[27074]_ ;
  assign \new_[27079]_  = A202 & ~A201;
  assign \new_[27080]_  = ~A166 & \new_[27079]_ ;
  assign \new_[27081]_  = \new_[27080]_  & \new_[27075]_ ;
  assign \new_[27085]_  = A267 & ~A266;
  assign \new_[27086]_  = A265 & \new_[27085]_ ;
  assign \new_[27090]_  = ~A302 & ~A300;
  assign \new_[27091]_  = A268 & \new_[27090]_ ;
  assign \new_[27092]_  = \new_[27091]_  & \new_[27086]_ ;
  assign \new_[27096]_  = A167 & A168;
  assign \new_[27097]_  = A170 & \new_[27096]_ ;
  assign \new_[27101]_  = A202 & ~A201;
  assign \new_[27102]_  = ~A166 & \new_[27101]_ ;
  assign \new_[27103]_  = \new_[27102]_  & \new_[27097]_ ;
  assign \new_[27107]_  = A267 & ~A266;
  assign \new_[27108]_  = A265 & \new_[27107]_ ;
  assign \new_[27112]_  = A299 & A298;
  assign \new_[27113]_  = A268 & \new_[27112]_ ;
  assign \new_[27114]_  = \new_[27113]_  & \new_[27108]_ ;
  assign \new_[27118]_  = A167 & A168;
  assign \new_[27119]_  = A170 & \new_[27118]_ ;
  assign \new_[27123]_  = A202 & ~A201;
  assign \new_[27124]_  = ~A166 & \new_[27123]_ ;
  assign \new_[27125]_  = \new_[27124]_  & \new_[27119]_ ;
  assign \new_[27129]_  = A267 & ~A266;
  assign \new_[27130]_  = A265 & \new_[27129]_ ;
  assign \new_[27134]_  = ~A299 & ~A298;
  assign \new_[27135]_  = A268 & \new_[27134]_ ;
  assign \new_[27136]_  = \new_[27135]_  & \new_[27130]_ ;
  assign \new_[27140]_  = A167 & A168;
  assign \new_[27141]_  = A170 & \new_[27140]_ ;
  assign \new_[27145]_  = A202 & ~A201;
  assign \new_[27146]_  = ~A166 & \new_[27145]_ ;
  assign \new_[27147]_  = \new_[27146]_  & \new_[27141]_ ;
  assign \new_[27151]_  = A267 & ~A266;
  assign \new_[27152]_  = A265 & \new_[27151]_ ;
  assign \new_[27156]_  = A301 & ~A300;
  assign \new_[27157]_  = ~A269 & \new_[27156]_ ;
  assign \new_[27158]_  = \new_[27157]_  & \new_[27152]_ ;
  assign \new_[27162]_  = A167 & A168;
  assign \new_[27163]_  = A170 & \new_[27162]_ ;
  assign \new_[27167]_  = A202 & ~A201;
  assign \new_[27168]_  = ~A166 & \new_[27167]_ ;
  assign \new_[27169]_  = \new_[27168]_  & \new_[27163]_ ;
  assign \new_[27173]_  = A267 & ~A266;
  assign \new_[27174]_  = A265 & \new_[27173]_ ;
  assign \new_[27178]_  = ~A302 & ~A300;
  assign \new_[27179]_  = ~A269 & \new_[27178]_ ;
  assign \new_[27180]_  = \new_[27179]_  & \new_[27174]_ ;
  assign \new_[27184]_  = A167 & A168;
  assign \new_[27185]_  = A170 & \new_[27184]_ ;
  assign \new_[27189]_  = A202 & ~A201;
  assign \new_[27190]_  = ~A166 & \new_[27189]_ ;
  assign \new_[27191]_  = \new_[27190]_  & \new_[27185]_ ;
  assign \new_[27195]_  = A267 & ~A266;
  assign \new_[27196]_  = A265 & \new_[27195]_ ;
  assign \new_[27200]_  = A299 & A298;
  assign \new_[27201]_  = ~A269 & \new_[27200]_ ;
  assign \new_[27202]_  = \new_[27201]_  & \new_[27196]_ ;
  assign \new_[27206]_  = A167 & A168;
  assign \new_[27207]_  = A170 & \new_[27206]_ ;
  assign \new_[27211]_  = A202 & ~A201;
  assign \new_[27212]_  = ~A166 & \new_[27211]_ ;
  assign \new_[27213]_  = \new_[27212]_  & \new_[27207]_ ;
  assign \new_[27217]_  = A267 & ~A266;
  assign \new_[27218]_  = A265 & \new_[27217]_ ;
  assign \new_[27222]_  = ~A299 & ~A298;
  assign \new_[27223]_  = ~A269 & \new_[27222]_ ;
  assign \new_[27224]_  = \new_[27223]_  & \new_[27218]_ ;
  assign \new_[27228]_  = A167 & A168;
  assign \new_[27229]_  = A170 & \new_[27228]_ ;
  assign \new_[27233]_  = A202 & ~A201;
  assign \new_[27234]_  = ~A166 & \new_[27233]_ ;
  assign \new_[27235]_  = \new_[27234]_  & \new_[27229]_ ;
  assign \new_[27239]_  = A298 & ~A266;
  assign \new_[27240]_  = ~A265 & \new_[27239]_ ;
  assign \new_[27244]_  = A301 & A300;
  assign \new_[27245]_  = ~A299 & \new_[27244]_ ;
  assign \new_[27246]_  = \new_[27245]_  & \new_[27240]_ ;
  assign \new_[27250]_  = A167 & A168;
  assign \new_[27251]_  = A170 & \new_[27250]_ ;
  assign \new_[27255]_  = A202 & ~A201;
  assign \new_[27256]_  = ~A166 & \new_[27255]_ ;
  assign \new_[27257]_  = \new_[27256]_  & \new_[27251]_ ;
  assign \new_[27261]_  = A298 & ~A266;
  assign \new_[27262]_  = ~A265 & \new_[27261]_ ;
  assign \new_[27266]_  = ~A302 & A300;
  assign \new_[27267]_  = ~A299 & \new_[27266]_ ;
  assign \new_[27268]_  = \new_[27267]_  & \new_[27262]_ ;
  assign \new_[27272]_  = A167 & A168;
  assign \new_[27273]_  = A170 & \new_[27272]_ ;
  assign \new_[27277]_  = A202 & ~A201;
  assign \new_[27278]_  = ~A166 & \new_[27277]_ ;
  assign \new_[27279]_  = \new_[27278]_  & \new_[27273]_ ;
  assign \new_[27283]_  = ~A298 & ~A266;
  assign \new_[27284]_  = ~A265 & \new_[27283]_ ;
  assign \new_[27288]_  = A301 & A300;
  assign \new_[27289]_  = A299 & \new_[27288]_ ;
  assign \new_[27290]_  = \new_[27289]_  & \new_[27284]_ ;
  assign \new_[27294]_  = A167 & A168;
  assign \new_[27295]_  = A170 & \new_[27294]_ ;
  assign \new_[27299]_  = A202 & ~A201;
  assign \new_[27300]_  = ~A166 & \new_[27299]_ ;
  assign \new_[27301]_  = \new_[27300]_  & \new_[27295]_ ;
  assign \new_[27305]_  = ~A298 & ~A266;
  assign \new_[27306]_  = ~A265 & \new_[27305]_ ;
  assign \new_[27310]_  = ~A302 & A300;
  assign \new_[27311]_  = A299 & \new_[27310]_ ;
  assign \new_[27312]_  = \new_[27311]_  & \new_[27306]_ ;
  assign \new_[27316]_  = A167 & A168;
  assign \new_[27317]_  = A170 & \new_[27316]_ ;
  assign \new_[27321]_  = ~A203 & ~A201;
  assign \new_[27322]_  = ~A166 & \new_[27321]_ ;
  assign \new_[27323]_  = \new_[27322]_  & \new_[27317]_ ;
  assign \new_[27327]_  = A298 & A268;
  assign \new_[27328]_  = ~A267 & \new_[27327]_ ;
  assign \new_[27332]_  = A301 & A300;
  assign \new_[27333]_  = ~A299 & \new_[27332]_ ;
  assign \new_[27334]_  = \new_[27333]_  & \new_[27328]_ ;
  assign \new_[27338]_  = A167 & A168;
  assign \new_[27339]_  = A170 & \new_[27338]_ ;
  assign \new_[27343]_  = ~A203 & ~A201;
  assign \new_[27344]_  = ~A166 & \new_[27343]_ ;
  assign \new_[27345]_  = \new_[27344]_  & \new_[27339]_ ;
  assign \new_[27349]_  = A298 & A268;
  assign \new_[27350]_  = ~A267 & \new_[27349]_ ;
  assign \new_[27354]_  = ~A302 & A300;
  assign \new_[27355]_  = ~A299 & \new_[27354]_ ;
  assign \new_[27356]_  = \new_[27355]_  & \new_[27350]_ ;
  assign \new_[27360]_  = A167 & A168;
  assign \new_[27361]_  = A170 & \new_[27360]_ ;
  assign \new_[27365]_  = ~A203 & ~A201;
  assign \new_[27366]_  = ~A166 & \new_[27365]_ ;
  assign \new_[27367]_  = \new_[27366]_  & \new_[27361]_ ;
  assign \new_[27371]_  = ~A298 & A268;
  assign \new_[27372]_  = ~A267 & \new_[27371]_ ;
  assign \new_[27376]_  = A301 & A300;
  assign \new_[27377]_  = A299 & \new_[27376]_ ;
  assign \new_[27378]_  = \new_[27377]_  & \new_[27372]_ ;
  assign \new_[27382]_  = A167 & A168;
  assign \new_[27383]_  = A170 & \new_[27382]_ ;
  assign \new_[27387]_  = ~A203 & ~A201;
  assign \new_[27388]_  = ~A166 & \new_[27387]_ ;
  assign \new_[27389]_  = \new_[27388]_  & \new_[27383]_ ;
  assign \new_[27393]_  = ~A298 & A268;
  assign \new_[27394]_  = ~A267 & \new_[27393]_ ;
  assign \new_[27398]_  = ~A302 & A300;
  assign \new_[27399]_  = A299 & \new_[27398]_ ;
  assign \new_[27400]_  = \new_[27399]_  & \new_[27394]_ ;
  assign \new_[27404]_  = A167 & A168;
  assign \new_[27405]_  = A170 & \new_[27404]_ ;
  assign \new_[27409]_  = ~A203 & ~A201;
  assign \new_[27410]_  = ~A166 & \new_[27409]_ ;
  assign \new_[27411]_  = \new_[27410]_  & \new_[27405]_ ;
  assign \new_[27415]_  = A298 & ~A269;
  assign \new_[27416]_  = ~A267 & \new_[27415]_ ;
  assign \new_[27420]_  = A301 & A300;
  assign \new_[27421]_  = ~A299 & \new_[27420]_ ;
  assign \new_[27422]_  = \new_[27421]_  & \new_[27416]_ ;
  assign \new_[27426]_  = A167 & A168;
  assign \new_[27427]_  = A170 & \new_[27426]_ ;
  assign \new_[27431]_  = ~A203 & ~A201;
  assign \new_[27432]_  = ~A166 & \new_[27431]_ ;
  assign \new_[27433]_  = \new_[27432]_  & \new_[27427]_ ;
  assign \new_[27437]_  = A298 & ~A269;
  assign \new_[27438]_  = ~A267 & \new_[27437]_ ;
  assign \new_[27442]_  = ~A302 & A300;
  assign \new_[27443]_  = ~A299 & \new_[27442]_ ;
  assign \new_[27444]_  = \new_[27443]_  & \new_[27438]_ ;
  assign \new_[27448]_  = A167 & A168;
  assign \new_[27449]_  = A170 & \new_[27448]_ ;
  assign \new_[27453]_  = ~A203 & ~A201;
  assign \new_[27454]_  = ~A166 & \new_[27453]_ ;
  assign \new_[27455]_  = \new_[27454]_  & \new_[27449]_ ;
  assign \new_[27459]_  = ~A298 & ~A269;
  assign \new_[27460]_  = ~A267 & \new_[27459]_ ;
  assign \new_[27464]_  = A301 & A300;
  assign \new_[27465]_  = A299 & \new_[27464]_ ;
  assign \new_[27466]_  = \new_[27465]_  & \new_[27460]_ ;
  assign \new_[27470]_  = A167 & A168;
  assign \new_[27471]_  = A170 & \new_[27470]_ ;
  assign \new_[27475]_  = ~A203 & ~A201;
  assign \new_[27476]_  = ~A166 & \new_[27475]_ ;
  assign \new_[27477]_  = \new_[27476]_  & \new_[27471]_ ;
  assign \new_[27481]_  = ~A298 & ~A269;
  assign \new_[27482]_  = ~A267 & \new_[27481]_ ;
  assign \new_[27486]_  = ~A302 & A300;
  assign \new_[27487]_  = A299 & \new_[27486]_ ;
  assign \new_[27488]_  = \new_[27487]_  & \new_[27482]_ ;
  assign \new_[27492]_  = A167 & A168;
  assign \new_[27493]_  = A170 & \new_[27492]_ ;
  assign \new_[27497]_  = ~A203 & ~A201;
  assign \new_[27498]_  = ~A166 & \new_[27497]_ ;
  assign \new_[27499]_  = \new_[27498]_  & \new_[27493]_ ;
  assign \new_[27503]_  = A298 & A266;
  assign \new_[27504]_  = A265 & \new_[27503]_ ;
  assign \new_[27508]_  = A301 & A300;
  assign \new_[27509]_  = ~A299 & \new_[27508]_ ;
  assign \new_[27510]_  = \new_[27509]_  & \new_[27504]_ ;
  assign \new_[27514]_  = A167 & A168;
  assign \new_[27515]_  = A170 & \new_[27514]_ ;
  assign \new_[27519]_  = ~A203 & ~A201;
  assign \new_[27520]_  = ~A166 & \new_[27519]_ ;
  assign \new_[27521]_  = \new_[27520]_  & \new_[27515]_ ;
  assign \new_[27525]_  = A298 & A266;
  assign \new_[27526]_  = A265 & \new_[27525]_ ;
  assign \new_[27530]_  = ~A302 & A300;
  assign \new_[27531]_  = ~A299 & \new_[27530]_ ;
  assign \new_[27532]_  = \new_[27531]_  & \new_[27526]_ ;
  assign \new_[27536]_  = A167 & A168;
  assign \new_[27537]_  = A170 & \new_[27536]_ ;
  assign \new_[27541]_  = ~A203 & ~A201;
  assign \new_[27542]_  = ~A166 & \new_[27541]_ ;
  assign \new_[27543]_  = \new_[27542]_  & \new_[27537]_ ;
  assign \new_[27547]_  = ~A298 & A266;
  assign \new_[27548]_  = A265 & \new_[27547]_ ;
  assign \new_[27552]_  = A301 & A300;
  assign \new_[27553]_  = A299 & \new_[27552]_ ;
  assign \new_[27554]_  = \new_[27553]_  & \new_[27548]_ ;
  assign \new_[27558]_  = A167 & A168;
  assign \new_[27559]_  = A170 & \new_[27558]_ ;
  assign \new_[27563]_  = ~A203 & ~A201;
  assign \new_[27564]_  = ~A166 & \new_[27563]_ ;
  assign \new_[27565]_  = \new_[27564]_  & \new_[27559]_ ;
  assign \new_[27569]_  = ~A298 & A266;
  assign \new_[27570]_  = A265 & \new_[27569]_ ;
  assign \new_[27574]_  = ~A302 & A300;
  assign \new_[27575]_  = A299 & \new_[27574]_ ;
  assign \new_[27576]_  = \new_[27575]_  & \new_[27570]_ ;
  assign \new_[27580]_  = A167 & A168;
  assign \new_[27581]_  = A170 & \new_[27580]_ ;
  assign \new_[27585]_  = ~A203 & ~A201;
  assign \new_[27586]_  = ~A166 & \new_[27585]_ ;
  assign \new_[27587]_  = \new_[27586]_  & \new_[27581]_ ;
  assign \new_[27591]_  = A267 & A266;
  assign \new_[27592]_  = ~A265 & \new_[27591]_ ;
  assign \new_[27596]_  = A301 & ~A300;
  assign \new_[27597]_  = A268 & \new_[27596]_ ;
  assign \new_[27598]_  = \new_[27597]_  & \new_[27592]_ ;
  assign \new_[27602]_  = A167 & A168;
  assign \new_[27603]_  = A170 & \new_[27602]_ ;
  assign \new_[27607]_  = ~A203 & ~A201;
  assign \new_[27608]_  = ~A166 & \new_[27607]_ ;
  assign \new_[27609]_  = \new_[27608]_  & \new_[27603]_ ;
  assign \new_[27613]_  = A267 & A266;
  assign \new_[27614]_  = ~A265 & \new_[27613]_ ;
  assign \new_[27618]_  = ~A302 & ~A300;
  assign \new_[27619]_  = A268 & \new_[27618]_ ;
  assign \new_[27620]_  = \new_[27619]_  & \new_[27614]_ ;
  assign \new_[27624]_  = A167 & A168;
  assign \new_[27625]_  = A170 & \new_[27624]_ ;
  assign \new_[27629]_  = ~A203 & ~A201;
  assign \new_[27630]_  = ~A166 & \new_[27629]_ ;
  assign \new_[27631]_  = \new_[27630]_  & \new_[27625]_ ;
  assign \new_[27635]_  = A267 & A266;
  assign \new_[27636]_  = ~A265 & \new_[27635]_ ;
  assign \new_[27640]_  = A299 & A298;
  assign \new_[27641]_  = A268 & \new_[27640]_ ;
  assign \new_[27642]_  = \new_[27641]_  & \new_[27636]_ ;
  assign \new_[27646]_  = A167 & A168;
  assign \new_[27647]_  = A170 & \new_[27646]_ ;
  assign \new_[27651]_  = ~A203 & ~A201;
  assign \new_[27652]_  = ~A166 & \new_[27651]_ ;
  assign \new_[27653]_  = \new_[27652]_  & \new_[27647]_ ;
  assign \new_[27657]_  = A267 & A266;
  assign \new_[27658]_  = ~A265 & \new_[27657]_ ;
  assign \new_[27662]_  = ~A299 & ~A298;
  assign \new_[27663]_  = A268 & \new_[27662]_ ;
  assign \new_[27664]_  = \new_[27663]_  & \new_[27658]_ ;
  assign \new_[27668]_  = A167 & A168;
  assign \new_[27669]_  = A170 & \new_[27668]_ ;
  assign \new_[27673]_  = ~A203 & ~A201;
  assign \new_[27674]_  = ~A166 & \new_[27673]_ ;
  assign \new_[27675]_  = \new_[27674]_  & \new_[27669]_ ;
  assign \new_[27679]_  = A267 & A266;
  assign \new_[27680]_  = ~A265 & \new_[27679]_ ;
  assign \new_[27684]_  = A301 & ~A300;
  assign \new_[27685]_  = ~A269 & \new_[27684]_ ;
  assign \new_[27686]_  = \new_[27685]_  & \new_[27680]_ ;
  assign \new_[27690]_  = A167 & A168;
  assign \new_[27691]_  = A170 & \new_[27690]_ ;
  assign \new_[27695]_  = ~A203 & ~A201;
  assign \new_[27696]_  = ~A166 & \new_[27695]_ ;
  assign \new_[27697]_  = \new_[27696]_  & \new_[27691]_ ;
  assign \new_[27701]_  = A267 & A266;
  assign \new_[27702]_  = ~A265 & \new_[27701]_ ;
  assign \new_[27706]_  = ~A302 & ~A300;
  assign \new_[27707]_  = ~A269 & \new_[27706]_ ;
  assign \new_[27708]_  = \new_[27707]_  & \new_[27702]_ ;
  assign \new_[27712]_  = A167 & A168;
  assign \new_[27713]_  = A170 & \new_[27712]_ ;
  assign \new_[27717]_  = ~A203 & ~A201;
  assign \new_[27718]_  = ~A166 & \new_[27717]_ ;
  assign \new_[27719]_  = \new_[27718]_  & \new_[27713]_ ;
  assign \new_[27723]_  = A267 & A266;
  assign \new_[27724]_  = ~A265 & \new_[27723]_ ;
  assign \new_[27728]_  = A299 & A298;
  assign \new_[27729]_  = ~A269 & \new_[27728]_ ;
  assign \new_[27730]_  = \new_[27729]_  & \new_[27724]_ ;
  assign \new_[27734]_  = A167 & A168;
  assign \new_[27735]_  = A170 & \new_[27734]_ ;
  assign \new_[27739]_  = ~A203 & ~A201;
  assign \new_[27740]_  = ~A166 & \new_[27739]_ ;
  assign \new_[27741]_  = \new_[27740]_  & \new_[27735]_ ;
  assign \new_[27745]_  = A267 & A266;
  assign \new_[27746]_  = ~A265 & \new_[27745]_ ;
  assign \new_[27750]_  = ~A299 & ~A298;
  assign \new_[27751]_  = ~A269 & \new_[27750]_ ;
  assign \new_[27752]_  = \new_[27751]_  & \new_[27746]_ ;
  assign \new_[27756]_  = A167 & A168;
  assign \new_[27757]_  = A170 & \new_[27756]_ ;
  assign \new_[27761]_  = ~A203 & ~A201;
  assign \new_[27762]_  = ~A166 & \new_[27761]_ ;
  assign \new_[27763]_  = \new_[27762]_  & \new_[27757]_ ;
  assign \new_[27767]_  = A267 & ~A266;
  assign \new_[27768]_  = A265 & \new_[27767]_ ;
  assign \new_[27772]_  = A301 & ~A300;
  assign \new_[27773]_  = A268 & \new_[27772]_ ;
  assign \new_[27774]_  = \new_[27773]_  & \new_[27768]_ ;
  assign \new_[27778]_  = A167 & A168;
  assign \new_[27779]_  = A170 & \new_[27778]_ ;
  assign \new_[27783]_  = ~A203 & ~A201;
  assign \new_[27784]_  = ~A166 & \new_[27783]_ ;
  assign \new_[27785]_  = \new_[27784]_  & \new_[27779]_ ;
  assign \new_[27789]_  = A267 & ~A266;
  assign \new_[27790]_  = A265 & \new_[27789]_ ;
  assign \new_[27794]_  = ~A302 & ~A300;
  assign \new_[27795]_  = A268 & \new_[27794]_ ;
  assign \new_[27796]_  = \new_[27795]_  & \new_[27790]_ ;
  assign \new_[27800]_  = A167 & A168;
  assign \new_[27801]_  = A170 & \new_[27800]_ ;
  assign \new_[27805]_  = ~A203 & ~A201;
  assign \new_[27806]_  = ~A166 & \new_[27805]_ ;
  assign \new_[27807]_  = \new_[27806]_  & \new_[27801]_ ;
  assign \new_[27811]_  = A267 & ~A266;
  assign \new_[27812]_  = A265 & \new_[27811]_ ;
  assign \new_[27816]_  = A299 & A298;
  assign \new_[27817]_  = A268 & \new_[27816]_ ;
  assign \new_[27818]_  = \new_[27817]_  & \new_[27812]_ ;
  assign \new_[27822]_  = A167 & A168;
  assign \new_[27823]_  = A170 & \new_[27822]_ ;
  assign \new_[27827]_  = ~A203 & ~A201;
  assign \new_[27828]_  = ~A166 & \new_[27827]_ ;
  assign \new_[27829]_  = \new_[27828]_  & \new_[27823]_ ;
  assign \new_[27833]_  = A267 & ~A266;
  assign \new_[27834]_  = A265 & \new_[27833]_ ;
  assign \new_[27838]_  = ~A299 & ~A298;
  assign \new_[27839]_  = A268 & \new_[27838]_ ;
  assign \new_[27840]_  = \new_[27839]_  & \new_[27834]_ ;
  assign \new_[27844]_  = A167 & A168;
  assign \new_[27845]_  = A170 & \new_[27844]_ ;
  assign \new_[27849]_  = ~A203 & ~A201;
  assign \new_[27850]_  = ~A166 & \new_[27849]_ ;
  assign \new_[27851]_  = \new_[27850]_  & \new_[27845]_ ;
  assign \new_[27855]_  = A267 & ~A266;
  assign \new_[27856]_  = A265 & \new_[27855]_ ;
  assign \new_[27860]_  = A301 & ~A300;
  assign \new_[27861]_  = ~A269 & \new_[27860]_ ;
  assign \new_[27862]_  = \new_[27861]_  & \new_[27856]_ ;
  assign \new_[27866]_  = A167 & A168;
  assign \new_[27867]_  = A170 & \new_[27866]_ ;
  assign \new_[27871]_  = ~A203 & ~A201;
  assign \new_[27872]_  = ~A166 & \new_[27871]_ ;
  assign \new_[27873]_  = \new_[27872]_  & \new_[27867]_ ;
  assign \new_[27877]_  = A267 & ~A266;
  assign \new_[27878]_  = A265 & \new_[27877]_ ;
  assign \new_[27882]_  = ~A302 & ~A300;
  assign \new_[27883]_  = ~A269 & \new_[27882]_ ;
  assign \new_[27884]_  = \new_[27883]_  & \new_[27878]_ ;
  assign \new_[27888]_  = A167 & A168;
  assign \new_[27889]_  = A170 & \new_[27888]_ ;
  assign \new_[27893]_  = ~A203 & ~A201;
  assign \new_[27894]_  = ~A166 & \new_[27893]_ ;
  assign \new_[27895]_  = \new_[27894]_  & \new_[27889]_ ;
  assign \new_[27899]_  = A267 & ~A266;
  assign \new_[27900]_  = A265 & \new_[27899]_ ;
  assign \new_[27904]_  = A299 & A298;
  assign \new_[27905]_  = ~A269 & \new_[27904]_ ;
  assign \new_[27906]_  = \new_[27905]_  & \new_[27900]_ ;
  assign \new_[27910]_  = A167 & A168;
  assign \new_[27911]_  = A170 & \new_[27910]_ ;
  assign \new_[27915]_  = ~A203 & ~A201;
  assign \new_[27916]_  = ~A166 & \new_[27915]_ ;
  assign \new_[27917]_  = \new_[27916]_  & \new_[27911]_ ;
  assign \new_[27921]_  = A267 & ~A266;
  assign \new_[27922]_  = A265 & \new_[27921]_ ;
  assign \new_[27926]_  = ~A299 & ~A298;
  assign \new_[27927]_  = ~A269 & \new_[27926]_ ;
  assign \new_[27928]_  = \new_[27927]_  & \new_[27922]_ ;
  assign \new_[27932]_  = A167 & A168;
  assign \new_[27933]_  = A170 & \new_[27932]_ ;
  assign \new_[27937]_  = ~A203 & ~A201;
  assign \new_[27938]_  = ~A166 & \new_[27937]_ ;
  assign \new_[27939]_  = \new_[27938]_  & \new_[27933]_ ;
  assign \new_[27943]_  = A298 & ~A266;
  assign \new_[27944]_  = ~A265 & \new_[27943]_ ;
  assign \new_[27948]_  = A301 & A300;
  assign \new_[27949]_  = ~A299 & \new_[27948]_ ;
  assign \new_[27950]_  = \new_[27949]_  & \new_[27944]_ ;
  assign \new_[27954]_  = A167 & A168;
  assign \new_[27955]_  = A170 & \new_[27954]_ ;
  assign \new_[27959]_  = ~A203 & ~A201;
  assign \new_[27960]_  = ~A166 & \new_[27959]_ ;
  assign \new_[27961]_  = \new_[27960]_  & \new_[27955]_ ;
  assign \new_[27965]_  = A298 & ~A266;
  assign \new_[27966]_  = ~A265 & \new_[27965]_ ;
  assign \new_[27970]_  = ~A302 & A300;
  assign \new_[27971]_  = ~A299 & \new_[27970]_ ;
  assign \new_[27972]_  = \new_[27971]_  & \new_[27966]_ ;
  assign \new_[27976]_  = A167 & A168;
  assign \new_[27977]_  = A170 & \new_[27976]_ ;
  assign \new_[27981]_  = ~A203 & ~A201;
  assign \new_[27982]_  = ~A166 & \new_[27981]_ ;
  assign \new_[27983]_  = \new_[27982]_  & \new_[27977]_ ;
  assign \new_[27987]_  = ~A298 & ~A266;
  assign \new_[27988]_  = ~A265 & \new_[27987]_ ;
  assign \new_[27992]_  = A301 & A300;
  assign \new_[27993]_  = A299 & \new_[27992]_ ;
  assign \new_[27994]_  = \new_[27993]_  & \new_[27988]_ ;
  assign \new_[27998]_  = A167 & A168;
  assign \new_[27999]_  = A170 & \new_[27998]_ ;
  assign \new_[28003]_  = ~A203 & ~A201;
  assign \new_[28004]_  = ~A166 & \new_[28003]_ ;
  assign \new_[28005]_  = \new_[28004]_  & \new_[27999]_ ;
  assign \new_[28009]_  = ~A298 & ~A266;
  assign \new_[28010]_  = ~A265 & \new_[28009]_ ;
  assign \new_[28014]_  = ~A302 & A300;
  assign \new_[28015]_  = A299 & \new_[28014]_ ;
  assign \new_[28016]_  = \new_[28015]_  & \new_[28010]_ ;
  assign \new_[28020]_  = A167 & A168;
  assign \new_[28021]_  = A170 & \new_[28020]_ ;
  assign \new_[28025]_  = A200 & A199;
  assign \new_[28026]_  = ~A166 & \new_[28025]_ ;
  assign \new_[28027]_  = \new_[28026]_  & \new_[28021]_ ;
  assign \new_[28031]_  = A298 & A268;
  assign \new_[28032]_  = ~A267 & \new_[28031]_ ;
  assign \new_[28036]_  = A301 & A300;
  assign \new_[28037]_  = ~A299 & \new_[28036]_ ;
  assign \new_[28038]_  = \new_[28037]_  & \new_[28032]_ ;
  assign \new_[28042]_  = A167 & A168;
  assign \new_[28043]_  = A170 & \new_[28042]_ ;
  assign \new_[28047]_  = A200 & A199;
  assign \new_[28048]_  = ~A166 & \new_[28047]_ ;
  assign \new_[28049]_  = \new_[28048]_  & \new_[28043]_ ;
  assign \new_[28053]_  = A298 & A268;
  assign \new_[28054]_  = ~A267 & \new_[28053]_ ;
  assign \new_[28058]_  = ~A302 & A300;
  assign \new_[28059]_  = ~A299 & \new_[28058]_ ;
  assign \new_[28060]_  = \new_[28059]_  & \new_[28054]_ ;
  assign \new_[28064]_  = A167 & A168;
  assign \new_[28065]_  = A170 & \new_[28064]_ ;
  assign \new_[28069]_  = A200 & A199;
  assign \new_[28070]_  = ~A166 & \new_[28069]_ ;
  assign \new_[28071]_  = \new_[28070]_  & \new_[28065]_ ;
  assign \new_[28075]_  = ~A298 & A268;
  assign \new_[28076]_  = ~A267 & \new_[28075]_ ;
  assign \new_[28080]_  = A301 & A300;
  assign \new_[28081]_  = A299 & \new_[28080]_ ;
  assign \new_[28082]_  = \new_[28081]_  & \new_[28076]_ ;
  assign \new_[28086]_  = A167 & A168;
  assign \new_[28087]_  = A170 & \new_[28086]_ ;
  assign \new_[28091]_  = A200 & A199;
  assign \new_[28092]_  = ~A166 & \new_[28091]_ ;
  assign \new_[28093]_  = \new_[28092]_  & \new_[28087]_ ;
  assign \new_[28097]_  = ~A298 & A268;
  assign \new_[28098]_  = ~A267 & \new_[28097]_ ;
  assign \new_[28102]_  = ~A302 & A300;
  assign \new_[28103]_  = A299 & \new_[28102]_ ;
  assign \new_[28104]_  = \new_[28103]_  & \new_[28098]_ ;
  assign \new_[28108]_  = A167 & A168;
  assign \new_[28109]_  = A170 & \new_[28108]_ ;
  assign \new_[28113]_  = A200 & A199;
  assign \new_[28114]_  = ~A166 & \new_[28113]_ ;
  assign \new_[28115]_  = \new_[28114]_  & \new_[28109]_ ;
  assign \new_[28119]_  = A298 & ~A269;
  assign \new_[28120]_  = ~A267 & \new_[28119]_ ;
  assign \new_[28124]_  = A301 & A300;
  assign \new_[28125]_  = ~A299 & \new_[28124]_ ;
  assign \new_[28126]_  = \new_[28125]_  & \new_[28120]_ ;
  assign \new_[28130]_  = A167 & A168;
  assign \new_[28131]_  = A170 & \new_[28130]_ ;
  assign \new_[28135]_  = A200 & A199;
  assign \new_[28136]_  = ~A166 & \new_[28135]_ ;
  assign \new_[28137]_  = \new_[28136]_  & \new_[28131]_ ;
  assign \new_[28141]_  = A298 & ~A269;
  assign \new_[28142]_  = ~A267 & \new_[28141]_ ;
  assign \new_[28146]_  = ~A302 & A300;
  assign \new_[28147]_  = ~A299 & \new_[28146]_ ;
  assign \new_[28148]_  = \new_[28147]_  & \new_[28142]_ ;
  assign \new_[28152]_  = A167 & A168;
  assign \new_[28153]_  = A170 & \new_[28152]_ ;
  assign \new_[28157]_  = A200 & A199;
  assign \new_[28158]_  = ~A166 & \new_[28157]_ ;
  assign \new_[28159]_  = \new_[28158]_  & \new_[28153]_ ;
  assign \new_[28163]_  = ~A298 & ~A269;
  assign \new_[28164]_  = ~A267 & \new_[28163]_ ;
  assign \new_[28168]_  = A301 & A300;
  assign \new_[28169]_  = A299 & \new_[28168]_ ;
  assign \new_[28170]_  = \new_[28169]_  & \new_[28164]_ ;
  assign \new_[28174]_  = A167 & A168;
  assign \new_[28175]_  = A170 & \new_[28174]_ ;
  assign \new_[28179]_  = A200 & A199;
  assign \new_[28180]_  = ~A166 & \new_[28179]_ ;
  assign \new_[28181]_  = \new_[28180]_  & \new_[28175]_ ;
  assign \new_[28185]_  = ~A298 & ~A269;
  assign \new_[28186]_  = ~A267 & \new_[28185]_ ;
  assign \new_[28190]_  = ~A302 & A300;
  assign \new_[28191]_  = A299 & \new_[28190]_ ;
  assign \new_[28192]_  = \new_[28191]_  & \new_[28186]_ ;
  assign \new_[28196]_  = A167 & A168;
  assign \new_[28197]_  = A170 & \new_[28196]_ ;
  assign \new_[28201]_  = A200 & A199;
  assign \new_[28202]_  = ~A166 & \new_[28201]_ ;
  assign \new_[28203]_  = \new_[28202]_  & \new_[28197]_ ;
  assign \new_[28207]_  = A298 & A266;
  assign \new_[28208]_  = A265 & \new_[28207]_ ;
  assign \new_[28212]_  = A301 & A300;
  assign \new_[28213]_  = ~A299 & \new_[28212]_ ;
  assign \new_[28214]_  = \new_[28213]_  & \new_[28208]_ ;
  assign \new_[28218]_  = A167 & A168;
  assign \new_[28219]_  = A170 & \new_[28218]_ ;
  assign \new_[28223]_  = A200 & A199;
  assign \new_[28224]_  = ~A166 & \new_[28223]_ ;
  assign \new_[28225]_  = \new_[28224]_  & \new_[28219]_ ;
  assign \new_[28229]_  = A298 & A266;
  assign \new_[28230]_  = A265 & \new_[28229]_ ;
  assign \new_[28234]_  = ~A302 & A300;
  assign \new_[28235]_  = ~A299 & \new_[28234]_ ;
  assign \new_[28236]_  = \new_[28235]_  & \new_[28230]_ ;
  assign \new_[28240]_  = A167 & A168;
  assign \new_[28241]_  = A170 & \new_[28240]_ ;
  assign \new_[28245]_  = A200 & A199;
  assign \new_[28246]_  = ~A166 & \new_[28245]_ ;
  assign \new_[28247]_  = \new_[28246]_  & \new_[28241]_ ;
  assign \new_[28251]_  = ~A298 & A266;
  assign \new_[28252]_  = A265 & \new_[28251]_ ;
  assign \new_[28256]_  = A301 & A300;
  assign \new_[28257]_  = A299 & \new_[28256]_ ;
  assign \new_[28258]_  = \new_[28257]_  & \new_[28252]_ ;
  assign \new_[28262]_  = A167 & A168;
  assign \new_[28263]_  = A170 & \new_[28262]_ ;
  assign \new_[28267]_  = A200 & A199;
  assign \new_[28268]_  = ~A166 & \new_[28267]_ ;
  assign \new_[28269]_  = \new_[28268]_  & \new_[28263]_ ;
  assign \new_[28273]_  = ~A298 & A266;
  assign \new_[28274]_  = A265 & \new_[28273]_ ;
  assign \new_[28278]_  = ~A302 & A300;
  assign \new_[28279]_  = A299 & \new_[28278]_ ;
  assign \new_[28280]_  = \new_[28279]_  & \new_[28274]_ ;
  assign \new_[28284]_  = A167 & A168;
  assign \new_[28285]_  = A170 & \new_[28284]_ ;
  assign \new_[28289]_  = A200 & A199;
  assign \new_[28290]_  = ~A166 & \new_[28289]_ ;
  assign \new_[28291]_  = \new_[28290]_  & \new_[28285]_ ;
  assign \new_[28295]_  = A267 & A266;
  assign \new_[28296]_  = ~A265 & \new_[28295]_ ;
  assign \new_[28300]_  = A301 & ~A300;
  assign \new_[28301]_  = A268 & \new_[28300]_ ;
  assign \new_[28302]_  = \new_[28301]_  & \new_[28296]_ ;
  assign \new_[28306]_  = A167 & A168;
  assign \new_[28307]_  = A170 & \new_[28306]_ ;
  assign \new_[28311]_  = A200 & A199;
  assign \new_[28312]_  = ~A166 & \new_[28311]_ ;
  assign \new_[28313]_  = \new_[28312]_  & \new_[28307]_ ;
  assign \new_[28317]_  = A267 & A266;
  assign \new_[28318]_  = ~A265 & \new_[28317]_ ;
  assign \new_[28322]_  = ~A302 & ~A300;
  assign \new_[28323]_  = A268 & \new_[28322]_ ;
  assign \new_[28324]_  = \new_[28323]_  & \new_[28318]_ ;
  assign \new_[28328]_  = A167 & A168;
  assign \new_[28329]_  = A170 & \new_[28328]_ ;
  assign \new_[28333]_  = A200 & A199;
  assign \new_[28334]_  = ~A166 & \new_[28333]_ ;
  assign \new_[28335]_  = \new_[28334]_  & \new_[28329]_ ;
  assign \new_[28339]_  = A267 & A266;
  assign \new_[28340]_  = ~A265 & \new_[28339]_ ;
  assign \new_[28344]_  = A299 & A298;
  assign \new_[28345]_  = A268 & \new_[28344]_ ;
  assign \new_[28346]_  = \new_[28345]_  & \new_[28340]_ ;
  assign \new_[28350]_  = A167 & A168;
  assign \new_[28351]_  = A170 & \new_[28350]_ ;
  assign \new_[28355]_  = A200 & A199;
  assign \new_[28356]_  = ~A166 & \new_[28355]_ ;
  assign \new_[28357]_  = \new_[28356]_  & \new_[28351]_ ;
  assign \new_[28361]_  = A267 & A266;
  assign \new_[28362]_  = ~A265 & \new_[28361]_ ;
  assign \new_[28366]_  = ~A299 & ~A298;
  assign \new_[28367]_  = A268 & \new_[28366]_ ;
  assign \new_[28368]_  = \new_[28367]_  & \new_[28362]_ ;
  assign \new_[28372]_  = A167 & A168;
  assign \new_[28373]_  = A170 & \new_[28372]_ ;
  assign \new_[28377]_  = A200 & A199;
  assign \new_[28378]_  = ~A166 & \new_[28377]_ ;
  assign \new_[28379]_  = \new_[28378]_  & \new_[28373]_ ;
  assign \new_[28383]_  = A267 & A266;
  assign \new_[28384]_  = ~A265 & \new_[28383]_ ;
  assign \new_[28388]_  = A301 & ~A300;
  assign \new_[28389]_  = ~A269 & \new_[28388]_ ;
  assign \new_[28390]_  = \new_[28389]_  & \new_[28384]_ ;
  assign \new_[28394]_  = A167 & A168;
  assign \new_[28395]_  = A170 & \new_[28394]_ ;
  assign \new_[28399]_  = A200 & A199;
  assign \new_[28400]_  = ~A166 & \new_[28399]_ ;
  assign \new_[28401]_  = \new_[28400]_  & \new_[28395]_ ;
  assign \new_[28405]_  = A267 & A266;
  assign \new_[28406]_  = ~A265 & \new_[28405]_ ;
  assign \new_[28410]_  = ~A302 & ~A300;
  assign \new_[28411]_  = ~A269 & \new_[28410]_ ;
  assign \new_[28412]_  = \new_[28411]_  & \new_[28406]_ ;
  assign \new_[28416]_  = A167 & A168;
  assign \new_[28417]_  = A170 & \new_[28416]_ ;
  assign \new_[28421]_  = A200 & A199;
  assign \new_[28422]_  = ~A166 & \new_[28421]_ ;
  assign \new_[28423]_  = \new_[28422]_  & \new_[28417]_ ;
  assign \new_[28427]_  = A267 & A266;
  assign \new_[28428]_  = ~A265 & \new_[28427]_ ;
  assign \new_[28432]_  = A299 & A298;
  assign \new_[28433]_  = ~A269 & \new_[28432]_ ;
  assign \new_[28434]_  = \new_[28433]_  & \new_[28428]_ ;
  assign \new_[28438]_  = A167 & A168;
  assign \new_[28439]_  = A170 & \new_[28438]_ ;
  assign \new_[28443]_  = A200 & A199;
  assign \new_[28444]_  = ~A166 & \new_[28443]_ ;
  assign \new_[28445]_  = \new_[28444]_  & \new_[28439]_ ;
  assign \new_[28449]_  = A267 & A266;
  assign \new_[28450]_  = ~A265 & \new_[28449]_ ;
  assign \new_[28454]_  = ~A299 & ~A298;
  assign \new_[28455]_  = ~A269 & \new_[28454]_ ;
  assign \new_[28456]_  = \new_[28455]_  & \new_[28450]_ ;
  assign \new_[28460]_  = A167 & A168;
  assign \new_[28461]_  = A170 & \new_[28460]_ ;
  assign \new_[28465]_  = A200 & A199;
  assign \new_[28466]_  = ~A166 & \new_[28465]_ ;
  assign \new_[28467]_  = \new_[28466]_  & \new_[28461]_ ;
  assign \new_[28471]_  = A267 & ~A266;
  assign \new_[28472]_  = A265 & \new_[28471]_ ;
  assign \new_[28476]_  = A301 & ~A300;
  assign \new_[28477]_  = A268 & \new_[28476]_ ;
  assign \new_[28478]_  = \new_[28477]_  & \new_[28472]_ ;
  assign \new_[28482]_  = A167 & A168;
  assign \new_[28483]_  = A170 & \new_[28482]_ ;
  assign \new_[28487]_  = A200 & A199;
  assign \new_[28488]_  = ~A166 & \new_[28487]_ ;
  assign \new_[28489]_  = \new_[28488]_  & \new_[28483]_ ;
  assign \new_[28493]_  = A267 & ~A266;
  assign \new_[28494]_  = A265 & \new_[28493]_ ;
  assign \new_[28498]_  = ~A302 & ~A300;
  assign \new_[28499]_  = A268 & \new_[28498]_ ;
  assign \new_[28500]_  = \new_[28499]_  & \new_[28494]_ ;
  assign \new_[28504]_  = A167 & A168;
  assign \new_[28505]_  = A170 & \new_[28504]_ ;
  assign \new_[28509]_  = A200 & A199;
  assign \new_[28510]_  = ~A166 & \new_[28509]_ ;
  assign \new_[28511]_  = \new_[28510]_  & \new_[28505]_ ;
  assign \new_[28515]_  = A267 & ~A266;
  assign \new_[28516]_  = A265 & \new_[28515]_ ;
  assign \new_[28520]_  = A299 & A298;
  assign \new_[28521]_  = A268 & \new_[28520]_ ;
  assign \new_[28522]_  = \new_[28521]_  & \new_[28516]_ ;
  assign \new_[28526]_  = A167 & A168;
  assign \new_[28527]_  = A170 & \new_[28526]_ ;
  assign \new_[28531]_  = A200 & A199;
  assign \new_[28532]_  = ~A166 & \new_[28531]_ ;
  assign \new_[28533]_  = \new_[28532]_  & \new_[28527]_ ;
  assign \new_[28537]_  = A267 & ~A266;
  assign \new_[28538]_  = A265 & \new_[28537]_ ;
  assign \new_[28542]_  = ~A299 & ~A298;
  assign \new_[28543]_  = A268 & \new_[28542]_ ;
  assign \new_[28544]_  = \new_[28543]_  & \new_[28538]_ ;
  assign \new_[28548]_  = A167 & A168;
  assign \new_[28549]_  = A170 & \new_[28548]_ ;
  assign \new_[28553]_  = A200 & A199;
  assign \new_[28554]_  = ~A166 & \new_[28553]_ ;
  assign \new_[28555]_  = \new_[28554]_  & \new_[28549]_ ;
  assign \new_[28559]_  = A267 & ~A266;
  assign \new_[28560]_  = A265 & \new_[28559]_ ;
  assign \new_[28564]_  = A301 & ~A300;
  assign \new_[28565]_  = ~A269 & \new_[28564]_ ;
  assign \new_[28566]_  = \new_[28565]_  & \new_[28560]_ ;
  assign \new_[28570]_  = A167 & A168;
  assign \new_[28571]_  = A170 & \new_[28570]_ ;
  assign \new_[28575]_  = A200 & A199;
  assign \new_[28576]_  = ~A166 & \new_[28575]_ ;
  assign \new_[28577]_  = \new_[28576]_  & \new_[28571]_ ;
  assign \new_[28581]_  = A267 & ~A266;
  assign \new_[28582]_  = A265 & \new_[28581]_ ;
  assign \new_[28586]_  = ~A302 & ~A300;
  assign \new_[28587]_  = ~A269 & \new_[28586]_ ;
  assign \new_[28588]_  = \new_[28587]_  & \new_[28582]_ ;
  assign \new_[28592]_  = A167 & A168;
  assign \new_[28593]_  = A170 & \new_[28592]_ ;
  assign \new_[28597]_  = A200 & A199;
  assign \new_[28598]_  = ~A166 & \new_[28597]_ ;
  assign \new_[28599]_  = \new_[28598]_  & \new_[28593]_ ;
  assign \new_[28603]_  = A267 & ~A266;
  assign \new_[28604]_  = A265 & \new_[28603]_ ;
  assign \new_[28608]_  = A299 & A298;
  assign \new_[28609]_  = ~A269 & \new_[28608]_ ;
  assign \new_[28610]_  = \new_[28609]_  & \new_[28604]_ ;
  assign \new_[28614]_  = A167 & A168;
  assign \new_[28615]_  = A170 & \new_[28614]_ ;
  assign \new_[28619]_  = A200 & A199;
  assign \new_[28620]_  = ~A166 & \new_[28619]_ ;
  assign \new_[28621]_  = \new_[28620]_  & \new_[28615]_ ;
  assign \new_[28625]_  = A267 & ~A266;
  assign \new_[28626]_  = A265 & \new_[28625]_ ;
  assign \new_[28630]_  = ~A299 & ~A298;
  assign \new_[28631]_  = ~A269 & \new_[28630]_ ;
  assign \new_[28632]_  = \new_[28631]_  & \new_[28626]_ ;
  assign \new_[28636]_  = A167 & A168;
  assign \new_[28637]_  = A170 & \new_[28636]_ ;
  assign \new_[28641]_  = A200 & A199;
  assign \new_[28642]_  = ~A166 & \new_[28641]_ ;
  assign \new_[28643]_  = \new_[28642]_  & \new_[28637]_ ;
  assign \new_[28647]_  = A298 & ~A266;
  assign \new_[28648]_  = ~A265 & \new_[28647]_ ;
  assign \new_[28652]_  = A301 & A300;
  assign \new_[28653]_  = ~A299 & \new_[28652]_ ;
  assign \new_[28654]_  = \new_[28653]_  & \new_[28648]_ ;
  assign \new_[28658]_  = A167 & A168;
  assign \new_[28659]_  = A170 & \new_[28658]_ ;
  assign \new_[28663]_  = A200 & A199;
  assign \new_[28664]_  = ~A166 & \new_[28663]_ ;
  assign \new_[28665]_  = \new_[28664]_  & \new_[28659]_ ;
  assign \new_[28669]_  = A298 & ~A266;
  assign \new_[28670]_  = ~A265 & \new_[28669]_ ;
  assign \new_[28674]_  = ~A302 & A300;
  assign \new_[28675]_  = ~A299 & \new_[28674]_ ;
  assign \new_[28676]_  = \new_[28675]_  & \new_[28670]_ ;
  assign \new_[28680]_  = A167 & A168;
  assign \new_[28681]_  = A170 & \new_[28680]_ ;
  assign \new_[28685]_  = A200 & A199;
  assign \new_[28686]_  = ~A166 & \new_[28685]_ ;
  assign \new_[28687]_  = \new_[28686]_  & \new_[28681]_ ;
  assign \new_[28691]_  = ~A298 & ~A266;
  assign \new_[28692]_  = ~A265 & \new_[28691]_ ;
  assign \new_[28696]_  = A301 & A300;
  assign \new_[28697]_  = A299 & \new_[28696]_ ;
  assign \new_[28698]_  = \new_[28697]_  & \new_[28692]_ ;
  assign \new_[28702]_  = A167 & A168;
  assign \new_[28703]_  = A170 & \new_[28702]_ ;
  assign \new_[28707]_  = A200 & A199;
  assign \new_[28708]_  = ~A166 & \new_[28707]_ ;
  assign \new_[28709]_  = \new_[28708]_  & \new_[28703]_ ;
  assign \new_[28713]_  = ~A298 & ~A266;
  assign \new_[28714]_  = ~A265 & \new_[28713]_ ;
  assign \new_[28718]_  = ~A302 & A300;
  assign \new_[28719]_  = A299 & \new_[28718]_ ;
  assign \new_[28720]_  = \new_[28719]_  & \new_[28714]_ ;
  assign \new_[28724]_  = A167 & A168;
  assign \new_[28725]_  = A170 & \new_[28724]_ ;
  assign \new_[28729]_  = ~A200 & ~A199;
  assign \new_[28730]_  = ~A166 & \new_[28729]_ ;
  assign \new_[28731]_  = \new_[28730]_  & \new_[28725]_ ;
  assign \new_[28735]_  = A298 & A268;
  assign \new_[28736]_  = ~A267 & \new_[28735]_ ;
  assign \new_[28740]_  = A301 & A300;
  assign \new_[28741]_  = ~A299 & \new_[28740]_ ;
  assign \new_[28742]_  = \new_[28741]_  & \new_[28736]_ ;
  assign \new_[28746]_  = A167 & A168;
  assign \new_[28747]_  = A170 & \new_[28746]_ ;
  assign \new_[28751]_  = ~A200 & ~A199;
  assign \new_[28752]_  = ~A166 & \new_[28751]_ ;
  assign \new_[28753]_  = \new_[28752]_  & \new_[28747]_ ;
  assign \new_[28757]_  = A298 & A268;
  assign \new_[28758]_  = ~A267 & \new_[28757]_ ;
  assign \new_[28762]_  = ~A302 & A300;
  assign \new_[28763]_  = ~A299 & \new_[28762]_ ;
  assign \new_[28764]_  = \new_[28763]_  & \new_[28758]_ ;
  assign \new_[28768]_  = A167 & A168;
  assign \new_[28769]_  = A170 & \new_[28768]_ ;
  assign \new_[28773]_  = ~A200 & ~A199;
  assign \new_[28774]_  = ~A166 & \new_[28773]_ ;
  assign \new_[28775]_  = \new_[28774]_  & \new_[28769]_ ;
  assign \new_[28779]_  = ~A298 & A268;
  assign \new_[28780]_  = ~A267 & \new_[28779]_ ;
  assign \new_[28784]_  = A301 & A300;
  assign \new_[28785]_  = A299 & \new_[28784]_ ;
  assign \new_[28786]_  = \new_[28785]_  & \new_[28780]_ ;
  assign \new_[28790]_  = A167 & A168;
  assign \new_[28791]_  = A170 & \new_[28790]_ ;
  assign \new_[28795]_  = ~A200 & ~A199;
  assign \new_[28796]_  = ~A166 & \new_[28795]_ ;
  assign \new_[28797]_  = \new_[28796]_  & \new_[28791]_ ;
  assign \new_[28801]_  = ~A298 & A268;
  assign \new_[28802]_  = ~A267 & \new_[28801]_ ;
  assign \new_[28806]_  = ~A302 & A300;
  assign \new_[28807]_  = A299 & \new_[28806]_ ;
  assign \new_[28808]_  = \new_[28807]_  & \new_[28802]_ ;
  assign \new_[28812]_  = A167 & A168;
  assign \new_[28813]_  = A170 & \new_[28812]_ ;
  assign \new_[28817]_  = ~A200 & ~A199;
  assign \new_[28818]_  = ~A166 & \new_[28817]_ ;
  assign \new_[28819]_  = \new_[28818]_  & \new_[28813]_ ;
  assign \new_[28823]_  = A298 & ~A269;
  assign \new_[28824]_  = ~A267 & \new_[28823]_ ;
  assign \new_[28828]_  = A301 & A300;
  assign \new_[28829]_  = ~A299 & \new_[28828]_ ;
  assign \new_[28830]_  = \new_[28829]_  & \new_[28824]_ ;
  assign \new_[28834]_  = A167 & A168;
  assign \new_[28835]_  = A170 & \new_[28834]_ ;
  assign \new_[28839]_  = ~A200 & ~A199;
  assign \new_[28840]_  = ~A166 & \new_[28839]_ ;
  assign \new_[28841]_  = \new_[28840]_  & \new_[28835]_ ;
  assign \new_[28845]_  = A298 & ~A269;
  assign \new_[28846]_  = ~A267 & \new_[28845]_ ;
  assign \new_[28850]_  = ~A302 & A300;
  assign \new_[28851]_  = ~A299 & \new_[28850]_ ;
  assign \new_[28852]_  = \new_[28851]_  & \new_[28846]_ ;
  assign \new_[28856]_  = A167 & A168;
  assign \new_[28857]_  = A170 & \new_[28856]_ ;
  assign \new_[28861]_  = ~A200 & ~A199;
  assign \new_[28862]_  = ~A166 & \new_[28861]_ ;
  assign \new_[28863]_  = \new_[28862]_  & \new_[28857]_ ;
  assign \new_[28867]_  = ~A298 & ~A269;
  assign \new_[28868]_  = ~A267 & \new_[28867]_ ;
  assign \new_[28872]_  = A301 & A300;
  assign \new_[28873]_  = A299 & \new_[28872]_ ;
  assign \new_[28874]_  = \new_[28873]_  & \new_[28868]_ ;
  assign \new_[28878]_  = A167 & A168;
  assign \new_[28879]_  = A170 & \new_[28878]_ ;
  assign \new_[28883]_  = ~A200 & ~A199;
  assign \new_[28884]_  = ~A166 & \new_[28883]_ ;
  assign \new_[28885]_  = \new_[28884]_  & \new_[28879]_ ;
  assign \new_[28889]_  = ~A298 & ~A269;
  assign \new_[28890]_  = ~A267 & \new_[28889]_ ;
  assign \new_[28894]_  = ~A302 & A300;
  assign \new_[28895]_  = A299 & \new_[28894]_ ;
  assign \new_[28896]_  = \new_[28895]_  & \new_[28890]_ ;
  assign \new_[28900]_  = A167 & A168;
  assign \new_[28901]_  = A170 & \new_[28900]_ ;
  assign \new_[28905]_  = ~A200 & ~A199;
  assign \new_[28906]_  = ~A166 & \new_[28905]_ ;
  assign \new_[28907]_  = \new_[28906]_  & \new_[28901]_ ;
  assign \new_[28911]_  = A298 & A266;
  assign \new_[28912]_  = A265 & \new_[28911]_ ;
  assign \new_[28916]_  = A301 & A300;
  assign \new_[28917]_  = ~A299 & \new_[28916]_ ;
  assign \new_[28918]_  = \new_[28917]_  & \new_[28912]_ ;
  assign \new_[28922]_  = A167 & A168;
  assign \new_[28923]_  = A170 & \new_[28922]_ ;
  assign \new_[28927]_  = ~A200 & ~A199;
  assign \new_[28928]_  = ~A166 & \new_[28927]_ ;
  assign \new_[28929]_  = \new_[28928]_  & \new_[28923]_ ;
  assign \new_[28933]_  = A298 & A266;
  assign \new_[28934]_  = A265 & \new_[28933]_ ;
  assign \new_[28938]_  = ~A302 & A300;
  assign \new_[28939]_  = ~A299 & \new_[28938]_ ;
  assign \new_[28940]_  = \new_[28939]_  & \new_[28934]_ ;
  assign \new_[28944]_  = A167 & A168;
  assign \new_[28945]_  = A170 & \new_[28944]_ ;
  assign \new_[28949]_  = ~A200 & ~A199;
  assign \new_[28950]_  = ~A166 & \new_[28949]_ ;
  assign \new_[28951]_  = \new_[28950]_  & \new_[28945]_ ;
  assign \new_[28955]_  = ~A298 & A266;
  assign \new_[28956]_  = A265 & \new_[28955]_ ;
  assign \new_[28960]_  = A301 & A300;
  assign \new_[28961]_  = A299 & \new_[28960]_ ;
  assign \new_[28962]_  = \new_[28961]_  & \new_[28956]_ ;
  assign \new_[28966]_  = A167 & A168;
  assign \new_[28967]_  = A170 & \new_[28966]_ ;
  assign \new_[28971]_  = ~A200 & ~A199;
  assign \new_[28972]_  = ~A166 & \new_[28971]_ ;
  assign \new_[28973]_  = \new_[28972]_  & \new_[28967]_ ;
  assign \new_[28977]_  = ~A298 & A266;
  assign \new_[28978]_  = A265 & \new_[28977]_ ;
  assign \new_[28982]_  = ~A302 & A300;
  assign \new_[28983]_  = A299 & \new_[28982]_ ;
  assign \new_[28984]_  = \new_[28983]_  & \new_[28978]_ ;
  assign \new_[28988]_  = A167 & A168;
  assign \new_[28989]_  = A170 & \new_[28988]_ ;
  assign \new_[28993]_  = ~A200 & ~A199;
  assign \new_[28994]_  = ~A166 & \new_[28993]_ ;
  assign \new_[28995]_  = \new_[28994]_  & \new_[28989]_ ;
  assign \new_[28999]_  = A267 & A266;
  assign \new_[29000]_  = ~A265 & \new_[28999]_ ;
  assign \new_[29004]_  = A301 & ~A300;
  assign \new_[29005]_  = A268 & \new_[29004]_ ;
  assign \new_[29006]_  = \new_[29005]_  & \new_[29000]_ ;
  assign \new_[29010]_  = A167 & A168;
  assign \new_[29011]_  = A170 & \new_[29010]_ ;
  assign \new_[29015]_  = ~A200 & ~A199;
  assign \new_[29016]_  = ~A166 & \new_[29015]_ ;
  assign \new_[29017]_  = \new_[29016]_  & \new_[29011]_ ;
  assign \new_[29021]_  = A267 & A266;
  assign \new_[29022]_  = ~A265 & \new_[29021]_ ;
  assign \new_[29026]_  = ~A302 & ~A300;
  assign \new_[29027]_  = A268 & \new_[29026]_ ;
  assign \new_[29028]_  = \new_[29027]_  & \new_[29022]_ ;
  assign \new_[29032]_  = A167 & A168;
  assign \new_[29033]_  = A170 & \new_[29032]_ ;
  assign \new_[29037]_  = ~A200 & ~A199;
  assign \new_[29038]_  = ~A166 & \new_[29037]_ ;
  assign \new_[29039]_  = \new_[29038]_  & \new_[29033]_ ;
  assign \new_[29043]_  = A267 & A266;
  assign \new_[29044]_  = ~A265 & \new_[29043]_ ;
  assign \new_[29048]_  = A299 & A298;
  assign \new_[29049]_  = A268 & \new_[29048]_ ;
  assign \new_[29050]_  = \new_[29049]_  & \new_[29044]_ ;
  assign \new_[29054]_  = A167 & A168;
  assign \new_[29055]_  = A170 & \new_[29054]_ ;
  assign \new_[29059]_  = ~A200 & ~A199;
  assign \new_[29060]_  = ~A166 & \new_[29059]_ ;
  assign \new_[29061]_  = \new_[29060]_  & \new_[29055]_ ;
  assign \new_[29065]_  = A267 & A266;
  assign \new_[29066]_  = ~A265 & \new_[29065]_ ;
  assign \new_[29070]_  = ~A299 & ~A298;
  assign \new_[29071]_  = A268 & \new_[29070]_ ;
  assign \new_[29072]_  = \new_[29071]_  & \new_[29066]_ ;
  assign \new_[29076]_  = A167 & A168;
  assign \new_[29077]_  = A170 & \new_[29076]_ ;
  assign \new_[29081]_  = ~A200 & ~A199;
  assign \new_[29082]_  = ~A166 & \new_[29081]_ ;
  assign \new_[29083]_  = \new_[29082]_  & \new_[29077]_ ;
  assign \new_[29087]_  = A267 & A266;
  assign \new_[29088]_  = ~A265 & \new_[29087]_ ;
  assign \new_[29092]_  = A301 & ~A300;
  assign \new_[29093]_  = ~A269 & \new_[29092]_ ;
  assign \new_[29094]_  = \new_[29093]_  & \new_[29088]_ ;
  assign \new_[29098]_  = A167 & A168;
  assign \new_[29099]_  = A170 & \new_[29098]_ ;
  assign \new_[29103]_  = ~A200 & ~A199;
  assign \new_[29104]_  = ~A166 & \new_[29103]_ ;
  assign \new_[29105]_  = \new_[29104]_  & \new_[29099]_ ;
  assign \new_[29109]_  = A267 & A266;
  assign \new_[29110]_  = ~A265 & \new_[29109]_ ;
  assign \new_[29114]_  = ~A302 & ~A300;
  assign \new_[29115]_  = ~A269 & \new_[29114]_ ;
  assign \new_[29116]_  = \new_[29115]_  & \new_[29110]_ ;
  assign \new_[29120]_  = A167 & A168;
  assign \new_[29121]_  = A170 & \new_[29120]_ ;
  assign \new_[29125]_  = ~A200 & ~A199;
  assign \new_[29126]_  = ~A166 & \new_[29125]_ ;
  assign \new_[29127]_  = \new_[29126]_  & \new_[29121]_ ;
  assign \new_[29131]_  = A267 & A266;
  assign \new_[29132]_  = ~A265 & \new_[29131]_ ;
  assign \new_[29136]_  = A299 & A298;
  assign \new_[29137]_  = ~A269 & \new_[29136]_ ;
  assign \new_[29138]_  = \new_[29137]_  & \new_[29132]_ ;
  assign \new_[29142]_  = A167 & A168;
  assign \new_[29143]_  = A170 & \new_[29142]_ ;
  assign \new_[29147]_  = ~A200 & ~A199;
  assign \new_[29148]_  = ~A166 & \new_[29147]_ ;
  assign \new_[29149]_  = \new_[29148]_  & \new_[29143]_ ;
  assign \new_[29153]_  = A267 & A266;
  assign \new_[29154]_  = ~A265 & \new_[29153]_ ;
  assign \new_[29158]_  = ~A299 & ~A298;
  assign \new_[29159]_  = ~A269 & \new_[29158]_ ;
  assign \new_[29160]_  = \new_[29159]_  & \new_[29154]_ ;
  assign \new_[29164]_  = A167 & A168;
  assign \new_[29165]_  = A170 & \new_[29164]_ ;
  assign \new_[29169]_  = ~A200 & ~A199;
  assign \new_[29170]_  = ~A166 & \new_[29169]_ ;
  assign \new_[29171]_  = \new_[29170]_  & \new_[29165]_ ;
  assign \new_[29175]_  = A267 & ~A266;
  assign \new_[29176]_  = A265 & \new_[29175]_ ;
  assign \new_[29180]_  = A301 & ~A300;
  assign \new_[29181]_  = A268 & \new_[29180]_ ;
  assign \new_[29182]_  = \new_[29181]_  & \new_[29176]_ ;
  assign \new_[29186]_  = A167 & A168;
  assign \new_[29187]_  = A170 & \new_[29186]_ ;
  assign \new_[29191]_  = ~A200 & ~A199;
  assign \new_[29192]_  = ~A166 & \new_[29191]_ ;
  assign \new_[29193]_  = \new_[29192]_  & \new_[29187]_ ;
  assign \new_[29197]_  = A267 & ~A266;
  assign \new_[29198]_  = A265 & \new_[29197]_ ;
  assign \new_[29202]_  = ~A302 & ~A300;
  assign \new_[29203]_  = A268 & \new_[29202]_ ;
  assign \new_[29204]_  = \new_[29203]_  & \new_[29198]_ ;
  assign \new_[29208]_  = A167 & A168;
  assign \new_[29209]_  = A170 & \new_[29208]_ ;
  assign \new_[29213]_  = ~A200 & ~A199;
  assign \new_[29214]_  = ~A166 & \new_[29213]_ ;
  assign \new_[29215]_  = \new_[29214]_  & \new_[29209]_ ;
  assign \new_[29219]_  = A267 & ~A266;
  assign \new_[29220]_  = A265 & \new_[29219]_ ;
  assign \new_[29224]_  = A299 & A298;
  assign \new_[29225]_  = A268 & \new_[29224]_ ;
  assign \new_[29226]_  = \new_[29225]_  & \new_[29220]_ ;
  assign \new_[29230]_  = A167 & A168;
  assign \new_[29231]_  = A170 & \new_[29230]_ ;
  assign \new_[29235]_  = ~A200 & ~A199;
  assign \new_[29236]_  = ~A166 & \new_[29235]_ ;
  assign \new_[29237]_  = \new_[29236]_  & \new_[29231]_ ;
  assign \new_[29241]_  = A267 & ~A266;
  assign \new_[29242]_  = A265 & \new_[29241]_ ;
  assign \new_[29246]_  = ~A299 & ~A298;
  assign \new_[29247]_  = A268 & \new_[29246]_ ;
  assign \new_[29248]_  = \new_[29247]_  & \new_[29242]_ ;
  assign \new_[29252]_  = A167 & A168;
  assign \new_[29253]_  = A170 & \new_[29252]_ ;
  assign \new_[29257]_  = ~A200 & ~A199;
  assign \new_[29258]_  = ~A166 & \new_[29257]_ ;
  assign \new_[29259]_  = \new_[29258]_  & \new_[29253]_ ;
  assign \new_[29263]_  = A267 & ~A266;
  assign \new_[29264]_  = A265 & \new_[29263]_ ;
  assign \new_[29268]_  = A301 & ~A300;
  assign \new_[29269]_  = ~A269 & \new_[29268]_ ;
  assign \new_[29270]_  = \new_[29269]_  & \new_[29264]_ ;
  assign \new_[29274]_  = A167 & A168;
  assign \new_[29275]_  = A170 & \new_[29274]_ ;
  assign \new_[29279]_  = ~A200 & ~A199;
  assign \new_[29280]_  = ~A166 & \new_[29279]_ ;
  assign \new_[29281]_  = \new_[29280]_  & \new_[29275]_ ;
  assign \new_[29285]_  = A267 & ~A266;
  assign \new_[29286]_  = A265 & \new_[29285]_ ;
  assign \new_[29290]_  = ~A302 & ~A300;
  assign \new_[29291]_  = ~A269 & \new_[29290]_ ;
  assign \new_[29292]_  = \new_[29291]_  & \new_[29286]_ ;
  assign \new_[29296]_  = A167 & A168;
  assign \new_[29297]_  = A170 & \new_[29296]_ ;
  assign \new_[29301]_  = ~A200 & ~A199;
  assign \new_[29302]_  = ~A166 & \new_[29301]_ ;
  assign \new_[29303]_  = \new_[29302]_  & \new_[29297]_ ;
  assign \new_[29307]_  = A267 & ~A266;
  assign \new_[29308]_  = A265 & \new_[29307]_ ;
  assign \new_[29312]_  = A299 & A298;
  assign \new_[29313]_  = ~A269 & \new_[29312]_ ;
  assign \new_[29314]_  = \new_[29313]_  & \new_[29308]_ ;
  assign \new_[29318]_  = A167 & A168;
  assign \new_[29319]_  = A170 & \new_[29318]_ ;
  assign \new_[29323]_  = ~A200 & ~A199;
  assign \new_[29324]_  = ~A166 & \new_[29323]_ ;
  assign \new_[29325]_  = \new_[29324]_  & \new_[29319]_ ;
  assign \new_[29329]_  = A267 & ~A266;
  assign \new_[29330]_  = A265 & \new_[29329]_ ;
  assign \new_[29334]_  = ~A299 & ~A298;
  assign \new_[29335]_  = ~A269 & \new_[29334]_ ;
  assign \new_[29336]_  = \new_[29335]_  & \new_[29330]_ ;
  assign \new_[29340]_  = A167 & A168;
  assign \new_[29341]_  = A170 & \new_[29340]_ ;
  assign \new_[29345]_  = ~A200 & ~A199;
  assign \new_[29346]_  = ~A166 & \new_[29345]_ ;
  assign \new_[29347]_  = \new_[29346]_  & \new_[29341]_ ;
  assign \new_[29351]_  = A298 & ~A266;
  assign \new_[29352]_  = ~A265 & \new_[29351]_ ;
  assign \new_[29356]_  = A301 & A300;
  assign \new_[29357]_  = ~A299 & \new_[29356]_ ;
  assign \new_[29358]_  = \new_[29357]_  & \new_[29352]_ ;
  assign \new_[29362]_  = A167 & A168;
  assign \new_[29363]_  = A170 & \new_[29362]_ ;
  assign \new_[29367]_  = ~A200 & ~A199;
  assign \new_[29368]_  = ~A166 & \new_[29367]_ ;
  assign \new_[29369]_  = \new_[29368]_  & \new_[29363]_ ;
  assign \new_[29373]_  = A298 & ~A266;
  assign \new_[29374]_  = ~A265 & \new_[29373]_ ;
  assign \new_[29378]_  = ~A302 & A300;
  assign \new_[29379]_  = ~A299 & \new_[29378]_ ;
  assign \new_[29380]_  = \new_[29379]_  & \new_[29374]_ ;
  assign \new_[29384]_  = A167 & A168;
  assign \new_[29385]_  = A170 & \new_[29384]_ ;
  assign \new_[29389]_  = ~A200 & ~A199;
  assign \new_[29390]_  = ~A166 & \new_[29389]_ ;
  assign \new_[29391]_  = \new_[29390]_  & \new_[29385]_ ;
  assign \new_[29395]_  = ~A298 & ~A266;
  assign \new_[29396]_  = ~A265 & \new_[29395]_ ;
  assign \new_[29400]_  = A301 & A300;
  assign \new_[29401]_  = A299 & \new_[29400]_ ;
  assign \new_[29402]_  = \new_[29401]_  & \new_[29396]_ ;
  assign \new_[29406]_  = A167 & A168;
  assign \new_[29407]_  = A170 & \new_[29406]_ ;
  assign \new_[29411]_  = ~A200 & ~A199;
  assign \new_[29412]_  = ~A166 & \new_[29411]_ ;
  assign \new_[29413]_  = \new_[29412]_  & \new_[29407]_ ;
  assign \new_[29417]_  = ~A298 & ~A266;
  assign \new_[29418]_  = ~A265 & \new_[29417]_ ;
  assign \new_[29422]_  = ~A302 & A300;
  assign \new_[29423]_  = A299 & \new_[29422]_ ;
  assign \new_[29424]_  = \new_[29423]_  & \new_[29418]_ ;
  assign \new_[29428]_  = ~A167 & A168;
  assign \new_[29429]_  = A170 & \new_[29428]_ ;
  assign \new_[29433]_  = A202 & ~A201;
  assign \new_[29434]_  = A166 & \new_[29433]_ ;
  assign \new_[29435]_  = \new_[29434]_  & \new_[29429]_ ;
  assign \new_[29439]_  = A298 & A268;
  assign \new_[29440]_  = ~A267 & \new_[29439]_ ;
  assign \new_[29444]_  = A301 & A300;
  assign \new_[29445]_  = ~A299 & \new_[29444]_ ;
  assign \new_[29446]_  = \new_[29445]_  & \new_[29440]_ ;
  assign \new_[29450]_  = ~A167 & A168;
  assign \new_[29451]_  = A170 & \new_[29450]_ ;
  assign \new_[29455]_  = A202 & ~A201;
  assign \new_[29456]_  = A166 & \new_[29455]_ ;
  assign \new_[29457]_  = \new_[29456]_  & \new_[29451]_ ;
  assign \new_[29461]_  = A298 & A268;
  assign \new_[29462]_  = ~A267 & \new_[29461]_ ;
  assign \new_[29466]_  = ~A302 & A300;
  assign \new_[29467]_  = ~A299 & \new_[29466]_ ;
  assign \new_[29468]_  = \new_[29467]_  & \new_[29462]_ ;
  assign \new_[29472]_  = ~A167 & A168;
  assign \new_[29473]_  = A170 & \new_[29472]_ ;
  assign \new_[29477]_  = A202 & ~A201;
  assign \new_[29478]_  = A166 & \new_[29477]_ ;
  assign \new_[29479]_  = \new_[29478]_  & \new_[29473]_ ;
  assign \new_[29483]_  = ~A298 & A268;
  assign \new_[29484]_  = ~A267 & \new_[29483]_ ;
  assign \new_[29488]_  = A301 & A300;
  assign \new_[29489]_  = A299 & \new_[29488]_ ;
  assign \new_[29490]_  = \new_[29489]_  & \new_[29484]_ ;
  assign \new_[29494]_  = ~A167 & A168;
  assign \new_[29495]_  = A170 & \new_[29494]_ ;
  assign \new_[29499]_  = A202 & ~A201;
  assign \new_[29500]_  = A166 & \new_[29499]_ ;
  assign \new_[29501]_  = \new_[29500]_  & \new_[29495]_ ;
  assign \new_[29505]_  = ~A298 & A268;
  assign \new_[29506]_  = ~A267 & \new_[29505]_ ;
  assign \new_[29510]_  = ~A302 & A300;
  assign \new_[29511]_  = A299 & \new_[29510]_ ;
  assign \new_[29512]_  = \new_[29511]_  & \new_[29506]_ ;
  assign \new_[29516]_  = ~A167 & A168;
  assign \new_[29517]_  = A170 & \new_[29516]_ ;
  assign \new_[29521]_  = A202 & ~A201;
  assign \new_[29522]_  = A166 & \new_[29521]_ ;
  assign \new_[29523]_  = \new_[29522]_  & \new_[29517]_ ;
  assign \new_[29527]_  = A298 & ~A269;
  assign \new_[29528]_  = ~A267 & \new_[29527]_ ;
  assign \new_[29532]_  = A301 & A300;
  assign \new_[29533]_  = ~A299 & \new_[29532]_ ;
  assign \new_[29534]_  = \new_[29533]_  & \new_[29528]_ ;
  assign \new_[29538]_  = ~A167 & A168;
  assign \new_[29539]_  = A170 & \new_[29538]_ ;
  assign \new_[29543]_  = A202 & ~A201;
  assign \new_[29544]_  = A166 & \new_[29543]_ ;
  assign \new_[29545]_  = \new_[29544]_  & \new_[29539]_ ;
  assign \new_[29549]_  = A298 & ~A269;
  assign \new_[29550]_  = ~A267 & \new_[29549]_ ;
  assign \new_[29554]_  = ~A302 & A300;
  assign \new_[29555]_  = ~A299 & \new_[29554]_ ;
  assign \new_[29556]_  = \new_[29555]_  & \new_[29550]_ ;
  assign \new_[29560]_  = ~A167 & A168;
  assign \new_[29561]_  = A170 & \new_[29560]_ ;
  assign \new_[29565]_  = A202 & ~A201;
  assign \new_[29566]_  = A166 & \new_[29565]_ ;
  assign \new_[29567]_  = \new_[29566]_  & \new_[29561]_ ;
  assign \new_[29571]_  = ~A298 & ~A269;
  assign \new_[29572]_  = ~A267 & \new_[29571]_ ;
  assign \new_[29576]_  = A301 & A300;
  assign \new_[29577]_  = A299 & \new_[29576]_ ;
  assign \new_[29578]_  = \new_[29577]_  & \new_[29572]_ ;
  assign \new_[29582]_  = ~A167 & A168;
  assign \new_[29583]_  = A170 & \new_[29582]_ ;
  assign \new_[29587]_  = A202 & ~A201;
  assign \new_[29588]_  = A166 & \new_[29587]_ ;
  assign \new_[29589]_  = \new_[29588]_  & \new_[29583]_ ;
  assign \new_[29593]_  = ~A298 & ~A269;
  assign \new_[29594]_  = ~A267 & \new_[29593]_ ;
  assign \new_[29598]_  = ~A302 & A300;
  assign \new_[29599]_  = A299 & \new_[29598]_ ;
  assign \new_[29600]_  = \new_[29599]_  & \new_[29594]_ ;
  assign \new_[29604]_  = ~A167 & A168;
  assign \new_[29605]_  = A170 & \new_[29604]_ ;
  assign \new_[29609]_  = A202 & ~A201;
  assign \new_[29610]_  = A166 & \new_[29609]_ ;
  assign \new_[29611]_  = \new_[29610]_  & \new_[29605]_ ;
  assign \new_[29615]_  = A298 & A266;
  assign \new_[29616]_  = A265 & \new_[29615]_ ;
  assign \new_[29620]_  = A301 & A300;
  assign \new_[29621]_  = ~A299 & \new_[29620]_ ;
  assign \new_[29622]_  = \new_[29621]_  & \new_[29616]_ ;
  assign \new_[29626]_  = ~A167 & A168;
  assign \new_[29627]_  = A170 & \new_[29626]_ ;
  assign \new_[29631]_  = A202 & ~A201;
  assign \new_[29632]_  = A166 & \new_[29631]_ ;
  assign \new_[29633]_  = \new_[29632]_  & \new_[29627]_ ;
  assign \new_[29637]_  = A298 & A266;
  assign \new_[29638]_  = A265 & \new_[29637]_ ;
  assign \new_[29642]_  = ~A302 & A300;
  assign \new_[29643]_  = ~A299 & \new_[29642]_ ;
  assign \new_[29644]_  = \new_[29643]_  & \new_[29638]_ ;
  assign \new_[29648]_  = ~A167 & A168;
  assign \new_[29649]_  = A170 & \new_[29648]_ ;
  assign \new_[29653]_  = A202 & ~A201;
  assign \new_[29654]_  = A166 & \new_[29653]_ ;
  assign \new_[29655]_  = \new_[29654]_  & \new_[29649]_ ;
  assign \new_[29659]_  = ~A298 & A266;
  assign \new_[29660]_  = A265 & \new_[29659]_ ;
  assign \new_[29664]_  = A301 & A300;
  assign \new_[29665]_  = A299 & \new_[29664]_ ;
  assign \new_[29666]_  = \new_[29665]_  & \new_[29660]_ ;
  assign \new_[29670]_  = ~A167 & A168;
  assign \new_[29671]_  = A170 & \new_[29670]_ ;
  assign \new_[29675]_  = A202 & ~A201;
  assign \new_[29676]_  = A166 & \new_[29675]_ ;
  assign \new_[29677]_  = \new_[29676]_  & \new_[29671]_ ;
  assign \new_[29681]_  = ~A298 & A266;
  assign \new_[29682]_  = A265 & \new_[29681]_ ;
  assign \new_[29686]_  = ~A302 & A300;
  assign \new_[29687]_  = A299 & \new_[29686]_ ;
  assign \new_[29688]_  = \new_[29687]_  & \new_[29682]_ ;
  assign \new_[29692]_  = ~A167 & A168;
  assign \new_[29693]_  = A170 & \new_[29692]_ ;
  assign \new_[29697]_  = A202 & ~A201;
  assign \new_[29698]_  = A166 & \new_[29697]_ ;
  assign \new_[29699]_  = \new_[29698]_  & \new_[29693]_ ;
  assign \new_[29703]_  = A267 & A266;
  assign \new_[29704]_  = ~A265 & \new_[29703]_ ;
  assign \new_[29708]_  = A301 & ~A300;
  assign \new_[29709]_  = A268 & \new_[29708]_ ;
  assign \new_[29710]_  = \new_[29709]_  & \new_[29704]_ ;
  assign \new_[29714]_  = ~A167 & A168;
  assign \new_[29715]_  = A170 & \new_[29714]_ ;
  assign \new_[29719]_  = A202 & ~A201;
  assign \new_[29720]_  = A166 & \new_[29719]_ ;
  assign \new_[29721]_  = \new_[29720]_  & \new_[29715]_ ;
  assign \new_[29725]_  = A267 & A266;
  assign \new_[29726]_  = ~A265 & \new_[29725]_ ;
  assign \new_[29730]_  = ~A302 & ~A300;
  assign \new_[29731]_  = A268 & \new_[29730]_ ;
  assign \new_[29732]_  = \new_[29731]_  & \new_[29726]_ ;
  assign \new_[29736]_  = ~A167 & A168;
  assign \new_[29737]_  = A170 & \new_[29736]_ ;
  assign \new_[29741]_  = A202 & ~A201;
  assign \new_[29742]_  = A166 & \new_[29741]_ ;
  assign \new_[29743]_  = \new_[29742]_  & \new_[29737]_ ;
  assign \new_[29747]_  = A267 & A266;
  assign \new_[29748]_  = ~A265 & \new_[29747]_ ;
  assign \new_[29752]_  = A299 & A298;
  assign \new_[29753]_  = A268 & \new_[29752]_ ;
  assign \new_[29754]_  = \new_[29753]_  & \new_[29748]_ ;
  assign \new_[29758]_  = ~A167 & A168;
  assign \new_[29759]_  = A170 & \new_[29758]_ ;
  assign \new_[29763]_  = A202 & ~A201;
  assign \new_[29764]_  = A166 & \new_[29763]_ ;
  assign \new_[29765]_  = \new_[29764]_  & \new_[29759]_ ;
  assign \new_[29769]_  = A267 & A266;
  assign \new_[29770]_  = ~A265 & \new_[29769]_ ;
  assign \new_[29774]_  = ~A299 & ~A298;
  assign \new_[29775]_  = A268 & \new_[29774]_ ;
  assign \new_[29776]_  = \new_[29775]_  & \new_[29770]_ ;
  assign \new_[29780]_  = ~A167 & A168;
  assign \new_[29781]_  = A170 & \new_[29780]_ ;
  assign \new_[29785]_  = A202 & ~A201;
  assign \new_[29786]_  = A166 & \new_[29785]_ ;
  assign \new_[29787]_  = \new_[29786]_  & \new_[29781]_ ;
  assign \new_[29791]_  = A267 & A266;
  assign \new_[29792]_  = ~A265 & \new_[29791]_ ;
  assign \new_[29796]_  = A301 & ~A300;
  assign \new_[29797]_  = ~A269 & \new_[29796]_ ;
  assign \new_[29798]_  = \new_[29797]_  & \new_[29792]_ ;
  assign \new_[29802]_  = ~A167 & A168;
  assign \new_[29803]_  = A170 & \new_[29802]_ ;
  assign \new_[29807]_  = A202 & ~A201;
  assign \new_[29808]_  = A166 & \new_[29807]_ ;
  assign \new_[29809]_  = \new_[29808]_  & \new_[29803]_ ;
  assign \new_[29813]_  = A267 & A266;
  assign \new_[29814]_  = ~A265 & \new_[29813]_ ;
  assign \new_[29818]_  = ~A302 & ~A300;
  assign \new_[29819]_  = ~A269 & \new_[29818]_ ;
  assign \new_[29820]_  = \new_[29819]_  & \new_[29814]_ ;
  assign \new_[29824]_  = ~A167 & A168;
  assign \new_[29825]_  = A170 & \new_[29824]_ ;
  assign \new_[29829]_  = A202 & ~A201;
  assign \new_[29830]_  = A166 & \new_[29829]_ ;
  assign \new_[29831]_  = \new_[29830]_  & \new_[29825]_ ;
  assign \new_[29835]_  = A267 & A266;
  assign \new_[29836]_  = ~A265 & \new_[29835]_ ;
  assign \new_[29840]_  = A299 & A298;
  assign \new_[29841]_  = ~A269 & \new_[29840]_ ;
  assign \new_[29842]_  = \new_[29841]_  & \new_[29836]_ ;
  assign \new_[29846]_  = ~A167 & A168;
  assign \new_[29847]_  = A170 & \new_[29846]_ ;
  assign \new_[29851]_  = A202 & ~A201;
  assign \new_[29852]_  = A166 & \new_[29851]_ ;
  assign \new_[29853]_  = \new_[29852]_  & \new_[29847]_ ;
  assign \new_[29857]_  = A267 & A266;
  assign \new_[29858]_  = ~A265 & \new_[29857]_ ;
  assign \new_[29862]_  = ~A299 & ~A298;
  assign \new_[29863]_  = ~A269 & \new_[29862]_ ;
  assign \new_[29864]_  = \new_[29863]_  & \new_[29858]_ ;
  assign \new_[29868]_  = ~A167 & A168;
  assign \new_[29869]_  = A170 & \new_[29868]_ ;
  assign \new_[29873]_  = A202 & ~A201;
  assign \new_[29874]_  = A166 & \new_[29873]_ ;
  assign \new_[29875]_  = \new_[29874]_  & \new_[29869]_ ;
  assign \new_[29879]_  = A267 & ~A266;
  assign \new_[29880]_  = A265 & \new_[29879]_ ;
  assign \new_[29884]_  = A301 & ~A300;
  assign \new_[29885]_  = A268 & \new_[29884]_ ;
  assign \new_[29886]_  = \new_[29885]_  & \new_[29880]_ ;
  assign \new_[29890]_  = ~A167 & A168;
  assign \new_[29891]_  = A170 & \new_[29890]_ ;
  assign \new_[29895]_  = A202 & ~A201;
  assign \new_[29896]_  = A166 & \new_[29895]_ ;
  assign \new_[29897]_  = \new_[29896]_  & \new_[29891]_ ;
  assign \new_[29901]_  = A267 & ~A266;
  assign \new_[29902]_  = A265 & \new_[29901]_ ;
  assign \new_[29906]_  = ~A302 & ~A300;
  assign \new_[29907]_  = A268 & \new_[29906]_ ;
  assign \new_[29908]_  = \new_[29907]_  & \new_[29902]_ ;
  assign \new_[29912]_  = ~A167 & A168;
  assign \new_[29913]_  = A170 & \new_[29912]_ ;
  assign \new_[29917]_  = A202 & ~A201;
  assign \new_[29918]_  = A166 & \new_[29917]_ ;
  assign \new_[29919]_  = \new_[29918]_  & \new_[29913]_ ;
  assign \new_[29923]_  = A267 & ~A266;
  assign \new_[29924]_  = A265 & \new_[29923]_ ;
  assign \new_[29928]_  = A299 & A298;
  assign \new_[29929]_  = A268 & \new_[29928]_ ;
  assign \new_[29930]_  = \new_[29929]_  & \new_[29924]_ ;
  assign \new_[29934]_  = ~A167 & A168;
  assign \new_[29935]_  = A170 & \new_[29934]_ ;
  assign \new_[29939]_  = A202 & ~A201;
  assign \new_[29940]_  = A166 & \new_[29939]_ ;
  assign \new_[29941]_  = \new_[29940]_  & \new_[29935]_ ;
  assign \new_[29945]_  = A267 & ~A266;
  assign \new_[29946]_  = A265 & \new_[29945]_ ;
  assign \new_[29950]_  = ~A299 & ~A298;
  assign \new_[29951]_  = A268 & \new_[29950]_ ;
  assign \new_[29952]_  = \new_[29951]_  & \new_[29946]_ ;
  assign \new_[29956]_  = ~A167 & A168;
  assign \new_[29957]_  = A170 & \new_[29956]_ ;
  assign \new_[29961]_  = A202 & ~A201;
  assign \new_[29962]_  = A166 & \new_[29961]_ ;
  assign \new_[29963]_  = \new_[29962]_  & \new_[29957]_ ;
  assign \new_[29967]_  = A267 & ~A266;
  assign \new_[29968]_  = A265 & \new_[29967]_ ;
  assign \new_[29972]_  = A301 & ~A300;
  assign \new_[29973]_  = ~A269 & \new_[29972]_ ;
  assign \new_[29974]_  = \new_[29973]_  & \new_[29968]_ ;
  assign \new_[29978]_  = ~A167 & A168;
  assign \new_[29979]_  = A170 & \new_[29978]_ ;
  assign \new_[29983]_  = A202 & ~A201;
  assign \new_[29984]_  = A166 & \new_[29983]_ ;
  assign \new_[29985]_  = \new_[29984]_  & \new_[29979]_ ;
  assign \new_[29989]_  = A267 & ~A266;
  assign \new_[29990]_  = A265 & \new_[29989]_ ;
  assign \new_[29994]_  = ~A302 & ~A300;
  assign \new_[29995]_  = ~A269 & \new_[29994]_ ;
  assign \new_[29996]_  = \new_[29995]_  & \new_[29990]_ ;
  assign \new_[30000]_  = ~A167 & A168;
  assign \new_[30001]_  = A170 & \new_[30000]_ ;
  assign \new_[30005]_  = A202 & ~A201;
  assign \new_[30006]_  = A166 & \new_[30005]_ ;
  assign \new_[30007]_  = \new_[30006]_  & \new_[30001]_ ;
  assign \new_[30011]_  = A267 & ~A266;
  assign \new_[30012]_  = A265 & \new_[30011]_ ;
  assign \new_[30016]_  = A299 & A298;
  assign \new_[30017]_  = ~A269 & \new_[30016]_ ;
  assign \new_[30018]_  = \new_[30017]_  & \new_[30012]_ ;
  assign \new_[30022]_  = ~A167 & A168;
  assign \new_[30023]_  = A170 & \new_[30022]_ ;
  assign \new_[30027]_  = A202 & ~A201;
  assign \new_[30028]_  = A166 & \new_[30027]_ ;
  assign \new_[30029]_  = \new_[30028]_  & \new_[30023]_ ;
  assign \new_[30033]_  = A267 & ~A266;
  assign \new_[30034]_  = A265 & \new_[30033]_ ;
  assign \new_[30038]_  = ~A299 & ~A298;
  assign \new_[30039]_  = ~A269 & \new_[30038]_ ;
  assign \new_[30040]_  = \new_[30039]_  & \new_[30034]_ ;
  assign \new_[30044]_  = ~A167 & A168;
  assign \new_[30045]_  = A170 & \new_[30044]_ ;
  assign \new_[30049]_  = A202 & ~A201;
  assign \new_[30050]_  = A166 & \new_[30049]_ ;
  assign \new_[30051]_  = \new_[30050]_  & \new_[30045]_ ;
  assign \new_[30055]_  = A298 & ~A266;
  assign \new_[30056]_  = ~A265 & \new_[30055]_ ;
  assign \new_[30060]_  = A301 & A300;
  assign \new_[30061]_  = ~A299 & \new_[30060]_ ;
  assign \new_[30062]_  = \new_[30061]_  & \new_[30056]_ ;
  assign \new_[30066]_  = ~A167 & A168;
  assign \new_[30067]_  = A170 & \new_[30066]_ ;
  assign \new_[30071]_  = A202 & ~A201;
  assign \new_[30072]_  = A166 & \new_[30071]_ ;
  assign \new_[30073]_  = \new_[30072]_  & \new_[30067]_ ;
  assign \new_[30077]_  = A298 & ~A266;
  assign \new_[30078]_  = ~A265 & \new_[30077]_ ;
  assign \new_[30082]_  = ~A302 & A300;
  assign \new_[30083]_  = ~A299 & \new_[30082]_ ;
  assign \new_[30084]_  = \new_[30083]_  & \new_[30078]_ ;
  assign \new_[30088]_  = ~A167 & A168;
  assign \new_[30089]_  = A170 & \new_[30088]_ ;
  assign \new_[30093]_  = A202 & ~A201;
  assign \new_[30094]_  = A166 & \new_[30093]_ ;
  assign \new_[30095]_  = \new_[30094]_  & \new_[30089]_ ;
  assign \new_[30099]_  = ~A298 & ~A266;
  assign \new_[30100]_  = ~A265 & \new_[30099]_ ;
  assign \new_[30104]_  = A301 & A300;
  assign \new_[30105]_  = A299 & \new_[30104]_ ;
  assign \new_[30106]_  = \new_[30105]_  & \new_[30100]_ ;
  assign \new_[30110]_  = ~A167 & A168;
  assign \new_[30111]_  = A170 & \new_[30110]_ ;
  assign \new_[30115]_  = A202 & ~A201;
  assign \new_[30116]_  = A166 & \new_[30115]_ ;
  assign \new_[30117]_  = \new_[30116]_  & \new_[30111]_ ;
  assign \new_[30121]_  = ~A298 & ~A266;
  assign \new_[30122]_  = ~A265 & \new_[30121]_ ;
  assign \new_[30126]_  = ~A302 & A300;
  assign \new_[30127]_  = A299 & \new_[30126]_ ;
  assign \new_[30128]_  = \new_[30127]_  & \new_[30122]_ ;
  assign \new_[30132]_  = ~A167 & A168;
  assign \new_[30133]_  = A170 & \new_[30132]_ ;
  assign \new_[30137]_  = ~A203 & ~A201;
  assign \new_[30138]_  = A166 & \new_[30137]_ ;
  assign \new_[30139]_  = \new_[30138]_  & \new_[30133]_ ;
  assign \new_[30143]_  = A298 & A268;
  assign \new_[30144]_  = ~A267 & \new_[30143]_ ;
  assign \new_[30148]_  = A301 & A300;
  assign \new_[30149]_  = ~A299 & \new_[30148]_ ;
  assign \new_[30150]_  = \new_[30149]_  & \new_[30144]_ ;
  assign \new_[30154]_  = ~A167 & A168;
  assign \new_[30155]_  = A170 & \new_[30154]_ ;
  assign \new_[30159]_  = ~A203 & ~A201;
  assign \new_[30160]_  = A166 & \new_[30159]_ ;
  assign \new_[30161]_  = \new_[30160]_  & \new_[30155]_ ;
  assign \new_[30165]_  = A298 & A268;
  assign \new_[30166]_  = ~A267 & \new_[30165]_ ;
  assign \new_[30170]_  = ~A302 & A300;
  assign \new_[30171]_  = ~A299 & \new_[30170]_ ;
  assign \new_[30172]_  = \new_[30171]_  & \new_[30166]_ ;
  assign \new_[30176]_  = ~A167 & A168;
  assign \new_[30177]_  = A170 & \new_[30176]_ ;
  assign \new_[30181]_  = ~A203 & ~A201;
  assign \new_[30182]_  = A166 & \new_[30181]_ ;
  assign \new_[30183]_  = \new_[30182]_  & \new_[30177]_ ;
  assign \new_[30187]_  = ~A298 & A268;
  assign \new_[30188]_  = ~A267 & \new_[30187]_ ;
  assign \new_[30192]_  = A301 & A300;
  assign \new_[30193]_  = A299 & \new_[30192]_ ;
  assign \new_[30194]_  = \new_[30193]_  & \new_[30188]_ ;
  assign \new_[30198]_  = ~A167 & A168;
  assign \new_[30199]_  = A170 & \new_[30198]_ ;
  assign \new_[30203]_  = ~A203 & ~A201;
  assign \new_[30204]_  = A166 & \new_[30203]_ ;
  assign \new_[30205]_  = \new_[30204]_  & \new_[30199]_ ;
  assign \new_[30209]_  = ~A298 & A268;
  assign \new_[30210]_  = ~A267 & \new_[30209]_ ;
  assign \new_[30214]_  = ~A302 & A300;
  assign \new_[30215]_  = A299 & \new_[30214]_ ;
  assign \new_[30216]_  = \new_[30215]_  & \new_[30210]_ ;
  assign \new_[30220]_  = ~A167 & A168;
  assign \new_[30221]_  = A170 & \new_[30220]_ ;
  assign \new_[30225]_  = ~A203 & ~A201;
  assign \new_[30226]_  = A166 & \new_[30225]_ ;
  assign \new_[30227]_  = \new_[30226]_  & \new_[30221]_ ;
  assign \new_[30231]_  = A298 & ~A269;
  assign \new_[30232]_  = ~A267 & \new_[30231]_ ;
  assign \new_[30236]_  = A301 & A300;
  assign \new_[30237]_  = ~A299 & \new_[30236]_ ;
  assign \new_[30238]_  = \new_[30237]_  & \new_[30232]_ ;
  assign \new_[30242]_  = ~A167 & A168;
  assign \new_[30243]_  = A170 & \new_[30242]_ ;
  assign \new_[30247]_  = ~A203 & ~A201;
  assign \new_[30248]_  = A166 & \new_[30247]_ ;
  assign \new_[30249]_  = \new_[30248]_  & \new_[30243]_ ;
  assign \new_[30253]_  = A298 & ~A269;
  assign \new_[30254]_  = ~A267 & \new_[30253]_ ;
  assign \new_[30258]_  = ~A302 & A300;
  assign \new_[30259]_  = ~A299 & \new_[30258]_ ;
  assign \new_[30260]_  = \new_[30259]_  & \new_[30254]_ ;
  assign \new_[30264]_  = ~A167 & A168;
  assign \new_[30265]_  = A170 & \new_[30264]_ ;
  assign \new_[30269]_  = ~A203 & ~A201;
  assign \new_[30270]_  = A166 & \new_[30269]_ ;
  assign \new_[30271]_  = \new_[30270]_  & \new_[30265]_ ;
  assign \new_[30275]_  = ~A298 & ~A269;
  assign \new_[30276]_  = ~A267 & \new_[30275]_ ;
  assign \new_[30280]_  = A301 & A300;
  assign \new_[30281]_  = A299 & \new_[30280]_ ;
  assign \new_[30282]_  = \new_[30281]_  & \new_[30276]_ ;
  assign \new_[30286]_  = ~A167 & A168;
  assign \new_[30287]_  = A170 & \new_[30286]_ ;
  assign \new_[30291]_  = ~A203 & ~A201;
  assign \new_[30292]_  = A166 & \new_[30291]_ ;
  assign \new_[30293]_  = \new_[30292]_  & \new_[30287]_ ;
  assign \new_[30297]_  = ~A298 & ~A269;
  assign \new_[30298]_  = ~A267 & \new_[30297]_ ;
  assign \new_[30302]_  = ~A302 & A300;
  assign \new_[30303]_  = A299 & \new_[30302]_ ;
  assign \new_[30304]_  = \new_[30303]_  & \new_[30298]_ ;
  assign \new_[30308]_  = ~A167 & A168;
  assign \new_[30309]_  = A170 & \new_[30308]_ ;
  assign \new_[30313]_  = ~A203 & ~A201;
  assign \new_[30314]_  = A166 & \new_[30313]_ ;
  assign \new_[30315]_  = \new_[30314]_  & \new_[30309]_ ;
  assign \new_[30319]_  = A298 & A266;
  assign \new_[30320]_  = A265 & \new_[30319]_ ;
  assign \new_[30324]_  = A301 & A300;
  assign \new_[30325]_  = ~A299 & \new_[30324]_ ;
  assign \new_[30326]_  = \new_[30325]_  & \new_[30320]_ ;
  assign \new_[30330]_  = ~A167 & A168;
  assign \new_[30331]_  = A170 & \new_[30330]_ ;
  assign \new_[30335]_  = ~A203 & ~A201;
  assign \new_[30336]_  = A166 & \new_[30335]_ ;
  assign \new_[30337]_  = \new_[30336]_  & \new_[30331]_ ;
  assign \new_[30341]_  = A298 & A266;
  assign \new_[30342]_  = A265 & \new_[30341]_ ;
  assign \new_[30346]_  = ~A302 & A300;
  assign \new_[30347]_  = ~A299 & \new_[30346]_ ;
  assign \new_[30348]_  = \new_[30347]_  & \new_[30342]_ ;
  assign \new_[30352]_  = ~A167 & A168;
  assign \new_[30353]_  = A170 & \new_[30352]_ ;
  assign \new_[30357]_  = ~A203 & ~A201;
  assign \new_[30358]_  = A166 & \new_[30357]_ ;
  assign \new_[30359]_  = \new_[30358]_  & \new_[30353]_ ;
  assign \new_[30363]_  = ~A298 & A266;
  assign \new_[30364]_  = A265 & \new_[30363]_ ;
  assign \new_[30368]_  = A301 & A300;
  assign \new_[30369]_  = A299 & \new_[30368]_ ;
  assign \new_[30370]_  = \new_[30369]_  & \new_[30364]_ ;
  assign \new_[30374]_  = ~A167 & A168;
  assign \new_[30375]_  = A170 & \new_[30374]_ ;
  assign \new_[30379]_  = ~A203 & ~A201;
  assign \new_[30380]_  = A166 & \new_[30379]_ ;
  assign \new_[30381]_  = \new_[30380]_  & \new_[30375]_ ;
  assign \new_[30385]_  = ~A298 & A266;
  assign \new_[30386]_  = A265 & \new_[30385]_ ;
  assign \new_[30390]_  = ~A302 & A300;
  assign \new_[30391]_  = A299 & \new_[30390]_ ;
  assign \new_[30392]_  = \new_[30391]_  & \new_[30386]_ ;
  assign \new_[30396]_  = ~A167 & A168;
  assign \new_[30397]_  = A170 & \new_[30396]_ ;
  assign \new_[30401]_  = ~A203 & ~A201;
  assign \new_[30402]_  = A166 & \new_[30401]_ ;
  assign \new_[30403]_  = \new_[30402]_  & \new_[30397]_ ;
  assign \new_[30407]_  = A267 & A266;
  assign \new_[30408]_  = ~A265 & \new_[30407]_ ;
  assign \new_[30412]_  = A301 & ~A300;
  assign \new_[30413]_  = A268 & \new_[30412]_ ;
  assign \new_[30414]_  = \new_[30413]_  & \new_[30408]_ ;
  assign \new_[30418]_  = ~A167 & A168;
  assign \new_[30419]_  = A170 & \new_[30418]_ ;
  assign \new_[30423]_  = ~A203 & ~A201;
  assign \new_[30424]_  = A166 & \new_[30423]_ ;
  assign \new_[30425]_  = \new_[30424]_  & \new_[30419]_ ;
  assign \new_[30429]_  = A267 & A266;
  assign \new_[30430]_  = ~A265 & \new_[30429]_ ;
  assign \new_[30434]_  = ~A302 & ~A300;
  assign \new_[30435]_  = A268 & \new_[30434]_ ;
  assign \new_[30436]_  = \new_[30435]_  & \new_[30430]_ ;
  assign \new_[30440]_  = ~A167 & A168;
  assign \new_[30441]_  = A170 & \new_[30440]_ ;
  assign \new_[30445]_  = ~A203 & ~A201;
  assign \new_[30446]_  = A166 & \new_[30445]_ ;
  assign \new_[30447]_  = \new_[30446]_  & \new_[30441]_ ;
  assign \new_[30451]_  = A267 & A266;
  assign \new_[30452]_  = ~A265 & \new_[30451]_ ;
  assign \new_[30456]_  = A299 & A298;
  assign \new_[30457]_  = A268 & \new_[30456]_ ;
  assign \new_[30458]_  = \new_[30457]_  & \new_[30452]_ ;
  assign \new_[30462]_  = ~A167 & A168;
  assign \new_[30463]_  = A170 & \new_[30462]_ ;
  assign \new_[30467]_  = ~A203 & ~A201;
  assign \new_[30468]_  = A166 & \new_[30467]_ ;
  assign \new_[30469]_  = \new_[30468]_  & \new_[30463]_ ;
  assign \new_[30473]_  = A267 & A266;
  assign \new_[30474]_  = ~A265 & \new_[30473]_ ;
  assign \new_[30478]_  = ~A299 & ~A298;
  assign \new_[30479]_  = A268 & \new_[30478]_ ;
  assign \new_[30480]_  = \new_[30479]_  & \new_[30474]_ ;
  assign \new_[30484]_  = ~A167 & A168;
  assign \new_[30485]_  = A170 & \new_[30484]_ ;
  assign \new_[30489]_  = ~A203 & ~A201;
  assign \new_[30490]_  = A166 & \new_[30489]_ ;
  assign \new_[30491]_  = \new_[30490]_  & \new_[30485]_ ;
  assign \new_[30495]_  = A267 & A266;
  assign \new_[30496]_  = ~A265 & \new_[30495]_ ;
  assign \new_[30500]_  = A301 & ~A300;
  assign \new_[30501]_  = ~A269 & \new_[30500]_ ;
  assign \new_[30502]_  = \new_[30501]_  & \new_[30496]_ ;
  assign \new_[30506]_  = ~A167 & A168;
  assign \new_[30507]_  = A170 & \new_[30506]_ ;
  assign \new_[30511]_  = ~A203 & ~A201;
  assign \new_[30512]_  = A166 & \new_[30511]_ ;
  assign \new_[30513]_  = \new_[30512]_  & \new_[30507]_ ;
  assign \new_[30517]_  = A267 & A266;
  assign \new_[30518]_  = ~A265 & \new_[30517]_ ;
  assign \new_[30522]_  = ~A302 & ~A300;
  assign \new_[30523]_  = ~A269 & \new_[30522]_ ;
  assign \new_[30524]_  = \new_[30523]_  & \new_[30518]_ ;
  assign \new_[30528]_  = ~A167 & A168;
  assign \new_[30529]_  = A170 & \new_[30528]_ ;
  assign \new_[30533]_  = ~A203 & ~A201;
  assign \new_[30534]_  = A166 & \new_[30533]_ ;
  assign \new_[30535]_  = \new_[30534]_  & \new_[30529]_ ;
  assign \new_[30539]_  = A267 & A266;
  assign \new_[30540]_  = ~A265 & \new_[30539]_ ;
  assign \new_[30544]_  = A299 & A298;
  assign \new_[30545]_  = ~A269 & \new_[30544]_ ;
  assign \new_[30546]_  = \new_[30545]_  & \new_[30540]_ ;
  assign \new_[30550]_  = ~A167 & A168;
  assign \new_[30551]_  = A170 & \new_[30550]_ ;
  assign \new_[30555]_  = ~A203 & ~A201;
  assign \new_[30556]_  = A166 & \new_[30555]_ ;
  assign \new_[30557]_  = \new_[30556]_  & \new_[30551]_ ;
  assign \new_[30561]_  = A267 & A266;
  assign \new_[30562]_  = ~A265 & \new_[30561]_ ;
  assign \new_[30566]_  = ~A299 & ~A298;
  assign \new_[30567]_  = ~A269 & \new_[30566]_ ;
  assign \new_[30568]_  = \new_[30567]_  & \new_[30562]_ ;
  assign \new_[30572]_  = ~A167 & A168;
  assign \new_[30573]_  = A170 & \new_[30572]_ ;
  assign \new_[30577]_  = ~A203 & ~A201;
  assign \new_[30578]_  = A166 & \new_[30577]_ ;
  assign \new_[30579]_  = \new_[30578]_  & \new_[30573]_ ;
  assign \new_[30583]_  = A267 & ~A266;
  assign \new_[30584]_  = A265 & \new_[30583]_ ;
  assign \new_[30588]_  = A301 & ~A300;
  assign \new_[30589]_  = A268 & \new_[30588]_ ;
  assign \new_[30590]_  = \new_[30589]_  & \new_[30584]_ ;
  assign \new_[30594]_  = ~A167 & A168;
  assign \new_[30595]_  = A170 & \new_[30594]_ ;
  assign \new_[30599]_  = ~A203 & ~A201;
  assign \new_[30600]_  = A166 & \new_[30599]_ ;
  assign \new_[30601]_  = \new_[30600]_  & \new_[30595]_ ;
  assign \new_[30605]_  = A267 & ~A266;
  assign \new_[30606]_  = A265 & \new_[30605]_ ;
  assign \new_[30610]_  = ~A302 & ~A300;
  assign \new_[30611]_  = A268 & \new_[30610]_ ;
  assign \new_[30612]_  = \new_[30611]_  & \new_[30606]_ ;
  assign \new_[30616]_  = ~A167 & A168;
  assign \new_[30617]_  = A170 & \new_[30616]_ ;
  assign \new_[30621]_  = ~A203 & ~A201;
  assign \new_[30622]_  = A166 & \new_[30621]_ ;
  assign \new_[30623]_  = \new_[30622]_  & \new_[30617]_ ;
  assign \new_[30627]_  = A267 & ~A266;
  assign \new_[30628]_  = A265 & \new_[30627]_ ;
  assign \new_[30632]_  = A299 & A298;
  assign \new_[30633]_  = A268 & \new_[30632]_ ;
  assign \new_[30634]_  = \new_[30633]_  & \new_[30628]_ ;
  assign \new_[30638]_  = ~A167 & A168;
  assign \new_[30639]_  = A170 & \new_[30638]_ ;
  assign \new_[30643]_  = ~A203 & ~A201;
  assign \new_[30644]_  = A166 & \new_[30643]_ ;
  assign \new_[30645]_  = \new_[30644]_  & \new_[30639]_ ;
  assign \new_[30649]_  = A267 & ~A266;
  assign \new_[30650]_  = A265 & \new_[30649]_ ;
  assign \new_[30654]_  = ~A299 & ~A298;
  assign \new_[30655]_  = A268 & \new_[30654]_ ;
  assign \new_[30656]_  = \new_[30655]_  & \new_[30650]_ ;
  assign \new_[30660]_  = ~A167 & A168;
  assign \new_[30661]_  = A170 & \new_[30660]_ ;
  assign \new_[30665]_  = ~A203 & ~A201;
  assign \new_[30666]_  = A166 & \new_[30665]_ ;
  assign \new_[30667]_  = \new_[30666]_  & \new_[30661]_ ;
  assign \new_[30671]_  = A267 & ~A266;
  assign \new_[30672]_  = A265 & \new_[30671]_ ;
  assign \new_[30676]_  = A301 & ~A300;
  assign \new_[30677]_  = ~A269 & \new_[30676]_ ;
  assign \new_[30678]_  = \new_[30677]_  & \new_[30672]_ ;
  assign \new_[30682]_  = ~A167 & A168;
  assign \new_[30683]_  = A170 & \new_[30682]_ ;
  assign \new_[30687]_  = ~A203 & ~A201;
  assign \new_[30688]_  = A166 & \new_[30687]_ ;
  assign \new_[30689]_  = \new_[30688]_  & \new_[30683]_ ;
  assign \new_[30693]_  = A267 & ~A266;
  assign \new_[30694]_  = A265 & \new_[30693]_ ;
  assign \new_[30698]_  = ~A302 & ~A300;
  assign \new_[30699]_  = ~A269 & \new_[30698]_ ;
  assign \new_[30700]_  = \new_[30699]_  & \new_[30694]_ ;
  assign \new_[30704]_  = ~A167 & A168;
  assign \new_[30705]_  = A170 & \new_[30704]_ ;
  assign \new_[30709]_  = ~A203 & ~A201;
  assign \new_[30710]_  = A166 & \new_[30709]_ ;
  assign \new_[30711]_  = \new_[30710]_  & \new_[30705]_ ;
  assign \new_[30715]_  = A267 & ~A266;
  assign \new_[30716]_  = A265 & \new_[30715]_ ;
  assign \new_[30720]_  = A299 & A298;
  assign \new_[30721]_  = ~A269 & \new_[30720]_ ;
  assign \new_[30722]_  = \new_[30721]_  & \new_[30716]_ ;
  assign \new_[30726]_  = ~A167 & A168;
  assign \new_[30727]_  = A170 & \new_[30726]_ ;
  assign \new_[30731]_  = ~A203 & ~A201;
  assign \new_[30732]_  = A166 & \new_[30731]_ ;
  assign \new_[30733]_  = \new_[30732]_  & \new_[30727]_ ;
  assign \new_[30737]_  = A267 & ~A266;
  assign \new_[30738]_  = A265 & \new_[30737]_ ;
  assign \new_[30742]_  = ~A299 & ~A298;
  assign \new_[30743]_  = ~A269 & \new_[30742]_ ;
  assign \new_[30744]_  = \new_[30743]_  & \new_[30738]_ ;
  assign \new_[30748]_  = ~A167 & A168;
  assign \new_[30749]_  = A170 & \new_[30748]_ ;
  assign \new_[30753]_  = ~A203 & ~A201;
  assign \new_[30754]_  = A166 & \new_[30753]_ ;
  assign \new_[30755]_  = \new_[30754]_  & \new_[30749]_ ;
  assign \new_[30759]_  = A298 & ~A266;
  assign \new_[30760]_  = ~A265 & \new_[30759]_ ;
  assign \new_[30764]_  = A301 & A300;
  assign \new_[30765]_  = ~A299 & \new_[30764]_ ;
  assign \new_[30766]_  = \new_[30765]_  & \new_[30760]_ ;
  assign \new_[30770]_  = ~A167 & A168;
  assign \new_[30771]_  = A170 & \new_[30770]_ ;
  assign \new_[30775]_  = ~A203 & ~A201;
  assign \new_[30776]_  = A166 & \new_[30775]_ ;
  assign \new_[30777]_  = \new_[30776]_  & \new_[30771]_ ;
  assign \new_[30781]_  = A298 & ~A266;
  assign \new_[30782]_  = ~A265 & \new_[30781]_ ;
  assign \new_[30786]_  = ~A302 & A300;
  assign \new_[30787]_  = ~A299 & \new_[30786]_ ;
  assign \new_[30788]_  = \new_[30787]_  & \new_[30782]_ ;
  assign \new_[30792]_  = ~A167 & A168;
  assign \new_[30793]_  = A170 & \new_[30792]_ ;
  assign \new_[30797]_  = ~A203 & ~A201;
  assign \new_[30798]_  = A166 & \new_[30797]_ ;
  assign \new_[30799]_  = \new_[30798]_  & \new_[30793]_ ;
  assign \new_[30803]_  = ~A298 & ~A266;
  assign \new_[30804]_  = ~A265 & \new_[30803]_ ;
  assign \new_[30808]_  = A301 & A300;
  assign \new_[30809]_  = A299 & \new_[30808]_ ;
  assign \new_[30810]_  = \new_[30809]_  & \new_[30804]_ ;
  assign \new_[30814]_  = ~A167 & A168;
  assign \new_[30815]_  = A170 & \new_[30814]_ ;
  assign \new_[30819]_  = ~A203 & ~A201;
  assign \new_[30820]_  = A166 & \new_[30819]_ ;
  assign \new_[30821]_  = \new_[30820]_  & \new_[30815]_ ;
  assign \new_[30825]_  = ~A298 & ~A266;
  assign \new_[30826]_  = ~A265 & \new_[30825]_ ;
  assign \new_[30830]_  = ~A302 & A300;
  assign \new_[30831]_  = A299 & \new_[30830]_ ;
  assign \new_[30832]_  = \new_[30831]_  & \new_[30826]_ ;
  assign \new_[30836]_  = ~A167 & A168;
  assign \new_[30837]_  = A170 & \new_[30836]_ ;
  assign \new_[30841]_  = A200 & A199;
  assign \new_[30842]_  = A166 & \new_[30841]_ ;
  assign \new_[30843]_  = \new_[30842]_  & \new_[30837]_ ;
  assign \new_[30847]_  = A298 & A268;
  assign \new_[30848]_  = ~A267 & \new_[30847]_ ;
  assign \new_[30852]_  = A301 & A300;
  assign \new_[30853]_  = ~A299 & \new_[30852]_ ;
  assign \new_[30854]_  = \new_[30853]_  & \new_[30848]_ ;
  assign \new_[30858]_  = ~A167 & A168;
  assign \new_[30859]_  = A170 & \new_[30858]_ ;
  assign \new_[30863]_  = A200 & A199;
  assign \new_[30864]_  = A166 & \new_[30863]_ ;
  assign \new_[30865]_  = \new_[30864]_  & \new_[30859]_ ;
  assign \new_[30869]_  = A298 & A268;
  assign \new_[30870]_  = ~A267 & \new_[30869]_ ;
  assign \new_[30874]_  = ~A302 & A300;
  assign \new_[30875]_  = ~A299 & \new_[30874]_ ;
  assign \new_[30876]_  = \new_[30875]_  & \new_[30870]_ ;
  assign \new_[30880]_  = ~A167 & A168;
  assign \new_[30881]_  = A170 & \new_[30880]_ ;
  assign \new_[30885]_  = A200 & A199;
  assign \new_[30886]_  = A166 & \new_[30885]_ ;
  assign \new_[30887]_  = \new_[30886]_  & \new_[30881]_ ;
  assign \new_[30891]_  = ~A298 & A268;
  assign \new_[30892]_  = ~A267 & \new_[30891]_ ;
  assign \new_[30896]_  = A301 & A300;
  assign \new_[30897]_  = A299 & \new_[30896]_ ;
  assign \new_[30898]_  = \new_[30897]_  & \new_[30892]_ ;
  assign \new_[30902]_  = ~A167 & A168;
  assign \new_[30903]_  = A170 & \new_[30902]_ ;
  assign \new_[30907]_  = A200 & A199;
  assign \new_[30908]_  = A166 & \new_[30907]_ ;
  assign \new_[30909]_  = \new_[30908]_  & \new_[30903]_ ;
  assign \new_[30913]_  = ~A298 & A268;
  assign \new_[30914]_  = ~A267 & \new_[30913]_ ;
  assign \new_[30918]_  = ~A302 & A300;
  assign \new_[30919]_  = A299 & \new_[30918]_ ;
  assign \new_[30920]_  = \new_[30919]_  & \new_[30914]_ ;
  assign \new_[30924]_  = ~A167 & A168;
  assign \new_[30925]_  = A170 & \new_[30924]_ ;
  assign \new_[30929]_  = A200 & A199;
  assign \new_[30930]_  = A166 & \new_[30929]_ ;
  assign \new_[30931]_  = \new_[30930]_  & \new_[30925]_ ;
  assign \new_[30935]_  = A298 & ~A269;
  assign \new_[30936]_  = ~A267 & \new_[30935]_ ;
  assign \new_[30940]_  = A301 & A300;
  assign \new_[30941]_  = ~A299 & \new_[30940]_ ;
  assign \new_[30942]_  = \new_[30941]_  & \new_[30936]_ ;
  assign \new_[30946]_  = ~A167 & A168;
  assign \new_[30947]_  = A170 & \new_[30946]_ ;
  assign \new_[30951]_  = A200 & A199;
  assign \new_[30952]_  = A166 & \new_[30951]_ ;
  assign \new_[30953]_  = \new_[30952]_  & \new_[30947]_ ;
  assign \new_[30957]_  = A298 & ~A269;
  assign \new_[30958]_  = ~A267 & \new_[30957]_ ;
  assign \new_[30962]_  = ~A302 & A300;
  assign \new_[30963]_  = ~A299 & \new_[30962]_ ;
  assign \new_[30964]_  = \new_[30963]_  & \new_[30958]_ ;
  assign \new_[30968]_  = ~A167 & A168;
  assign \new_[30969]_  = A170 & \new_[30968]_ ;
  assign \new_[30973]_  = A200 & A199;
  assign \new_[30974]_  = A166 & \new_[30973]_ ;
  assign \new_[30975]_  = \new_[30974]_  & \new_[30969]_ ;
  assign \new_[30979]_  = ~A298 & ~A269;
  assign \new_[30980]_  = ~A267 & \new_[30979]_ ;
  assign \new_[30984]_  = A301 & A300;
  assign \new_[30985]_  = A299 & \new_[30984]_ ;
  assign \new_[30986]_  = \new_[30985]_  & \new_[30980]_ ;
  assign \new_[30990]_  = ~A167 & A168;
  assign \new_[30991]_  = A170 & \new_[30990]_ ;
  assign \new_[30995]_  = A200 & A199;
  assign \new_[30996]_  = A166 & \new_[30995]_ ;
  assign \new_[30997]_  = \new_[30996]_  & \new_[30991]_ ;
  assign \new_[31001]_  = ~A298 & ~A269;
  assign \new_[31002]_  = ~A267 & \new_[31001]_ ;
  assign \new_[31006]_  = ~A302 & A300;
  assign \new_[31007]_  = A299 & \new_[31006]_ ;
  assign \new_[31008]_  = \new_[31007]_  & \new_[31002]_ ;
  assign \new_[31012]_  = ~A167 & A168;
  assign \new_[31013]_  = A170 & \new_[31012]_ ;
  assign \new_[31017]_  = A200 & A199;
  assign \new_[31018]_  = A166 & \new_[31017]_ ;
  assign \new_[31019]_  = \new_[31018]_  & \new_[31013]_ ;
  assign \new_[31023]_  = A298 & A266;
  assign \new_[31024]_  = A265 & \new_[31023]_ ;
  assign \new_[31028]_  = A301 & A300;
  assign \new_[31029]_  = ~A299 & \new_[31028]_ ;
  assign \new_[31030]_  = \new_[31029]_  & \new_[31024]_ ;
  assign \new_[31034]_  = ~A167 & A168;
  assign \new_[31035]_  = A170 & \new_[31034]_ ;
  assign \new_[31039]_  = A200 & A199;
  assign \new_[31040]_  = A166 & \new_[31039]_ ;
  assign \new_[31041]_  = \new_[31040]_  & \new_[31035]_ ;
  assign \new_[31045]_  = A298 & A266;
  assign \new_[31046]_  = A265 & \new_[31045]_ ;
  assign \new_[31050]_  = ~A302 & A300;
  assign \new_[31051]_  = ~A299 & \new_[31050]_ ;
  assign \new_[31052]_  = \new_[31051]_  & \new_[31046]_ ;
  assign \new_[31056]_  = ~A167 & A168;
  assign \new_[31057]_  = A170 & \new_[31056]_ ;
  assign \new_[31061]_  = A200 & A199;
  assign \new_[31062]_  = A166 & \new_[31061]_ ;
  assign \new_[31063]_  = \new_[31062]_  & \new_[31057]_ ;
  assign \new_[31067]_  = ~A298 & A266;
  assign \new_[31068]_  = A265 & \new_[31067]_ ;
  assign \new_[31072]_  = A301 & A300;
  assign \new_[31073]_  = A299 & \new_[31072]_ ;
  assign \new_[31074]_  = \new_[31073]_  & \new_[31068]_ ;
  assign \new_[31078]_  = ~A167 & A168;
  assign \new_[31079]_  = A170 & \new_[31078]_ ;
  assign \new_[31083]_  = A200 & A199;
  assign \new_[31084]_  = A166 & \new_[31083]_ ;
  assign \new_[31085]_  = \new_[31084]_  & \new_[31079]_ ;
  assign \new_[31089]_  = ~A298 & A266;
  assign \new_[31090]_  = A265 & \new_[31089]_ ;
  assign \new_[31094]_  = ~A302 & A300;
  assign \new_[31095]_  = A299 & \new_[31094]_ ;
  assign \new_[31096]_  = \new_[31095]_  & \new_[31090]_ ;
  assign \new_[31100]_  = ~A167 & A168;
  assign \new_[31101]_  = A170 & \new_[31100]_ ;
  assign \new_[31105]_  = A200 & A199;
  assign \new_[31106]_  = A166 & \new_[31105]_ ;
  assign \new_[31107]_  = \new_[31106]_  & \new_[31101]_ ;
  assign \new_[31111]_  = A267 & A266;
  assign \new_[31112]_  = ~A265 & \new_[31111]_ ;
  assign \new_[31116]_  = A301 & ~A300;
  assign \new_[31117]_  = A268 & \new_[31116]_ ;
  assign \new_[31118]_  = \new_[31117]_  & \new_[31112]_ ;
  assign \new_[31122]_  = ~A167 & A168;
  assign \new_[31123]_  = A170 & \new_[31122]_ ;
  assign \new_[31127]_  = A200 & A199;
  assign \new_[31128]_  = A166 & \new_[31127]_ ;
  assign \new_[31129]_  = \new_[31128]_  & \new_[31123]_ ;
  assign \new_[31133]_  = A267 & A266;
  assign \new_[31134]_  = ~A265 & \new_[31133]_ ;
  assign \new_[31138]_  = ~A302 & ~A300;
  assign \new_[31139]_  = A268 & \new_[31138]_ ;
  assign \new_[31140]_  = \new_[31139]_  & \new_[31134]_ ;
  assign \new_[31144]_  = ~A167 & A168;
  assign \new_[31145]_  = A170 & \new_[31144]_ ;
  assign \new_[31149]_  = A200 & A199;
  assign \new_[31150]_  = A166 & \new_[31149]_ ;
  assign \new_[31151]_  = \new_[31150]_  & \new_[31145]_ ;
  assign \new_[31155]_  = A267 & A266;
  assign \new_[31156]_  = ~A265 & \new_[31155]_ ;
  assign \new_[31160]_  = A299 & A298;
  assign \new_[31161]_  = A268 & \new_[31160]_ ;
  assign \new_[31162]_  = \new_[31161]_  & \new_[31156]_ ;
  assign \new_[31166]_  = ~A167 & A168;
  assign \new_[31167]_  = A170 & \new_[31166]_ ;
  assign \new_[31171]_  = A200 & A199;
  assign \new_[31172]_  = A166 & \new_[31171]_ ;
  assign \new_[31173]_  = \new_[31172]_  & \new_[31167]_ ;
  assign \new_[31177]_  = A267 & A266;
  assign \new_[31178]_  = ~A265 & \new_[31177]_ ;
  assign \new_[31182]_  = ~A299 & ~A298;
  assign \new_[31183]_  = A268 & \new_[31182]_ ;
  assign \new_[31184]_  = \new_[31183]_  & \new_[31178]_ ;
  assign \new_[31188]_  = ~A167 & A168;
  assign \new_[31189]_  = A170 & \new_[31188]_ ;
  assign \new_[31193]_  = A200 & A199;
  assign \new_[31194]_  = A166 & \new_[31193]_ ;
  assign \new_[31195]_  = \new_[31194]_  & \new_[31189]_ ;
  assign \new_[31199]_  = A267 & A266;
  assign \new_[31200]_  = ~A265 & \new_[31199]_ ;
  assign \new_[31204]_  = A301 & ~A300;
  assign \new_[31205]_  = ~A269 & \new_[31204]_ ;
  assign \new_[31206]_  = \new_[31205]_  & \new_[31200]_ ;
  assign \new_[31210]_  = ~A167 & A168;
  assign \new_[31211]_  = A170 & \new_[31210]_ ;
  assign \new_[31215]_  = A200 & A199;
  assign \new_[31216]_  = A166 & \new_[31215]_ ;
  assign \new_[31217]_  = \new_[31216]_  & \new_[31211]_ ;
  assign \new_[31221]_  = A267 & A266;
  assign \new_[31222]_  = ~A265 & \new_[31221]_ ;
  assign \new_[31226]_  = ~A302 & ~A300;
  assign \new_[31227]_  = ~A269 & \new_[31226]_ ;
  assign \new_[31228]_  = \new_[31227]_  & \new_[31222]_ ;
  assign \new_[31232]_  = ~A167 & A168;
  assign \new_[31233]_  = A170 & \new_[31232]_ ;
  assign \new_[31237]_  = A200 & A199;
  assign \new_[31238]_  = A166 & \new_[31237]_ ;
  assign \new_[31239]_  = \new_[31238]_  & \new_[31233]_ ;
  assign \new_[31243]_  = A267 & A266;
  assign \new_[31244]_  = ~A265 & \new_[31243]_ ;
  assign \new_[31248]_  = A299 & A298;
  assign \new_[31249]_  = ~A269 & \new_[31248]_ ;
  assign \new_[31250]_  = \new_[31249]_  & \new_[31244]_ ;
  assign \new_[31254]_  = ~A167 & A168;
  assign \new_[31255]_  = A170 & \new_[31254]_ ;
  assign \new_[31259]_  = A200 & A199;
  assign \new_[31260]_  = A166 & \new_[31259]_ ;
  assign \new_[31261]_  = \new_[31260]_  & \new_[31255]_ ;
  assign \new_[31265]_  = A267 & A266;
  assign \new_[31266]_  = ~A265 & \new_[31265]_ ;
  assign \new_[31270]_  = ~A299 & ~A298;
  assign \new_[31271]_  = ~A269 & \new_[31270]_ ;
  assign \new_[31272]_  = \new_[31271]_  & \new_[31266]_ ;
  assign \new_[31276]_  = ~A167 & A168;
  assign \new_[31277]_  = A170 & \new_[31276]_ ;
  assign \new_[31281]_  = A200 & A199;
  assign \new_[31282]_  = A166 & \new_[31281]_ ;
  assign \new_[31283]_  = \new_[31282]_  & \new_[31277]_ ;
  assign \new_[31287]_  = A267 & ~A266;
  assign \new_[31288]_  = A265 & \new_[31287]_ ;
  assign \new_[31292]_  = A301 & ~A300;
  assign \new_[31293]_  = A268 & \new_[31292]_ ;
  assign \new_[31294]_  = \new_[31293]_  & \new_[31288]_ ;
  assign \new_[31298]_  = ~A167 & A168;
  assign \new_[31299]_  = A170 & \new_[31298]_ ;
  assign \new_[31303]_  = A200 & A199;
  assign \new_[31304]_  = A166 & \new_[31303]_ ;
  assign \new_[31305]_  = \new_[31304]_  & \new_[31299]_ ;
  assign \new_[31309]_  = A267 & ~A266;
  assign \new_[31310]_  = A265 & \new_[31309]_ ;
  assign \new_[31314]_  = ~A302 & ~A300;
  assign \new_[31315]_  = A268 & \new_[31314]_ ;
  assign \new_[31316]_  = \new_[31315]_  & \new_[31310]_ ;
  assign \new_[31320]_  = ~A167 & A168;
  assign \new_[31321]_  = A170 & \new_[31320]_ ;
  assign \new_[31325]_  = A200 & A199;
  assign \new_[31326]_  = A166 & \new_[31325]_ ;
  assign \new_[31327]_  = \new_[31326]_  & \new_[31321]_ ;
  assign \new_[31331]_  = A267 & ~A266;
  assign \new_[31332]_  = A265 & \new_[31331]_ ;
  assign \new_[31336]_  = A299 & A298;
  assign \new_[31337]_  = A268 & \new_[31336]_ ;
  assign \new_[31338]_  = \new_[31337]_  & \new_[31332]_ ;
  assign \new_[31342]_  = ~A167 & A168;
  assign \new_[31343]_  = A170 & \new_[31342]_ ;
  assign \new_[31347]_  = A200 & A199;
  assign \new_[31348]_  = A166 & \new_[31347]_ ;
  assign \new_[31349]_  = \new_[31348]_  & \new_[31343]_ ;
  assign \new_[31353]_  = A267 & ~A266;
  assign \new_[31354]_  = A265 & \new_[31353]_ ;
  assign \new_[31358]_  = ~A299 & ~A298;
  assign \new_[31359]_  = A268 & \new_[31358]_ ;
  assign \new_[31360]_  = \new_[31359]_  & \new_[31354]_ ;
  assign \new_[31364]_  = ~A167 & A168;
  assign \new_[31365]_  = A170 & \new_[31364]_ ;
  assign \new_[31369]_  = A200 & A199;
  assign \new_[31370]_  = A166 & \new_[31369]_ ;
  assign \new_[31371]_  = \new_[31370]_  & \new_[31365]_ ;
  assign \new_[31375]_  = A267 & ~A266;
  assign \new_[31376]_  = A265 & \new_[31375]_ ;
  assign \new_[31380]_  = A301 & ~A300;
  assign \new_[31381]_  = ~A269 & \new_[31380]_ ;
  assign \new_[31382]_  = \new_[31381]_  & \new_[31376]_ ;
  assign \new_[31386]_  = ~A167 & A168;
  assign \new_[31387]_  = A170 & \new_[31386]_ ;
  assign \new_[31391]_  = A200 & A199;
  assign \new_[31392]_  = A166 & \new_[31391]_ ;
  assign \new_[31393]_  = \new_[31392]_  & \new_[31387]_ ;
  assign \new_[31397]_  = A267 & ~A266;
  assign \new_[31398]_  = A265 & \new_[31397]_ ;
  assign \new_[31402]_  = ~A302 & ~A300;
  assign \new_[31403]_  = ~A269 & \new_[31402]_ ;
  assign \new_[31404]_  = \new_[31403]_  & \new_[31398]_ ;
  assign \new_[31408]_  = ~A167 & A168;
  assign \new_[31409]_  = A170 & \new_[31408]_ ;
  assign \new_[31413]_  = A200 & A199;
  assign \new_[31414]_  = A166 & \new_[31413]_ ;
  assign \new_[31415]_  = \new_[31414]_  & \new_[31409]_ ;
  assign \new_[31419]_  = A267 & ~A266;
  assign \new_[31420]_  = A265 & \new_[31419]_ ;
  assign \new_[31424]_  = A299 & A298;
  assign \new_[31425]_  = ~A269 & \new_[31424]_ ;
  assign \new_[31426]_  = \new_[31425]_  & \new_[31420]_ ;
  assign \new_[31430]_  = ~A167 & A168;
  assign \new_[31431]_  = A170 & \new_[31430]_ ;
  assign \new_[31435]_  = A200 & A199;
  assign \new_[31436]_  = A166 & \new_[31435]_ ;
  assign \new_[31437]_  = \new_[31436]_  & \new_[31431]_ ;
  assign \new_[31441]_  = A267 & ~A266;
  assign \new_[31442]_  = A265 & \new_[31441]_ ;
  assign \new_[31446]_  = ~A299 & ~A298;
  assign \new_[31447]_  = ~A269 & \new_[31446]_ ;
  assign \new_[31448]_  = \new_[31447]_  & \new_[31442]_ ;
  assign \new_[31452]_  = ~A167 & A168;
  assign \new_[31453]_  = A170 & \new_[31452]_ ;
  assign \new_[31457]_  = A200 & A199;
  assign \new_[31458]_  = A166 & \new_[31457]_ ;
  assign \new_[31459]_  = \new_[31458]_  & \new_[31453]_ ;
  assign \new_[31463]_  = A298 & ~A266;
  assign \new_[31464]_  = ~A265 & \new_[31463]_ ;
  assign \new_[31468]_  = A301 & A300;
  assign \new_[31469]_  = ~A299 & \new_[31468]_ ;
  assign \new_[31470]_  = \new_[31469]_  & \new_[31464]_ ;
  assign \new_[31474]_  = ~A167 & A168;
  assign \new_[31475]_  = A170 & \new_[31474]_ ;
  assign \new_[31479]_  = A200 & A199;
  assign \new_[31480]_  = A166 & \new_[31479]_ ;
  assign \new_[31481]_  = \new_[31480]_  & \new_[31475]_ ;
  assign \new_[31485]_  = A298 & ~A266;
  assign \new_[31486]_  = ~A265 & \new_[31485]_ ;
  assign \new_[31490]_  = ~A302 & A300;
  assign \new_[31491]_  = ~A299 & \new_[31490]_ ;
  assign \new_[31492]_  = \new_[31491]_  & \new_[31486]_ ;
  assign \new_[31496]_  = ~A167 & A168;
  assign \new_[31497]_  = A170 & \new_[31496]_ ;
  assign \new_[31501]_  = A200 & A199;
  assign \new_[31502]_  = A166 & \new_[31501]_ ;
  assign \new_[31503]_  = \new_[31502]_  & \new_[31497]_ ;
  assign \new_[31507]_  = ~A298 & ~A266;
  assign \new_[31508]_  = ~A265 & \new_[31507]_ ;
  assign \new_[31512]_  = A301 & A300;
  assign \new_[31513]_  = A299 & \new_[31512]_ ;
  assign \new_[31514]_  = \new_[31513]_  & \new_[31508]_ ;
  assign \new_[31518]_  = ~A167 & A168;
  assign \new_[31519]_  = A170 & \new_[31518]_ ;
  assign \new_[31523]_  = A200 & A199;
  assign \new_[31524]_  = A166 & \new_[31523]_ ;
  assign \new_[31525]_  = \new_[31524]_  & \new_[31519]_ ;
  assign \new_[31529]_  = ~A298 & ~A266;
  assign \new_[31530]_  = ~A265 & \new_[31529]_ ;
  assign \new_[31534]_  = ~A302 & A300;
  assign \new_[31535]_  = A299 & \new_[31534]_ ;
  assign \new_[31536]_  = \new_[31535]_  & \new_[31530]_ ;
  assign \new_[31540]_  = ~A167 & A168;
  assign \new_[31541]_  = A170 & \new_[31540]_ ;
  assign \new_[31545]_  = ~A200 & ~A199;
  assign \new_[31546]_  = A166 & \new_[31545]_ ;
  assign \new_[31547]_  = \new_[31546]_  & \new_[31541]_ ;
  assign \new_[31551]_  = A298 & A268;
  assign \new_[31552]_  = ~A267 & \new_[31551]_ ;
  assign \new_[31556]_  = A301 & A300;
  assign \new_[31557]_  = ~A299 & \new_[31556]_ ;
  assign \new_[31558]_  = \new_[31557]_  & \new_[31552]_ ;
  assign \new_[31562]_  = ~A167 & A168;
  assign \new_[31563]_  = A170 & \new_[31562]_ ;
  assign \new_[31567]_  = ~A200 & ~A199;
  assign \new_[31568]_  = A166 & \new_[31567]_ ;
  assign \new_[31569]_  = \new_[31568]_  & \new_[31563]_ ;
  assign \new_[31573]_  = A298 & A268;
  assign \new_[31574]_  = ~A267 & \new_[31573]_ ;
  assign \new_[31578]_  = ~A302 & A300;
  assign \new_[31579]_  = ~A299 & \new_[31578]_ ;
  assign \new_[31580]_  = \new_[31579]_  & \new_[31574]_ ;
  assign \new_[31584]_  = ~A167 & A168;
  assign \new_[31585]_  = A170 & \new_[31584]_ ;
  assign \new_[31589]_  = ~A200 & ~A199;
  assign \new_[31590]_  = A166 & \new_[31589]_ ;
  assign \new_[31591]_  = \new_[31590]_  & \new_[31585]_ ;
  assign \new_[31595]_  = ~A298 & A268;
  assign \new_[31596]_  = ~A267 & \new_[31595]_ ;
  assign \new_[31600]_  = A301 & A300;
  assign \new_[31601]_  = A299 & \new_[31600]_ ;
  assign \new_[31602]_  = \new_[31601]_  & \new_[31596]_ ;
  assign \new_[31606]_  = ~A167 & A168;
  assign \new_[31607]_  = A170 & \new_[31606]_ ;
  assign \new_[31611]_  = ~A200 & ~A199;
  assign \new_[31612]_  = A166 & \new_[31611]_ ;
  assign \new_[31613]_  = \new_[31612]_  & \new_[31607]_ ;
  assign \new_[31617]_  = ~A298 & A268;
  assign \new_[31618]_  = ~A267 & \new_[31617]_ ;
  assign \new_[31622]_  = ~A302 & A300;
  assign \new_[31623]_  = A299 & \new_[31622]_ ;
  assign \new_[31624]_  = \new_[31623]_  & \new_[31618]_ ;
  assign \new_[31628]_  = ~A167 & A168;
  assign \new_[31629]_  = A170 & \new_[31628]_ ;
  assign \new_[31633]_  = ~A200 & ~A199;
  assign \new_[31634]_  = A166 & \new_[31633]_ ;
  assign \new_[31635]_  = \new_[31634]_  & \new_[31629]_ ;
  assign \new_[31639]_  = A298 & ~A269;
  assign \new_[31640]_  = ~A267 & \new_[31639]_ ;
  assign \new_[31644]_  = A301 & A300;
  assign \new_[31645]_  = ~A299 & \new_[31644]_ ;
  assign \new_[31646]_  = \new_[31645]_  & \new_[31640]_ ;
  assign \new_[31650]_  = ~A167 & A168;
  assign \new_[31651]_  = A170 & \new_[31650]_ ;
  assign \new_[31655]_  = ~A200 & ~A199;
  assign \new_[31656]_  = A166 & \new_[31655]_ ;
  assign \new_[31657]_  = \new_[31656]_  & \new_[31651]_ ;
  assign \new_[31661]_  = A298 & ~A269;
  assign \new_[31662]_  = ~A267 & \new_[31661]_ ;
  assign \new_[31666]_  = ~A302 & A300;
  assign \new_[31667]_  = ~A299 & \new_[31666]_ ;
  assign \new_[31668]_  = \new_[31667]_  & \new_[31662]_ ;
  assign \new_[31672]_  = ~A167 & A168;
  assign \new_[31673]_  = A170 & \new_[31672]_ ;
  assign \new_[31677]_  = ~A200 & ~A199;
  assign \new_[31678]_  = A166 & \new_[31677]_ ;
  assign \new_[31679]_  = \new_[31678]_  & \new_[31673]_ ;
  assign \new_[31683]_  = ~A298 & ~A269;
  assign \new_[31684]_  = ~A267 & \new_[31683]_ ;
  assign \new_[31688]_  = A301 & A300;
  assign \new_[31689]_  = A299 & \new_[31688]_ ;
  assign \new_[31690]_  = \new_[31689]_  & \new_[31684]_ ;
  assign \new_[31694]_  = ~A167 & A168;
  assign \new_[31695]_  = A170 & \new_[31694]_ ;
  assign \new_[31699]_  = ~A200 & ~A199;
  assign \new_[31700]_  = A166 & \new_[31699]_ ;
  assign \new_[31701]_  = \new_[31700]_  & \new_[31695]_ ;
  assign \new_[31705]_  = ~A298 & ~A269;
  assign \new_[31706]_  = ~A267 & \new_[31705]_ ;
  assign \new_[31710]_  = ~A302 & A300;
  assign \new_[31711]_  = A299 & \new_[31710]_ ;
  assign \new_[31712]_  = \new_[31711]_  & \new_[31706]_ ;
  assign \new_[31716]_  = ~A167 & A168;
  assign \new_[31717]_  = A170 & \new_[31716]_ ;
  assign \new_[31721]_  = ~A200 & ~A199;
  assign \new_[31722]_  = A166 & \new_[31721]_ ;
  assign \new_[31723]_  = \new_[31722]_  & \new_[31717]_ ;
  assign \new_[31727]_  = A298 & A266;
  assign \new_[31728]_  = A265 & \new_[31727]_ ;
  assign \new_[31732]_  = A301 & A300;
  assign \new_[31733]_  = ~A299 & \new_[31732]_ ;
  assign \new_[31734]_  = \new_[31733]_  & \new_[31728]_ ;
  assign \new_[31738]_  = ~A167 & A168;
  assign \new_[31739]_  = A170 & \new_[31738]_ ;
  assign \new_[31743]_  = ~A200 & ~A199;
  assign \new_[31744]_  = A166 & \new_[31743]_ ;
  assign \new_[31745]_  = \new_[31744]_  & \new_[31739]_ ;
  assign \new_[31749]_  = A298 & A266;
  assign \new_[31750]_  = A265 & \new_[31749]_ ;
  assign \new_[31754]_  = ~A302 & A300;
  assign \new_[31755]_  = ~A299 & \new_[31754]_ ;
  assign \new_[31756]_  = \new_[31755]_  & \new_[31750]_ ;
  assign \new_[31760]_  = ~A167 & A168;
  assign \new_[31761]_  = A170 & \new_[31760]_ ;
  assign \new_[31765]_  = ~A200 & ~A199;
  assign \new_[31766]_  = A166 & \new_[31765]_ ;
  assign \new_[31767]_  = \new_[31766]_  & \new_[31761]_ ;
  assign \new_[31771]_  = ~A298 & A266;
  assign \new_[31772]_  = A265 & \new_[31771]_ ;
  assign \new_[31776]_  = A301 & A300;
  assign \new_[31777]_  = A299 & \new_[31776]_ ;
  assign \new_[31778]_  = \new_[31777]_  & \new_[31772]_ ;
  assign \new_[31782]_  = ~A167 & A168;
  assign \new_[31783]_  = A170 & \new_[31782]_ ;
  assign \new_[31787]_  = ~A200 & ~A199;
  assign \new_[31788]_  = A166 & \new_[31787]_ ;
  assign \new_[31789]_  = \new_[31788]_  & \new_[31783]_ ;
  assign \new_[31793]_  = ~A298 & A266;
  assign \new_[31794]_  = A265 & \new_[31793]_ ;
  assign \new_[31798]_  = ~A302 & A300;
  assign \new_[31799]_  = A299 & \new_[31798]_ ;
  assign \new_[31800]_  = \new_[31799]_  & \new_[31794]_ ;
  assign \new_[31804]_  = ~A167 & A168;
  assign \new_[31805]_  = A170 & \new_[31804]_ ;
  assign \new_[31809]_  = ~A200 & ~A199;
  assign \new_[31810]_  = A166 & \new_[31809]_ ;
  assign \new_[31811]_  = \new_[31810]_  & \new_[31805]_ ;
  assign \new_[31815]_  = A267 & A266;
  assign \new_[31816]_  = ~A265 & \new_[31815]_ ;
  assign \new_[31820]_  = A301 & ~A300;
  assign \new_[31821]_  = A268 & \new_[31820]_ ;
  assign \new_[31822]_  = \new_[31821]_  & \new_[31816]_ ;
  assign \new_[31826]_  = ~A167 & A168;
  assign \new_[31827]_  = A170 & \new_[31826]_ ;
  assign \new_[31831]_  = ~A200 & ~A199;
  assign \new_[31832]_  = A166 & \new_[31831]_ ;
  assign \new_[31833]_  = \new_[31832]_  & \new_[31827]_ ;
  assign \new_[31837]_  = A267 & A266;
  assign \new_[31838]_  = ~A265 & \new_[31837]_ ;
  assign \new_[31842]_  = ~A302 & ~A300;
  assign \new_[31843]_  = A268 & \new_[31842]_ ;
  assign \new_[31844]_  = \new_[31843]_  & \new_[31838]_ ;
  assign \new_[31848]_  = ~A167 & A168;
  assign \new_[31849]_  = A170 & \new_[31848]_ ;
  assign \new_[31853]_  = ~A200 & ~A199;
  assign \new_[31854]_  = A166 & \new_[31853]_ ;
  assign \new_[31855]_  = \new_[31854]_  & \new_[31849]_ ;
  assign \new_[31859]_  = A267 & A266;
  assign \new_[31860]_  = ~A265 & \new_[31859]_ ;
  assign \new_[31864]_  = A299 & A298;
  assign \new_[31865]_  = A268 & \new_[31864]_ ;
  assign \new_[31866]_  = \new_[31865]_  & \new_[31860]_ ;
  assign \new_[31870]_  = ~A167 & A168;
  assign \new_[31871]_  = A170 & \new_[31870]_ ;
  assign \new_[31875]_  = ~A200 & ~A199;
  assign \new_[31876]_  = A166 & \new_[31875]_ ;
  assign \new_[31877]_  = \new_[31876]_  & \new_[31871]_ ;
  assign \new_[31881]_  = A267 & A266;
  assign \new_[31882]_  = ~A265 & \new_[31881]_ ;
  assign \new_[31886]_  = ~A299 & ~A298;
  assign \new_[31887]_  = A268 & \new_[31886]_ ;
  assign \new_[31888]_  = \new_[31887]_  & \new_[31882]_ ;
  assign \new_[31892]_  = ~A167 & A168;
  assign \new_[31893]_  = A170 & \new_[31892]_ ;
  assign \new_[31897]_  = ~A200 & ~A199;
  assign \new_[31898]_  = A166 & \new_[31897]_ ;
  assign \new_[31899]_  = \new_[31898]_  & \new_[31893]_ ;
  assign \new_[31903]_  = A267 & A266;
  assign \new_[31904]_  = ~A265 & \new_[31903]_ ;
  assign \new_[31908]_  = A301 & ~A300;
  assign \new_[31909]_  = ~A269 & \new_[31908]_ ;
  assign \new_[31910]_  = \new_[31909]_  & \new_[31904]_ ;
  assign \new_[31914]_  = ~A167 & A168;
  assign \new_[31915]_  = A170 & \new_[31914]_ ;
  assign \new_[31919]_  = ~A200 & ~A199;
  assign \new_[31920]_  = A166 & \new_[31919]_ ;
  assign \new_[31921]_  = \new_[31920]_  & \new_[31915]_ ;
  assign \new_[31925]_  = A267 & A266;
  assign \new_[31926]_  = ~A265 & \new_[31925]_ ;
  assign \new_[31930]_  = ~A302 & ~A300;
  assign \new_[31931]_  = ~A269 & \new_[31930]_ ;
  assign \new_[31932]_  = \new_[31931]_  & \new_[31926]_ ;
  assign \new_[31936]_  = ~A167 & A168;
  assign \new_[31937]_  = A170 & \new_[31936]_ ;
  assign \new_[31941]_  = ~A200 & ~A199;
  assign \new_[31942]_  = A166 & \new_[31941]_ ;
  assign \new_[31943]_  = \new_[31942]_  & \new_[31937]_ ;
  assign \new_[31947]_  = A267 & A266;
  assign \new_[31948]_  = ~A265 & \new_[31947]_ ;
  assign \new_[31952]_  = A299 & A298;
  assign \new_[31953]_  = ~A269 & \new_[31952]_ ;
  assign \new_[31954]_  = \new_[31953]_  & \new_[31948]_ ;
  assign \new_[31958]_  = ~A167 & A168;
  assign \new_[31959]_  = A170 & \new_[31958]_ ;
  assign \new_[31963]_  = ~A200 & ~A199;
  assign \new_[31964]_  = A166 & \new_[31963]_ ;
  assign \new_[31965]_  = \new_[31964]_  & \new_[31959]_ ;
  assign \new_[31969]_  = A267 & A266;
  assign \new_[31970]_  = ~A265 & \new_[31969]_ ;
  assign \new_[31974]_  = ~A299 & ~A298;
  assign \new_[31975]_  = ~A269 & \new_[31974]_ ;
  assign \new_[31976]_  = \new_[31975]_  & \new_[31970]_ ;
  assign \new_[31980]_  = ~A167 & A168;
  assign \new_[31981]_  = A170 & \new_[31980]_ ;
  assign \new_[31985]_  = ~A200 & ~A199;
  assign \new_[31986]_  = A166 & \new_[31985]_ ;
  assign \new_[31987]_  = \new_[31986]_  & \new_[31981]_ ;
  assign \new_[31991]_  = A267 & ~A266;
  assign \new_[31992]_  = A265 & \new_[31991]_ ;
  assign \new_[31996]_  = A301 & ~A300;
  assign \new_[31997]_  = A268 & \new_[31996]_ ;
  assign \new_[31998]_  = \new_[31997]_  & \new_[31992]_ ;
  assign \new_[32002]_  = ~A167 & A168;
  assign \new_[32003]_  = A170 & \new_[32002]_ ;
  assign \new_[32007]_  = ~A200 & ~A199;
  assign \new_[32008]_  = A166 & \new_[32007]_ ;
  assign \new_[32009]_  = \new_[32008]_  & \new_[32003]_ ;
  assign \new_[32013]_  = A267 & ~A266;
  assign \new_[32014]_  = A265 & \new_[32013]_ ;
  assign \new_[32018]_  = ~A302 & ~A300;
  assign \new_[32019]_  = A268 & \new_[32018]_ ;
  assign \new_[32020]_  = \new_[32019]_  & \new_[32014]_ ;
  assign \new_[32024]_  = ~A167 & A168;
  assign \new_[32025]_  = A170 & \new_[32024]_ ;
  assign \new_[32029]_  = ~A200 & ~A199;
  assign \new_[32030]_  = A166 & \new_[32029]_ ;
  assign \new_[32031]_  = \new_[32030]_  & \new_[32025]_ ;
  assign \new_[32035]_  = A267 & ~A266;
  assign \new_[32036]_  = A265 & \new_[32035]_ ;
  assign \new_[32040]_  = A299 & A298;
  assign \new_[32041]_  = A268 & \new_[32040]_ ;
  assign \new_[32042]_  = \new_[32041]_  & \new_[32036]_ ;
  assign \new_[32046]_  = ~A167 & A168;
  assign \new_[32047]_  = A170 & \new_[32046]_ ;
  assign \new_[32051]_  = ~A200 & ~A199;
  assign \new_[32052]_  = A166 & \new_[32051]_ ;
  assign \new_[32053]_  = \new_[32052]_  & \new_[32047]_ ;
  assign \new_[32057]_  = A267 & ~A266;
  assign \new_[32058]_  = A265 & \new_[32057]_ ;
  assign \new_[32062]_  = ~A299 & ~A298;
  assign \new_[32063]_  = A268 & \new_[32062]_ ;
  assign \new_[32064]_  = \new_[32063]_  & \new_[32058]_ ;
  assign \new_[32068]_  = ~A167 & A168;
  assign \new_[32069]_  = A170 & \new_[32068]_ ;
  assign \new_[32073]_  = ~A200 & ~A199;
  assign \new_[32074]_  = A166 & \new_[32073]_ ;
  assign \new_[32075]_  = \new_[32074]_  & \new_[32069]_ ;
  assign \new_[32079]_  = A267 & ~A266;
  assign \new_[32080]_  = A265 & \new_[32079]_ ;
  assign \new_[32084]_  = A301 & ~A300;
  assign \new_[32085]_  = ~A269 & \new_[32084]_ ;
  assign \new_[32086]_  = \new_[32085]_  & \new_[32080]_ ;
  assign \new_[32090]_  = ~A167 & A168;
  assign \new_[32091]_  = A170 & \new_[32090]_ ;
  assign \new_[32095]_  = ~A200 & ~A199;
  assign \new_[32096]_  = A166 & \new_[32095]_ ;
  assign \new_[32097]_  = \new_[32096]_  & \new_[32091]_ ;
  assign \new_[32101]_  = A267 & ~A266;
  assign \new_[32102]_  = A265 & \new_[32101]_ ;
  assign \new_[32106]_  = ~A302 & ~A300;
  assign \new_[32107]_  = ~A269 & \new_[32106]_ ;
  assign \new_[32108]_  = \new_[32107]_  & \new_[32102]_ ;
  assign \new_[32112]_  = ~A167 & A168;
  assign \new_[32113]_  = A170 & \new_[32112]_ ;
  assign \new_[32117]_  = ~A200 & ~A199;
  assign \new_[32118]_  = A166 & \new_[32117]_ ;
  assign \new_[32119]_  = \new_[32118]_  & \new_[32113]_ ;
  assign \new_[32123]_  = A267 & ~A266;
  assign \new_[32124]_  = A265 & \new_[32123]_ ;
  assign \new_[32128]_  = A299 & A298;
  assign \new_[32129]_  = ~A269 & \new_[32128]_ ;
  assign \new_[32130]_  = \new_[32129]_  & \new_[32124]_ ;
  assign \new_[32134]_  = ~A167 & A168;
  assign \new_[32135]_  = A170 & \new_[32134]_ ;
  assign \new_[32139]_  = ~A200 & ~A199;
  assign \new_[32140]_  = A166 & \new_[32139]_ ;
  assign \new_[32141]_  = \new_[32140]_  & \new_[32135]_ ;
  assign \new_[32145]_  = A267 & ~A266;
  assign \new_[32146]_  = A265 & \new_[32145]_ ;
  assign \new_[32150]_  = ~A299 & ~A298;
  assign \new_[32151]_  = ~A269 & \new_[32150]_ ;
  assign \new_[32152]_  = \new_[32151]_  & \new_[32146]_ ;
  assign \new_[32156]_  = ~A167 & A168;
  assign \new_[32157]_  = A170 & \new_[32156]_ ;
  assign \new_[32161]_  = ~A200 & ~A199;
  assign \new_[32162]_  = A166 & \new_[32161]_ ;
  assign \new_[32163]_  = \new_[32162]_  & \new_[32157]_ ;
  assign \new_[32167]_  = A298 & ~A266;
  assign \new_[32168]_  = ~A265 & \new_[32167]_ ;
  assign \new_[32172]_  = A301 & A300;
  assign \new_[32173]_  = ~A299 & \new_[32172]_ ;
  assign \new_[32174]_  = \new_[32173]_  & \new_[32168]_ ;
  assign \new_[32178]_  = ~A167 & A168;
  assign \new_[32179]_  = A170 & \new_[32178]_ ;
  assign \new_[32183]_  = ~A200 & ~A199;
  assign \new_[32184]_  = A166 & \new_[32183]_ ;
  assign \new_[32185]_  = \new_[32184]_  & \new_[32179]_ ;
  assign \new_[32189]_  = A298 & ~A266;
  assign \new_[32190]_  = ~A265 & \new_[32189]_ ;
  assign \new_[32194]_  = ~A302 & A300;
  assign \new_[32195]_  = ~A299 & \new_[32194]_ ;
  assign \new_[32196]_  = \new_[32195]_  & \new_[32190]_ ;
  assign \new_[32200]_  = ~A167 & A168;
  assign \new_[32201]_  = A170 & \new_[32200]_ ;
  assign \new_[32205]_  = ~A200 & ~A199;
  assign \new_[32206]_  = A166 & \new_[32205]_ ;
  assign \new_[32207]_  = \new_[32206]_  & \new_[32201]_ ;
  assign \new_[32211]_  = ~A298 & ~A266;
  assign \new_[32212]_  = ~A265 & \new_[32211]_ ;
  assign \new_[32216]_  = A301 & A300;
  assign \new_[32217]_  = A299 & \new_[32216]_ ;
  assign \new_[32218]_  = \new_[32217]_  & \new_[32212]_ ;
  assign \new_[32222]_  = ~A167 & A168;
  assign \new_[32223]_  = A170 & \new_[32222]_ ;
  assign \new_[32227]_  = ~A200 & ~A199;
  assign \new_[32228]_  = A166 & \new_[32227]_ ;
  assign \new_[32229]_  = \new_[32228]_  & \new_[32223]_ ;
  assign \new_[32233]_  = ~A298 & ~A266;
  assign \new_[32234]_  = ~A265 & \new_[32233]_ ;
  assign \new_[32238]_  = ~A302 & A300;
  assign \new_[32239]_  = A299 & \new_[32238]_ ;
  assign \new_[32240]_  = \new_[32239]_  & \new_[32234]_ ;
  assign \new_[32244]_  = ~A232 & ~A168;
  assign \new_[32245]_  = A170 & \new_[32244]_ ;
  assign \new_[32249]_  = ~A235 & ~A234;
  assign \new_[32250]_  = A233 & \new_[32249]_ ;
  assign \new_[32251]_  = \new_[32250]_  & \new_[32245]_ ;
  assign \new_[32255]_  = A266 & ~A265;
  assign \new_[32256]_  = A236 & \new_[32255]_ ;
  assign \new_[32260]_  = A269 & ~A268;
  assign \new_[32261]_  = ~A267 & \new_[32260]_ ;
  assign \new_[32262]_  = \new_[32261]_  & \new_[32256]_ ;
  assign \new_[32266]_  = ~A232 & ~A168;
  assign \new_[32267]_  = A170 & \new_[32266]_ ;
  assign \new_[32271]_  = ~A235 & ~A234;
  assign \new_[32272]_  = A233 & \new_[32271]_ ;
  assign \new_[32273]_  = \new_[32272]_  & \new_[32267]_ ;
  assign \new_[32277]_  = ~A266 & A265;
  assign \new_[32278]_  = A236 & \new_[32277]_ ;
  assign \new_[32282]_  = A269 & ~A268;
  assign \new_[32283]_  = ~A267 & \new_[32282]_ ;
  assign \new_[32284]_  = \new_[32283]_  & \new_[32278]_ ;
  assign \new_[32288]_  = A232 & ~A168;
  assign \new_[32289]_  = A170 & \new_[32288]_ ;
  assign \new_[32293]_  = ~A235 & ~A234;
  assign \new_[32294]_  = ~A233 & \new_[32293]_ ;
  assign \new_[32295]_  = \new_[32294]_  & \new_[32289]_ ;
  assign \new_[32299]_  = A266 & ~A265;
  assign \new_[32300]_  = A236 & \new_[32299]_ ;
  assign \new_[32304]_  = A269 & ~A268;
  assign \new_[32305]_  = ~A267 & \new_[32304]_ ;
  assign \new_[32306]_  = \new_[32305]_  & \new_[32300]_ ;
  assign \new_[32310]_  = A232 & ~A168;
  assign \new_[32311]_  = A170 & \new_[32310]_ ;
  assign \new_[32315]_  = ~A235 & ~A234;
  assign \new_[32316]_  = ~A233 & \new_[32315]_ ;
  assign \new_[32317]_  = \new_[32316]_  & \new_[32311]_ ;
  assign \new_[32321]_  = ~A266 & A265;
  assign \new_[32322]_  = A236 & \new_[32321]_ ;
  assign \new_[32326]_  = A269 & ~A268;
  assign \new_[32327]_  = ~A267 & \new_[32326]_ ;
  assign \new_[32328]_  = \new_[32327]_  & \new_[32322]_ ;
  assign \new_[32332]_  = ~A199 & ~A168;
  assign \new_[32333]_  = A170 & \new_[32332]_ ;
  assign \new_[32337]_  = A202 & A201;
  assign \new_[32338]_  = A200 & \new_[32337]_ ;
  assign \new_[32339]_  = \new_[32338]_  & \new_[32333]_ ;
  assign \new_[32343]_  = A269 & ~A268;
  assign \new_[32344]_  = A267 & \new_[32343]_ ;
  assign \new_[32348]_  = A302 & ~A301;
  assign \new_[32349]_  = A300 & \new_[32348]_ ;
  assign \new_[32350]_  = \new_[32349]_  & \new_[32344]_ ;
  assign \new_[32354]_  = ~A199 & ~A168;
  assign \new_[32355]_  = A170 & \new_[32354]_ ;
  assign \new_[32359]_  = ~A203 & A201;
  assign \new_[32360]_  = A200 & \new_[32359]_ ;
  assign \new_[32361]_  = \new_[32360]_  & \new_[32355]_ ;
  assign \new_[32365]_  = A269 & ~A268;
  assign \new_[32366]_  = A267 & \new_[32365]_ ;
  assign \new_[32370]_  = A302 & ~A301;
  assign \new_[32371]_  = A300 & \new_[32370]_ ;
  assign \new_[32372]_  = \new_[32371]_  & \new_[32366]_ ;
  assign \new_[32376]_  = ~A199 & ~A168;
  assign \new_[32377]_  = A170 & \new_[32376]_ ;
  assign \new_[32381]_  = ~A202 & ~A201;
  assign \new_[32382]_  = A200 & \new_[32381]_ ;
  assign \new_[32383]_  = \new_[32382]_  & \new_[32377]_ ;
  assign \new_[32387]_  = ~A268 & A267;
  assign \new_[32388]_  = A203 & \new_[32387]_ ;
  assign \new_[32392]_  = A301 & ~A300;
  assign \new_[32393]_  = A269 & \new_[32392]_ ;
  assign \new_[32394]_  = \new_[32393]_  & \new_[32388]_ ;
  assign \new_[32398]_  = ~A199 & ~A168;
  assign \new_[32399]_  = A170 & \new_[32398]_ ;
  assign \new_[32403]_  = ~A202 & ~A201;
  assign \new_[32404]_  = A200 & \new_[32403]_ ;
  assign \new_[32405]_  = \new_[32404]_  & \new_[32399]_ ;
  assign \new_[32409]_  = ~A268 & A267;
  assign \new_[32410]_  = A203 & \new_[32409]_ ;
  assign \new_[32414]_  = ~A302 & ~A300;
  assign \new_[32415]_  = A269 & \new_[32414]_ ;
  assign \new_[32416]_  = \new_[32415]_  & \new_[32410]_ ;
  assign \new_[32420]_  = ~A199 & ~A168;
  assign \new_[32421]_  = A170 & \new_[32420]_ ;
  assign \new_[32425]_  = ~A202 & ~A201;
  assign \new_[32426]_  = A200 & \new_[32425]_ ;
  assign \new_[32427]_  = \new_[32426]_  & \new_[32421]_ ;
  assign \new_[32431]_  = ~A268 & A267;
  assign \new_[32432]_  = A203 & \new_[32431]_ ;
  assign \new_[32436]_  = A299 & A298;
  assign \new_[32437]_  = A269 & \new_[32436]_ ;
  assign \new_[32438]_  = \new_[32437]_  & \new_[32432]_ ;
  assign \new_[32442]_  = ~A199 & ~A168;
  assign \new_[32443]_  = A170 & \new_[32442]_ ;
  assign \new_[32447]_  = ~A202 & ~A201;
  assign \new_[32448]_  = A200 & \new_[32447]_ ;
  assign \new_[32449]_  = \new_[32448]_  & \new_[32443]_ ;
  assign \new_[32453]_  = ~A268 & A267;
  assign \new_[32454]_  = A203 & \new_[32453]_ ;
  assign \new_[32458]_  = ~A299 & ~A298;
  assign \new_[32459]_  = A269 & \new_[32458]_ ;
  assign \new_[32460]_  = \new_[32459]_  & \new_[32454]_ ;
  assign \new_[32464]_  = ~A199 & ~A168;
  assign \new_[32465]_  = A170 & \new_[32464]_ ;
  assign \new_[32469]_  = ~A202 & ~A201;
  assign \new_[32470]_  = A200 & \new_[32469]_ ;
  assign \new_[32471]_  = \new_[32470]_  & \new_[32465]_ ;
  assign \new_[32475]_  = A268 & ~A267;
  assign \new_[32476]_  = A203 & \new_[32475]_ ;
  assign \new_[32480]_  = A302 & ~A301;
  assign \new_[32481]_  = A300 & \new_[32480]_ ;
  assign \new_[32482]_  = \new_[32481]_  & \new_[32476]_ ;
  assign \new_[32486]_  = ~A199 & ~A168;
  assign \new_[32487]_  = A170 & \new_[32486]_ ;
  assign \new_[32491]_  = ~A202 & ~A201;
  assign \new_[32492]_  = A200 & \new_[32491]_ ;
  assign \new_[32493]_  = \new_[32492]_  & \new_[32487]_ ;
  assign \new_[32497]_  = ~A269 & ~A267;
  assign \new_[32498]_  = A203 & \new_[32497]_ ;
  assign \new_[32502]_  = A302 & ~A301;
  assign \new_[32503]_  = A300 & \new_[32502]_ ;
  assign \new_[32504]_  = \new_[32503]_  & \new_[32498]_ ;
  assign \new_[32508]_  = ~A199 & ~A168;
  assign \new_[32509]_  = A170 & \new_[32508]_ ;
  assign \new_[32513]_  = ~A202 & ~A201;
  assign \new_[32514]_  = A200 & \new_[32513]_ ;
  assign \new_[32515]_  = \new_[32514]_  & \new_[32509]_ ;
  assign \new_[32519]_  = A266 & A265;
  assign \new_[32520]_  = A203 & \new_[32519]_ ;
  assign \new_[32524]_  = A302 & ~A301;
  assign \new_[32525]_  = A300 & \new_[32524]_ ;
  assign \new_[32526]_  = \new_[32525]_  & \new_[32520]_ ;
  assign \new_[32530]_  = ~A199 & ~A168;
  assign \new_[32531]_  = A170 & \new_[32530]_ ;
  assign \new_[32535]_  = ~A202 & ~A201;
  assign \new_[32536]_  = A200 & \new_[32535]_ ;
  assign \new_[32537]_  = \new_[32536]_  & \new_[32531]_ ;
  assign \new_[32541]_  = ~A266 & ~A265;
  assign \new_[32542]_  = A203 & \new_[32541]_ ;
  assign \new_[32546]_  = A302 & ~A301;
  assign \new_[32547]_  = A300 & \new_[32546]_ ;
  assign \new_[32548]_  = \new_[32547]_  & \new_[32542]_ ;
  assign \new_[32552]_  = A199 & ~A168;
  assign \new_[32553]_  = A170 & \new_[32552]_ ;
  assign \new_[32557]_  = A202 & A201;
  assign \new_[32558]_  = ~A200 & \new_[32557]_ ;
  assign \new_[32559]_  = \new_[32558]_  & \new_[32553]_ ;
  assign \new_[32563]_  = A269 & ~A268;
  assign \new_[32564]_  = A267 & \new_[32563]_ ;
  assign \new_[32568]_  = A302 & ~A301;
  assign \new_[32569]_  = A300 & \new_[32568]_ ;
  assign \new_[32570]_  = \new_[32569]_  & \new_[32564]_ ;
  assign \new_[32574]_  = A199 & ~A168;
  assign \new_[32575]_  = A170 & \new_[32574]_ ;
  assign \new_[32579]_  = ~A203 & A201;
  assign \new_[32580]_  = ~A200 & \new_[32579]_ ;
  assign \new_[32581]_  = \new_[32580]_  & \new_[32575]_ ;
  assign \new_[32585]_  = A269 & ~A268;
  assign \new_[32586]_  = A267 & \new_[32585]_ ;
  assign \new_[32590]_  = A302 & ~A301;
  assign \new_[32591]_  = A300 & \new_[32590]_ ;
  assign \new_[32592]_  = \new_[32591]_  & \new_[32586]_ ;
  assign \new_[32596]_  = A199 & ~A168;
  assign \new_[32597]_  = A170 & \new_[32596]_ ;
  assign \new_[32601]_  = ~A202 & ~A201;
  assign \new_[32602]_  = ~A200 & \new_[32601]_ ;
  assign \new_[32603]_  = \new_[32602]_  & \new_[32597]_ ;
  assign \new_[32607]_  = ~A268 & A267;
  assign \new_[32608]_  = A203 & \new_[32607]_ ;
  assign \new_[32612]_  = A301 & ~A300;
  assign \new_[32613]_  = A269 & \new_[32612]_ ;
  assign \new_[32614]_  = \new_[32613]_  & \new_[32608]_ ;
  assign \new_[32618]_  = A199 & ~A168;
  assign \new_[32619]_  = A170 & \new_[32618]_ ;
  assign \new_[32623]_  = ~A202 & ~A201;
  assign \new_[32624]_  = ~A200 & \new_[32623]_ ;
  assign \new_[32625]_  = \new_[32624]_  & \new_[32619]_ ;
  assign \new_[32629]_  = ~A268 & A267;
  assign \new_[32630]_  = A203 & \new_[32629]_ ;
  assign \new_[32634]_  = ~A302 & ~A300;
  assign \new_[32635]_  = A269 & \new_[32634]_ ;
  assign \new_[32636]_  = \new_[32635]_  & \new_[32630]_ ;
  assign \new_[32640]_  = A199 & ~A168;
  assign \new_[32641]_  = A170 & \new_[32640]_ ;
  assign \new_[32645]_  = ~A202 & ~A201;
  assign \new_[32646]_  = ~A200 & \new_[32645]_ ;
  assign \new_[32647]_  = \new_[32646]_  & \new_[32641]_ ;
  assign \new_[32651]_  = ~A268 & A267;
  assign \new_[32652]_  = A203 & \new_[32651]_ ;
  assign \new_[32656]_  = A299 & A298;
  assign \new_[32657]_  = A269 & \new_[32656]_ ;
  assign \new_[32658]_  = \new_[32657]_  & \new_[32652]_ ;
  assign \new_[32662]_  = A199 & ~A168;
  assign \new_[32663]_  = A170 & \new_[32662]_ ;
  assign \new_[32667]_  = ~A202 & ~A201;
  assign \new_[32668]_  = ~A200 & \new_[32667]_ ;
  assign \new_[32669]_  = \new_[32668]_  & \new_[32663]_ ;
  assign \new_[32673]_  = ~A268 & A267;
  assign \new_[32674]_  = A203 & \new_[32673]_ ;
  assign \new_[32678]_  = ~A299 & ~A298;
  assign \new_[32679]_  = A269 & \new_[32678]_ ;
  assign \new_[32680]_  = \new_[32679]_  & \new_[32674]_ ;
  assign \new_[32684]_  = A199 & ~A168;
  assign \new_[32685]_  = A170 & \new_[32684]_ ;
  assign \new_[32689]_  = ~A202 & ~A201;
  assign \new_[32690]_  = ~A200 & \new_[32689]_ ;
  assign \new_[32691]_  = \new_[32690]_  & \new_[32685]_ ;
  assign \new_[32695]_  = A268 & ~A267;
  assign \new_[32696]_  = A203 & \new_[32695]_ ;
  assign \new_[32700]_  = A302 & ~A301;
  assign \new_[32701]_  = A300 & \new_[32700]_ ;
  assign \new_[32702]_  = \new_[32701]_  & \new_[32696]_ ;
  assign \new_[32706]_  = A199 & ~A168;
  assign \new_[32707]_  = A170 & \new_[32706]_ ;
  assign \new_[32711]_  = ~A202 & ~A201;
  assign \new_[32712]_  = ~A200 & \new_[32711]_ ;
  assign \new_[32713]_  = \new_[32712]_  & \new_[32707]_ ;
  assign \new_[32717]_  = ~A269 & ~A267;
  assign \new_[32718]_  = A203 & \new_[32717]_ ;
  assign \new_[32722]_  = A302 & ~A301;
  assign \new_[32723]_  = A300 & \new_[32722]_ ;
  assign \new_[32724]_  = \new_[32723]_  & \new_[32718]_ ;
  assign \new_[32728]_  = A199 & ~A168;
  assign \new_[32729]_  = A170 & \new_[32728]_ ;
  assign \new_[32733]_  = ~A202 & ~A201;
  assign \new_[32734]_  = ~A200 & \new_[32733]_ ;
  assign \new_[32735]_  = \new_[32734]_  & \new_[32729]_ ;
  assign \new_[32739]_  = A266 & A265;
  assign \new_[32740]_  = A203 & \new_[32739]_ ;
  assign \new_[32744]_  = A302 & ~A301;
  assign \new_[32745]_  = A300 & \new_[32744]_ ;
  assign \new_[32746]_  = \new_[32745]_  & \new_[32740]_ ;
  assign \new_[32750]_  = A199 & ~A168;
  assign \new_[32751]_  = A170 & \new_[32750]_ ;
  assign \new_[32755]_  = ~A202 & ~A201;
  assign \new_[32756]_  = ~A200 & \new_[32755]_ ;
  assign \new_[32757]_  = \new_[32756]_  & \new_[32751]_ ;
  assign \new_[32761]_  = ~A266 & ~A265;
  assign \new_[32762]_  = A203 & \new_[32761]_ ;
  assign \new_[32766]_  = A302 & ~A301;
  assign \new_[32767]_  = A300 & \new_[32766]_ ;
  assign \new_[32768]_  = \new_[32767]_  & \new_[32762]_ ;
  assign \new_[32772]_  = A167 & A168;
  assign \new_[32773]_  = A169 & \new_[32772]_ ;
  assign \new_[32777]_  = A202 & ~A201;
  assign \new_[32778]_  = ~A166 & \new_[32777]_ ;
  assign \new_[32779]_  = \new_[32778]_  & \new_[32773]_ ;
  assign \new_[32783]_  = A298 & A268;
  assign \new_[32784]_  = ~A267 & \new_[32783]_ ;
  assign \new_[32788]_  = A301 & A300;
  assign \new_[32789]_  = ~A299 & \new_[32788]_ ;
  assign \new_[32790]_  = \new_[32789]_  & \new_[32784]_ ;
  assign \new_[32794]_  = A167 & A168;
  assign \new_[32795]_  = A169 & \new_[32794]_ ;
  assign \new_[32799]_  = A202 & ~A201;
  assign \new_[32800]_  = ~A166 & \new_[32799]_ ;
  assign \new_[32801]_  = \new_[32800]_  & \new_[32795]_ ;
  assign \new_[32805]_  = A298 & A268;
  assign \new_[32806]_  = ~A267 & \new_[32805]_ ;
  assign \new_[32810]_  = ~A302 & A300;
  assign \new_[32811]_  = ~A299 & \new_[32810]_ ;
  assign \new_[32812]_  = \new_[32811]_  & \new_[32806]_ ;
  assign \new_[32816]_  = A167 & A168;
  assign \new_[32817]_  = A169 & \new_[32816]_ ;
  assign \new_[32821]_  = A202 & ~A201;
  assign \new_[32822]_  = ~A166 & \new_[32821]_ ;
  assign \new_[32823]_  = \new_[32822]_  & \new_[32817]_ ;
  assign \new_[32827]_  = ~A298 & A268;
  assign \new_[32828]_  = ~A267 & \new_[32827]_ ;
  assign \new_[32832]_  = A301 & A300;
  assign \new_[32833]_  = A299 & \new_[32832]_ ;
  assign \new_[32834]_  = \new_[32833]_  & \new_[32828]_ ;
  assign \new_[32838]_  = A167 & A168;
  assign \new_[32839]_  = A169 & \new_[32838]_ ;
  assign \new_[32843]_  = A202 & ~A201;
  assign \new_[32844]_  = ~A166 & \new_[32843]_ ;
  assign \new_[32845]_  = \new_[32844]_  & \new_[32839]_ ;
  assign \new_[32849]_  = ~A298 & A268;
  assign \new_[32850]_  = ~A267 & \new_[32849]_ ;
  assign \new_[32854]_  = ~A302 & A300;
  assign \new_[32855]_  = A299 & \new_[32854]_ ;
  assign \new_[32856]_  = \new_[32855]_  & \new_[32850]_ ;
  assign \new_[32860]_  = A167 & A168;
  assign \new_[32861]_  = A169 & \new_[32860]_ ;
  assign \new_[32865]_  = A202 & ~A201;
  assign \new_[32866]_  = ~A166 & \new_[32865]_ ;
  assign \new_[32867]_  = \new_[32866]_  & \new_[32861]_ ;
  assign \new_[32871]_  = A298 & ~A269;
  assign \new_[32872]_  = ~A267 & \new_[32871]_ ;
  assign \new_[32876]_  = A301 & A300;
  assign \new_[32877]_  = ~A299 & \new_[32876]_ ;
  assign \new_[32878]_  = \new_[32877]_  & \new_[32872]_ ;
  assign \new_[32882]_  = A167 & A168;
  assign \new_[32883]_  = A169 & \new_[32882]_ ;
  assign \new_[32887]_  = A202 & ~A201;
  assign \new_[32888]_  = ~A166 & \new_[32887]_ ;
  assign \new_[32889]_  = \new_[32888]_  & \new_[32883]_ ;
  assign \new_[32893]_  = A298 & ~A269;
  assign \new_[32894]_  = ~A267 & \new_[32893]_ ;
  assign \new_[32898]_  = ~A302 & A300;
  assign \new_[32899]_  = ~A299 & \new_[32898]_ ;
  assign \new_[32900]_  = \new_[32899]_  & \new_[32894]_ ;
  assign \new_[32904]_  = A167 & A168;
  assign \new_[32905]_  = A169 & \new_[32904]_ ;
  assign \new_[32909]_  = A202 & ~A201;
  assign \new_[32910]_  = ~A166 & \new_[32909]_ ;
  assign \new_[32911]_  = \new_[32910]_  & \new_[32905]_ ;
  assign \new_[32915]_  = ~A298 & ~A269;
  assign \new_[32916]_  = ~A267 & \new_[32915]_ ;
  assign \new_[32920]_  = A301 & A300;
  assign \new_[32921]_  = A299 & \new_[32920]_ ;
  assign \new_[32922]_  = \new_[32921]_  & \new_[32916]_ ;
  assign \new_[32926]_  = A167 & A168;
  assign \new_[32927]_  = A169 & \new_[32926]_ ;
  assign \new_[32931]_  = A202 & ~A201;
  assign \new_[32932]_  = ~A166 & \new_[32931]_ ;
  assign \new_[32933]_  = \new_[32932]_  & \new_[32927]_ ;
  assign \new_[32937]_  = ~A298 & ~A269;
  assign \new_[32938]_  = ~A267 & \new_[32937]_ ;
  assign \new_[32942]_  = ~A302 & A300;
  assign \new_[32943]_  = A299 & \new_[32942]_ ;
  assign \new_[32944]_  = \new_[32943]_  & \new_[32938]_ ;
  assign \new_[32948]_  = A167 & A168;
  assign \new_[32949]_  = A169 & \new_[32948]_ ;
  assign \new_[32953]_  = A202 & ~A201;
  assign \new_[32954]_  = ~A166 & \new_[32953]_ ;
  assign \new_[32955]_  = \new_[32954]_  & \new_[32949]_ ;
  assign \new_[32959]_  = A298 & A266;
  assign \new_[32960]_  = A265 & \new_[32959]_ ;
  assign \new_[32964]_  = A301 & A300;
  assign \new_[32965]_  = ~A299 & \new_[32964]_ ;
  assign \new_[32966]_  = \new_[32965]_  & \new_[32960]_ ;
  assign \new_[32970]_  = A167 & A168;
  assign \new_[32971]_  = A169 & \new_[32970]_ ;
  assign \new_[32975]_  = A202 & ~A201;
  assign \new_[32976]_  = ~A166 & \new_[32975]_ ;
  assign \new_[32977]_  = \new_[32976]_  & \new_[32971]_ ;
  assign \new_[32981]_  = A298 & A266;
  assign \new_[32982]_  = A265 & \new_[32981]_ ;
  assign \new_[32986]_  = ~A302 & A300;
  assign \new_[32987]_  = ~A299 & \new_[32986]_ ;
  assign \new_[32988]_  = \new_[32987]_  & \new_[32982]_ ;
  assign \new_[32992]_  = A167 & A168;
  assign \new_[32993]_  = A169 & \new_[32992]_ ;
  assign \new_[32997]_  = A202 & ~A201;
  assign \new_[32998]_  = ~A166 & \new_[32997]_ ;
  assign \new_[32999]_  = \new_[32998]_  & \new_[32993]_ ;
  assign \new_[33003]_  = ~A298 & A266;
  assign \new_[33004]_  = A265 & \new_[33003]_ ;
  assign \new_[33008]_  = A301 & A300;
  assign \new_[33009]_  = A299 & \new_[33008]_ ;
  assign \new_[33010]_  = \new_[33009]_  & \new_[33004]_ ;
  assign \new_[33014]_  = A167 & A168;
  assign \new_[33015]_  = A169 & \new_[33014]_ ;
  assign \new_[33019]_  = A202 & ~A201;
  assign \new_[33020]_  = ~A166 & \new_[33019]_ ;
  assign \new_[33021]_  = \new_[33020]_  & \new_[33015]_ ;
  assign \new_[33025]_  = ~A298 & A266;
  assign \new_[33026]_  = A265 & \new_[33025]_ ;
  assign \new_[33030]_  = ~A302 & A300;
  assign \new_[33031]_  = A299 & \new_[33030]_ ;
  assign \new_[33032]_  = \new_[33031]_  & \new_[33026]_ ;
  assign \new_[33036]_  = A167 & A168;
  assign \new_[33037]_  = A169 & \new_[33036]_ ;
  assign \new_[33041]_  = A202 & ~A201;
  assign \new_[33042]_  = ~A166 & \new_[33041]_ ;
  assign \new_[33043]_  = \new_[33042]_  & \new_[33037]_ ;
  assign \new_[33047]_  = A267 & A266;
  assign \new_[33048]_  = ~A265 & \new_[33047]_ ;
  assign \new_[33052]_  = A301 & ~A300;
  assign \new_[33053]_  = A268 & \new_[33052]_ ;
  assign \new_[33054]_  = \new_[33053]_  & \new_[33048]_ ;
  assign \new_[33058]_  = A167 & A168;
  assign \new_[33059]_  = A169 & \new_[33058]_ ;
  assign \new_[33063]_  = A202 & ~A201;
  assign \new_[33064]_  = ~A166 & \new_[33063]_ ;
  assign \new_[33065]_  = \new_[33064]_  & \new_[33059]_ ;
  assign \new_[33069]_  = A267 & A266;
  assign \new_[33070]_  = ~A265 & \new_[33069]_ ;
  assign \new_[33074]_  = ~A302 & ~A300;
  assign \new_[33075]_  = A268 & \new_[33074]_ ;
  assign \new_[33076]_  = \new_[33075]_  & \new_[33070]_ ;
  assign \new_[33080]_  = A167 & A168;
  assign \new_[33081]_  = A169 & \new_[33080]_ ;
  assign \new_[33085]_  = A202 & ~A201;
  assign \new_[33086]_  = ~A166 & \new_[33085]_ ;
  assign \new_[33087]_  = \new_[33086]_  & \new_[33081]_ ;
  assign \new_[33091]_  = A267 & A266;
  assign \new_[33092]_  = ~A265 & \new_[33091]_ ;
  assign \new_[33096]_  = A299 & A298;
  assign \new_[33097]_  = A268 & \new_[33096]_ ;
  assign \new_[33098]_  = \new_[33097]_  & \new_[33092]_ ;
  assign \new_[33102]_  = A167 & A168;
  assign \new_[33103]_  = A169 & \new_[33102]_ ;
  assign \new_[33107]_  = A202 & ~A201;
  assign \new_[33108]_  = ~A166 & \new_[33107]_ ;
  assign \new_[33109]_  = \new_[33108]_  & \new_[33103]_ ;
  assign \new_[33113]_  = A267 & A266;
  assign \new_[33114]_  = ~A265 & \new_[33113]_ ;
  assign \new_[33118]_  = ~A299 & ~A298;
  assign \new_[33119]_  = A268 & \new_[33118]_ ;
  assign \new_[33120]_  = \new_[33119]_  & \new_[33114]_ ;
  assign \new_[33124]_  = A167 & A168;
  assign \new_[33125]_  = A169 & \new_[33124]_ ;
  assign \new_[33129]_  = A202 & ~A201;
  assign \new_[33130]_  = ~A166 & \new_[33129]_ ;
  assign \new_[33131]_  = \new_[33130]_  & \new_[33125]_ ;
  assign \new_[33135]_  = A267 & A266;
  assign \new_[33136]_  = ~A265 & \new_[33135]_ ;
  assign \new_[33140]_  = A301 & ~A300;
  assign \new_[33141]_  = ~A269 & \new_[33140]_ ;
  assign \new_[33142]_  = \new_[33141]_  & \new_[33136]_ ;
  assign \new_[33146]_  = A167 & A168;
  assign \new_[33147]_  = A169 & \new_[33146]_ ;
  assign \new_[33151]_  = A202 & ~A201;
  assign \new_[33152]_  = ~A166 & \new_[33151]_ ;
  assign \new_[33153]_  = \new_[33152]_  & \new_[33147]_ ;
  assign \new_[33157]_  = A267 & A266;
  assign \new_[33158]_  = ~A265 & \new_[33157]_ ;
  assign \new_[33162]_  = ~A302 & ~A300;
  assign \new_[33163]_  = ~A269 & \new_[33162]_ ;
  assign \new_[33164]_  = \new_[33163]_  & \new_[33158]_ ;
  assign \new_[33168]_  = A167 & A168;
  assign \new_[33169]_  = A169 & \new_[33168]_ ;
  assign \new_[33173]_  = A202 & ~A201;
  assign \new_[33174]_  = ~A166 & \new_[33173]_ ;
  assign \new_[33175]_  = \new_[33174]_  & \new_[33169]_ ;
  assign \new_[33179]_  = A267 & A266;
  assign \new_[33180]_  = ~A265 & \new_[33179]_ ;
  assign \new_[33184]_  = A299 & A298;
  assign \new_[33185]_  = ~A269 & \new_[33184]_ ;
  assign \new_[33186]_  = \new_[33185]_  & \new_[33180]_ ;
  assign \new_[33190]_  = A167 & A168;
  assign \new_[33191]_  = A169 & \new_[33190]_ ;
  assign \new_[33195]_  = A202 & ~A201;
  assign \new_[33196]_  = ~A166 & \new_[33195]_ ;
  assign \new_[33197]_  = \new_[33196]_  & \new_[33191]_ ;
  assign \new_[33201]_  = A267 & A266;
  assign \new_[33202]_  = ~A265 & \new_[33201]_ ;
  assign \new_[33206]_  = ~A299 & ~A298;
  assign \new_[33207]_  = ~A269 & \new_[33206]_ ;
  assign \new_[33208]_  = \new_[33207]_  & \new_[33202]_ ;
  assign \new_[33212]_  = A167 & A168;
  assign \new_[33213]_  = A169 & \new_[33212]_ ;
  assign \new_[33217]_  = A202 & ~A201;
  assign \new_[33218]_  = ~A166 & \new_[33217]_ ;
  assign \new_[33219]_  = \new_[33218]_  & \new_[33213]_ ;
  assign \new_[33223]_  = A267 & ~A266;
  assign \new_[33224]_  = A265 & \new_[33223]_ ;
  assign \new_[33228]_  = A301 & ~A300;
  assign \new_[33229]_  = A268 & \new_[33228]_ ;
  assign \new_[33230]_  = \new_[33229]_  & \new_[33224]_ ;
  assign \new_[33234]_  = A167 & A168;
  assign \new_[33235]_  = A169 & \new_[33234]_ ;
  assign \new_[33239]_  = A202 & ~A201;
  assign \new_[33240]_  = ~A166 & \new_[33239]_ ;
  assign \new_[33241]_  = \new_[33240]_  & \new_[33235]_ ;
  assign \new_[33245]_  = A267 & ~A266;
  assign \new_[33246]_  = A265 & \new_[33245]_ ;
  assign \new_[33250]_  = ~A302 & ~A300;
  assign \new_[33251]_  = A268 & \new_[33250]_ ;
  assign \new_[33252]_  = \new_[33251]_  & \new_[33246]_ ;
  assign \new_[33256]_  = A167 & A168;
  assign \new_[33257]_  = A169 & \new_[33256]_ ;
  assign \new_[33261]_  = A202 & ~A201;
  assign \new_[33262]_  = ~A166 & \new_[33261]_ ;
  assign \new_[33263]_  = \new_[33262]_  & \new_[33257]_ ;
  assign \new_[33267]_  = A267 & ~A266;
  assign \new_[33268]_  = A265 & \new_[33267]_ ;
  assign \new_[33272]_  = A299 & A298;
  assign \new_[33273]_  = A268 & \new_[33272]_ ;
  assign \new_[33274]_  = \new_[33273]_  & \new_[33268]_ ;
  assign \new_[33278]_  = A167 & A168;
  assign \new_[33279]_  = A169 & \new_[33278]_ ;
  assign \new_[33283]_  = A202 & ~A201;
  assign \new_[33284]_  = ~A166 & \new_[33283]_ ;
  assign \new_[33285]_  = \new_[33284]_  & \new_[33279]_ ;
  assign \new_[33289]_  = A267 & ~A266;
  assign \new_[33290]_  = A265 & \new_[33289]_ ;
  assign \new_[33294]_  = ~A299 & ~A298;
  assign \new_[33295]_  = A268 & \new_[33294]_ ;
  assign \new_[33296]_  = \new_[33295]_  & \new_[33290]_ ;
  assign \new_[33300]_  = A167 & A168;
  assign \new_[33301]_  = A169 & \new_[33300]_ ;
  assign \new_[33305]_  = A202 & ~A201;
  assign \new_[33306]_  = ~A166 & \new_[33305]_ ;
  assign \new_[33307]_  = \new_[33306]_  & \new_[33301]_ ;
  assign \new_[33311]_  = A267 & ~A266;
  assign \new_[33312]_  = A265 & \new_[33311]_ ;
  assign \new_[33316]_  = A301 & ~A300;
  assign \new_[33317]_  = ~A269 & \new_[33316]_ ;
  assign \new_[33318]_  = \new_[33317]_  & \new_[33312]_ ;
  assign \new_[33322]_  = A167 & A168;
  assign \new_[33323]_  = A169 & \new_[33322]_ ;
  assign \new_[33327]_  = A202 & ~A201;
  assign \new_[33328]_  = ~A166 & \new_[33327]_ ;
  assign \new_[33329]_  = \new_[33328]_  & \new_[33323]_ ;
  assign \new_[33333]_  = A267 & ~A266;
  assign \new_[33334]_  = A265 & \new_[33333]_ ;
  assign \new_[33338]_  = ~A302 & ~A300;
  assign \new_[33339]_  = ~A269 & \new_[33338]_ ;
  assign \new_[33340]_  = \new_[33339]_  & \new_[33334]_ ;
  assign \new_[33344]_  = A167 & A168;
  assign \new_[33345]_  = A169 & \new_[33344]_ ;
  assign \new_[33349]_  = A202 & ~A201;
  assign \new_[33350]_  = ~A166 & \new_[33349]_ ;
  assign \new_[33351]_  = \new_[33350]_  & \new_[33345]_ ;
  assign \new_[33355]_  = A267 & ~A266;
  assign \new_[33356]_  = A265 & \new_[33355]_ ;
  assign \new_[33360]_  = A299 & A298;
  assign \new_[33361]_  = ~A269 & \new_[33360]_ ;
  assign \new_[33362]_  = \new_[33361]_  & \new_[33356]_ ;
  assign \new_[33366]_  = A167 & A168;
  assign \new_[33367]_  = A169 & \new_[33366]_ ;
  assign \new_[33371]_  = A202 & ~A201;
  assign \new_[33372]_  = ~A166 & \new_[33371]_ ;
  assign \new_[33373]_  = \new_[33372]_  & \new_[33367]_ ;
  assign \new_[33377]_  = A267 & ~A266;
  assign \new_[33378]_  = A265 & \new_[33377]_ ;
  assign \new_[33382]_  = ~A299 & ~A298;
  assign \new_[33383]_  = ~A269 & \new_[33382]_ ;
  assign \new_[33384]_  = \new_[33383]_  & \new_[33378]_ ;
  assign \new_[33388]_  = A167 & A168;
  assign \new_[33389]_  = A169 & \new_[33388]_ ;
  assign \new_[33393]_  = A202 & ~A201;
  assign \new_[33394]_  = ~A166 & \new_[33393]_ ;
  assign \new_[33395]_  = \new_[33394]_  & \new_[33389]_ ;
  assign \new_[33399]_  = A298 & ~A266;
  assign \new_[33400]_  = ~A265 & \new_[33399]_ ;
  assign \new_[33404]_  = A301 & A300;
  assign \new_[33405]_  = ~A299 & \new_[33404]_ ;
  assign \new_[33406]_  = \new_[33405]_  & \new_[33400]_ ;
  assign \new_[33410]_  = A167 & A168;
  assign \new_[33411]_  = A169 & \new_[33410]_ ;
  assign \new_[33415]_  = A202 & ~A201;
  assign \new_[33416]_  = ~A166 & \new_[33415]_ ;
  assign \new_[33417]_  = \new_[33416]_  & \new_[33411]_ ;
  assign \new_[33421]_  = A298 & ~A266;
  assign \new_[33422]_  = ~A265 & \new_[33421]_ ;
  assign \new_[33426]_  = ~A302 & A300;
  assign \new_[33427]_  = ~A299 & \new_[33426]_ ;
  assign \new_[33428]_  = \new_[33427]_  & \new_[33422]_ ;
  assign \new_[33432]_  = A167 & A168;
  assign \new_[33433]_  = A169 & \new_[33432]_ ;
  assign \new_[33437]_  = A202 & ~A201;
  assign \new_[33438]_  = ~A166 & \new_[33437]_ ;
  assign \new_[33439]_  = \new_[33438]_  & \new_[33433]_ ;
  assign \new_[33443]_  = ~A298 & ~A266;
  assign \new_[33444]_  = ~A265 & \new_[33443]_ ;
  assign \new_[33448]_  = A301 & A300;
  assign \new_[33449]_  = A299 & \new_[33448]_ ;
  assign \new_[33450]_  = \new_[33449]_  & \new_[33444]_ ;
  assign \new_[33454]_  = A167 & A168;
  assign \new_[33455]_  = A169 & \new_[33454]_ ;
  assign \new_[33459]_  = A202 & ~A201;
  assign \new_[33460]_  = ~A166 & \new_[33459]_ ;
  assign \new_[33461]_  = \new_[33460]_  & \new_[33455]_ ;
  assign \new_[33465]_  = ~A298 & ~A266;
  assign \new_[33466]_  = ~A265 & \new_[33465]_ ;
  assign \new_[33470]_  = ~A302 & A300;
  assign \new_[33471]_  = A299 & \new_[33470]_ ;
  assign \new_[33472]_  = \new_[33471]_  & \new_[33466]_ ;
  assign \new_[33476]_  = A167 & A168;
  assign \new_[33477]_  = A169 & \new_[33476]_ ;
  assign \new_[33481]_  = ~A203 & ~A201;
  assign \new_[33482]_  = ~A166 & \new_[33481]_ ;
  assign \new_[33483]_  = \new_[33482]_  & \new_[33477]_ ;
  assign \new_[33487]_  = A298 & A268;
  assign \new_[33488]_  = ~A267 & \new_[33487]_ ;
  assign \new_[33492]_  = A301 & A300;
  assign \new_[33493]_  = ~A299 & \new_[33492]_ ;
  assign \new_[33494]_  = \new_[33493]_  & \new_[33488]_ ;
  assign \new_[33498]_  = A167 & A168;
  assign \new_[33499]_  = A169 & \new_[33498]_ ;
  assign \new_[33503]_  = ~A203 & ~A201;
  assign \new_[33504]_  = ~A166 & \new_[33503]_ ;
  assign \new_[33505]_  = \new_[33504]_  & \new_[33499]_ ;
  assign \new_[33509]_  = A298 & A268;
  assign \new_[33510]_  = ~A267 & \new_[33509]_ ;
  assign \new_[33514]_  = ~A302 & A300;
  assign \new_[33515]_  = ~A299 & \new_[33514]_ ;
  assign \new_[33516]_  = \new_[33515]_  & \new_[33510]_ ;
  assign \new_[33520]_  = A167 & A168;
  assign \new_[33521]_  = A169 & \new_[33520]_ ;
  assign \new_[33525]_  = ~A203 & ~A201;
  assign \new_[33526]_  = ~A166 & \new_[33525]_ ;
  assign \new_[33527]_  = \new_[33526]_  & \new_[33521]_ ;
  assign \new_[33531]_  = ~A298 & A268;
  assign \new_[33532]_  = ~A267 & \new_[33531]_ ;
  assign \new_[33536]_  = A301 & A300;
  assign \new_[33537]_  = A299 & \new_[33536]_ ;
  assign \new_[33538]_  = \new_[33537]_  & \new_[33532]_ ;
  assign \new_[33542]_  = A167 & A168;
  assign \new_[33543]_  = A169 & \new_[33542]_ ;
  assign \new_[33547]_  = ~A203 & ~A201;
  assign \new_[33548]_  = ~A166 & \new_[33547]_ ;
  assign \new_[33549]_  = \new_[33548]_  & \new_[33543]_ ;
  assign \new_[33553]_  = ~A298 & A268;
  assign \new_[33554]_  = ~A267 & \new_[33553]_ ;
  assign \new_[33558]_  = ~A302 & A300;
  assign \new_[33559]_  = A299 & \new_[33558]_ ;
  assign \new_[33560]_  = \new_[33559]_  & \new_[33554]_ ;
  assign \new_[33564]_  = A167 & A168;
  assign \new_[33565]_  = A169 & \new_[33564]_ ;
  assign \new_[33569]_  = ~A203 & ~A201;
  assign \new_[33570]_  = ~A166 & \new_[33569]_ ;
  assign \new_[33571]_  = \new_[33570]_  & \new_[33565]_ ;
  assign \new_[33575]_  = A298 & ~A269;
  assign \new_[33576]_  = ~A267 & \new_[33575]_ ;
  assign \new_[33580]_  = A301 & A300;
  assign \new_[33581]_  = ~A299 & \new_[33580]_ ;
  assign \new_[33582]_  = \new_[33581]_  & \new_[33576]_ ;
  assign \new_[33586]_  = A167 & A168;
  assign \new_[33587]_  = A169 & \new_[33586]_ ;
  assign \new_[33591]_  = ~A203 & ~A201;
  assign \new_[33592]_  = ~A166 & \new_[33591]_ ;
  assign \new_[33593]_  = \new_[33592]_  & \new_[33587]_ ;
  assign \new_[33597]_  = A298 & ~A269;
  assign \new_[33598]_  = ~A267 & \new_[33597]_ ;
  assign \new_[33602]_  = ~A302 & A300;
  assign \new_[33603]_  = ~A299 & \new_[33602]_ ;
  assign \new_[33604]_  = \new_[33603]_  & \new_[33598]_ ;
  assign \new_[33608]_  = A167 & A168;
  assign \new_[33609]_  = A169 & \new_[33608]_ ;
  assign \new_[33613]_  = ~A203 & ~A201;
  assign \new_[33614]_  = ~A166 & \new_[33613]_ ;
  assign \new_[33615]_  = \new_[33614]_  & \new_[33609]_ ;
  assign \new_[33619]_  = ~A298 & ~A269;
  assign \new_[33620]_  = ~A267 & \new_[33619]_ ;
  assign \new_[33624]_  = A301 & A300;
  assign \new_[33625]_  = A299 & \new_[33624]_ ;
  assign \new_[33626]_  = \new_[33625]_  & \new_[33620]_ ;
  assign \new_[33630]_  = A167 & A168;
  assign \new_[33631]_  = A169 & \new_[33630]_ ;
  assign \new_[33635]_  = ~A203 & ~A201;
  assign \new_[33636]_  = ~A166 & \new_[33635]_ ;
  assign \new_[33637]_  = \new_[33636]_  & \new_[33631]_ ;
  assign \new_[33641]_  = ~A298 & ~A269;
  assign \new_[33642]_  = ~A267 & \new_[33641]_ ;
  assign \new_[33646]_  = ~A302 & A300;
  assign \new_[33647]_  = A299 & \new_[33646]_ ;
  assign \new_[33648]_  = \new_[33647]_  & \new_[33642]_ ;
  assign \new_[33652]_  = A167 & A168;
  assign \new_[33653]_  = A169 & \new_[33652]_ ;
  assign \new_[33657]_  = ~A203 & ~A201;
  assign \new_[33658]_  = ~A166 & \new_[33657]_ ;
  assign \new_[33659]_  = \new_[33658]_  & \new_[33653]_ ;
  assign \new_[33663]_  = A298 & A266;
  assign \new_[33664]_  = A265 & \new_[33663]_ ;
  assign \new_[33668]_  = A301 & A300;
  assign \new_[33669]_  = ~A299 & \new_[33668]_ ;
  assign \new_[33670]_  = \new_[33669]_  & \new_[33664]_ ;
  assign \new_[33674]_  = A167 & A168;
  assign \new_[33675]_  = A169 & \new_[33674]_ ;
  assign \new_[33679]_  = ~A203 & ~A201;
  assign \new_[33680]_  = ~A166 & \new_[33679]_ ;
  assign \new_[33681]_  = \new_[33680]_  & \new_[33675]_ ;
  assign \new_[33685]_  = A298 & A266;
  assign \new_[33686]_  = A265 & \new_[33685]_ ;
  assign \new_[33690]_  = ~A302 & A300;
  assign \new_[33691]_  = ~A299 & \new_[33690]_ ;
  assign \new_[33692]_  = \new_[33691]_  & \new_[33686]_ ;
  assign \new_[33696]_  = A167 & A168;
  assign \new_[33697]_  = A169 & \new_[33696]_ ;
  assign \new_[33701]_  = ~A203 & ~A201;
  assign \new_[33702]_  = ~A166 & \new_[33701]_ ;
  assign \new_[33703]_  = \new_[33702]_  & \new_[33697]_ ;
  assign \new_[33707]_  = ~A298 & A266;
  assign \new_[33708]_  = A265 & \new_[33707]_ ;
  assign \new_[33712]_  = A301 & A300;
  assign \new_[33713]_  = A299 & \new_[33712]_ ;
  assign \new_[33714]_  = \new_[33713]_  & \new_[33708]_ ;
  assign \new_[33718]_  = A167 & A168;
  assign \new_[33719]_  = A169 & \new_[33718]_ ;
  assign \new_[33723]_  = ~A203 & ~A201;
  assign \new_[33724]_  = ~A166 & \new_[33723]_ ;
  assign \new_[33725]_  = \new_[33724]_  & \new_[33719]_ ;
  assign \new_[33729]_  = ~A298 & A266;
  assign \new_[33730]_  = A265 & \new_[33729]_ ;
  assign \new_[33734]_  = ~A302 & A300;
  assign \new_[33735]_  = A299 & \new_[33734]_ ;
  assign \new_[33736]_  = \new_[33735]_  & \new_[33730]_ ;
  assign \new_[33740]_  = A167 & A168;
  assign \new_[33741]_  = A169 & \new_[33740]_ ;
  assign \new_[33745]_  = ~A203 & ~A201;
  assign \new_[33746]_  = ~A166 & \new_[33745]_ ;
  assign \new_[33747]_  = \new_[33746]_  & \new_[33741]_ ;
  assign \new_[33751]_  = A267 & A266;
  assign \new_[33752]_  = ~A265 & \new_[33751]_ ;
  assign \new_[33756]_  = A301 & ~A300;
  assign \new_[33757]_  = A268 & \new_[33756]_ ;
  assign \new_[33758]_  = \new_[33757]_  & \new_[33752]_ ;
  assign \new_[33762]_  = A167 & A168;
  assign \new_[33763]_  = A169 & \new_[33762]_ ;
  assign \new_[33767]_  = ~A203 & ~A201;
  assign \new_[33768]_  = ~A166 & \new_[33767]_ ;
  assign \new_[33769]_  = \new_[33768]_  & \new_[33763]_ ;
  assign \new_[33773]_  = A267 & A266;
  assign \new_[33774]_  = ~A265 & \new_[33773]_ ;
  assign \new_[33778]_  = ~A302 & ~A300;
  assign \new_[33779]_  = A268 & \new_[33778]_ ;
  assign \new_[33780]_  = \new_[33779]_  & \new_[33774]_ ;
  assign \new_[33784]_  = A167 & A168;
  assign \new_[33785]_  = A169 & \new_[33784]_ ;
  assign \new_[33789]_  = ~A203 & ~A201;
  assign \new_[33790]_  = ~A166 & \new_[33789]_ ;
  assign \new_[33791]_  = \new_[33790]_  & \new_[33785]_ ;
  assign \new_[33795]_  = A267 & A266;
  assign \new_[33796]_  = ~A265 & \new_[33795]_ ;
  assign \new_[33800]_  = A299 & A298;
  assign \new_[33801]_  = A268 & \new_[33800]_ ;
  assign \new_[33802]_  = \new_[33801]_  & \new_[33796]_ ;
  assign \new_[33806]_  = A167 & A168;
  assign \new_[33807]_  = A169 & \new_[33806]_ ;
  assign \new_[33811]_  = ~A203 & ~A201;
  assign \new_[33812]_  = ~A166 & \new_[33811]_ ;
  assign \new_[33813]_  = \new_[33812]_  & \new_[33807]_ ;
  assign \new_[33817]_  = A267 & A266;
  assign \new_[33818]_  = ~A265 & \new_[33817]_ ;
  assign \new_[33822]_  = ~A299 & ~A298;
  assign \new_[33823]_  = A268 & \new_[33822]_ ;
  assign \new_[33824]_  = \new_[33823]_  & \new_[33818]_ ;
  assign \new_[33828]_  = A167 & A168;
  assign \new_[33829]_  = A169 & \new_[33828]_ ;
  assign \new_[33833]_  = ~A203 & ~A201;
  assign \new_[33834]_  = ~A166 & \new_[33833]_ ;
  assign \new_[33835]_  = \new_[33834]_  & \new_[33829]_ ;
  assign \new_[33839]_  = A267 & A266;
  assign \new_[33840]_  = ~A265 & \new_[33839]_ ;
  assign \new_[33844]_  = A301 & ~A300;
  assign \new_[33845]_  = ~A269 & \new_[33844]_ ;
  assign \new_[33846]_  = \new_[33845]_  & \new_[33840]_ ;
  assign \new_[33850]_  = A167 & A168;
  assign \new_[33851]_  = A169 & \new_[33850]_ ;
  assign \new_[33855]_  = ~A203 & ~A201;
  assign \new_[33856]_  = ~A166 & \new_[33855]_ ;
  assign \new_[33857]_  = \new_[33856]_  & \new_[33851]_ ;
  assign \new_[33861]_  = A267 & A266;
  assign \new_[33862]_  = ~A265 & \new_[33861]_ ;
  assign \new_[33866]_  = ~A302 & ~A300;
  assign \new_[33867]_  = ~A269 & \new_[33866]_ ;
  assign \new_[33868]_  = \new_[33867]_  & \new_[33862]_ ;
  assign \new_[33872]_  = A167 & A168;
  assign \new_[33873]_  = A169 & \new_[33872]_ ;
  assign \new_[33877]_  = ~A203 & ~A201;
  assign \new_[33878]_  = ~A166 & \new_[33877]_ ;
  assign \new_[33879]_  = \new_[33878]_  & \new_[33873]_ ;
  assign \new_[33883]_  = A267 & A266;
  assign \new_[33884]_  = ~A265 & \new_[33883]_ ;
  assign \new_[33888]_  = A299 & A298;
  assign \new_[33889]_  = ~A269 & \new_[33888]_ ;
  assign \new_[33890]_  = \new_[33889]_  & \new_[33884]_ ;
  assign \new_[33894]_  = A167 & A168;
  assign \new_[33895]_  = A169 & \new_[33894]_ ;
  assign \new_[33899]_  = ~A203 & ~A201;
  assign \new_[33900]_  = ~A166 & \new_[33899]_ ;
  assign \new_[33901]_  = \new_[33900]_  & \new_[33895]_ ;
  assign \new_[33905]_  = A267 & A266;
  assign \new_[33906]_  = ~A265 & \new_[33905]_ ;
  assign \new_[33910]_  = ~A299 & ~A298;
  assign \new_[33911]_  = ~A269 & \new_[33910]_ ;
  assign \new_[33912]_  = \new_[33911]_  & \new_[33906]_ ;
  assign \new_[33916]_  = A167 & A168;
  assign \new_[33917]_  = A169 & \new_[33916]_ ;
  assign \new_[33921]_  = ~A203 & ~A201;
  assign \new_[33922]_  = ~A166 & \new_[33921]_ ;
  assign \new_[33923]_  = \new_[33922]_  & \new_[33917]_ ;
  assign \new_[33927]_  = A267 & ~A266;
  assign \new_[33928]_  = A265 & \new_[33927]_ ;
  assign \new_[33932]_  = A301 & ~A300;
  assign \new_[33933]_  = A268 & \new_[33932]_ ;
  assign \new_[33934]_  = \new_[33933]_  & \new_[33928]_ ;
  assign \new_[33938]_  = A167 & A168;
  assign \new_[33939]_  = A169 & \new_[33938]_ ;
  assign \new_[33943]_  = ~A203 & ~A201;
  assign \new_[33944]_  = ~A166 & \new_[33943]_ ;
  assign \new_[33945]_  = \new_[33944]_  & \new_[33939]_ ;
  assign \new_[33949]_  = A267 & ~A266;
  assign \new_[33950]_  = A265 & \new_[33949]_ ;
  assign \new_[33954]_  = ~A302 & ~A300;
  assign \new_[33955]_  = A268 & \new_[33954]_ ;
  assign \new_[33956]_  = \new_[33955]_  & \new_[33950]_ ;
  assign \new_[33960]_  = A167 & A168;
  assign \new_[33961]_  = A169 & \new_[33960]_ ;
  assign \new_[33965]_  = ~A203 & ~A201;
  assign \new_[33966]_  = ~A166 & \new_[33965]_ ;
  assign \new_[33967]_  = \new_[33966]_  & \new_[33961]_ ;
  assign \new_[33971]_  = A267 & ~A266;
  assign \new_[33972]_  = A265 & \new_[33971]_ ;
  assign \new_[33976]_  = A299 & A298;
  assign \new_[33977]_  = A268 & \new_[33976]_ ;
  assign \new_[33978]_  = \new_[33977]_  & \new_[33972]_ ;
  assign \new_[33982]_  = A167 & A168;
  assign \new_[33983]_  = A169 & \new_[33982]_ ;
  assign \new_[33987]_  = ~A203 & ~A201;
  assign \new_[33988]_  = ~A166 & \new_[33987]_ ;
  assign \new_[33989]_  = \new_[33988]_  & \new_[33983]_ ;
  assign \new_[33993]_  = A267 & ~A266;
  assign \new_[33994]_  = A265 & \new_[33993]_ ;
  assign \new_[33998]_  = ~A299 & ~A298;
  assign \new_[33999]_  = A268 & \new_[33998]_ ;
  assign \new_[34000]_  = \new_[33999]_  & \new_[33994]_ ;
  assign \new_[34004]_  = A167 & A168;
  assign \new_[34005]_  = A169 & \new_[34004]_ ;
  assign \new_[34009]_  = ~A203 & ~A201;
  assign \new_[34010]_  = ~A166 & \new_[34009]_ ;
  assign \new_[34011]_  = \new_[34010]_  & \new_[34005]_ ;
  assign \new_[34015]_  = A267 & ~A266;
  assign \new_[34016]_  = A265 & \new_[34015]_ ;
  assign \new_[34020]_  = A301 & ~A300;
  assign \new_[34021]_  = ~A269 & \new_[34020]_ ;
  assign \new_[34022]_  = \new_[34021]_  & \new_[34016]_ ;
  assign \new_[34026]_  = A167 & A168;
  assign \new_[34027]_  = A169 & \new_[34026]_ ;
  assign \new_[34031]_  = ~A203 & ~A201;
  assign \new_[34032]_  = ~A166 & \new_[34031]_ ;
  assign \new_[34033]_  = \new_[34032]_  & \new_[34027]_ ;
  assign \new_[34037]_  = A267 & ~A266;
  assign \new_[34038]_  = A265 & \new_[34037]_ ;
  assign \new_[34042]_  = ~A302 & ~A300;
  assign \new_[34043]_  = ~A269 & \new_[34042]_ ;
  assign \new_[34044]_  = \new_[34043]_  & \new_[34038]_ ;
  assign \new_[34048]_  = A167 & A168;
  assign \new_[34049]_  = A169 & \new_[34048]_ ;
  assign \new_[34053]_  = ~A203 & ~A201;
  assign \new_[34054]_  = ~A166 & \new_[34053]_ ;
  assign \new_[34055]_  = \new_[34054]_  & \new_[34049]_ ;
  assign \new_[34059]_  = A267 & ~A266;
  assign \new_[34060]_  = A265 & \new_[34059]_ ;
  assign \new_[34064]_  = A299 & A298;
  assign \new_[34065]_  = ~A269 & \new_[34064]_ ;
  assign \new_[34066]_  = \new_[34065]_  & \new_[34060]_ ;
  assign \new_[34070]_  = A167 & A168;
  assign \new_[34071]_  = A169 & \new_[34070]_ ;
  assign \new_[34075]_  = ~A203 & ~A201;
  assign \new_[34076]_  = ~A166 & \new_[34075]_ ;
  assign \new_[34077]_  = \new_[34076]_  & \new_[34071]_ ;
  assign \new_[34081]_  = A267 & ~A266;
  assign \new_[34082]_  = A265 & \new_[34081]_ ;
  assign \new_[34086]_  = ~A299 & ~A298;
  assign \new_[34087]_  = ~A269 & \new_[34086]_ ;
  assign \new_[34088]_  = \new_[34087]_  & \new_[34082]_ ;
  assign \new_[34092]_  = A167 & A168;
  assign \new_[34093]_  = A169 & \new_[34092]_ ;
  assign \new_[34097]_  = ~A203 & ~A201;
  assign \new_[34098]_  = ~A166 & \new_[34097]_ ;
  assign \new_[34099]_  = \new_[34098]_  & \new_[34093]_ ;
  assign \new_[34103]_  = A298 & ~A266;
  assign \new_[34104]_  = ~A265 & \new_[34103]_ ;
  assign \new_[34108]_  = A301 & A300;
  assign \new_[34109]_  = ~A299 & \new_[34108]_ ;
  assign \new_[34110]_  = \new_[34109]_  & \new_[34104]_ ;
  assign \new_[34114]_  = A167 & A168;
  assign \new_[34115]_  = A169 & \new_[34114]_ ;
  assign \new_[34119]_  = ~A203 & ~A201;
  assign \new_[34120]_  = ~A166 & \new_[34119]_ ;
  assign \new_[34121]_  = \new_[34120]_  & \new_[34115]_ ;
  assign \new_[34125]_  = A298 & ~A266;
  assign \new_[34126]_  = ~A265 & \new_[34125]_ ;
  assign \new_[34130]_  = ~A302 & A300;
  assign \new_[34131]_  = ~A299 & \new_[34130]_ ;
  assign \new_[34132]_  = \new_[34131]_  & \new_[34126]_ ;
  assign \new_[34136]_  = A167 & A168;
  assign \new_[34137]_  = A169 & \new_[34136]_ ;
  assign \new_[34141]_  = ~A203 & ~A201;
  assign \new_[34142]_  = ~A166 & \new_[34141]_ ;
  assign \new_[34143]_  = \new_[34142]_  & \new_[34137]_ ;
  assign \new_[34147]_  = ~A298 & ~A266;
  assign \new_[34148]_  = ~A265 & \new_[34147]_ ;
  assign \new_[34152]_  = A301 & A300;
  assign \new_[34153]_  = A299 & \new_[34152]_ ;
  assign \new_[34154]_  = \new_[34153]_  & \new_[34148]_ ;
  assign \new_[34158]_  = A167 & A168;
  assign \new_[34159]_  = A169 & \new_[34158]_ ;
  assign \new_[34163]_  = ~A203 & ~A201;
  assign \new_[34164]_  = ~A166 & \new_[34163]_ ;
  assign \new_[34165]_  = \new_[34164]_  & \new_[34159]_ ;
  assign \new_[34169]_  = ~A298 & ~A266;
  assign \new_[34170]_  = ~A265 & \new_[34169]_ ;
  assign \new_[34174]_  = ~A302 & A300;
  assign \new_[34175]_  = A299 & \new_[34174]_ ;
  assign \new_[34176]_  = \new_[34175]_  & \new_[34170]_ ;
  assign \new_[34180]_  = A167 & A168;
  assign \new_[34181]_  = A169 & \new_[34180]_ ;
  assign \new_[34185]_  = A200 & A199;
  assign \new_[34186]_  = ~A166 & \new_[34185]_ ;
  assign \new_[34187]_  = \new_[34186]_  & \new_[34181]_ ;
  assign \new_[34191]_  = A298 & A268;
  assign \new_[34192]_  = ~A267 & \new_[34191]_ ;
  assign \new_[34196]_  = A301 & A300;
  assign \new_[34197]_  = ~A299 & \new_[34196]_ ;
  assign \new_[34198]_  = \new_[34197]_  & \new_[34192]_ ;
  assign \new_[34202]_  = A167 & A168;
  assign \new_[34203]_  = A169 & \new_[34202]_ ;
  assign \new_[34207]_  = A200 & A199;
  assign \new_[34208]_  = ~A166 & \new_[34207]_ ;
  assign \new_[34209]_  = \new_[34208]_  & \new_[34203]_ ;
  assign \new_[34213]_  = A298 & A268;
  assign \new_[34214]_  = ~A267 & \new_[34213]_ ;
  assign \new_[34218]_  = ~A302 & A300;
  assign \new_[34219]_  = ~A299 & \new_[34218]_ ;
  assign \new_[34220]_  = \new_[34219]_  & \new_[34214]_ ;
  assign \new_[34224]_  = A167 & A168;
  assign \new_[34225]_  = A169 & \new_[34224]_ ;
  assign \new_[34229]_  = A200 & A199;
  assign \new_[34230]_  = ~A166 & \new_[34229]_ ;
  assign \new_[34231]_  = \new_[34230]_  & \new_[34225]_ ;
  assign \new_[34235]_  = ~A298 & A268;
  assign \new_[34236]_  = ~A267 & \new_[34235]_ ;
  assign \new_[34240]_  = A301 & A300;
  assign \new_[34241]_  = A299 & \new_[34240]_ ;
  assign \new_[34242]_  = \new_[34241]_  & \new_[34236]_ ;
  assign \new_[34246]_  = A167 & A168;
  assign \new_[34247]_  = A169 & \new_[34246]_ ;
  assign \new_[34251]_  = A200 & A199;
  assign \new_[34252]_  = ~A166 & \new_[34251]_ ;
  assign \new_[34253]_  = \new_[34252]_  & \new_[34247]_ ;
  assign \new_[34257]_  = ~A298 & A268;
  assign \new_[34258]_  = ~A267 & \new_[34257]_ ;
  assign \new_[34262]_  = ~A302 & A300;
  assign \new_[34263]_  = A299 & \new_[34262]_ ;
  assign \new_[34264]_  = \new_[34263]_  & \new_[34258]_ ;
  assign \new_[34268]_  = A167 & A168;
  assign \new_[34269]_  = A169 & \new_[34268]_ ;
  assign \new_[34273]_  = A200 & A199;
  assign \new_[34274]_  = ~A166 & \new_[34273]_ ;
  assign \new_[34275]_  = \new_[34274]_  & \new_[34269]_ ;
  assign \new_[34279]_  = A298 & ~A269;
  assign \new_[34280]_  = ~A267 & \new_[34279]_ ;
  assign \new_[34284]_  = A301 & A300;
  assign \new_[34285]_  = ~A299 & \new_[34284]_ ;
  assign \new_[34286]_  = \new_[34285]_  & \new_[34280]_ ;
  assign \new_[34290]_  = A167 & A168;
  assign \new_[34291]_  = A169 & \new_[34290]_ ;
  assign \new_[34295]_  = A200 & A199;
  assign \new_[34296]_  = ~A166 & \new_[34295]_ ;
  assign \new_[34297]_  = \new_[34296]_  & \new_[34291]_ ;
  assign \new_[34301]_  = A298 & ~A269;
  assign \new_[34302]_  = ~A267 & \new_[34301]_ ;
  assign \new_[34306]_  = ~A302 & A300;
  assign \new_[34307]_  = ~A299 & \new_[34306]_ ;
  assign \new_[34308]_  = \new_[34307]_  & \new_[34302]_ ;
  assign \new_[34312]_  = A167 & A168;
  assign \new_[34313]_  = A169 & \new_[34312]_ ;
  assign \new_[34317]_  = A200 & A199;
  assign \new_[34318]_  = ~A166 & \new_[34317]_ ;
  assign \new_[34319]_  = \new_[34318]_  & \new_[34313]_ ;
  assign \new_[34323]_  = ~A298 & ~A269;
  assign \new_[34324]_  = ~A267 & \new_[34323]_ ;
  assign \new_[34328]_  = A301 & A300;
  assign \new_[34329]_  = A299 & \new_[34328]_ ;
  assign \new_[34330]_  = \new_[34329]_  & \new_[34324]_ ;
  assign \new_[34334]_  = A167 & A168;
  assign \new_[34335]_  = A169 & \new_[34334]_ ;
  assign \new_[34339]_  = A200 & A199;
  assign \new_[34340]_  = ~A166 & \new_[34339]_ ;
  assign \new_[34341]_  = \new_[34340]_  & \new_[34335]_ ;
  assign \new_[34345]_  = ~A298 & ~A269;
  assign \new_[34346]_  = ~A267 & \new_[34345]_ ;
  assign \new_[34350]_  = ~A302 & A300;
  assign \new_[34351]_  = A299 & \new_[34350]_ ;
  assign \new_[34352]_  = \new_[34351]_  & \new_[34346]_ ;
  assign \new_[34356]_  = A167 & A168;
  assign \new_[34357]_  = A169 & \new_[34356]_ ;
  assign \new_[34361]_  = A200 & A199;
  assign \new_[34362]_  = ~A166 & \new_[34361]_ ;
  assign \new_[34363]_  = \new_[34362]_  & \new_[34357]_ ;
  assign \new_[34367]_  = A298 & A266;
  assign \new_[34368]_  = A265 & \new_[34367]_ ;
  assign \new_[34372]_  = A301 & A300;
  assign \new_[34373]_  = ~A299 & \new_[34372]_ ;
  assign \new_[34374]_  = \new_[34373]_  & \new_[34368]_ ;
  assign \new_[34378]_  = A167 & A168;
  assign \new_[34379]_  = A169 & \new_[34378]_ ;
  assign \new_[34383]_  = A200 & A199;
  assign \new_[34384]_  = ~A166 & \new_[34383]_ ;
  assign \new_[34385]_  = \new_[34384]_  & \new_[34379]_ ;
  assign \new_[34389]_  = A298 & A266;
  assign \new_[34390]_  = A265 & \new_[34389]_ ;
  assign \new_[34394]_  = ~A302 & A300;
  assign \new_[34395]_  = ~A299 & \new_[34394]_ ;
  assign \new_[34396]_  = \new_[34395]_  & \new_[34390]_ ;
  assign \new_[34400]_  = A167 & A168;
  assign \new_[34401]_  = A169 & \new_[34400]_ ;
  assign \new_[34405]_  = A200 & A199;
  assign \new_[34406]_  = ~A166 & \new_[34405]_ ;
  assign \new_[34407]_  = \new_[34406]_  & \new_[34401]_ ;
  assign \new_[34411]_  = ~A298 & A266;
  assign \new_[34412]_  = A265 & \new_[34411]_ ;
  assign \new_[34416]_  = A301 & A300;
  assign \new_[34417]_  = A299 & \new_[34416]_ ;
  assign \new_[34418]_  = \new_[34417]_  & \new_[34412]_ ;
  assign \new_[34422]_  = A167 & A168;
  assign \new_[34423]_  = A169 & \new_[34422]_ ;
  assign \new_[34427]_  = A200 & A199;
  assign \new_[34428]_  = ~A166 & \new_[34427]_ ;
  assign \new_[34429]_  = \new_[34428]_  & \new_[34423]_ ;
  assign \new_[34433]_  = ~A298 & A266;
  assign \new_[34434]_  = A265 & \new_[34433]_ ;
  assign \new_[34438]_  = ~A302 & A300;
  assign \new_[34439]_  = A299 & \new_[34438]_ ;
  assign \new_[34440]_  = \new_[34439]_  & \new_[34434]_ ;
  assign \new_[34444]_  = A167 & A168;
  assign \new_[34445]_  = A169 & \new_[34444]_ ;
  assign \new_[34449]_  = A200 & A199;
  assign \new_[34450]_  = ~A166 & \new_[34449]_ ;
  assign \new_[34451]_  = \new_[34450]_  & \new_[34445]_ ;
  assign \new_[34455]_  = A267 & A266;
  assign \new_[34456]_  = ~A265 & \new_[34455]_ ;
  assign \new_[34460]_  = A301 & ~A300;
  assign \new_[34461]_  = A268 & \new_[34460]_ ;
  assign \new_[34462]_  = \new_[34461]_  & \new_[34456]_ ;
  assign \new_[34466]_  = A167 & A168;
  assign \new_[34467]_  = A169 & \new_[34466]_ ;
  assign \new_[34471]_  = A200 & A199;
  assign \new_[34472]_  = ~A166 & \new_[34471]_ ;
  assign \new_[34473]_  = \new_[34472]_  & \new_[34467]_ ;
  assign \new_[34477]_  = A267 & A266;
  assign \new_[34478]_  = ~A265 & \new_[34477]_ ;
  assign \new_[34482]_  = ~A302 & ~A300;
  assign \new_[34483]_  = A268 & \new_[34482]_ ;
  assign \new_[34484]_  = \new_[34483]_  & \new_[34478]_ ;
  assign \new_[34488]_  = A167 & A168;
  assign \new_[34489]_  = A169 & \new_[34488]_ ;
  assign \new_[34493]_  = A200 & A199;
  assign \new_[34494]_  = ~A166 & \new_[34493]_ ;
  assign \new_[34495]_  = \new_[34494]_  & \new_[34489]_ ;
  assign \new_[34499]_  = A267 & A266;
  assign \new_[34500]_  = ~A265 & \new_[34499]_ ;
  assign \new_[34504]_  = A299 & A298;
  assign \new_[34505]_  = A268 & \new_[34504]_ ;
  assign \new_[34506]_  = \new_[34505]_  & \new_[34500]_ ;
  assign \new_[34510]_  = A167 & A168;
  assign \new_[34511]_  = A169 & \new_[34510]_ ;
  assign \new_[34515]_  = A200 & A199;
  assign \new_[34516]_  = ~A166 & \new_[34515]_ ;
  assign \new_[34517]_  = \new_[34516]_  & \new_[34511]_ ;
  assign \new_[34521]_  = A267 & A266;
  assign \new_[34522]_  = ~A265 & \new_[34521]_ ;
  assign \new_[34526]_  = ~A299 & ~A298;
  assign \new_[34527]_  = A268 & \new_[34526]_ ;
  assign \new_[34528]_  = \new_[34527]_  & \new_[34522]_ ;
  assign \new_[34532]_  = A167 & A168;
  assign \new_[34533]_  = A169 & \new_[34532]_ ;
  assign \new_[34537]_  = A200 & A199;
  assign \new_[34538]_  = ~A166 & \new_[34537]_ ;
  assign \new_[34539]_  = \new_[34538]_  & \new_[34533]_ ;
  assign \new_[34543]_  = A267 & A266;
  assign \new_[34544]_  = ~A265 & \new_[34543]_ ;
  assign \new_[34548]_  = A301 & ~A300;
  assign \new_[34549]_  = ~A269 & \new_[34548]_ ;
  assign \new_[34550]_  = \new_[34549]_  & \new_[34544]_ ;
  assign \new_[34554]_  = A167 & A168;
  assign \new_[34555]_  = A169 & \new_[34554]_ ;
  assign \new_[34559]_  = A200 & A199;
  assign \new_[34560]_  = ~A166 & \new_[34559]_ ;
  assign \new_[34561]_  = \new_[34560]_  & \new_[34555]_ ;
  assign \new_[34565]_  = A267 & A266;
  assign \new_[34566]_  = ~A265 & \new_[34565]_ ;
  assign \new_[34570]_  = ~A302 & ~A300;
  assign \new_[34571]_  = ~A269 & \new_[34570]_ ;
  assign \new_[34572]_  = \new_[34571]_  & \new_[34566]_ ;
  assign \new_[34576]_  = A167 & A168;
  assign \new_[34577]_  = A169 & \new_[34576]_ ;
  assign \new_[34581]_  = A200 & A199;
  assign \new_[34582]_  = ~A166 & \new_[34581]_ ;
  assign \new_[34583]_  = \new_[34582]_  & \new_[34577]_ ;
  assign \new_[34587]_  = A267 & A266;
  assign \new_[34588]_  = ~A265 & \new_[34587]_ ;
  assign \new_[34592]_  = A299 & A298;
  assign \new_[34593]_  = ~A269 & \new_[34592]_ ;
  assign \new_[34594]_  = \new_[34593]_  & \new_[34588]_ ;
  assign \new_[34598]_  = A167 & A168;
  assign \new_[34599]_  = A169 & \new_[34598]_ ;
  assign \new_[34603]_  = A200 & A199;
  assign \new_[34604]_  = ~A166 & \new_[34603]_ ;
  assign \new_[34605]_  = \new_[34604]_  & \new_[34599]_ ;
  assign \new_[34609]_  = A267 & A266;
  assign \new_[34610]_  = ~A265 & \new_[34609]_ ;
  assign \new_[34614]_  = ~A299 & ~A298;
  assign \new_[34615]_  = ~A269 & \new_[34614]_ ;
  assign \new_[34616]_  = \new_[34615]_  & \new_[34610]_ ;
  assign \new_[34620]_  = A167 & A168;
  assign \new_[34621]_  = A169 & \new_[34620]_ ;
  assign \new_[34625]_  = A200 & A199;
  assign \new_[34626]_  = ~A166 & \new_[34625]_ ;
  assign \new_[34627]_  = \new_[34626]_  & \new_[34621]_ ;
  assign \new_[34631]_  = A267 & ~A266;
  assign \new_[34632]_  = A265 & \new_[34631]_ ;
  assign \new_[34636]_  = A301 & ~A300;
  assign \new_[34637]_  = A268 & \new_[34636]_ ;
  assign \new_[34638]_  = \new_[34637]_  & \new_[34632]_ ;
  assign \new_[34642]_  = A167 & A168;
  assign \new_[34643]_  = A169 & \new_[34642]_ ;
  assign \new_[34647]_  = A200 & A199;
  assign \new_[34648]_  = ~A166 & \new_[34647]_ ;
  assign \new_[34649]_  = \new_[34648]_  & \new_[34643]_ ;
  assign \new_[34653]_  = A267 & ~A266;
  assign \new_[34654]_  = A265 & \new_[34653]_ ;
  assign \new_[34658]_  = ~A302 & ~A300;
  assign \new_[34659]_  = A268 & \new_[34658]_ ;
  assign \new_[34660]_  = \new_[34659]_  & \new_[34654]_ ;
  assign \new_[34664]_  = A167 & A168;
  assign \new_[34665]_  = A169 & \new_[34664]_ ;
  assign \new_[34669]_  = A200 & A199;
  assign \new_[34670]_  = ~A166 & \new_[34669]_ ;
  assign \new_[34671]_  = \new_[34670]_  & \new_[34665]_ ;
  assign \new_[34675]_  = A267 & ~A266;
  assign \new_[34676]_  = A265 & \new_[34675]_ ;
  assign \new_[34680]_  = A299 & A298;
  assign \new_[34681]_  = A268 & \new_[34680]_ ;
  assign \new_[34682]_  = \new_[34681]_  & \new_[34676]_ ;
  assign \new_[34686]_  = A167 & A168;
  assign \new_[34687]_  = A169 & \new_[34686]_ ;
  assign \new_[34691]_  = A200 & A199;
  assign \new_[34692]_  = ~A166 & \new_[34691]_ ;
  assign \new_[34693]_  = \new_[34692]_  & \new_[34687]_ ;
  assign \new_[34697]_  = A267 & ~A266;
  assign \new_[34698]_  = A265 & \new_[34697]_ ;
  assign \new_[34702]_  = ~A299 & ~A298;
  assign \new_[34703]_  = A268 & \new_[34702]_ ;
  assign \new_[34704]_  = \new_[34703]_  & \new_[34698]_ ;
  assign \new_[34708]_  = A167 & A168;
  assign \new_[34709]_  = A169 & \new_[34708]_ ;
  assign \new_[34713]_  = A200 & A199;
  assign \new_[34714]_  = ~A166 & \new_[34713]_ ;
  assign \new_[34715]_  = \new_[34714]_  & \new_[34709]_ ;
  assign \new_[34719]_  = A267 & ~A266;
  assign \new_[34720]_  = A265 & \new_[34719]_ ;
  assign \new_[34724]_  = A301 & ~A300;
  assign \new_[34725]_  = ~A269 & \new_[34724]_ ;
  assign \new_[34726]_  = \new_[34725]_  & \new_[34720]_ ;
  assign \new_[34730]_  = A167 & A168;
  assign \new_[34731]_  = A169 & \new_[34730]_ ;
  assign \new_[34735]_  = A200 & A199;
  assign \new_[34736]_  = ~A166 & \new_[34735]_ ;
  assign \new_[34737]_  = \new_[34736]_  & \new_[34731]_ ;
  assign \new_[34741]_  = A267 & ~A266;
  assign \new_[34742]_  = A265 & \new_[34741]_ ;
  assign \new_[34746]_  = ~A302 & ~A300;
  assign \new_[34747]_  = ~A269 & \new_[34746]_ ;
  assign \new_[34748]_  = \new_[34747]_  & \new_[34742]_ ;
  assign \new_[34752]_  = A167 & A168;
  assign \new_[34753]_  = A169 & \new_[34752]_ ;
  assign \new_[34757]_  = A200 & A199;
  assign \new_[34758]_  = ~A166 & \new_[34757]_ ;
  assign \new_[34759]_  = \new_[34758]_  & \new_[34753]_ ;
  assign \new_[34763]_  = A267 & ~A266;
  assign \new_[34764]_  = A265 & \new_[34763]_ ;
  assign \new_[34768]_  = A299 & A298;
  assign \new_[34769]_  = ~A269 & \new_[34768]_ ;
  assign \new_[34770]_  = \new_[34769]_  & \new_[34764]_ ;
  assign \new_[34774]_  = A167 & A168;
  assign \new_[34775]_  = A169 & \new_[34774]_ ;
  assign \new_[34779]_  = A200 & A199;
  assign \new_[34780]_  = ~A166 & \new_[34779]_ ;
  assign \new_[34781]_  = \new_[34780]_  & \new_[34775]_ ;
  assign \new_[34785]_  = A267 & ~A266;
  assign \new_[34786]_  = A265 & \new_[34785]_ ;
  assign \new_[34790]_  = ~A299 & ~A298;
  assign \new_[34791]_  = ~A269 & \new_[34790]_ ;
  assign \new_[34792]_  = \new_[34791]_  & \new_[34786]_ ;
  assign \new_[34796]_  = A167 & A168;
  assign \new_[34797]_  = A169 & \new_[34796]_ ;
  assign \new_[34801]_  = A200 & A199;
  assign \new_[34802]_  = ~A166 & \new_[34801]_ ;
  assign \new_[34803]_  = \new_[34802]_  & \new_[34797]_ ;
  assign \new_[34807]_  = A298 & ~A266;
  assign \new_[34808]_  = ~A265 & \new_[34807]_ ;
  assign \new_[34812]_  = A301 & A300;
  assign \new_[34813]_  = ~A299 & \new_[34812]_ ;
  assign \new_[34814]_  = \new_[34813]_  & \new_[34808]_ ;
  assign \new_[34818]_  = A167 & A168;
  assign \new_[34819]_  = A169 & \new_[34818]_ ;
  assign \new_[34823]_  = A200 & A199;
  assign \new_[34824]_  = ~A166 & \new_[34823]_ ;
  assign \new_[34825]_  = \new_[34824]_  & \new_[34819]_ ;
  assign \new_[34829]_  = A298 & ~A266;
  assign \new_[34830]_  = ~A265 & \new_[34829]_ ;
  assign \new_[34834]_  = ~A302 & A300;
  assign \new_[34835]_  = ~A299 & \new_[34834]_ ;
  assign \new_[34836]_  = \new_[34835]_  & \new_[34830]_ ;
  assign \new_[34840]_  = A167 & A168;
  assign \new_[34841]_  = A169 & \new_[34840]_ ;
  assign \new_[34845]_  = A200 & A199;
  assign \new_[34846]_  = ~A166 & \new_[34845]_ ;
  assign \new_[34847]_  = \new_[34846]_  & \new_[34841]_ ;
  assign \new_[34851]_  = ~A298 & ~A266;
  assign \new_[34852]_  = ~A265 & \new_[34851]_ ;
  assign \new_[34856]_  = A301 & A300;
  assign \new_[34857]_  = A299 & \new_[34856]_ ;
  assign \new_[34858]_  = \new_[34857]_  & \new_[34852]_ ;
  assign \new_[34862]_  = A167 & A168;
  assign \new_[34863]_  = A169 & \new_[34862]_ ;
  assign \new_[34867]_  = A200 & A199;
  assign \new_[34868]_  = ~A166 & \new_[34867]_ ;
  assign \new_[34869]_  = \new_[34868]_  & \new_[34863]_ ;
  assign \new_[34873]_  = ~A298 & ~A266;
  assign \new_[34874]_  = ~A265 & \new_[34873]_ ;
  assign \new_[34878]_  = ~A302 & A300;
  assign \new_[34879]_  = A299 & \new_[34878]_ ;
  assign \new_[34880]_  = \new_[34879]_  & \new_[34874]_ ;
  assign \new_[34884]_  = A167 & A168;
  assign \new_[34885]_  = A169 & \new_[34884]_ ;
  assign \new_[34889]_  = ~A200 & ~A199;
  assign \new_[34890]_  = ~A166 & \new_[34889]_ ;
  assign \new_[34891]_  = \new_[34890]_  & \new_[34885]_ ;
  assign \new_[34895]_  = A298 & A268;
  assign \new_[34896]_  = ~A267 & \new_[34895]_ ;
  assign \new_[34900]_  = A301 & A300;
  assign \new_[34901]_  = ~A299 & \new_[34900]_ ;
  assign \new_[34902]_  = \new_[34901]_  & \new_[34896]_ ;
  assign \new_[34906]_  = A167 & A168;
  assign \new_[34907]_  = A169 & \new_[34906]_ ;
  assign \new_[34911]_  = ~A200 & ~A199;
  assign \new_[34912]_  = ~A166 & \new_[34911]_ ;
  assign \new_[34913]_  = \new_[34912]_  & \new_[34907]_ ;
  assign \new_[34917]_  = A298 & A268;
  assign \new_[34918]_  = ~A267 & \new_[34917]_ ;
  assign \new_[34922]_  = ~A302 & A300;
  assign \new_[34923]_  = ~A299 & \new_[34922]_ ;
  assign \new_[34924]_  = \new_[34923]_  & \new_[34918]_ ;
  assign \new_[34928]_  = A167 & A168;
  assign \new_[34929]_  = A169 & \new_[34928]_ ;
  assign \new_[34933]_  = ~A200 & ~A199;
  assign \new_[34934]_  = ~A166 & \new_[34933]_ ;
  assign \new_[34935]_  = \new_[34934]_  & \new_[34929]_ ;
  assign \new_[34939]_  = ~A298 & A268;
  assign \new_[34940]_  = ~A267 & \new_[34939]_ ;
  assign \new_[34944]_  = A301 & A300;
  assign \new_[34945]_  = A299 & \new_[34944]_ ;
  assign \new_[34946]_  = \new_[34945]_  & \new_[34940]_ ;
  assign \new_[34950]_  = A167 & A168;
  assign \new_[34951]_  = A169 & \new_[34950]_ ;
  assign \new_[34955]_  = ~A200 & ~A199;
  assign \new_[34956]_  = ~A166 & \new_[34955]_ ;
  assign \new_[34957]_  = \new_[34956]_  & \new_[34951]_ ;
  assign \new_[34961]_  = ~A298 & A268;
  assign \new_[34962]_  = ~A267 & \new_[34961]_ ;
  assign \new_[34966]_  = ~A302 & A300;
  assign \new_[34967]_  = A299 & \new_[34966]_ ;
  assign \new_[34968]_  = \new_[34967]_  & \new_[34962]_ ;
  assign \new_[34972]_  = A167 & A168;
  assign \new_[34973]_  = A169 & \new_[34972]_ ;
  assign \new_[34977]_  = ~A200 & ~A199;
  assign \new_[34978]_  = ~A166 & \new_[34977]_ ;
  assign \new_[34979]_  = \new_[34978]_  & \new_[34973]_ ;
  assign \new_[34983]_  = A298 & ~A269;
  assign \new_[34984]_  = ~A267 & \new_[34983]_ ;
  assign \new_[34988]_  = A301 & A300;
  assign \new_[34989]_  = ~A299 & \new_[34988]_ ;
  assign \new_[34990]_  = \new_[34989]_  & \new_[34984]_ ;
  assign \new_[34994]_  = A167 & A168;
  assign \new_[34995]_  = A169 & \new_[34994]_ ;
  assign \new_[34999]_  = ~A200 & ~A199;
  assign \new_[35000]_  = ~A166 & \new_[34999]_ ;
  assign \new_[35001]_  = \new_[35000]_  & \new_[34995]_ ;
  assign \new_[35005]_  = A298 & ~A269;
  assign \new_[35006]_  = ~A267 & \new_[35005]_ ;
  assign \new_[35010]_  = ~A302 & A300;
  assign \new_[35011]_  = ~A299 & \new_[35010]_ ;
  assign \new_[35012]_  = \new_[35011]_  & \new_[35006]_ ;
  assign \new_[35016]_  = A167 & A168;
  assign \new_[35017]_  = A169 & \new_[35016]_ ;
  assign \new_[35021]_  = ~A200 & ~A199;
  assign \new_[35022]_  = ~A166 & \new_[35021]_ ;
  assign \new_[35023]_  = \new_[35022]_  & \new_[35017]_ ;
  assign \new_[35027]_  = ~A298 & ~A269;
  assign \new_[35028]_  = ~A267 & \new_[35027]_ ;
  assign \new_[35032]_  = A301 & A300;
  assign \new_[35033]_  = A299 & \new_[35032]_ ;
  assign \new_[35034]_  = \new_[35033]_  & \new_[35028]_ ;
  assign \new_[35038]_  = A167 & A168;
  assign \new_[35039]_  = A169 & \new_[35038]_ ;
  assign \new_[35043]_  = ~A200 & ~A199;
  assign \new_[35044]_  = ~A166 & \new_[35043]_ ;
  assign \new_[35045]_  = \new_[35044]_  & \new_[35039]_ ;
  assign \new_[35049]_  = ~A298 & ~A269;
  assign \new_[35050]_  = ~A267 & \new_[35049]_ ;
  assign \new_[35054]_  = ~A302 & A300;
  assign \new_[35055]_  = A299 & \new_[35054]_ ;
  assign \new_[35056]_  = \new_[35055]_  & \new_[35050]_ ;
  assign \new_[35060]_  = A167 & A168;
  assign \new_[35061]_  = A169 & \new_[35060]_ ;
  assign \new_[35065]_  = ~A200 & ~A199;
  assign \new_[35066]_  = ~A166 & \new_[35065]_ ;
  assign \new_[35067]_  = \new_[35066]_  & \new_[35061]_ ;
  assign \new_[35071]_  = A298 & A266;
  assign \new_[35072]_  = A265 & \new_[35071]_ ;
  assign \new_[35076]_  = A301 & A300;
  assign \new_[35077]_  = ~A299 & \new_[35076]_ ;
  assign \new_[35078]_  = \new_[35077]_  & \new_[35072]_ ;
  assign \new_[35082]_  = A167 & A168;
  assign \new_[35083]_  = A169 & \new_[35082]_ ;
  assign \new_[35087]_  = ~A200 & ~A199;
  assign \new_[35088]_  = ~A166 & \new_[35087]_ ;
  assign \new_[35089]_  = \new_[35088]_  & \new_[35083]_ ;
  assign \new_[35093]_  = A298 & A266;
  assign \new_[35094]_  = A265 & \new_[35093]_ ;
  assign \new_[35098]_  = ~A302 & A300;
  assign \new_[35099]_  = ~A299 & \new_[35098]_ ;
  assign \new_[35100]_  = \new_[35099]_  & \new_[35094]_ ;
  assign \new_[35104]_  = A167 & A168;
  assign \new_[35105]_  = A169 & \new_[35104]_ ;
  assign \new_[35109]_  = ~A200 & ~A199;
  assign \new_[35110]_  = ~A166 & \new_[35109]_ ;
  assign \new_[35111]_  = \new_[35110]_  & \new_[35105]_ ;
  assign \new_[35115]_  = ~A298 & A266;
  assign \new_[35116]_  = A265 & \new_[35115]_ ;
  assign \new_[35120]_  = A301 & A300;
  assign \new_[35121]_  = A299 & \new_[35120]_ ;
  assign \new_[35122]_  = \new_[35121]_  & \new_[35116]_ ;
  assign \new_[35126]_  = A167 & A168;
  assign \new_[35127]_  = A169 & \new_[35126]_ ;
  assign \new_[35131]_  = ~A200 & ~A199;
  assign \new_[35132]_  = ~A166 & \new_[35131]_ ;
  assign \new_[35133]_  = \new_[35132]_  & \new_[35127]_ ;
  assign \new_[35137]_  = ~A298 & A266;
  assign \new_[35138]_  = A265 & \new_[35137]_ ;
  assign \new_[35142]_  = ~A302 & A300;
  assign \new_[35143]_  = A299 & \new_[35142]_ ;
  assign \new_[35144]_  = \new_[35143]_  & \new_[35138]_ ;
  assign \new_[35148]_  = A167 & A168;
  assign \new_[35149]_  = A169 & \new_[35148]_ ;
  assign \new_[35153]_  = ~A200 & ~A199;
  assign \new_[35154]_  = ~A166 & \new_[35153]_ ;
  assign \new_[35155]_  = \new_[35154]_  & \new_[35149]_ ;
  assign \new_[35159]_  = A267 & A266;
  assign \new_[35160]_  = ~A265 & \new_[35159]_ ;
  assign \new_[35164]_  = A301 & ~A300;
  assign \new_[35165]_  = A268 & \new_[35164]_ ;
  assign \new_[35166]_  = \new_[35165]_  & \new_[35160]_ ;
  assign \new_[35170]_  = A167 & A168;
  assign \new_[35171]_  = A169 & \new_[35170]_ ;
  assign \new_[35175]_  = ~A200 & ~A199;
  assign \new_[35176]_  = ~A166 & \new_[35175]_ ;
  assign \new_[35177]_  = \new_[35176]_  & \new_[35171]_ ;
  assign \new_[35181]_  = A267 & A266;
  assign \new_[35182]_  = ~A265 & \new_[35181]_ ;
  assign \new_[35186]_  = ~A302 & ~A300;
  assign \new_[35187]_  = A268 & \new_[35186]_ ;
  assign \new_[35188]_  = \new_[35187]_  & \new_[35182]_ ;
  assign \new_[35192]_  = A167 & A168;
  assign \new_[35193]_  = A169 & \new_[35192]_ ;
  assign \new_[35197]_  = ~A200 & ~A199;
  assign \new_[35198]_  = ~A166 & \new_[35197]_ ;
  assign \new_[35199]_  = \new_[35198]_  & \new_[35193]_ ;
  assign \new_[35203]_  = A267 & A266;
  assign \new_[35204]_  = ~A265 & \new_[35203]_ ;
  assign \new_[35208]_  = A299 & A298;
  assign \new_[35209]_  = A268 & \new_[35208]_ ;
  assign \new_[35210]_  = \new_[35209]_  & \new_[35204]_ ;
  assign \new_[35214]_  = A167 & A168;
  assign \new_[35215]_  = A169 & \new_[35214]_ ;
  assign \new_[35219]_  = ~A200 & ~A199;
  assign \new_[35220]_  = ~A166 & \new_[35219]_ ;
  assign \new_[35221]_  = \new_[35220]_  & \new_[35215]_ ;
  assign \new_[35225]_  = A267 & A266;
  assign \new_[35226]_  = ~A265 & \new_[35225]_ ;
  assign \new_[35230]_  = ~A299 & ~A298;
  assign \new_[35231]_  = A268 & \new_[35230]_ ;
  assign \new_[35232]_  = \new_[35231]_  & \new_[35226]_ ;
  assign \new_[35236]_  = A167 & A168;
  assign \new_[35237]_  = A169 & \new_[35236]_ ;
  assign \new_[35241]_  = ~A200 & ~A199;
  assign \new_[35242]_  = ~A166 & \new_[35241]_ ;
  assign \new_[35243]_  = \new_[35242]_  & \new_[35237]_ ;
  assign \new_[35247]_  = A267 & A266;
  assign \new_[35248]_  = ~A265 & \new_[35247]_ ;
  assign \new_[35252]_  = A301 & ~A300;
  assign \new_[35253]_  = ~A269 & \new_[35252]_ ;
  assign \new_[35254]_  = \new_[35253]_  & \new_[35248]_ ;
  assign \new_[35258]_  = A167 & A168;
  assign \new_[35259]_  = A169 & \new_[35258]_ ;
  assign \new_[35263]_  = ~A200 & ~A199;
  assign \new_[35264]_  = ~A166 & \new_[35263]_ ;
  assign \new_[35265]_  = \new_[35264]_  & \new_[35259]_ ;
  assign \new_[35269]_  = A267 & A266;
  assign \new_[35270]_  = ~A265 & \new_[35269]_ ;
  assign \new_[35274]_  = ~A302 & ~A300;
  assign \new_[35275]_  = ~A269 & \new_[35274]_ ;
  assign \new_[35276]_  = \new_[35275]_  & \new_[35270]_ ;
  assign \new_[35280]_  = A167 & A168;
  assign \new_[35281]_  = A169 & \new_[35280]_ ;
  assign \new_[35285]_  = ~A200 & ~A199;
  assign \new_[35286]_  = ~A166 & \new_[35285]_ ;
  assign \new_[35287]_  = \new_[35286]_  & \new_[35281]_ ;
  assign \new_[35291]_  = A267 & A266;
  assign \new_[35292]_  = ~A265 & \new_[35291]_ ;
  assign \new_[35296]_  = A299 & A298;
  assign \new_[35297]_  = ~A269 & \new_[35296]_ ;
  assign \new_[35298]_  = \new_[35297]_  & \new_[35292]_ ;
  assign \new_[35302]_  = A167 & A168;
  assign \new_[35303]_  = A169 & \new_[35302]_ ;
  assign \new_[35307]_  = ~A200 & ~A199;
  assign \new_[35308]_  = ~A166 & \new_[35307]_ ;
  assign \new_[35309]_  = \new_[35308]_  & \new_[35303]_ ;
  assign \new_[35313]_  = A267 & A266;
  assign \new_[35314]_  = ~A265 & \new_[35313]_ ;
  assign \new_[35318]_  = ~A299 & ~A298;
  assign \new_[35319]_  = ~A269 & \new_[35318]_ ;
  assign \new_[35320]_  = \new_[35319]_  & \new_[35314]_ ;
  assign \new_[35324]_  = A167 & A168;
  assign \new_[35325]_  = A169 & \new_[35324]_ ;
  assign \new_[35329]_  = ~A200 & ~A199;
  assign \new_[35330]_  = ~A166 & \new_[35329]_ ;
  assign \new_[35331]_  = \new_[35330]_  & \new_[35325]_ ;
  assign \new_[35335]_  = A267 & ~A266;
  assign \new_[35336]_  = A265 & \new_[35335]_ ;
  assign \new_[35340]_  = A301 & ~A300;
  assign \new_[35341]_  = A268 & \new_[35340]_ ;
  assign \new_[35342]_  = \new_[35341]_  & \new_[35336]_ ;
  assign \new_[35346]_  = A167 & A168;
  assign \new_[35347]_  = A169 & \new_[35346]_ ;
  assign \new_[35351]_  = ~A200 & ~A199;
  assign \new_[35352]_  = ~A166 & \new_[35351]_ ;
  assign \new_[35353]_  = \new_[35352]_  & \new_[35347]_ ;
  assign \new_[35357]_  = A267 & ~A266;
  assign \new_[35358]_  = A265 & \new_[35357]_ ;
  assign \new_[35362]_  = ~A302 & ~A300;
  assign \new_[35363]_  = A268 & \new_[35362]_ ;
  assign \new_[35364]_  = \new_[35363]_  & \new_[35358]_ ;
  assign \new_[35368]_  = A167 & A168;
  assign \new_[35369]_  = A169 & \new_[35368]_ ;
  assign \new_[35373]_  = ~A200 & ~A199;
  assign \new_[35374]_  = ~A166 & \new_[35373]_ ;
  assign \new_[35375]_  = \new_[35374]_  & \new_[35369]_ ;
  assign \new_[35379]_  = A267 & ~A266;
  assign \new_[35380]_  = A265 & \new_[35379]_ ;
  assign \new_[35384]_  = A299 & A298;
  assign \new_[35385]_  = A268 & \new_[35384]_ ;
  assign \new_[35386]_  = \new_[35385]_  & \new_[35380]_ ;
  assign \new_[35390]_  = A167 & A168;
  assign \new_[35391]_  = A169 & \new_[35390]_ ;
  assign \new_[35395]_  = ~A200 & ~A199;
  assign \new_[35396]_  = ~A166 & \new_[35395]_ ;
  assign \new_[35397]_  = \new_[35396]_  & \new_[35391]_ ;
  assign \new_[35401]_  = A267 & ~A266;
  assign \new_[35402]_  = A265 & \new_[35401]_ ;
  assign \new_[35406]_  = ~A299 & ~A298;
  assign \new_[35407]_  = A268 & \new_[35406]_ ;
  assign \new_[35408]_  = \new_[35407]_  & \new_[35402]_ ;
  assign \new_[35412]_  = A167 & A168;
  assign \new_[35413]_  = A169 & \new_[35412]_ ;
  assign \new_[35417]_  = ~A200 & ~A199;
  assign \new_[35418]_  = ~A166 & \new_[35417]_ ;
  assign \new_[35419]_  = \new_[35418]_  & \new_[35413]_ ;
  assign \new_[35423]_  = A267 & ~A266;
  assign \new_[35424]_  = A265 & \new_[35423]_ ;
  assign \new_[35428]_  = A301 & ~A300;
  assign \new_[35429]_  = ~A269 & \new_[35428]_ ;
  assign \new_[35430]_  = \new_[35429]_  & \new_[35424]_ ;
  assign \new_[35434]_  = A167 & A168;
  assign \new_[35435]_  = A169 & \new_[35434]_ ;
  assign \new_[35439]_  = ~A200 & ~A199;
  assign \new_[35440]_  = ~A166 & \new_[35439]_ ;
  assign \new_[35441]_  = \new_[35440]_  & \new_[35435]_ ;
  assign \new_[35445]_  = A267 & ~A266;
  assign \new_[35446]_  = A265 & \new_[35445]_ ;
  assign \new_[35450]_  = ~A302 & ~A300;
  assign \new_[35451]_  = ~A269 & \new_[35450]_ ;
  assign \new_[35452]_  = \new_[35451]_  & \new_[35446]_ ;
  assign \new_[35456]_  = A167 & A168;
  assign \new_[35457]_  = A169 & \new_[35456]_ ;
  assign \new_[35461]_  = ~A200 & ~A199;
  assign \new_[35462]_  = ~A166 & \new_[35461]_ ;
  assign \new_[35463]_  = \new_[35462]_  & \new_[35457]_ ;
  assign \new_[35467]_  = A267 & ~A266;
  assign \new_[35468]_  = A265 & \new_[35467]_ ;
  assign \new_[35472]_  = A299 & A298;
  assign \new_[35473]_  = ~A269 & \new_[35472]_ ;
  assign \new_[35474]_  = \new_[35473]_  & \new_[35468]_ ;
  assign \new_[35478]_  = A167 & A168;
  assign \new_[35479]_  = A169 & \new_[35478]_ ;
  assign \new_[35483]_  = ~A200 & ~A199;
  assign \new_[35484]_  = ~A166 & \new_[35483]_ ;
  assign \new_[35485]_  = \new_[35484]_  & \new_[35479]_ ;
  assign \new_[35489]_  = A267 & ~A266;
  assign \new_[35490]_  = A265 & \new_[35489]_ ;
  assign \new_[35494]_  = ~A299 & ~A298;
  assign \new_[35495]_  = ~A269 & \new_[35494]_ ;
  assign \new_[35496]_  = \new_[35495]_  & \new_[35490]_ ;
  assign \new_[35500]_  = A167 & A168;
  assign \new_[35501]_  = A169 & \new_[35500]_ ;
  assign \new_[35505]_  = ~A200 & ~A199;
  assign \new_[35506]_  = ~A166 & \new_[35505]_ ;
  assign \new_[35507]_  = \new_[35506]_  & \new_[35501]_ ;
  assign \new_[35511]_  = A298 & ~A266;
  assign \new_[35512]_  = ~A265 & \new_[35511]_ ;
  assign \new_[35516]_  = A301 & A300;
  assign \new_[35517]_  = ~A299 & \new_[35516]_ ;
  assign \new_[35518]_  = \new_[35517]_  & \new_[35512]_ ;
  assign \new_[35522]_  = A167 & A168;
  assign \new_[35523]_  = A169 & \new_[35522]_ ;
  assign \new_[35527]_  = ~A200 & ~A199;
  assign \new_[35528]_  = ~A166 & \new_[35527]_ ;
  assign \new_[35529]_  = \new_[35528]_  & \new_[35523]_ ;
  assign \new_[35533]_  = A298 & ~A266;
  assign \new_[35534]_  = ~A265 & \new_[35533]_ ;
  assign \new_[35538]_  = ~A302 & A300;
  assign \new_[35539]_  = ~A299 & \new_[35538]_ ;
  assign \new_[35540]_  = \new_[35539]_  & \new_[35534]_ ;
  assign \new_[35544]_  = A167 & A168;
  assign \new_[35545]_  = A169 & \new_[35544]_ ;
  assign \new_[35549]_  = ~A200 & ~A199;
  assign \new_[35550]_  = ~A166 & \new_[35549]_ ;
  assign \new_[35551]_  = \new_[35550]_  & \new_[35545]_ ;
  assign \new_[35555]_  = ~A298 & ~A266;
  assign \new_[35556]_  = ~A265 & \new_[35555]_ ;
  assign \new_[35560]_  = A301 & A300;
  assign \new_[35561]_  = A299 & \new_[35560]_ ;
  assign \new_[35562]_  = \new_[35561]_  & \new_[35556]_ ;
  assign \new_[35566]_  = A167 & A168;
  assign \new_[35567]_  = A169 & \new_[35566]_ ;
  assign \new_[35571]_  = ~A200 & ~A199;
  assign \new_[35572]_  = ~A166 & \new_[35571]_ ;
  assign \new_[35573]_  = \new_[35572]_  & \new_[35567]_ ;
  assign \new_[35577]_  = ~A298 & ~A266;
  assign \new_[35578]_  = ~A265 & \new_[35577]_ ;
  assign \new_[35582]_  = ~A302 & A300;
  assign \new_[35583]_  = A299 & \new_[35582]_ ;
  assign \new_[35584]_  = \new_[35583]_  & \new_[35578]_ ;
  assign \new_[35588]_  = ~A167 & A168;
  assign \new_[35589]_  = A169 & \new_[35588]_ ;
  assign \new_[35593]_  = A202 & ~A201;
  assign \new_[35594]_  = A166 & \new_[35593]_ ;
  assign \new_[35595]_  = \new_[35594]_  & \new_[35589]_ ;
  assign \new_[35599]_  = A298 & A268;
  assign \new_[35600]_  = ~A267 & \new_[35599]_ ;
  assign \new_[35604]_  = A301 & A300;
  assign \new_[35605]_  = ~A299 & \new_[35604]_ ;
  assign \new_[35606]_  = \new_[35605]_  & \new_[35600]_ ;
  assign \new_[35610]_  = ~A167 & A168;
  assign \new_[35611]_  = A169 & \new_[35610]_ ;
  assign \new_[35615]_  = A202 & ~A201;
  assign \new_[35616]_  = A166 & \new_[35615]_ ;
  assign \new_[35617]_  = \new_[35616]_  & \new_[35611]_ ;
  assign \new_[35621]_  = A298 & A268;
  assign \new_[35622]_  = ~A267 & \new_[35621]_ ;
  assign \new_[35626]_  = ~A302 & A300;
  assign \new_[35627]_  = ~A299 & \new_[35626]_ ;
  assign \new_[35628]_  = \new_[35627]_  & \new_[35622]_ ;
  assign \new_[35632]_  = ~A167 & A168;
  assign \new_[35633]_  = A169 & \new_[35632]_ ;
  assign \new_[35637]_  = A202 & ~A201;
  assign \new_[35638]_  = A166 & \new_[35637]_ ;
  assign \new_[35639]_  = \new_[35638]_  & \new_[35633]_ ;
  assign \new_[35643]_  = ~A298 & A268;
  assign \new_[35644]_  = ~A267 & \new_[35643]_ ;
  assign \new_[35648]_  = A301 & A300;
  assign \new_[35649]_  = A299 & \new_[35648]_ ;
  assign \new_[35650]_  = \new_[35649]_  & \new_[35644]_ ;
  assign \new_[35654]_  = ~A167 & A168;
  assign \new_[35655]_  = A169 & \new_[35654]_ ;
  assign \new_[35659]_  = A202 & ~A201;
  assign \new_[35660]_  = A166 & \new_[35659]_ ;
  assign \new_[35661]_  = \new_[35660]_  & \new_[35655]_ ;
  assign \new_[35665]_  = ~A298 & A268;
  assign \new_[35666]_  = ~A267 & \new_[35665]_ ;
  assign \new_[35670]_  = ~A302 & A300;
  assign \new_[35671]_  = A299 & \new_[35670]_ ;
  assign \new_[35672]_  = \new_[35671]_  & \new_[35666]_ ;
  assign \new_[35676]_  = ~A167 & A168;
  assign \new_[35677]_  = A169 & \new_[35676]_ ;
  assign \new_[35681]_  = A202 & ~A201;
  assign \new_[35682]_  = A166 & \new_[35681]_ ;
  assign \new_[35683]_  = \new_[35682]_  & \new_[35677]_ ;
  assign \new_[35687]_  = A298 & ~A269;
  assign \new_[35688]_  = ~A267 & \new_[35687]_ ;
  assign \new_[35692]_  = A301 & A300;
  assign \new_[35693]_  = ~A299 & \new_[35692]_ ;
  assign \new_[35694]_  = \new_[35693]_  & \new_[35688]_ ;
  assign \new_[35698]_  = ~A167 & A168;
  assign \new_[35699]_  = A169 & \new_[35698]_ ;
  assign \new_[35703]_  = A202 & ~A201;
  assign \new_[35704]_  = A166 & \new_[35703]_ ;
  assign \new_[35705]_  = \new_[35704]_  & \new_[35699]_ ;
  assign \new_[35709]_  = A298 & ~A269;
  assign \new_[35710]_  = ~A267 & \new_[35709]_ ;
  assign \new_[35714]_  = ~A302 & A300;
  assign \new_[35715]_  = ~A299 & \new_[35714]_ ;
  assign \new_[35716]_  = \new_[35715]_  & \new_[35710]_ ;
  assign \new_[35720]_  = ~A167 & A168;
  assign \new_[35721]_  = A169 & \new_[35720]_ ;
  assign \new_[35725]_  = A202 & ~A201;
  assign \new_[35726]_  = A166 & \new_[35725]_ ;
  assign \new_[35727]_  = \new_[35726]_  & \new_[35721]_ ;
  assign \new_[35731]_  = ~A298 & ~A269;
  assign \new_[35732]_  = ~A267 & \new_[35731]_ ;
  assign \new_[35736]_  = A301 & A300;
  assign \new_[35737]_  = A299 & \new_[35736]_ ;
  assign \new_[35738]_  = \new_[35737]_  & \new_[35732]_ ;
  assign \new_[35742]_  = ~A167 & A168;
  assign \new_[35743]_  = A169 & \new_[35742]_ ;
  assign \new_[35747]_  = A202 & ~A201;
  assign \new_[35748]_  = A166 & \new_[35747]_ ;
  assign \new_[35749]_  = \new_[35748]_  & \new_[35743]_ ;
  assign \new_[35753]_  = ~A298 & ~A269;
  assign \new_[35754]_  = ~A267 & \new_[35753]_ ;
  assign \new_[35758]_  = ~A302 & A300;
  assign \new_[35759]_  = A299 & \new_[35758]_ ;
  assign \new_[35760]_  = \new_[35759]_  & \new_[35754]_ ;
  assign \new_[35764]_  = ~A167 & A168;
  assign \new_[35765]_  = A169 & \new_[35764]_ ;
  assign \new_[35769]_  = A202 & ~A201;
  assign \new_[35770]_  = A166 & \new_[35769]_ ;
  assign \new_[35771]_  = \new_[35770]_  & \new_[35765]_ ;
  assign \new_[35775]_  = A298 & A266;
  assign \new_[35776]_  = A265 & \new_[35775]_ ;
  assign \new_[35780]_  = A301 & A300;
  assign \new_[35781]_  = ~A299 & \new_[35780]_ ;
  assign \new_[35782]_  = \new_[35781]_  & \new_[35776]_ ;
  assign \new_[35786]_  = ~A167 & A168;
  assign \new_[35787]_  = A169 & \new_[35786]_ ;
  assign \new_[35791]_  = A202 & ~A201;
  assign \new_[35792]_  = A166 & \new_[35791]_ ;
  assign \new_[35793]_  = \new_[35792]_  & \new_[35787]_ ;
  assign \new_[35797]_  = A298 & A266;
  assign \new_[35798]_  = A265 & \new_[35797]_ ;
  assign \new_[35802]_  = ~A302 & A300;
  assign \new_[35803]_  = ~A299 & \new_[35802]_ ;
  assign \new_[35804]_  = \new_[35803]_  & \new_[35798]_ ;
  assign \new_[35808]_  = ~A167 & A168;
  assign \new_[35809]_  = A169 & \new_[35808]_ ;
  assign \new_[35813]_  = A202 & ~A201;
  assign \new_[35814]_  = A166 & \new_[35813]_ ;
  assign \new_[35815]_  = \new_[35814]_  & \new_[35809]_ ;
  assign \new_[35819]_  = ~A298 & A266;
  assign \new_[35820]_  = A265 & \new_[35819]_ ;
  assign \new_[35824]_  = A301 & A300;
  assign \new_[35825]_  = A299 & \new_[35824]_ ;
  assign \new_[35826]_  = \new_[35825]_  & \new_[35820]_ ;
  assign \new_[35830]_  = ~A167 & A168;
  assign \new_[35831]_  = A169 & \new_[35830]_ ;
  assign \new_[35835]_  = A202 & ~A201;
  assign \new_[35836]_  = A166 & \new_[35835]_ ;
  assign \new_[35837]_  = \new_[35836]_  & \new_[35831]_ ;
  assign \new_[35841]_  = ~A298 & A266;
  assign \new_[35842]_  = A265 & \new_[35841]_ ;
  assign \new_[35846]_  = ~A302 & A300;
  assign \new_[35847]_  = A299 & \new_[35846]_ ;
  assign \new_[35848]_  = \new_[35847]_  & \new_[35842]_ ;
  assign \new_[35852]_  = ~A167 & A168;
  assign \new_[35853]_  = A169 & \new_[35852]_ ;
  assign \new_[35857]_  = A202 & ~A201;
  assign \new_[35858]_  = A166 & \new_[35857]_ ;
  assign \new_[35859]_  = \new_[35858]_  & \new_[35853]_ ;
  assign \new_[35863]_  = A267 & A266;
  assign \new_[35864]_  = ~A265 & \new_[35863]_ ;
  assign \new_[35868]_  = A301 & ~A300;
  assign \new_[35869]_  = A268 & \new_[35868]_ ;
  assign \new_[35870]_  = \new_[35869]_  & \new_[35864]_ ;
  assign \new_[35874]_  = ~A167 & A168;
  assign \new_[35875]_  = A169 & \new_[35874]_ ;
  assign \new_[35879]_  = A202 & ~A201;
  assign \new_[35880]_  = A166 & \new_[35879]_ ;
  assign \new_[35881]_  = \new_[35880]_  & \new_[35875]_ ;
  assign \new_[35885]_  = A267 & A266;
  assign \new_[35886]_  = ~A265 & \new_[35885]_ ;
  assign \new_[35890]_  = ~A302 & ~A300;
  assign \new_[35891]_  = A268 & \new_[35890]_ ;
  assign \new_[35892]_  = \new_[35891]_  & \new_[35886]_ ;
  assign \new_[35896]_  = ~A167 & A168;
  assign \new_[35897]_  = A169 & \new_[35896]_ ;
  assign \new_[35901]_  = A202 & ~A201;
  assign \new_[35902]_  = A166 & \new_[35901]_ ;
  assign \new_[35903]_  = \new_[35902]_  & \new_[35897]_ ;
  assign \new_[35907]_  = A267 & A266;
  assign \new_[35908]_  = ~A265 & \new_[35907]_ ;
  assign \new_[35912]_  = A299 & A298;
  assign \new_[35913]_  = A268 & \new_[35912]_ ;
  assign \new_[35914]_  = \new_[35913]_  & \new_[35908]_ ;
  assign \new_[35918]_  = ~A167 & A168;
  assign \new_[35919]_  = A169 & \new_[35918]_ ;
  assign \new_[35923]_  = A202 & ~A201;
  assign \new_[35924]_  = A166 & \new_[35923]_ ;
  assign \new_[35925]_  = \new_[35924]_  & \new_[35919]_ ;
  assign \new_[35929]_  = A267 & A266;
  assign \new_[35930]_  = ~A265 & \new_[35929]_ ;
  assign \new_[35934]_  = ~A299 & ~A298;
  assign \new_[35935]_  = A268 & \new_[35934]_ ;
  assign \new_[35936]_  = \new_[35935]_  & \new_[35930]_ ;
  assign \new_[35940]_  = ~A167 & A168;
  assign \new_[35941]_  = A169 & \new_[35940]_ ;
  assign \new_[35945]_  = A202 & ~A201;
  assign \new_[35946]_  = A166 & \new_[35945]_ ;
  assign \new_[35947]_  = \new_[35946]_  & \new_[35941]_ ;
  assign \new_[35951]_  = A267 & A266;
  assign \new_[35952]_  = ~A265 & \new_[35951]_ ;
  assign \new_[35956]_  = A301 & ~A300;
  assign \new_[35957]_  = ~A269 & \new_[35956]_ ;
  assign \new_[35958]_  = \new_[35957]_  & \new_[35952]_ ;
  assign \new_[35962]_  = ~A167 & A168;
  assign \new_[35963]_  = A169 & \new_[35962]_ ;
  assign \new_[35967]_  = A202 & ~A201;
  assign \new_[35968]_  = A166 & \new_[35967]_ ;
  assign \new_[35969]_  = \new_[35968]_  & \new_[35963]_ ;
  assign \new_[35973]_  = A267 & A266;
  assign \new_[35974]_  = ~A265 & \new_[35973]_ ;
  assign \new_[35978]_  = ~A302 & ~A300;
  assign \new_[35979]_  = ~A269 & \new_[35978]_ ;
  assign \new_[35980]_  = \new_[35979]_  & \new_[35974]_ ;
  assign \new_[35984]_  = ~A167 & A168;
  assign \new_[35985]_  = A169 & \new_[35984]_ ;
  assign \new_[35989]_  = A202 & ~A201;
  assign \new_[35990]_  = A166 & \new_[35989]_ ;
  assign \new_[35991]_  = \new_[35990]_  & \new_[35985]_ ;
  assign \new_[35995]_  = A267 & A266;
  assign \new_[35996]_  = ~A265 & \new_[35995]_ ;
  assign \new_[36000]_  = A299 & A298;
  assign \new_[36001]_  = ~A269 & \new_[36000]_ ;
  assign \new_[36002]_  = \new_[36001]_  & \new_[35996]_ ;
  assign \new_[36006]_  = ~A167 & A168;
  assign \new_[36007]_  = A169 & \new_[36006]_ ;
  assign \new_[36011]_  = A202 & ~A201;
  assign \new_[36012]_  = A166 & \new_[36011]_ ;
  assign \new_[36013]_  = \new_[36012]_  & \new_[36007]_ ;
  assign \new_[36017]_  = A267 & A266;
  assign \new_[36018]_  = ~A265 & \new_[36017]_ ;
  assign \new_[36022]_  = ~A299 & ~A298;
  assign \new_[36023]_  = ~A269 & \new_[36022]_ ;
  assign \new_[36024]_  = \new_[36023]_  & \new_[36018]_ ;
  assign \new_[36028]_  = ~A167 & A168;
  assign \new_[36029]_  = A169 & \new_[36028]_ ;
  assign \new_[36033]_  = A202 & ~A201;
  assign \new_[36034]_  = A166 & \new_[36033]_ ;
  assign \new_[36035]_  = \new_[36034]_  & \new_[36029]_ ;
  assign \new_[36039]_  = A267 & ~A266;
  assign \new_[36040]_  = A265 & \new_[36039]_ ;
  assign \new_[36044]_  = A301 & ~A300;
  assign \new_[36045]_  = A268 & \new_[36044]_ ;
  assign \new_[36046]_  = \new_[36045]_  & \new_[36040]_ ;
  assign \new_[36050]_  = ~A167 & A168;
  assign \new_[36051]_  = A169 & \new_[36050]_ ;
  assign \new_[36055]_  = A202 & ~A201;
  assign \new_[36056]_  = A166 & \new_[36055]_ ;
  assign \new_[36057]_  = \new_[36056]_  & \new_[36051]_ ;
  assign \new_[36061]_  = A267 & ~A266;
  assign \new_[36062]_  = A265 & \new_[36061]_ ;
  assign \new_[36066]_  = ~A302 & ~A300;
  assign \new_[36067]_  = A268 & \new_[36066]_ ;
  assign \new_[36068]_  = \new_[36067]_  & \new_[36062]_ ;
  assign \new_[36072]_  = ~A167 & A168;
  assign \new_[36073]_  = A169 & \new_[36072]_ ;
  assign \new_[36077]_  = A202 & ~A201;
  assign \new_[36078]_  = A166 & \new_[36077]_ ;
  assign \new_[36079]_  = \new_[36078]_  & \new_[36073]_ ;
  assign \new_[36083]_  = A267 & ~A266;
  assign \new_[36084]_  = A265 & \new_[36083]_ ;
  assign \new_[36088]_  = A299 & A298;
  assign \new_[36089]_  = A268 & \new_[36088]_ ;
  assign \new_[36090]_  = \new_[36089]_  & \new_[36084]_ ;
  assign \new_[36094]_  = ~A167 & A168;
  assign \new_[36095]_  = A169 & \new_[36094]_ ;
  assign \new_[36099]_  = A202 & ~A201;
  assign \new_[36100]_  = A166 & \new_[36099]_ ;
  assign \new_[36101]_  = \new_[36100]_  & \new_[36095]_ ;
  assign \new_[36105]_  = A267 & ~A266;
  assign \new_[36106]_  = A265 & \new_[36105]_ ;
  assign \new_[36110]_  = ~A299 & ~A298;
  assign \new_[36111]_  = A268 & \new_[36110]_ ;
  assign \new_[36112]_  = \new_[36111]_  & \new_[36106]_ ;
  assign \new_[36116]_  = ~A167 & A168;
  assign \new_[36117]_  = A169 & \new_[36116]_ ;
  assign \new_[36121]_  = A202 & ~A201;
  assign \new_[36122]_  = A166 & \new_[36121]_ ;
  assign \new_[36123]_  = \new_[36122]_  & \new_[36117]_ ;
  assign \new_[36127]_  = A267 & ~A266;
  assign \new_[36128]_  = A265 & \new_[36127]_ ;
  assign \new_[36132]_  = A301 & ~A300;
  assign \new_[36133]_  = ~A269 & \new_[36132]_ ;
  assign \new_[36134]_  = \new_[36133]_  & \new_[36128]_ ;
  assign \new_[36138]_  = ~A167 & A168;
  assign \new_[36139]_  = A169 & \new_[36138]_ ;
  assign \new_[36143]_  = A202 & ~A201;
  assign \new_[36144]_  = A166 & \new_[36143]_ ;
  assign \new_[36145]_  = \new_[36144]_  & \new_[36139]_ ;
  assign \new_[36149]_  = A267 & ~A266;
  assign \new_[36150]_  = A265 & \new_[36149]_ ;
  assign \new_[36154]_  = ~A302 & ~A300;
  assign \new_[36155]_  = ~A269 & \new_[36154]_ ;
  assign \new_[36156]_  = \new_[36155]_  & \new_[36150]_ ;
  assign \new_[36160]_  = ~A167 & A168;
  assign \new_[36161]_  = A169 & \new_[36160]_ ;
  assign \new_[36165]_  = A202 & ~A201;
  assign \new_[36166]_  = A166 & \new_[36165]_ ;
  assign \new_[36167]_  = \new_[36166]_  & \new_[36161]_ ;
  assign \new_[36171]_  = A267 & ~A266;
  assign \new_[36172]_  = A265 & \new_[36171]_ ;
  assign \new_[36176]_  = A299 & A298;
  assign \new_[36177]_  = ~A269 & \new_[36176]_ ;
  assign \new_[36178]_  = \new_[36177]_  & \new_[36172]_ ;
  assign \new_[36182]_  = ~A167 & A168;
  assign \new_[36183]_  = A169 & \new_[36182]_ ;
  assign \new_[36187]_  = A202 & ~A201;
  assign \new_[36188]_  = A166 & \new_[36187]_ ;
  assign \new_[36189]_  = \new_[36188]_  & \new_[36183]_ ;
  assign \new_[36193]_  = A267 & ~A266;
  assign \new_[36194]_  = A265 & \new_[36193]_ ;
  assign \new_[36198]_  = ~A299 & ~A298;
  assign \new_[36199]_  = ~A269 & \new_[36198]_ ;
  assign \new_[36200]_  = \new_[36199]_  & \new_[36194]_ ;
  assign \new_[36204]_  = ~A167 & A168;
  assign \new_[36205]_  = A169 & \new_[36204]_ ;
  assign \new_[36209]_  = A202 & ~A201;
  assign \new_[36210]_  = A166 & \new_[36209]_ ;
  assign \new_[36211]_  = \new_[36210]_  & \new_[36205]_ ;
  assign \new_[36215]_  = A298 & ~A266;
  assign \new_[36216]_  = ~A265 & \new_[36215]_ ;
  assign \new_[36220]_  = A301 & A300;
  assign \new_[36221]_  = ~A299 & \new_[36220]_ ;
  assign \new_[36222]_  = \new_[36221]_  & \new_[36216]_ ;
  assign \new_[36226]_  = ~A167 & A168;
  assign \new_[36227]_  = A169 & \new_[36226]_ ;
  assign \new_[36231]_  = A202 & ~A201;
  assign \new_[36232]_  = A166 & \new_[36231]_ ;
  assign \new_[36233]_  = \new_[36232]_  & \new_[36227]_ ;
  assign \new_[36237]_  = A298 & ~A266;
  assign \new_[36238]_  = ~A265 & \new_[36237]_ ;
  assign \new_[36242]_  = ~A302 & A300;
  assign \new_[36243]_  = ~A299 & \new_[36242]_ ;
  assign \new_[36244]_  = \new_[36243]_  & \new_[36238]_ ;
  assign \new_[36248]_  = ~A167 & A168;
  assign \new_[36249]_  = A169 & \new_[36248]_ ;
  assign \new_[36253]_  = A202 & ~A201;
  assign \new_[36254]_  = A166 & \new_[36253]_ ;
  assign \new_[36255]_  = \new_[36254]_  & \new_[36249]_ ;
  assign \new_[36259]_  = ~A298 & ~A266;
  assign \new_[36260]_  = ~A265 & \new_[36259]_ ;
  assign \new_[36264]_  = A301 & A300;
  assign \new_[36265]_  = A299 & \new_[36264]_ ;
  assign \new_[36266]_  = \new_[36265]_  & \new_[36260]_ ;
  assign \new_[36270]_  = ~A167 & A168;
  assign \new_[36271]_  = A169 & \new_[36270]_ ;
  assign \new_[36275]_  = A202 & ~A201;
  assign \new_[36276]_  = A166 & \new_[36275]_ ;
  assign \new_[36277]_  = \new_[36276]_  & \new_[36271]_ ;
  assign \new_[36281]_  = ~A298 & ~A266;
  assign \new_[36282]_  = ~A265 & \new_[36281]_ ;
  assign \new_[36286]_  = ~A302 & A300;
  assign \new_[36287]_  = A299 & \new_[36286]_ ;
  assign \new_[36288]_  = \new_[36287]_  & \new_[36282]_ ;
  assign \new_[36292]_  = ~A167 & A168;
  assign \new_[36293]_  = A169 & \new_[36292]_ ;
  assign \new_[36297]_  = ~A203 & ~A201;
  assign \new_[36298]_  = A166 & \new_[36297]_ ;
  assign \new_[36299]_  = \new_[36298]_  & \new_[36293]_ ;
  assign \new_[36303]_  = A298 & A268;
  assign \new_[36304]_  = ~A267 & \new_[36303]_ ;
  assign \new_[36308]_  = A301 & A300;
  assign \new_[36309]_  = ~A299 & \new_[36308]_ ;
  assign \new_[36310]_  = \new_[36309]_  & \new_[36304]_ ;
  assign \new_[36314]_  = ~A167 & A168;
  assign \new_[36315]_  = A169 & \new_[36314]_ ;
  assign \new_[36319]_  = ~A203 & ~A201;
  assign \new_[36320]_  = A166 & \new_[36319]_ ;
  assign \new_[36321]_  = \new_[36320]_  & \new_[36315]_ ;
  assign \new_[36325]_  = A298 & A268;
  assign \new_[36326]_  = ~A267 & \new_[36325]_ ;
  assign \new_[36330]_  = ~A302 & A300;
  assign \new_[36331]_  = ~A299 & \new_[36330]_ ;
  assign \new_[36332]_  = \new_[36331]_  & \new_[36326]_ ;
  assign \new_[36336]_  = ~A167 & A168;
  assign \new_[36337]_  = A169 & \new_[36336]_ ;
  assign \new_[36341]_  = ~A203 & ~A201;
  assign \new_[36342]_  = A166 & \new_[36341]_ ;
  assign \new_[36343]_  = \new_[36342]_  & \new_[36337]_ ;
  assign \new_[36347]_  = ~A298 & A268;
  assign \new_[36348]_  = ~A267 & \new_[36347]_ ;
  assign \new_[36352]_  = A301 & A300;
  assign \new_[36353]_  = A299 & \new_[36352]_ ;
  assign \new_[36354]_  = \new_[36353]_  & \new_[36348]_ ;
  assign \new_[36358]_  = ~A167 & A168;
  assign \new_[36359]_  = A169 & \new_[36358]_ ;
  assign \new_[36363]_  = ~A203 & ~A201;
  assign \new_[36364]_  = A166 & \new_[36363]_ ;
  assign \new_[36365]_  = \new_[36364]_  & \new_[36359]_ ;
  assign \new_[36369]_  = ~A298 & A268;
  assign \new_[36370]_  = ~A267 & \new_[36369]_ ;
  assign \new_[36374]_  = ~A302 & A300;
  assign \new_[36375]_  = A299 & \new_[36374]_ ;
  assign \new_[36376]_  = \new_[36375]_  & \new_[36370]_ ;
  assign \new_[36380]_  = ~A167 & A168;
  assign \new_[36381]_  = A169 & \new_[36380]_ ;
  assign \new_[36385]_  = ~A203 & ~A201;
  assign \new_[36386]_  = A166 & \new_[36385]_ ;
  assign \new_[36387]_  = \new_[36386]_  & \new_[36381]_ ;
  assign \new_[36391]_  = A298 & ~A269;
  assign \new_[36392]_  = ~A267 & \new_[36391]_ ;
  assign \new_[36396]_  = A301 & A300;
  assign \new_[36397]_  = ~A299 & \new_[36396]_ ;
  assign \new_[36398]_  = \new_[36397]_  & \new_[36392]_ ;
  assign \new_[36402]_  = ~A167 & A168;
  assign \new_[36403]_  = A169 & \new_[36402]_ ;
  assign \new_[36407]_  = ~A203 & ~A201;
  assign \new_[36408]_  = A166 & \new_[36407]_ ;
  assign \new_[36409]_  = \new_[36408]_  & \new_[36403]_ ;
  assign \new_[36413]_  = A298 & ~A269;
  assign \new_[36414]_  = ~A267 & \new_[36413]_ ;
  assign \new_[36418]_  = ~A302 & A300;
  assign \new_[36419]_  = ~A299 & \new_[36418]_ ;
  assign \new_[36420]_  = \new_[36419]_  & \new_[36414]_ ;
  assign \new_[36424]_  = ~A167 & A168;
  assign \new_[36425]_  = A169 & \new_[36424]_ ;
  assign \new_[36429]_  = ~A203 & ~A201;
  assign \new_[36430]_  = A166 & \new_[36429]_ ;
  assign \new_[36431]_  = \new_[36430]_  & \new_[36425]_ ;
  assign \new_[36435]_  = ~A298 & ~A269;
  assign \new_[36436]_  = ~A267 & \new_[36435]_ ;
  assign \new_[36440]_  = A301 & A300;
  assign \new_[36441]_  = A299 & \new_[36440]_ ;
  assign \new_[36442]_  = \new_[36441]_  & \new_[36436]_ ;
  assign \new_[36446]_  = ~A167 & A168;
  assign \new_[36447]_  = A169 & \new_[36446]_ ;
  assign \new_[36451]_  = ~A203 & ~A201;
  assign \new_[36452]_  = A166 & \new_[36451]_ ;
  assign \new_[36453]_  = \new_[36452]_  & \new_[36447]_ ;
  assign \new_[36457]_  = ~A298 & ~A269;
  assign \new_[36458]_  = ~A267 & \new_[36457]_ ;
  assign \new_[36462]_  = ~A302 & A300;
  assign \new_[36463]_  = A299 & \new_[36462]_ ;
  assign \new_[36464]_  = \new_[36463]_  & \new_[36458]_ ;
  assign \new_[36468]_  = ~A167 & A168;
  assign \new_[36469]_  = A169 & \new_[36468]_ ;
  assign \new_[36473]_  = ~A203 & ~A201;
  assign \new_[36474]_  = A166 & \new_[36473]_ ;
  assign \new_[36475]_  = \new_[36474]_  & \new_[36469]_ ;
  assign \new_[36479]_  = A298 & A266;
  assign \new_[36480]_  = A265 & \new_[36479]_ ;
  assign \new_[36484]_  = A301 & A300;
  assign \new_[36485]_  = ~A299 & \new_[36484]_ ;
  assign \new_[36486]_  = \new_[36485]_  & \new_[36480]_ ;
  assign \new_[36490]_  = ~A167 & A168;
  assign \new_[36491]_  = A169 & \new_[36490]_ ;
  assign \new_[36495]_  = ~A203 & ~A201;
  assign \new_[36496]_  = A166 & \new_[36495]_ ;
  assign \new_[36497]_  = \new_[36496]_  & \new_[36491]_ ;
  assign \new_[36501]_  = A298 & A266;
  assign \new_[36502]_  = A265 & \new_[36501]_ ;
  assign \new_[36506]_  = ~A302 & A300;
  assign \new_[36507]_  = ~A299 & \new_[36506]_ ;
  assign \new_[36508]_  = \new_[36507]_  & \new_[36502]_ ;
  assign \new_[36512]_  = ~A167 & A168;
  assign \new_[36513]_  = A169 & \new_[36512]_ ;
  assign \new_[36517]_  = ~A203 & ~A201;
  assign \new_[36518]_  = A166 & \new_[36517]_ ;
  assign \new_[36519]_  = \new_[36518]_  & \new_[36513]_ ;
  assign \new_[36523]_  = ~A298 & A266;
  assign \new_[36524]_  = A265 & \new_[36523]_ ;
  assign \new_[36528]_  = A301 & A300;
  assign \new_[36529]_  = A299 & \new_[36528]_ ;
  assign \new_[36530]_  = \new_[36529]_  & \new_[36524]_ ;
  assign \new_[36534]_  = ~A167 & A168;
  assign \new_[36535]_  = A169 & \new_[36534]_ ;
  assign \new_[36539]_  = ~A203 & ~A201;
  assign \new_[36540]_  = A166 & \new_[36539]_ ;
  assign \new_[36541]_  = \new_[36540]_  & \new_[36535]_ ;
  assign \new_[36545]_  = ~A298 & A266;
  assign \new_[36546]_  = A265 & \new_[36545]_ ;
  assign \new_[36550]_  = ~A302 & A300;
  assign \new_[36551]_  = A299 & \new_[36550]_ ;
  assign \new_[36552]_  = \new_[36551]_  & \new_[36546]_ ;
  assign \new_[36556]_  = ~A167 & A168;
  assign \new_[36557]_  = A169 & \new_[36556]_ ;
  assign \new_[36561]_  = ~A203 & ~A201;
  assign \new_[36562]_  = A166 & \new_[36561]_ ;
  assign \new_[36563]_  = \new_[36562]_  & \new_[36557]_ ;
  assign \new_[36567]_  = A267 & A266;
  assign \new_[36568]_  = ~A265 & \new_[36567]_ ;
  assign \new_[36572]_  = A301 & ~A300;
  assign \new_[36573]_  = A268 & \new_[36572]_ ;
  assign \new_[36574]_  = \new_[36573]_  & \new_[36568]_ ;
  assign \new_[36578]_  = ~A167 & A168;
  assign \new_[36579]_  = A169 & \new_[36578]_ ;
  assign \new_[36583]_  = ~A203 & ~A201;
  assign \new_[36584]_  = A166 & \new_[36583]_ ;
  assign \new_[36585]_  = \new_[36584]_  & \new_[36579]_ ;
  assign \new_[36589]_  = A267 & A266;
  assign \new_[36590]_  = ~A265 & \new_[36589]_ ;
  assign \new_[36594]_  = ~A302 & ~A300;
  assign \new_[36595]_  = A268 & \new_[36594]_ ;
  assign \new_[36596]_  = \new_[36595]_  & \new_[36590]_ ;
  assign \new_[36600]_  = ~A167 & A168;
  assign \new_[36601]_  = A169 & \new_[36600]_ ;
  assign \new_[36605]_  = ~A203 & ~A201;
  assign \new_[36606]_  = A166 & \new_[36605]_ ;
  assign \new_[36607]_  = \new_[36606]_  & \new_[36601]_ ;
  assign \new_[36611]_  = A267 & A266;
  assign \new_[36612]_  = ~A265 & \new_[36611]_ ;
  assign \new_[36616]_  = A299 & A298;
  assign \new_[36617]_  = A268 & \new_[36616]_ ;
  assign \new_[36618]_  = \new_[36617]_  & \new_[36612]_ ;
  assign \new_[36622]_  = ~A167 & A168;
  assign \new_[36623]_  = A169 & \new_[36622]_ ;
  assign \new_[36627]_  = ~A203 & ~A201;
  assign \new_[36628]_  = A166 & \new_[36627]_ ;
  assign \new_[36629]_  = \new_[36628]_  & \new_[36623]_ ;
  assign \new_[36633]_  = A267 & A266;
  assign \new_[36634]_  = ~A265 & \new_[36633]_ ;
  assign \new_[36638]_  = ~A299 & ~A298;
  assign \new_[36639]_  = A268 & \new_[36638]_ ;
  assign \new_[36640]_  = \new_[36639]_  & \new_[36634]_ ;
  assign \new_[36644]_  = ~A167 & A168;
  assign \new_[36645]_  = A169 & \new_[36644]_ ;
  assign \new_[36649]_  = ~A203 & ~A201;
  assign \new_[36650]_  = A166 & \new_[36649]_ ;
  assign \new_[36651]_  = \new_[36650]_  & \new_[36645]_ ;
  assign \new_[36655]_  = A267 & A266;
  assign \new_[36656]_  = ~A265 & \new_[36655]_ ;
  assign \new_[36660]_  = A301 & ~A300;
  assign \new_[36661]_  = ~A269 & \new_[36660]_ ;
  assign \new_[36662]_  = \new_[36661]_  & \new_[36656]_ ;
  assign \new_[36666]_  = ~A167 & A168;
  assign \new_[36667]_  = A169 & \new_[36666]_ ;
  assign \new_[36671]_  = ~A203 & ~A201;
  assign \new_[36672]_  = A166 & \new_[36671]_ ;
  assign \new_[36673]_  = \new_[36672]_  & \new_[36667]_ ;
  assign \new_[36677]_  = A267 & A266;
  assign \new_[36678]_  = ~A265 & \new_[36677]_ ;
  assign \new_[36682]_  = ~A302 & ~A300;
  assign \new_[36683]_  = ~A269 & \new_[36682]_ ;
  assign \new_[36684]_  = \new_[36683]_  & \new_[36678]_ ;
  assign \new_[36688]_  = ~A167 & A168;
  assign \new_[36689]_  = A169 & \new_[36688]_ ;
  assign \new_[36693]_  = ~A203 & ~A201;
  assign \new_[36694]_  = A166 & \new_[36693]_ ;
  assign \new_[36695]_  = \new_[36694]_  & \new_[36689]_ ;
  assign \new_[36699]_  = A267 & A266;
  assign \new_[36700]_  = ~A265 & \new_[36699]_ ;
  assign \new_[36704]_  = A299 & A298;
  assign \new_[36705]_  = ~A269 & \new_[36704]_ ;
  assign \new_[36706]_  = \new_[36705]_  & \new_[36700]_ ;
  assign \new_[36710]_  = ~A167 & A168;
  assign \new_[36711]_  = A169 & \new_[36710]_ ;
  assign \new_[36715]_  = ~A203 & ~A201;
  assign \new_[36716]_  = A166 & \new_[36715]_ ;
  assign \new_[36717]_  = \new_[36716]_  & \new_[36711]_ ;
  assign \new_[36721]_  = A267 & A266;
  assign \new_[36722]_  = ~A265 & \new_[36721]_ ;
  assign \new_[36726]_  = ~A299 & ~A298;
  assign \new_[36727]_  = ~A269 & \new_[36726]_ ;
  assign \new_[36728]_  = \new_[36727]_  & \new_[36722]_ ;
  assign \new_[36732]_  = ~A167 & A168;
  assign \new_[36733]_  = A169 & \new_[36732]_ ;
  assign \new_[36737]_  = ~A203 & ~A201;
  assign \new_[36738]_  = A166 & \new_[36737]_ ;
  assign \new_[36739]_  = \new_[36738]_  & \new_[36733]_ ;
  assign \new_[36743]_  = A267 & ~A266;
  assign \new_[36744]_  = A265 & \new_[36743]_ ;
  assign \new_[36748]_  = A301 & ~A300;
  assign \new_[36749]_  = A268 & \new_[36748]_ ;
  assign \new_[36750]_  = \new_[36749]_  & \new_[36744]_ ;
  assign \new_[36754]_  = ~A167 & A168;
  assign \new_[36755]_  = A169 & \new_[36754]_ ;
  assign \new_[36759]_  = ~A203 & ~A201;
  assign \new_[36760]_  = A166 & \new_[36759]_ ;
  assign \new_[36761]_  = \new_[36760]_  & \new_[36755]_ ;
  assign \new_[36765]_  = A267 & ~A266;
  assign \new_[36766]_  = A265 & \new_[36765]_ ;
  assign \new_[36770]_  = ~A302 & ~A300;
  assign \new_[36771]_  = A268 & \new_[36770]_ ;
  assign \new_[36772]_  = \new_[36771]_  & \new_[36766]_ ;
  assign \new_[36776]_  = ~A167 & A168;
  assign \new_[36777]_  = A169 & \new_[36776]_ ;
  assign \new_[36781]_  = ~A203 & ~A201;
  assign \new_[36782]_  = A166 & \new_[36781]_ ;
  assign \new_[36783]_  = \new_[36782]_  & \new_[36777]_ ;
  assign \new_[36787]_  = A267 & ~A266;
  assign \new_[36788]_  = A265 & \new_[36787]_ ;
  assign \new_[36792]_  = A299 & A298;
  assign \new_[36793]_  = A268 & \new_[36792]_ ;
  assign \new_[36794]_  = \new_[36793]_  & \new_[36788]_ ;
  assign \new_[36798]_  = ~A167 & A168;
  assign \new_[36799]_  = A169 & \new_[36798]_ ;
  assign \new_[36803]_  = ~A203 & ~A201;
  assign \new_[36804]_  = A166 & \new_[36803]_ ;
  assign \new_[36805]_  = \new_[36804]_  & \new_[36799]_ ;
  assign \new_[36809]_  = A267 & ~A266;
  assign \new_[36810]_  = A265 & \new_[36809]_ ;
  assign \new_[36814]_  = ~A299 & ~A298;
  assign \new_[36815]_  = A268 & \new_[36814]_ ;
  assign \new_[36816]_  = \new_[36815]_  & \new_[36810]_ ;
  assign \new_[36820]_  = ~A167 & A168;
  assign \new_[36821]_  = A169 & \new_[36820]_ ;
  assign \new_[36825]_  = ~A203 & ~A201;
  assign \new_[36826]_  = A166 & \new_[36825]_ ;
  assign \new_[36827]_  = \new_[36826]_  & \new_[36821]_ ;
  assign \new_[36831]_  = A267 & ~A266;
  assign \new_[36832]_  = A265 & \new_[36831]_ ;
  assign \new_[36836]_  = A301 & ~A300;
  assign \new_[36837]_  = ~A269 & \new_[36836]_ ;
  assign \new_[36838]_  = \new_[36837]_  & \new_[36832]_ ;
  assign \new_[36842]_  = ~A167 & A168;
  assign \new_[36843]_  = A169 & \new_[36842]_ ;
  assign \new_[36847]_  = ~A203 & ~A201;
  assign \new_[36848]_  = A166 & \new_[36847]_ ;
  assign \new_[36849]_  = \new_[36848]_  & \new_[36843]_ ;
  assign \new_[36853]_  = A267 & ~A266;
  assign \new_[36854]_  = A265 & \new_[36853]_ ;
  assign \new_[36858]_  = ~A302 & ~A300;
  assign \new_[36859]_  = ~A269 & \new_[36858]_ ;
  assign \new_[36860]_  = \new_[36859]_  & \new_[36854]_ ;
  assign \new_[36864]_  = ~A167 & A168;
  assign \new_[36865]_  = A169 & \new_[36864]_ ;
  assign \new_[36869]_  = ~A203 & ~A201;
  assign \new_[36870]_  = A166 & \new_[36869]_ ;
  assign \new_[36871]_  = \new_[36870]_  & \new_[36865]_ ;
  assign \new_[36875]_  = A267 & ~A266;
  assign \new_[36876]_  = A265 & \new_[36875]_ ;
  assign \new_[36880]_  = A299 & A298;
  assign \new_[36881]_  = ~A269 & \new_[36880]_ ;
  assign \new_[36882]_  = \new_[36881]_  & \new_[36876]_ ;
  assign \new_[36886]_  = ~A167 & A168;
  assign \new_[36887]_  = A169 & \new_[36886]_ ;
  assign \new_[36891]_  = ~A203 & ~A201;
  assign \new_[36892]_  = A166 & \new_[36891]_ ;
  assign \new_[36893]_  = \new_[36892]_  & \new_[36887]_ ;
  assign \new_[36897]_  = A267 & ~A266;
  assign \new_[36898]_  = A265 & \new_[36897]_ ;
  assign \new_[36902]_  = ~A299 & ~A298;
  assign \new_[36903]_  = ~A269 & \new_[36902]_ ;
  assign \new_[36904]_  = \new_[36903]_  & \new_[36898]_ ;
  assign \new_[36908]_  = ~A167 & A168;
  assign \new_[36909]_  = A169 & \new_[36908]_ ;
  assign \new_[36913]_  = ~A203 & ~A201;
  assign \new_[36914]_  = A166 & \new_[36913]_ ;
  assign \new_[36915]_  = \new_[36914]_  & \new_[36909]_ ;
  assign \new_[36919]_  = A298 & ~A266;
  assign \new_[36920]_  = ~A265 & \new_[36919]_ ;
  assign \new_[36924]_  = A301 & A300;
  assign \new_[36925]_  = ~A299 & \new_[36924]_ ;
  assign \new_[36926]_  = \new_[36925]_  & \new_[36920]_ ;
  assign \new_[36930]_  = ~A167 & A168;
  assign \new_[36931]_  = A169 & \new_[36930]_ ;
  assign \new_[36935]_  = ~A203 & ~A201;
  assign \new_[36936]_  = A166 & \new_[36935]_ ;
  assign \new_[36937]_  = \new_[36936]_  & \new_[36931]_ ;
  assign \new_[36941]_  = A298 & ~A266;
  assign \new_[36942]_  = ~A265 & \new_[36941]_ ;
  assign \new_[36946]_  = ~A302 & A300;
  assign \new_[36947]_  = ~A299 & \new_[36946]_ ;
  assign \new_[36948]_  = \new_[36947]_  & \new_[36942]_ ;
  assign \new_[36952]_  = ~A167 & A168;
  assign \new_[36953]_  = A169 & \new_[36952]_ ;
  assign \new_[36957]_  = ~A203 & ~A201;
  assign \new_[36958]_  = A166 & \new_[36957]_ ;
  assign \new_[36959]_  = \new_[36958]_  & \new_[36953]_ ;
  assign \new_[36963]_  = ~A298 & ~A266;
  assign \new_[36964]_  = ~A265 & \new_[36963]_ ;
  assign \new_[36968]_  = A301 & A300;
  assign \new_[36969]_  = A299 & \new_[36968]_ ;
  assign \new_[36970]_  = \new_[36969]_  & \new_[36964]_ ;
  assign \new_[36974]_  = ~A167 & A168;
  assign \new_[36975]_  = A169 & \new_[36974]_ ;
  assign \new_[36979]_  = ~A203 & ~A201;
  assign \new_[36980]_  = A166 & \new_[36979]_ ;
  assign \new_[36981]_  = \new_[36980]_  & \new_[36975]_ ;
  assign \new_[36985]_  = ~A298 & ~A266;
  assign \new_[36986]_  = ~A265 & \new_[36985]_ ;
  assign \new_[36990]_  = ~A302 & A300;
  assign \new_[36991]_  = A299 & \new_[36990]_ ;
  assign \new_[36992]_  = \new_[36991]_  & \new_[36986]_ ;
  assign \new_[36996]_  = ~A167 & A168;
  assign \new_[36997]_  = A169 & \new_[36996]_ ;
  assign \new_[37001]_  = A200 & A199;
  assign \new_[37002]_  = A166 & \new_[37001]_ ;
  assign \new_[37003]_  = \new_[37002]_  & \new_[36997]_ ;
  assign \new_[37007]_  = A298 & A268;
  assign \new_[37008]_  = ~A267 & \new_[37007]_ ;
  assign \new_[37012]_  = A301 & A300;
  assign \new_[37013]_  = ~A299 & \new_[37012]_ ;
  assign \new_[37014]_  = \new_[37013]_  & \new_[37008]_ ;
  assign \new_[37018]_  = ~A167 & A168;
  assign \new_[37019]_  = A169 & \new_[37018]_ ;
  assign \new_[37023]_  = A200 & A199;
  assign \new_[37024]_  = A166 & \new_[37023]_ ;
  assign \new_[37025]_  = \new_[37024]_  & \new_[37019]_ ;
  assign \new_[37029]_  = A298 & A268;
  assign \new_[37030]_  = ~A267 & \new_[37029]_ ;
  assign \new_[37034]_  = ~A302 & A300;
  assign \new_[37035]_  = ~A299 & \new_[37034]_ ;
  assign \new_[37036]_  = \new_[37035]_  & \new_[37030]_ ;
  assign \new_[37040]_  = ~A167 & A168;
  assign \new_[37041]_  = A169 & \new_[37040]_ ;
  assign \new_[37045]_  = A200 & A199;
  assign \new_[37046]_  = A166 & \new_[37045]_ ;
  assign \new_[37047]_  = \new_[37046]_  & \new_[37041]_ ;
  assign \new_[37051]_  = ~A298 & A268;
  assign \new_[37052]_  = ~A267 & \new_[37051]_ ;
  assign \new_[37056]_  = A301 & A300;
  assign \new_[37057]_  = A299 & \new_[37056]_ ;
  assign \new_[37058]_  = \new_[37057]_  & \new_[37052]_ ;
  assign \new_[37062]_  = ~A167 & A168;
  assign \new_[37063]_  = A169 & \new_[37062]_ ;
  assign \new_[37067]_  = A200 & A199;
  assign \new_[37068]_  = A166 & \new_[37067]_ ;
  assign \new_[37069]_  = \new_[37068]_  & \new_[37063]_ ;
  assign \new_[37073]_  = ~A298 & A268;
  assign \new_[37074]_  = ~A267 & \new_[37073]_ ;
  assign \new_[37078]_  = ~A302 & A300;
  assign \new_[37079]_  = A299 & \new_[37078]_ ;
  assign \new_[37080]_  = \new_[37079]_  & \new_[37074]_ ;
  assign \new_[37084]_  = ~A167 & A168;
  assign \new_[37085]_  = A169 & \new_[37084]_ ;
  assign \new_[37089]_  = A200 & A199;
  assign \new_[37090]_  = A166 & \new_[37089]_ ;
  assign \new_[37091]_  = \new_[37090]_  & \new_[37085]_ ;
  assign \new_[37095]_  = A298 & ~A269;
  assign \new_[37096]_  = ~A267 & \new_[37095]_ ;
  assign \new_[37100]_  = A301 & A300;
  assign \new_[37101]_  = ~A299 & \new_[37100]_ ;
  assign \new_[37102]_  = \new_[37101]_  & \new_[37096]_ ;
  assign \new_[37106]_  = ~A167 & A168;
  assign \new_[37107]_  = A169 & \new_[37106]_ ;
  assign \new_[37111]_  = A200 & A199;
  assign \new_[37112]_  = A166 & \new_[37111]_ ;
  assign \new_[37113]_  = \new_[37112]_  & \new_[37107]_ ;
  assign \new_[37117]_  = A298 & ~A269;
  assign \new_[37118]_  = ~A267 & \new_[37117]_ ;
  assign \new_[37122]_  = ~A302 & A300;
  assign \new_[37123]_  = ~A299 & \new_[37122]_ ;
  assign \new_[37124]_  = \new_[37123]_  & \new_[37118]_ ;
  assign \new_[37128]_  = ~A167 & A168;
  assign \new_[37129]_  = A169 & \new_[37128]_ ;
  assign \new_[37133]_  = A200 & A199;
  assign \new_[37134]_  = A166 & \new_[37133]_ ;
  assign \new_[37135]_  = \new_[37134]_  & \new_[37129]_ ;
  assign \new_[37139]_  = ~A298 & ~A269;
  assign \new_[37140]_  = ~A267 & \new_[37139]_ ;
  assign \new_[37144]_  = A301 & A300;
  assign \new_[37145]_  = A299 & \new_[37144]_ ;
  assign \new_[37146]_  = \new_[37145]_  & \new_[37140]_ ;
  assign \new_[37150]_  = ~A167 & A168;
  assign \new_[37151]_  = A169 & \new_[37150]_ ;
  assign \new_[37155]_  = A200 & A199;
  assign \new_[37156]_  = A166 & \new_[37155]_ ;
  assign \new_[37157]_  = \new_[37156]_  & \new_[37151]_ ;
  assign \new_[37161]_  = ~A298 & ~A269;
  assign \new_[37162]_  = ~A267 & \new_[37161]_ ;
  assign \new_[37166]_  = ~A302 & A300;
  assign \new_[37167]_  = A299 & \new_[37166]_ ;
  assign \new_[37168]_  = \new_[37167]_  & \new_[37162]_ ;
  assign \new_[37172]_  = ~A167 & A168;
  assign \new_[37173]_  = A169 & \new_[37172]_ ;
  assign \new_[37177]_  = A200 & A199;
  assign \new_[37178]_  = A166 & \new_[37177]_ ;
  assign \new_[37179]_  = \new_[37178]_  & \new_[37173]_ ;
  assign \new_[37183]_  = A298 & A266;
  assign \new_[37184]_  = A265 & \new_[37183]_ ;
  assign \new_[37188]_  = A301 & A300;
  assign \new_[37189]_  = ~A299 & \new_[37188]_ ;
  assign \new_[37190]_  = \new_[37189]_  & \new_[37184]_ ;
  assign \new_[37194]_  = ~A167 & A168;
  assign \new_[37195]_  = A169 & \new_[37194]_ ;
  assign \new_[37199]_  = A200 & A199;
  assign \new_[37200]_  = A166 & \new_[37199]_ ;
  assign \new_[37201]_  = \new_[37200]_  & \new_[37195]_ ;
  assign \new_[37205]_  = A298 & A266;
  assign \new_[37206]_  = A265 & \new_[37205]_ ;
  assign \new_[37210]_  = ~A302 & A300;
  assign \new_[37211]_  = ~A299 & \new_[37210]_ ;
  assign \new_[37212]_  = \new_[37211]_  & \new_[37206]_ ;
  assign \new_[37216]_  = ~A167 & A168;
  assign \new_[37217]_  = A169 & \new_[37216]_ ;
  assign \new_[37221]_  = A200 & A199;
  assign \new_[37222]_  = A166 & \new_[37221]_ ;
  assign \new_[37223]_  = \new_[37222]_  & \new_[37217]_ ;
  assign \new_[37227]_  = ~A298 & A266;
  assign \new_[37228]_  = A265 & \new_[37227]_ ;
  assign \new_[37232]_  = A301 & A300;
  assign \new_[37233]_  = A299 & \new_[37232]_ ;
  assign \new_[37234]_  = \new_[37233]_  & \new_[37228]_ ;
  assign \new_[37238]_  = ~A167 & A168;
  assign \new_[37239]_  = A169 & \new_[37238]_ ;
  assign \new_[37243]_  = A200 & A199;
  assign \new_[37244]_  = A166 & \new_[37243]_ ;
  assign \new_[37245]_  = \new_[37244]_  & \new_[37239]_ ;
  assign \new_[37249]_  = ~A298 & A266;
  assign \new_[37250]_  = A265 & \new_[37249]_ ;
  assign \new_[37254]_  = ~A302 & A300;
  assign \new_[37255]_  = A299 & \new_[37254]_ ;
  assign \new_[37256]_  = \new_[37255]_  & \new_[37250]_ ;
  assign \new_[37260]_  = ~A167 & A168;
  assign \new_[37261]_  = A169 & \new_[37260]_ ;
  assign \new_[37265]_  = A200 & A199;
  assign \new_[37266]_  = A166 & \new_[37265]_ ;
  assign \new_[37267]_  = \new_[37266]_  & \new_[37261]_ ;
  assign \new_[37271]_  = A267 & A266;
  assign \new_[37272]_  = ~A265 & \new_[37271]_ ;
  assign \new_[37276]_  = A301 & ~A300;
  assign \new_[37277]_  = A268 & \new_[37276]_ ;
  assign \new_[37278]_  = \new_[37277]_  & \new_[37272]_ ;
  assign \new_[37282]_  = ~A167 & A168;
  assign \new_[37283]_  = A169 & \new_[37282]_ ;
  assign \new_[37287]_  = A200 & A199;
  assign \new_[37288]_  = A166 & \new_[37287]_ ;
  assign \new_[37289]_  = \new_[37288]_  & \new_[37283]_ ;
  assign \new_[37293]_  = A267 & A266;
  assign \new_[37294]_  = ~A265 & \new_[37293]_ ;
  assign \new_[37298]_  = ~A302 & ~A300;
  assign \new_[37299]_  = A268 & \new_[37298]_ ;
  assign \new_[37300]_  = \new_[37299]_  & \new_[37294]_ ;
  assign \new_[37304]_  = ~A167 & A168;
  assign \new_[37305]_  = A169 & \new_[37304]_ ;
  assign \new_[37309]_  = A200 & A199;
  assign \new_[37310]_  = A166 & \new_[37309]_ ;
  assign \new_[37311]_  = \new_[37310]_  & \new_[37305]_ ;
  assign \new_[37315]_  = A267 & A266;
  assign \new_[37316]_  = ~A265 & \new_[37315]_ ;
  assign \new_[37320]_  = A299 & A298;
  assign \new_[37321]_  = A268 & \new_[37320]_ ;
  assign \new_[37322]_  = \new_[37321]_  & \new_[37316]_ ;
  assign \new_[37326]_  = ~A167 & A168;
  assign \new_[37327]_  = A169 & \new_[37326]_ ;
  assign \new_[37331]_  = A200 & A199;
  assign \new_[37332]_  = A166 & \new_[37331]_ ;
  assign \new_[37333]_  = \new_[37332]_  & \new_[37327]_ ;
  assign \new_[37337]_  = A267 & A266;
  assign \new_[37338]_  = ~A265 & \new_[37337]_ ;
  assign \new_[37342]_  = ~A299 & ~A298;
  assign \new_[37343]_  = A268 & \new_[37342]_ ;
  assign \new_[37344]_  = \new_[37343]_  & \new_[37338]_ ;
  assign \new_[37348]_  = ~A167 & A168;
  assign \new_[37349]_  = A169 & \new_[37348]_ ;
  assign \new_[37353]_  = A200 & A199;
  assign \new_[37354]_  = A166 & \new_[37353]_ ;
  assign \new_[37355]_  = \new_[37354]_  & \new_[37349]_ ;
  assign \new_[37359]_  = A267 & A266;
  assign \new_[37360]_  = ~A265 & \new_[37359]_ ;
  assign \new_[37364]_  = A301 & ~A300;
  assign \new_[37365]_  = ~A269 & \new_[37364]_ ;
  assign \new_[37366]_  = \new_[37365]_  & \new_[37360]_ ;
  assign \new_[37370]_  = ~A167 & A168;
  assign \new_[37371]_  = A169 & \new_[37370]_ ;
  assign \new_[37375]_  = A200 & A199;
  assign \new_[37376]_  = A166 & \new_[37375]_ ;
  assign \new_[37377]_  = \new_[37376]_  & \new_[37371]_ ;
  assign \new_[37381]_  = A267 & A266;
  assign \new_[37382]_  = ~A265 & \new_[37381]_ ;
  assign \new_[37386]_  = ~A302 & ~A300;
  assign \new_[37387]_  = ~A269 & \new_[37386]_ ;
  assign \new_[37388]_  = \new_[37387]_  & \new_[37382]_ ;
  assign \new_[37392]_  = ~A167 & A168;
  assign \new_[37393]_  = A169 & \new_[37392]_ ;
  assign \new_[37397]_  = A200 & A199;
  assign \new_[37398]_  = A166 & \new_[37397]_ ;
  assign \new_[37399]_  = \new_[37398]_  & \new_[37393]_ ;
  assign \new_[37403]_  = A267 & A266;
  assign \new_[37404]_  = ~A265 & \new_[37403]_ ;
  assign \new_[37408]_  = A299 & A298;
  assign \new_[37409]_  = ~A269 & \new_[37408]_ ;
  assign \new_[37410]_  = \new_[37409]_  & \new_[37404]_ ;
  assign \new_[37414]_  = ~A167 & A168;
  assign \new_[37415]_  = A169 & \new_[37414]_ ;
  assign \new_[37419]_  = A200 & A199;
  assign \new_[37420]_  = A166 & \new_[37419]_ ;
  assign \new_[37421]_  = \new_[37420]_  & \new_[37415]_ ;
  assign \new_[37425]_  = A267 & A266;
  assign \new_[37426]_  = ~A265 & \new_[37425]_ ;
  assign \new_[37430]_  = ~A299 & ~A298;
  assign \new_[37431]_  = ~A269 & \new_[37430]_ ;
  assign \new_[37432]_  = \new_[37431]_  & \new_[37426]_ ;
  assign \new_[37436]_  = ~A167 & A168;
  assign \new_[37437]_  = A169 & \new_[37436]_ ;
  assign \new_[37441]_  = A200 & A199;
  assign \new_[37442]_  = A166 & \new_[37441]_ ;
  assign \new_[37443]_  = \new_[37442]_  & \new_[37437]_ ;
  assign \new_[37447]_  = A267 & ~A266;
  assign \new_[37448]_  = A265 & \new_[37447]_ ;
  assign \new_[37452]_  = A301 & ~A300;
  assign \new_[37453]_  = A268 & \new_[37452]_ ;
  assign \new_[37454]_  = \new_[37453]_  & \new_[37448]_ ;
  assign \new_[37458]_  = ~A167 & A168;
  assign \new_[37459]_  = A169 & \new_[37458]_ ;
  assign \new_[37463]_  = A200 & A199;
  assign \new_[37464]_  = A166 & \new_[37463]_ ;
  assign \new_[37465]_  = \new_[37464]_  & \new_[37459]_ ;
  assign \new_[37469]_  = A267 & ~A266;
  assign \new_[37470]_  = A265 & \new_[37469]_ ;
  assign \new_[37474]_  = ~A302 & ~A300;
  assign \new_[37475]_  = A268 & \new_[37474]_ ;
  assign \new_[37476]_  = \new_[37475]_  & \new_[37470]_ ;
  assign \new_[37480]_  = ~A167 & A168;
  assign \new_[37481]_  = A169 & \new_[37480]_ ;
  assign \new_[37485]_  = A200 & A199;
  assign \new_[37486]_  = A166 & \new_[37485]_ ;
  assign \new_[37487]_  = \new_[37486]_  & \new_[37481]_ ;
  assign \new_[37491]_  = A267 & ~A266;
  assign \new_[37492]_  = A265 & \new_[37491]_ ;
  assign \new_[37496]_  = A299 & A298;
  assign \new_[37497]_  = A268 & \new_[37496]_ ;
  assign \new_[37498]_  = \new_[37497]_  & \new_[37492]_ ;
  assign \new_[37502]_  = ~A167 & A168;
  assign \new_[37503]_  = A169 & \new_[37502]_ ;
  assign \new_[37507]_  = A200 & A199;
  assign \new_[37508]_  = A166 & \new_[37507]_ ;
  assign \new_[37509]_  = \new_[37508]_  & \new_[37503]_ ;
  assign \new_[37513]_  = A267 & ~A266;
  assign \new_[37514]_  = A265 & \new_[37513]_ ;
  assign \new_[37518]_  = ~A299 & ~A298;
  assign \new_[37519]_  = A268 & \new_[37518]_ ;
  assign \new_[37520]_  = \new_[37519]_  & \new_[37514]_ ;
  assign \new_[37524]_  = ~A167 & A168;
  assign \new_[37525]_  = A169 & \new_[37524]_ ;
  assign \new_[37529]_  = A200 & A199;
  assign \new_[37530]_  = A166 & \new_[37529]_ ;
  assign \new_[37531]_  = \new_[37530]_  & \new_[37525]_ ;
  assign \new_[37535]_  = A267 & ~A266;
  assign \new_[37536]_  = A265 & \new_[37535]_ ;
  assign \new_[37540]_  = A301 & ~A300;
  assign \new_[37541]_  = ~A269 & \new_[37540]_ ;
  assign \new_[37542]_  = \new_[37541]_  & \new_[37536]_ ;
  assign \new_[37546]_  = ~A167 & A168;
  assign \new_[37547]_  = A169 & \new_[37546]_ ;
  assign \new_[37551]_  = A200 & A199;
  assign \new_[37552]_  = A166 & \new_[37551]_ ;
  assign \new_[37553]_  = \new_[37552]_  & \new_[37547]_ ;
  assign \new_[37557]_  = A267 & ~A266;
  assign \new_[37558]_  = A265 & \new_[37557]_ ;
  assign \new_[37562]_  = ~A302 & ~A300;
  assign \new_[37563]_  = ~A269 & \new_[37562]_ ;
  assign \new_[37564]_  = \new_[37563]_  & \new_[37558]_ ;
  assign \new_[37568]_  = ~A167 & A168;
  assign \new_[37569]_  = A169 & \new_[37568]_ ;
  assign \new_[37573]_  = A200 & A199;
  assign \new_[37574]_  = A166 & \new_[37573]_ ;
  assign \new_[37575]_  = \new_[37574]_  & \new_[37569]_ ;
  assign \new_[37579]_  = A267 & ~A266;
  assign \new_[37580]_  = A265 & \new_[37579]_ ;
  assign \new_[37584]_  = A299 & A298;
  assign \new_[37585]_  = ~A269 & \new_[37584]_ ;
  assign \new_[37586]_  = \new_[37585]_  & \new_[37580]_ ;
  assign \new_[37590]_  = ~A167 & A168;
  assign \new_[37591]_  = A169 & \new_[37590]_ ;
  assign \new_[37595]_  = A200 & A199;
  assign \new_[37596]_  = A166 & \new_[37595]_ ;
  assign \new_[37597]_  = \new_[37596]_  & \new_[37591]_ ;
  assign \new_[37601]_  = A267 & ~A266;
  assign \new_[37602]_  = A265 & \new_[37601]_ ;
  assign \new_[37606]_  = ~A299 & ~A298;
  assign \new_[37607]_  = ~A269 & \new_[37606]_ ;
  assign \new_[37608]_  = \new_[37607]_  & \new_[37602]_ ;
  assign \new_[37612]_  = ~A167 & A168;
  assign \new_[37613]_  = A169 & \new_[37612]_ ;
  assign \new_[37617]_  = A200 & A199;
  assign \new_[37618]_  = A166 & \new_[37617]_ ;
  assign \new_[37619]_  = \new_[37618]_  & \new_[37613]_ ;
  assign \new_[37623]_  = A298 & ~A266;
  assign \new_[37624]_  = ~A265 & \new_[37623]_ ;
  assign \new_[37628]_  = A301 & A300;
  assign \new_[37629]_  = ~A299 & \new_[37628]_ ;
  assign \new_[37630]_  = \new_[37629]_  & \new_[37624]_ ;
  assign \new_[37634]_  = ~A167 & A168;
  assign \new_[37635]_  = A169 & \new_[37634]_ ;
  assign \new_[37639]_  = A200 & A199;
  assign \new_[37640]_  = A166 & \new_[37639]_ ;
  assign \new_[37641]_  = \new_[37640]_  & \new_[37635]_ ;
  assign \new_[37645]_  = A298 & ~A266;
  assign \new_[37646]_  = ~A265 & \new_[37645]_ ;
  assign \new_[37650]_  = ~A302 & A300;
  assign \new_[37651]_  = ~A299 & \new_[37650]_ ;
  assign \new_[37652]_  = \new_[37651]_  & \new_[37646]_ ;
  assign \new_[37656]_  = ~A167 & A168;
  assign \new_[37657]_  = A169 & \new_[37656]_ ;
  assign \new_[37661]_  = A200 & A199;
  assign \new_[37662]_  = A166 & \new_[37661]_ ;
  assign \new_[37663]_  = \new_[37662]_  & \new_[37657]_ ;
  assign \new_[37667]_  = ~A298 & ~A266;
  assign \new_[37668]_  = ~A265 & \new_[37667]_ ;
  assign \new_[37672]_  = A301 & A300;
  assign \new_[37673]_  = A299 & \new_[37672]_ ;
  assign \new_[37674]_  = \new_[37673]_  & \new_[37668]_ ;
  assign \new_[37678]_  = ~A167 & A168;
  assign \new_[37679]_  = A169 & \new_[37678]_ ;
  assign \new_[37683]_  = A200 & A199;
  assign \new_[37684]_  = A166 & \new_[37683]_ ;
  assign \new_[37685]_  = \new_[37684]_  & \new_[37679]_ ;
  assign \new_[37689]_  = ~A298 & ~A266;
  assign \new_[37690]_  = ~A265 & \new_[37689]_ ;
  assign \new_[37694]_  = ~A302 & A300;
  assign \new_[37695]_  = A299 & \new_[37694]_ ;
  assign \new_[37696]_  = \new_[37695]_  & \new_[37690]_ ;
  assign \new_[37700]_  = ~A167 & A168;
  assign \new_[37701]_  = A169 & \new_[37700]_ ;
  assign \new_[37705]_  = ~A200 & ~A199;
  assign \new_[37706]_  = A166 & \new_[37705]_ ;
  assign \new_[37707]_  = \new_[37706]_  & \new_[37701]_ ;
  assign \new_[37711]_  = A298 & A268;
  assign \new_[37712]_  = ~A267 & \new_[37711]_ ;
  assign \new_[37716]_  = A301 & A300;
  assign \new_[37717]_  = ~A299 & \new_[37716]_ ;
  assign \new_[37718]_  = \new_[37717]_  & \new_[37712]_ ;
  assign \new_[37722]_  = ~A167 & A168;
  assign \new_[37723]_  = A169 & \new_[37722]_ ;
  assign \new_[37727]_  = ~A200 & ~A199;
  assign \new_[37728]_  = A166 & \new_[37727]_ ;
  assign \new_[37729]_  = \new_[37728]_  & \new_[37723]_ ;
  assign \new_[37733]_  = A298 & A268;
  assign \new_[37734]_  = ~A267 & \new_[37733]_ ;
  assign \new_[37738]_  = ~A302 & A300;
  assign \new_[37739]_  = ~A299 & \new_[37738]_ ;
  assign \new_[37740]_  = \new_[37739]_  & \new_[37734]_ ;
  assign \new_[37744]_  = ~A167 & A168;
  assign \new_[37745]_  = A169 & \new_[37744]_ ;
  assign \new_[37749]_  = ~A200 & ~A199;
  assign \new_[37750]_  = A166 & \new_[37749]_ ;
  assign \new_[37751]_  = \new_[37750]_  & \new_[37745]_ ;
  assign \new_[37755]_  = ~A298 & A268;
  assign \new_[37756]_  = ~A267 & \new_[37755]_ ;
  assign \new_[37760]_  = A301 & A300;
  assign \new_[37761]_  = A299 & \new_[37760]_ ;
  assign \new_[37762]_  = \new_[37761]_  & \new_[37756]_ ;
  assign \new_[37766]_  = ~A167 & A168;
  assign \new_[37767]_  = A169 & \new_[37766]_ ;
  assign \new_[37771]_  = ~A200 & ~A199;
  assign \new_[37772]_  = A166 & \new_[37771]_ ;
  assign \new_[37773]_  = \new_[37772]_  & \new_[37767]_ ;
  assign \new_[37777]_  = ~A298 & A268;
  assign \new_[37778]_  = ~A267 & \new_[37777]_ ;
  assign \new_[37782]_  = ~A302 & A300;
  assign \new_[37783]_  = A299 & \new_[37782]_ ;
  assign \new_[37784]_  = \new_[37783]_  & \new_[37778]_ ;
  assign \new_[37788]_  = ~A167 & A168;
  assign \new_[37789]_  = A169 & \new_[37788]_ ;
  assign \new_[37793]_  = ~A200 & ~A199;
  assign \new_[37794]_  = A166 & \new_[37793]_ ;
  assign \new_[37795]_  = \new_[37794]_  & \new_[37789]_ ;
  assign \new_[37799]_  = A298 & ~A269;
  assign \new_[37800]_  = ~A267 & \new_[37799]_ ;
  assign \new_[37804]_  = A301 & A300;
  assign \new_[37805]_  = ~A299 & \new_[37804]_ ;
  assign \new_[37806]_  = \new_[37805]_  & \new_[37800]_ ;
  assign \new_[37810]_  = ~A167 & A168;
  assign \new_[37811]_  = A169 & \new_[37810]_ ;
  assign \new_[37815]_  = ~A200 & ~A199;
  assign \new_[37816]_  = A166 & \new_[37815]_ ;
  assign \new_[37817]_  = \new_[37816]_  & \new_[37811]_ ;
  assign \new_[37821]_  = A298 & ~A269;
  assign \new_[37822]_  = ~A267 & \new_[37821]_ ;
  assign \new_[37826]_  = ~A302 & A300;
  assign \new_[37827]_  = ~A299 & \new_[37826]_ ;
  assign \new_[37828]_  = \new_[37827]_  & \new_[37822]_ ;
  assign \new_[37832]_  = ~A167 & A168;
  assign \new_[37833]_  = A169 & \new_[37832]_ ;
  assign \new_[37837]_  = ~A200 & ~A199;
  assign \new_[37838]_  = A166 & \new_[37837]_ ;
  assign \new_[37839]_  = \new_[37838]_  & \new_[37833]_ ;
  assign \new_[37843]_  = ~A298 & ~A269;
  assign \new_[37844]_  = ~A267 & \new_[37843]_ ;
  assign \new_[37848]_  = A301 & A300;
  assign \new_[37849]_  = A299 & \new_[37848]_ ;
  assign \new_[37850]_  = \new_[37849]_  & \new_[37844]_ ;
  assign \new_[37854]_  = ~A167 & A168;
  assign \new_[37855]_  = A169 & \new_[37854]_ ;
  assign \new_[37859]_  = ~A200 & ~A199;
  assign \new_[37860]_  = A166 & \new_[37859]_ ;
  assign \new_[37861]_  = \new_[37860]_  & \new_[37855]_ ;
  assign \new_[37865]_  = ~A298 & ~A269;
  assign \new_[37866]_  = ~A267 & \new_[37865]_ ;
  assign \new_[37870]_  = ~A302 & A300;
  assign \new_[37871]_  = A299 & \new_[37870]_ ;
  assign \new_[37872]_  = \new_[37871]_  & \new_[37866]_ ;
  assign \new_[37876]_  = ~A167 & A168;
  assign \new_[37877]_  = A169 & \new_[37876]_ ;
  assign \new_[37881]_  = ~A200 & ~A199;
  assign \new_[37882]_  = A166 & \new_[37881]_ ;
  assign \new_[37883]_  = \new_[37882]_  & \new_[37877]_ ;
  assign \new_[37887]_  = A298 & A266;
  assign \new_[37888]_  = A265 & \new_[37887]_ ;
  assign \new_[37892]_  = A301 & A300;
  assign \new_[37893]_  = ~A299 & \new_[37892]_ ;
  assign \new_[37894]_  = \new_[37893]_  & \new_[37888]_ ;
  assign \new_[37898]_  = ~A167 & A168;
  assign \new_[37899]_  = A169 & \new_[37898]_ ;
  assign \new_[37903]_  = ~A200 & ~A199;
  assign \new_[37904]_  = A166 & \new_[37903]_ ;
  assign \new_[37905]_  = \new_[37904]_  & \new_[37899]_ ;
  assign \new_[37909]_  = A298 & A266;
  assign \new_[37910]_  = A265 & \new_[37909]_ ;
  assign \new_[37914]_  = ~A302 & A300;
  assign \new_[37915]_  = ~A299 & \new_[37914]_ ;
  assign \new_[37916]_  = \new_[37915]_  & \new_[37910]_ ;
  assign \new_[37920]_  = ~A167 & A168;
  assign \new_[37921]_  = A169 & \new_[37920]_ ;
  assign \new_[37925]_  = ~A200 & ~A199;
  assign \new_[37926]_  = A166 & \new_[37925]_ ;
  assign \new_[37927]_  = \new_[37926]_  & \new_[37921]_ ;
  assign \new_[37931]_  = ~A298 & A266;
  assign \new_[37932]_  = A265 & \new_[37931]_ ;
  assign \new_[37936]_  = A301 & A300;
  assign \new_[37937]_  = A299 & \new_[37936]_ ;
  assign \new_[37938]_  = \new_[37937]_  & \new_[37932]_ ;
  assign \new_[37942]_  = ~A167 & A168;
  assign \new_[37943]_  = A169 & \new_[37942]_ ;
  assign \new_[37947]_  = ~A200 & ~A199;
  assign \new_[37948]_  = A166 & \new_[37947]_ ;
  assign \new_[37949]_  = \new_[37948]_  & \new_[37943]_ ;
  assign \new_[37953]_  = ~A298 & A266;
  assign \new_[37954]_  = A265 & \new_[37953]_ ;
  assign \new_[37958]_  = ~A302 & A300;
  assign \new_[37959]_  = A299 & \new_[37958]_ ;
  assign \new_[37960]_  = \new_[37959]_  & \new_[37954]_ ;
  assign \new_[37964]_  = ~A167 & A168;
  assign \new_[37965]_  = A169 & \new_[37964]_ ;
  assign \new_[37969]_  = ~A200 & ~A199;
  assign \new_[37970]_  = A166 & \new_[37969]_ ;
  assign \new_[37971]_  = \new_[37970]_  & \new_[37965]_ ;
  assign \new_[37975]_  = A267 & A266;
  assign \new_[37976]_  = ~A265 & \new_[37975]_ ;
  assign \new_[37980]_  = A301 & ~A300;
  assign \new_[37981]_  = A268 & \new_[37980]_ ;
  assign \new_[37982]_  = \new_[37981]_  & \new_[37976]_ ;
  assign \new_[37986]_  = ~A167 & A168;
  assign \new_[37987]_  = A169 & \new_[37986]_ ;
  assign \new_[37991]_  = ~A200 & ~A199;
  assign \new_[37992]_  = A166 & \new_[37991]_ ;
  assign \new_[37993]_  = \new_[37992]_  & \new_[37987]_ ;
  assign \new_[37997]_  = A267 & A266;
  assign \new_[37998]_  = ~A265 & \new_[37997]_ ;
  assign \new_[38002]_  = ~A302 & ~A300;
  assign \new_[38003]_  = A268 & \new_[38002]_ ;
  assign \new_[38004]_  = \new_[38003]_  & \new_[37998]_ ;
  assign \new_[38008]_  = ~A167 & A168;
  assign \new_[38009]_  = A169 & \new_[38008]_ ;
  assign \new_[38013]_  = ~A200 & ~A199;
  assign \new_[38014]_  = A166 & \new_[38013]_ ;
  assign \new_[38015]_  = \new_[38014]_  & \new_[38009]_ ;
  assign \new_[38019]_  = A267 & A266;
  assign \new_[38020]_  = ~A265 & \new_[38019]_ ;
  assign \new_[38024]_  = A299 & A298;
  assign \new_[38025]_  = A268 & \new_[38024]_ ;
  assign \new_[38026]_  = \new_[38025]_  & \new_[38020]_ ;
  assign \new_[38030]_  = ~A167 & A168;
  assign \new_[38031]_  = A169 & \new_[38030]_ ;
  assign \new_[38035]_  = ~A200 & ~A199;
  assign \new_[38036]_  = A166 & \new_[38035]_ ;
  assign \new_[38037]_  = \new_[38036]_  & \new_[38031]_ ;
  assign \new_[38041]_  = A267 & A266;
  assign \new_[38042]_  = ~A265 & \new_[38041]_ ;
  assign \new_[38046]_  = ~A299 & ~A298;
  assign \new_[38047]_  = A268 & \new_[38046]_ ;
  assign \new_[38048]_  = \new_[38047]_  & \new_[38042]_ ;
  assign \new_[38052]_  = ~A167 & A168;
  assign \new_[38053]_  = A169 & \new_[38052]_ ;
  assign \new_[38057]_  = ~A200 & ~A199;
  assign \new_[38058]_  = A166 & \new_[38057]_ ;
  assign \new_[38059]_  = \new_[38058]_  & \new_[38053]_ ;
  assign \new_[38063]_  = A267 & A266;
  assign \new_[38064]_  = ~A265 & \new_[38063]_ ;
  assign \new_[38068]_  = A301 & ~A300;
  assign \new_[38069]_  = ~A269 & \new_[38068]_ ;
  assign \new_[38070]_  = \new_[38069]_  & \new_[38064]_ ;
  assign \new_[38074]_  = ~A167 & A168;
  assign \new_[38075]_  = A169 & \new_[38074]_ ;
  assign \new_[38079]_  = ~A200 & ~A199;
  assign \new_[38080]_  = A166 & \new_[38079]_ ;
  assign \new_[38081]_  = \new_[38080]_  & \new_[38075]_ ;
  assign \new_[38085]_  = A267 & A266;
  assign \new_[38086]_  = ~A265 & \new_[38085]_ ;
  assign \new_[38090]_  = ~A302 & ~A300;
  assign \new_[38091]_  = ~A269 & \new_[38090]_ ;
  assign \new_[38092]_  = \new_[38091]_  & \new_[38086]_ ;
  assign \new_[38096]_  = ~A167 & A168;
  assign \new_[38097]_  = A169 & \new_[38096]_ ;
  assign \new_[38101]_  = ~A200 & ~A199;
  assign \new_[38102]_  = A166 & \new_[38101]_ ;
  assign \new_[38103]_  = \new_[38102]_  & \new_[38097]_ ;
  assign \new_[38107]_  = A267 & A266;
  assign \new_[38108]_  = ~A265 & \new_[38107]_ ;
  assign \new_[38112]_  = A299 & A298;
  assign \new_[38113]_  = ~A269 & \new_[38112]_ ;
  assign \new_[38114]_  = \new_[38113]_  & \new_[38108]_ ;
  assign \new_[38118]_  = ~A167 & A168;
  assign \new_[38119]_  = A169 & \new_[38118]_ ;
  assign \new_[38123]_  = ~A200 & ~A199;
  assign \new_[38124]_  = A166 & \new_[38123]_ ;
  assign \new_[38125]_  = \new_[38124]_  & \new_[38119]_ ;
  assign \new_[38129]_  = A267 & A266;
  assign \new_[38130]_  = ~A265 & \new_[38129]_ ;
  assign \new_[38134]_  = ~A299 & ~A298;
  assign \new_[38135]_  = ~A269 & \new_[38134]_ ;
  assign \new_[38136]_  = \new_[38135]_  & \new_[38130]_ ;
  assign \new_[38140]_  = ~A167 & A168;
  assign \new_[38141]_  = A169 & \new_[38140]_ ;
  assign \new_[38145]_  = ~A200 & ~A199;
  assign \new_[38146]_  = A166 & \new_[38145]_ ;
  assign \new_[38147]_  = \new_[38146]_  & \new_[38141]_ ;
  assign \new_[38151]_  = A267 & ~A266;
  assign \new_[38152]_  = A265 & \new_[38151]_ ;
  assign \new_[38156]_  = A301 & ~A300;
  assign \new_[38157]_  = A268 & \new_[38156]_ ;
  assign \new_[38158]_  = \new_[38157]_  & \new_[38152]_ ;
  assign \new_[38162]_  = ~A167 & A168;
  assign \new_[38163]_  = A169 & \new_[38162]_ ;
  assign \new_[38167]_  = ~A200 & ~A199;
  assign \new_[38168]_  = A166 & \new_[38167]_ ;
  assign \new_[38169]_  = \new_[38168]_  & \new_[38163]_ ;
  assign \new_[38173]_  = A267 & ~A266;
  assign \new_[38174]_  = A265 & \new_[38173]_ ;
  assign \new_[38178]_  = ~A302 & ~A300;
  assign \new_[38179]_  = A268 & \new_[38178]_ ;
  assign \new_[38180]_  = \new_[38179]_  & \new_[38174]_ ;
  assign \new_[38184]_  = ~A167 & A168;
  assign \new_[38185]_  = A169 & \new_[38184]_ ;
  assign \new_[38189]_  = ~A200 & ~A199;
  assign \new_[38190]_  = A166 & \new_[38189]_ ;
  assign \new_[38191]_  = \new_[38190]_  & \new_[38185]_ ;
  assign \new_[38195]_  = A267 & ~A266;
  assign \new_[38196]_  = A265 & \new_[38195]_ ;
  assign \new_[38200]_  = A299 & A298;
  assign \new_[38201]_  = A268 & \new_[38200]_ ;
  assign \new_[38202]_  = \new_[38201]_  & \new_[38196]_ ;
  assign \new_[38206]_  = ~A167 & A168;
  assign \new_[38207]_  = A169 & \new_[38206]_ ;
  assign \new_[38211]_  = ~A200 & ~A199;
  assign \new_[38212]_  = A166 & \new_[38211]_ ;
  assign \new_[38213]_  = \new_[38212]_  & \new_[38207]_ ;
  assign \new_[38217]_  = A267 & ~A266;
  assign \new_[38218]_  = A265 & \new_[38217]_ ;
  assign \new_[38222]_  = ~A299 & ~A298;
  assign \new_[38223]_  = A268 & \new_[38222]_ ;
  assign \new_[38224]_  = \new_[38223]_  & \new_[38218]_ ;
  assign \new_[38228]_  = ~A167 & A168;
  assign \new_[38229]_  = A169 & \new_[38228]_ ;
  assign \new_[38233]_  = ~A200 & ~A199;
  assign \new_[38234]_  = A166 & \new_[38233]_ ;
  assign \new_[38235]_  = \new_[38234]_  & \new_[38229]_ ;
  assign \new_[38239]_  = A267 & ~A266;
  assign \new_[38240]_  = A265 & \new_[38239]_ ;
  assign \new_[38244]_  = A301 & ~A300;
  assign \new_[38245]_  = ~A269 & \new_[38244]_ ;
  assign \new_[38246]_  = \new_[38245]_  & \new_[38240]_ ;
  assign \new_[38250]_  = ~A167 & A168;
  assign \new_[38251]_  = A169 & \new_[38250]_ ;
  assign \new_[38255]_  = ~A200 & ~A199;
  assign \new_[38256]_  = A166 & \new_[38255]_ ;
  assign \new_[38257]_  = \new_[38256]_  & \new_[38251]_ ;
  assign \new_[38261]_  = A267 & ~A266;
  assign \new_[38262]_  = A265 & \new_[38261]_ ;
  assign \new_[38266]_  = ~A302 & ~A300;
  assign \new_[38267]_  = ~A269 & \new_[38266]_ ;
  assign \new_[38268]_  = \new_[38267]_  & \new_[38262]_ ;
  assign \new_[38272]_  = ~A167 & A168;
  assign \new_[38273]_  = A169 & \new_[38272]_ ;
  assign \new_[38277]_  = ~A200 & ~A199;
  assign \new_[38278]_  = A166 & \new_[38277]_ ;
  assign \new_[38279]_  = \new_[38278]_  & \new_[38273]_ ;
  assign \new_[38283]_  = A267 & ~A266;
  assign \new_[38284]_  = A265 & \new_[38283]_ ;
  assign \new_[38288]_  = A299 & A298;
  assign \new_[38289]_  = ~A269 & \new_[38288]_ ;
  assign \new_[38290]_  = \new_[38289]_  & \new_[38284]_ ;
  assign \new_[38294]_  = ~A167 & A168;
  assign \new_[38295]_  = A169 & \new_[38294]_ ;
  assign \new_[38299]_  = ~A200 & ~A199;
  assign \new_[38300]_  = A166 & \new_[38299]_ ;
  assign \new_[38301]_  = \new_[38300]_  & \new_[38295]_ ;
  assign \new_[38305]_  = A267 & ~A266;
  assign \new_[38306]_  = A265 & \new_[38305]_ ;
  assign \new_[38310]_  = ~A299 & ~A298;
  assign \new_[38311]_  = ~A269 & \new_[38310]_ ;
  assign \new_[38312]_  = \new_[38311]_  & \new_[38306]_ ;
  assign \new_[38316]_  = ~A167 & A168;
  assign \new_[38317]_  = A169 & \new_[38316]_ ;
  assign \new_[38321]_  = ~A200 & ~A199;
  assign \new_[38322]_  = A166 & \new_[38321]_ ;
  assign \new_[38323]_  = \new_[38322]_  & \new_[38317]_ ;
  assign \new_[38327]_  = A298 & ~A266;
  assign \new_[38328]_  = ~A265 & \new_[38327]_ ;
  assign \new_[38332]_  = A301 & A300;
  assign \new_[38333]_  = ~A299 & \new_[38332]_ ;
  assign \new_[38334]_  = \new_[38333]_  & \new_[38328]_ ;
  assign \new_[38338]_  = ~A167 & A168;
  assign \new_[38339]_  = A169 & \new_[38338]_ ;
  assign \new_[38343]_  = ~A200 & ~A199;
  assign \new_[38344]_  = A166 & \new_[38343]_ ;
  assign \new_[38345]_  = \new_[38344]_  & \new_[38339]_ ;
  assign \new_[38349]_  = A298 & ~A266;
  assign \new_[38350]_  = ~A265 & \new_[38349]_ ;
  assign \new_[38354]_  = ~A302 & A300;
  assign \new_[38355]_  = ~A299 & \new_[38354]_ ;
  assign \new_[38356]_  = \new_[38355]_  & \new_[38350]_ ;
  assign \new_[38360]_  = ~A167 & A168;
  assign \new_[38361]_  = A169 & \new_[38360]_ ;
  assign \new_[38365]_  = ~A200 & ~A199;
  assign \new_[38366]_  = A166 & \new_[38365]_ ;
  assign \new_[38367]_  = \new_[38366]_  & \new_[38361]_ ;
  assign \new_[38371]_  = ~A298 & ~A266;
  assign \new_[38372]_  = ~A265 & \new_[38371]_ ;
  assign \new_[38376]_  = A301 & A300;
  assign \new_[38377]_  = A299 & \new_[38376]_ ;
  assign \new_[38378]_  = \new_[38377]_  & \new_[38372]_ ;
  assign \new_[38382]_  = ~A167 & A168;
  assign \new_[38383]_  = A169 & \new_[38382]_ ;
  assign \new_[38387]_  = ~A200 & ~A199;
  assign \new_[38388]_  = A166 & \new_[38387]_ ;
  assign \new_[38389]_  = \new_[38388]_  & \new_[38383]_ ;
  assign \new_[38393]_  = ~A298 & ~A266;
  assign \new_[38394]_  = ~A265 & \new_[38393]_ ;
  assign \new_[38398]_  = ~A302 & A300;
  assign \new_[38399]_  = A299 & \new_[38398]_ ;
  assign \new_[38400]_  = \new_[38399]_  & \new_[38394]_ ;
  assign \new_[38404]_  = ~A232 & ~A168;
  assign \new_[38405]_  = A169 & \new_[38404]_ ;
  assign \new_[38409]_  = ~A235 & ~A234;
  assign \new_[38410]_  = A233 & \new_[38409]_ ;
  assign \new_[38411]_  = \new_[38410]_  & \new_[38405]_ ;
  assign \new_[38415]_  = A266 & ~A265;
  assign \new_[38416]_  = A236 & \new_[38415]_ ;
  assign \new_[38420]_  = A269 & ~A268;
  assign \new_[38421]_  = ~A267 & \new_[38420]_ ;
  assign \new_[38422]_  = \new_[38421]_  & \new_[38416]_ ;
  assign \new_[38426]_  = ~A232 & ~A168;
  assign \new_[38427]_  = A169 & \new_[38426]_ ;
  assign \new_[38431]_  = ~A235 & ~A234;
  assign \new_[38432]_  = A233 & \new_[38431]_ ;
  assign \new_[38433]_  = \new_[38432]_  & \new_[38427]_ ;
  assign \new_[38437]_  = ~A266 & A265;
  assign \new_[38438]_  = A236 & \new_[38437]_ ;
  assign \new_[38442]_  = A269 & ~A268;
  assign \new_[38443]_  = ~A267 & \new_[38442]_ ;
  assign \new_[38444]_  = \new_[38443]_  & \new_[38438]_ ;
  assign \new_[38448]_  = A232 & ~A168;
  assign \new_[38449]_  = A169 & \new_[38448]_ ;
  assign \new_[38453]_  = ~A235 & ~A234;
  assign \new_[38454]_  = ~A233 & \new_[38453]_ ;
  assign \new_[38455]_  = \new_[38454]_  & \new_[38449]_ ;
  assign \new_[38459]_  = A266 & ~A265;
  assign \new_[38460]_  = A236 & \new_[38459]_ ;
  assign \new_[38464]_  = A269 & ~A268;
  assign \new_[38465]_  = ~A267 & \new_[38464]_ ;
  assign \new_[38466]_  = \new_[38465]_  & \new_[38460]_ ;
  assign \new_[38470]_  = A232 & ~A168;
  assign \new_[38471]_  = A169 & \new_[38470]_ ;
  assign \new_[38475]_  = ~A235 & ~A234;
  assign \new_[38476]_  = ~A233 & \new_[38475]_ ;
  assign \new_[38477]_  = \new_[38476]_  & \new_[38471]_ ;
  assign \new_[38481]_  = ~A266 & A265;
  assign \new_[38482]_  = A236 & \new_[38481]_ ;
  assign \new_[38486]_  = A269 & ~A268;
  assign \new_[38487]_  = ~A267 & \new_[38486]_ ;
  assign \new_[38488]_  = \new_[38487]_  & \new_[38482]_ ;
  assign \new_[38492]_  = ~A199 & ~A168;
  assign \new_[38493]_  = A169 & \new_[38492]_ ;
  assign \new_[38497]_  = A202 & A201;
  assign \new_[38498]_  = A200 & \new_[38497]_ ;
  assign \new_[38499]_  = \new_[38498]_  & \new_[38493]_ ;
  assign \new_[38503]_  = A269 & ~A268;
  assign \new_[38504]_  = A267 & \new_[38503]_ ;
  assign \new_[38508]_  = A302 & ~A301;
  assign \new_[38509]_  = A300 & \new_[38508]_ ;
  assign \new_[38510]_  = \new_[38509]_  & \new_[38504]_ ;
  assign \new_[38514]_  = ~A199 & ~A168;
  assign \new_[38515]_  = A169 & \new_[38514]_ ;
  assign \new_[38519]_  = ~A203 & A201;
  assign \new_[38520]_  = A200 & \new_[38519]_ ;
  assign \new_[38521]_  = \new_[38520]_  & \new_[38515]_ ;
  assign \new_[38525]_  = A269 & ~A268;
  assign \new_[38526]_  = A267 & \new_[38525]_ ;
  assign \new_[38530]_  = A302 & ~A301;
  assign \new_[38531]_  = A300 & \new_[38530]_ ;
  assign \new_[38532]_  = \new_[38531]_  & \new_[38526]_ ;
  assign \new_[38536]_  = ~A199 & ~A168;
  assign \new_[38537]_  = A169 & \new_[38536]_ ;
  assign \new_[38541]_  = ~A202 & ~A201;
  assign \new_[38542]_  = A200 & \new_[38541]_ ;
  assign \new_[38543]_  = \new_[38542]_  & \new_[38537]_ ;
  assign \new_[38547]_  = ~A268 & A267;
  assign \new_[38548]_  = A203 & \new_[38547]_ ;
  assign \new_[38552]_  = A301 & ~A300;
  assign \new_[38553]_  = A269 & \new_[38552]_ ;
  assign \new_[38554]_  = \new_[38553]_  & \new_[38548]_ ;
  assign \new_[38558]_  = ~A199 & ~A168;
  assign \new_[38559]_  = A169 & \new_[38558]_ ;
  assign \new_[38563]_  = ~A202 & ~A201;
  assign \new_[38564]_  = A200 & \new_[38563]_ ;
  assign \new_[38565]_  = \new_[38564]_  & \new_[38559]_ ;
  assign \new_[38569]_  = ~A268 & A267;
  assign \new_[38570]_  = A203 & \new_[38569]_ ;
  assign \new_[38574]_  = ~A302 & ~A300;
  assign \new_[38575]_  = A269 & \new_[38574]_ ;
  assign \new_[38576]_  = \new_[38575]_  & \new_[38570]_ ;
  assign \new_[38580]_  = ~A199 & ~A168;
  assign \new_[38581]_  = A169 & \new_[38580]_ ;
  assign \new_[38585]_  = ~A202 & ~A201;
  assign \new_[38586]_  = A200 & \new_[38585]_ ;
  assign \new_[38587]_  = \new_[38586]_  & \new_[38581]_ ;
  assign \new_[38591]_  = ~A268 & A267;
  assign \new_[38592]_  = A203 & \new_[38591]_ ;
  assign \new_[38596]_  = A299 & A298;
  assign \new_[38597]_  = A269 & \new_[38596]_ ;
  assign \new_[38598]_  = \new_[38597]_  & \new_[38592]_ ;
  assign \new_[38602]_  = ~A199 & ~A168;
  assign \new_[38603]_  = A169 & \new_[38602]_ ;
  assign \new_[38607]_  = ~A202 & ~A201;
  assign \new_[38608]_  = A200 & \new_[38607]_ ;
  assign \new_[38609]_  = \new_[38608]_  & \new_[38603]_ ;
  assign \new_[38613]_  = ~A268 & A267;
  assign \new_[38614]_  = A203 & \new_[38613]_ ;
  assign \new_[38618]_  = ~A299 & ~A298;
  assign \new_[38619]_  = A269 & \new_[38618]_ ;
  assign \new_[38620]_  = \new_[38619]_  & \new_[38614]_ ;
  assign \new_[38624]_  = ~A199 & ~A168;
  assign \new_[38625]_  = A169 & \new_[38624]_ ;
  assign \new_[38629]_  = ~A202 & ~A201;
  assign \new_[38630]_  = A200 & \new_[38629]_ ;
  assign \new_[38631]_  = \new_[38630]_  & \new_[38625]_ ;
  assign \new_[38635]_  = A268 & ~A267;
  assign \new_[38636]_  = A203 & \new_[38635]_ ;
  assign \new_[38640]_  = A302 & ~A301;
  assign \new_[38641]_  = A300 & \new_[38640]_ ;
  assign \new_[38642]_  = \new_[38641]_  & \new_[38636]_ ;
  assign \new_[38646]_  = ~A199 & ~A168;
  assign \new_[38647]_  = A169 & \new_[38646]_ ;
  assign \new_[38651]_  = ~A202 & ~A201;
  assign \new_[38652]_  = A200 & \new_[38651]_ ;
  assign \new_[38653]_  = \new_[38652]_  & \new_[38647]_ ;
  assign \new_[38657]_  = ~A269 & ~A267;
  assign \new_[38658]_  = A203 & \new_[38657]_ ;
  assign \new_[38662]_  = A302 & ~A301;
  assign \new_[38663]_  = A300 & \new_[38662]_ ;
  assign \new_[38664]_  = \new_[38663]_  & \new_[38658]_ ;
  assign \new_[38668]_  = ~A199 & ~A168;
  assign \new_[38669]_  = A169 & \new_[38668]_ ;
  assign \new_[38673]_  = ~A202 & ~A201;
  assign \new_[38674]_  = A200 & \new_[38673]_ ;
  assign \new_[38675]_  = \new_[38674]_  & \new_[38669]_ ;
  assign \new_[38679]_  = A266 & A265;
  assign \new_[38680]_  = A203 & \new_[38679]_ ;
  assign \new_[38684]_  = A302 & ~A301;
  assign \new_[38685]_  = A300 & \new_[38684]_ ;
  assign \new_[38686]_  = \new_[38685]_  & \new_[38680]_ ;
  assign \new_[38690]_  = ~A199 & ~A168;
  assign \new_[38691]_  = A169 & \new_[38690]_ ;
  assign \new_[38695]_  = ~A202 & ~A201;
  assign \new_[38696]_  = A200 & \new_[38695]_ ;
  assign \new_[38697]_  = \new_[38696]_  & \new_[38691]_ ;
  assign \new_[38701]_  = ~A266 & ~A265;
  assign \new_[38702]_  = A203 & \new_[38701]_ ;
  assign \new_[38706]_  = A302 & ~A301;
  assign \new_[38707]_  = A300 & \new_[38706]_ ;
  assign \new_[38708]_  = \new_[38707]_  & \new_[38702]_ ;
  assign \new_[38712]_  = A199 & ~A168;
  assign \new_[38713]_  = A169 & \new_[38712]_ ;
  assign \new_[38717]_  = A202 & A201;
  assign \new_[38718]_  = ~A200 & \new_[38717]_ ;
  assign \new_[38719]_  = \new_[38718]_  & \new_[38713]_ ;
  assign \new_[38723]_  = A269 & ~A268;
  assign \new_[38724]_  = A267 & \new_[38723]_ ;
  assign \new_[38728]_  = A302 & ~A301;
  assign \new_[38729]_  = A300 & \new_[38728]_ ;
  assign \new_[38730]_  = \new_[38729]_  & \new_[38724]_ ;
  assign \new_[38734]_  = A199 & ~A168;
  assign \new_[38735]_  = A169 & \new_[38734]_ ;
  assign \new_[38739]_  = ~A203 & A201;
  assign \new_[38740]_  = ~A200 & \new_[38739]_ ;
  assign \new_[38741]_  = \new_[38740]_  & \new_[38735]_ ;
  assign \new_[38745]_  = A269 & ~A268;
  assign \new_[38746]_  = A267 & \new_[38745]_ ;
  assign \new_[38750]_  = A302 & ~A301;
  assign \new_[38751]_  = A300 & \new_[38750]_ ;
  assign \new_[38752]_  = \new_[38751]_  & \new_[38746]_ ;
  assign \new_[38756]_  = A199 & ~A168;
  assign \new_[38757]_  = A169 & \new_[38756]_ ;
  assign \new_[38761]_  = ~A202 & ~A201;
  assign \new_[38762]_  = ~A200 & \new_[38761]_ ;
  assign \new_[38763]_  = \new_[38762]_  & \new_[38757]_ ;
  assign \new_[38767]_  = ~A268 & A267;
  assign \new_[38768]_  = A203 & \new_[38767]_ ;
  assign \new_[38772]_  = A301 & ~A300;
  assign \new_[38773]_  = A269 & \new_[38772]_ ;
  assign \new_[38774]_  = \new_[38773]_  & \new_[38768]_ ;
  assign \new_[38778]_  = A199 & ~A168;
  assign \new_[38779]_  = A169 & \new_[38778]_ ;
  assign \new_[38783]_  = ~A202 & ~A201;
  assign \new_[38784]_  = ~A200 & \new_[38783]_ ;
  assign \new_[38785]_  = \new_[38784]_  & \new_[38779]_ ;
  assign \new_[38789]_  = ~A268 & A267;
  assign \new_[38790]_  = A203 & \new_[38789]_ ;
  assign \new_[38794]_  = ~A302 & ~A300;
  assign \new_[38795]_  = A269 & \new_[38794]_ ;
  assign \new_[38796]_  = \new_[38795]_  & \new_[38790]_ ;
  assign \new_[38800]_  = A199 & ~A168;
  assign \new_[38801]_  = A169 & \new_[38800]_ ;
  assign \new_[38805]_  = ~A202 & ~A201;
  assign \new_[38806]_  = ~A200 & \new_[38805]_ ;
  assign \new_[38807]_  = \new_[38806]_  & \new_[38801]_ ;
  assign \new_[38811]_  = ~A268 & A267;
  assign \new_[38812]_  = A203 & \new_[38811]_ ;
  assign \new_[38816]_  = A299 & A298;
  assign \new_[38817]_  = A269 & \new_[38816]_ ;
  assign \new_[38818]_  = \new_[38817]_  & \new_[38812]_ ;
  assign \new_[38822]_  = A199 & ~A168;
  assign \new_[38823]_  = A169 & \new_[38822]_ ;
  assign \new_[38827]_  = ~A202 & ~A201;
  assign \new_[38828]_  = ~A200 & \new_[38827]_ ;
  assign \new_[38829]_  = \new_[38828]_  & \new_[38823]_ ;
  assign \new_[38833]_  = ~A268 & A267;
  assign \new_[38834]_  = A203 & \new_[38833]_ ;
  assign \new_[38838]_  = ~A299 & ~A298;
  assign \new_[38839]_  = A269 & \new_[38838]_ ;
  assign \new_[38840]_  = \new_[38839]_  & \new_[38834]_ ;
  assign \new_[38844]_  = A199 & ~A168;
  assign \new_[38845]_  = A169 & \new_[38844]_ ;
  assign \new_[38849]_  = ~A202 & ~A201;
  assign \new_[38850]_  = ~A200 & \new_[38849]_ ;
  assign \new_[38851]_  = \new_[38850]_  & \new_[38845]_ ;
  assign \new_[38855]_  = A268 & ~A267;
  assign \new_[38856]_  = A203 & \new_[38855]_ ;
  assign \new_[38860]_  = A302 & ~A301;
  assign \new_[38861]_  = A300 & \new_[38860]_ ;
  assign \new_[38862]_  = \new_[38861]_  & \new_[38856]_ ;
  assign \new_[38866]_  = A199 & ~A168;
  assign \new_[38867]_  = A169 & \new_[38866]_ ;
  assign \new_[38871]_  = ~A202 & ~A201;
  assign \new_[38872]_  = ~A200 & \new_[38871]_ ;
  assign \new_[38873]_  = \new_[38872]_  & \new_[38867]_ ;
  assign \new_[38877]_  = ~A269 & ~A267;
  assign \new_[38878]_  = A203 & \new_[38877]_ ;
  assign \new_[38882]_  = A302 & ~A301;
  assign \new_[38883]_  = A300 & \new_[38882]_ ;
  assign \new_[38884]_  = \new_[38883]_  & \new_[38878]_ ;
  assign \new_[38888]_  = A199 & ~A168;
  assign \new_[38889]_  = A169 & \new_[38888]_ ;
  assign \new_[38893]_  = ~A202 & ~A201;
  assign \new_[38894]_  = ~A200 & \new_[38893]_ ;
  assign \new_[38895]_  = \new_[38894]_  & \new_[38889]_ ;
  assign \new_[38899]_  = A266 & A265;
  assign \new_[38900]_  = A203 & \new_[38899]_ ;
  assign \new_[38904]_  = A302 & ~A301;
  assign \new_[38905]_  = A300 & \new_[38904]_ ;
  assign \new_[38906]_  = \new_[38905]_  & \new_[38900]_ ;
  assign \new_[38910]_  = A199 & ~A168;
  assign \new_[38911]_  = A169 & \new_[38910]_ ;
  assign \new_[38915]_  = ~A202 & ~A201;
  assign \new_[38916]_  = ~A200 & \new_[38915]_ ;
  assign \new_[38917]_  = \new_[38916]_  & \new_[38911]_ ;
  assign \new_[38921]_  = ~A266 & ~A265;
  assign \new_[38922]_  = A203 & \new_[38921]_ ;
  assign \new_[38926]_  = A302 & ~A301;
  assign \new_[38927]_  = A300 & \new_[38926]_ ;
  assign \new_[38928]_  = \new_[38927]_  & \new_[38922]_ ;
  assign \new_[38932]_  = A168 & ~A169;
  assign \new_[38933]_  = ~A170 & \new_[38932]_ ;
  assign \new_[38937]_  = A201 & A200;
  assign \new_[38938]_  = ~A199 & \new_[38937]_ ;
  assign \new_[38939]_  = \new_[38938]_  & \new_[38933]_ ;
  assign \new_[38943]_  = ~A268 & A267;
  assign \new_[38944]_  = A202 & \new_[38943]_ ;
  assign \new_[38948]_  = A301 & ~A300;
  assign \new_[38949]_  = A269 & \new_[38948]_ ;
  assign \new_[38950]_  = \new_[38949]_  & \new_[38944]_ ;
  assign \new_[38954]_  = A168 & ~A169;
  assign \new_[38955]_  = ~A170 & \new_[38954]_ ;
  assign \new_[38959]_  = A201 & A200;
  assign \new_[38960]_  = ~A199 & \new_[38959]_ ;
  assign \new_[38961]_  = \new_[38960]_  & \new_[38955]_ ;
  assign \new_[38965]_  = ~A268 & A267;
  assign \new_[38966]_  = A202 & \new_[38965]_ ;
  assign \new_[38970]_  = ~A302 & ~A300;
  assign \new_[38971]_  = A269 & \new_[38970]_ ;
  assign \new_[38972]_  = \new_[38971]_  & \new_[38966]_ ;
  assign \new_[38976]_  = A168 & ~A169;
  assign \new_[38977]_  = ~A170 & \new_[38976]_ ;
  assign \new_[38981]_  = A201 & A200;
  assign \new_[38982]_  = ~A199 & \new_[38981]_ ;
  assign \new_[38983]_  = \new_[38982]_  & \new_[38977]_ ;
  assign \new_[38987]_  = ~A268 & A267;
  assign \new_[38988]_  = A202 & \new_[38987]_ ;
  assign \new_[38992]_  = A299 & A298;
  assign \new_[38993]_  = A269 & \new_[38992]_ ;
  assign \new_[38994]_  = \new_[38993]_  & \new_[38988]_ ;
  assign \new_[38998]_  = A168 & ~A169;
  assign \new_[38999]_  = ~A170 & \new_[38998]_ ;
  assign \new_[39003]_  = A201 & A200;
  assign \new_[39004]_  = ~A199 & \new_[39003]_ ;
  assign \new_[39005]_  = \new_[39004]_  & \new_[38999]_ ;
  assign \new_[39009]_  = ~A268 & A267;
  assign \new_[39010]_  = A202 & \new_[39009]_ ;
  assign \new_[39014]_  = ~A299 & ~A298;
  assign \new_[39015]_  = A269 & \new_[39014]_ ;
  assign \new_[39016]_  = \new_[39015]_  & \new_[39010]_ ;
  assign \new_[39020]_  = A168 & ~A169;
  assign \new_[39021]_  = ~A170 & \new_[39020]_ ;
  assign \new_[39025]_  = A201 & A200;
  assign \new_[39026]_  = ~A199 & \new_[39025]_ ;
  assign \new_[39027]_  = \new_[39026]_  & \new_[39021]_ ;
  assign \new_[39031]_  = A268 & ~A267;
  assign \new_[39032]_  = A202 & \new_[39031]_ ;
  assign \new_[39036]_  = A302 & ~A301;
  assign \new_[39037]_  = A300 & \new_[39036]_ ;
  assign \new_[39038]_  = \new_[39037]_  & \new_[39032]_ ;
  assign \new_[39042]_  = A168 & ~A169;
  assign \new_[39043]_  = ~A170 & \new_[39042]_ ;
  assign \new_[39047]_  = A201 & A200;
  assign \new_[39048]_  = ~A199 & \new_[39047]_ ;
  assign \new_[39049]_  = \new_[39048]_  & \new_[39043]_ ;
  assign \new_[39053]_  = ~A269 & ~A267;
  assign \new_[39054]_  = A202 & \new_[39053]_ ;
  assign \new_[39058]_  = A302 & ~A301;
  assign \new_[39059]_  = A300 & \new_[39058]_ ;
  assign \new_[39060]_  = \new_[39059]_  & \new_[39054]_ ;
  assign \new_[39064]_  = A168 & ~A169;
  assign \new_[39065]_  = ~A170 & \new_[39064]_ ;
  assign \new_[39069]_  = A201 & A200;
  assign \new_[39070]_  = ~A199 & \new_[39069]_ ;
  assign \new_[39071]_  = \new_[39070]_  & \new_[39065]_ ;
  assign \new_[39075]_  = A266 & A265;
  assign \new_[39076]_  = A202 & \new_[39075]_ ;
  assign \new_[39080]_  = A302 & ~A301;
  assign \new_[39081]_  = A300 & \new_[39080]_ ;
  assign \new_[39082]_  = \new_[39081]_  & \new_[39076]_ ;
  assign \new_[39086]_  = A168 & ~A169;
  assign \new_[39087]_  = ~A170 & \new_[39086]_ ;
  assign \new_[39091]_  = A201 & A200;
  assign \new_[39092]_  = ~A199 & \new_[39091]_ ;
  assign \new_[39093]_  = \new_[39092]_  & \new_[39087]_ ;
  assign \new_[39097]_  = ~A266 & ~A265;
  assign \new_[39098]_  = A202 & \new_[39097]_ ;
  assign \new_[39102]_  = A302 & ~A301;
  assign \new_[39103]_  = A300 & \new_[39102]_ ;
  assign \new_[39104]_  = \new_[39103]_  & \new_[39098]_ ;
  assign \new_[39108]_  = A168 & ~A169;
  assign \new_[39109]_  = ~A170 & \new_[39108]_ ;
  assign \new_[39113]_  = A201 & A200;
  assign \new_[39114]_  = ~A199 & \new_[39113]_ ;
  assign \new_[39115]_  = \new_[39114]_  & \new_[39109]_ ;
  assign \new_[39119]_  = ~A268 & A267;
  assign \new_[39120]_  = ~A203 & \new_[39119]_ ;
  assign \new_[39124]_  = A301 & ~A300;
  assign \new_[39125]_  = A269 & \new_[39124]_ ;
  assign \new_[39126]_  = \new_[39125]_  & \new_[39120]_ ;
  assign \new_[39130]_  = A168 & ~A169;
  assign \new_[39131]_  = ~A170 & \new_[39130]_ ;
  assign \new_[39135]_  = A201 & A200;
  assign \new_[39136]_  = ~A199 & \new_[39135]_ ;
  assign \new_[39137]_  = \new_[39136]_  & \new_[39131]_ ;
  assign \new_[39141]_  = ~A268 & A267;
  assign \new_[39142]_  = ~A203 & \new_[39141]_ ;
  assign \new_[39146]_  = ~A302 & ~A300;
  assign \new_[39147]_  = A269 & \new_[39146]_ ;
  assign \new_[39148]_  = \new_[39147]_  & \new_[39142]_ ;
  assign \new_[39152]_  = A168 & ~A169;
  assign \new_[39153]_  = ~A170 & \new_[39152]_ ;
  assign \new_[39157]_  = A201 & A200;
  assign \new_[39158]_  = ~A199 & \new_[39157]_ ;
  assign \new_[39159]_  = \new_[39158]_  & \new_[39153]_ ;
  assign \new_[39163]_  = ~A268 & A267;
  assign \new_[39164]_  = ~A203 & \new_[39163]_ ;
  assign \new_[39168]_  = A299 & A298;
  assign \new_[39169]_  = A269 & \new_[39168]_ ;
  assign \new_[39170]_  = \new_[39169]_  & \new_[39164]_ ;
  assign \new_[39174]_  = A168 & ~A169;
  assign \new_[39175]_  = ~A170 & \new_[39174]_ ;
  assign \new_[39179]_  = A201 & A200;
  assign \new_[39180]_  = ~A199 & \new_[39179]_ ;
  assign \new_[39181]_  = \new_[39180]_  & \new_[39175]_ ;
  assign \new_[39185]_  = ~A268 & A267;
  assign \new_[39186]_  = ~A203 & \new_[39185]_ ;
  assign \new_[39190]_  = ~A299 & ~A298;
  assign \new_[39191]_  = A269 & \new_[39190]_ ;
  assign \new_[39192]_  = \new_[39191]_  & \new_[39186]_ ;
  assign \new_[39196]_  = A168 & ~A169;
  assign \new_[39197]_  = ~A170 & \new_[39196]_ ;
  assign \new_[39201]_  = A201 & A200;
  assign \new_[39202]_  = ~A199 & \new_[39201]_ ;
  assign \new_[39203]_  = \new_[39202]_  & \new_[39197]_ ;
  assign \new_[39207]_  = A268 & ~A267;
  assign \new_[39208]_  = ~A203 & \new_[39207]_ ;
  assign \new_[39212]_  = A302 & ~A301;
  assign \new_[39213]_  = A300 & \new_[39212]_ ;
  assign \new_[39214]_  = \new_[39213]_  & \new_[39208]_ ;
  assign \new_[39218]_  = A168 & ~A169;
  assign \new_[39219]_  = ~A170 & \new_[39218]_ ;
  assign \new_[39223]_  = A201 & A200;
  assign \new_[39224]_  = ~A199 & \new_[39223]_ ;
  assign \new_[39225]_  = \new_[39224]_  & \new_[39219]_ ;
  assign \new_[39229]_  = ~A269 & ~A267;
  assign \new_[39230]_  = ~A203 & \new_[39229]_ ;
  assign \new_[39234]_  = A302 & ~A301;
  assign \new_[39235]_  = A300 & \new_[39234]_ ;
  assign \new_[39236]_  = \new_[39235]_  & \new_[39230]_ ;
  assign \new_[39240]_  = A168 & ~A169;
  assign \new_[39241]_  = ~A170 & \new_[39240]_ ;
  assign \new_[39245]_  = A201 & A200;
  assign \new_[39246]_  = ~A199 & \new_[39245]_ ;
  assign \new_[39247]_  = \new_[39246]_  & \new_[39241]_ ;
  assign \new_[39251]_  = A266 & A265;
  assign \new_[39252]_  = ~A203 & \new_[39251]_ ;
  assign \new_[39256]_  = A302 & ~A301;
  assign \new_[39257]_  = A300 & \new_[39256]_ ;
  assign \new_[39258]_  = \new_[39257]_  & \new_[39252]_ ;
  assign \new_[39262]_  = A168 & ~A169;
  assign \new_[39263]_  = ~A170 & \new_[39262]_ ;
  assign \new_[39267]_  = A201 & A200;
  assign \new_[39268]_  = ~A199 & \new_[39267]_ ;
  assign \new_[39269]_  = \new_[39268]_  & \new_[39263]_ ;
  assign \new_[39273]_  = ~A266 & ~A265;
  assign \new_[39274]_  = ~A203 & \new_[39273]_ ;
  assign \new_[39278]_  = A302 & ~A301;
  assign \new_[39279]_  = A300 & \new_[39278]_ ;
  assign \new_[39280]_  = \new_[39279]_  & \new_[39274]_ ;
  assign \new_[39284]_  = A168 & ~A169;
  assign \new_[39285]_  = ~A170 & \new_[39284]_ ;
  assign \new_[39289]_  = ~A201 & A200;
  assign \new_[39290]_  = ~A199 & \new_[39289]_ ;
  assign \new_[39291]_  = \new_[39290]_  & \new_[39285]_ ;
  assign \new_[39295]_  = ~A267 & A203;
  assign \new_[39296]_  = ~A202 & \new_[39295]_ ;
  assign \new_[39300]_  = A301 & ~A300;
  assign \new_[39301]_  = A268 & \new_[39300]_ ;
  assign \new_[39302]_  = \new_[39301]_  & \new_[39296]_ ;
  assign \new_[39306]_  = A168 & ~A169;
  assign \new_[39307]_  = ~A170 & \new_[39306]_ ;
  assign \new_[39311]_  = ~A201 & A200;
  assign \new_[39312]_  = ~A199 & \new_[39311]_ ;
  assign \new_[39313]_  = \new_[39312]_  & \new_[39307]_ ;
  assign \new_[39317]_  = ~A267 & A203;
  assign \new_[39318]_  = ~A202 & \new_[39317]_ ;
  assign \new_[39322]_  = ~A302 & ~A300;
  assign \new_[39323]_  = A268 & \new_[39322]_ ;
  assign \new_[39324]_  = \new_[39323]_  & \new_[39318]_ ;
  assign \new_[39328]_  = A168 & ~A169;
  assign \new_[39329]_  = ~A170 & \new_[39328]_ ;
  assign \new_[39333]_  = ~A201 & A200;
  assign \new_[39334]_  = ~A199 & \new_[39333]_ ;
  assign \new_[39335]_  = \new_[39334]_  & \new_[39329]_ ;
  assign \new_[39339]_  = ~A267 & A203;
  assign \new_[39340]_  = ~A202 & \new_[39339]_ ;
  assign \new_[39344]_  = A299 & A298;
  assign \new_[39345]_  = A268 & \new_[39344]_ ;
  assign \new_[39346]_  = \new_[39345]_  & \new_[39340]_ ;
  assign \new_[39350]_  = A168 & ~A169;
  assign \new_[39351]_  = ~A170 & \new_[39350]_ ;
  assign \new_[39355]_  = ~A201 & A200;
  assign \new_[39356]_  = ~A199 & \new_[39355]_ ;
  assign \new_[39357]_  = \new_[39356]_  & \new_[39351]_ ;
  assign \new_[39361]_  = ~A267 & A203;
  assign \new_[39362]_  = ~A202 & \new_[39361]_ ;
  assign \new_[39366]_  = ~A299 & ~A298;
  assign \new_[39367]_  = A268 & \new_[39366]_ ;
  assign \new_[39368]_  = \new_[39367]_  & \new_[39362]_ ;
  assign \new_[39372]_  = A168 & ~A169;
  assign \new_[39373]_  = ~A170 & \new_[39372]_ ;
  assign \new_[39377]_  = ~A201 & A200;
  assign \new_[39378]_  = ~A199 & \new_[39377]_ ;
  assign \new_[39379]_  = \new_[39378]_  & \new_[39373]_ ;
  assign \new_[39383]_  = ~A267 & A203;
  assign \new_[39384]_  = ~A202 & \new_[39383]_ ;
  assign \new_[39388]_  = A301 & ~A300;
  assign \new_[39389]_  = ~A269 & \new_[39388]_ ;
  assign \new_[39390]_  = \new_[39389]_  & \new_[39384]_ ;
  assign \new_[39394]_  = A168 & ~A169;
  assign \new_[39395]_  = ~A170 & \new_[39394]_ ;
  assign \new_[39399]_  = ~A201 & A200;
  assign \new_[39400]_  = ~A199 & \new_[39399]_ ;
  assign \new_[39401]_  = \new_[39400]_  & \new_[39395]_ ;
  assign \new_[39405]_  = ~A267 & A203;
  assign \new_[39406]_  = ~A202 & \new_[39405]_ ;
  assign \new_[39410]_  = ~A302 & ~A300;
  assign \new_[39411]_  = ~A269 & \new_[39410]_ ;
  assign \new_[39412]_  = \new_[39411]_  & \new_[39406]_ ;
  assign \new_[39416]_  = A168 & ~A169;
  assign \new_[39417]_  = ~A170 & \new_[39416]_ ;
  assign \new_[39421]_  = ~A201 & A200;
  assign \new_[39422]_  = ~A199 & \new_[39421]_ ;
  assign \new_[39423]_  = \new_[39422]_  & \new_[39417]_ ;
  assign \new_[39427]_  = ~A267 & A203;
  assign \new_[39428]_  = ~A202 & \new_[39427]_ ;
  assign \new_[39432]_  = A299 & A298;
  assign \new_[39433]_  = ~A269 & \new_[39432]_ ;
  assign \new_[39434]_  = \new_[39433]_  & \new_[39428]_ ;
  assign \new_[39438]_  = A168 & ~A169;
  assign \new_[39439]_  = ~A170 & \new_[39438]_ ;
  assign \new_[39443]_  = ~A201 & A200;
  assign \new_[39444]_  = ~A199 & \new_[39443]_ ;
  assign \new_[39445]_  = \new_[39444]_  & \new_[39439]_ ;
  assign \new_[39449]_  = ~A267 & A203;
  assign \new_[39450]_  = ~A202 & \new_[39449]_ ;
  assign \new_[39454]_  = ~A299 & ~A298;
  assign \new_[39455]_  = ~A269 & \new_[39454]_ ;
  assign \new_[39456]_  = \new_[39455]_  & \new_[39450]_ ;
  assign \new_[39460]_  = A168 & ~A169;
  assign \new_[39461]_  = ~A170 & \new_[39460]_ ;
  assign \new_[39465]_  = ~A201 & A200;
  assign \new_[39466]_  = ~A199 & \new_[39465]_ ;
  assign \new_[39467]_  = \new_[39466]_  & \new_[39461]_ ;
  assign \new_[39471]_  = A265 & A203;
  assign \new_[39472]_  = ~A202 & \new_[39471]_ ;
  assign \new_[39476]_  = A301 & ~A300;
  assign \new_[39477]_  = A266 & \new_[39476]_ ;
  assign \new_[39478]_  = \new_[39477]_  & \new_[39472]_ ;
  assign \new_[39482]_  = A168 & ~A169;
  assign \new_[39483]_  = ~A170 & \new_[39482]_ ;
  assign \new_[39487]_  = ~A201 & A200;
  assign \new_[39488]_  = ~A199 & \new_[39487]_ ;
  assign \new_[39489]_  = \new_[39488]_  & \new_[39483]_ ;
  assign \new_[39493]_  = A265 & A203;
  assign \new_[39494]_  = ~A202 & \new_[39493]_ ;
  assign \new_[39498]_  = ~A302 & ~A300;
  assign \new_[39499]_  = A266 & \new_[39498]_ ;
  assign \new_[39500]_  = \new_[39499]_  & \new_[39494]_ ;
  assign \new_[39504]_  = A168 & ~A169;
  assign \new_[39505]_  = ~A170 & \new_[39504]_ ;
  assign \new_[39509]_  = ~A201 & A200;
  assign \new_[39510]_  = ~A199 & \new_[39509]_ ;
  assign \new_[39511]_  = \new_[39510]_  & \new_[39505]_ ;
  assign \new_[39515]_  = A265 & A203;
  assign \new_[39516]_  = ~A202 & \new_[39515]_ ;
  assign \new_[39520]_  = A299 & A298;
  assign \new_[39521]_  = A266 & \new_[39520]_ ;
  assign \new_[39522]_  = \new_[39521]_  & \new_[39516]_ ;
  assign \new_[39526]_  = A168 & ~A169;
  assign \new_[39527]_  = ~A170 & \new_[39526]_ ;
  assign \new_[39531]_  = ~A201 & A200;
  assign \new_[39532]_  = ~A199 & \new_[39531]_ ;
  assign \new_[39533]_  = \new_[39532]_  & \new_[39527]_ ;
  assign \new_[39537]_  = A265 & A203;
  assign \new_[39538]_  = ~A202 & \new_[39537]_ ;
  assign \new_[39542]_  = ~A299 & ~A298;
  assign \new_[39543]_  = A266 & \new_[39542]_ ;
  assign \new_[39544]_  = \new_[39543]_  & \new_[39538]_ ;
  assign \new_[39548]_  = A168 & ~A169;
  assign \new_[39549]_  = ~A170 & \new_[39548]_ ;
  assign \new_[39553]_  = ~A201 & A200;
  assign \new_[39554]_  = ~A199 & \new_[39553]_ ;
  assign \new_[39555]_  = \new_[39554]_  & \new_[39549]_ ;
  assign \new_[39559]_  = ~A265 & A203;
  assign \new_[39560]_  = ~A202 & \new_[39559]_ ;
  assign \new_[39564]_  = A301 & ~A300;
  assign \new_[39565]_  = ~A266 & \new_[39564]_ ;
  assign \new_[39566]_  = \new_[39565]_  & \new_[39560]_ ;
  assign \new_[39570]_  = A168 & ~A169;
  assign \new_[39571]_  = ~A170 & \new_[39570]_ ;
  assign \new_[39575]_  = ~A201 & A200;
  assign \new_[39576]_  = ~A199 & \new_[39575]_ ;
  assign \new_[39577]_  = \new_[39576]_  & \new_[39571]_ ;
  assign \new_[39581]_  = ~A265 & A203;
  assign \new_[39582]_  = ~A202 & \new_[39581]_ ;
  assign \new_[39586]_  = ~A302 & ~A300;
  assign \new_[39587]_  = ~A266 & \new_[39586]_ ;
  assign \new_[39588]_  = \new_[39587]_  & \new_[39582]_ ;
  assign \new_[39592]_  = A168 & ~A169;
  assign \new_[39593]_  = ~A170 & \new_[39592]_ ;
  assign \new_[39597]_  = ~A201 & A200;
  assign \new_[39598]_  = ~A199 & \new_[39597]_ ;
  assign \new_[39599]_  = \new_[39598]_  & \new_[39593]_ ;
  assign \new_[39603]_  = ~A265 & A203;
  assign \new_[39604]_  = ~A202 & \new_[39603]_ ;
  assign \new_[39608]_  = A299 & A298;
  assign \new_[39609]_  = ~A266 & \new_[39608]_ ;
  assign \new_[39610]_  = \new_[39609]_  & \new_[39604]_ ;
  assign \new_[39614]_  = A168 & ~A169;
  assign \new_[39615]_  = ~A170 & \new_[39614]_ ;
  assign \new_[39619]_  = ~A201 & A200;
  assign \new_[39620]_  = ~A199 & \new_[39619]_ ;
  assign \new_[39621]_  = \new_[39620]_  & \new_[39615]_ ;
  assign \new_[39625]_  = ~A265 & A203;
  assign \new_[39626]_  = ~A202 & \new_[39625]_ ;
  assign \new_[39630]_  = ~A299 & ~A298;
  assign \new_[39631]_  = ~A266 & \new_[39630]_ ;
  assign \new_[39632]_  = \new_[39631]_  & \new_[39626]_ ;
  assign \new_[39636]_  = A168 & ~A169;
  assign \new_[39637]_  = ~A170 & \new_[39636]_ ;
  assign \new_[39641]_  = A201 & ~A200;
  assign \new_[39642]_  = A199 & \new_[39641]_ ;
  assign \new_[39643]_  = \new_[39642]_  & \new_[39637]_ ;
  assign \new_[39647]_  = ~A268 & A267;
  assign \new_[39648]_  = A202 & \new_[39647]_ ;
  assign \new_[39652]_  = A301 & ~A300;
  assign \new_[39653]_  = A269 & \new_[39652]_ ;
  assign \new_[39654]_  = \new_[39653]_  & \new_[39648]_ ;
  assign \new_[39658]_  = A168 & ~A169;
  assign \new_[39659]_  = ~A170 & \new_[39658]_ ;
  assign \new_[39663]_  = A201 & ~A200;
  assign \new_[39664]_  = A199 & \new_[39663]_ ;
  assign \new_[39665]_  = \new_[39664]_  & \new_[39659]_ ;
  assign \new_[39669]_  = ~A268 & A267;
  assign \new_[39670]_  = A202 & \new_[39669]_ ;
  assign \new_[39674]_  = ~A302 & ~A300;
  assign \new_[39675]_  = A269 & \new_[39674]_ ;
  assign \new_[39676]_  = \new_[39675]_  & \new_[39670]_ ;
  assign \new_[39680]_  = A168 & ~A169;
  assign \new_[39681]_  = ~A170 & \new_[39680]_ ;
  assign \new_[39685]_  = A201 & ~A200;
  assign \new_[39686]_  = A199 & \new_[39685]_ ;
  assign \new_[39687]_  = \new_[39686]_  & \new_[39681]_ ;
  assign \new_[39691]_  = ~A268 & A267;
  assign \new_[39692]_  = A202 & \new_[39691]_ ;
  assign \new_[39696]_  = A299 & A298;
  assign \new_[39697]_  = A269 & \new_[39696]_ ;
  assign \new_[39698]_  = \new_[39697]_  & \new_[39692]_ ;
  assign \new_[39702]_  = A168 & ~A169;
  assign \new_[39703]_  = ~A170 & \new_[39702]_ ;
  assign \new_[39707]_  = A201 & ~A200;
  assign \new_[39708]_  = A199 & \new_[39707]_ ;
  assign \new_[39709]_  = \new_[39708]_  & \new_[39703]_ ;
  assign \new_[39713]_  = ~A268 & A267;
  assign \new_[39714]_  = A202 & \new_[39713]_ ;
  assign \new_[39718]_  = ~A299 & ~A298;
  assign \new_[39719]_  = A269 & \new_[39718]_ ;
  assign \new_[39720]_  = \new_[39719]_  & \new_[39714]_ ;
  assign \new_[39724]_  = A168 & ~A169;
  assign \new_[39725]_  = ~A170 & \new_[39724]_ ;
  assign \new_[39729]_  = A201 & ~A200;
  assign \new_[39730]_  = A199 & \new_[39729]_ ;
  assign \new_[39731]_  = \new_[39730]_  & \new_[39725]_ ;
  assign \new_[39735]_  = A268 & ~A267;
  assign \new_[39736]_  = A202 & \new_[39735]_ ;
  assign \new_[39740]_  = A302 & ~A301;
  assign \new_[39741]_  = A300 & \new_[39740]_ ;
  assign \new_[39742]_  = \new_[39741]_  & \new_[39736]_ ;
  assign \new_[39746]_  = A168 & ~A169;
  assign \new_[39747]_  = ~A170 & \new_[39746]_ ;
  assign \new_[39751]_  = A201 & ~A200;
  assign \new_[39752]_  = A199 & \new_[39751]_ ;
  assign \new_[39753]_  = \new_[39752]_  & \new_[39747]_ ;
  assign \new_[39757]_  = ~A269 & ~A267;
  assign \new_[39758]_  = A202 & \new_[39757]_ ;
  assign \new_[39762]_  = A302 & ~A301;
  assign \new_[39763]_  = A300 & \new_[39762]_ ;
  assign \new_[39764]_  = \new_[39763]_  & \new_[39758]_ ;
  assign \new_[39768]_  = A168 & ~A169;
  assign \new_[39769]_  = ~A170 & \new_[39768]_ ;
  assign \new_[39773]_  = A201 & ~A200;
  assign \new_[39774]_  = A199 & \new_[39773]_ ;
  assign \new_[39775]_  = \new_[39774]_  & \new_[39769]_ ;
  assign \new_[39779]_  = A266 & A265;
  assign \new_[39780]_  = A202 & \new_[39779]_ ;
  assign \new_[39784]_  = A302 & ~A301;
  assign \new_[39785]_  = A300 & \new_[39784]_ ;
  assign \new_[39786]_  = \new_[39785]_  & \new_[39780]_ ;
  assign \new_[39790]_  = A168 & ~A169;
  assign \new_[39791]_  = ~A170 & \new_[39790]_ ;
  assign \new_[39795]_  = A201 & ~A200;
  assign \new_[39796]_  = A199 & \new_[39795]_ ;
  assign \new_[39797]_  = \new_[39796]_  & \new_[39791]_ ;
  assign \new_[39801]_  = ~A266 & ~A265;
  assign \new_[39802]_  = A202 & \new_[39801]_ ;
  assign \new_[39806]_  = A302 & ~A301;
  assign \new_[39807]_  = A300 & \new_[39806]_ ;
  assign \new_[39808]_  = \new_[39807]_  & \new_[39802]_ ;
  assign \new_[39812]_  = A168 & ~A169;
  assign \new_[39813]_  = ~A170 & \new_[39812]_ ;
  assign \new_[39817]_  = A201 & ~A200;
  assign \new_[39818]_  = A199 & \new_[39817]_ ;
  assign \new_[39819]_  = \new_[39818]_  & \new_[39813]_ ;
  assign \new_[39823]_  = ~A268 & A267;
  assign \new_[39824]_  = ~A203 & \new_[39823]_ ;
  assign \new_[39828]_  = A301 & ~A300;
  assign \new_[39829]_  = A269 & \new_[39828]_ ;
  assign \new_[39830]_  = \new_[39829]_  & \new_[39824]_ ;
  assign \new_[39834]_  = A168 & ~A169;
  assign \new_[39835]_  = ~A170 & \new_[39834]_ ;
  assign \new_[39839]_  = A201 & ~A200;
  assign \new_[39840]_  = A199 & \new_[39839]_ ;
  assign \new_[39841]_  = \new_[39840]_  & \new_[39835]_ ;
  assign \new_[39845]_  = ~A268 & A267;
  assign \new_[39846]_  = ~A203 & \new_[39845]_ ;
  assign \new_[39850]_  = ~A302 & ~A300;
  assign \new_[39851]_  = A269 & \new_[39850]_ ;
  assign \new_[39852]_  = \new_[39851]_  & \new_[39846]_ ;
  assign \new_[39856]_  = A168 & ~A169;
  assign \new_[39857]_  = ~A170 & \new_[39856]_ ;
  assign \new_[39861]_  = A201 & ~A200;
  assign \new_[39862]_  = A199 & \new_[39861]_ ;
  assign \new_[39863]_  = \new_[39862]_  & \new_[39857]_ ;
  assign \new_[39867]_  = ~A268 & A267;
  assign \new_[39868]_  = ~A203 & \new_[39867]_ ;
  assign \new_[39872]_  = A299 & A298;
  assign \new_[39873]_  = A269 & \new_[39872]_ ;
  assign \new_[39874]_  = \new_[39873]_  & \new_[39868]_ ;
  assign \new_[39878]_  = A168 & ~A169;
  assign \new_[39879]_  = ~A170 & \new_[39878]_ ;
  assign \new_[39883]_  = A201 & ~A200;
  assign \new_[39884]_  = A199 & \new_[39883]_ ;
  assign \new_[39885]_  = \new_[39884]_  & \new_[39879]_ ;
  assign \new_[39889]_  = ~A268 & A267;
  assign \new_[39890]_  = ~A203 & \new_[39889]_ ;
  assign \new_[39894]_  = ~A299 & ~A298;
  assign \new_[39895]_  = A269 & \new_[39894]_ ;
  assign \new_[39896]_  = \new_[39895]_  & \new_[39890]_ ;
  assign \new_[39900]_  = A168 & ~A169;
  assign \new_[39901]_  = ~A170 & \new_[39900]_ ;
  assign \new_[39905]_  = A201 & ~A200;
  assign \new_[39906]_  = A199 & \new_[39905]_ ;
  assign \new_[39907]_  = \new_[39906]_  & \new_[39901]_ ;
  assign \new_[39911]_  = A268 & ~A267;
  assign \new_[39912]_  = ~A203 & \new_[39911]_ ;
  assign \new_[39916]_  = A302 & ~A301;
  assign \new_[39917]_  = A300 & \new_[39916]_ ;
  assign \new_[39918]_  = \new_[39917]_  & \new_[39912]_ ;
  assign \new_[39922]_  = A168 & ~A169;
  assign \new_[39923]_  = ~A170 & \new_[39922]_ ;
  assign \new_[39927]_  = A201 & ~A200;
  assign \new_[39928]_  = A199 & \new_[39927]_ ;
  assign \new_[39929]_  = \new_[39928]_  & \new_[39923]_ ;
  assign \new_[39933]_  = ~A269 & ~A267;
  assign \new_[39934]_  = ~A203 & \new_[39933]_ ;
  assign \new_[39938]_  = A302 & ~A301;
  assign \new_[39939]_  = A300 & \new_[39938]_ ;
  assign \new_[39940]_  = \new_[39939]_  & \new_[39934]_ ;
  assign \new_[39944]_  = A168 & ~A169;
  assign \new_[39945]_  = ~A170 & \new_[39944]_ ;
  assign \new_[39949]_  = A201 & ~A200;
  assign \new_[39950]_  = A199 & \new_[39949]_ ;
  assign \new_[39951]_  = \new_[39950]_  & \new_[39945]_ ;
  assign \new_[39955]_  = A266 & A265;
  assign \new_[39956]_  = ~A203 & \new_[39955]_ ;
  assign \new_[39960]_  = A302 & ~A301;
  assign \new_[39961]_  = A300 & \new_[39960]_ ;
  assign \new_[39962]_  = \new_[39961]_  & \new_[39956]_ ;
  assign \new_[39966]_  = A168 & ~A169;
  assign \new_[39967]_  = ~A170 & \new_[39966]_ ;
  assign \new_[39971]_  = A201 & ~A200;
  assign \new_[39972]_  = A199 & \new_[39971]_ ;
  assign \new_[39973]_  = \new_[39972]_  & \new_[39967]_ ;
  assign \new_[39977]_  = ~A266 & ~A265;
  assign \new_[39978]_  = ~A203 & \new_[39977]_ ;
  assign \new_[39982]_  = A302 & ~A301;
  assign \new_[39983]_  = A300 & \new_[39982]_ ;
  assign \new_[39984]_  = \new_[39983]_  & \new_[39978]_ ;
  assign \new_[39988]_  = A168 & ~A169;
  assign \new_[39989]_  = ~A170 & \new_[39988]_ ;
  assign \new_[39993]_  = ~A201 & ~A200;
  assign \new_[39994]_  = A199 & \new_[39993]_ ;
  assign \new_[39995]_  = \new_[39994]_  & \new_[39989]_ ;
  assign \new_[39999]_  = ~A267 & A203;
  assign \new_[40000]_  = ~A202 & \new_[39999]_ ;
  assign \new_[40004]_  = A301 & ~A300;
  assign \new_[40005]_  = A268 & \new_[40004]_ ;
  assign \new_[40006]_  = \new_[40005]_  & \new_[40000]_ ;
  assign \new_[40010]_  = A168 & ~A169;
  assign \new_[40011]_  = ~A170 & \new_[40010]_ ;
  assign \new_[40015]_  = ~A201 & ~A200;
  assign \new_[40016]_  = A199 & \new_[40015]_ ;
  assign \new_[40017]_  = \new_[40016]_  & \new_[40011]_ ;
  assign \new_[40021]_  = ~A267 & A203;
  assign \new_[40022]_  = ~A202 & \new_[40021]_ ;
  assign \new_[40026]_  = ~A302 & ~A300;
  assign \new_[40027]_  = A268 & \new_[40026]_ ;
  assign \new_[40028]_  = \new_[40027]_  & \new_[40022]_ ;
  assign \new_[40032]_  = A168 & ~A169;
  assign \new_[40033]_  = ~A170 & \new_[40032]_ ;
  assign \new_[40037]_  = ~A201 & ~A200;
  assign \new_[40038]_  = A199 & \new_[40037]_ ;
  assign \new_[40039]_  = \new_[40038]_  & \new_[40033]_ ;
  assign \new_[40043]_  = ~A267 & A203;
  assign \new_[40044]_  = ~A202 & \new_[40043]_ ;
  assign \new_[40048]_  = A299 & A298;
  assign \new_[40049]_  = A268 & \new_[40048]_ ;
  assign \new_[40050]_  = \new_[40049]_  & \new_[40044]_ ;
  assign \new_[40054]_  = A168 & ~A169;
  assign \new_[40055]_  = ~A170 & \new_[40054]_ ;
  assign \new_[40059]_  = ~A201 & ~A200;
  assign \new_[40060]_  = A199 & \new_[40059]_ ;
  assign \new_[40061]_  = \new_[40060]_  & \new_[40055]_ ;
  assign \new_[40065]_  = ~A267 & A203;
  assign \new_[40066]_  = ~A202 & \new_[40065]_ ;
  assign \new_[40070]_  = ~A299 & ~A298;
  assign \new_[40071]_  = A268 & \new_[40070]_ ;
  assign \new_[40072]_  = \new_[40071]_  & \new_[40066]_ ;
  assign \new_[40076]_  = A168 & ~A169;
  assign \new_[40077]_  = ~A170 & \new_[40076]_ ;
  assign \new_[40081]_  = ~A201 & ~A200;
  assign \new_[40082]_  = A199 & \new_[40081]_ ;
  assign \new_[40083]_  = \new_[40082]_  & \new_[40077]_ ;
  assign \new_[40087]_  = ~A267 & A203;
  assign \new_[40088]_  = ~A202 & \new_[40087]_ ;
  assign \new_[40092]_  = A301 & ~A300;
  assign \new_[40093]_  = ~A269 & \new_[40092]_ ;
  assign \new_[40094]_  = \new_[40093]_  & \new_[40088]_ ;
  assign \new_[40098]_  = A168 & ~A169;
  assign \new_[40099]_  = ~A170 & \new_[40098]_ ;
  assign \new_[40103]_  = ~A201 & ~A200;
  assign \new_[40104]_  = A199 & \new_[40103]_ ;
  assign \new_[40105]_  = \new_[40104]_  & \new_[40099]_ ;
  assign \new_[40109]_  = ~A267 & A203;
  assign \new_[40110]_  = ~A202 & \new_[40109]_ ;
  assign \new_[40114]_  = ~A302 & ~A300;
  assign \new_[40115]_  = ~A269 & \new_[40114]_ ;
  assign \new_[40116]_  = \new_[40115]_  & \new_[40110]_ ;
  assign \new_[40120]_  = A168 & ~A169;
  assign \new_[40121]_  = ~A170 & \new_[40120]_ ;
  assign \new_[40125]_  = ~A201 & ~A200;
  assign \new_[40126]_  = A199 & \new_[40125]_ ;
  assign \new_[40127]_  = \new_[40126]_  & \new_[40121]_ ;
  assign \new_[40131]_  = ~A267 & A203;
  assign \new_[40132]_  = ~A202 & \new_[40131]_ ;
  assign \new_[40136]_  = A299 & A298;
  assign \new_[40137]_  = ~A269 & \new_[40136]_ ;
  assign \new_[40138]_  = \new_[40137]_  & \new_[40132]_ ;
  assign \new_[40142]_  = A168 & ~A169;
  assign \new_[40143]_  = ~A170 & \new_[40142]_ ;
  assign \new_[40147]_  = ~A201 & ~A200;
  assign \new_[40148]_  = A199 & \new_[40147]_ ;
  assign \new_[40149]_  = \new_[40148]_  & \new_[40143]_ ;
  assign \new_[40153]_  = ~A267 & A203;
  assign \new_[40154]_  = ~A202 & \new_[40153]_ ;
  assign \new_[40158]_  = ~A299 & ~A298;
  assign \new_[40159]_  = ~A269 & \new_[40158]_ ;
  assign \new_[40160]_  = \new_[40159]_  & \new_[40154]_ ;
  assign \new_[40164]_  = A168 & ~A169;
  assign \new_[40165]_  = ~A170 & \new_[40164]_ ;
  assign \new_[40169]_  = ~A201 & ~A200;
  assign \new_[40170]_  = A199 & \new_[40169]_ ;
  assign \new_[40171]_  = \new_[40170]_  & \new_[40165]_ ;
  assign \new_[40175]_  = A265 & A203;
  assign \new_[40176]_  = ~A202 & \new_[40175]_ ;
  assign \new_[40180]_  = A301 & ~A300;
  assign \new_[40181]_  = A266 & \new_[40180]_ ;
  assign \new_[40182]_  = \new_[40181]_  & \new_[40176]_ ;
  assign \new_[40186]_  = A168 & ~A169;
  assign \new_[40187]_  = ~A170 & \new_[40186]_ ;
  assign \new_[40191]_  = ~A201 & ~A200;
  assign \new_[40192]_  = A199 & \new_[40191]_ ;
  assign \new_[40193]_  = \new_[40192]_  & \new_[40187]_ ;
  assign \new_[40197]_  = A265 & A203;
  assign \new_[40198]_  = ~A202 & \new_[40197]_ ;
  assign \new_[40202]_  = ~A302 & ~A300;
  assign \new_[40203]_  = A266 & \new_[40202]_ ;
  assign \new_[40204]_  = \new_[40203]_  & \new_[40198]_ ;
  assign \new_[40208]_  = A168 & ~A169;
  assign \new_[40209]_  = ~A170 & \new_[40208]_ ;
  assign \new_[40213]_  = ~A201 & ~A200;
  assign \new_[40214]_  = A199 & \new_[40213]_ ;
  assign \new_[40215]_  = \new_[40214]_  & \new_[40209]_ ;
  assign \new_[40219]_  = A265 & A203;
  assign \new_[40220]_  = ~A202 & \new_[40219]_ ;
  assign \new_[40224]_  = A299 & A298;
  assign \new_[40225]_  = A266 & \new_[40224]_ ;
  assign \new_[40226]_  = \new_[40225]_  & \new_[40220]_ ;
  assign \new_[40230]_  = A168 & ~A169;
  assign \new_[40231]_  = ~A170 & \new_[40230]_ ;
  assign \new_[40235]_  = ~A201 & ~A200;
  assign \new_[40236]_  = A199 & \new_[40235]_ ;
  assign \new_[40237]_  = \new_[40236]_  & \new_[40231]_ ;
  assign \new_[40241]_  = A265 & A203;
  assign \new_[40242]_  = ~A202 & \new_[40241]_ ;
  assign \new_[40246]_  = ~A299 & ~A298;
  assign \new_[40247]_  = A266 & \new_[40246]_ ;
  assign \new_[40248]_  = \new_[40247]_  & \new_[40242]_ ;
  assign \new_[40252]_  = A168 & ~A169;
  assign \new_[40253]_  = ~A170 & \new_[40252]_ ;
  assign \new_[40257]_  = ~A201 & ~A200;
  assign \new_[40258]_  = A199 & \new_[40257]_ ;
  assign \new_[40259]_  = \new_[40258]_  & \new_[40253]_ ;
  assign \new_[40263]_  = ~A265 & A203;
  assign \new_[40264]_  = ~A202 & \new_[40263]_ ;
  assign \new_[40268]_  = A301 & ~A300;
  assign \new_[40269]_  = ~A266 & \new_[40268]_ ;
  assign \new_[40270]_  = \new_[40269]_  & \new_[40264]_ ;
  assign \new_[40274]_  = A168 & ~A169;
  assign \new_[40275]_  = ~A170 & \new_[40274]_ ;
  assign \new_[40279]_  = ~A201 & ~A200;
  assign \new_[40280]_  = A199 & \new_[40279]_ ;
  assign \new_[40281]_  = \new_[40280]_  & \new_[40275]_ ;
  assign \new_[40285]_  = ~A265 & A203;
  assign \new_[40286]_  = ~A202 & \new_[40285]_ ;
  assign \new_[40290]_  = ~A302 & ~A300;
  assign \new_[40291]_  = ~A266 & \new_[40290]_ ;
  assign \new_[40292]_  = \new_[40291]_  & \new_[40286]_ ;
  assign \new_[40296]_  = A168 & ~A169;
  assign \new_[40297]_  = ~A170 & \new_[40296]_ ;
  assign \new_[40301]_  = ~A201 & ~A200;
  assign \new_[40302]_  = A199 & \new_[40301]_ ;
  assign \new_[40303]_  = \new_[40302]_  & \new_[40297]_ ;
  assign \new_[40307]_  = ~A265 & A203;
  assign \new_[40308]_  = ~A202 & \new_[40307]_ ;
  assign \new_[40312]_  = A299 & A298;
  assign \new_[40313]_  = ~A266 & \new_[40312]_ ;
  assign \new_[40314]_  = \new_[40313]_  & \new_[40308]_ ;
  assign \new_[40318]_  = A168 & ~A169;
  assign \new_[40319]_  = ~A170 & \new_[40318]_ ;
  assign \new_[40323]_  = ~A201 & ~A200;
  assign \new_[40324]_  = A199 & \new_[40323]_ ;
  assign \new_[40325]_  = \new_[40324]_  & \new_[40319]_ ;
  assign \new_[40329]_  = ~A265 & A203;
  assign \new_[40330]_  = ~A202 & \new_[40329]_ ;
  assign \new_[40334]_  = ~A299 & ~A298;
  assign \new_[40335]_  = ~A266 & \new_[40334]_ ;
  assign \new_[40336]_  = \new_[40335]_  & \new_[40330]_ ;
  assign \new_[40340]_  = A202 & A200;
  assign \new_[40341]_  = ~A199 & \new_[40340]_ ;
  assign \new_[40345]_  = ~A234 & A233;
  assign \new_[40346]_  = ~A232 & \new_[40345]_ ;
  assign \new_[40347]_  = \new_[40346]_  & \new_[40341]_ ;
  assign \new_[40351]_  = ~A265 & A236;
  assign \new_[40352]_  = ~A235 & \new_[40351]_ ;
  assign \new_[40355]_  = ~A267 & A266;
  assign \new_[40358]_  = A269 & ~A268;
  assign \new_[40359]_  = \new_[40358]_  & \new_[40355]_ ;
  assign \new_[40360]_  = \new_[40359]_  & \new_[40352]_ ;
  assign \new_[40364]_  = A202 & A200;
  assign \new_[40365]_  = ~A199 & \new_[40364]_ ;
  assign \new_[40369]_  = ~A234 & A233;
  assign \new_[40370]_  = ~A232 & \new_[40369]_ ;
  assign \new_[40371]_  = \new_[40370]_  & \new_[40365]_ ;
  assign \new_[40375]_  = A265 & A236;
  assign \new_[40376]_  = ~A235 & \new_[40375]_ ;
  assign \new_[40379]_  = ~A267 & ~A266;
  assign \new_[40382]_  = A269 & ~A268;
  assign \new_[40383]_  = \new_[40382]_  & \new_[40379]_ ;
  assign \new_[40384]_  = \new_[40383]_  & \new_[40376]_ ;
  assign \new_[40388]_  = A202 & A200;
  assign \new_[40389]_  = ~A199 & \new_[40388]_ ;
  assign \new_[40393]_  = ~A234 & ~A233;
  assign \new_[40394]_  = A232 & \new_[40393]_ ;
  assign \new_[40395]_  = \new_[40394]_  & \new_[40389]_ ;
  assign \new_[40399]_  = ~A265 & A236;
  assign \new_[40400]_  = ~A235 & \new_[40399]_ ;
  assign \new_[40403]_  = ~A267 & A266;
  assign \new_[40406]_  = A269 & ~A268;
  assign \new_[40407]_  = \new_[40406]_  & \new_[40403]_ ;
  assign \new_[40408]_  = \new_[40407]_  & \new_[40400]_ ;
  assign \new_[40412]_  = A202 & A200;
  assign \new_[40413]_  = ~A199 & \new_[40412]_ ;
  assign \new_[40417]_  = ~A234 & ~A233;
  assign \new_[40418]_  = A232 & \new_[40417]_ ;
  assign \new_[40419]_  = \new_[40418]_  & \new_[40413]_ ;
  assign \new_[40423]_  = A265 & A236;
  assign \new_[40424]_  = ~A235 & \new_[40423]_ ;
  assign \new_[40427]_  = ~A267 & ~A266;
  assign \new_[40430]_  = A269 & ~A268;
  assign \new_[40431]_  = \new_[40430]_  & \new_[40427]_ ;
  assign \new_[40432]_  = \new_[40431]_  & \new_[40424]_ ;
  assign \new_[40436]_  = ~A203 & A200;
  assign \new_[40437]_  = ~A199 & \new_[40436]_ ;
  assign \new_[40441]_  = ~A234 & A233;
  assign \new_[40442]_  = ~A232 & \new_[40441]_ ;
  assign \new_[40443]_  = \new_[40442]_  & \new_[40437]_ ;
  assign \new_[40447]_  = ~A265 & A236;
  assign \new_[40448]_  = ~A235 & \new_[40447]_ ;
  assign \new_[40451]_  = ~A267 & A266;
  assign \new_[40454]_  = A269 & ~A268;
  assign \new_[40455]_  = \new_[40454]_  & \new_[40451]_ ;
  assign \new_[40456]_  = \new_[40455]_  & \new_[40448]_ ;
  assign \new_[40460]_  = ~A203 & A200;
  assign \new_[40461]_  = ~A199 & \new_[40460]_ ;
  assign \new_[40465]_  = ~A234 & A233;
  assign \new_[40466]_  = ~A232 & \new_[40465]_ ;
  assign \new_[40467]_  = \new_[40466]_  & \new_[40461]_ ;
  assign \new_[40471]_  = A265 & A236;
  assign \new_[40472]_  = ~A235 & \new_[40471]_ ;
  assign \new_[40475]_  = ~A267 & ~A266;
  assign \new_[40478]_  = A269 & ~A268;
  assign \new_[40479]_  = \new_[40478]_  & \new_[40475]_ ;
  assign \new_[40480]_  = \new_[40479]_  & \new_[40472]_ ;
  assign \new_[40484]_  = ~A203 & A200;
  assign \new_[40485]_  = ~A199 & \new_[40484]_ ;
  assign \new_[40489]_  = ~A234 & ~A233;
  assign \new_[40490]_  = A232 & \new_[40489]_ ;
  assign \new_[40491]_  = \new_[40490]_  & \new_[40485]_ ;
  assign \new_[40495]_  = ~A265 & A236;
  assign \new_[40496]_  = ~A235 & \new_[40495]_ ;
  assign \new_[40499]_  = ~A267 & A266;
  assign \new_[40502]_  = A269 & ~A268;
  assign \new_[40503]_  = \new_[40502]_  & \new_[40499]_ ;
  assign \new_[40504]_  = \new_[40503]_  & \new_[40496]_ ;
  assign \new_[40508]_  = ~A203 & A200;
  assign \new_[40509]_  = ~A199 & \new_[40508]_ ;
  assign \new_[40513]_  = ~A234 & ~A233;
  assign \new_[40514]_  = A232 & \new_[40513]_ ;
  assign \new_[40515]_  = \new_[40514]_  & \new_[40509]_ ;
  assign \new_[40519]_  = A265 & A236;
  assign \new_[40520]_  = ~A235 & \new_[40519]_ ;
  assign \new_[40523]_  = ~A267 & ~A266;
  assign \new_[40526]_  = A269 & ~A268;
  assign \new_[40527]_  = \new_[40526]_  & \new_[40523]_ ;
  assign \new_[40528]_  = \new_[40527]_  & \new_[40520]_ ;
  assign \new_[40532]_  = A202 & ~A200;
  assign \new_[40533]_  = A199 & \new_[40532]_ ;
  assign \new_[40537]_  = ~A234 & A233;
  assign \new_[40538]_  = ~A232 & \new_[40537]_ ;
  assign \new_[40539]_  = \new_[40538]_  & \new_[40533]_ ;
  assign \new_[40543]_  = ~A265 & A236;
  assign \new_[40544]_  = ~A235 & \new_[40543]_ ;
  assign \new_[40547]_  = ~A267 & A266;
  assign \new_[40550]_  = A269 & ~A268;
  assign \new_[40551]_  = \new_[40550]_  & \new_[40547]_ ;
  assign \new_[40552]_  = \new_[40551]_  & \new_[40544]_ ;
  assign \new_[40556]_  = A202 & ~A200;
  assign \new_[40557]_  = A199 & \new_[40556]_ ;
  assign \new_[40561]_  = ~A234 & A233;
  assign \new_[40562]_  = ~A232 & \new_[40561]_ ;
  assign \new_[40563]_  = \new_[40562]_  & \new_[40557]_ ;
  assign \new_[40567]_  = A265 & A236;
  assign \new_[40568]_  = ~A235 & \new_[40567]_ ;
  assign \new_[40571]_  = ~A267 & ~A266;
  assign \new_[40574]_  = A269 & ~A268;
  assign \new_[40575]_  = \new_[40574]_  & \new_[40571]_ ;
  assign \new_[40576]_  = \new_[40575]_  & \new_[40568]_ ;
  assign \new_[40580]_  = A202 & ~A200;
  assign \new_[40581]_  = A199 & \new_[40580]_ ;
  assign \new_[40585]_  = ~A234 & ~A233;
  assign \new_[40586]_  = A232 & \new_[40585]_ ;
  assign \new_[40587]_  = \new_[40586]_  & \new_[40581]_ ;
  assign \new_[40591]_  = ~A265 & A236;
  assign \new_[40592]_  = ~A235 & \new_[40591]_ ;
  assign \new_[40595]_  = ~A267 & A266;
  assign \new_[40598]_  = A269 & ~A268;
  assign \new_[40599]_  = \new_[40598]_  & \new_[40595]_ ;
  assign \new_[40600]_  = \new_[40599]_  & \new_[40592]_ ;
  assign \new_[40604]_  = A202 & ~A200;
  assign \new_[40605]_  = A199 & \new_[40604]_ ;
  assign \new_[40609]_  = ~A234 & ~A233;
  assign \new_[40610]_  = A232 & \new_[40609]_ ;
  assign \new_[40611]_  = \new_[40610]_  & \new_[40605]_ ;
  assign \new_[40615]_  = A265 & A236;
  assign \new_[40616]_  = ~A235 & \new_[40615]_ ;
  assign \new_[40619]_  = ~A267 & ~A266;
  assign \new_[40622]_  = A269 & ~A268;
  assign \new_[40623]_  = \new_[40622]_  & \new_[40619]_ ;
  assign \new_[40624]_  = \new_[40623]_  & \new_[40616]_ ;
  assign \new_[40628]_  = ~A203 & ~A200;
  assign \new_[40629]_  = A199 & \new_[40628]_ ;
  assign \new_[40633]_  = ~A234 & A233;
  assign \new_[40634]_  = ~A232 & \new_[40633]_ ;
  assign \new_[40635]_  = \new_[40634]_  & \new_[40629]_ ;
  assign \new_[40639]_  = ~A265 & A236;
  assign \new_[40640]_  = ~A235 & \new_[40639]_ ;
  assign \new_[40643]_  = ~A267 & A266;
  assign \new_[40646]_  = A269 & ~A268;
  assign \new_[40647]_  = \new_[40646]_  & \new_[40643]_ ;
  assign \new_[40648]_  = \new_[40647]_  & \new_[40640]_ ;
  assign \new_[40652]_  = ~A203 & ~A200;
  assign \new_[40653]_  = A199 & \new_[40652]_ ;
  assign \new_[40657]_  = ~A234 & A233;
  assign \new_[40658]_  = ~A232 & \new_[40657]_ ;
  assign \new_[40659]_  = \new_[40658]_  & \new_[40653]_ ;
  assign \new_[40663]_  = A265 & A236;
  assign \new_[40664]_  = ~A235 & \new_[40663]_ ;
  assign \new_[40667]_  = ~A267 & ~A266;
  assign \new_[40670]_  = A269 & ~A268;
  assign \new_[40671]_  = \new_[40670]_  & \new_[40667]_ ;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40664]_ ;
  assign \new_[40676]_  = ~A203 & ~A200;
  assign \new_[40677]_  = A199 & \new_[40676]_ ;
  assign \new_[40681]_  = ~A234 & ~A233;
  assign \new_[40682]_  = A232 & \new_[40681]_ ;
  assign \new_[40683]_  = \new_[40682]_  & \new_[40677]_ ;
  assign \new_[40687]_  = ~A265 & A236;
  assign \new_[40688]_  = ~A235 & \new_[40687]_ ;
  assign \new_[40691]_  = ~A267 & A266;
  assign \new_[40694]_  = A269 & ~A268;
  assign \new_[40695]_  = \new_[40694]_  & \new_[40691]_ ;
  assign \new_[40696]_  = \new_[40695]_  & \new_[40688]_ ;
  assign \new_[40700]_  = ~A203 & ~A200;
  assign \new_[40701]_  = A199 & \new_[40700]_ ;
  assign \new_[40705]_  = ~A234 & ~A233;
  assign \new_[40706]_  = A232 & \new_[40705]_ ;
  assign \new_[40707]_  = \new_[40706]_  & \new_[40701]_ ;
  assign \new_[40711]_  = A265 & A236;
  assign \new_[40712]_  = ~A235 & \new_[40711]_ ;
  assign \new_[40715]_  = ~A267 & ~A266;
  assign \new_[40718]_  = A269 & ~A268;
  assign \new_[40719]_  = \new_[40718]_  & \new_[40715]_ ;
  assign \new_[40720]_  = \new_[40719]_  & \new_[40712]_ ;
  assign \new_[40724]_  = ~A199 & A166;
  assign \new_[40725]_  = A167 & \new_[40724]_ ;
  assign \new_[40729]_  = ~A202 & ~A201;
  assign \new_[40730]_  = A200 & \new_[40729]_ ;
  assign \new_[40731]_  = \new_[40730]_  & \new_[40725]_ ;
  assign \new_[40735]_  = ~A268 & A267;
  assign \new_[40736]_  = A203 & \new_[40735]_ ;
  assign \new_[40739]_  = A300 & A269;
  assign \new_[40742]_  = A302 & ~A301;
  assign \new_[40743]_  = \new_[40742]_  & \new_[40739]_ ;
  assign \new_[40744]_  = \new_[40743]_  & \new_[40736]_ ;
  assign \new_[40748]_  = A199 & A166;
  assign \new_[40749]_  = A167 & \new_[40748]_ ;
  assign \new_[40753]_  = ~A202 & ~A201;
  assign \new_[40754]_  = ~A200 & \new_[40753]_ ;
  assign \new_[40755]_  = \new_[40754]_  & \new_[40749]_ ;
  assign \new_[40759]_  = ~A268 & A267;
  assign \new_[40760]_  = A203 & \new_[40759]_ ;
  assign \new_[40763]_  = A300 & A269;
  assign \new_[40766]_  = A302 & ~A301;
  assign \new_[40767]_  = \new_[40766]_  & \new_[40763]_ ;
  assign \new_[40768]_  = \new_[40767]_  & \new_[40760]_ ;
  assign \new_[40772]_  = ~A199 & ~A166;
  assign \new_[40773]_  = ~A167 & \new_[40772]_ ;
  assign \new_[40777]_  = ~A202 & ~A201;
  assign \new_[40778]_  = A200 & \new_[40777]_ ;
  assign \new_[40779]_  = \new_[40778]_  & \new_[40773]_ ;
  assign \new_[40783]_  = ~A268 & A267;
  assign \new_[40784]_  = A203 & \new_[40783]_ ;
  assign \new_[40787]_  = A300 & A269;
  assign \new_[40790]_  = A302 & ~A301;
  assign \new_[40791]_  = \new_[40790]_  & \new_[40787]_ ;
  assign \new_[40792]_  = \new_[40791]_  & \new_[40784]_ ;
  assign \new_[40796]_  = A199 & ~A166;
  assign \new_[40797]_  = ~A167 & \new_[40796]_ ;
  assign \new_[40801]_  = ~A202 & ~A201;
  assign \new_[40802]_  = ~A200 & \new_[40801]_ ;
  assign \new_[40803]_  = \new_[40802]_  & \new_[40797]_ ;
  assign \new_[40807]_  = ~A268 & A267;
  assign \new_[40808]_  = A203 & \new_[40807]_ ;
  assign \new_[40811]_  = A300 & A269;
  assign \new_[40814]_  = A302 & ~A301;
  assign \new_[40815]_  = \new_[40814]_  & \new_[40811]_ ;
  assign \new_[40816]_  = \new_[40815]_  & \new_[40808]_ ;
  assign \new_[40820]_  = A200 & ~A199;
  assign \new_[40821]_  = A170 & \new_[40820]_ ;
  assign \new_[40825]_  = ~A234 & A233;
  assign \new_[40826]_  = ~A232 & \new_[40825]_ ;
  assign \new_[40827]_  = \new_[40826]_  & \new_[40821]_ ;
  assign \new_[40831]_  = ~A265 & A236;
  assign \new_[40832]_  = ~A235 & \new_[40831]_ ;
  assign \new_[40835]_  = ~A267 & A266;
  assign \new_[40838]_  = A269 & ~A268;
  assign \new_[40839]_  = \new_[40838]_  & \new_[40835]_ ;
  assign \new_[40840]_  = \new_[40839]_  & \new_[40832]_ ;
  assign \new_[40844]_  = A200 & ~A199;
  assign \new_[40845]_  = A170 & \new_[40844]_ ;
  assign \new_[40849]_  = ~A234 & A233;
  assign \new_[40850]_  = ~A232 & \new_[40849]_ ;
  assign \new_[40851]_  = \new_[40850]_  & \new_[40845]_ ;
  assign \new_[40855]_  = A265 & A236;
  assign \new_[40856]_  = ~A235 & \new_[40855]_ ;
  assign \new_[40859]_  = ~A267 & ~A266;
  assign \new_[40862]_  = A269 & ~A268;
  assign \new_[40863]_  = \new_[40862]_  & \new_[40859]_ ;
  assign \new_[40864]_  = \new_[40863]_  & \new_[40856]_ ;
  assign \new_[40868]_  = A200 & ~A199;
  assign \new_[40869]_  = A170 & \new_[40868]_ ;
  assign \new_[40873]_  = ~A234 & ~A233;
  assign \new_[40874]_  = A232 & \new_[40873]_ ;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40869]_ ;
  assign \new_[40879]_  = ~A265 & A236;
  assign \new_[40880]_  = ~A235 & \new_[40879]_ ;
  assign \new_[40883]_  = ~A267 & A266;
  assign \new_[40886]_  = A269 & ~A268;
  assign \new_[40887]_  = \new_[40886]_  & \new_[40883]_ ;
  assign \new_[40888]_  = \new_[40887]_  & \new_[40880]_ ;
  assign \new_[40892]_  = A200 & ~A199;
  assign \new_[40893]_  = A170 & \new_[40892]_ ;
  assign \new_[40897]_  = ~A234 & ~A233;
  assign \new_[40898]_  = A232 & \new_[40897]_ ;
  assign \new_[40899]_  = \new_[40898]_  & \new_[40893]_ ;
  assign \new_[40903]_  = A265 & A236;
  assign \new_[40904]_  = ~A235 & \new_[40903]_ ;
  assign \new_[40907]_  = ~A267 & ~A266;
  assign \new_[40910]_  = A269 & ~A268;
  assign \new_[40911]_  = \new_[40910]_  & \new_[40907]_ ;
  assign \new_[40912]_  = \new_[40911]_  & \new_[40904]_ ;
  assign \new_[40916]_  = ~A200 & A199;
  assign \new_[40917]_  = A170 & \new_[40916]_ ;
  assign \new_[40921]_  = ~A234 & A233;
  assign \new_[40922]_  = ~A232 & \new_[40921]_ ;
  assign \new_[40923]_  = \new_[40922]_  & \new_[40917]_ ;
  assign \new_[40927]_  = ~A265 & A236;
  assign \new_[40928]_  = ~A235 & \new_[40927]_ ;
  assign \new_[40931]_  = ~A267 & A266;
  assign \new_[40934]_  = A269 & ~A268;
  assign \new_[40935]_  = \new_[40934]_  & \new_[40931]_ ;
  assign \new_[40936]_  = \new_[40935]_  & \new_[40928]_ ;
  assign \new_[40940]_  = ~A200 & A199;
  assign \new_[40941]_  = A170 & \new_[40940]_ ;
  assign \new_[40945]_  = ~A234 & A233;
  assign \new_[40946]_  = ~A232 & \new_[40945]_ ;
  assign \new_[40947]_  = \new_[40946]_  & \new_[40941]_ ;
  assign \new_[40951]_  = A265 & A236;
  assign \new_[40952]_  = ~A235 & \new_[40951]_ ;
  assign \new_[40955]_  = ~A267 & ~A266;
  assign \new_[40958]_  = A269 & ~A268;
  assign \new_[40959]_  = \new_[40958]_  & \new_[40955]_ ;
  assign \new_[40960]_  = \new_[40959]_  & \new_[40952]_ ;
  assign \new_[40964]_  = ~A200 & A199;
  assign \new_[40965]_  = A170 & \new_[40964]_ ;
  assign \new_[40969]_  = ~A234 & ~A233;
  assign \new_[40970]_  = A232 & \new_[40969]_ ;
  assign \new_[40971]_  = \new_[40970]_  & \new_[40965]_ ;
  assign \new_[40975]_  = ~A265 & A236;
  assign \new_[40976]_  = ~A235 & \new_[40975]_ ;
  assign \new_[40979]_  = ~A267 & A266;
  assign \new_[40982]_  = A269 & ~A268;
  assign \new_[40983]_  = \new_[40982]_  & \new_[40979]_ ;
  assign \new_[40984]_  = \new_[40983]_  & \new_[40976]_ ;
  assign \new_[40988]_  = ~A200 & A199;
  assign \new_[40989]_  = A170 & \new_[40988]_ ;
  assign \new_[40993]_  = ~A234 & ~A233;
  assign \new_[40994]_  = A232 & \new_[40993]_ ;
  assign \new_[40995]_  = \new_[40994]_  & \new_[40989]_ ;
  assign \new_[40999]_  = A265 & A236;
  assign \new_[41000]_  = ~A235 & \new_[40999]_ ;
  assign \new_[41003]_  = ~A267 & ~A266;
  assign \new_[41006]_  = A269 & ~A268;
  assign \new_[41007]_  = \new_[41006]_  & \new_[41003]_ ;
  assign \new_[41008]_  = \new_[41007]_  & \new_[41000]_ ;
  assign \new_[41012]_  = A167 & A168;
  assign \new_[41013]_  = A170 & \new_[41012]_ ;
  assign \new_[41017]_  = ~A202 & A201;
  assign \new_[41018]_  = ~A166 & \new_[41017]_ ;
  assign \new_[41019]_  = \new_[41018]_  & \new_[41013]_ ;
  assign \new_[41023]_  = A268 & ~A267;
  assign \new_[41024]_  = A203 & \new_[41023]_ ;
  assign \new_[41027]_  = ~A299 & A298;
  assign \new_[41030]_  = A301 & A300;
  assign \new_[41031]_  = \new_[41030]_  & \new_[41027]_ ;
  assign \new_[41032]_  = \new_[41031]_  & \new_[41024]_ ;
  assign \new_[41036]_  = A167 & A168;
  assign \new_[41037]_  = A170 & \new_[41036]_ ;
  assign \new_[41041]_  = ~A202 & A201;
  assign \new_[41042]_  = ~A166 & \new_[41041]_ ;
  assign \new_[41043]_  = \new_[41042]_  & \new_[41037]_ ;
  assign \new_[41047]_  = A268 & ~A267;
  assign \new_[41048]_  = A203 & \new_[41047]_ ;
  assign \new_[41051]_  = ~A299 & A298;
  assign \new_[41054]_  = ~A302 & A300;
  assign \new_[41055]_  = \new_[41054]_  & \new_[41051]_ ;
  assign \new_[41056]_  = \new_[41055]_  & \new_[41048]_ ;
  assign \new_[41060]_  = A167 & A168;
  assign \new_[41061]_  = A170 & \new_[41060]_ ;
  assign \new_[41065]_  = ~A202 & A201;
  assign \new_[41066]_  = ~A166 & \new_[41065]_ ;
  assign \new_[41067]_  = \new_[41066]_  & \new_[41061]_ ;
  assign \new_[41071]_  = A268 & ~A267;
  assign \new_[41072]_  = A203 & \new_[41071]_ ;
  assign \new_[41075]_  = A299 & ~A298;
  assign \new_[41078]_  = A301 & A300;
  assign \new_[41079]_  = \new_[41078]_  & \new_[41075]_ ;
  assign \new_[41080]_  = \new_[41079]_  & \new_[41072]_ ;
  assign \new_[41084]_  = A167 & A168;
  assign \new_[41085]_  = A170 & \new_[41084]_ ;
  assign \new_[41089]_  = ~A202 & A201;
  assign \new_[41090]_  = ~A166 & \new_[41089]_ ;
  assign \new_[41091]_  = \new_[41090]_  & \new_[41085]_ ;
  assign \new_[41095]_  = A268 & ~A267;
  assign \new_[41096]_  = A203 & \new_[41095]_ ;
  assign \new_[41099]_  = A299 & ~A298;
  assign \new_[41102]_  = ~A302 & A300;
  assign \new_[41103]_  = \new_[41102]_  & \new_[41099]_ ;
  assign \new_[41104]_  = \new_[41103]_  & \new_[41096]_ ;
  assign \new_[41108]_  = A167 & A168;
  assign \new_[41109]_  = A170 & \new_[41108]_ ;
  assign \new_[41113]_  = ~A202 & A201;
  assign \new_[41114]_  = ~A166 & \new_[41113]_ ;
  assign \new_[41115]_  = \new_[41114]_  & \new_[41109]_ ;
  assign \new_[41119]_  = ~A269 & ~A267;
  assign \new_[41120]_  = A203 & \new_[41119]_ ;
  assign \new_[41123]_  = ~A299 & A298;
  assign \new_[41126]_  = A301 & A300;
  assign \new_[41127]_  = \new_[41126]_  & \new_[41123]_ ;
  assign \new_[41128]_  = \new_[41127]_  & \new_[41120]_ ;
  assign \new_[41132]_  = A167 & A168;
  assign \new_[41133]_  = A170 & \new_[41132]_ ;
  assign \new_[41137]_  = ~A202 & A201;
  assign \new_[41138]_  = ~A166 & \new_[41137]_ ;
  assign \new_[41139]_  = \new_[41138]_  & \new_[41133]_ ;
  assign \new_[41143]_  = ~A269 & ~A267;
  assign \new_[41144]_  = A203 & \new_[41143]_ ;
  assign \new_[41147]_  = ~A299 & A298;
  assign \new_[41150]_  = ~A302 & A300;
  assign \new_[41151]_  = \new_[41150]_  & \new_[41147]_ ;
  assign \new_[41152]_  = \new_[41151]_  & \new_[41144]_ ;
  assign \new_[41156]_  = A167 & A168;
  assign \new_[41157]_  = A170 & \new_[41156]_ ;
  assign \new_[41161]_  = ~A202 & A201;
  assign \new_[41162]_  = ~A166 & \new_[41161]_ ;
  assign \new_[41163]_  = \new_[41162]_  & \new_[41157]_ ;
  assign \new_[41167]_  = ~A269 & ~A267;
  assign \new_[41168]_  = A203 & \new_[41167]_ ;
  assign \new_[41171]_  = A299 & ~A298;
  assign \new_[41174]_  = A301 & A300;
  assign \new_[41175]_  = \new_[41174]_  & \new_[41171]_ ;
  assign \new_[41176]_  = \new_[41175]_  & \new_[41168]_ ;
  assign \new_[41180]_  = A167 & A168;
  assign \new_[41181]_  = A170 & \new_[41180]_ ;
  assign \new_[41185]_  = ~A202 & A201;
  assign \new_[41186]_  = ~A166 & \new_[41185]_ ;
  assign \new_[41187]_  = \new_[41186]_  & \new_[41181]_ ;
  assign \new_[41191]_  = ~A269 & ~A267;
  assign \new_[41192]_  = A203 & \new_[41191]_ ;
  assign \new_[41195]_  = A299 & ~A298;
  assign \new_[41198]_  = ~A302 & A300;
  assign \new_[41199]_  = \new_[41198]_  & \new_[41195]_ ;
  assign \new_[41200]_  = \new_[41199]_  & \new_[41192]_ ;
  assign \new_[41204]_  = A167 & A168;
  assign \new_[41205]_  = A170 & \new_[41204]_ ;
  assign \new_[41209]_  = ~A202 & A201;
  assign \new_[41210]_  = ~A166 & \new_[41209]_ ;
  assign \new_[41211]_  = \new_[41210]_  & \new_[41205]_ ;
  assign \new_[41215]_  = A266 & A265;
  assign \new_[41216]_  = A203 & \new_[41215]_ ;
  assign \new_[41219]_  = ~A299 & A298;
  assign \new_[41222]_  = A301 & A300;
  assign \new_[41223]_  = \new_[41222]_  & \new_[41219]_ ;
  assign \new_[41224]_  = \new_[41223]_  & \new_[41216]_ ;
  assign \new_[41228]_  = A167 & A168;
  assign \new_[41229]_  = A170 & \new_[41228]_ ;
  assign \new_[41233]_  = ~A202 & A201;
  assign \new_[41234]_  = ~A166 & \new_[41233]_ ;
  assign \new_[41235]_  = \new_[41234]_  & \new_[41229]_ ;
  assign \new_[41239]_  = A266 & A265;
  assign \new_[41240]_  = A203 & \new_[41239]_ ;
  assign \new_[41243]_  = ~A299 & A298;
  assign \new_[41246]_  = ~A302 & A300;
  assign \new_[41247]_  = \new_[41246]_  & \new_[41243]_ ;
  assign \new_[41248]_  = \new_[41247]_  & \new_[41240]_ ;
  assign \new_[41252]_  = A167 & A168;
  assign \new_[41253]_  = A170 & \new_[41252]_ ;
  assign \new_[41257]_  = ~A202 & A201;
  assign \new_[41258]_  = ~A166 & \new_[41257]_ ;
  assign \new_[41259]_  = \new_[41258]_  & \new_[41253]_ ;
  assign \new_[41263]_  = A266 & A265;
  assign \new_[41264]_  = A203 & \new_[41263]_ ;
  assign \new_[41267]_  = A299 & ~A298;
  assign \new_[41270]_  = A301 & A300;
  assign \new_[41271]_  = \new_[41270]_  & \new_[41267]_ ;
  assign \new_[41272]_  = \new_[41271]_  & \new_[41264]_ ;
  assign \new_[41276]_  = A167 & A168;
  assign \new_[41277]_  = A170 & \new_[41276]_ ;
  assign \new_[41281]_  = ~A202 & A201;
  assign \new_[41282]_  = ~A166 & \new_[41281]_ ;
  assign \new_[41283]_  = \new_[41282]_  & \new_[41277]_ ;
  assign \new_[41287]_  = A266 & A265;
  assign \new_[41288]_  = A203 & \new_[41287]_ ;
  assign \new_[41291]_  = A299 & ~A298;
  assign \new_[41294]_  = ~A302 & A300;
  assign \new_[41295]_  = \new_[41294]_  & \new_[41291]_ ;
  assign \new_[41296]_  = \new_[41295]_  & \new_[41288]_ ;
  assign \new_[41300]_  = A167 & A168;
  assign \new_[41301]_  = A170 & \new_[41300]_ ;
  assign \new_[41305]_  = ~A202 & A201;
  assign \new_[41306]_  = ~A166 & \new_[41305]_ ;
  assign \new_[41307]_  = \new_[41306]_  & \new_[41301]_ ;
  assign \new_[41311]_  = A266 & ~A265;
  assign \new_[41312]_  = A203 & \new_[41311]_ ;
  assign \new_[41315]_  = A268 & A267;
  assign \new_[41318]_  = A301 & ~A300;
  assign \new_[41319]_  = \new_[41318]_  & \new_[41315]_ ;
  assign \new_[41320]_  = \new_[41319]_  & \new_[41312]_ ;
  assign \new_[41324]_  = A167 & A168;
  assign \new_[41325]_  = A170 & \new_[41324]_ ;
  assign \new_[41329]_  = ~A202 & A201;
  assign \new_[41330]_  = ~A166 & \new_[41329]_ ;
  assign \new_[41331]_  = \new_[41330]_  & \new_[41325]_ ;
  assign \new_[41335]_  = A266 & ~A265;
  assign \new_[41336]_  = A203 & \new_[41335]_ ;
  assign \new_[41339]_  = A268 & A267;
  assign \new_[41342]_  = ~A302 & ~A300;
  assign \new_[41343]_  = \new_[41342]_  & \new_[41339]_ ;
  assign \new_[41344]_  = \new_[41343]_  & \new_[41336]_ ;
  assign \new_[41348]_  = A167 & A168;
  assign \new_[41349]_  = A170 & \new_[41348]_ ;
  assign \new_[41353]_  = ~A202 & A201;
  assign \new_[41354]_  = ~A166 & \new_[41353]_ ;
  assign \new_[41355]_  = \new_[41354]_  & \new_[41349]_ ;
  assign \new_[41359]_  = A266 & ~A265;
  assign \new_[41360]_  = A203 & \new_[41359]_ ;
  assign \new_[41363]_  = A268 & A267;
  assign \new_[41366]_  = A299 & A298;
  assign \new_[41367]_  = \new_[41366]_  & \new_[41363]_ ;
  assign \new_[41368]_  = \new_[41367]_  & \new_[41360]_ ;
  assign \new_[41372]_  = A167 & A168;
  assign \new_[41373]_  = A170 & \new_[41372]_ ;
  assign \new_[41377]_  = ~A202 & A201;
  assign \new_[41378]_  = ~A166 & \new_[41377]_ ;
  assign \new_[41379]_  = \new_[41378]_  & \new_[41373]_ ;
  assign \new_[41383]_  = A266 & ~A265;
  assign \new_[41384]_  = A203 & \new_[41383]_ ;
  assign \new_[41387]_  = A268 & A267;
  assign \new_[41390]_  = ~A299 & ~A298;
  assign \new_[41391]_  = \new_[41390]_  & \new_[41387]_ ;
  assign \new_[41392]_  = \new_[41391]_  & \new_[41384]_ ;
  assign \new_[41396]_  = A167 & A168;
  assign \new_[41397]_  = A170 & \new_[41396]_ ;
  assign \new_[41401]_  = ~A202 & A201;
  assign \new_[41402]_  = ~A166 & \new_[41401]_ ;
  assign \new_[41403]_  = \new_[41402]_  & \new_[41397]_ ;
  assign \new_[41407]_  = A266 & ~A265;
  assign \new_[41408]_  = A203 & \new_[41407]_ ;
  assign \new_[41411]_  = ~A269 & A267;
  assign \new_[41414]_  = A301 & ~A300;
  assign \new_[41415]_  = \new_[41414]_  & \new_[41411]_ ;
  assign \new_[41416]_  = \new_[41415]_  & \new_[41408]_ ;
  assign \new_[41420]_  = A167 & A168;
  assign \new_[41421]_  = A170 & \new_[41420]_ ;
  assign \new_[41425]_  = ~A202 & A201;
  assign \new_[41426]_  = ~A166 & \new_[41425]_ ;
  assign \new_[41427]_  = \new_[41426]_  & \new_[41421]_ ;
  assign \new_[41431]_  = A266 & ~A265;
  assign \new_[41432]_  = A203 & \new_[41431]_ ;
  assign \new_[41435]_  = ~A269 & A267;
  assign \new_[41438]_  = ~A302 & ~A300;
  assign \new_[41439]_  = \new_[41438]_  & \new_[41435]_ ;
  assign \new_[41440]_  = \new_[41439]_  & \new_[41432]_ ;
  assign \new_[41444]_  = A167 & A168;
  assign \new_[41445]_  = A170 & \new_[41444]_ ;
  assign \new_[41449]_  = ~A202 & A201;
  assign \new_[41450]_  = ~A166 & \new_[41449]_ ;
  assign \new_[41451]_  = \new_[41450]_  & \new_[41445]_ ;
  assign \new_[41455]_  = A266 & ~A265;
  assign \new_[41456]_  = A203 & \new_[41455]_ ;
  assign \new_[41459]_  = ~A269 & A267;
  assign \new_[41462]_  = A299 & A298;
  assign \new_[41463]_  = \new_[41462]_  & \new_[41459]_ ;
  assign \new_[41464]_  = \new_[41463]_  & \new_[41456]_ ;
  assign \new_[41468]_  = A167 & A168;
  assign \new_[41469]_  = A170 & \new_[41468]_ ;
  assign \new_[41473]_  = ~A202 & A201;
  assign \new_[41474]_  = ~A166 & \new_[41473]_ ;
  assign \new_[41475]_  = \new_[41474]_  & \new_[41469]_ ;
  assign \new_[41479]_  = A266 & ~A265;
  assign \new_[41480]_  = A203 & \new_[41479]_ ;
  assign \new_[41483]_  = ~A269 & A267;
  assign \new_[41486]_  = ~A299 & ~A298;
  assign \new_[41487]_  = \new_[41486]_  & \new_[41483]_ ;
  assign \new_[41488]_  = \new_[41487]_  & \new_[41480]_ ;
  assign \new_[41492]_  = A167 & A168;
  assign \new_[41493]_  = A170 & \new_[41492]_ ;
  assign \new_[41497]_  = ~A202 & A201;
  assign \new_[41498]_  = ~A166 & \new_[41497]_ ;
  assign \new_[41499]_  = \new_[41498]_  & \new_[41493]_ ;
  assign \new_[41503]_  = ~A266 & A265;
  assign \new_[41504]_  = A203 & \new_[41503]_ ;
  assign \new_[41507]_  = A268 & A267;
  assign \new_[41510]_  = A301 & ~A300;
  assign \new_[41511]_  = \new_[41510]_  & \new_[41507]_ ;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41504]_ ;
  assign \new_[41516]_  = A167 & A168;
  assign \new_[41517]_  = A170 & \new_[41516]_ ;
  assign \new_[41521]_  = ~A202 & A201;
  assign \new_[41522]_  = ~A166 & \new_[41521]_ ;
  assign \new_[41523]_  = \new_[41522]_  & \new_[41517]_ ;
  assign \new_[41527]_  = ~A266 & A265;
  assign \new_[41528]_  = A203 & \new_[41527]_ ;
  assign \new_[41531]_  = A268 & A267;
  assign \new_[41534]_  = ~A302 & ~A300;
  assign \new_[41535]_  = \new_[41534]_  & \new_[41531]_ ;
  assign \new_[41536]_  = \new_[41535]_  & \new_[41528]_ ;
  assign \new_[41540]_  = A167 & A168;
  assign \new_[41541]_  = A170 & \new_[41540]_ ;
  assign \new_[41545]_  = ~A202 & A201;
  assign \new_[41546]_  = ~A166 & \new_[41545]_ ;
  assign \new_[41547]_  = \new_[41546]_  & \new_[41541]_ ;
  assign \new_[41551]_  = ~A266 & A265;
  assign \new_[41552]_  = A203 & \new_[41551]_ ;
  assign \new_[41555]_  = A268 & A267;
  assign \new_[41558]_  = A299 & A298;
  assign \new_[41559]_  = \new_[41558]_  & \new_[41555]_ ;
  assign \new_[41560]_  = \new_[41559]_  & \new_[41552]_ ;
  assign \new_[41564]_  = A167 & A168;
  assign \new_[41565]_  = A170 & \new_[41564]_ ;
  assign \new_[41569]_  = ~A202 & A201;
  assign \new_[41570]_  = ~A166 & \new_[41569]_ ;
  assign \new_[41571]_  = \new_[41570]_  & \new_[41565]_ ;
  assign \new_[41575]_  = ~A266 & A265;
  assign \new_[41576]_  = A203 & \new_[41575]_ ;
  assign \new_[41579]_  = A268 & A267;
  assign \new_[41582]_  = ~A299 & ~A298;
  assign \new_[41583]_  = \new_[41582]_  & \new_[41579]_ ;
  assign \new_[41584]_  = \new_[41583]_  & \new_[41576]_ ;
  assign \new_[41588]_  = A167 & A168;
  assign \new_[41589]_  = A170 & \new_[41588]_ ;
  assign \new_[41593]_  = ~A202 & A201;
  assign \new_[41594]_  = ~A166 & \new_[41593]_ ;
  assign \new_[41595]_  = \new_[41594]_  & \new_[41589]_ ;
  assign \new_[41599]_  = ~A266 & A265;
  assign \new_[41600]_  = A203 & \new_[41599]_ ;
  assign \new_[41603]_  = ~A269 & A267;
  assign \new_[41606]_  = A301 & ~A300;
  assign \new_[41607]_  = \new_[41606]_  & \new_[41603]_ ;
  assign \new_[41608]_  = \new_[41607]_  & \new_[41600]_ ;
  assign \new_[41612]_  = A167 & A168;
  assign \new_[41613]_  = A170 & \new_[41612]_ ;
  assign \new_[41617]_  = ~A202 & A201;
  assign \new_[41618]_  = ~A166 & \new_[41617]_ ;
  assign \new_[41619]_  = \new_[41618]_  & \new_[41613]_ ;
  assign \new_[41623]_  = ~A266 & A265;
  assign \new_[41624]_  = A203 & \new_[41623]_ ;
  assign \new_[41627]_  = ~A269 & A267;
  assign \new_[41630]_  = ~A302 & ~A300;
  assign \new_[41631]_  = \new_[41630]_  & \new_[41627]_ ;
  assign \new_[41632]_  = \new_[41631]_  & \new_[41624]_ ;
  assign \new_[41636]_  = A167 & A168;
  assign \new_[41637]_  = A170 & \new_[41636]_ ;
  assign \new_[41641]_  = ~A202 & A201;
  assign \new_[41642]_  = ~A166 & \new_[41641]_ ;
  assign \new_[41643]_  = \new_[41642]_  & \new_[41637]_ ;
  assign \new_[41647]_  = ~A266 & A265;
  assign \new_[41648]_  = A203 & \new_[41647]_ ;
  assign \new_[41651]_  = ~A269 & A267;
  assign \new_[41654]_  = A299 & A298;
  assign \new_[41655]_  = \new_[41654]_  & \new_[41651]_ ;
  assign \new_[41656]_  = \new_[41655]_  & \new_[41648]_ ;
  assign \new_[41660]_  = A167 & A168;
  assign \new_[41661]_  = A170 & \new_[41660]_ ;
  assign \new_[41665]_  = ~A202 & A201;
  assign \new_[41666]_  = ~A166 & \new_[41665]_ ;
  assign \new_[41667]_  = \new_[41666]_  & \new_[41661]_ ;
  assign \new_[41671]_  = ~A266 & A265;
  assign \new_[41672]_  = A203 & \new_[41671]_ ;
  assign \new_[41675]_  = ~A269 & A267;
  assign \new_[41678]_  = ~A299 & ~A298;
  assign \new_[41679]_  = \new_[41678]_  & \new_[41675]_ ;
  assign \new_[41680]_  = \new_[41679]_  & \new_[41672]_ ;
  assign \new_[41684]_  = A167 & A168;
  assign \new_[41685]_  = A170 & \new_[41684]_ ;
  assign \new_[41689]_  = ~A202 & A201;
  assign \new_[41690]_  = ~A166 & \new_[41689]_ ;
  assign \new_[41691]_  = \new_[41690]_  & \new_[41685]_ ;
  assign \new_[41695]_  = ~A266 & ~A265;
  assign \new_[41696]_  = A203 & \new_[41695]_ ;
  assign \new_[41699]_  = ~A299 & A298;
  assign \new_[41702]_  = A301 & A300;
  assign \new_[41703]_  = \new_[41702]_  & \new_[41699]_ ;
  assign \new_[41704]_  = \new_[41703]_  & \new_[41696]_ ;
  assign \new_[41708]_  = A167 & A168;
  assign \new_[41709]_  = A170 & \new_[41708]_ ;
  assign \new_[41713]_  = ~A202 & A201;
  assign \new_[41714]_  = ~A166 & \new_[41713]_ ;
  assign \new_[41715]_  = \new_[41714]_  & \new_[41709]_ ;
  assign \new_[41719]_  = ~A266 & ~A265;
  assign \new_[41720]_  = A203 & \new_[41719]_ ;
  assign \new_[41723]_  = ~A299 & A298;
  assign \new_[41726]_  = ~A302 & A300;
  assign \new_[41727]_  = \new_[41726]_  & \new_[41723]_ ;
  assign \new_[41728]_  = \new_[41727]_  & \new_[41720]_ ;
  assign \new_[41732]_  = A167 & A168;
  assign \new_[41733]_  = A170 & \new_[41732]_ ;
  assign \new_[41737]_  = ~A202 & A201;
  assign \new_[41738]_  = ~A166 & \new_[41737]_ ;
  assign \new_[41739]_  = \new_[41738]_  & \new_[41733]_ ;
  assign \new_[41743]_  = ~A266 & ~A265;
  assign \new_[41744]_  = A203 & \new_[41743]_ ;
  assign \new_[41747]_  = A299 & ~A298;
  assign \new_[41750]_  = A301 & A300;
  assign \new_[41751]_  = \new_[41750]_  & \new_[41747]_ ;
  assign \new_[41752]_  = \new_[41751]_  & \new_[41744]_ ;
  assign \new_[41756]_  = A167 & A168;
  assign \new_[41757]_  = A170 & \new_[41756]_ ;
  assign \new_[41761]_  = ~A202 & A201;
  assign \new_[41762]_  = ~A166 & \new_[41761]_ ;
  assign \new_[41763]_  = \new_[41762]_  & \new_[41757]_ ;
  assign \new_[41767]_  = ~A266 & ~A265;
  assign \new_[41768]_  = A203 & \new_[41767]_ ;
  assign \new_[41771]_  = A299 & ~A298;
  assign \new_[41774]_  = ~A302 & A300;
  assign \new_[41775]_  = \new_[41774]_  & \new_[41771]_ ;
  assign \new_[41776]_  = \new_[41775]_  & \new_[41768]_ ;
  assign \new_[41780]_  = A167 & A168;
  assign \new_[41781]_  = A170 & \new_[41780]_ ;
  assign \new_[41785]_  = A202 & ~A201;
  assign \new_[41786]_  = ~A166 & \new_[41785]_ ;
  assign \new_[41787]_  = \new_[41786]_  & \new_[41781]_ ;
  assign \new_[41791]_  = A269 & ~A268;
  assign \new_[41792]_  = A267 & \new_[41791]_ ;
  assign \new_[41795]_  = ~A299 & A298;
  assign \new_[41798]_  = A301 & A300;
  assign \new_[41799]_  = \new_[41798]_  & \new_[41795]_ ;
  assign \new_[41800]_  = \new_[41799]_  & \new_[41792]_ ;
  assign \new_[41804]_  = A167 & A168;
  assign \new_[41805]_  = A170 & \new_[41804]_ ;
  assign \new_[41809]_  = A202 & ~A201;
  assign \new_[41810]_  = ~A166 & \new_[41809]_ ;
  assign \new_[41811]_  = \new_[41810]_  & \new_[41805]_ ;
  assign \new_[41815]_  = A269 & ~A268;
  assign \new_[41816]_  = A267 & \new_[41815]_ ;
  assign \new_[41819]_  = ~A299 & A298;
  assign \new_[41822]_  = ~A302 & A300;
  assign \new_[41823]_  = \new_[41822]_  & \new_[41819]_ ;
  assign \new_[41824]_  = \new_[41823]_  & \new_[41816]_ ;
  assign \new_[41828]_  = A167 & A168;
  assign \new_[41829]_  = A170 & \new_[41828]_ ;
  assign \new_[41833]_  = A202 & ~A201;
  assign \new_[41834]_  = ~A166 & \new_[41833]_ ;
  assign \new_[41835]_  = \new_[41834]_  & \new_[41829]_ ;
  assign \new_[41839]_  = A269 & ~A268;
  assign \new_[41840]_  = A267 & \new_[41839]_ ;
  assign \new_[41843]_  = A299 & ~A298;
  assign \new_[41846]_  = A301 & A300;
  assign \new_[41847]_  = \new_[41846]_  & \new_[41843]_ ;
  assign \new_[41848]_  = \new_[41847]_  & \new_[41840]_ ;
  assign \new_[41852]_  = A167 & A168;
  assign \new_[41853]_  = A170 & \new_[41852]_ ;
  assign \new_[41857]_  = A202 & ~A201;
  assign \new_[41858]_  = ~A166 & \new_[41857]_ ;
  assign \new_[41859]_  = \new_[41858]_  & \new_[41853]_ ;
  assign \new_[41863]_  = A269 & ~A268;
  assign \new_[41864]_  = A267 & \new_[41863]_ ;
  assign \new_[41867]_  = A299 & ~A298;
  assign \new_[41870]_  = ~A302 & A300;
  assign \new_[41871]_  = \new_[41870]_  & \new_[41867]_ ;
  assign \new_[41872]_  = \new_[41871]_  & \new_[41864]_ ;
  assign \new_[41876]_  = A167 & A168;
  assign \new_[41877]_  = A170 & \new_[41876]_ ;
  assign \new_[41881]_  = A202 & ~A201;
  assign \new_[41882]_  = ~A166 & \new_[41881]_ ;
  assign \new_[41883]_  = \new_[41882]_  & \new_[41877]_ ;
  assign \new_[41887]_  = A298 & A268;
  assign \new_[41888]_  = ~A267 & \new_[41887]_ ;
  assign \new_[41891]_  = ~A300 & ~A299;
  assign \new_[41894]_  = A302 & ~A301;
  assign \new_[41895]_  = \new_[41894]_  & \new_[41891]_ ;
  assign \new_[41896]_  = \new_[41895]_  & \new_[41888]_ ;
  assign \new_[41900]_  = A167 & A168;
  assign \new_[41901]_  = A170 & \new_[41900]_ ;
  assign \new_[41905]_  = A202 & ~A201;
  assign \new_[41906]_  = ~A166 & \new_[41905]_ ;
  assign \new_[41907]_  = \new_[41906]_  & \new_[41901]_ ;
  assign \new_[41911]_  = ~A298 & A268;
  assign \new_[41912]_  = ~A267 & \new_[41911]_ ;
  assign \new_[41915]_  = ~A300 & A299;
  assign \new_[41918]_  = A302 & ~A301;
  assign \new_[41919]_  = \new_[41918]_  & \new_[41915]_ ;
  assign \new_[41920]_  = \new_[41919]_  & \new_[41912]_ ;
  assign \new_[41924]_  = A167 & A168;
  assign \new_[41925]_  = A170 & \new_[41924]_ ;
  assign \new_[41929]_  = A202 & ~A201;
  assign \new_[41930]_  = ~A166 & \new_[41929]_ ;
  assign \new_[41931]_  = \new_[41930]_  & \new_[41925]_ ;
  assign \new_[41935]_  = A298 & ~A269;
  assign \new_[41936]_  = ~A267 & \new_[41935]_ ;
  assign \new_[41939]_  = ~A300 & ~A299;
  assign \new_[41942]_  = A302 & ~A301;
  assign \new_[41943]_  = \new_[41942]_  & \new_[41939]_ ;
  assign \new_[41944]_  = \new_[41943]_  & \new_[41936]_ ;
  assign \new_[41948]_  = A167 & A168;
  assign \new_[41949]_  = A170 & \new_[41948]_ ;
  assign \new_[41953]_  = A202 & ~A201;
  assign \new_[41954]_  = ~A166 & \new_[41953]_ ;
  assign \new_[41955]_  = \new_[41954]_  & \new_[41949]_ ;
  assign \new_[41959]_  = ~A298 & ~A269;
  assign \new_[41960]_  = ~A267 & \new_[41959]_ ;
  assign \new_[41963]_  = ~A300 & A299;
  assign \new_[41966]_  = A302 & ~A301;
  assign \new_[41967]_  = \new_[41966]_  & \new_[41963]_ ;
  assign \new_[41968]_  = \new_[41967]_  & \new_[41960]_ ;
  assign \new_[41972]_  = A167 & A168;
  assign \new_[41973]_  = A170 & \new_[41972]_ ;
  assign \new_[41977]_  = A202 & ~A201;
  assign \new_[41978]_  = ~A166 & \new_[41977]_ ;
  assign \new_[41979]_  = \new_[41978]_  & \new_[41973]_ ;
  assign \new_[41983]_  = A298 & A266;
  assign \new_[41984]_  = A265 & \new_[41983]_ ;
  assign \new_[41987]_  = ~A300 & ~A299;
  assign \new_[41990]_  = A302 & ~A301;
  assign \new_[41991]_  = \new_[41990]_  & \new_[41987]_ ;
  assign \new_[41992]_  = \new_[41991]_  & \new_[41984]_ ;
  assign \new_[41996]_  = A167 & A168;
  assign \new_[41997]_  = A170 & \new_[41996]_ ;
  assign \new_[42001]_  = A202 & ~A201;
  assign \new_[42002]_  = ~A166 & \new_[42001]_ ;
  assign \new_[42003]_  = \new_[42002]_  & \new_[41997]_ ;
  assign \new_[42007]_  = ~A298 & A266;
  assign \new_[42008]_  = A265 & \new_[42007]_ ;
  assign \new_[42011]_  = ~A300 & A299;
  assign \new_[42014]_  = A302 & ~A301;
  assign \new_[42015]_  = \new_[42014]_  & \new_[42011]_ ;
  assign \new_[42016]_  = \new_[42015]_  & \new_[42008]_ ;
  assign \new_[42020]_  = A167 & A168;
  assign \new_[42021]_  = A170 & \new_[42020]_ ;
  assign \new_[42025]_  = A202 & ~A201;
  assign \new_[42026]_  = ~A166 & \new_[42025]_ ;
  assign \new_[42027]_  = \new_[42026]_  & \new_[42021]_ ;
  assign \new_[42031]_  = A267 & A266;
  assign \new_[42032]_  = ~A265 & \new_[42031]_ ;
  assign \new_[42035]_  = A300 & A268;
  assign \new_[42038]_  = A302 & ~A301;
  assign \new_[42039]_  = \new_[42038]_  & \new_[42035]_ ;
  assign \new_[42040]_  = \new_[42039]_  & \new_[42032]_ ;
  assign \new_[42044]_  = A167 & A168;
  assign \new_[42045]_  = A170 & \new_[42044]_ ;
  assign \new_[42049]_  = A202 & ~A201;
  assign \new_[42050]_  = ~A166 & \new_[42049]_ ;
  assign \new_[42051]_  = \new_[42050]_  & \new_[42045]_ ;
  assign \new_[42055]_  = A267 & A266;
  assign \new_[42056]_  = ~A265 & \new_[42055]_ ;
  assign \new_[42059]_  = A300 & ~A269;
  assign \new_[42062]_  = A302 & ~A301;
  assign \new_[42063]_  = \new_[42062]_  & \new_[42059]_ ;
  assign \new_[42064]_  = \new_[42063]_  & \new_[42056]_ ;
  assign \new_[42068]_  = A167 & A168;
  assign \new_[42069]_  = A170 & \new_[42068]_ ;
  assign \new_[42073]_  = A202 & ~A201;
  assign \new_[42074]_  = ~A166 & \new_[42073]_ ;
  assign \new_[42075]_  = \new_[42074]_  & \new_[42069]_ ;
  assign \new_[42079]_  = ~A267 & A266;
  assign \new_[42080]_  = ~A265 & \new_[42079]_ ;
  assign \new_[42083]_  = A269 & ~A268;
  assign \new_[42086]_  = A301 & ~A300;
  assign \new_[42087]_  = \new_[42086]_  & \new_[42083]_ ;
  assign \new_[42088]_  = \new_[42087]_  & \new_[42080]_ ;
  assign \new_[42092]_  = A167 & A168;
  assign \new_[42093]_  = A170 & \new_[42092]_ ;
  assign \new_[42097]_  = A202 & ~A201;
  assign \new_[42098]_  = ~A166 & \new_[42097]_ ;
  assign \new_[42099]_  = \new_[42098]_  & \new_[42093]_ ;
  assign \new_[42103]_  = ~A267 & A266;
  assign \new_[42104]_  = ~A265 & \new_[42103]_ ;
  assign \new_[42107]_  = A269 & ~A268;
  assign \new_[42110]_  = ~A302 & ~A300;
  assign \new_[42111]_  = \new_[42110]_  & \new_[42107]_ ;
  assign \new_[42112]_  = \new_[42111]_  & \new_[42104]_ ;
  assign \new_[42116]_  = A167 & A168;
  assign \new_[42117]_  = A170 & \new_[42116]_ ;
  assign \new_[42121]_  = A202 & ~A201;
  assign \new_[42122]_  = ~A166 & \new_[42121]_ ;
  assign \new_[42123]_  = \new_[42122]_  & \new_[42117]_ ;
  assign \new_[42127]_  = ~A267 & A266;
  assign \new_[42128]_  = ~A265 & \new_[42127]_ ;
  assign \new_[42131]_  = A269 & ~A268;
  assign \new_[42134]_  = A299 & A298;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42136]_  = \new_[42135]_  & \new_[42128]_ ;
  assign \new_[42140]_  = A167 & A168;
  assign \new_[42141]_  = A170 & \new_[42140]_ ;
  assign \new_[42145]_  = A202 & ~A201;
  assign \new_[42146]_  = ~A166 & \new_[42145]_ ;
  assign \new_[42147]_  = \new_[42146]_  & \new_[42141]_ ;
  assign \new_[42151]_  = ~A267 & A266;
  assign \new_[42152]_  = ~A265 & \new_[42151]_ ;
  assign \new_[42155]_  = A269 & ~A268;
  assign \new_[42158]_  = ~A299 & ~A298;
  assign \new_[42159]_  = \new_[42158]_  & \new_[42155]_ ;
  assign \new_[42160]_  = \new_[42159]_  & \new_[42152]_ ;
  assign \new_[42164]_  = A167 & A168;
  assign \new_[42165]_  = A170 & \new_[42164]_ ;
  assign \new_[42169]_  = A202 & ~A201;
  assign \new_[42170]_  = ~A166 & \new_[42169]_ ;
  assign \new_[42171]_  = \new_[42170]_  & \new_[42165]_ ;
  assign \new_[42175]_  = A267 & ~A266;
  assign \new_[42176]_  = A265 & \new_[42175]_ ;
  assign \new_[42179]_  = A300 & A268;
  assign \new_[42182]_  = A302 & ~A301;
  assign \new_[42183]_  = \new_[42182]_  & \new_[42179]_ ;
  assign \new_[42184]_  = \new_[42183]_  & \new_[42176]_ ;
  assign \new_[42188]_  = A167 & A168;
  assign \new_[42189]_  = A170 & \new_[42188]_ ;
  assign \new_[42193]_  = A202 & ~A201;
  assign \new_[42194]_  = ~A166 & \new_[42193]_ ;
  assign \new_[42195]_  = \new_[42194]_  & \new_[42189]_ ;
  assign \new_[42199]_  = A267 & ~A266;
  assign \new_[42200]_  = A265 & \new_[42199]_ ;
  assign \new_[42203]_  = A300 & ~A269;
  assign \new_[42206]_  = A302 & ~A301;
  assign \new_[42207]_  = \new_[42206]_  & \new_[42203]_ ;
  assign \new_[42208]_  = \new_[42207]_  & \new_[42200]_ ;
  assign \new_[42212]_  = A167 & A168;
  assign \new_[42213]_  = A170 & \new_[42212]_ ;
  assign \new_[42217]_  = A202 & ~A201;
  assign \new_[42218]_  = ~A166 & \new_[42217]_ ;
  assign \new_[42219]_  = \new_[42218]_  & \new_[42213]_ ;
  assign \new_[42223]_  = ~A267 & ~A266;
  assign \new_[42224]_  = A265 & \new_[42223]_ ;
  assign \new_[42227]_  = A269 & ~A268;
  assign \new_[42230]_  = A301 & ~A300;
  assign \new_[42231]_  = \new_[42230]_  & \new_[42227]_ ;
  assign \new_[42232]_  = \new_[42231]_  & \new_[42224]_ ;
  assign \new_[42236]_  = A167 & A168;
  assign \new_[42237]_  = A170 & \new_[42236]_ ;
  assign \new_[42241]_  = A202 & ~A201;
  assign \new_[42242]_  = ~A166 & \new_[42241]_ ;
  assign \new_[42243]_  = \new_[42242]_  & \new_[42237]_ ;
  assign \new_[42247]_  = ~A267 & ~A266;
  assign \new_[42248]_  = A265 & \new_[42247]_ ;
  assign \new_[42251]_  = A269 & ~A268;
  assign \new_[42254]_  = ~A302 & ~A300;
  assign \new_[42255]_  = \new_[42254]_  & \new_[42251]_ ;
  assign \new_[42256]_  = \new_[42255]_  & \new_[42248]_ ;
  assign \new_[42260]_  = A167 & A168;
  assign \new_[42261]_  = A170 & \new_[42260]_ ;
  assign \new_[42265]_  = A202 & ~A201;
  assign \new_[42266]_  = ~A166 & \new_[42265]_ ;
  assign \new_[42267]_  = \new_[42266]_  & \new_[42261]_ ;
  assign \new_[42271]_  = ~A267 & ~A266;
  assign \new_[42272]_  = A265 & \new_[42271]_ ;
  assign \new_[42275]_  = A269 & ~A268;
  assign \new_[42278]_  = A299 & A298;
  assign \new_[42279]_  = \new_[42278]_  & \new_[42275]_ ;
  assign \new_[42280]_  = \new_[42279]_  & \new_[42272]_ ;
  assign \new_[42284]_  = A167 & A168;
  assign \new_[42285]_  = A170 & \new_[42284]_ ;
  assign \new_[42289]_  = A202 & ~A201;
  assign \new_[42290]_  = ~A166 & \new_[42289]_ ;
  assign \new_[42291]_  = \new_[42290]_  & \new_[42285]_ ;
  assign \new_[42295]_  = ~A267 & ~A266;
  assign \new_[42296]_  = A265 & \new_[42295]_ ;
  assign \new_[42299]_  = A269 & ~A268;
  assign \new_[42302]_  = ~A299 & ~A298;
  assign \new_[42303]_  = \new_[42302]_  & \new_[42299]_ ;
  assign \new_[42304]_  = \new_[42303]_  & \new_[42296]_ ;
  assign \new_[42308]_  = A167 & A168;
  assign \new_[42309]_  = A170 & \new_[42308]_ ;
  assign \new_[42313]_  = A202 & ~A201;
  assign \new_[42314]_  = ~A166 & \new_[42313]_ ;
  assign \new_[42315]_  = \new_[42314]_  & \new_[42309]_ ;
  assign \new_[42319]_  = A298 & ~A266;
  assign \new_[42320]_  = ~A265 & \new_[42319]_ ;
  assign \new_[42323]_  = ~A300 & ~A299;
  assign \new_[42326]_  = A302 & ~A301;
  assign \new_[42327]_  = \new_[42326]_  & \new_[42323]_ ;
  assign \new_[42328]_  = \new_[42327]_  & \new_[42320]_ ;
  assign \new_[42332]_  = A167 & A168;
  assign \new_[42333]_  = A170 & \new_[42332]_ ;
  assign \new_[42337]_  = A202 & ~A201;
  assign \new_[42338]_  = ~A166 & \new_[42337]_ ;
  assign \new_[42339]_  = \new_[42338]_  & \new_[42333]_ ;
  assign \new_[42343]_  = ~A298 & ~A266;
  assign \new_[42344]_  = ~A265 & \new_[42343]_ ;
  assign \new_[42347]_  = ~A300 & A299;
  assign \new_[42350]_  = A302 & ~A301;
  assign \new_[42351]_  = \new_[42350]_  & \new_[42347]_ ;
  assign \new_[42352]_  = \new_[42351]_  & \new_[42344]_ ;
  assign \new_[42356]_  = A167 & A168;
  assign \new_[42357]_  = A170 & \new_[42356]_ ;
  assign \new_[42361]_  = ~A203 & ~A201;
  assign \new_[42362]_  = ~A166 & \new_[42361]_ ;
  assign \new_[42363]_  = \new_[42362]_  & \new_[42357]_ ;
  assign \new_[42367]_  = A269 & ~A268;
  assign \new_[42368]_  = A267 & \new_[42367]_ ;
  assign \new_[42371]_  = ~A299 & A298;
  assign \new_[42374]_  = A301 & A300;
  assign \new_[42375]_  = \new_[42374]_  & \new_[42371]_ ;
  assign \new_[42376]_  = \new_[42375]_  & \new_[42368]_ ;
  assign \new_[42380]_  = A167 & A168;
  assign \new_[42381]_  = A170 & \new_[42380]_ ;
  assign \new_[42385]_  = ~A203 & ~A201;
  assign \new_[42386]_  = ~A166 & \new_[42385]_ ;
  assign \new_[42387]_  = \new_[42386]_  & \new_[42381]_ ;
  assign \new_[42391]_  = A269 & ~A268;
  assign \new_[42392]_  = A267 & \new_[42391]_ ;
  assign \new_[42395]_  = ~A299 & A298;
  assign \new_[42398]_  = ~A302 & A300;
  assign \new_[42399]_  = \new_[42398]_  & \new_[42395]_ ;
  assign \new_[42400]_  = \new_[42399]_  & \new_[42392]_ ;
  assign \new_[42404]_  = A167 & A168;
  assign \new_[42405]_  = A170 & \new_[42404]_ ;
  assign \new_[42409]_  = ~A203 & ~A201;
  assign \new_[42410]_  = ~A166 & \new_[42409]_ ;
  assign \new_[42411]_  = \new_[42410]_  & \new_[42405]_ ;
  assign \new_[42415]_  = A269 & ~A268;
  assign \new_[42416]_  = A267 & \new_[42415]_ ;
  assign \new_[42419]_  = A299 & ~A298;
  assign \new_[42422]_  = A301 & A300;
  assign \new_[42423]_  = \new_[42422]_  & \new_[42419]_ ;
  assign \new_[42424]_  = \new_[42423]_  & \new_[42416]_ ;
  assign \new_[42428]_  = A167 & A168;
  assign \new_[42429]_  = A170 & \new_[42428]_ ;
  assign \new_[42433]_  = ~A203 & ~A201;
  assign \new_[42434]_  = ~A166 & \new_[42433]_ ;
  assign \new_[42435]_  = \new_[42434]_  & \new_[42429]_ ;
  assign \new_[42439]_  = A269 & ~A268;
  assign \new_[42440]_  = A267 & \new_[42439]_ ;
  assign \new_[42443]_  = A299 & ~A298;
  assign \new_[42446]_  = ~A302 & A300;
  assign \new_[42447]_  = \new_[42446]_  & \new_[42443]_ ;
  assign \new_[42448]_  = \new_[42447]_  & \new_[42440]_ ;
  assign \new_[42452]_  = A167 & A168;
  assign \new_[42453]_  = A170 & \new_[42452]_ ;
  assign \new_[42457]_  = ~A203 & ~A201;
  assign \new_[42458]_  = ~A166 & \new_[42457]_ ;
  assign \new_[42459]_  = \new_[42458]_  & \new_[42453]_ ;
  assign \new_[42463]_  = A298 & A268;
  assign \new_[42464]_  = ~A267 & \new_[42463]_ ;
  assign \new_[42467]_  = ~A300 & ~A299;
  assign \new_[42470]_  = A302 & ~A301;
  assign \new_[42471]_  = \new_[42470]_  & \new_[42467]_ ;
  assign \new_[42472]_  = \new_[42471]_  & \new_[42464]_ ;
  assign \new_[42476]_  = A167 & A168;
  assign \new_[42477]_  = A170 & \new_[42476]_ ;
  assign \new_[42481]_  = ~A203 & ~A201;
  assign \new_[42482]_  = ~A166 & \new_[42481]_ ;
  assign \new_[42483]_  = \new_[42482]_  & \new_[42477]_ ;
  assign \new_[42487]_  = ~A298 & A268;
  assign \new_[42488]_  = ~A267 & \new_[42487]_ ;
  assign \new_[42491]_  = ~A300 & A299;
  assign \new_[42494]_  = A302 & ~A301;
  assign \new_[42495]_  = \new_[42494]_  & \new_[42491]_ ;
  assign \new_[42496]_  = \new_[42495]_  & \new_[42488]_ ;
  assign \new_[42500]_  = A167 & A168;
  assign \new_[42501]_  = A170 & \new_[42500]_ ;
  assign \new_[42505]_  = ~A203 & ~A201;
  assign \new_[42506]_  = ~A166 & \new_[42505]_ ;
  assign \new_[42507]_  = \new_[42506]_  & \new_[42501]_ ;
  assign \new_[42511]_  = A298 & ~A269;
  assign \new_[42512]_  = ~A267 & \new_[42511]_ ;
  assign \new_[42515]_  = ~A300 & ~A299;
  assign \new_[42518]_  = A302 & ~A301;
  assign \new_[42519]_  = \new_[42518]_  & \new_[42515]_ ;
  assign \new_[42520]_  = \new_[42519]_  & \new_[42512]_ ;
  assign \new_[42524]_  = A167 & A168;
  assign \new_[42525]_  = A170 & \new_[42524]_ ;
  assign \new_[42529]_  = ~A203 & ~A201;
  assign \new_[42530]_  = ~A166 & \new_[42529]_ ;
  assign \new_[42531]_  = \new_[42530]_  & \new_[42525]_ ;
  assign \new_[42535]_  = ~A298 & ~A269;
  assign \new_[42536]_  = ~A267 & \new_[42535]_ ;
  assign \new_[42539]_  = ~A300 & A299;
  assign \new_[42542]_  = A302 & ~A301;
  assign \new_[42543]_  = \new_[42542]_  & \new_[42539]_ ;
  assign \new_[42544]_  = \new_[42543]_  & \new_[42536]_ ;
  assign \new_[42548]_  = A167 & A168;
  assign \new_[42549]_  = A170 & \new_[42548]_ ;
  assign \new_[42553]_  = ~A203 & ~A201;
  assign \new_[42554]_  = ~A166 & \new_[42553]_ ;
  assign \new_[42555]_  = \new_[42554]_  & \new_[42549]_ ;
  assign \new_[42559]_  = A298 & A266;
  assign \new_[42560]_  = A265 & \new_[42559]_ ;
  assign \new_[42563]_  = ~A300 & ~A299;
  assign \new_[42566]_  = A302 & ~A301;
  assign \new_[42567]_  = \new_[42566]_  & \new_[42563]_ ;
  assign \new_[42568]_  = \new_[42567]_  & \new_[42560]_ ;
  assign \new_[42572]_  = A167 & A168;
  assign \new_[42573]_  = A170 & \new_[42572]_ ;
  assign \new_[42577]_  = ~A203 & ~A201;
  assign \new_[42578]_  = ~A166 & \new_[42577]_ ;
  assign \new_[42579]_  = \new_[42578]_  & \new_[42573]_ ;
  assign \new_[42583]_  = ~A298 & A266;
  assign \new_[42584]_  = A265 & \new_[42583]_ ;
  assign \new_[42587]_  = ~A300 & A299;
  assign \new_[42590]_  = A302 & ~A301;
  assign \new_[42591]_  = \new_[42590]_  & \new_[42587]_ ;
  assign \new_[42592]_  = \new_[42591]_  & \new_[42584]_ ;
  assign \new_[42596]_  = A167 & A168;
  assign \new_[42597]_  = A170 & \new_[42596]_ ;
  assign \new_[42601]_  = ~A203 & ~A201;
  assign \new_[42602]_  = ~A166 & \new_[42601]_ ;
  assign \new_[42603]_  = \new_[42602]_  & \new_[42597]_ ;
  assign \new_[42607]_  = A267 & A266;
  assign \new_[42608]_  = ~A265 & \new_[42607]_ ;
  assign \new_[42611]_  = A300 & A268;
  assign \new_[42614]_  = A302 & ~A301;
  assign \new_[42615]_  = \new_[42614]_  & \new_[42611]_ ;
  assign \new_[42616]_  = \new_[42615]_  & \new_[42608]_ ;
  assign \new_[42620]_  = A167 & A168;
  assign \new_[42621]_  = A170 & \new_[42620]_ ;
  assign \new_[42625]_  = ~A203 & ~A201;
  assign \new_[42626]_  = ~A166 & \new_[42625]_ ;
  assign \new_[42627]_  = \new_[42626]_  & \new_[42621]_ ;
  assign \new_[42631]_  = A267 & A266;
  assign \new_[42632]_  = ~A265 & \new_[42631]_ ;
  assign \new_[42635]_  = A300 & ~A269;
  assign \new_[42638]_  = A302 & ~A301;
  assign \new_[42639]_  = \new_[42638]_  & \new_[42635]_ ;
  assign \new_[42640]_  = \new_[42639]_  & \new_[42632]_ ;
  assign \new_[42644]_  = A167 & A168;
  assign \new_[42645]_  = A170 & \new_[42644]_ ;
  assign \new_[42649]_  = ~A203 & ~A201;
  assign \new_[42650]_  = ~A166 & \new_[42649]_ ;
  assign \new_[42651]_  = \new_[42650]_  & \new_[42645]_ ;
  assign \new_[42655]_  = ~A267 & A266;
  assign \new_[42656]_  = ~A265 & \new_[42655]_ ;
  assign \new_[42659]_  = A269 & ~A268;
  assign \new_[42662]_  = A301 & ~A300;
  assign \new_[42663]_  = \new_[42662]_  & \new_[42659]_ ;
  assign \new_[42664]_  = \new_[42663]_  & \new_[42656]_ ;
  assign \new_[42668]_  = A167 & A168;
  assign \new_[42669]_  = A170 & \new_[42668]_ ;
  assign \new_[42673]_  = ~A203 & ~A201;
  assign \new_[42674]_  = ~A166 & \new_[42673]_ ;
  assign \new_[42675]_  = \new_[42674]_  & \new_[42669]_ ;
  assign \new_[42679]_  = ~A267 & A266;
  assign \new_[42680]_  = ~A265 & \new_[42679]_ ;
  assign \new_[42683]_  = A269 & ~A268;
  assign \new_[42686]_  = ~A302 & ~A300;
  assign \new_[42687]_  = \new_[42686]_  & \new_[42683]_ ;
  assign \new_[42688]_  = \new_[42687]_  & \new_[42680]_ ;
  assign \new_[42692]_  = A167 & A168;
  assign \new_[42693]_  = A170 & \new_[42692]_ ;
  assign \new_[42697]_  = ~A203 & ~A201;
  assign \new_[42698]_  = ~A166 & \new_[42697]_ ;
  assign \new_[42699]_  = \new_[42698]_  & \new_[42693]_ ;
  assign \new_[42703]_  = ~A267 & A266;
  assign \new_[42704]_  = ~A265 & \new_[42703]_ ;
  assign \new_[42707]_  = A269 & ~A268;
  assign \new_[42710]_  = A299 & A298;
  assign \new_[42711]_  = \new_[42710]_  & \new_[42707]_ ;
  assign \new_[42712]_  = \new_[42711]_  & \new_[42704]_ ;
  assign \new_[42716]_  = A167 & A168;
  assign \new_[42717]_  = A170 & \new_[42716]_ ;
  assign \new_[42721]_  = ~A203 & ~A201;
  assign \new_[42722]_  = ~A166 & \new_[42721]_ ;
  assign \new_[42723]_  = \new_[42722]_  & \new_[42717]_ ;
  assign \new_[42727]_  = ~A267 & A266;
  assign \new_[42728]_  = ~A265 & \new_[42727]_ ;
  assign \new_[42731]_  = A269 & ~A268;
  assign \new_[42734]_  = ~A299 & ~A298;
  assign \new_[42735]_  = \new_[42734]_  & \new_[42731]_ ;
  assign \new_[42736]_  = \new_[42735]_  & \new_[42728]_ ;
  assign \new_[42740]_  = A167 & A168;
  assign \new_[42741]_  = A170 & \new_[42740]_ ;
  assign \new_[42745]_  = ~A203 & ~A201;
  assign \new_[42746]_  = ~A166 & \new_[42745]_ ;
  assign \new_[42747]_  = \new_[42746]_  & \new_[42741]_ ;
  assign \new_[42751]_  = A267 & ~A266;
  assign \new_[42752]_  = A265 & \new_[42751]_ ;
  assign \new_[42755]_  = A300 & A268;
  assign \new_[42758]_  = A302 & ~A301;
  assign \new_[42759]_  = \new_[42758]_  & \new_[42755]_ ;
  assign \new_[42760]_  = \new_[42759]_  & \new_[42752]_ ;
  assign \new_[42764]_  = A167 & A168;
  assign \new_[42765]_  = A170 & \new_[42764]_ ;
  assign \new_[42769]_  = ~A203 & ~A201;
  assign \new_[42770]_  = ~A166 & \new_[42769]_ ;
  assign \new_[42771]_  = \new_[42770]_  & \new_[42765]_ ;
  assign \new_[42775]_  = A267 & ~A266;
  assign \new_[42776]_  = A265 & \new_[42775]_ ;
  assign \new_[42779]_  = A300 & ~A269;
  assign \new_[42782]_  = A302 & ~A301;
  assign \new_[42783]_  = \new_[42782]_  & \new_[42779]_ ;
  assign \new_[42784]_  = \new_[42783]_  & \new_[42776]_ ;
  assign \new_[42788]_  = A167 & A168;
  assign \new_[42789]_  = A170 & \new_[42788]_ ;
  assign \new_[42793]_  = ~A203 & ~A201;
  assign \new_[42794]_  = ~A166 & \new_[42793]_ ;
  assign \new_[42795]_  = \new_[42794]_  & \new_[42789]_ ;
  assign \new_[42799]_  = ~A267 & ~A266;
  assign \new_[42800]_  = A265 & \new_[42799]_ ;
  assign \new_[42803]_  = A269 & ~A268;
  assign \new_[42806]_  = A301 & ~A300;
  assign \new_[42807]_  = \new_[42806]_  & \new_[42803]_ ;
  assign \new_[42808]_  = \new_[42807]_  & \new_[42800]_ ;
  assign \new_[42812]_  = A167 & A168;
  assign \new_[42813]_  = A170 & \new_[42812]_ ;
  assign \new_[42817]_  = ~A203 & ~A201;
  assign \new_[42818]_  = ~A166 & \new_[42817]_ ;
  assign \new_[42819]_  = \new_[42818]_  & \new_[42813]_ ;
  assign \new_[42823]_  = ~A267 & ~A266;
  assign \new_[42824]_  = A265 & \new_[42823]_ ;
  assign \new_[42827]_  = A269 & ~A268;
  assign \new_[42830]_  = ~A302 & ~A300;
  assign \new_[42831]_  = \new_[42830]_  & \new_[42827]_ ;
  assign \new_[42832]_  = \new_[42831]_  & \new_[42824]_ ;
  assign \new_[42836]_  = A167 & A168;
  assign \new_[42837]_  = A170 & \new_[42836]_ ;
  assign \new_[42841]_  = ~A203 & ~A201;
  assign \new_[42842]_  = ~A166 & \new_[42841]_ ;
  assign \new_[42843]_  = \new_[42842]_  & \new_[42837]_ ;
  assign \new_[42847]_  = ~A267 & ~A266;
  assign \new_[42848]_  = A265 & \new_[42847]_ ;
  assign \new_[42851]_  = A269 & ~A268;
  assign \new_[42854]_  = A299 & A298;
  assign \new_[42855]_  = \new_[42854]_  & \new_[42851]_ ;
  assign \new_[42856]_  = \new_[42855]_  & \new_[42848]_ ;
  assign \new_[42860]_  = A167 & A168;
  assign \new_[42861]_  = A170 & \new_[42860]_ ;
  assign \new_[42865]_  = ~A203 & ~A201;
  assign \new_[42866]_  = ~A166 & \new_[42865]_ ;
  assign \new_[42867]_  = \new_[42866]_  & \new_[42861]_ ;
  assign \new_[42871]_  = ~A267 & ~A266;
  assign \new_[42872]_  = A265 & \new_[42871]_ ;
  assign \new_[42875]_  = A269 & ~A268;
  assign \new_[42878]_  = ~A299 & ~A298;
  assign \new_[42879]_  = \new_[42878]_  & \new_[42875]_ ;
  assign \new_[42880]_  = \new_[42879]_  & \new_[42872]_ ;
  assign \new_[42884]_  = A167 & A168;
  assign \new_[42885]_  = A170 & \new_[42884]_ ;
  assign \new_[42889]_  = ~A203 & ~A201;
  assign \new_[42890]_  = ~A166 & \new_[42889]_ ;
  assign \new_[42891]_  = \new_[42890]_  & \new_[42885]_ ;
  assign \new_[42895]_  = A298 & ~A266;
  assign \new_[42896]_  = ~A265 & \new_[42895]_ ;
  assign \new_[42899]_  = ~A300 & ~A299;
  assign \new_[42902]_  = A302 & ~A301;
  assign \new_[42903]_  = \new_[42902]_  & \new_[42899]_ ;
  assign \new_[42904]_  = \new_[42903]_  & \new_[42896]_ ;
  assign \new_[42908]_  = A167 & A168;
  assign \new_[42909]_  = A170 & \new_[42908]_ ;
  assign \new_[42913]_  = ~A203 & ~A201;
  assign \new_[42914]_  = ~A166 & \new_[42913]_ ;
  assign \new_[42915]_  = \new_[42914]_  & \new_[42909]_ ;
  assign \new_[42919]_  = ~A298 & ~A266;
  assign \new_[42920]_  = ~A265 & \new_[42919]_ ;
  assign \new_[42923]_  = ~A300 & A299;
  assign \new_[42926]_  = A302 & ~A301;
  assign \new_[42927]_  = \new_[42926]_  & \new_[42923]_ ;
  assign \new_[42928]_  = \new_[42927]_  & \new_[42920]_ ;
  assign \new_[42932]_  = A167 & A168;
  assign \new_[42933]_  = A170 & \new_[42932]_ ;
  assign \new_[42937]_  = A200 & A199;
  assign \new_[42938]_  = ~A166 & \new_[42937]_ ;
  assign \new_[42939]_  = \new_[42938]_  & \new_[42933]_ ;
  assign \new_[42943]_  = A269 & ~A268;
  assign \new_[42944]_  = A267 & \new_[42943]_ ;
  assign \new_[42947]_  = ~A299 & A298;
  assign \new_[42950]_  = A301 & A300;
  assign \new_[42951]_  = \new_[42950]_  & \new_[42947]_ ;
  assign \new_[42952]_  = \new_[42951]_  & \new_[42944]_ ;
  assign \new_[42956]_  = A167 & A168;
  assign \new_[42957]_  = A170 & \new_[42956]_ ;
  assign \new_[42961]_  = A200 & A199;
  assign \new_[42962]_  = ~A166 & \new_[42961]_ ;
  assign \new_[42963]_  = \new_[42962]_  & \new_[42957]_ ;
  assign \new_[42967]_  = A269 & ~A268;
  assign \new_[42968]_  = A267 & \new_[42967]_ ;
  assign \new_[42971]_  = ~A299 & A298;
  assign \new_[42974]_  = ~A302 & A300;
  assign \new_[42975]_  = \new_[42974]_  & \new_[42971]_ ;
  assign \new_[42976]_  = \new_[42975]_  & \new_[42968]_ ;
  assign \new_[42980]_  = A167 & A168;
  assign \new_[42981]_  = A170 & \new_[42980]_ ;
  assign \new_[42985]_  = A200 & A199;
  assign \new_[42986]_  = ~A166 & \new_[42985]_ ;
  assign \new_[42987]_  = \new_[42986]_  & \new_[42981]_ ;
  assign \new_[42991]_  = A269 & ~A268;
  assign \new_[42992]_  = A267 & \new_[42991]_ ;
  assign \new_[42995]_  = A299 & ~A298;
  assign \new_[42998]_  = A301 & A300;
  assign \new_[42999]_  = \new_[42998]_  & \new_[42995]_ ;
  assign \new_[43000]_  = \new_[42999]_  & \new_[42992]_ ;
  assign \new_[43004]_  = A167 & A168;
  assign \new_[43005]_  = A170 & \new_[43004]_ ;
  assign \new_[43009]_  = A200 & A199;
  assign \new_[43010]_  = ~A166 & \new_[43009]_ ;
  assign \new_[43011]_  = \new_[43010]_  & \new_[43005]_ ;
  assign \new_[43015]_  = A269 & ~A268;
  assign \new_[43016]_  = A267 & \new_[43015]_ ;
  assign \new_[43019]_  = A299 & ~A298;
  assign \new_[43022]_  = ~A302 & A300;
  assign \new_[43023]_  = \new_[43022]_  & \new_[43019]_ ;
  assign \new_[43024]_  = \new_[43023]_  & \new_[43016]_ ;
  assign \new_[43028]_  = A167 & A168;
  assign \new_[43029]_  = A170 & \new_[43028]_ ;
  assign \new_[43033]_  = A200 & A199;
  assign \new_[43034]_  = ~A166 & \new_[43033]_ ;
  assign \new_[43035]_  = \new_[43034]_  & \new_[43029]_ ;
  assign \new_[43039]_  = A298 & A268;
  assign \new_[43040]_  = ~A267 & \new_[43039]_ ;
  assign \new_[43043]_  = ~A300 & ~A299;
  assign \new_[43046]_  = A302 & ~A301;
  assign \new_[43047]_  = \new_[43046]_  & \new_[43043]_ ;
  assign \new_[43048]_  = \new_[43047]_  & \new_[43040]_ ;
  assign \new_[43052]_  = A167 & A168;
  assign \new_[43053]_  = A170 & \new_[43052]_ ;
  assign \new_[43057]_  = A200 & A199;
  assign \new_[43058]_  = ~A166 & \new_[43057]_ ;
  assign \new_[43059]_  = \new_[43058]_  & \new_[43053]_ ;
  assign \new_[43063]_  = ~A298 & A268;
  assign \new_[43064]_  = ~A267 & \new_[43063]_ ;
  assign \new_[43067]_  = ~A300 & A299;
  assign \new_[43070]_  = A302 & ~A301;
  assign \new_[43071]_  = \new_[43070]_  & \new_[43067]_ ;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43064]_ ;
  assign \new_[43076]_  = A167 & A168;
  assign \new_[43077]_  = A170 & \new_[43076]_ ;
  assign \new_[43081]_  = A200 & A199;
  assign \new_[43082]_  = ~A166 & \new_[43081]_ ;
  assign \new_[43083]_  = \new_[43082]_  & \new_[43077]_ ;
  assign \new_[43087]_  = A298 & ~A269;
  assign \new_[43088]_  = ~A267 & \new_[43087]_ ;
  assign \new_[43091]_  = ~A300 & ~A299;
  assign \new_[43094]_  = A302 & ~A301;
  assign \new_[43095]_  = \new_[43094]_  & \new_[43091]_ ;
  assign \new_[43096]_  = \new_[43095]_  & \new_[43088]_ ;
  assign \new_[43100]_  = A167 & A168;
  assign \new_[43101]_  = A170 & \new_[43100]_ ;
  assign \new_[43105]_  = A200 & A199;
  assign \new_[43106]_  = ~A166 & \new_[43105]_ ;
  assign \new_[43107]_  = \new_[43106]_  & \new_[43101]_ ;
  assign \new_[43111]_  = ~A298 & ~A269;
  assign \new_[43112]_  = ~A267 & \new_[43111]_ ;
  assign \new_[43115]_  = ~A300 & A299;
  assign \new_[43118]_  = A302 & ~A301;
  assign \new_[43119]_  = \new_[43118]_  & \new_[43115]_ ;
  assign \new_[43120]_  = \new_[43119]_  & \new_[43112]_ ;
  assign \new_[43124]_  = A167 & A168;
  assign \new_[43125]_  = A170 & \new_[43124]_ ;
  assign \new_[43129]_  = A200 & A199;
  assign \new_[43130]_  = ~A166 & \new_[43129]_ ;
  assign \new_[43131]_  = \new_[43130]_  & \new_[43125]_ ;
  assign \new_[43135]_  = A298 & A266;
  assign \new_[43136]_  = A265 & \new_[43135]_ ;
  assign \new_[43139]_  = ~A300 & ~A299;
  assign \new_[43142]_  = A302 & ~A301;
  assign \new_[43143]_  = \new_[43142]_  & \new_[43139]_ ;
  assign \new_[43144]_  = \new_[43143]_  & \new_[43136]_ ;
  assign \new_[43148]_  = A167 & A168;
  assign \new_[43149]_  = A170 & \new_[43148]_ ;
  assign \new_[43153]_  = A200 & A199;
  assign \new_[43154]_  = ~A166 & \new_[43153]_ ;
  assign \new_[43155]_  = \new_[43154]_  & \new_[43149]_ ;
  assign \new_[43159]_  = ~A298 & A266;
  assign \new_[43160]_  = A265 & \new_[43159]_ ;
  assign \new_[43163]_  = ~A300 & A299;
  assign \new_[43166]_  = A302 & ~A301;
  assign \new_[43167]_  = \new_[43166]_  & \new_[43163]_ ;
  assign \new_[43168]_  = \new_[43167]_  & \new_[43160]_ ;
  assign \new_[43172]_  = A167 & A168;
  assign \new_[43173]_  = A170 & \new_[43172]_ ;
  assign \new_[43177]_  = A200 & A199;
  assign \new_[43178]_  = ~A166 & \new_[43177]_ ;
  assign \new_[43179]_  = \new_[43178]_  & \new_[43173]_ ;
  assign \new_[43183]_  = A267 & A266;
  assign \new_[43184]_  = ~A265 & \new_[43183]_ ;
  assign \new_[43187]_  = A300 & A268;
  assign \new_[43190]_  = A302 & ~A301;
  assign \new_[43191]_  = \new_[43190]_  & \new_[43187]_ ;
  assign \new_[43192]_  = \new_[43191]_  & \new_[43184]_ ;
  assign \new_[43196]_  = A167 & A168;
  assign \new_[43197]_  = A170 & \new_[43196]_ ;
  assign \new_[43201]_  = A200 & A199;
  assign \new_[43202]_  = ~A166 & \new_[43201]_ ;
  assign \new_[43203]_  = \new_[43202]_  & \new_[43197]_ ;
  assign \new_[43207]_  = A267 & A266;
  assign \new_[43208]_  = ~A265 & \new_[43207]_ ;
  assign \new_[43211]_  = A300 & ~A269;
  assign \new_[43214]_  = A302 & ~A301;
  assign \new_[43215]_  = \new_[43214]_  & \new_[43211]_ ;
  assign \new_[43216]_  = \new_[43215]_  & \new_[43208]_ ;
  assign \new_[43220]_  = A167 & A168;
  assign \new_[43221]_  = A170 & \new_[43220]_ ;
  assign \new_[43225]_  = A200 & A199;
  assign \new_[43226]_  = ~A166 & \new_[43225]_ ;
  assign \new_[43227]_  = \new_[43226]_  & \new_[43221]_ ;
  assign \new_[43231]_  = ~A267 & A266;
  assign \new_[43232]_  = ~A265 & \new_[43231]_ ;
  assign \new_[43235]_  = A269 & ~A268;
  assign \new_[43238]_  = A301 & ~A300;
  assign \new_[43239]_  = \new_[43238]_  & \new_[43235]_ ;
  assign \new_[43240]_  = \new_[43239]_  & \new_[43232]_ ;
  assign \new_[43244]_  = A167 & A168;
  assign \new_[43245]_  = A170 & \new_[43244]_ ;
  assign \new_[43249]_  = A200 & A199;
  assign \new_[43250]_  = ~A166 & \new_[43249]_ ;
  assign \new_[43251]_  = \new_[43250]_  & \new_[43245]_ ;
  assign \new_[43255]_  = ~A267 & A266;
  assign \new_[43256]_  = ~A265 & \new_[43255]_ ;
  assign \new_[43259]_  = A269 & ~A268;
  assign \new_[43262]_  = ~A302 & ~A300;
  assign \new_[43263]_  = \new_[43262]_  & \new_[43259]_ ;
  assign \new_[43264]_  = \new_[43263]_  & \new_[43256]_ ;
  assign \new_[43268]_  = A167 & A168;
  assign \new_[43269]_  = A170 & \new_[43268]_ ;
  assign \new_[43273]_  = A200 & A199;
  assign \new_[43274]_  = ~A166 & \new_[43273]_ ;
  assign \new_[43275]_  = \new_[43274]_  & \new_[43269]_ ;
  assign \new_[43279]_  = ~A267 & A266;
  assign \new_[43280]_  = ~A265 & \new_[43279]_ ;
  assign \new_[43283]_  = A269 & ~A268;
  assign \new_[43286]_  = A299 & A298;
  assign \new_[43287]_  = \new_[43286]_  & \new_[43283]_ ;
  assign \new_[43288]_  = \new_[43287]_  & \new_[43280]_ ;
  assign \new_[43292]_  = A167 & A168;
  assign \new_[43293]_  = A170 & \new_[43292]_ ;
  assign \new_[43297]_  = A200 & A199;
  assign \new_[43298]_  = ~A166 & \new_[43297]_ ;
  assign \new_[43299]_  = \new_[43298]_  & \new_[43293]_ ;
  assign \new_[43303]_  = ~A267 & A266;
  assign \new_[43304]_  = ~A265 & \new_[43303]_ ;
  assign \new_[43307]_  = A269 & ~A268;
  assign \new_[43310]_  = ~A299 & ~A298;
  assign \new_[43311]_  = \new_[43310]_  & \new_[43307]_ ;
  assign \new_[43312]_  = \new_[43311]_  & \new_[43304]_ ;
  assign \new_[43316]_  = A167 & A168;
  assign \new_[43317]_  = A170 & \new_[43316]_ ;
  assign \new_[43321]_  = A200 & A199;
  assign \new_[43322]_  = ~A166 & \new_[43321]_ ;
  assign \new_[43323]_  = \new_[43322]_  & \new_[43317]_ ;
  assign \new_[43327]_  = A267 & ~A266;
  assign \new_[43328]_  = A265 & \new_[43327]_ ;
  assign \new_[43331]_  = A300 & A268;
  assign \new_[43334]_  = A302 & ~A301;
  assign \new_[43335]_  = \new_[43334]_  & \new_[43331]_ ;
  assign \new_[43336]_  = \new_[43335]_  & \new_[43328]_ ;
  assign \new_[43340]_  = A167 & A168;
  assign \new_[43341]_  = A170 & \new_[43340]_ ;
  assign \new_[43345]_  = A200 & A199;
  assign \new_[43346]_  = ~A166 & \new_[43345]_ ;
  assign \new_[43347]_  = \new_[43346]_  & \new_[43341]_ ;
  assign \new_[43351]_  = A267 & ~A266;
  assign \new_[43352]_  = A265 & \new_[43351]_ ;
  assign \new_[43355]_  = A300 & ~A269;
  assign \new_[43358]_  = A302 & ~A301;
  assign \new_[43359]_  = \new_[43358]_  & \new_[43355]_ ;
  assign \new_[43360]_  = \new_[43359]_  & \new_[43352]_ ;
  assign \new_[43364]_  = A167 & A168;
  assign \new_[43365]_  = A170 & \new_[43364]_ ;
  assign \new_[43369]_  = A200 & A199;
  assign \new_[43370]_  = ~A166 & \new_[43369]_ ;
  assign \new_[43371]_  = \new_[43370]_  & \new_[43365]_ ;
  assign \new_[43375]_  = ~A267 & ~A266;
  assign \new_[43376]_  = A265 & \new_[43375]_ ;
  assign \new_[43379]_  = A269 & ~A268;
  assign \new_[43382]_  = A301 & ~A300;
  assign \new_[43383]_  = \new_[43382]_  & \new_[43379]_ ;
  assign \new_[43384]_  = \new_[43383]_  & \new_[43376]_ ;
  assign \new_[43388]_  = A167 & A168;
  assign \new_[43389]_  = A170 & \new_[43388]_ ;
  assign \new_[43393]_  = A200 & A199;
  assign \new_[43394]_  = ~A166 & \new_[43393]_ ;
  assign \new_[43395]_  = \new_[43394]_  & \new_[43389]_ ;
  assign \new_[43399]_  = ~A267 & ~A266;
  assign \new_[43400]_  = A265 & \new_[43399]_ ;
  assign \new_[43403]_  = A269 & ~A268;
  assign \new_[43406]_  = ~A302 & ~A300;
  assign \new_[43407]_  = \new_[43406]_  & \new_[43403]_ ;
  assign \new_[43408]_  = \new_[43407]_  & \new_[43400]_ ;
  assign \new_[43412]_  = A167 & A168;
  assign \new_[43413]_  = A170 & \new_[43412]_ ;
  assign \new_[43417]_  = A200 & A199;
  assign \new_[43418]_  = ~A166 & \new_[43417]_ ;
  assign \new_[43419]_  = \new_[43418]_  & \new_[43413]_ ;
  assign \new_[43423]_  = ~A267 & ~A266;
  assign \new_[43424]_  = A265 & \new_[43423]_ ;
  assign \new_[43427]_  = A269 & ~A268;
  assign \new_[43430]_  = A299 & A298;
  assign \new_[43431]_  = \new_[43430]_  & \new_[43427]_ ;
  assign \new_[43432]_  = \new_[43431]_  & \new_[43424]_ ;
  assign \new_[43436]_  = A167 & A168;
  assign \new_[43437]_  = A170 & \new_[43436]_ ;
  assign \new_[43441]_  = A200 & A199;
  assign \new_[43442]_  = ~A166 & \new_[43441]_ ;
  assign \new_[43443]_  = \new_[43442]_  & \new_[43437]_ ;
  assign \new_[43447]_  = ~A267 & ~A266;
  assign \new_[43448]_  = A265 & \new_[43447]_ ;
  assign \new_[43451]_  = A269 & ~A268;
  assign \new_[43454]_  = ~A299 & ~A298;
  assign \new_[43455]_  = \new_[43454]_  & \new_[43451]_ ;
  assign \new_[43456]_  = \new_[43455]_  & \new_[43448]_ ;
  assign \new_[43460]_  = A167 & A168;
  assign \new_[43461]_  = A170 & \new_[43460]_ ;
  assign \new_[43465]_  = A200 & A199;
  assign \new_[43466]_  = ~A166 & \new_[43465]_ ;
  assign \new_[43467]_  = \new_[43466]_  & \new_[43461]_ ;
  assign \new_[43471]_  = A298 & ~A266;
  assign \new_[43472]_  = ~A265 & \new_[43471]_ ;
  assign \new_[43475]_  = ~A300 & ~A299;
  assign \new_[43478]_  = A302 & ~A301;
  assign \new_[43479]_  = \new_[43478]_  & \new_[43475]_ ;
  assign \new_[43480]_  = \new_[43479]_  & \new_[43472]_ ;
  assign \new_[43484]_  = A167 & A168;
  assign \new_[43485]_  = A170 & \new_[43484]_ ;
  assign \new_[43489]_  = A200 & A199;
  assign \new_[43490]_  = ~A166 & \new_[43489]_ ;
  assign \new_[43491]_  = \new_[43490]_  & \new_[43485]_ ;
  assign \new_[43495]_  = ~A298 & ~A266;
  assign \new_[43496]_  = ~A265 & \new_[43495]_ ;
  assign \new_[43499]_  = ~A300 & A299;
  assign \new_[43502]_  = A302 & ~A301;
  assign \new_[43503]_  = \new_[43502]_  & \new_[43499]_ ;
  assign \new_[43504]_  = \new_[43503]_  & \new_[43496]_ ;
  assign \new_[43508]_  = A167 & A168;
  assign \new_[43509]_  = A170 & \new_[43508]_ ;
  assign \new_[43513]_  = ~A200 & ~A199;
  assign \new_[43514]_  = ~A166 & \new_[43513]_ ;
  assign \new_[43515]_  = \new_[43514]_  & \new_[43509]_ ;
  assign \new_[43519]_  = A269 & ~A268;
  assign \new_[43520]_  = A267 & \new_[43519]_ ;
  assign \new_[43523]_  = ~A299 & A298;
  assign \new_[43526]_  = A301 & A300;
  assign \new_[43527]_  = \new_[43526]_  & \new_[43523]_ ;
  assign \new_[43528]_  = \new_[43527]_  & \new_[43520]_ ;
  assign \new_[43532]_  = A167 & A168;
  assign \new_[43533]_  = A170 & \new_[43532]_ ;
  assign \new_[43537]_  = ~A200 & ~A199;
  assign \new_[43538]_  = ~A166 & \new_[43537]_ ;
  assign \new_[43539]_  = \new_[43538]_  & \new_[43533]_ ;
  assign \new_[43543]_  = A269 & ~A268;
  assign \new_[43544]_  = A267 & \new_[43543]_ ;
  assign \new_[43547]_  = ~A299 & A298;
  assign \new_[43550]_  = ~A302 & A300;
  assign \new_[43551]_  = \new_[43550]_  & \new_[43547]_ ;
  assign \new_[43552]_  = \new_[43551]_  & \new_[43544]_ ;
  assign \new_[43556]_  = A167 & A168;
  assign \new_[43557]_  = A170 & \new_[43556]_ ;
  assign \new_[43561]_  = ~A200 & ~A199;
  assign \new_[43562]_  = ~A166 & \new_[43561]_ ;
  assign \new_[43563]_  = \new_[43562]_  & \new_[43557]_ ;
  assign \new_[43567]_  = A269 & ~A268;
  assign \new_[43568]_  = A267 & \new_[43567]_ ;
  assign \new_[43571]_  = A299 & ~A298;
  assign \new_[43574]_  = A301 & A300;
  assign \new_[43575]_  = \new_[43574]_  & \new_[43571]_ ;
  assign \new_[43576]_  = \new_[43575]_  & \new_[43568]_ ;
  assign \new_[43580]_  = A167 & A168;
  assign \new_[43581]_  = A170 & \new_[43580]_ ;
  assign \new_[43585]_  = ~A200 & ~A199;
  assign \new_[43586]_  = ~A166 & \new_[43585]_ ;
  assign \new_[43587]_  = \new_[43586]_  & \new_[43581]_ ;
  assign \new_[43591]_  = A269 & ~A268;
  assign \new_[43592]_  = A267 & \new_[43591]_ ;
  assign \new_[43595]_  = A299 & ~A298;
  assign \new_[43598]_  = ~A302 & A300;
  assign \new_[43599]_  = \new_[43598]_  & \new_[43595]_ ;
  assign \new_[43600]_  = \new_[43599]_  & \new_[43592]_ ;
  assign \new_[43604]_  = A167 & A168;
  assign \new_[43605]_  = A170 & \new_[43604]_ ;
  assign \new_[43609]_  = ~A200 & ~A199;
  assign \new_[43610]_  = ~A166 & \new_[43609]_ ;
  assign \new_[43611]_  = \new_[43610]_  & \new_[43605]_ ;
  assign \new_[43615]_  = A298 & A268;
  assign \new_[43616]_  = ~A267 & \new_[43615]_ ;
  assign \new_[43619]_  = ~A300 & ~A299;
  assign \new_[43622]_  = A302 & ~A301;
  assign \new_[43623]_  = \new_[43622]_  & \new_[43619]_ ;
  assign \new_[43624]_  = \new_[43623]_  & \new_[43616]_ ;
  assign \new_[43628]_  = A167 & A168;
  assign \new_[43629]_  = A170 & \new_[43628]_ ;
  assign \new_[43633]_  = ~A200 & ~A199;
  assign \new_[43634]_  = ~A166 & \new_[43633]_ ;
  assign \new_[43635]_  = \new_[43634]_  & \new_[43629]_ ;
  assign \new_[43639]_  = ~A298 & A268;
  assign \new_[43640]_  = ~A267 & \new_[43639]_ ;
  assign \new_[43643]_  = ~A300 & A299;
  assign \new_[43646]_  = A302 & ~A301;
  assign \new_[43647]_  = \new_[43646]_  & \new_[43643]_ ;
  assign \new_[43648]_  = \new_[43647]_  & \new_[43640]_ ;
  assign \new_[43652]_  = A167 & A168;
  assign \new_[43653]_  = A170 & \new_[43652]_ ;
  assign \new_[43657]_  = ~A200 & ~A199;
  assign \new_[43658]_  = ~A166 & \new_[43657]_ ;
  assign \new_[43659]_  = \new_[43658]_  & \new_[43653]_ ;
  assign \new_[43663]_  = A298 & ~A269;
  assign \new_[43664]_  = ~A267 & \new_[43663]_ ;
  assign \new_[43667]_  = ~A300 & ~A299;
  assign \new_[43670]_  = A302 & ~A301;
  assign \new_[43671]_  = \new_[43670]_  & \new_[43667]_ ;
  assign \new_[43672]_  = \new_[43671]_  & \new_[43664]_ ;
  assign \new_[43676]_  = A167 & A168;
  assign \new_[43677]_  = A170 & \new_[43676]_ ;
  assign \new_[43681]_  = ~A200 & ~A199;
  assign \new_[43682]_  = ~A166 & \new_[43681]_ ;
  assign \new_[43683]_  = \new_[43682]_  & \new_[43677]_ ;
  assign \new_[43687]_  = ~A298 & ~A269;
  assign \new_[43688]_  = ~A267 & \new_[43687]_ ;
  assign \new_[43691]_  = ~A300 & A299;
  assign \new_[43694]_  = A302 & ~A301;
  assign \new_[43695]_  = \new_[43694]_  & \new_[43691]_ ;
  assign \new_[43696]_  = \new_[43695]_  & \new_[43688]_ ;
  assign \new_[43700]_  = A167 & A168;
  assign \new_[43701]_  = A170 & \new_[43700]_ ;
  assign \new_[43705]_  = ~A200 & ~A199;
  assign \new_[43706]_  = ~A166 & \new_[43705]_ ;
  assign \new_[43707]_  = \new_[43706]_  & \new_[43701]_ ;
  assign \new_[43711]_  = A298 & A266;
  assign \new_[43712]_  = A265 & \new_[43711]_ ;
  assign \new_[43715]_  = ~A300 & ~A299;
  assign \new_[43718]_  = A302 & ~A301;
  assign \new_[43719]_  = \new_[43718]_  & \new_[43715]_ ;
  assign \new_[43720]_  = \new_[43719]_  & \new_[43712]_ ;
  assign \new_[43724]_  = A167 & A168;
  assign \new_[43725]_  = A170 & \new_[43724]_ ;
  assign \new_[43729]_  = ~A200 & ~A199;
  assign \new_[43730]_  = ~A166 & \new_[43729]_ ;
  assign \new_[43731]_  = \new_[43730]_  & \new_[43725]_ ;
  assign \new_[43735]_  = ~A298 & A266;
  assign \new_[43736]_  = A265 & \new_[43735]_ ;
  assign \new_[43739]_  = ~A300 & A299;
  assign \new_[43742]_  = A302 & ~A301;
  assign \new_[43743]_  = \new_[43742]_  & \new_[43739]_ ;
  assign \new_[43744]_  = \new_[43743]_  & \new_[43736]_ ;
  assign \new_[43748]_  = A167 & A168;
  assign \new_[43749]_  = A170 & \new_[43748]_ ;
  assign \new_[43753]_  = ~A200 & ~A199;
  assign \new_[43754]_  = ~A166 & \new_[43753]_ ;
  assign \new_[43755]_  = \new_[43754]_  & \new_[43749]_ ;
  assign \new_[43759]_  = A267 & A266;
  assign \new_[43760]_  = ~A265 & \new_[43759]_ ;
  assign \new_[43763]_  = A300 & A268;
  assign \new_[43766]_  = A302 & ~A301;
  assign \new_[43767]_  = \new_[43766]_  & \new_[43763]_ ;
  assign \new_[43768]_  = \new_[43767]_  & \new_[43760]_ ;
  assign \new_[43772]_  = A167 & A168;
  assign \new_[43773]_  = A170 & \new_[43772]_ ;
  assign \new_[43777]_  = ~A200 & ~A199;
  assign \new_[43778]_  = ~A166 & \new_[43777]_ ;
  assign \new_[43779]_  = \new_[43778]_  & \new_[43773]_ ;
  assign \new_[43783]_  = A267 & A266;
  assign \new_[43784]_  = ~A265 & \new_[43783]_ ;
  assign \new_[43787]_  = A300 & ~A269;
  assign \new_[43790]_  = A302 & ~A301;
  assign \new_[43791]_  = \new_[43790]_  & \new_[43787]_ ;
  assign \new_[43792]_  = \new_[43791]_  & \new_[43784]_ ;
  assign \new_[43796]_  = A167 & A168;
  assign \new_[43797]_  = A170 & \new_[43796]_ ;
  assign \new_[43801]_  = ~A200 & ~A199;
  assign \new_[43802]_  = ~A166 & \new_[43801]_ ;
  assign \new_[43803]_  = \new_[43802]_  & \new_[43797]_ ;
  assign \new_[43807]_  = ~A267 & A266;
  assign \new_[43808]_  = ~A265 & \new_[43807]_ ;
  assign \new_[43811]_  = A269 & ~A268;
  assign \new_[43814]_  = A301 & ~A300;
  assign \new_[43815]_  = \new_[43814]_  & \new_[43811]_ ;
  assign \new_[43816]_  = \new_[43815]_  & \new_[43808]_ ;
  assign \new_[43820]_  = A167 & A168;
  assign \new_[43821]_  = A170 & \new_[43820]_ ;
  assign \new_[43825]_  = ~A200 & ~A199;
  assign \new_[43826]_  = ~A166 & \new_[43825]_ ;
  assign \new_[43827]_  = \new_[43826]_  & \new_[43821]_ ;
  assign \new_[43831]_  = ~A267 & A266;
  assign \new_[43832]_  = ~A265 & \new_[43831]_ ;
  assign \new_[43835]_  = A269 & ~A268;
  assign \new_[43838]_  = ~A302 & ~A300;
  assign \new_[43839]_  = \new_[43838]_  & \new_[43835]_ ;
  assign \new_[43840]_  = \new_[43839]_  & \new_[43832]_ ;
  assign \new_[43844]_  = A167 & A168;
  assign \new_[43845]_  = A170 & \new_[43844]_ ;
  assign \new_[43849]_  = ~A200 & ~A199;
  assign \new_[43850]_  = ~A166 & \new_[43849]_ ;
  assign \new_[43851]_  = \new_[43850]_  & \new_[43845]_ ;
  assign \new_[43855]_  = ~A267 & A266;
  assign \new_[43856]_  = ~A265 & \new_[43855]_ ;
  assign \new_[43859]_  = A269 & ~A268;
  assign \new_[43862]_  = A299 & A298;
  assign \new_[43863]_  = \new_[43862]_  & \new_[43859]_ ;
  assign \new_[43864]_  = \new_[43863]_  & \new_[43856]_ ;
  assign \new_[43868]_  = A167 & A168;
  assign \new_[43869]_  = A170 & \new_[43868]_ ;
  assign \new_[43873]_  = ~A200 & ~A199;
  assign \new_[43874]_  = ~A166 & \new_[43873]_ ;
  assign \new_[43875]_  = \new_[43874]_  & \new_[43869]_ ;
  assign \new_[43879]_  = ~A267 & A266;
  assign \new_[43880]_  = ~A265 & \new_[43879]_ ;
  assign \new_[43883]_  = A269 & ~A268;
  assign \new_[43886]_  = ~A299 & ~A298;
  assign \new_[43887]_  = \new_[43886]_  & \new_[43883]_ ;
  assign \new_[43888]_  = \new_[43887]_  & \new_[43880]_ ;
  assign \new_[43892]_  = A167 & A168;
  assign \new_[43893]_  = A170 & \new_[43892]_ ;
  assign \new_[43897]_  = ~A200 & ~A199;
  assign \new_[43898]_  = ~A166 & \new_[43897]_ ;
  assign \new_[43899]_  = \new_[43898]_  & \new_[43893]_ ;
  assign \new_[43903]_  = A267 & ~A266;
  assign \new_[43904]_  = A265 & \new_[43903]_ ;
  assign \new_[43907]_  = A300 & A268;
  assign \new_[43910]_  = A302 & ~A301;
  assign \new_[43911]_  = \new_[43910]_  & \new_[43907]_ ;
  assign \new_[43912]_  = \new_[43911]_  & \new_[43904]_ ;
  assign \new_[43916]_  = A167 & A168;
  assign \new_[43917]_  = A170 & \new_[43916]_ ;
  assign \new_[43921]_  = ~A200 & ~A199;
  assign \new_[43922]_  = ~A166 & \new_[43921]_ ;
  assign \new_[43923]_  = \new_[43922]_  & \new_[43917]_ ;
  assign \new_[43927]_  = A267 & ~A266;
  assign \new_[43928]_  = A265 & \new_[43927]_ ;
  assign \new_[43931]_  = A300 & ~A269;
  assign \new_[43934]_  = A302 & ~A301;
  assign \new_[43935]_  = \new_[43934]_  & \new_[43931]_ ;
  assign \new_[43936]_  = \new_[43935]_  & \new_[43928]_ ;
  assign \new_[43940]_  = A167 & A168;
  assign \new_[43941]_  = A170 & \new_[43940]_ ;
  assign \new_[43945]_  = ~A200 & ~A199;
  assign \new_[43946]_  = ~A166 & \new_[43945]_ ;
  assign \new_[43947]_  = \new_[43946]_  & \new_[43941]_ ;
  assign \new_[43951]_  = ~A267 & ~A266;
  assign \new_[43952]_  = A265 & \new_[43951]_ ;
  assign \new_[43955]_  = A269 & ~A268;
  assign \new_[43958]_  = A301 & ~A300;
  assign \new_[43959]_  = \new_[43958]_  & \new_[43955]_ ;
  assign \new_[43960]_  = \new_[43959]_  & \new_[43952]_ ;
  assign \new_[43964]_  = A167 & A168;
  assign \new_[43965]_  = A170 & \new_[43964]_ ;
  assign \new_[43969]_  = ~A200 & ~A199;
  assign \new_[43970]_  = ~A166 & \new_[43969]_ ;
  assign \new_[43971]_  = \new_[43970]_  & \new_[43965]_ ;
  assign \new_[43975]_  = ~A267 & ~A266;
  assign \new_[43976]_  = A265 & \new_[43975]_ ;
  assign \new_[43979]_  = A269 & ~A268;
  assign \new_[43982]_  = ~A302 & ~A300;
  assign \new_[43983]_  = \new_[43982]_  & \new_[43979]_ ;
  assign \new_[43984]_  = \new_[43983]_  & \new_[43976]_ ;
  assign \new_[43988]_  = A167 & A168;
  assign \new_[43989]_  = A170 & \new_[43988]_ ;
  assign \new_[43993]_  = ~A200 & ~A199;
  assign \new_[43994]_  = ~A166 & \new_[43993]_ ;
  assign \new_[43995]_  = \new_[43994]_  & \new_[43989]_ ;
  assign \new_[43999]_  = ~A267 & ~A266;
  assign \new_[44000]_  = A265 & \new_[43999]_ ;
  assign \new_[44003]_  = A269 & ~A268;
  assign \new_[44006]_  = A299 & A298;
  assign \new_[44007]_  = \new_[44006]_  & \new_[44003]_ ;
  assign \new_[44008]_  = \new_[44007]_  & \new_[44000]_ ;
  assign \new_[44012]_  = A167 & A168;
  assign \new_[44013]_  = A170 & \new_[44012]_ ;
  assign \new_[44017]_  = ~A200 & ~A199;
  assign \new_[44018]_  = ~A166 & \new_[44017]_ ;
  assign \new_[44019]_  = \new_[44018]_  & \new_[44013]_ ;
  assign \new_[44023]_  = ~A267 & ~A266;
  assign \new_[44024]_  = A265 & \new_[44023]_ ;
  assign \new_[44027]_  = A269 & ~A268;
  assign \new_[44030]_  = ~A299 & ~A298;
  assign \new_[44031]_  = \new_[44030]_  & \new_[44027]_ ;
  assign \new_[44032]_  = \new_[44031]_  & \new_[44024]_ ;
  assign \new_[44036]_  = A167 & A168;
  assign \new_[44037]_  = A170 & \new_[44036]_ ;
  assign \new_[44041]_  = ~A200 & ~A199;
  assign \new_[44042]_  = ~A166 & \new_[44041]_ ;
  assign \new_[44043]_  = \new_[44042]_  & \new_[44037]_ ;
  assign \new_[44047]_  = A298 & ~A266;
  assign \new_[44048]_  = ~A265 & \new_[44047]_ ;
  assign \new_[44051]_  = ~A300 & ~A299;
  assign \new_[44054]_  = A302 & ~A301;
  assign \new_[44055]_  = \new_[44054]_  & \new_[44051]_ ;
  assign \new_[44056]_  = \new_[44055]_  & \new_[44048]_ ;
  assign \new_[44060]_  = A167 & A168;
  assign \new_[44061]_  = A170 & \new_[44060]_ ;
  assign \new_[44065]_  = ~A200 & ~A199;
  assign \new_[44066]_  = ~A166 & \new_[44065]_ ;
  assign \new_[44067]_  = \new_[44066]_  & \new_[44061]_ ;
  assign \new_[44071]_  = ~A298 & ~A266;
  assign \new_[44072]_  = ~A265 & \new_[44071]_ ;
  assign \new_[44075]_  = ~A300 & A299;
  assign \new_[44078]_  = A302 & ~A301;
  assign \new_[44079]_  = \new_[44078]_  & \new_[44075]_ ;
  assign \new_[44080]_  = \new_[44079]_  & \new_[44072]_ ;
  assign \new_[44084]_  = ~A167 & A168;
  assign \new_[44085]_  = A170 & \new_[44084]_ ;
  assign \new_[44089]_  = ~A202 & A201;
  assign \new_[44090]_  = A166 & \new_[44089]_ ;
  assign \new_[44091]_  = \new_[44090]_  & \new_[44085]_ ;
  assign \new_[44095]_  = A268 & ~A267;
  assign \new_[44096]_  = A203 & \new_[44095]_ ;
  assign \new_[44099]_  = ~A299 & A298;
  assign \new_[44102]_  = A301 & A300;
  assign \new_[44103]_  = \new_[44102]_  & \new_[44099]_ ;
  assign \new_[44104]_  = \new_[44103]_  & \new_[44096]_ ;
  assign \new_[44108]_  = ~A167 & A168;
  assign \new_[44109]_  = A170 & \new_[44108]_ ;
  assign \new_[44113]_  = ~A202 & A201;
  assign \new_[44114]_  = A166 & \new_[44113]_ ;
  assign \new_[44115]_  = \new_[44114]_  & \new_[44109]_ ;
  assign \new_[44119]_  = A268 & ~A267;
  assign \new_[44120]_  = A203 & \new_[44119]_ ;
  assign \new_[44123]_  = ~A299 & A298;
  assign \new_[44126]_  = ~A302 & A300;
  assign \new_[44127]_  = \new_[44126]_  & \new_[44123]_ ;
  assign \new_[44128]_  = \new_[44127]_  & \new_[44120]_ ;
  assign \new_[44132]_  = ~A167 & A168;
  assign \new_[44133]_  = A170 & \new_[44132]_ ;
  assign \new_[44137]_  = ~A202 & A201;
  assign \new_[44138]_  = A166 & \new_[44137]_ ;
  assign \new_[44139]_  = \new_[44138]_  & \new_[44133]_ ;
  assign \new_[44143]_  = A268 & ~A267;
  assign \new_[44144]_  = A203 & \new_[44143]_ ;
  assign \new_[44147]_  = A299 & ~A298;
  assign \new_[44150]_  = A301 & A300;
  assign \new_[44151]_  = \new_[44150]_  & \new_[44147]_ ;
  assign \new_[44152]_  = \new_[44151]_  & \new_[44144]_ ;
  assign \new_[44156]_  = ~A167 & A168;
  assign \new_[44157]_  = A170 & \new_[44156]_ ;
  assign \new_[44161]_  = ~A202 & A201;
  assign \new_[44162]_  = A166 & \new_[44161]_ ;
  assign \new_[44163]_  = \new_[44162]_  & \new_[44157]_ ;
  assign \new_[44167]_  = A268 & ~A267;
  assign \new_[44168]_  = A203 & \new_[44167]_ ;
  assign \new_[44171]_  = A299 & ~A298;
  assign \new_[44174]_  = ~A302 & A300;
  assign \new_[44175]_  = \new_[44174]_  & \new_[44171]_ ;
  assign \new_[44176]_  = \new_[44175]_  & \new_[44168]_ ;
  assign \new_[44180]_  = ~A167 & A168;
  assign \new_[44181]_  = A170 & \new_[44180]_ ;
  assign \new_[44185]_  = ~A202 & A201;
  assign \new_[44186]_  = A166 & \new_[44185]_ ;
  assign \new_[44187]_  = \new_[44186]_  & \new_[44181]_ ;
  assign \new_[44191]_  = ~A269 & ~A267;
  assign \new_[44192]_  = A203 & \new_[44191]_ ;
  assign \new_[44195]_  = ~A299 & A298;
  assign \new_[44198]_  = A301 & A300;
  assign \new_[44199]_  = \new_[44198]_  & \new_[44195]_ ;
  assign \new_[44200]_  = \new_[44199]_  & \new_[44192]_ ;
  assign \new_[44204]_  = ~A167 & A168;
  assign \new_[44205]_  = A170 & \new_[44204]_ ;
  assign \new_[44209]_  = ~A202 & A201;
  assign \new_[44210]_  = A166 & \new_[44209]_ ;
  assign \new_[44211]_  = \new_[44210]_  & \new_[44205]_ ;
  assign \new_[44215]_  = ~A269 & ~A267;
  assign \new_[44216]_  = A203 & \new_[44215]_ ;
  assign \new_[44219]_  = ~A299 & A298;
  assign \new_[44222]_  = ~A302 & A300;
  assign \new_[44223]_  = \new_[44222]_  & \new_[44219]_ ;
  assign \new_[44224]_  = \new_[44223]_  & \new_[44216]_ ;
  assign \new_[44228]_  = ~A167 & A168;
  assign \new_[44229]_  = A170 & \new_[44228]_ ;
  assign \new_[44233]_  = ~A202 & A201;
  assign \new_[44234]_  = A166 & \new_[44233]_ ;
  assign \new_[44235]_  = \new_[44234]_  & \new_[44229]_ ;
  assign \new_[44239]_  = ~A269 & ~A267;
  assign \new_[44240]_  = A203 & \new_[44239]_ ;
  assign \new_[44243]_  = A299 & ~A298;
  assign \new_[44246]_  = A301 & A300;
  assign \new_[44247]_  = \new_[44246]_  & \new_[44243]_ ;
  assign \new_[44248]_  = \new_[44247]_  & \new_[44240]_ ;
  assign \new_[44252]_  = ~A167 & A168;
  assign \new_[44253]_  = A170 & \new_[44252]_ ;
  assign \new_[44257]_  = ~A202 & A201;
  assign \new_[44258]_  = A166 & \new_[44257]_ ;
  assign \new_[44259]_  = \new_[44258]_  & \new_[44253]_ ;
  assign \new_[44263]_  = ~A269 & ~A267;
  assign \new_[44264]_  = A203 & \new_[44263]_ ;
  assign \new_[44267]_  = A299 & ~A298;
  assign \new_[44270]_  = ~A302 & A300;
  assign \new_[44271]_  = \new_[44270]_  & \new_[44267]_ ;
  assign \new_[44272]_  = \new_[44271]_  & \new_[44264]_ ;
  assign \new_[44276]_  = ~A167 & A168;
  assign \new_[44277]_  = A170 & \new_[44276]_ ;
  assign \new_[44281]_  = ~A202 & A201;
  assign \new_[44282]_  = A166 & \new_[44281]_ ;
  assign \new_[44283]_  = \new_[44282]_  & \new_[44277]_ ;
  assign \new_[44287]_  = A266 & A265;
  assign \new_[44288]_  = A203 & \new_[44287]_ ;
  assign \new_[44291]_  = ~A299 & A298;
  assign \new_[44294]_  = A301 & A300;
  assign \new_[44295]_  = \new_[44294]_  & \new_[44291]_ ;
  assign \new_[44296]_  = \new_[44295]_  & \new_[44288]_ ;
  assign \new_[44300]_  = ~A167 & A168;
  assign \new_[44301]_  = A170 & \new_[44300]_ ;
  assign \new_[44305]_  = ~A202 & A201;
  assign \new_[44306]_  = A166 & \new_[44305]_ ;
  assign \new_[44307]_  = \new_[44306]_  & \new_[44301]_ ;
  assign \new_[44311]_  = A266 & A265;
  assign \new_[44312]_  = A203 & \new_[44311]_ ;
  assign \new_[44315]_  = ~A299 & A298;
  assign \new_[44318]_  = ~A302 & A300;
  assign \new_[44319]_  = \new_[44318]_  & \new_[44315]_ ;
  assign \new_[44320]_  = \new_[44319]_  & \new_[44312]_ ;
  assign \new_[44324]_  = ~A167 & A168;
  assign \new_[44325]_  = A170 & \new_[44324]_ ;
  assign \new_[44329]_  = ~A202 & A201;
  assign \new_[44330]_  = A166 & \new_[44329]_ ;
  assign \new_[44331]_  = \new_[44330]_  & \new_[44325]_ ;
  assign \new_[44335]_  = A266 & A265;
  assign \new_[44336]_  = A203 & \new_[44335]_ ;
  assign \new_[44339]_  = A299 & ~A298;
  assign \new_[44342]_  = A301 & A300;
  assign \new_[44343]_  = \new_[44342]_  & \new_[44339]_ ;
  assign \new_[44344]_  = \new_[44343]_  & \new_[44336]_ ;
  assign \new_[44348]_  = ~A167 & A168;
  assign \new_[44349]_  = A170 & \new_[44348]_ ;
  assign \new_[44353]_  = ~A202 & A201;
  assign \new_[44354]_  = A166 & \new_[44353]_ ;
  assign \new_[44355]_  = \new_[44354]_  & \new_[44349]_ ;
  assign \new_[44359]_  = A266 & A265;
  assign \new_[44360]_  = A203 & \new_[44359]_ ;
  assign \new_[44363]_  = A299 & ~A298;
  assign \new_[44366]_  = ~A302 & A300;
  assign \new_[44367]_  = \new_[44366]_  & \new_[44363]_ ;
  assign \new_[44368]_  = \new_[44367]_  & \new_[44360]_ ;
  assign \new_[44372]_  = ~A167 & A168;
  assign \new_[44373]_  = A170 & \new_[44372]_ ;
  assign \new_[44377]_  = ~A202 & A201;
  assign \new_[44378]_  = A166 & \new_[44377]_ ;
  assign \new_[44379]_  = \new_[44378]_  & \new_[44373]_ ;
  assign \new_[44383]_  = A266 & ~A265;
  assign \new_[44384]_  = A203 & \new_[44383]_ ;
  assign \new_[44387]_  = A268 & A267;
  assign \new_[44390]_  = A301 & ~A300;
  assign \new_[44391]_  = \new_[44390]_  & \new_[44387]_ ;
  assign \new_[44392]_  = \new_[44391]_  & \new_[44384]_ ;
  assign \new_[44396]_  = ~A167 & A168;
  assign \new_[44397]_  = A170 & \new_[44396]_ ;
  assign \new_[44401]_  = ~A202 & A201;
  assign \new_[44402]_  = A166 & \new_[44401]_ ;
  assign \new_[44403]_  = \new_[44402]_  & \new_[44397]_ ;
  assign \new_[44407]_  = A266 & ~A265;
  assign \new_[44408]_  = A203 & \new_[44407]_ ;
  assign \new_[44411]_  = A268 & A267;
  assign \new_[44414]_  = ~A302 & ~A300;
  assign \new_[44415]_  = \new_[44414]_  & \new_[44411]_ ;
  assign \new_[44416]_  = \new_[44415]_  & \new_[44408]_ ;
  assign \new_[44420]_  = ~A167 & A168;
  assign \new_[44421]_  = A170 & \new_[44420]_ ;
  assign \new_[44425]_  = ~A202 & A201;
  assign \new_[44426]_  = A166 & \new_[44425]_ ;
  assign \new_[44427]_  = \new_[44426]_  & \new_[44421]_ ;
  assign \new_[44431]_  = A266 & ~A265;
  assign \new_[44432]_  = A203 & \new_[44431]_ ;
  assign \new_[44435]_  = A268 & A267;
  assign \new_[44438]_  = A299 & A298;
  assign \new_[44439]_  = \new_[44438]_  & \new_[44435]_ ;
  assign \new_[44440]_  = \new_[44439]_  & \new_[44432]_ ;
  assign \new_[44444]_  = ~A167 & A168;
  assign \new_[44445]_  = A170 & \new_[44444]_ ;
  assign \new_[44449]_  = ~A202 & A201;
  assign \new_[44450]_  = A166 & \new_[44449]_ ;
  assign \new_[44451]_  = \new_[44450]_  & \new_[44445]_ ;
  assign \new_[44455]_  = A266 & ~A265;
  assign \new_[44456]_  = A203 & \new_[44455]_ ;
  assign \new_[44459]_  = A268 & A267;
  assign \new_[44462]_  = ~A299 & ~A298;
  assign \new_[44463]_  = \new_[44462]_  & \new_[44459]_ ;
  assign \new_[44464]_  = \new_[44463]_  & \new_[44456]_ ;
  assign \new_[44468]_  = ~A167 & A168;
  assign \new_[44469]_  = A170 & \new_[44468]_ ;
  assign \new_[44473]_  = ~A202 & A201;
  assign \new_[44474]_  = A166 & \new_[44473]_ ;
  assign \new_[44475]_  = \new_[44474]_  & \new_[44469]_ ;
  assign \new_[44479]_  = A266 & ~A265;
  assign \new_[44480]_  = A203 & \new_[44479]_ ;
  assign \new_[44483]_  = ~A269 & A267;
  assign \new_[44486]_  = A301 & ~A300;
  assign \new_[44487]_  = \new_[44486]_  & \new_[44483]_ ;
  assign \new_[44488]_  = \new_[44487]_  & \new_[44480]_ ;
  assign \new_[44492]_  = ~A167 & A168;
  assign \new_[44493]_  = A170 & \new_[44492]_ ;
  assign \new_[44497]_  = ~A202 & A201;
  assign \new_[44498]_  = A166 & \new_[44497]_ ;
  assign \new_[44499]_  = \new_[44498]_  & \new_[44493]_ ;
  assign \new_[44503]_  = A266 & ~A265;
  assign \new_[44504]_  = A203 & \new_[44503]_ ;
  assign \new_[44507]_  = ~A269 & A267;
  assign \new_[44510]_  = ~A302 & ~A300;
  assign \new_[44511]_  = \new_[44510]_  & \new_[44507]_ ;
  assign \new_[44512]_  = \new_[44511]_  & \new_[44504]_ ;
  assign \new_[44516]_  = ~A167 & A168;
  assign \new_[44517]_  = A170 & \new_[44516]_ ;
  assign \new_[44521]_  = ~A202 & A201;
  assign \new_[44522]_  = A166 & \new_[44521]_ ;
  assign \new_[44523]_  = \new_[44522]_  & \new_[44517]_ ;
  assign \new_[44527]_  = A266 & ~A265;
  assign \new_[44528]_  = A203 & \new_[44527]_ ;
  assign \new_[44531]_  = ~A269 & A267;
  assign \new_[44534]_  = A299 & A298;
  assign \new_[44535]_  = \new_[44534]_  & \new_[44531]_ ;
  assign \new_[44536]_  = \new_[44535]_  & \new_[44528]_ ;
  assign \new_[44540]_  = ~A167 & A168;
  assign \new_[44541]_  = A170 & \new_[44540]_ ;
  assign \new_[44545]_  = ~A202 & A201;
  assign \new_[44546]_  = A166 & \new_[44545]_ ;
  assign \new_[44547]_  = \new_[44546]_  & \new_[44541]_ ;
  assign \new_[44551]_  = A266 & ~A265;
  assign \new_[44552]_  = A203 & \new_[44551]_ ;
  assign \new_[44555]_  = ~A269 & A267;
  assign \new_[44558]_  = ~A299 & ~A298;
  assign \new_[44559]_  = \new_[44558]_  & \new_[44555]_ ;
  assign \new_[44560]_  = \new_[44559]_  & \new_[44552]_ ;
  assign \new_[44564]_  = ~A167 & A168;
  assign \new_[44565]_  = A170 & \new_[44564]_ ;
  assign \new_[44569]_  = ~A202 & A201;
  assign \new_[44570]_  = A166 & \new_[44569]_ ;
  assign \new_[44571]_  = \new_[44570]_  & \new_[44565]_ ;
  assign \new_[44575]_  = ~A266 & A265;
  assign \new_[44576]_  = A203 & \new_[44575]_ ;
  assign \new_[44579]_  = A268 & A267;
  assign \new_[44582]_  = A301 & ~A300;
  assign \new_[44583]_  = \new_[44582]_  & \new_[44579]_ ;
  assign \new_[44584]_  = \new_[44583]_  & \new_[44576]_ ;
  assign \new_[44588]_  = ~A167 & A168;
  assign \new_[44589]_  = A170 & \new_[44588]_ ;
  assign \new_[44593]_  = ~A202 & A201;
  assign \new_[44594]_  = A166 & \new_[44593]_ ;
  assign \new_[44595]_  = \new_[44594]_  & \new_[44589]_ ;
  assign \new_[44599]_  = ~A266 & A265;
  assign \new_[44600]_  = A203 & \new_[44599]_ ;
  assign \new_[44603]_  = A268 & A267;
  assign \new_[44606]_  = ~A302 & ~A300;
  assign \new_[44607]_  = \new_[44606]_  & \new_[44603]_ ;
  assign \new_[44608]_  = \new_[44607]_  & \new_[44600]_ ;
  assign \new_[44612]_  = ~A167 & A168;
  assign \new_[44613]_  = A170 & \new_[44612]_ ;
  assign \new_[44617]_  = ~A202 & A201;
  assign \new_[44618]_  = A166 & \new_[44617]_ ;
  assign \new_[44619]_  = \new_[44618]_  & \new_[44613]_ ;
  assign \new_[44623]_  = ~A266 & A265;
  assign \new_[44624]_  = A203 & \new_[44623]_ ;
  assign \new_[44627]_  = A268 & A267;
  assign \new_[44630]_  = A299 & A298;
  assign \new_[44631]_  = \new_[44630]_  & \new_[44627]_ ;
  assign \new_[44632]_  = \new_[44631]_  & \new_[44624]_ ;
  assign \new_[44636]_  = ~A167 & A168;
  assign \new_[44637]_  = A170 & \new_[44636]_ ;
  assign \new_[44641]_  = ~A202 & A201;
  assign \new_[44642]_  = A166 & \new_[44641]_ ;
  assign \new_[44643]_  = \new_[44642]_  & \new_[44637]_ ;
  assign \new_[44647]_  = ~A266 & A265;
  assign \new_[44648]_  = A203 & \new_[44647]_ ;
  assign \new_[44651]_  = A268 & A267;
  assign \new_[44654]_  = ~A299 & ~A298;
  assign \new_[44655]_  = \new_[44654]_  & \new_[44651]_ ;
  assign \new_[44656]_  = \new_[44655]_  & \new_[44648]_ ;
  assign \new_[44660]_  = ~A167 & A168;
  assign \new_[44661]_  = A170 & \new_[44660]_ ;
  assign \new_[44665]_  = ~A202 & A201;
  assign \new_[44666]_  = A166 & \new_[44665]_ ;
  assign \new_[44667]_  = \new_[44666]_  & \new_[44661]_ ;
  assign \new_[44671]_  = ~A266 & A265;
  assign \new_[44672]_  = A203 & \new_[44671]_ ;
  assign \new_[44675]_  = ~A269 & A267;
  assign \new_[44678]_  = A301 & ~A300;
  assign \new_[44679]_  = \new_[44678]_  & \new_[44675]_ ;
  assign \new_[44680]_  = \new_[44679]_  & \new_[44672]_ ;
  assign \new_[44684]_  = ~A167 & A168;
  assign \new_[44685]_  = A170 & \new_[44684]_ ;
  assign \new_[44689]_  = ~A202 & A201;
  assign \new_[44690]_  = A166 & \new_[44689]_ ;
  assign \new_[44691]_  = \new_[44690]_  & \new_[44685]_ ;
  assign \new_[44695]_  = ~A266 & A265;
  assign \new_[44696]_  = A203 & \new_[44695]_ ;
  assign \new_[44699]_  = ~A269 & A267;
  assign \new_[44702]_  = ~A302 & ~A300;
  assign \new_[44703]_  = \new_[44702]_  & \new_[44699]_ ;
  assign \new_[44704]_  = \new_[44703]_  & \new_[44696]_ ;
  assign \new_[44708]_  = ~A167 & A168;
  assign \new_[44709]_  = A170 & \new_[44708]_ ;
  assign \new_[44713]_  = ~A202 & A201;
  assign \new_[44714]_  = A166 & \new_[44713]_ ;
  assign \new_[44715]_  = \new_[44714]_  & \new_[44709]_ ;
  assign \new_[44719]_  = ~A266 & A265;
  assign \new_[44720]_  = A203 & \new_[44719]_ ;
  assign \new_[44723]_  = ~A269 & A267;
  assign \new_[44726]_  = A299 & A298;
  assign \new_[44727]_  = \new_[44726]_  & \new_[44723]_ ;
  assign \new_[44728]_  = \new_[44727]_  & \new_[44720]_ ;
  assign \new_[44732]_  = ~A167 & A168;
  assign \new_[44733]_  = A170 & \new_[44732]_ ;
  assign \new_[44737]_  = ~A202 & A201;
  assign \new_[44738]_  = A166 & \new_[44737]_ ;
  assign \new_[44739]_  = \new_[44738]_  & \new_[44733]_ ;
  assign \new_[44743]_  = ~A266 & A265;
  assign \new_[44744]_  = A203 & \new_[44743]_ ;
  assign \new_[44747]_  = ~A269 & A267;
  assign \new_[44750]_  = ~A299 & ~A298;
  assign \new_[44751]_  = \new_[44750]_  & \new_[44747]_ ;
  assign \new_[44752]_  = \new_[44751]_  & \new_[44744]_ ;
  assign \new_[44756]_  = ~A167 & A168;
  assign \new_[44757]_  = A170 & \new_[44756]_ ;
  assign \new_[44761]_  = ~A202 & A201;
  assign \new_[44762]_  = A166 & \new_[44761]_ ;
  assign \new_[44763]_  = \new_[44762]_  & \new_[44757]_ ;
  assign \new_[44767]_  = ~A266 & ~A265;
  assign \new_[44768]_  = A203 & \new_[44767]_ ;
  assign \new_[44771]_  = ~A299 & A298;
  assign \new_[44774]_  = A301 & A300;
  assign \new_[44775]_  = \new_[44774]_  & \new_[44771]_ ;
  assign \new_[44776]_  = \new_[44775]_  & \new_[44768]_ ;
  assign \new_[44780]_  = ~A167 & A168;
  assign \new_[44781]_  = A170 & \new_[44780]_ ;
  assign \new_[44785]_  = ~A202 & A201;
  assign \new_[44786]_  = A166 & \new_[44785]_ ;
  assign \new_[44787]_  = \new_[44786]_  & \new_[44781]_ ;
  assign \new_[44791]_  = ~A266 & ~A265;
  assign \new_[44792]_  = A203 & \new_[44791]_ ;
  assign \new_[44795]_  = ~A299 & A298;
  assign \new_[44798]_  = ~A302 & A300;
  assign \new_[44799]_  = \new_[44798]_  & \new_[44795]_ ;
  assign \new_[44800]_  = \new_[44799]_  & \new_[44792]_ ;
  assign \new_[44804]_  = ~A167 & A168;
  assign \new_[44805]_  = A170 & \new_[44804]_ ;
  assign \new_[44809]_  = ~A202 & A201;
  assign \new_[44810]_  = A166 & \new_[44809]_ ;
  assign \new_[44811]_  = \new_[44810]_  & \new_[44805]_ ;
  assign \new_[44815]_  = ~A266 & ~A265;
  assign \new_[44816]_  = A203 & \new_[44815]_ ;
  assign \new_[44819]_  = A299 & ~A298;
  assign \new_[44822]_  = A301 & A300;
  assign \new_[44823]_  = \new_[44822]_  & \new_[44819]_ ;
  assign \new_[44824]_  = \new_[44823]_  & \new_[44816]_ ;
  assign \new_[44828]_  = ~A167 & A168;
  assign \new_[44829]_  = A170 & \new_[44828]_ ;
  assign \new_[44833]_  = ~A202 & A201;
  assign \new_[44834]_  = A166 & \new_[44833]_ ;
  assign \new_[44835]_  = \new_[44834]_  & \new_[44829]_ ;
  assign \new_[44839]_  = ~A266 & ~A265;
  assign \new_[44840]_  = A203 & \new_[44839]_ ;
  assign \new_[44843]_  = A299 & ~A298;
  assign \new_[44846]_  = ~A302 & A300;
  assign \new_[44847]_  = \new_[44846]_  & \new_[44843]_ ;
  assign \new_[44848]_  = \new_[44847]_  & \new_[44840]_ ;
  assign \new_[44852]_  = ~A167 & A168;
  assign \new_[44853]_  = A170 & \new_[44852]_ ;
  assign \new_[44857]_  = A202 & ~A201;
  assign \new_[44858]_  = A166 & \new_[44857]_ ;
  assign \new_[44859]_  = \new_[44858]_  & \new_[44853]_ ;
  assign \new_[44863]_  = A269 & ~A268;
  assign \new_[44864]_  = A267 & \new_[44863]_ ;
  assign \new_[44867]_  = ~A299 & A298;
  assign \new_[44870]_  = A301 & A300;
  assign \new_[44871]_  = \new_[44870]_  & \new_[44867]_ ;
  assign \new_[44872]_  = \new_[44871]_  & \new_[44864]_ ;
  assign \new_[44876]_  = ~A167 & A168;
  assign \new_[44877]_  = A170 & \new_[44876]_ ;
  assign \new_[44881]_  = A202 & ~A201;
  assign \new_[44882]_  = A166 & \new_[44881]_ ;
  assign \new_[44883]_  = \new_[44882]_  & \new_[44877]_ ;
  assign \new_[44887]_  = A269 & ~A268;
  assign \new_[44888]_  = A267 & \new_[44887]_ ;
  assign \new_[44891]_  = ~A299 & A298;
  assign \new_[44894]_  = ~A302 & A300;
  assign \new_[44895]_  = \new_[44894]_  & \new_[44891]_ ;
  assign \new_[44896]_  = \new_[44895]_  & \new_[44888]_ ;
  assign \new_[44900]_  = ~A167 & A168;
  assign \new_[44901]_  = A170 & \new_[44900]_ ;
  assign \new_[44905]_  = A202 & ~A201;
  assign \new_[44906]_  = A166 & \new_[44905]_ ;
  assign \new_[44907]_  = \new_[44906]_  & \new_[44901]_ ;
  assign \new_[44911]_  = A269 & ~A268;
  assign \new_[44912]_  = A267 & \new_[44911]_ ;
  assign \new_[44915]_  = A299 & ~A298;
  assign \new_[44918]_  = A301 & A300;
  assign \new_[44919]_  = \new_[44918]_  & \new_[44915]_ ;
  assign \new_[44920]_  = \new_[44919]_  & \new_[44912]_ ;
  assign \new_[44924]_  = ~A167 & A168;
  assign \new_[44925]_  = A170 & \new_[44924]_ ;
  assign \new_[44929]_  = A202 & ~A201;
  assign \new_[44930]_  = A166 & \new_[44929]_ ;
  assign \new_[44931]_  = \new_[44930]_  & \new_[44925]_ ;
  assign \new_[44935]_  = A269 & ~A268;
  assign \new_[44936]_  = A267 & \new_[44935]_ ;
  assign \new_[44939]_  = A299 & ~A298;
  assign \new_[44942]_  = ~A302 & A300;
  assign \new_[44943]_  = \new_[44942]_  & \new_[44939]_ ;
  assign \new_[44944]_  = \new_[44943]_  & \new_[44936]_ ;
  assign \new_[44948]_  = ~A167 & A168;
  assign \new_[44949]_  = A170 & \new_[44948]_ ;
  assign \new_[44953]_  = A202 & ~A201;
  assign \new_[44954]_  = A166 & \new_[44953]_ ;
  assign \new_[44955]_  = \new_[44954]_  & \new_[44949]_ ;
  assign \new_[44959]_  = A298 & A268;
  assign \new_[44960]_  = ~A267 & \new_[44959]_ ;
  assign \new_[44963]_  = ~A300 & ~A299;
  assign \new_[44966]_  = A302 & ~A301;
  assign \new_[44967]_  = \new_[44966]_  & \new_[44963]_ ;
  assign \new_[44968]_  = \new_[44967]_  & \new_[44960]_ ;
  assign \new_[44972]_  = ~A167 & A168;
  assign \new_[44973]_  = A170 & \new_[44972]_ ;
  assign \new_[44977]_  = A202 & ~A201;
  assign \new_[44978]_  = A166 & \new_[44977]_ ;
  assign \new_[44979]_  = \new_[44978]_  & \new_[44973]_ ;
  assign \new_[44983]_  = ~A298 & A268;
  assign \new_[44984]_  = ~A267 & \new_[44983]_ ;
  assign \new_[44987]_  = ~A300 & A299;
  assign \new_[44990]_  = A302 & ~A301;
  assign \new_[44991]_  = \new_[44990]_  & \new_[44987]_ ;
  assign \new_[44992]_  = \new_[44991]_  & \new_[44984]_ ;
  assign \new_[44996]_  = ~A167 & A168;
  assign \new_[44997]_  = A170 & \new_[44996]_ ;
  assign \new_[45001]_  = A202 & ~A201;
  assign \new_[45002]_  = A166 & \new_[45001]_ ;
  assign \new_[45003]_  = \new_[45002]_  & \new_[44997]_ ;
  assign \new_[45007]_  = A298 & ~A269;
  assign \new_[45008]_  = ~A267 & \new_[45007]_ ;
  assign \new_[45011]_  = ~A300 & ~A299;
  assign \new_[45014]_  = A302 & ~A301;
  assign \new_[45015]_  = \new_[45014]_  & \new_[45011]_ ;
  assign \new_[45016]_  = \new_[45015]_  & \new_[45008]_ ;
  assign \new_[45020]_  = ~A167 & A168;
  assign \new_[45021]_  = A170 & \new_[45020]_ ;
  assign \new_[45025]_  = A202 & ~A201;
  assign \new_[45026]_  = A166 & \new_[45025]_ ;
  assign \new_[45027]_  = \new_[45026]_  & \new_[45021]_ ;
  assign \new_[45031]_  = ~A298 & ~A269;
  assign \new_[45032]_  = ~A267 & \new_[45031]_ ;
  assign \new_[45035]_  = ~A300 & A299;
  assign \new_[45038]_  = A302 & ~A301;
  assign \new_[45039]_  = \new_[45038]_  & \new_[45035]_ ;
  assign \new_[45040]_  = \new_[45039]_  & \new_[45032]_ ;
  assign \new_[45044]_  = ~A167 & A168;
  assign \new_[45045]_  = A170 & \new_[45044]_ ;
  assign \new_[45049]_  = A202 & ~A201;
  assign \new_[45050]_  = A166 & \new_[45049]_ ;
  assign \new_[45051]_  = \new_[45050]_  & \new_[45045]_ ;
  assign \new_[45055]_  = A298 & A266;
  assign \new_[45056]_  = A265 & \new_[45055]_ ;
  assign \new_[45059]_  = ~A300 & ~A299;
  assign \new_[45062]_  = A302 & ~A301;
  assign \new_[45063]_  = \new_[45062]_  & \new_[45059]_ ;
  assign \new_[45064]_  = \new_[45063]_  & \new_[45056]_ ;
  assign \new_[45068]_  = ~A167 & A168;
  assign \new_[45069]_  = A170 & \new_[45068]_ ;
  assign \new_[45073]_  = A202 & ~A201;
  assign \new_[45074]_  = A166 & \new_[45073]_ ;
  assign \new_[45075]_  = \new_[45074]_  & \new_[45069]_ ;
  assign \new_[45079]_  = ~A298 & A266;
  assign \new_[45080]_  = A265 & \new_[45079]_ ;
  assign \new_[45083]_  = ~A300 & A299;
  assign \new_[45086]_  = A302 & ~A301;
  assign \new_[45087]_  = \new_[45086]_  & \new_[45083]_ ;
  assign \new_[45088]_  = \new_[45087]_  & \new_[45080]_ ;
  assign \new_[45092]_  = ~A167 & A168;
  assign \new_[45093]_  = A170 & \new_[45092]_ ;
  assign \new_[45097]_  = A202 & ~A201;
  assign \new_[45098]_  = A166 & \new_[45097]_ ;
  assign \new_[45099]_  = \new_[45098]_  & \new_[45093]_ ;
  assign \new_[45103]_  = A267 & A266;
  assign \new_[45104]_  = ~A265 & \new_[45103]_ ;
  assign \new_[45107]_  = A300 & A268;
  assign \new_[45110]_  = A302 & ~A301;
  assign \new_[45111]_  = \new_[45110]_  & \new_[45107]_ ;
  assign \new_[45112]_  = \new_[45111]_  & \new_[45104]_ ;
  assign \new_[45116]_  = ~A167 & A168;
  assign \new_[45117]_  = A170 & \new_[45116]_ ;
  assign \new_[45121]_  = A202 & ~A201;
  assign \new_[45122]_  = A166 & \new_[45121]_ ;
  assign \new_[45123]_  = \new_[45122]_  & \new_[45117]_ ;
  assign \new_[45127]_  = A267 & A266;
  assign \new_[45128]_  = ~A265 & \new_[45127]_ ;
  assign \new_[45131]_  = A300 & ~A269;
  assign \new_[45134]_  = A302 & ~A301;
  assign \new_[45135]_  = \new_[45134]_  & \new_[45131]_ ;
  assign \new_[45136]_  = \new_[45135]_  & \new_[45128]_ ;
  assign \new_[45140]_  = ~A167 & A168;
  assign \new_[45141]_  = A170 & \new_[45140]_ ;
  assign \new_[45145]_  = A202 & ~A201;
  assign \new_[45146]_  = A166 & \new_[45145]_ ;
  assign \new_[45147]_  = \new_[45146]_  & \new_[45141]_ ;
  assign \new_[45151]_  = ~A267 & A266;
  assign \new_[45152]_  = ~A265 & \new_[45151]_ ;
  assign \new_[45155]_  = A269 & ~A268;
  assign \new_[45158]_  = A301 & ~A300;
  assign \new_[45159]_  = \new_[45158]_  & \new_[45155]_ ;
  assign \new_[45160]_  = \new_[45159]_  & \new_[45152]_ ;
  assign \new_[45164]_  = ~A167 & A168;
  assign \new_[45165]_  = A170 & \new_[45164]_ ;
  assign \new_[45169]_  = A202 & ~A201;
  assign \new_[45170]_  = A166 & \new_[45169]_ ;
  assign \new_[45171]_  = \new_[45170]_  & \new_[45165]_ ;
  assign \new_[45175]_  = ~A267 & A266;
  assign \new_[45176]_  = ~A265 & \new_[45175]_ ;
  assign \new_[45179]_  = A269 & ~A268;
  assign \new_[45182]_  = ~A302 & ~A300;
  assign \new_[45183]_  = \new_[45182]_  & \new_[45179]_ ;
  assign \new_[45184]_  = \new_[45183]_  & \new_[45176]_ ;
  assign \new_[45188]_  = ~A167 & A168;
  assign \new_[45189]_  = A170 & \new_[45188]_ ;
  assign \new_[45193]_  = A202 & ~A201;
  assign \new_[45194]_  = A166 & \new_[45193]_ ;
  assign \new_[45195]_  = \new_[45194]_  & \new_[45189]_ ;
  assign \new_[45199]_  = ~A267 & A266;
  assign \new_[45200]_  = ~A265 & \new_[45199]_ ;
  assign \new_[45203]_  = A269 & ~A268;
  assign \new_[45206]_  = A299 & A298;
  assign \new_[45207]_  = \new_[45206]_  & \new_[45203]_ ;
  assign \new_[45208]_  = \new_[45207]_  & \new_[45200]_ ;
  assign \new_[45212]_  = ~A167 & A168;
  assign \new_[45213]_  = A170 & \new_[45212]_ ;
  assign \new_[45217]_  = A202 & ~A201;
  assign \new_[45218]_  = A166 & \new_[45217]_ ;
  assign \new_[45219]_  = \new_[45218]_  & \new_[45213]_ ;
  assign \new_[45223]_  = ~A267 & A266;
  assign \new_[45224]_  = ~A265 & \new_[45223]_ ;
  assign \new_[45227]_  = A269 & ~A268;
  assign \new_[45230]_  = ~A299 & ~A298;
  assign \new_[45231]_  = \new_[45230]_  & \new_[45227]_ ;
  assign \new_[45232]_  = \new_[45231]_  & \new_[45224]_ ;
  assign \new_[45236]_  = ~A167 & A168;
  assign \new_[45237]_  = A170 & \new_[45236]_ ;
  assign \new_[45241]_  = A202 & ~A201;
  assign \new_[45242]_  = A166 & \new_[45241]_ ;
  assign \new_[45243]_  = \new_[45242]_  & \new_[45237]_ ;
  assign \new_[45247]_  = A267 & ~A266;
  assign \new_[45248]_  = A265 & \new_[45247]_ ;
  assign \new_[45251]_  = A300 & A268;
  assign \new_[45254]_  = A302 & ~A301;
  assign \new_[45255]_  = \new_[45254]_  & \new_[45251]_ ;
  assign \new_[45256]_  = \new_[45255]_  & \new_[45248]_ ;
  assign \new_[45260]_  = ~A167 & A168;
  assign \new_[45261]_  = A170 & \new_[45260]_ ;
  assign \new_[45265]_  = A202 & ~A201;
  assign \new_[45266]_  = A166 & \new_[45265]_ ;
  assign \new_[45267]_  = \new_[45266]_  & \new_[45261]_ ;
  assign \new_[45271]_  = A267 & ~A266;
  assign \new_[45272]_  = A265 & \new_[45271]_ ;
  assign \new_[45275]_  = A300 & ~A269;
  assign \new_[45278]_  = A302 & ~A301;
  assign \new_[45279]_  = \new_[45278]_  & \new_[45275]_ ;
  assign \new_[45280]_  = \new_[45279]_  & \new_[45272]_ ;
  assign \new_[45284]_  = ~A167 & A168;
  assign \new_[45285]_  = A170 & \new_[45284]_ ;
  assign \new_[45289]_  = A202 & ~A201;
  assign \new_[45290]_  = A166 & \new_[45289]_ ;
  assign \new_[45291]_  = \new_[45290]_  & \new_[45285]_ ;
  assign \new_[45295]_  = ~A267 & ~A266;
  assign \new_[45296]_  = A265 & \new_[45295]_ ;
  assign \new_[45299]_  = A269 & ~A268;
  assign \new_[45302]_  = A301 & ~A300;
  assign \new_[45303]_  = \new_[45302]_  & \new_[45299]_ ;
  assign \new_[45304]_  = \new_[45303]_  & \new_[45296]_ ;
  assign \new_[45308]_  = ~A167 & A168;
  assign \new_[45309]_  = A170 & \new_[45308]_ ;
  assign \new_[45313]_  = A202 & ~A201;
  assign \new_[45314]_  = A166 & \new_[45313]_ ;
  assign \new_[45315]_  = \new_[45314]_  & \new_[45309]_ ;
  assign \new_[45319]_  = ~A267 & ~A266;
  assign \new_[45320]_  = A265 & \new_[45319]_ ;
  assign \new_[45323]_  = A269 & ~A268;
  assign \new_[45326]_  = ~A302 & ~A300;
  assign \new_[45327]_  = \new_[45326]_  & \new_[45323]_ ;
  assign \new_[45328]_  = \new_[45327]_  & \new_[45320]_ ;
  assign \new_[45332]_  = ~A167 & A168;
  assign \new_[45333]_  = A170 & \new_[45332]_ ;
  assign \new_[45337]_  = A202 & ~A201;
  assign \new_[45338]_  = A166 & \new_[45337]_ ;
  assign \new_[45339]_  = \new_[45338]_  & \new_[45333]_ ;
  assign \new_[45343]_  = ~A267 & ~A266;
  assign \new_[45344]_  = A265 & \new_[45343]_ ;
  assign \new_[45347]_  = A269 & ~A268;
  assign \new_[45350]_  = A299 & A298;
  assign \new_[45351]_  = \new_[45350]_  & \new_[45347]_ ;
  assign \new_[45352]_  = \new_[45351]_  & \new_[45344]_ ;
  assign \new_[45356]_  = ~A167 & A168;
  assign \new_[45357]_  = A170 & \new_[45356]_ ;
  assign \new_[45361]_  = A202 & ~A201;
  assign \new_[45362]_  = A166 & \new_[45361]_ ;
  assign \new_[45363]_  = \new_[45362]_  & \new_[45357]_ ;
  assign \new_[45367]_  = ~A267 & ~A266;
  assign \new_[45368]_  = A265 & \new_[45367]_ ;
  assign \new_[45371]_  = A269 & ~A268;
  assign \new_[45374]_  = ~A299 & ~A298;
  assign \new_[45375]_  = \new_[45374]_  & \new_[45371]_ ;
  assign \new_[45376]_  = \new_[45375]_  & \new_[45368]_ ;
  assign \new_[45380]_  = ~A167 & A168;
  assign \new_[45381]_  = A170 & \new_[45380]_ ;
  assign \new_[45385]_  = A202 & ~A201;
  assign \new_[45386]_  = A166 & \new_[45385]_ ;
  assign \new_[45387]_  = \new_[45386]_  & \new_[45381]_ ;
  assign \new_[45391]_  = A298 & ~A266;
  assign \new_[45392]_  = ~A265 & \new_[45391]_ ;
  assign \new_[45395]_  = ~A300 & ~A299;
  assign \new_[45398]_  = A302 & ~A301;
  assign \new_[45399]_  = \new_[45398]_  & \new_[45395]_ ;
  assign \new_[45400]_  = \new_[45399]_  & \new_[45392]_ ;
  assign \new_[45404]_  = ~A167 & A168;
  assign \new_[45405]_  = A170 & \new_[45404]_ ;
  assign \new_[45409]_  = A202 & ~A201;
  assign \new_[45410]_  = A166 & \new_[45409]_ ;
  assign \new_[45411]_  = \new_[45410]_  & \new_[45405]_ ;
  assign \new_[45415]_  = ~A298 & ~A266;
  assign \new_[45416]_  = ~A265 & \new_[45415]_ ;
  assign \new_[45419]_  = ~A300 & A299;
  assign \new_[45422]_  = A302 & ~A301;
  assign \new_[45423]_  = \new_[45422]_  & \new_[45419]_ ;
  assign \new_[45424]_  = \new_[45423]_  & \new_[45416]_ ;
  assign \new_[45428]_  = ~A167 & A168;
  assign \new_[45429]_  = A170 & \new_[45428]_ ;
  assign \new_[45433]_  = ~A203 & ~A201;
  assign \new_[45434]_  = A166 & \new_[45433]_ ;
  assign \new_[45435]_  = \new_[45434]_  & \new_[45429]_ ;
  assign \new_[45439]_  = A269 & ~A268;
  assign \new_[45440]_  = A267 & \new_[45439]_ ;
  assign \new_[45443]_  = ~A299 & A298;
  assign \new_[45446]_  = A301 & A300;
  assign \new_[45447]_  = \new_[45446]_  & \new_[45443]_ ;
  assign \new_[45448]_  = \new_[45447]_  & \new_[45440]_ ;
  assign \new_[45452]_  = ~A167 & A168;
  assign \new_[45453]_  = A170 & \new_[45452]_ ;
  assign \new_[45457]_  = ~A203 & ~A201;
  assign \new_[45458]_  = A166 & \new_[45457]_ ;
  assign \new_[45459]_  = \new_[45458]_  & \new_[45453]_ ;
  assign \new_[45463]_  = A269 & ~A268;
  assign \new_[45464]_  = A267 & \new_[45463]_ ;
  assign \new_[45467]_  = ~A299 & A298;
  assign \new_[45470]_  = ~A302 & A300;
  assign \new_[45471]_  = \new_[45470]_  & \new_[45467]_ ;
  assign \new_[45472]_  = \new_[45471]_  & \new_[45464]_ ;
  assign \new_[45476]_  = ~A167 & A168;
  assign \new_[45477]_  = A170 & \new_[45476]_ ;
  assign \new_[45481]_  = ~A203 & ~A201;
  assign \new_[45482]_  = A166 & \new_[45481]_ ;
  assign \new_[45483]_  = \new_[45482]_  & \new_[45477]_ ;
  assign \new_[45487]_  = A269 & ~A268;
  assign \new_[45488]_  = A267 & \new_[45487]_ ;
  assign \new_[45491]_  = A299 & ~A298;
  assign \new_[45494]_  = A301 & A300;
  assign \new_[45495]_  = \new_[45494]_  & \new_[45491]_ ;
  assign \new_[45496]_  = \new_[45495]_  & \new_[45488]_ ;
  assign \new_[45500]_  = ~A167 & A168;
  assign \new_[45501]_  = A170 & \new_[45500]_ ;
  assign \new_[45505]_  = ~A203 & ~A201;
  assign \new_[45506]_  = A166 & \new_[45505]_ ;
  assign \new_[45507]_  = \new_[45506]_  & \new_[45501]_ ;
  assign \new_[45511]_  = A269 & ~A268;
  assign \new_[45512]_  = A267 & \new_[45511]_ ;
  assign \new_[45515]_  = A299 & ~A298;
  assign \new_[45518]_  = ~A302 & A300;
  assign \new_[45519]_  = \new_[45518]_  & \new_[45515]_ ;
  assign \new_[45520]_  = \new_[45519]_  & \new_[45512]_ ;
  assign \new_[45524]_  = ~A167 & A168;
  assign \new_[45525]_  = A170 & \new_[45524]_ ;
  assign \new_[45529]_  = ~A203 & ~A201;
  assign \new_[45530]_  = A166 & \new_[45529]_ ;
  assign \new_[45531]_  = \new_[45530]_  & \new_[45525]_ ;
  assign \new_[45535]_  = A298 & A268;
  assign \new_[45536]_  = ~A267 & \new_[45535]_ ;
  assign \new_[45539]_  = ~A300 & ~A299;
  assign \new_[45542]_  = A302 & ~A301;
  assign \new_[45543]_  = \new_[45542]_  & \new_[45539]_ ;
  assign \new_[45544]_  = \new_[45543]_  & \new_[45536]_ ;
  assign \new_[45548]_  = ~A167 & A168;
  assign \new_[45549]_  = A170 & \new_[45548]_ ;
  assign \new_[45553]_  = ~A203 & ~A201;
  assign \new_[45554]_  = A166 & \new_[45553]_ ;
  assign \new_[45555]_  = \new_[45554]_  & \new_[45549]_ ;
  assign \new_[45559]_  = ~A298 & A268;
  assign \new_[45560]_  = ~A267 & \new_[45559]_ ;
  assign \new_[45563]_  = ~A300 & A299;
  assign \new_[45566]_  = A302 & ~A301;
  assign \new_[45567]_  = \new_[45566]_  & \new_[45563]_ ;
  assign \new_[45568]_  = \new_[45567]_  & \new_[45560]_ ;
  assign \new_[45572]_  = ~A167 & A168;
  assign \new_[45573]_  = A170 & \new_[45572]_ ;
  assign \new_[45577]_  = ~A203 & ~A201;
  assign \new_[45578]_  = A166 & \new_[45577]_ ;
  assign \new_[45579]_  = \new_[45578]_  & \new_[45573]_ ;
  assign \new_[45583]_  = A298 & ~A269;
  assign \new_[45584]_  = ~A267 & \new_[45583]_ ;
  assign \new_[45587]_  = ~A300 & ~A299;
  assign \new_[45590]_  = A302 & ~A301;
  assign \new_[45591]_  = \new_[45590]_  & \new_[45587]_ ;
  assign \new_[45592]_  = \new_[45591]_  & \new_[45584]_ ;
  assign \new_[45596]_  = ~A167 & A168;
  assign \new_[45597]_  = A170 & \new_[45596]_ ;
  assign \new_[45601]_  = ~A203 & ~A201;
  assign \new_[45602]_  = A166 & \new_[45601]_ ;
  assign \new_[45603]_  = \new_[45602]_  & \new_[45597]_ ;
  assign \new_[45607]_  = ~A298 & ~A269;
  assign \new_[45608]_  = ~A267 & \new_[45607]_ ;
  assign \new_[45611]_  = ~A300 & A299;
  assign \new_[45614]_  = A302 & ~A301;
  assign \new_[45615]_  = \new_[45614]_  & \new_[45611]_ ;
  assign \new_[45616]_  = \new_[45615]_  & \new_[45608]_ ;
  assign \new_[45620]_  = ~A167 & A168;
  assign \new_[45621]_  = A170 & \new_[45620]_ ;
  assign \new_[45625]_  = ~A203 & ~A201;
  assign \new_[45626]_  = A166 & \new_[45625]_ ;
  assign \new_[45627]_  = \new_[45626]_  & \new_[45621]_ ;
  assign \new_[45631]_  = A298 & A266;
  assign \new_[45632]_  = A265 & \new_[45631]_ ;
  assign \new_[45635]_  = ~A300 & ~A299;
  assign \new_[45638]_  = A302 & ~A301;
  assign \new_[45639]_  = \new_[45638]_  & \new_[45635]_ ;
  assign \new_[45640]_  = \new_[45639]_  & \new_[45632]_ ;
  assign \new_[45644]_  = ~A167 & A168;
  assign \new_[45645]_  = A170 & \new_[45644]_ ;
  assign \new_[45649]_  = ~A203 & ~A201;
  assign \new_[45650]_  = A166 & \new_[45649]_ ;
  assign \new_[45651]_  = \new_[45650]_  & \new_[45645]_ ;
  assign \new_[45655]_  = ~A298 & A266;
  assign \new_[45656]_  = A265 & \new_[45655]_ ;
  assign \new_[45659]_  = ~A300 & A299;
  assign \new_[45662]_  = A302 & ~A301;
  assign \new_[45663]_  = \new_[45662]_  & \new_[45659]_ ;
  assign \new_[45664]_  = \new_[45663]_  & \new_[45656]_ ;
  assign \new_[45668]_  = ~A167 & A168;
  assign \new_[45669]_  = A170 & \new_[45668]_ ;
  assign \new_[45673]_  = ~A203 & ~A201;
  assign \new_[45674]_  = A166 & \new_[45673]_ ;
  assign \new_[45675]_  = \new_[45674]_  & \new_[45669]_ ;
  assign \new_[45679]_  = A267 & A266;
  assign \new_[45680]_  = ~A265 & \new_[45679]_ ;
  assign \new_[45683]_  = A300 & A268;
  assign \new_[45686]_  = A302 & ~A301;
  assign \new_[45687]_  = \new_[45686]_  & \new_[45683]_ ;
  assign \new_[45688]_  = \new_[45687]_  & \new_[45680]_ ;
  assign \new_[45692]_  = ~A167 & A168;
  assign \new_[45693]_  = A170 & \new_[45692]_ ;
  assign \new_[45697]_  = ~A203 & ~A201;
  assign \new_[45698]_  = A166 & \new_[45697]_ ;
  assign \new_[45699]_  = \new_[45698]_  & \new_[45693]_ ;
  assign \new_[45703]_  = A267 & A266;
  assign \new_[45704]_  = ~A265 & \new_[45703]_ ;
  assign \new_[45707]_  = A300 & ~A269;
  assign \new_[45710]_  = A302 & ~A301;
  assign \new_[45711]_  = \new_[45710]_  & \new_[45707]_ ;
  assign \new_[45712]_  = \new_[45711]_  & \new_[45704]_ ;
  assign \new_[45716]_  = ~A167 & A168;
  assign \new_[45717]_  = A170 & \new_[45716]_ ;
  assign \new_[45721]_  = ~A203 & ~A201;
  assign \new_[45722]_  = A166 & \new_[45721]_ ;
  assign \new_[45723]_  = \new_[45722]_  & \new_[45717]_ ;
  assign \new_[45727]_  = ~A267 & A266;
  assign \new_[45728]_  = ~A265 & \new_[45727]_ ;
  assign \new_[45731]_  = A269 & ~A268;
  assign \new_[45734]_  = A301 & ~A300;
  assign \new_[45735]_  = \new_[45734]_  & \new_[45731]_ ;
  assign \new_[45736]_  = \new_[45735]_  & \new_[45728]_ ;
  assign \new_[45740]_  = ~A167 & A168;
  assign \new_[45741]_  = A170 & \new_[45740]_ ;
  assign \new_[45745]_  = ~A203 & ~A201;
  assign \new_[45746]_  = A166 & \new_[45745]_ ;
  assign \new_[45747]_  = \new_[45746]_  & \new_[45741]_ ;
  assign \new_[45751]_  = ~A267 & A266;
  assign \new_[45752]_  = ~A265 & \new_[45751]_ ;
  assign \new_[45755]_  = A269 & ~A268;
  assign \new_[45758]_  = ~A302 & ~A300;
  assign \new_[45759]_  = \new_[45758]_  & \new_[45755]_ ;
  assign \new_[45760]_  = \new_[45759]_  & \new_[45752]_ ;
  assign \new_[45764]_  = ~A167 & A168;
  assign \new_[45765]_  = A170 & \new_[45764]_ ;
  assign \new_[45769]_  = ~A203 & ~A201;
  assign \new_[45770]_  = A166 & \new_[45769]_ ;
  assign \new_[45771]_  = \new_[45770]_  & \new_[45765]_ ;
  assign \new_[45775]_  = ~A267 & A266;
  assign \new_[45776]_  = ~A265 & \new_[45775]_ ;
  assign \new_[45779]_  = A269 & ~A268;
  assign \new_[45782]_  = A299 & A298;
  assign \new_[45783]_  = \new_[45782]_  & \new_[45779]_ ;
  assign \new_[45784]_  = \new_[45783]_  & \new_[45776]_ ;
  assign \new_[45788]_  = ~A167 & A168;
  assign \new_[45789]_  = A170 & \new_[45788]_ ;
  assign \new_[45793]_  = ~A203 & ~A201;
  assign \new_[45794]_  = A166 & \new_[45793]_ ;
  assign \new_[45795]_  = \new_[45794]_  & \new_[45789]_ ;
  assign \new_[45799]_  = ~A267 & A266;
  assign \new_[45800]_  = ~A265 & \new_[45799]_ ;
  assign \new_[45803]_  = A269 & ~A268;
  assign \new_[45806]_  = ~A299 & ~A298;
  assign \new_[45807]_  = \new_[45806]_  & \new_[45803]_ ;
  assign \new_[45808]_  = \new_[45807]_  & \new_[45800]_ ;
  assign \new_[45812]_  = ~A167 & A168;
  assign \new_[45813]_  = A170 & \new_[45812]_ ;
  assign \new_[45817]_  = ~A203 & ~A201;
  assign \new_[45818]_  = A166 & \new_[45817]_ ;
  assign \new_[45819]_  = \new_[45818]_  & \new_[45813]_ ;
  assign \new_[45823]_  = A267 & ~A266;
  assign \new_[45824]_  = A265 & \new_[45823]_ ;
  assign \new_[45827]_  = A300 & A268;
  assign \new_[45830]_  = A302 & ~A301;
  assign \new_[45831]_  = \new_[45830]_  & \new_[45827]_ ;
  assign \new_[45832]_  = \new_[45831]_  & \new_[45824]_ ;
  assign \new_[45836]_  = ~A167 & A168;
  assign \new_[45837]_  = A170 & \new_[45836]_ ;
  assign \new_[45841]_  = ~A203 & ~A201;
  assign \new_[45842]_  = A166 & \new_[45841]_ ;
  assign \new_[45843]_  = \new_[45842]_  & \new_[45837]_ ;
  assign \new_[45847]_  = A267 & ~A266;
  assign \new_[45848]_  = A265 & \new_[45847]_ ;
  assign \new_[45851]_  = A300 & ~A269;
  assign \new_[45854]_  = A302 & ~A301;
  assign \new_[45855]_  = \new_[45854]_  & \new_[45851]_ ;
  assign \new_[45856]_  = \new_[45855]_  & \new_[45848]_ ;
  assign \new_[45860]_  = ~A167 & A168;
  assign \new_[45861]_  = A170 & \new_[45860]_ ;
  assign \new_[45865]_  = ~A203 & ~A201;
  assign \new_[45866]_  = A166 & \new_[45865]_ ;
  assign \new_[45867]_  = \new_[45866]_  & \new_[45861]_ ;
  assign \new_[45871]_  = ~A267 & ~A266;
  assign \new_[45872]_  = A265 & \new_[45871]_ ;
  assign \new_[45875]_  = A269 & ~A268;
  assign \new_[45878]_  = A301 & ~A300;
  assign \new_[45879]_  = \new_[45878]_  & \new_[45875]_ ;
  assign \new_[45880]_  = \new_[45879]_  & \new_[45872]_ ;
  assign \new_[45884]_  = ~A167 & A168;
  assign \new_[45885]_  = A170 & \new_[45884]_ ;
  assign \new_[45889]_  = ~A203 & ~A201;
  assign \new_[45890]_  = A166 & \new_[45889]_ ;
  assign \new_[45891]_  = \new_[45890]_  & \new_[45885]_ ;
  assign \new_[45895]_  = ~A267 & ~A266;
  assign \new_[45896]_  = A265 & \new_[45895]_ ;
  assign \new_[45899]_  = A269 & ~A268;
  assign \new_[45902]_  = ~A302 & ~A300;
  assign \new_[45903]_  = \new_[45902]_  & \new_[45899]_ ;
  assign \new_[45904]_  = \new_[45903]_  & \new_[45896]_ ;
  assign \new_[45908]_  = ~A167 & A168;
  assign \new_[45909]_  = A170 & \new_[45908]_ ;
  assign \new_[45913]_  = ~A203 & ~A201;
  assign \new_[45914]_  = A166 & \new_[45913]_ ;
  assign \new_[45915]_  = \new_[45914]_  & \new_[45909]_ ;
  assign \new_[45919]_  = ~A267 & ~A266;
  assign \new_[45920]_  = A265 & \new_[45919]_ ;
  assign \new_[45923]_  = A269 & ~A268;
  assign \new_[45926]_  = A299 & A298;
  assign \new_[45927]_  = \new_[45926]_  & \new_[45923]_ ;
  assign \new_[45928]_  = \new_[45927]_  & \new_[45920]_ ;
  assign \new_[45932]_  = ~A167 & A168;
  assign \new_[45933]_  = A170 & \new_[45932]_ ;
  assign \new_[45937]_  = ~A203 & ~A201;
  assign \new_[45938]_  = A166 & \new_[45937]_ ;
  assign \new_[45939]_  = \new_[45938]_  & \new_[45933]_ ;
  assign \new_[45943]_  = ~A267 & ~A266;
  assign \new_[45944]_  = A265 & \new_[45943]_ ;
  assign \new_[45947]_  = A269 & ~A268;
  assign \new_[45950]_  = ~A299 & ~A298;
  assign \new_[45951]_  = \new_[45950]_  & \new_[45947]_ ;
  assign \new_[45952]_  = \new_[45951]_  & \new_[45944]_ ;
  assign \new_[45956]_  = ~A167 & A168;
  assign \new_[45957]_  = A170 & \new_[45956]_ ;
  assign \new_[45961]_  = ~A203 & ~A201;
  assign \new_[45962]_  = A166 & \new_[45961]_ ;
  assign \new_[45963]_  = \new_[45962]_  & \new_[45957]_ ;
  assign \new_[45967]_  = A298 & ~A266;
  assign \new_[45968]_  = ~A265 & \new_[45967]_ ;
  assign \new_[45971]_  = ~A300 & ~A299;
  assign \new_[45974]_  = A302 & ~A301;
  assign \new_[45975]_  = \new_[45974]_  & \new_[45971]_ ;
  assign \new_[45976]_  = \new_[45975]_  & \new_[45968]_ ;
  assign \new_[45980]_  = ~A167 & A168;
  assign \new_[45981]_  = A170 & \new_[45980]_ ;
  assign \new_[45985]_  = ~A203 & ~A201;
  assign \new_[45986]_  = A166 & \new_[45985]_ ;
  assign \new_[45987]_  = \new_[45986]_  & \new_[45981]_ ;
  assign \new_[45991]_  = ~A298 & ~A266;
  assign \new_[45992]_  = ~A265 & \new_[45991]_ ;
  assign \new_[45995]_  = ~A300 & A299;
  assign \new_[45998]_  = A302 & ~A301;
  assign \new_[45999]_  = \new_[45998]_  & \new_[45995]_ ;
  assign \new_[46000]_  = \new_[45999]_  & \new_[45992]_ ;
  assign \new_[46004]_  = ~A167 & A168;
  assign \new_[46005]_  = A170 & \new_[46004]_ ;
  assign \new_[46009]_  = A200 & A199;
  assign \new_[46010]_  = A166 & \new_[46009]_ ;
  assign \new_[46011]_  = \new_[46010]_  & \new_[46005]_ ;
  assign \new_[46015]_  = A269 & ~A268;
  assign \new_[46016]_  = A267 & \new_[46015]_ ;
  assign \new_[46019]_  = ~A299 & A298;
  assign \new_[46022]_  = A301 & A300;
  assign \new_[46023]_  = \new_[46022]_  & \new_[46019]_ ;
  assign \new_[46024]_  = \new_[46023]_  & \new_[46016]_ ;
  assign \new_[46028]_  = ~A167 & A168;
  assign \new_[46029]_  = A170 & \new_[46028]_ ;
  assign \new_[46033]_  = A200 & A199;
  assign \new_[46034]_  = A166 & \new_[46033]_ ;
  assign \new_[46035]_  = \new_[46034]_  & \new_[46029]_ ;
  assign \new_[46039]_  = A269 & ~A268;
  assign \new_[46040]_  = A267 & \new_[46039]_ ;
  assign \new_[46043]_  = ~A299 & A298;
  assign \new_[46046]_  = ~A302 & A300;
  assign \new_[46047]_  = \new_[46046]_  & \new_[46043]_ ;
  assign \new_[46048]_  = \new_[46047]_  & \new_[46040]_ ;
  assign \new_[46052]_  = ~A167 & A168;
  assign \new_[46053]_  = A170 & \new_[46052]_ ;
  assign \new_[46057]_  = A200 & A199;
  assign \new_[46058]_  = A166 & \new_[46057]_ ;
  assign \new_[46059]_  = \new_[46058]_  & \new_[46053]_ ;
  assign \new_[46063]_  = A269 & ~A268;
  assign \new_[46064]_  = A267 & \new_[46063]_ ;
  assign \new_[46067]_  = A299 & ~A298;
  assign \new_[46070]_  = A301 & A300;
  assign \new_[46071]_  = \new_[46070]_  & \new_[46067]_ ;
  assign \new_[46072]_  = \new_[46071]_  & \new_[46064]_ ;
  assign \new_[46076]_  = ~A167 & A168;
  assign \new_[46077]_  = A170 & \new_[46076]_ ;
  assign \new_[46081]_  = A200 & A199;
  assign \new_[46082]_  = A166 & \new_[46081]_ ;
  assign \new_[46083]_  = \new_[46082]_  & \new_[46077]_ ;
  assign \new_[46087]_  = A269 & ~A268;
  assign \new_[46088]_  = A267 & \new_[46087]_ ;
  assign \new_[46091]_  = A299 & ~A298;
  assign \new_[46094]_  = ~A302 & A300;
  assign \new_[46095]_  = \new_[46094]_  & \new_[46091]_ ;
  assign \new_[46096]_  = \new_[46095]_  & \new_[46088]_ ;
  assign \new_[46100]_  = ~A167 & A168;
  assign \new_[46101]_  = A170 & \new_[46100]_ ;
  assign \new_[46105]_  = A200 & A199;
  assign \new_[46106]_  = A166 & \new_[46105]_ ;
  assign \new_[46107]_  = \new_[46106]_  & \new_[46101]_ ;
  assign \new_[46111]_  = A298 & A268;
  assign \new_[46112]_  = ~A267 & \new_[46111]_ ;
  assign \new_[46115]_  = ~A300 & ~A299;
  assign \new_[46118]_  = A302 & ~A301;
  assign \new_[46119]_  = \new_[46118]_  & \new_[46115]_ ;
  assign \new_[46120]_  = \new_[46119]_  & \new_[46112]_ ;
  assign \new_[46124]_  = ~A167 & A168;
  assign \new_[46125]_  = A170 & \new_[46124]_ ;
  assign \new_[46129]_  = A200 & A199;
  assign \new_[46130]_  = A166 & \new_[46129]_ ;
  assign \new_[46131]_  = \new_[46130]_  & \new_[46125]_ ;
  assign \new_[46135]_  = ~A298 & A268;
  assign \new_[46136]_  = ~A267 & \new_[46135]_ ;
  assign \new_[46139]_  = ~A300 & A299;
  assign \new_[46142]_  = A302 & ~A301;
  assign \new_[46143]_  = \new_[46142]_  & \new_[46139]_ ;
  assign \new_[46144]_  = \new_[46143]_  & \new_[46136]_ ;
  assign \new_[46148]_  = ~A167 & A168;
  assign \new_[46149]_  = A170 & \new_[46148]_ ;
  assign \new_[46153]_  = A200 & A199;
  assign \new_[46154]_  = A166 & \new_[46153]_ ;
  assign \new_[46155]_  = \new_[46154]_  & \new_[46149]_ ;
  assign \new_[46159]_  = A298 & ~A269;
  assign \new_[46160]_  = ~A267 & \new_[46159]_ ;
  assign \new_[46163]_  = ~A300 & ~A299;
  assign \new_[46166]_  = A302 & ~A301;
  assign \new_[46167]_  = \new_[46166]_  & \new_[46163]_ ;
  assign \new_[46168]_  = \new_[46167]_  & \new_[46160]_ ;
  assign \new_[46172]_  = ~A167 & A168;
  assign \new_[46173]_  = A170 & \new_[46172]_ ;
  assign \new_[46177]_  = A200 & A199;
  assign \new_[46178]_  = A166 & \new_[46177]_ ;
  assign \new_[46179]_  = \new_[46178]_  & \new_[46173]_ ;
  assign \new_[46183]_  = ~A298 & ~A269;
  assign \new_[46184]_  = ~A267 & \new_[46183]_ ;
  assign \new_[46187]_  = ~A300 & A299;
  assign \new_[46190]_  = A302 & ~A301;
  assign \new_[46191]_  = \new_[46190]_  & \new_[46187]_ ;
  assign \new_[46192]_  = \new_[46191]_  & \new_[46184]_ ;
  assign \new_[46196]_  = ~A167 & A168;
  assign \new_[46197]_  = A170 & \new_[46196]_ ;
  assign \new_[46201]_  = A200 & A199;
  assign \new_[46202]_  = A166 & \new_[46201]_ ;
  assign \new_[46203]_  = \new_[46202]_  & \new_[46197]_ ;
  assign \new_[46207]_  = A298 & A266;
  assign \new_[46208]_  = A265 & \new_[46207]_ ;
  assign \new_[46211]_  = ~A300 & ~A299;
  assign \new_[46214]_  = A302 & ~A301;
  assign \new_[46215]_  = \new_[46214]_  & \new_[46211]_ ;
  assign \new_[46216]_  = \new_[46215]_  & \new_[46208]_ ;
  assign \new_[46220]_  = ~A167 & A168;
  assign \new_[46221]_  = A170 & \new_[46220]_ ;
  assign \new_[46225]_  = A200 & A199;
  assign \new_[46226]_  = A166 & \new_[46225]_ ;
  assign \new_[46227]_  = \new_[46226]_  & \new_[46221]_ ;
  assign \new_[46231]_  = ~A298 & A266;
  assign \new_[46232]_  = A265 & \new_[46231]_ ;
  assign \new_[46235]_  = ~A300 & A299;
  assign \new_[46238]_  = A302 & ~A301;
  assign \new_[46239]_  = \new_[46238]_  & \new_[46235]_ ;
  assign \new_[46240]_  = \new_[46239]_  & \new_[46232]_ ;
  assign \new_[46244]_  = ~A167 & A168;
  assign \new_[46245]_  = A170 & \new_[46244]_ ;
  assign \new_[46249]_  = A200 & A199;
  assign \new_[46250]_  = A166 & \new_[46249]_ ;
  assign \new_[46251]_  = \new_[46250]_  & \new_[46245]_ ;
  assign \new_[46255]_  = A267 & A266;
  assign \new_[46256]_  = ~A265 & \new_[46255]_ ;
  assign \new_[46259]_  = A300 & A268;
  assign \new_[46262]_  = A302 & ~A301;
  assign \new_[46263]_  = \new_[46262]_  & \new_[46259]_ ;
  assign \new_[46264]_  = \new_[46263]_  & \new_[46256]_ ;
  assign \new_[46268]_  = ~A167 & A168;
  assign \new_[46269]_  = A170 & \new_[46268]_ ;
  assign \new_[46273]_  = A200 & A199;
  assign \new_[46274]_  = A166 & \new_[46273]_ ;
  assign \new_[46275]_  = \new_[46274]_  & \new_[46269]_ ;
  assign \new_[46279]_  = A267 & A266;
  assign \new_[46280]_  = ~A265 & \new_[46279]_ ;
  assign \new_[46283]_  = A300 & ~A269;
  assign \new_[46286]_  = A302 & ~A301;
  assign \new_[46287]_  = \new_[46286]_  & \new_[46283]_ ;
  assign \new_[46288]_  = \new_[46287]_  & \new_[46280]_ ;
  assign \new_[46292]_  = ~A167 & A168;
  assign \new_[46293]_  = A170 & \new_[46292]_ ;
  assign \new_[46297]_  = A200 & A199;
  assign \new_[46298]_  = A166 & \new_[46297]_ ;
  assign \new_[46299]_  = \new_[46298]_  & \new_[46293]_ ;
  assign \new_[46303]_  = ~A267 & A266;
  assign \new_[46304]_  = ~A265 & \new_[46303]_ ;
  assign \new_[46307]_  = A269 & ~A268;
  assign \new_[46310]_  = A301 & ~A300;
  assign \new_[46311]_  = \new_[46310]_  & \new_[46307]_ ;
  assign \new_[46312]_  = \new_[46311]_  & \new_[46304]_ ;
  assign \new_[46316]_  = ~A167 & A168;
  assign \new_[46317]_  = A170 & \new_[46316]_ ;
  assign \new_[46321]_  = A200 & A199;
  assign \new_[46322]_  = A166 & \new_[46321]_ ;
  assign \new_[46323]_  = \new_[46322]_  & \new_[46317]_ ;
  assign \new_[46327]_  = ~A267 & A266;
  assign \new_[46328]_  = ~A265 & \new_[46327]_ ;
  assign \new_[46331]_  = A269 & ~A268;
  assign \new_[46334]_  = ~A302 & ~A300;
  assign \new_[46335]_  = \new_[46334]_  & \new_[46331]_ ;
  assign \new_[46336]_  = \new_[46335]_  & \new_[46328]_ ;
  assign \new_[46340]_  = ~A167 & A168;
  assign \new_[46341]_  = A170 & \new_[46340]_ ;
  assign \new_[46345]_  = A200 & A199;
  assign \new_[46346]_  = A166 & \new_[46345]_ ;
  assign \new_[46347]_  = \new_[46346]_  & \new_[46341]_ ;
  assign \new_[46351]_  = ~A267 & A266;
  assign \new_[46352]_  = ~A265 & \new_[46351]_ ;
  assign \new_[46355]_  = A269 & ~A268;
  assign \new_[46358]_  = A299 & A298;
  assign \new_[46359]_  = \new_[46358]_  & \new_[46355]_ ;
  assign \new_[46360]_  = \new_[46359]_  & \new_[46352]_ ;
  assign \new_[46364]_  = ~A167 & A168;
  assign \new_[46365]_  = A170 & \new_[46364]_ ;
  assign \new_[46369]_  = A200 & A199;
  assign \new_[46370]_  = A166 & \new_[46369]_ ;
  assign \new_[46371]_  = \new_[46370]_  & \new_[46365]_ ;
  assign \new_[46375]_  = ~A267 & A266;
  assign \new_[46376]_  = ~A265 & \new_[46375]_ ;
  assign \new_[46379]_  = A269 & ~A268;
  assign \new_[46382]_  = ~A299 & ~A298;
  assign \new_[46383]_  = \new_[46382]_  & \new_[46379]_ ;
  assign \new_[46384]_  = \new_[46383]_  & \new_[46376]_ ;
  assign \new_[46388]_  = ~A167 & A168;
  assign \new_[46389]_  = A170 & \new_[46388]_ ;
  assign \new_[46393]_  = A200 & A199;
  assign \new_[46394]_  = A166 & \new_[46393]_ ;
  assign \new_[46395]_  = \new_[46394]_  & \new_[46389]_ ;
  assign \new_[46399]_  = A267 & ~A266;
  assign \new_[46400]_  = A265 & \new_[46399]_ ;
  assign \new_[46403]_  = A300 & A268;
  assign \new_[46406]_  = A302 & ~A301;
  assign \new_[46407]_  = \new_[46406]_  & \new_[46403]_ ;
  assign \new_[46408]_  = \new_[46407]_  & \new_[46400]_ ;
  assign \new_[46412]_  = ~A167 & A168;
  assign \new_[46413]_  = A170 & \new_[46412]_ ;
  assign \new_[46417]_  = A200 & A199;
  assign \new_[46418]_  = A166 & \new_[46417]_ ;
  assign \new_[46419]_  = \new_[46418]_  & \new_[46413]_ ;
  assign \new_[46423]_  = A267 & ~A266;
  assign \new_[46424]_  = A265 & \new_[46423]_ ;
  assign \new_[46427]_  = A300 & ~A269;
  assign \new_[46430]_  = A302 & ~A301;
  assign \new_[46431]_  = \new_[46430]_  & \new_[46427]_ ;
  assign \new_[46432]_  = \new_[46431]_  & \new_[46424]_ ;
  assign \new_[46436]_  = ~A167 & A168;
  assign \new_[46437]_  = A170 & \new_[46436]_ ;
  assign \new_[46441]_  = A200 & A199;
  assign \new_[46442]_  = A166 & \new_[46441]_ ;
  assign \new_[46443]_  = \new_[46442]_  & \new_[46437]_ ;
  assign \new_[46447]_  = ~A267 & ~A266;
  assign \new_[46448]_  = A265 & \new_[46447]_ ;
  assign \new_[46451]_  = A269 & ~A268;
  assign \new_[46454]_  = A301 & ~A300;
  assign \new_[46455]_  = \new_[46454]_  & \new_[46451]_ ;
  assign \new_[46456]_  = \new_[46455]_  & \new_[46448]_ ;
  assign \new_[46460]_  = ~A167 & A168;
  assign \new_[46461]_  = A170 & \new_[46460]_ ;
  assign \new_[46465]_  = A200 & A199;
  assign \new_[46466]_  = A166 & \new_[46465]_ ;
  assign \new_[46467]_  = \new_[46466]_  & \new_[46461]_ ;
  assign \new_[46471]_  = ~A267 & ~A266;
  assign \new_[46472]_  = A265 & \new_[46471]_ ;
  assign \new_[46475]_  = A269 & ~A268;
  assign \new_[46478]_  = ~A302 & ~A300;
  assign \new_[46479]_  = \new_[46478]_  & \new_[46475]_ ;
  assign \new_[46480]_  = \new_[46479]_  & \new_[46472]_ ;
  assign \new_[46484]_  = ~A167 & A168;
  assign \new_[46485]_  = A170 & \new_[46484]_ ;
  assign \new_[46489]_  = A200 & A199;
  assign \new_[46490]_  = A166 & \new_[46489]_ ;
  assign \new_[46491]_  = \new_[46490]_  & \new_[46485]_ ;
  assign \new_[46495]_  = ~A267 & ~A266;
  assign \new_[46496]_  = A265 & \new_[46495]_ ;
  assign \new_[46499]_  = A269 & ~A268;
  assign \new_[46502]_  = A299 & A298;
  assign \new_[46503]_  = \new_[46502]_  & \new_[46499]_ ;
  assign \new_[46504]_  = \new_[46503]_  & \new_[46496]_ ;
  assign \new_[46508]_  = ~A167 & A168;
  assign \new_[46509]_  = A170 & \new_[46508]_ ;
  assign \new_[46513]_  = A200 & A199;
  assign \new_[46514]_  = A166 & \new_[46513]_ ;
  assign \new_[46515]_  = \new_[46514]_  & \new_[46509]_ ;
  assign \new_[46519]_  = ~A267 & ~A266;
  assign \new_[46520]_  = A265 & \new_[46519]_ ;
  assign \new_[46523]_  = A269 & ~A268;
  assign \new_[46526]_  = ~A299 & ~A298;
  assign \new_[46527]_  = \new_[46526]_  & \new_[46523]_ ;
  assign \new_[46528]_  = \new_[46527]_  & \new_[46520]_ ;
  assign \new_[46532]_  = ~A167 & A168;
  assign \new_[46533]_  = A170 & \new_[46532]_ ;
  assign \new_[46537]_  = A200 & A199;
  assign \new_[46538]_  = A166 & \new_[46537]_ ;
  assign \new_[46539]_  = \new_[46538]_  & \new_[46533]_ ;
  assign \new_[46543]_  = A298 & ~A266;
  assign \new_[46544]_  = ~A265 & \new_[46543]_ ;
  assign \new_[46547]_  = ~A300 & ~A299;
  assign \new_[46550]_  = A302 & ~A301;
  assign \new_[46551]_  = \new_[46550]_  & \new_[46547]_ ;
  assign \new_[46552]_  = \new_[46551]_  & \new_[46544]_ ;
  assign \new_[46556]_  = ~A167 & A168;
  assign \new_[46557]_  = A170 & \new_[46556]_ ;
  assign \new_[46561]_  = A200 & A199;
  assign \new_[46562]_  = A166 & \new_[46561]_ ;
  assign \new_[46563]_  = \new_[46562]_  & \new_[46557]_ ;
  assign \new_[46567]_  = ~A298 & ~A266;
  assign \new_[46568]_  = ~A265 & \new_[46567]_ ;
  assign \new_[46571]_  = ~A300 & A299;
  assign \new_[46574]_  = A302 & ~A301;
  assign \new_[46575]_  = \new_[46574]_  & \new_[46571]_ ;
  assign \new_[46576]_  = \new_[46575]_  & \new_[46568]_ ;
  assign \new_[46580]_  = ~A167 & A168;
  assign \new_[46581]_  = A170 & \new_[46580]_ ;
  assign \new_[46585]_  = ~A200 & ~A199;
  assign \new_[46586]_  = A166 & \new_[46585]_ ;
  assign \new_[46587]_  = \new_[46586]_  & \new_[46581]_ ;
  assign \new_[46591]_  = A269 & ~A268;
  assign \new_[46592]_  = A267 & \new_[46591]_ ;
  assign \new_[46595]_  = ~A299 & A298;
  assign \new_[46598]_  = A301 & A300;
  assign \new_[46599]_  = \new_[46598]_  & \new_[46595]_ ;
  assign \new_[46600]_  = \new_[46599]_  & \new_[46592]_ ;
  assign \new_[46604]_  = ~A167 & A168;
  assign \new_[46605]_  = A170 & \new_[46604]_ ;
  assign \new_[46609]_  = ~A200 & ~A199;
  assign \new_[46610]_  = A166 & \new_[46609]_ ;
  assign \new_[46611]_  = \new_[46610]_  & \new_[46605]_ ;
  assign \new_[46615]_  = A269 & ~A268;
  assign \new_[46616]_  = A267 & \new_[46615]_ ;
  assign \new_[46619]_  = ~A299 & A298;
  assign \new_[46622]_  = ~A302 & A300;
  assign \new_[46623]_  = \new_[46622]_  & \new_[46619]_ ;
  assign \new_[46624]_  = \new_[46623]_  & \new_[46616]_ ;
  assign \new_[46628]_  = ~A167 & A168;
  assign \new_[46629]_  = A170 & \new_[46628]_ ;
  assign \new_[46633]_  = ~A200 & ~A199;
  assign \new_[46634]_  = A166 & \new_[46633]_ ;
  assign \new_[46635]_  = \new_[46634]_  & \new_[46629]_ ;
  assign \new_[46639]_  = A269 & ~A268;
  assign \new_[46640]_  = A267 & \new_[46639]_ ;
  assign \new_[46643]_  = A299 & ~A298;
  assign \new_[46646]_  = A301 & A300;
  assign \new_[46647]_  = \new_[46646]_  & \new_[46643]_ ;
  assign \new_[46648]_  = \new_[46647]_  & \new_[46640]_ ;
  assign \new_[46652]_  = ~A167 & A168;
  assign \new_[46653]_  = A170 & \new_[46652]_ ;
  assign \new_[46657]_  = ~A200 & ~A199;
  assign \new_[46658]_  = A166 & \new_[46657]_ ;
  assign \new_[46659]_  = \new_[46658]_  & \new_[46653]_ ;
  assign \new_[46663]_  = A269 & ~A268;
  assign \new_[46664]_  = A267 & \new_[46663]_ ;
  assign \new_[46667]_  = A299 & ~A298;
  assign \new_[46670]_  = ~A302 & A300;
  assign \new_[46671]_  = \new_[46670]_  & \new_[46667]_ ;
  assign \new_[46672]_  = \new_[46671]_  & \new_[46664]_ ;
  assign \new_[46676]_  = ~A167 & A168;
  assign \new_[46677]_  = A170 & \new_[46676]_ ;
  assign \new_[46681]_  = ~A200 & ~A199;
  assign \new_[46682]_  = A166 & \new_[46681]_ ;
  assign \new_[46683]_  = \new_[46682]_  & \new_[46677]_ ;
  assign \new_[46687]_  = A298 & A268;
  assign \new_[46688]_  = ~A267 & \new_[46687]_ ;
  assign \new_[46691]_  = ~A300 & ~A299;
  assign \new_[46694]_  = A302 & ~A301;
  assign \new_[46695]_  = \new_[46694]_  & \new_[46691]_ ;
  assign \new_[46696]_  = \new_[46695]_  & \new_[46688]_ ;
  assign \new_[46700]_  = ~A167 & A168;
  assign \new_[46701]_  = A170 & \new_[46700]_ ;
  assign \new_[46705]_  = ~A200 & ~A199;
  assign \new_[46706]_  = A166 & \new_[46705]_ ;
  assign \new_[46707]_  = \new_[46706]_  & \new_[46701]_ ;
  assign \new_[46711]_  = ~A298 & A268;
  assign \new_[46712]_  = ~A267 & \new_[46711]_ ;
  assign \new_[46715]_  = ~A300 & A299;
  assign \new_[46718]_  = A302 & ~A301;
  assign \new_[46719]_  = \new_[46718]_  & \new_[46715]_ ;
  assign \new_[46720]_  = \new_[46719]_  & \new_[46712]_ ;
  assign \new_[46724]_  = ~A167 & A168;
  assign \new_[46725]_  = A170 & \new_[46724]_ ;
  assign \new_[46729]_  = ~A200 & ~A199;
  assign \new_[46730]_  = A166 & \new_[46729]_ ;
  assign \new_[46731]_  = \new_[46730]_  & \new_[46725]_ ;
  assign \new_[46735]_  = A298 & ~A269;
  assign \new_[46736]_  = ~A267 & \new_[46735]_ ;
  assign \new_[46739]_  = ~A300 & ~A299;
  assign \new_[46742]_  = A302 & ~A301;
  assign \new_[46743]_  = \new_[46742]_  & \new_[46739]_ ;
  assign \new_[46744]_  = \new_[46743]_  & \new_[46736]_ ;
  assign \new_[46748]_  = ~A167 & A168;
  assign \new_[46749]_  = A170 & \new_[46748]_ ;
  assign \new_[46753]_  = ~A200 & ~A199;
  assign \new_[46754]_  = A166 & \new_[46753]_ ;
  assign \new_[46755]_  = \new_[46754]_  & \new_[46749]_ ;
  assign \new_[46759]_  = ~A298 & ~A269;
  assign \new_[46760]_  = ~A267 & \new_[46759]_ ;
  assign \new_[46763]_  = ~A300 & A299;
  assign \new_[46766]_  = A302 & ~A301;
  assign \new_[46767]_  = \new_[46766]_  & \new_[46763]_ ;
  assign \new_[46768]_  = \new_[46767]_  & \new_[46760]_ ;
  assign \new_[46772]_  = ~A167 & A168;
  assign \new_[46773]_  = A170 & \new_[46772]_ ;
  assign \new_[46777]_  = ~A200 & ~A199;
  assign \new_[46778]_  = A166 & \new_[46777]_ ;
  assign \new_[46779]_  = \new_[46778]_  & \new_[46773]_ ;
  assign \new_[46783]_  = A298 & A266;
  assign \new_[46784]_  = A265 & \new_[46783]_ ;
  assign \new_[46787]_  = ~A300 & ~A299;
  assign \new_[46790]_  = A302 & ~A301;
  assign \new_[46791]_  = \new_[46790]_  & \new_[46787]_ ;
  assign \new_[46792]_  = \new_[46791]_  & \new_[46784]_ ;
  assign \new_[46796]_  = ~A167 & A168;
  assign \new_[46797]_  = A170 & \new_[46796]_ ;
  assign \new_[46801]_  = ~A200 & ~A199;
  assign \new_[46802]_  = A166 & \new_[46801]_ ;
  assign \new_[46803]_  = \new_[46802]_  & \new_[46797]_ ;
  assign \new_[46807]_  = ~A298 & A266;
  assign \new_[46808]_  = A265 & \new_[46807]_ ;
  assign \new_[46811]_  = ~A300 & A299;
  assign \new_[46814]_  = A302 & ~A301;
  assign \new_[46815]_  = \new_[46814]_  & \new_[46811]_ ;
  assign \new_[46816]_  = \new_[46815]_  & \new_[46808]_ ;
  assign \new_[46820]_  = ~A167 & A168;
  assign \new_[46821]_  = A170 & \new_[46820]_ ;
  assign \new_[46825]_  = ~A200 & ~A199;
  assign \new_[46826]_  = A166 & \new_[46825]_ ;
  assign \new_[46827]_  = \new_[46826]_  & \new_[46821]_ ;
  assign \new_[46831]_  = A267 & A266;
  assign \new_[46832]_  = ~A265 & \new_[46831]_ ;
  assign \new_[46835]_  = A300 & A268;
  assign \new_[46838]_  = A302 & ~A301;
  assign \new_[46839]_  = \new_[46838]_  & \new_[46835]_ ;
  assign \new_[46840]_  = \new_[46839]_  & \new_[46832]_ ;
  assign \new_[46844]_  = ~A167 & A168;
  assign \new_[46845]_  = A170 & \new_[46844]_ ;
  assign \new_[46849]_  = ~A200 & ~A199;
  assign \new_[46850]_  = A166 & \new_[46849]_ ;
  assign \new_[46851]_  = \new_[46850]_  & \new_[46845]_ ;
  assign \new_[46855]_  = A267 & A266;
  assign \new_[46856]_  = ~A265 & \new_[46855]_ ;
  assign \new_[46859]_  = A300 & ~A269;
  assign \new_[46862]_  = A302 & ~A301;
  assign \new_[46863]_  = \new_[46862]_  & \new_[46859]_ ;
  assign \new_[46864]_  = \new_[46863]_  & \new_[46856]_ ;
  assign \new_[46868]_  = ~A167 & A168;
  assign \new_[46869]_  = A170 & \new_[46868]_ ;
  assign \new_[46873]_  = ~A200 & ~A199;
  assign \new_[46874]_  = A166 & \new_[46873]_ ;
  assign \new_[46875]_  = \new_[46874]_  & \new_[46869]_ ;
  assign \new_[46879]_  = ~A267 & A266;
  assign \new_[46880]_  = ~A265 & \new_[46879]_ ;
  assign \new_[46883]_  = A269 & ~A268;
  assign \new_[46886]_  = A301 & ~A300;
  assign \new_[46887]_  = \new_[46886]_  & \new_[46883]_ ;
  assign \new_[46888]_  = \new_[46887]_  & \new_[46880]_ ;
  assign \new_[46892]_  = ~A167 & A168;
  assign \new_[46893]_  = A170 & \new_[46892]_ ;
  assign \new_[46897]_  = ~A200 & ~A199;
  assign \new_[46898]_  = A166 & \new_[46897]_ ;
  assign \new_[46899]_  = \new_[46898]_  & \new_[46893]_ ;
  assign \new_[46903]_  = ~A267 & A266;
  assign \new_[46904]_  = ~A265 & \new_[46903]_ ;
  assign \new_[46907]_  = A269 & ~A268;
  assign \new_[46910]_  = ~A302 & ~A300;
  assign \new_[46911]_  = \new_[46910]_  & \new_[46907]_ ;
  assign \new_[46912]_  = \new_[46911]_  & \new_[46904]_ ;
  assign \new_[46916]_  = ~A167 & A168;
  assign \new_[46917]_  = A170 & \new_[46916]_ ;
  assign \new_[46921]_  = ~A200 & ~A199;
  assign \new_[46922]_  = A166 & \new_[46921]_ ;
  assign \new_[46923]_  = \new_[46922]_  & \new_[46917]_ ;
  assign \new_[46927]_  = ~A267 & A266;
  assign \new_[46928]_  = ~A265 & \new_[46927]_ ;
  assign \new_[46931]_  = A269 & ~A268;
  assign \new_[46934]_  = A299 & A298;
  assign \new_[46935]_  = \new_[46934]_  & \new_[46931]_ ;
  assign \new_[46936]_  = \new_[46935]_  & \new_[46928]_ ;
  assign \new_[46940]_  = ~A167 & A168;
  assign \new_[46941]_  = A170 & \new_[46940]_ ;
  assign \new_[46945]_  = ~A200 & ~A199;
  assign \new_[46946]_  = A166 & \new_[46945]_ ;
  assign \new_[46947]_  = \new_[46946]_  & \new_[46941]_ ;
  assign \new_[46951]_  = ~A267 & A266;
  assign \new_[46952]_  = ~A265 & \new_[46951]_ ;
  assign \new_[46955]_  = A269 & ~A268;
  assign \new_[46958]_  = ~A299 & ~A298;
  assign \new_[46959]_  = \new_[46958]_  & \new_[46955]_ ;
  assign \new_[46960]_  = \new_[46959]_  & \new_[46952]_ ;
  assign \new_[46964]_  = ~A167 & A168;
  assign \new_[46965]_  = A170 & \new_[46964]_ ;
  assign \new_[46969]_  = ~A200 & ~A199;
  assign \new_[46970]_  = A166 & \new_[46969]_ ;
  assign \new_[46971]_  = \new_[46970]_  & \new_[46965]_ ;
  assign \new_[46975]_  = A267 & ~A266;
  assign \new_[46976]_  = A265 & \new_[46975]_ ;
  assign \new_[46979]_  = A300 & A268;
  assign \new_[46982]_  = A302 & ~A301;
  assign \new_[46983]_  = \new_[46982]_  & \new_[46979]_ ;
  assign \new_[46984]_  = \new_[46983]_  & \new_[46976]_ ;
  assign \new_[46988]_  = ~A167 & A168;
  assign \new_[46989]_  = A170 & \new_[46988]_ ;
  assign \new_[46993]_  = ~A200 & ~A199;
  assign \new_[46994]_  = A166 & \new_[46993]_ ;
  assign \new_[46995]_  = \new_[46994]_  & \new_[46989]_ ;
  assign \new_[46999]_  = A267 & ~A266;
  assign \new_[47000]_  = A265 & \new_[46999]_ ;
  assign \new_[47003]_  = A300 & ~A269;
  assign \new_[47006]_  = A302 & ~A301;
  assign \new_[47007]_  = \new_[47006]_  & \new_[47003]_ ;
  assign \new_[47008]_  = \new_[47007]_  & \new_[47000]_ ;
  assign \new_[47012]_  = ~A167 & A168;
  assign \new_[47013]_  = A170 & \new_[47012]_ ;
  assign \new_[47017]_  = ~A200 & ~A199;
  assign \new_[47018]_  = A166 & \new_[47017]_ ;
  assign \new_[47019]_  = \new_[47018]_  & \new_[47013]_ ;
  assign \new_[47023]_  = ~A267 & ~A266;
  assign \new_[47024]_  = A265 & \new_[47023]_ ;
  assign \new_[47027]_  = A269 & ~A268;
  assign \new_[47030]_  = A301 & ~A300;
  assign \new_[47031]_  = \new_[47030]_  & \new_[47027]_ ;
  assign \new_[47032]_  = \new_[47031]_  & \new_[47024]_ ;
  assign \new_[47036]_  = ~A167 & A168;
  assign \new_[47037]_  = A170 & \new_[47036]_ ;
  assign \new_[47041]_  = ~A200 & ~A199;
  assign \new_[47042]_  = A166 & \new_[47041]_ ;
  assign \new_[47043]_  = \new_[47042]_  & \new_[47037]_ ;
  assign \new_[47047]_  = ~A267 & ~A266;
  assign \new_[47048]_  = A265 & \new_[47047]_ ;
  assign \new_[47051]_  = A269 & ~A268;
  assign \new_[47054]_  = ~A302 & ~A300;
  assign \new_[47055]_  = \new_[47054]_  & \new_[47051]_ ;
  assign \new_[47056]_  = \new_[47055]_  & \new_[47048]_ ;
  assign \new_[47060]_  = ~A167 & A168;
  assign \new_[47061]_  = A170 & \new_[47060]_ ;
  assign \new_[47065]_  = ~A200 & ~A199;
  assign \new_[47066]_  = A166 & \new_[47065]_ ;
  assign \new_[47067]_  = \new_[47066]_  & \new_[47061]_ ;
  assign \new_[47071]_  = ~A267 & ~A266;
  assign \new_[47072]_  = A265 & \new_[47071]_ ;
  assign \new_[47075]_  = A269 & ~A268;
  assign \new_[47078]_  = A299 & A298;
  assign \new_[47079]_  = \new_[47078]_  & \new_[47075]_ ;
  assign \new_[47080]_  = \new_[47079]_  & \new_[47072]_ ;
  assign \new_[47084]_  = ~A167 & A168;
  assign \new_[47085]_  = A170 & \new_[47084]_ ;
  assign \new_[47089]_  = ~A200 & ~A199;
  assign \new_[47090]_  = A166 & \new_[47089]_ ;
  assign \new_[47091]_  = \new_[47090]_  & \new_[47085]_ ;
  assign \new_[47095]_  = ~A267 & ~A266;
  assign \new_[47096]_  = A265 & \new_[47095]_ ;
  assign \new_[47099]_  = A269 & ~A268;
  assign \new_[47102]_  = ~A299 & ~A298;
  assign \new_[47103]_  = \new_[47102]_  & \new_[47099]_ ;
  assign \new_[47104]_  = \new_[47103]_  & \new_[47096]_ ;
  assign \new_[47108]_  = ~A167 & A168;
  assign \new_[47109]_  = A170 & \new_[47108]_ ;
  assign \new_[47113]_  = ~A200 & ~A199;
  assign \new_[47114]_  = A166 & \new_[47113]_ ;
  assign \new_[47115]_  = \new_[47114]_  & \new_[47109]_ ;
  assign \new_[47119]_  = A298 & ~A266;
  assign \new_[47120]_  = ~A265 & \new_[47119]_ ;
  assign \new_[47123]_  = ~A300 & ~A299;
  assign \new_[47126]_  = A302 & ~A301;
  assign \new_[47127]_  = \new_[47126]_  & \new_[47123]_ ;
  assign \new_[47128]_  = \new_[47127]_  & \new_[47120]_ ;
  assign \new_[47132]_  = ~A167 & A168;
  assign \new_[47133]_  = A170 & \new_[47132]_ ;
  assign \new_[47137]_  = ~A200 & ~A199;
  assign \new_[47138]_  = A166 & \new_[47137]_ ;
  assign \new_[47139]_  = \new_[47138]_  & \new_[47133]_ ;
  assign \new_[47143]_  = ~A298 & ~A266;
  assign \new_[47144]_  = ~A265 & \new_[47143]_ ;
  assign \new_[47147]_  = ~A300 & A299;
  assign \new_[47150]_  = A302 & ~A301;
  assign \new_[47151]_  = \new_[47150]_  & \new_[47147]_ ;
  assign \new_[47152]_  = \new_[47151]_  & \new_[47144]_ ;
  assign \new_[47156]_  = ~A199 & ~A168;
  assign \new_[47157]_  = A170 & \new_[47156]_ ;
  assign \new_[47161]_  = ~A202 & ~A201;
  assign \new_[47162]_  = A200 & \new_[47161]_ ;
  assign \new_[47163]_  = \new_[47162]_  & \new_[47157]_ ;
  assign \new_[47167]_  = ~A268 & A267;
  assign \new_[47168]_  = A203 & \new_[47167]_ ;
  assign \new_[47171]_  = A300 & A269;
  assign \new_[47174]_  = A302 & ~A301;
  assign \new_[47175]_  = \new_[47174]_  & \new_[47171]_ ;
  assign \new_[47176]_  = \new_[47175]_  & \new_[47168]_ ;
  assign \new_[47180]_  = A199 & ~A168;
  assign \new_[47181]_  = A170 & \new_[47180]_ ;
  assign \new_[47185]_  = ~A202 & ~A201;
  assign \new_[47186]_  = ~A200 & \new_[47185]_ ;
  assign \new_[47187]_  = \new_[47186]_  & \new_[47181]_ ;
  assign \new_[47191]_  = ~A268 & A267;
  assign \new_[47192]_  = A203 & \new_[47191]_ ;
  assign \new_[47195]_  = A300 & A269;
  assign \new_[47198]_  = A302 & ~A301;
  assign \new_[47199]_  = \new_[47198]_  & \new_[47195]_ ;
  assign \new_[47200]_  = \new_[47199]_  & \new_[47192]_ ;
  assign \new_[47204]_  = A167 & A168;
  assign \new_[47205]_  = A169 & \new_[47204]_ ;
  assign \new_[47209]_  = ~A202 & A201;
  assign \new_[47210]_  = ~A166 & \new_[47209]_ ;
  assign \new_[47211]_  = \new_[47210]_  & \new_[47205]_ ;
  assign \new_[47215]_  = A268 & ~A267;
  assign \new_[47216]_  = A203 & \new_[47215]_ ;
  assign \new_[47219]_  = ~A299 & A298;
  assign \new_[47222]_  = A301 & A300;
  assign \new_[47223]_  = \new_[47222]_  & \new_[47219]_ ;
  assign \new_[47224]_  = \new_[47223]_  & \new_[47216]_ ;
  assign \new_[47228]_  = A167 & A168;
  assign \new_[47229]_  = A169 & \new_[47228]_ ;
  assign \new_[47233]_  = ~A202 & A201;
  assign \new_[47234]_  = ~A166 & \new_[47233]_ ;
  assign \new_[47235]_  = \new_[47234]_  & \new_[47229]_ ;
  assign \new_[47239]_  = A268 & ~A267;
  assign \new_[47240]_  = A203 & \new_[47239]_ ;
  assign \new_[47243]_  = ~A299 & A298;
  assign \new_[47246]_  = ~A302 & A300;
  assign \new_[47247]_  = \new_[47246]_  & \new_[47243]_ ;
  assign \new_[47248]_  = \new_[47247]_  & \new_[47240]_ ;
  assign \new_[47252]_  = A167 & A168;
  assign \new_[47253]_  = A169 & \new_[47252]_ ;
  assign \new_[47257]_  = ~A202 & A201;
  assign \new_[47258]_  = ~A166 & \new_[47257]_ ;
  assign \new_[47259]_  = \new_[47258]_  & \new_[47253]_ ;
  assign \new_[47263]_  = A268 & ~A267;
  assign \new_[47264]_  = A203 & \new_[47263]_ ;
  assign \new_[47267]_  = A299 & ~A298;
  assign \new_[47270]_  = A301 & A300;
  assign \new_[47271]_  = \new_[47270]_  & \new_[47267]_ ;
  assign \new_[47272]_  = \new_[47271]_  & \new_[47264]_ ;
  assign \new_[47276]_  = A167 & A168;
  assign \new_[47277]_  = A169 & \new_[47276]_ ;
  assign \new_[47281]_  = ~A202 & A201;
  assign \new_[47282]_  = ~A166 & \new_[47281]_ ;
  assign \new_[47283]_  = \new_[47282]_  & \new_[47277]_ ;
  assign \new_[47287]_  = A268 & ~A267;
  assign \new_[47288]_  = A203 & \new_[47287]_ ;
  assign \new_[47291]_  = A299 & ~A298;
  assign \new_[47294]_  = ~A302 & A300;
  assign \new_[47295]_  = \new_[47294]_  & \new_[47291]_ ;
  assign \new_[47296]_  = \new_[47295]_  & \new_[47288]_ ;
  assign \new_[47300]_  = A167 & A168;
  assign \new_[47301]_  = A169 & \new_[47300]_ ;
  assign \new_[47305]_  = ~A202 & A201;
  assign \new_[47306]_  = ~A166 & \new_[47305]_ ;
  assign \new_[47307]_  = \new_[47306]_  & \new_[47301]_ ;
  assign \new_[47311]_  = ~A269 & ~A267;
  assign \new_[47312]_  = A203 & \new_[47311]_ ;
  assign \new_[47315]_  = ~A299 & A298;
  assign \new_[47318]_  = A301 & A300;
  assign \new_[47319]_  = \new_[47318]_  & \new_[47315]_ ;
  assign \new_[47320]_  = \new_[47319]_  & \new_[47312]_ ;
  assign \new_[47324]_  = A167 & A168;
  assign \new_[47325]_  = A169 & \new_[47324]_ ;
  assign \new_[47329]_  = ~A202 & A201;
  assign \new_[47330]_  = ~A166 & \new_[47329]_ ;
  assign \new_[47331]_  = \new_[47330]_  & \new_[47325]_ ;
  assign \new_[47335]_  = ~A269 & ~A267;
  assign \new_[47336]_  = A203 & \new_[47335]_ ;
  assign \new_[47339]_  = ~A299 & A298;
  assign \new_[47342]_  = ~A302 & A300;
  assign \new_[47343]_  = \new_[47342]_  & \new_[47339]_ ;
  assign \new_[47344]_  = \new_[47343]_  & \new_[47336]_ ;
  assign \new_[47348]_  = A167 & A168;
  assign \new_[47349]_  = A169 & \new_[47348]_ ;
  assign \new_[47353]_  = ~A202 & A201;
  assign \new_[47354]_  = ~A166 & \new_[47353]_ ;
  assign \new_[47355]_  = \new_[47354]_  & \new_[47349]_ ;
  assign \new_[47359]_  = ~A269 & ~A267;
  assign \new_[47360]_  = A203 & \new_[47359]_ ;
  assign \new_[47363]_  = A299 & ~A298;
  assign \new_[47366]_  = A301 & A300;
  assign \new_[47367]_  = \new_[47366]_  & \new_[47363]_ ;
  assign \new_[47368]_  = \new_[47367]_  & \new_[47360]_ ;
  assign \new_[47372]_  = A167 & A168;
  assign \new_[47373]_  = A169 & \new_[47372]_ ;
  assign \new_[47377]_  = ~A202 & A201;
  assign \new_[47378]_  = ~A166 & \new_[47377]_ ;
  assign \new_[47379]_  = \new_[47378]_  & \new_[47373]_ ;
  assign \new_[47383]_  = ~A269 & ~A267;
  assign \new_[47384]_  = A203 & \new_[47383]_ ;
  assign \new_[47387]_  = A299 & ~A298;
  assign \new_[47390]_  = ~A302 & A300;
  assign \new_[47391]_  = \new_[47390]_  & \new_[47387]_ ;
  assign \new_[47392]_  = \new_[47391]_  & \new_[47384]_ ;
  assign \new_[47396]_  = A167 & A168;
  assign \new_[47397]_  = A169 & \new_[47396]_ ;
  assign \new_[47401]_  = ~A202 & A201;
  assign \new_[47402]_  = ~A166 & \new_[47401]_ ;
  assign \new_[47403]_  = \new_[47402]_  & \new_[47397]_ ;
  assign \new_[47407]_  = A266 & A265;
  assign \new_[47408]_  = A203 & \new_[47407]_ ;
  assign \new_[47411]_  = ~A299 & A298;
  assign \new_[47414]_  = A301 & A300;
  assign \new_[47415]_  = \new_[47414]_  & \new_[47411]_ ;
  assign \new_[47416]_  = \new_[47415]_  & \new_[47408]_ ;
  assign \new_[47420]_  = A167 & A168;
  assign \new_[47421]_  = A169 & \new_[47420]_ ;
  assign \new_[47425]_  = ~A202 & A201;
  assign \new_[47426]_  = ~A166 & \new_[47425]_ ;
  assign \new_[47427]_  = \new_[47426]_  & \new_[47421]_ ;
  assign \new_[47431]_  = A266 & A265;
  assign \new_[47432]_  = A203 & \new_[47431]_ ;
  assign \new_[47435]_  = ~A299 & A298;
  assign \new_[47438]_  = ~A302 & A300;
  assign \new_[47439]_  = \new_[47438]_  & \new_[47435]_ ;
  assign \new_[47440]_  = \new_[47439]_  & \new_[47432]_ ;
  assign \new_[47444]_  = A167 & A168;
  assign \new_[47445]_  = A169 & \new_[47444]_ ;
  assign \new_[47449]_  = ~A202 & A201;
  assign \new_[47450]_  = ~A166 & \new_[47449]_ ;
  assign \new_[47451]_  = \new_[47450]_  & \new_[47445]_ ;
  assign \new_[47455]_  = A266 & A265;
  assign \new_[47456]_  = A203 & \new_[47455]_ ;
  assign \new_[47459]_  = A299 & ~A298;
  assign \new_[47462]_  = A301 & A300;
  assign \new_[47463]_  = \new_[47462]_  & \new_[47459]_ ;
  assign \new_[47464]_  = \new_[47463]_  & \new_[47456]_ ;
  assign \new_[47468]_  = A167 & A168;
  assign \new_[47469]_  = A169 & \new_[47468]_ ;
  assign \new_[47473]_  = ~A202 & A201;
  assign \new_[47474]_  = ~A166 & \new_[47473]_ ;
  assign \new_[47475]_  = \new_[47474]_  & \new_[47469]_ ;
  assign \new_[47479]_  = A266 & A265;
  assign \new_[47480]_  = A203 & \new_[47479]_ ;
  assign \new_[47483]_  = A299 & ~A298;
  assign \new_[47486]_  = ~A302 & A300;
  assign \new_[47487]_  = \new_[47486]_  & \new_[47483]_ ;
  assign \new_[47488]_  = \new_[47487]_  & \new_[47480]_ ;
  assign \new_[47492]_  = A167 & A168;
  assign \new_[47493]_  = A169 & \new_[47492]_ ;
  assign \new_[47497]_  = ~A202 & A201;
  assign \new_[47498]_  = ~A166 & \new_[47497]_ ;
  assign \new_[47499]_  = \new_[47498]_  & \new_[47493]_ ;
  assign \new_[47503]_  = A266 & ~A265;
  assign \new_[47504]_  = A203 & \new_[47503]_ ;
  assign \new_[47507]_  = A268 & A267;
  assign \new_[47510]_  = A301 & ~A300;
  assign \new_[47511]_  = \new_[47510]_  & \new_[47507]_ ;
  assign \new_[47512]_  = \new_[47511]_  & \new_[47504]_ ;
  assign \new_[47516]_  = A167 & A168;
  assign \new_[47517]_  = A169 & \new_[47516]_ ;
  assign \new_[47521]_  = ~A202 & A201;
  assign \new_[47522]_  = ~A166 & \new_[47521]_ ;
  assign \new_[47523]_  = \new_[47522]_  & \new_[47517]_ ;
  assign \new_[47527]_  = A266 & ~A265;
  assign \new_[47528]_  = A203 & \new_[47527]_ ;
  assign \new_[47531]_  = A268 & A267;
  assign \new_[47534]_  = ~A302 & ~A300;
  assign \new_[47535]_  = \new_[47534]_  & \new_[47531]_ ;
  assign \new_[47536]_  = \new_[47535]_  & \new_[47528]_ ;
  assign \new_[47540]_  = A167 & A168;
  assign \new_[47541]_  = A169 & \new_[47540]_ ;
  assign \new_[47545]_  = ~A202 & A201;
  assign \new_[47546]_  = ~A166 & \new_[47545]_ ;
  assign \new_[47547]_  = \new_[47546]_  & \new_[47541]_ ;
  assign \new_[47551]_  = A266 & ~A265;
  assign \new_[47552]_  = A203 & \new_[47551]_ ;
  assign \new_[47555]_  = A268 & A267;
  assign \new_[47558]_  = A299 & A298;
  assign \new_[47559]_  = \new_[47558]_  & \new_[47555]_ ;
  assign \new_[47560]_  = \new_[47559]_  & \new_[47552]_ ;
  assign \new_[47564]_  = A167 & A168;
  assign \new_[47565]_  = A169 & \new_[47564]_ ;
  assign \new_[47569]_  = ~A202 & A201;
  assign \new_[47570]_  = ~A166 & \new_[47569]_ ;
  assign \new_[47571]_  = \new_[47570]_  & \new_[47565]_ ;
  assign \new_[47575]_  = A266 & ~A265;
  assign \new_[47576]_  = A203 & \new_[47575]_ ;
  assign \new_[47579]_  = A268 & A267;
  assign \new_[47582]_  = ~A299 & ~A298;
  assign \new_[47583]_  = \new_[47582]_  & \new_[47579]_ ;
  assign \new_[47584]_  = \new_[47583]_  & \new_[47576]_ ;
  assign \new_[47588]_  = A167 & A168;
  assign \new_[47589]_  = A169 & \new_[47588]_ ;
  assign \new_[47593]_  = ~A202 & A201;
  assign \new_[47594]_  = ~A166 & \new_[47593]_ ;
  assign \new_[47595]_  = \new_[47594]_  & \new_[47589]_ ;
  assign \new_[47599]_  = A266 & ~A265;
  assign \new_[47600]_  = A203 & \new_[47599]_ ;
  assign \new_[47603]_  = ~A269 & A267;
  assign \new_[47606]_  = A301 & ~A300;
  assign \new_[47607]_  = \new_[47606]_  & \new_[47603]_ ;
  assign \new_[47608]_  = \new_[47607]_  & \new_[47600]_ ;
  assign \new_[47612]_  = A167 & A168;
  assign \new_[47613]_  = A169 & \new_[47612]_ ;
  assign \new_[47617]_  = ~A202 & A201;
  assign \new_[47618]_  = ~A166 & \new_[47617]_ ;
  assign \new_[47619]_  = \new_[47618]_  & \new_[47613]_ ;
  assign \new_[47623]_  = A266 & ~A265;
  assign \new_[47624]_  = A203 & \new_[47623]_ ;
  assign \new_[47627]_  = ~A269 & A267;
  assign \new_[47630]_  = ~A302 & ~A300;
  assign \new_[47631]_  = \new_[47630]_  & \new_[47627]_ ;
  assign \new_[47632]_  = \new_[47631]_  & \new_[47624]_ ;
  assign \new_[47636]_  = A167 & A168;
  assign \new_[47637]_  = A169 & \new_[47636]_ ;
  assign \new_[47641]_  = ~A202 & A201;
  assign \new_[47642]_  = ~A166 & \new_[47641]_ ;
  assign \new_[47643]_  = \new_[47642]_  & \new_[47637]_ ;
  assign \new_[47647]_  = A266 & ~A265;
  assign \new_[47648]_  = A203 & \new_[47647]_ ;
  assign \new_[47651]_  = ~A269 & A267;
  assign \new_[47654]_  = A299 & A298;
  assign \new_[47655]_  = \new_[47654]_  & \new_[47651]_ ;
  assign \new_[47656]_  = \new_[47655]_  & \new_[47648]_ ;
  assign \new_[47660]_  = A167 & A168;
  assign \new_[47661]_  = A169 & \new_[47660]_ ;
  assign \new_[47665]_  = ~A202 & A201;
  assign \new_[47666]_  = ~A166 & \new_[47665]_ ;
  assign \new_[47667]_  = \new_[47666]_  & \new_[47661]_ ;
  assign \new_[47671]_  = A266 & ~A265;
  assign \new_[47672]_  = A203 & \new_[47671]_ ;
  assign \new_[47675]_  = ~A269 & A267;
  assign \new_[47678]_  = ~A299 & ~A298;
  assign \new_[47679]_  = \new_[47678]_  & \new_[47675]_ ;
  assign \new_[47680]_  = \new_[47679]_  & \new_[47672]_ ;
  assign \new_[47684]_  = A167 & A168;
  assign \new_[47685]_  = A169 & \new_[47684]_ ;
  assign \new_[47689]_  = ~A202 & A201;
  assign \new_[47690]_  = ~A166 & \new_[47689]_ ;
  assign \new_[47691]_  = \new_[47690]_  & \new_[47685]_ ;
  assign \new_[47695]_  = ~A266 & A265;
  assign \new_[47696]_  = A203 & \new_[47695]_ ;
  assign \new_[47699]_  = A268 & A267;
  assign \new_[47702]_  = A301 & ~A300;
  assign \new_[47703]_  = \new_[47702]_  & \new_[47699]_ ;
  assign \new_[47704]_  = \new_[47703]_  & \new_[47696]_ ;
  assign \new_[47708]_  = A167 & A168;
  assign \new_[47709]_  = A169 & \new_[47708]_ ;
  assign \new_[47713]_  = ~A202 & A201;
  assign \new_[47714]_  = ~A166 & \new_[47713]_ ;
  assign \new_[47715]_  = \new_[47714]_  & \new_[47709]_ ;
  assign \new_[47719]_  = ~A266 & A265;
  assign \new_[47720]_  = A203 & \new_[47719]_ ;
  assign \new_[47723]_  = A268 & A267;
  assign \new_[47726]_  = ~A302 & ~A300;
  assign \new_[47727]_  = \new_[47726]_  & \new_[47723]_ ;
  assign \new_[47728]_  = \new_[47727]_  & \new_[47720]_ ;
  assign \new_[47732]_  = A167 & A168;
  assign \new_[47733]_  = A169 & \new_[47732]_ ;
  assign \new_[47737]_  = ~A202 & A201;
  assign \new_[47738]_  = ~A166 & \new_[47737]_ ;
  assign \new_[47739]_  = \new_[47738]_  & \new_[47733]_ ;
  assign \new_[47743]_  = ~A266 & A265;
  assign \new_[47744]_  = A203 & \new_[47743]_ ;
  assign \new_[47747]_  = A268 & A267;
  assign \new_[47750]_  = A299 & A298;
  assign \new_[47751]_  = \new_[47750]_  & \new_[47747]_ ;
  assign \new_[47752]_  = \new_[47751]_  & \new_[47744]_ ;
  assign \new_[47756]_  = A167 & A168;
  assign \new_[47757]_  = A169 & \new_[47756]_ ;
  assign \new_[47761]_  = ~A202 & A201;
  assign \new_[47762]_  = ~A166 & \new_[47761]_ ;
  assign \new_[47763]_  = \new_[47762]_  & \new_[47757]_ ;
  assign \new_[47767]_  = ~A266 & A265;
  assign \new_[47768]_  = A203 & \new_[47767]_ ;
  assign \new_[47771]_  = A268 & A267;
  assign \new_[47774]_  = ~A299 & ~A298;
  assign \new_[47775]_  = \new_[47774]_  & \new_[47771]_ ;
  assign \new_[47776]_  = \new_[47775]_  & \new_[47768]_ ;
  assign \new_[47780]_  = A167 & A168;
  assign \new_[47781]_  = A169 & \new_[47780]_ ;
  assign \new_[47785]_  = ~A202 & A201;
  assign \new_[47786]_  = ~A166 & \new_[47785]_ ;
  assign \new_[47787]_  = \new_[47786]_  & \new_[47781]_ ;
  assign \new_[47791]_  = ~A266 & A265;
  assign \new_[47792]_  = A203 & \new_[47791]_ ;
  assign \new_[47795]_  = ~A269 & A267;
  assign \new_[47798]_  = A301 & ~A300;
  assign \new_[47799]_  = \new_[47798]_  & \new_[47795]_ ;
  assign \new_[47800]_  = \new_[47799]_  & \new_[47792]_ ;
  assign \new_[47804]_  = A167 & A168;
  assign \new_[47805]_  = A169 & \new_[47804]_ ;
  assign \new_[47809]_  = ~A202 & A201;
  assign \new_[47810]_  = ~A166 & \new_[47809]_ ;
  assign \new_[47811]_  = \new_[47810]_  & \new_[47805]_ ;
  assign \new_[47815]_  = ~A266 & A265;
  assign \new_[47816]_  = A203 & \new_[47815]_ ;
  assign \new_[47819]_  = ~A269 & A267;
  assign \new_[47822]_  = ~A302 & ~A300;
  assign \new_[47823]_  = \new_[47822]_  & \new_[47819]_ ;
  assign \new_[47824]_  = \new_[47823]_  & \new_[47816]_ ;
  assign \new_[47828]_  = A167 & A168;
  assign \new_[47829]_  = A169 & \new_[47828]_ ;
  assign \new_[47833]_  = ~A202 & A201;
  assign \new_[47834]_  = ~A166 & \new_[47833]_ ;
  assign \new_[47835]_  = \new_[47834]_  & \new_[47829]_ ;
  assign \new_[47839]_  = ~A266 & A265;
  assign \new_[47840]_  = A203 & \new_[47839]_ ;
  assign \new_[47843]_  = ~A269 & A267;
  assign \new_[47846]_  = A299 & A298;
  assign \new_[47847]_  = \new_[47846]_  & \new_[47843]_ ;
  assign \new_[47848]_  = \new_[47847]_  & \new_[47840]_ ;
  assign \new_[47852]_  = A167 & A168;
  assign \new_[47853]_  = A169 & \new_[47852]_ ;
  assign \new_[47857]_  = ~A202 & A201;
  assign \new_[47858]_  = ~A166 & \new_[47857]_ ;
  assign \new_[47859]_  = \new_[47858]_  & \new_[47853]_ ;
  assign \new_[47863]_  = ~A266 & A265;
  assign \new_[47864]_  = A203 & \new_[47863]_ ;
  assign \new_[47867]_  = ~A269 & A267;
  assign \new_[47870]_  = ~A299 & ~A298;
  assign \new_[47871]_  = \new_[47870]_  & \new_[47867]_ ;
  assign \new_[47872]_  = \new_[47871]_  & \new_[47864]_ ;
  assign \new_[47876]_  = A167 & A168;
  assign \new_[47877]_  = A169 & \new_[47876]_ ;
  assign \new_[47881]_  = ~A202 & A201;
  assign \new_[47882]_  = ~A166 & \new_[47881]_ ;
  assign \new_[47883]_  = \new_[47882]_  & \new_[47877]_ ;
  assign \new_[47887]_  = ~A266 & ~A265;
  assign \new_[47888]_  = A203 & \new_[47887]_ ;
  assign \new_[47891]_  = ~A299 & A298;
  assign \new_[47894]_  = A301 & A300;
  assign \new_[47895]_  = \new_[47894]_  & \new_[47891]_ ;
  assign \new_[47896]_  = \new_[47895]_  & \new_[47888]_ ;
  assign \new_[47900]_  = A167 & A168;
  assign \new_[47901]_  = A169 & \new_[47900]_ ;
  assign \new_[47905]_  = ~A202 & A201;
  assign \new_[47906]_  = ~A166 & \new_[47905]_ ;
  assign \new_[47907]_  = \new_[47906]_  & \new_[47901]_ ;
  assign \new_[47911]_  = ~A266 & ~A265;
  assign \new_[47912]_  = A203 & \new_[47911]_ ;
  assign \new_[47915]_  = ~A299 & A298;
  assign \new_[47918]_  = ~A302 & A300;
  assign \new_[47919]_  = \new_[47918]_  & \new_[47915]_ ;
  assign \new_[47920]_  = \new_[47919]_  & \new_[47912]_ ;
  assign \new_[47924]_  = A167 & A168;
  assign \new_[47925]_  = A169 & \new_[47924]_ ;
  assign \new_[47929]_  = ~A202 & A201;
  assign \new_[47930]_  = ~A166 & \new_[47929]_ ;
  assign \new_[47931]_  = \new_[47930]_  & \new_[47925]_ ;
  assign \new_[47935]_  = ~A266 & ~A265;
  assign \new_[47936]_  = A203 & \new_[47935]_ ;
  assign \new_[47939]_  = A299 & ~A298;
  assign \new_[47942]_  = A301 & A300;
  assign \new_[47943]_  = \new_[47942]_  & \new_[47939]_ ;
  assign \new_[47944]_  = \new_[47943]_  & \new_[47936]_ ;
  assign \new_[47948]_  = A167 & A168;
  assign \new_[47949]_  = A169 & \new_[47948]_ ;
  assign \new_[47953]_  = ~A202 & A201;
  assign \new_[47954]_  = ~A166 & \new_[47953]_ ;
  assign \new_[47955]_  = \new_[47954]_  & \new_[47949]_ ;
  assign \new_[47959]_  = ~A266 & ~A265;
  assign \new_[47960]_  = A203 & \new_[47959]_ ;
  assign \new_[47963]_  = A299 & ~A298;
  assign \new_[47966]_  = ~A302 & A300;
  assign \new_[47967]_  = \new_[47966]_  & \new_[47963]_ ;
  assign \new_[47968]_  = \new_[47967]_  & \new_[47960]_ ;
  assign \new_[47972]_  = A167 & A168;
  assign \new_[47973]_  = A169 & \new_[47972]_ ;
  assign \new_[47977]_  = A202 & ~A201;
  assign \new_[47978]_  = ~A166 & \new_[47977]_ ;
  assign \new_[47979]_  = \new_[47978]_  & \new_[47973]_ ;
  assign \new_[47983]_  = A269 & ~A268;
  assign \new_[47984]_  = A267 & \new_[47983]_ ;
  assign \new_[47987]_  = ~A299 & A298;
  assign \new_[47990]_  = A301 & A300;
  assign \new_[47991]_  = \new_[47990]_  & \new_[47987]_ ;
  assign \new_[47992]_  = \new_[47991]_  & \new_[47984]_ ;
  assign \new_[47996]_  = A167 & A168;
  assign \new_[47997]_  = A169 & \new_[47996]_ ;
  assign \new_[48001]_  = A202 & ~A201;
  assign \new_[48002]_  = ~A166 & \new_[48001]_ ;
  assign \new_[48003]_  = \new_[48002]_  & \new_[47997]_ ;
  assign \new_[48007]_  = A269 & ~A268;
  assign \new_[48008]_  = A267 & \new_[48007]_ ;
  assign \new_[48011]_  = ~A299 & A298;
  assign \new_[48014]_  = ~A302 & A300;
  assign \new_[48015]_  = \new_[48014]_  & \new_[48011]_ ;
  assign \new_[48016]_  = \new_[48015]_  & \new_[48008]_ ;
  assign \new_[48020]_  = A167 & A168;
  assign \new_[48021]_  = A169 & \new_[48020]_ ;
  assign \new_[48025]_  = A202 & ~A201;
  assign \new_[48026]_  = ~A166 & \new_[48025]_ ;
  assign \new_[48027]_  = \new_[48026]_  & \new_[48021]_ ;
  assign \new_[48031]_  = A269 & ~A268;
  assign \new_[48032]_  = A267 & \new_[48031]_ ;
  assign \new_[48035]_  = A299 & ~A298;
  assign \new_[48038]_  = A301 & A300;
  assign \new_[48039]_  = \new_[48038]_  & \new_[48035]_ ;
  assign \new_[48040]_  = \new_[48039]_  & \new_[48032]_ ;
  assign \new_[48044]_  = A167 & A168;
  assign \new_[48045]_  = A169 & \new_[48044]_ ;
  assign \new_[48049]_  = A202 & ~A201;
  assign \new_[48050]_  = ~A166 & \new_[48049]_ ;
  assign \new_[48051]_  = \new_[48050]_  & \new_[48045]_ ;
  assign \new_[48055]_  = A269 & ~A268;
  assign \new_[48056]_  = A267 & \new_[48055]_ ;
  assign \new_[48059]_  = A299 & ~A298;
  assign \new_[48062]_  = ~A302 & A300;
  assign \new_[48063]_  = \new_[48062]_  & \new_[48059]_ ;
  assign \new_[48064]_  = \new_[48063]_  & \new_[48056]_ ;
  assign \new_[48068]_  = A167 & A168;
  assign \new_[48069]_  = A169 & \new_[48068]_ ;
  assign \new_[48073]_  = A202 & ~A201;
  assign \new_[48074]_  = ~A166 & \new_[48073]_ ;
  assign \new_[48075]_  = \new_[48074]_  & \new_[48069]_ ;
  assign \new_[48079]_  = A298 & A268;
  assign \new_[48080]_  = ~A267 & \new_[48079]_ ;
  assign \new_[48083]_  = ~A300 & ~A299;
  assign \new_[48086]_  = A302 & ~A301;
  assign \new_[48087]_  = \new_[48086]_  & \new_[48083]_ ;
  assign \new_[48088]_  = \new_[48087]_  & \new_[48080]_ ;
  assign \new_[48092]_  = A167 & A168;
  assign \new_[48093]_  = A169 & \new_[48092]_ ;
  assign \new_[48097]_  = A202 & ~A201;
  assign \new_[48098]_  = ~A166 & \new_[48097]_ ;
  assign \new_[48099]_  = \new_[48098]_  & \new_[48093]_ ;
  assign \new_[48103]_  = ~A298 & A268;
  assign \new_[48104]_  = ~A267 & \new_[48103]_ ;
  assign \new_[48107]_  = ~A300 & A299;
  assign \new_[48110]_  = A302 & ~A301;
  assign \new_[48111]_  = \new_[48110]_  & \new_[48107]_ ;
  assign \new_[48112]_  = \new_[48111]_  & \new_[48104]_ ;
  assign \new_[48116]_  = A167 & A168;
  assign \new_[48117]_  = A169 & \new_[48116]_ ;
  assign \new_[48121]_  = A202 & ~A201;
  assign \new_[48122]_  = ~A166 & \new_[48121]_ ;
  assign \new_[48123]_  = \new_[48122]_  & \new_[48117]_ ;
  assign \new_[48127]_  = A298 & ~A269;
  assign \new_[48128]_  = ~A267 & \new_[48127]_ ;
  assign \new_[48131]_  = ~A300 & ~A299;
  assign \new_[48134]_  = A302 & ~A301;
  assign \new_[48135]_  = \new_[48134]_  & \new_[48131]_ ;
  assign \new_[48136]_  = \new_[48135]_  & \new_[48128]_ ;
  assign \new_[48140]_  = A167 & A168;
  assign \new_[48141]_  = A169 & \new_[48140]_ ;
  assign \new_[48145]_  = A202 & ~A201;
  assign \new_[48146]_  = ~A166 & \new_[48145]_ ;
  assign \new_[48147]_  = \new_[48146]_  & \new_[48141]_ ;
  assign \new_[48151]_  = ~A298 & ~A269;
  assign \new_[48152]_  = ~A267 & \new_[48151]_ ;
  assign \new_[48155]_  = ~A300 & A299;
  assign \new_[48158]_  = A302 & ~A301;
  assign \new_[48159]_  = \new_[48158]_  & \new_[48155]_ ;
  assign \new_[48160]_  = \new_[48159]_  & \new_[48152]_ ;
  assign \new_[48164]_  = A167 & A168;
  assign \new_[48165]_  = A169 & \new_[48164]_ ;
  assign \new_[48169]_  = A202 & ~A201;
  assign \new_[48170]_  = ~A166 & \new_[48169]_ ;
  assign \new_[48171]_  = \new_[48170]_  & \new_[48165]_ ;
  assign \new_[48175]_  = A298 & A266;
  assign \new_[48176]_  = A265 & \new_[48175]_ ;
  assign \new_[48179]_  = ~A300 & ~A299;
  assign \new_[48182]_  = A302 & ~A301;
  assign \new_[48183]_  = \new_[48182]_  & \new_[48179]_ ;
  assign \new_[48184]_  = \new_[48183]_  & \new_[48176]_ ;
  assign \new_[48188]_  = A167 & A168;
  assign \new_[48189]_  = A169 & \new_[48188]_ ;
  assign \new_[48193]_  = A202 & ~A201;
  assign \new_[48194]_  = ~A166 & \new_[48193]_ ;
  assign \new_[48195]_  = \new_[48194]_  & \new_[48189]_ ;
  assign \new_[48199]_  = ~A298 & A266;
  assign \new_[48200]_  = A265 & \new_[48199]_ ;
  assign \new_[48203]_  = ~A300 & A299;
  assign \new_[48206]_  = A302 & ~A301;
  assign \new_[48207]_  = \new_[48206]_  & \new_[48203]_ ;
  assign \new_[48208]_  = \new_[48207]_  & \new_[48200]_ ;
  assign \new_[48212]_  = A167 & A168;
  assign \new_[48213]_  = A169 & \new_[48212]_ ;
  assign \new_[48217]_  = A202 & ~A201;
  assign \new_[48218]_  = ~A166 & \new_[48217]_ ;
  assign \new_[48219]_  = \new_[48218]_  & \new_[48213]_ ;
  assign \new_[48223]_  = A267 & A266;
  assign \new_[48224]_  = ~A265 & \new_[48223]_ ;
  assign \new_[48227]_  = A300 & A268;
  assign \new_[48230]_  = A302 & ~A301;
  assign \new_[48231]_  = \new_[48230]_  & \new_[48227]_ ;
  assign \new_[48232]_  = \new_[48231]_  & \new_[48224]_ ;
  assign \new_[48236]_  = A167 & A168;
  assign \new_[48237]_  = A169 & \new_[48236]_ ;
  assign \new_[48241]_  = A202 & ~A201;
  assign \new_[48242]_  = ~A166 & \new_[48241]_ ;
  assign \new_[48243]_  = \new_[48242]_  & \new_[48237]_ ;
  assign \new_[48247]_  = A267 & A266;
  assign \new_[48248]_  = ~A265 & \new_[48247]_ ;
  assign \new_[48251]_  = A300 & ~A269;
  assign \new_[48254]_  = A302 & ~A301;
  assign \new_[48255]_  = \new_[48254]_  & \new_[48251]_ ;
  assign \new_[48256]_  = \new_[48255]_  & \new_[48248]_ ;
  assign \new_[48260]_  = A167 & A168;
  assign \new_[48261]_  = A169 & \new_[48260]_ ;
  assign \new_[48265]_  = A202 & ~A201;
  assign \new_[48266]_  = ~A166 & \new_[48265]_ ;
  assign \new_[48267]_  = \new_[48266]_  & \new_[48261]_ ;
  assign \new_[48271]_  = ~A267 & A266;
  assign \new_[48272]_  = ~A265 & \new_[48271]_ ;
  assign \new_[48275]_  = A269 & ~A268;
  assign \new_[48278]_  = A301 & ~A300;
  assign \new_[48279]_  = \new_[48278]_  & \new_[48275]_ ;
  assign \new_[48280]_  = \new_[48279]_  & \new_[48272]_ ;
  assign \new_[48284]_  = A167 & A168;
  assign \new_[48285]_  = A169 & \new_[48284]_ ;
  assign \new_[48289]_  = A202 & ~A201;
  assign \new_[48290]_  = ~A166 & \new_[48289]_ ;
  assign \new_[48291]_  = \new_[48290]_  & \new_[48285]_ ;
  assign \new_[48295]_  = ~A267 & A266;
  assign \new_[48296]_  = ~A265 & \new_[48295]_ ;
  assign \new_[48299]_  = A269 & ~A268;
  assign \new_[48302]_  = ~A302 & ~A300;
  assign \new_[48303]_  = \new_[48302]_  & \new_[48299]_ ;
  assign \new_[48304]_  = \new_[48303]_  & \new_[48296]_ ;
  assign \new_[48308]_  = A167 & A168;
  assign \new_[48309]_  = A169 & \new_[48308]_ ;
  assign \new_[48313]_  = A202 & ~A201;
  assign \new_[48314]_  = ~A166 & \new_[48313]_ ;
  assign \new_[48315]_  = \new_[48314]_  & \new_[48309]_ ;
  assign \new_[48319]_  = ~A267 & A266;
  assign \new_[48320]_  = ~A265 & \new_[48319]_ ;
  assign \new_[48323]_  = A269 & ~A268;
  assign \new_[48326]_  = A299 & A298;
  assign \new_[48327]_  = \new_[48326]_  & \new_[48323]_ ;
  assign \new_[48328]_  = \new_[48327]_  & \new_[48320]_ ;
  assign \new_[48332]_  = A167 & A168;
  assign \new_[48333]_  = A169 & \new_[48332]_ ;
  assign \new_[48337]_  = A202 & ~A201;
  assign \new_[48338]_  = ~A166 & \new_[48337]_ ;
  assign \new_[48339]_  = \new_[48338]_  & \new_[48333]_ ;
  assign \new_[48343]_  = ~A267 & A266;
  assign \new_[48344]_  = ~A265 & \new_[48343]_ ;
  assign \new_[48347]_  = A269 & ~A268;
  assign \new_[48350]_  = ~A299 & ~A298;
  assign \new_[48351]_  = \new_[48350]_  & \new_[48347]_ ;
  assign \new_[48352]_  = \new_[48351]_  & \new_[48344]_ ;
  assign \new_[48356]_  = A167 & A168;
  assign \new_[48357]_  = A169 & \new_[48356]_ ;
  assign \new_[48361]_  = A202 & ~A201;
  assign \new_[48362]_  = ~A166 & \new_[48361]_ ;
  assign \new_[48363]_  = \new_[48362]_  & \new_[48357]_ ;
  assign \new_[48367]_  = A267 & ~A266;
  assign \new_[48368]_  = A265 & \new_[48367]_ ;
  assign \new_[48371]_  = A300 & A268;
  assign \new_[48374]_  = A302 & ~A301;
  assign \new_[48375]_  = \new_[48374]_  & \new_[48371]_ ;
  assign \new_[48376]_  = \new_[48375]_  & \new_[48368]_ ;
  assign \new_[48380]_  = A167 & A168;
  assign \new_[48381]_  = A169 & \new_[48380]_ ;
  assign \new_[48385]_  = A202 & ~A201;
  assign \new_[48386]_  = ~A166 & \new_[48385]_ ;
  assign \new_[48387]_  = \new_[48386]_  & \new_[48381]_ ;
  assign \new_[48391]_  = A267 & ~A266;
  assign \new_[48392]_  = A265 & \new_[48391]_ ;
  assign \new_[48395]_  = A300 & ~A269;
  assign \new_[48398]_  = A302 & ~A301;
  assign \new_[48399]_  = \new_[48398]_  & \new_[48395]_ ;
  assign \new_[48400]_  = \new_[48399]_  & \new_[48392]_ ;
  assign \new_[48404]_  = A167 & A168;
  assign \new_[48405]_  = A169 & \new_[48404]_ ;
  assign \new_[48409]_  = A202 & ~A201;
  assign \new_[48410]_  = ~A166 & \new_[48409]_ ;
  assign \new_[48411]_  = \new_[48410]_  & \new_[48405]_ ;
  assign \new_[48415]_  = ~A267 & ~A266;
  assign \new_[48416]_  = A265 & \new_[48415]_ ;
  assign \new_[48419]_  = A269 & ~A268;
  assign \new_[48422]_  = A301 & ~A300;
  assign \new_[48423]_  = \new_[48422]_  & \new_[48419]_ ;
  assign \new_[48424]_  = \new_[48423]_  & \new_[48416]_ ;
  assign \new_[48428]_  = A167 & A168;
  assign \new_[48429]_  = A169 & \new_[48428]_ ;
  assign \new_[48433]_  = A202 & ~A201;
  assign \new_[48434]_  = ~A166 & \new_[48433]_ ;
  assign \new_[48435]_  = \new_[48434]_  & \new_[48429]_ ;
  assign \new_[48439]_  = ~A267 & ~A266;
  assign \new_[48440]_  = A265 & \new_[48439]_ ;
  assign \new_[48443]_  = A269 & ~A268;
  assign \new_[48446]_  = ~A302 & ~A300;
  assign \new_[48447]_  = \new_[48446]_  & \new_[48443]_ ;
  assign \new_[48448]_  = \new_[48447]_  & \new_[48440]_ ;
  assign \new_[48452]_  = A167 & A168;
  assign \new_[48453]_  = A169 & \new_[48452]_ ;
  assign \new_[48457]_  = A202 & ~A201;
  assign \new_[48458]_  = ~A166 & \new_[48457]_ ;
  assign \new_[48459]_  = \new_[48458]_  & \new_[48453]_ ;
  assign \new_[48463]_  = ~A267 & ~A266;
  assign \new_[48464]_  = A265 & \new_[48463]_ ;
  assign \new_[48467]_  = A269 & ~A268;
  assign \new_[48470]_  = A299 & A298;
  assign \new_[48471]_  = \new_[48470]_  & \new_[48467]_ ;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48464]_ ;
  assign \new_[48476]_  = A167 & A168;
  assign \new_[48477]_  = A169 & \new_[48476]_ ;
  assign \new_[48481]_  = A202 & ~A201;
  assign \new_[48482]_  = ~A166 & \new_[48481]_ ;
  assign \new_[48483]_  = \new_[48482]_  & \new_[48477]_ ;
  assign \new_[48487]_  = ~A267 & ~A266;
  assign \new_[48488]_  = A265 & \new_[48487]_ ;
  assign \new_[48491]_  = A269 & ~A268;
  assign \new_[48494]_  = ~A299 & ~A298;
  assign \new_[48495]_  = \new_[48494]_  & \new_[48491]_ ;
  assign \new_[48496]_  = \new_[48495]_  & \new_[48488]_ ;
  assign \new_[48500]_  = A167 & A168;
  assign \new_[48501]_  = A169 & \new_[48500]_ ;
  assign \new_[48505]_  = A202 & ~A201;
  assign \new_[48506]_  = ~A166 & \new_[48505]_ ;
  assign \new_[48507]_  = \new_[48506]_  & \new_[48501]_ ;
  assign \new_[48511]_  = A298 & ~A266;
  assign \new_[48512]_  = ~A265 & \new_[48511]_ ;
  assign \new_[48515]_  = ~A300 & ~A299;
  assign \new_[48518]_  = A302 & ~A301;
  assign \new_[48519]_  = \new_[48518]_  & \new_[48515]_ ;
  assign \new_[48520]_  = \new_[48519]_  & \new_[48512]_ ;
  assign \new_[48524]_  = A167 & A168;
  assign \new_[48525]_  = A169 & \new_[48524]_ ;
  assign \new_[48529]_  = A202 & ~A201;
  assign \new_[48530]_  = ~A166 & \new_[48529]_ ;
  assign \new_[48531]_  = \new_[48530]_  & \new_[48525]_ ;
  assign \new_[48535]_  = ~A298 & ~A266;
  assign \new_[48536]_  = ~A265 & \new_[48535]_ ;
  assign \new_[48539]_  = ~A300 & A299;
  assign \new_[48542]_  = A302 & ~A301;
  assign \new_[48543]_  = \new_[48542]_  & \new_[48539]_ ;
  assign \new_[48544]_  = \new_[48543]_  & \new_[48536]_ ;
  assign \new_[48548]_  = A167 & A168;
  assign \new_[48549]_  = A169 & \new_[48548]_ ;
  assign \new_[48553]_  = ~A203 & ~A201;
  assign \new_[48554]_  = ~A166 & \new_[48553]_ ;
  assign \new_[48555]_  = \new_[48554]_  & \new_[48549]_ ;
  assign \new_[48559]_  = A269 & ~A268;
  assign \new_[48560]_  = A267 & \new_[48559]_ ;
  assign \new_[48563]_  = ~A299 & A298;
  assign \new_[48566]_  = A301 & A300;
  assign \new_[48567]_  = \new_[48566]_  & \new_[48563]_ ;
  assign \new_[48568]_  = \new_[48567]_  & \new_[48560]_ ;
  assign \new_[48572]_  = A167 & A168;
  assign \new_[48573]_  = A169 & \new_[48572]_ ;
  assign \new_[48577]_  = ~A203 & ~A201;
  assign \new_[48578]_  = ~A166 & \new_[48577]_ ;
  assign \new_[48579]_  = \new_[48578]_  & \new_[48573]_ ;
  assign \new_[48583]_  = A269 & ~A268;
  assign \new_[48584]_  = A267 & \new_[48583]_ ;
  assign \new_[48587]_  = ~A299 & A298;
  assign \new_[48590]_  = ~A302 & A300;
  assign \new_[48591]_  = \new_[48590]_  & \new_[48587]_ ;
  assign \new_[48592]_  = \new_[48591]_  & \new_[48584]_ ;
  assign \new_[48596]_  = A167 & A168;
  assign \new_[48597]_  = A169 & \new_[48596]_ ;
  assign \new_[48601]_  = ~A203 & ~A201;
  assign \new_[48602]_  = ~A166 & \new_[48601]_ ;
  assign \new_[48603]_  = \new_[48602]_  & \new_[48597]_ ;
  assign \new_[48607]_  = A269 & ~A268;
  assign \new_[48608]_  = A267 & \new_[48607]_ ;
  assign \new_[48611]_  = A299 & ~A298;
  assign \new_[48614]_  = A301 & A300;
  assign \new_[48615]_  = \new_[48614]_  & \new_[48611]_ ;
  assign \new_[48616]_  = \new_[48615]_  & \new_[48608]_ ;
  assign \new_[48620]_  = A167 & A168;
  assign \new_[48621]_  = A169 & \new_[48620]_ ;
  assign \new_[48625]_  = ~A203 & ~A201;
  assign \new_[48626]_  = ~A166 & \new_[48625]_ ;
  assign \new_[48627]_  = \new_[48626]_  & \new_[48621]_ ;
  assign \new_[48631]_  = A269 & ~A268;
  assign \new_[48632]_  = A267 & \new_[48631]_ ;
  assign \new_[48635]_  = A299 & ~A298;
  assign \new_[48638]_  = ~A302 & A300;
  assign \new_[48639]_  = \new_[48638]_  & \new_[48635]_ ;
  assign \new_[48640]_  = \new_[48639]_  & \new_[48632]_ ;
  assign \new_[48644]_  = A167 & A168;
  assign \new_[48645]_  = A169 & \new_[48644]_ ;
  assign \new_[48649]_  = ~A203 & ~A201;
  assign \new_[48650]_  = ~A166 & \new_[48649]_ ;
  assign \new_[48651]_  = \new_[48650]_  & \new_[48645]_ ;
  assign \new_[48655]_  = A298 & A268;
  assign \new_[48656]_  = ~A267 & \new_[48655]_ ;
  assign \new_[48659]_  = ~A300 & ~A299;
  assign \new_[48662]_  = A302 & ~A301;
  assign \new_[48663]_  = \new_[48662]_  & \new_[48659]_ ;
  assign \new_[48664]_  = \new_[48663]_  & \new_[48656]_ ;
  assign \new_[48668]_  = A167 & A168;
  assign \new_[48669]_  = A169 & \new_[48668]_ ;
  assign \new_[48673]_  = ~A203 & ~A201;
  assign \new_[48674]_  = ~A166 & \new_[48673]_ ;
  assign \new_[48675]_  = \new_[48674]_  & \new_[48669]_ ;
  assign \new_[48679]_  = ~A298 & A268;
  assign \new_[48680]_  = ~A267 & \new_[48679]_ ;
  assign \new_[48683]_  = ~A300 & A299;
  assign \new_[48686]_  = A302 & ~A301;
  assign \new_[48687]_  = \new_[48686]_  & \new_[48683]_ ;
  assign \new_[48688]_  = \new_[48687]_  & \new_[48680]_ ;
  assign \new_[48692]_  = A167 & A168;
  assign \new_[48693]_  = A169 & \new_[48692]_ ;
  assign \new_[48697]_  = ~A203 & ~A201;
  assign \new_[48698]_  = ~A166 & \new_[48697]_ ;
  assign \new_[48699]_  = \new_[48698]_  & \new_[48693]_ ;
  assign \new_[48703]_  = A298 & ~A269;
  assign \new_[48704]_  = ~A267 & \new_[48703]_ ;
  assign \new_[48707]_  = ~A300 & ~A299;
  assign \new_[48710]_  = A302 & ~A301;
  assign \new_[48711]_  = \new_[48710]_  & \new_[48707]_ ;
  assign \new_[48712]_  = \new_[48711]_  & \new_[48704]_ ;
  assign \new_[48716]_  = A167 & A168;
  assign \new_[48717]_  = A169 & \new_[48716]_ ;
  assign \new_[48721]_  = ~A203 & ~A201;
  assign \new_[48722]_  = ~A166 & \new_[48721]_ ;
  assign \new_[48723]_  = \new_[48722]_  & \new_[48717]_ ;
  assign \new_[48727]_  = ~A298 & ~A269;
  assign \new_[48728]_  = ~A267 & \new_[48727]_ ;
  assign \new_[48731]_  = ~A300 & A299;
  assign \new_[48734]_  = A302 & ~A301;
  assign \new_[48735]_  = \new_[48734]_  & \new_[48731]_ ;
  assign \new_[48736]_  = \new_[48735]_  & \new_[48728]_ ;
  assign \new_[48740]_  = A167 & A168;
  assign \new_[48741]_  = A169 & \new_[48740]_ ;
  assign \new_[48745]_  = ~A203 & ~A201;
  assign \new_[48746]_  = ~A166 & \new_[48745]_ ;
  assign \new_[48747]_  = \new_[48746]_  & \new_[48741]_ ;
  assign \new_[48751]_  = A298 & A266;
  assign \new_[48752]_  = A265 & \new_[48751]_ ;
  assign \new_[48755]_  = ~A300 & ~A299;
  assign \new_[48758]_  = A302 & ~A301;
  assign \new_[48759]_  = \new_[48758]_  & \new_[48755]_ ;
  assign \new_[48760]_  = \new_[48759]_  & \new_[48752]_ ;
  assign \new_[48764]_  = A167 & A168;
  assign \new_[48765]_  = A169 & \new_[48764]_ ;
  assign \new_[48769]_  = ~A203 & ~A201;
  assign \new_[48770]_  = ~A166 & \new_[48769]_ ;
  assign \new_[48771]_  = \new_[48770]_  & \new_[48765]_ ;
  assign \new_[48775]_  = ~A298 & A266;
  assign \new_[48776]_  = A265 & \new_[48775]_ ;
  assign \new_[48779]_  = ~A300 & A299;
  assign \new_[48782]_  = A302 & ~A301;
  assign \new_[48783]_  = \new_[48782]_  & \new_[48779]_ ;
  assign \new_[48784]_  = \new_[48783]_  & \new_[48776]_ ;
  assign \new_[48788]_  = A167 & A168;
  assign \new_[48789]_  = A169 & \new_[48788]_ ;
  assign \new_[48793]_  = ~A203 & ~A201;
  assign \new_[48794]_  = ~A166 & \new_[48793]_ ;
  assign \new_[48795]_  = \new_[48794]_  & \new_[48789]_ ;
  assign \new_[48799]_  = A267 & A266;
  assign \new_[48800]_  = ~A265 & \new_[48799]_ ;
  assign \new_[48803]_  = A300 & A268;
  assign \new_[48806]_  = A302 & ~A301;
  assign \new_[48807]_  = \new_[48806]_  & \new_[48803]_ ;
  assign \new_[48808]_  = \new_[48807]_  & \new_[48800]_ ;
  assign \new_[48812]_  = A167 & A168;
  assign \new_[48813]_  = A169 & \new_[48812]_ ;
  assign \new_[48817]_  = ~A203 & ~A201;
  assign \new_[48818]_  = ~A166 & \new_[48817]_ ;
  assign \new_[48819]_  = \new_[48818]_  & \new_[48813]_ ;
  assign \new_[48823]_  = A267 & A266;
  assign \new_[48824]_  = ~A265 & \new_[48823]_ ;
  assign \new_[48827]_  = A300 & ~A269;
  assign \new_[48830]_  = A302 & ~A301;
  assign \new_[48831]_  = \new_[48830]_  & \new_[48827]_ ;
  assign \new_[48832]_  = \new_[48831]_  & \new_[48824]_ ;
  assign \new_[48836]_  = A167 & A168;
  assign \new_[48837]_  = A169 & \new_[48836]_ ;
  assign \new_[48841]_  = ~A203 & ~A201;
  assign \new_[48842]_  = ~A166 & \new_[48841]_ ;
  assign \new_[48843]_  = \new_[48842]_  & \new_[48837]_ ;
  assign \new_[48847]_  = ~A267 & A266;
  assign \new_[48848]_  = ~A265 & \new_[48847]_ ;
  assign \new_[48851]_  = A269 & ~A268;
  assign \new_[48854]_  = A301 & ~A300;
  assign \new_[48855]_  = \new_[48854]_  & \new_[48851]_ ;
  assign \new_[48856]_  = \new_[48855]_  & \new_[48848]_ ;
  assign \new_[48860]_  = A167 & A168;
  assign \new_[48861]_  = A169 & \new_[48860]_ ;
  assign \new_[48865]_  = ~A203 & ~A201;
  assign \new_[48866]_  = ~A166 & \new_[48865]_ ;
  assign \new_[48867]_  = \new_[48866]_  & \new_[48861]_ ;
  assign \new_[48871]_  = ~A267 & A266;
  assign \new_[48872]_  = ~A265 & \new_[48871]_ ;
  assign \new_[48875]_  = A269 & ~A268;
  assign \new_[48878]_  = ~A302 & ~A300;
  assign \new_[48879]_  = \new_[48878]_  & \new_[48875]_ ;
  assign \new_[48880]_  = \new_[48879]_  & \new_[48872]_ ;
  assign \new_[48884]_  = A167 & A168;
  assign \new_[48885]_  = A169 & \new_[48884]_ ;
  assign \new_[48889]_  = ~A203 & ~A201;
  assign \new_[48890]_  = ~A166 & \new_[48889]_ ;
  assign \new_[48891]_  = \new_[48890]_  & \new_[48885]_ ;
  assign \new_[48895]_  = ~A267 & A266;
  assign \new_[48896]_  = ~A265 & \new_[48895]_ ;
  assign \new_[48899]_  = A269 & ~A268;
  assign \new_[48902]_  = A299 & A298;
  assign \new_[48903]_  = \new_[48902]_  & \new_[48899]_ ;
  assign \new_[48904]_  = \new_[48903]_  & \new_[48896]_ ;
  assign \new_[48908]_  = A167 & A168;
  assign \new_[48909]_  = A169 & \new_[48908]_ ;
  assign \new_[48913]_  = ~A203 & ~A201;
  assign \new_[48914]_  = ~A166 & \new_[48913]_ ;
  assign \new_[48915]_  = \new_[48914]_  & \new_[48909]_ ;
  assign \new_[48919]_  = ~A267 & A266;
  assign \new_[48920]_  = ~A265 & \new_[48919]_ ;
  assign \new_[48923]_  = A269 & ~A268;
  assign \new_[48926]_  = ~A299 & ~A298;
  assign \new_[48927]_  = \new_[48926]_  & \new_[48923]_ ;
  assign \new_[48928]_  = \new_[48927]_  & \new_[48920]_ ;
  assign \new_[48932]_  = A167 & A168;
  assign \new_[48933]_  = A169 & \new_[48932]_ ;
  assign \new_[48937]_  = ~A203 & ~A201;
  assign \new_[48938]_  = ~A166 & \new_[48937]_ ;
  assign \new_[48939]_  = \new_[48938]_  & \new_[48933]_ ;
  assign \new_[48943]_  = A267 & ~A266;
  assign \new_[48944]_  = A265 & \new_[48943]_ ;
  assign \new_[48947]_  = A300 & A268;
  assign \new_[48950]_  = A302 & ~A301;
  assign \new_[48951]_  = \new_[48950]_  & \new_[48947]_ ;
  assign \new_[48952]_  = \new_[48951]_  & \new_[48944]_ ;
  assign \new_[48956]_  = A167 & A168;
  assign \new_[48957]_  = A169 & \new_[48956]_ ;
  assign \new_[48961]_  = ~A203 & ~A201;
  assign \new_[48962]_  = ~A166 & \new_[48961]_ ;
  assign \new_[48963]_  = \new_[48962]_  & \new_[48957]_ ;
  assign \new_[48967]_  = A267 & ~A266;
  assign \new_[48968]_  = A265 & \new_[48967]_ ;
  assign \new_[48971]_  = A300 & ~A269;
  assign \new_[48974]_  = A302 & ~A301;
  assign \new_[48975]_  = \new_[48974]_  & \new_[48971]_ ;
  assign \new_[48976]_  = \new_[48975]_  & \new_[48968]_ ;
  assign \new_[48980]_  = A167 & A168;
  assign \new_[48981]_  = A169 & \new_[48980]_ ;
  assign \new_[48985]_  = ~A203 & ~A201;
  assign \new_[48986]_  = ~A166 & \new_[48985]_ ;
  assign \new_[48987]_  = \new_[48986]_  & \new_[48981]_ ;
  assign \new_[48991]_  = ~A267 & ~A266;
  assign \new_[48992]_  = A265 & \new_[48991]_ ;
  assign \new_[48995]_  = A269 & ~A268;
  assign \new_[48998]_  = A301 & ~A300;
  assign \new_[48999]_  = \new_[48998]_  & \new_[48995]_ ;
  assign \new_[49000]_  = \new_[48999]_  & \new_[48992]_ ;
  assign \new_[49004]_  = A167 & A168;
  assign \new_[49005]_  = A169 & \new_[49004]_ ;
  assign \new_[49009]_  = ~A203 & ~A201;
  assign \new_[49010]_  = ~A166 & \new_[49009]_ ;
  assign \new_[49011]_  = \new_[49010]_  & \new_[49005]_ ;
  assign \new_[49015]_  = ~A267 & ~A266;
  assign \new_[49016]_  = A265 & \new_[49015]_ ;
  assign \new_[49019]_  = A269 & ~A268;
  assign \new_[49022]_  = ~A302 & ~A300;
  assign \new_[49023]_  = \new_[49022]_  & \new_[49019]_ ;
  assign \new_[49024]_  = \new_[49023]_  & \new_[49016]_ ;
  assign \new_[49028]_  = A167 & A168;
  assign \new_[49029]_  = A169 & \new_[49028]_ ;
  assign \new_[49033]_  = ~A203 & ~A201;
  assign \new_[49034]_  = ~A166 & \new_[49033]_ ;
  assign \new_[49035]_  = \new_[49034]_  & \new_[49029]_ ;
  assign \new_[49039]_  = ~A267 & ~A266;
  assign \new_[49040]_  = A265 & \new_[49039]_ ;
  assign \new_[49043]_  = A269 & ~A268;
  assign \new_[49046]_  = A299 & A298;
  assign \new_[49047]_  = \new_[49046]_  & \new_[49043]_ ;
  assign \new_[49048]_  = \new_[49047]_  & \new_[49040]_ ;
  assign \new_[49052]_  = A167 & A168;
  assign \new_[49053]_  = A169 & \new_[49052]_ ;
  assign \new_[49057]_  = ~A203 & ~A201;
  assign \new_[49058]_  = ~A166 & \new_[49057]_ ;
  assign \new_[49059]_  = \new_[49058]_  & \new_[49053]_ ;
  assign \new_[49063]_  = ~A267 & ~A266;
  assign \new_[49064]_  = A265 & \new_[49063]_ ;
  assign \new_[49067]_  = A269 & ~A268;
  assign \new_[49070]_  = ~A299 & ~A298;
  assign \new_[49071]_  = \new_[49070]_  & \new_[49067]_ ;
  assign \new_[49072]_  = \new_[49071]_  & \new_[49064]_ ;
  assign \new_[49076]_  = A167 & A168;
  assign \new_[49077]_  = A169 & \new_[49076]_ ;
  assign \new_[49081]_  = ~A203 & ~A201;
  assign \new_[49082]_  = ~A166 & \new_[49081]_ ;
  assign \new_[49083]_  = \new_[49082]_  & \new_[49077]_ ;
  assign \new_[49087]_  = A298 & ~A266;
  assign \new_[49088]_  = ~A265 & \new_[49087]_ ;
  assign \new_[49091]_  = ~A300 & ~A299;
  assign \new_[49094]_  = A302 & ~A301;
  assign \new_[49095]_  = \new_[49094]_  & \new_[49091]_ ;
  assign \new_[49096]_  = \new_[49095]_  & \new_[49088]_ ;
  assign \new_[49100]_  = A167 & A168;
  assign \new_[49101]_  = A169 & \new_[49100]_ ;
  assign \new_[49105]_  = ~A203 & ~A201;
  assign \new_[49106]_  = ~A166 & \new_[49105]_ ;
  assign \new_[49107]_  = \new_[49106]_  & \new_[49101]_ ;
  assign \new_[49111]_  = ~A298 & ~A266;
  assign \new_[49112]_  = ~A265 & \new_[49111]_ ;
  assign \new_[49115]_  = ~A300 & A299;
  assign \new_[49118]_  = A302 & ~A301;
  assign \new_[49119]_  = \new_[49118]_  & \new_[49115]_ ;
  assign \new_[49120]_  = \new_[49119]_  & \new_[49112]_ ;
  assign \new_[49124]_  = A167 & A168;
  assign \new_[49125]_  = A169 & \new_[49124]_ ;
  assign \new_[49129]_  = A200 & A199;
  assign \new_[49130]_  = ~A166 & \new_[49129]_ ;
  assign \new_[49131]_  = \new_[49130]_  & \new_[49125]_ ;
  assign \new_[49135]_  = A269 & ~A268;
  assign \new_[49136]_  = A267 & \new_[49135]_ ;
  assign \new_[49139]_  = ~A299 & A298;
  assign \new_[49142]_  = A301 & A300;
  assign \new_[49143]_  = \new_[49142]_  & \new_[49139]_ ;
  assign \new_[49144]_  = \new_[49143]_  & \new_[49136]_ ;
  assign \new_[49148]_  = A167 & A168;
  assign \new_[49149]_  = A169 & \new_[49148]_ ;
  assign \new_[49153]_  = A200 & A199;
  assign \new_[49154]_  = ~A166 & \new_[49153]_ ;
  assign \new_[49155]_  = \new_[49154]_  & \new_[49149]_ ;
  assign \new_[49159]_  = A269 & ~A268;
  assign \new_[49160]_  = A267 & \new_[49159]_ ;
  assign \new_[49163]_  = ~A299 & A298;
  assign \new_[49166]_  = ~A302 & A300;
  assign \new_[49167]_  = \new_[49166]_  & \new_[49163]_ ;
  assign \new_[49168]_  = \new_[49167]_  & \new_[49160]_ ;
  assign \new_[49172]_  = A167 & A168;
  assign \new_[49173]_  = A169 & \new_[49172]_ ;
  assign \new_[49177]_  = A200 & A199;
  assign \new_[49178]_  = ~A166 & \new_[49177]_ ;
  assign \new_[49179]_  = \new_[49178]_  & \new_[49173]_ ;
  assign \new_[49183]_  = A269 & ~A268;
  assign \new_[49184]_  = A267 & \new_[49183]_ ;
  assign \new_[49187]_  = A299 & ~A298;
  assign \new_[49190]_  = A301 & A300;
  assign \new_[49191]_  = \new_[49190]_  & \new_[49187]_ ;
  assign \new_[49192]_  = \new_[49191]_  & \new_[49184]_ ;
  assign \new_[49196]_  = A167 & A168;
  assign \new_[49197]_  = A169 & \new_[49196]_ ;
  assign \new_[49201]_  = A200 & A199;
  assign \new_[49202]_  = ~A166 & \new_[49201]_ ;
  assign \new_[49203]_  = \new_[49202]_  & \new_[49197]_ ;
  assign \new_[49207]_  = A269 & ~A268;
  assign \new_[49208]_  = A267 & \new_[49207]_ ;
  assign \new_[49211]_  = A299 & ~A298;
  assign \new_[49214]_  = ~A302 & A300;
  assign \new_[49215]_  = \new_[49214]_  & \new_[49211]_ ;
  assign \new_[49216]_  = \new_[49215]_  & \new_[49208]_ ;
  assign \new_[49220]_  = A167 & A168;
  assign \new_[49221]_  = A169 & \new_[49220]_ ;
  assign \new_[49225]_  = A200 & A199;
  assign \new_[49226]_  = ~A166 & \new_[49225]_ ;
  assign \new_[49227]_  = \new_[49226]_  & \new_[49221]_ ;
  assign \new_[49231]_  = A298 & A268;
  assign \new_[49232]_  = ~A267 & \new_[49231]_ ;
  assign \new_[49235]_  = ~A300 & ~A299;
  assign \new_[49238]_  = A302 & ~A301;
  assign \new_[49239]_  = \new_[49238]_  & \new_[49235]_ ;
  assign \new_[49240]_  = \new_[49239]_  & \new_[49232]_ ;
  assign \new_[49244]_  = A167 & A168;
  assign \new_[49245]_  = A169 & \new_[49244]_ ;
  assign \new_[49249]_  = A200 & A199;
  assign \new_[49250]_  = ~A166 & \new_[49249]_ ;
  assign \new_[49251]_  = \new_[49250]_  & \new_[49245]_ ;
  assign \new_[49255]_  = ~A298 & A268;
  assign \new_[49256]_  = ~A267 & \new_[49255]_ ;
  assign \new_[49259]_  = ~A300 & A299;
  assign \new_[49262]_  = A302 & ~A301;
  assign \new_[49263]_  = \new_[49262]_  & \new_[49259]_ ;
  assign \new_[49264]_  = \new_[49263]_  & \new_[49256]_ ;
  assign \new_[49268]_  = A167 & A168;
  assign \new_[49269]_  = A169 & \new_[49268]_ ;
  assign \new_[49273]_  = A200 & A199;
  assign \new_[49274]_  = ~A166 & \new_[49273]_ ;
  assign \new_[49275]_  = \new_[49274]_  & \new_[49269]_ ;
  assign \new_[49279]_  = A298 & ~A269;
  assign \new_[49280]_  = ~A267 & \new_[49279]_ ;
  assign \new_[49283]_  = ~A300 & ~A299;
  assign \new_[49286]_  = A302 & ~A301;
  assign \new_[49287]_  = \new_[49286]_  & \new_[49283]_ ;
  assign \new_[49288]_  = \new_[49287]_  & \new_[49280]_ ;
  assign \new_[49292]_  = A167 & A168;
  assign \new_[49293]_  = A169 & \new_[49292]_ ;
  assign \new_[49297]_  = A200 & A199;
  assign \new_[49298]_  = ~A166 & \new_[49297]_ ;
  assign \new_[49299]_  = \new_[49298]_  & \new_[49293]_ ;
  assign \new_[49303]_  = ~A298 & ~A269;
  assign \new_[49304]_  = ~A267 & \new_[49303]_ ;
  assign \new_[49307]_  = ~A300 & A299;
  assign \new_[49310]_  = A302 & ~A301;
  assign \new_[49311]_  = \new_[49310]_  & \new_[49307]_ ;
  assign \new_[49312]_  = \new_[49311]_  & \new_[49304]_ ;
  assign \new_[49316]_  = A167 & A168;
  assign \new_[49317]_  = A169 & \new_[49316]_ ;
  assign \new_[49321]_  = A200 & A199;
  assign \new_[49322]_  = ~A166 & \new_[49321]_ ;
  assign \new_[49323]_  = \new_[49322]_  & \new_[49317]_ ;
  assign \new_[49327]_  = A298 & A266;
  assign \new_[49328]_  = A265 & \new_[49327]_ ;
  assign \new_[49331]_  = ~A300 & ~A299;
  assign \new_[49334]_  = A302 & ~A301;
  assign \new_[49335]_  = \new_[49334]_  & \new_[49331]_ ;
  assign \new_[49336]_  = \new_[49335]_  & \new_[49328]_ ;
  assign \new_[49340]_  = A167 & A168;
  assign \new_[49341]_  = A169 & \new_[49340]_ ;
  assign \new_[49345]_  = A200 & A199;
  assign \new_[49346]_  = ~A166 & \new_[49345]_ ;
  assign \new_[49347]_  = \new_[49346]_  & \new_[49341]_ ;
  assign \new_[49351]_  = ~A298 & A266;
  assign \new_[49352]_  = A265 & \new_[49351]_ ;
  assign \new_[49355]_  = ~A300 & A299;
  assign \new_[49358]_  = A302 & ~A301;
  assign \new_[49359]_  = \new_[49358]_  & \new_[49355]_ ;
  assign \new_[49360]_  = \new_[49359]_  & \new_[49352]_ ;
  assign \new_[49364]_  = A167 & A168;
  assign \new_[49365]_  = A169 & \new_[49364]_ ;
  assign \new_[49369]_  = A200 & A199;
  assign \new_[49370]_  = ~A166 & \new_[49369]_ ;
  assign \new_[49371]_  = \new_[49370]_  & \new_[49365]_ ;
  assign \new_[49375]_  = A267 & A266;
  assign \new_[49376]_  = ~A265 & \new_[49375]_ ;
  assign \new_[49379]_  = A300 & A268;
  assign \new_[49382]_  = A302 & ~A301;
  assign \new_[49383]_  = \new_[49382]_  & \new_[49379]_ ;
  assign \new_[49384]_  = \new_[49383]_  & \new_[49376]_ ;
  assign \new_[49388]_  = A167 & A168;
  assign \new_[49389]_  = A169 & \new_[49388]_ ;
  assign \new_[49393]_  = A200 & A199;
  assign \new_[49394]_  = ~A166 & \new_[49393]_ ;
  assign \new_[49395]_  = \new_[49394]_  & \new_[49389]_ ;
  assign \new_[49399]_  = A267 & A266;
  assign \new_[49400]_  = ~A265 & \new_[49399]_ ;
  assign \new_[49403]_  = A300 & ~A269;
  assign \new_[49406]_  = A302 & ~A301;
  assign \new_[49407]_  = \new_[49406]_  & \new_[49403]_ ;
  assign \new_[49408]_  = \new_[49407]_  & \new_[49400]_ ;
  assign \new_[49412]_  = A167 & A168;
  assign \new_[49413]_  = A169 & \new_[49412]_ ;
  assign \new_[49417]_  = A200 & A199;
  assign \new_[49418]_  = ~A166 & \new_[49417]_ ;
  assign \new_[49419]_  = \new_[49418]_  & \new_[49413]_ ;
  assign \new_[49423]_  = ~A267 & A266;
  assign \new_[49424]_  = ~A265 & \new_[49423]_ ;
  assign \new_[49427]_  = A269 & ~A268;
  assign \new_[49430]_  = A301 & ~A300;
  assign \new_[49431]_  = \new_[49430]_  & \new_[49427]_ ;
  assign \new_[49432]_  = \new_[49431]_  & \new_[49424]_ ;
  assign \new_[49436]_  = A167 & A168;
  assign \new_[49437]_  = A169 & \new_[49436]_ ;
  assign \new_[49441]_  = A200 & A199;
  assign \new_[49442]_  = ~A166 & \new_[49441]_ ;
  assign \new_[49443]_  = \new_[49442]_  & \new_[49437]_ ;
  assign \new_[49447]_  = ~A267 & A266;
  assign \new_[49448]_  = ~A265 & \new_[49447]_ ;
  assign \new_[49451]_  = A269 & ~A268;
  assign \new_[49454]_  = ~A302 & ~A300;
  assign \new_[49455]_  = \new_[49454]_  & \new_[49451]_ ;
  assign \new_[49456]_  = \new_[49455]_  & \new_[49448]_ ;
  assign \new_[49460]_  = A167 & A168;
  assign \new_[49461]_  = A169 & \new_[49460]_ ;
  assign \new_[49465]_  = A200 & A199;
  assign \new_[49466]_  = ~A166 & \new_[49465]_ ;
  assign \new_[49467]_  = \new_[49466]_  & \new_[49461]_ ;
  assign \new_[49471]_  = ~A267 & A266;
  assign \new_[49472]_  = ~A265 & \new_[49471]_ ;
  assign \new_[49475]_  = A269 & ~A268;
  assign \new_[49478]_  = A299 & A298;
  assign \new_[49479]_  = \new_[49478]_  & \new_[49475]_ ;
  assign \new_[49480]_  = \new_[49479]_  & \new_[49472]_ ;
  assign \new_[49484]_  = A167 & A168;
  assign \new_[49485]_  = A169 & \new_[49484]_ ;
  assign \new_[49489]_  = A200 & A199;
  assign \new_[49490]_  = ~A166 & \new_[49489]_ ;
  assign \new_[49491]_  = \new_[49490]_  & \new_[49485]_ ;
  assign \new_[49495]_  = ~A267 & A266;
  assign \new_[49496]_  = ~A265 & \new_[49495]_ ;
  assign \new_[49499]_  = A269 & ~A268;
  assign \new_[49502]_  = ~A299 & ~A298;
  assign \new_[49503]_  = \new_[49502]_  & \new_[49499]_ ;
  assign \new_[49504]_  = \new_[49503]_  & \new_[49496]_ ;
  assign \new_[49508]_  = A167 & A168;
  assign \new_[49509]_  = A169 & \new_[49508]_ ;
  assign \new_[49513]_  = A200 & A199;
  assign \new_[49514]_  = ~A166 & \new_[49513]_ ;
  assign \new_[49515]_  = \new_[49514]_  & \new_[49509]_ ;
  assign \new_[49519]_  = A267 & ~A266;
  assign \new_[49520]_  = A265 & \new_[49519]_ ;
  assign \new_[49523]_  = A300 & A268;
  assign \new_[49526]_  = A302 & ~A301;
  assign \new_[49527]_  = \new_[49526]_  & \new_[49523]_ ;
  assign \new_[49528]_  = \new_[49527]_  & \new_[49520]_ ;
  assign \new_[49532]_  = A167 & A168;
  assign \new_[49533]_  = A169 & \new_[49532]_ ;
  assign \new_[49537]_  = A200 & A199;
  assign \new_[49538]_  = ~A166 & \new_[49537]_ ;
  assign \new_[49539]_  = \new_[49538]_  & \new_[49533]_ ;
  assign \new_[49543]_  = A267 & ~A266;
  assign \new_[49544]_  = A265 & \new_[49543]_ ;
  assign \new_[49547]_  = A300 & ~A269;
  assign \new_[49550]_  = A302 & ~A301;
  assign \new_[49551]_  = \new_[49550]_  & \new_[49547]_ ;
  assign \new_[49552]_  = \new_[49551]_  & \new_[49544]_ ;
  assign \new_[49556]_  = A167 & A168;
  assign \new_[49557]_  = A169 & \new_[49556]_ ;
  assign \new_[49561]_  = A200 & A199;
  assign \new_[49562]_  = ~A166 & \new_[49561]_ ;
  assign \new_[49563]_  = \new_[49562]_  & \new_[49557]_ ;
  assign \new_[49567]_  = ~A267 & ~A266;
  assign \new_[49568]_  = A265 & \new_[49567]_ ;
  assign \new_[49571]_  = A269 & ~A268;
  assign \new_[49574]_  = A301 & ~A300;
  assign \new_[49575]_  = \new_[49574]_  & \new_[49571]_ ;
  assign \new_[49576]_  = \new_[49575]_  & \new_[49568]_ ;
  assign \new_[49580]_  = A167 & A168;
  assign \new_[49581]_  = A169 & \new_[49580]_ ;
  assign \new_[49585]_  = A200 & A199;
  assign \new_[49586]_  = ~A166 & \new_[49585]_ ;
  assign \new_[49587]_  = \new_[49586]_  & \new_[49581]_ ;
  assign \new_[49591]_  = ~A267 & ~A266;
  assign \new_[49592]_  = A265 & \new_[49591]_ ;
  assign \new_[49595]_  = A269 & ~A268;
  assign \new_[49598]_  = ~A302 & ~A300;
  assign \new_[49599]_  = \new_[49598]_  & \new_[49595]_ ;
  assign \new_[49600]_  = \new_[49599]_  & \new_[49592]_ ;
  assign \new_[49604]_  = A167 & A168;
  assign \new_[49605]_  = A169 & \new_[49604]_ ;
  assign \new_[49609]_  = A200 & A199;
  assign \new_[49610]_  = ~A166 & \new_[49609]_ ;
  assign \new_[49611]_  = \new_[49610]_  & \new_[49605]_ ;
  assign \new_[49615]_  = ~A267 & ~A266;
  assign \new_[49616]_  = A265 & \new_[49615]_ ;
  assign \new_[49619]_  = A269 & ~A268;
  assign \new_[49622]_  = A299 & A298;
  assign \new_[49623]_  = \new_[49622]_  & \new_[49619]_ ;
  assign \new_[49624]_  = \new_[49623]_  & \new_[49616]_ ;
  assign \new_[49628]_  = A167 & A168;
  assign \new_[49629]_  = A169 & \new_[49628]_ ;
  assign \new_[49633]_  = A200 & A199;
  assign \new_[49634]_  = ~A166 & \new_[49633]_ ;
  assign \new_[49635]_  = \new_[49634]_  & \new_[49629]_ ;
  assign \new_[49639]_  = ~A267 & ~A266;
  assign \new_[49640]_  = A265 & \new_[49639]_ ;
  assign \new_[49643]_  = A269 & ~A268;
  assign \new_[49646]_  = ~A299 & ~A298;
  assign \new_[49647]_  = \new_[49646]_  & \new_[49643]_ ;
  assign \new_[49648]_  = \new_[49647]_  & \new_[49640]_ ;
  assign \new_[49652]_  = A167 & A168;
  assign \new_[49653]_  = A169 & \new_[49652]_ ;
  assign \new_[49657]_  = A200 & A199;
  assign \new_[49658]_  = ~A166 & \new_[49657]_ ;
  assign \new_[49659]_  = \new_[49658]_  & \new_[49653]_ ;
  assign \new_[49663]_  = A298 & ~A266;
  assign \new_[49664]_  = ~A265 & \new_[49663]_ ;
  assign \new_[49667]_  = ~A300 & ~A299;
  assign \new_[49670]_  = A302 & ~A301;
  assign \new_[49671]_  = \new_[49670]_  & \new_[49667]_ ;
  assign \new_[49672]_  = \new_[49671]_  & \new_[49664]_ ;
  assign \new_[49676]_  = A167 & A168;
  assign \new_[49677]_  = A169 & \new_[49676]_ ;
  assign \new_[49681]_  = A200 & A199;
  assign \new_[49682]_  = ~A166 & \new_[49681]_ ;
  assign \new_[49683]_  = \new_[49682]_  & \new_[49677]_ ;
  assign \new_[49687]_  = ~A298 & ~A266;
  assign \new_[49688]_  = ~A265 & \new_[49687]_ ;
  assign \new_[49691]_  = ~A300 & A299;
  assign \new_[49694]_  = A302 & ~A301;
  assign \new_[49695]_  = \new_[49694]_  & \new_[49691]_ ;
  assign \new_[49696]_  = \new_[49695]_  & \new_[49688]_ ;
  assign \new_[49700]_  = A167 & A168;
  assign \new_[49701]_  = A169 & \new_[49700]_ ;
  assign \new_[49705]_  = ~A200 & ~A199;
  assign \new_[49706]_  = ~A166 & \new_[49705]_ ;
  assign \new_[49707]_  = \new_[49706]_  & \new_[49701]_ ;
  assign \new_[49711]_  = A269 & ~A268;
  assign \new_[49712]_  = A267 & \new_[49711]_ ;
  assign \new_[49715]_  = ~A299 & A298;
  assign \new_[49718]_  = A301 & A300;
  assign \new_[49719]_  = \new_[49718]_  & \new_[49715]_ ;
  assign \new_[49720]_  = \new_[49719]_  & \new_[49712]_ ;
  assign \new_[49724]_  = A167 & A168;
  assign \new_[49725]_  = A169 & \new_[49724]_ ;
  assign \new_[49729]_  = ~A200 & ~A199;
  assign \new_[49730]_  = ~A166 & \new_[49729]_ ;
  assign \new_[49731]_  = \new_[49730]_  & \new_[49725]_ ;
  assign \new_[49735]_  = A269 & ~A268;
  assign \new_[49736]_  = A267 & \new_[49735]_ ;
  assign \new_[49739]_  = ~A299 & A298;
  assign \new_[49742]_  = ~A302 & A300;
  assign \new_[49743]_  = \new_[49742]_  & \new_[49739]_ ;
  assign \new_[49744]_  = \new_[49743]_  & \new_[49736]_ ;
  assign \new_[49748]_  = A167 & A168;
  assign \new_[49749]_  = A169 & \new_[49748]_ ;
  assign \new_[49753]_  = ~A200 & ~A199;
  assign \new_[49754]_  = ~A166 & \new_[49753]_ ;
  assign \new_[49755]_  = \new_[49754]_  & \new_[49749]_ ;
  assign \new_[49759]_  = A269 & ~A268;
  assign \new_[49760]_  = A267 & \new_[49759]_ ;
  assign \new_[49763]_  = A299 & ~A298;
  assign \new_[49766]_  = A301 & A300;
  assign \new_[49767]_  = \new_[49766]_  & \new_[49763]_ ;
  assign \new_[49768]_  = \new_[49767]_  & \new_[49760]_ ;
  assign \new_[49772]_  = A167 & A168;
  assign \new_[49773]_  = A169 & \new_[49772]_ ;
  assign \new_[49777]_  = ~A200 & ~A199;
  assign \new_[49778]_  = ~A166 & \new_[49777]_ ;
  assign \new_[49779]_  = \new_[49778]_  & \new_[49773]_ ;
  assign \new_[49783]_  = A269 & ~A268;
  assign \new_[49784]_  = A267 & \new_[49783]_ ;
  assign \new_[49787]_  = A299 & ~A298;
  assign \new_[49790]_  = ~A302 & A300;
  assign \new_[49791]_  = \new_[49790]_  & \new_[49787]_ ;
  assign \new_[49792]_  = \new_[49791]_  & \new_[49784]_ ;
  assign \new_[49796]_  = A167 & A168;
  assign \new_[49797]_  = A169 & \new_[49796]_ ;
  assign \new_[49801]_  = ~A200 & ~A199;
  assign \new_[49802]_  = ~A166 & \new_[49801]_ ;
  assign \new_[49803]_  = \new_[49802]_  & \new_[49797]_ ;
  assign \new_[49807]_  = A298 & A268;
  assign \new_[49808]_  = ~A267 & \new_[49807]_ ;
  assign \new_[49811]_  = ~A300 & ~A299;
  assign \new_[49814]_  = A302 & ~A301;
  assign \new_[49815]_  = \new_[49814]_  & \new_[49811]_ ;
  assign \new_[49816]_  = \new_[49815]_  & \new_[49808]_ ;
  assign \new_[49820]_  = A167 & A168;
  assign \new_[49821]_  = A169 & \new_[49820]_ ;
  assign \new_[49825]_  = ~A200 & ~A199;
  assign \new_[49826]_  = ~A166 & \new_[49825]_ ;
  assign \new_[49827]_  = \new_[49826]_  & \new_[49821]_ ;
  assign \new_[49831]_  = ~A298 & A268;
  assign \new_[49832]_  = ~A267 & \new_[49831]_ ;
  assign \new_[49835]_  = ~A300 & A299;
  assign \new_[49838]_  = A302 & ~A301;
  assign \new_[49839]_  = \new_[49838]_  & \new_[49835]_ ;
  assign \new_[49840]_  = \new_[49839]_  & \new_[49832]_ ;
  assign \new_[49844]_  = A167 & A168;
  assign \new_[49845]_  = A169 & \new_[49844]_ ;
  assign \new_[49849]_  = ~A200 & ~A199;
  assign \new_[49850]_  = ~A166 & \new_[49849]_ ;
  assign \new_[49851]_  = \new_[49850]_  & \new_[49845]_ ;
  assign \new_[49855]_  = A298 & ~A269;
  assign \new_[49856]_  = ~A267 & \new_[49855]_ ;
  assign \new_[49859]_  = ~A300 & ~A299;
  assign \new_[49862]_  = A302 & ~A301;
  assign \new_[49863]_  = \new_[49862]_  & \new_[49859]_ ;
  assign \new_[49864]_  = \new_[49863]_  & \new_[49856]_ ;
  assign \new_[49868]_  = A167 & A168;
  assign \new_[49869]_  = A169 & \new_[49868]_ ;
  assign \new_[49873]_  = ~A200 & ~A199;
  assign \new_[49874]_  = ~A166 & \new_[49873]_ ;
  assign \new_[49875]_  = \new_[49874]_  & \new_[49869]_ ;
  assign \new_[49879]_  = ~A298 & ~A269;
  assign \new_[49880]_  = ~A267 & \new_[49879]_ ;
  assign \new_[49883]_  = ~A300 & A299;
  assign \new_[49886]_  = A302 & ~A301;
  assign \new_[49887]_  = \new_[49886]_  & \new_[49883]_ ;
  assign \new_[49888]_  = \new_[49887]_  & \new_[49880]_ ;
  assign \new_[49892]_  = A167 & A168;
  assign \new_[49893]_  = A169 & \new_[49892]_ ;
  assign \new_[49897]_  = ~A200 & ~A199;
  assign \new_[49898]_  = ~A166 & \new_[49897]_ ;
  assign \new_[49899]_  = \new_[49898]_  & \new_[49893]_ ;
  assign \new_[49903]_  = A298 & A266;
  assign \new_[49904]_  = A265 & \new_[49903]_ ;
  assign \new_[49907]_  = ~A300 & ~A299;
  assign \new_[49910]_  = A302 & ~A301;
  assign \new_[49911]_  = \new_[49910]_  & \new_[49907]_ ;
  assign \new_[49912]_  = \new_[49911]_  & \new_[49904]_ ;
  assign \new_[49916]_  = A167 & A168;
  assign \new_[49917]_  = A169 & \new_[49916]_ ;
  assign \new_[49921]_  = ~A200 & ~A199;
  assign \new_[49922]_  = ~A166 & \new_[49921]_ ;
  assign \new_[49923]_  = \new_[49922]_  & \new_[49917]_ ;
  assign \new_[49927]_  = ~A298 & A266;
  assign \new_[49928]_  = A265 & \new_[49927]_ ;
  assign \new_[49931]_  = ~A300 & A299;
  assign \new_[49934]_  = A302 & ~A301;
  assign \new_[49935]_  = \new_[49934]_  & \new_[49931]_ ;
  assign \new_[49936]_  = \new_[49935]_  & \new_[49928]_ ;
  assign \new_[49940]_  = A167 & A168;
  assign \new_[49941]_  = A169 & \new_[49940]_ ;
  assign \new_[49945]_  = ~A200 & ~A199;
  assign \new_[49946]_  = ~A166 & \new_[49945]_ ;
  assign \new_[49947]_  = \new_[49946]_  & \new_[49941]_ ;
  assign \new_[49951]_  = A267 & A266;
  assign \new_[49952]_  = ~A265 & \new_[49951]_ ;
  assign \new_[49955]_  = A300 & A268;
  assign \new_[49958]_  = A302 & ~A301;
  assign \new_[49959]_  = \new_[49958]_  & \new_[49955]_ ;
  assign \new_[49960]_  = \new_[49959]_  & \new_[49952]_ ;
  assign \new_[49964]_  = A167 & A168;
  assign \new_[49965]_  = A169 & \new_[49964]_ ;
  assign \new_[49969]_  = ~A200 & ~A199;
  assign \new_[49970]_  = ~A166 & \new_[49969]_ ;
  assign \new_[49971]_  = \new_[49970]_  & \new_[49965]_ ;
  assign \new_[49975]_  = A267 & A266;
  assign \new_[49976]_  = ~A265 & \new_[49975]_ ;
  assign \new_[49979]_  = A300 & ~A269;
  assign \new_[49982]_  = A302 & ~A301;
  assign \new_[49983]_  = \new_[49982]_  & \new_[49979]_ ;
  assign \new_[49984]_  = \new_[49983]_  & \new_[49976]_ ;
  assign \new_[49988]_  = A167 & A168;
  assign \new_[49989]_  = A169 & \new_[49988]_ ;
  assign \new_[49993]_  = ~A200 & ~A199;
  assign \new_[49994]_  = ~A166 & \new_[49993]_ ;
  assign \new_[49995]_  = \new_[49994]_  & \new_[49989]_ ;
  assign \new_[49999]_  = ~A267 & A266;
  assign \new_[50000]_  = ~A265 & \new_[49999]_ ;
  assign \new_[50003]_  = A269 & ~A268;
  assign \new_[50006]_  = A301 & ~A300;
  assign \new_[50007]_  = \new_[50006]_  & \new_[50003]_ ;
  assign \new_[50008]_  = \new_[50007]_  & \new_[50000]_ ;
  assign \new_[50012]_  = A167 & A168;
  assign \new_[50013]_  = A169 & \new_[50012]_ ;
  assign \new_[50017]_  = ~A200 & ~A199;
  assign \new_[50018]_  = ~A166 & \new_[50017]_ ;
  assign \new_[50019]_  = \new_[50018]_  & \new_[50013]_ ;
  assign \new_[50023]_  = ~A267 & A266;
  assign \new_[50024]_  = ~A265 & \new_[50023]_ ;
  assign \new_[50027]_  = A269 & ~A268;
  assign \new_[50030]_  = ~A302 & ~A300;
  assign \new_[50031]_  = \new_[50030]_  & \new_[50027]_ ;
  assign \new_[50032]_  = \new_[50031]_  & \new_[50024]_ ;
  assign \new_[50036]_  = A167 & A168;
  assign \new_[50037]_  = A169 & \new_[50036]_ ;
  assign \new_[50041]_  = ~A200 & ~A199;
  assign \new_[50042]_  = ~A166 & \new_[50041]_ ;
  assign \new_[50043]_  = \new_[50042]_  & \new_[50037]_ ;
  assign \new_[50047]_  = ~A267 & A266;
  assign \new_[50048]_  = ~A265 & \new_[50047]_ ;
  assign \new_[50051]_  = A269 & ~A268;
  assign \new_[50054]_  = A299 & A298;
  assign \new_[50055]_  = \new_[50054]_  & \new_[50051]_ ;
  assign \new_[50056]_  = \new_[50055]_  & \new_[50048]_ ;
  assign \new_[50060]_  = A167 & A168;
  assign \new_[50061]_  = A169 & \new_[50060]_ ;
  assign \new_[50065]_  = ~A200 & ~A199;
  assign \new_[50066]_  = ~A166 & \new_[50065]_ ;
  assign \new_[50067]_  = \new_[50066]_  & \new_[50061]_ ;
  assign \new_[50071]_  = ~A267 & A266;
  assign \new_[50072]_  = ~A265 & \new_[50071]_ ;
  assign \new_[50075]_  = A269 & ~A268;
  assign \new_[50078]_  = ~A299 & ~A298;
  assign \new_[50079]_  = \new_[50078]_  & \new_[50075]_ ;
  assign \new_[50080]_  = \new_[50079]_  & \new_[50072]_ ;
  assign \new_[50084]_  = A167 & A168;
  assign \new_[50085]_  = A169 & \new_[50084]_ ;
  assign \new_[50089]_  = ~A200 & ~A199;
  assign \new_[50090]_  = ~A166 & \new_[50089]_ ;
  assign \new_[50091]_  = \new_[50090]_  & \new_[50085]_ ;
  assign \new_[50095]_  = A267 & ~A266;
  assign \new_[50096]_  = A265 & \new_[50095]_ ;
  assign \new_[50099]_  = A300 & A268;
  assign \new_[50102]_  = A302 & ~A301;
  assign \new_[50103]_  = \new_[50102]_  & \new_[50099]_ ;
  assign \new_[50104]_  = \new_[50103]_  & \new_[50096]_ ;
  assign \new_[50108]_  = A167 & A168;
  assign \new_[50109]_  = A169 & \new_[50108]_ ;
  assign \new_[50113]_  = ~A200 & ~A199;
  assign \new_[50114]_  = ~A166 & \new_[50113]_ ;
  assign \new_[50115]_  = \new_[50114]_  & \new_[50109]_ ;
  assign \new_[50119]_  = A267 & ~A266;
  assign \new_[50120]_  = A265 & \new_[50119]_ ;
  assign \new_[50123]_  = A300 & ~A269;
  assign \new_[50126]_  = A302 & ~A301;
  assign \new_[50127]_  = \new_[50126]_  & \new_[50123]_ ;
  assign \new_[50128]_  = \new_[50127]_  & \new_[50120]_ ;
  assign \new_[50132]_  = A167 & A168;
  assign \new_[50133]_  = A169 & \new_[50132]_ ;
  assign \new_[50137]_  = ~A200 & ~A199;
  assign \new_[50138]_  = ~A166 & \new_[50137]_ ;
  assign \new_[50139]_  = \new_[50138]_  & \new_[50133]_ ;
  assign \new_[50143]_  = ~A267 & ~A266;
  assign \new_[50144]_  = A265 & \new_[50143]_ ;
  assign \new_[50147]_  = A269 & ~A268;
  assign \new_[50150]_  = A301 & ~A300;
  assign \new_[50151]_  = \new_[50150]_  & \new_[50147]_ ;
  assign \new_[50152]_  = \new_[50151]_  & \new_[50144]_ ;
  assign \new_[50156]_  = A167 & A168;
  assign \new_[50157]_  = A169 & \new_[50156]_ ;
  assign \new_[50161]_  = ~A200 & ~A199;
  assign \new_[50162]_  = ~A166 & \new_[50161]_ ;
  assign \new_[50163]_  = \new_[50162]_  & \new_[50157]_ ;
  assign \new_[50167]_  = ~A267 & ~A266;
  assign \new_[50168]_  = A265 & \new_[50167]_ ;
  assign \new_[50171]_  = A269 & ~A268;
  assign \new_[50174]_  = ~A302 & ~A300;
  assign \new_[50175]_  = \new_[50174]_  & \new_[50171]_ ;
  assign \new_[50176]_  = \new_[50175]_  & \new_[50168]_ ;
  assign \new_[50180]_  = A167 & A168;
  assign \new_[50181]_  = A169 & \new_[50180]_ ;
  assign \new_[50185]_  = ~A200 & ~A199;
  assign \new_[50186]_  = ~A166 & \new_[50185]_ ;
  assign \new_[50187]_  = \new_[50186]_  & \new_[50181]_ ;
  assign \new_[50191]_  = ~A267 & ~A266;
  assign \new_[50192]_  = A265 & \new_[50191]_ ;
  assign \new_[50195]_  = A269 & ~A268;
  assign \new_[50198]_  = A299 & A298;
  assign \new_[50199]_  = \new_[50198]_  & \new_[50195]_ ;
  assign \new_[50200]_  = \new_[50199]_  & \new_[50192]_ ;
  assign \new_[50204]_  = A167 & A168;
  assign \new_[50205]_  = A169 & \new_[50204]_ ;
  assign \new_[50209]_  = ~A200 & ~A199;
  assign \new_[50210]_  = ~A166 & \new_[50209]_ ;
  assign \new_[50211]_  = \new_[50210]_  & \new_[50205]_ ;
  assign \new_[50215]_  = ~A267 & ~A266;
  assign \new_[50216]_  = A265 & \new_[50215]_ ;
  assign \new_[50219]_  = A269 & ~A268;
  assign \new_[50222]_  = ~A299 & ~A298;
  assign \new_[50223]_  = \new_[50222]_  & \new_[50219]_ ;
  assign \new_[50224]_  = \new_[50223]_  & \new_[50216]_ ;
  assign \new_[50228]_  = A167 & A168;
  assign \new_[50229]_  = A169 & \new_[50228]_ ;
  assign \new_[50233]_  = ~A200 & ~A199;
  assign \new_[50234]_  = ~A166 & \new_[50233]_ ;
  assign \new_[50235]_  = \new_[50234]_  & \new_[50229]_ ;
  assign \new_[50239]_  = A298 & ~A266;
  assign \new_[50240]_  = ~A265 & \new_[50239]_ ;
  assign \new_[50243]_  = ~A300 & ~A299;
  assign \new_[50246]_  = A302 & ~A301;
  assign \new_[50247]_  = \new_[50246]_  & \new_[50243]_ ;
  assign \new_[50248]_  = \new_[50247]_  & \new_[50240]_ ;
  assign \new_[50252]_  = A167 & A168;
  assign \new_[50253]_  = A169 & \new_[50252]_ ;
  assign \new_[50257]_  = ~A200 & ~A199;
  assign \new_[50258]_  = ~A166 & \new_[50257]_ ;
  assign \new_[50259]_  = \new_[50258]_  & \new_[50253]_ ;
  assign \new_[50263]_  = ~A298 & ~A266;
  assign \new_[50264]_  = ~A265 & \new_[50263]_ ;
  assign \new_[50267]_  = ~A300 & A299;
  assign \new_[50270]_  = A302 & ~A301;
  assign \new_[50271]_  = \new_[50270]_  & \new_[50267]_ ;
  assign \new_[50272]_  = \new_[50271]_  & \new_[50264]_ ;
  assign \new_[50276]_  = ~A167 & A168;
  assign \new_[50277]_  = A169 & \new_[50276]_ ;
  assign \new_[50281]_  = ~A202 & A201;
  assign \new_[50282]_  = A166 & \new_[50281]_ ;
  assign \new_[50283]_  = \new_[50282]_  & \new_[50277]_ ;
  assign \new_[50287]_  = A268 & ~A267;
  assign \new_[50288]_  = A203 & \new_[50287]_ ;
  assign \new_[50291]_  = ~A299 & A298;
  assign \new_[50294]_  = A301 & A300;
  assign \new_[50295]_  = \new_[50294]_  & \new_[50291]_ ;
  assign \new_[50296]_  = \new_[50295]_  & \new_[50288]_ ;
  assign \new_[50300]_  = ~A167 & A168;
  assign \new_[50301]_  = A169 & \new_[50300]_ ;
  assign \new_[50305]_  = ~A202 & A201;
  assign \new_[50306]_  = A166 & \new_[50305]_ ;
  assign \new_[50307]_  = \new_[50306]_  & \new_[50301]_ ;
  assign \new_[50311]_  = A268 & ~A267;
  assign \new_[50312]_  = A203 & \new_[50311]_ ;
  assign \new_[50315]_  = ~A299 & A298;
  assign \new_[50318]_  = ~A302 & A300;
  assign \new_[50319]_  = \new_[50318]_  & \new_[50315]_ ;
  assign \new_[50320]_  = \new_[50319]_  & \new_[50312]_ ;
  assign \new_[50324]_  = ~A167 & A168;
  assign \new_[50325]_  = A169 & \new_[50324]_ ;
  assign \new_[50329]_  = ~A202 & A201;
  assign \new_[50330]_  = A166 & \new_[50329]_ ;
  assign \new_[50331]_  = \new_[50330]_  & \new_[50325]_ ;
  assign \new_[50335]_  = A268 & ~A267;
  assign \new_[50336]_  = A203 & \new_[50335]_ ;
  assign \new_[50339]_  = A299 & ~A298;
  assign \new_[50342]_  = A301 & A300;
  assign \new_[50343]_  = \new_[50342]_  & \new_[50339]_ ;
  assign \new_[50344]_  = \new_[50343]_  & \new_[50336]_ ;
  assign \new_[50348]_  = ~A167 & A168;
  assign \new_[50349]_  = A169 & \new_[50348]_ ;
  assign \new_[50353]_  = ~A202 & A201;
  assign \new_[50354]_  = A166 & \new_[50353]_ ;
  assign \new_[50355]_  = \new_[50354]_  & \new_[50349]_ ;
  assign \new_[50359]_  = A268 & ~A267;
  assign \new_[50360]_  = A203 & \new_[50359]_ ;
  assign \new_[50363]_  = A299 & ~A298;
  assign \new_[50366]_  = ~A302 & A300;
  assign \new_[50367]_  = \new_[50366]_  & \new_[50363]_ ;
  assign \new_[50368]_  = \new_[50367]_  & \new_[50360]_ ;
  assign \new_[50372]_  = ~A167 & A168;
  assign \new_[50373]_  = A169 & \new_[50372]_ ;
  assign \new_[50377]_  = ~A202 & A201;
  assign \new_[50378]_  = A166 & \new_[50377]_ ;
  assign \new_[50379]_  = \new_[50378]_  & \new_[50373]_ ;
  assign \new_[50383]_  = ~A269 & ~A267;
  assign \new_[50384]_  = A203 & \new_[50383]_ ;
  assign \new_[50387]_  = ~A299 & A298;
  assign \new_[50390]_  = A301 & A300;
  assign \new_[50391]_  = \new_[50390]_  & \new_[50387]_ ;
  assign \new_[50392]_  = \new_[50391]_  & \new_[50384]_ ;
  assign \new_[50396]_  = ~A167 & A168;
  assign \new_[50397]_  = A169 & \new_[50396]_ ;
  assign \new_[50401]_  = ~A202 & A201;
  assign \new_[50402]_  = A166 & \new_[50401]_ ;
  assign \new_[50403]_  = \new_[50402]_  & \new_[50397]_ ;
  assign \new_[50407]_  = ~A269 & ~A267;
  assign \new_[50408]_  = A203 & \new_[50407]_ ;
  assign \new_[50411]_  = ~A299 & A298;
  assign \new_[50414]_  = ~A302 & A300;
  assign \new_[50415]_  = \new_[50414]_  & \new_[50411]_ ;
  assign \new_[50416]_  = \new_[50415]_  & \new_[50408]_ ;
  assign \new_[50420]_  = ~A167 & A168;
  assign \new_[50421]_  = A169 & \new_[50420]_ ;
  assign \new_[50425]_  = ~A202 & A201;
  assign \new_[50426]_  = A166 & \new_[50425]_ ;
  assign \new_[50427]_  = \new_[50426]_  & \new_[50421]_ ;
  assign \new_[50431]_  = ~A269 & ~A267;
  assign \new_[50432]_  = A203 & \new_[50431]_ ;
  assign \new_[50435]_  = A299 & ~A298;
  assign \new_[50438]_  = A301 & A300;
  assign \new_[50439]_  = \new_[50438]_  & \new_[50435]_ ;
  assign \new_[50440]_  = \new_[50439]_  & \new_[50432]_ ;
  assign \new_[50444]_  = ~A167 & A168;
  assign \new_[50445]_  = A169 & \new_[50444]_ ;
  assign \new_[50449]_  = ~A202 & A201;
  assign \new_[50450]_  = A166 & \new_[50449]_ ;
  assign \new_[50451]_  = \new_[50450]_  & \new_[50445]_ ;
  assign \new_[50455]_  = ~A269 & ~A267;
  assign \new_[50456]_  = A203 & \new_[50455]_ ;
  assign \new_[50459]_  = A299 & ~A298;
  assign \new_[50462]_  = ~A302 & A300;
  assign \new_[50463]_  = \new_[50462]_  & \new_[50459]_ ;
  assign \new_[50464]_  = \new_[50463]_  & \new_[50456]_ ;
  assign \new_[50468]_  = ~A167 & A168;
  assign \new_[50469]_  = A169 & \new_[50468]_ ;
  assign \new_[50473]_  = ~A202 & A201;
  assign \new_[50474]_  = A166 & \new_[50473]_ ;
  assign \new_[50475]_  = \new_[50474]_  & \new_[50469]_ ;
  assign \new_[50479]_  = A266 & A265;
  assign \new_[50480]_  = A203 & \new_[50479]_ ;
  assign \new_[50483]_  = ~A299 & A298;
  assign \new_[50486]_  = A301 & A300;
  assign \new_[50487]_  = \new_[50486]_  & \new_[50483]_ ;
  assign \new_[50488]_  = \new_[50487]_  & \new_[50480]_ ;
  assign \new_[50492]_  = ~A167 & A168;
  assign \new_[50493]_  = A169 & \new_[50492]_ ;
  assign \new_[50497]_  = ~A202 & A201;
  assign \new_[50498]_  = A166 & \new_[50497]_ ;
  assign \new_[50499]_  = \new_[50498]_  & \new_[50493]_ ;
  assign \new_[50503]_  = A266 & A265;
  assign \new_[50504]_  = A203 & \new_[50503]_ ;
  assign \new_[50507]_  = ~A299 & A298;
  assign \new_[50510]_  = ~A302 & A300;
  assign \new_[50511]_  = \new_[50510]_  & \new_[50507]_ ;
  assign \new_[50512]_  = \new_[50511]_  & \new_[50504]_ ;
  assign \new_[50516]_  = ~A167 & A168;
  assign \new_[50517]_  = A169 & \new_[50516]_ ;
  assign \new_[50521]_  = ~A202 & A201;
  assign \new_[50522]_  = A166 & \new_[50521]_ ;
  assign \new_[50523]_  = \new_[50522]_  & \new_[50517]_ ;
  assign \new_[50527]_  = A266 & A265;
  assign \new_[50528]_  = A203 & \new_[50527]_ ;
  assign \new_[50531]_  = A299 & ~A298;
  assign \new_[50534]_  = A301 & A300;
  assign \new_[50535]_  = \new_[50534]_  & \new_[50531]_ ;
  assign \new_[50536]_  = \new_[50535]_  & \new_[50528]_ ;
  assign \new_[50540]_  = ~A167 & A168;
  assign \new_[50541]_  = A169 & \new_[50540]_ ;
  assign \new_[50545]_  = ~A202 & A201;
  assign \new_[50546]_  = A166 & \new_[50545]_ ;
  assign \new_[50547]_  = \new_[50546]_  & \new_[50541]_ ;
  assign \new_[50551]_  = A266 & A265;
  assign \new_[50552]_  = A203 & \new_[50551]_ ;
  assign \new_[50555]_  = A299 & ~A298;
  assign \new_[50558]_  = ~A302 & A300;
  assign \new_[50559]_  = \new_[50558]_  & \new_[50555]_ ;
  assign \new_[50560]_  = \new_[50559]_  & \new_[50552]_ ;
  assign \new_[50564]_  = ~A167 & A168;
  assign \new_[50565]_  = A169 & \new_[50564]_ ;
  assign \new_[50569]_  = ~A202 & A201;
  assign \new_[50570]_  = A166 & \new_[50569]_ ;
  assign \new_[50571]_  = \new_[50570]_  & \new_[50565]_ ;
  assign \new_[50575]_  = A266 & ~A265;
  assign \new_[50576]_  = A203 & \new_[50575]_ ;
  assign \new_[50579]_  = A268 & A267;
  assign \new_[50582]_  = A301 & ~A300;
  assign \new_[50583]_  = \new_[50582]_  & \new_[50579]_ ;
  assign \new_[50584]_  = \new_[50583]_  & \new_[50576]_ ;
  assign \new_[50588]_  = ~A167 & A168;
  assign \new_[50589]_  = A169 & \new_[50588]_ ;
  assign \new_[50593]_  = ~A202 & A201;
  assign \new_[50594]_  = A166 & \new_[50593]_ ;
  assign \new_[50595]_  = \new_[50594]_  & \new_[50589]_ ;
  assign \new_[50599]_  = A266 & ~A265;
  assign \new_[50600]_  = A203 & \new_[50599]_ ;
  assign \new_[50603]_  = A268 & A267;
  assign \new_[50606]_  = ~A302 & ~A300;
  assign \new_[50607]_  = \new_[50606]_  & \new_[50603]_ ;
  assign \new_[50608]_  = \new_[50607]_  & \new_[50600]_ ;
  assign \new_[50612]_  = ~A167 & A168;
  assign \new_[50613]_  = A169 & \new_[50612]_ ;
  assign \new_[50617]_  = ~A202 & A201;
  assign \new_[50618]_  = A166 & \new_[50617]_ ;
  assign \new_[50619]_  = \new_[50618]_  & \new_[50613]_ ;
  assign \new_[50623]_  = A266 & ~A265;
  assign \new_[50624]_  = A203 & \new_[50623]_ ;
  assign \new_[50627]_  = A268 & A267;
  assign \new_[50630]_  = A299 & A298;
  assign \new_[50631]_  = \new_[50630]_  & \new_[50627]_ ;
  assign \new_[50632]_  = \new_[50631]_  & \new_[50624]_ ;
  assign \new_[50636]_  = ~A167 & A168;
  assign \new_[50637]_  = A169 & \new_[50636]_ ;
  assign \new_[50641]_  = ~A202 & A201;
  assign \new_[50642]_  = A166 & \new_[50641]_ ;
  assign \new_[50643]_  = \new_[50642]_  & \new_[50637]_ ;
  assign \new_[50647]_  = A266 & ~A265;
  assign \new_[50648]_  = A203 & \new_[50647]_ ;
  assign \new_[50651]_  = A268 & A267;
  assign \new_[50654]_  = ~A299 & ~A298;
  assign \new_[50655]_  = \new_[50654]_  & \new_[50651]_ ;
  assign \new_[50656]_  = \new_[50655]_  & \new_[50648]_ ;
  assign \new_[50660]_  = ~A167 & A168;
  assign \new_[50661]_  = A169 & \new_[50660]_ ;
  assign \new_[50665]_  = ~A202 & A201;
  assign \new_[50666]_  = A166 & \new_[50665]_ ;
  assign \new_[50667]_  = \new_[50666]_  & \new_[50661]_ ;
  assign \new_[50671]_  = A266 & ~A265;
  assign \new_[50672]_  = A203 & \new_[50671]_ ;
  assign \new_[50675]_  = ~A269 & A267;
  assign \new_[50678]_  = A301 & ~A300;
  assign \new_[50679]_  = \new_[50678]_  & \new_[50675]_ ;
  assign \new_[50680]_  = \new_[50679]_  & \new_[50672]_ ;
  assign \new_[50684]_  = ~A167 & A168;
  assign \new_[50685]_  = A169 & \new_[50684]_ ;
  assign \new_[50689]_  = ~A202 & A201;
  assign \new_[50690]_  = A166 & \new_[50689]_ ;
  assign \new_[50691]_  = \new_[50690]_  & \new_[50685]_ ;
  assign \new_[50695]_  = A266 & ~A265;
  assign \new_[50696]_  = A203 & \new_[50695]_ ;
  assign \new_[50699]_  = ~A269 & A267;
  assign \new_[50702]_  = ~A302 & ~A300;
  assign \new_[50703]_  = \new_[50702]_  & \new_[50699]_ ;
  assign \new_[50704]_  = \new_[50703]_  & \new_[50696]_ ;
  assign \new_[50708]_  = ~A167 & A168;
  assign \new_[50709]_  = A169 & \new_[50708]_ ;
  assign \new_[50713]_  = ~A202 & A201;
  assign \new_[50714]_  = A166 & \new_[50713]_ ;
  assign \new_[50715]_  = \new_[50714]_  & \new_[50709]_ ;
  assign \new_[50719]_  = A266 & ~A265;
  assign \new_[50720]_  = A203 & \new_[50719]_ ;
  assign \new_[50723]_  = ~A269 & A267;
  assign \new_[50726]_  = A299 & A298;
  assign \new_[50727]_  = \new_[50726]_  & \new_[50723]_ ;
  assign \new_[50728]_  = \new_[50727]_  & \new_[50720]_ ;
  assign \new_[50732]_  = ~A167 & A168;
  assign \new_[50733]_  = A169 & \new_[50732]_ ;
  assign \new_[50737]_  = ~A202 & A201;
  assign \new_[50738]_  = A166 & \new_[50737]_ ;
  assign \new_[50739]_  = \new_[50738]_  & \new_[50733]_ ;
  assign \new_[50743]_  = A266 & ~A265;
  assign \new_[50744]_  = A203 & \new_[50743]_ ;
  assign \new_[50747]_  = ~A269 & A267;
  assign \new_[50750]_  = ~A299 & ~A298;
  assign \new_[50751]_  = \new_[50750]_  & \new_[50747]_ ;
  assign \new_[50752]_  = \new_[50751]_  & \new_[50744]_ ;
  assign \new_[50756]_  = ~A167 & A168;
  assign \new_[50757]_  = A169 & \new_[50756]_ ;
  assign \new_[50761]_  = ~A202 & A201;
  assign \new_[50762]_  = A166 & \new_[50761]_ ;
  assign \new_[50763]_  = \new_[50762]_  & \new_[50757]_ ;
  assign \new_[50767]_  = ~A266 & A265;
  assign \new_[50768]_  = A203 & \new_[50767]_ ;
  assign \new_[50771]_  = A268 & A267;
  assign \new_[50774]_  = A301 & ~A300;
  assign \new_[50775]_  = \new_[50774]_  & \new_[50771]_ ;
  assign \new_[50776]_  = \new_[50775]_  & \new_[50768]_ ;
  assign \new_[50780]_  = ~A167 & A168;
  assign \new_[50781]_  = A169 & \new_[50780]_ ;
  assign \new_[50785]_  = ~A202 & A201;
  assign \new_[50786]_  = A166 & \new_[50785]_ ;
  assign \new_[50787]_  = \new_[50786]_  & \new_[50781]_ ;
  assign \new_[50791]_  = ~A266 & A265;
  assign \new_[50792]_  = A203 & \new_[50791]_ ;
  assign \new_[50795]_  = A268 & A267;
  assign \new_[50798]_  = ~A302 & ~A300;
  assign \new_[50799]_  = \new_[50798]_  & \new_[50795]_ ;
  assign \new_[50800]_  = \new_[50799]_  & \new_[50792]_ ;
  assign \new_[50804]_  = ~A167 & A168;
  assign \new_[50805]_  = A169 & \new_[50804]_ ;
  assign \new_[50809]_  = ~A202 & A201;
  assign \new_[50810]_  = A166 & \new_[50809]_ ;
  assign \new_[50811]_  = \new_[50810]_  & \new_[50805]_ ;
  assign \new_[50815]_  = ~A266 & A265;
  assign \new_[50816]_  = A203 & \new_[50815]_ ;
  assign \new_[50819]_  = A268 & A267;
  assign \new_[50822]_  = A299 & A298;
  assign \new_[50823]_  = \new_[50822]_  & \new_[50819]_ ;
  assign \new_[50824]_  = \new_[50823]_  & \new_[50816]_ ;
  assign \new_[50828]_  = ~A167 & A168;
  assign \new_[50829]_  = A169 & \new_[50828]_ ;
  assign \new_[50833]_  = ~A202 & A201;
  assign \new_[50834]_  = A166 & \new_[50833]_ ;
  assign \new_[50835]_  = \new_[50834]_  & \new_[50829]_ ;
  assign \new_[50839]_  = ~A266 & A265;
  assign \new_[50840]_  = A203 & \new_[50839]_ ;
  assign \new_[50843]_  = A268 & A267;
  assign \new_[50846]_  = ~A299 & ~A298;
  assign \new_[50847]_  = \new_[50846]_  & \new_[50843]_ ;
  assign \new_[50848]_  = \new_[50847]_  & \new_[50840]_ ;
  assign \new_[50852]_  = ~A167 & A168;
  assign \new_[50853]_  = A169 & \new_[50852]_ ;
  assign \new_[50857]_  = ~A202 & A201;
  assign \new_[50858]_  = A166 & \new_[50857]_ ;
  assign \new_[50859]_  = \new_[50858]_  & \new_[50853]_ ;
  assign \new_[50863]_  = ~A266 & A265;
  assign \new_[50864]_  = A203 & \new_[50863]_ ;
  assign \new_[50867]_  = ~A269 & A267;
  assign \new_[50870]_  = A301 & ~A300;
  assign \new_[50871]_  = \new_[50870]_  & \new_[50867]_ ;
  assign \new_[50872]_  = \new_[50871]_  & \new_[50864]_ ;
  assign \new_[50876]_  = ~A167 & A168;
  assign \new_[50877]_  = A169 & \new_[50876]_ ;
  assign \new_[50881]_  = ~A202 & A201;
  assign \new_[50882]_  = A166 & \new_[50881]_ ;
  assign \new_[50883]_  = \new_[50882]_  & \new_[50877]_ ;
  assign \new_[50887]_  = ~A266 & A265;
  assign \new_[50888]_  = A203 & \new_[50887]_ ;
  assign \new_[50891]_  = ~A269 & A267;
  assign \new_[50894]_  = ~A302 & ~A300;
  assign \new_[50895]_  = \new_[50894]_  & \new_[50891]_ ;
  assign \new_[50896]_  = \new_[50895]_  & \new_[50888]_ ;
  assign \new_[50900]_  = ~A167 & A168;
  assign \new_[50901]_  = A169 & \new_[50900]_ ;
  assign \new_[50905]_  = ~A202 & A201;
  assign \new_[50906]_  = A166 & \new_[50905]_ ;
  assign \new_[50907]_  = \new_[50906]_  & \new_[50901]_ ;
  assign \new_[50911]_  = ~A266 & A265;
  assign \new_[50912]_  = A203 & \new_[50911]_ ;
  assign \new_[50915]_  = ~A269 & A267;
  assign \new_[50918]_  = A299 & A298;
  assign \new_[50919]_  = \new_[50918]_  & \new_[50915]_ ;
  assign \new_[50920]_  = \new_[50919]_  & \new_[50912]_ ;
  assign \new_[50924]_  = ~A167 & A168;
  assign \new_[50925]_  = A169 & \new_[50924]_ ;
  assign \new_[50929]_  = ~A202 & A201;
  assign \new_[50930]_  = A166 & \new_[50929]_ ;
  assign \new_[50931]_  = \new_[50930]_  & \new_[50925]_ ;
  assign \new_[50935]_  = ~A266 & A265;
  assign \new_[50936]_  = A203 & \new_[50935]_ ;
  assign \new_[50939]_  = ~A269 & A267;
  assign \new_[50942]_  = ~A299 & ~A298;
  assign \new_[50943]_  = \new_[50942]_  & \new_[50939]_ ;
  assign \new_[50944]_  = \new_[50943]_  & \new_[50936]_ ;
  assign \new_[50948]_  = ~A167 & A168;
  assign \new_[50949]_  = A169 & \new_[50948]_ ;
  assign \new_[50953]_  = ~A202 & A201;
  assign \new_[50954]_  = A166 & \new_[50953]_ ;
  assign \new_[50955]_  = \new_[50954]_  & \new_[50949]_ ;
  assign \new_[50959]_  = ~A266 & ~A265;
  assign \new_[50960]_  = A203 & \new_[50959]_ ;
  assign \new_[50963]_  = ~A299 & A298;
  assign \new_[50966]_  = A301 & A300;
  assign \new_[50967]_  = \new_[50966]_  & \new_[50963]_ ;
  assign \new_[50968]_  = \new_[50967]_  & \new_[50960]_ ;
  assign \new_[50972]_  = ~A167 & A168;
  assign \new_[50973]_  = A169 & \new_[50972]_ ;
  assign \new_[50977]_  = ~A202 & A201;
  assign \new_[50978]_  = A166 & \new_[50977]_ ;
  assign \new_[50979]_  = \new_[50978]_  & \new_[50973]_ ;
  assign \new_[50983]_  = ~A266 & ~A265;
  assign \new_[50984]_  = A203 & \new_[50983]_ ;
  assign \new_[50987]_  = ~A299 & A298;
  assign \new_[50990]_  = ~A302 & A300;
  assign \new_[50991]_  = \new_[50990]_  & \new_[50987]_ ;
  assign \new_[50992]_  = \new_[50991]_  & \new_[50984]_ ;
  assign \new_[50996]_  = ~A167 & A168;
  assign \new_[50997]_  = A169 & \new_[50996]_ ;
  assign \new_[51001]_  = ~A202 & A201;
  assign \new_[51002]_  = A166 & \new_[51001]_ ;
  assign \new_[51003]_  = \new_[51002]_  & \new_[50997]_ ;
  assign \new_[51007]_  = ~A266 & ~A265;
  assign \new_[51008]_  = A203 & \new_[51007]_ ;
  assign \new_[51011]_  = A299 & ~A298;
  assign \new_[51014]_  = A301 & A300;
  assign \new_[51015]_  = \new_[51014]_  & \new_[51011]_ ;
  assign \new_[51016]_  = \new_[51015]_  & \new_[51008]_ ;
  assign \new_[51020]_  = ~A167 & A168;
  assign \new_[51021]_  = A169 & \new_[51020]_ ;
  assign \new_[51025]_  = ~A202 & A201;
  assign \new_[51026]_  = A166 & \new_[51025]_ ;
  assign \new_[51027]_  = \new_[51026]_  & \new_[51021]_ ;
  assign \new_[51031]_  = ~A266 & ~A265;
  assign \new_[51032]_  = A203 & \new_[51031]_ ;
  assign \new_[51035]_  = A299 & ~A298;
  assign \new_[51038]_  = ~A302 & A300;
  assign \new_[51039]_  = \new_[51038]_  & \new_[51035]_ ;
  assign \new_[51040]_  = \new_[51039]_  & \new_[51032]_ ;
  assign \new_[51044]_  = ~A167 & A168;
  assign \new_[51045]_  = A169 & \new_[51044]_ ;
  assign \new_[51049]_  = A202 & ~A201;
  assign \new_[51050]_  = A166 & \new_[51049]_ ;
  assign \new_[51051]_  = \new_[51050]_  & \new_[51045]_ ;
  assign \new_[51055]_  = A269 & ~A268;
  assign \new_[51056]_  = A267 & \new_[51055]_ ;
  assign \new_[51059]_  = ~A299 & A298;
  assign \new_[51062]_  = A301 & A300;
  assign \new_[51063]_  = \new_[51062]_  & \new_[51059]_ ;
  assign \new_[51064]_  = \new_[51063]_  & \new_[51056]_ ;
  assign \new_[51068]_  = ~A167 & A168;
  assign \new_[51069]_  = A169 & \new_[51068]_ ;
  assign \new_[51073]_  = A202 & ~A201;
  assign \new_[51074]_  = A166 & \new_[51073]_ ;
  assign \new_[51075]_  = \new_[51074]_  & \new_[51069]_ ;
  assign \new_[51079]_  = A269 & ~A268;
  assign \new_[51080]_  = A267 & \new_[51079]_ ;
  assign \new_[51083]_  = ~A299 & A298;
  assign \new_[51086]_  = ~A302 & A300;
  assign \new_[51087]_  = \new_[51086]_  & \new_[51083]_ ;
  assign \new_[51088]_  = \new_[51087]_  & \new_[51080]_ ;
  assign \new_[51092]_  = ~A167 & A168;
  assign \new_[51093]_  = A169 & \new_[51092]_ ;
  assign \new_[51097]_  = A202 & ~A201;
  assign \new_[51098]_  = A166 & \new_[51097]_ ;
  assign \new_[51099]_  = \new_[51098]_  & \new_[51093]_ ;
  assign \new_[51103]_  = A269 & ~A268;
  assign \new_[51104]_  = A267 & \new_[51103]_ ;
  assign \new_[51107]_  = A299 & ~A298;
  assign \new_[51110]_  = A301 & A300;
  assign \new_[51111]_  = \new_[51110]_  & \new_[51107]_ ;
  assign \new_[51112]_  = \new_[51111]_  & \new_[51104]_ ;
  assign \new_[51116]_  = ~A167 & A168;
  assign \new_[51117]_  = A169 & \new_[51116]_ ;
  assign \new_[51121]_  = A202 & ~A201;
  assign \new_[51122]_  = A166 & \new_[51121]_ ;
  assign \new_[51123]_  = \new_[51122]_  & \new_[51117]_ ;
  assign \new_[51127]_  = A269 & ~A268;
  assign \new_[51128]_  = A267 & \new_[51127]_ ;
  assign \new_[51131]_  = A299 & ~A298;
  assign \new_[51134]_  = ~A302 & A300;
  assign \new_[51135]_  = \new_[51134]_  & \new_[51131]_ ;
  assign \new_[51136]_  = \new_[51135]_  & \new_[51128]_ ;
  assign \new_[51140]_  = ~A167 & A168;
  assign \new_[51141]_  = A169 & \new_[51140]_ ;
  assign \new_[51145]_  = A202 & ~A201;
  assign \new_[51146]_  = A166 & \new_[51145]_ ;
  assign \new_[51147]_  = \new_[51146]_  & \new_[51141]_ ;
  assign \new_[51151]_  = A298 & A268;
  assign \new_[51152]_  = ~A267 & \new_[51151]_ ;
  assign \new_[51155]_  = ~A300 & ~A299;
  assign \new_[51158]_  = A302 & ~A301;
  assign \new_[51159]_  = \new_[51158]_  & \new_[51155]_ ;
  assign \new_[51160]_  = \new_[51159]_  & \new_[51152]_ ;
  assign \new_[51164]_  = ~A167 & A168;
  assign \new_[51165]_  = A169 & \new_[51164]_ ;
  assign \new_[51169]_  = A202 & ~A201;
  assign \new_[51170]_  = A166 & \new_[51169]_ ;
  assign \new_[51171]_  = \new_[51170]_  & \new_[51165]_ ;
  assign \new_[51175]_  = ~A298 & A268;
  assign \new_[51176]_  = ~A267 & \new_[51175]_ ;
  assign \new_[51179]_  = ~A300 & A299;
  assign \new_[51182]_  = A302 & ~A301;
  assign \new_[51183]_  = \new_[51182]_  & \new_[51179]_ ;
  assign \new_[51184]_  = \new_[51183]_  & \new_[51176]_ ;
  assign \new_[51188]_  = ~A167 & A168;
  assign \new_[51189]_  = A169 & \new_[51188]_ ;
  assign \new_[51193]_  = A202 & ~A201;
  assign \new_[51194]_  = A166 & \new_[51193]_ ;
  assign \new_[51195]_  = \new_[51194]_  & \new_[51189]_ ;
  assign \new_[51199]_  = A298 & ~A269;
  assign \new_[51200]_  = ~A267 & \new_[51199]_ ;
  assign \new_[51203]_  = ~A300 & ~A299;
  assign \new_[51206]_  = A302 & ~A301;
  assign \new_[51207]_  = \new_[51206]_  & \new_[51203]_ ;
  assign \new_[51208]_  = \new_[51207]_  & \new_[51200]_ ;
  assign \new_[51212]_  = ~A167 & A168;
  assign \new_[51213]_  = A169 & \new_[51212]_ ;
  assign \new_[51217]_  = A202 & ~A201;
  assign \new_[51218]_  = A166 & \new_[51217]_ ;
  assign \new_[51219]_  = \new_[51218]_  & \new_[51213]_ ;
  assign \new_[51223]_  = ~A298 & ~A269;
  assign \new_[51224]_  = ~A267 & \new_[51223]_ ;
  assign \new_[51227]_  = ~A300 & A299;
  assign \new_[51230]_  = A302 & ~A301;
  assign \new_[51231]_  = \new_[51230]_  & \new_[51227]_ ;
  assign \new_[51232]_  = \new_[51231]_  & \new_[51224]_ ;
  assign \new_[51236]_  = ~A167 & A168;
  assign \new_[51237]_  = A169 & \new_[51236]_ ;
  assign \new_[51241]_  = A202 & ~A201;
  assign \new_[51242]_  = A166 & \new_[51241]_ ;
  assign \new_[51243]_  = \new_[51242]_  & \new_[51237]_ ;
  assign \new_[51247]_  = A298 & A266;
  assign \new_[51248]_  = A265 & \new_[51247]_ ;
  assign \new_[51251]_  = ~A300 & ~A299;
  assign \new_[51254]_  = A302 & ~A301;
  assign \new_[51255]_  = \new_[51254]_  & \new_[51251]_ ;
  assign \new_[51256]_  = \new_[51255]_  & \new_[51248]_ ;
  assign \new_[51260]_  = ~A167 & A168;
  assign \new_[51261]_  = A169 & \new_[51260]_ ;
  assign \new_[51265]_  = A202 & ~A201;
  assign \new_[51266]_  = A166 & \new_[51265]_ ;
  assign \new_[51267]_  = \new_[51266]_  & \new_[51261]_ ;
  assign \new_[51271]_  = ~A298 & A266;
  assign \new_[51272]_  = A265 & \new_[51271]_ ;
  assign \new_[51275]_  = ~A300 & A299;
  assign \new_[51278]_  = A302 & ~A301;
  assign \new_[51279]_  = \new_[51278]_  & \new_[51275]_ ;
  assign \new_[51280]_  = \new_[51279]_  & \new_[51272]_ ;
  assign \new_[51284]_  = ~A167 & A168;
  assign \new_[51285]_  = A169 & \new_[51284]_ ;
  assign \new_[51289]_  = A202 & ~A201;
  assign \new_[51290]_  = A166 & \new_[51289]_ ;
  assign \new_[51291]_  = \new_[51290]_  & \new_[51285]_ ;
  assign \new_[51295]_  = A267 & A266;
  assign \new_[51296]_  = ~A265 & \new_[51295]_ ;
  assign \new_[51299]_  = A300 & A268;
  assign \new_[51302]_  = A302 & ~A301;
  assign \new_[51303]_  = \new_[51302]_  & \new_[51299]_ ;
  assign \new_[51304]_  = \new_[51303]_  & \new_[51296]_ ;
  assign \new_[51308]_  = ~A167 & A168;
  assign \new_[51309]_  = A169 & \new_[51308]_ ;
  assign \new_[51313]_  = A202 & ~A201;
  assign \new_[51314]_  = A166 & \new_[51313]_ ;
  assign \new_[51315]_  = \new_[51314]_  & \new_[51309]_ ;
  assign \new_[51319]_  = A267 & A266;
  assign \new_[51320]_  = ~A265 & \new_[51319]_ ;
  assign \new_[51323]_  = A300 & ~A269;
  assign \new_[51326]_  = A302 & ~A301;
  assign \new_[51327]_  = \new_[51326]_  & \new_[51323]_ ;
  assign \new_[51328]_  = \new_[51327]_  & \new_[51320]_ ;
  assign \new_[51332]_  = ~A167 & A168;
  assign \new_[51333]_  = A169 & \new_[51332]_ ;
  assign \new_[51337]_  = A202 & ~A201;
  assign \new_[51338]_  = A166 & \new_[51337]_ ;
  assign \new_[51339]_  = \new_[51338]_  & \new_[51333]_ ;
  assign \new_[51343]_  = ~A267 & A266;
  assign \new_[51344]_  = ~A265 & \new_[51343]_ ;
  assign \new_[51347]_  = A269 & ~A268;
  assign \new_[51350]_  = A301 & ~A300;
  assign \new_[51351]_  = \new_[51350]_  & \new_[51347]_ ;
  assign \new_[51352]_  = \new_[51351]_  & \new_[51344]_ ;
  assign \new_[51356]_  = ~A167 & A168;
  assign \new_[51357]_  = A169 & \new_[51356]_ ;
  assign \new_[51361]_  = A202 & ~A201;
  assign \new_[51362]_  = A166 & \new_[51361]_ ;
  assign \new_[51363]_  = \new_[51362]_  & \new_[51357]_ ;
  assign \new_[51367]_  = ~A267 & A266;
  assign \new_[51368]_  = ~A265 & \new_[51367]_ ;
  assign \new_[51371]_  = A269 & ~A268;
  assign \new_[51374]_  = ~A302 & ~A300;
  assign \new_[51375]_  = \new_[51374]_  & \new_[51371]_ ;
  assign \new_[51376]_  = \new_[51375]_  & \new_[51368]_ ;
  assign \new_[51380]_  = ~A167 & A168;
  assign \new_[51381]_  = A169 & \new_[51380]_ ;
  assign \new_[51385]_  = A202 & ~A201;
  assign \new_[51386]_  = A166 & \new_[51385]_ ;
  assign \new_[51387]_  = \new_[51386]_  & \new_[51381]_ ;
  assign \new_[51391]_  = ~A267 & A266;
  assign \new_[51392]_  = ~A265 & \new_[51391]_ ;
  assign \new_[51395]_  = A269 & ~A268;
  assign \new_[51398]_  = A299 & A298;
  assign \new_[51399]_  = \new_[51398]_  & \new_[51395]_ ;
  assign \new_[51400]_  = \new_[51399]_  & \new_[51392]_ ;
  assign \new_[51404]_  = ~A167 & A168;
  assign \new_[51405]_  = A169 & \new_[51404]_ ;
  assign \new_[51409]_  = A202 & ~A201;
  assign \new_[51410]_  = A166 & \new_[51409]_ ;
  assign \new_[51411]_  = \new_[51410]_  & \new_[51405]_ ;
  assign \new_[51415]_  = ~A267 & A266;
  assign \new_[51416]_  = ~A265 & \new_[51415]_ ;
  assign \new_[51419]_  = A269 & ~A268;
  assign \new_[51422]_  = ~A299 & ~A298;
  assign \new_[51423]_  = \new_[51422]_  & \new_[51419]_ ;
  assign \new_[51424]_  = \new_[51423]_  & \new_[51416]_ ;
  assign \new_[51428]_  = ~A167 & A168;
  assign \new_[51429]_  = A169 & \new_[51428]_ ;
  assign \new_[51433]_  = A202 & ~A201;
  assign \new_[51434]_  = A166 & \new_[51433]_ ;
  assign \new_[51435]_  = \new_[51434]_  & \new_[51429]_ ;
  assign \new_[51439]_  = A267 & ~A266;
  assign \new_[51440]_  = A265 & \new_[51439]_ ;
  assign \new_[51443]_  = A300 & A268;
  assign \new_[51446]_  = A302 & ~A301;
  assign \new_[51447]_  = \new_[51446]_  & \new_[51443]_ ;
  assign \new_[51448]_  = \new_[51447]_  & \new_[51440]_ ;
  assign \new_[51452]_  = ~A167 & A168;
  assign \new_[51453]_  = A169 & \new_[51452]_ ;
  assign \new_[51457]_  = A202 & ~A201;
  assign \new_[51458]_  = A166 & \new_[51457]_ ;
  assign \new_[51459]_  = \new_[51458]_  & \new_[51453]_ ;
  assign \new_[51463]_  = A267 & ~A266;
  assign \new_[51464]_  = A265 & \new_[51463]_ ;
  assign \new_[51467]_  = A300 & ~A269;
  assign \new_[51470]_  = A302 & ~A301;
  assign \new_[51471]_  = \new_[51470]_  & \new_[51467]_ ;
  assign \new_[51472]_  = \new_[51471]_  & \new_[51464]_ ;
  assign \new_[51476]_  = ~A167 & A168;
  assign \new_[51477]_  = A169 & \new_[51476]_ ;
  assign \new_[51481]_  = A202 & ~A201;
  assign \new_[51482]_  = A166 & \new_[51481]_ ;
  assign \new_[51483]_  = \new_[51482]_  & \new_[51477]_ ;
  assign \new_[51487]_  = ~A267 & ~A266;
  assign \new_[51488]_  = A265 & \new_[51487]_ ;
  assign \new_[51491]_  = A269 & ~A268;
  assign \new_[51494]_  = A301 & ~A300;
  assign \new_[51495]_  = \new_[51494]_  & \new_[51491]_ ;
  assign \new_[51496]_  = \new_[51495]_  & \new_[51488]_ ;
  assign \new_[51500]_  = ~A167 & A168;
  assign \new_[51501]_  = A169 & \new_[51500]_ ;
  assign \new_[51505]_  = A202 & ~A201;
  assign \new_[51506]_  = A166 & \new_[51505]_ ;
  assign \new_[51507]_  = \new_[51506]_  & \new_[51501]_ ;
  assign \new_[51511]_  = ~A267 & ~A266;
  assign \new_[51512]_  = A265 & \new_[51511]_ ;
  assign \new_[51515]_  = A269 & ~A268;
  assign \new_[51518]_  = ~A302 & ~A300;
  assign \new_[51519]_  = \new_[51518]_  & \new_[51515]_ ;
  assign \new_[51520]_  = \new_[51519]_  & \new_[51512]_ ;
  assign \new_[51524]_  = ~A167 & A168;
  assign \new_[51525]_  = A169 & \new_[51524]_ ;
  assign \new_[51529]_  = A202 & ~A201;
  assign \new_[51530]_  = A166 & \new_[51529]_ ;
  assign \new_[51531]_  = \new_[51530]_  & \new_[51525]_ ;
  assign \new_[51535]_  = ~A267 & ~A266;
  assign \new_[51536]_  = A265 & \new_[51535]_ ;
  assign \new_[51539]_  = A269 & ~A268;
  assign \new_[51542]_  = A299 & A298;
  assign \new_[51543]_  = \new_[51542]_  & \new_[51539]_ ;
  assign \new_[51544]_  = \new_[51543]_  & \new_[51536]_ ;
  assign \new_[51548]_  = ~A167 & A168;
  assign \new_[51549]_  = A169 & \new_[51548]_ ;
  assign \new_[51553]_  = A202 & ~A201;
  assign \new_[51554]_  = A166 & \new_[51553]_ ;
  assign \new_[51555]_  = \new_[51554]_  & \new_[51549]_ ;
  assign \new_[51559]_  = ~A267 & ~A266;
  assign \new_[51560]_  = A265 & \new_[51559]_ ;
  assign \new_[51563]_  = A269 & ~A268;
  assign \new_[51566]_  = ~A299 & ~A298;
  assign \new_[51567]_  = \new_[51566]_  & \new_[51563]_ ;
  assign \new_[51568]_  = \new_[51567]_  & \new_[51560]_ ;
  assign \new_[51572]_  = ~A167 & A168;
  assign \new_[51573]_  = A169 & \new_[51572]_ ;
  assign \new_[51577]_  = A202 & ~A201;
  assign \new_[51578]_  = A166 & \new_[51577]_ ;
  assign \new_[51579]_  = \new_[51578]_  & \new_[51573]_ ;
  assign \new_[51583]_  = A298 & ~A266;
  assign \new_[51584]_  = ~A265 & \new_[51583]_ ;
  assign \new_[51587]_  = ~A300 & ~A299;
  assign \new_[51590]_  = A302 & ~A301;
  assign \new_[51591]_  = \new_[51590]_  & \new_[51587]_ ;
  assign \new_[51592]_  = \new_[51591]_  & \new_[51584]_ ;
  assign \new_[51596]_  = ~A167 & A168;
  assign \new_[51597]_  = A169 & \new_[51596]_ ;
  assign \new_[51601]_  = A202 & ~A201;
  assign \new_[51602]_  = A166 & \new_[51601]_ ;
  assign \new_[51603]_  = \new_[51602]_  & \new_[51597]_ ;
  assign \new_[51607]_  = ~A298 & ~A266;
  assign \new_[51608]_  = ~A265 & \new_[51607]_ ;
  assign \new_[51611]_  = ~A300 & A299;
  assign \new_[51614]_  = A302 & ~A301;
  assign \new_[51615]_  = \new_[51614]_  & \new_[51611]_ ;
  assign \new_[51616]_  = \new_[51615]_  & \new_[51608]_ ;
  assign \new_[51620]_  = ~A167 & A168;
  assign \new_[51621]_  = A169 & \new_[51620]_ ;
  assign \new_[51625]_  = ~A203 & ~A201;
  assign \new_[51626]_  = A166 & \new_[51625]_ ;
  assign \new_[51627]_  = \new_[51626]_  & \new_[51621]_ ;
  assign \new_[51631]_  = A269 & ~A268;
  assign \new_[51632]_  = A267 & \new_[51631]_ ;
  assign \new_[51635]_  = ~A299 & A298;
  assign \new_[51638]_  = A301 & A300;
  assign \new_[51639]_  = \new_[51638]_  & \new_[51635]_ ;
  assign \new_[51640]_  = \new_[51639]_  & \new_[51632]_ ;
  assign \new_[51644]_  = ~A167 & A168;
  assign \new_[51645]_  = A169 & \new_[51644]_ ;
  assign \new_[51649]_  = ~A203 & ~A201;
  assign \new_[51650]_  = A166 & \new_[51649]_ ;
  assign \new_[51651]_  = \new_[51650]_  & \new_[51645]_ ;
  assign \new_[51655]_  = A269 & ~A268;
  assign \new_[51656]_  = A267 & \new_[51655]_ ;
  assign \new_[51659]_  = ~A299 & A298;
  assign \new_[51662]_  = ~A302 & A300;
  assign \new_[51663]_  = \new_[51662]_  & \new_[51659]_ ;
  assign \new_[51664]_  = \new_[51663]_  & \new_[51656]_ ;
  assign \new_[51668]_  = ~A167 & A168;
  assign \new_[51669]_  = A169 & \new_[51668]_ ;
  assign \new_[51673]_  = ~A203 & ~A201;
  assign \new_[51674]_  = A166 & \new_[51673]_ ;
  assign \new_[51675]_  = \new_[51674]_  & \new_[51669]_ ;
  assign \new_[51679]_  = A269 & ~A268;
  assign \new_[51680]_  = A267 & \new_[51679]_ ;
  assign \new_[51683]_  = A299 & ~A298;
  assign \new_[51686]_  = A301 & A300;
  assign \new_[51687]_  = \new_[51686]_  & \new_[51683]_ ;
  assign \new_[51688]_  = \new_[51687]_  & \new_[51680]_ ;
  assign \new_[51692]_  = ~A167 & A168;
  assign \new_[51693]_  = A169 & \new_[51692]_ ;
  assign \new_[51697]_  = ~A203 & ~A201;
  assign \new_[51698]_  = A166 & \new_[51697]_ ;
  assign \new_[51699]_  = \new_[51698]_  & \new_[51693]_ ;
  assign \new_[51703]_  = A269 & ~A268;
  assign \new_[51704]_  = A267 & \new_[51703]_ ;
  assign \new_[51707]_  = A299 & ~A298;
  assign \new_[51710]_  = ~A302 & A300;
  assign \new_[51711]_  = \new_[51710]_  & \new_[51707]_ ;
  assign \new_[51712]_  = \new_[51711]_  & \new_[51704]_ ;
  assign \new_[51716]_  = ~A167 & A168;
  assign \new_[51717]_  = A169 & \new_[51716]_ ;
  assign \new_[51721]_  = ~A203 & ~A201;
  assign \new_[51722]_  = A166 & \new_[51721]_ ;
  assign \new_[51723]_  = \new_[51722]_  & \new_[51717]_ ;
  assign \new_[51727]_  = A298 & A268;
  assign \new_[51728]_  = ~A267 & \new_[51727]_ ;
  assign \new_[51731]_  = ~A300 & ~A299;
  assign \new_[51734]_  = A302 & ~A301;
  assign \new_[51735]_  = \new_[51734]_  & \new_[51731]_ ;
  assign \new_[51736]_  = \new_[51735]_  & \new_[51728]_ ;
  assign \new_[51740]_  = ~A167 & A168;
  assign \new_[51741]_  = A169 & \new_[51740]_ ;
  assign \new_[51745]_  = ~A203 & ~A201;
  assign \new_[51746]_  = A166 & \new_[51745]_ ;
  assign \new_[51747]_  = \new_[51746]_  & \new_[51741]_ ;
  assign \new_[51751]_  = ~A298 & A268;
  assign \new_[51752]_  = ~A267 & \new_[51751]_ ;
  assign \new_[51755]_  = ~A300 & A299;
  assign \new_[51758]_  = A302 & ~A301;
  assign \new_[51759]_  = \new_[51758]_  & \new_[51755]_ ;
  assign \new_[51760]_  = \new_[51759]_  & \new_[51752]_ ;
  assign \new_[51764]_  = ~A167 & A168;
  assign \new_[51765]_  = A169 & \new_[51764]_ ;
  assign \new_[51769]_  = ~A203 & ~A201;
  assign \new_[51770]_  = A166 & \new_[51769]_ ;
  assign \new_[51771]_  = \new_[51770]_  & \new_[51765]_ ;
  assign \new_[51775]_  = A298 & ~A269;
  assign \new_[51776]_  = ~A267 & \new_[51775]_ ;
  assign \new_[51779]_  = ~A300 & ~A299;
  assign \new_[51782]_  = A302 & ~A301;
  assign \new_[51783]_  = \new_[51782]_  & \new_[51779]_ ;
  assign \new_[51784]_  = \new_[51783]_  & \new_[51776]_ ;
  assign \new_[51788]_  = ~A167 & A168;
  assign \new_[51789]_  = A169 & \new_[51788]_ ;
  assign \new_[51793]_  = ~A203 & ~A201;
  assign \new_[51794]_  = A166 & \new_[51793]_ ;
  assign \new_[51795]_  = \new_[51794]_  & \new_[51789]_ ;
  assign \new_[51799]_  = ~A298 & ~A269;
  assign \new_[51800]_  = ~A267 & \new_[51799]_ ;
  assign \new_[51803]_  = ~A300 & A299;
  assign \new_[51806]_  = A302 & ~A301;
  assign \new_[51807]_  = \new_[51806]_  & \new_[51803]_ ;
  assign \new_[51808]_  = \new_[51807]_  & \new_[51800]_ ;
  assign \new_[51812]_  = ~A167 & A168;
  assign \new_[51813]_  = A169 & \new_[51812]_ ;
  assign \new_[51817]_  = ~A203 & ~A201;
  assign \new_[51818]_  = A166 & \new_[51817]_ ;
  assign \new_[51819]_  = \new_[51818]_  & \new_[51813]_ ;
  assign \new_[51823]_  = A298 & A266;
  assign \new_[51824]_  = A265 & \new_[51823]_ ;
  assign \new_[51827]_  = ~A300 & ~A299;
  assign \new_[51830]_  = A302 & ~A301;
  assign \new_[51831]_  = \new_[51830]_  & \new_[51827]_ ;
  assign \new_[51832]_  = \new_[51831]_  & \new_[51824]_ ;
  assign \new_[51836]_  = ~A167 & A168;
  assign \new_[51837]_  = A169 & \new_[51836]_ ;
  assign \new_[51841]_  = ~A203 & ~A201;
  assign \new_[51842]_  = A166 & \new_[51841]_ ;
  assign \new_[51843]_  = \new_[51842]_  & \new_[51837]_ ;
  assign \new_[51847]_  = ~A298 & A266;
  assign \new_[51848]_  = A265 & \new_[51847]_ ;
  assign \new_[51851]_  = ~A300 & A299;
  assign \new_[51854]_  = A302 & ~A301;
  assign \new_[51855]_  = \new_[51854]_  & \new_[51851]_ ;
  assign \new_[51856]_  = \new_[51855]_  & \new_[51848]_ ;
  assign \new_[51860]_  = ~A167 & A168;
  assign \new_[51861]_  = A169 & \new_[51860]_ ;
  assign \new_[51865]_  = ~A203 & ~A201;
  assign \new_[51866]_  = A166 & \new_[51865]_ ;
  assign \new_[51867]_  = \new_[51866]_  & \new_[51861]_ ;
  assign \new_[51871]_  = A267 & A266;
  assign \new_[51872]_  = ~A265 & \new_[51871]_ ;
  assign \new_[51875]_  = A300 & A268;
  assign \new_[51878]_  = A302 & ~A301;
  assign \new_[51879]_  = \new_[51878]_  & \new_[51875]_ ;
  assign \new_[51880]_  = \new_[51879]_  & \new_[51872]_ ;
  assign \new_[51884]_  = ~A167 & A168;
  assign \new_[51885]_  = A169 & \new_[51884]_ ;
  assign \new_[51889]_  = ~A203 & ~A201;
  assign \new_[51890]_  = A166 & \new_[51889]_ ;
  assign \new_[51891]_  = \new_[51890]_  & \new_[51885]_ ;
  assign \new_[51895]_  = A267 & A266;
  assign \new_[51896]_  = ~A265 & \new_[51895]_ ;
  assign \new_[51899]_  = A300 & ~A269;
  assign \new_[51902]_  = A302 & ~A301;
  assign \new_[51903]_  = \new_[51902]_  & \new_[51899]_ ;
  assign \new_[51904]_  = \new_[51903]_  & \new_[51896]_ ;
  assign \new_[51908]_  = ~A167 & A168;
  assign \new_[51909]_  = A169 & \new_[51908]_ ;
  assign \new_[51913]_  = ~A203 & ~A201;
  assign \new_[51914]_  = A166 & \new_[51913]_ ;
  assign \new_[51915]_  = \new_[51914]_  & \new_[51909]_ ;
  assign \new_[51919]_  = ~A267 & A266;
  assign \new_[51920]_  = ~A265 & \new_[51919]_ ;
  assign \new_[51923]_  = A269 & ~A268;
  assign \new_[51926]_  = A301 & ~A300;
  assign \new_[51927]_  = \new_[51926]_  & \new_[51923]_ ;
  assign \new_[51928]_  = \new_[51927]_  & \new_[51920]_ ;
  assign \new_[51932]_  = ~A167 & A168;
  assign \new_[51933]_  = A169 & \new_[51932]_ ;
  assign \new_[51937]_  = ~A203 & ~A201;
  assign \new_[51938]_  = A166 & \new_[51937]_ ;
  assign \new_[51939]_  = \new_[51938]_  & \new_[51933]_ ;
  assign \new_[51943]_  = ~A267 & A266;
  assign \new_[51944]_  = ~A265 & \new_[51943]_ ;
  assign \new_[51947]_  = A269 & ~A268;
  assign \new_[51950]_  = ~A302 & ~A300;
  assign \new_[51951]_  = \new_[51950]_  & \new_[51947]_ ;
  assign \new_[51952]_  = \new_[51951]_  & \new_[51944]_ ;
  assign \new_[51956]_  = ~A167 & A168;
  assign \new_[51957]_  = A169 & \new_[51956]_ ;
  assign \new_[51961]_  = ~A203 & ~A201;
  assign \new_[51962]_  = A166 & \new_[51961]_ ;
  assign \new_[51963]_  = \new_[51962]_  & \new_[51957]_ ;
  assign \new_[51967]_  = ~A267 & A266;
  assign \new_[51968]_  = ~A265 & \new_[51967]_ ;
  assign \new_[51971]_  = A269 & ~A268;
  assign \new_[51974]_  = A299 & A298;
  assign \new_[51975]_  = \new_[51974]_  & \new_[51971]_ ;
  assign \new_[51976]_  = \new_[51975]_  & \new_[51968]_ ;
  assign \new_[51980]_  = ~A167 & A168;
  assign \new_[51981]_  = A169 & \new_[51980]_ ;
  assign \new_[51985]_  = ~A203 & ~A201;
  assign \new_[51986]_  = A166 & \new_[51985]_ ;
  assign \new_[51987]_  = \new_[51986]_  & \new_[51981]_ ;
  assign \new_[51991]_  = ~A267 & A266;
  assign \new_[51992]_  = ~A265 & \new_[51991]_ ;
  assign \new_[51995]_  = A269 & ~A268;
  assign \new_[51998]_  = ~A299 & ~A298;
  assign \new_[51999]_  = \new_[51998]_  & \new_[51995]_ ;
  assign \new_[52000]_  = \new_[51999]_  & \new_[51992]_ ;
  assign \new_[52004]_  = ~A167 & A168;
  assign \new_[52005]_  = A169 & \new_[52004]_ ;
  assign \new_[52009]_  = ~A203 & ~A201;
  assign \new_[52010]_  = A166 & \new_[52009]_ ;
  assign \new_[52011]_  = \new_[52010]_  & \new_[52005]_ ;
  assign \new_[52015]_  = A267 & ~A266;
  assign \new_[52016]_  = A265 & \new_[52015]_ ;
  assign \new_[52019]_  = A300 & A268;
  assign \new_[52022]_  = A302 & ~A301;
  assign \new_[52023]_  = \new_[52022]_  & \new_[52019]_ ;
  assign \new_[52024]_  = \new_[52023]_  & \new_[52016]_ ;
  assign \new_[52028]_  = ~A167 & A168;
  assign \new_[52029]_  = A169 & \new_[52028]_ ;
  assign \new_[52033]_  = ~A203 & ~A201;
  assign \new_[52034]_  = A166 & \new_[52033]_ ;
  assign \new_[52035]_  = \new_[52034]_  & \new_[52029]_ ;
  assign \new_[52039]_  = A267 & ~A266;
  assign \new_[52040]_  = A265 & \new_[52039]_ ;
  assign \new_[52043]_  = A300 & ~A269;
  assign \new_[52046]_  = A302 & ~A301;
  assign \new_[52047]_  = \new_[52046]_  & \new_[52043]_ ;
  assign \new_[52048]_  = \new_[52047]_  & \new_[52040]_ ;
  assign \new_[52052]_  = ~A167 & A168;
  assign \new_[52053]_  = A169 & \new_[52052]_ ;
  assign \new_[52057]_  = ~A203 & ~A201;
  assign \new_[52058]_  = A166 & \new_[52057]_ ;
  assign \new_[52059]_  = \new_[52058]_  & \new_[52053]_ ;
  assign \new_[52063]_  = ~A267 & ~A266;
  assign \new_[52064]_  = A265 & \new_[52063]_ ;
  assign \new_[52067]_  = A269 & ~A268;
  assign \new_[52070]_  = A301 & ~A300;
  assign \new_[52071]_  = \new_[52070]_  & \new_[52067]_ ;
  assign \new_[52072]_  = \new_[52071]_  & \new_[52064]_ ;
  assign \new_[52076]_  = ~A167 & A168;
  assign \new_[52077]_  = A169 & \new_[52076]_ ;
  assign \new_[52081]_  = ~A203 & ~A201;
  assign \new_[52082]_  = A166 & \new_[52081]_ ;
  assign \new_[52083]_  = \new_[52082]_  & \new_[52077]_ ;
  assign \new_[52087]_  = ~A267 & ~A266;
  assign \new_[52088]_  = A265 & \new_[52087]_ ;
  assign \new_[52091]_  = A269 & ~A268;
  assign \new_[52094]_  = ~A302 & ~A300;
  assign \new_[52095]_  = \new_[52094]_  & \new_[52091]_ ;
  assign \new_[52096]_  = \new_[52095]_  & \new_[52088]_ ;
  assign \new_[52100]_  = ~A167 & A168;
  assign \new_[52101]_  = A169 & \new_[52100]_ ;
  assign \new_[52105]_  = ~A203 & ~A201;
  assign \new_[52106]_  = A166 & \new_[52105]_ ;
  assign \new_[52107]_  = \new_[52106]_  & \new_[52101]_ ;
  assign \new_[52111]_  = ~A267 & ~A266;
  assign \new_[52112]_  = A265 & \new_[52111]_ ;
  assign \new_[52115]_  = A269 & ~A268;
  assign \new_[52118]_  = A299 & A298;
  assign \new_[52119]_  = \new_[52118]_  & \new_[52115]_ ;
  assign \new_[52120]_  = \new_[52119]_  & \new_[52112]_ ;
  assign \new_[52124]_  = ~A167 & A168;
  assign \new_[52125]_  = A169 & \new_[52124]_ ;
  assign \new_[52129]_  = ~A203 & ~A201;
  assign \new_[52130]_  = A166 & \new_[52129]_ ;
  assign \new_[52131]_  = \new_[52130]_  & \new_[52125]_ ;
  assign \new_[52135]_  = ~A267 & ~A266;
  assign \new_[52136]_  = A265 & \new_[52135]_ ;
  assign \new_[52139]_  = A269 & ~A268;
  assign \new_[52142]_  = ~A299 & ~A298;
  assign \new_[52143]_  = \new_[52142]_  & \new_[52139]_ ;
  assign \new_[52144]_  = \new_[52143]_  & \new_[52136]_ ;
  assign \new_[52148]_  = ~A167 & A168;
  assign \new_[52149]_  = A169 & \new_[52148]_ ;
  assign \new_[52153]_  = ~A203 & ~A201;
  assign \new_[52154]_  = A166 & \new_[52153]_ ;
  assign \new_[52155]_  = \new_[52154]_  & \new_[52149]_ ;
  assign \new_[52159]_  = A298 & ~A266;
  assign \new_[52160]_  = ~A265 & \new_[52159]_ ;
  assign \new_[52163]_  = ~A300 & ~A299;
  assign \new_[52166]_  = A302 & ~A301;
  assign \new_[52167]_  = \new_[52166]_  & \new_[52163]_ ;
  assign \new_[52168]_  = \new_[52167]_  & \new_[52160]_ ;
  assign \new_[52172]_  = ~A167 & A168;
  assign \new_[52173]_  = A169 & \new_[52172]_ ;
  assign \new_[52177]_  = ~A203 & ~A201;
  assign \new_[52178]_  = A166 & \new_[52177]_ ;
  assign \new_[52179]_  = \new_[52178]_  & \new_[52173]_ ;
  assign \new_[52183]_  = ~A298 & ~A266;
  assign \new_[52184]_  = ~A265 & \new_[52183]_ ;
  assign \new_[52187]_  = ~A300 & A299;
  assign \new_[52190]_  = A302 & ~A301;
  assign \new_[52191]_  = \new_[52190]_  & \new_[52187]_ ;
  assign \new_[52192]_  = \new_[52191]_  & \new_[52184]_ ;
  assign \new_[52196]_  = ~A167 & A168;
  assign \new_[52197]_  = A169 & \new_[52196]_ ;
  assign \new_[52201]_  = A200 & A199;
  assign \new_[52202]_  = A166 & \new_[52201]_ ;
  assign \new_[52203]_  = \new_[52202]_  & \new_[52197]_ ;
  assign \new_[52207]_  = A269 & ~A268;
  assign \new_[52208]_  = A267 & \new_[52207]_ ;
  assign \new_[52211]_  = ~A299 & A298;
  assign \new_[52214]_  = A301 & A300;
  assign \new_[52215]_  = \new_[52214]_  & \new_[52211]_ ;
  assign \new_[52216]_  = \new_[52215]_  & \new_[52208]_ ;
  assign \new_[52220]_  = ~A167 & A168;
  assign \new_[52221]_  = A169 & \new_[52220]_ ;
  assign \new_[52225]_  = A200 & A199;
  assign \new_[52226]_  = A166 & \new_[52225]_ ;
  assign \new_[52227]_  = \new_[52226]_  & \new_[52221]_ ;
  assign \new_[52231]_  = A269 & ~A268;
  assign \new_[52232]_  = A267 & \new_[52231]_ ;
  assign \new_[52235]_  = ~A299 & A298;
  assign \new_[52238]_  = ~A302 & A300;
  assign \new_[52239]_  = \new_[52238]_  & \new_[52235]_ ;
  assign \new_[52240]_  = \new_[52239]_  & \new_[52232]_ ;
  assign \new_[52244]_  = ~A167 & A168;
  assign \new_[52245]_  = A169 & \new_[52244]_ ;
  assign \new_[52249]_  = A200 & A199;
  assign \new_[52250]_  = A166 & \new_[52249]_ ;
  assign \new_[52251]_  = \new_[52250]_  & \new_[52245]_ ;
  assign \new_[52255]_  = A269 & ~A268;
  assign \new_[52256]_  = A267 & \new_[52255]_ ;
  assign \new_[52259]_  = A299 & ~A298;
  assign \new_[52262]_  = A301 & A300;
  assign \new_[52263]_  = \new_[52262]_  & \new_[52259]_ ;
  assign \new_[52264]_  = \new_[52263]_  & \new_[52256]_ ;
  assign \new_[52268]_  = ~A167 & A168;
  assign \new_[52269]_  = A169 & \new_[52268]_ ;
  assign \new_[52273]_  = A200 & A199;
  assign \new_[52274]_  = A166 & \new_[52273]_ ;
  assign \new_[52275]_  = \new_[52274]_  & \new_[52269]_ ;
  assign \new_[52279]_  = A269 & ~A268;
  assign \new_[52280]_  = A267 & \new_[52279]_ ;
  assign \new_[52283]_  = A299 & ~A298;
  assign \new_[52286]_  = ~A302 & A300;
  assign \new_[52287]_  = \new_[52286]_  & \new_[52283]_ ;
  assign \new_[52288]_  = \new_[52287]_  & \new_[52280]_ ;
  assign \new_[52292]_  = ~A167 & A168;
  assign \new_[52293]_  = A169 & \new_[52292]_ ;
  assign \new_[52297]_  = A200 & A199;
  assign \new_[52298]_  = A166 & \new_[52297]_ ;
  assign \new_[52299]_  = \new_[52298]_  & \new_[52293]_ ;
  assign \new_[52303]_  = A298 & A268;
  assign \new_[52304]_  = ~A267 & \new_[52303]_ ;
  assign \new_[52307]_  = ~A300 & ~A299;
  assign \new_[52310]_  = A302 & ~A301;
  assign \new_[52311]_  = \new_[52310]_  & \new_[52307]_ ;
  assign \new_[52312]_  = \new_[52311]_  & \new_[52304]_ ;
  assign \new_[52316]_  = ~A167 & A168;
  assign \new_[52317]_  = A169 & \new_[52316]_ ;
  assign \new_[52321]_  = A200 & A199;
  assign \new_[52322]_  = A166 & \new_[52321]_ ;
  assign \new_[52323]_  = \new_[52322]_  & \new_[52317]_ ;
  assign \new_[52327]_  = ~A298 & A268;
  assign \new_[52328]_  = ~A267 & \new_[52327]_ ;
  assign \new_[52331]_  = ~A300 & A299;
  assign \new_[52334]_  = A302 & ~A301;
  assign \new_[52335]_  = \new_[52334]_  & \new_[52331]_ ;
  assign \new_[52336]_  = \new_[52335]_  & \new_[52328]_ ;
  assign \new_[52340]_  = ~A167 & A168;
  assign \new_[52341]_  = A169 & \new_[52340]_ ;
  assign \new_[52345]_  = A200 & A199;
  assign \new_[52346]_  = A166 & \new_[52345]_ ;
  assign \new_[52347]_  = \new_[52346]_  & \new_[52341]_ ;
  assign \new_[52351]_  = A298 & ~A269;
  assign \new_[52352]_  = ~A267 & \new_[52351]_ ;
  assign \new_[52355]_  = ~A300 & ~A299;
  assign \new_[52358]_  = A302 & ~A301;
  assign \new_[52359]_  = \new_[52358]_  & \new_[52355]_ ;
  assign \new_[52360]_  = \new_[52359]_  & \new_[52352]_ ;
  assign \new_[52364]_  = ~A167 & A168;
  assign \new_[52365]_  = A169 & \new_[52364]_ ;
  assign \new_[52369]_  = A200 & A199;
  assign \new_[52370]_  = A166 & \new_[52369]_ ;
  assign \new_[52371]_  = \new_[52370]_  & \new_[52365]_ ;
  assign \new_[52375]_  = ~A298 & ~A269;
  assign \new_[52376]_  = ~A267 & \new_[52375]_ ;
  assign \new_[52379]_  = ~A300 & A299;
  assign \new_[52382]_  = A302 & ~A301;
  assign \new_[52383]_  = \new_[52382]_  & \new_[52379]_ ;
  assign \new_[52384]_  = \new_[52383]_  & \new_[52376]_ ;
  assign \new_[52388]_  = ~A167 & A168;
  assign \new_[52389]_  = A169 & \new_[52388]_ ;
  assign \new_[52393]_  = A200 & A199;
  assign \new_[52394]_  = A166 & \new_[52393]_ ;
  assign \new_[52395]_  = \new_[52394]_  & \new_[52389]_ ;
  assign \new_[52399]_  = A298 & A266;
  assign \new_[52400]_  = A265 & \new_[52399]_ ;
  assign \new_[52403]_  = ~A300 & ~A299;
  assign \new_[52406]_  = A302 & ~A301;
  assign \new_[52407]_  = \new_[52406]_  & \new_[52403]_ ;
  assign \new_[52408]_  = \new_[52407]_  & \new_[52400]_ ;
  assign \new_[52412]_  = ~A167 & A168;
  assign \new_[52413]_  = A169 & \new_[52412]_ ;
  assign \new_[52417]_  = A200 & A199;
  assign \new_[52418]_  = A166 & \new_[52417]_ ;
  assign \new_[52419]_  = \new_[52418]_  & \new_[52413]_ ;
  assign \new_[52423]_  = ~A298 & A266;
  assign \new_[52424]_  = A265 & \new_[52423]_ ;
  assign \new_[52427]_  = ~A300 & A299;
  assign \new_[52430]_  = A302 & ~A301;
  assign \new_[52431]_  = \new_[52430]_  & \new_[52427]_ ;
  assign \new_[52432]_  = \new_[52431]_  & \new_[52424]_ ;
  assign \new_[52436]_  = ~A167 & A168;
  assign \new_[52437]_  = A169 & \new_[52436]_ ;
  assign \new_[52441]_  = A200 & A199;
  assign \new_[52442]_  = A166 & \new_[52441]_ ;
  assign \new_[52443]_  = \new_[52442]_  & \new_[52437]_ ;
  assign \new_[52447]_  = A267 & A266;
  assign \new_[52448]_  = ~A265 & \new_[52447]_ ;
  assign \new_[52451]_  = A300 & A268;
  assign \new_[52454]_  = A302 & ~A301;
  assign \new_[52455]_  = \new_[52454]_  & \new_[52451]_ ;
  assign \new_[52456]_  = \new_[52455]_  & \new_[52448]_ ;
  assign \new_[52460]_  = ~A167 & A168;
  assign \new_[52461]_  = A169 & \new_[52460]_ ;
  assign \new_[52465]_  = A200 & A199;
  assign \new_[52466]_  = A166 & \new_[52465]_ ;
  assign \new_[52467]_  = \new_[52466]_  & \new_[52461]_ ;
  assign \new_[52471]_  = A267 & A266;
  assign \new_[52472]_  = ~A265 & \new_[52471]_ ;
  assign \new_[52475]_  = A300 & ~A269;
  assign \new_[52478]_  = A302 & ~A301;
  assign \new_[52479]_  = \new_[52478]_  & \new_[52475]_ ;
  assign \new_[52480]_  = \new_[52479]_  & \new_[52472]_ ;
  assign \new_[52484]_  = ~A167 & A168;
  assign \new_[52485]_  = A169 & \new_[52484]_ ;
  assign \new_[52489]_  = A200 & A199;
  assign \new_[52490]_  = A166 & \new_[52489]_ ;
  assign \new_[52491]_  = \new_[52490]_  & \new_[52485]_ ;
  assign \new_[52495]_  = ~A267 & A266;
  assign \new_[52496]_  = ~A265 & \new_[52495]_ ;
  assign \new_[52499]_  = A269 & ~A268;
  assign \new_[52502]_  = A301 & ~A300;
  assign \new_[52503]_  = \new_[52502]_  & \new_[52499]_ ;
  assign \new_[52504]_  = \new_[52503]_  & \new_[52496]_ ;
  assign \new_[52508]_  = ~A167 & A168;
  assign \new_[52509]_  = A169 & \new_[52508]_ ;
  assign \new_[52513]_  = A200 & A199;
  assign \new_[52514]_  = A166 & \new_[52513]_ ;
  assign \new_[52515]_  = \new_[52514]_  & \new_[52509]_ ;
  assign \new_[52519]_  = ~A267 & A266;
  assign \new_[52520]_  = ~A265 & \new_[52519]_ ;
  assign \new_[52523]_  = A269 & ~A268;
  assign \new_[52526]_  = ~A302 & ~A300;
  assign \new_[52527]_  = \new_[52526]_  & \new_[52523]_ ;
  assign \new_[52528]_  = \new_[52527]_  & \new_[52520]_ ;
  assign \new_[52532]_  = ~A167 & A168;
  assign \new_[52533]_  = A169 & \new_[52532]_ ;
  assign \new_[52537]_  = A200 & A199;
  assign \new_[52538]_  = A166 & \new_[52537]_ ;
  assign \new_[52539]_  = \new_[52538]_  & \new_[52533]_ ;
  assign \new_[52543]_  = ~A267 & A266;
  assign \new_[52544]_  = ~A265 & \new_[52543]_ ;
  assign \new_[52547]_  = A269 & ~A268;
  assign \new_[52550]_  = A299 & A298;
  assign \new_[52551]_  = \new_[52550]_  & \new_[52547]_ ;
  assign \new_[52552]_  = \new_[52551]_  & \new_[52544]_ ;
  assign \new_[52556]_  = ~A167 & A168;
  assign \new_[52557]_  = A169 & \new_[52556]_ ;
  assign \new_[52561]_  = A200 & A199;
  assign \new_[52562]_  = A166 & \new_[52561]_ ;
  assign \new_[52563]_  = \new_[52562]_  & \new_[52557]_ ;
  assign \new_[52567]_  = ~A267 & A266;
  assign \new_[52568]_  = ~A265 & \new_[52567]_ ;
  assign \new_[52571]_  = A269 & ~A268;
  assign \new_[52574]_  = ~A299 & ~A298;
  assign \new_[52575]_  = \new_[52574]_  & \new_[52571]_ ;
  assign \new_[52576]_  = \new_[52575]_  & \new_[52568]_ ;
  assign \new_[52580]_  = ~A167 & A168;
  assign \new_[52581]_  = A169 & \new_[52580]_ ;
  assign \new_[52585]_  = A200 & A199;
  assign \new_[52586]_  = A166 & \new_[52585]_ ;
  assign \new_[52587]_  = \new_[52586]_  & \new_[52581]_ ;
  assign \new_[52591]_  = A267 & ~A266;
  assign \new_[52592]_  = A265 & \new_[52591]_ ;
  assign \new_[52595]_  = A300 & A268;
  assign \new_[52598]_  = A302 & ~A301;
  assign \new_[52599]_  = \new_[52598]_  & \new_[52595]_ ;
  assign \new_[52600]_  = \new_[52599]_  & \new_[52592]_ ;
  assign \new_[52604]_  = ~A167 & A168;
  assign \new_[52605]_  = A169 & \new_[52604]_ ;
  assign \new_[52609]_  = A200 & A199;
  assign \new_[52610]_  = A166 & \new_[52609]_ ;
  assign \new_[52611]_  = \new_[52610]_  & \new_[52605]_ ;
  assign \new_[52615]_  = A267 & ~A266;
  assign \new_[52616]_  = A265 & \new_[52615]_ ;
  assign \new_[52619]_  = A300 & ~A269;
  assign \new_[52622]_  = A302 & ~A301;
  assign \new_[52623]_  = \new_[52622]_  & \new_[52619]_ ;
  assign \new_[52624]_  = \new_[52623]_  & \new_[52616]_ ;
  assign \new_[52628]_  = ~A167 & A168;
  assign \new_[52629]_  = A169 & \new_[52628]_ ;
  assign \new_[52633]_  = A200 & A199;
  assign \new_[52634]_  = A166 & \new_[52633]_ ;
  assign \new_[52635]_  = \new_[52634]_  & \new_[52629]_ ;
  assign \new_[52639]_  = ~A267 & ~A266;
  assign \new_[52640]_  = A265 & \new_[52639]_ ;
  assign \new_[52643]_  = A269 & ~A268;
  assign \new_[52646]_  = A301 & ~A300;
  assign \new_[52647]_  = \new_[52646]_  & \new_[52643]_ ;
  assign \new_[52648]_  = \new_[52647]_  & \new_[52640]_ ;
  assign \new_[52652]_  = ~A167 & A168;
  assign \new_[52653]_  = A169 & \new_[52652]_ ;
  assign \new_[52657]_  = A200 & A199;
  assign \new_[52658]_  = A166 & \new_[52657]_ ;
  assign \new_[52659]_  = \new_[52658]_  & \new_[52653]_ ;
  assign \new_[52663]_  = ~A267 & ~A266;
  assign \new_[52664]_  = A265 & \new_[52663]_ ;
  assign \new_[52667]_  = A269 & ~A268;
  assign \new_[52670]_  = ~A302 & ~A300;
  assign \new_[52671]_  = \new_[52670]_  & \new_[52667]_ ;
  assign \new_[52672]_  = \new_[52671]_  & \new_[52664]_ ;
  assign \new_[52676]_  = ~A167 & A168;
  assign \new_[52677]_  = A169 & \new_[52676]_ ;
  assign \new_[52681]_  = A200 & A199;
  assign \new_[52682]_  = A166 & \new_[52681]_ ;
  assign \new_[52683]_  = \new_[52682]_  & \new_[52677]_ ;
  assign \new_[52687]_  = ~A267 & ~A266;
  assign \new_[52688]_  = A265 & \new_[52687]_ ;
  assign \new_[52691]_  = A269 & ~A268;
  assign \new_[52694]_  = A299 & A298;
  assign \new_[52695]_  = \new_[52694]_  & \new_[52691]_ ;
  assign \new_[52696]_  = \new_[52695]_  & \new_[52688]_ ;
  assign \new_[52700]_  = ~A167 & A168;
  assign \new_[52701]_  = A169 & \new_[52700]_ ;
  assign \new_[52705]_  = A200 & A199;
  assign \new_[52706]_  = A166 & \new_[52705]_ ;
  assign \new_[52707]_  = \new_[52706]_  & \new_[52701]_ ;
  assign \new_[52711]_  = ~A267 & ~A266;
  assign \new_[52712]_  = A265 & \new_[52711]_ ;
  assign \new_[52715]_  = A269 & ~A268;
  assign \new_[52718]_  = ~A299 & ~A298;
  assign \new_[52719]_  = \new_[52718]_  & \new_[52715]_ ;
  assign \new_[52720]_  = \new_[52719]_  & \new_[52712]_ ;
  assign \new_[52724]_  = ~A167 & A168;
  assign \new_[52725]_  = A169 & \new_[52724]_ ;
  assign \new_[52729]_  = A200 & A199;
  assign \new_[52730]_  = A166 & \new_[52729]_ ;
  assign \new_[52731]_  = \new_[52730]_  & \new_[52725]_ ;
  assign \new_[52735]_  = A298 & ~A266;
  assign \new_[52736]_  = ~A265 & \new_[52735]_ ;
  assign \new_[52739]_  = ~A300 & ~A299;
  assign \new_[52742]_  = A302 & ~A301;
  assign \new_[52743]_  = \new_[52742]_  & \new_[52739]_ ;
  assign \new_[52744]_  = \new_[52743]_  & \new_[52736]_ ;
  assign \new_[52748]_  = ~A167 & A168;
  assign \new_[52749]_  = A169 & \new_[52748]_ ;
  assign \new_[52753]_  = A200 & A199;
  assign \new_[52754]_  = A166 & \new_[52753]_ ;
  assign \new_[52755]_  = \new_[52754]_  & \new_[52749]_ ;
  assign \new_[52759]_  = ~A298 & ~A266;
  assign \new_[52760]_  = ~A265 & \new_[52759]_ ;
  assign \new_[52763]_  = ~A300 & A299;
  assign \new_[52766]_  = A302 & ~A301;
  assign \new_[52767]_  = \new_[52766]_  & \new_[52763]_ ;
  assign \new_[52768]_  = \new_[52767]_  & \new_[52760]_ ;
  assign \new_[52772]_  = ~A167 & A168;
  assign \new_[52773]_  = A169 & \new_[52772]_ ;
  assign \new_[52777]_  = ~A200 & ~A199;
  assign \new_[52778]_  = A166 & \new_[52777]_ ;
  assign \new_[52779]_  = \new_[52778]_  & \new_[52773]_ ;
  assign \new_[52783]_  = A269 & ~A268;
  assign \new_[52784]_  = A267 & \new_[52783]_ ;
  assign \new_[52787]_  = ~A299 & A298;
  assign \new_[52790]_  = A301 & A300;
  assign \new_[52791]_  = \new_[52790]_  & \new_[52787]_ ;
  assign \new_[52792]_  = \new_[52791]_  & \new_[52784]_ ;
  assign \new_[52796]_  = ~A167 & A168;
  assign \new_[52797]_  = A169 & \new_[52796]_ ;
  assign \new_[52801]_  = ~A200 & ~A199;
  assign \new_[52802]_  = A166 & \new_[52801]_ ;
  assign \new_[52803]_  = \new_[52802]_  & \new_[52797]_ ;
  assign \new_[52807]_  = A269 & ~A268;
  assign \new_[52808]_  = A267 & \new_[52807]_ ;
  assign \new_[52811]_  = ~A299 & A298;
  assign \new_[52814]_  = ~A302 & A300;
  assign \new_[52815]_  = \new_[52814]_  & \new_[52811]_ ;
  assign \new_[52816]_  = \new_[52815]_  & \new_[52808]_ ;
  assign \new_[52820]_  = ~A167 & A168;
  assign \new_[52821]_  = A169 & \new_[52820]_ ;
  assign \new_[52825]_  = ~A200 & ~A199;
  assign \new_[52826]_  = A166 & \new_[52825]_ ;
  assign \new_[52827]_  = \new_[52826]_  & \new_[52821]_ ;
  assign \new_[52831]_  = A269 & ~A268;
  assign \new_[52832]_  = A267 & \new_[52831]_ ;
  assign \new_[52835]_  = A299 & ~A298;
  assign \new_[52838]_  = A301 & A300;
  assign \new_[52839]_  = \new_[52838]_  & \new_[52835]_ ;
  assign \new_[52840]_  = \new_[52839]_  & \new_[52832]_ ;
  assign \new_[52844]_  = ~A167 & A168;
  assign \new_[52845]_  = A169 & \new_[52844]_ ;
  assign \new_[52849]_  = ~A200 & ~A199;
  assign \new_[52850]_  = A166 & \new_[52849]_ ;
  assign \new_[52851]_  = \new_[52850]_  & \new_[52845]_ ;
  assign \new_[52855]_  = A269 & ~A268;
  assign \new_[52856]_  = A267 & \new_[52855]_ ;
  assign \new_[52859]_  = A299 & ~A298;
  assign \new_[52862]_  = ~A302 & A300;
  assign \new_[52863]_  = \new_[52862]_  & \new_[52859]_ ;
  assign \new_[52864]_  = \new_[52863]_  & \new_[52856]_ ;
  assign \new_[52868]_  = ~A167 & A168;
  assign \new_[52869]_  = A169 & \new_[52868]_ ;
  assign \new_[52873]_  = ~A200 & ~A199;
  assign \new_[52874]_  = A166 & \new_[52873]_ ;
  assign \new_[52875]_  = \new_[52874]_  & \new_[52869]_ ;
  assign \new_[52879]_  = A298 & A268;
  assign \new_[52880]_  = ~A267 & \new_[52879]_ ;
  assign \new_[52883]_  = ~A300 & ~A299;
  assign \new_[52886]_  = A302 & ~A301;
  assign \new_[52887]_  = \new_[52886]_  & \new_[52883]_ ;
  assign \new_[52888]_  = \new_[52887]_  & \new_[52880]_ ;
  assign \new_[52892]_  = ~A167 & A168;
  assign \new_[52893]_  = A169 & \new_[52892]_ ;
  assign \new_[52897]_  = ~A200 & ~A199;
  assign \new_[52898]_  = A166 & \new_[52897]_ ;
  assign \new_[52899]_  = \new_[52898]_  & \new_[52893]_ ;
  assign \new_[52903]_  = ~A298 & A268;
  assign \new_[52904]_  = ~A267 & \new_[52903]_ ;
  assign \new_[52907]_  = ~A300 & A299;
  assign \new_[52910]_  = A302 & ~A301;
  assign \new_[52911]_  = \new_[52910]_  & \new_[52907]_ ;
  assign \new_[52912]_  = \new_[52911]_  & \new_[52904]_ ;
  assign \new_[52916]_  = ~A167 & A168;
  assign \new_[52917]_  = A169 & \new_[52916]_ ;
  assign \new_[52921]_  = ~A200 & ~A199;
  assign \new_[52922]_  = A166 & \new_[52921]_ ;
  assign \new_[52923]_  = \new_[52922]_  & \new_[52917]_ ;
  assign \new_[52927]_  = A298 & ~A269;
  assign \new_[52928]_  = ~A267 & \new_[52927]_ ;
  assign \new_[52931]_  = ~A300 & ~A299;
  assign \new_[52934]_  = A302 & ~A301;
  assign \new_[52935]_  = \new_[52934]_  & \new_[52931]_ ;
  assign \new_[52936]_  = \new_[52935]_  & \new_[52928]_ ;
  assign \new_[52940]_  = ~A167 & A168;
  assign \new_[52941]_  = A169 & \new_[52940]_ ;
  assign \new_[52945]_  = ~A200 & ~A199;
  assign \new_[52946]_  = A166 & \new_[52945]_ ;
  assign \new_[52947]_  = \new_[52946]_  & \new_[52941]_ ;
  assign \new_[52951]_  = ~A298 & ~A269;
  assign \new_[52952]_  = ~A267 & \new_[52951]_ ;
  assign \new_[52955]_  = ~A300 & A299;
  assign \new_[52958]_  = A302 & ~A301;
  assign \new_[52959]_  = \new_[52958]_  & \new_[52955]_ ;
  assign \new_[52960]_  = \new_[52959]_  & \new_[52952]_ ;
  assign \new_[52964]_  = ~A167 & A168;
  assign \new_[52965]_  = A169 & \new_[52964]_ ;
  assign \new_[52969]_  = ~A200 & ~A199;
  assign \new_[52970]_  = A166 & \new_[52969]_ ;
  assign \new_[52971]_  = \new_[52970]_  & \new_[52965]_ ;
  assign \new_[52975]_  = A298 & A266;
  assign \new_[52976]_  = A265 & \new_[52975]_ ;
  assign \new_[52979]_  = ~A300 & ~A299;
  assign \new_[52982]_  = A302 & ~A301;
  assign \new_[52983]_  = \new_[52982]_  & \new_[52979]_ ;
  assign \new_[52984]_  = \new_[52983]_  & \new_[52976]_ ;
  assign \new_[52988]_  = ~A167 & A168;
  assign \new_[52989]_  = A169 & \new_[52988]_ ;
  assign \new_[52993]_  = ~A200 & ~A199;
  assign \new_[52994]_  = A166 & \new_[52993]_ ;
  assign \new_[52995]_  = \new_[52994]_  & \new_[52989]_ ;
  assign \new_[52999]_  = ~A298 & A266;
  assign \new_[53000]_  = A265 & \new_[52999]_ ;
  assign \new_[53003]_  = ~A300 & A299;
  assign \new_[53006]_  = A302 & ~A301;
  assign \new_[53007]_  = \new_[53006]_  & \new_[53003]_ ;
  assign \new_[53008]_  = \new_[53007]_  & \new_[53000]_ ;
  assign \new_[53012]_  = ~A167 & A168;
  assign \new_[53013]_  = A169 & \new_[53012]_ ;
  assign \new_[53017]_  = ~A200 & ~A199;
  assign \new_[53018]_  = A166 & \new_[53017]_ ;
  assign \new_[53019]_  = \new_[53018]_  & \new_[53013]_ ;
  assign \new_[53023]_  = A267 & A266;
  assign \new_[53024]_  = ~A265 & \new_[53023]_ ;
  assign \new_[53027]_  = A300 & A268;
  assign \new_[53030]_  = A302 & ~A301;
  assign \new_[53031]_  = \new_[53030]_  & \new_[53027]_ ;
  assign \new_[53032]_  = \new_[53031]_  & \new_[53024]_ ;
  assign \new_[53036]_  = ~A167 & A168;
  assign \new_[53037]_  = A169 & \new_[53036]_ ;
  assign \new_[53041]_  = ~A200 & ~A199;
  assign \new_[53042]_  = A166 & \new_[53041]_ ;
  assign \new_[53043]_  = \new_[53042]_  & \new_[53037]_ ;
  assign \new_[53047]_  = A267 & A266;
  assign \new_[53048]_  = ~A265 & \new_[53047]_ ;
  assign \new_[53051]_  = A300 & ~A269;
  assign \new_[53054]_  = A302 & ~A301;
  assign \new_[53055]_  = \new_[53054]_  & \new_[53051]_ ;
  assign \new_[53056]_  = \new_[53055]_  & \new_[53048]_ ;
  assign \new_[53060]_  = ~A167 & A168;
  assign \new_[53061]_  = A169 & \new_[53060]_ ;
  assign \new_[53065]_  = ~A200 & ~A199;
  assign \new_[53066]_  = A166 & \new_[53065]_ ;
  assign \new_[53067]_  = \new_[53066]_  & \new_[53061]_ ;
  assign \new_[53071]_  = ~A267 & A266;
  assign \new_[53072]_  = ~A265 & \new_[53071]_ ;
  assign \new_[53075]_  = A269 & ~A268;
  assign \new_[53078]_  = A301 & ~A300;
  assign \new_[53079]_  = \new_[53078]_  & \new_[53075]_ ;
  assign \new_[53080]_  = \new_[53079]_  & \new_[53072]_ ;
  assign \new_[53084]_  = ~A167 & A168;
  assign \new_[53085]_  = A169 & \new_[53084]_ ;
  assign \new_[53089]_  = ~A200 & ~A199;
  assign \new_[53090]_  = A166 & \new_[53089]_ ;
  assign \new_[53091]_  = \new_[53090]_  & \new_[53085]_ ;
  assign \new_[53095]_  = ~A267 & A266;
  assign \new_[53096]_  = ~A265 & \new_[53095]_ ;
  assign \new_[53099]_  = A269 & ~A268;
  assign \new_[53102]_  = ~A302 & ~A300;
  assign \new_[53103]_  = \new_[53102]_  & \new_[53099]_ ;
  assign \new_[53104]_  = \new_[53103]_  & \new_[53096]_ ;
  assign \new_[53108]_  = ~A167 & A168;
  assign \new_[53109]_  = A169 & \new_[53108]_ ;
  assign \new_[53113]_  = ~A200 & ~A199;
  assign \new_[53114]_  = A166 & \new_[53113]_ ;
  assign \new_[53115]_  = \new_[53114]_  & \new_[53109]_ ;
  assign \new_[53119]_  = ~A267 & A266;
  assign \new_[53120]_  = ~A265 & \new_[53119]_ ;
  assign \new_[53123]_  = A269 & ~A268;
  assign \new_[53126]_  = A299 & A298;
  assign \new_[53127]_  = \new_[53126]_  & \new_[53123]_ ;
  assign \new_[53128]_  = \new_[53127]_  & \new_[53120]_ ;
  assign \new_[53132]_  = ~A167 & A168;
  assign \new_[53133]_  = A169 & \new_[53132]_ ;
  assign \new_[53137]_  = ~A200 & ~A199;
  assign \new_[53138]_  = A166 & \new_[53137]_ ;
  assign \new_[53139]_  = \new_[53138]_  & \new_[53133]_ ;
  assign \new_[53143]_  = ~A267 & A266;
  assign \new_[53144]_  = ~A265 & \new_[53143]_ ;
  assign \new_[53147]_  = A269 & ~A268;
  assign \new_[53150]_  = ~A299 & ~A298;
  assign \new_[53151]_  = \new_[53150]_  & \new_[53147]_ ;
  assign \new_[53152]_  = \new_[53151]_  & \new_[53144]_ ;
  assign \new_[53156]_  = ~A167 & A168;
  assign \new_[53157]_  = A169 & \new_[53156]_ ;
  assign \new_[53161]_  = ~A200 & ~A199;
  assign \new_[53162]_  = A166 & \new_[53161]_ ;
  assign \new_[53163]_  = \new_[53162]_  & \new_[53157]_ ;
  assign \new_[53167]_  = A267 & ~A266;
  assign \new_[53168]_  = A265 & \new_[53167]_ ;
  assign \new_[53171]_  = A300 & A268;
  assign \new_[53174]_  = A302 & ~A301;
  assign \new_[53175]_  = \new_[53174]_  & \new_[53171]_ ;
  assign \new_[53176]_  = \new_[53175]_  & \new_[53168]_ ;
  assign \new_[53180]_  = ~A167 & A168;
  assign \new_[53181]_  = A169 & \new_[53180]_ ;
  assign \new_[53185]_  = ~A200 & ~A199;
  assign \new_[53186]_  = A166 & \new_[53185]_ ;
  assign \new_[53187]_  = \new_[53186]_  & \new_[53181]_ ;
  assign \new_[53191]_  = A267 & ~A266;
  assign \new_[53192]_  = A265 & \new_[53191]_ ;
  assign \new_[53195]_  = A300 & ~A269;
  assign \new_[53198]_  = A302 & ~A301;
  assign \new_[53199]_  = \new_[53198]_  & \new_[53195]_ ;
  assign \new_[53200]_  = \new_[53199]_  & \new_[53192]_ ;
  assign \new_[53204]_  = ~A167 & A168;
  assign \new_[53205]_  = A169 & \new_[53204]_ ;
  assign \new_[53209]_  = ~A200 & ~A199;
  assign \new_[53210]_  = A166 & \new_[53209]_ ;
  assign \new_[53211]_  = \new_[53210]_  & \new_[53205]_ ;
  assign \new_[53215]_  = ~A267 & ~A266;
  assign \new_[53216]_  = A265 & \new_[53215]_ ;
  assign \new_[53219]_  = A269 & ~A268;
  assign \new_[53222]_  = A301 & ~A300;
  assign \new_[53223]_  = \new_[53222]_  & \new_[53219]_ ;
  assign \new_[53224]_  = \new_[53223]_  & \new_[53216]_ ;
  assign \new_[53228]_  = ~A167 & A168;
  assign \new_[53229]_  = A169 & \new_[53228]_ ;
  assign \new_[53233]_  = ~A200 & ~A199;
  assign \new_[53234]_  = A166 & \new_[53233]_ ;
  assign \new_[53235]_  = \new_[53234]_  & \new_[53229]_ ;
  assign \new_[53239]_  = ~A267 & ~A266;
  assign \new_[53240]_  = A265 & \new_[53239]_ ;
  assign \new_[53243]_  = A269 & ~A268;
  assign \new_[53246]_  = ~A302 & ~A300;
  assign \new_[53247]_  = \new_[53246]_  & \new_[53243]_ ;
  assign \new_[53248]_  = \new_[53247]_  & \new_[53240]_ ;
  assign \new_[53252]_  = ~A167 & A168;
  assign \new_[53253]_  = A169 & \new_[53252]_ ;
  assign \new_[53257]_  = ~A200 & ~A199;
  assign \new_[53258]_  = A166 & \new_[53257]_ ;
  assign \new_[53259]_  = \new_[53258]_  & \new_[53253]_ ;
  assign \new_[53263]_  = ~A267 & ~A266;
  assign \new_[53264]_  = A265 & \new_[53263]_ ;
  assign \new_[53267]_  = A269 & ~A268;
  assign \new_[53270]_  = A299 & A298;
  assign \new_[53271]_  = \new_[53270]_  & \new_[53267]_ ;
  assign \new_[53272]_  = \new_[53271]_  & \new_[53264]_ ;
  assign \new_[53276]_  = ~A167 & A168;
  assign \new_[53277]_  = A169 & \new_[53276]_ ;
  assign \new_[53281]_  = ~A200 & ~A199;
  assign \new_[53282]_  = A166 & \new_[53281]_ ;
  assign \new_[53283]_  = \new_[53282]_  & \new_[53277]_ ;
  assign \new_[53287]_  = ~A267 & ~A266;
  assign \new_[53288]_  = A265 & \new_[53287]_ ;
  assign \new_[53291]_  = A269 & ~A268;
  assign \new_[53294]_  = ~A299 & ~A298;
  assign \new_[53295]_  = \new_[53294]_  & \new_[53291]_ ;
  assign \new_[53296]_  = \new_[53295]_  & \new_[53288]_ ;
  assign \new_[53300]_  = ~A167 & A168;
  assign \new_[53301]_  = A169 & \new_[53300]_ ;
  assign \new_[53305]_  = ~A200 & ~A199;
  assign \new_[53306]_  = A166 & \new_[53305]_ ;
  assign \new_[53307]_  = \new_[53306]_  & \new_[53301]_ ;
  assign \new_[53311]_  = A298 & ~A266;
  assign \new_[53312]_  = ~A265 & \new_[53311]_ ;
  assign \new_[53315]_  = ~A300 & ~A299;
  assign \new_[53318]_  = A302 & ~A301;
  assign \new_[53319]_  = \new_[53318]_  & \new_[53315]_ ;
  assign \new_[53320]_  = \new_[53319]_  & \new_[53312]_ ;
  assign \new_[53324]_  = ~A167 & A168;
  assign \new_[53325]_  = A169 & \new_[53324]_ ;
  assign \new_[53329]_  = ~A200 & ~A199;
  assign \new_[53330]_  = A166 & \new_[53329]_ ;
  assign \new_[53331]_  = \new_[53330]_  & \new_[53325]_ ;
  assign \new_[53335]_  = ~A298 & ~A266;
  assign \new_[53336]_  = ~A265 & \new_[53335]_ ;
  assign \new_[53339]_  = ~A300 & A299;
  assign \new_[53342]_  = A302 & ~A301;
  assign \new_[53343]_  = \new_[53342]_  & \new_[53339]_ ;
  assign \new_[53344]_  = \new_[53343]_  & \new_[53336]_ ;
  assign \new_[53348]_  = ~A199 & ~A168;
  assign \new_[53349]_  = A169 & \new_[53348]_ ;
  assign \new_[53353]_  = ~A202 & ~A201;
  assign \new_[53354]_  = A200 & \new_[53353]_ ;
  assign \new_[53355]_  = \new_[53354]_  & \new_[53349]_ ;
  assign \new_[53359]_  = ~A268 & A267;
  assign \new_[53360]_  = A203 & \new_[53359]_ ;
  assign \new_[53363]_  = A300 & A269;
  assign \new_[53366]_  = A302 & ~A301;
  assign \new_[53367]_  = \new_[53366]_  & \new_[53363]_ ;
  assign \new_[53368]_  = \new_[53367]_  & \new_[53360]_ ;
  assign \new_[53372]_  = A199 & ~A168;
  assign \new_[53373]_  = A169 & \new_[53372]_ ;
  assign \new_[53377]_  = ~A202 & ~A201;
  assign \new_[53378]_  = ~A200 & \new_[53377]_ ;
  assign \new_[53379]_  = \new_[53378]_  & \new_[53373]_ ;
  assign \new_[53383]_  = ~A268 & A267;
  assign \new_[53384]_  = A203 & \new_[53383]_ ;
  assign \new_[53387]_  = A300 & A269;
  assign \new_[53390]_  = A302 & ~A301;
  assign \new_[53391]_  = \new_[53390]_  & \new_[53387]_ ;
  assign \new_[53392]_  = \new_[53391]_  & \new_[53384]_ ;
  assign \new_[53396]_  = A168 & ~A169;
  assign \new_[53397]_  = ~A170 & \new_[53396]_ ;
  assign \new_[53401]_  = ~A234 & A233;
  assign \new_[53402]_  = ~A232 & \new_[53401]_ ;
  assign \new_[53403]_  = \new_[53402]_  & \new_[53397]_ ;
  assign \new_[53407]_  = ~A265 & A236;
  assign \new_[53408]_  = ~A235 & \new_[53407]_ ;
  assign \new_[53411]_  = ~A267 & A266;
  assign \new_[53414]_  = A269 & ~A268;
  assign \new_[53415]_  = \new_[53414]_  & \new_[53411]_ ;
  assign \new_[53416]_  = \new_[53415]_  & \new_[53408]_ ;
  assign \new_[53420]_  = A168 & ~A169;
  assign \new_[53421]_  = ~A170 & \new_[53420]_ ;
  assign \new_[53425]_  = ~A234 & A233;
  assign \new_[53426]_  = ~A232 & \new_[53425]_ ;
  assign \new_[53427]_  = \new_[53426]_  & \new_[53421]_ ;
  assign \new_[53431]_  = A265 & A236;
  assign \new_[53432]_  = ~A235 & \new_[53431]_ ;
  assign \new_[53435]_  = ~A267 & ~A266;
  assign \new_[53438]_  = A269 & ~A268;
  assign \new_[53439]_  = \new_[53438]_  & \new_[53435]_ ;
  assign \new_[53440]_  = \new_[53439]_  & \new_[53432]_ ;
  assign \new_[53444]_  = A168 & ~A169;
  assign \new_[53445]_  = ~A170 & \new_[53444]_ ;
  assign \new_[53449]_  = ~A234 & ~A233;
  assign \new_[53450]_  = A232 & \new_[53449]_ ;
  assign \new_[53451]_  = \new_[53450]_  & \new_[53445]_ ;
  assign \new_[53455]_  = ~A265 & A236;
  assign \new_[53456]_  = ~A235 & \new_[53455]_ ;
  assign \new_[53459]_  = ~A267 & A266;
  assign \new_[53462]_  = A269 & ~A268;
  assign \new_[53463]_  = \new_[53462]_  & \new_[53459]_ ;
  assign \new_[53464]_  = \new_[53463]_  & \new_[53456]_ ;
  assign \new_[53468]_  = A168 & ~A169;
  assign \new_[53469]_  = ~A170 & \new_[53468]_ ;
  assign \new_[53473]_  = ~A234 & ~A233;
  assign \new_[53474]_  = A232 & \new_[53473]_ ;
  assign \new_[53475]_  = \new_[53474]_  & \new_[53469]_ ;
  assign \new_[53479]_  = A265 & A236;
  assign \new_[53480]_  = ~A235 & \new_[53479]_ ;
  assign \new_[53483]_  = ~A267 & ~A266;
  assign \new_[53486]_  = A269 & ~A268;
  assign \new_[53487]_  = \new_[53486]_  & \new_[53483]_ ;
  assign \new_[53488]_  = \new_[53487]_  & \new_[53480]_ ;
  assign \new_[53492]_  = A168 & ~A169;
  assign \new_[53493]_  = ~A170 & \new_[53492]_ ;
  assign \new_[53497]_  = A201 & A200;
  assign \new_[53498]_  = ~A199 & \new_[53497]_ ;
  assign \new_[53499]_  = \new_[53498]_  & \new_[53493]_ ;
  assign \new_[53503]_  = ~A268 & A267;
  assign \new_[53504]_  = A202 & \new_[53503]_ ;
  assign \new_[53507]_  = A300 & A269;
  assign \new_[53510]_  = A302 & ~A301;
  assign \new_[53511]_  = \new_[53510]_  & \new_[53507]_ ;
  assign \new_[53512]_  = \new_[53511]_  & \new_[53504]_ ;
  assign \new_[53516]_  = A168 & ~A169;
  assign \new_[53517]_  = ~A170 & \new_[53516]_ ;
  assign \new_[53521]_  = A201 & A200;
  assign \new_[53522]_  = ~A199 & \new_[53521]_ ;
  assign \new_[53523]_  = \new_[53522]_  & \new_[53517]_ ;
  assign \new_[53527]_  = ~A268 & A267;
  assign \new_[53528]_  = ~A203 & \new_[53527]_ ;
  assign \new_[53531]_  = A300 & A269;
  assign \new_[53534]_  = A302 & ~A301;
  assign \new_[53535]_  = \new_[53534]_  & \new_[53531]_ ;
  assign \new_[53536]_  = \new_[53535]_  & \new_[53528]_ ;
  assign \new_[53540]_  = A168 & ~A169;
  assign \new_[53541]_  = ~A170 & \new_[53540]_ ;
  assign \new_[53545]_  = ~A201 & A200;
  assign \new_[53546]_  = ~A199 & \new_[53545]_ ;
  assign \new_[53547]_  = \new_[53546]_  & \new_[53541]_ ;
  assign \new_[53551]_  = A267 & A203;
  assign \new_[53552]_  = ~A202 & \new_[53551]_ ;
  assign \new_[53555]_  = A269 & ~A268;
  assign \new_[53558]_  = A301 & ~A300;
  assign \new_[53559]_  = \new_[53558]_  & \new_[53555]_ ;
  assign \new_[53560]_  = \new_[53559]_  & \new_[53552]_ ;
  assign \new_[53564]_  = A168 & ~A169;
  assign \new_[53565]_  = ~A170 & \new_[53564]_ ;
  assign \new_[53569]_  = ~A201 & A200;
  assign \new_[53570]_  = ~A199 & \new_[53569]_ ;
  assign \new_[53571]_  = \new_[53570]_  & \new_[53565]_ ;
  assign \new_[53575]_  = A267 & A203;
  assign \new_[53576]_  = ~A202 & \new_[53575]_ ;
  assign \new_[53579]_  = A269 & ~A268;
  assign \new_[53582]_  = ~A302 & ~A300;
  assign \new_[53583]_  = \new_[53582]_  & \new_[53579]_ ;
  assign \new_[53584]_  = \new_[53583]_  & \new_[53576]_ ;
  assign \new_[53588]_  = A168 & ~A169;
  assign \new_[53589]_  = ~A170 & \new_[53588]_ ;
  assign \new_[53593]_  = ~A201 & A200;
  assign \new_[53594]_  = ~A199 & \new_[53593]_ ;
  assign \new_[53595]_  = \new_[53594]_  & \new_[53589]_ ;
  assign \new_[53599]_  = A267 & A203;
  assign \new_[53600]_  = ~A202 & \new_[53599]_ ;
  assign \new_[53603]_  = A269 & ~A268;
  assign \new_[53606]_  = A299 & A298;
  assign \new_[53607]_  = \new_[53606]_  & \new_[53603]_ ;
  assign \new_[53608]_  = \new_[53607]_  & \new_[53600]_ ;
  assign \new_[53612]_  = A168 & ~A169;
  assign \new_[53613]_  = ~A170 & \new_[53612]_ ;
  assign \new_[53617]_  = ~A201 & A200;
  assign \new_[53618]_  = ~A199 & \new_[53617]_ ;
  assign \new_[53619]_  = \new_[53618]_  & \new_[53613]_ ;
  assign \new_[53623]_  = A267 & A203;
  assign \new_[53624]_  = ~A202 & \new_[53623]_ ;
  assign \new_[53627]_  = A269 & ~A268;
  assign \new_[53630]_  = ~A299 & ~A298;
  assign \new_[53631]_  = \new_[53630]_  & \new_[53627]_ ;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53624]_ ;
  assign \new_[53636]_  = A168 & ~A169;
  assign \new_[53637]_  = ~A170 & \new_[53636]_ ;
  assign \new_[53641]_  = ~A201 & A200;
  assign \new_[53642]_  = ~A199 & \new_[53641]_ ;
  assign \new_[53643]_  = \new_[53642]_  & \new_[53637]_ ;
  assign \new_[53647]_  = ~A267 & A203;
  assign \new_[53648]_  = ~A202 & \new_[53647]_ ;
  assign \new_[53651]_  = A300 & A268;
  assign \new_[53654]_  = A302 & ~A301;
  assign \new_[53655]_  = \new_[53654]_  & \new_[53651]_ ;
  assign \new_[53656]_  = \new_[53655]_  & \new_[53648]_ ;
  assign \new_[53660]_  = A168 & ~A169;
  assign \new_[53661]_  = ~A170 & \new_[53660]_ ;
  assign \new_[53665]_  = ~A201 & A200;
  assign \new_[53666]_  = ~A199 & \new_[53665]_ ;
  assign \new_[53667]_  = \new_[53666]_  & \new_[53661]_ ;
  assign \new_[53671]_  = ~A267 & A203;
  assign \new_[53672]_  = ~A202 & \new_[53671]_ ;
  assign \new_[53675]_  = A300 & ~A269;
  assign \new_[53678]_  = A302 & ~A301;
  assign \new_[53679]_  = \new_[53678]_  & \new_[53675]_ ;
  assign \new_[53680]_  = \new_[53679]_  & \new_[53672]_ ;
  assign \new_[53684]_  = A168 & ~A169;
  assign \new_[53685]_  = ~A170 & \new_[53684]_ ;
  assign \new_[53689]_  = ~A201 & A200;
  assign \new_[53690]_  = ~A199 & \new_[53689]_ ;
  assign \new_[53691]_  = \new_[53690]_  & \new_[53685]_ ;
  assign \new_[53695]_  = A265 & A203;
  assign \new_[53696]_  = ~A202 & \new_[53695]_ ;
  assign \new_[53699]_  = A300 & A266;
  assign \new_[53702]_  = A302 & ~A301;
  assign \new_[53703]_  = \new_[53702]_  & \new_[53699]_ ;
  assign \new_[53704]_  = \new_[53703]_  & \new_[53696]_ ;
  assign \new_[53708]_  = A168 & ~A169;
  assign \new_[53709]_  = ~A170 & \new_[53708]_ ;
  assign \new_[53713]_  = ~A201 & A200;
  assign \new_[53714]_  = ~A199 & \new_[53713]_ ;
  assign \new_[53715]_  = \new_[53714]_  & \new_[53709]_ ;
  assign \new_[53719]_  = ~A265 & A203;
  assign \new_[53720]_  = ~A202 & \new_[53719]_ ;
  assign \new_[53723]_  = A300 & ~A266;
  assign \new_[53726]_  = A302 & ~A301;
  assign \new_[53727]_  = \new_[53726]_  & \new_[53723]_ ;
  assign \new_[53728]_  = \new_[53727]_  & \new_[53720]_ ;
  assign \new_[53732]_  = A168 & ~A169;
  assign \new_[53733]_  = ~A170 & \new_[53732]_ ;
  assign \new_[53737]_  = A201 & ~A200;
  assign \new_[53738]_  = A199 & \new_[53737]_ ;
  assign \new_[53739]_  = \new_[53738]_  & \new_[53733]_ ;
  assign \new_[53743]_  = ~A268 & A267;
  assign \new_[53744]_  = A202 & \new_[53743]_ ;
  assign \new_[53747]_  = A300 & A269;
  assign \new_[53750]_  = A302 & ~A301;
  assign \new_[53751]_  = \new_[53750]_  & \new_[53747]_ ;
  assign \new_[53752]_  = \new_[53751]_  & \new_[53744]_ ;
  assign \new_[53756]_  = A168 & ~A169;
  assign \new_[53757]_  = ~A170 & \new_[53756]_ ;
  assign \new_[53761]_  = A201 & ~A200;
  assign \new_[53762]_  = A199 & \new_[53761]_ ;
  assign \new_[53763]_  = \new_[53762]_  & \new_[53757]_ ;
  assign \new_[53767]_  = ~A268 & A267;
  assign \new_[53768]_  = ~A203 & \new_[53767]_ ;
  assign \new_[53771]_  = A300 & A269;
  assign \new_[53774]_  = A302 & ~A301;
  assign \new_[53775]_  = \new_[53774]_  & \new_[53771]_ ;
  assign \new_[53776]_  = \new_[53775]_  & \new_[53768]_ ;
  assign \new_[53780]_  = A168 & ~A169;
  assign \new_[53781]_  = ~A170 & \new_[53780]_ ;
  assign \new_[53785]_  = ~A201 & ~A200;
  assign \new_[53786]_  = A199 & \new_[53785]_ ;
  assign \new_[53787]_  = \new_[53786]_  & \new_[53781]_ ;
  assign \new_[53791]_  = A267 & A203;
  assign \new_[53792]_  = ~A202 & \new_[53791]_ ;
  assign \new_[53795]_  = A269 & ~A268;
  assign \new_[53798]_  = A301 & ~A300;
  assign \new_[53799]_  = \new_[53798]_  & \new_[53795]_ ;
  assign \new_[53800]_  = \new_[53799]_  & \new_[53792]_ ;
  assign \new_[53804]_  = A168 & ~A169;
  assign \new_[53805]_  = ~A170 & \new_[53804]_ ;
  assign \new_[53809]_  = ~A201 & ~A200;
  assign \new_[53810]_  = A199 & \new_[53809]_ ;
  assign \new_[53811]_  = \new_[53810]_  & \new_[53805]_ ;
  assign \new_[53815]_  = A267 & A203;
  assign \new_[53816]_  = ~A202 & \new_[53815]_ ;
  assign \new_[53819]_  = A269 & ~A268;
  assign \new_[53822]_  = ~A302 & ~A300;
  assign \new_[53823]_  = \new_[53822]_  & \new_[53819]_ ;
  assign \new_[53824]_  = \new_[53823]_  & \new_[53816]_ ;
  assign \new_[53828]_  = A168 & ~A169;
  assign \new_[53829]_  = ~A170 & \new_[53828]_ ;
  assign \new_[53833]_  = ~A201 & ~A200;
  assign \new_[53834]_  = A199 & \new_[53833]_ ;
  assign \new_[53835]_  = \new_[53834]_  & \new_[53829]_ ;
  assign \new_[53839]_  = A267 & A203;
  assign \new_[53840]_  = ~A202 & \new_[53839]_ ;
  assign \new_[53843]_  = A269 & ~A268;
  assign \new_[53846]_  = A299 & A298;
  assign \new_[53847]_  = \new_[53846]_  & \new_[53843]_ ;
  assign \new_[53848]_  = \new_[53847]_  & \new_[53840]_ ;
  assign \new_[53852]_  = A168 & ~A169;
  assign \new_[53853]_  = ~A170 & \new_[53852]_ ;
  assign \new_[53857]_  = ~A201 & ~A200;
  assign \new_[53858]_  = A199 & \new_[53857]_ ;
  assign \new_[53859]_  = \new_[53858]_  & \new_[53853]_ ;
  assign \new_[53863]_  = A267 & A203;
  assign \new_[53864]_  = ~A202 & \new_[53863]_ ;
  assign \new_[53867]_  = A269 & ~A268;
  assign \new_[53870]_  = ~A299 & ~A298;
  assign \new_[53871]_  = \new_[53870]_  & \new_[53867]_ ;
  assign \new_[53872]_  = \new_[53871]_  & \new_[53864]_ ;
  assign \new_[53876]_  = A168 & ~A169;
  assign \new_[53877]_  = ~A170 & \new_[53876]_ ;
  assign \new_[53881]_  = ~A201 & ~A200;
  assign \new_[53882]_  = A199 & \new_[53881]_ ;
  assign \new_[53883]_  = \new_[53882]_  & \new_[53877]_ ;
  assign \new_[53887]_  = ~A267 & A203;
  assign \new_[53888]_  = ~A202 & \new_[53887]_ ;
  assign \new_[53891]_  = A300 & A268;
  assign \new_[53894]_  = A302 & ~A301;
  assign \new_[53895]_  = \new_[53894]_  & \new_[53891]_ ;
  assign \new_[53896]_  = \new_[53895]_  & \new_[53888]_ ;
  assign \new_[53900]_  = A168 & ~A169;
  assign \new_[53901]_  = ~A170 & \new_[53900]_ ;
  assign \new_[53905]_  = ~A201 & ~A200;
  assign \new_[53906]_  = A199 & \new_[53905]_ ;
  assign \new_[53907]_  = \new_[53906]_  & \new_[53901]_ ;
  assign \new_[53911]_  = ~A267 & A203;
  assign \new_[53912]_  = ~A202 & \new_[53911]_ ;
  assign \new_[53915]_  = A300 & ~A269;
  assign \new_[53918]_  = A302 & ~A301;
  assign \new_[53919]_  = \new_[53918]_  & \new_[53915]_ ;
  assign \new_[53920]_  = \new_[53919]_  & \new_[53912]_ ;
  assign \new_[53924]_  = A168 & ~A169;
  assign \new_[53925]_  = ~A170 & \new_[53924]_ ;
  assign \new_[53929]_  = ~A201 & ~A200;
  assign \new_[53930]_  = A199 & \new_[53929]_ ;
  assign \new_[53931]_  = \new_[53930]_  & \new_[53925]_ ;
  assign \new_[53935]_  = A265 & A203;
  assign \new_[53936]_  = ~A202 & \new_[53935]_ ;
  assign \new_[53939]_  = A300 & A266;
  assign \new_[53942]_  = A302 & ~A301;
  assign \new_[53943]_  = \new_[53942]_  & \new_[53939]_ ;
  assign \new_[53944]_  = \new_[53943]_  & \new_[53936]_ ;
  assign \new_[53948]_  = A168 & ~A169;
  assign \new_[53949]_  = ~A170 & \new_[53948]_ ;
  assign \new_[53953]_  = ~A201 & ~A200;
  assign \new_[53954]_  = A199 & \new_[53953]_ ;
  assign \new_[53955]_  = \new_[53954]_  & \new_[53949]_ ;
  assign \new_[53959]_  = ~A265 & A203;
  assign \new_[53960]_  = ~A202 & \new_[53959]_ ;
  assign \new_[53963]_  = A300 & ~A266;
  assign \new_[53966]_  = A302 & ~A301;
  assign \new_[53967]_  = \new_[53966]_  & \new_[53963]_ ;
  assign \new_[53968]_  = \new_[53967]_  & \new_[53960]_ ;
  assign \new_[53972]_  = ~A168 & ~A169;
  assign \new_[53973]_  = ~A170 & \new_[53972]_ ;
  assign \new_[53977]_  = ~A201 & ~A166;
  assign \new_[53978]_  = A167 & \new_[53977]_ ;
  assign \new_[53979]_  = \new_[53978]_  & \new_[53973]_ ;
  assign \new_[53983]_  = A268 & ~A267;
  assign \new_[53984]_  = A202 & \new_[53983]_ ;
  assign \new_[53987]_  = ~A299 & A298;
  assign \new_[53990]_  = A301 & A300;
  assign \new_[53991]_  = \new_[53990]_  & \new_[53987]_ ;
  assign \new_[53992]_  = \new_[53991]_  & \new_[53984]_ ;
  assign \new_[53996]_  = ~A168 & ~A169;
  assign \new_[53997]_  = ~A170 & \new_[53996]_ ;
  assign \new_[54001]_  = ~A201 & ~A166;
  assign \new_[54002]_  = A167 & \new_[54001]_ ;
  assign \new_[54003]_  = \new_[54002]_  & \new_[53997]_ ;
  assign \new_[54007]_  = A268 & ~A267;
  assign \new_[54008]_  = A202 & \new_[54007]_ ;
  assign \new_[54011]_  = ~A299 & A298;
  assign \new_[54014]_  = ~A302 & A300;
  assign \new_[54015]_  = \new_[54014]_  & \new_[54011]_ ;
  assign \new_[54016]_  = \new_[54015]_  & \new_[54008]_ ;
  assign \new_[54020]_  = ~A168 & ~A169;
  assign \new_[54021]_  = ~A170 & \new_[54020]_ ;
  assign \new_[54025]_  = ~A201 & ~A166;
  assign \new_[54026]_  = A167 & \new_[54025]_ ;
  assign \new_[54027]_  = \new_[54026]_  & \new_[54021]_ ;
  assign \new_[54031]_  = A268 & ~A267;
  assign \new_[54032]_  = A202 & \new_[54031]_ ;
  assign \new_[54035]_  = A299 & ~A298;
  assign \new_[54038]_  = A301 & A300;
  assign \new_[54039]_  = \new_[54038]_  & \new_[54035]_ ;
  assign \new_[54040]_  = \new_[54039]_  & \new_[54032]_ ;
  assign \new_[54044]_  = ~A168 & ~A169;
  assign \new_[54045]_  = ~A170 & \new_[54044]_ ;
  assign \new_[54049]_  = ~A201 & ~A166;
  assign \new_[54050]_  = A167 & \new_[54049]_ ;
  assign \new_[54051]_  = \new_[54050]_  & \new_[54045]_ ;
  assign \new_[54055]_  = A268 & ~A267;
  assign \new_[54056]_  = A202 & \new_[54055]_ ;
  assign \new_[54059]_  = A299 & ~A298;
  assign \new_[54062]_  = ~A302 & A300;
  assign \new_[54063]_  = \new_[54062]_  & \new_[54059]_ ;
  assign \new_[54064]_  = \new_[54063]_  & \new_[54056]_ ;
  assign \new_[54068]_  = ~A168 & ~A169;
  assign \new_[54069]_  = ~A170 & \new_[54068]_ ;
  assign \new_[54073]_  = ~A201 & ~A166;
  assign \new_[54074]_  = A167 & \new_[54073]_ ;
  assign \new_[54075]_  = \new_[54074]_  & \new_[54069]_ ;
  assign \new_[54079]_  = ~A269 & ~A267;
  assign \new_[54080]_  = A202 & \new_[54079]_ ;
  assign \new_[54083]_  = ~A299 & A298;
  assign \new_[54086]_  = A301 & A300;
  assign \new_[54087]_  = \new_[54086]_  & \new_[54083]_ ;
  assign \new_[54088]_  = \new_[54087]_  & \new_[54080]_ ;
  assign \new_[54092]_  = ~A168 & ~A169;
  assign \new_[54093]_  = ~A170 & \new_[54092]_ ;
  assign \new_[54097]_  = ~A201 & ~A166;
  assign \new_[54098]_  = A167 & \new_[54097]_ ;
  assign \new_[54099]_  = \new_[54098]_  & \new_[54093]_ ;
  assign \new_[54103]_  = ~A269 & ~A267;
  assign \new_[54104]_  = A202 & \new_[54103]_ ;
  assign \new_[54107]_  = ~A299 & A298;
  assign \new_[54110]_  = ~A302 & A300;
  assign \new_[54111]_  = \new_[54110]_  & \new_[54107]_ ;
  assign \new_[54112]_  = \new_[54111]_  & \new_[54104]_ ;
  assign \new_[54116]_  = ~A168 & ~A169;
  assign \new_[54117]_  = ~A170 & \new_[54116]_ ;
  assign \new_[54121]_  = ~A201 & ~A166;
  assign \new_[54122]_  = A167 & \new_[54121]_ ;
  assign \new_[54123]_  = \new_[54122]_  & \new_[54117]_ ;
  assign \new_[54127]_  = ~A269 & ~A267;
  assign \new_[54128]_  = A202 & \new_[54127]_ ;
  assign \new_[54131]_  = A299 & ~A298;
  assign \new_[54134]_  = A301 & A300;
  assign \new_[54135]_  = \new_[54134]_  & \new_[54131]_ ;
  assign \new_[54136]_  = \new_[54135]_  & \new_[54128]_ ;
  assign \new_[54140]_  = ~A168 & ~A169;
  assign \new_[54141]_  = ~A170 & \new_[54140]_ ;
  assign \new_[54145]_  = ~A201 & ~A166;
  assign \new_[54146]_  = A167 & \new_[54145]_ ;
  assign \new_[54147]_  = \new_[54146]_  & \new_[54141]_ ;
  assign \new_[54151]_  = ~A269 & ~A267;
  assign \new_[54152]_  = A202 & \new_[54151]_ ;
  assign \new_[54155]_  = A299 & ~A298;
  assign \new_[54158]_  = ~A302 & A300;
  assign \new_[54159]_  = \new_[54158]_  & \new_[54155]_ ;
  assign \new_[54160]_  = \new_[54159]_  & \new_[54152]_ ;
  assign \new_[54164]_  = ~A168 & ~A169;
  assign \new_[54165]_  = ~A170 & \new_[54164]_ ;
  assign \new_[54169]_  = ~A201 & ~A166;
  assign \new_[54170]_  = A167 & \new_[54169]_ ;
  assign \new_[54171]_  = \new_[54170]_  & \new_[54165]_ ;
  assign \new_[54175]_  = A266 & A265;
  assign \new_[54176]_  = A202 & \new_[54175]_ ;
  assign \new_[54179]_  = ~A299 & A298;
  assign \new_[54182]_  = A301 & A300;
  assign \new_[54183]_  = \new_[54182]_  & \new_[54179]_ ;
  assign \new_[54184]_  = \new_[54183]_  & \new_[54176]_ ;
  assign \new_[54188]_  = ~A168 & ~A169;
  assign \new_[54189]_  = ~A170 & \new_[54188]_ ;
  assign \new_[54193]_  = ~A201 & ~A166;
  assign \new_[54194]_  = A167 & \new_[54193]_ ;
  assign \new_[54195]_  = \new_[54194]_  & \new_[54189]_ ;
  assign \new_[54199]_  = A266 & A265;
  assign \new_[54200]_  = A202 & \new_[54199]_ ;
  assign \new_[54203]_  = ~A299 & A298;
  assign \new_[54206]_  = ~A302 & A300;
  assign \new_[54207]_  = \new_[54206]_  & \new_[54203]_ ;
  assign \new_[54208]_  = \new_[54207]_  & \new_[54200]_ ;
  assign \new_[54212]_  = ~A168 & ~A169;
  assign \new_[54213]_  = ~A170 & \new_[54212]_ ;
  assign \new_[54217]_  = ~A201 & ~A166;
  assign \new_[54218]_  = A167 & \new_[54217]_ ;
  assign \new_[54219]_  = \new_[54218]_  & \new_[54213]_ ;
  assign \new_[54223]_  = A266 & A265;
  assign \new_[54224]_  = A202 & \new_[54223]_ ;
  assign \new_[54227]_  = A299 & ~A298;
  assign \new_[54230]_  = A301 & A300;
  assign \new_[54231]_  = \new_[54230]_  & \new_[54227]_ ;
  assign \new_[54232]_  = \new_[54231]_  & \new_[54224]_ ;
  assign \new_[54236]_  = ~A168 & ~A169;
  assign \new_[54237]_  = ~A170 & \new_[54236]_ ;
  assign \new_[54241]_  = ~A201 & ~A166;
  assign \new_[54242]_  = A167 & \new_[54241]_ ;
  assign \new_[54243]_  = \new_[54242]_  & \new_[54237]_ ;
  assign \new_[54247]_  = A266 & A265;
  assign \new_[54248]_  = A202 & \new_[54247]_ ;
  assign \new_[54251]_  = A299 & ~A298;
  assign \new_[54254]_  = ~A302 & A300;
  assign \new_[54255]_  = \new_[54254]_  & \new_[54251]_ ;
  assign \new_[54256]_  = \new_[54255]_  & \new_[54248]_ ;
  assign \new_[54260]_  = ~A168 & ~A169;
  assign \new_[54261]_  = ~A170 & \new_[54260]_ ;
  assign \new_[54265]_  = ~A201 & ~A166;
  assign \new_[54266]_  = A167 & \new_[54265]_ ;
  assign \new_[54267]_  = \new_[54266]_  & \new_[54261]_ ;
  assign \new_[54271]_  = A266 & ~A265;
  assign \new_[54272]_  = A202 & \new_[54271]_ ;
  assign \new_[54275]_  = A268 & A267;
  assign \new_[54278]_  = A301 & ~A300;
  assign \new_[54279]_  = \new_[54278]_  & \new_[54275]_ ;
  assign \new_[54280]_  = \new_[54279]_  & \new_[54272]_ ;
  assign \new_[54284]_  = ~A168 & ~A169;
  assign \new_[54285]_  = ~A170 & \new_[54284]_ ;
  assign \new_[54289]_  = ~A201 & ~A166;
  assign \new_[54290]_  = A167 & \new_[54289]_ ;
  assign \new_[54291]_  = \new_[54290]_  & \new_[54285]_ ;
  assign \new_[54295]_  = A266 & ~A265;
  assign \new_[54296]_  = A202 & \new_[54295]_ ;
  assign \new_[54299]_  = A268 & A267;
  assign \new_[54302]_  = ~A302 & ~A300;
  assign \new_[54303]_  = \new_[54302]_  & \new_[54299]_ ;
  assign \new_[54304]_  = \new_[54303]_  & \new_[54296]_ ;
  assign \new_[54308]_  = ~A168 & ~A169;
  assign \new_[54309]_  = ~A170 & \new_[54308]_ ;
  assign \new_[54313]_  = ~A201 & ~A166;
  assign \new_[54314]_  = A167 & \new_[54313]_ ;
  assign \new_[54315]_  = \new_[54314]_  & \new_[54309]_ ;
  assign \new_[54319]_  = A266 & ~A265;
  assign \new_[54320]_  = A202 & \new_[54319]_ ;
  assign \new_[54323]_  = A268 & A267;
  assign \new_[54326]_  = A299 & A298;
  assign \new_[54327]_  = \new_[54326]_  & \new_[54323]_ ;
  assign \new_[54328]_  = \new_[54327]_  & \new_[54320]_ ;
  assign \new_[54332]_  = ~A168 & ~A169;
  assign \new_[54333]_  = ~A170 & \new_[54332]_ ;
  assign \new_[54337]_  = ~A201 & ~A166;
  assign \new_[54338]_  = A167 & \new_[54337]_ ;
  assign \new_[54339]_  = \new_[54338]_  & \new_[54333]_ ;
  assign \new_[54343]_  = A266 & ~A265;
  assign \new_[54344]_  = A202 & \new_[54343]_ ;
  assign \new_[54347]_  = A268 & A267;
  assign \new_[54350]_  = ~A299 & ~A298;
  assign \new_[54351]_  = \new_[54350]_  & \new_[54347]_ ;
  assign \new_[54352]_  = \new_[54351]_  & \new_[54344]_ ;
  assign \new_[54356]_  = ~A168 & ~A169;
  assign \new_[54357]_  = ~A170 & \new_[54356]_ ;
  assign \new_[54361]_  = ~A201 & ~A166;
  assign \new_[54362]_  = A167 & \new_[54361]_ ;
  assign \new_[54363]_  = \new_[54362]_  & \new_[54357]_ ;
  assign \new_[54367]_  = A266 & ~A265;
  assign \new_[54368]_  = A202 & \new_[54367]_ ;
  assign \new_[54371]_  = ~A269 & A267;
  assign \new_[54374]_  = A301 & ~A300;
  assign \new_[54375]_  = \new_[54374]_  & \new_[54371]_ ;
  assign \new_[54376]_  = \new_[54375]_  & \new_[54368]_ ;
  assign \new_[54380]_  = ~A168 & ~A169;
  assign \new_[54381]_  = ~A170 & \new_[54380]_ ;
  assign \new_[54385]_  = ~A201 & ~A166;
  assign \new_[54386]_  = A167 & \new_[54385]_ ;
  assign \new_[54387]_  = \new_[54386]_  & \new_[54381]_ ;
  assign \new_[54391]_  = A266 & ~A265;
  assign \new_[54392]_  = A202 & \new_[54391]_ ;
  assign \new_[54395]_  = ~A269 & A267;
  assign \new_[54398]_  = ~A302 & ~A300;
  assign \new_[54399]_  = \new_[54398]_  & \new_[54395]_ ;
  assign \new_[54400]_  = \new_[54399]_  & \new_[54392]_ ;
  assign \new_[54404]_  = ~A168 & ~A169;
  assign \new_[54405]_  = ~A170 & \new_[54404]_ ;
  assign \new_[54409]_  = ~A201 & ~A166;
  assign \new_[54410]_  = A167 & \new_[54409]_ ;
  assign \new_[54411]_  = \new_[54410]_  & \new_[54405]_ ;
  assign \new_[54415]_  = A266 & ~A265;
  assign \new_[54416]_  = A202 & \new_[54415]_ ;
  assign \new_[54419]_  = ~A269 & A267;
  assign \new_[54422]_  = A299 & A298;
  assign \new_[54423]_  = \new_[54422]_  & \new_[54419]_ ;
  assign \new_[54424]_  = \new_[54423]_  & \new_[54416]_ ;
  assign \new_[54428]_  = ~A168 & ~A169;
  assign \new_[54429]_  = ~A170 & \new_[54428]_ ;
  assign \new_[54433]_  = ~A201 & ~A166;
  assign \new_[54434]_  = A167 & \new_[54433]_ ;
  assign \new_[54435]_  = \new_[54434]_  & \new_[54429]_ ;
  assign \new_[54439]_  = A266 & ~A265;
  assign \new_[54440]_  = A202 & \new_[54439]_ ;
  assign \new_[54443]_  = ~A269 & A267;
  assign \new_[54446]_  = ~A299 & ~A298;
  assign \new_[54447]_  = \new_[54446]_  & \new_[54443]_ ;
  assign \new_[54448]_  = \new_[54447]_  & \new_[54440]_ ;
  assign \new_[54452]_  = ~A168 & ~A169;
  assign \new_[54453]_  = ~A170 & \new_[54452]_ ;
  assign \new_[54457]_  = ~A201 & ~A166;
  assign \new_[54458]_  = A167 & \new_[54457]_ ;
  assign \new_[54459]_  = \new_[54458]_  & \new_[54453]_ ;
  assign \new_[54463]_  = ~A266 & A265;
  assign \new_[54464]_  = A202 & \new_[54463]_ ;
  assign \new_[54467]_  = A268 & A267;
  assign \new_[54470]_  = A301 & ~A300;
  assign \new_[54471]_  = \new_[54470]_  & \new_[54467]_ ;
  assign \new_[54472]_  = \new_[54471]_  & \new_[54464]_ ;
  assign \new_[54476]_  = ~A168 & ~A169;
  assign \new_[54477]_  = ~A170 & \new_[54476]_ ;
  assign \new_[54481]_  = ~A201 & ~A166;
  assign \new_[54482]_  = A167 & \new_[54481]_ ;
  assign \new_[54483]_  = \new_[54482]_  & \new_[54477]_ ;
  assign \new_[54487]_  = ~A266 & A265;
  assign \new_[54488]_  = A202 & \new_[54487]_ ;
  assign \new_[54491]_  = A268 & A267;
  assign \new_[54494]_  = ~A302 & ~A300;
  assign \new_[54495]_  = \new_[54494]_  & \new_[54491]_ ;
  assign \new_[54496]_  = \new_[54495]_  & \new_[54488]_ ;
  assign \new_[54500]_  = ~A168 & ~A169;
  assign \new_[54501]_  = ~A170 & \new_[54500]_ ;
  assign \new_[54505]_  = ~A201 & ~A166;
  assign \new_[54506]_  = A167 & \new_[54505]_ ;
  assign \new_[54507]_  = \new_[54506]_  & \new_[54501]_ ;
  assign \new_[54511]_  = ~A266 & A265;
  assign \new_[54512]_  = A202 & \new_[54511]_ ;
  assign \new_[54515]_  = A268 & A267;
  assign \new_[54518]_  = A299 & A298;
  assign \new_[54519]_  = \new_[54518]_  & \new_[54515]_ ;
  assign \new_[54520]_  = \new_[54519]_  & \new_[54512]_ ;
  assign \new_[54524]_  = ~A168 & ~A169;
  assign \new_[54525]_  = ~A170 & \new_[54524]_ ;
  assign \new_[54529]_  = ~A201 & ~A166;
  assign \new_[54530]_  = A167 & \new_[54529]_ ;
  assign \new_[54531]_  = \new_[54530]_  & \new_[54525]_ ;
  assign \new_[54535]_  = ~A266 & A265;
  assign \new_[54536]_  = A202 & \new_[54535]_ ;
  assign \new_[54539]_  = A268 & A267;
  assign \new_[54542]_  = ~A299 & ~A298;
  assign \new_[54543]_  = \new_[54542]_  & \new_[54539]_ ;
  assign \new_[54544]_  = \new_[54543]_  & \new_[54536]_ ;
  assign \new_[54548]_  = ~A168 & ~A169;
  assign \new_[54549]_  = ~A170 & \new_[54548]_ ;
  assign \new_[54553]_  = ~A201 & ~A166;
  assign \new_[54554]_  = A167 & \new_[54553]_ ;
  assign \new_[54555]_  = \new_[54554]_  & \new_[54549]_ ;
  assign \new_[54559]_  = ~A266 & A265;
  assign \new_[54560]_  = A202 & \new_[54559]_ ;
  assign \new_[54563]_  = ~A269 & A267;
  assign \new_[54566]_  = A301 & ~A300;
  assign \new_[54567]_  = \new_[54566]_  & \new_[54563]_ ;
  assign \new_[54568]_  = \new_[54567]_  & \new_[54560]_ ;
  assign \new_[54572]_  = ~A168 & ~A169;
  assign \new_[54573]_  = ~A170 & \new_[54572]_ ;
  assign \new_[54577]_  = ~A201 & ~A166;
  assign \new_[54578]_  = A167 & \new_[54577]_ ;
  assign \new_[54579]_  = \new_[54578]_  & \new_[54573]_ ;
  assign \new_[54583]_  = ~A266 & A265;
  assign \new_[54584]_  = A202 & \new_[54583]_ ;
  assign \new_[54587]_  = ~A269 & A267;
  assign \new_[54590]_  = ~A302 & ~A300;
  assign \new_[54591]_  = \new_[54590]_  & \new_[54587]_ ;
  assign \new_[54592]_  = \new_[54591]_  & \new_[54584]_ ;
  assign \new_[54596]_  = ~A168 & ~A169;
  assign \new_[54597]_  = ~A170 & \new_[54596]_ ;
  assign \new_[54601]_  = ~A201 & ~A166;
  assign \new_[54602]_  = A167 & \new_[54601]_ ;
  assign \new_[54603]_  = \new_[54602]_  & \new_[54597]_ ;
  assign \new_[54607]_  = ~A266 & A265;
  assign \new_[54608]_  = A202 & \new_[54607]_ ;
  assign \new_[54611]_  = ~A269 & A267;
  assign \new_[54614]_  = A299 & A298;
  assign \new_[54615]_  = \new_[54614]_  & \new_[54611]_ ;
  assign \new_[54616]_  = \new_[54615]_  & \new_[54608]_ ;
  assign \new_[54620]_  = ~A168 & ~A169;
  assign \new_[54621]_  = ~A170 & \new_[54620]_ ;
  assign \new_[54625]_  = ~A201 & ~A166;
  assign \new_[54626]_  = A167 & \new_[54625]_ ;
  assign \new_[54627]_  = \new_[54626]_  & \new_[54621]_ ;
  assign \new_[54631]_  = ~A266 & A265;
  assign \new_[54632]_  = A202 & \new_[54631]_ ;
  assign \new_[54635]_  = ~A269 & A267;
  assign \new_[54638]_  = ~A299 & ~A298;
  assign \new_[54639]_  = \new_[54638]_  & \new_[54635]_ ;
  assign \new_[54640]_  = \new_[54639]_  & \new_[54632]_ ;
  assign \new_[54644]_  = ~A168 & ~A169;
  assign \new_[54645]_  = ~A170 & \new_[54644]_ ;
  assign \new_[54649]_  = ~A201 & ~A166;
  assign \new_[54650]_  = A167 & \new_[54649]_ ;
  assign \new_[54651]_  = \new_[54650]_  & \new_[54645]_ ;
  assign \new_[54655]_  = ~A266 & ~A265;
  assign \new_[54656]_  = A202 & \new_[54655]_ ;
  assign \new_[54659]_  = ~A299 & A298;
  assign \new_[54662]_  = A301 & A300;
  assign \new_[54663]_  = \new_[54662]_  & \new_[54659]_ ;
  assign \new_[54664]_  = \new_[54663]_  & \new_[54656]_ ;
  assign \new_[54668]_  = ~A168 & ~A169;
  assign \new_[54669]_  = ~A170 & \new_[54668]_ ;
  assign \new_[54673]_  = ~A201 & ~A166;
  assign \new_[54674]_  = A167 & \new_[54673]_ ;
  assign \new_[54675]_  = \new_[54674]_  & \new_[54669]_ ;
  assign \new_[54679]_  = ~A266 & ~A265;
  assign \new_[54680]_  = A202 & \new_[54679]_ ;
  assign \new_[54683]_  = ~A299 & A298;
  assign \new_[54686]_  = ~A302 & A300;
  assign \new_[54687]_  = \new_[54686]_  & \new_[54683]_ ;
  assign \new_[54688]_  = \new_[54687]_  & \new_[54680]_ ;
  assign \new_[54692]_  = ~A168 & ~A169;
  assign \new_[54693]_  = ~A170 & \new_[54692]_ ;
  assign \new_[54697]_  = ~A201 & ~A166;
  assign \new_[54698]_  = A167 & \new_[54697]_ ;
  assign \new_[54699]_  = \new_[54698]_  & \new_[54693]_ ;
  assign \new_[54703]_  = ~A266 & ~A265;
  assign \new_[54704]_  = A202 & \new_[54703]_ ;
  assign \new_[54707]_  = A299 & ~A298;
  assign \new_[54710]_  = A301 & A300;
  assign \new_[54711]_  = \new_[54710]_  & \new_[54707]_ ;
  assign \new_[54712]_  = \new_[54711]_  & \new_[54704]_ ;
  assign \new_[54716]_  = ~A168 & ~A169;
  assign \new_[54717]_  = ~A170 & \new_[54716]_ ;
  assign \new_[54721]_  = ~A201 & ~A166;
  assign \new_[54722]_  = A167 & \new_[54721]_ ;
  assign \new_[54723]_  = \new_[54722]_  & \new_[54717]_ ;
  assign \new_[54727]_  = ~A266 & ~A265;
  assign \new_[54728]_  = A202 & \new_[54727]_ ;
  assign \new_[54731]_  = A299 & ~A298;
  assign \new_[54734]_  = ~A302 & A300;
  assign \new_[54735]_  = \new_[54734]_  & \new_[54731]_ ;
  assign \new_[54736]_  = \new_[54735]_  & \new_[54728]_ ;
  assign \new_[54740]_  = ~A168 & ~A169;
  assign \new_[54741]_  = ~A170 & \new_[54740]_ ;
  assign \new_[54745]_  = ~A201 & ~A166;
  assign \new_[54746]_  = A167 & \new_[54745]_ ;
  assign \new_[54747]_  = \new_[54746]_  & \new_[54741]_ ;
  assign \new_[54751]_  = A268 & ~A267;
  assign \new_[54752]_  = ~A203 & \new_[54751]_ ;
  assign \new_[54755]_  = ~A299 & A298;
  assign \new_[54758]_  = A301 & A300;
  assign \new_[54759]_  = \new_[54758]_  & \new_[54755]_ ;
  assign \new_[54760]_  = \new_[54759]_  & \new_[54752]_ ;
  assign \new_[54764]_  = ~A168 & ~A169;
  assign \new_[54765]_  = ~A170 & \new_[54764]_ ;
  assign \new_[54769]_  = ~A201 & ~A166;
  assign \new_[54770]_  = A167 & \new_[54769]_ ;
  assign \new_[54771]_  = \new_[54770]_  & \new_[54765]_ ;
  assign \new_[54775]_  = A268 & ~A267;
  assign \new_[54776]_  = ~A203 & \new_[54775]_ ;
  assign \new_[54779]_  = ~A299 & A298;
  assign \new_[54782]_  = ~A302 & A300;
  assign \new_[54783]_  = \new_[54782]_  & \new_[54779]_ ;
  assign \new_[54784]_  = \new_[54783]_  & \new_[54776]_ ;
  assign \new_[54788]_  = ~A168 & ~A169;
  assign \new_[54789]_  = ~A170 & \new_[54788]_ ;
  assign \new_[54793]_  = ~A201 & ~A166;
  assign \new_[54794]_  = A167 & \new_[54793]_ ;
  assign \new_[54795]_  = \new_[54794]_  & \new_[54789]_ ;
  assign \new_[54799]_  = A268 & ~A267;
  assign \new_[54800]_  = ~A203 & \new_[54799]_ ;
  assign \new_[54803]_  = A299 & ~A298;
  assign \new_[54806]_  = A301 & A300;
  assign \new_[54807]_  = \new_[54806]_  & \new_[54803]_ ;
  assign \new_[54808]_  = \new_[54807]_  & \new_[54800]_ ;
  assign \new_[54812]_  = ~A168 & ~A169;
  assign \new_[54813]_  = ~A170 & \new_[54812]_ ;
  assign \new_[54817]_  = ~A201 & ~A166;
  assign \new_[54818]_  = A167 & \new_[54817]_ ;
  assign \new_[54819]_  = \new_[54818]_  & \new_[54813]_ ;
  assign \new_[54823]_  = A268 & ~A267;
  assign \new_[54824]_  = ~A203 & \new_[54823]_ ;
  assign \new_[54827]_  = A299 & ~A298;
  assign \new_[54830]_  = ~A302 & A300;
  assign \new_[54831]_  = \new_[54830]_  & \new_[54827]_ ;
  assign \new_[54832]_  = \new_[54831]_  & \new_[54824]_ ;
  assign \new_[54836]_  = ~A168 & ~A169;
  assign \new_[54837]_  = ~A170 & \new_[54836]_ ;
  assign \new_[54841]_  = ~A201 & ~A166;
  assign \new_[54842]_  = A167 & \new_[54841]_ ;
  assign \new_[54843]_  = \new_[54842]_  & \new_[54837]_ ;
  assign \new_[54847]_  = ~A269 & ~A267;
  assign \new_[54848]_  = ~A203 & \new_[54847]_ ;
  assign \new_[54851]_  = ~A299 & A298;
  assign \new_[54854]_  = A301 & A300;
  assign \new_[54855]_  = \new_[54854]_  & \new_[54851]_ ;
  assign \new_[54856]_  = \new_[54855]_  & \new_[54848]_ ;
  assign \new_[54860]_  = ~A168 & ~A169;
  assign \new_[54861]_  = ~A170 & \new_[54860]_ ;
  assign \new_[54865]_  = ~A201 & ~A166;
  assign \new_[54866]_  = A167 & \new_[54865]_ ;
  assign \new_[54867]_  = \new_[54866]_  & \new_[54861]_ ;
  assign \new_[54871]_  = ~A269 & ~A267;
  assign \new_[54872]_  = ~A203 & \new_[54871]_ ;
  assign \new_[54875]_  = ~A299 & A298;
  assign \new_[54878]_  = ~A302 & A300;
  assign \new_[54879]_  = \new_[54878]_  & \new_[54875]_ ;
  assign \new_[54880]_  = \new_[54879]_  & \new_[54872]_ ;
  assign \new_[54884]_  = ~A168 & ~A169;
  assign \new_[54885]_  = ~A170 & \new_[54884]_ ;
  assign \new_[54889]_  = ~A201 & ~A166;
  assign \new_[54890]_  = A167 & \new_[54889]_ ;
  assign \new_[54891]_  = \new_[54890]_  & \new_[54885]_ ;
  assign \new_[54895]_  = ~A269 & ~A267;
  assign \new_[54896]_  = ~A203 & \new_[54895]_ ;
  assign \new_[54899]_  = A299 & ~A298;
  assign \new_[54902]_  = A301 & A300;
  assign \new_[54903]_  = \new_[54902]_  & \new_[54899]_ ;
  assign \new_[54904]_  = \new_[54903]_  & \new_[54896]_ ;
  assign \new_[54908]_  = ~A168 & ~A169;
  assign \new_[54909]_  = ~A170 & \new_[54908]_ ;
  assign \new_[54913]_  = ~A201 & ~A166;
  assign \new_[54914]_  = A167 & \new_[54913]_ ;
  assign \new_[54915]_  = \new_[54914]_  & \new_[54909]_ ;
  assign \new_[54919]_  = ~A269 & ~A267;
  assign \new_[54920]_  = ~A203 & \new_[54919]_ ;
  assign \new_[54923]_  = A299 & ~A298;
  assign \new_[54926]_  = ~A302 & A300;
  assign \new_[54927]_  = \new_[54926]_  & \new_[54923]_ ;
  assign \new_[54928]_  = \new_[54927]_  & \new_[54920]_ ;
  assign \new_[54932]_  = ~A168 & ~A169;
  assign \new_[54933]_  = ~A170 & \new_[54932]_ ;
  assign \new_[54937]_  = ~A201 & ~A166;
  assign \new_[54938]_  = A167 & \new_[54937]_ ;
  assign \new_[54939]_  = \new_[54938]_  & \new_[54933]_ ;
  assign \new_[54943]_  = A266 & A265;
  assign \new_[54944]_  = ~A203 & \new_[54943]_ ;
  assign \new_[54947]_  = ~A299 & A298;
  assign \new_[54950]_  = A301 & A300;
  assign \new_[54951]_  = \new_[54950]_  & \new_[54947]_ ;
  assign \new_[54952]_  = \new_[54951]_  & \new_[54944]_ ;
  assign \new_[54956]_  = ~A168 & ~A169;
  assign \new_[54957]_  = ~A170 & \new_[54956]_ ;
  assign \new_[54961]_  = ~A201 & ~A166;
  assign \new_[54962]_  = A167 & \new_[54961]_ ;
  assign \new_[54963]_  = \new_[54962]_  & \new_[54957]_ ;
  assign \new_[54967]_  = A266 & A265;
  assign \new_[54968]_  = ~A203 & \new_[54967]_ ;
  assign \new_[54971]_  = ~A299 & A298;
  assign \new_[54974]_  = ~A302 & A300;
  assign \new_[54975]_  = \new_[54974]_  & \new_[54971]_ ;
  assign \new_[54976]_  = \new_[54975]_  & \new_[54968]_ ;
  assign \new_[54980]_  = ~A168 & ~A169;
  assign \new_[54981]_  = ~A170 & \new_[54980]_ ;
  assign \new_[54985]_  = ~A201 & ~A166;
  assign \new_[54986]_  = A167 & \new_[54985]_ ;
  assign \new_[54987]_  = \new_[54986]_  & \new_[54981]_ ;
  assign \new_[54991]_  = A266 & A265;
  assign \new_[54992]_  = ~A203 & \new_[54991]_ ;
  assign \new_[54995]_  = A299 & ~A298;
  assign \new_[54998]_  = A301 & A300;
  assign \new_[54999]_  = \new_[54998]_  & \new_[54995]_ ;
  assign \new_[55000]_  = \new_[54999]_  & \new_[54992]_ ;
  assign \new_[55004]_  = ~A168 & ~A169;
  assign \new_[55005]_  = ~A170 & \new_[55004]_ ;
  assign \new_[55009]_  = ~A201 & ~A166;
  assign \new_[55010]_  = A167 & \new_[55009]_ ;
  assign \new_[55011]_  = \new_[55010]_  & \new_[55005]_ ;
  assign \new_[55015]_  = A266 & A265;
  assign \new_[55016]_  = ~A203 & \new_[55015]_ ;
  assign \new_[55019]_  = A299 & ~A298;
  assign \new_[55022]_  = ~A302 & A300;
  assign \new_[55023]_  = \new_[55022]_  & \new_[55019]_ ;
  assign \new_[55024]_  = \new_[55023]_  & \new_[55016]_ ;
  assign \new_[55028]_  = ~A168 & ~A169;
  assign \new_[55029]_  = ~A170 & \new_[55028]_ ;
  assign \new_[55033]_  = ~A201 & ~A166;
  assign \new_[55034]_  = A167 & \new_[55033]_ ;
  assign \new_[55035]_  = \new_[55034]_  & \new_[55029]_ ;
  assign \new_[55039]_  = A266 & ~A265;
  assign \new_[55040]_  = ~A203 & \new_[55039]_ ;
  assign \new_[55043]_  = A268 & A267;
  assign \new_[55046]_  = A301 & ~A300;
  assign \new_[55047]_  = \new_[55046]_  & \new_[55043]_ ;
  assign \new_[55048]_  = \new_[55047]_  & \new_[55040]_ ;
  assign \new_[55052]_  = ~A168 & ~A169;
  assign \new_[55053]_  = ~A170 & \new_[55052]_ ;
  assign \new_[55057]_  = ~A201 & ~A166;
  assign \new_[55058]_  = A167 & \new_[55057]_ ;
  assign \new_[55059]_  = \new_[55058]_  & \new_[55053]_ ;
  assign \new_[55063]_  = A266 & ~A265;
  assign \new_[55064]_  = ~A203 & \new_[55063]_ ;
  assign \new_[55067]_  = A268 & A267;
  assign \new_[55070]_  = ~A302 & ~A300;
  assign \new_[55071]_  = \new_[55070]_  & \new_[55067]_ ;
  assign \new_[55072]_  = \new_[55071]_  & \new_[55064]_ ;
  assign \new_[55076]_  = ~A168 & ~A169;
  assign \new_[55077]_  = ~A170 & \new_[55076]_ ;
  assign \new_[55081]_  = ~A201 & ~A166;
  assign \new_[55082]_  = A167 & \new_[55081]_ ;
  assign \new_[55083]_  = \new_[55082]_  & \new_[55077]_ ;
  assign \new_[55087]_  = A266 & ~A265;
  assign \new_[55088]_  = ~A203 & \new_[55087]_ ;
  assign \new_[55091]_  = A268 & A267;
  assign \new_[55094]_  = A299 & A298;
  assign \new_[55095]_  = \new_[55094]_  & \new_[55091]_ ;
  assign \new_[55096]_  = \new_[55095]_  & \new_[55088]_ ;
  assign \new_[55100]_  = ~A168 & ~A169;
  assign \new_[55101]_  = ~A170 & \new_[55100]_ ;
  assign \new_[55105]_  = ~A201 & ~A166;
  assign \new_[55106]_  = A167 & \new_[55105]_ ;
  assign \new_[55107]_  = \new_[55106]_  & \new_[55101]_ ;
  assign \new_[55111]_  = A266 & ~A265;
  assign \new_[55112]_  = ~A203 & \new_[55111]_ ;
  assign \new_[55115]_  = A268 & A267;
  assign \new_[55118]_  = ~A299 & ~A298;
  assign \new_[55119]_  = \new_[55118]_  & \new_[55115]_ ;
  assign \new_[55120]_  = \new_[55119]_  & \new_[55112]_ ;
  assign \new_[55124]_  = ~A168 & ~A169;
  assign \new_[55125]_  = ~A170 & \new_[55124]_ ;
  assign \new_[55129]_  = ~A201 & ~A166;
  assign \new_[55130]_  = A167 & \new_[55129]_ ;
  assign \new_[55131]_  = \new_[55130]_  & \new_[55125]_ ;
  assign \new_[55135]_  = A266 & ~A265;
  assign \new_[55136]_  = ~A203 & \new_[55135]_ ;
  assign \new_[55139]_  = ~A269 & A267;
  assign \new_[55142]_  = A301 & ~A300;
  assign \new_[55143]_  = \new_[55142]_  & \new_[55139]_ ;
  assign \new_[55144]_  = \new_[55143]_  & \new_[55136]_ ;
  assign \new_[55148]_  = ~A168 & ~A169;
  assign \new_[55149]_  = ~A170 & \new_[55148]_ ;
  assign \new_[55153]_  = ~A201 & ~A166;
  assign \new_[55154]_  = A167 & \new_[55153]_ ;
  assign \new_[55155]_  = \new_[55154]_  & \new_[55149]_ ;
  assign \new_[55159]_  = A266 & ~A265;
  assign \new_[55160]_  = ~A203 & \new_[55159]_ ;
  assign \new_[55163]_  = ~A269 & A267;
  assign \new_[55166]_  = ~A302 & ~A300;
  assign \new_[55167]_  = \new_[55166]_  & \new_[55163]_ ;
  assign \new_[55168]_  = \new_[55167]_  & \new_[55160]_ ;
  assign \new_[55172]_  = ~A168 & ~A169;
  assign \new_[55173]_  = ~A170 & \new_[55172]_ ;
  assign \new_[55177]_  = ~A201 & ~A166;
  assign \new_[55178]_  = A167 & \new_[55177]_ ;
  assign \new_[55179]_  = \new_[55178]_  & \new_[55173]_ ;
  assign \new_[55183]_  = A266 & ~A265;
  assign \new_[55184]_  = ~A203 & \new_[55183]_ ;
  assign \new_[55187]_  = ~A269 & A267;
  assign \new_[55190]_  = A299 & A298;
  assign \new_[55191]_  = \new_[55190]_  & \new_[55187]_ ;
  assign \new_[55192]_  = \new_[55191]_  & \new_[55184]_ ;
  assign \new_[55196]_  = ~A168 & ~A169;
  assign \new_[55197]_  = ~A170 & \new_[55196]_ ;
  assign \new_[55201]_  = ~A201 & ~A166;
  assign \new_[55202]_  = A167 & \new_[55201]_ ;
  assign \new_[55203]_  = \new_[55202]_  & \new_[55197]_ ;
  assign \new_[55207]_  = A266 & ~A265;
  assign \new_[55208]_  = ~A203 & \new_[55207]_ ;
  assign \new_[55211]_  = ~A269 & A267;
  assign \new_[55214]_  = ~A299 & ~A298;
  assign \new_[55215]_  = \new_[55214]_  & \new_[55211]_ ;
  assign \new_[55216]_  = \new_[55215]_  & \new_[55208]_ ;
  assign \new_[55220]_  = ~A168 & ~A169;
  assign \new_[55221]_  = ~A170 & \new_[55220]_ ;
  assign \new_[55225]_  = ~A201 & ~A166;
  assign \new_[55226]_  = A167 & \new_[55225]_ ;
  assign \new_[55227]_  = \new_[55226]_  & \new_[55221]_ ;
  assign \new_[55231]_  = ~A266 & A265;
  assign \new_[55232]_  = ~A203 & \new_[55231]_ ;
  assign \new_[55235]_  = A268 & A267;
  assign \new_[55238]_  = A301 & ~A300;
  assign \new_[55239]_  = \new_[55238]_  & \new_[55235]_ ;
  assign \new_[55240]_  = \new_[55239]_  & \new_[55232]_ ;
  assign \new_[55244]_  = ~A168 & ~A169;
  assign \new_[55245]_  = ~A170 & \new_[55244]_ ;
  assign \new_[55249]_  = ~A201 & ~A166;
  assign \new_[55250]_  = A167 & \new_[55249]_ ;
  assign \new_[55251]_  = \new_[55250]_  & \new_[55245]_ ;
  assign \new_[55255]_  = ~A266 & A265;
  assign \new_[55256]_  = ~A203 & \new_[55255]_ ;
  assign \new_[55259]_  = A268 & A267;
  assign \new_[55262]_  = ~A302 & ~A300;
  assign \new_[55263]_  = \new_[55262]_  & \new_[55259]_ ;
  assign \new_[55264]_  = \new_[55263]_  & \new_[55256]_ ;
  assign \new_[55268]_  = ~A168 & ~A169;
  assign \new_[55269]_  = ~A170 & \new_[55268]_ ;
  assign \new_[55273]_  = ~A201 & ~A166;
  assign \new_[55274]_  = A167 & \new_[55273]_ ;
  assign \new_[55275]_  = \new_[55274]_  & \new_[55269]_ ;
  assign \new_[55279]_  = ~A266 & A265;
  assign \new_[55280]_  = ~A203 & \new_[55279]_ ;
  assign \new_[55283]_  = A268 & A267;
  assign \new_[55286]_  = A299 & A298;
  assign \new_[55287]_  = \new_[55286]_  & \new_[55283]_ ;
  assign \new_[55288]_  = \new_[55287]_  & \new_[55280]_ ;
  assign \new_[55292]_  = ~A168 & ~A169;
  assign \new_[55293]_  = ~A170 & \new_[55292]_ ;
  assign \new_[55297]_  = ~A201 & ~A166;
  assign \new_[55298]_  = A167 & \new_[55297]_ ;
  assign \new_[55299]_  = \new_[55298]_  & \new_[55293]_ ;
  assign \new_[55303]_  = ~A266 & A265;
  assign \new_[55304]_  = ~A203 & \new_[55303]_ ;
  assign \new_[55307]_  = A268 & A267;
  assign \new_[55310]_  = ~A299 & ~A298;
  assign \new_[55311]_  = \new_[55310]_  & \new_[55307]_ ;
  assign \new_[55312]_  = \new_[55311]_  & \new_[55304]_ ;
  assign \new_[55316]_  = ~A168 & ~A169;
  assign \new_[55317]_  = ~A170 & \new_[55316]_ ;
  assign \new_[55321]_  = ~A201 & ~A166;
  assign \new_[55322]_  = A167 & \new_[55321]_ ;
  assign \new_[55323]_  = \new_[55322]_  & \new_[55317]_ ;
  assign \new_[55327]_  = ~A266 & A265;
  assign \new_[55328]_  = ~A203 & \new_[55327]_ ;
  assign \new_[55331]_  = ~A269 & A267;
  assign \new_[55334]_  = A301 & ~A300;
  assign \new_[55335]_  = \new_[55334]_  & \new_[55331]_ ;
  assign \new_[55336]_  = \new_[55335]_  & \new_[55328]_ ;
  assign \new_[55340]_  = ~A168 & ~A169;
  assign \new_[55341]_  = ~A170 & \new_[55340]_ ;
  assign \new_[55345]_  = ~A201 & ~A166;
  assign \new_[55346]_  = A167 & \new_[55345]_ ;
  assign \new_[55347]_  = \new_[55346]_  & \new_[55341]_ ;
  assign \new_[55351]_  = ~A266 & A265;
  assign \new_[55352]_  = ~A203 & \new_[55351]_ ;
  assign \new_[55355]_  = ~A269 & A267;
  assign \new_[55358]_  = ~A302 & ~A300;
  assign \new_[55359]_  = \new_[55358]_  & \new_[55355]_ ;
  assign \new_[55360]_  = \new_[55359]_  & \new_[55352]_ ;
  assign \new_[55364]_  = ~A168 & ~A169;
  assign \new_[55365]_  = ~A170 & \new_[55364]_ ;
  assign \new_[55369]_  = ~A201 & ~A166;
  assign \new_[55370]_  = A167 & \new_[55369]_ ;
  assign \new_[55371]_  = \new_[55370]_  & \new_[55365]_ ;
  assign \new_[55375]_  = ~A266 & A265;
  assign \new_[55376]_  = ~A203 & \new_[55375]_ ;
  assign \new_[55379]_  = ~A269 & A267;
  assign \new_[55382]_  = A299 & A298;
  assign \new_[55383]_  = \new_[55382]_  & \new_[55379]_ ;
  assign \new_[55384]_  = \new_[55383]_  & \new_[55376]_ ;
  assign \new_[55388]_  = ~A168 & ~A169;
  assign \new_[55389]_  = ~A170 & \new_[55388]_ ;
  assign \new_[55393]_  = ~A201 & ~A166;
  assign \new_[55394]_  = A167 & \new_[55393]_ ;
  assign \new_[55395]_  = \new_[55394]_  & \new_[55389]_ ;
  assign \new_[55399]_  = ~A266 & A265;
  assign \new_[55400]_  = ~A203 & \new_[55399]_ ;
  assign \new_[55403]_  = ~A269 & A267;
  assign \new_[55406]_  = ~A299 & ~A298;
  assign \new_[55407]_  = \new_[55406]_  & \new_[55403]_ ;
  assign \new_[55408]_  = \new_[55407]_  & \new_[55400]_ ;
  assign \new_[55412]_  = ~A168 & ~A169;
  assign \new_[55413]_  = ~A170 & \new_[55412]_ ;
  assign \new_[55417]_  = ~A201 & ~A166;
  assign \new_[55418]_  = A167 & \new_[55417]_ ;
  assign \new_[55419]_  = \new_[55418]_  & \new_[55413]_ ;
  assign \new_[55423]_  = ~A266 & ~A265;
  assign \new_[55424]_  = ~A203 & \new_[55423]_ ;
  assign \new_[55427]_  = ~A299 & A298;
  assign \new_[55430]_  = A301 & A300;
  assign \new_[55431]_  = \new_[55430]_  & \new_[55427]_ ;
  assign \new_[55432]_  = \new_[55431]_  & \new_[55424]_ ;
  assign \new_[55436]_  = ~A168 & ~A169;
  assign \new_[55437]_  = ~A170 & \new_[55436]_ ;
  assign \new_[55441]_  = ~A201 & ~A166;
  assign \new_[55442]_  = A167 & \new_[55441]_ ;
  assign \new_[55443]_  = \new_[55442]_  & \new_[55437]_ ;
  assign \new_[55447]_  = ~A266 & ~A265;
  assign \new_[55448]_  = ~A203 & \new_[55447]_ ;
  assign \new_[55451]_  = ~A299 & A298;
  assign \new_[55454]_  = ~A302 & A300;
  assign \new_[55455]_  = \new_[55454]_  & \new_[55451]_ ;
  assign \new_[55456]_  = \new_[55455]_  & \new_[55448]_ ;
  assign \new_[55460]_  = ~A168 & ~A169;
  assign \new_[55461]_  = ~A170 & \new_[55460]_ ;
  assign \new_[55465]_  = ~A201 & ~A166;
  assign \new_[55466]_  = A167 & \new_[55465]_ ;
  assign \new_[55467]_  = \new_[55466]_  & \new_[55461]_ ;
  assign \new_[55471]_  = ~A266 & ~A265;
  assign \new_[55472]_  = ~A203 & \new_[55471]_ ;
  assign \new_[55475]_  = A299 & ~A298;
  assign \new_[55478]_  = A301 & A300;
  assign \new_[55479]_  = \new_[55478]_  & \new_[55475]_ ;
  assign \new_[55480]_  = \new_[55479]_  & \new_[55472]_ ;
  assign \new_[55484]_  = ~A168 & ~A169;
  assign \new_[55485]_  = ~A170 & \new_[55484]_ ;
  assign \new_[55489]_  = ~A201 & ~A166;
  assign \new_[55490]_  = A167 & \new_[55489]_ ;
  assign \new_[55491]_  = \new_[55490]_  & \new_[55485]_ ;
  assign \new_[55495]_  = ~A266 & ~A265;
  assign \new_[55496]_  = ~A203 & \new_[55495]_ ;
  assign \new_[55499]_  = A299 & ~A298;
  assign \new_[55502]_  = ~A302 & A300;
  assign \new_[55503]_  = \new_[55502]_  & \new_[55499]_ ;
  assign \new_[55504]_  = \new_[55503]_  & \new_[55496]_ ;
  assign \new_[55508]_  = ~A168 & ~A169;
  assign \new_[55509]_  = ~A170 & \new_[55508]_ ;
  assign \new_[55513]_  = A199 & ~A166;
  assign \new_[55514]_  = A167 & \new_[55513]_ ;
  assign \new_[55515]_  = \new_[55514]_  & \new_[55509]_ ;
  assign \new_[55519]_  = A268 & ~A267;
  assign \new_[55520]_  = A200 & \new_[55519]_ ;
  assign \new_[55523]_  = ~A299 & A298;
  assign \new_[55526]_  = A301 & A300;
  assign \new_[55527]_  = \new_[55526]_  & \new_[55523]_ ;
  assign \new_[55528]_  = \new_[55527]_  & \new_[55520]_ ;
  assign \new_[55532]_  = ~A168 & ~A169;
  assign \new_[55533]_  = ~A170 & \new_[55532]_ ;
  assign \new_[55537]_  = A199 & ~A166;
  assign \new_[55538]_  = A167 & \new_[55537]_ ;
  assign \new_[55539]_  = \new_[55538]_  & \new_[55533]_ ;
  assign \new_[55543]_  = A268 & ~A267;
  assign \new_[55544]_  = A200 & \new_[55543]_ ;
  assign \new_[55547]_  = ~A299 & A298;
  assign \new_[55550]_  = ~A302 & A300;
  assign \new_[55551]_  = \new_[55550]_  & \new_[55547]_ ;
  assign \new_[55552]_  = \new_[55551]_  & \new_[55544]_ ;
  assign \new_[55556]_  = ~A168 & ~A169;
  assign \new_[55557]_  = ~A170 & \new_[55556]_ ;
  assign \new_[55561]_  = A199 & ~A166;
  assign \new_[55562]_  = A167 & \new_[55561]_ ;
  assign \new_[55563]_  = \new_[55562]_  & \new_[55557]_ ;
  assign \new_[55567]_  = A268 & ~A267;
  assign \new_[55568]_  = A200 & \new_[55567]_ ;
  assign \new_[55571]_  = A299 & ~A298;
  assign \new_[55574]_  = A301 & A300;
  assign \new_[55575]_  = \new_[55574]_  & \new_[55571]_ ;
  assign \new_[55576]_  = \new_[55575]_  & \new_[55568]_ ;
  assign \new_[55580]_  = ~A168 & ~A169;
  assign \new_[55581]_  = ~A170 & \new_[55580]_ ;
  assign \new_[55585]_  = A199 & ~A166;
  assign \new_[55586]_  = A167 & \new_[55585]_ ;
  assign \new_[55587]_  = \new_[55586]_  & \new_[55581]_ ;
  assign \new_[55591]_  = A268 & ~A267;
  assign \new_[55592]_  = A200 & \new_[55591]_ ;
  assign \new_[55595]_  = A299 & ~A298;
  assign \new_[55598]_  = ~A302 & A300;
  assign \new_[55599]_  = \new_[55598]_  & \new_[55595]_ ;
  assign \new_[55600]_  = \new_[55599]_  & \new_[55592]_ ;
  assign \new_[55604]_  = ~A168 & ~A169;
  assign \new_[55605]_  = ~A170 & \new_[55604]_ ;
  assign \new_[55609]_  = A199 & ~A166;
  assign \new_[55610]_  = A167 & \new_[55609]_ ;
  assign \new_[55611]_  = \new_[55610]_  & \new_[55605]_ ;
  assign \new_[55615]_  = ~A269 & ~A267;
  assign \new_[55616]_  = A200 & \new_[55615]_ ;
  assign \new_[55619]_  = ~A299 & A298;
  assign \new_[55622]_  = A301 & A300;
  assign \new_[55623]_  = \new_[55622]_  & \new_[55619]_ ;
  assign \new_[55624]_  = \new_[55623]_  & \new_[55616]_ ;
  assign \new_[55628]_  = ~A168 & ~A169;
  assign \new_[55629]_  = ~A170 & \new_[55628]_ ;
  assign \new_[55633]_  = A199 & ~A166;
  assign \new_[55634]_  = A167 & \new_[55633]_ ;
  assign \new_[55635]_  = \new_[55634]_  & \new_[55629]_ ;
  assign \new_[55639]_  = ~A269 & ~A267;
  assign \new_[55640]_  = A200 & \new_[55639]_ ;
  assign \new_[55643]_  = ~A299 & A298;
  assign \new_[55646]_  = ~A302 & A300;
  assign \new_[55647]_  = \new_[55646]_  & \new_[55643]_ ;
  assign \new_[55648]_  = \new_[55647]_  & \new_[55640]_ ;
  assign \new_[55652]_  = ~A168 & ~A169;
  assign \new_[55653]_  = ~A170 & \new_[55652]_ ;
  assign \new_[55657]_  = A199 & ~A166;
  assign \new_[55658]_  = A167 & \new_[55657]_ ;
  assign \new_[55659]_  = \new_[55658]_  & \new_[55653]_ ;
  assign \new_[55663]_  = ~A269 & ~A267;
  assign \new_[55664]_  = A200 & \new_[55663]_ ;
  assign \new_[55667]_  = A299 & ~A298;
  assign \new_[55670]_  = A301 & A300;
  assign \new_[55671]_  = \new_[55670]_  & \new_[55667]_ ;
  assign \new_[55672]_  = \new_[55671]_  & \new_[55664]_ ;
  assign \new_[55676]_  = ~A168 & ~A169;
  assign \new_[55677]_  = ~A170 & \new_[55676]_ ;
  assign \new_[55681]_  = A199 & ~A166;
  assign \new_[55682]_  = A167 & \new_[55681]_ ;
  assign \new_[55683]_  = \new_[55682]_  & \new_[55677]_ ;
  assign \new_[55687]_  = ~A269 & ~A267;
  assign \new_[55688]_  = A200 & \new_[55687]_ ;
  assign \new_[55691]_  = A299 & ~A298;
  assign \new_[55694]_  = ~A302 & A300;
  assign \new_[55695]_  = \new_[55694]_  & \new_[55691]_ ;
  assign \new_[55696]_  = \new_[55695]_  & \new_[55688]_ ;
  assign \new_[55700]_  = ~A168 & ~A169;
  assign \new_[55701]_  = ~A170 & \new_[55700]_ ;
  assign \new_[55705]_  = A199 & ~A166;
  assign \new_[55706]_  = A167 & \new_[55705]_ ;
  assign \new_[55707]_  = \new_[55706]_  & \new_[55701]_ ;
  assign \new_[55711]_  = A266 & A265;
  assign \new_[55712]_  = A200 & \new_[55711]_ ;
  assign \new_[55715]_  = ~A299 & A298;
  assign \new_[55718]_  = A301 & A300;
  assign \new_[55719]_  = \new_[55718]_  & \new_[55715]_ ;
  assign \new_[55720]_  = \new_[55719]_  & \new_[55712]_ ;
  assign \new_[55724]_  = ~A168 & ~A169;
  assign \new_[55725]_  = ~A170 & \new_[55724]_ ;
  assign \new_[55729]_  = A199 & ~A166;
  assign \new_[55730]_  = A167 & \new_[55729]_ ;
  assign \new_[55731]_  = \new_[55730]_  & \new_[55725]_ ;
  assign \new_[55735]_  = A266 & A265;
  assign \new_[55736]_  = A200 & \new_[55735]_ ;
  assign \new_[55739]_  = ~A299 & A298;
  assign \new_[55742]_  = ~A302 & A300;
  assign \new_[55743]_  = \new_[55742]_  & \new_[55739]_ ;
  assign \new_[55744]_  = \new_[55743]_  & \new_[55736]_ ;
  assign \new_[55748]_  = ~A168 & ~A169;
  assign \new_[55749]_  = ~A170 & \new_[55748]_ ;
  assign \new_[55753]_  = A199 & ~A166;
  assign \new_[55754]_  = A167 & \new_[55753]_ ;
  assign \new_[55755]_  = \new_[55754]_  & \new_[55749]_ ;
  assign \new_[55759]_  = A266 & A265;
  assign \new_[55760]_  = A200 & \new_[55759]_ ;
  assign \new_[55763]_  = A299 & ~A298;
  assign \new_[55766]_  = A301 & A300;
  assign \new_[55767]_  = \new_[55766]_  & \new_[55763]_ ;
  assign \new_[55768]_  = \new_[55767]_  & \new_[55760]_ ;
  assign \new_[55772]_  = ~A168 & ~A169;
  assign \new_[55773]_  = ~A170 & \new_[55772]_ ;
  assign \new_[55777]_  = A199 & ~A166;
  assign \new_[55778]_  = A167 & \new_[55777]_ ;
  assign \new_[55779]_  = \new_[55778]_  & \new_[55773]_ ;
  assign \new_[55783]_  = A266 & A265;
  assign \new_[55784]_  = A200 & \new_[55783]_ ;
  assign \new_[55787]_  = A299 & ~A298;
  assign \new_[55790]_  = ~A302 & A300;
  assign \new_[55791]_  = \new_[55790]_  & \new_[55787]_ ;
  assign \new_[55792]_  = \new_[55791]_  & \new_[55784]_ ;
  assign \new_[55796]_  = ~A168 & ~A169;
  assign \new_[55797]_  = ~A170 & \new_[55796]_ ;
  assign \new_[55801]_  = A199 & ~A166;
  assign \new_[55802]_  = A167 & \new_[55801]_ ;
  assign \new_[55803]_  = \new_[55802]_  & \new_[55797]_ ;
  assign \new_[55807]_  = A266 & ~A265;
  assign \new_[55808]_  = A200 & \new_[55807]_ ;
  assign \new_[55811]_  = A268 & A267;
  assign \new_[55814]_  = A301 & ~A300;
  assign \new_[55815]_  = \new_[55814]_  & \new_[55811]_ ;
  assign \new_[55816]_  = \new_[55815]_  & \new_[55808]_ ;
  assign \new_[55820]_  = ~A168 & ~A169;
  assign \new_[55821]_  = ~A170 & \new_[55820]_ ;
  assign \new_[55825]_  = A199 & ~A166;
  assign \new_[55826]_  = A167 & \new_[55825]_ ;
  assign \new_[55827]_  = \new_[55826]_  & \new_[55821]_ ;
  assign \new_[55831]_  = A266 & ~A265;
  assign \new_[55832]_  = A200 & \new_[55831]_ ;
  assign \new_[55835]_  = A268 & A267;
  assign \new_[55838]_  = ~A302 & ~A300;
  assign \new_[55839]_  = \new_[55838]_  & \new_[55835]_ ;
  assign \new_[55840]_  = \new_[55839]_  & \new_[55832]_ ;
  assign \new_[55844]_  = ~A168 & ~A169;
  assign \new_[55845]_  = ~A170 & \new_[55844]_ ;
  assign \new_[55849]_  = A199 & ~A166;
  assign \new_[55850]_  = A167 & \new_[55849]_ ;
  assign \new_[55851]_  = \new_[55850]_  & \new_[55845]_ ;
  assign \new_[55855]_  = A266 & ~A265;
  assign \new_[55856]_  = A200 & \new_[55855]_ ;
  assign \new_[55859]_  = A268 & A267;
  assign \new_[55862]_  = A299 & A298;
  assign \new_[55863]_  = \new_[55862]_  & \new_[55859]_ ;
  assign \new_[55864]_  = \new_[55863]_  & \new_[55856]_ ;
  assign \new_[55868]_  = ~A168 & ~A169;
  assign \new_[55869]_  = ~A170 & \new_[55868]_ ;
  assign \new_[55873]_  = A199 & ~A166;
  assign \new_[55874]_  = A167 & \new_[55873]_ ;
  assign \new_[55875]_  = \new_[55874]_  & \new_[55869]_ ;
  assign \new_[55879]_  = A266 & ~A265;
  assign \new_[55880]_  = A200 & \new_[55879]_ ;
  assign \new_[55883]_  = A268 & A267;
  assign \new_[55886]_  = ~A299 & ~A298;
  assign \new_[55887]_  = \new_[55886]_  & \new_[55883]_ ;
  assign \new_[55888]_  = \new_[55887]_  & \new_[55880]_ ;
  assign \new_[55892]_  = ~A168 & ~A169;
  assign \new_[55893]_  = ~A170 & \new_[55892]_ ;
  assign \new_[55897]_  = A199 & ~A166;
  assign \new_[55898]_  = A167 & \new_[55897]_ ;
  assign \new_[55899]_  = \new_[55898]_  & \new_[55893]_ ;
  assign \new_[55903]_  = A266 & ~A265;
  assign \new_[55904]_  = A200 & \new_[55903]_ ;
  assign \new_[55907]_  = ~A269 & A267;
  assign \new_[55910]_  = A301 & ~A300;
  assign \new_[55911]_  = \new_[55910]_  & \new_[55907]_ ;
  assign \new_[55912]_  = \new_[55911]_  & \new_[55904]_ ;
  assign \new_[55916]_  = ~A168 & ~A169;
  assign \new_[55917]_  = ~A170 & \new_[55916]_ ;
  assign \new_[55921]_  = A199 & ~A166;
  assign \new_[55922]_  = A167 & \new_[55921]_ ;
  assign \new_[55923]_  = \new_[55922]_  & \new_[55917]_ ;
  assign \new_[55927]_  = A266 & ~A265;
  assign \new_[55928]_  = A200 & \new_[55927]_ ;
  assign \new_[55931]_  = ~A269 & A267;
  assign \new_[55934]_  = ~A302 & ~A300;
  assign \new_[55935]_  = \new_[55934]_  & \new_[55931]_ ;
  assign \new_[55936]_  = \new_[55935]_  & \new_[55928]_ ;
  assign \new_[55940]_  = ~A168 & ~A169;
  assign \new_[55941]_  = ~A170 & \new_[55940]_ ;
  assign \new_[55945]_  = A199 & ~A166;
  assign \new_[55946]_  = A167 & \new_[55945]_ ;
  assign \new_[55947]_  = \new_[55946]_  & \new_[55941]_ ;
  assign \new_[55951]_  = A266 & ~A265;
  assign \new_[55952]_  = A200 & \new_[55951]_ ;
  assign \new_[55955]_  = ~A269 & A267;
  assign \new_[55958]_  = A299 & A298;
  assign \new_[55959]_  = \new_[55958]_  & \new_[55955]_ ;
  assign \new_[55960]_  = \new_[55959]_  & \new_[55952]_ ;
  assign \new_[55964]_  = ~A168 & ~A169;
  assign \new_[55965]_  = ~A170 & \new_[55964]_ ;
  assign \new_[55969]_  = A199 & ~A166;
  assign \new_[55970]_  = A167 & \new_[55969]_ ;
  assign \new_[55971]_  = \new_[55970]_  & \new_[55965]_ ;
  assign \new_[55975]_  = A266 & ~A265;
  assign \new_[55976]_  = A200 & \new_[55975]_ ;
  assign \new_[55979]_  = ~A269 & A267;
  assign \new_[55982]_  = ~A299 & ~A298;
  assign \new_[55983]_  = \new_[55982]_  & \new_[55979]_ ;
  assign \new_[55984]_  = \new_[55983]_  & \new_[55976]_ ;
  assign \new_[55988]_  = ~A168 & ~A169;
  assign \new_[55989]_  = ~A170 & \new_[55988]_ ;
  assign \new_[55993]_  = A199 & ~A166;
  assign \new_[55994]_  = A167 & \new_[55993]_ ;
  assign \new_[55995]_  = \new_[55994]_  & \new_[55989]_ ;
  assign \new_[55999]_  = ~A266 & A265;
  assign \new_[56000]_  = A200 & \new_[55999]_ ;
  assign \new_[56003]_  = A268 & A267;
  assign \new_[56006]_  = A301 & ~A300;
  assign \new_[56007]_  = \new_[56006]_  & \new_[56003]_ ;
  assign \new_[56008]_  = \new_[56007]_  & \new_[56000]_ ;
  assign \new_[56012]_  = ~A168 & ~A169;
  assign \new_[56013]_  = ~A170 & \new_[56012]_ ;
  assign \new_[56017]_  = A199 & ~A166;
  assign \new_[56018]_  = A167 & \new_[56017]_ ;
  assign \new_[56019]_  = \new_[56018]_  & \new_[56013]_ ;
  assign \new_[56023]_  = ~A266 & A265;
  assign \new_[56024]_  = A200 & \new_[56023]_ ;
  assign \new_[56027]_  = A268 & A267;
  assign \new_[56030]_  = ~A302 & ~A300;
  assign \new_[56031]_  = \new_[56030]_  & \new_[56027]_ ;
  assign \new_[56032]_  = \new_[56031]_  & \new_[56024]_ ;
  assign \new_[56036]_  = ~A168 & ~A169;
  assign \new_[56037]_  = ~A170 & \new_[56036]_ ;
  assign \new_[56041]_  = A199 & ~A166;
  assign \new_[56042]_  = A167 & \new_[56041]_ ;
  assign \new_[56043]_  = \new_[56042]_  & \new_[56037]_ ;
  assign \new_[56047]_  = ~A266 & A265;
  assign \new_[56048]_  = A200 & \new_[56047]_ ;
  assign \new_[56051]_  = A268 & A267;
  assign \new_[56054]_  = A299 & A298;
  assign \new_[56055]_  = \new_[56054]_  & \new_[56051]_ ;
  assign \new_[56056]_  = \new_[56055]_  & \new_[56048]_ ;
  assign \new_[56060]_  = ~A168 & ~A169;
  assign \new_[56061]_  = ~A170 & \new_[56060]_ ;
  assign \new_[56065]_  = A199 & ~A166;
  assign \new_[56066]_  = A167 & \new_[56065]_ ;
  assign \new_[56067]_  = \new_[56066]_  & \new_[56061]_ ;
  assign \new_[56071]_  = ~A266 & A265;
  assign \new_[56072]_  = A200 & \new_[56071]_ ;
  assign \new_[56075]_  = A268 & A267;
  assign \new_[56078]_  = ~A299 & ~A298;
  assign \new_[56079]_  = \new_[56078]_  & \new_[56075]_ ;
  assign \new_[56080]_  = \new_[56079]_  & \new_[56072]_ ;
  assign \new_[56084]_  = ~A168 & ~A169;
  assign \new_[56085]_  = ~A170 & \new_[56084]_ ;
  assign \new_[56089]_  = A199 & ~A166;
  assign \new_[56090]_  = A167 & \new_[56089]_ ;
  assign \new_[56091]_  = \new_[56090]_  & \new_[56085]_ ;
  assign \new_[56095]_  = ~A266 & A265;
  assign \new_[56096]_  = A200 & \new_[56095]_ ;
  assign \new_[56099]_  = ~A269 & A267;
  assign \new_[56102]_  = A301 & ~A300;
  assign \new_[56103]_  = \new_[56102]_  & \new_[56099]_ ;
  assign \new_[56104]_  = \new_[56103]_  & \new_[56096]_ ;
  assign \new_[56108]_  = ~A168 & ~A169;
  assign \new_[56109]_  = ~A170 & \new_[56108]_ ;
  assign \new_[56113]_  = A199 & ~A166;
  assign \new_[56114]_  = A167 & \new_[56113]_ ;
  assign \new_[56115]_  = \new_[56114]_  & \new_[56109]_ ;
  assign \new_[56119]_  = ~A266 & A265;
  assign \new_[56120]_  = A200 & \new_[56119]_ ;
  assign \new_[56123]_  = ~A269 & A267;
  assign \new_[56126]_  = ~A302 & ~A300;
  assign \new_[56127]_  = \new_[56126]_  & \new_[56123]_ ;
  assign \new_[56128]_  = \new_[56127]_  & \new_[56120]_ ;
  assign \new_[56132]_  = ~A168 & ~A169;
  assign \new_[56133]_  = ~A170 & \new_[56132]_ ;
  assign \new_[56137]_  = A199 & ~A166;
  assign \new_[56138]_  = A167 & \new_[56137]_ ;
  assign \new_[56139]_  = \new_[56138]_  & \new_[56133]_ ;
  assign \new_[56143]_  = ~A266 & A265;
  assign \new_[56144]_  = A200 & \new_[56143]_ ;
  assign \new_[56147]_  = ~A269 & A267;
  assign \new_[56150]_  = A299 & A298;
  assign \new_[56151]_  = \new_[56150]_  & \new_[56147]_ ;
  assign \new_[56152]_  = \new_[56151]_  & \new_[56144]_ ;
  assign \new_[56156]_  = ~A168 & ~A169;
  assign \new_[56157]_  = ~A170 & \new_[56156]_ ;
  assign \new_[56161]_  = A199 & ~A166;
  assign \new_[56162]_  = A167 & \new_[56161]_ ;
  assign \new_[56163]_  = \new_[56162]_  & \new_[56157]_ ;
  assign \new_[56167]_  = ~A266 & A265;
  assign \new_[56168]_  = A200 & \new_[56167]_ ;
  assign \new_[56171]_  = ~A269 & A267;
  assign \new_[56174]_  = ~A299 & ~A298;
  assign \new_[56175]_  = \new_[56174]_  & \new_[56171]_ ;
  assign \new_[56176]_  = \new_[56175]_  & \new_[56168]_ ;
  assign \new_[56180]_  = ~A168 & ~A169;
  assign \new_[56181]_  = ~A170 & \new_[56180]_ ;
  assign \new_[56185]_  = A199 & ~A166;
  assign \new_[56186]_  = A167 & \new_[56185]_ ;
  assign \new_[56187]_  = \new_[56186]_  & \new_[56181]_ ;
  assign \new_[56191]_  = ~A266 & ~A265;
  assign \new_[56192]_  = A200 & \new_[56191]_ ;
  assign \new_[56195]_  = ~A299 & A298;
  assign \new_[56198]_  = A301 & A300;
  assign \new_[56199]_  = \new_[56198]_  & \new_[56195]_ ;
  assign \new_[56200]_  = \new_[56199]_  & \new_[56192]_ ;
  assign \new_[56204]_  = ~A168 & ~A169;
  assign \new_[56205]_  = ~A170 & \new_[56204]_ ;
  assign \new_[56209]_  = A199 & ~A166;
  assign \new_[56210]_  = A167 & \new_[56209]_ ;
  assign \new_[56211]_  = \new_[56210]_  & \new_[56205]_ ;
  assign \new_[56215]_  = ~A266 & ~A265;
  assign \new_[56216]_  = A200 & \new_[56215]_ ;
  assign \new_[56219]_  = ~A299 & A298;
  assign \new_[56222]_  = ~A302 & A300;
  assign \new_[56223]_  = \new_[56222]_  & \new_[56219]_ ;
  assign \new_[56224]_  = \new_[56223]_  & \new_[56216]_ ;
  assign \new_[56228]_  = ~A168 & ~A169;
  assign \new_[56229]_  = ~A170 & \new_[56228]_ ;
  assign \new_[56233]_  = A199 & ~A166;
  assign \new_[56234]_  = A167 & \new_[56233]_ ;
  assign \new_[56235]_  = \new_[56234]_  & \new_[56229]_ ;
  assign \new_[56239]_  = ~A266 & ~A265;
  assign \new_[56240]_  = A200 & \new_[56239]_ ;
  assign \new_[56243]_  = A299 & ~A298;
  assign \new_[56246]_  = A301 & A300;
  assign \new_[56247]_  = \new_[56246]_  & \new_[56243]_ ;
  assign \new_[56248]_  = \new_[56247]_  & \new_[56240]_ ;
  assign \new_[56252]_  = ~A168 & ~A169;
  assign \new_[56253]_  = ~A170 & \new_[56252]_ ;
  assign \new_[56257]_  = A199 & ~A166;
  assign \new_[56258]_  = A167 & \new_[56257]_ ;
  assign \new_[56259]_  = \new_[56258]_  & \new_[56253]_ ;
  assign \new_[56263]_  = ~A266 & ~A265;
  assign \new_[56264]_  = A200 & \new_[56263]_ ;
  assign \new_[56267]_  = A299 & ~A298;
  assign \new_[56270]_  = ~A302 & A300;
  assign \new_[56271]_  = \new_[56270]_  & \new_[56267]_ ;
  assign \new_[56272]_  = \new_[56271]_  & \new_[56264]_ ;
  assign \new_[56276]_  = ~A168 & ~A169;
  assign \new_[56277]_  = ~A170 & \new_[56276]_ ;
  assign \new_[56281]_  = ~A199 & ~A166;
  assign \new_[56282]_  = A167 & \new_[56281]_ ;
  assign \new_[56283]_  = \new_[56282]_  & \new_[56277]_ ;
  assign \new_[56287]_  = A268 & ~A267;
  assign \new_[56288]_  = ~A200 & \new_[56287]_ ;
  assign \new_[56291]_  = ~A299 & A298;
  assign \new_[56294]_  = A301 & A300;
  assign \new_[56295]_  = \new_[56294]_  & \new_[56291]_ ;
  assign \new_[56296]_  = \new_[56295]_  & \new_[56288]_ ;
  assign \new_[56300]_  = ~A168 & ~A169;
  assign \new_[56301]_  = ~A170 & \new_[56300]_ ;
  assign \new_[56305]_  = ~A199 & ~A166;
  assign \new_[56306]_  = A167 & \new_[56305]_ ;
  assign \new_[56307]_  = \new_[56306]_  & \new_[56301]_ ;
  assign \new_[56311]_  = A268 & ~A267;
  assign \new_[56312]_  = ~A200 & \new_[56311]_ ;
  assign \new_[56315]_  = ~A299 & A298;
  assign \new_[56318]_  = ~A302 & A300;
  assign \new_[56319]_  = \new_[56318]_  & \new_[56315]_ ;
  assign \new_[56320]_  = \new_[56319]_  & \new_[56312]_ ;
  assign \new_[56324]_  = ~A168 & ~A169;
  assign \new_[56325]_  = ~A170 & \new_[56324]_ ;
  assign \new_[56329]_  = ~A199 & ~A166;
  assign \new_[56330]_  = A167 & \new_[56329]_ ;
  assign \new_[56331]_  = \new_[56330]_  & \new_[56325]_ ;
  assign \new_[56335]_  = A268 & ~A267;
  assign \new_[56336]_  = ~A200 & \new_[56335]_ ;
  assign \new_[56339]_  = A299 & ~A298;
  assign \new_[56342]_  = A301 & A300;
  assign \new_[56343]_  = \new_[56342]_  & \new_[56339]_ ;
  assign \new_[56344]_  = \new_[56343]_  & \new_[56336]_ ;
  assign \new_[56348]_  = ~A168 & ~A169;
  assign \new_[56349]_  = ~A170 & \new_[56348]_ ;
  assign \new_[56353]_  = ~A199 & ~A166;
  assign \new_[56354]_  = A167 & \new_[56353]_ ;
  assign \new_[56355]_  = \new_[56354]_  & \new_[56349]_ ;
  assign \new_[56359]_  = A268 & ~A267;
  assign \new_[56360]_  = ~A200 & \new_[56359]_ ;
  assign \new_[56363]_  = A299 & ~A298;
  assign \new_[56366]_  = ~A302 & A300;
  assign \new_[56367]_  = \new_[56366]_  & \new_[56363]_ ;
  assign \new_[56368]_  = \new_[56367]_  & \new_[56360]_ ;
  assign \new_[56372]_  = ~A168 & ~A169;
  assign \new_[56373]_  = ~A170 & \new_[56372]_ ;
  assign \new_[56377]_  = ~A199 & ~A166;
  assign \new_[56378]_  = A167 & \new_[56377]_ ;
  assign \new_[56379]_  = \new_[56378]_  & \new_[56373]_ ;
  assign \new_[56383]_  = ~A269 & ~A267;
  assign \new_[56384]_  = ~A200 & \new_[56383]_ ;
  assign \new_[56387]_  = ~A299 & A298;
  assign \new_[56390]_  = A301 & A300;
  assign \new_[56391]_  = \new_[56390]_  & \new_[56387]_ ;
  assign \new_[56392]_  = \new_[56391]_  & \new_[56384]_ ;
  assign \new_[56396]_  = ~A168 & ~A169;
  assign \new_[56397]_  = ~A170 & \new_[56396]_ ;
  assign \new_[56401]_  = ~A199 & ~A166;
  assign \new_[56402]_  = A167 & \new_[56401]_ ;
  assign \new_[56403]_  = \new_[56402]_  & \new_[56397]_ ;
  assign \new_[56407]_  = ~A269 & ~A267;
  assign \new_[56408]_  = ~A200 & \new_[56407]_ ;
  assign \new_[56411]_  = ~A299 & A298;
  assign \new_[56414]_  = ~A302 & A300;
  assign \new_[56415]_  = \new_[56414]_  & \new_[56411]_ ;
  assign \new_[56416]_  = \new_[56415]_  & \new_[56408]_ ;
  assign \new_[56420]_  = ~A168 & ~A169;
  assign \new_[56421]_  = ~A170 & \new_[56420]_ ;
  assign \new_[56425]_  = ~A199 & ~A166;
  assign \new_[56426]_  = A167 & \new_[56425]_ ;
  assign \new_[56427]_  = \new_[56426]_  & \new_[56421]_ ;
  assign \new_[56431]_  = ~A269 & ~A267;
  assign \new_[56432]_  = ~A200 & \new_[56431]_ ;
  assign \new_[56435]_  = A299 & ~A298;
  assign \new_[56438]_  = A301 & A300;
  assign \new_[56439]_  = \new_[56438]_  & \new_[56435]_ ;
  assign \new_[56440]_  = \new_[56439]_  & \new_[56432]_ ;
  assign \new_[56444]_  = ~A168 & ~A169;
  assign \new_[56445]_  = ~A170 & \new_[56444]_ ;
  assign \new_[56449]_  = ~A199 & ~A166;
  assign \new_[56450]_  = A167 & \new_[56449]_ ;
  assign \new_[56451]_  = \new_[56450]_  & \new_[56445]_ ;
  assign \new_[56455]_  = ~A269 & ~A267;
  assign \new_[56456]_  = ~A200 & \new_[56455]_ ;
  assign \new_[56459]_  = A299 & ~A298;
  assign \new_[56462]_  = ~A302 & A300;
  assign \new_[56463]_  = \new_[56462]_  & \new_[56459]_ ;
  assign \new_[56464]_  = \new_[56463]_  & \new_[56456]_ ;
  assign \new_[56468]_  = ~A168 & ~A169;
  assign \new_[56469]_  = ~A170 & \new_[56468]_ ;
  assign \new_[56473]_  = ~A199 & ~A166;
  assign \new_[56474]_  = A167 & \new_[56473]_ ;
  assign \new_[56475]_  = \new_[56474]_  & \new_[56469]_ ;
  assign \new_[56479]_  = A266 & A265;
  assign \new_[56480]_  = ~A200 & \new_[56479]_ ;
  assign \new_[56483]_  = ~A299 & A298;
  assign \new_[56486]_  = A301 & A300;
  assign \new_[56487]_  = \new_[56486]_  & \new_[56483]_ ;
  assign \new_[56488]_  = \new_[56487]_  & \new_[56480]_ ;
  assign \new_[56492]_  = ~A168 & ~A169;
  assign \new_[56493]_  = ~A170 & \new_[56492]_ ;
  assign \new_[56497]_  = ~A199 & ~A166;
  assign \new_[56498]_  = A167 & \new_[56497]_ ;
  assign \new_[56499]_  = \new_[56498]_  & \new_[56493]_ ;
  assign \new_[56503]_  = A266 & A265;
  assign \new_[56504]_  = ~A200 & \new_[56503]_ ;
  assign \new_[56507]_  = ~A299 & A298;
  assign \new_[56510]_  = ~A302 & A300;
  assign \new_[56511]_  = \new_[56510]_  & \new_[56507]_ ;
  assign \new_[56512]_  = \new_[56511]_  & \new_[56504]_ ;
  assign \new_[56516]_  = ~A168 & ~A169;
  assign \new_[56517]_  = ~A170 & \new_[56516]_ ;
  assign \new_[56521]_  = ~A199 & ~A166;
  assign \new_[56522]_  = A167 & \new_[56521]_ ;
  assign \new_[56523]_  = \new_[56522]_  & \new_[56517]_ ;
  assign \new_[56527]_  = A266 & A265;
  assign \new_[56528]_  = ~A200 & \new_[56527]_ ;
  assign \new_[56531]_  = A299 & ~A298;
  assign \new_[56534]_  = A301 & A300;
  assign \new_[56535]_  = \new_[56534]_  & \new_[56531]_ ;
  assign \new_[56536]_  = \new_[56535]_  & \new_[56528]_ ;
  assign \new_[56540]_  = ~A168 & ~A169;
  assign \new_[56541]_  = ~A170 & \new_[56540]_ ;
  assign \new_[56545]_  = ~A199 & ~A166;
  assign \new_[56546]_  = A167 & \new_[56545]_ ;
  assign \new_[56547]_  = \new_[56546]_  & \new_[56541]_ ;
  assign \new_[56551]_  = A266 & A265;
  assign \new_[56552]_  = ~A200 & \new_[56551]_ ;
  assign \new_[56555]_  = A299 & ~A298;
  assign \new_[56558]_  = ~A302 & A300;
  assign \new_[56559]_  = \new_[56558]_  & \new_[56555]_ ;
  assign \new_[56560]_  = \new_[56559]_  & \new_[56552]_ ;
  assign \new_[56564]_  = ~A168 & ~A169;
  assign \new_[56565]_  = ~A170 & \new_[56564]_ ;
  assign \new_[56569]_  = ~A199 & ~A166;
  assign \new_[56570]_  = A167 & \new_[56569]_ ;
  assign \new_[56571]_  = \new_[56570]_  & \new_[56565]_ ;
  assign \new_[56575]_  = A266 & ~A265;
  assign \new_[56576]_  = ~A200 & \new_[56575]_ ;
  assign \new_[56579]_  = A268 & A267;
  assign \new_[56582]_  = A301 & ~A300;
  assign \new_[56583]_  = \new_[56582]_  & \new_[56579]_ ;
  assign \new_[56584]_  = \new_[56583]_  & \new_[56576]_ ;
  assign \new_[56588]_  = ~A168 & ~A169;
  assign \new_[56589]_  = ~A170 & \new_[56588]_ ;
  assign \new_[56593]_  = ~A199 & ~A166;
  assign \new_[56594]_  = A167 & \new_[56593]_ ;
  assign \new_[56595]_  = \new_[56594]_  & \new_[56589]_ ;
  assign \new_[56599]_  = A266 & ~A265;
  assign \new_[56600]_  = ~A200 & \new_[56599]_ ;
  assign \new_[56603]_  = A268 & A267;
  assign \new_[56606]_  = ~A302 & ~A300;
  assign \new_[56607]_  = \new_[56606]_  & \new_[56603]_ ;
  assign \new_[56608]_  = \new_[56607]_  & \new_[56600]_ ;
  assign \new_[56612]_  = ~A168 & ~A169;
  assign \new_[56613]_  = ~A170 & \new_[56612]_ ;
  assign \new_[56617]_  = ~A199 & ~A166;
  assign \new_[56618]_  = A167 & \new_[56617]_ ;
  assign \new_[56619]_  = \new_[56618]_  & \new_[56613]_ ;
  assign \new_[56623]_  = A266 & ~A265;
  assign \new_[56624]_  = ~A200 & \new_[56623]_ ;
  assign \new_[56627]_  = A268 & A267;
  assign \new_[56630]_  = A299 & A298;
  assign \new_[56631]_  = \new_[56630]_  & \new_[56627]_ ;
  assign \new_[56632]_  = \new_[56631]_  & \new_[56624]_ ;
  assign \new_[56636]_  = ~A168 & ~A169;
  assign \new_[56637]_  = ~A170 & \new_[56636]_ ;
  assign \new_[56641]_  = ~A199 & ~A166;
  assign \new_[56642]_  = A167 & \new_[56641]_ ;
  assign \new_[56643]_  = \new_[56642]_  & \new_[56637]_ ;
  assign \new_[56647]_  = A266 & ~A265;
  assign \new_[56648]_  = ~A200 & \new_[56647]_ ;
  assign \new_[56651]_  = A268 & A267;
  assign \new_[56654]_  = ~A299 & ~A298;
  assign \new_[56655]_  = \new_[56654]_  & \new_[56651]_ ;
  assign \new_[56656]_  = \new_[56655]_  & \new_[56648]_ ;
  assign \new_[56660]_  = ~A168 & ~A169;
  assign \new_[56661]_  = ~A170 & \new_[56660]_ ;
  assign \new_[56665]_  = ~A199 & ~A166;
  assign \new_[56666]_  = A167 & \new_[56665]_ ;
  assign \new_[56667]_  = \new_[56666]_  & \new_[56661]_ ;
  assign \new_[56671]_  = A266 & ~A265;
  assign \new_[56672]_  = ~A200 & \new_[56671]_ ;
  assign \new_[56675]_  = ~A269 & A267;
  assign \new_[56678]_  = A301 & ~A300;
  assign \new_[56679]_  = \new_[56678]_  & \new_[56675]_ ;
  assign \new_[56680]_  = \new_[56679]_  & \new_[56672]_ ;
  assign \new_[56684]_  = ~A168 & ~A169;
  assign \new_[56685]_  = ~A170 & \new_[56684]_ ;
  assign \new_[56689]_  = ~A199 & ~A166;
  assign \new_[56690]_  = A167 & \new_[56689]_ ;
  assign \new_[56691]_  = \new_[56690]_  & \new_[56685]_ ;
  assign \new_[56695]_  = A266 & ~A265;
  assign \new_[56696]_  = ~A200 & \new_[56695]_ ;
  assign \new_[56699]_  = ~A269 & A267;
  assign \new_[56702]_  = ~A302 & ~A300;
  assign \new_[56703]_  = \new_[56702]_  & \new_[56699]_ ;
  assign \new_[56704]_  = \new_[56703]_  & \new_[56696]_ ;
  assign \new_[56708]_  = ~A168 & ~A169;
  assign \new_[56709]_  = ~A170 & \new_[56708]_ ;
  assign \new_[56713]_  = ~A199 & ~A166;
  assign \new_[56714]_  = A167 & \new_[56713]_ ;
  assign \new_[56715]_  = \new_[56714]_  & \new_[56709]_ ;
  assign \new_[56719]_  = A266 & ~A265;
  assign \new_[56720]_  = ~A200 & \new_[56719]_ ;
  assign \new_[56723]_  = ~A269 & A267;
  assign \new_[56726]_  = A299 & A298;
  assign \new_[56727]_  = \new_[56726]_  & \new_[56723]_ ;
  assign \new_[56728]_  = \new_[56727]_  & \new_[56720]_ ;
  assign \new_[56732]_  = ~A168 & ~A169;
  assign \new_[56733]_  = ~A170 & \new_[56732]_ ;
  assign \new_[56737]_  = ~A199 & ~A166;
  assign \new_[56738]_  = A167 & \new_[56737]_ ;
  assign \new_[56739]_  = \new_[56738]_  & \new_[56733]_ ;
  assign \new_[56743]_  = A266 & ~A265;
  assign \new_[56744]_  = ~A200 & \new_[56743]_ ;
  assign \new_[56747]_  = ~A269 & A267;
  assign \new_[56750]_  = ~A299 & ~A298;
  assign \new_[56751]_  = \new_[56750]_  & \new_[56747]_ ;
  assign \new_[56752]_  = \new_[56751]_  & \new_[56744]_ ;
  assign \new_[56756]_  = ~A168 & ~A169;
  assign \new_[56757]_  = ~A170 & \new_[56756]_ ;
  assign \new_[56761]_  = ~A199 & ~A166;
  assign \new_[56762]_  = A167 & \new_[56761]_ ;
  assign \new_[56763]_  = \new_[56762]_  & \new_[56757]_ ;
  assign \new_[56767]_  = ~A266 & A265;
  assign \new_[56768]_  = ~A200 & \new_[56767]_ ;
  assign \new_[56771]_  = A268 & A267;
  assign \new_[56774]_  = A301 & ~A300;
  assign \new_[56775]_  = \new_[56774]_  & \new_[56771]_ ;
  assign \new_[56776]_  = \new_[56775]_  & \new_[56768]_ ;
  assign \new_[56780]_  = ~A168 & ~A169;
  assign \new_[56781]_  = ~A170 & \new_[56780]_ ;
  assign \new_[56785]_  = ~A199 & ~A166;
  assign \new_[56786]_  = A167 & \new_[56785]_ ;
  assign \new_[56787]_  = \new_[56786]_  & \new_[56781]_ ;
  assign \new_[56791]_  = ~A266 & A265;
  assign \new_[56792]_  = ~A200 & \new_[56791]_ ;
  assign \new_[56795]_  = A268 & A267;
  assign \new_[56798]_  = ~A302 & ~A300;
  assign \new_[56799]_  = \new_[56798]_  & \new_[56795]_ ;
  assign \new_[56800]_  = \new_[56799]_  & \new_[56792]_ ;
  assign \new_[56804]_  = ~A168 & ~A169;
  assign \new_[56805]_  = ~A170 & \new_[56804]_ ;
  assign \new_[56809]_  = ~A199 & ~A166;
  assign \new_[56810]_  = A167 & \new_[56809]_ ;
  assign \new_[56811]_  = \new_[56810]_  & \new_[56805]_ ;
  assign \new_[56815]_  = ~A266 & A265;
  assign \new_[56816]_  = ~A200 & \new_[56815]_ ;
  assign \new_[56819]_  = A268 & A267;
  assign \new_[56822]_  = A299 & A298;
  assign \new_[56823]_  = \new_[56822]_  & \new_[56819]_ ;
  assign \new_[56824]_  = \new_[56823]_  & \new_[56816]_ ;
  assign \new_[56828]_  = ~A168 & ~A169;
  assign \new_[56829]_  = ~A170 & \new_[56828]_ ;
  assign \new_[56833]_  = ~A199 & ~A166;
  assign \new_[56834]_  = A167 & \new_[56833]_ ;
  assign \new_[56835]_  = \new_[56834]_  & \new_[56829]_ ;
  assign \new_[56839]_  = ~A266 & A265;
  assign \new_[56840]_  = ~A200 & \new_[56839]_ ;
  assign \new_[56843]_  = A268 & A267;
  assign \new_[56846]_  = ~A299 & ~A298;
  assign \new_[56847]_  = \new_[56846]_  & \new_[56843]_ ;
  assign \new_[56848]_  = \new_[56847]_  & \new_[56840]_ ;
  assign \new_[56852]_  = ~A168 & ~A169;
  assign \new_[56853]_  = ~A170 & \new_[56852]_ ;
  assign \new_[56857]_  = ~A199 & ~A166;
  assign \new_[56858]_  = A167 & \new_[56857]_ ;
  assign \new_[56859]_  = \new_[56858]_  & \new_[56853]_ ;
  assign \new_[56863]_  = ~A266 & A265;
  assign \new_[56864]_  = ~A200 & \new_[56863]_ ;
  assign \new_[56867]_  = ~A269 & A267;
  assign \new_[56870]_  = A301 & ~A300;
  assign \new_[56871]_  = \new_[56870]_  & \new_[56867]_ ;
  assign \new_[56872]_  = \new_[56871]_  & \new_[56864]_ ;
  assign \new_[56876]_  = ~A168 & ~A169;
  assign \new_[56877]_  = ~A170 & \new_[56876]_ ;
  assign \new_[56881]_  = ~A199 & ~A166;
  assign \new_[56882]_  = A167 & \new_[56881]_ ;
  assign \new_[56883]_  = \new_[56882]_  & \new_[56877]_ ;
  assign \new_[56887]_  = ~A266 & A265;
  assign \new_[56888]_  = ~A200 & \new_[56887]_ ;
  assign \new_[56891]_  = ~A269 & A267;
  assign \new_[56894]_  = ~A302 & ~A300;
  assign \new_[56895]_  = \new_[56894]_  & \new_[56891]_ ;
  assign \new_[56896]_  = \new_[56895]_  & \new_[56888]_ ;
  assign \new_[56900]_  = ~A168 & ~A169;
  assign \new_[56901]_  = ~A170 & \new_[56900]_ ;
  assign \new_[56905]_  = ~A199 & ~A166;
  assign \new_[56906]_  = A167 & \new_[56905]_ ;
  assign \new_[56907]_  = \new_[56906]_  & \new_[56901]_ ;
  assign \new_[56911]_  = ~A266 & A265;
  assign \new_[56912]_  = ~A200 & \new_[56911]_ ;
  assign \new_[56915]_  = ~A269 & A267;
  assign \new_[56918]_  = A299 & A298;
  assign \new_[56919]_  = \new_[56918]_  & \new_[56915]_ ;
  assign \new_[56920]_  = \new_[56919]_  & \new_[56912]_ ;
  assign \new_[56924]_  = ~A168 & ~A169;
  assign \new_[56925]_  = ~A170 & \new_[56924]_ ;
  assign \new_[56929]_  = ~A199 & ~A166;
  assign \new_[56930]_  = A167 & \new_[56929]_ ;
  assign \new_[56931]_  = \new_[56930]_  & \new_[56925]_ ;
  assign \new_[56935]_  = ~A266 & A265;
  assign \new_[56936]_  = ~A200 & \new_[56935]_ ;
  assign \new_[56939]_  = ~A269 & A267;
  assign \new_[56942]_  = ~A299 & ~A298;
  assign \new_[56943]_  = \new_[56942]_  & \new_[56939]_ ;
  assign \new_[56944]_  = \new_[56943]_  & \new_[56936]_ ;
  assign \new_[56948]_  = ~A168 & ~A169;
  assign \new_[56949]_  = ~A170 & \new_[56948]_ ;
  assign \new_[56953]_  = ~A199 & ~A166;
  assign \new_[56954]_  = A167 & \new_[56953]_ ;
  assign \new_[56955]_  = \new_[56954]_  & \new_[56949]_ ;
  assign \new_[56959]_  = ~A266 & ~A265;
  assign \new_[56960]_  = ~A200 & \new_[56959]_ ;
  assign \new_[56963]_  = ~A299 & A298;
  assign \new_[56966]_  = A301 & A300;
  assign \new_[56967]_  = \new_[56966]_  & \new_[56963]_ ;
  assign \new_[56968]_  = \new_[56967]_  & \new_[56960]_ ;
  assign \new_[56972]_  = ~A168 & ~A169;
  assign \new_[56973]_  = ~A170 & \new_[56972]_ ;
  assign \new_[56977]_  = ~A199 & ~A166;
  assign \new_[56978]_  = A167 & \new_[56977]_ ;
  assign \new_[56979]_  = \new_[56978]_  & \new_[56973]_ ;
  assign \new_[56983]_  = ~A266 & ~A265;
  assign \new_[56984]_  = ~A200 & \new_[56983]_ ;
  assign \new_[56987]_  = ~A299 & A298;
  assign \new_[56990]_  = ~A302 & A300;
  assign \new_[56991]_  = \new_[56990]_  & \new_[56987]_ ;
  assign \new_[56992]_  = \new_[56991]_  & \new_[56984]_ ;
  assign \new_[56996]_  = ~A168 & ~A169;
  assign \new_[56997]_  = ~A170 & \new_[56996]_ ;
  assign \new_[57001]_  = ~A199 & ~A166;
  assign \new_[57002]_  = A167 & \new_[57001]_ ;
  assign \new_[57003]_  = \new_[57002]_  & \new_[56997]_ ;
  assign \new_[57007]_  = ~A266 & ~A265;
  assign \new_[57008]_  = ~A200 & \new_[57007]_ ;
  assign \new_[57011]_  = A299 & ~A298;
  assign \new_[57014]_  = A301 & A300;
  assign \new_[57015]_  = \new_[57014]_  & \new_[57011]_ ;
  assign \new_[57016]_  = \new_[57015]_  & \new_[57008]_ ;
  assign \new_[57020]_  = ~A168 & ~A169;
  assign \new_[57021]_  = ~A170 & \new_[57020]_ ;
  assign \new_[57025]_  = ~A199 & ~A166;
  assign \new_[57026]_  = A167 & \new_[57025]_ ;
  assign \new_[57027]_  = \new_[57026]_  & \new_[57021]_ ;
  assign \new_[57031]_  = ~A266 & ~A265;
  assign \new_[57032]_  = ~A200 & \new_[57031]_ ;
  assign \new_[57035]_  = A299 & ~A298;
  assign \new_[57038]_  = ~A302 & A300;
  assign \new_[57039]_  = \new_[57038]_  & \new_[57035]_ ;
  assign \new_[57040]_  = \new_[57039]_  & \new_[57032]_ ;
  assign \new_[57044]_  = ~A168 & ~A169;
  assign \new_[57045]_  = ~A170 & \new_[57044]_ ;
  assign \new_[57049]_  = ~A201 & A166;
  assign \new_[57050]_  = ~A167 & \new_[57049]_ ;
  assign \new_[57051]_  = \new_[57050]_  & \new_[57045]_ ;
  assign \new_[57055]_  = A268 & ~A267;
  assign \new_[57056]_  = A202 & \new_[57055]_ ;
  assign \new_[57059]_  = ~A299 & A298;
  assign \new_[57062]_  = A301 & A300;
  assign \new_[57063]_  = \new_[57062]_  & \new_[57059]_ ;
  assign \new_[57064]_  = \new_[57063]_  & \new_[57056]_ ;
  assign \new_[57068]_  = ~A168 & ~A169;
  assign \new_[57069]_  = ~A170 & \new_[57068]_ ;
  assign \new_[57073]_  = ~A201 & A166;
  assign \new_[57074]_  = ~A167 & \new_[57073]_ ;
  assign \new_[57075]_  = \new_[57074]_  & \new_[57069]_ ;
  assign \new_[57079]_  = A268 & ~A267;
  assign \new_[57080]_  = A202 & \new_[57079]_ ;
  assign \new_[57083]_  = ~A299 & A298;
  assign \new_[57086]_  = ~A302 & A300;
  assign \new_[57087]_  = \new_[57086]_  & \new_[57083]_ ;
  assign \new_[57088]_  = \new_[57087]_  & \new_[57080]_ ;
  assign \new_[57092]_  = ~A168 & ~A169;
  assign \new_[57093]_  = ~A170 & \new_[57092]_ ;
  assign \new_[57097]_  = ~A201 & A166;
  assign \new_[57098]_  = ~A167 & \new_[57097]_ ;
  assign \new_[57099]_  = \new_[57098]_  & \new_[57093]_ ;
  assign \new_[57103]_  = A268 & ~A267;
  assign \new_[57104]_  = A202 & \new_[57103]_ ;
  assign \new_[57107]_  = A299 & ~A298;
  assign \new_[57110]_  = A301 & A300;
  assign \new_[57111]_  = \new_[57110]_  & \new_[57107]_ ;
  assign \new_[57112]_  = \new_[57111]_  & \new_[57104]_ ;
  assign \new_[57116]_  = ~A168 & ~A169;
  assign \new_[57117]_  = ~A170 & \new_[57116]_ ;
  assign \new_[57121]_  = ~A201 & A166;
  assign \new_[57122]_  = ~A167 & \new_[57121]_ ;
  assign \new_[57123]_  = \new_[57122]_  & \new_[57117]_ ;
  assign \new_[57127]_  = A268 & ~A267;
  assign \new_[57128]_  = A202 & \new_[57127]_ ;
  assign \new_[57131]_  = A299 & ~A298;
  assign \new_[57134]_  = ~A302 & A300;
  assign \new_[57135]_  = \new_[57134]_  & \new_[57131]_ ;
  assign \new_[57136]_  = \new_[57135]_  & \new_[57128]_ ;
  assign \new_[57140]_  = ~A168 & ~A169;
  assign \new_[57141]_  = ~A170 & \new_[57140]_ ;
  assign \new_[57145]_  = ~A201 & A166;
  assign \new_[57146]_  = ~A167 & \new_[57145]_ ;
  assign \new_[57147]_  = \new_[57146]_  & \new_[57141]_ ;
  assign \new_[57151]_  = ~A269 & ~A267;
  assign \new_[57152]_  = A202 & \new_[57151]_ ;
  assign \new_[57155]_  = ~A299 & A298;
  assign \new_[57158]_  = A301 & A300;
  assign \new_[57159]_  = \new_[57158]_  & \new_[57155]_ ;
  assign \new_[57160]_  = \new_[57159]_  & \new_[57152]_ ;
  assign \new_[57164]_  = ~A168 & ~A169;
  assign \new_[57165]_  = ~A170 & \new_[57164]_ ;
  assign \new_[57169]_  = ~A201 & A166;
  assign \new_[57170]_  = ~A167 & \new_[57169]_ ;
  assign \new_[57171]_  = \new_[57170]_  & \new_[57165]_ ;
  assign \new_[57175]_  = ~A269 & ~A267;
  assign \new_[57176]_  = A202 & \new_[57175]_ ;
  assign \new_[57179]_  = ~A299 & A298;
  assign \new_[57182]_  = ~A302 & A300;
  assign \new_[57183]_  = \new_[57182]_  & \new_[57179]_ ;
  assign \new_[57184]_  = \new_[57183]_  & \new_[57176]_ ;
  assign \new_[57188]_  = ~A168 & ~A169;
  assign \new_[57189]_  = ~A170 & \new_[57188]_ ;
  assign \new_[57193]_  = ~A201 & A166;
  assign \new_[57194]_  = ~A167 & \new_[57193]_ ;
  assign \new_[57195]_  = \new_[57194]_  & \new_[57189]_ ;
  assign \new_[57199]_  = ~A269 & ~A267;
  assign \new_[57200]_  = A202 & \new_[57199]_ ;
  assign \new_[57203]_  = A299 & ~A298;
  assign \new_[57206]_  = A301 & A300;
  assign \new_[57207]_  = \new_[57206]_  & \new_[57203]_ ;
  assign \new_[57208]_  = \new_[57207]_  & \new_[57200]_ ;
  assign \new_[57212]_  = ~A168 & ~A169;
  assign \new_[57213]_  = ~A170 & \new_[57212]_ ;
  assign \new_[57217]_  = ~A201 & A166;
  assign \new_[57218]_  = ~A167 & \new_[57217]_ ;
  assign \new_[57219]_  = \new_[57218]_  & \new_[57213]_ ;
  assign \new_[57223]_  = ~A269 & ~A267;
  assign \new_[57224]_  = A202 & \new_[57223]_ ;
  assign \new_[57227]_  = A299 & ~A298;
  assign \new_[57230]_  = ~A302 & A300;
  assign \new_[57231]_  = \new_[57230]_  & \new_[57227]_ ;
  assign \new_[57232]_  = \new_[57231]_  & \new_[57224]_ ;
  assign \new_[57236]_  = ~A168 & ~A169;
  assign \new_[57237]_  = ~A170 & \new_[57236]_ ;
  assign \new_[57241]_  = ~A201 & A166;
  assign \new_[57242]_  = ~A167 & \new_[57241]_ ;
  assign \new_[57243]_  = \new_[57242]_  & \new_[57237]_ ;
  assign \new_[57247]_  = A266 & A265;
  assign \new_[57248]_  = A202 & \new_[57247]_ ;
  assign \new_[57251]_  = ~A299 & A298;
  assign \new_[57254]_  = A301 & A300;
  assign \new_[57255]_  = \new_[57254]_  & \new_[57251]_ ;
  assign \new_[57256]_  = \new_[57255]_  & \new_[57248]_ ;
  assign \new_[57260]_  = ~A168 & ~A169;
  assign \new_[57261]_  = ~A170 & \new_[57260]_ ;
  assign \new_[57265]_  = ~A201 & A166;
  assign \new_[57266]_  = ~A167 & \new_[57265]_ ;
  assign \new_[57267]_  = \new_[57266]_  & \new_[57261]_ ;
  assign \new_[57271]_  = A266 & A265;
  assign \new_[57272]_  = A202 & \new_[57271]_ ;
  assign \new_[57275]_  = ~A299 & A298;
  assign \new_[57278]_  = ~A302 & A300;
  assign \new_[57279]_  = \new_[57278]_  & \new_[57275]_ ;
  assign \new_[57280]_  = \new_[57279]_  & \new_[57272]_ ;
  assign \new_[57284]_  = ~A168 & ~A169;
  assign \new_[57285]_  = ~A170 & \new_[57284]_ ;
  assign \new_[57289]_  = ~A201 & A166;
  assign \new_[57290]_  = ~A167 & \new_[57289]_ ;
  assign \new_[57291]_  = \new_[57290]_  & \new_[57285]_ ;
  assign \new_[57295]_  = A266 & A265;
  assign \new_[57296]_  = A202 & \new_[57295]_ ;
  assign \new_[57299]_  = A299 & ~A298;
  assign \new_[57302]_  = A301 & A300;
  assign \new_[57303]_  = \new_[57302]_  & \new_[57299]_ ;
  assign \new_[57304]_  = \new_[57303]_  & \new_[57296]_ ;
  assign \new_[57308]_  = ~A168 & ~A169;
  assign \new_[57309]_  = ~A170 & \new_[57308]_ ;
  assign \new_[57313]_  = ~A201 & A166;
  assign \new_[57314]_  = ~A167 & \new_[57313]_ ;
  assign \new_[57315]_  = \new_[57314]_  & \new_[57309]_ ;
  assign \new_[57319]_  = A266 & A265;
  assign \new_[57320]_  = A202 & \new_[57319]_ ;
  assign \new_[57323]_  = A299 & ~A298;
  assign \new_[57326]_  = ~A302 & A300;
  assign \new_[57327]_  = \new_[57326]_  & \new_[57323]_ ;
  assign \new_[57328]_  = \new_[57327]_  & \new_[57320]_ ;
  assign \new_[57332]_  = ~A168 & ~A169;
  assign \new_[57333]_  = ~A170 & \new_[57332]_ ;
  assign \new_[57337]_  = ~A201 & A166;
  assign \new_[57338]_  = ~A167 & \new_[57337]_ ;
  assign \new_[57339]_  = \new_[57338]_  & \new_[57333]_ ;
  assign \new_[57343]_  = A266 & ~A265;
  assign \new_[57344]_  = A202 & \new_[57343]_ ;
  assign \new_[57347]_  = A268 & A267;
  assign \new_[57350]_  = A301 & ~A300;
  assign \new_[57351]_  = \new_[57350]_  & \new_[57347]_ ;
  assign \new_[57352]_  = \new_[57351]_  & \new_[57344]_ ;
  assign \new_[57356]_  = ~A168 & ~A169;
  assign \new_[57357]_  = ~A170 & \new_[57356]_ ;
  assign \new_[57361]_  = ~A201 & A166;
  assign \new_[57362]_  = ~A167 & \new_[57361]_ ;
  assign \new_[57363]_  = \new_[57362]_  & \new_[57357]_ ;
  assign \new_[57367]_  = A266 & ~A265;
  assign \new_[57368]_  = A202 & \new_[57367]_ ;
  assign \new_[57371]_  = A268 & A267;
  assign \new_[57374]_  = ~A302 & ~A300;
  assign \new_[57375]_  = \new_[57374]_  & \new_[57371]_ ;
  assign \new_[57376]_  = \new_[57375]_  & \new_[57368]_ ;
  assign \new_[57380]_  = ~A168 & ~A169;
  assign \new_[57381]_  = ~A170 & \new_[57380]_ ;
  assign \new_[57385]_  = ~A201 & A166;
  assign \new_[57386]_  = ~A167 & \new_[57385]_ ;
  assign \new_[57387]_  = \new_[57386]_  & \new_[57381]_ ;
  assign \new_[57391]_  = A266 & ~A265;
  assign \new_[57392]_  = A202 & \new_[57391]_ ;
  assign \new_[57395]_  = A268 & A267;
  assign \new_[57398]_  = A299 & A298;
  assign \new_[57399]_  = \new_[57398]_  & \new_[57395]_ ;
  assign \new_[57400]_  = \new_[57399]_  & \new_[57392]_ ;
  assign \new_[57404]_  = ~A168 & ~A169;
  assign \new_[57405]_  = ~A170 & \new_[57404]_ ;
  assign \new_[57409]_  = ~A201 & A166;
  assign \new_[57410]_  = ~A167 & \new_[57409]_ ;
  assign \new_[57411]_  = \new_[57410]_  & \new_[57405]_ ;
  assign \new_[57415]_  = A266 & ~A265;
  assign \new_[57416]_  = A202 & \new_[57415]_ ;
  assign \new_[57419]_  = A268 & A267;
  assign \new_[57422]_  = ~A299 & ~A298;
  assign \new_[57423]_  = \new_[57422]_  & \new_[57419]_ ;
  assign \new_[57424]_  = \new_[57423]_  & \new_[57416]_ ;
  assign \new_[57428]_  = ~A168 & ~A169;
  assign \new_[57429]_  = ~A170 & \new_[57428]_ ;
  assign \new_[57433]_  = ~A201 & A166;
  assign \new_[57434]_  = ~A167 & \new_[57433]_ ;
  assign \new_[57435]_  = \new_[57434]_  & \new_[57429]_ ;
  assign \new_[57439]_  = A266 & ~A265;
  assign \new_[57440]_  = A202 & \new_[57439]_ ;
  assign \new_[57443]_  = ~A269 & A267;
  assign \new_[57446]_  = A301 & ~A300;
  assign \new_[57447]_  = \new_[57446]_  & \new_[57443]_ ;
  assign \new_[57448]_  = \new_[57447]_  & \new_[57440]_ ;
  assign \new_[57452]_  = ~A168 & ~A169;
  assign \new_[57453]_  = ~A170 & \new_[57452]_ ;
  assign \new_[57457]_  = ~A201 & A166;
  assign \new_[57458]_  = ~A167 & \new_[57457]_ ;
  assign \new_[57459]_  = \new_[57458]_  & \new_[57453]_ ;
  assign \new_[57463]_  = A266 & ~A265;
  assign \new_[57464]_  = A202 & \new_[57463]_ ;
  assign \new_[57467]_  = ~A269 & A267;
  assign \new_[57470]_  = ~A302 & ~A300;
  assign \new_[57471]_  = \new_[57470]_  & \new_[57467]_ ;
  assign \new_[57472]_  = \new_[57471]_  & \new_[57464]_ ;
  assign \new_[57476]_  = ~A168 & ~A169;
  assign \new_[57477]_  = ~A170 & \new_[57476]_ ;
  assign \new_[57481]_  = ~A201 & A166;
  assign \new_[57482]_  = ~A167 & \new_[57481]_ ;
  assign \new_[57483]_  = \new_[57482]_  & \new_[57477]_ ;
  assign \new_[57487]_  = A266 & ~A265;
  assign \new_[57488]_  = A202 & \new_[57487]_ ;
  assign \new_[57491]_  = ~A269 & A267;
  assign \new_[57494]_  = A299 & A298;
  assign \new_[57495]_  = \new_[57494]_  & \new_[57491]_ ;
  assign \new_[57496]_  = \new_[57495]_  & \new_[57488]_ ;
  assign \new_[57500]_  = ~A168 & ~A169;
  assign \new_[57501]_  = ~A170 & \new_[57500]_ ;
  assign \new_[57505]_  = ~A201 & A166;
  assign \new_[57506]_  = ~A167 & \new_[57505]_ ;
  assign \new_[57507]_  = \new_[57506]_  & \new_[57501]_ ;
  assign \new_[57511]_  = A266 & ~A265;
  assign \new_[57512]_  = A202 & \new_[57511]_ ;
  assign \new_[57515]_  = ~A269 & A267;
  assign \new_[57518]_  = ~A299 & ~A298;
  assign \new_[57519]_  = \new_[57518]_  & \new_[57515]_ ;
  assign \new_[57520]_  = \new_[57519]_  & \new_[57512]_ ;
  assign \new_[57524]_  = ~A168 & ~A169;
  assign \new_[57525]_  = ~A170 & \new_[57524]_ ;
  assign \new_[57529]_  = ~A201 & A166;
  assign \new_[57530]_  = ~A167 & \new_[57529]_ ;
  assign \new_[57531]_  = \new_[57530]_  & \new_[57525]_ ;
  assign \new_[57535]_  = ~A266 & A265;
  assign \new_[57536]_  = A202 & \new_[57535]_ ;
  assign \new_[57539]_  = A268 & A267;
  assign \new_[57542]_  = A301 & ~A300;
  assign \new_[57543]_  = \new_[57542]_  & \new_[57539]_ ;
  assign \new_[57544]_  = \new_[57543]_  & \new_[57536]_ ;
  assign \new_[57548]_  = ~A168 & ~A169;
  assign \new_[57549]_  = ~A170 & \new_[57548]_ ;
  assign \new_[57553]_  = ~A201 & A166;
  assign \new_[57554]_  = ~A167 & \new_[57553]_ ;
  assign \new_[57555]_  = \new_[57554]_  & \new_[57549]_ ;
  assign \new_[57559]_  = ~A266 & A265;
  assign \new_[57560]_  = A202 & \new_[57559]_ ;
  assign \new_[57563]_  = A268 & A267;
  assign \new_[57566]_  = ~A302 & ~A300;
  assign \new_[57567]_  = \new_[57566]_  & \new_[57563]_ ;
  assign \new_[57568]_  = \new_[57567]_  & \new_[57560]_ ;
  assign \new_[57572]_  = ~A168 & ~A169;
  assign \new_[57573]_  = ~A170 & \new_[57572]_ ;
  assign \new_[57577]_  = ~A201 & A166;
  assign \new_[57578]_  = ~A167 & \new_[57577]_ ;
  assign \new_[57579]_  = \new_[57578]_  & \new_[57573]_ ;
  assign \new_[57583]_  = ~A266 & A265;
  assign \new_[57584]_  = A202 & \new_[57583]_ ;
  assign \new_[57587]_  = A268 & A267;
  assign \new_[57590]_  = A299 & A298;
  assign \new_[57591]_  = \new_[57590]_  & \new_[57587]_ ;
  assign \new_[57592]_  = \new_[57591]_  & \new_[57584]_ ;
  assign \new_[57596]_  = ~A168 & ~A169;
  assign \new_[57597]_  = ~A170 & \new_[57596]_ ;
  assign \new_[57601]_  = ~A201 & A166;
  assign \new_[57602]_  = ~A167 & \new_[57601]_ ;
  assign \new_[57603]_  = \new_[57602]_  & \new_[57597]_ ;
  assign \new_[57607]_  = ~A266 & A265;
  assign \new_[57608]_  = A202 & \new_[57607]_ ;
  assign \new_[57611]_  = A268 & A267;
  assign \new_[57614]_  = ~A299 & ~A298;
  assign \new_[57615]_  = \new_[57614]_  & \new_[57611]_ ;
  assign \new_[57616]_  = \new_[57615]_  & \new_[57608]_ ;
  assign \new_[57620]_  = ~A168 & ~A169;
  assign \new_[57621]_  = ~A170 & \new_[57620]_ ;
  assign \new_[57625]_  = ~A201 & A166;
  assign \new_[57626]_  = ~A167 & \new_[57625]_ ;
  assign \new_[57627]_  = \new_[57626]_  & \new_[57621]_ ;
  assign \new_[57631]_  = ~A266 & A265;
  assign \new_[57632]_  = A202 & \new_[57631]_ ;
  assign \new_[57635]_  = ~A269 & A267;
  assign \new_[57638]_  = A301 & ~A300;
  assign \new_[57639]_  = \new_[57638]_  & \new_[57635]_ ;
  assign \new_[57640]_  = \new_[57639]_  & \new_[57632]_ ;
  assign \new_[57644]_  = ~A168 & ~A169;
  assign \new_[57645]_  = ~A170 & \new_[57644]_ ;
  assign \new_[57649]_  = ~A201 & A166;
  assign \new_[57650]_  = ~A167 & \new_[57649]_ ;
  assign \new_[57651]_  = \new_[57650]_  & \new_[57645]_ ;
  assign \new_[57655]_  = ~A266 & A265;
  assign \new_[57656]_  = A202 & \new_[57655]_ ;
  assign \new_[57659]_  = ~A269 & A267;
  assign \new_[57662]_  = ~A302 & ~A300;
  assign \new_[57663]_  = \new_[57662]_  & \new_[57659]_ ;
  assign \new_[57664]_  = \new_[57663]_  & \new_[57656]_ ;
  assign \new_[57668]_  = ~A168 & ~A169;
  assign \new_[57669]_  = ~A170 & \new_[57668]_ ;
  assign \new_[57673]_  = ~A201 & A166;
  assign \new_[57674]_  = ~A167 & \new_[57673]_ ;
  assign \new_[57675]_  = \new_[57674]_  & \new_[57669]_ ;
  assign \new_[57679]_  = ~A266 & A265;
  assign \new_[57680]_  = A202 & \new_[57679]_ ;
  assign \new_[57683]_  = ~A269 & A267;
  assign \new_[57686]_  = A299 & A298;
  assign \new_[57687]_  = \new_[57686]_  & \new_[57683]_ ;
  assign \new_[57688]_  = \new_[57687]_  & \new_[57680]_ ;
  assign \new_[57692]_  = ~A168 & ~A169;
  assign \new_[57693]_  = ~A170 & \new_[57692]_ ;
  assign \new_[57697]_  = ~A201 & A166;
  assign \new_[57698]_  = ~A167 & \new_[57697]_ ;
  assign \new_[57699]_  = \new_[57698]_  & \new_[57693]_ ;
  assign \new_[57703]_  = ~A266 & A265;
  assign \new_[57704]_  = A202 & \new_[57703]_ ;
  assign \new_[57707]_  = ~A269 & A267;
  assign \new_[57710]_  = ~A299 & ~A298;
  assign \new_[57711]_  = \new_[57710]_  & \new_[57707]_ ;
  assign \new_[57712]_  = \new_[57711]_  & \new_[57704]_ ;
  assign \new_[57716]_  = ~A168 & ~A169;
  assign \new_[57717]_  = ~A170 & \new_[57716]_ ;
  assign \new_[57721]_  = ~A201 & A166;
  assign \new_[57722]_  = ~A167 & \new_[57721]_ ;
  assign \new_[57723]_  = \new_[57722]_  & \new_[57717]_ ;
  assign \new_[57727]_  = ~A266 & ~A265;
  assign \new_[57728]_  = A202 & \new_[57727]_ ;
  assign \new_[57731]_  = ~A299 & A298;
  assign \new_[57734]_  = A301 & A300;
  assign \new_[57735]_  = \new_[57734]_  & \new_[57731]_ ;
  assign \new_[57736]_  = \new_[57735]_  & \new_[57728]_ ;
  assign \new_[57740]_  = ~A168 & ~A169;
  assign \new_[57741]_  = ~A170 & \new_[57740]_ ;
  assign \new_[57745]_  = ~A201 & A166;
  assign \new_[57746]_  = ~A167 & \new_[57745]_ ;
  assign \new_[57747]_  = \new_[57746]_  & \new_[57741]_ ;
  assign \new_[57751]_  = ~A266 & ~A265;
  assign \new_[57752]_  = A202 & \new_[57751]_ ;
  assign \new_[57755]_  = ~A299 & A298;
  assign \new_[57758]_  = ~A302 & A300;
  assign \new_[57759]_  = \new_[57758]_  & \new_[57755]_ ;
  assign \new_[57760]_  = \new_[57759]_  & \new_[57752]_ ;
  assign \new_[57764]_  = ~A168 & ~A169;
  assign \new_[57765]_  = ~A170 & \new_[57764]_ ;
  assign \new_[57769]_  = ~A201 & A166;
  assign \new_[57770]_  = ~A167 & \new_[57769]_ ;
  assign \new_[57771]_  = \new_[57770]_  & \new_[57765]_ ;
  assign \new_[57775]_  = ~A266 & ~A265;
  assign \new_[57776]_  = A202 & \new_[57775]_ ;
  assign \new_[57779]_  = A299 & ~A298;
  assign \new_[57782]_  = A301 & A300;
  assign \new_[57783]_  = \new_[57782]_  & \new_[57779]_ ;
  assign \new_[57784]_  = \new_[57783]_  & \new_[57776]_ ;
  assign \new_[57788]_  = ~A168 & ~A169;
  assign \new_[57789]_  = ~A170 & \new_[57788]_ ;
  assign \new_[57793]_  = ~A201 & A166;
  assign \new_[57794]_  = ~A167 & \new_[57793]_ ;
  assign \new_[57795]_  = \new_[57794]_  & \new_[57789]_ ;
  assign \new_[57799]_  = ~A266 & ~A265;
  assign \new_[57800]_  = A202 & \new_[57799]_ ;
  assign \new_[57803]_  = A299 & ~A298;
  assign \new_[57806]_  = ~A302 & A300;
  assign \new_[57807]_  = \new_[57806]_  & \new_[57803]_ ;
  assign \new_[57808]_  = \new_[57807]_  & \new_[57800]_ ;
  assign \new_[57812]_  = ~A168 & ~A169;
  assign \new_[57813]_  = ~A170 & \new_[57812]_ ;
  assign \new_[57817]_  = ~A201 & A166;
  assign \new_[57818]_  = ~A167 & \new_[57817]_ ;
  assign \new_[57819]_  = \new_[57818]_  & \new_[57813]_ ;
  assign \new_[57823]_  = A268 & ~A267;
  assign \new_[57824]_  = ~A203 & \new_[57823]_ ;
  assign \new_[57827]_  = ~A299 & A298;
  assign \new_[57830]_  = A301 & A300;
  assign \new_[57831]_  = \new_[57830]_  & \new_[57827]_ ;
  assign \new_[57832]_  = \new_[57831]_  & \new_[57824]_ ;
  assign \new_[57836]_  = ~A168 & ~A169;
  assign \new_[57837]_  = ~A170 & \new_[57836]_ ;
  assign \new_[57841]_  = ~A201 & A166;
  assign \new_[57842]_  = ~A167 & \new_[57841]_ ;
  assign \new_[57843]_  = \new_[57842]_  & \new_[57837]_ ;
  assign \new_[57847]_  = A268 & ~A267;
  assign \new_[57848]_  = ~A203 & \new_[57847]_ ;
  assign \new_[57851]_  = ~A299 & A298;
  assign \new_[57854]_  = ~A302 & A300;
  assign \new_[57855]_  = \new_[57854]_  & \new_[57851]_ ;
  assign \new_[57856]_  = \new_[57855]_  & \new_[57848]_ ;
  assign \new_[57860]_  = ~A168 & ~A169;
  assign \new_[57861]_  = ~A170 & \new_[57860]_ ;
  assign \new_[57865]_  = ~A201 & A166;
  assign \new_[57866]_  = ~A167 & \new_[57865]_ ;
  assign \new_[57867]_  = \new_[57866]_  & \new_[57861]_ ;
  assign \new_[57871]_  = A268 & ~A267;
  assign \new_[57872]_  = ~A203 & \new_[57871]_ ;
  assign \new_[57875]_  = A299 & ~A298;
  assign \new_[57878]_  = A301 & A300;
  assign \new_[57879]_  = \new_[57878]_  & \new_[57875]_ ;
  assign \new_[57880]_  = \new_[57879]_  & \new_[57872]_ ;
  assign \new_[57884]_  = ~A168 & ~A169;
  assign \new_[57885]_  = ~A170 & \new_[57884]_ ;
  assign \new_[57889]_  = ~A201 & A166;
  assign \new_[57890]_  = ~A167 & \new_[57889]_ ;
  assign \new_[57891]_  = \new_[57890]_  & \new_[57885]_ ;
  assign \new_[57895]_  = A268 & ~A267;
  assign \new_[57896]_  = ~A203 & \new_[57895]_ ;
  assign \new_[57899]_  = A299 & ~A298;
  assign \new_[57902]_  = ~A302 & A300;
  assign \new_[57903]_  = \new_[57902]_  & \new_[57899]_ ;
  assign \new_[57904]_  = \new_[57903]_  & \new_[57896]_ ;
  assign \new_[57908]_  = ~A168 & ~A169;
  assign \new_[57909]_  = ~A170 & \new_[57908]_ ;
  assign \new_[57913]_  = ~A201 & A166;
  assign \new_[57914]_  = ~A167 & \new_[57913]_ ;
  assign \new_[57915]_  = \new_[57914]_  & \new_[57909]_ ;
  assign \new_[57919]_  = ~A269 & ~A267;
  assign \new_[57920]_  = ~A203 & \new_[57919]_ ;
  assign \new_[57923]_  = ~A299 & A298;
  assign \new_[57926]_  = A301 & A300;
  assign \new_[57927]_  = \new_[57926]_  & \new_[57923]_ ;
  assign \new_[57928]_  = \new_[57927]_  & \new_[57920]_ ;
  assign \new_[57932]_  = ~A168 & ~A169;
  assign \new_[57933]_  = ~A170 & \new_[57932]_ ;
  assign \new_[57937]_  = ~A201 & A166;
  assign \new_[57938]_  = ~A167 & \new_[57937]_ ;
  assign \new_[57939]_  = \new_[57938]_  & \new_[57933]_ ;
  assign \new_[57943]_  = ~A269 & ~A267;
  assign \new_[57944]_  = ~A203 & \new_[57943]_ ;
  assign \new_[57947]_  = ~A299 & A298;
  assign \new_[57950]_  = ~A302 & A300;
  assign \new_[57951]_  = \new_[57950]_  & \new_[57947]_ ;
  assign \new_[57952]_  = \new_[57951]_  & \new_[57944]_ ;
  assign \new_[57956]_  = ~A168 & ~A169;
  assign \new_[57957]_  = ~A170 & \new_[57956]_ ;
  assign \new_[57961]_  = ~A201 & A166;
  assign \new_[57962]_  = ~A167 & \new_[57961]_ ;
  assign \new_[57963]_  = \new_[57962]_  & \new_[57957]_ ;
  assign \new_[57967]_  = ~A269 & ~A267;
  assign \new_[57968]_  = ~A203 & \new_[57967]_ ;
  assign \new_[57971]_  = A299 & ~A298;
  assign \new_[57974]_  = A301 & A300;
  assign \new_[57975]_  = \new_[57974]_  & \new_[57971]_ ;
  assign \new_[57976]_  = \new_[57975]_  & \new_[57968]_ ;
  assign \new_[57980]_  = ~A168 & ~A169;
  assign \new_[57981]_  = ~A170 & \new_[57980]_ ;
  assign \new_[57985]_  = ~A201 & A166;
  assign \new_[57986]_  = ~A167 & \new_[57985]_ ;
  assign \new_[57987]_  = \new_[57986]_  & \new_[57981]_ ;
  assign \new_[57991]_  = ~A269 & ~A267;
  assign \new_[57992]_  = ~A203 & \new_[57991]_ ;
  assign \new_[57995]_  = A299 & ~A298;
  assign \new_[57998]_  = ~A302 & A300;
  assign \new_[57999]_  = \new_[57998]_  & \new_[57995]_ ;
  assign \new_[58000]_  = \new_[57999]_  & \new_[57992]_ ;
  assign \new_[58004]_  = ~A168 & ~A169;
  assign \new_[58005]_  = ~A170 & \new_[58004]_ ;
  assign \new_[58009]_  = ~A201 & A166;
  assign \new_[58010]_  = ~A167 & \new_[58009]_ ;
  assign \new_[58011]_  = \new_[58010]_  & \new_[58005]_ ;
  assign \new_[58015]_  = A266 & A265;
  assign \new_[58016]_  = ~A203 & \new_[58015]_ ;
  assign \new_[58019]_  = ~A299 & A298;
  assign \new_[58022]_  = A301 & A300;
  assign \new_[58023]_  = \new_[58022]_  & \new_[58019]_ ;
  assign \new_[58024]_  = \new_[58023]_  & \new_[58016]_ ;
  assign \new_[58028]_  = ~A168 & ~A169;
  assign \new_[58029]_  = ~A170 & \new_[58028]_ ;
  assign \new_[58033]_  = ~A201 & A166;
  assign \new_[58034]_  = ~A167 & \new_[58033]_ ;
  assign \new_[58035]_  = \new_[58034]_  & \new_[58029]_ ;
  assign \new_[58039]_  = A266 & A265;
  assign \new_[58040]_  = ~A203 & \new_[58039]_ ;
  assign \new_[58043]_  = ~A299 & A298;
  assign \new_[58046]_  = ~A302 & A300;
  assign \new_[58047]_  = \new_[58046]_  & \new_[58043]_ ;
  assign \new_[58048]_  = \new_[58047]_  & \new_[58040]_ ;
  assign \new_[58052]_  = ~A168 & ~A169;
  assign \new_[58053]_  = ~A170 & \new_[58052]_ ;
  assign \new_[58057]_  = ~A201 & A166;
  assign \new_[58058]_  = ~A167 & \new_[58057]_ ;
  assign \new_[58059]_  = \new_[58058]_  & \new_[58053]_ ;
  assign \new_[58063]_  = A266 & A265;
  assign \new_[58064]_  = ~A203 & \new_[58063]_ ;
  assign \new_[58067]_  = A299 & ~A298;
  assign \new_[58070]_  = A301 & A300;
  assign \new_[58071]_  = \new_[58070]_  & \new_[58067]_ ;
  assign \new_[58072]_  = \new_[58071]_  & \new_[58064]_ ;
  assign \new_[58076]_  = ~A168 & ~A169;
  assign \new_[58077]_  = ~A170 & \new_[58076]_ ;
  assign \new_[58081]_  = ~A201 & A166;
  assign \new_[58082]_  = ~A167 & \new_[58081]_ ;
  assign \new_[58083]_  = \new_[58082]_  & \new_[58077]_ ;
  assign \new_[58087]_  = A266 & A265;
  assign \new_[58088]_  = ~A203 & \new_[58087]_ ;
  assign \new_[58091]_  = A299 & ~A298;
  assign \new_[58094]_  = ~A302 & A300;
  assign \new_[58095]_  = \new_[58094]_  & \new_[58091]_ ;
  assign \new_[58096]_  = \new_[58095]_  & \new_[58088]_ ;
  assign \new_[58100]_  = ~A168 & ~A169;
  assign \new_[58101]_  = ~A170 & \new_[58100]_ ;
  assign \new_[58105]_  = ~A201 & A166;
  assign \new_[58106]_  = ~A167 & \new_[58105]_ ;
  assign \new_[58107]_  = \new_[58106]_  & \new_[58101]_ ;
  assign \new_[58111]_  = A266 & ~A265;
  assign \new_[58112]_  = ~A203 & \new_[58111]_ ;
  assign \new_[58115]_  = A268 & A267;
  assign \new_[58118]_  = A301 & ~A300;
  assign \new_[58119]_  = \new_[58118]_  & \new_[58115]_ ;
  assign \new_[58120]_  = \new_[58119]_  & \new_[58112]_ ;
  assign \new_[58124]_  = ~A168 & ~A169;
  assign \new_[58125]_  = ~A170 & \new_[58124]_ ;
  assign \new_[58129]_  = ~A201 & A166;
  assign \new_[58130]_  = ~A167 & \new_[58129]_ ;
  assign \new_[58131]_  = \new_[58130]_  & \new_[58125]_ ;
  assign \new_[58135]_  = A266 & ~A265;
  assign \new_[58136]_  = ~A203 & \new_[58135]_ ;
  assign \new_[58139]_  = A268 & A267;
  assign \new_[58142]_  = ~A302 & ~A300;
  assign \new_[58143]_  = \new_[58142]_  & \new_[58139]_ ;
  assign \new_[58144]_  = \new_[58143]_  & \new_[58136]_ ;
  assign \new_[58148]_  = ~A168 & ~A169;
  assign \new_[58149]_  = ~A170 & \new_[58148]_ ;
  assign \new_[58153]_  = ~A201 & A166;
  assign \new_[58154]_  = ~A167 & \new_[58153]_ ;
  assign \new_[58155]_  = \new_[58154]_  & \new_[58149]_ ;
  assign \new_[58159]_  = A266 & ~A265;
  assign \new_[58160]_  = ~A203 & \new_[58159]_ ;
  assign \new_[58163]_  = A268 & A267;
  assign \new_[58166]_  = A299 & A298;
  assign \new_[58167]_  = \new_[58166]_  & \new_[58163]_ ;
  assign \new_[58168]_  = \new_[58167]_  & \new_[58160]_ ;
  assign \new_[58172]_  = ~A168 & ~A169;
  assign \new_[58173]_  = ~A170 & \new_[58172]_ ;
  assign \new_[58177]_  = ~A201 & A166;
  assign \new_[58178]_  = ~A167 & \new_[58177]_ ;
  assign \new_[58179]_  = \new_[58178]_  & \new_[58173]_ ;
  assign \new_[58183]_  = A266 & ~A265;
  assign \new_[58184]_  = ~A203 & \new_[58183]_ ;
  assign \new_[58187]_  = A268 & A267;
  assign \new_[58190]_  = ~A299 & ~A298;
  assign \new_[58191]_  = \new_[58190]_  & \new_[58187]_ ;
  assign \new_[58192]_  = \new_[58191]_  & \new_[58184]_ ;
  assign \new_[58196]_  = ~A168 & ~A169;
  assign \new_[58197]_  = ~A170 & \new_[58196]_ ;
  assign \new_[58201]_  = ~A201 & A166;
  assign \new_[58202]_  = ~A167 & \new_[58201]_ ;
  assign \new_[58203]_  = \new_[58202]_  & \new_[58197]_ ;
  assign \new_[58207]_  = A266 & ~A265;
  assign \new_[58208]_  = ~A203 & \new_[58207]_ ;
  assign \new_[58211]_  = ~A269 & A267;
  assign \new_[58214]_  = A301 & ~A300;
  assign \new_[58215]_  = \new_[58214]_  & \new_[58211]_ ;
  assign \new_[58216]_  = \new_[58215]_  & \new_[58208]_ ;
  assign \new_[58220]_  = ~A168 & ~A169;
  assign \new_[58221]_  = ~A170 & \new_[58220]_ ;
  assign \new_[58225]_  = ~A201 & A166;
  assign \new_[58226]_  = ~A167 & \new_[58225]_ ;
  assign \new_[58227]_  = \new_[58226]_  & \new_[58221]_ ;
  assign \new_[58231]_  = A266 & ~A265;
  assign \new_[58232]_  = ~A203 & \new_[58231]_ ;
  assign \new_[58235]_  = ~A269 & A267;
  assign \new_[58238]_  = ~A302 & ~A300;
  assign \new_[58239]_  = \new_[58238]_  & \new_[58235]_ ;
  assign \new_[58240]_  = \new_[58239]_  & \new_[58232]_ ;
  assign \new_[58244]_  = ~A168 & ~A169;
  assign \new_[58245]_  = ~A170 & \new_[58244]_ ;
  assign \new_[58249]_  = ~A201 & A166;
  assign \new_[58250]_  = ~A167 & \new_[58249]_ ;
  assign \new_[58251]_  = \new_[58250]_  & \new_[58245]_ ;
  assign \new_[58255]_  = A266 & ~A265;
  assign \new_[58256]_  = ~A203 & \new_[58255]_ ;
  assign \new_[58259]_  = ~A269 & A267;
  assign \new_[58262]_  = A299 & A298;
  assign \new_[58263]_  = \new_[58262]_  & \new_[58259]_ ;
  assign \new_[58264]_  = \new_[58263]_  & \new_[58256]_ ;
  assign \new_[58268]_  = ~A168 & ~A169;
  assign \new_[58269]_  = ~A170 & \new_[58268]_ ;
  assign \new_[58273]_  = ~A201 & A166;
  assign \new_[58274]_  = ~A167 & \new_[58273]_ ;
  assign \new_[58275]_  = \new_[58274]_  & \new_[58269]_ ;
  assign \new_[58279]_  = A266 & ~A265;
  assign \new_[58280]_  = ~A203 & \new_[58279]_ ;
  assign \new_[58283]_  = ~A269 & A267;
  assign \new_[58286]_  = ~A299 & ~A298;
  assign \new_[58287]_  = \new_[58286]_  & \new_[58283]_ ;
  assign \new_[58288]_  = \new_[58287]_  & \new_[58280]_ ;
  assign \new_[58292]_  = ~A168 & ~A169;
  assign \new_[58293]_  = ~A170 & \new_[58292]_ ;
  assign \new_[58297]_  = ~A201 & A166;
  assign \new_[58298]_  = ~A167 & \new_[58297]_ ;
  assign \new_[58299]_  = \new_[58298]_  & \new_[58293]_ ;
  assign \new_[58303]_  = ~A266 & A265;
  assign \new_[58304]_  = ~A203 & \new_[58303]_ ;
  assign \new_[58307]_  = A268 & A267;
  assign \new_[58310]_  = A301 & ~A300;
  assign \new_[58311]_  = \new_[58310]_  & \new_[58307]_ ;
  assign \new_[58312]_  = \new_[58311]_  & \new_[58304]_ ;
  assign \new_[58316]_  = ~A168 & ~A169;
  assign \new_[58317]_  = ~A170 & \new_[58316]_ ;
  assign \new_[58321]_  = ~A201 & A166;
  assign \new_[58322]_  = ~A167 & \new_[58321]_ ;
  assign \new_[58323]_  = \new_[58322]_  & \new_[58317]_ ;
  assign \new_[58327]_  = ~A266 & A265;
  assign \new_[58328]_  = ~A203 & \new_[58327]_ ;
  assign \new_[58331]_  = A268 & A267;
  assign \new_[58334]_  = ~A302 & ~A300;
  assign \new_[58335]_  = \new_[58334]_  & \new_[58331]_ ;
  assign \new_[58336]_  = \new_[58335]_  & \new_[58328]_ ;
  assign \new_[58340]_  = ~A168 & ~A169;
  assign \new_[58341]_  = ~A170 & \new_[58340]_ ;
  assign \new_[58345]_  = ~A201 & A166;
  assign \new_[58346]_  = ~A167 & \new_[58345]_ ;
  assign \new_[58347]_  = \new_[58346]_  & \new_[58341]_ ;
  assign \new_[58351]_  = ~A266 & A265;
  assign \new_[58352]_  = ~A203 & \new_[58351]_ ;
  assign \new_[58355]_  = A268 & A267;
  assign \new_[58358]_  = A299 & A298;
  assign \new_[58359]_  = \new_[58358]_  & \new_[58355]_ ;
  assign \new_[58360]_  = \new_[58359]_  & \new_[58352]_ ;
  assign \new_[58364]_  = ~A168 & ~A169;
  assign \new_[58365]_  = ~A170 & \new_[58364]_ ;
  assign \new_[58369]_  = ~A201 & A166;
  assign \new_[58370]_  = ~A167 & \new_[58369]_ ;
  assign \new_[58371]_  = \new_[58370]_  & \new_[58365]_ ;
  assign \new_[58375]_  = ~A266 & A265;
  assign \new_[58376]_  = ~A203 & \new_[58375]_ ;
  assign \new_[58379]_  = A268 & A267;
  assign \new_[58382]_  = ~A299 & ~A298;
  assign \new_[58383]_  = \new_[58382]_  & \new_[58379]_ ;
  assign \new_[58384]_  = \new_[58383]_  & \new_[58376]_ ;
  assign \new_[58388]_  = ~A168 & ~A169;
  assign \new_[58389]_  = ~A170 & \new_[58388]_ ;
  assign \new_[58393]_  = ~A201 & A166;
  assign \new_[58394]_  = ~A167 & \new_[58393]_ ;
  assign \new_[58395]_  = \new_[58394]_  & \new_[58389]_ ;
  assign \new_[58399]_  = ~A266 & A265;
  assign \new_[58400]_  = ~A203 & \new_[58399]_ ;
  assign \new_[58403]_  = ~A269 & A267;
  assign \new_[58406]_  = A301 & ~A300;
  assign \new_[58407]_  = \new_[58406]_  & \new_[58403]_ ;
  assign \new_[58408]_  = \new_[58407]_  & \new_[58400]_ ;
  assign \new_[58412]_  = ~A168 & ~A169;
  assign \new_[58413]_  = ~A170 & \new_[58412]_ ;
  assign \new_[58417]_  = ~A201 & A166;
  assign \new_[58418]_  = ~A167 & \new_[58417]_ ;
  assign \new_[58419]_  = \new_[58418]_  & \new_[58413]_ ;
  assign \new_[58423]_  = ~A266 & A265;
  assign \new_[58424]_  = ~A203 & \new_[58423]_ ;
  assign \new_[58427]_  = ~A269 & A267;
  assign \new_[58430]_  = ~A302 & ~A300;
  assign \new_[58431]_  = \new_[58430]_  & \new_[58427]_ ;
  assign \new_[58432]_  = \new_[58431]_  & \new_[58424]_ ;
  assign \new_[58436]_  = ~A168 & ~A169;
  assign \new_[58437]_  = ~A170 & \new_[58436]_ ;
  assign \new_[58441]_  = ~A201 & A166;
  assign \new_[58442]_  = ~A167 & \new_[58441]_ ;
  assign \new_[58443]_  = \new_[58442]_  & \new_[58437]_ ;
  assign \new_[58447]_  = ~A266 & A265;
  assign \new_[58448]_  = ~A203 & \new_[58447]_ ;
  assign \new_[58451]_  = ~A269 & A267;
  assign \new_[58454]_  = A299 & A298;
  assign \new_[58455]_  = \new_[58454]_  & \new_[58451]_ ;
  assign \new_[58456]_  = \new_[58455]_  & \new_[58448]_ ;
  assign \new_[58460]_  = ~A168 & ~A169;
  assign \new_[58461]_  = ~A170 & \new_[58460]_ ;
  assign \new_[58465]_  = ~A201 & A166;
  assign \new_[58466]_  = ~A167 & \new_[58465]_ ;
  assign \new_[58467]_  = \new_[58466]_  & \new_[58461]_ ;
  assign \new_[58471]_  = ~A266 & A265;
  assign \new_[58472]_  = ~A203 & \new_[58471]_ ;
  assign \new_[58475]_  = ~A269 & A267;
  assign \new_[58478]_  = ~A299 & ~A298;
  assign \new_[58479]_  = \new_[58478]_  & \new_[58475]_ ;
  assign \new_[58480]_  = \new_[58479]_  & \new_[58472]_ ;
  assign \new_[58484]_  = ~A168 & ~A169;
  assign \new_[58485]_  = ~A170 & \new_[58484]_ ;
  assign \new_[58489]_  = ~A201 & A166;
  assign \new_[58490]_  = ~A167 & \new_[58489]_ ;
  assign \new_[58491]_  = \new_[58490]_  & \new_[58485]_ ;
  assign \new_[58495]_  = ~A266 & ~A265;
  assign \new_[58496]_  = ~A203 & \new_[58495]_ ;
  assign \new_[58499]_  = ~A299 & A298;
  assign \new_[58502]_  = A301 & A300;
  assign \new_[58503]_  = \new_[58502]_  & \new_[58499]_ ;
  assign \new_[58504]_  = \new_[58503]_  & \new_[58496]_ ;
  assign \new_[58508]_  = ~A168 & ~A169;
  assign \new_[58509]_  = ~A170 & \new_[58508]_ ;
  assign \new_[58513]_  = ~A201 & A166;
  assign \new_[58514]_  = ~A167 & \new_[58513]_ ;
  assign \new_[58515]_  = \new_[58514]_  & \new_[58509]_ ;
  assign \new_[58519]_  = ~A266 & ~A265;
  assign \new_[58520]_  = ~A203 & \new_[58519]_ ;
  assign \new_[58523]_  = ~A299 & A298;
  assign \new_[58526]_  = ~A302 & A300;
  assign \new_[58527]_  = \new_[58526]_  & \new_[58523]_ ;
  assign \new_[58528]_  = \new_[58527]_  & \new_[58520]_ ;
  assign \new_[58532]_  = ~A168 & ~A169;
  assign \new_[58533]_  = ~A170 & \new_[58532]_ ;
  assign \new_[58537]_  = ~A201 & A166;
  assign \new_[58538]_  = ~A167 & \new_[58537]_ ;
  assign \new_[58539]_  = \new_[58538]_  & \new_[58533]_ ;
  assign \new_[58543]_  = ~A266 & ~A265;
  assign \new_[58544]_  = ~A203 & \new_[58543]_ ;
  assign \new_[58547]_  = A299 & ~A298;
  assign \new_[58550]_  = A301 & A300;
  assign \new_[58551]_  = \new_[58550]_  & \new_[58547]_ ;
  assign \new_[58552]_  = \new_[58551]_  & \new_[58544]_ ;
  assign \new_[58556]_  = ~A168 & ~A169;
  assign \new_[58557]_  = ~A170 & \new_[58556]_ ;
  assign \new_[58561]_  = ~A201 & A166;
  assign \new_[58562]_  = ~A167 & \new_[58561]_ ;
  assign \new_[58563]_  = \new_[58562]_  & \new_[58557]_ ;
  assign \new_[58567]_  = ~A266 & ~A265;
  assign \new_[58568]_  = ~A203 & \new_[58567]_ ;
  assign \new_[58571]_  = A299 & ~A298;
  assign \new_[58574]_  = ~A302 & A300;
  assign \new_[58575]_  = \new_[58574]_  & \new_[58571]_ ;
  assign \new_[58576]_  = \new_[58575]_  & \new_[58568]_ ;
  assign \new_[58580]_  = ~A168 & ~A169;
  assign \new_[58581]_  = ~A170 & \new_[58580]_ ;
  assign \new_[58585]_  = A199 & A166;
  assign \new_[58586]_  = ~A167 & \new_[58585]_ ;
  assign \new_[58587]_  = \new_[58586]_  & \new_[58581]_ ;
  assign \new_[58591]_  = A268 & ~A267;
  assign \new_[58592]_  = A200 & \new_[58591]_ ;
  assign \new_[58595]_  = ~A299 & A298;
  assign \new_[58598]_  = A301 & A300;
  assign \new_[58599]_  = \new_[58598]_  & \new_[58595]_ ;
  assign \new_[58600]_  = \new_[58599]_  & \new_[58592]_ ;
  assign \new_[58604]_  = ~A168 & ~A169;
  assign \new_[58605]_  = ~A170 & \new_[58604]_ ;
  assign \new_[58609]_  = A199 & A166;
  assign \new_[58610]_  = ~A167 & \new_[58609]_ ;
  assign \new_[58611]_  = \new_[58610]_  & \new_[58605]_ ;
  assign \new_[58615]_  = A268 & ~A267;
  assign \new_[58616]_  = A200 & \new_[58615]_ ;
  assign \new_[58619]_  = ~A299 & A298;
  assign \new_[58622]_  = ~A302 & A300;
  assign \new_[58623]_  = \new_[58622]_  & \new_[58619]_ ;
  assign \new_[58624]_  = \new_[58623]_  & \new_[58616]_ ;
  assign \new_[58628]_  = ~A168 & ~A169;
  assign \new_[58629]_  = ~A170 & \new_[58628]_ ;
  assign \new_[58633]_  = A199 & A166;
  assign \new_[58634]_  = ~A167 & \new_[58633]_ ;
  assign \new_[58635]_  = \new_[58634]_  & \new_[58629]_ ;
  assign \new_[58639]_  = A268 & ~A267;
  assign \new_[58640]_  = A200 & \new_[58639]_ ;
  assign \new_[58643]_  = A299 & ~A298;
  assign \new_[58646]_  = A301 & A300;
  assign \new_[58647]_  = \new_[58646]_  & \new_[58643]_ ;
  assign \new_[58648]_  = \new_[58647]_  & \new_[58640]_ ;
  assign \new_[58652]_  = ~A168 & ~A169;
  assign \new_[58653]_  = ~A170 & \new_[58652]_ ;
  assign \new_[58657]_  = A199 & A166;
  assign \new_[58658]_  = ~A167 & \new_[58657]_ ;
  assign \new_[58659]_  = \new_[58658]_  & \new_[58653]_ ;
  assign \new_[58663]_  = A268 & ~A267;
  assign \new_[58664]_  = A200 & \new_[58663]_ ;
  assign \new_[58667]_  = A299 & ~A298;
  assign \new_[58670]_  = ~A302 & A300;
  assign \new_[58671]_  = \new_[58670]_  & \new_[58667]_ ;
  assign \new_[58672]_  = \new_[58671]_  & \new_[58664]_ ;
  assign \new_[58676]_  = ~A168 & ~A169;
  assign \new_[58677]_  = ~A170 & \new_[58676]_ ;
  assign \new_[58681]_  = A199 & A166;
  assign \new_[58682]_  = ~A167 & \new_[58681]_ ;
  assign \new_[58683]_  = \new_[58682]_  & \new_[58677]_ ;
  assign \new_[58687]_  = ~A269 & ~A267;
  assign \new_[58688]_  = A200 & \new_[58687]_ ;
  assign \new_[58691]_  = ~A299 & A298;
  assign \new_[58694]_  = A301 & A300;
  assign \new_[58695]_  = \new_[58694]_  & \new_[58691]_ ;
  assign \new_[58696]_  = \new_[58695]_  & \new_[58688]_ ;
  assign \new_[58700]_  = ~A168 & ~A169;
  assign \new_[58701]_  = ~A170 & \new_[58700]_ ;
  assign \new_[58705]_  = A199 & A166;
  assign \new_[58706]_  = ~A167 & \new_[58705]_ ;
  assign \new_[58707]_  = \new_[58706]_  & \new_[58701]_ ;
  assign \new_[58711]_  = ~A269 & ~A267;
  assign \new_[58712]_  = A200 & \new_[58711]_ ;
  assign \new_[58715]_  = ~A299 & A298;
  assign \new_[58718]_  = ~A302 & A300;
  assign \new_[58719]_  = \new_[58718]_  & \new_[58715]_ ;
  assign \new_[58720]_  = \new_[58719]_  & \new_[58712]_ ;
  assign \new_[58724]_  = ~A168 & ~A169;
  assign \new_[58725]_  = ~A170 & \new_[58724]_ ;
  assign \new_[58729]_  = A199 & A166;
  assign \new_[58730]_  = ~A167 & \new_[58729]_ ;
  assign \new_[58731]_  = \new_[58730]_  & \new_[58725]_ ;
  assign \new_[58735]_  = ~A269 & ~A267;
  assign \new_[58736]_  = A200 & \new_[58735]_ ;
  assign \new_[58739]_  = A299 & ~A298;
  assign \new_[58742]_  = A301 & A300;
  assign \new_[58743]_  = \new_[58742]_  & \new_[58739]_ ;
  assign \new_[58744]_  = \new_[58743]_  & \new_[58736]_ ;
  assign \new_[58748]_  = ~A168 & ~A169;
  assign \new_[58749]_  = ~A170 & \new_[58748]_ ;
  assign \new_[58753]_  = A199 & A166;
  assign \new_[58754]_  = ~A167 & \new_[58753]_ ;
  assign \new_[58755]_  = \new_[58754]_  & \new_[58749]_ ;
  assign \new_[58759]_  = ~A269 & ~A267;
  assign \new_[58760]_  = A200 & \new_[58759]_ ;
  assign \new_[58763]_  = A299 & ~A298;
  assign \new_[58766]_  = ~A302 & A300;
  assign \new_[58767]_  = \new_[58766]_  & \new_[58763]_ ;
  assign \new_[58768]_  = \new_[58767]_  & \new_[58760]_ ;
  assign \new_[58772]_  = ~A168 & ~A169;
  assign \new_[58773]_  = ~A170 & \new_[58772]_ ;
  assign \new_[58777]_  = A199 & A166;
  assign \new_[58778]_  = ~A167 & \new_[58777]_ ;
  assign \new_[58779]_  = \new_[58778]_  & \new_[58773]_ ;
  assign \new_[58783]_  = A266 & A265;
  assign \new_[58784]_  = A200 & \new_[58783]_ ;
  assign \new_[58787]_  = ~A299 & A298;
  assign \new_[58790]_  = A301 & A300;
  assign \new_[58791]_  = \new_[58790]_  & \new_[58787]_ ;
  assign \new_[58792]_  = \new_[58791]_  & \new_[58784]_ ;
  assign \new_[58796]_  = ~A168 & ~A169;
  assign \new_[58797]_  = ~A170 & \new_[58796]_ ;
  assign \new_[58801]_  = A199 & A166;
  assign \new_[58802]_  = ~A167 & \new_[58801]_ ;
  assign \new_[58803]_  = \new_[58802]_  & \new_[58797]_ ;
  assign \new_[58807]_  = A266 & A265;
  assign \new_[58808]_  = A200 & \new_[58807]_ ;
  assign \new_[58811]_  = ~A299 & A298;
  assign \new_[58814]_  = ~A302 & A300;
  assign \new_[58815]_  = \new_[58814]_  & \new_[58811]_ ;
  assign \new_[58816]_  = \new_[58815]_  & \new_[58808]_ ;
  assign \new_[58820]_  = ~A168 & ~A169;
  assign \new_[58821]_  = ~A170 & \new_[58820]_ ;
  assign \new_[58825]_  = A199 & A166;
  assign \new_[58826]_  = ~A167 & \new_[58825]_ ;
  assign \new_[58827]_  = \new_[58826]_  & \new_[58821]_ ;
  assign \new_[58831]_  = A266 & A265;
  assign \new_[58832]_  = A200 & \new_[58831]_ ;
  assign \new_[58835]_  = A299 & ~A298;
  assign \new_[58838]_  = A301 & A300;
  assign \new_[58839]_  = \new_[58838]_  & \new_[58835]_ ;
  assign \new_[58840]_  = \new_[58839]_  & \new_[58832]_ ;
  assign \new_[58844]_  = ~A168 & ~A169;
  assign \new_[58845]_  = ~A170 & \new_[58844]_ ;
  assign \new_[58849]_  = A199 & A166;
  assign \new_[58850]_  = ~A167 & \new_[58849]_ ;
  assign \new_[58851]_  = \new_[58850]_  & \new_[58845]_ ;
  assign \new_[58855]_  = A266 & A265;
  assign \new_[58856]_  = A200 & \new_[58855]_ ;
  assign \new_[58859]_  = A299 & ~A298;
  assign \new_[58862]_  = ~A302 & A300;
  assign \new_[58863]_  = \new_[58862]_  & \new_[58859]_ ;
  assign \new_[58864]_  = \new_[58863]_  & \new_[58856]_ ;
  assign \new_[58868]_  = ~A168 & ~A169;
  assign \new_[58869]_  = ~A170 & \new_[58868]_ ;
  assign \new_[58873]_  = A199 & A166;
  assign \new_[58874]_  = ~A167 & \new_[58873]_ ;
  assign \new_[58875]_  = \new_[58874]_  & \new_[58869]_ ;
  assign \new_[58879]_  = A266 & ~A265;
  assign \new_[58880]_  = A200 & \new_[58879]_ ;
  assign \new_[58883]_  = A268 & A267;
  assign \new_[58886]_  = A301 & ~A300;
  assign \new_[58887]_  = \new_[58886]_  & \new_[58883]_ ;
  assign \new_[58888]_  = \new_[58887]_  & \new_[58880]_ ;
  assign \new_[58892]_  = ~A168 & ~A169;
  assign \new_[58893]_  = ~A170 & \new_[58892]_ ;
  assign \new_[58897]_  = A199 & A166;
  assign \new_[58898]_  = ~A167 & \new_[58897]_ ;
  assign \new_[58899]_  = \new_[58898]_  & \new_[58893]_ ;
  assign \new_[58903]_  = A266 & ~A265;
  assign \new_[58904]_  = A200 & \new_[58903]_ ;
  assign \new_[58907]_  = A268 & A267;
  assign \new_[58910]_  = ~A302 & ~A300;
  assign \new_[58911]_  = \new_[58910]_  & \new_[58907]_ ;
  assign \new_[58912]_  = \new_[58911]_  & \new_[58904]_ ;
  assign \new_[58916]_  = ~A168 & ~A169;
  assign \new_[58917]_  = ~A170 & \new_[58916]_ ;
  assign \new_[58921]_  = A199 & A166;
  assign \new_[58922]_  = ~A167 & \new_[58921]_ ;
  assign \new_[58923]_  = \new_[58922]_  & \new_[58917]_ ;
  assign \new_[58927]_  = A266 & ~A265;
  assign \new_[58928]_  = A200 & \new_[58927]_ ;
  assign \new_[58931]_  = A268 & A267;
  assign \new_[58934]_  = A299 & A298;
  assign \new_[58935]_  = \new_[58934]_  & \new_[58931]_ ;
  assign \new_[58936]_  = \new_[58935]_  & \new_[58928]_ ;
  assign \new_[58940]_  = ~A168 & ~A169;
  assign \new_[58941]_  = ~A170 & \new_[58940]_ ;
  assign \new_[58945]_  = A199 & A166;
  assign \new_[58946]_  = ~A167 & \new_[58945]_ ;
  assign \new_[58947]_  = \new_[58946]_  & \new_[58941]_ ;
  assign \new_[58951]_  = A266 & ~A265;
  assign \new_[58952]_  = A200 & \new_[58951]_ ;
  assign \new_[58955]_  = A268 & A267;
  assign \new_[58958]_  = ~A299 & ~A298;
  assign \new_[58959]_  = \new_[58958]_  & \new_[58955]_ ;
  assign \new_[58960]_  = \new_[58959]_  & \new_[58952]_ ;
  assign \new_[58964]_  = ~A168 & ~A169;
  assign \new_[58965]_  = ~A170 & \new_[58964]_ ;
  assign \new_[58969]_  = A199 & A166;
  assign \new_[58970]_  = ~A167 & \new_[58969]_ ;
  assign \new_[58971]_  = \new_[58970]_  & \new_[58965]_ ;
  assign \new_[58975]_  = A266 & ~A265;
  assign \new_[58976]_  = A200 & \new_[58975]_ ;
  assign \new_[58979]_  = ~A269 & A267;
  assign \new_[58982]_  = A301 & ~A300;
  assign \new_[58983]_  = \new_[58982]_  & \new_[58979]_ ;
  assign \new_[58984]_  = \new_[58983]_  & \new_[58976]_ ;
  assign \new_[58988]_  = ~A168 & ~A169;
  assign \new_[58989]_  = ~A170 & \new_[58988]_ ;
  assign \new_[58993]_  = A199 & A166;
  assign \new_[58994]_  = ~A167 & \new_[58993]_ ;
  assign \new_[58995]_  = \new_[58994]_  & \new_[58989]_ ;
  assign \new_[58999]_  = A266 & ~A265;
  assign \new_[59000]_  = A200 & \new_[58999]_ ;
  assign \new_[59003]_  = ~A269 & A267;
  assign \new_[59006]_  = ~A302 & ~A300;
  assign \new_[59007]_  = \new_[59006]_  & \new_[59003]_ ;
  assign \new_[59008]_  = \new_[59007]_  & \new_[59000]_ ;
  assign \new_[59012]_  = ~A168 & ~A169;
  assign \new_[59013]_  = ~A170 & \new_[59012]_ ;
  assign \new_[59017]_  = A199 & A166;
  assign \new_[59018]_  = ~A167 & \new_[59017]_ ;
  assign \new_[59019]_  = \new_[59018]_  & \new_[59013]_ ;
  assign \new_[59023]_  = A266 & ~A265;
  assign \new_[59024]_  = A200 & \new_[59023]_ ;
  assign \new_[59027]_  = ~A269 & A267;
  assign \new_[59030]_  = A299 & A298;
  assign \new_[59031]_  = \new_[59030]_  & \new_[59027]_ ;
  assign \new_[59032]_  = \new_[59031]_  & \new_[59024]_ ;
  assign \new_[59036]_  = ~A168 & ~A169;
  assign \new_[59037]_  = ~A170 & \new_[59036]_ ;
  assign \new_[59041]_  = A199 & A166;
  assign \new_[59042]_  = ~A167 & \new_[59041]_ ;
  assign \new_[59043]_  = \new_[59042]_  & \new_[59037]_ ;
  assign \new_[59047]_  = A266 & ~A265;
  assign \new_[59048]_  = A200 & \new_[59047]_ ;
  assign \new_[59051]_  = ~A269 & A267;
  assign \new_[59054]_  = ~A299 & ~A298;
  assign \new_[59055]_  = \new_[59054]_  & \new_[59051]_ ;
  assign \new_[59056]_  = \new_[59055]_  & \new_[59048]_ ;
  assign \new_[59060]_  = ~A168 & ~A169;
  assign \new_[59061]_  = ~A170 & \new_[59060]_ ;
  assign \new_[59065]_  = A199 & A166;
  assign \new_[59066]_  = ~A167 & \new_[59065]_ ;
  assign \new_[59067]_  = \new_[59066]_  & \new_[59061]_ ;
  assign \new_[59071]_  = ~A266 & A265;
  assign \new_[59072]_  = A200 & \new_[59071]_ ;
  assign \new_[59075]_  = A268 & A267;
  assign \new_[59078]_  = A301 & ~A300;
  assign \new_[59079]_  = \new_[59078]_  & \new_[59075]_ ;
  assign \new_[59080]_  = \new_[59079]_  & \new_[59072]_ ;
  assign \new_[59084]_  = ~A168 & ~A169;
  assign \new_[59085]_  = ~A170 & \new_[59084]_ ;
  assign \new_[59089]_  = A199 & A166;
  assign \new_[59090]_  = ~A167 & \new_[59089]_ ;
  assign \new_[59091]_  = \new_[59090]_  & \new_[59085]_ ;
  assign \new_[59095]_  = ~A266 & A265;
  assign \new_[59096]_  = A200 & \new_[59095]_ ;
  assign \new_[59099]_  = A268 & A267;
  assign \new_[59102]_  = ~A302 & ~A300;
  assign \new_[59103]_  = \new_[59102]_  & \new_[59099]_ ;
  assign \new_[59104]_  = \new_[59103]_  & \new_[59096]_ ;
  assign \new_[59108]_  = ~A168 & ~A169;
  assign \new_[59109]_  = ~A170 & \new_[59108]_ ;
  assign \new_[59113]_  = A199 & A166;
  assign \new_[59114]_  = ~A167 & \new_[59113]_ ;
  assign \new_[59115]_  = \new_[59114]_  & \new_[59109]_ ;
  assign \new_[59119]_  = ~A266 & A265;
  assign \new_[59120]_  = A200 & \new_[59119]_ ;
  assign \new_[59123]_  = A268 & A267;
  assign \new_[59126]_  = A299 & A298;
  assign \new_[59127]_  = \new_[59126]_  & \new_[59123]_ ;
  assign \new_[59128]_  = \new_[59127]_  & \new_[59120]_ ;
  assign \new_[59132]_  = ~A168 & ~A169;
  assign \new_[59133]_  = ~A170 & \new_[59132]_ ;
  assign \new_[59137]_  = A199 & A166;
  assign \new_[59138]_  = ~A167 & \new_[59137]_ ;
  assign \new_[59139]_  = \new_[59138]_  & \new_[59133]_ ;
  assign \new_[59143]_  = ~A266 & A265;
  assign \new_[59144]_  = A200 & \new_[59143]_ ;
  assign \new_[59147]_  = A268 & A267;
  assign \new_[59150]_  = ~A299 & ~A298;
  assign \new_[59151]_  = \new_[59150]_  & \new_[59147]_ ;
  assign \new_[59152]_  = \new_[59151]_  & \new_[59144]_ ;
  assign \new_[59156]_  = ~A168 & ~A169;
  assign \new_[59157]_  = ~A170 & \new_[59156]_ ;
  assign \new_[59161]_  = A199 & A166;
  assign \new_[59162]_  = ~A167 & \new_[59161]_ ;
  assign \new_[59163]_  = \new_[59162]_  & \new_[59157]_ ;
  assign \new_[59167]_  = ~A266 & A265;
  assign \new_[59168]_  = A200 & \new_[59167]_ ;
  assign \new_[59171]_  = ~A269 & A267;
  assign \new_[59174]_  = A301 & ~A300;
  assign \new_[59175]_  = \new_[59174]_  & \new_[59171]_ ;
  assign \new_[59176]_  = \new_[59175]_  & \new_[59168]_ ;
  assign \new_[59180]_  = ~A168 & ~A169;
  assign \new_[59181]_  = ~A170 & \new_[59180]_ ;
  assign \new_[59185]_  = A199 & A166;
  assign \new_[59186]_  = ~A167 & \new_[59185]_ ;
  assign \new_[59187]_  = \new_[59186]_  & \new_[59181]_ ;
  assign \new_[59191]_  = ~A266 & A265;
  assign \new_[59192]_  = A200 & \new_[59191]_ ;
  assign \new_[59195]_  = ~A269 & A267;
  assign \new_[59198]_  = ~A302 & ~A300;
  assign \new_[59199]_  = \new_[59198]_  & \new_[59195]_ ;
  assign \new_[59200]_  = \new_[59199]_  & \new_[59192]_ ;
  assign \new_[59204]_  = ~A168 & ~A169;
  assign \new_[59205]_  = ~A170 & \new_[59204]_ ;
  assign \new_[59209]_  = A199 & A166;
  assign \new_[59210]_  = ~A167 & \new_[59209]_ ;
  assign \new_[59211]_  = \new_[59210]_  & \new_[59205]_ ;
  assign \new_[59215]_  = ~A266 & A265;
  assign \new_[59216]_  = A200 & \new_[59215]_ ;
  assign \new_[59219]_  = ~A269 & A267;
  assign \new_[59222]_  = A299 & A298;
  assign \new_[59223]_  = \new_[59222]_  & \new_[59219]_ ;
  assign \new_[59224]_  = \new_[59223]_  & \new_[59216]_ ;
  assign \new_[59228]_  = ~A168 & ~A169;
  assign \new_[59229]_  = ~A170 & \new_[59228]_ ;
  assign \new_[59233]_  = A199 & A166;
  assign \new_[59234]_  = ~A167 & \new_[59233]_ ;
  assign \new_[59235]_  = \new_[59234]_  & \new_[59229]_ ;
  assign \new_[59239]_  = ~A266 & A265;
  assign \new_[59240]_  = A200 & \new_[59239]_ ;
  assign \new_[59243]_  = ~A269 & A267;
  assign \new_[59246]_  = ~A299 & ~A298;
  assign \new_[59247]_  = \new_[59246]_  & \new_[59243]_ ;
  assign \new_[59248]_  = \new_[59247]_  & \new_[59240]_ ;
  assign \new_[59252]_  = ~A168 & ~A169;
  assign \new_[59253]_  = ~A170 & \new_[59252]_ ;
  assign \new_[59257]_  = A199 & A166;
  assign \new_[59258]_  = ~A167 & \new_[59257]_ ;
  assign \new_[59259]_  = \new_[59258]_  & \new_[59253]_ ;
  assign \new_[59263]_  = ~A266 & ~A265;
  assign \new_[59264]_  = A200 & \new_[59263]_ ;
  assign \new_[59267]_  = ~A299 & A298;
  assign \new_[59270]_  = A301 & A300;
  assign \new_[59271]_  = \new_[59270]_  & \new_[59267]_ ;
  assign \new_[59272]_  = \new_[59271]_  & \new_[59264]_ ;
  assign \new_[59276]_  = ~A168 & ~A169;
  assign \new_[59277]_  = ~A170 & \new_[59276]_ ;
  assign \new_[59281]_  = A199 & A166;
  assign \new_[59282]_  = ~A167 & \new_[59281]_ ;
  assign \new_[59283]_  = \new_[59282]_  & \new_[59277]_ ;
  assign \new_[59287]_  = ~A266 & ~A265;
  assign \new_[59288]_  = A200 & \new_[59287]_ ;
  assign \new_[59291]_  = ~A299 & A298;
  assign \new_[59294]_  = ~A302 & A300;
  assign \new_[59295]_  = \new_[59294]_  & \new_[59291]_ ;
  assign \new_[59296]_  = \new_[59295]_  & \new_[59288]_ ;
  assign \new_[59300]_  = ~A168 & ~A169;
  assign \new_[59301]_  = ~A170 & \new_[59300]_ ;
  assign \new_[59305]_  = A199 & A166;
  assign \new_[59306]_  = ~A167 & \new_[59305]_ ;
  assign \new_[59307]_  = \new_[59306]_  & \new_[59301]_ ;
  assign \new_[59311]_  = ~A266 & ~A265;
  assign \new_[59312]_  = A200 & \new_[59311]_ ;
  assign \new_[59315]_  = A299 & ~A298;
  assign \new_[59318]_  = A301 & A300;
  assign \new_[59319]_  = \new_[59318]_  & \new_[59315]_ ;
  assign \new_[59320]_  = \new_[59319]_  & \new_[59312]_ ;
  assign \new_[59324]_  = ~A168 & ~A169;
  assign \new_[59325]_  = ~A170 & \new_[59324]_ ;
  assign \new_[59329]_  = A199 & A166;
  assign \new_[59330]_  = ~A167 & \new_[59329]_ ;
  assign \new_[59331]_  = \new_[59330]_  & \new_[59325]_ ;
  assign \new_[59335]_  = ~A266 & ~A265;
  assign \new_[59336]_  = A200 & \new_[59335]_ ;
  assign \new_[59339]_  = A299 & ~A298;
  assign \new_[59342]_  = ~A302 & A300;
  assign \new_[59343]_  = \new_[59342]_  & \new_[59339]_ ;
  assign \new_[59344]_  = \new_[59343]_  & \new_[59336]_ ;
  assign \new_[59348]_  = ~A168 & ~A169;
  assign \new_[59349]_  = ~A170 & \new_[59348]_ ;
  assign \new_[59353]_  = ~A199 & A166;
  assign \new_[59354]_  = ~A167 & \new_[59353]_ ;
  assign \new_[59355]_  = \new_[59354]_  & \new_[59349]_ ;
  assign \new_[59359]_  = A268 & ~A267;
  assign \new_[59360]_  = ~A200 & \new_[59359]_ ;
  assign \new_[59363]_  = ~A299 & A298;
  assign \new_[59366]_  = A301 & A300;
  assign \new_[59367]_  = \new_[59366]_  & \new_[59363]_ ;
  assign \new_[59368]_  = \new_[59367]_  & \new_[59360]_ ;
  assign \new_[59372]_  = ~A168 & ~A169;
  assign \new_[59373]_  = ~A170 & \new_[59372]_ ;
  assign \new_[59377]_  = ~A199 & A166;
  assign \new_[59378]_  = ~A167 & \new_[59377]_ ;
  assign \new_[59379]_  = \new_[59378]_  & \new_[59373]_ ;
  assign \new_[59383]_  = A268 & ~A267;
  assign \new_[59384]_  = ~A200 & \new_[59383]_ ;
  assign \new_[59387]_  = ~A299 & A298;
  assign \new_[59390]_  = ~A302 & A300;
  assign \new_[59391]_  = \new_[59390]_  & \new_[59387]_ ;
  assign \new_[59392]_  = \new_[59391]_  & \new_[59384]_ ;
  assign \new_[59396]_  = ~A168 & ~A169;
  assign \new_[59397]_  = ~A170 & \new_[59396]_ ;
  assign \new_[59401]_  = ~A199 & A166;
  assign \new_[59402]_  = ~A167 & \new_[59401]_ ;
  assign \new_[59403]_  = \new_[59402]_  & \new_[59397]_ ;
  assign \new_[59407]_  = A268 & ~A267;
  assign \new_[59408]_  = ~A200 & \new_[59407]_ ;
  assign \new_[59411]_  = A299 & ~A298;
  assign \new_[59414]_  = A301 & A300;
  assign \new_[59415]_  = \new_[59414]_  & \new_[59411]_ ;
  assign \new_[59416]_  = \new_[59415]_  & \new_[59408]_ ;
  assign \new_[59420]_  = ~A168 & ~A169;
  assign \new_[59421]_  = ~A170 & \new_[59420]_ ;
  assign \new_[59425]_  = ~A199 & A166;
  assign \new_[59426]_  = ~A167 & \new_[59425]_ ;
  assign \new_[59427]_  = \new_[59426]_  & \new_[59421]_ ;
  assign \new_[59431]_  = A268 & ~A267;
  assign \new_[59432]_  = ~A200 & \new_[59431]_ ;
  assign \new_[59435]_  = A299 & ~A298;
  assign \new_[59438]_  = ~A302 & A300;
  assign \new_[59439]_  = \new_[59438]_  & \new_[59435]_ ;
  assign \new_[59440]_  = \new_[59439]_  & \new_[59432]_ ;
  assign \new_[59444]_  = ~A168 & ~A169;
  assign \new_[59445]_  = ~A170 & \new_[59444]_ ;
  assign \new_[59449]_  = ~A199 & A166;
  assign \new_[59450]_  = ~A167 & \new_[59449]_ ;
  assign \new_[59451]_  = \new_[59450]_  & \new_[59445]_ ;
  assign \new_[59455]_  = ~A269 & ~A267;
  assign \new_[59456]_  = ~A200 & \new_[59455]_ ;
  assign \new_[59459]_  = ~A299 & A298;
  assign \new_[59462]_  = A301 & A300;
  assign \new_[59463]_  = \new_[59462]_  & \new_[59459]_ ;
  assign \new_[59464]_  = \new_[59463]_  & \new_[59456]_ ;
  assign \new_[59468]_  = ~A168 & ~A169;
  assign \new_[59469]_  = ~A170 & \new_[59468]_ ;
  assign \new_[59473]_  = ~A199 & A166;
  assign \new_[59474]_  = ~A167 & \new_[59473]_ ;
  assign \new_[59475]_  = \new_[59474]_  & \new_[59469]_ ;
  assign \new_[59479]_  = ~A269 & ~A267;
  assign \new_[59480]_  = ~A200 & \new_[59479]_ ;
  assign \new_[59483]_  = ~A299 & A298;
  assign \new_[59486]_  = ~A302 & A300;
  assign \new_[59487]_  = \new_[59486]_  & \new_[59483]_ ;
  assign \new_[59488]_  = \new_[59487]_  & \new_[59480]_ ;
  assign \new_[59492]_  = ~A168 & ~A169;
  assign \new_[59493]_  = ~A170 & \new_[59492]_ ;
  assign \new_[59497]_  = ~A199 & A166;
  assign \new_[59498]_  = ~A167 & \new_[59497]_ ;
  assign \new_[59499]_  = \new_[59498]_  & \new_[59493]_ ;
  assign \new_[59503]_  = ~A269 & ~A267;
  assign \new_[59504]_  = ~A200 & \new_[59503]_ ;
  assign \new_[59507]_  = A299 & ~A298;
  assign \new_[59510]_  = A301 & A300;
  assign \new_[59511]_  = \new_[59510]_  & \new_[59507]_ ;
  assign \new_[59512]_  = \new_[59511]_  & \new_[59504]_ ;
  assign \new_[59516]_  = ~A168 & ~A169;
  assign \new_[59517]_  = ~A170 & \new_[59516]_ ;
  assign \new_[59521]_  = ~A199 & A166;
  assign \new_[59522]_  = ~A167 & \new_[59521]_ ;
  assign \new_[59523]_  = \new_[59522]_  & \new_[59517]_ ;
  assign \new_[59527]_  = ~A269 & ~A267;
  assign \new_[59528]_  = ~A200 & \new_[59527]_ ;
  assign \new_[59531]_  = A299 & ~A298;
  assign \new_[59534]_  = ~A302 & A300;
  assign \new_[59535]_  = \new_[59534]_  & \new_[59531]_ ;
  assign \new_[59536]_  = \new_[59535]_  & \new_[59528]_ ;
  assign \new_[59540]_  = ~A168 & ~A169;
  assign \new_[59541]_  = ~A170 & \new_[59540]_ ;
  assign \new_[59545]_  = ~A199 & A166;
  assign \new_[59546]_  = ~A167 & \new_[59545]_ ;
  assign \new_[59547]_  = \new_[59546]_  & \new_[59541]_ ;
  assign \new_[59551]_  = A266 & A265;
  assign \new_[59552]_  = ~A200 & \new_[59551]_ ;
  assign \new_[59555]_  = ~A299 & A298;
  assign \new_[59558]_  = A301 & A300;
  assign \new_[59559]_  = \new_[59558]_  & \new_[59555]_ ;
  assign \new_[59560]_  = \new_[59559]_  & \new_[59552]_ ;
  assign \new_[59564]_  = ~A168 & ~A169;
  assign \new_[59565]_  = ~A170 & \new_[59564]_ ;
  assign \new_[59569]_  = ~A199 & A166;
  assign \new_[59570]_  = ~A167 & \new_[59569]_ ;
  assign \new_[59571]_  = \new_[59570]_  & \new_[59565]_ ;
  assign \new_[59575]_  = A266 & A265;
  assign \new_[59576]_  = ~A200 & \new_[59575]_ ;
  assign \new_[59579]_  = ~A299 & A298;
  assign \new_[59582]_  = ~A302 & A300;
  assign \new_[59583]_  = \new_[59582]_  & \new_[59579]_ ;
  assign \new_[59584]_  = \new_[59583]_  & \new_[59576]_ ;
  assign \new_[59588]_  = ~A168 & ~A169;
  assign \new_[59589]_  = ~A170 & \new_[59588]_ ;
  assign \new_[59593]_  = ~A199 & A166;
  assign \new_[59594]_  = ~A167 & \new_[59593]_ ;
  assign \new_[59595]_  = \new_[59594]_  & \new_[59589]_ ;
  assign \new_[59599]_  = A266 & A265;
  assign \new_[59600]_  = ~A200 & \new_[59599]_ ;
  assign \new_[59603]_  = A299 & ~A298;
  assign \new_[59606]_  = A301 & A300;
  assign \new_[59607]_  = \new_[59606]_  & \new_[59603]_ ;
  assign \new_[59608]_  = \new_[59607]_  & \new_[59600]_ ;
  assign \new_[59612]_  = ~A168 & ~A169;
  assign \new_[59613]_  = ~A170 & \new_[59612]_ ;
  assign \new_[59617]_  = ~A199 & A166;
  assign \new_[59618]_  = ~A167 & \new_[59617]_ ;
  assign \new_[59619]_  = \new_[59618]_  & \new_[59613]_ ;
  assign \new_[59623]_  = A266 & A265;
  assign \new_[59624]_  = ~A200 & \new_[59623]_ ;
  assign \new_[59627]_  = A299 & ~A298;
  assign \new_[59630]_  = ~A302 & A300;
  assign \new_[59631]_  = \new_[59630]_  & \new_[59627]_ ;
  assign \new_[59632]_  = \new_[59631]_  & \new_[59624]_ ;
  assign \new_[59636]_  = ~A168 & ~A169;
  assign \new_[59637]_  = ~A170 & \new_[59636]_ ;
  assign \new_[59641]_  = ~A199 & A166;
  assign \new_[59642]_  = ~A167 & \new_[59641]_ ;
  assign \new_[59643]_  = \new_[59642]_  & \new_[59637]_ ;
  assign \new_[59647]_  = A266 & ~A265;
  assign \new_[59648]_  = ~A200 & \new_[59647]_ ;
  assign \new_[59651]_  = A268 & A267;
  assign \new_[59654]_  = A301 & ~A300;
  assign \new_[59655]_  = \new_[59654]_  & \new_[59651]_ ;
  assign \new_[59656]_  = \new_[59655]_  & \new_[59648]_ ;
  assign \new_[59660]_  = ~A168 & ~A169;
  assign \new_[59661]_  = ~A170 & \new_[59660]_ ;
  assign \new_[59665]_  = ~A199 & A166;
  assign \new_[59666]_  = ~A167 & \new_[59665]_ ;
  assign \new_[59667]_  = \new_[59666]_  & \new_[59661]_ ;
  assign \new_[59671]_  = A266 & ~A265;
  assign \new_[59672]_  = ~A200 & \new_[59671]_ ;
  assign \new_[59675]_  = A268 & A267;
  assign \new_[59678]_  = ~A302 & ~A300;
  assign \new_[59679]_  = \new_[59678]_  & \new_[59675]_ ;
  assign \new_[59680]_  = \new_[59679]_  & \new_[59672]_ ;
  assign \new_[59684]_  = ~A168 & ~A169;
  assign \new_[59685]_  = ~A170 & \new_[59684]_ ;
  assign \new_[59689]_  = ~A199 & A166;
  assign \new_[59690]_  = ~A167 & \new_[59689]_ ;
  assign \new_[59691]_  = \new_[59690]_  & \new_[59685]_ ;
  assign \new_[59695]_  = A266 & ~A265;
  assign \new_[59696]_  = ~A200 & \new_[59695]_ ;
  assign \new_[59699]_  = A268 & A267;
  assign \new_[59702]_  = A299 & A298;
  assign \new_[59703]_  = \new_[59702]_  & \new_[59699]_ ;
  assign \new_[59704]_  = \new_[59703]_  & \new_[59696]_ ;
  assign \new_[59708]_  = ~A168 & ~A169;
  assign \new_[59709]_  = ~A170 & \new_[59708]_ ;
  assign \new_[59713]_  = ~A199 & A166;
  assign \new_[59714]_  = ~A167 & \new_[59713]_ ;
  assign \new_[59715]_  = \new_[59714]_  & \new_[59709]_ ;
  assign \new_[59719]_  = A266 & ~A265;
  assign \new_[59720]_  = ~A200 & \new_[59719]_ ;
  assign \new_[59723]_  = A268 & A267;
  assign \new_[59726]_  = ~A299 & ~A298;
  assign \new_[59727]_  = \new_[59726]_  & \new_[59723]_ ;
  assign \new_[59728]_  = \new_[59727]_  & \new_[59720]_ ;
  assign \new_[59732]_  = ~A168 & ~A169;
  assign \new_[59733]_  = ~A170 & \new_[59732]_ ;
  assign \new_[59737]_  = ~A199 & A166;
  assign \new_[59738]_  = ~A167 & \new_[59737]_ ;
  assign \new_[59739]_  = \new_[59738]_  & \new_[59733]_ ;
  assign \new_[59743]_  = A266 & ~A265;
  assign \new_[59744]_  = ~A200 & \new_[59743]_ ;
  assign \new_[59747]_  = ~A269 & A267;
  assign \new_[59750]_  = A301 & ~A300;
  assign \new_[59751]_  = \new_[59750]_  & \new_[59747]_ ;
  assign \new_[59752]_  = \new_[59751]_  & \new_[59744]_ ;
  assign \new_[59756]_  = ~A168 & ~A169;
  assign \new_[59757]_  = ~A170 & \new_[59756]_ ;
  assign \new_[59761]_  = ~A199 & A166;
  assign \new_[59762]_  = ~A167 & \new_[59761]_ ;
  assign \new_[59763]_  = \new_[59762]_  & \new_[59757]_ ;
  assign \new_[59767]_  = A266 & ~A265;
  assign \new_[59768]_  = ~A200 & \new_[59767]_ ;
  assign \new_[59771]_  = ~A269 & A267;
  assign \new_[59774]_  = ~A302 & ~A300;
  assign \new_[59775]_  = \new_[59774]_  & \new_[59771]_ ;
  assign \new_[59776]_  = \new_[59775]_  & \new_[59768]_ ;
  assign \new_[59780]_  = ~A168 & ~A169;
  assign \new_[59781]_  = ~A170 & \new_[59780]_ ;
  assign \new_[59785]_  = ~A199 & A166;
  assign \new_[59786]_  = ~A167 & \new_[59785]_ ;
  assign \new_[59787]_  = \new_[59786]_  & \new_[59781]_ ;
  assign \new_[59791]_  = A266 & ~A265;
  assign \new_[59792]_  = ~A200 & \new_[59791]_ ;
  assign \new_[59795]_  = ~A269 & A267;
  assign \new_[59798]_  = A299 & A298;
  assign \new_[59799]_  = \new_[59798]_  & \new_[59795]_ ;
  assign \new_[59800]_  = \new_[59799]_  & \new_[59792]_ ;
  assign \new_[59804]_  = ~A168 & ~A169;
  assign \new_[59805]_  = ~A170 & \new_[59804]_ ;
  assign \new_[59809]_  = ~A199 & A166;
  assign \new_[59810]_  = ~A167 & \new_[59809]_ ;
  assign \new_[59811]_  = \new_[59810]_  & \new_[59805]_ ;
  assign \new_[59815]_  = A266 & ~A265;
  assign \new_[59816]_  = ~A200 & \new_[59815]_ ;
  assign \new_[59819]_  = ~A269 & A267;
  assign \new_[59822]_  = ~A299 & ~A298;
  assign \new_[59823]_  = \new_[59822]_  & \new_[59819]_ ;
  assign \new_[59824]_  = \new_[59823]_  & \new_[59816]_ ;
  assign \new_[59828]_  = ~A168 & ~A169;
  assign \new_[59829]_  = ~A170 & \new_[59828]_ ;
  assign \new_[59833]_  = ~A199 & A166;
  assign \new_[59834]_  = ~A167 & \new_[59833]_ ;
  assign \new_[59835]_  = \new_[59834]_  & \new_[59829]_ ;
  assign \new_[59839]_  = ~A266 & A265;
  assign \new_[59840]_  = ~A200 & \new_[59839]_ ;
  assign \new_[59843]_  = A268 & A267;
  assign \new_[59846]_  = A301 & ~A300;
  assign \new_[59847]_  = \new_[59846]_  & \new_[59843]_ ;
  assign \new_[59848]_  = \new_[59847]_  & \new_[59840]_ ;
  assign \new_[59852]_  = ~A168 & ~A169;
  assign \new_[59853]_  = ~A170 & \new_[59852]_ ;
  assign \new_[59857]_  = ~A199 & A166;
  assign \new_[59858]_  = ~A167 & \new_[59857]_ ;
  assign \new_[59859]_  = \new_[59858]_  & \new_[59853]_ ;
  assign \new_[59863]_  = ~A266 & A265;
  assign \new_[59864]_  = ~A200 & \new_[59863]_ ;
  assign \new_[59867]_  = A268 & A267;
  assign \new_[59870]_  = ~A302 & ~A300;
  assign \new_[59871]_  = \new_[59870]_  & \new_[59867]_ ;
  assign \new_[59872]_  = \new_[59871]_  & \new_[59864]_ ;
  assign \new_[59876]_  = ~A168 & ~A169;
  assign \new_[59877]_  = ~A170 & \new_[59876]_ ;
  assign \new_[59881]_  = ~A199 & A166;
  assign \new_[59882]_  = ~A167 & \new_[59881]_ ;
  assign \new_[59883]_  = \new_[59882]_  & \new_[59877]_ ;
  assign \new_[59887]_  = ~A266 & A265;
  assign \new_[59888]_  = ~A200 & \new_[59887]_ ;
  assign \new_[59891]_  = A268 & A267;
  assign \new_[59894]_  = A299 & A298;
  assign \new_[59895]_  = \new_[59894]_  & \new_[59891]_ ;
  assign \new_[59896]_  = \new_[59895]_  & \new_[59888]_ ;
  assign \new_[59900]_  = ~A168 & ~A169;
  assign \new_[59901]_  = ~A170 & \new_[59900]_ ;
  assign \new_[59905]_  = ~A199 & A166;
  assign \new_[59906]_  = ~A167 & \new_[59905]_ ;
  assign \new_[59907]_  = \new_[59906]_  & \new_[59901]_ ;
  assign \new_[59911]_  = ~A266 & A265;
  assign \new_[59912]_  = ~A200 & \new_[59911]_ ;
  assign \new_[59915]_  = A268 & A267;
  assign \new_[59918]_  = ~A299 & ~A298;
  assign \new_[59919]_  = \new_[59918]_  & \new_[59915]_ ;
  assign \new_[59920]_  = \new_[59919]_  & \new_[59912]_ ;
  assign \new_[59924]_  = ~A168 & ~A169;
  assign \new_[59925]_  = ~A170 & \new_[59924]_ ;
  assign \new_[59929]_  = ~A199 & A166;
  assign \new_[59930]_  = ~A167 & \new_[59929]_ ;
  assign \new_[59931]_  = \new_[59930]_  & \new_[59925]_ ;
  assign \new_[59935]_  = ~A266 & A265;
  assign \new_[59936]_  = ~A200 & \new_[59935]_ ;
  assign \new_[59939]_  = ~A269 & A267;
  assign \new_[59942]_  = A301 & ~A300;
  assign \new_[59943]_  = \new_[59942]_  & \new_[59939]_ ;
  assign \new_[59944]_  = \new_[59943]_  & \new_[59936]_ ;
  assign \new_[59948]_  = ~A168 & ~A169;
  assign \new_[59949]_  = ~A170 & \new_[59948]_ ;
  assign \new_[59953]_  = ~A199 & A166;
  assign \new_[59954]_  = ~A167 & \new_[59953]_ ;
  assign \new_[59955]_  = \new_[59954]_  & \new_[59949]_ ;
  assign \new_[59959]_  = ~A266 & A265;
  assign \new_[59960]_  = ~A200 & \new_[59959]_ ;
  assign \new_[59963]_  = ~A269 & A267;
  assign \new_[59966]_  = ~A302 & ~A300;
  assign \new_[59967]_  = \new_[59966]_  & \new_[59963]_ ;
  assign \new_[59968]_  = \new_[59967]_  & \new_[59960]_ ;
  assign \new_[59972]_  = ~A168 & ~A169;
  assign \new_[59973]_  = ~A170 & \new_[59972]_ ;
  assign \new_[59977]_  = ~A199 & A166;
  assign \new_[59978]_  = ~A167 & \new_[59977]_ ;
  assign \new_[59979]_  = \new_[59978]_  & \new_[59973]_ ;
  assign \new_[59983]_  = ~A266 & A265;
  assign \new_[59984]_  = ~A200 & \new_[59983]_ ;
  assign \new_[59987]_  = ~A269 & A267;
  assign \new_[59990]_  = A299 & A298;
  assign \new_[59991]_  = \new_[59990]_  & \new_[59987]_ ;
  assign \new_[59992]_  = \new_[59991]_  & \new_[59984]_ ;
  assign \new_[59996]_  = ~A168 & ~A169;
  assign \new_[59997]_  = ~A170 & \new_[59996]_ ;
  assign \new_[60001]_  = ~A199 & A166;
  assign \new_[60002]_  = ~A167 & \new_[60001]_ ;
  assign \new_[60003]_  = \new_[60002]_  & \new_[59997]_ ;
  assign \new_[60007]_  = ~A266 & A265;
  assign \new_[60008]_  = ~A200 & \new_[60007]_ ;
  assign \new_[60011]_  = ~A269 & A267;
  assign \new_[60014]_  = ~A299 & ~A298;
  assign \new_[60015]_  = \new_[60014]_  & \new_[60011]_ ;
  assign \new_[60016]_  = \new_[60015]_  & \new_[60008]_ ;
  assign \new_[60020]_  = ~A168 & ~A169;
  assign \new_[60021]_  = ~A170 & \new_[60020]_ ;
  assign \new_[60025]_  = ~A199 & A166;
  assign \new_[60026]_  = ~A167 & \new_[60025]_ ;
  assign \new_[60027]_  = \new_[60026]_  & \new_[60021]_ ;
  assign \new_[60031]_  = ~A266 & ~A265;
  assign \new_[60032]_  = ~A200 & \new_[60031]_ ;
  assign \new_[60035]_  = ~A299 & A298;
  assign \new_[60038]_  = A301 & A300;
  assign \new_[60039]_  = \new_[60038]_  & \new_[60035]_ ;
  assign \new_[60040]_  = \new_[60039]_  & \new_[60032]_ ;
  assign \new_[60044]_  = ~A168 & ~A169;
  assign \new_[60045]_  = ~A170 & \new_[60044]_ ;
  assign \new_[60049]_  = ~A199 & A166;
  assign \new_[60050]_  = ~A167 & \new_[60049]_ ;
  assign \new_[60051]_  = \new_[60050]_  & \new_[60045]_ ;
  assign \new_[60055]_  = ~A266 & ~A265;
  assign \new_[60056]_  = ~A200 & \new_[60055]_ ;
  assign \new_[60059]_  = ~A299 & A298;
  assign \new_[60062]_  = ~A302 & A300;
  assign \new_[60063]_  = \new_[60062]_  & \new_[60059]_ ;
  assign \new_[60064]_  = \new_[60063]_  & \new_[60056]_ ;
  assign \new_[60068]_  = ~A168 & ~A169;
  assign \new_[60069]_  = ~A170 & \new_[60068]_ ;
  assign \new_[60073]_  = ~A199 & A166;
  assign \new_[60074]_  = ~A167 & \new_[60073]_ ;
  assign \new_[60075]_  = \new_[60074]_  & \new_[60069]_ ;
  assign \new_[60079]_  = ~A266 & ~A265;
  assign \new_[60080]_  = ~A200 & \new_[60079]_ ;
  assign \new_[60083]_  = A299 & ~A298;
  assign \new_[60086]_  = A301 & A300;
  assign \new_[60087]_  = \new_[60086]_  & \new_[60083]_ ;
  assign \new_[60088]_  = \new_[60087]_  & \new_[60080]_ ;
  assign \new_[60092]_  = ~A168 & ~A169;
  assign \new_[60093]_  = ~A170 & \new_[60092]_ ;
  assign \new_[60097]_  = ~A199 & A166;
  assign \new_[60098]_  = ~A167 & \new_[60097]_ ;
  assign \new_[60099]_  = \new_[60098]_  & \new_[60093]_ ;
  assign \new_[60103]_  = ~A266 & ~A265;
  assign \new_[60104]_  = ~A200 & \new_[60103]_ ;
  assign \new_[60107]_  = A299 & ~A298;
  assign \new_[60110]_  = ~A302 & A300;
  assign \new_[60111]_  = \new_[60110]_  & \new_[60107]_ ;
  assign \new_[60112]_  = \new_[60111]_  & \new_[60104]_ ;
  assign \new_[60116]_  = ~A199 & A166;
  assign \new_[60117]_  = A167 & \new_[60116]_ ;
  assign \new_[60120]_  = A201 & A200;
  assign \new_[60123]_  = ~A265 & A202;
  assign \new_[60124]_  = \new_[60123]_  & \new_[60120]_ ;
  assign \new_[60125]_  = \new_[60124]_  & \new_[60117]_ ;
  assign \new_[60129]_  = A268 & A267;
  assign \new_[60130]_  = A266 & \new_[60129]_ ;
  assign \new_[60133]_  = ~A299 & A298;
  assign \new_[60136]_  = A301 & A300;
  assign \new_[60137]_  = \new_[60136]_  & \new_[60133]_ ;
  assign \new_[60138]_  = \new_[60137]_  & \new_[60130]_ ;
  assign \new_[60142]_  = ~A199 & A166;
  assign \new_[60143]_  = A167 & \new_[60142]_ ;
  assign \new_[60146]_  = A201 & A200;
  assign \new_[60149]_  = ~A265 & A202;
  assign \new_[60150]_  = \new_[60149]_  & \new_[60146]_ ;
  assign \new_[60151]_  = \new_[60150]_  & \new_[60143]_ ;
  assign \new_[60155]_  = A268 & A267;
  assign \new_[60156]_  = A266 & \new_[60155]_ ;
  assign \new_[60159]_  = ~A299 & A298;
  assign \new_[60162]_  = ~A302 & A300;
  assign \new_[60163]_  = \new_[60162]_  & \new_[60159]_ ;
  assign \new_[60164]_  = \new_[60163]_  & \new_[60156]_ ;
  assign \new_[60168]_  = ~A199 & A166;
  assign \new_[60169]_  = A167 & \new_[60168]_ ;
  assign \new_[60172]_  = A201 & A200;
  assign \new_[60175]_  = ~A265 & A202;
  assign \new_[60176]_  = \new_[60175]_  & \new_[60172]_ ;
  assign \new_[60177]_  = \new_[60176]_  & \new_[60169]_ ;
  assign \new_[60181]_  = A268 & A267;
  assign \new_[60182]_  = A266 & \new_[60181]_ ;
  assign \new_[60185]_  = A299 & ~A298;
  assign \new_[60188]_  = A301 & A300;
  assign \new_[60189]_  = \new_[60188]_  & \new_[60185]_ ;
  assign \new_[60190]_  = \new_[60189]_  & \new_[60182]_ ;
  assign \new_[60194]_  = ~A199 & A166;
  assign \new_[60195]_  = A167 & \new_[60194]_ ;
  assign \new_[60198]_  = A201 & A200;
  assign \new_[60201]_  = ~A265 & A202;
  assign \new_[60202]_  = \new_[60201]_  & \new_[60198]_ ;
  assign \new_[60203]_  = \new_[60202]_  & \new_[60195]_ ;
  assign \new_[60207]_  = A268 & A267;
  assign \new_[60208]_  = A266 & \new_[60207]_ ;
  assign \new_[60211]_  = A299 & ~A298;
  assign \new_[60214]_  = ~A302 & A300;
  assign \new_[60215]_  = \new_[60214]_  & \new_[60211]_ ;
  assign \new_[60216]_  = \new_[60215]_  & \new_[60208]_ ;
  assign \new_[60220]_  = ~A199 & A166;
  assign \new_[60221]_  = A167 & \new_[60220]_ ;
  assign \new_[60224]_  = A201 & A200;
  assign \new_[60227]_  = ~A265 & A202;
  assign \new_[60228]_  = \new_[60227]_  & \new_[60224]_ ;
  assign \new_[60229]_  = \new_[60228]_  & \new_[60221]_ ;
  assign \new_[60233]_  = ~A269 & A267;
  assign \new_[60234]_  = A266 & \new_[60233]_ ;
  assign \new_[60237]_  = ~A299 & A298;
  assign \new_[60240]_  = A301 & A300;
  assign \new_[60241]_  = \new_[60240]_  & \new_[60237]_ ;
  assign \new_[60242]_  = \new_[60241]_  & \new_[60234]_ ;
  assign \new_[60246]_  = ~A199 & A166;
  assign \new_[60247]_  = A167 & \new_[60246]_ ;
  assign \new_[60250]_  = A201 & A200;
  assign \new_[60253]_  = ~A265 & A202;
  assign \new_[60254]_  = \new_[60253]_  & \new_[60250]_ ;
  assign \new_[60255]_  = \new_[60254]_  & \new_[60247]_ ;
  assign \new_[60259]_  = ~A269 & A267;
  assign \new_[60260]_  = A266 & \new_[60259]_ ;
  assign \new_[60263]_  = ~A299 & A298;
  assign \new_[60266]_  = ~A302 & A300;
  assign \new_[60267]_  = \new_[60266]_  & \new_[60263]_ ;
  assign \new_[60268]_  = \new_[60267]_  & \new_[60260]_ ;
  assign \new_[60272]_  = ~A199 & A166;
  assign \new_[60273]_  = A167 & \new_[60272]_ ;
  assign \new_[60276]_  = A201 & A200;
  assign \new_[60279]_  = ~A265 & A202;
  assign \new_[60280]_  = \new_[60279]_  & \new_[60276]_ ;
  assign \new_[60281]_  = \new_[60280]_  & \new_[60273]_ ;
  assign \new_[60285]_  = ~A269 & A267;
  assign \new_[60286]_  = A266 & \new_[60285]_ ;
  assign \new_[60289]_  = A299 & ~A298;
  assign \new_[60292]_  = A301 & A300;
  assign \new_[60293]_  = \new_[60292]_  & \new_[60289]_ ;
  assign \new_[60294]_  = \new_[60293]_  & \new_[60286]_ ;
  assign \new_[60298]_  = ~A199 & A166;
  assign \new_[60299]_  = A167 & \new_[60298]_ ;
  assign \new_[60302]_  = A201 & A200;
  assign \new_[60305]_  = ~A265 & A202;
  assign \new_[60306]_  = \new_[60305]_  & \new_[60302]_ ;
  assign \new_[60307]_  = \new_[60306]_  & \new_[60299]_ ;
  assign \new_[60311]_  = ~A269 & A267;
  assign \new_[60312]_  = A266 & \new_[60311]_ ;
  assign \new_[60315]_  = A299 & ~A298;
  assign \new_[60318]_  = ~A302 & A300;
  assign \new_[60319]_  = \new_[60318]_  & \new_[60315]_ ;
  assign \new_[60320]_  = \new_[60319]_  & \new_[60312]_ ;
  assign \new_[60324]_  = ~A199 & A166;
  assign \new_[60325]_  = A167 & \new_[60324]_ ;
  assign \new_[60328]_  = A201 & A200;
  assign \new_[60331]_  = A265 & A202;
  assign \new_[60332]_  = \new_[60331]_  & \new_[60328]_ ;
  assign \new_[60333]_  = \new_[60332]_  & \new_[60325]_ ;
  assign \new_[60337]_  = A268 & A267;
  assign \new_[60338]_  = ~A266 & \new_[60337]_ ;
  assign \new_[60341]_  = ~A299 & A298;
  assign \new_[60344]_  = A301 & A300;
  assign \new_[60345]_  = \new_[60344]_  & \new_[60341]_ ;
  assign \new_[60346]_  = \new_[60345]_  & \new_[60338]_ ;
  assign \new_[60350]_  = ~A199 & A166;
  assign \new_[60351]_  = A167 & \new_[60350]_ ;
  assign \new_[60354]_  = A201 & A200;
  assign \new_[60357]_  = A265 & A202;
  assign \new_[60358]_  = \new_[60357]_  & \new_[60354]_ ;
  assign \new_[60359]_  = \new_[60358]_  & \new_[60351]_ ;
  assign \new_[60363]_  = A268 & A267;
  assign \new_[60364]_  = ~A266 & \new_[60363]_ ;
  assign \new_[60367]_  = ~A299 & A298;
  assign \new_[60370]_  = ~A302 & A300;
  assign \new_[60371]_  = \new_[60370]_  & \new_[60367]_ ;
  assign \new_[60372]_  = \new_[60371]_  & \new_[60364]_ ;
  assign \new_[60376]_  = ~A199 & A166;
  assign \new_[60377]_  = A167 & \new_[60376]_ ;
  assign \new_[60380]_  = A201 & A200;
  assign \new_[60383]_  = A265 & A202;
  assign \new_[60384]_  = \new_[60383]_  & \new_[60380]_ ;
  assign \new_[60385]_  = \new_[60384]_  & \new_[60377]_ ;
  assign \new_[60389]_  = A268 & A267;
  assign \new_[60390]_  = ~A266 & \new_[60389]_ ;
  assign \new_[60393]_  = A299 & ~A298;
  assign \new_[60396]_  = A301 & A300;
  assign \new_[60397]_  = \new_[60396]_  & \new_[60393]_ ;
  assign \new_[60398]_  = \new_[60397]_  & \new_[60390]_ ;
  assign \new_[60402]_  = ~A199 & A166;
  assign \new_[60403]_  = A167 & \new_[60402]_ ;
  assign \new_[60406]_  = A201 & A200;
  assign \new_[60409]_  = A265 & A202;
  assign \new_[60410]_  = \new_[60409]_  & \new_[60406]_ ;
  assign \new_[60411]_  = \new_[60410]_  & \new_[60403]_ ;
  assign \new_[60415]_  = A268 & A267;
  assign \new_[60416]_  = ~A266 & \new_[60415]_ ;
  assign \new_[60419]_  = A299 & ~A298;
  assign \new_[60422]_  = ~A302 & A300;
  assign \new_[60423]_  = \new_[60422]_  & \new_[60419]_ ;
  assign \new_[60424]_  = \new_[60423]_  & \new_[60416]_ ;
  assign \new_[60428]_  = ~A199 & A166;
  assign \new_[60429]_  = A167 & \new_[60428]_ ;
  assign \new_[60432]_  = A201 & A200;
  assign \new_[60435]_  = A265 & A202;
  assign \new_[60436]_  = \new_[60435]_  & \new_[60432]_ ;
  assign \new_[60437]_  = \new_[60436]_  & \new_[60429]_ ;
  assign \new_[60441]_  = ~A269 & A267;
  assign \new_[60442]_  = ~A266 & \new_[60441]_ ;
  assign \new_[60445]_  = ~A299 & A298;
  assign \new_[60448]_  = A301 & A300;
  assign \new_[60449]_  = \new_[60448]_  & \new_[60445]_ ;
  assign \new_[60450]_  = \new_[60449]_  & \new_[60442]_ ;
  assign \new_[60454]_  = ~A199 & A166;
  assign \new_[60455]_  = A167 & \new_[60454]_ ;
  assign \new_[60458]_  = A201 & A200;
  assign \new_[60461]_  = A265 & A202;
  assign \new_[60462]_  = \new_[60461]_  & \new_[60458]_ ;
  assign \new_[60463]_  = \new_[60462]_  & \new_[60455]_ ;
  assign \new_[60467]_  = ~A269 & A267;
  assign \new_[60468]_  = ~A266 & \new_[60467]_ ;
  assign \new_[60471]_  = ~A299 & A298;
  assign \new_[60474]_  = ~A302 & A300;
  assign \new_[60475]_  = \new_[60474]_  & \new_[60471]_ ;
  assign \new_[60476]_  = \new_[60475]_  & \new_[60468]_ ;
  assign \new_[60480]_  = ~A199 & A166;
  assign \new_[60481]_  = A167 & \new_[60480]_ ;
  assign \new_[60484]_  = A201 & A200;
  assign \new_[60487]_  = A265 & A202;
  assign \new_[60488]_  = \new_[60487]_  & \new_[60484]_ ;
  assign \new_[60489]_  = \new_[60488]_  & \new_[60481]_ ;
  assign \new_[60493]_  = ~A269 & A267;
  assign \new_[60494]_  = ~A266 & \new_[60493]_ ;
  assign \new_[60497]_  = A299 & ~A298;
  assign \new_[60500]_  = A301 & A300;
  assign \new_[60501]_  = \new_[60500]_  & \new_[60497]_ ;
  assign \new_[60502]_  = \new_[60501]_  & \new_[60494]_ ;
  assign \new_[60506]_  = ~A199 & A166;
  assign \new_[60507]_  = A167 & \new_[60506]_ ;
  assign \new_[60510]_  = A201 & A200;
  assign \new_[60513]_  = A265 & A202;
  assign \new_[60514]_  = \new_[60513]_  & \new_[60510]_ ;
  assign \new_[60515]_  = \new_[60514]_  & \new_[60507]_ ;
  assign \new_[60519]_  = ~A269 & A267;
  assign \new_[60520]_  = ~A266 & \new_[60519]_ ;
  assign \new_[60523]_  = A299 & ~A298;
  assign \new_[60526]_  = ~A302 & A300;
  assign \new_[60527]_  = \new_[60526]_  & \new_[60523]_ ;
  assign \new_[60528]_  = \new_[60527]_  & \new_[60520]_ ;
  assign \new_[60532]_  = ~A199 & A166;
  assign \new_[60533]_  = A167 & \new_[60532]_ ;
  assign \new_[60536]_  = A201 & A200;
  assign \new_[60539]_  = ~A265 & ~A203;
  assign \new_[60540]_  = \new_[60539]_  & \new_[60536]_ ;
  assign \new_[60541]_  = \new_[60540]_  & \new_[60533]_ ;
  assign \new_[60545]_  = A268 & A267;
  assign \new_[60546]_  = A266 & \new_[60545]_ ;
  assign \new_[60549]_  = ~A299 & A298;
  assign \new_[60552]_  = A301 & A300;
  assign \new_[60553]_  = \new_[60552]_  & \new_[60549]_ ;
  assign \new_[60554]_  = \new_[60553]_  & \new_[60546]_ ;
  assign \new_[60558]_  = ~A199 & A166;
  assign \new_[60559]_  = A167 & \new_[60558]_ ;
  assign \new_[60562]_  = A201 & A200;
  assign \new_[60565]_  = ~A265 & ~A203;
  assign \new_[60566]_  = \new_[60565]_  & \new_[60562]_ ;
  assign \new_[60567]_  = \new_[60566]_  & \new_[60559]_ ;
  assign \new_[60571]_  = A268 & A267;
  assign \new_[60572]_  = A266 & \new_[60571]_ ;
  assign \new_[60575]_  = ~A299 & A298;
  assign \new_[60578]_  = ~A302 & A300;
  assign \new_[60579]_  = \new_[60578]_  & \new_[60575]_ ;
  assign \new_[60580]_  = \new_[60579]_  & \new_[60572]_ ;
  assign \new_[60584]_  = ~A199 & A166;
  assign \new_[60585]_  = A167 & \new_[60584]_ ;
  assign \new_[60588]_  = A201 & A200;
  assign \new_[60591]_  = ~A265 & ~A203;
  assign \new_[60592]_  = \new_[60591]_  & \new_[60588]_ ;
  assign \new_[60593]_  = \new_[60592]_  & \new_[60585]_ ;
  assign \new_[60597]_  = A268 & A267;
  assign \new_[60598]_  = A266 & \new_[60597]_ ;
  assign \new_[60601]_  = A299 & ~A298;
  assign \new_[60604]_  = A301 & A300;
  assign \new_[60605]_  = \new_[60604]_  & \new_[60601]_ ;
  assign \new_[60606]_  = \new_[60605]_  & \new_[60598]_ ;
  assign \new_[60610]_  = ~A199 & A166;
  assign \new_[60611]_  = A167 & \new_[60610]_ ;
  assign \new_[60614]_  = A201 & A200;
  assign \new_[60617]_  = ~A265 & ~A203;
  assign \new_[60618]_  = \new_[60617]_  & \new_[60614]_ ;
  assign \new_[60619]_  = \new_[60618]_  & \new_[60611]_ ;
  assign \new_[60623]_  = A268 & A267;
  assign \new_[60624]_  = A266 & \new_[60623]_ ;
  assign \new_[60627]_  = A299 & ~A298;
  assign \new_[60630]_  = ~A302 & A300;
  assign \new_[60631]_  = \new_[60630]_  & \new_[60627]_ ;
  assign \new_[60632]_  = \new_[60631]_  & \new_[60624]_ ;
  assign \new_[60636]_  = ~A199 & A166;
  assign \new_[60637]_  = A167 & \new_[60636]_ ;
  assign \new_[60640]_  = A201 & A200;
  assign \new_[60643]_  = ~A265 & ~A203;
  assign \new_[60644]_  = \new_[60643]_  & \new_[60640]_ ;
  assign \new_[60645]_  = \new_[60644]_  & \new_[60637]_ ;
  assign \new_[60649]_  = ~A269 & A267;
  assign \new_[60650]_  = A266 & \new_[60649]_ ;
  assign \new_[60653]_  = ~A299 & A298;
  assign \new_[60656]_  = A301 & A300;
  assign \new_[60657]_  = \new_[60656]_  & \new_[60653]_ ;
  assign \new_[60658]_  = \new_[60657]_  & \new_[60650]_ ;
  assign \new_[60662]_  = ~A199 & A166;
  assign \new_[60663]_  = A167 & \new_[60662]_ ;
  assign \new_[60666]_  = A201 & A200;
  assign \new_[60669]_  = ~A265 & ~A203;
  assign \new_[60670]_  = \new_[60669]_  & \new_[60666]_ ;
  assign \new_[60671]_  = \new_[60670]_  & \new_[60663]_ ;
  assign \new_[60675]_  = ~A269 & A267;
  assign \new_[60676]_  = A266 & \new_[60675]_ ;
  assign \new_[60679]_  = ~A299 & A298;
  assign \new_[60682]_  = ~A302 & A300;
  assign \new_[60683]_  = \new_[60682]_  & \new_[60679]_ ;
  assign \new_[60684]_  = \new_[60683]_  & \new_[60676]_ ;
  assign \new_[60688]_  = ~A199 & A166;
  assign \new_[60689]_  = A167 & \new_[60688]_ ;
  assign \new_[60692]_  = A201 & A200;
  assign \new_[60695]_  = ~A265 & ~A203;
  assign \new_[60696]_  = \new_[60695]_  & \new_[60692]_ ;
  assign \new_[60697]_  = \new_[60696]_  & \new_[60689]_ ;
  assign \new_[60701]_  = ~A269 & A267;
  assign \new_[60702]_  = A266 & \new_[60701]_ ;
  assign \new_[60705]_  = A299 & ~A298;
  assign \new_[60708]_  = A301 & A300;
  assign \new_[60709]_  = \new_[60708]_  & \new_[60705]_ ;
  assign \new_[60710]_  = \new_[60709]_  & \new_[60702]_ ;
  assign \new_[60714]_  = ~A199 & A166;
  assign \new_[60715]_  = A167 & \new_[60714]_ ;
  assign \new_[60718]_  = A201 & A200;
  assign \new_[60721]_  = ~A265 & ~A203;
  assign \new_[60722]_  = \new_[60721]_  & \new_[60718]_ ;
  assign \new_[60723]_  = \new_[60722]_  & \new_[60715]_ ;
  assign \new_[60727]_  = ~A269 & A267;
  assign \new_[60728]_  = A266 & \new_[60727]_ ;
  assign \new_[60731]_  = A299 & ~A298;
  assign \new_[60734]_  = ~A302 & A300;
  assign \new_[60735]_  = \new_[60734]_  & \new_[60731]_ ;
  assign \new_[60736]_  = \new_[60735]_  & \new_[60728]_ ;
  assign \new_[60740]_  = ~A199 & A166;
  assign \new_[60741]_  = A167 & \new_[60740]_ ;
  assign \new_[60744]_  = A201 & A200;
  assign \new_[60747]_  = A265 & ~A203;
  assign \new_[60748]_  = \new_[60747]_  & \new_[60744]_ ;
  assign \new_[60749]_  = \new_[60748]_  & \new_[60741]_ ;
  assign \new_[60753]_  = A268 & A267;
  assign \new_[60754]_  = ~A266 & \new_[60753]_ ;
  assign \new_[60757]_  = ~A299 & A298;
  assign \new_[60760]_  = A301 & A300;
  assign \new_[60761]_  = \new_[60760]_  & \new_[60757]_ ;
  assign \new_[60762]_  = \new_[60761]_  & \new_[60754]_ ;
  assign \new_[60766]_  = ~A199 & A166;
  assign \new_[60767]_  = A167 & \new_[60766]_ ;
  assign \new_[60770]_  = A201 & A200;
  assign \new_[60773]_  = A265 & ~A203;
  assign \new_[60774]_  = \new_[60773]_  & \new_[60770]_ ;
  assign \new_[60775]_  = \new_[60774]_  & \new_[60767]_ ;
  assign \new_[60779]_  = A268 & A267;
  assign \new_[60780]_  = ~A266 & \new_[60779]_ ;
  assign \new_[60783]_  = ~A299 & A298;
  assign \new_[60786]_  = ~A302 & A300;
  assign \new_[60787]_  = \new_[60786]_  & \new_[60783]_ ;
  assign \new_[60788]_  = \new_[60787]_  & \new_[60780]_ ;
  assign \new_[60792]_  = ~A199 & A166;
  assign \new_[60793]_  = A167 & \new_[60792]_ ;
  assign \new_[60796]_  = A201 & A200;
  assign \new_[60799]_  = A265 & ~A203;
  assign \new_[60800]_  = \new_[60799]_  & \new_[60796]_ ;
  assign \new_[60801]_  = \new_[60800]_  & \new_[60793]_ ;
  assign \new_[60805]_  = A268 & A267;
  assign \new_[60806]_  = ~A266 & \new_[60805]_ ;
  assign \new_[60809]_  = A299 & ~A298;
  assign \new_[60812]_  = A301 & A300;
  assign \new_[60813]_  = \new_[60812]_  & \new_[60809]_ ;
  assign \new_[60814]_  = \new_[60813]_  & \new_[60806]_ ;
  assign \new_[60818]_  = ~A199 & A166;
  assign \new_[60819]_  = A167 & \new_[60818]_ ;
  assign \new_[60822]_  = A201 & A200;
  assign \new_[60825]_  = A265 & ~A203;
  assign \new_[60826]_  = \new_[60825]_  & \new_[60822]_ ;
  assign \new_[60827]_  = \new_[60826]_  & \new_[60819]_ ;
  assign \new_[60831]_  = A268 & A267;
  assign \new_[60832]_  = ~A266 & \new_[60831]_ ;
  assign \new_[60835]_  = A299 & ~A298;
  assign \new_[60838]_  = ~A302 & A300;
  assign \new_[60839]_  = \new_[60838]_  & \new_[60835]_ ;
  assign \new_[60840]_  = \new_[60839]_  & \new_[60832]_ ;
  assign \new_[60844]_  = ~A199 & A166;
  assign \new_[60845]_  = A167 & \new_[60844]_ ;
  assign \new_[60848]_  = A201 & A200;
  assign \new_[60851]_  = A265 & ~A203;
  assign \new_[60852]_  = \new_[60851]_  & \new_[60848]_ ;
  assign \new_[60853]_  = \new_[60852]_  & \new_[60845]_ ;
  assign \new_[60857]_  = ~A269 & A267;
  assign \new_[60858]_  = ~A266 & \new_[60857]_ ;
  assign \new_[60861]_  = ~A299 & A298;
  assign \new_[60864]_  = A301 & A300;
  assign \new_[60865]_  = \new_[60864]_  & \new_[60861]_ ;
  assign \new_[60866]_  = \new_[60865]_  & \new_[60858]_ ;
  assign \new_[60870]_  = ~A199 & A166;
  assign \new_[60871]_  = A167 & \new_[60870]_ ;
  assign \new_[60874]_  = A201 & A200;
  assign \new_[60877]_  = A265 & ~A203;
  assign \new_[60878]_  = \new_[60877]_  & \new_[60874]_ ;
  assign \new_[60879]_  = \new_[60878]_  & \new_[60871]_ ;
  assign \new_[60883]_  = ~A269 & A267;
  assign \new_[60884]_  = ~A266 & \new_[60883]_ ;
  assign \new_[60887]_  = ~A299 & A298;
  assign \new_[60890]_  = ~A302 & A300;
  assign \new_[60891]_  = \new_[60890]_  & \new_[60887]_ ;
  assign \new_[60892]_  = \new_[60891]_  & \new_[60884]_ ;
  assign \new_[60896]_  = ~A199 & A166;
  assign \new_[60897]_  = A167 & \new_[60896]_ ;
  assign \new_[60900]_  = A201 & A200;
  assign \new_[60903]_  = A265 & ~A203;
  assign \new_[60904]_  = \new_[60903]_  & \new_[60900]_ ;
  assign \new_[60905]_  = \new_[60904]_  & \new_[60897]_ ;
  assign \new_[60909]_  = ~A269 & A267;
  assign \new_[60910]_  = ~A266 & \new_[60909]_ ;
  assign \new_[60913]_  = A299 & ~A298;
  assign \new_[60916]_  = A301 & A300;
  assign \new_[60917]_  = \new_[60916]_  & \new_[60913]_ ;
  assign \new_[60918]_  = \new_[60917]_  & \new_[60910]_ ;
  assign \new_[60922]_  = ~A199 & A166;
  assign \new_[60923]_  = A167 & \new_[60922]_ ;
  assign \new_[60926]_  = A201 & A200;
  assign \new_[60929]_  = A265 & ~A203;
  assign \new_[60930]_  = \new_[60929]_  & \new_[60926]_ ;
  assign \new_[60931]_  = \new_[60930]_  & \new_[60923]_ ;
  assign \new_[60935]_  = ~A269 & A267;
  assign \new_[60936]_  = ~A266 & \new_[60935]_ ;
  assign \new_[60939]_  = A299 & ~A298;
  assign \new_[60942]_  = ~A302 & A300;
  assign \new_[60943]_  = \new_[60942]_  & \new_[60939]_ ;
  assign \new_[60944]_  = \new_[60943]_  & \new_[60936]_ ;
  assign \new_[60948]_  = A199 & A166;
  assign \new_[60949]_  = A167 & \new_[60948]_ ;
  assign \new_[60952]_  = A201 & ~A200;
  assign \new_[60955]_  = ~A265 & A202;
  assign \new_[60956]_  = \new_[60955]_  & \new_[60952]_ ;
  assign \new_[60957]_  = \new_[60956]_  & \new_[60949]_ ;
  assign \new_[60961]_  = A268 & A267;
  assign \new_[60962]_  = A266 & \new_[60961]_ ;
  assign \new_[60965]_  = ~A299 & A298;
  assign \new_[60968]_  = A301 & A300;
  assign \new_[60969]_  = \new_[60968]_  & \new_[60965]_ ;
  assign \new_[60970]_  = \new_[60969]_  & \new_[60962]_ ;
  assign \new_[60974]_  = A199 & A166;
  assign \new_[60975]_  = A167 & \new_[60974]_ ;
  assign \new_[60978]_  = A201 & ~A200;
  assign \new_[60981]_  = ~A265 & A202;
  assign \new_[60982]_  = \new_[60981]_  & \new_[60978]_ ;
  assign \new_[60983]_  = \new_[60982]_  & \new_[60975]_ ;
  assign \new_[60987]_  = A268 & A267;
  assign \new_[60988]_  = A266 & \new_[60987]_ ;
  assign \new_[60991]_  = ~A299 & A298;
  assign \new_[60994]_  = ~A302 & A300;
  assign \new_[60995]_  = \new_[60994]_  & \new_[60991]_ ;
  assign \new_[60996]_  = \new_[60995]_  & \new_[60988]_ ;
  assign \new_[61000]_  = A199 & A166;
  assign \new_[61001]_  = A167 & \new_[61000]_ ;
  assign \new_[61004]_  = A201 & ~A200;
  assign \new_[61007]_  = ~A265 & A202;
  assign \new_[61008]_  = \new_[61007]_  & \new_[61004]_ ;
  assign \new_[61009]_  = \new_[61008]_  & \new_[61001]_ ;
  assign \new_[61013]_  = A268 & A267;
  assign \new_[61014]_  = A266 & \new_[61013]_ ;
  assign \new_[61017]_  = A299 & ~A298;
  assign \new_[61020]_  = A301 & A300;
  assign \new_[61021]_  = \new_[61020]_  & \new_[61017]_ ;
  assign \new_[61022]_  = \new_[61021]_  & \new_[61014]_ ;
  assign \new_[61026]_  = A199 & A166;
  assign \new_[61027]_  = A167 & \new_[61026]_ ;
  assign \new_[61030]_  = A201 & ~A200;
  assign \new_[61033]_  = ~A265 & A202;
  assign \new_[61034]_  = \new_[61033]_  & \new_[61030]_ ;
  assign \new_[61035]_  = \new_[61034]_  & \new_[61027]_ ;
  assign \new_[61039]_  = A268 & A267;
  assign \new_[61040]_  = A266 & \new_[61039]_ ;
  assign \new_[61043]_  = A299 & ~A298;
  assign \new_[61046]_  = ~A302 & A300;
  assign \new_[61047]_  = \new_[61046]_  & \new_[61043]_ ;
  assign \new_[61048]_  = \new_[61047]_  & \new_[61040]_ ;
  assign \new_[61052]_  = A199 & A166;
  assign \new_[61053]_  = A167 & \new_[61052]_ ;
  assign \new_[61056]_  = A201 & ~A200;
  assign \new_[61059]_  = ~A265 & A202;
  assign \new_[61060]_  = \new_[61059]_  & \new_[61056]_ ;
  assign \new_[61061]_  = \new_[61060]_  & \new_[61053]_ ;
  assign \new_[61065]_  = ~A269 & A267;
  assign \new_[61066]_  = A266 & \new_[61065]_ ;
  assign \new_[61069]_  = ~A299 & A298;
  assign \new_[61072]_  = A301 & A300;
  assign \new_[61073]_  = \new_[61072]_  & \new_[61069]_ ;
  assign \new_[61074]_  = \new_[61073]_  & \new_[61066]_ ;
  assign \new_[61078]_  = A199 & A166;
  assign \new_[61079]_  = A167 & \new_[61078]_ ;
  assign \new_[61082]_  = A201 & ~A200;
  assign \new_[61085]_  = ~A265 & A202;
  assign \new_[61086]_  = \new_[61085]_  & \new_[61082]_ ;
  assign \new_[61087]_  = \new_[61086]_  & \new_[61079]_ ;
  assign \new_[61091]_  = ~A269 & A267;
  assign \new_[61092]_  = A266 & \new_[61091]_ ;
  assign \new_[61095]_  = ~A299 & A298;
  assign \new_[61098]_  = ~A302 & A300;
  assign \new_[61099]_  = \new_[61098]_  & \new_[61095]_ ;
  assign \new_[61100]_  = \new_[61099]_  & \new_[61092]_ ;
  assign \new_[61104]_  = A199 & A166;
  assign \new_[61105]_  = A167 & \new_[61104]_ ;
  assign \new_[61108]_  = A201 & ~A200;
  assign \new_[61111]_  = ~A265 & A202;
  assign \new_[61112]_  = \new_[61111]_  & \new_[61108]_ ;
  assign \new_[61113]_  = \new_[61112]_  & \new_[61105]_ ;
  assign \new_[61117]_  = ~A269 & A267;
  assign \new_[61118]_  = A266 & \new_[61117]_ ;
  assign \new_[61121]_  = A299 & ~A298;
  assign \new_[61124]_  = A301 & A300;
  assign \new_[61125]_  = \new_[61124]_  & \new_[61121]_ ;
  assign \new_[61126]_  = \new_[61125]_  & \new_[61118]_ ;
  assign \new_[61130]_  = A199 & A166;
  assign \new_[61131]_  = A167 & \new_[61130]_ ;
  assign \new_[61134]_  = A201 & ~A200;
  assign \new_[61137]_  = ~A265 & A202;
  assign \new_[61138]_  = \new_[61137]_  & \new_[61134]_ ;
  assign \new_[61139]_  = \new_[61138]_  & \new_[61131]_ ;
  assign \new_[61143]_  = ~A269 & A267;
  assign \new_[61144]_  = A266 & \new_[61143]_ ;
  assign \new_[61147]_  = A299 & ~A298;
  assign \new_[61150]_  = ~A302 & A300;
  assign \new_[61151]_  = \new_[61150]_  & \new_[61147]_ ;
  assign \new_[61152]_  = \new_[61151]_  & \new_[61144]_ ;
  assign \new_[61156]_  = A199 & A166;
  assign \new_[61157]_  = A167 & \new_[61156]_ ;
  assign \new_[61160]_  = A201 & ~A200;
  assign \new_[61163]_  = A265 & A202;
  assign \new_[61164]_  = \new_[61163]_  & \new_[61160]_ ;
  assign \new_[61165]_  = \new_[61164]_  & \new_[61157]_ ;
  assign \new_[61169]_  = A268 & A267;
  assign \new_[61170]_  = ~A266 & \new_[61169]_ ;
  assign \new_[61173]_  = ~A299 & A298;
  assign \new_[61176]_  = A301 & A300;
  assign \new_[61177]_  = \new_[61176]_  & \new_[61173]_ ;
  assign \new_[61178]_  = \new_[61177]_  & \new_[61170]_ ;
  assign \new_[61182]_  = A199 & A166;
  assign \new_[61183]_  = A167 & \new_[61182]_ ;
  assign \new_[61186]_  = A201 & ~A200;
  assign \new_[61189]_  = A265 & A202;
  assign \new_[61190]_  = \new_[61189]_  & \new_[61186]_ ;
  assign \new_[61191]_  = \new_[61190]_  & \new_[61183]_ ;
  assign \new_[61195]_  = A268 & A267;
  assign \new_[61196]_  = ~A266 & \new_[61195]_ ;
  assign \new_[61199]_  = ~A299 & A298;
  assign \new_[61202]_  = ~A302 & A300;
  assign \new_[61203]_  = \new_[61202]_  & \new_[61199]_ ;
  assign \new_[61204]_  = \new_[61203]_  & \new_[61196]_ ;
  assign \new_[61208]_  = A199 & A166;
  assign \new_[61209]_  = A167 & \new_[61208]_ ;
  assign \new_[61212]_  = A201 & ~A200;
  assign \new_[61215]_  = A265 & A202;
  assign \new_[61216]_  = \new_[61215]_  & \new_[61212]_ ;
  assign \new_[61217]_  = \new_[61216]_  & \new_[61209]_ ;
  assign \new_[61221]_  = A268 & A267;
  assign \new_[61222]_  = ~A266 & \new_[61221]_ ;
  assign \new_[61225]_  = A299 & ~A298;
  assign \new_[61228]_  = A301 & A300;
  assign \new_[61229]_  = \new_[61228]_  & \new_[61225]_ ;
  assign \new_[61230]_  = \new_[61229]_  & \new_[61222]_ ;
  assign \new_[61234]_  = A199 & A166;
  assign \new_[61235]_  = A167 & \new_[61234]_ ;
  assign \new_[61238]_  = A201 & ~A200;
  assign \new_[61241]_  = A265 & A202;
  assign \new_[61242]_  = \new_[61241]_  & \new_[61238]_ ;
  assign \new_[61243]_  = \new_[61242]_  & \new_[61235]_ ;
  assign \new_[61247]_  = A268 & A267;
  assign \new_[61248]_  = ~A266 & \new_[61247]_ ;
  assign \new_[61251]_  = A299 & ~A298;
  assign \new_[61254]_  = ~A302 & A300;
  assign \new_[61255]_  = \new_[61254]_  & \new_[61251]_ ;
  assign \new_[61256]_  = \new_[61255]_  & \new_[61248]_ ;
  assign \new_[61260]_  = A199 & A166;
  assign \new_[61261]_  = A167 & \new_[61260]_ ;
  assign \new_[61264]_  = A201 & ~A200;
  assign \new_[61267]_  = A265 & A202;
  assign \new_[61268]_  = \new_[61267]_  & \new_[61264]_ ;
  assign \new_[61269]_  = \new_[61268]_  & \new_[61261]_ ;
  assign \new_[61273]_  = ~A269 & A267;
  assign \new_[61274]_  = ~A266 & \new_[61273]_ ;
  assign \new_[61277]_  = ~A299 & A298;
  assign \new_[61280]_  = A301 & A300;
  assign \new_[61281]_  = \new_[61280]_  & \new_[61277]_ ;
  assign \new_[61282]_  = \new_[61281]_  & \new_[61274]_ ;
  assign \new_[61286]_  = A199 & A166;
  assign \new_[61287]_  = A167 & \new_[61286]_ ;
  assign \new_[61290]_  = A201 & ~A200;
  assign \new_[61293]_  = A265 & A202;
  assign \new_[61294]_  = \new_[61293]_  & \new_[61290]_ ;
  assign \new_[61295]_  = \new_[61294]_  & \new_[61287]_ ;
  assign \new_[61299]_  = ~A269 & A267;
  assign \new_[61300]_  = ~A266 & \new_[61299]_ ;
  assign \new_[61303]_  = ~A299 & A298;
  assign \new_[61306]_  = ~A302 & A300;
  assign \new_[61307]_  = \new_[61306]_  & \new_[61303]_ ;
  assign \new_[61308]_  = \new_[61307]_  & \new_[61300]_ ;
  assign \new_[61312]_  = A199 & A166;
  assign \new_[61313]_  = A167 & \new_[61312]_ ;
  assign \new_[61316]_  = A201 & ~A200;
  assign \new_[61319]_  = A265 & A202;
  assign \new_[61320]_  = \new_[61319]_  & \new_[61316]_ ;
  assign \new_[61321]_  = \new_[61320]_  & \new_[61313]_ ;
  assign \new_[61325]_  = ~A269 & A267;
  assign \new_[61326]_  = ~A266 & \new_[61325]_ ;
  assign \new_[61329]_  = A299 & ~A298;
  assign \new_[61332]_  = A301 & A300;
  assign \new_[61333]_  = \new_[61332]_  & \new_[61329]_ ;
  assign \new_[61334]_  = \new_[61333]_  & \new_[61326]_ ;
  assign \new_[61338]_  = A199 & A166;
  assign \new_[61339]_  = A167 & \new_[61338]_ ;
  assign \new_[61342]_  = A201 & ~A200;
  assign \new_[61345]_  = A265 & A202;
  assign \new_[61346]_  = \new_[61345]_  & \new_[61342]_ ;
  assign \new_[61347]_  = \new_[61346]_  & \new_[61339]_ ;
  assign \new_[61351]_  = ~A269 & A267;
  assign \new_[61352]_  = ~A266 & \new_[61351]_ ;
  assign \new_[61355]_  = A299 & ~A298;
  assign \new_[61358]_  = ~A302 & A300;
  assign \new_[61359]_  = \new_[61358]_  & \new_[61355]_ ;
  assign \new_[61360]_  = \new_[61359]_  & \new_[61352]_ ;
  assign \new_[61364]_  = A199 & A166;
  assign \new_[61365]_  = A167 & \new_[61364]_ ;
  assign \new_[61368]_  = A201 & ~A200;
  assign \new_[61371]_  = ~A265 & ~A203;
  assign \new_[61372]_  = \new_[61371]_  & \new_[61368]_ ;
  assign \new_[61373]_  = \new_[61372]_  & \new_[61365]_ ;
  assign \new_[61377]_  = A268 & A267;
  assign \new_[61378]_  = A266 & \new_[61377]_ ;
  assign \new_[61381]_  = ~A299 & A298;
  assign \new_[61384]_  = A301 & A300;
  assign \new_[61385]_  = \new_[61384]_  & \new_[61381]_ ;
  assign \new_[61386]_  = \new_[61385]_  & \new_[61378]_ ;
  assign \new_[61390]_  = A199 & A166;
  assign \new_[61391]_  = A167 & \new_[61390]_ ;
  assign \new_[61394]_  = A201 & ~A200;
  assign \new_[61397]_  = ~A265 & ~A203;
  assign \new_[61398]_  = \new_[61397]_  & \new_[61394]_ ;
  assign \new_[61399]_  = \new_[61398]_  & \new_[61391]_ ;
  assign \new_[61403]_  = A268 & A267;
  assign \new_[61404]_  = A266 & \new_[61403]_ ;
  assign \new_[61407]_  = ~A299 & A298;
  assign \new_[61410]_  = ~A302 & A300;
  assign \new_[61411]_  = \new_[61410]_  & \new_[61407]_ ;
  assign \new_[61412]_  = \new_[61411]_  & \new_[61404]_ ;
  assign \new_[61416]_  = A199 & A166;
  assign \new_[61417]_  = A167 & \new_[61416]_ ;
  assign \new_[61420]_  = A201 & ~A200;
  assign \new_[61423]_  = ~A265 & ~A203;
  assign \new_[61424]_  = \new_[61423]_  & \new_[61420]_ ;
  assign \new_[61425]_  = \new_[61424]_  & \new_[61417]_ ;
  assign \new_[61429]_  = A268 & A267;
  assign \new_[61430]_  = A266 & \new_[61429]_ ;
  assign \new_[61433]_  = A299 & ~A298;
  assign \new_[61436]_  = A301 & A300;
  assign \new_[61437]_  = \new_[61436]_  & \new_[61433]_ ;
  assign \new_[61438]_  = \new_[61437]_  & \new_[61430]_ ;
  assign \new_[61442]_  = A199 & A166;
  assign \new_[61443]_  = A167 & \new_[61442]_ ;
  assign \new_[61446]_  = A201 & ~A200;
  assign \new_[61449]_  = ~A265 & ~A203;
  assign \new_[61450]_  = \new_[61449]_  & \new_[61446]_ ;
  assign \new_[61451]_  = \new_[61450]_  & \new_[61443]_ ;
  assign \new_[61455]_  = A268 & A267;
  assign \new_[61456]_  = A266 & \new_[61455]_ ;
  assign \new_[61459]_  = A299 & ~A298;
  assign \new_[61462]_  = ~A302 & A300;
  assign \new_[61463]_  = \new_[61462]_  & \new_[61459]_ ;
  assign \new_[61464]_  = \new_[61463]_  & \new_[61456]_ ;
  assign \new_[61468]_  = A199 & A166;
  assign \new_[61469]_  = A167 & \new_[61468]_ ;
  assign \new_[61472]_  = A201 & ~A200;
  assign \new_[61475]_  = ~A265 & ~A203;
  assign \new_[61476]_  = \new_[61475]_  & \new_[61472]_ ;
  assign \new_[61477]_  = \new_[61476]_  & \new_[61469]_ ;
  assign \new_[61481]_  = ~A269 & A267;
  assign \new_[61482]_  = A266 & \new_[61481]_ ;
  assign \new_[61485]_  = ~A299 & A298;
  assign \new_[61488]_  = A301 & A300;
  assign \new_[61489]_  = \new_[61488]_  & \new_[61485]_ ;
  assign \new_[61490]_  = \new_[61489]_  & \new_[61482]_ ;
  assign \new_[61494]_  = A199 & A166;
  assign \new_[61495]_  = A167 & \new_[61494]_ ;
  assign \new_[61498]_  = A201 & ~A200;
  assign \new_[61501]_  = ~A265 & ~A203;
  assign \new_[61502]_  = \new_[61501]_  & \new_[61498]_ ;
  assign \new_[61503]_  = \new_[61502]_  & \new_[61495]_ ;
  assign \new_[61507]_  = ~A269 & A267;
  assign \new_[61508]_  = A266 & \new_[61507]_ ;
  assign \new_[61511]_  = ~A299 & A298;
  assign \new_[61514]_  = ~A302 & A300;
  assign \new_[61515]_  = \new_[61514]_  & \new_[61511]_ ;
  assign \new_[61516]_  = \new_[61515]_  & \new_[61508]_ ;
  assign \new_[61520]_  = A199 & A166;
  assign \new_[61521]_  = A167 & \new_[61520]_ ;
  assign \new_[61524]_  = A201 & ~A200;
  assign \new_[61527]_  = ~A265 & ~A203;
  assign \new_[61528]_  = \new_[61527]_  & \new_[61524]_ ;
  assign \new_[61529]_  = \new_[61528]_  & \new_[61521]_ ;
  assign \new_[61533]_  = ~A269 & A267;
  assign \new_[61534]_  = A266 & \new_[61533]_ ;
  assign \new_[61537]_  = A299 & ~A298;
  assign \new_[61540]_  = A301 & A300;
  assign \new_[61541]_  = \new_[61540]_  & \new_[61537]_ ;
  assign \new_[61542]_  = \new_[61541]_  & \new_[61534]_ ;
  assign \new_[61546]_  = A199 & A166;
  assign \new_[61547]_  = A167 & \new_[61546]_ ;
  assign \new_[61550]_  = A201 & ~A200;
  assign \new_[61553]_  = ~A265 & ~A203;
  assign \new_[61554]_  = \new_[61553]_  & \new_[61550]_ ;
  assign \new_[61555]_  = \new_[61554]_  & \new_[61547]_ ;
  assign \new_[61559]_  = ~A269 & A267;
  assign \new_[61560]_  = A266 & \new_[61559]_ ;
  assign \new_[61563]_  = A299 & ~A298;
  assign \new_[61566]_  = ~A302 & A300;
  assign \new_[61567]_  = \new_[61566]_  & \new_[61563]_ ;
  assign \new_[61568]_  = \new_[61567]_  & \new_[61560]_ ;
  assign \new_[61572]_  = A199 & A166;
  assign \new_[61573]_  = A167 & \new_[61572]_ ;
  assign \new_[61576]_  = A201 & ~A200;
  assign \new_[61579]_  = A265 & ~A203;
  assign \new_[61580]_  = \new_[61579]_  & \new_[61576]_ ;
  assign \new_[61581]_  = \new_[61580]_  & \new_[61573]_ ;
  assign \new_[61585]_  = A268 & A267;
  assign \new_[61586]_  = ~A266 & \new_[61585]_ ;
  assign \new_[61589]_  = ~A299 & A298;
  assign \new_[61592]_  = A301 & A300;
  assign \new_[61593]_  = \new_[61592]_  & \new_[61589]_ ;
  assign \new_[61594]_  = \new_[61593]_  & \new_[61586]_ ;
  assign \new_[61598]_  = A199 & A166;
  assign \new_[61599]_  = A167 & \new_[61598]_ ;
  assign \new_[61602]_  = A201 & ~A200;
  assign \new_[61605]_  = A265 & ~A203;
  assign \new_[61606]_  = \new_[61605]_  & \new_[61602]_ ;
  assign \new_[61607]_  = \new_[61606]_  & \new_[61599]_ ;
  assign \new_[61611]_  = A268 & A267;
  assign \new_[61612]_  = ~A266 & \new_[61611]_ ;
  assign \new_[61615]_  = ~A299 & A298;
  assign \new_[61618]_  = ~A302 & A300;
  assign \new_[61619]_  = \new_[61618]_  & \new_[61615]_ ;
  assign \new_[61620]_  = \new_[61619]_  & \new_[61612]_ ;
  assign \new_[61624]_  = A199 & A166;
  assign \new_[61625]_  = A167 & \new_[61624]_ ;
  assign \new_[61628]_  = A201 & ~A200;
  assign \new_[61631]_  = A265 & ~A203;
  assign \new_[61632]_  = \new_[61631]_  & \new_[61628]_ ;
  assign \new_[61633]_  = \new_[61632]_  & \new_[61625]_ ;
  assign \new_[61637]_  = A268 & A267;
  assign \new_[61638]_  = ~A266 & \new_[61637]_ ;
  assign \new_[61641]_  = A299 & ~A298;
  assign \new_[61644]_  = A301 & A300;
  assign \new_[61645]_  = \new_[61644]_  & \new_[61641]_ ;
  assign \new_[61646]_  = \new_[61645]_  & \new_[61638]_ ;
  assign \new_[61650]_  = A199 & A166;
  assign \new_[61651]_  = A167 & \new_[61650]_ ;
  assign \new_[61654]_  = A201 & ~A200;
  assign \new_[61657]_  = A265 & ~A203;
  assign \new_[61658]_  = \new_[61657]_  & \new_[61654]_ ;
  assign \new_[61659]_  = \new_[61658]_  & \new_[61651]_ ;
  assign \new_[61663]_  = A268 & A267;
  assign \new_[61664]_  = ~A266 & \new_[61663]_ ;
  assign \new_[61667]_  = A299 & ~A298;
  assign \new_[61670]_  = ~A302 & A300;
  assign \new_[61671]_  = \new_[61670]_  & \new_[61667]_ ;
  assign \new_[61672]_  = \new_[61671]_  & \new_[61664]_ ;
  assign \new_[61676]_  = A199 & A166;
  assign \new_[61677]_  = A167 & \new_[61676]_ ;
  assign \new_[61680]_  = A201 & ~A200;
  assign \new_[61683]_  = A265 & ~A203;
  assign \new_[61684]_  = \new_[61683]_  & \new_[61680]_ ;
  assign \new_[61685]_  = \new_[61684]_  & \new_[61677]_ ;
  assign \new_[61689]_  = ~A269 & A267;
  assign \new_[61690]_  = ~A266 & \new_[61689]_ ;
  assign \new_[61693]_  = ~A299 & A298;
  assign \new_[61696]_  = A301 & A300;
  assign \new_[61697]_  = \new_[61696]_  & \new_[61693]_ ;
  assign \new_[61698]_  = \new_[61697]_  & \new_[61690]_ ;
  assign \new_[61702]_  = A199 & A166;
  assign \new_[61703]_  = A167 & \new_[61702]_ ;
  assign \new_[61706]_  = A201 & ~A200;
  assign \new_[61709]_  = A265 & ~A203;
  assign \new_[61710]_  = \new_[61709]_  & \new_[61706]_ ;
  assign \new_[61711]_  = \new_[61710]_  & \new_[61703]_ ;
  assign \new_[61715]_  = ~A269 & A267;
  assign \new_[61716]_  = ~A266 & \new_[61715]_ ;
  assign \new_[61719]_  = ~A299 & A298;
  assign \new_[61722]_  = ~A302 & A300;
  assign \new_[61723]_  = \new_[61722]_  & \new_[61719]_ ;
  assign \new_[61724]_  = \new_[61723]_  & \new_[61716]_ ;
  assign \new_[61728]_  = A199 & A166;
  assign \new_[61729]_  = A167 & \new_[61728]_ ;
  assign \new_[61732]_  = A201 & ~A200;
  assign \new_[61735]_  = A265 & ~A203;
  assign \new_[61736]_  = \new_[61735]_  & \new_[61732]_ ;
  assign \new_[61737]_  = \new_[61736]_  & \new_[61729]_ ;
  assign \new_[61741]_  = ~A269 & A267;
  assign \new_[61742]_  = ~A266 & \new_[61741]_ ;
  assign \new_[61745]_  = A299 & ~A298;
  assign \new_[61748]_  = A301 & A300;
  assign \new_[61749]_  = \new_[61748]_  & \new_[61745]_ ;
  assign \new_[61750]_  = \new_[61749]_  & \new_[61742]_ ;
  assign \new_[61754]_  = A199 & A166;
  assign \new_[61755]_  = A167 & \new_[61754]_ ;
  assign \new_[61758]_  = A201 & ~A200;
  assign \new_[61761]_  = A265 & ~A203;
  assign \new_[61762]_  = \new_[61761]_  & \new_[61758]_ ;
  assign \new_[61763]_  = \new_[61762]_  & \new_[61755]_ ;
  assign \new_[61767]_  = ~A269 & A267;
  assign \new_[61768]_  = ~A266 & \new_[61767]_ ;
  assign \new_[61771]_  = A299 & ~A298;
  assign \new_[61774]_  = ~A302 & A300;
  assign \new_[61775]_  = \new_[61774]_  & \new_[61771]_ ;
  assign \new_[61776]_  = \new_[61775]_  & \new_[61768]_ ;
  assign \new_[61780]_  = ~A199 & ~A166;
  assign \new_[61781]_  = ~A167 & \new_[61780]_ ;
  assign \new_[61784]_  = A201 & A200;
  assign \new_[61787]_  = ~A265 & A202;
  assign \new_[61788]_  = \new_[61787]_  & \new_[61784]_ ;
  assign \new_[61789]_  = \new_[61788]_  & \new_[61781]_ ;
  assign \new_[61793]_  = A268 & A267;
  assign \new_[61794]_  = A266 & \new_[61793]_ ;
  assign \new_[61797]_  = ~A299 & A298;
  assign \new_[61800]_  = A301 & A300;
  assign \new_[61801]_  = \new_[61800]_  & \new_[61797]_ ;
  assign \new_[61802]_  = \new_[61801]_  & \new_[61794]_ ;
  assign \new_[61806]_  = ~A199 & ~A166;
  assign \new_[61807]_  = ~A167 & \new_[61806]_ ;
  assign \new_[61810]_  = A201 & A200;
  assign \new_[61813]_  = ~A265 & A202;
  assign \new_[61814]_  = \new_[61813]_  & \new_[61810]_ ;
  assign \new_[61815]_  = \new_[61814]_  & \new_[61807]_ ;
  assign \new_[61819]_  = A268 & A267;
  assign \new_[61820]_  = A266 & \new_[61819]_ ;
  assign \new_[61823]_  = ~A299 & A298;
  assign \new_[61826]_  = ~A302 & A300;
  assign \new_[61827]_  = \new_[61826]_  & \new_[61823]_ ;
  assign \new_[61828]_  = \new_[61827]_  & \new_[61820]_ ;
  assign \new_[61832]_  = ~A199 & ~A166;
  assign \new_[61833]_  = ~A167 & \new_[61832]_ ;
  assign \new_[61836]_  = A201 & A200;
  assign \new_[61839]_  = ~A265 & A202;
  assign \new_[61840]_  = \new_[61839]_  & \new_[61836]_ ;
  assign \new_[61841]_  = \new_[61840]_  & \new_[61833]_ ;
  assign \new_[61845]_  = A268 & A267;
  assign \new_[61846]_  = A266 & \new_[61845]_ ;
  assign \new_[61849]_  = A299 & ~A298;
  assign \new_[61852]_  = A301 & A300;
  assign \new_[61853]_  = \new_[61852]_  & \new_[61849]_ ;
  assign \new_[61854]_  = \new_[61853]_  & \new_[61846]_ ;
  assign \new_[61858]_  = ~A199 & ~A166;
  assign \new_[61859]_  = ~A167 & \new_[61858]_ ;
  assign \new_[61862]_  = A201 & A200;
  assign \new_[61865]_  = ~A265 & A202;
  assign \new_[61866]_  = \new_[61865]_  & \new_[61862]_ ;
  assign \new_[61867]_  = \new_[61866]_  & \new_[61859]_ ;
  assign \new_[61871]_  = A268 & A267;
  assign \new_[61872]_  = A266 & \new_[61871]_ ;
  assign \new_[61875]_  = A299 & ~A298;
  assign \new_[61878]_  = ~A302 & A300;
  assign \new_[61879]_  = \new_[61878]_  & \new_[61875]_ ;
  assign \new_[61880]_  = \new_[61879]_  & \new_[61872]_ ;
  assign \new_[61884]_  = ~A199 & ~A166;
  assign \new_[61885]_  = ~A167 & \new_[61884]_ ;
  assign \new_[61888]_  = A201 & A200;
  assign \new_[61891]_  = ~A265 & A202;
  assign \new_[61892]_  = \new_[61891]_  & \new_[61888]_ ;
  assign \new_[61893]_  = \new_[61892]_  & \new_[61885]_ ;
  assign \new_[61897]_  = ~A269 & A267;
  assign \new_[61898]_  = A266 & \new_[61897]_ ;
  assign \new_[61901]_  = ~A299 & A298;
  assign \new_[61904]_  = A301 & A300;
  assign \new_[61905]_  = \new_[61904]_  & \new_[61901]_ ;
  assign \new_[61906]_  = \new_[61905]_  & \new_[61898]_ ;
  assign \new_[61910]_  = ~A199 & ~A166;
  assign \new_[61911]_  = ~A167 & \new_[61910]_ ;
  assign \new_[61914]_  = A201 & A200;
  assign \new_[61917]_  = ~A265 & A202;
  assign \new_[61918]_  = \new_[61917]_  & \new_[61914]_ ;
  assign \new_[61919]_  = \new_[61918]_  & \new_[61911]_ ;
  assign \new_[61923]_  = ~A269 & A267;
  assign \new_[61924]_  = A266 & \new_[61923]_ ;
  assign \new_[61927]_  = ~A299 & A298;
  assign \new_[61930]_  = ~A302 & A300;
  assign \new_[61931]_  = \new_[61930]_  & \new_[61927]_ ;
  assign \new_[61932]_  = \new_[61931]_  & \new_[61924]_ ;
  assign \new_[61936]_  = ~A199 & ~A166;
  assign \new_[61937]_  = ~A167 & \new_[61936]_ ;
  assign \new_[61940]_  = A201 & A200;
  assign \new_[61943]_  = ~A265 & A202;
  assign \new_[61944]_  = \new_[61943]_  & \new_[61940]_ ;
  assign \new_[61945]_  = \new_[61944]_  & \new_[61937]_ ;
  assign \new_[61949]_  = ~A269 & A267;
  assign \new_[61950]_  = A266 & \new_[61949]_ ;
  assign \new_[61953]_  = A299 & ~A298;
  assign \new_[61956]_  = A301 & A300;
  assign \new_[61957]_  = \new_[61956]_  & \new_[61953]_ ;
  assign \new_[61958]_  = \new_[61957]_  & \new_[61950]_ ;
  assign \new_[61962]_  = ~A199 & ~A166;
  assign \new_[61963]_  = ~A167 & \new_[61962]_ ;
  assign \new_[61966]_  = A201 & A200;
  assign \new_[61969]_  = ~A265 & A202;
  assign \new_[61970]_  = \new_[61969]_  & \new_[61966]_ ;
  assign \new_[61971]_  = \new_[61970]_  & \new_[61963]_ ;
  assign \new_[61975]_  = ~A269 & A267;
  assign \new_[61976]_  = A266 & \new_[61975]_ ;
  assign \new_[61979]_  = A299 & ~A298;
  assign \new_[61982]_  = ~A302 & A300;
  assign \new_[61983]_  = \new_[61982]_  & \new_[61979]_ ;
  assign \new_[61984]_  = \new_[61983]_  & \new_[61976]_ ;
  assign \new_[61988]_  = ~A199 & ~A166;
  assign \new_[61989]_  = ~A167 & \new_[61988]_ ;
  assign \new_[61992]_  = A201 & A200;
  assign \new_[61995]_  = A265 & A202;
  assign \new_[61996]_  = \new_[61995]_  & \new_[61992]_ ;
  assign \new_[61997]_  = \new_[61996]_  & \new_[61989]_ ;
  assign \new_[62001]_  = A268 & A267;
  assign \new_[62002]_  = ~A266 & \new_[62001]_ ;
  assign \new_[62005]_  = ~A299 & A298;
  assign \new_[62008]_  = A301 & A300;
  assign \new_[62009]_  = \new_[62008]_  & \new_[62005]_ ;
  assign \new_[62010]_  = \new_[62009]_  & \new_[62002]_ ;
  assign \new_[62014]_  = ~A199 & ~A166;
  assign \new_[62015]_  = ~A167 & \new_[62014]_ ;
  assign \new_[62018]_  = A201 & A200;
  assign \new_[62021]_  = A265 & A202;
  assign \new_[62022]_  = \new_[62021]_  & \new_[62018]_ ;
  assign \new_[62023]_  = \new_[62022]_  & \new_[62015]_ ;
  assign \new_[62027]_  = A268 & A267;
  assign \new_[62028]_  = ~A266 & \new_[62027]_ ;
  assign \new_[62031]_  = ~A299 & A298;
  assign \new_[62034]_  = ~A302 & A300;
  assign \new_[62035]_  = \new_[62034]_  & \new_[62031]_ ;
  assign \new_[62036]_  = \new_[62035]_  & \new_[62028]_ ;
  assign \new_[62040]_  = ~A199 & ~A166;
  assign \new_[62041]_  = ~A167 & \new_[62040]_ ;
  assign \new_[62044]_  = A201 & A200;
  assign \new_[62047]_  = A265 & A202;
  assign \new_[62048]_  = \new_[62047]_  & \new_[62044]_ ;
  assign \new_[62049]_  = \new_[62048]_  & \new_[62041]_ ;
  assign \new_[62053]_  = A268 & A267;
  assign \new_[62054]_  = ~A266 & \new_[62053]_ ;
  assign \new_[62057]_  = A299 & ~A298;
  assign \new_[62060]_  = A301 & A300;
  assign \new_[62061]_  = \new_[62060]_  & \new_[62057]_ ;
  assign \new_[62062]_  = \new_[62061]_  & \new_[62054]_ ;
  assign \new_[62066]_  = ~A199 & ~A166;
  assign \new_[62067]_  = ~A167 & \new_[62066]_ ;
  assign \new_[62070]_  = A201 & A200;
  assign \new_[62073]_  = A265 & A202;
  assign \new_[62074]_  = \new_[62073]_  & \new_[62070]_ ;
  assign \new_[62075]_  = \new_[62074]_  & \new_[62067]_ ;
  assign \new_[62079]_  = A268 & A267;
  assign \new_[62080]_  = ~A266 & \new_[62079]_ ;
  assign \new_[62083]_  = A299 & ~A298;
  assign \new_[62086]_  = ~A302 & A300;
  assign \new_[62087]_  = \new_[62086]_  & \new_[62083]_ ;
  assign \new_[62088]_  = \new_[62087]_  & \new_[62080]_ ;
  assign \new_[62092]_  = ~A199 & ~A166;
  assign \new_[62093]_  = ~A167 & \new_[62092]_ ;
  assign \new_[62096]_  = A201 & A200;
  assign \new_[62099]_  = A265 & A202;
  assign \new_[62100]_  = \new_[62099]_  & \new_[62096]_ ;
  assign \new_[62101]_  = \new_[62100]_  & \new_[62093]_ ;
  assign \new_[62105]_  = ~A269 & A267;
  assign \new_[62106]_  = ~A266 & \new_[62105]_ ;
  assign \new_[62109]_  = ~A299 & A298;
  assign \new_[62112]_  = A301 & A300;
  assign \new_[62113]_  = \new_[62112]_  & \new_[62109]_ ;
  assign \new_[62114]_  = \new_[62113]_  & \new_[62106]_ ;
  assign \new_[62118]_  = ~A199 & ~A166;
  assign \new_[62119]_  = ~A167 & \new_[62118]_ ;
  assign \new_[62122]_  = A201 & A200;
  assign \new_[62125]_  = A265 & A202;
  assign \new_[62126]_  = \new_[62125]_  & \new_[62122]_ ;
  assign \new_[62127]_  = \new_[62126]_  & \new_[62119]_ ;
  assign \new_[62131]_  = ~A269 & A267;
  assign \new_[62132]_  = ~A266 & \new_[62131]_ ;
  assign \new_[62135]_  = ~A299 & A298;
  assign \new_[62138]_  = ~A302 & A300;
  assign \new_[62139]_  = \new_[62138]_  & \new_[62135]_ ;
  assign \new_[62140]_  = \new_[62139]_  & \new_[62132]_ ;
  assign \new_[62144]_  = ~A199 & ~A166;
  assign \new_[62145]_  = ~A167 & \new_[62144]_ ;
  assign \new_[62148]_  = A201 & A200;
  assign \new_[62151]_  = A265 & A202;
  assign \new_[62152]_  = \new_[62151]_  & \new_[62148]_ ;
  assign \new_[62153]_  = \new_[62152]_  & \new_[62145]_ ;
  assign \new_[62157]_  = ~A269 & A267;
  assign \new_[62158]_  = ~A266 & \new_[62157]_ ;
  assign \new_[62161]_  = A299 & ~A298;
  assign \new_[62164]_  = A301 & A300;
  assign \new_[62165]_  = \new_[62164]_  & \new_[62161]_ ;
  assign \new_[62166]_  = \new_[62165]_  & \new_[62158]_ ;
  assign \new_[62170]_  = ~A199 & ~A166;
  assign \new_[62171]_  = ~A167 & \new_[62170]_ ;
  assign \new_[62174]_  = A201 & A200;
  assign \new_[62177]_  = A265 & A202;
  assign \new_[62178]_  = \new_[62177]_  & \new_[62174]_ ;
  assign \new_[62179]_  = \new_[62178]_  & \new_[62171]_ ;
  assign \new_[62183]_  = ~A269 & A267;
  assign \new_[62184]_  = ~A266 & \new_[62183]_ ;
  assign \new_[62187]_  = A299 & ~A298;
  assign \new_[62190]_  = ~A302 & A300;
  assign \new_[62191]_  = \new_[62190]_  & \new_[62187]_ ;
  assign \new_[62192]_  = \new_[62191]_  & \new_[62184]_ ;
  assign \new_[62196]_  = ~A199 & ~A166;
  assign \new_[62197]_  = ~A167 & \new_[62196]_ ;
  assign \new_[62200]_  = A201 & A200;
  assign \new_[62203]_  = ~A265 & ~A203;
  assign \new_[62204]_  = \new_[62203]_  & \new_[62200]_ ;
  assign \new_[62205]_  = \new_[62204]_  & \new_[62197]_ ;
  assign \new_[62209]_  = A268 & A267;
  assign \new_[62210]_  = A266 & \new_[62209]_ ;
  assign \new_[62213]_  = ~A299 & A298;
  assign \new_[62216]_  = A301 & A300;
  assign \new_[62217]_  = \new_[62216]_  & \new_[62213]_ ;
  assign \new_[62218]_  = \new_[62217]_  & \new_[62210]_ ;
  assign \new_[62222]_  = ~A199 & ~A166;
  assign \new_[62223]_  = ~A167 & \new_[62222]_ ;
  assign \new_[62226]_  = A201 & A200;
  assign \new_[62229]_  = ~A265 & ~A203;
  assign \new_[62230]_  = \new_[62229]_  & \new_[62226]_ ;
  assign \new_[62231]_  = \new_[62230]_  & \new_[62223]_ ;
  assign \new_[62235]_  = A268 & A267;
  assign \new_[62236]_  = A266 & \new_[62235]_ ;
  assign \new_[62239]_  = ~A299 & A298;
  assign \new_[62242]_  = ~A302 & A300;
  assign \new_[62243]_  = \new_[62242]_  & \new_[62239]_ ;
  assign \new_[62244]_  = \new_[62243]_  & \new_[62236]_ ;
  assign \new_[62248]_  = ~A199 & ~A166;
  assign \new_[62249]_  = ~A167 & \new_[62248]_ ;
  assign \new_[62252]_  = A201 & A200;
  assign \new_[62255]_  = ~A265 & ~A203;
  assign \new_[62256]_  = \new_[62255]_  & \new_[62252]_ ;
  assign \new_[62257]_  = \new_[62256]_  & \new_[62249]_ ;
  assign \new_[62261]_  = A268 & A267;
  assign \new_[62262]_  = A266 & \new_[62261]_ ;
  assign \new_[62265]_  = A299 & ~A298;
  assign \new_[62268]_  = A301 & A300;
  assign \new_[62269]_  = \new_[62268]_  & \new_[62265]_ ;
  assign \new_[62270]_  = \new_[62269]_  & \new_[62262]_ ;
  assign \new_[62274]_  = ~A199 & ~A166;
  assign \new_[62275]_  = ~A167 & \new_[62274]_ ;
  assign \new_[62278]_  = A201 & A200;
  assign \new_[62281]_  = ~A265 & ~A203;
  assign \new_[62282]_  = \new_[62281]_  & \new_[62278]_ ;
  assign \new_[62283]_  = \new_[62282]_  & \new_[62275]_ ;
  assign \new_[62287]_  = A268 & A267;
  assign \new_[62288]_  = A266 & \new_[62287]_ ;
  assign \new_[62291]_  = A299 & ~A298;
  assign \new_[62294]_  = ~A302 & A300;
  assign \new_[62295]_  = \new_[62294]_  & \new_[62291]_ ;
  assign \new_[62296]_  = \new_[62295]_  & \new_[62288]_ ;
  assign \new_[62300]_  = ~A199 & ~A166;
  assign \new_[62301]_  = ~A167 & \new_[62300]_ ;
  assign \new_[62304]_  = A201 & A200;
  assign \new_[62307]_  = ~A265 & ~A203;
  assign \new_[62308]_  = \new_[62307]_  & \new_[62304]_ ;
  assign \new_[62309]_  = \new_[62308]_  & \new_[62301]_ ;
  assign \new_[62313]_  = ~A269 & A267;
  assign \new_[62314]_  = A266 & \new_[62313]_ ;
  assign \new_[62317]_  = ~A299 & A298;
  assign \new_[62320]_  = A301 & A300;
  assign \new_[62321]_  = \new_[62320]_  & \new_[62317]_ ;
  assign \new_[62322]_  = \new_[62321]_  & \new_[62314]_ ;
  assign \new_[62326]_  = ~A199 & ~A166;
  assign \new_[62327]_  = ~A167 & \new_[62326]_ ;
  assign \new_[62330]_  = A201 & A200;
  assign \new_[62333]_  = ~A265 & ~A203;
  assign \new_[62334]_  = \new_[62333]_  & \new_[62330]_ ;
  assign \new_[62335]_  = \new_[62334]_  & \new_[62327]_ ;
  assign \new_[62339]_  = ~A269 & A267;
  assign \new_[62340]_  = A266 & \new_[62339]_ ;
  assign \new_[62343]_  = ~A299 & A298;
  assign \new_[62346]_  = ~A302 & A300;
  assign \new_[62347]_  = \new_[62346]_  & \new_[62343]_ ;
  assign \new_[62348]_  = \new_[62347]_  & \new_[62340]_ ;
  assign \new_[62352]_  = ~A199 & ~A166;
  assign \new_[62353]_  = ~A167 & \new_[62352]_ ;
  assign \new_[62356]_  = A201 & A200;
  assign \new_[62359]_  = ~A265 & ~A203;
  assign \new_[62360]_  = \new_[62359]_  & \new_[62356]_ ;
  assign \new_[62361]_  = \new_[62360]_  & \new_[62353]_ ;
  assign \new_[62365]_  = ~A269 & A267;
  assign \new_[62366]_  = A266 & \new_[62365]_ ;
  assign \new_[62369]_  = A299 & ~A298;
  assign \new_[62372]_  = A301 & A300;
  assign \new_[62373]_  = \new_[62372]_  & \new_[62369]_ ;
  assign \new_[62374]_  = \new_[62373]_  & \new_[62366]_ ;
  assign \new_[62378]_  = ~A199 & ~A166;
  assign \new_[62379]_  = ~A167 & \new_[62378]_ ;
  assign \new_[62382]_  = A201 & A200;
  assign \new_[62385]_  = ~A265 & ~A203;
  assign \new_[62386]_  = \new_[62385]_  & \new_[62382]_ ;
  assign \new_[62387]_  = \new_[62386]_  & \new_[62379]_ ;
  assign \new_[62391]_  = ~A269 & A267;
  assign \new_[62392]_  = A266 & \new_[62391]_ ;
  assign \new_[62395]_  = A299 & ~A298;
  assign \new_[62398]_  = ~A302 & A300;
  assign \new_[62399]_  = \new_[62398]_  & \new_[62395]_ ;
  assign \new_[62400]_  = \new_[62399]_  & \new_[62392]_ ;
  assign \new_[62404]_  = ~A199 & ~A166;
  assign \new_[62405]_  = ~A167 & \new_[62404]_ ;
  assign \new_[62408]_  = A201 & A200;
  assign \new_[62411]_  = A265 & ~A203;
  assign \new_[62412]_  = \new_[62411]_  & \new_[62408]_ ;
  assign \new_[62413]_  = \new_[62412]_  & \new_[62405]_ ;
  assign \new_[62417]_  = A268 & A267;
  assign \new_[62418]_  = ~A266 & \new_[62417]_ ;
  assign \new_[62421]_  = ~A299 & A298;
  assign \new_[62424]_  = A301 & A300;
  assign \new_[62425]_  = \new_[62424]_  & \new_[62421]_ ;
  assign \new_[62426]_  = \new_[62425]_  & \new_[62418]_ ;
  assign \new_[62430]_  = ~A199 & ~A166;
  assign \new_[62431]_  = ~A167 & \new_[62430]_ ;
  assign \new_[62434]_  = A201 & A200;
  assign \new_[62437]_  = A265 & ~A203;
  assign \new_[62438]_  = \new_[62437]_  & \new_[62434]_ ;
  assign \new_[62439]_  = \new_[62438]_  & \new_[62431]_ ;
  assign \new_[62443]_  = A268 & A267;
  assign \new_[62444]_  = ~A266 & \new_[62443]_ ;
  assign \new_[62447]_  = ~A299 & A298;
  assign \new_[62450]_  = ~A302 & A300;
  assign \new_[62451]_  = \new_[62450]_  & \new_[62447]_ ;
  assign \new_[62452]_  = \new_[62451]_  & \new_[62444]_ ;
  assign \new_[62456]_  = ~A199 & ~A166;
  assign \new_[62457]_  = ~A167 & \new_[62456]_ ;
  assign \new_[62460]_  = A201 & A200;
  assign \new_[62463]_  = A265 & ~A203;
  assign \new_[62464]_  = \new_[62463]_  & \new_[62460]_ ;
  assign \new_[62465]_  = \new_[62464]_  & \new_[62457]_ ;
  assign \new_[62469]_  = A268 & A267;
  assign \new_[62470]_  = ~A266 & \new_[62469]_ ;
  assign \new_[62473]_  = A299 & ~A298;
  assign \new_[62476]_  = A301 & A300;
  assign \new_[62477]_  = \new_[62476]_  & \new_[62473]_ ;
  assign \new_[62478]_  = \new_[62477]_  & \new_[62470]_ ;
  assign \new_[62482]_  = ~A199 & ~A166;
  assign \new_[62483]_  = ~A167 & \new_[62482]_ ;
  assign \new_[62486]_  = A201 & A200;
  assign \new_[62489]_  = A265 & ~A203;
  assign \new_[62490]_  = \new_[62489]_  & \new_[62486]_ ;
  assign \new_[62491]_  = \new_[62490]_  & \new_[62483]_ ;
  assign \new_[62495]_  = A268 & A267;
  assign \new_[62496]_  = ~A266 & \new_[62495]_ ;
  assign \new_[62499]_  = A299 & ~A298;
  assign \new_[62502]_  = ~A302 & A300;
  assign \new_[62503]_  = \new_[62502]_  & \new_[62499]_ ;
  assign \new_[62504]_  = \new_[62503]_  & \new_[62496]_ ;
  assign \new_[62508]_  = ~A199 & ~A166;
  assign \new_[62509]_  = ~A167 & \new_[62508]_ ;
  assign \new_[62512]_  = A201 & A200;
  assign \new_[62515]_  = A265 & ~A203;
  assign \new_[62516]_  = \new_[62515]_  & \new_[62512]_ ;
  assign \new_[62517]_  = \new_[62516]_  & \new_[62509]_ ;
  assign \new_[62521]_  = ~A269 & A267;
  assign \new_[62522]_  = ~A266 & \new_[62521]_ ;
  assign \new_[62525]_  = ~A299 & A298;
  assign \new_[62528]_  = A301 & A300;
  assign \new_[62529]_  = \new_[62528]_  & \new_[62525]_ ;
  assign \new_[62530]_  = \new_[62529]_  & \new_[62522]_ ;
  assign \new_[62534]_  = ~A199 & ~A166;
  assign \new_[62535]_  = ~A167 & \new_[62534]_ ;
  assign \new_[62538]_  = A201 & A200;
  assign \new_[62541]_  = A265 & ~A203;
  assign \new_[62542]_  = \new_[62541]_  & \new_[62538]_ ;
  assign \new_[62543]_  = \new_[62542]_  & \new_[62535]_ ;
  assign \new_[62547]_  = ~A269 & A267;
  assign \new_[62548]_  = ~A266 & \new_[62547]_ ;
  assign \new_[62551]_  = ~A299 & A298;
  assign \new_[62554]_  = ~A302 & A300;
  assign \new_[62555]_  = \new_[62554]_  & \new_[62551]_ ;
  assign \new_[62556]_  = \new_[62555]_  & \new_[62548]_ ;
  assign \new_[62560]_  = ~A199 & ~A166;
  assign \new_[62561]_  = ~A167 & \new_[62560]_ ;
  assign \new_[62564]_  = A201 & A200;
  assign \new_[62567]_  = A265 & ~A203;
  assign \new_[62568]_  = \new_[62567]_  & \new_[62564]_ ;
  assign \new_[62569]_  = \new_[62568]_  & \new_[62561]_ ;
  assign \new_[62573]_  = ~A269 & A267;
  assign \new_[62574]_  = ~A266 & \new_[62573]_ ;
  assign \new_[62577]_  = A299 & ~A298;
  assign \new_[62580]_  = A301 & A300;
  assign \new_[62581]_  = \new_[62580]_  & \new_[62577]_ ;
  assign \new_[62582]_  = \new_[62581]_  & \new_[62574]_ ;
  assign \new_[62586]_  = ~A199 & ~A166;
  assign \new_[62587]_  = ~A167 & \new_[62586]_ ;
  assign \new_[62590]_  = A201 & A200;
  assign \new_[62593]_  = A265 & ~A203;
  assign \new_[62594]_  = \new_[62593]_  & \new_[62590]_ ;
  assign \new_[62595]_  = \new_[62594]_  & \new_[62587]_ ;
  assign \new_[62599]_  = ~A269 & A267;
  assign \new_[62600]_  = ~A266 & \new_[62599]_ ;
  assign \new_[62603]_  = A299 & ~A298;
  assign \new_[62606]_  = ~A302 & A300;
  assign \new_[62607]_  = \new_[62606]_  & \new_[62603]_ ;
  assign \new_[62608]_  = \new_[62607]_  & \new_[62600]_ ;
  assign \new_[62612]_  = A199 & ~A166;
  assign \new_[62613]_  = ~A167 & \new_[62612]_ ;
  assign \new_[62616]_  = A201 & ~A200;
  assign \new_[62619]_  = ~A265 & A202;
  assign \new_[62620]_  = \new_[62619]_  & \new_[62616]_ ;
  assign \new_[62621]_  = \new_[62620]_  & \new_[62613]_ ;
  assign \new_[62625]_  = A268 & A267;
  assign \new_[62626]_  = A266 & \new_[62625]_ ;
  assign \new_[62629]_  = ~A299 & A298;
  assign \new_[62632]_  = A301 & A300;
  assign \new_[62633]_  = \new_[62632]_  & \new_[62629]_ ;
  assign \new_[62634]_  = \new_[62633]_  & \new_[62626]_ ;
  assign \new_[62638]_  = A199 & ~A166;
  assign \new_[62639]_  = ~A167 & \new_[62638]_ ;
  assign \new_[62642]_  = A201 & ~A200;
  assign \new_[62645]_  = ~A265 & A202;
  assign \new_[62646]_  = \new_[62645]_  & \new_[62642]_ ;
  assign \new_[62647]_  = \new_[62646]_  & \new_[62639]_ ;
  assign \new_[62651]_  = A268 & A267;
  assign \new_[62652]_  = A266 & \new_[62651]_ ;
  assign \new_[62655]_  = ~A299 & A298;
  assign \new_[62658]_  = ~A302 & A300;
  assign \new_[62659]_  = \new_[62658]_  & \new_[62655]_ ;
  assign \new_[62660]_  = \new_[62659]_  & \new_[62652]_ ;
  assign \new_[62664]_  = A199 & ~A166;
  assign \new_[62665]_  = ~A167 & \new_[62664]_ ;
  assign \new_[62668]_  = A201 & ~A200;
  assign \new_[62671]_  = ~A265 & A202;
  assign \new_[62672]_  = \new_[62671]_  & \new_[62668]_ ;
  assign \new_[62673]_  = \new_[62672]_  & \new_[62665]_ ;
  assign \new_[62677]_  = A268 & A267;
  assign \new_[62678]_  = A266 & \new_[62677]_ ;
  assign \new_[62681]_  = A299 & ~A298;
  assign \new_[62684]_  = A301 & A300;
  assign \new_[62685]_  = \new_[62684]_  & \new_[62681]_ ;
  assign \new_[62686]_  = \new_[62685]_  & \new_[62678]_ ;
  assign \new_[62690]_  = A199 & ~A166;
  assign \new_[62691]_  = ~A167 & \new_[62690]_ ;
  assign \new_[62694]_  = A201 & ~A200;
  assign \new_[62697]_  = ~A265 & A202;
  assign \new_[62698]_  = \new_[62697]_  & \new_[62694]_ ;
  assign \new_[62699]_  = \new_[62698]_  & \new_[62691]_ ;
  assign \new_[62703]_  = A268 & A267;
  assign \new_[62704]_  = A266 & \new_[62703]_ ;
  assign \new_[62707]_  = A299 & ~A298;
  assign \new_[62710]_  = ~A302 & A300;
  assign \new_[62711]_  = \new_[62710]_  & \new_[62707]_ ;
  assign \new_[62712]_  = \new_[62711]_  & \new_[62704]_ ;
  assign \new_[62716]_  = A199 & ~A166;
  assign \new_[62717]_  = ~A167 & \new_[62716]_ ;
  assign \new_[62720]_  = A201 & ~A200;
  assign \new_[62723]_  = ~A265 & A202;
  assign \new_[62724]_  = \new_[62723]_  & \new_[62720]_ ;
  assign \new_[62725]_  = \new_[62724]_  & \new_[62717]_ ;
  assign \new_[62729]_  = ~A269 & A267;
  assign \new_[62730]_  = A266 & \new_[62729]_ ;
  assign \new_[62733]_  = ~A299 & A298;
  assign \new_[62736]_  = A301 & A300;
  assign \new_[62737]_  = \new_[62736]_  & \new_[62733]_ ;
  assign \new_[62738]_  = \new_[62737]_  & \new_[62730]_ ;
  assign \new_[62742]_  = A199 & ~A166;
  assign \new_[62743]_  = ~A167 & \new_[62742]_ ;
  assign \new_[62746]_  = A201 & ~A200;
  assign \new_[62749]_  = ~A265 & A202;
  assign \new_[62750]_  = \new_[62749]_  & \new_[62746]_ ;
  assign \new_[62751]_  = \new_[62750]_  & \new_[62743]_ ;
  assign \new_[62755]_  = ~A269 & A267;
  assign \new_[62756]_  = A266 & \new_[62755]_ ;
  assign \new_[62759]_  = ~A299 & A298;
  assign \new_[62762]_  = ~A302 & A300;
  assign \new_[62763]_  = \new_[62762]_  & \new_[62759]_ ;
  assign \new_[62764]_  = \new_[62763]_  & \new_[62756]_ ;
  assign \new_[62768]_  = A199 & ~A166;
  assign \new_[62769]_  = ~A167 & \new_[62768]_ ;
  assign \new_[62772]_  = A201 & ~A200;
  assign \new_[62775]_  = ~A265 & A202;
  assign \new_[62776]_  = \new_[62775]_  & \new_[62772]_ ;
  assign \new_[62777]_  = \new_[62776]_  & \new_[62769]_ ;
  assign \new_[62781]_  = ~A269 & A267;
  assign \new_[62782]_  = A266 & \new_[62781]_ ;
  assign \new_[62785]_  = A299 & ~A298;
  assign \new_[62788]_  = A301 & A300;
  assign \new_[62789]_  = \new_[62788]_  & \new_[62785]_ ;
  assign \new_[62790]_  = \new_[62789]_  & \new_[62782]_ ;
  assign \new_[62794]_  = A199 & ~A166;
  assign \new_[62795]_  = ~A167 & \new_[62794]_ ;
  assign \new_[62798]_  = A201 & ~A200;
  assign \new_[62801]_  = ~A265 & A202;
  assign \new_[62802]_  = \new_[62801]_  & \new_[62798]_ ;
  assign \new_[62803]_  = \new_[62802]_  & \new_[62795]_ ;
  assign \new_[62807]_  = ~A269 & A267;
  assign \new_[62808]_  = A266 & \new_[62807]_ ;
  assign \new_[62811]_  = A299 & ~A298;
  assign \new_[62814]_  = ~A302 & A300;
  assign \new_[62815]_  = \new_[62814]_  & \new_[62811]_ ;
  assign \new_[62816]_  = \new_[62815]_  & \new_[62808]_ ;
  assign \new_[62820]_  = A199 & ~A166;
  assign \new_[62821]_  = ~A167 & \new_[62820]_ ;
  assign \new_[62824]_  = A201 & ~A200;
  assign \new_[62827]_  = A265 & A202;
  assign \new_[62828]_  = \new_[62827]_  & \new_[62824]_ ;
  assign \new_[62829]_  = \new_[62828]_  & \new_[62821]_ ;
  assign \new_[62833]_  = A268 & A267;
  assign \new_[62834]_  = ~A266 & \new_[62833]_ ;
  assign \new_[62837]_  = ~A299 & A298;
  assign \new_[62840]_  = A301 & A300;
  assign \new_[62841]_  = \new_[62840]_  & \new_[62837]_ ;
  assign \new_[62842]_  = \new_[62841]_  & \new_[62834]_ ;
  assign \new_[62846]_  = A199 & ~A166;
  assign \new_[62847]_  = ~A167 & \new_[62846]_ ;
  assign \new_[62850]_  = A201 & ~A200;
  assign \new_[62853]_  = A265 & A202;
  assign \new_[62854]_  = \new_[62853]_  & \new_[62850]_ ;
  assign \new_[62855]_  = \new_[62854]_  & \new_[62847]_ ;
  assign \new_[62859]_  = A268 & A267;
  assign \new_[62860]_  = ~A266 & \new_[62859]_ ;
  assign \new_[62863]_  = ~A299 & A298;
  assign \new_[62866]_  = ~A302 & A300;
  assign \new_[62867]_  = \new_[62866]_  & \new_[62863]_ ;
  assign \new_[62868]_  = \new_[62867]_  & \new_[62860]_ ;
  assign \new_[62872]_  = A199 & ~A166;
  assign \new_[62873]_  = ~A167 & \new_[62872]_ ;
  assign \new_[62876]_  = A201 & ~A200;
  assign \new_[62879]_  = A265 & A202;
  assign \new_[62880]_  = \new_[62879]_  & \new_[62876]_ ;
  assign \new_[62881]_  = \new_[62880]_  & \new_[62873]_ ;
  assign \new_[62885]_  = A268 & A267;
  assign \new_[62886]_  = ~A266 & \new_[62885]_ ;
  assign \new_[62889]_  = A299 & ~A298;
  assign \new_[62892]_  = A301 & A300;
  assign \new_[62893]_  = \new_[62892]_  & \new_[62889]_ ;
  assign \new_[62894]_  = \new_[62893]_  & \new_[62886]_ ;
  assign \new_[62898]_  = A199 & ~A166;
  assign \new_[62899]_  = ~A167 & \new_[62898]_ ;
  assign \new_[62902]_  = A201 & ~A200;
  assign \new_[62905]_  = A265 & A202;
  assign \new_[62906]_  = \new_[62905]_  & \new_[62902]_ ;
  assign \new_[62907]_  = \new_[62906]_  & \new_[62899]_ ;
  assign \new_[62911]_  = A268 & A267;
  assign \new_[62912]_  = ~A266 & \new_[62911]_ ;
  assign \new_[62915]_  = A299 & ~A298;
  assign \new_[62918]_  = ~A302 & A300;
  assign \new_[62919]_  = \new_[62918]_  & \new_[62915]_ ;
  assign \new_[62920]_  = \new_[62919]_  & \new_[62912]_ ;
  assign \new_[62924]_  = A199 & ~A166;
  assign \new_[62925]_  = ~A167 & \new_[62924]_ ;
  assign \new_[62928]_  = A201 & ~A200;
  assign \new_[62931]_  = A265 & A202;
  assign \new_[62932]_  = \new_[62931]_  & \new_[62928]_ ;
  assign \new_[62933]_  = \new_[62932]_  & \new_[62925]_ ;
  assign \new_[62937]_  = ~A269 & A267;
  assign \new_[62938]_  = ~A266 & \new_[62937]_ ;
  assign \new_[62941]_  = ~A299 & A298;
  assign \new_[62944]_  = A301 & A300;
  assign \new_[62945]_  = \new_[62944]_  & \new_[62941]_ ;
  assign \new_[62946]_  = \new_[62945]_  & \new_[62938]_ ;
  assign \new_[62950]_  = A199 & ~A166;
  assign \new_[62951]_  = ~A167 & \new_[62950]_ ;
  assign \new_[62954]_  = A201 & ~A200;
  assign \new_[62957]_  = A265 & A202;
  assign \new_[62958]_  = \new_[62957]_  & \new_[62954]_ ;
  assign \new_[62959]_  = \new_[62958]_  & \new_[62951]_ ;
  assign \new_[62963]_  = ~A269 & A267;
  assign \new_[62964]_  = ~A266 & \new_[62963]_ ;
  assign \new_[62967]_  = ~A299 & A298;
  assign \new_[62970]_  = ~A302 & A300;
  assign \new_[62971]_  = \new_[62970]_  & \new_[62967]_ ;
  assign \new_[62972]_  = \new_[62971]_  & \new_[62964]_ ;
  assign \new_[62976]_  = A199 & ~A166;
  assign \new_[62977]_  = ~A167 & \new_[62976]_ ;
  assign \new_[62980]_  = A201 & ~A200;
  assign \new_[62983]_  = A265 & A202;
  assign \new_[62984]_  = \new_[62983]_  & \new_[62980]_ ;
  assign \new_[62985]_  = \new_[62984]_  & \new_[62977]_ ;
  assign \new_[62989]_  = ~A269 & A267;
  assign \new_[62990]_  = ~A266 & \new_[62989]_ ;
  assign \new_[62993]_  = A299 & ~A298;
  assign \new_[62996]_  = A301 & A300;
  assign \new_[62997]_  = \new_[62996]_  & \new_[62993]_ ;
  assign \new_[62998]_  = \new_[62997]_  & \new_[62990]_ ;
  assign \new_[63002]_  = A199 & ~A166;
  assign \new_[63003]_  = ~A167 & \new_[63002]_ ;
  assign \new_[63006]_  = A201 & ~A200;
  assign \new_[63009]_  = A265 & A202;
  assign \new_[63010]_  = \new_[63009]_  & \new_[63006]_ ;
  assign \new_[63011]_  = \new_[63010]_  & \new_[63003]_ ;
  assign \new_[63015]_  = ~A269 & A267;
  assign \new_[63016]_  = ~A266 & \new_[63015]_ ;
  assign \new_[63019]_  = A299 & ~A298;
  assign \new_[63022]_  = ~A302 & A300;
  assign \new_[63023]_  = \new_[63022]_  & \new_[63019]_ ;
  assign \new_[63024]_  = \new_[63023]_  & \new_[63016]_ ;
  assign \new_[63028]_  = A199 & ~A166;
  assign \new_[63029]_  = ~A167 & \new_[63028]_ ;
  assign \new_[63032]_  = A201 & ~A200;
  assign \new_[63035]_  = ~A265 & ~A203;
  assign \new_[63036]_  = \new_[63035]_  & \new_[63032]_ ;
  assign \new_[63037]_  = \new_[63036]_  & \new_[63029]_ ;
  assign \new_[63041]_  = A268 & A267;
  assign \new_[63042]_  = A266 & \new_[63041]_ ;
  assign \new_[63045]_  = ~A299 & A298;
  assign \new_[63048]_  = A301 & A300;
  assign \new_[63049]_  = \new_[63048]_  & \new_[63045]_ ;
  assign \new_[63050]_  = \new_[63049]_  & \new_[63042]_ ;
  assign \new_[63054]_  = A199 & ~A166;
  assign \new_[63055]_  = ~A167 & \new_[63054]_ ;
  assign \new_[63058]_  = A201 & ~A200;
  assign \new_[63061]_  = ~A265 & ~A203;
  assign \new_[63062]_  = \new_[63061]_  & \new_[63058]_ ;
  assign \new_[63063]_  = \new_[63062]_  & \new_[63055]_ ;
  assign \new_[63067]_  = A268 & A267;
  assign \new_[63068]_  = A266 & \new_[63067]_ ;
  assign \new_[63071]_  = ~A299 & A298;
  assign \new_[63074]_  = ~A302 & A300;
  assign \new_[63075]_  = \new_[63074]_  & \new_[63071]_ ;
  assign \new_[63076]_  = \new_[63075]_  & \new_[63068]_ ;
  assign \new_[63080]_  = A199 & ~A166;
  assign \new_[63081]_  = ~A167 & \new_[63080]_ ;
  assign \new_[63084]_  = A201 & ~A200;
  assign \new_[63087]_  = ~A265 & ~A203;
  assign \new_[63088]_  = \new_[63087]_  & \new_[63084]_ ;
  assign \new_[63089]_  = \new_[63088]_  & \new_[63081]_ ;
  assign \new_[63093]_  = A268 & A267;
  assign \new_[63094]_  = A266 & \new_[63093]_ ;
  assign \new_[63097]_  = A299 & ~A298;
  assign \new_[63100]_  = A301 & A300;
  assign \new_[63101]_  = \new_[63100]_  & \new_[63097]_ ;
  assign \new_[63102]_  = \new_[63101]_  & \new_[63094]_ ;
  assign \new_[63106]_  = A199 & ~A166;
  assign \new_[63107]_  = ~A167 & \new_[63106]_ ;
  assign \new_[63110]_  = A201 & ~A200;
  assign \new_[63113]_  = ~A265 & ~A203;
  assign \new_[63114]_  = \new_[63113]_  & \new_[63110]_ ;
  assign \new_[63115]_  = \new_[63114]_  & \new_[63107]_ ;
  assign \new_[63119]_  = A268 & A267;
  assign \new_[63120]_  = A266 & \new_[63119]_ ;
  assign \new_[63123]_  = A299 & ~A298;
  assign \new_[63126]_  = ~A302 & A300;
  assign \new_[63127]_  = \new_[63126]_  & \new_[63123]_ ;
  assign \new_[63128]_  = \new_[63127]_  & \new_[63120]_ ;
  assign \new_[63132]_  = A199 & ~A166;
  assign \new_[63133]_  = ~A167 & \new_[63132]_ ;
  assign \new_[63136]_  = A201 & ~A200;
  assign \new_[63139]_  = ~A265 & ~A203;
  assign \new_[63140]_  = \new_[63139]_  & \new_[63136]_ ;
  assign \new_[63141]_  = \new_[63140]_  & \new_[63133]_ ;
  assign \new_[63145]_  = ~A269 & A267;
  assign \new_[63146]_  = A266 & \new_[63145]_ ;
  assign \new_[63149]_  = ~A299 & A298;
  assign \new_[63152]_  = A301 & A300;
  assign \new_[63153]_  = \new_[63152]_  & \new_[63149]_ ;
  assign \new_[63154]_  = \new_[63153]_  & \new_[63146]_ ;
  assign \new_[63158]_  = A199 & ~A166;
  assign \new_[63159]_  = ~A167 & \new_[63158]_ ;
  assign \new_[63162]_  = A201 & ~A200;
  assign \new_[63165]_  = ~A265 & ~A203;
  assign \new_[63166]_  = \new_[63165]_  & \new_[63162]_ ;
  assign \new_[63167]_  = \new_[63166]_  & \new_[63159]_ ;
  assign \new_[63171]_  = ~A269 & A267;
  assign \new_[63172]_  = A266 & \new_[63171]_ ;
  assign \new_[63175]_  = ~A299 & A298;
  assign \new_[63178]_  = ~A302 & A300;
  assign \new_[63179]_  = \new_[63178]_  & \new_[63175]_ ;
  assign \new_[63180]_  = \new_[63179]_  & \new_[63172]_ ;
  assign \new_[63184]_  = A199 & ~A166;
  assign \new_[63185]_  = ~A167 & \new_[63184]_ ;
  assign \new_[63188]_  = A201 & ~A200;
  assign \new_[63191]_  = ~A265 & ~A203;
  assign \new_[63192]_  = \new_[63191]_  & \new_[63188]_ ;
  assign \new_[63193]_  = \new_[63192]_  & \new_[63185]_ ;
  assign \new_[63197]_  = ~A269 & A267;
  assign \new_[63198]_  = A266 & \new_[63197]_ ;
  assign \new_[63201]_  = A299 & ~A298;
  assign \new_[63204]_  = A301 & A300;
  assign \new_[63205]_  = \new_[63204]_  & \new_[63201]_ ;
  assign \new_[63206]_  = \new_[63205]_  & \new_[63198]_ ;
  assign \new_[63210]_  = A199 & ~A166;
  assign \new_[63211]_  = ~A167 & \new_[63210]_ ;
  assign \new_[63214]_  = A201 & ~A200;
  assign \new_[63217]_  = ~A265 & ~A203;
  assign \new_[63218]_  = \new_[63217]_  & \new_[63214]_ ;
  assign \new_[63219]_  = \new_[63218]_  & \new_[63211]_ ;
  assign \new_[63223]_  = ~A269 & A267;
  assign \new_[63224]_  = A266 & \new_[63223]_ ;
  assign \new_[63227]_  = A299 & ~A298;
  assign \new_[63230]_  = ~A302 & A300;
  assign \new_[63231]_  = \new_[63230]_  & \new_[63227]_ ;
  assign \new_[63232]_  = \new_[63231]_  & \new_[63224]_ ;
  assign \new_[63236]_  = A199 & ~A166;
  assign \new_[63237]_  = ~A167 & \new_[63236]_ ;
  assign \new_[63240]_  = A201 & ~A200;
  assign \new_[63243]_  = A265 & ~A203;
  assign \new_[63244]_  = \new_[63243]_  & \new_[63240]_ ;
  assign \new_[63245]_  = \new_[63244]_  & \new_[63237]_ ;
  assign \new_[63249]_  = A268 & A267;
  assign \new_[63250]_  = ~A266 & \new_[63249]_ ;
  assign \new_[63253]_  = ~A299 & A298;
  assign \new_[63256]_  = A301 & A300;
  assign \new_[63257]_  = \new_[63256]_  & \new_[63253]_ ;
  assign \new_[63258]_  = \new_[63257]_  & \new_[63250]_ ;
  assign \new_[63262]_  = A199 & ~A166;
  assign \new_[63263]_  = ~A167 & \new_[63262]_ ;
  assign \new_[63266]_  = A201 & ~A200;
  assign \new_[63269]_  = A265 & ~A203;
  assign \new_[63270]_  = \new_[63269]_  & \new_[63266]_ ;
  assign \new_[63271]_  = \new_[63270]_  & \new_[63263]_ ;
  assign \new_[63275]_  = A268 & A267;
  assign \new_[63276]_  = ~A266 & \new_[63275]_ ;
  assign \new_[63279]_  = ~A299 & A298;
  assign \new_[63282]_  = ~A302 & A300;
  assign \new_[63283]_  = \new_[63282]_  & \new_[63279]_ ;
  assign \new_[63284]_  = \new_[63283]_  & \new_[63276]_ ;
  assign \new_[63288]_  = A199 & ~A166;
  assign \new_[63289]_  = ~A167 & \new_[63288]_ ;
  assign \new_[63292]_  = A201 & ~A200;
  assign \new_[63295]_  = A265 & ~A203;
  assign \new_[63296]_  = \new_[63295]_  & \new_[63292]_ ;
  assign \new_[63297]_  = \new_[63296]_  & \new_[63289]_ ;
  assign \new_[63301]_  = A268 & A267;
  assign \new_[63302]_  = ~A266 & \new_[63301]_ ;
  assign \new_[63305]_  = A299 & ~A298;
  assign \new_[63308]_  = A301 & A300;
  assign \new_[63309]_  = \new_[63308]_  & \new_[63305]_ ;
  assign \new_[63310]_  = \new_[63309]_  & \new_[63302]_ ;
  assign \new_[63314]_  = A199 & ~A166;
  assign \new_[63315]_  = ~A167 & \new_[63314]_ ;
  assign \new_[63318]_  = A201 & ~A200;
  assign \new_[63321]_  = A265 & ~A203;
  assign \new_[63322]_  = \new_[63321]_  & \new_[63318]_ ;
  assign \new_[63323]_  = \new_[63322]_  & \new_[63315]_ ;
  assign \new_[63327]_  = A268 & A267;
  assign \new_[63328]_  = ~A266 & \new_[63327]_ ;
  assign \new_[63331]_  = A299 & ~A298;
  assign \new_[63334]_  = ~A302 & A300;
  assign \new_[63335]_  = \new_[63334]_  & \new_[63331]_ ;
  assign \new_[63336]_  = \new_[63335]_  & \new_[63328]_ ;
  assign \new_[63340]_  = A199 & ~A166;
  assign \new_[63341]_  = ~A167 & \new_[63340]_ ;
  assign \new_[63344]_  = A201 & ~A200;
  assign \new_[63347]_  = A265 & ~A203;
  assign \new_[63348]_  = \new_[63347]_  & \new_[63344]_ ;
  assign \new_[63349]_  = \new_[63348]_  & \new_[63341]_ ;
  assign \new_[63353]_  = ~A269 & A267;
  assign \new_[63354]_  = ~A266 & \new_[63353]_ ;
  assign \new_[63357]_  = ~A299 & A298;
  assign \new_[63360]_  = A301 & A300;
  assign \new_[63361]_  = \new_[63360]_  & \new_[63357]_ ;
  assign \new_[63362]_  = \new_[63361]_  & \new_[63354]_ ;
  assign \new_[63366]_  = A199 & ~A166;
  assign \new_[63367]_  = ~A167 & \new_[63366]_ ;
  assign \new_[63370]_  = A201 & ~A200;
  assign \new_[63373]_  = A265 & ~A203;
  assign \new_[63374]_  = \new_[63373]_  & \new_[63370]_ ;
  assign \new_[63375]_  = \new_[63374]_  & \new_[63367]_ ;
  assign \new_[63379]_  = ~A269 & A267;
  assign \new_[63380]_  = ~A266 & \new_[63379]_ ;
  assign \new_[63383]_  = ~A299 & A298;
  assign \new_[63386]_  = ~A302 & A300;
  assign \new_[63387]_  = \new_[63386]_  & \new_[63383]_ ;
  assign \new_[63388]_  = \new_[63387]_  & \new_[63380]_ ;
  assign \new_[63392]_  = A199 & ~A166;
  assign \new_[63393]_  = ~A167 & \new_[63392]_ ;
  assign \new_[63396]_  = A201 & ~A200;
  assign \new_[63399]_  = A265 & ~A203;
  assign \new_[63400]_  = \new_[63399]_  & \new_[63396]_ ;
  assign \new_[63401]_  = \new_[63400]_  & \new_[63393]_ ;
  assign \new_[63405]_  = ~A269 & A267;
  assign \new_[63406]_  = ~A266 & \new_[63405]_ ;
  assign \new_[63409]_  = A299 & ~A298;
  assign \new_[63412]_  = A301 & A300;
  assign \new_[63413]_  = \new_[63412]_  & \new_[63409]_ ;
  assign \new_[63414]_  = \new_[63413]_  & \new_[63406]_ ;
  assign \new_[63418]_  = A199 & ~A166;
  assign \new_[63419]_  = ~A167 & \new_[63418]_ ;
  assign \new_[63422]_  = A201 & ~A200;
  assign \new_[63425]_  = A265 & ~A203;
  assign \new_[63426]_  = \new_[63425]_  & \new_[63422]_ ;
  assign \new_[63427]_  = \new_[63426]_  & \new_[63419]_ ;
  assign \new_[63431]_  = ~A269 & A267;
  assign \new_[63432]_  = ~A266 & \new_[63431]_ ;
  assign \new_[63435]_  = A299 & ~A298;
  assign \new_[63438]_  = ~A302 & A300;
  assign \new_[63439]_  = \new_[63438]_  & \new_[63435]_ ;
  assign \new_[63440]_  = \new_[63439]_  & \new_[63432]_ ;
  assign \new_[63444]_  = A167 & A168;
  assign \new_[63445]_  = A170 & \new_[63444]_ ;
  assign \new_[63448]_  = A201 & ~A166;
  assign \new_[63451]_  = A203 & ~A202;
  assign \new_[63452]_  = \new_[63451]_  & \new_[63448]_ ;
  assign \new_[63453]_  = \new_[63452]_  & \new_[63445]_ ;
  assign \new_[63457]_  = A269 & ~A268;
  assign \new_[63458]_  = A267 & \new_[63457]_ ;
  assign \new_[63461]_  = ~A299 & A298;
  assign \new_[63464]_  = A301 & A300;
  assign \new_[63465]_  = \new_[63464]_  & \new_[63461]_ ;
  assign \new_[63466]_  = \new_[63465]_  & \new_[63458]_ ;
  assign \new_[63470]_  = A167 & A168;
  assign \new_[63471]_  = A170 & \new_[63470]_ ;
  assign \new_[63474]_  = A201 & ~A166;
  assign \new_[63477]_  = A203 & ~A202;
  assign \new_[63478]_  = \new_[63477]_  & \new_[63474]_ ;
  assign \new_[63479]_  = \new_[63478]_  & \new_[63471]_ ;
  assign \new_[63483]_  = A269 & ~A268;
  assign \new_[63484]_  = A267 & \new_[63483]_ ;
  assign \new_[63487]_  = ~A299 & A298;
  assign \new_[63490]_  = ~A302 & A300;
  assign \new_[63491]_  = \new_[63490]_  & \new_[63487]_ ;
  assign \new_[63492]_  = \new_[63491]_  & \new_[63484]_ ;
  assign \new_[63496]_  = A167 & A168;
  assign \new_[63497]_  = A170 & \new_[63496]_ ;
  assign \new_[63500]_  = A201 & ~A166;
  assign \new_[63503]_  = A203 & ~A202;
  assign \new_[63504]_  = \new_[63503]_  & \new_[63500]_ ;
  assign \new_[63505]_  = \new_[63504]_  & \new_[63497]_ ;
  assign \new_[63509]_  = A269 & ~A268;
  assign \new_[63510]_  = A267 & \new_[63509]_ ;
  assign \new_[63513]_  = A299 & ~A298;
  assign \new_[63516]_  = A301 & A300;
  assign \new_[63517]_  = \new_[63516]_  & \new_[63513]_ ;
  assign \new_[63518]_  = \new_[63517]_  & \new_[63510]_ ;
  assign \new_[63522]_  = A167 & A168;
  assign \new_[63523]_  = A170 & \new_[63522]_ ;
  assign \new_[63526]_  = A201 & ~A166;
  assign \new_[63529]_  = A203 & ~A202;
  assign \new_[63530]_  = \new_[63529]_  & \new_[63526]_ ;
  assign \new_[63531]_  = \new_[63530]_  & \new_[63523]_ ;
  assign \new_[63535]_  = A269 & ~A268;
  assign \new_[63536]_  = A267 & \new_[63535]_ ;
  assign \new_[63539]_  = A299 & ~A298;
  assign \new_[63542]_  = ~A302 & A300;
  assign \new_[63543]_  = \new_[63542]_  & \new_[63539]_ ;
  assign \new_[63544]_  = \new_[63543]_  & \new_[63536]_ ;
  assign \new_[63548]_  = A167 & A168;
  assign \new_[63549]_  = A170 & \new_[63548]_ ;
  assign \new_[63552]_  = A201 & ~A166;
  assign \new_[63555]_  = A203 & ~A202;
  assign \new_[63556]_  = \new_[63555]_  & \new_[63552]_ ;
  assign \new_[63557]_  = \new_[63556]_  & \new_[63549]_ ;
  assign \new_[63561]_  = A298 & A268;
  assign \new_[63562]_  = ~A267 & \new_[63561]_ ;
  assign \new_[63565]_  = ~A300 & ~A299;
  assign \new_[63568]_  = A302 & ~A301;
  assign \new_[63569]_  = \new_[63568]_  & \new_[63565]_ ;
  assign \new_[63570]_  = \new_[63569]_  & \new_[63562]_ ;
  assign \new_[63574]_  = A167 & A168;
  assign \new_[63575]_  = A170 & \new_[63574]_ ;
  assign \new_[63578]_  = A201 & ~A166;
  assign \new_[63581]_  = A203 & ~A202;
  assign \new_[63582]_  = \new_[63581]_  & \new_[63578]_ ;
  assign \new_[63583]_  = \new_[63582]_  & \new_[63575]_ ;
  assign \new_[63587]_  = ~A298 & A268;
  assign \new_[63588]_  = ~A267 & \new_[63587]_ ;
  assign \new_[63591]_  = ~A300 & A299;
  assign \new_[63594]_  = A302 & ~A301;
  assign \new_[63595]_  = \new_[63594]_  & \new_[63591]_ ;
  assign \new_[63596]_  = \new_[63595]_  & \new_[63588]_ ;
  assign \new_[63600]_  = A167 & A168;
  assign \new_[63601]_  = A170 & \new_[63600]_ ;
  assign \new_[63604]_  = A201 & ~A166;
  assign \new_[63607]_  = A203 & ~A202;
  assign \new_[63608]_  = \new_[63607]_  & \new_[63604]_ ;
  assign \new_[63609]_  = \new_[63608]_  & \new_[63601]_ ;
  assign \new_[63613]_  = A298 & ~A269;
  assign \new_[63614]_  = ~A267 & \new_[63613]_ ;
  assign \new_[63617]_  = ~A300 & ~A299;
  assign \new_[63620]_  = A302 & ~A301;
  assign \new_[63621]_  = \new_[63620]_  & \new_[63617]_ ;
  assign \new_[63622]_  = \new_[63621]_  & \new_[63614]_ ;
  assign \new_[63626]_  = A167 & A168;
  assign \new_[63627]_  = A170 & \new_[63626]_ ;
  assign \new_[63630]_  = A201 & ~A166;
  assign \new_[63633]_  = A203 & ~A202;
  assign \new_[63634]_  = \new_[63633]_  & \new_[63630]_ ;
  assign \new_[63635]_  = \new_[63634]_  & \new_[63627]_ ;
  assign \new_[63639]_  = ~A298 & ~A269;
  assign \new_[63640]_  = ~A267 & \new_[63639]_ ;
  assign \new_[63643]_  = ~A300 & A299;
  assign \new_[63646]_  = A302 & ~A301;
  assign \new_[63647]_  = \new_[63646]_  & \new_[63643]_ ;
  assign \new_[63648]_  = \new_[63647]_  & \new_[63640]_ ;
  assign \new_[63652]_  = A167 & A168;
  assign \new_[63653]_  = A170 & \new_[63652]_ ;
  assign \new_[63656]_  = A201 & ~A166;
  assign \new_[63659]_  = A203 & ~A202;
  assign \new_[63660]_  = \new_[63659]_  & \new_[63656]_ ;
  assign \new_[63661]_  = \new_[63660]_  & \new_[63653]_ ;
  assign \new_[63665]_  = A298 & A266;
  assign \new_[63666]_  = A265 & \new_[63665]_ ;
  assign \new_[63669]_  = ~A300 & ~A299;
  assign \new_[63672]_  = A302 & ~A301;
  assign \new_[63673]_  = \new_[63672]_  & \new_[63669]_ ;
  assign \new_[63674]_  = \new_[63673]_  & \new_[63666]_ ;
  assign \new_[63678]_  = A167 & A168;
  assign \new_[63679]_  = A170 & \new_[63678]_ ;
  assign \new_[63682]_  = A201 & ~A166;
  assign \new_[63685]_  = A203 & ~A202;
  assign \new_[63686]_  = \new_[63685]_  & \new_[63682]_ ;
  assign \new_[63687]_  = \new_[63686]_  & \new_[63679]_ ;
  assign \new_[63691]_  = ~A298 & A266;
  assign \new_[63692]_  = A265 & \new_[63691]_ ;
  assign \new_[63695]_  = ~A300 & A299;
  assign \new_[63698]_  = A302 & ~A301;
  assign \new_[63699]_  = \new_[63698]_  & \new_[63695]_ ;
  assign \new_[63700]_  = \new_[63699]_  & \new_[63692]_ ;
  assign \new_[63704]_  = A167 & A168;
  assign \new_[63705]_  = A170 & \new_[63704]_ ;
  assign \new_[63708]_  = A201 & ~A166;
  assign \new_[63711]_  = A203 & ~A202;
  assign \new_[63712]_  = \new_[63711]_  & \new_[63708]_ ;
  assign \new_[63713]_  = \new_[63712]_  & \new_[63705]_ ;
  assign \new_[63717]_  = A267 & A266;
  assign \new_[63718]_  = ~A265 & \new_[63717]_ ;
  assign \new_[63721]_  = A300 & A268;
  assign \new_[63724]_  = A302 & ~A301;
  assign \new_[63725]_  = \new_[63724]_  & \new_[63721]_ ;
  assign \new_[63726]_  = \new_[63725]_  & \new_[63718]_ ;
  assign \new_[63730]_  = A167 & A168;
  assign \new_[63731]_  = A170 & \new_[63730]_ ;
  assign \new_[63734]_  = A201 & ~A166;
  assign \new_[63737]_  = A203 & ~A202;
  assign \new_[63738]_  = \new_[63737]_  & \new_[63734]_ ;
  assign \new_[63739]_  = \new_[63738]_  & \new_[63731]_ ;
  assign \new_[63743]_  = A267 & A266;
  assign \new_[63744]_  = ~A265 & \new_[63743]_ ;
  assign \new_[63747]_  = A300 & ~A269;
  assign \new_[63750]_  = A302 & ~A301;
  assign \new_[63751]_  = \new_[63750]_  & \new_[63747]_ ;
  assign \new_[63752]_  = \new_[63751]_  & \new_[63744]_ ;
  assign \new_[63756]_  = A167 & A168;
  assign \new_[63757]_  = A170 & \new_[63756]_ ;
  assign \new_[63760]_  = A201 & ~A166;
  assign \new_[63763]_  = A203 & ~A202;
  assign \new_[63764]_  = \new_[63763]_  & \new_[63760]_ ;
  assign \new_[63765]_  = \new_[63764]_  & \new_[63757]_ ;
  assign \new_[63769]_  = ~A267 & A266;
  assign \new_[63770]_  = ~A265 & \new_[63769]_ ;
  assign \new_[63773]_  = A269 & ~A268;
  assign \new_[63776]_  = A301 & ~A300;
  assign \new_[63777]_  = \new_[63776]_  & \new_[63773]_ ;
  assign \new_[63778]_  = \new_[63777]_  & \new_[63770]_ ;
  assign \new_[63782]_  = A167 & A168;
  assign \new_[63783]_  = A170 & \new_[63782]_ ;
  assign \new_[63786]_  = A201 & ~A166;
  assign \new_[63789]_  = A203 & ~A202;
  assign \new_[63790]_  = \new_[63789]_  & \new_[63786]_ ;
  assign \new_[63791]_  = \new_[63790]_  & \new_[63783]_ ;
  assign \new_[63795]_  = ~A267 & A266;
  assign \new_[63796]_  = ~A265 & \new_[63795]_ ;
  assign \new_[63799]_  = A269 & ~A268;
  assign \new_[63802]_  = ~A302 & ~A300;
  assign \new_[63803]_  = \new_[63802]_  & \new_[63799]_ ;
  assign \new_[63804]_  = \new_[63803]_  & \new_[63796]_ ;
  assign \new_[63808]_  = A167 & A168;
  assign \new_[63809]_  = A170 & \new_[63808]_ ;
  assign \new_[63812]_  = A201 & ~A166;
  assign \new_[63815]_  = A203 & ~A202;
  assign \new_[63816]_  = \new_[63815]_  & \new_[63812]_ ;
  assign \new_[63817]_  = \new_[63816]_  & \new_[63809]_ ;
  assign \new_[63821]_  = ~A267 & A266;
  assign \new_[63822]_  = ~A265 & \new_[63821]_ ;
  assign \new_[63825]_  = A269 & ~A268;
  assign \new_[63828]_  = A299 & A298;
  assign \new_[63829]_  = \new_[63828]_  & \new_[63825]_ ;
  assign \new_[63830]_  = \new_[63829]_  & \new_[63822]_ ;
  assign \new_[63834]_  = A167 & A168;
  assign \new_[63835]_  = A170 & \new_[63834]_ ;
  assign \new_[63838]_  = A201 & ~A166;
  assign \new_[63841]_  = A203 & ~A202;
  assign \new_[63842]_  = \new_[63841]_  & \new_[63838]_ ;
  assign \new_[63843]_  = \new_[63842]_  & \new_[63835]_ ;
  assign \new_[63847]_  = ~A267 & A266;
  assign \new_[63848]_  = ~A265 & \new_[63847]_ ;
  assign \new_[63851]_  = A269 & ~A268;
  assign \new_[63854]_  = ~A299 & ~A298;
  assign \new_[63855]_  = \new_[63854]_  & \new_[63851]_ ;
  assign \new_[63856]_  = \new_[63855]_  & \new_[63848]_ ;
  assign \new_[63860]_  = A167 & A168;
  assign \new_[63861]_  = A170 & \new_[63860]_ ;
  assign \new_[63864]_  = A201 & ~A166;
  assign \new_[63867]_  = A203 & ~A202;
  assign \new_[63868]_  = \new_[63867]_  & \new_[63864]_ ;
  assign \new_[63869]_  = \new_[63868]_  & \new_[63861]_ ;
  assign \new_[63873]_  = A267 & ~A266;
  assign \new_[63874]_  = A265 & \new_[63873]_ ;
  assign \new_[63877]_  = A300 & A268;
  assign \new_[63880]_  = A302 & ~A301;
  assign \new_[63881]_  = \new_[63880]_  & \new_[63877]_ ;
  assign \new_[63882]_  = \new_[63881]_  & \new_[63874]_ ;
  assign \new_[63886]_  = A167 & A168;
  assign \new_[63887]_  = A170 & \new_[63886]_ ;
  assign \new_[63890]_  = A201 & ~A166;
  assign \new_[63893]_  = A203 & ~A202;
  assign \new_[63894]_  = \new_[63893]_  & \new_[63890]_ ;
  assign \new_[63895]_  = \new_[63894]_  & \new_[63887]_ ;
  assign \new_[63899]_  = A267 & ~A266;
  assign \new_[63900]_  = A265 & \new_[63899]_ ;
  assign \new_[63903]_  = A300 & ~A269;
  assign \new_[63906]_  = A302 & ~A301;
  assign \new_[63907]_  = \new_[63906]_  & \new_[63903]_ ;
  assign \new_[63908]_  = \new_[63907]_  & \new_[63900]_ ;
  assign \new_[63912]_  = A167 & A168;
  assign \new_[63913]_  = A170 & \new_[63912]_ ;
  assign \new_[63916]_  = A201 & ~A166;
  assign \new_[63919]_  = A203 & ~A202;
  assign \new_[63920]_  = \new_[63919]_  & \new_[63916]_ ;
  assign \new_[63921]_  = \new_[63920]_  & \new_[63913]_ ;
  assign \new_[63925]_  = ~A267 & ~A266;
  assign \new_[63926]_  = A265 & \new_[63925]_ ;
  assign \new_[63929]_  = A269 & ~A268;
  assign \new_[63932]_  = A301 & ~A300;
  assign \new_[63933]_  = \new_[63932]_  & \new_[63929]_ ;
  assign \new_[63934]_  = \new_[63933]_  & \new_[63926]_ ;
  assign \new_[63938]_  = A167 & A168;
  assign \new_[63939]_  = A170 & \new_[63938]_ ;
  assign \new_[63942]_  = A201 & ~A166;
  assign \new_[63945]_  = A203 & ~A202;
  assign \new_[63946]_  = \new_[63945]_  & \new_[63942]_ ;
  assign \new_[63947]_  = \new_[63946]_  & \new_[63939]_ ;
  assign \new_[63951]_  = ~A267 & ~A266;
  assign \new_[63952]_  = A265 & \new_[63951]_ ;
  assign \new_[63955]_  = A269 & ~A268;
  assign \new_[63958]_  = ~A302 & ~A300;
  assign \new_[63959]_  = \new_[63958]_  & \new_[63955]_ ;
  assign \new_[63960]_  = \new_[63959]_  & \new_[63952]_ ;
  assign \new_[63964]_  = A167 & A168;
  assign \new_[63965]_  = A170 & \new_[63964]_ ;
  assign \new_[63968]_  = A201 & ~A166;
  assign \new_[63971]_  = A203 & ~A202;
  assign \new_[63972]_  = \new_[63971]_  & \new_[63968]_ ;
  assign \new_[63973]_  = \new_[63972]_  & \new_[63965]_ ;
  assign \new_[63977]_  = ~A267 & ~A266;
  assign \new_[63978]_  = A265 & \new_[63977]_ ;
  assign \new_[63981]_  = A269 & ~A268;
  assign \new_[63984]_  = A299 & A298;
  assign \new_[63985]_  = \new_[63984]_  & \new_[63981]_ ;
  assign \new_[63986]_  = \new_[63985]_  & \new_[63978]_ ;
  assign \new_[63990]_  = A167 & A168;
  assign \new_[63991]_  = A170 & \new_[63990]_ ;
  assign \new_[63994]_  = A201 & ~A166;
  assign \new_[63997]_  = A203 & ~A202;
  assign \new_[63998]_  = \new_[63997]_  & \new_[63994]_ ;
  assign \new_[63999]_  = \new_[63998]_  & \new_[63991]_ ;
  assign \new_[64003]_  = ~A267 & ~A266;
  assign \new_[64004]_  = A265 & \new_[64003]_ ;
  assign \new_[64007]_  = A269 & ~A268;
  assign \new_[64010]_  = ~A299 & ~A298;
  assign \new_[64011]_  = \new_[64010]_  & \new_[64007]_ ;
  assign \new_[64012]_  = \new_[64011]_  & \new_[64004]_ ;
  assign \new_[64016]_  = A167 & A168;
  assign \new_[64017]_  = A170 & \new_[64016]_ ;
  assign \new_[64020]_  = A201 & ~A166;
  assign \new_[64023]_  = A203 & ~A202;
  assign \new_[64024]_  = \new_[64023]_  & \new_[64020]_ ;
  assign \new_[64025]_  = \new_[64024]_  & \new_[64017]_ ;
  assign \new_[64029]_  = A298 & ~A266;
  assign \new_[64030]_  = ~A265 & \new_[64029]_ ;
  assign \new_[64033]_  = ~A300 & ~A299;
  assign \new_[64036]_  = A302 & ~A301;
  assign \new_[64037]_  = \new_[64036]_  & \new_[64033]_ ;
  assign \new_[64038]_  = \new_[64037]_  & \new_[64030]_ ;
  assign \new_[64042]_  = A167 & A168;
  assign \new_[64043]_  = A170 & \new_[64042]_ ;
  assign \new_[64046]_  = A201 & ~A166;
  assign \new_[64049]_  = A203 & ~A202;
  assign \new_[64050]_  = \new_[64049]_  & \new_[64046]_ ;
  assign \new_[64051]_  = \new_[64050]_  & \new_[64043]_ ;
  assign \new_[64055]_  = ~A298 & ~A266;
  assign \new_[64056]_  = ~A265 & \new_[64055]_ ;
  assign \new_[64059]_  = ~A300 & A299;
  assign \new_[64062]_  = A302 & ~A301;
  assign \new_[64063]_  = \new_[64062]_  & \new_[64059]_ ;
  assign \new_[64064]_  = \new_[64063]_  & \new_[64056]_ ;
  assign \new_[64068]_  = A167 & A168;
  assign \new_[64069]_  = A170 & \new_[64068]_ ;
  assign \new_[64072]_  = ~A201 & ~A166;
  assign \new_[64075]_  = A267 & A202;
  assign \new_[64076]_  = \new_[64075]_  & \new_[64072]_ ;
  assign \new_[64077]_  = \new_[64076]_  & \new_[64069]_ ;
  assign \new_[64081]_  = A298 & A269;
  assign \new_[64082]_  = ~A268 & \new_[64081]_ ;
  assign \new_[64085]_  = ~A300 & ~A299;
  assign \new_[64088]_  = A302 & ~A301;
  assign \new_[64089]_  = \new_[64088]_  & \new_[64085]_ ;
  assign \new_[64090]_  = \new_[64089]_  & \new_[64082]_ ;
  assign \new_[64094]_  = A167 & A168;
  assign \new_[64095]_  = A170 & \new_[64094]_ ;
  assign \new_[64098]_  = ~A201 & ~A166;
  assign \new_[64101]_  = A267 & A202;
  assign \new_[64102]_  = \new_[64101]_  & \new_[64098]_ ;
  assign \new_[64103]_  = \new_[64102]_  & \new_[64095]_ ;
  assign \new_[64107]_  = ~A298 & A269;
  assign \new_[64108]_  = ~A268 & \new_[64107]_ ;
  assign \new_[64111]_  = ~A300 & A299;
  assign \new_[64114]_  = A302 & ~A301;
  assign \new_[64115]_  = \new_[64114]_  & \new_[64111]_ ;
  assign \new_[64116]_  = \new_[64115]_  & \new_[64108]_ ;
  assign \new_[64120]_  = A167 & A168;
  assign \new_[64121]_  = A170 & \new_[64120]_ ;
  assign \new_[64124]_  = ~A201 & ~A166;
  assign \new_[64127]_  = ~A265 & A202;
  assign \new_[64128]_  = \new_[64127]_  & \new_[64124]_ ;
  assign \new_[64129]_  = \new_[64128]_  & \new_[64121]_ ;
  assign \new_[64133]_  = ~A268 & ~A267;
  assign \new_[64134]_  = A266 & \new_[64133]_ ;
  assign \new_[64137]_  = A300 & A269;
  assign \new_[64140]_  = A302 & ~A301;
  assign \new_[64141]_  = \new_[64140]_  & \new_[64137]_ ;
  assign \new_[64142]_  = \new_[64141]_  & \new_[64134]_ ;
  assign \new_[64146]_  = A167 & A168;
  assign \new_[64147]_  = A170 & \new_[64146]_ ;
  assign \new_[64150]_  = ~A201 & ~A166;
  assign \new_[64153]_  = A265 & A202;
  assign \new_[64154]_  = \new_[64153]_  & \new_[64150]_ ;
  assign \new_[64155]_  = \new_[64154]_  & \new_[64147]_ ;
  assign \new_[64159]_  = ~A268 & ~A267;
  assign \new_[64160]_  = ~A266 & \new_[64159]_ ;
  assign \new_[64163]_  = A300 & A269;
  assign \new_[64166]_  = A302 & ~A301;
  assign \new_[64167]_  = \new_[64166]_  & \new_[64163]_ ;
  assign \new_[64168]_  = \new_[64167]_  & \new_[64160]_ ;
  assign \new_[64172]_  = A167 & A168;
  assign \new_[64173]_  = A170 & \new_[64172]_ ;
  assign \new_[64176]_  = ~A201 & ~A166;
  assign \new_[64179]_  = A267 & ~A203;
  assign \new_[64180]_  = \new_[64179]_  & \new_[64176]_ ;
  assign \new_[64181]_  = \new_[64180]_  & \new_[64173]_ ;
  assign \new_[64185]_  = A298 & A269;
  assign \new_[64186]_  = ~A268 & \new_[64185]_ ;
  assign \new_[64189]_  = ~A300 & ~A299;
  assign \new_[64192]_  = A302 & ~A301;
  assign \new_[64193]_  = \new_[64192]_  & \new_[64189]_ ;
  assign \new_[64194]_  = \new_[64193]_  & \new_[64186]_ ;
  assign \new_[64198]_  = A167 & A168;
  assign \new_[64199]_  = A170 & \new_[64198]_ ;
  assign \new_[64202]_  = ~A201 & ~A166;
  assign \new_[64205]_  = A267 & ~A203;
  assign \new_[64206]_  = \new_[64205]_  & \new_[64202]_ ;
  assign \new_[64207]_  = \new_[64206]_  & \new_[64199]_ ;
  assign \new_[64211]_  = ~A298 & A269;
  assign \new_[64212]_  = ~A268 & \new_[64211]_ ;
  assign \new_[64215]_  = ~A300 & A299;
  assign \new_[64218]_  = A302 & ~A301;
  assign \new_[64219]_  = \new_[64218]_  & \new_[64215]_ ;
  assign \new_[64220]_  = \new_[64219]_  & \new_[64212]_ ;
  assign \new_[64224]_  = A167 & A168;
  assign \new_[64225]_  = A170 & \new_[64224]_ ;
  assign \new_[64228]_  = ~A201 & ~A166;
  assign \new_[64231]_  = ~A265 & ~A203;
  assign \new_[64232]_  = \new_[64231]_  & \new_[64228]_ ;
  assign \new_[64233]_  = \new_[64232]_  & \new_[64225]_ ;
  assign \new_[64237]_  = ~A268 & ~A267;
  assign \new_[64238]_  = A266 & \new_[64237]_ ;
  assign \new_[64241]_  = A300 & A269;
  assign \new_[64244]_  = A302 & ~A301;
  assign \new_[64245]_  = \new_[64244]_  & \new_[64241]_ ;
  assign \new_[64246]_  = \new_[64245]_  & \new_[64238]_ ;
  assign \new_[64250]_  = A167 & A168;
  assign \new_[64251]_  = A170 & \new_[64250]_ ;
  assign \new_[64254]_  = ~A201 & ~A166;
  assign \new_[64257]_  = A265 & ~A203;
  assign \new_[64258]_  = \new_[64257]_  & \new_[64254]_ ;
  assign \new_[64259]_  = \new_[64258]_  & \new_[64251]_ ;
  assign \new_[64263]_  = ~A268 & ~A267;
  assign \new_[64264]_  = ~A266 & \new_[64263]_ ;
  assign \new_[64267]_  = A300 & A269;
  assign \new_[64270]_  = A302 & ~A301;
  assign \new_[64271]_  = \new_[64270]_  & \new_[64267]_ ;
  assign \new_[64272]_  = \new_[64271]_  & \new_[64264]_ ;
  assign \new_[64276]_  = A167 & A168;
  assign \new_[64277]_  = A170 & \new_[64276]_ ;
  assign \new_[64280]_  = A199 & ~A166;
  assign \new_[64283]_  = A267 & A200;
  assign \new_[64284]_  = \new_[64283]_  & \new_[64280]_ ;
  assign \new_[64285]_  = \new_[64284]_  & \new_[64277]_ ;
  assign \new_[64289]_  = A298 & A269;
  assign \new_[64290]_  = ~A268 & \new_[64289]_ ;
  assign \new_[64293]_  = ~A300 & ~A299;
  assign \new_[64296]_  = A302 & ~A301;
  assign \new_[64297]_  = \new_[64296]_  & \new_[64293]_ ;
  assign \new_[64298]_  = \new_[64297]_  & \new_[64290]_ ;
  assign \new_[64302]_  = A167 & A168;
  assign \new_[64303]_  = A170 & \new_[64302]_ ;
  assign \new_[64306]_  = A199 & ~A166;
  assign \new_[64309]_  = A267 & A200;
  assign \new_[64310]_  = \new_[64309]_  & \new_[64306]_ ;
  assign \new_[64311]_  = \new_[64310]_  & \new_[64303]_ ;
  assign \new_[64315]_  = ~A298 & A269;
  assign \new_[64316]_  = ~A268 & \new_[64315]_ ;
  assign \new_[64319]_  = ~A300 & A299;
  assign \new_[64322]_  = A302 & ~A301;
  assign \new_[64323]_  = \new_[64322]_  & \new_[64319]_ ;
  assign \new_[64324]_  = \new_[64323]_  & \new_[64316]_ ;
  assign \new_[64328]_  = A167 & A168;
  assign \new_[64329]_  = A170 & \new_[64328]_ ;
  assign \new_[64332]_  = A199 & ~A166;
  assign \new_[64335]_  = ~A265 & A200;
  assign \new_[64336]_  = \new_[64335]_  & \new_[64332]_ ;
  assign \new_[64337]_  = \new_[64336]_  & \new_[64329]_ ;
  assign \new_[64341]_  = ~A268 & ~A267;
  assign \new_[64342]_  = A266 & \new_[64341]_ ;
  assign \new_[64345]_  = A300 & A269;
  assign \new_[64348]_  = A302 & ~A301;
  assign \new_[64349]_  = \new_[64348]_  & \new_[64345]_ ;
  assign \new_[64350]_  = \new_[64349]_  & \new_[64342]_ ;
  assign \new_[64354]_  = A167 & A168;
  assign \new_[64355]_  = A170 & \new_[64354]_ ;
  assign \new_[64358]_  = A199 & ~A166;
  assign \new_[64361]_  = A265 & A200;
  assign \new_[64362]_  = \new_[64361]_  & \new_[64358]_ ;
  assign \new_[64363]_  = \new_[64362]_  & \new_[64355]_ ;
  assign \new_[64367]_  = ~A268 & ~A267;
  assign \new_[64368]_  = ~A266 & \new_[64367]_ ;
  assign \new_[64371]_  = A300 & A269;
  assign \new_[64374]_  = A302 & ~A301;
  assign \new_[64375]_  = \new_[64374]_  & \new_[64371]_ ;
  assign \new_[64376]_  = \new_[64375]_  & \new_[64368]_ ;
  assign \new_[64380]_  = A167 & A168;
  assign \new_[64381]_  = A170 & \new_[64380]_ ;
  assign \new_[64384]_  = ~A199 & ~A166;
  assign \new_[64387]_  = A267 & ~A200;
  assign \new_[64388]_  = \new_[64387]_  & \new_[64384]_ ;
  assign \new_[64389]_  = \new_[64388]_  & \new_[64381]_ ;
  assign \new_[64393]_  = A298 & A269;
  assign \new_[64394]_  = ~A268 & \new_[64393]_ ;
  assign \new_[64397]_  = ~A300 & ~A299;
  assign \new_[64400]_  = A302 & ~A301;
  assign \new_[64401]_  = \new_[64400]_  & \new_[64397]_ ;
  assign \new_[64402]_  = \new_[64401]_  & \new_[64394]_ ;
  assign \new_[64406]_  = A167 & A168;
  assign \new_[64407]_  = A170 & \new_[64406]_ ;
  assign \new_[64410]_  = ~A199 & ~A166;
  assign \new_[64413]_  = A267 & ~A200;
  assign \new_[64414]_  = \new_[64413]_  & \new_[64410]_ ;
  assign \new_[64415]_  = \new_[64414]_  & \new_[64407]_ ;
  assign \new_[64419]_  = ~A298 & A269;
  assign \new_[64420]_  = ~A268 & \new_[64419]_ ;
  assign \new_[64423]_  = ~A300 & A299;
  assign \new_[64426]_  = A302 & ~A301;
  assign \new_[64427]_  = \new_[64426]_  & \new_[64423]_ ;
  assign \new_[64428]_  = \new_[64427]_  & \new_[64420]_ ;
  assign \new_[64432]_  = A167 & A168;
  assign \new_[64433]_  = A170 & \new_[64432]_ ;
  assign \new_[64436]_  = ~A199 & ~A166;
  assign \new_[64439]_  = ~A265 & ~A200;
  assign \new_[64440]_  = \new_[64439]_  & \new_[64436]_ ;
  assign \new_[64441]_  = \new_[64440]_  & \new_[64433]_ ;
  assign \new_[64445]_  = ~A268 & ~A267;
  assign \new_[64446]_  = A266 & \new_[64445]_ ;
  assign \new_[64449]_  = A300 & A269;
  assign \new_[64452]_  = A302 & ~A301;
  assign \new_[64453]_  = \new_[64452]_  & \new_[64449]_ ;
  assign \new_[64454]_  = \new_[64453]_  & \new_[64446]_ ;
  assign \new_[64458]_  = A167 & A168;
  assign \new_[64459]_  = A170 & \new_[64458]_ ;
  assign \new_[64462]_  = ~A199 & ~A166;
  assign \new_[64465]_  = A265 & ~A200;
  assign \new_[64466]_  = \new_[64465]_  & \new_[64462]_ ;
  assign \new_[64467]_  = \new_[64466]_  & \new_[64459]_ ;
  assign \new_[64471]_  = ~A268 & ~A267;
  assign \new_[64472]_  = ~A266 & \new_[64471]_ ;
  assign \new_[64475]_  = A300 & A269;
  assign \new_[64478]_  = A302 & ~A301;
  assign \new_[64479]_  = \new_[64478]_  & \new_[64475]_ ;
  assign \new_[64480]_  = \new_[64479]_  & \new_[64472]_ ;
  assign \new_[64484]_  = ~A167 & A168;
  assign \new_[64485]_  = A170 & \new_[64484]_ ;
  assign \new_[64488]_  = A201 & A166;
  assign \new_[64491]_  = A203 & ~A202;
  assign \new_[64492]_  = \new_[64491]_  & \new_[64488]_ ;
  assign \new_[64493]_  = \new_[64492]_  & \new_[64485]_ ;
  assign \new_[64497]_  = A269 & ~A268;
  assign \new_[64498]_  = A267 & \new_[64497]_ ;
  assign \new_[64501]_  = ~A299 & A298;
  assign \new_[64504]_  = A301 & A300;
  assign \new_[64505]_  = \new_[64504]_  & \new_[64501]_ ;
  assign \new_[64506]_  = \new_[64505]_  & \new_[64498]_ ;
  assign \new_[64510]_  = ~A167 & A168;
  assign \new_[64511]_  = A170 & \new_[64510]_ ;
  assign \new_[64514]_  = A201 & A166;
  assign \new_[64517]_  = A203 & ~A202;
  assign \new_[64518]_  = \new_[64517]_  & \new_[64514]_ ;
  assign \new_[64519]_  = \new_[64518]_  & \new_[64511]_ ;
  assign \new_[64523]_  = A269 & ~A268;
  assign \new_[64524]_  = A267 & \new_[64523]_ ;
  assign \new_[64527]_  = ~A299 & A298;
  assign \new_[64530]_  = ~A302 & A300;
  assign \new_[64531]_  = \new_[64530]_  & \new_[64527]_ ;
  assign \new_[64532]_  = \new_[64531]_  & \new_[64524]_ ;
  assign \new_[64536]_  = ~A167 & A168;
  assign \new_[64537]_  = A170 & \new_[64536]_ ;
  assign \new_[64540]_  = A201 & A166;
  assign \new_[64543]_  = A203 & ~A202;
  assign \new_[64544]_  = \new_[64543]_  & \new_[64540]_ ;
  assign \new_[64545]_  = \new_[64544]_  & \new_[64537]_ ;
  assign \new_[64549]_  = A269 & ~A268;
  assign \new_[64550]_  = A267 & \new_[64549]_ ;
  assign \new_[64553]_  = A299 & ~A298;
  assign \new_[64556]_  = A301 & A300;
  assign \new_[64557]_  = \new_[64556]_  & \new_[64553]_ ;
  assign \new_[64558]_  = \new_[64557]_  & \new_[64550]_ ;
  assign \new_[64562]_  = ~A167 & A168;
  assign \new_[64563]_  = A170 & \new_[64562]_ ;
  assign \new_[64566]_  = A201 & A166;
  assign \new_[64569]_  = A203 & ~A202;
  assign \new_[64570]_  = \new_[64569]_  & \new_[64566]_ ;
  assign \new_[64571]_  = \new_[64570]_  & \new_[64563]_ ;
  assign \new_[64575]_  = A269 & ~A268;
  assign \new_[64576]_  = A267 & \new_[64575]_ ;
  assign \new_[64579]_  = A299 & ~A298;
  assign \new_[64582]_  = ~A302 & A300;
  assign \new_[64583]_  = \new_[64582]_  & \new_[64579]_ ;
  assign \new_[64584]_  = \new_[64583]_  & \new_[64576]_ ;
  assign \new_[64588]_  = ~A167 & A168;
  assign \new_[64589]_  = A170 & \new_[64588]_ ;
  assign \new_[64592]_  = A201 & A166;
  assign \new_[64595]_  = A203 & ~A202;
  assign \new_[64596]_  = \new_[64595]_  & \new_[64592]_ ;
  assign \new_[64597]_  = \new_[64596]_  & \new_[64589]_ ;
  assign \new_[64601]_  = A298 & A268;
  assign \new_[64602]_  = ~A267 & \new_[64601]_ ;
  assign \new_[64605]_  = ~A300 & ~A299;
  assign \new_[64608]_  = A302 & ~A301;
  assign \new_[64609]_  = \new_[64608]_  & \new_[64605]_ ;
  assign \new_[64610]_  = \new_[64609]_  & \new_[64602]_ ;
  assign \new_[64614]_  = ~A167 & A168;
  assign \new_[64615]_  = A170 & \new_[64614]_ ;
  assign \new_[64618]_  = A201 & A166;
  assign \new_[64621]_  = A203 & ~A202;
  assign \new_[64622]_  = \new_[64621]_  & \new_[64618]_ ;
  assign \new_[64623]_  = \new_[64622]_  & \new_[64615]_ ;
  assign \new_[64627]_  = ~A298 & A268;
  assign \new_[64628]_  = ~A267 & \new_[64627]_ ;
  assign \new_[64631]_  = ~A300 & A299;
  assign \new_[64634]_  = A302 & ~A301;
  assign \new_[64635]_  = \new_[64634]_  & \new_[64631]_ ;
  assign \new_[64636]_  = \new_[64635]_  & \new_[64628]_ ;
  assign \new_[64640]_  = ~A167 & A168;
  assign \new_[64641]_  = A170 & \new_[64640]_ ;
  assign \new_[64644]_  = A201 & A166;
  assign \new_[64647]_  = A203 & ~A202;
  assign \new_[64648]_  = \new_[64647]_  & \new_[64644]_ ;
  assign \new_[64649]_  = \new_[64648]_  & \new_[64641]_ ;
  assign \new_[64653]_  = A298 & ~A269;
  assign \new_[64654]_  = ~A267 & \new_[64653]_ ;
  assign \new_[64657]_  = ~A300 & ~A299;
  assign \new_[64660]_  = A302 & ~A301;
  assign \new_[64661]_  = \new_[64660]_  & \new_[64657]_ ;
  assign \new_[64662]_  = \new_[64661]_  & \new_[64654]_ ;
  assign \new_[64666]_  = ~A167 & A168;
  assign \new_[64667]_  = A170 & \new_[64666]_ ;
  assign \new_[64670]_  = A201 & A166;
  assign \new_[64673]_  = A203 & ~A202;
  assign \new_[64674]_  = \new_[64673]_  & \new_[64670]_ ;
  assign \new_[64675]_  = \new_[64674]_  & \new_[64667]_ ;
  assign \new_[64679]_  = ~A298 & ~A269;
  assign \new_[64680]_  = ~A267 & \new_[64679]_ ;
  assign \new_[64683]_  = ~A300 & A299;
  assign \new_[64686]_  = A302 & ~A301;
  assign \new_[64687]_  = \new_[64686]_  & \new_[64683]_ ;
  assign \new_[64688]_  = \new_[64687]_  & \new_[64680]_ ;
  assign \new_[64692]_  = ~A167 & A168;
  assign \new_[64693]_  = A170 & \new_[64692]_ ;
  assign \new_[64696]_  = A201 & A166;
  assign \new_[64699]_  = A203 & ~A202;
  assign \new_[64700]_  = \new_[64699]_  & \new_[64696]_ ;
  assign \new_[64701]_  = \new_[64700]_  & \new_[64693]_ ;
  assign \new_[64705]_  = A298 & A266;
  assign \new_[64706]_  = A265 & \new_[64705]_ ;
  assign \new_[64709]_  = ~A300 & ~A299;
  assign \new_[64712]_  = A302 & ~A301;
  assign \new_[64713]_  = \new_[64712]_  & \new_[64709]_ ;
  assign \new_[64714]_  = \new_[64713]_  & \new_[64706]_ ;
  assign \new_[64718]_  = ~A167 & A168;
  assign \new_[64719]_  = A170 & \new_[64718]_ ;
  assign \new_[64722]_  = A201 & A166;
  assign \new_[64725]_  = A203 & ~A202;
  assign \new_[64726]_  = \new_[64725]_  & \new_[64722]_ ;
  assign \new_[64727]_  = \new_[64726]_  & \new_[64719]_ ;
  assign \new_[64731]_  = ~A298 & A266;
  assign \new_[64732]_  = A265 & \new_[64731]_ ;
  assign \new_[64735]_  = ~A300 & A299;
  assign \new_[64738]_  = A302 & ~A301;
  assign \new_[64739]_  = \new_[64738]_  & \new_[64735]_ ;
  assign \new_[64740]_  = \new_[64739]_  & \new_[64732]_ ;
  assign \new_[64744]_  = ~A167 & A168;
  assign \new_[64745]_  = A170 & \new_[64744]_ ;
  assign \new_[64748]_  = A201 & A166;
  assign \new_[64751]_  = A203 & ~A202;
  assign \new_[64752]_  = \new_[64751]_  & \new_[64748]_ ;
  assign \new_[64753]_  = \new_[64752]_  & \new_[64745]_ ;
  assign \new_[64757]_  = A267 & A266;
  assign \new_[64758]_  = ~A265 & \new_[64757]_ ;
  assign \new_[64761]_  = A300 & A268;
  assign \new_[64764]_  = A302 & ~A301;
  assign \new_[64765]_  = \new_[64764]_  & \new_[64761]_ ;
  assign \new_[64766]_  = \new_[64765]_  & \new_[64758]_ ;
  assign \new_[64770]_  = ~A167 & A168;
  assign \new_[64771]_  = A170 & \new_[64770]_ ;
  assign \new_[64774]_  = A201 & A166;
  assign \new_[64777]_  = A203 & ~A202;
  assign \new_[64778]_  = \new_[64777]_  & \new_[64774]_ ;
  assign \new_[64779]_  = \new_[64778]_  & \new_[64771]_ ;
  assign \new_[64783]_  = A267 & A266;
  assign \new_[64784]_  = ~A265 & \new_[64783]_ ;
  assign \new_[64787]_  = A300 & ~A269;
  assign \new_[64790]_  = A302 & ~A301;
  assign \new_[64791]_  = \new_[64790]_  & \new_[64787]_ ;
  assign \new_[64792]_  = \new_[64791]_  & \new_[64784]_ ;
  assign \new_[64796]_  = ~A167 & A168;
  assign \new_[64797]_  = A170 & \new_[64796]_ ;
  assign \new_[64800]_  = A201 & A166;
  assign \new_[64803]_  = A203 & ~A202;
  assign \new_[64804]_  = \new_[64803]_  & \new_[64800]_ ;
  assign \new_[64805]_  = \new_[64804]_  & \new_[64797]_ ;
  assign \new_[64809]_  = ~A267 & A266;
  assign \new_[64810]_  = ~A265 & \new_[64809]_ ;
  assign \new_[64813]_  = A269 & ~A268;
  assign \new_[64816]_  = A301 & ~A300;
  assign \new_[64817]_  = \new_[64816]_  & \new_[64813]_ ;
  assign \new_[64818]_  = \new_[64817]_  & \new_[64810]_ ;
  assign \new_[64822]_  = ~A167 & A168;
  assign \new_[64823]_  = A170 & \new_[64822]_ ;
  assign \new_[64826]_  = A201 & A166;
  assign \new_[64829]_  = A203 & ~A202;
  assign \new_[64830]_  = \new_[64829]_  & \new_[64826]_ ;
  assign \new_[64831]_  = \new_[64830]_  & \new_[64823]_ ;
  assign \new_[64835]_  = ~A267 & A266;
  assign \new_[64836]_  = ~A265 & \new_[64835]_ ;
  assign \new_[64839]_  = A269 & ~A268;
  assign \new_[64842]_  = ~A302 & ~A300;
  assign \new_[64843]_  = \new_[64842]_  & \new_[64839]_ ;
  assign \new_[64844]_  = \new_[64843]_  & \new_[64836]_ ;
  assign \new_[64848]_  = ~A167 & A168;
  assign \new_[64849]_  = A170 & \new_[64848]_ ;
  assign \new_[64852]_  = A201 & A166;
  assign \new_[64855]_  = A203 & ~A202;
  assign \new_[64856]_  = \new_[64855]_  & \new_[64852]_ ;
  assign \new_[64857]_  = \new_[64856]_  & \new_[64849]_ ;
  assign \new_[64861]_  = ~A267 & A266;
  assign \new_[64862]_  = ~A265 & \new_[64861]_ ;
  assign \new_[64865]_  = A269 & ~A268;
  assign \new_[64868]_  = A299 & A298;
  assign \new_[64869]_  = \new_[64868]_  & \new_[64865]_ ;
  assign \new_[64870]_  = \new_[64869]_  & \new_[64862]_ ;
  assign \new_[64874]_  = ~A167 & A168;
  assign \new_[64875]_  = A170 & \new_[64874]_ ;
  assign \new_[64878]_  = A201 & A166;
  assign \new_[64881]_  = A203 & ~A202;
  assign \new_[64882]_  = \new_[64881]_  & \new_[64878]_ ;
  assign \new_[64883]_  = \new_[64882]_  & \new_[64875]_ ;
  assign \new_[64887]_  = ~A267 & A266;
  assign \new_[64888]_  = ~A265 & \new_[64887]_ ;
  assign \new_[64891]_  = A269 & ~A268;
  assign \new_[64894]_  = ~A299 & ~A298;
  assign \new_[64895]_  = \new_[64894]_  & \new_[64891]_ ;
  assign \new_[64896]_  = \new_[64895]_  & \new_[64888]_ ;
  assign \new_[64900]_  = ~A167 & A168;
  assign \new_[64901]_  = A170 & \new_[64900]_ ;
  assign \new_[64904]_  = A201 & A166;
  assign \new_[64907]_  = A203 & ~A202;
  assign \new_[64908]_  = \new_[64907]_  & \new_[64904]_ ;
  assign \new_[64909]_  = \new_[64908]_  & \new_[64901]_ ;
  assign \new_[64913]_  = A267 & ~A266;
  assign \new_[64914]_  = A265 & \new_[64913]_ ;
  assign \new_[64917]_  = A300 & A268;
  assign \new_[64920]_  = A302 & ~A301;
  assign \new_[64921]_  = \new_[64920]_  & \new_[64917]_ ;
  assign \new_[64922]_  = \new_[64921]_  & \new_[64914]_ ;
  assign \new_[64926]_  = ~A167 & A168;
  assign \new_[64927]_  = A170 & \new_[64926]_ ;
  assign \new_[64930]_  = A201 & A166;
  assign \new_[64933]_  = A203 & ~A202;
  assign \new_[64934]_  = \new_[64933]_  & \new_[64930]_ ;
  assign \new_[64935]_  = \new_[64934]_  & \new_[64927]_ ;
  assign \new_[64939]_  = A267 & ~A266;
  assign \new_[64940]_  = A265 & \new_[64939]_ ;
  assign \new_[64943]_  = A300 & ~A269;
  assign \new_[64946]_  = A302 & ~A301;
  assign \new_[64947]_  = \new_[64946]_  & \new_[64943]_ ;
  assign \new_[64948]_  = \new_[64947]_  & \new_[64940]_ ;
  assign \new_[64952]_  = ~A167 & A168;
  assign \new_[64953]_  = A170 & \new_[64952]_ ;
  assign \new_[64956]_  = A201 & A166;
  assign \new_[64959]_  = A203 & ~A202;
  assign \new_[64960]_  = \new_[64959]_  & \new_[64956]_ ;
  assign \new_[64961]_  = \new_[64960]_  & \new_[64953]_ ;
  assign \new_[64965]_  = ~A267 & ~A266;
  assign \new_[64966]_  = A265 & \new_[64965]_ ;
  assign \new_[64969]_  = A269 & ~A268;
  assign \new_[64972]_  = A301 & ~A300;
  assign \new_[64973]_  = \new_[64972]_  & \new_[64969]_ ;
  assign \new_[64974]_  = \new_[64973]_  & \new_[64966]_ ;
  assign \new_[64978]_  = ~A167 & A168;
  assign \new_[64979]_  = A170 & \new_[64978]_ ;
  assign \new_[64982]_  = A201 & A166;
  assign \new_[64985]_  = A203 & ~A202;
  assign \new_[64986]_  = \new_[64985]_  & \new_[64982]_ ;
  assign \new_[64987]_  = \new_[64986]_  & \new_[64979]_ ;
  assign \new_[64991]_  = ~A267 & ~A266;
  assign \new_[64992]_  = A265 & \new_[64991]_ ;
  assign \new_[64995]_  = A269 & ~A268;
  assign \new_[64998]_  = ~A302 & ~A300;
  assign \new_[64999]_  = \new_[64998]_  & \new_[64995]_ ;
  assign \new_[65000]_  = \new_[64999]_  & \new_[64992]_ ;
  assign \new_[65004]_  = ~A167 & A168;
  assign \new_[65005]_  = A170 & \new_[65004]_ ;
  assign \new_[65008]_  = A201 & A166;
  assign \new_[65011]_  = A203 & ~A202;
  assign \new_[65012]_  = \new_[65011]_  & \new_[65008]_ ;
  assign \new_[65013]_  = \new_[65012]_  & \new_[65005]_ ;
  assign \new_[65017]_  = ~A267 & ~A266;
  assign \new_[65018]_  = A265 & \new_[65017]_ ;
  assign \new_[65021]_  = A269 & ~A268;
  assign \new_[65024]_  = A299 & A298;
  assign \new_[65025]_  = \new_[65024]_  & \new_[65021]_ ;
  assign \new_[65026]_  = \new_[65025]_  & \new_[65018]_ ;
  assign \new_[65030]_  = ~A167 & A168;
  assign \new_[65031]_  = A170 & \new_[65030]_ ;
  assign \new_[65034]_  = A201 & A166;
  assign \new_[65037]_  = A203 & ~A202;
  assign \new_[65038]_  = \new_[65037]_  & \new_[65034]_ ;
  assign \new_[65039]_  = \new_[65038]_  & \new_[65031]_ ;
  assign \new_[65043]_  = ~A267 & ~A266;
  assign \new_[65044]_  = A265 & \new_[65043]_ ;
  assign \new_[65047]_  = A269 & ~A268;
  assign \new_[65050]_  = ~A299 & ~A298;
  assign \new_[65051]_  = \new_[65050]_  & \new_[65047]_ ;
  assign \new_[65052]_  = \new_[65051]_  & \new_[65044]_ ;
  assign \new_[65056]_  = ~A167 & A168;
  assign \new_[65057]_  = A170 & \new_[65056]_ ;
  assign \new_[65060]_  = A201 & A166;
  assign \new_[65063]_  = A203 & ~A202;
  assign \new_[65064]_  = \new_[65063]_  & \new_[65060]_ ;
  assign \new_[65065]_  = \new_[65064]_  & \new_[65057]_ ;
  assign \new_[65069]_  = A298 & ~A266;
  assign \new_[65070]_  = ~A265 & \new_[65069]_ ;
  assign \new_[65073]_  = ~A300 & ~A299;
  assign \new_[65076]_  = A302 & ~A301;
  assign \new_[65077]_  = \new_[65076]_  & \new_[65073]_ ;
  assign \new_[65078]_  = \new_[65077]_  & \new_[65070]_ ;
  assign \new_[65082]_  = ~A167 & A168;
  assign \new_[65083]_  = A170 & \new_[65082]_ ;
  assign \new_[65086]_  = A201 & A166;
  assign \new_[65089]_  = A203 & ~A202;
  assign \new_[65090]_  = \new_[65089]_  & \new_[65086]_ ;
  assign \new_[65091]_  = \new_[65090]_  & \new_[65083]_ ;
  assign \new_[65095]_  = ~A298 & ~A266;
  assign \new_[65096]_  = ~A265 & \new_[65095]_ ;
  assign \new_[65099]_  = ~A300 & A299;
  assign \new_[65102]_  = A302 & ~A301;
  assign \new_[65103]_  = \new_[65102]_  & \new_[65099]_ ;
  assign \new_[65104]_  = \new_[65103]_  & \new_[65096]_ ;
  assign \new_[65108]_  = ~A167 & A168;
  assign \new_[65109]_  = A170 & \new_[65108]_ ;
  assign \new_[65112]_  = ~A201 & A166;
  assign \new_[65115]_  = A267 & A202;
  assign \new_[65116]_  = \new_[65115]_  & \new_[65112]_ ;
  assign \new_[65117]_  = \new_[65116]_  & \new_[65109]_ ;
  assign \new_[65121]_  = A298 & A269;
  assign \new_[65122]_  = ~A268 & \new_[65121]_ ;
  assign \new_[65125]_  = ~A300 & ~A299;
  assign \new_[65128]_  = A302 & ~A301;
  assign \new_[65129]_  = \new_[65128]_  & \new_[65125]_ ;
  assign \new_[65130]_  = \new_[65129]_  & \new_[65122]_ ;
  assign \new_[65134]_  = ~A167 & A168;
  assign \new_[65135]_  = A170 & \new_[65134]_ ;
  assign \new_[65138]_  = ~A201 & A166;
  assign \new_[65141]_  = A267 & A202;
  assign \new_[65142]_  = \new_[65141]_  & \new_[65138]_ ;
  assign \new_[65143]_  = \new_[65142]_  & \new_[65135]_ ;
  assign \new_[65147]_  = ~A298 & A269;
  assign \new_[65148]_  = ~A268 & \new_[65147]_ ;
  assign \new_[65151]_  = ~A300 & A299;
  assign \new_[65154]_  = A302 & ~A301;
  assign \new_[65155]_  = \new_[65154]_  & \new_[65151]_ ;
  assign \new_[65156]_  = \new_[65155]_  & \new_[65148]_ ;
  assign \new_[65160]_  = ~A167 & A168;
  assign \new_[65161]_  = A170 & \new_[65160]_ ;
  assign \new_[65164]_  = ~A201 & A166;
  assign \new_[65167]_  = ~A265 & A202;
  assign \new_[65168]_  = \new_[65167]_  & \new_[65164]_ ;
  assign \new_[65169]_  = \new_[65168]_  & \new_[65161]_ ;
  assign \new_[65173]_  = ~A268 & ~A267;
  assign \new_[65174]_  = A266 & \new_[65173]_ ;
  assign \new_[65177]_  = A300 & A269;
  assign \new_[65180]_  = A302 & ~A301;
  assign \new_[65181]_  = \new_[65180]_  & \new_[65177]_ ;
  assign \new_[65182]_  = \new_[65181]_  & \new_[65174]_ ;
  assign \new_[65186]_  = ~A167 & A168;
  assign \new_[65187]_  = A170 & \new_[65186]_ ;
  assign \new_[65190]_  = ~A201 & A166;
  assign \new_[65193]_  = A265 & A202;
  assign \new_[65194]_  = \new_[65193]_  & \new_[65190]_ ;
  assign \new_[65195]_  = \new_[65194]_  & \new_[65187]_ ;
  assign \new_[65199]_  = ~A268 & ~A267;
  assign \new_[65200]_  = ~A266 & \new_[65199]_ ;
  assign \new_[65203]_  = A300 & A269;
  assign \new_[65206]_  = A302 & ~A301;
  assign \new_[65207]_  = \new_[65206]_  & \new_[65203]_ ;
  assign \new_[65208]_  = \new_[65207]_  & \new_[65200]_ ;
  assign \new_[65212]_  = ~A167 & A168;
  assign \new_[65213]_  = A170 & \new_[65212]_ ;
  assign \new_[65216]_  = ~A201 & A166;
  assign \new_[65219]_  = A267 & ~A203;
  assign \new_[65220]_  = \new_[65219]_  & \new_[65216]_ ;
  assign \new_[65221]_  = \new_[65220]_  & \new_[65213]_ ;
  assign \new_[65225]_  = A298 & A269;
  assign \new_[65226]_  = ~A268 & \new_[65225]_ ;
  assign \new_[65229]_  = ~A300 & ~A299;
  assign \new_[65232]_  = A302 & ~A301;
  assign \new_[65233]_  = \new_[65232]_  & \new_[65229]_ ;
  assign \new_[65234]_  = \new_[65233]_  & \new_[65226]_ ;
  assign \new_[65238]_  = ~A167 & A168;
  assign \new_[65239]_  = A170 & \new_[65238]_ ;
  assign \new_[65242]_  = ~A201 & A166;
  assign \new_[65245]_  = A267 & ~A203;
  assign \new_[65246]_  = \new_[65245]_  & \new_[65242]_ ;
  assign \new_[65247]_  = \new_[65246]_  & \new_[65239]_ ;
  assign \new_[65251]_  = ~A298 & A269;
  assign \new_[65252]_  = ~A268 & \new_[65251]_ ;
  assign \new_[65255]_  = ~A300 & A299;
  assign \new_[65258]_  = A302 & ~A301;
  assign \new_[65259]_  = \new_[65258]_  & \new_[65255]_ ;
  assign \new_[65260]_  = \new_[65259]_  & \new_[65252]_ ;
  assign \new_[65264]_  = ~A167 & A168;
  assign \new_[65265]_  = A170 & \new_[65264]_ ;
  assign \new_[65268]_  = ~A201 & A166;
  assign \new_[65271]_  = ~A265 & ~A203;
  assign \new_[65272]_  = \new_[65271]_  & \new_[65268]_ ;
  assign \new_[65273]_  = \new_[65272]_  & \new_[65265]_ ;
  assign \new_[65277]_  = ~A268 & ~A267;
  assign \new_[65278]_  = A266 & \new_[65277]_ ;
  assign \new_[65281]_  = A300 & A269;
  assign \new_[65284]_  = A302 & ~A301;
  assign \new_[65285]_  = \new_[65284]_  & \new_[65281]_ ;
  assign \new_[65286]_  = \new_[65285]_  & \new_[65278]_ ;
  assign \new_[65290]_  = ~A167 & A168;
  assign \new_[65291]_  = A170 & \new_[65290]_ ;
  assign \new_[65294]_  = ~A201 & A166;
  assign \new_[65297]_  = A265 & ~A203;
  assign \new_[65298]_  = \new_[65297]_  & \new_[65294]_ ;
  assign \new_[65299]_  = \new_[65298]_  & \new_[65291]_ ;
  assign \new_[65303]_  = ~A268 & ~A267;
  assign \new_[65304]_  = ~A266 & \new_[65303]_ ;
  assign \new_[65307]_  = A300 & A269;
  assign \new_[65310]_  = A302 & ~A301;
  assign \new_[65311]_  = \new_[65310]_  & \new_[65307]_ ;
  assign \new_[65312]_  = \new_[65311]_  & \new_[65304]_ ;
  assign \new_[65316]_  = ~A167 & A168;
  assign \new_[65317]_  = A170 & \new_[65316]_ ;
  assign \new_[65320]_  = A199 & A166;
  assign \new_[65323]_  = A267 & A200;
  assign \new_[65324]_  = \new_[65323]_  & \new_[65320]_ ;
  assign \new_[65325]_  = \new_[65324]_  & \new_[65317]_ ;
  assign \new_[65329]_  = A298 & A269;
  assign \new_[65330]_  = ~A268 & \new_[65329]_ ;
  assign \new_[65333]_  = ~A300 & ~A299;
  assign \new_[65336]_  = A302 & ~A301;
  assign \new_[65337]_  = \new_[65336]_  & \new_[65333]_ ;
  assign \new_[65338]_  = \new_[65337]_  & \new_[65330]_ ;
  assign \new_[65342]_  = ~A167 & A168;
  assign \new_[65343]_  = A170 & \new_[65342]_ ;
  assign \new_[65346]_  = A199 & A166;
  assign \new_[65349]_  = A267 & A200;
  assign \new_[65350]_  = \new_[65349]_  & \new_[65346]_ ;
  assign \new_[65351]_  = \new_[65350]_  & \new_[65343]_ ;
  assign \new_[65355]_  = ~A298 & A269;
  assign \new_[65356]_  = ~A268 & \new_[65355]_ ;
  assign \new_[65359]_  = ~A300 & A299;
  assign \new_[65362]_  = A302 & ~A301;
  assign \new_[65363]_  = \new_[65362]_  & \new_[65359]_ ;
  assign \new_[65364]_  = \new_[65363]_  & \new_[65356]_ ;
  assign \new_[65368]_  = ~A167 & A168;
  assign \new_[65369]_  = A170 & \new_[65368]_ ;
  assign \new_[65372]_  = A199 & A166;
  assign \new_[65375]_  = ~A265 & A200;
  assign \new_[65376]_  = \new_[65375]_  & \new_[65372]_ ;
  assign \new_[65377]_  = \new_[65376]_  & \new_[65369]_ ;
  assign \new_[65381]_  = ~A268 & ~A267;
  assign \new_[65382]_  = A266 & \new_[65381]_ ;
  assign \new_[65385]_  = A300 & A269;
  assign \new_[65388]_  = A302 & ~A301;
  assign \new_[65389]_  = \new_[65388]_  & \new_[65385]_ ;
  assign \new_[65390]_  = \new_[65389]_  & \new_[65382]_ ;
  assign \new_[65394]_  = ~A167 & A168;
  assign \new_[65395]_  = A170 & \new_[65394]_ ;
  assign \new_[65398]_  = A199 & A166;
  assign \new_[65401]_  = A265 & A200;
  assign \new_[65402]_  = \new_[65401]_  & \new_[65398]_ ;
  assign \new_[65403]_  = \new_[65402]_  & \new_[65395]_ ;
  assign \new_[65407]_  = ~A268 & ~A267;
  assign \new_[65408]_  = ~A266 & \new_[65407]_ ;
  assign \new_[65411]_  = A300 & A269;
  assign \new_[65414]_  = A302 & ~A301;
  assign \new_[65415]_  = \new_[65414]_  & \new_[65411]_ ;
  assign \new_[65416]_  = \new_[65415]_  & \new_[65408]_ ;
  assign \new_[65420]_  = ~A167 & A168;
  assign \new_[65421]_  = A170 & \new_[65420]_ ;
  assign \new_[65424]_  = ~A199 & A166;
  assign \new_[65427]_  = A267 & ~A200;
  assign \new_[65428]_  = \new_[65427]_  & \new_[65424]_ ;
  assign \new_[65429]_  = \new_[65428]_  & \new_[65421]_ ;
  assign \new_[65433]_  = A298 & A269;
  assign \new_[65434]_  = ~A268 & \new_[65433]_ ;
  assign \new_[65437]_  = ~A300 & ~A299;
  assign \new_[65440]_  = A302 & ~A301;
  assign \new_[65441]_  = \new_[65440]_  & \new_[65437]_ ;
  assign \new_[65442]_  = \new_[65441]_  & \new_[65434]_ ;
  assign \new_[65446]_  = ~A167 & A168;
  assign \new_[65447]_  = A170 & \new_[65446]_ ;
  assign \new_[65450]_  = ~A199 & A166;
  assign \new_[65453]_  = A267 & ~A200;
  assign \new_[65454]_  = \new_[65453]_  & \new_[65450]_ ;
  assign \new_[65455]_  = \new_[65454]_  & \new_[65447]_ ;
  assign \new_[65459]_  = ~A298 & A269;
  assign \new_[65460]_  = ~A268 & \new_[65459]_ ;
  assign \new_[65463]_  = ~A300 & A299;
  assign \new_[65466]_  = A302 & ~A301;
  assign \new_[65467]_  = \new_[65466]_  & \new_[65463]_ ;
  assign \new_[65468]_  = \new_[65467]_  & \new_[65460]_ ;
  assign \new_[65472]_  = ~A167 & A168;
  assign \new_[65473]_  = A170 & \new_[65472]_ ;
  assign \new_[65476]_  = ~A199 & A166;
  assign \new_[65479]_  = ~A265 & ~A200;
  assign \new_[65480]_  = \new_[65479]_  & \new_[65476]_ ;
  assign \new_[65481]_  = \new_[65480]_  & \new_[65473]_ ;
  assign \new_[65485]_  = ~A268 & ~A267;
  assign \new_[65486]_  = A266 & \new_[65485]_ ;
  assign \new_[65489]_  = A300 & A269;
  assign \new_[65492]_  = A302 & ~A301;
  assign \new_[65493]_  = \new_[65492]_  & \new_[65489]_ ;
  assign \new_[65494]_  = \new_[65493]_  & \new_[65486]_ ;
  assign \new_[65498]_  = ~A167 & A168;
  assign \new_[65499]_  = A170 & \new_[65498]_ ;
  assign \new_[65502]_  = ~A199 & A166;
  assign \new_[65505]_  = A265 & ~A200;
  assign \new_[65506]_  = \new_[65505]_  & \new_[65502]_ ;
  assign \new_[65507]_  = \new_[65506]_  & \new_[65499]_ ;
  assign \new_[65511]_  = ~A268 & ~A267;
  assign \new_[65512]_  = ~A266 & \new_[65511]_ ;
  assign \new_[65515]_  = A300 & A269;
  assign \new_[65518]_  = A302 & ~A301;
  assign \new_[65519]_  = \new_[65518]_  & \new_[65515]_ ;
  assign \new_[65520]_  = \new_[65519]_  & \new_[65512]_ ;
  assign \new_[65524]_  = ~A199 & ~A168;
  assign \new_[65525]_  = A170 & \new_[65524]_ ;
  assign \new_[65528]_  = A201 & A200;
  assign \new_[65531]_  = ~A265 & A202;
  assign \new_[65532]_  = \new_[65531]_  & \new_[65528]_ ;
  assign \new_[65533]_  = \new_[65532]_  & \new_[65525]_ ;
  assign \new_[65537]_  = A268 & A267;
  assign \new_[65538]_  = A266 & \new_[65537]_ ;
  assign \new_[65541]_  = ~A299 & A298;
  assign \new_[65544]_  = A301 & A300;
  assign \new_[65545]_  = \new_[65544]_  & \new_[65541]_ ;
  assign \new_[65546]_  = \new_[65545]_  & \new_[65538]_ ;
  assign \new_[65550]_  = ~A199 & ~A168;
  assign \new_[65551]_  = A170 & \new_[65550]_ ;
  assign \new_[65554]_  = A201 & A200;
  assign \new_[65557]_  = ~A265 & A202;
  assign \new_[65558]_  = \new_[65557]_  & \new_[65554]_ ;
  assign \new_[65559]_  = \new_[65558]_  & \new_[65551]_ ;
  assign \new_[65563]_  = A268 & A267;
  assign \new_[65564]_  = A266 & \new_[65563]_ ;
  assign \new_[65567]_  = ~A299 & A298;
  assign \new_[65570]_  = ~A302 & A300;
  assign \new_[65571]_  = \new_[65570]_  & \new_[65567]_ ;
  assign \new_[65572]_  = \new_[65571]_  & \new_[65564]_ ;
  assign \new_[65576]_  = ~A199 & ~A168;
  assign \new_[65577]_  = A170 & \new_[65576]_ ;
  assign \new_[65580]_  = A201 & A200;
  assign \new_[65583]_  = ~A265 & A202;
  assign \new_[65584]_  = \new_[65583]_  & \new_[65580]_ ;
  assign \new_[65585]_  = \new_[65584]_  & \new_[65577]_ ;
  assign \new_[65589]_  = A268 & A267;
  assign \new_[65590]_  = A266 & \new_[65589]_ ;
  assign \new_[65593]_  = A299 & ~A298;
  assign \new_[65596]_  = A301 & A300;
  assign \new_[65597]_  = \new_[65596]_  & \new_[65593]_ ;
  assign \new_[65598]_  = \new_[65597]_  & \new_[65590]_ ;
  assign \new_[65602]_  = ~A199 & ~A168;
  assign \new_[65603]_  = A170 & \new_[65602]_ ;
  assign \new_[65606]_  = A201 & A200;
  assign \new_[65609]_  = ~A265 & A202;
  assign \new_[65610]_  = \new_[65609]_  & \new_[65606]_ ;
  assign \new_[65611]_  = \new_[65610]_  & \new_[65603]_ ;
  assign \new_[65615]_  = A268 & A267;
  assign \new_[65616]_  = A266 & \new_[65615]_ ;
  assign \new_[65619]_  = A299 & ~A298;
  assign \new_[65622]_  = ~A302 & A300;
  assign \new_[65623]_  = \new_[65622]_  & \new_[65619]_ ;
  assign \new_[65624]_  = \new_[65623]_  & \new_[65616]_ ;
  assign \new_[65628]_  = ~A199 & ~A168;
  assign \new_[65629]_  = A170 & \new_[65628]_ ;
  assign \new_[65632]_  = A201 & A200;
  assign \new_[65635]_  = ~A265 & A202;
  assign \new_[65636]_  = \new_[65635]_  & \new_[65632]_ ;
  assign \new_[65637]_  = \new_[65636]_  & \new_[65629]_ ;
  assign \new_[65641]_  = ~A269 & A267;
  assign \new_[65642]_  = A266 & \new_[65641]_ ;
  assign \new_[65645]_  = ~A299 & A298;
  assign \new_[65648]_  = A301 & A300;
  assign \new_[65649]_  = \new_[65648]_  & \new_[65645]_ ;
  assign \new_[65650]_  = \new_[65649]_  & \new_[65642]_ ;
  assign \new_[65654]_  = ~A199 & ~A168;
  assign \new_[65655]_  = A170 & \new_[65654]_ ;
  assign \new_[65658]_  = A201 & A200;
  assign \new_[65661]_  = ~A265 & A202;
  assign \new_[65662]_  = \new_[65661]_  & \new_[65658]_ ;
  assign \new_[65663]_  = \new_[65662]_  & \new_[65655]_ ;
  assign \new_[65667]_  = ~A269 & A267;
  assign \new_[65668]_  = A266 & \new_[65667]_ ;
  assign \new_[65671]_  = ~A299 & A298;
  assign \new_[65674]_  = ~A302 & A300;
  assign \new_[65675]_  = \new_[65674]_  & \new_[65671]_ ;
  assign \new_[65676]_  = \new_[65675]_  & \new_[65668]_ ;
  assign \new_[65680]_  = ~A199 & ~A168;
  assign \new_[65681]_  = A170 & \new_[65680]_ ;
  assign \new_[65684]_  = A201 & A200;
  assign \new_[65687]_  = ~A265 & A202;
  assign \new_[65688]_  = \new_[65687]_  & \new_[65684]_ ;
  assign \new_[65689]_  = \new_[65688]_  & \new_[65681]_ ;
  assign \new_[65693]_  = ~A269 & A267;
  assign \new_[65694]_  = A266 & \new_[65693]_ ;
  assign \new_[65697]_  = A299 & ~A298;
  assign \new_[65700]_  = A301 & A300;
  assign \new_[65701]_  = \new_[65700]_  & \new_[65697]_ ;
  assign \new_[65702]_  = \new_[65701]_  & \new_[65694]_ ;
  assign \new_[65706]_  = ~A199 & ~A168;
  assign \new_[65707]_  = A170 & \new_[65706]_ ;
  assign \new_[65710]_  = A201 & A200;
  assign \new_[65713]_  = ~A265 & A202;
  assign \new_[65714]_  = \new_[65713]_  & \new_[65710]_ ;
  assign \new_[65715]_  = \new_[65714]_  & \new_[65707]_ ;
  assign \new_[65719]_  = ~A269 & A267;
  assign \new_[65720]_  = A266 & \new_[65719]_ ;
  assign \new_[65723]_  = A299 & ~A298;
  assign \new_[65726]_  = ~A302 & A300;
  assign \new_[65727]_  = \new_[65726]_  & \new_[65723]_ ;
  assign \new_[65728]_  = \new_[65727]_  & \new_[65720]_ ;
  assign \new_[65732]_  = ~A199 & ~A168;
  assign \new_[65733]_  = A170 & \new_[65732]_ ;
  assign \new_[65736]_  = A201 & A200;
  assign \new_[65739]_  = A265 & A202;
  assign \new_[65740]_  = \new_[65739]_  & \new_[65736]_ ;
  assign \new_[65741]_  = \new_[65740]_  & \new_[65733]_ ;
  assign \new_[65745]_  = A268 & A267;
  assign \new_[65746]_  = ~A266 & \new_[65745]_ ;
  assign \new_[65749]_  = ~A299 & A298;
  assign \new_[65752]_  = A301 & A300;
  assign \new_[65753]_  = \new_[65752]_  & \new_[65749]_ ;
  assign \new_[65754]_  = \new_[65753]_  & \new_[65746]_ ;
  assign \new_[65758]_  = ~A199 & ~A168;
  assign \new_[65759]_  = A170 & \new_[65758]_ ;
  assign \new_[65762]_  = A201 & A200;
  assign \new_[65765]_  = A265 & A202;
  assign \new_[65766]_  = \new_[65765]_  & \new_[65762]_ ;
  assign \new_[65767]_  = \new_[65766]_  & \new_[65759]_ ;
  assign \new_[65771]_  = A268 & A267;
  assign \new_[65772]_  = ~A266 & \new_[65771]_ ;
  assign \new_[65775]_  = ~A299 & A298;
  assign \new_[65778]_  = ~A302 & A300;
  assign \new_[65779]_  = \new_[65778]_  & \new_[65775]_ ;
  assign \new_[65780]_  = \new_[65779]_  & \new_[65772]_ ;
  assign \new_[65784]_  = ~A199 & ~A168;
  assign \new_[65785]_  = A170 & \new_[65784]_ ;
  assign \new_[65788]_  = A201 & A200;
  assign \new_[65791]_  = A265 & A202;
  assign \new_[65792]_  = \new_[65791]_  & \new_[65788]_ ;
  assign \new_[65793]_  = \new_[65792]_  & \new_[65785]_ ;
  assign \new_[65797]_  = A268 & A267;
  assign \new_[65798]_  = ~A266 & \new_[65797]_ ;
  assign \new_[65801]_  = A299 & ~A298;
  assign \new_[65804]_  = A301 & A300;
  assign \new_[65805]_  = \new_[65804]_  & \new_[65801]_ ;
  assign \new_[65806]_  = \new_[65805]_  & \new_[65798]_ ;
  assign \new_[65810]_  = ~A199 & ~A168;
  assign \new_[65811]_  = A170 & \new_[65810]_ ;
  assign \new_[65814]_  = A201 & A200;
  assign \new_[65817]_  = A265 & A202;
  assign \new_[65818]_  = \new_[65817]_  & \new_[65814]_ ;
  assign \new_[65819]_  = \new_[65818]_  & \new_[65811]_ ;
  assign \new_[65823]_  = A268 & A267;
  assign \new_[65824]_  = ~A266 & \new_[65823]_ ;
  assign \new_[65827]_  = A299 & ~A298;
  assign \new_[65830]_  = ~A302 & A300;
  assign \new_[65831]_  = \new_[65830]_  & \new_[65827]_ ;
  assign \new_[65832]_  = \new_[65831]_  & \new_[65824]_ ;
  assign \new_[65836]_  = ~A199 & ~A168;
  assign \new_[65837]_  = A170 & \new_[65836]_ ;
  assign \new_[65840]_  = A201 & A200;
  assign \new_[65843]_  = A265 & A202;
  assign \new_[65844]_  = \new_[65843]_  & \new_[65840]_ ;
  assign \new_[65845]_  = \new_[65844]_  & \new_[65837]_ ;
  assign \new_[65849]_  = ~A269 & A267;
  assign \new_[65850]_  = ~A266 & \new_[65849]_ ;
  assign \new_[65853]_  = ~A299 & A298;
  assign \new_[65856]_  = A301 & A300;
  assign \new_[65857]_  = \new_[65856]_  & \new_[65853]_ ;
  assign \new_[65858]_  = \new_[65857]_  & \new_[65850]_ ;
  assign \new_[65862]_  = ~A199 & ~A168;
  assign \new_[65863]_  = A170 & \new_[65862]_ ;
  assign \new_[65866]_  = A201 & A200;
  assign \new_[65869]_  = A265 & A202;
  assign \new_[65870]_  = \new_[65869]_  & \new_[65866]_ ;
  assign \new_[65871]_  = \new_[65870]_  & \new_[65863]_ ;
  assign \new_[65875]_  = ~A269 & A267;
  assign \new_[65876]_  = ~A266 & \new_[65875]_ ;
  assign \new_[65879]_  = ~A299 & A298;
  assign \new_[65882]_  = ~A302 & A300;
  assign \new_[65883]_  = \new_[65882]_  & \new_[65879]_ ;
  assign \new_[65884]_  = \new_[65883]_  & \new_[65876]_ ;
  assign \new_[65888]_  = ~A199 & ~A168;
  assign \new_[65889]_  = A170 & \new_[65888]_ ;
  assign \new_[65892]_  = A201 & A200;
  assign \new_[65895]_  = A265 & A202;
  assign \new_[65896]_  = \new_[65895]_  & \new_[65892]_ ;
  assign \new_[65897]_  = \new_[65896]_  & \new_[65889]_ ;
  assign \new_[65901]_  = ~A269 & A267;
  assign \new_[65902]_  = ~A266 & \new_[65901]_ ;
  assign \new_[65905]_  = A299 & ~A298;
  assign \new_[65908]_  = A301 & A300;
  assign \new_[65909]_  = \new_[65908]_  & \new_[65905]_ ;
  assign \new_[65910]_  = \new_[65909]_  & \new_[65902]_ ;
  assign \new_[65914]_  = ~A199 & ~A168;
  assign \new_[65915]_  = A170 & \new_[65914]_ ;
  assign \new_[65918]_  = A201 & A200;
  assign \new_[65921]_  = A265 & A202;
  assign \new_[65922]_  = \new_[65921]_  & \new_[65918]_ ;
  assign \new_[65923]_  = \new_[65922]_  & \new_[65915]_ ;
  assign \new_[65927]_  = ~A269 & A267;
  assign \new_[65928]_  = ~A266 & \new_[65927]_ ;
  assign \new_[65931]_  = A299 & ~A298;
  assign \new_[65934]_  = ~A302 & A300;
  assign \new_[65935]_  = \new_[65934]_  & \new_[65931]_ ;
  assign \new_[65936]_  = \new_[65935]_  & \new_[65928]_ ;
  assign \new_[65940]_  = ~A199 & ~A168;
  assign \new_[65941]_  = A170 & \new_[65940]_ ;
  assign \new_[65944]_  = A201 & A200;
  assign \new_[65947]_  = ~A265 & ~A203;
  assign \new_[65948]_  = \new_[65947]_  & \new_[65944]_ ;
  assign \new_[65949]_  = \new_[65948]_  & \new_[65941]_ ;
  assign \new_[65953]_  = A268 & A267;
  assign \new_[65954]_  = A266 & \new_[65953]_ ;
  assign \new_[65957]_  = ~A299 & A298;
  assign \new_[65960]_  = A301 & A300;
  assign \new_[65961]_  = \new_[65960]_  & \new_[65957]_ ;
  assign \new_[65962]_  = \new_[65961]_  & \new_[65954]_ ;
  assign \new_[65966]_  = ~A199 & ~A168;
  assign \new_[65967]_  = A170 & \new_[65966]_ ;
  assign \new_[65970]_  = A201 & A200;
  assign \new_[65973]_  = ~A265 & ~A203;
  assign \new_[65974]_  = \new_[65973]_  & \new_[65970]_ ;
  assign \new_[65975]_  = \new_[65974]_  & \new_[65967]_ ;
  assign \new_[65979]_  = A268 & A267;
  assign \new_[65980]_  = A266 & \new_[65979]_ ;
  assign \new_[65983]_  = ~A299 & A298;
  assign \new_[65986]_  = ~A302 & A300;
  assign \new_[65987]_  = \new_[65986]_  & \new_[65983]_ ;
  assign \new_[65988]_  = \new_[65987]_  & \new_[65980]_ ;
  assign \new_[65992]_  = ~A199 & ~A168;
  assign \new_[65993]_  = A170 & \new_[65992]_ ;
  assign \new_[65996]_  = A201 & A200;
  assign \new_[65999]_  = ~A265 & ~A203;
  assign \new_[66000]_  = \new_[65999]_  & \new_[65996]_ ;
  assign \new_[66001]_  = \new_[66000]_  & \new_[65993]_ ;
  assign \new_[66005]_  = A268 & A267;
  assign \new_[66006]_  = A266 & \new_[66005]_ ;
  assign \new_[66009]_  = A299 & ~A298;
  assign \new_[66012]_  = A301 & A300;
  assign \new_[66013]_  = \new_[66012]_  & \new_[66009]_ ;
  assign \new_[66014]_  = \new_[66013]_  & \new_[66006]_ ;
  assign \new_[66018]_  = ~A199 & ~A168;
  assign \new_[66019]_  = A170 & \new_[66018]_ ;
  assign \new_[66022]_  = A201 & A200;
  assign \new_[66025]_  = ~A265 & ~A203;
  assign \new_[66026]_  = \new_[66025]_  & \new_[66022]_ ;
  assign \new_[66027]_  = \new_[66026]_  & \new_[66019]_ ;
  assign \new_[66031]_  = A268 & A267;
  assign \new_[66032]_  = A266 & \new_[66031]_ ;
  assign \new_[66035]_  = A299 & ~A298;
  assign \new_[66038]_  = ~A302 & A300;
  assign \new_[66039]_  = \new_[66038]_  & \new_[66035]_ ;
  assign \new_[66040]_  = \new_[66039]_  & \new_[66032]_ ;
  assign \new_[66044]_  = ~A199 & ~A168;
  assign \new_[66045]_  = A170 & \new_[66044]_ ;
  assign \new_[66048]_  = A201 & A200;
  assign \new_[66051]_  = ~A265 & ~A203;
  assign \new_[66052]_  = \new_[66051]_  & \new_[66048]_ ;
  assign \new_[66053]_  = \new_[66052]_  & \new_[66045]_ ;
  assign \new_[66057]_  = ~A269 & A267;
  assign \new_[66058]_  = A266 & \new_[66057]_ ;
  assign \new_[66061]_  = ~A299 & A298;
  assign \new_[66064]_  = A301 & A300;
  assign \new_[66065]_  = \new_[66064]_  & \new_[66061]_ ;
  assign \new_[66066]_  = \new_[66065]_  & \new_[66058]_ ;
  assign \new_[66070]_  = ~A199 & ~A168;
  assign \new_[66071]_  = A170 & \new_[66070]_ ;
  assign \new_[66074]_  = A201 & A200;
  assign \new_[66077]_  = ~A265 & ~A203;
  assign \new_[66078]_  = \new_[66077]_  & \new_[66074]_ ;
  assign \new_[66079]_  = \new_[66078]_  & \new_[66071]_ ;
  assign \new_[66083]_  = ~A269 & A267;
  assign \new_[66084]_  = A266 & \new_[66083]_ ;
  assign \new_[66087]_  = ~A299 & A298;
  assign \new_[66090]_  = ~A302 & A300;
  assign \new_[66091]_  = \new_[66090]_  & \new_[66087]_ ;
  assign \new_[66092]_  = \new_[66091]_  & \new_[66084]_ ;
  assign \new_[66096]_  = ~A199 & ~A168;
  assign \new_[66097]_  = A170 & \new_[66096]_ ;
  assign \new_[66100]_  = A201 & A200;
  assign \new_[66103]_  = ~A265 & ~A203;
  assign \new_[66104]_  = \new_[66103]_  & \new_[66100]_ ;
  assign \new_[66105]_  = \new_[66104]_  & \new_[66097]_ ;
  assign \new_[66109]_  = ~A269 & A267;
  assign \new_[66110]_  = A266 & \new_[66109]_ ;
  assign \new_[66113]_  = A299 & ~A298;
  assign \new_[66116]_  = A301 & A300;
  assign \new_[66117]_  = \new_[66116]_  & \new_[66113]_ ;
  assign \new_[66118]_  = \new_[66117]_  & \new_[66110]_ ;
  assign \new_[66122]_  = ~A199 & ~A168;
  assign \new_[66123]_  = A170 & \new_[66122]_ ;
  assign \new_[66126]_  = A201 & A200;
  assign \new_[66129]_  = ~A265 & ~A203;
  assign \new_[66130]_  = \new_[66129]_  & \new_[66126]_ ;
  assign \new_[66131]_  = \new_[66130]_  & \new_[66123]_ ;
  assign \new_[66135]_  = ~A269 & A267;
  assign \new_[66136]_  = A266 & \new_[66135]_ ;
  assign \new_[66139]_  = A299 & ~A298;
  assign \new_[66142]_  = ~A302 & A300;
  assign \new_[66143]_  = \new_[66142]_  & \new_[66139]_ ;
  assign \new_[66144]_  = \new_[66143]_  & \new_[66136]_ ;
  assign \new_[66148]_  = ~A199 & ~A168;
  assign \new_[66149]_  = A170 & \new_[66148]_ ;
  assign \new_[66152]_  = A201 & A200;
  assign \new_[66155]_  = A265 & ~A203;
  assign \new_[66156]_  = \new_[66155]_  & \new_[66152]_ ;
  assign \new_[66157]_  = \new_[66156]_  & \new_[66149]_ ;
  assign \new_[66161]_  = A268 & A267;
  assign \new_[66162]_  = ~A266 & \new_[66161]_ ;
  assign \new_[66165]_  = ~A299 & A298;
  assign \new_[66168]_  = A301 & A300;
  assign \new_[66169]_  = \new_[66168]_  & \new_[66165]_ ;
  assign \new_[66170]_  = \new_[66169]_  & \new_[66162]_ ;
  assign \new_[66174]_  = ~A199 & ~A168;
  assign \new_[66175]_  = A170 & \new_[66174]_ ;
  assign \new_[66178]_  = A201 & A200;
  assign \new_[66181]_  = A265 & ~A203;
  assign \new_[66182]_  = \new_[66181]_  & \new_[66178]_ ;
  assign \new_[66183]_  = \new_[66182]_  & \new_[66175]_ ;
  assign \new_[66187]_  = A268 & A267;
  assign \new_[66188]_  = ~A266 & \new_[66187]_ ;
  assign \new_[66191]_  = ~A299 & A298;
  assign \new_[66194]_  = ~A302 & A300;
  assign \new_[66195]_  = \new_[66194]_  & \new_[66191]_ ;
  assign \new_[66196]_  = \new_[66195]_  & \new_[66188]_ ;
  assign \new_[66200]_  = ~A199 & ~A168;
  assign \new_[66201]_  = A170 & \new_[66200]_ ;
  assign \new_[66204]_  = A201 & A200;
  assign \new_[66207]_  = A265 & ~A203;
  assign \new_[66208]_  = \new_[66207]_  & \new_[66204]_ ;
  assign \new_[66209]_  = \new_[66208]_  & \new_[66201]_ ;
  assign \new_[66213]_  = A268 & A267;
  assign \new_[66214]_  = ~A266 & \new_[66213]_ ;
  assign \new_[66217]_  = A299 & ~A298;
  assign \new_[66220]_  = A301 & A300;
  assign \new_[66221]_  = \new_[66220]_  & \new_[66217]_ ;
  assign \new_[66222]_  = \new_[66221]_  & \new_[66214]_ ;
  assign \new_[66226]_  = ~A199 & ~A168;
  assign \new_[66227]_  = A170 & \new_[66226]_ ;
  assign \new_[66230]_  = A201 & A200;
  assign \new_[66233]_  = A265 & ~A203;
  assign \new_[66234]_  = \new_[66233]_  & \new_[66230]_ ;
  assign \new_[66235]_  = \new_[66234]_  & \new_[66227]_ ;
  assign \new_[66239]_  = A268 & A267;
  assign \new_[66240]_  = ~A266 & \new_[66239]_ ;
  assign \new_[66243]_  = A299 & ~A298;
  assign \new_[66246]_  = ~A302 & A300;
  assign \new_[66247]_  = \new_[66246]_  & \new_[66243]_ ;
  assign \new_[66248]_  = \new_[66247]_  & \new_[66240]_ ;
  assign \new_[66252]_  = ~A199 & ~A168;
  assign \new_[66253]_  = A170 & \new_[66252]_ ;
  assign \new_[66256]_  = A201 & A200;
  assign \new_[66259]_  = A265 & ~A203;
  assign \new_[66260]_  = \new_[66259]_  & \new_[66256]_ ;
  assign \new_[66261]_  = \new_[66260]_  & \new_[66253]_ ;
  assign \new_[66265]_  = ~A269 & A267;
  assign \new_[66266]_  = ~A266 & \new_[66265]_ ;
  assign \new_[66269]_  = ~A299 & A298;
  assign \new_[66272]_  = A301 & A300;
  assign \new_[66273]_  = \new_[66272]_  & \new_[66269]_ ;
  assign \new_[66274]_  = \new_[66273]_  & \new_[66266]_ ;
  assign \new_[66278]_  = ~A199 & ~A168;
  assign \new_[66279]_  = A170 & \new_[66278]_ ;
  assign \new_[66282]_  = A201 & A200;
  assign \new_[66285]_  = A265 & ~A203;
  assign \new_[66286]_  = \new_[66285]_  & \new_[66282]_ ;
  assign \new_[66287]_  = \new_[66286]_  & \new_[66279]_ ;
  assign \new_[66291]_  = ~A269 & A267;
  assign \new_[66292]_  = ~A266 & \new_[66291]_ ;
  assign \new_[66295]_  = ~A299 & A298;
  assign \new_[66298]_  = ~A302 & A300;
  assign \new_[66299]_  = \new_[66298]_  & \new_[66295]_ ;
  assign \new_[66300]_  = \new_[66299]_  & \new_[66292]_ ;
  assign \new_[66304]_  = ~A199 & ~A168;
  assign \new_[66305]_  = A170 & \new_[66304]_ ;
  assign \new_[66308]_  = A201 & A200;
  assign \new_[66311]_  = A265 & ~A203;
  assign \new_[66312]_  = \new_[66311]_  & \new_[66308]_ ;
  assign \new_[66313]_  = \new_[66312]_  & \new_[66305]_ ;
  assign \new_[66317]_  = ~A269 & A267;
  assign \new_[66318]_  = ~A266 & \new_[66317]_ ;
  assign \new_[66321]_  = A299 & ~A298;
  assign \new_[66324]_  = A301 & A300;
  assign \new_[66325]_  = \new_[66324]_  & \new_[66321]_ ;
  assign \new_[66326]_  = \new_[66325]_  & \new_[66318]_ ;
  assign \new_[66330]_  = ~A199 & ~A168;
  assign \new_[66331]_  = A170 & \new_[66330]_ ;
  assign \new_[66334]_  = A201 & A200;
  assign \new_[66337]_  = A265 & ~A203;
  assign \new_[66338]_  = \new_[66337]_  & \new_[66334]_ ;
  assign \new_[66339]_  = \new_[66338]_  & \new_[66331]_ ;
  assign \new_[66343]_  = ~A269 & A267;
  assign \new_[66344]_  = ~A266 & \new_[66343]_ ;
  assign \new_[66347]_  = A299 & ~A298;
  assign \new_[66350]_  = ~A302 & A300;
  assign \new_[66351]_  = \new_[66350]_  & \new_[66347]_ ;
  assign \new_[66352]_  = \new_[66351]_  & \new_[66344]_ ;
  assign \new_[66356]_  = A199 & ~A168;
  assign \new_[66357]_  = A170 & \new_[66356]_ ;
  assign \new_[66360]_  = A201 & ~A200;
  assign \new_[66363]_  = ~A265 & A202;
  assign \new_[66364]_  = \new_[66363]_  & \new_[66360]_ ;
  assign \new_[66365]_  = \new_[66364]_  & \new_[66357]_ ;
  assign \new_[66369]_  = A268 & A267;
  assign \new_[66370]_  = A266 & \new_[66369]_ ;
  assign \new_[66373]_  = ~A299 & A298;
  assign \new_[66376]_  = A301 & A300;
  assign \new_[66377]_  = \new_[66376]_  & \new_[66373]_ ;
  assign \new_[66378]_  = \new_[66377]_  & \new_[66370]_ ;
  assign \new_[66382]_  = A199 & ~A168;
  assign \new_[66383]_  = A170 & \new_[66382]_ ;
  assign \new_[66386]_  = A201 & ~A200;
  assign \new_[66389]_  = ~A265 & A202;
  assign \new_[66390]_  = \new_[66389]_  & \new_[66386]_ ;
  assign \new_[66391]_  = \new_[66390]_  & \new_[66383]_ ;
  assign \new_[66395]_  = A268 & A267;
  assign \new_[66396]_  = A266 & \new_[66395]_ ;
  assign \new_[66399]_  = ~A299 & A298;
  assign \new_[66402]_  = ~A302 & A300;
  assign \new_[66403]_  = \new_[66402]_  & \new_[66399]_ ;
  assign \new_[66404]_  = \new_[66403]_  & \new_[66396]_ ;
  assign \new_[66408]_  = A199 & ~A168;
  assign \new_[66409]_  = A170 & \new_[66408]_ ;
  assign \new_[66412]_  = A201 & ~A200;
  assign \new_[66415]_  = ~A265 & A202;
  assign \new_[66416]_  = \new_[66415]_  & \new_[66412]_ ;
  assign \new_[66417]_  = \new_[66416]_  & \new_[66409]_ ;
  assign \new_[66421]_  = A268 & A267;
  assign \new_[66422]_  = A266 & \new_[66421]_ ;
  assign \new_[66425]_  = A299 & ~A298;
  assign \new_[66428]_  = A301 & A300;
  assign \new_[66429]_  = \new_[66428]_  & \new_[66425]_ ;
  assign \new_[66430]_  = \new_[66429]_  & \new_[66422]_ ;
  assign \new_[66434]_  = A199 & ~A168;
  assign \new_[66435]_  = A170 & \new_[66434]_ ;
  assign \new_[66438]_  = A201 & ~A200;
  assign \new_[66441]_  = ~A265 & A202;
  assign \new_[66442]_  = \new_[66441]_  & \new_[66438]_ ;
  assign \new_[66443]_  = \new_[66442]_  & \new_[66435]_ ;
  assign \new_[66447]_  = A268 & A267;
  assign \new_[66448]_  = A266 & \new_[66447]_ ;
  assign \new_[66451]_  = A299 & ~A298;
  assign \new_[66454]_  = ~A302 & A300;
  assign \new_[66455]_  = \new_[66454]_  & \new_[66451]_ ;
  assign \new_[66456]_  = \new_[66455]_  & \new_[66448]_ ;
  assign \new_[66460]_  = A199 & ~A168;
  assign \new_[66461]_  = A170 & \new_[66460]_ ;
  assign \new_[66464]_  = A201 & ~A200;
  assign \new_[66467]_  = ~A265 & A202;
  assign \new_[66468]_  = \new_[66467]_  & \new_[66464]_ ;
  assign \new_[66469]_  = \new_[66468]_  & \new_[66461]_ ;
  assign \new_[66473]_  = ~A269 & A267;
  assign \new_[66474]_  = A266 & \new_[66473]_ ;
  assign \new_[66477]_  = ~A299 & A298;
  assign \new_[66480]_  = A301 & A300;
  assign \new_[66481]_  = \new_[66480]_  & \new_[66477]_ ;
  assign \new_[66482]_  = \new_[66481]_  & \new_[66474]_ ;
  assign \new_[66486]_  = A199 & ~A168;
  assign \new_[66487]_  = A170 & \new_[66486]_ ;
  assign \new_[66490]_  = A201 & ~A200;
  assign \new_[66493]_  = ~A265 & A202;
  assign \new_[66494]_  = \new_[66493]_  & \new_[66490]_ ;
  assign \new_[66495]_  = \new_[66494]_  & \new_[66487]_ ;
  assign \new_[66499]_  = ~A269 & A267;
  assign \new_[66500]_  = A266 & \new_[66499]_ ;
  assign \new_[66503]_  = ~A299 & A298;
  assign \new_[66506]_  = ~A302 & A300;
  assign \new_[66507]_  = \new_[66506]_  & \new_[66503]_ ;
  assign \new_[66508]_  = \new_[66507]_  & \new_[66500]_ ;
  assign \new_[66512]_  = A199 & ~A168;
  assign \new_[66513]_  = A170 & \new_[66512]_ ;
  assign \new_[66516]_  = A201 & ~A200;
  assign \new_[66519]_  = ~A265 & A202;
  assign \new_[66520]_  = \new_[66519]_  & \new_[66516]_ ;
  assign \new_[66521]_  = \new_[66520]_  & \new_[66513]_ ;
  assign \new_[66525]_  = ~A269 & A267;
  assign \new_[66526]_  = A266 & \new_[66525]_ ;
  assign \new_[66529]_  = A299 & ~A298;
  assign \new_[66532]_  = A301 & A300;
  assign \new_[66533]_  = \new_[66532]_  & \new_[66529]_ ;
  assign \new_[66534]_  = \new_[66533]_  & \new_[66526]_ ;
  assign \new_[66538]_  = A199 & ~A168;
  assign \new_[66539]_  = A170 & \new_[66538]_ ;
  assign \new_[66542]_  = A201 & ~A200;
  assign \new_[66545]_  = ~A265 & A202;
  assign \new_[66546]_  = \new_[66545]_  & \new_[66542]_ ;
  assign \new_[66547]_  = \new_[66546]_  & \new_[66539]_ ;
  assign \new_[66551]_  = ~A269 & A267;
  assign \new_[66552]_  = A266 & \new_[66551]_ ;
  assign \new_[66555]_  = A299 & ~A298;
  assign \new_[66558]_  = ~A302 & A300;
  assign \new_[66559]_  = \new_[66558]_  & \new_[66555]_ ;
  assign \new_[66560]_  = \new_[66559]_  & \new_[66552]_ ;
  assign \new_[66564]_  = A199 & ~A168;
  assign \new_[66565]_  = A170 & \new_[66564]_ ;
  assign \new_[66568]_  = A201 & ~A200;
  assign \new_[66571]_  = A265 & A202;
  assign \new_[66572]_  = \new_[66571]_  & \new_[66568]_ ;
  assign \new_[66573]_  = \new_[66572]_  & \new_[66565]_ ;
  assign \new_[66577]_  = A268 & A267;
  assign \new_[66578]_  = ~A266 & \new_[66577]_ ;
  assign \new_[66581]_  = ~A299 & A298;
  assign \new_[66584]_  = A301 & A300;
  assign \new_[66585]_  = \new_[66584]_  & \new_[66581]_ ;
  assign \new_[66586]_  = \new_[66585]_  & \new_[66578]_ ;
  assign \new_[66590]_  = A199 & ~A168;
  assign \new_[66591]_  = A170 & \new_[66590]_ ;
  assign \new_[66594]_  = A201 & ~A200;
  assign \new_[66597]_  = A265 & A202;
  assign \new_[66598]_  = \new_[66597]_  & \new_[66594]_ ;
  assign \new_[66599]_  = \new_[66598]_  & \new_[66591]_ ;
  assign \new_[66603]_  = A268 & A267;
  assign \new_[66604]_  = ~A266 & \new_[66603]_ ;
  assign \new_[66607]_  = ~A299 & A298;
  assign \new_[66610]_  = ~A302 & A300;
  assign \new_[66611]_  = \new_[66610]_  & \new_[66607]_ ;
  assign \new_[66612]_  = \new_[66611]_  & \new_[66604]_ ;
  assign \new_[66616]_  = A199 & ~A168;
  assign \new_[66617]_  = A170 & \new_[66616]_ ;
  assign \new_[66620]_  = A201 & ~A200;
  assign \new_[66623]_  = A265 & A202;
  assign \new_[66624]_  = \new_[66623]_  & \new_[66620]_ ;
  assign \new_[66625]_  = \new_[66624]_  & \new_[66617]_ ;
  assign \new_[66629]_  = A268 & A267;
  assign \new_[66630]_  = ~A266 & \new_[66629]_ ;
  assign \new_[66633]_  = A299 & ~A298;
  assign \new_[66636]_  = A301 & A300;
  assign \new_[66637]_  = \new_[66636]_  & \new_[66633]_ ;
  assign \new_[66638]_  = \new_[66637]_  & \new_[66630]_ ;
  assign \new_[66642]_  = A199 & ~A168;
  assign \new_[66643]_  = A170 & \new_[66642]_ ;
  assign \new_[66646]_  = A201 & ~A200;
  assign \new_[66649]_  = A265 & A202;
  assign \new_[66650]_  = \new_[66649]_  & \new_[66646]_ ;
  assign \new_[66651]_  = \new_[66650]_  & \new_[66643]_ ;
  assign \new_[66655]_  = A268 & A267;
  assign \new_[66656]_  = ~A266 & \new_[66655]_ ;
  assign \new_[66659]_  = A299 & ~A298;
  assign \new_[66662]_  = ~A302 & A300;
  assign \new_[66663]_  = \new_[66662]_  & \new_[66659]_ ;
  assign \new_[66664]_  = \new_[66663]_  & \new_[66656]_ ;
  assign \new_[66668]_  = A199 & ~A168;
  assign \new_[66669]_  = A170 & \new_[66668]_ ;
  assign \new_[66672]_  = A201 & ~A200;
  assign \new_[66675]_  = A265 & A202;
  assign \new_[66676]_  = \new_[66675]_  & \new_[66672]_ ;
  assign \new_[66677]_  = \new_[66676]_  & \new_[66669]_ ;
  assign \new_[66681]_  = ~A269 & A267;
  assign \new_[66682]_  = ~A266 & \new_[66681]_ ;
  assign \new_[66685]_  = ~A299 & A298;
  assign \new_[66688]_  = A301 & A300;
  assign \new_[66689]_  = \new_[66688]_  & \new_[66685]_ ;
  assign \new_[66690]_  = \new_[66689]_  & \new_[66682]_ ;
  assign \new_[66694]_  = A199 & ~A168;
  assign \new_[66695]_  = A170 & \new_[66694]_ ;
  assign \new_[66698]_  = A201 & ~A200;
  assign \new_[66701]_  = A265 & A202;
  assign \new_[66702]_  = \new_[66701]_  & \new_[66698]_ ;
  assign \new_[66703]_  = \new_[66702]_  & \new_[66695]_ ;
  assign \new_[66707]_  = ~A269 & A267;
  assign \new_[66708]_  = ~A266 & \new_[66707]_ ;
  assign \new_[66711]_  = ~A299 & A298;
  assign \new_[66714]_  = ~A302 & A300;
  assign \new_[66715]_  = \new_[66714]_  & \new_[66711]_ ;
  assign \new_[66716]_  = \new_[66715]_  & \new_[66708]_ ;
  assign \new_[66720]_  = A199 & ~A168;
  assign \new_[66721]_  = A170 & \new_[66720]_ ;
  assign \new_[66724]_  = A201 & ~A200;
  assign \new_[66727]_  = A265 & A202;
  assign \new_[66728]_  = \new_[66727]_  & \new_[66724]_ ;
  assign \new_[66729]_  = \new_[66728]_  & \new_[66721]_ ;
  assign \new_[66733]_  = ~A269 & A267;
  assign \new_[66734]_  = ~A266 & \new_[66733]_ ;
  assign \new_[66737]_  = A299 & ~A298;
  assign \new_[66740]_  = A301 & A300;
  assign \new_[66741]_  = \new_[66740]_  & \new_[66737]_ ;
  assign \new_[66742]_  = \new_[66741]_  & \new_[66734]_ ;
  assign \new_[66746]_  = A199 & ~A168;
  assign \new_[66747]_  = A170 & \new_[66746]_ ;
  assign \new_[66750]_  = A201 & ~A200;
  assign \new_[66753]_  = A265 & A202;
  assign \new_[66754]_  = \new_[66753]_  & \new_[66750]_ ;
  assign \new_[66755]_  = \new_[66754]_  & \new_[66747]_ ;
  assign \new_[66759]_  = ~A269 & A267;
  assign \new_[66760]_  = ~A266 & \new_[66759]_ ;
  assign \new_[66763]_  = A299 & ~A298;
  assign \new_[66766]_  = ~A302 & A300;
  assign \new_[66767]_  = \new_[66766]_  & \new_[66763]_ ;
  assign \new_[66768]_  = \new_[66767]_  & \new_[66760]_ ;
  assign \new_[66772]_  = A199 & ~A168;
  assign \new_[66773]_  = A170 & \new_[66772]_ ;
  assign \new_[66776]_  = A201 & ~A200;
  assign \new_[66779]_  = ~A265 & ~A203;
  assign \new_[66780]_  = \new_[66779]_  & \new_[66776]_ ;
  assign \new_[66781]_  = \new_[66780]_  & \new_[66773]_ ;
  assign \new_[66785]_  = A268 & A267;
  assign \new_[66786]_  = A266 & \new_[66785]_ ;
  assign \new_[66789]_  = ~A299 & A298;
  assign \new_[66792]_  = A301 & A300;
  assign \new_[66793]_  = \new_[66792]_  & \new_[66789]_ ;
  assign \new_[66794]_  = \new_[66793]_  & \new_[66786]_ ;
  assign \new_[66798]_  = A199 & ~A168;
  assign \new_[66799]_  = A170 & \new_[66798]_ ;
  assign \new_[66802]_  = A201 & ~A200;
  assign \new_[66805]_  = ~A265 & ~A203;
  assign \new_[66806]_  = \new_[66805]_  & \new_[66802]_ ;
  assign \new_[66807]_  = \new_[66806]_  & \new_[66799]_ ;
  assign \new_[66811]_  = A268 & A267;
  assign \new_[66812]_  = A266 & \new_[66811]_ ;
  assign \new_[66815]_  = ~A299 & A298;
  assign \new_[66818]_  = ~A302 & A300;
  assign \new_[66819]_  = \new_[66818]_  & \new_[66815]_ ;
  assign \new_[66820]_  = \new_[66819]_  & \new_[66812]_ ;
  assign \new_[66824]_  = A199 & ~A168;
  assign \new_[66825]_  = A170 & \new_[66824]_ ;
  assign \new_[66828]_  = A201 & ~A200;
  assign \new_[66831]_  = ~A265 & ~A203;
  assign \new_[66832]_  = \new_[66831]_  & \new_[66828]_ ;
  assign \new_[66833]_  = \new_[66832]_  & \new_[66825]_ ;
  assign \new_[66837]_  = A268 & A267;
  assign \new_[66838]_  = A266 & \new_[66837]_ ;
  assign \new_[66841]_  = A299 & ~A298;
  assign \new_[66844]_  = A301 & A300;
  assign \new_[66845]_  = \new_[66844]_  & \new_[66841]_ ;
  assign \new_[66846]_  = \new_[66845]_  & \new_[66838]_ ;
  assign \new_[66850]_  = A199 & ~A168;
  assign \new_[66851]_  = A170 & \new_[66850]_ ;
  assign \new_[66854]_  = A201 & ~A200;
  assign \new_[66857]_  = ~A265 & ~A203;
  assign \new_[66858]_  = \new_[66857]_  & \new_[66854]_ ;
  assign \new_[66859]_  = \new_[66858]_  & \new_[66851]_ ;
  assign \new_[66863]_  = A268 & A267;
  assign \new_[66864]_  = A266 & \new_[66863]_ ;
  assign \new_[66867]_  = A299 & ~A298;
  assign \new_[66870]_  = ~A302 & A300;
  assign \new_[66871]_  = \new_[66870]_  & \new_[66867]_ ;
  assign \new_[66872]_  = \new_[66871]_  & \new_[66864]_ ;
  assign \new_[66876]_  = A199 & ~A168;
  assign \new_[66877]_  = A170 & \new_[66876]_ ;
  assign \new_[66880]_  = A201 & ~A200;
  assign \new_[66883]_  = ~A265 & ~A203;
  assign \new_[66884]_  = \new_[66883]_  & \new_[66880]_ ;
  assign \new_[66885]_  = \new_[66884]_  & \new_[66877]_ ;
  assign \new_[66889]_  = ~A269 & A267;
  assign \new_[66890]_  = A266 & \new_[66889]_ ;
  assign \new_[66893]_  = ~A299 & A298;
  assign \new_[66896]_  = A301 & A300;
  assign \new_[66897]_  = \new_[66896]_  & \new_[66893]_ ;
  assign \new_[66898]_  = \new_[66897]_  & \new_[66890]_ ;
  assign \new_[66902]_  = A199 & ~A168;
  assign \new_[66903]_  = A170 & \new_[66902]_ ;
  assign \new_[66906]_  = A201 & ~A200;
  assign \new_[66909]_  = ~A265 & ~A203;
  assign \new_[66910]_  = \new_[66909]_  & \new_[66906]_ ;
  assign \new_[66911]_  = \new_[66910]_  & \new_[66903]_ ;
  assign \new_[66915]_  = ~A269 & A267;
  assign \new_[66916]_  = A266 & \new_[66915]_ ;
  assign \new_[66919]_  = ~A299 & A298;
  assign \new_[66922]_  = ~A302 & A300;
  assign \new_[66923]_  = \new_[66922]_  & \new_[66919]_ ;
  assign \new_[66924]_  = \new_[66923]_  & \new_[66916]_ ;
  assign \new_[66928]_  = A199 & ~A168;
  assign \new_[66929]_  = A170 & \new_[66928]_ ;
  assign \new_[66932]_  = A201 & ~A200;
  assign \new_[66935]_  = ~A265 & ~A203;
  assign \new_[66936]_  = \new_[66935]_  & \new_[66932]_ ;
  assign \new_[66937]_  = \new_[66936]_  & \new_[66929]_ ;
  assign \new_[66941]_  = ~A269 & A267;
  assign \new_[66942]_  = A266 & \new_[66941]_ ;
  assign \new_[66945]_  = A299 & ~A298;
  assign \new_[66948]_  = A301 & A300;
  assign \new_[66949]_  = \new_[66948]_  & \new_[66945]_ ;
  assign \new_[66950]_  = \new_[66949]_  & \new_[66942]_ ;
  assign \new_[66954]_  = A199 & ~A168;
  assign \new_[66955]_  = A170 & \new_[66954]_ ;
  assign \new_[66958]_  = A201 & ~A200;
  assign \new_[66961]_  = ~A265 & ~A203;
  assign \new_[66962]_  = \new_[66961]_  & \new_[66958]_ ;
  assign \new_[66963]_  = \new_[66962]_  & \new_[66955]_ ;
  assign \new_[66967]_  = ~A269 & A267;
  assign \new_[66968]_  = A266 & \new_[66967]_ ;
  assign \new_[66971]_  = A299 & ~A298;
  assign \new_[66974]_  = ~A302 & A300;
  assign \new_[66975]_  = \new_[66974]_  & \new_[66971]_ ;
  assign \new_[66976]_  = \new_[66975]_  & \new_[66968]_ ;
  assign \new_[66980]_  = A199 & ~A168;
  assign \new_[66981]_  = A170 & \new_[66980]_ ;
  assign \new_[66984]_  = A201 & ~A200;
  assign \new_[66987]_  = A265 & ~A203;
  assign \new_[66988]_  = \new_[66987]_  & \new_[66984]_ ;
  assign \new_[66989]_  = \new_[66988]_  & \new_[66981]_ ;
  assign \new_[66993]_  = A268 & A267;
  assign \new_[66994]_  = ~A266 & \new_[66993]_ ;
  assign \new_[66997]_  = ~A299 & A298;
  assign \new_[67000]_  = A301 & A300;
  assign \new_[67001]_  = \new_[67000]_  & \new_[66997]_ ;
  assign \new_[67002]_  = \new_[67001]_  & \new_[66994]_ ;
  assign \new_[67006]_  = A199 & ~A168;
  assign \new_[67007]_  = A170 & \new_[67006]_ ;
  assign \new_[67010]_  = A201 & ~A200;
  assign \new_[67013]_  = A265 & ~A203;
  assign \new_[67014]_  = \new_[67013]_  & \new_[67010]_ ;
  assign \new_[67015]_  = \new_[67014]_  & \new_[67007]_ ;
  assign \new_[67019]_  = A268 & A267;
  assign \new_[67020]_  = ~A266 & \new_[67019]_ ;
  assign \new_[67023]_  = ~A299 & A298;
  assign \new_[67026]_  = ~A302 & A300;
  assign \new_[67027]_  = \new_[67026]_  & \new_[67023]_ ;
  assign \new_[67028]_  = \new_[67027]_  & \new_[67020]_ ;
  assign \new_[67032]_  = A199 & ~A168;
  assign \new_[67033]_  = A170 & \new_[67032]_ ;
  assign \new_[67036]_  = A201 & ~A200;
  assign \new_[67039]_  = A265 & ~A203;
  assign \new_[67040]_  = \new_[67039]_  & \new_[67036]_ ;
  assign \new_[67041]_  = \new_[67040]_  & \new_[67033]_ ;
  assign \new_[67045]_  = A268 & A267;
  assign \new_[67046]_  = ~A266 & \new_[67045]_ ;
  assign \new_[67049]_  = A299 & ~A298;
  assign \new_[67052]_  = A301 & A300;
  assign \new_[67053]_  = \new_[67052]_  & \new_[67049]_ ;
  assign \new_[67054]_  = \new_[67053]_  & \new_[67046]_ ;
  assign \new_[67058]_  = A199 & ~A168;
  assign \new_[67059]_  = A170 & \new_[67058]_ ;
  assign \new_[67062]_  = A201 & ~A200;
  assign \new_[67065]_  = A265 & ~A203;
  assign \new_[67066]_  = \new_[67065]_  & \new_[67062]_ ;
  assign \new_[67067]_  = \new_[67066]_  & \new_[67059]_ ;
  assign \new_[67071]_  = A268 & A267;
  assign \new_[67072]_  = ~A266 & \new_[67071]_ ;
  assign \new_[67075]_  = A299 & ~A298;
  assign \new_[67078]_  = ~A302 & A300;
  assign \new_[67079]_  = \new_[67078]_  & \new_[67075]_ ;
  assign \new_[67080]_  = \new_[67079]_  & \new_[67072]_ ;
  assign \new_[67084]_  = A199 & ~A168;
  assign \new_[67085]_  = A170 & \new_[67084]_ ;
  assign \new_[67088]_  = A201 & ~A200;
  assign \new_[67091]_  = A265 & ~A203;
  assign \new_[67092]_  = \new_[67091]_  & \new_[67088]_ ;
  assign \new_[67093]_  = \new_[67092]_  & \new_[67085]_ ;
  assign \new_[67097]_  = ~A269 & A267;
  assign \new_[67098]_  = ~A266 & \new_[67097]_ ;
  assign \new_[67101]_  = ~A299 & A298;
  assign \new_[67104]_  = A301 & A300;
  assign \new_[67105]_  = \new_[67104]_  & \new_[67101]_ ;
  assign \new_[67106]_  = \new_[67105]_  & \new_[67098]_ ;
  assign \new_[67110]_  = A199 & ~A168;
  assign \new_[67111]_  = A170 & \new_[67110]_ ;
  assign \new_[67114]_  = A201 & ~A200;
  assign \new_[67117]_  = A265 & ~A203;
  assign \new_[67118]_  = \new_[67117]_  & \new_[67114]_ ;
  assign \new_[67119]_  = \new_[67118]_  & \new_[67111]_ ;
  assign \new_[67123]_  = ~A269 & A267;
  assign \new_[67124]_  = ~A266 & \new_[67123]_ ;
  assign \new_[67127]_  = ~A299 & A298;
  assign \new_[67130]_  = ~A302 & A300;
  assign \new_[67131]_  = \new_[67130]_  & \new_[67127]_ ;
  assign \new_[67132]_  = \new_[67131]_  & \new_[67124]_ ;
  assign \new_[67136]_  = A199 & ~A168;
  assign \new_[67137]_  = A170 & \new_[67136]_ ;
  assign \new_[67140]_  = A201 & ~A200;
  assign \new_[67143]_  = A265 & ~A203;
  assign \new_[67144]_  = \new_[67143]_  & \new_[67140]_ ;
  assign \new_[67145]_  = \new_[67144]_  & \new_[67137]_ ;
  assign \new_[67149]_  = ~A269 & A267;
  assign \new_[67150]_  = ~A266 & \new_[67149]_ ;
  assign \new_[67153]_  = A299 & ~A298;
  assign \new_[67156]_  = A301 & A300;
  assign \new_[67157]_  = \new_[67156]_  & \new_[67153]_ ;
  assign \new_[67158]_  = \new_[67157]_  & \new_[67150]_ ;
  assign \new_[67162]_  = A199 & ~A168;
  assign \new_[67163]_  = A170 & \new_[67162]_ ;
  assign \new_[67166]_  = A201 & ~A200;
  assign \new_[67169]_  = A265 & ~A203;
  assign \new_[67170]_  = \new_[67169]_  & \new_[67166]_ ;
  assign \new_[67171]_  = \new_[67170]_  & \new_[67163]_ ;
  assign \new_[67175]_  = ~A269 & A267;
  assign \new_[67176]_  = ~A266 & \new_[67175]_ ;
  assign \new_[67179]_  = A299 & ~A298;
  assign \new_[67182]_  = ~A302 & A300;
  assign \new_[67183]_  = \new_[67182]_  & \new_[67179]_ ;
  assign \new_[67184]_  = \new_[67183]_  & \new_[67176]_ ;
  assign \new_[67188]_  = A167 & A168;
  assign \new_[67189]_  = A169 & \new_[67188]_ ;
  assign \new_[67192]_  = A201 & ~A166;
  assign \new_[67195]_  = A203 & ~A202;
  assign \new_[67196]_  = \new_[67195]_  & \new_[67192]_ ;
  assign \new_[67197]_  = \new_[67196]_  & \new_[67189]_ ;
  assign \new_[67201]_  = A269 & ~A268;
  assign \new_[67202]_  = A267 & \new_[67201]_ ;
  assign \new_[67205]_  = ~A299 & A298;
  assign \new_[67208]_  = A301 & A300;
  assign \new_[67209]_  = \new_[67208]_  & \new_[67205]_ ;
  assign \new_[67210]_  = \new_[67209]_  & \new_[67202]_ ;
  assign \new_[67214]_  = A167 & A168;
  assign \new_[67215]_  = A169 & \new_[67214]_ ;
  assign \new_[67218]_  = A201 & ~A166;
  assign \new_[67221]_  = A203 & ~A202;
  assign \new_[67222]_  = \new_[67221]_  & \new_[67218]_ ;
  assign \new_[67223]_  = \new_[67222]_  & \new_[67215]_ ;
  assign \new_[67227]_  = A269 & ~A268;
  assign \new_[67228]_  = A267 & \new_[67227]_ ;
  assign \new_[67231]_  = ~A299 & A298;
  assign \new_[67234]_  = ~A302 & A300;
  assign \new_[67235]_  = \new_[67234]_  & \new_[67231]_ ;
  assign \new_[67236]_  = \new_[67235]_  & \new_[67228]_ ;
  assign \new_[67240]_  = A167 & A168;
  assign \new_[67241]_  = A169 & \new_[67240]_ ;
  assign \new_[67244]_  = A201 & ~A166;
  assign \new_[67247]_  = A203 & ~A202;
  assign \new_[67248]_  = \new_[67247]_  & \new_[67244]_ ;
  assign \new_[67249]_  = \new_[67248]_  & \new_[67241]_ ;
  assign \new_[67253]_  = A269 & ~A268;
  assign \new_[67254]_  = A267 & \new_[67253]_ ;
  assign \new_[67257]_  = A299 & ~A298;
  assign \new_[67260]_  = A301 & A300;
  assign \new_[67261]_  = \new_[67260]_  & \new_[67257]_ ;
  assign \new_[67262]_  = \new_[67261]_  & \new_[67254]_ ;
  assign \new_[67266]_  = A167 & A168;
  assign \new_[67267]_  = A169 & \new_[67266]_ ;
  assign \new_[67270]_  = A201 & ~A166;
  assign \new_[67273]_  = A203 & ~A202;
  assign \new_[67274]_  = \new_[67273]_  & \new_[67270]_ ;
  assign \new_[67275]_  = \new_[67274]_  & \new_[67267]_ ;
  assign \new_[67279]_  = A269 & ~A268;
  assign \new_[67280]_  = A267 & \new_[67279]_ ;
  assign \new_[67283]_  = A299 & ~A298;
  assign \new_[67286]_  = ~A302 & A300;
  assign \new_[67287]_  = \new_[67286]_  & \new_[67283]_ ;
  assign \new_[67288]_  = \new_[67287]_  & \new_[67280]_ ;
  assign \new_[67292]_  = A167 & A168;
  assign \new_[67293]_  = A169 & \new_[67292]_ ;
  assign \new_[67296]_  = A201 & ~A166;
  assign \new_[67299]_  = A203 & ~A202;
  assign \new_[67300]_  = \new_[67299]_  & \new_[67296]_ ;
  assign \new_[67301]_  = \new_[67300]_  & \new_[67293]_ ;
  assign \new_[67305]_  = A298 & A268;
  assign \new_[67306]_  = ~A267 & \new_[67305]_ ;
  assign \new_[67309]_  = ~A300 & ~A299;
  assign \new_[67312]_  = A302 & ~A301;
  assign \new_[67313]_  = \new_[67312]_  & \new_[67309]_ ;
  assign \new_[67314]_  = \new_[67313]_  & \new_[67306]_ ;
  assign \new_[67318]_  = A167 & A168;
  assign \new_[67319]_  = A169 & \new_[67318]_ ;
  assign \new_[67322]_  = A201 & ~A166;
  assign \new_[67325]_  = A203 & ~A202;
  assign \new_[67326]_  = \new_[67325]_  & \new_[67322]_ ;
  assign \new_[67327]_  = \new_[67326]_  & \new_[67319]_ ;
  assign \new_[67331]_  = ~A298 & A268;
  assign \new_[67332]_  = ~A267 & \new_[67331]_ ;
  assign \new_[67335]_  = ~A300 & A299;
  assign \new_[67338]_  = A302 & ~A301;
  assign \new_[67339]_  = \new_[67338]_  & \new_[67335]_ ;
  assign \new_[67340]_  = \new_[67339]_  & \new_[67332]_ ;
  assign \new_[67344]_  = A167 & A168;
  assign \new_[67345]_  = A169 & \new_[67344]_ ;
  assign \new_[67348]_  = A201 & ~A166;
  assign \new_[67351]_  = A203 & ~A202;
  assign \new_[67352]_  = \new_[67351]_  & \new_[67348]_ ;
  assign \new_[67353]_  = \new_[67352]_  & \new_[67345]_ ;
  assign \new_[67357]_  = A298 & ~A269;
  assign \new_[67358]_  = ~A267 & \new_[67357]_ ;
  assign \new_[67361]_  = ~A300 & ~A299;
  assign \new_[67364]_  = A302 & ~A301;
  assign \new_[67365]_  = \new_[67364]_  & \new_[67361]_ ;
  assign \new_[67366]_  = \new_[67365]_  & \new_[67358]_ ;
  assign \new_[67370]_  = A167 & A168;
  assign \new_[67371]_  = A169 & \new_[67370]_ ;
  assign \new_[67374]_  = A201 & ~A166;
  assign \new_[67377]_  = A203 & ~A202;
  assign \new_[67378]_  = \new_[67377]_  & \new_[67374]_ ;
  assign \new_[67379]_  = \new_[67378]_  & \new_[67371]_ ;
  assign \new_[67383]_  = ~A298 & ~A269;
  assign \new_[67384]_  = ~A267 & \new_[67383]_ ;
  assign \new_[67387]_  = ~A300 & A299;
  assign \new_[67390]_  = A302 & ~A301;
  assign \new_[67391]_  = \new_[67390]_  & \new_[67387]_ ;
  assign \new_[67392]_  = \new_[67391]_  & \new_[67384]_ ;
  assign \new_[67396]_  = A167 & A168;
  assign \new_[67397]_  = A169 & \new_[67396]_ ;
  assign \new_[67400]_  = A201 & ~A166;
  assign \new_[67403]_  = A203 & ~A202;
  assign \new_[67404]_  = \new_[67403]_  & \new_[67400]_ ;
  assign \new_[67405]_  = \new_[67404]_  & \new_[67397]_ ;
  assign \new_[67409]_  = A298 & A266;
  assign \new_[67410]_  = A265 & \new_[67409]_ ;
  assign \new_[67413]_  = ~A300 & ~A299;
  assign \new_[67416]_  = A302 & ~A301;
  assign \new_[67417]_  = \new_[67416]_  & \new_[67413]_ ;
  assign \new_[67418]_  = \new_[67417]_  & \new_[67410]_ ;
  assign \new_[67422]_  = A167 & A168;
  assign \new_[67423]_  = A169 & \new_[67422]_ ;
  assign \new_[67426]_  = A201 & ~A166;
  assign \new_[67429]_  = A203 & ~A202;
  assign \new_[67430]_  = \new_[67429]_  & \new_[67426]_ ;
  assign \new_[67431]_  = \new_[67430]_  & \new_[67423]_ ;
  assign \new_[67435]_  = ~A298 & A266;
  assign \new_[67436]_  = A265 & \new_[67435]_ ;
  assign \new_[67439]_  = ~A300 & A299;
  assign \new_[67442]_  = A302 & ~A301;
  assign \new_[67443]_  = \new_[67442]_  & \new_[67439]_ ;
  assign \new_[67444]_  = \new_[67443]_  & \new_[67436]_ ;
  assign \new_[67448]_  = A167 & A168;
  assign \new_[67449]_  = A169 & \new_[67448]_ ;
  assign \new_[67452]_  = A201 & ~A166;
  assign \new_[67455]_  = A203 & ~A202;
  assign \new_[67456]_  = \new_[67455]_  & \new_[67452]_ ;
  assign \new_[67457]_  = \new_[67456]_  & \new_[67449]_ ;
  assign \new_[67461]_  = A267 & A266;
  assign \new_[67462]_  = ~A265 & \new_[67461]_ ;
  assign \new_[67465]_  = A300 & A268;
  assign \new_[67468]_  = A302 & ~A301;
  assign \new_[67469]_  = \new_[67468]_  & \new_[67465]_ ;
  assign \new_[67470]_  = \new_[67469]_  & \new_[67462]_ ;
  assign \new_[67474]_  = A167 & A168;
  assign \new_[67475]_  = A169 & \new_[67474]_ ;
  assign \new_[67478]_  = A201 & ~A166;
  assign \new_[67481]_  = A203 & ~A202;
  assign \new_[67482]_  = \new_[67481]_  & \new_[67478]_ ;
  assign \new_[67483]_  = \new_[67482]_  & \new_[67475]_ ;
  assign \new_[67487]_  = A267 & A266;
  assign \new_[67488]_  = ~A265 & \new_[67487]_ ;
  assign \new_[67491]_  = A300 & ~A269;
  assign \new_[67494]_  = A302 & ~A301;
  assign \new_[67495]_  = \new_[67494]_  & \new_[67491]_ ;
  assign \new_[67496]_  = \new_[67495]_  & \new_[67488]_ ;
  assign \new_[67500]_  = A167 & A168;
  assign \new_[67501]_  = A169 & \new_[67500]_ ;
  assign \new_[67504]_  = A201 & ~A166;
  assign \new_[67507]_  = A203 & ~A202;
  assign \new_[67508]_  = \new_[67507]_  & \new_[67504]_ ;
  assign \new_[67509]_  = \new_[67508]_  & \new_[67501]_ ;
  assign \new_[67513]_  = ~A267 & A266;
  assign \new_[67514]_  = ~A265 & \new_[67513]_ ;
  assign \new_[67517]_  = A269 & ~A268;
  assign \new_[67520]_  = A301 & ~A300;
  assign \new_[67521]_  = \new_[67520]_  & \new_[67517]_ ;
  assign \new_[67522]_  = \new_[67521]_  & \new_[67514]_ ;
  assign \new_[67526]_  = A167 & A168;
  assign \new_[67527]_  = A169 & \new_[67526]_ ;
  assign \new_[67530]_  = A201 & ~A166;
  assign \new_[67533]_  = A203 & ~A202;
  assign \new_[67534]_  = \new_[67533]_  & \new_[67530]_ ;
  assign \new_[67535]_  = \new_[67534]_  & \new_[67527]_ ;
  assign \new_[67539]_  = ~A267 & A266;
  assign \new_[67540]_  = ~A265 & \new_[67539]_ ;
  assign \new_[67543]_  = A269 & ~A268;
  assign \new_[67546]_  = ~A302 & ~A300;
  assign \new_[67547]_  = \new_[67546]_  & \new_[67543]_ ;
  assign \new_[67548]_  = \new_[67547]_  & \new_[67540]_ ;
  assign \new_[67552]_  = A167 & A168;
  assign \new_[67553]_  = A169 & \new_[67552]_ ;
  assign \new_[67556]_  = A201 & ~A166;
  assign \new_[67559]_  = A203 & ~A202;
  assign \new_[67560]_  = \new_[67559]_  & \new_[67556]_ ;
  assign \new_[67561]_  = \new_[67560]_  & \new_[67553]_ ;
  assign \new_[67565]_  = ~A267 & A266;
  assign \new_[67566]_  = ~A265 & \new_[67565]_ ;
  assign \new_[67569]_  = A269 & ~A268;
  assign \new_[67572]_  = A299 & A298;
  assign \new_[67573]_  = \new_[67572]_  & \new_[67569]_ ;
  assign \new_[67574]_  = \new_[67573]_  & \new_[67566]_ ;
  assign \new_[67578]_  = A167 & A168;
  assign \new_[67579]_  = A169 & \new_[67578]_ ;
  assign \new_[67582]_  = A201 & ~A166;
  assign \new_[67585]_  = A203 & ~A202;
  assign \new_[67586]_  = \new_[67585]_  & \new_[67582]_ ;
  assign \new_[67587]_  = \new_[67586]_  & \new_[67579]_ ;
  assign \new_[67591]_  = ~A267 & A266;
  assign \new_[67592]_  = ~A265 & \new_[67591]_ ;
  assign \new_[67595]_  = A269 & ~A268;
  assign \new_[67598]_  = ~A299 & ~A298;
  assign \new_[67599]_  = \new_[67598]_  & \new_[67595]_ ;
  assign \new_[67600]_  = \new_[67599]_  & \new_[67592]_ ;
  assign \new_[67604]_  = A167 & A168;
  assign \new_[67605]_  = A169 & \new_[67604]_ ;
  assign \new_[67608]_  = A201 & ~A166;
  assign \new_[67611]_  = A203 & ~A202;
  assign \new_[67612]_  = \new_[67611]_  & \new_[67608]_ ;
  assign \new_[67613]_  = \new_[67612]_  & \new_[67605]_ ;
  assign \new_[67617]_  = A267 & ~A266;
  assign \new_[67618]_  = A265 & \new_[67617]_ ;
  assign \new_[67621]_  = A300 & A268;
  assign \new_[67624]_  = A302 & ~A301;
  assign \new_[67625]_  = \new_[67624]_  & \new_[67621]_ ;
  assign \new_[67626]_  = \new_[67625]_  & \new_[67618]_ ;
  assign \new_[67630]_  = A167 & A168;
  assign \new_[67631]_  = A169 & \new_[67630]_ ;
  assign \new_[67634]_  = A201 & ~A166;
  assign \new_[67637]_  = A203 & ~A202;
  assign \new_[67638]_  = \new_[67637]_  & \new_[67634]_ ;
  assign \new_[67639]_  = \new_[67638]_  & \new_[67631]_ ;
  assign \new_[67643]_  = A267 & ~A266;
  assign \new_[67644]_  = A265 & \new_[67643]_ ;
  assign \new_[67647]_  = A300 & ~A269;
  assign \new_[67650]_  = A302 & ~A301;
  assign \new_[67651]_  = \new_[67650]_  & \new_[67647]_ ;
  assign \new_[67652]_  = \new_[67651]_  & \new_[67644]_ ;
  assign \new_[67656]_  = A167 & A168;
  assign \new_[67657]_  = A169 & \new_[67656]_ ;
  assign \new_[67660]_  = A201 & ~A166;
  assign \new_[67663]_  = A203 & ~A202;
  assign \new_[67664]_  = \new_[67663]_  & \new_[67660]_ ;
  assign \new_[67665]_  = \new_[67664]_  & \new_[67657]_ ;
  assign \new_[67669]_  = ~A267 & ~A266;
  assign \new_[67670]_  = A265 & \new_[67669]_ ;
  assign \new_[67673]_  = A269 & ~A268;
  assign \new_[67676]_  = A301 & ~A300;
  assign \new_[67677]_  = \new_[67676]_  & \new_[67673]_ ;
  assign \new_[67678]_  = \new_[67677]_  & \new_[67670]_ ;
  assign \new_[67682]_  = A167 & A168;
  assign \new_[67683]_  = A169 & \new_[67682]_ ;
  assign \new_[67686]_  = A201 & ~A166;
  assign \new_[67689]_  = A203 & ~A202;
  assign \new_[67690]_  = \new_[67689]_  & \new_[67686]_ ;
  assign \new_[67691]_  = \new_[67690]_  & \new_[67683]_ ;
  assign \new_[67695]_  = ~A267 & ~A266;
  assign \new_[67696]_  = A265 & \new_[67695]_ ;
  assign \new_[67699]_  = A269 & ~A268;
  assign \new_[67702]_  = ~A302 & ~A300;
  assign \new_[67703]_  = \new_[67702]_  & \new_[67699]_ ;
  assign \new_[67704]_  = \new_[67703]_  & \new_[67696]_ ;
  assign \new_[67708]_  = A167 & A168;
  assign \new_[67709]_  = A169 & \new_[67708]_ ;
  assign \new_[67712]_  = A201 & ~A166;
  assign \new_[67715]_  = A203 & ~A202;
  assign \new_[67716]_  = \new_[67715]_  & \new_[67712]_ ;
  assign \new_[67717]_  = \new_[67716]_  & \new_[67709]_ ;
  assign \new_[67721]_  = ~A267 & ~A266;
  assign \new_[67722]_  = A265 & \new_[67721]_ ;
  assign \new_[67725]_  = A269 & ~A268;
  assign \new_[67728]_  = A299 & A298;
  assign \new_[67729]_  = \new_[67728]_  & \new_[67725]_ ;
  assign \new_[67730]_  = \new_[67729]_  & \new_[67722]_ ;
  assign \new_[67734]_  = A167 & A168;
  assign \new_[67735]_  = A169 & \new_[67734]_ ;
  assign \new_[67738]_  = A201 & ~A166;
  assign \new_[67741]_  = A203 & ~A202;
  assign \new_[67742]_  = \new_[67741]_  & \new_[67738]_ ;
  assign \new_[67743]_  = \new_[67742]_  & \new_[67735]_ ;
  assign \new_[67747]_  = ~A267 & ~A266;
  assign \new_[67748]_  = A265 & \new_[67747]_ ;
  assign \new_[67751]_  = A269 & ~A268;
  assign \new_[67754]_  = ~A299 & ~A298;
  assign \new_[67755]_  = \new_[67754]_  & \new_[67751]_ ;
  assign \new_[67756]_  = \new_[67755]_  & \new_[67748]_ ;
  assign \new_[67760]_  = A167 & A168;
  assign \new_[67761]_  = A169 & \new_[67760]_ ;
  assign \new_[67764]_  = A201 & ~A166;
  assign \new_[67767]_  = A203 & ~A202;
  assign \new_[67768]_  = \new_[67767]_  & \new_[67764]_ ;
  assign \new_[67769]_  = \new_[67768]_  & \new_[67761]_ ;
  assign \new_[67773]_  = A298 & ~A266;
  assign \new_[67774]_  = ~A265 & \new_[67773]_ ;
  assign \new_[67777]_  = ~A300 & ~A299;
  assign \new_[67780]_  = A302 & ~A301;
  assign \new_[67781]_  = \new_[67780]_  & \new_[67777]_ ;
  assign \new_[67782]_  = \new_[67781]_  & \new_[67774]_ ;
  assign \new_[67786]_  = A167 & A168;
  assign \new_[67787]_  = A169 & \new_[67786]_ ;
  assign \new_[67790]_  = A201 & ~A166;
  assign \new_[67793]_  = A203 & ~A202;
  assign \new_[67794]_  = \new_[67793]_  & \new_[67790]_ ;
  assign \new_[67795]_  = \new_[67794]_  & \new_[67787]_ ;
  assign \new_[67799]_  = ~A298 & ~A266;
  assign \new_[67800]_  = ~A265 & \new_[67799]_ ;
  assign \new_[67803]_  = ~A300 & A299;
  assign \new_[67806]_  = A302 & ~A301;
  assign \new_[67807]_  = \new_[67806]_  & \new_[67803]_ ;
  assign \new_[67808]_  = \new_[67807]_  & \new_[67800]_ ;
  assign \new_[67812]_  = A167 & A168;
  assign \new_[67813]_  = A169 & \new_[67812]_ ;
  assign \new_[67816]_  = ~A201 & ~A166;
  assign \new_[67819]_  = A267 & A202;
  assign \new_[67820]_  = \new_[67819]_  & \new_[67816]_ ;
  assign \new_[67821]_  = \new_[67820]_  & \new_[67813]_ ;
  assign \new_[67825]_  = A298 & A269;
  assign \new_[67826]_  = ~A268 & \new_[67825]_ ;
  assign \new_[67829]_  = ~A300 & ~A299;
  assign \new_[67832]_  = A302 & ~A301;
  assign \new_[67833]_  = \new_[67832]_  & \new_[67829]_ ;
  assign \new_[67834]_  = \new_[67833]_  & \new_[67826]_ ;
  assign \new_[67838]_  = A167 & A168;
  assign \new_[67839]_  = A169 & \new_[67838]_ ;
  assign \new_[67842]_  = ~A201 & ~A166;
  assign \new_[67845]_  = A267 & A202;
  assign \new_[67846]_  = \new_[67845]_  & \new_[67842]_ ;
  assign \new_[67847]_  = \new_[67846]_  & \new_[67839]_ ;
  assign \new_[67851]_  = ~A298 & A269;
  assign \new_[67852]_  = ~A268 & \new_[67851]_ ;
  assign \new_[67855]_  = ~A300 & A299;
  assign \new_[67858]_  = A302 & ~A301;
  assign \new_[67859]_  = \new_[67858]_  & \new_[67855]_ ;
  assign \new_[67860]_  = \new_[67859]_  & \new_[67852]_ ;
  assign \new_[67864]_  = A167 & A168;
  assign \new_[67865]_  = A169 & \new_[67864]_ ;
  assign \new_[67868]_  = ~A201 & ~A166;
  assign \new_[67871]_  = ~A265 & A202;
  assign \new_[67872]_  = \new_[67871]_  & \new_[67868]_ ;
  assign \new_[67873]_  = \new_[67872]_  & \new_[67865]_ ;
  assign \new_[67877]_  = ~A268 & ~A267;
  assign \new_[67878]_  = A266 & \new_[67877]_ ;
  assign \new_[67881]_  = A300 & A269;
  assign \new_[67884]_  = A302 & ~A301;
  assign \new_[67885]_  = \new_[67884]_  & \new_[67881]_ ;
  assign \new_[67886]_  = \new_[67885]_  & \new_[67878]_ ;
  assign \new_[67890]_  = A167 & A168;
  assign \new_[67891]_  = A169 & \new_[67890]_ ;
  assign \new_[67894]_  = ~A201 & ~A166;
  assign \new_[67897]_  = A265 & A202;
  assign \new_[67898]_  = \new_[67897]_  & \new_[67894]_ ;
  assign \new_[67899]_  = \new_[67898]_  & \new_[67891]_ ;
  assign \new_[67903]_  = ~A268 & ~A267;
  assign \new_[67904]_  = ~A266 & \new_[67903]_ ;
  assign \new_[67907]_  = A300 & A269;
  assign \new_[67910]_  = A302 & ~A301;
  assign \new_[67911]_  = \new_[67910]_  & \new_[67907]_ ;
  assign \new_[67912]_  = \new_[67911]_  & \new_[67904]_ ;
  assign \new_[67916]_  = A167 & A168;
  assign \new_[67917]_  = A169 & \new_[67916]_ ;
  assign \new_[67920]_  = ~A201 & ~A166;
  assign \new_[67923]_  = A267 & ~A203;
  assign \new_[67924]_  = \new_[67923]_  & \new_[67920]_ ;
  assign \new_[67925]_  = \new_[67924]_  & \new_[67917]_ ;
  assign \new_[67929]_  = A298 & A269;
  assign \new_[67930]_  = ~A268 & \new_[67929]_ ;
  assign \new_[67933]_  = ~A300 & ~A299;
  assign \new_[67936]_  = A302 & ~A301;
  assign \new_[67937]_  = \new_[67936]_  & \new_[67933]_ ;
  assign \new_[67938]_  = \new_[67937]_  & \new_[67930]_ ;
  assign \new_[67942]_  = A167 & A168;
  assign \new_[67943]_  = A169 & \new_[67942]_ ;
  assign \new_[67946]_  = ~A201 & ~A166;
  assign \new_[67949]_  = A267 & ~A203;
  assign \new_[67950]_  = \new_[67949]_  & \new_[67946]_ ;
  assign \new_[67951]_  = \new_[67950]_  & \new_[67943]_ ;
  assign \new_[67955]_  = ~A298 & A269;
  assign \new_[67956]_  = ~A268 & \new_[67955]_ ;
  assign \new_[67959]_  = ~A300 & A299;
  assign \new_[67962]_  = A302 & ~A301;
  assign \new_[67963]_  = \new_[67962]_  & \new_[67959]_ ;
  assign \new_[67964]_  = \new_[67963]_  & \new_[67956]_ ;
  assign \new_[67968]_  = A167 & A168;
  assign \new_[67969]_  = A169 & \new_[67968]_ ;
  assign \new_[67972]_  = ~A201 & ~A166;
  assign \new_[67975]_  = ~A265 & ~A203;
  assign \new_[67976]_  = \new_[67975]_  & \new_[67972]_ ;
  assign \new_[67977]_  = \new_[67976]_  & \new_[67969]_ ;
  assign \new_[67981]_  = ~A268 & ~A267;
  assign \new_[67982]_  = A266 & \new_[67981]_ ;
  assign \new_[67985]_  = A300 & A269;
  assign \new_[67988]_  = A302 & ~A301;
  assign \new_[67989]_  = \new_[67988]_  & \new_[67985]_ ;
  assign \new_[67990]_  = \new_[67989]_  & \new_[67982]_ ;
  assign \new_[67994]_  = A167 & A168;
  assign \new_[67995]_  = A169 & \new_[67994]_ ;
  assign \new_[67998]_  = ~A201 & ~A166;
  assign \new_[68001]_  = A265 & ~A203;
  assign \new_[68002]_  = \new_[68001]_  & \new_[67998]_ ;
  assign \new_[68003]_  = \new_[68002]_  & \new_[67995]_ ;
  assign \new_[68007]_  = ~A268 & ~A267;
  assign \new_[68008]_  = ~A266 & \new_[68007]_ ;
  assign \new_[68011]_  = A300 & A269;
  assign \new_[68014]_  = A302 & ~A301;
  assign \new_[68015]_  = \new_[68014]_  & \new_[68011]_ ;
  assign \new_[68016]_  = \new_[68015]_  & \new_[68008]_ ;
  assign \new_[68020]_  = A167 & A168;
  assign \new_[68021]_  = A169 & \new_[68020]_ ;
  assign \new_[68024]_  = A199 & ~A166;
  assign \new_[68027]_  = A267 & A200;
  assign \new_[68028]_  = \new_[68027]_  & \new_[68024]_ ;
  assign \new_[68029]_  = \new_[68028]_  & \new_[68021]_ ;
  assign \new_[68033]_  = A298 & A269;
  assign \new_[68034]_  = ~A268 & \new_[68033]_ ;
  assign \new_[68037]_  = ~A300 & ~A299;
  assign \new_[68040]_  = A302 & ~A301;
  assign \new_[68041]_  = \new_[68040]_  & \new_[68037]_ ;
  assign \new_[68042]_  = \new_[68041]_  & \new_[68034]_ ;
  assign \new_[68046]_  = A167 & A168;
  assign \new_[68047]_  = A169 & \new_[68046]_ ;
  assign \new_[68050]_  = A199 & ~A166;
  assign \new_[68053]_  = A267 & A200;
  assign \new_[68054]_  = \new_[68053]_  & \new_[68050]_ ;
  assign \new_[68055]_  = \new_[68054]_  & \new_[68047]_ ;
  assign \new_[68059]_  = ~A298 & A269;
  assign \new_[68060]_  = ~A268 & \new_[68059]_ ;
  assign \new_[68063]_  = ~A300 & A299;
  assign \new_[68066]_  = A302 & ~A301;
  assign \new_[68067]_  = \new_[68066]_  & \new_[68063]_ ;
  assign \new_[68068]_  = \new_[68067]_  & \new_[68060]_ ;
  assign \new_[68072]_  = A167 & A168;
  assign \new_[68073]_  = A169 & \new_[68072]_ ;
  assign \new_[68076]_  = A199 & ~A166;
  assign \new_[68079]_  = ~A265 & A200;
  assign \new_[68080]_  = \new_[68079]_  & \new_[68076]_ ;
  assign \new_[68081]_  = \new_[68080]_  & \new_[68073]_ ;
  assign \new_[68085]_  = ~A268 & ~A267;
  assign \new_[68086]_  = A266 & \new_[68085]_ ;
  assign \new_[68089]_  = A300 & A269;
  assign \new_[68092]_  = A302 & ~A301;
  assign \new_[68093]_  = \new_[68092]_  & \new_[68089]_ ;
  assign \new_[68094]_  = \new_[68093]_  & \new_[68086]_ ;
  assign \new_[68098]_  = A167 & A168;
  assign \new_[68099]_  = A169 & \new_[68098]_ ;
  assign \new_[68102]_  = A199 & ~A166;
  assign \new_[68105]_  = A265 & A200;
  assign \new_[68106]_  = \new_[68105]_  & \new_[68102]_ ;
  assign \new_[68107]_  = \new_[68106]_  & \new_[68099]_ ;
  assign \new_[68111]_  = ~A268 & ~A267;
  assign \new_[68112]_  = ~A266 & \new_[68111]_ ;
  assign \new_[68115]_  = A300 & A269;
  assign \new_[68118]_  = A302 & ~A301;
  assign \new_[68119]_  = \new_[68118]_  & \new_[68115]_ ;
  assign \new_[68120]_  = \new_[68119]_  & \new_[68112]_ ;
  assign \new_[68124]_  = A167 & A168;
  assign \new_[68125]_  = A169 & \new_[68124]_ ;
  assign \new_[68128]_  = ~A199 & ~A166;
  assign \new_[68131]_  = A267 & ~A200;
  assign \new_[68132]_  = \new_[68131]_  & \new_[68128]_ ;
  assign \new_[68133]_  = \new_[68132]_  & \new_[68125]_ ;
  assign \new_[68137]_  = A298 & A269;
  assign \new_[68138]_  = ~A268 & \new_[68137]_ ;
  assign \new_[68141]_  = ~A300 & ~A299;
  assign \new_[68144]_  = A302 & ~A301;
  assign \new_[68145]_  = \new_[68144]_  & \new_[68141]_ ;
  assign \new_[68146]_  = \new_[68145]_  & \new_[68138]_ ;
  assign \new_[68150]_  = A167 & A168;
  assign \new_[68151]_  = A169 & \new_[68150]_ ;
  assign \new_[68154]_  = ~A199 & ~A166;
  assign \new_[68157]_  = A267 & ~A200;
  assign \new_[68158]_  = \new_[68157]_  & \new_[68154]_ ;
  assign \new_[68159]_  = \new_[68158]_  & \new_[68151]_ ;
  assign \new_[68163]_  = ~A298 & A269;
  assign \new_[68164]_  = ~A268 & \new_[68163]_ ;
  assign \new_[68167]_  = ~A300 & A299;
  assign \new_[68170]_  = A302 & ~A301;
  assign \new_[68171]_  = \new_[68170]_  & \new_[68167]_ ;
  assign \new_[68172]_  = \new_[68171]_  & \new_[68164]_ ;
  assign \new_[68176]_  = A167 & A168;
  assign \new_[68177]_  = A169 & \new_[68176]_ ;
  assign \new_[68180]_  = ~A199 & ~A166;
  assign \new_[68183]_  = ~A265 & ~A200;
  assign \new_[68184]_  = \new_[68183]_  & \new_[68180]_ ;
  assign \new_[68185]_  = \new_[68184]_  & \new_[68177]_ ;
  assign \new_[68189]_  = ~A268 & ~A267;
  assign \new_[68190]_  = A266 & \new_[68189]_ ;
  assign \new_[68193]_  = A300 & A269;
  assign \new_[68196]_  = A302 & ~A301;
  assign \new_[68197]_  = \new_[68196]_  & \new_[68193]_ ;
  assign \new_[68198]_  = \new_[68197]_  & \new_[68190]_ ;
  assign \new_[68202]_  = A167 & A168;
  assign \new_[68203]_  = A169 & \new_[68202]_ ;
  assign \new_[68206]_  = ~A199 & ~A166;
  assign \new_[68209]_  = A265 & ~A200;
  assign \new_[68210]_  = \new_[68209]_  & \new_[68206]_ ;
  assign \new_[68211]_  = \new_[68210]_  & \new_[68203]_ ;
  assign \new_[68215]_  = ~A268 & ~A267;
  assign \new_[68216]_  = ~A266 & \new_[68215]_ ;
  assign \new_[68219]_  = A300 & A269;
  assign \new_[68222]_  = A302 & ~A301;
  assign \new_[68223]_  = \new_[68222]_  & \new_[68219]_ ;
  assign \new_[68224]_  = \new_[68223]_  & \new_[68216]_ ;
  assign \new_[68228]_  = ~A167 & A168;
  assign \new_[68229]_  = A169 & \new_[68228]_ ;
  assign \new_[68232]_  = A201 & A166;
  assign \new_[68235]_  = A203 & ~A202;
  assign \new_[68236]_  = \new_[68235]_  & \new_[68232]_ ;
  assign \new_[68237]_  = \new_[68236]_  & \new_[68229]_ ;
  assign \new_[68241]_  = A269 & ~A268;
  assign \new_[68242]_  = A267 & \new_[68241]_ ;
  assign \new_[68245]_  = ~A299 & A298;
  assign \new_[68248]_  = A301 & A300;
  assign \new_[68249]_  = \new_[68248]_  & \new_[68245]_ ;
  assign \new_[68250]_  = \new_[68249]_  & \new_[68242]_ ;
  assign \new_[68254]_  = ~A167 & A168;
  assign \new_[68255]_  = A169 & \new_[68254]_ ;
  assign \new_[68258]_  = A201 & A166;
  assign \new_[68261]_  = A203 & ~A202;
  assign \new_[68262]_  = \new_[68261]_  & \new_[68258]_ ;
  assign \new_[68263]_  = \new_[68262]_  & \new_[68255]_ ;
  assign \new_[68267]_  = A269 & ~A268;
  assign \new_[68268]_  = A267 & \new_[68267]_ ;
  assign \new_[68271]_  = ~A299 & A298;
  assign \new_[68274]_  = ~A302 & A300;
  assign \new_[68275]_  = \new_[68274]_  & \new_[68271]_ ;
  assign \new_[68276]_  = \new_[68275]_  & \new_[68268]_ ;
  assign \new_[68280]_  = ~A167 & A168;
  assign \new_[68281]_  = A169 & \new_[68280]_ ;
  assign \new_[68284]_  = A201 & A166;
  assign \new_[68287]_  = A203 & ~A202;
  assign \new_[68288]_  = \new_[68287]_  & \new_[68284]_ ;
  assign \new_[68289]_  = \new_[68288]_  & \new_[68281]_ ;
  assign \new_[68293]_  = A269 & ~A268;
  assign \new_[68294]_  = A267 & \new_[68293]_ ;
  assign \new_[68297]_  = A299 & ~A298;
  assign \new_[68300]_  = A301 & A300;
  assign \new_[68301]_  = \new_[68300]_  & \new_[68297]_ ;
  assign \new_[68302]_  = \new_[68301]_  & \new_[68294]_ ;
  assign \new_[68306]_  = ~A167 & A168;
  assign \new_[68307]_  = A169 & \new_[68306]_ ;
  assign \new_[68310]_  = A201 & A166;
  assign \new_[68313]_  = A203 & ~A202;
  assign \new_[68314]_  = \new_[68313]_  & \new_[68310]_ ;
  assign \new_[68315]_  = \new_[68314]_  & \new_[68307]_ ;
  assign \new_[68319]_  = A269 & ~A268;
  assign \new_[68320]_  = A267 & \new_[68319]_ ;
  assign \new_[68323]_  = A299 & ~A298;
  assign \new_[68326]_  = ~A302 & A300;
  assign \new_[68327]_  = \new_[68326]_  & \new_[68323]_ ;
  assign \new_[68328]_  = \new_[68327]_  & \new_[68320]_ ;
  assign \new_[68332]_  = ~A167 & A168;
  assign \new_[68333]_  = A169 & \new_[68332]_ ;
  assign \new_[68336]_  = A201 & A166;
  assign \new_[68339]_  = A203 & ~A202;
  assign \new_[68340]_  = \new_[68339]_  & \new_[68336]_ ;
  assign \new_[68341]_  = \new_[68340]_  & \new_[68333]_ ;
  assign \new_[68345]_  = A298 & A268;
  assign \new_[68346]_  = ~A267 & \new_[68345]_ ;
  assign \new_[68349]_  = ~A300 & ~A299;
  assign \new_[68352]_  = A302 & ~A301;
  assign \new_[68353]_  = \new_[68352]_  & \new_[68349]_ ;
  assign \new_[68354]_  = \new_[68353]_  & \new_[68346]_ ;
  assign \new_[68358]_  = ~A167 & A168;
  assign \new_[68359]_  = A169 & \new_[68358]_ ;
  assign \new_[68362]_  = A201 & A166;
  assign \new_[68365]_  = A203 & ~A202;
  assign \new_[68366]_  = \new_[68365]_  & \new_[68362]_ ;
  assign \new_[68367]_  = \new_[68366]_  & \new_[68359]_ ;
  assign \new_[68371]_  = ~A298 & A268;
  assign \new_[68372]_  = ~A267 & \new_[68371]_ ;
  assign \new_[68375]_  = ~A300 & A299;
  assign \new_[68378]_  = A302 & ~A301;
  assign \new_[68379]_  = \new_[68378]_  & \new_[68375]_ ;
  assign \new_[68380]_  = \new_[68379]_  & \new_[68372]_ ;
  assign \new_[68384]_  = ~A167 & A168;
  assign \new_[68385]_  = A169 & \new_[68384]_ ;
  assign \new_[68388]_  = A201 & A166;
  assign \new_[68391]_  = A203 & ~A202;
  assign \new_[68392]_  = \new_[68391]_  & \new_[68388]_ ;
  assign \new_[68393]_  = \new_[68392]_  & \new_[68385]_ ;
  assign \new_[68397]_  = A298 & ~A269;
  assign \new_[68398]_  = ~A267 & \new_[68397]_ ;
  assign \new_[68401]_  = ~A300 & ~A299;
  assign \new_[68404]_  = A302 & ~A301;
  assign \new_[68405]_  = \new_[68404]_  & \new_[68401]_ ;
  assign \new_[68406]_  = \new_[68405]_  & \new_[68398]_ ;
  assign \new_[68410]_  = ~A167 & A168;
  assign \new_[68411]_  = A169 & \new_[68410]_ ;
  assign \new_[68414]_  = A201 & A166;
  assign \new_[68417]_  = A203 & ~A202;
  assign \new_[68418]_  = \new_[68417]_  & \new_[68414]_ ;
  assign \new_[68419]_  = \new_[68418]_  & \new_[68411]_ ;
  assign \new_[68423]_  = ~A298 & ~A269;
  assign \new_[68424]_  = ~A267 & \new_[68423]_ ;
  assign \new_[68427]_  = ~A300 & A299;
  assign \new_[68430]_  = A302 & ~A301;
  assign \new_[68431]_  = \new_[68430]_  & \new_[68427]_ ;
  assign \new_[68432]_  = \new_[68431]_  & \new_[68424]_ ;
  assign \new_[68436]_  = ~A167 & A168;
  assign \new_[68437]_  = A169 & \new_[68436]_ ;
  assign \new_[68440]_  = A201 & A166;
  assign \new_[68443]_  = A203 & ~A202;
  assign \new_[68444]_  = \new_[68443]_  & \new_[68440]_ ;
  assign \new_[68445]_  = \new_[68444]_  & \new_[68437]_ ;
  assign \new_[68449]_  = A298 & A266;
  assign \new_[68450]_  = A265 & \new_[68449]_ ;
  assign \new_[68453]_  = ~A300 & ~A299;
  assign \new_[68456]_  = A302 & ~A301;
  assign \new_[68457]_  = \new_[68456]_  & \new_[68453]_ ;
  assign \new_[68458]_  = \new_[68457]_  & \new_[68450]_ ;
  assign \new_[68462]_  = ~A167 & A168;
  assign \new_[68463]_  = A169 & \new_[68462]_ ;
  assign \new_[68466]_  = A201 & A166;
  assign \new_[68469]_  = A203 & ~A202;
  assign \new_[68470]_  = \new_[68469]_  & \new_[68466]_ ;
  assign \new_[68471]_  = \new_[68470]_  & \new_[68463]_ ;
  assign \new_[68475]_  = ~A298 & A266;
  assign \new_[68476]_  = A265 & \new_[68475]_ ;
  assign \new_[68479]_  = ~A300 & A299;
  assign \new_[68482]_  = A302 & ~A301;
  assign \new_[68483]_  = \new_[68482]_  & \new_[68479]_ ;
  assign \new_[68484]_  = \new_[68483]_  & \new_[68476]_ ;
  assign \new_[68488]_  = ~A167 & A168;
  assign \new_[68489]_  = A169 & \new_[68488]_ ;
  assign \new_[68492]_  = A201 & A166;
  assign \new_[68495]_  = A203 & ~A202;
  assign \new_[68496]_  = \new_[68495]_  & \new_[68492]_ ;
  assign \new_[68497]_  = \new_[68496]_  & \new_[68489]_ ;
  assign \new_[68501]_  = A267 & A266;
  assign \new_[68502]_  = ~A265 & \new_[68501]_ ;
  assign \new_[68505]_  = A300 & A268;
  assign \new_[68508]_  = A302 & ~A301;
  assign \new_[68509]_  = \new_[68508]_  & \new_[68505]_ ;
  assign \new_[68510]_  = \new_[68509]_  & \new_[68502]_ ;
  assign \new_[68514]_  = ~A167 & A168;
  assign \new_[68515]_  = A169 & \new_[68514]_ ;
  assign \new_[68518]_  = A201 & A166;
  assign \new_[68521]_  = A203 & ~A202;
  assign \new_[68522]_  = \new_[68521]_  & \new_[68518]_ ;
  assign \new_[68523]_  = \new_[68522]_  & \new_[68515]_ ;
  assign \new_[68527]_  = A267 & A266;
  assign \new_[68528]_  = ~A265 & \new_[68527]_ ;
  assign \new_[68531]_  = A300 & ~A269;
  assign \new_[68534]_  = A302 & ~A301;
  assign \new_[68535]_  = \new_[68534]_  & \new_[68531]_ ;
  assign \new_[68536]_  = \new_[68535]_  & \new_[68528]_ ;
  assign \new_[68540]_  = ~A167 & A168;
  assign \new_[68541]_  = A169 & \new_[68540]_ ;
  assign \new_[68544]_  = A201 & A166;
  assign \new_[68547]_  = A203 & ~A202;
  assign \new_[68548]_  = \new_[68547]_  & \new_[68544]_ ;
  assign \new_[68549]_  = \new_[68548]_  & \new_[68541]_ ;
  assign \new_[68553]_  = ~A267 & A266;
  assign \new_[68554]_  = ~A265 & \new_[68553]_ ;
  assign \new_[68557]_  = A269 & ~A268;
  assign \new_[68560]_  = A301 & ~A300;
  assign \new_[68561]_  = \new_[68560]_  & \new_[68557]_ ;
  assign \new_[68562]_  = \new_[68561]_  & \new_[68554]_ ;
  assign \new_[68566]_  = ~A167 & A168;
  assign \new_[68567]_  = A169 & \new_[68566]_ ;
  assign \new_[68570]_  = A201 & A166;
  assign \new_[68573]_  = A203 & ~A202;
  assign \new_[68574]_  = \new_[68573]_  & \new_[68570]_ ;
  assign \new_[68575]_  = \new_[68574]_  & \new_[68567]_ ;
  assign \new_[68579]_  = ~A267 & A266;
  assign \new_[68580]_  = ~A265 & \new_[68579]_ ;
  assign \new_[68583]_  = A269 & ~A268;
  assign \new_[68586]_  = ~A302 & ~A300;
  assign \new_[68587]_  = \new_[68586]_  & \new_[68583]_ ;
  assign \new_[68588]_  = \new_[68587]_  & \new_[68580]_ ;
  assign \new_[68592]_  = ~A167 & A168;
  assign \new_[68593]_  = A169 & \new_[68592]_ ;
  assign \new_[68596]_  = A201 & A166;
  assign \new_[68599]_  = A203 & ~A202;
  assign \new_[68600]_  = \new_[68599]_  & \new_[68596]_ ;
  assign \new_[68601]_  = \new_[68600]_  & \new_[68593]_ ;
  assign \new_[68605]_  = ~A267 & A266;
  assign \new_[68606]_  = ~A265 & \new_[68605]_ ;
  assign \new_[68609]_  = A269 & ~A268;
  assign \new_[68612]_  = A299 & A298;
  assign \new_[68613]_  = \new_[68612]_  & \new_[68609]_ ;
  assign \new_[68614]_  = \new_[68613]_  & \new_[68606]_ ;
  assign \new_[68618]_  = ~A167 & A168;
  assign \new_[68619]_  = A169 & \new_[68618]_ ;
  assign \new_[68622]_  = A201 & A166;
  assign \new_[68625]_  = A203 & ~A202;
  assign \new_[68626]_  = \new_[68625]_  & \new_[68622]_ ;
  assign \new_[68627]_  = \new_[68626]_  & \new_[68619]_ ;
  assign \new_[68631]_  = ~A267 & A266;
  assign \new_[68632]_  = ~A265 & \new_[68631]_ ;
  assign \new_[68635]_  = A269 & ~A268;
  assign \new_[68638]_  = ~A299 & ~A298;
  assign \new_[68639]_  = \new_[68638]_  & \new_[68635]_ ;
  assign \new_[68640]_  = \new_[68639]_  & \new_[68632]_ ;
  assign \new_[68644]_  = ~A167 & A168;
  assign \new_[68645]_  = A169 & \new_[68644]_ ;
  assign \new_[68648]_  = A201 & A166;
  assign \new_[68651]_  = A203 & ~A202;
  assign \new_[68652]_  = \new_[68651]_  & \new_[68648]_ ;
  assign \new_[68653]_  = \new_[68652]_  & \new_[68645]_ ;
  assign \new_[68657]_  = A267 & ~A266;
  assign \new_[68658]_  = A265 & \new_[68657]_ ;
  assign \new_[68661]_  = A300 & A268;
  assign \new_[68664]_  = A302 & ~A301;
  assign \new_[68665]_  = \new_[68664]_  & \new_[68661]_ ;
  assign \new_[68666]_  = \new_[68665]_  & \new_[68658]_ ;
  assign \new_[68670]_  = ~A167 & A168;
  assign \new_[68671]_  = A169 & \new_[68670]_ ;
  assign \new_[68674]_  = A201 & A166;
  assign \new_[68677]_  = A203 & ~A202;
  assign \new_[68678]_  = \new_[68677]_  & \new_[68674]_ ;
  assign \new_[68679]_  = \new_[68678]_  & \new_[68671]_ ;
  assign \new_[68683]_  = A267 & ~A266;
  assign \new_[68684]_  = A265 & \new_[68683]_ ;
  assign \new_[68687]_  = A300 & ~A269;
  assign \new_[68690]_  = A302 & ~A301;
  assign \new_[68691]_  = \new_[68690]_  & \new_[68687]_ ;
  assign \new_[68692]_  = \new_[68691]_  & \new_[68684]_ ;
  assign \new_[68696]_  = ~A167 & A168;
  assign \new_[68697]_  = A169 & \new_[68696]_ ;
  assign \new_[68700]_  = A201 & A166;
  assign \new_[68703]_  = A203 & ~A202;
  assign \new_[68704]_  = \new_[68703]_  & \new_[68700]_ ;
  assign \new_[68705]_  = \new_[68704]_  & \new_[68697]_ ;
  assign \new_[68709]_  = ~A267 & ~A266;
  assign \new_[68710]_  = A265 & \new_[68709]_ ;
  assign \new_[68713]_  = A269 & ~A268;
  assign \new_[68716]_  = A301 & ~A300;
  assign \new_[68717]_  = \new_[68716]_  & \new_[68713]_ ;
  assign \new_[68718]_  = \new_[68717]_  & \new_[68710]_ ;
  assign \new_[68722]_  = ~A167 & A168;
  assign \new_[68723]_  = A169 & \new_[68722]_ ;
  assign \new_[68726]_  = A201 & A166;
  assign \new_[68729]_  = A203 & ~A202;
  assign \new_[68730]_  = \new_[68729]_  & \new_[68726]_ ;
  assign \new_[68731]_  = \new_[68730]_  & \new_[68723]_ ;
  assign \new_[68735]_  = ~A267 & ~A266;
  assign \new_[68736]_  = A265 & \new_[68735]_ ;
  assign \new_[68739]_  = A269 & ~A268;
  assign \new_[68742]_  = ~A302 & ~A300;
  assign \new_[68743]_  = \new_[68742]_  & \new_[68739]_ ;
  assign \new_[68744]_  = \new_[68743]_  & \new_[68736]_ ;
  assign \new_[68748]_  = ~A167 & A168;
  assign \new_[68749]_  = A169 & \new_[68748]_ ;
  assign \new_[68752]_  = A201 & A166;
  assign \new_[68755]_  = A203 & ~A202;
  assign \new_[68756]_  = \new_[68755]_  & \new_[68752]_ ;
  assign \new_[68757]_  = \new_[68756]_  & \new_[68749]_ ;
  assign \new_[68761]_  = ~A267 & ~A266;
  assign \new_[68762]_  = A265 & \new_[68761]_ ;
  assign \new_[68765]_  = A269 & ~A268;
  assign \new_[68768]_  = A299 & A298;
  assign \new_[68769]_  = \new_[68768]_  & \new_[68765]_ ;
  assign \new_[68770]_  = \new_[68769]_  & \new_[68762]_ ;
  assign \new_[68774]_  = ~A167 & A168;
  assign \new_[68775]_  = A169 & \new_[68774]_ ;
  assign \new_[68778]_  = A201 & A166;
  assign \new_[68781]_  = A203 & ~A202;
  assign \new_[68782]_  = \new_[68781]_  & \new_[68778]_ ;
  assign \new_[68783]_  = \new_[68782]_  & \new_[68775]_ ;
  assign \new_[68787]_  = ~A267 & ~A266;
  assign \new_[68788]_  = A265 & \new_[68787]_ ;
  assign \new_[68791]_  = A269 & ~A268;
  assign \new_[68794]_  = ~A299 & ~A298;
  assign \new_[68795]_  = \new_[68794]_  & \new_[68791]_ ;
  assign \new_[68796]_  = \new_[68795]_  & \new_[68788]_ ;
  assign \new_[68800]_  = ~A167 & A168;
  assign \new_[68801]_  = A169 & \new_[68800]_ ;
  assign \new_[68804]_  = A201 & A166;
  assign \new_[68807]_  = A203 & ~A202;
  assign \new_[68808]_  = \new_[68807]_  & \new_[68804]_ ;
  assign \new_[68809]_  = \new_[68808]_  & \new_[68801]_ ;
  assign \new_[68813]_  = A298 & ~A266;
  assign \new_[68814]_  = ~A265 & \new_[68813]_ ;
  assign \new_[68817]_  = ~A300 & ~A299;
  assign \new_[68820]_  = A302 & ~A301;
  assign \new_[68821]_  = \new_[68820]_  & \new_[68817]_ ;
  assign \new_[68822]_  = \new_[68821]_  & \new_[68814]_ ;
  assign \new_[68826]_  = ~A167 & A168;
  assign \new_[68827]_  = A169 & \new_[68826]_ ;
  assign \new_[68830]_  = A201 & A166;
  assign \new_[68833]_  = A203 & ~A202;
  assign \new_[68834]_  = \new_[68833]_  & \new_[68830]_ ;
  assign \new_[68835]_  = \new_[68834]_  & \new_[68827]_ ;
  assign \new_[68839]_  = ~A298 & ~A266;
  assign \new_[68840]_  = ~A265 & \new_[68839]_ ;
  assign \new_[68843]_  = ~A300 & A299;
  assign \new_[68846]_  = A302 & ~A301;
  assign \new_[68847]_  = \new_[68846]_  & \new_[68843]_ ;
  assign \new_[68848]_  = \new_[68847]_  & \new_[68840]_ ;
  assign \new_[68852]_  = ~A167 & A168;
  assign \new_[68853]_  = A169 & \new_[68852]_ ;
  assign \new_[68856]_  = ~A201 & A166;
  assign \new_[68859]_  = A267 & A202;
  assign \new_[68860]_  = \new_[68859]_  & \new_[68856]_ ;
  assign \new_[68861]_  = \new_[68860]_  & \new_[68853]_ ;
  assign \new_[68865]_  = A298 & A269;
  assign \new_[68866]_  = ~A268 & \new_[68865]_ ;
  assign \new_[68869]_  = ~A300 & ~A299;
  assign \new_[68872]_  = A302 & ~A301;
  assign \new_[68873]_  = \new_[68872]_  & \new_[68869]_ ;
  assign \new_[68874]_  = \new_[68873]_  & \new_[68866]_ ;
  assign \new_[68878]_  = ~A167 & A168;
  assign \new_[68879]_  = A169 & \new_[68878]_ ;
  assign \new_[68882]_  = ~A201 & A166;
  assign \new_[68885]_  = A267 & A202;
  assign \new_[68886]_  = \new_[68885]_  & \new_[68882]_ ;
  assign \new_[68887]_  = \new_[68886]_  & \new_[68879]_ ;
  assign \new_[68891]_  = ~A298 & A269;
  assign \new_[68892]_  = ~A268 & \new_[68891]_ ;
  assign \new_[68895]_  = ~A300 & A299;
  assign \new_[68898]_  = A302 & ~A301;
  assign \new_[68899]_  = \new_[68898]_  & \new_[68895]_ ;
  assign \new_[68900]_  = \new_[68899]_  & \new_[68892]_ ;
  assign \new_[68904]_  = ~A167 & A168;
  assign \new_[68905]_  = A169 & \new_[68904]_ ;
  assign \new_[68908]_  = ~A201 & A166;
  assign \new_[68911]_  = ~A265 & A202;
  assign \new_[68912]_  = \new_[68911]_  & \new_[68908]_ ;
  assign \new_[68913]_  = \new_[68912]_  & \new_[68905]_ ;
  assign \new_[68917]_  = ~A268 & ~A267;
  assign \new_[68918]_  = A266 & \new_[68917]_ ;
  assign \new_[68921]_  = A300 & A269;
  assign \new_[68924]_  = A302 & ~A301;
  assign \new_[68925]_  = \new_[68924]_  & \new_[68921]_ ;
  assign \new_[68926]_  = \new_[68925]_  & \new_[68918]_ ;
  assign \new_[68930]_  = ~A167 & A168;
  assign \new_[68931]_  = A169 & \new_[68930]_ ;
  assign \new_[68934]_  = ~A201 & A166;
  assign \new_[68937]_  = A265 & A202;
  assign \new_[68938]_  = \new_[68937]_  & \new_[68934]_ ;
  assign \new_[68939]_  = \new_[68938]_  & \new_[68931]_ ;
  assign \new_[68943]_  = ~A268 & ~A267;
  assign \new_[68944]_  = ~A266 & \new_[68943]_ ;
  assign \new_[68947]_  = A300 & A269;
  assign \new_[68950]_  = A302 & ~A301;
  assign \new_[68951]_  = \new_[68950]_  & \new_[68947]_ ;
  assign \new_[68952]_  = \new_[68951]_  & \new_[68944]_ ;
  assign \new_[68956]_  = ~A167 & A168;
  assign \new_[68957]_  = A169 & \new_[68956]_ ;
  assign \new_[68960]_  = ~A201 & A166;
  assign \new_[68963]_  = A267 & ~A203;
  assign \new_[68964]_  = \new_[68963]_  & \new_[68960]_ ;
  assign \new_[68965]_  = \new_[68964]_  & \new_[68957]_ ;
  assign \new_[68969]_  = A298 & A269;
  assign \new_[68970]_  = ~A268 & \new_[68969]_ ;
  assign \new_[68973]_  = ~A300 & ~A299;
  assign \new_[68976]_  = A302 & ~A301;
  assign \new_[68977]_  = \new_[68976]_  & \new_[68973]_ ;
  assign \new_[68978]_  = \new_[68977]_  & \new_[68970]_ ;
  assign \new_[68982]_  = ~A167 & A168;
  assign \new_[68983]_  = A169 & \new_[68982]_ ;
  assign \new_[68986]_  = ~A201 & A166;
  assign \new_[68989]_  = A267 & ~A203;
  assign \new_[68990]_  = \new_[68989]_  & \new_[68986]_ ;
  assign \new_[68991]_  = \new_[68990]_  & \new_[68983]_ ;
  assign \new_[68995]_  = ~A298 & A269;
  assign \new_[68996]_  = ~A268 & \new_[68995]_ ;
  assign \new_[68999]_  = ~A300 & A299;
  assign \new_[69002]_  = A302 & ~A301;
  assign \new_[69003]_  = \new_[69002]_  & \new_[68999]_ ;
  assign \new_[69004]_  = \new_[69003]_  & \new_[68996]_ ;
  assign \new_[69008]_  = ~A167 & A168;
  assign \new_[69009]_  = A169 & \new_[69008]_ ;
  assign \new_[69012]_  = ~A201 & A166;
  assign \new_[69015]_  = ~A265 & ~A203;
  assign \new_[69016]_  = \new_[69015]_  & \new_[69012]_ ;
  assign \new_[69017]_  = \new_[69016]_  & \new_[69009]_ ;
  assign \new_[69021]_  = ~A268 & ~A267;
  assign \new_[69022]_  = A266 & \new_[69021]_ ;
  assign \new_[69025]_  = A300 & A269;
  assign \new_[69028]_  = A302 & ~A301;
  assign \new_[69029]_  = \new_[69028]_  & \new_[69025]_ ;
  assign \new_[69030]_  = \new_[69029]_  & \new_[69022]_ ;
  assign \new_[69034]_  = ~A167 & A168;
  assign \new_[69035]_  = A169 & \new_[69034]_ ;
  assign \new_[69038]_  = ~A201 & A166;
  assign \new_[69041]_  = A265 & ~A203;
  assign \new_[69042]_  = \new_[69041]_  & \new_[69038]_ ;
  assign \new_[69043]_  = \new_[69042]_  & \new_[69035]_ ;
  assign \new_[69047]_  = ~A268 & ~A267;
  assign \new_[69048]_  = ~A266 & \new_[69047]_ ;
  assign \new_[69051]_  = A300 & A269;
  assign \new_[69054]_  = A302 & ~A301;
  assign \new_[69055]_  = \new_[69054]_  & \new_[69051]_ ;
  assign \new_[69056]_  = \new_[69055]_  & \new_[69048]_ ;
  assign \new_[69060]_  = ~A167 & A168;
  assign \new_[69061]_  = A169 & \new_[69060]_ ;
  assign \new_[69064]_  = A199 & A166;
  assign \new_[69067]_  = A267 & A200;
  assign \new_[69068]_  = \new_[69067]_  & \new_[69064]_ ;
  assign \new_[69069]_  = \new_[69068]_  & \new_[69061]_ ;
  assign \new_[69073]_  = A298 & A269;
  assign \new_[69074]_  = ~A268 & \new_[69073]_ ;
  assign \new_[69077]_  = ~A300 & ~A299;
  assign \new_[69080]_  = A302 & ~A301;
  assign \new_[69081]_  = \new_[69080]_  & \new_[69077]_ ;
  assign \new_[69082]_  = \new_[69081]_  & \new_[69074]_ ;
  assign \new_[69086]_  = ~A167 & A168;
  assign \new_[69087]_  = A169 & \new_[69086]_ ;
  assign \new_[69090]_  = A199 & A166;
  assign \new_[69093]_  = A267 & A200;
  assign \new_[69094]_  = \new_[69093]_  & \new_[69090]_ ;
  assign \new_[69095]_  = \new_[69094]_  & \new_[69087]_ ;
  assign \new_[69099]_  = ~A298 & A269;
  assign \new_[69100]_  = ~A268 & \new_[69099]_ ;
  assign \new_[69103]_  = ~A300 & A299;
  assign \new_[69106]_  = A302 & ~A301;
  assign \new_[69107]_  = \new_[69106]_  & \new_[69103]_ ;
  assign \new_[69108]_  = \new_[69107]_  & \new_[69100]_ ;
  assign \new_[69112]_  = ~A167 & A168;
  assign \new_[69113]_  = A169 & \new_[69112]_ ;
  assign \new_[69116]_  = A199 & A166;
  assign \new_[69119]_  = ~A265 & A200;
  assign \new_[69120]_  = \new_[69119]_  & \new_[69116]_ ;
  assign \new_[69121]_  = \new_[69120]_  & \new_[69113]_ ;
  assign \new_[69125]_  = ~A268 & ~A267;
  assign \new_[69126]_  = A266 & \new_[69125]_ ;
  assign \new_[69129]_  = A300 & A269;
  assign \new_[69132]_  = A302 & ~A301;
  assign \new_[69133]_  = \new_[69132]_  & \new_[69129]_ ;
  assign \new_[69134]_  = \new_[69133]_  & \new_[69126]_ ;
  assign \new_[69138]_  = ~A167 & A168;
  assign \new_[69139]_  = A169 & \new_[69138]_ ;
  assign \new_[69142]_  = A199 & A166;
  assign \new_[69145]_  = A265 & A200;
  assign \new_[69146]_  = \new_[69145]_  & \new_[69142]_ ;
  assign \new_[69147]_  = \new_[69146]_  & \new_[69139]_ ;
  assign \new_[69151]_  = ~A268 & ~A267;
  assign \new_[69152]_  = ~A266 & \new_[69151]_ ;
  assign \new_[69155]_  = A300 & A269;
  assign \new_[69158]_  = A302 & ~A301;
  assign \new_[69159]_  = \new_[69158]_  & \new_[69155]_ ;
  assign \new_[69160]_  = \new_[69159]_  & \new_[69152]_ ;
  assign \new_[69164]_  = ~A167 & A168;
  assign \new_[69165]_  = A169 & \new_[69164]_ ;
  assign \new_[69168]_  = ~A199 & A166;
  assign \new_[69171]_  = A267 & ~A200;
  assign \new_[69172]_  = \new_[69171]_  & \new_[69168]_ ;
  assign \new_[69173]_  = \new_[69172]_  & \new_[69165]_ ;
  assign \new_[69177]_  = A298 & A269;
  assign \new_[69178]_  = ~A268 & \new_[69177]_ ;
  assign \new_[69181]_  = ~A300 & ~A299;
  assign \new_[69184]_  = A302 & ~A301;
  assign \new_[69185]_  = \new_[69184]_  & \new_[69181]_ ;
  assign \new_[69186]_  = \new_[69185]_  & \new_[69178]_ ;
  assign \new_[69190]_  = ~A167 & A168;
  assign \new_[69191]_  = A169 & \new_[69190]_ ;
  assign \new_[69194]_  = ~A199 & A166;
  assign \new_[69197]_  = A267 & ~A200;
  assign \new_[69198]_  = \new_[69197]_  & \new_[69194]_ ;
  assign \new_[69199]_  = \new_[69198]_  & \new_[69191]_ ;
  assign \new_[69203]_  = ~A298 & A269;
  assign \new_[69204]_  = ~A268 & \new_[69203]_ ;
  assign \new_[69207]_  = ~A300 & A299;
  assign \new_[69210]_  = A302 & ~A301;
  assign \new_[69211]_  = \new_[69210]_  & \new_[69207]_ ;
  assign \new_[69212]_  = \new_[69211]_  & \new_[69204]_ ;
  assign \new_[69216]_  = ~A167 & A168;
  assign \new_[69217]_  = A169 & \new_[69216]_ ;
  assign \new_[69220]_  = ~A199 & A166;
  assign \new_[69223]_  = ~A265 & ~A200;
  assign \new_[69224]_  = \new_[69223]_  & \new_[69220]_ ;
  assign \new_[69225]_  = \new_[69224]_  & \new_[69217]_ ;
  assign \new_[69229]_  = ~A268 & ~A267;
  assign \new_[69230]_  = A266 & \new_[69229]_ ;
  assign \new_[69233]_  = A300 & A269;
  assign \new_[69236]_  = A302 & ~A301;
  assign \new_[69237]_  = \new_[69236]_  & \new_[69233]_ ;
  assign \new_[69238]_  = \new_[69237]_  & \new_[69230]_ ;
  assign \new_[69242]_  = ~A167 & A168;
  assign \new_[69243]_  = A169 & \new_[69242]_ ;
  assign \new_[69246]_  = ~A199 & A166;
  assign \new_[69249]_  = A265 & ~A200;
  assign \new_[69250]_  = \new_[69249]_  & \new_[69246]_ ;
  assign \new_[69251]_  = \new_[69250]_  & \new_[69243]_ ;
  assign \new_[69255]_  = ~A268 & ~A267;
  assign \new_[69256]_  = ~A266 & \new_[69255]_ ;
  assign \new_[69259]_  = A300 & A269;
  assign \new_[69262]_  = A302 & ~A301;
  assign \new_[69263]_  = \new_[69262]_  & \new_[69259]_ ;
  assign \new_[69264]_  = \new_[69263]_  & \new_[69256]_ ;
  assign \new_[69268]_  = ~A199 & ~A168;
  assign \new_[69269]_  = A169 & \new_[69268]_ ;
  assign \new_[69272]_  = A201 & A200;
  assign \new_[69275]_  = ~A265 & A202;
  assign \new_[69276]_  = \new_[69275]_  & \new_[69272]_ ;
  assign \new_[69277]_  = \new_[69276]_  & \new_[69269]_ ;
  assign \new_[69281]_  = A268 & A267;
  assign \new_[69282]_  = A266 & \new_[69281]_ ;
  assign \new_[69285]_  = ~A299 & A298;
  assign \new_[69288]_  = A301 & A300;
  assign \new_[69289]_  = \new_[69288]_  & \new_[69285]_ ;
  assign \new_[69290]_  = \new_[69289]_  & \new_[69282]_ ;
  assign \new_[69294]_  = ~A199 & ~A168;
  assign \new_[69295]_  = A169 & \new_[69294]_ ;
  assign \new_[69298]_  = A201 & A200;
  assign \new_[69301]_  = ~A265 & A202;
  assign \new_[69302]_  = \new_[69301]_  & \new_[69298]_ ;
  assign \new_[69303]_  = \new_[69302]_  & \new_[69295]_ ;
  assign \new_[69307]_  = A268 & A267;
  assign \new_[69308]_  = A266 & \new_[69307]_ ;
  assign \new_[69311]_  = ~A299 & A298;
  assign \new_[69314]_  = ~A302 & A300;
  assign \new_[69315]_  = \new_[69314]_  & \new_[69311]_ ;
  assign \new_[69316]_  = \new_[69315]_  & \new_[69308]_ ;
  assign \new_[69320]_  = ~A199 & ~A168;
  assign \new_[69321]_  = A169 & \new_[69320]_ ;
  assign \new_[69324]_  = A201 & A200;
  assign \new_[69327]_  = ~A265 & A202;
  assign \new_[69328]_  = \new_[69327]_  & \new_[69324]_ ;
  assign \new_[69329]_  = \new_[69328]_  & \new_[69321]_ ;
  assign \new_[69333]_  = A268 & A267;
  assign \new_[69334]_  = A266 & \new_[69333]_ ;
  assign \new_[69337]_  = A299 & ~A298;
  assign \new_[69340]_  = A301 & A300;
  assign \new_[69341]_  = \new_[69340]_  & \new_[69337]_ ;
  assign \new_[69342]_  = \new_[69341]_  & \new_[69334]_ ;
  assign \new_[69346]_  = ~A199 & ~A168;
  assign \new_[69347]_  = A169 & \new_[69346]_ ;
  assign \new_[69350]_  = A201 & A200;
  assign \new_[69353]_  = ~A265 & A202;
  assign \new_[69354]_  = \new_[69353]_  & \new_[69350]_ ;
  assign \new_[69355]_  = \new_[69354]_  & \new_[69347]_ ;
  assign \new_[69359]_  = A268 & A267;
  assign \new_[69360]_  = A266 & \new_[69359]_ ;
  assign \new_[69363]_  = A299 & ~A298;
  assign \new_[69366]_  = ~A302 & A300;
  assign \new_[69367]_  = \new_[69366]_  & \new_[69363]_ ;
  assign \new_[69368]_  = \new_[69367]_  & \new_[69360]_ ;
  assign \new_[69372]_  = ~A199 & ~A168;
  assign \new_[69373]_  = A169 & \new_[69372]_ ;
  assign \new_[69376]_  = A201 & A200;
  assign \new_[69379]_  = ~A265 & A202;
  assign \new_[69380]_  = \new_[69379]_  & \new_[69376]_ ;
  assign \new_[69381]_  = \new_[69380]_  & \new_[69373]_ ;
  assign \new_[69385]_  = ~A269 & A267;
  assign \new_[69386]_  = A266 & \new_[69385]_ ;
  assign \new_[69389]_  = ~A299 & A298;
  assign \new_[69392]_  = A301 & A300;
  assign \new_[69393]_  = \new_[69392]_  & \new_[69389]_ ;
  assign \new_[69394]_  = \new_[69393]_  & \new_[69386]_ ;
  assign \new_[69398]_  = ~A199 & ~A168;
  assign \new_[69399]_  = A169 & \new_[69398]_ ;
  assign \new_[69402]_  = A201 & A200;
  assign \new_[69405]_  = ~A265 & A202;
  assign \new_[69406]_  = \new_[69405]_  & \new_[69402]_ ;
  assign \new_[69407]_  = \new_[69406]_  & \new_[69399]_ ;
  assign \new_[69411]_  = ~A269 & A267;
  assign \new_[69412]_  = A266 & \new_[69411]_ ;
  assign \new_[69415]_  = ~A299 & A298;
  assign \new_[69418]_  = ~A302 & A300;
  assign \new_[69419]_  = \new_[69418]_  & \new_[69415]_ ;
  assign \new_[69420]_  = \new_[69419]_  & \new_[69412]_ ;
  assign \new_[69424]_  = ~A199 & ~A168;
  assign \new_[69425]_  = A169 & \new_[69424]_ ;
  assign \new_[69428]_  = A201 & A200;
  assign \new_[69431]_  = ~A265 & A202;
  assign \new_[69432]_  = \new_[69431]_  & \new_[69428]_ ;
  assign \new_[69433]_  = \new_[69432]_  & \new_[69425]_ ;
  assign \new_[69437]_  = ~A269 & A267;
  assign \new_[69438]_  = A266 & \new_[69437]_ ;
  assign \new_[69441]_  = A299 & ~A298;
  assign \new_[69444]_  = A301 & A300;
  assign \new_[69445]_  = \new_[69444]_  & \new_[69441]_ ;
  assign \new_[69446]_  = \new_[69445]_  & \new_[69438]_ ;
  assign \new_[69450]_  = ~A199 & ~A168;
  assign \new_[69451]_  = A169 & \new_[69450]_ ;
  assign \new_[69454]_  = A201 & A200;
  assign \new_[69457]_  = ~A265 & A202;
  assign \new_[69458]_  = \new_[69457]_  & \new_[69454]_ ;
  assign \new_[69459]_  = \new_[69458]_  & \new_[69451]_ ;
  assign \new_[69463]_  = ~A269 & A267;
  assign \new_[69464]_  = A266 & \new_[69463]_ ;
  assign \new_[69467]_  = A299 & ~A298;
  assign \new_[69470]_  = ~A302 & A300;
  assign \new_[69471]_  = \new_[69470]_  & \new_[69467]_ ;
  assign \new_[69472]_  = \new_[69471]_  & \new_[69464]_ ;
  assign \new_[69476]_  = ~A199 & ~A168;
  assign \new_[69477]_  = A169 & \new_[69476]_ ;
  assign \new_[69480]_  = A201 & A200;
  assign \new_[69483]_  = A265 & A202;
  assign \new_[69484]_  = \new_[69483]_  & \new_[69480]_ ;
  assign \new_[69485]_  = \new_[69484]_  & \new_[69477]_ ;
  assign \new_[69489]_  = A268 & A267;
  assign \new_[69490]_  = ~A266 & \new_[69489]_ ;
  assign \new_[69493]_  = ~A299 & A298;
  assign \new_[69496]_  = A301 & A300;
  assign \new_[69497]_  = \new_[69496]_  & \new_[69493]_ ;
  assign \new_[69498]_  = \new_[69497]_  & \new_[69490]_ ;
  assign \new_[69502]_  = ~A199 & ~A168;
  assign \new_[69503]_  = A169 & \new_[69502]_ ;
  assign \new_[69506]_  = A201 & A200;
  assign \new_[69509]_  = A265 & A202;
  assign \new_[69510]_  = \new_[69509]_  & \new_[69506]_ ;
  assign \new_[69511]_  = \new_[69510]_  & \new_[69503]_ ;
  assign \new_[69515]_  = A268 & A267;
  assign \new_[69516]_  = ~A266 & \new_[69515]_ ;
  assign \new_[69519]_  = ~A299 & A298;
  assign \new_[69522]_  = ~A302 & A300;
  assign \new_[69523]_  = \new_[69522]_  & \new_[69519]_ ;
  assign \new_[69524]_  = \new_[69523]_  & \new_[69516]_ ;
  assign \new_[69528]_  = ~A199 & ~A168;
  assign \new_[69529]_  = A169 & \new_[69528]_ ;
  assign \new_[69532]_  = A201 & A200;
  assign \new_[69535]_  = A265 & A202;
  assign \new_[69536]_  = \new_[69535]_  & \new_[69532]_ ;
  assign \new_[69537]_  = \new_[69536]_  & \new_[69529]_ ;
  assign \new_[69541]_  = A268 & A267;
  assign \new_[69542]_  = ~A266 & \new_[69541]_ ;
  assign \new_[69545]_  = A299 & ~A298;
  assign \new_[69548]_  = A301 & A300;
  assign \new_[69549]_  = \new_[69548]_  & \new_[69545]_ ;
  assign \new_[69550]_  = \new_[69549]_  & \new_[69542]_ ;
  assign \new_[69554]_  = ~A199 & ~A168;
  assign \new_[69555]_  = A169 & \new_[69554]_ ;
  assign \new_[69558]_  = A201 & A200;
  assign \new_[69561]_  = A265 & A202;
  assign \new_[69562]_  = \new_[69561]_  & \new_[69558]_ ;
  assign \new_[69563]_  = \new_[69562]_  & \new_[69555]_ ;
  assign \new_[69567]_  = A268 & A267;
  assign \new_[69568]_  = ~A266 & \new_[69567]_ ;
  assign \new_[69571]_  = A299 & ~A298;
  assign \new_[69574]_  = ~A302 & A300;
  assign \new_[69575]_  = \new_[69574]_  & \new_[69571]_ ;
  assign \new_[69576]_  = \new_[69575]_  & \new_[69568]_ ;
  assign \new_[69580]_  = ~A199 & ~A168;
  assign \new_[69581]_  = A169 & \new_[69580]_ ;
  assign \new_[69584]_  = A201 & A200;
  assign \new_[69587]_  = A265 & A202;
  assign \new_[69588]_  = \new_[69587]_  & \new_[69584]_ ;
  assign \new_[69589]_  = \new_[69588]_  & \new_[69581]_ ;
  assign \new_[69593]_  = ~A269 & A267;
  assign \new_[69594]_  = ~A266 & \new_[69593]_ ;
  assign \new_[69597]_  = ~A299 & A298;
  assign \new_[69600]_  = A301 & A300;
  assign \new_[69601]_  = \new_[69600]_  & \new_[69597]_ ;
  assign \new_[69602]_  = \new_[69601]_  & \new_[69594]_ ;
  assign \new_[69606]_  = ~A199 & ~A168;
  assign \new_[69607]_  = A169 & \new_[69606]_ ;
  assign \new_[69610]_  = A201 & A200;
  assign \new_[69613]_  = A265 & A202;
  assign \new_[69614]_  = \new_[69613]_  & \new_[69610]_ ;
  assign \new_[69615]_  = \new_[69614]_  & \new_[69607]_ ;
  assign \new_[69619]_  = ~A269 & A267;
  assign \new_[69620]_  = ~A266 & \new_[69619]_ ;
  assign \new_[69623]_  = ~A299 & A298;
  assign \new_[69626]_  = ~A302 & A300;
  assign \new_[69627]_  = \new_[69626]_  & \new_[69623]_ ;
  assign \new_[69628]_  = \new_[69627]_  & \new_[69620]_ ;
  assign \new_[69632]_  = ~A199 & ~A168;
  assign \new_[69633]_  = A169 & \new_[69632]_ ;
  assign \new_[69636]_  = A201 & A200;
  assign \new_[69639]_  = A265 & A202;
  assign \new_[69640]_  = \new_[69639]_  & \new_[69636]_ ;
  assign \new_[69641]_  = \new_[69640]_  & \new_[69633]_ ;
  assign \new_[69645]_  = ~A269 & A267;
  assign \new_[69646]_  = ~A266 & \new_[69645]_ ;
  assign \new_[69649]_  = A299 & ~A298;
  assign \new_[69652]_  = A301 & A300;
  assign \new_[69653]_  = \new_[69652]_  & \new_[69649]_ ;
  assign \new_[69654]_  = \new_[69653]_  & \new_[69646]_ ;
  assign \new_[69658]_  = ~A199 & ~A168;
  assign \new_[69659]_  = A169 & \new_[69658]_ ;
  assign \new_[69662]_  = A201 & A200;
  assign \new_[69665]_  = A265 & A202;
  assign \new_[69666]_  = \new_[69665]_  & \new_[69662]_ ;
  assign \new_[69667]_  = \new_[69666]_  & \new_[69659]_ ;
  assign \new_[69671]_  = ~A269 & A267;
  assign \new_[69672]_  = ~A266 & \new_[69671]_ ;
  assign \new_[69675]_  = A299 & ~A298;
  assign \new_[69678]_  = ~A302 & A300;
  assign \new_[69679]_  = \new_[69678]_  & \new_[69675]_ ;
  assign \new_[69680]_  = \new_[69679]_  & \new_[69672]_ ;
  assign \new_[69684]_  = ~A199 & ~A168;
  assign \new_[69685]_  = A169 & \new_[69684]_ ;
  assign \new_[69688]_  = A201 & A200;
  assign \new_[69691]_  = ~A265 & ~A203;
  assign \new_[69692]_  = \new_[69691]_  & \new_[69688]_ ;
  assign \new_[69693]_  = \new_[69692]_  & \new_[69685]_ ;
  assign \new_[69697]_  = A268 & A267;
  assign \new_[69698]_  = A266 & \new_[69697]_ ;
  assign \new_[69701]_  = ~A299 & A298;
  assign \new_[69704]_  = A301 & A300;
  assign \new_[69705]_  = \new_[69704]_  & \new_[69701]_ ;
  assign \new_[69706]_  = \new_[69705]_  & \new_[69698]_ ;
  assign \new_[69710]_  = ~A199 & ~A168;
  assign \new_[69711]_  = A169 & \new_[69710]_ ;
  assign \new_[69714]_  = A201 & A200;
  assign \new_[69717]_  = ~A265 & ~A203;
  assign \new_[69718]_  = \new_[69717]_  & \new_[69714]_ ;
  assign \new_[69719]_  = \new_[69718]_  & \new_[69711]_ ;
  assign \new_[69723]_  = A268 & A267;
  assign \new_[69724]_  = A266 & \new_[69723]_ ;
  assign \new_[69727]_  = ~A299 & A298;
  assign \new_[69730]_  = ~A302 & A300;
  assign \new_[69731]_  = \new_[69730]_  & \new_[69727]_ ;
  assign \new_[69732]_  = \new_[69731]_  & \new_[69724]_ ;
  assign \new_[69736]_  = ~A199 & ~A168;
  assign \new_[69737]_  = A169 & \new_[69736]_ ;
  assign \new_[69740]_  = A201 & A200;
  assign \new_[69743]_  = ~A265 & ~A203;
  assign \new_[69744]_  = \new_[69743]_  & \new_[69740]_ ;
  assign \new_[69745]_  = \new_[69744]_  & \new_[69737]_ ;
  assign \new_[69749]_  = A268 & A267;
  assign \new_[69750]_  = A266 & \new_[69749]_ ;
  assign \new_[69753]_  = A299 & ~A298;
  assign \new_[69756]_  = A301 & A300;
  assign \new_[69757]_  = \new_[69756]_  & \new_[69753]_ ;
  assign \new_[69758]_  = \new_[69757]_  & \new_[69750]_ ;
  assign \new_[69762]_  = ~A199 & ~A168;
  assign \new_[69763]_  = A169 & \new_[69762]_ ;
  assign \new_[69766]_  = A201 & A200;
  assign \new_[69769]_  = ~A265 & ~A203;
  assign \new_[69770]_  = \new_[69769]_  & \new_[69766]_ ;
  assign \new_[69771]_  = \new_[69770]_  & \new_[69763]_ ;
  assign \new_[69775]_  = A268 & A267;
  assign \new_[69776]_  = A266 & \new_[69775]_ ;
  assign \new_[69779]_  = A299 & ~A298;
  assign \new_[69782]_  = ~A302 & A300;
  assign \new_[69783]_  = \new_[69782]_  & \new_[69779]_ ;
  assign \new_[69784]_  = \new_[69783]_  & \new_[69776]_ ;
  assign \new_[69788]_  = ~A199 & ~A168;
  assign \new_[69789]_  = A169 & \new_[69788]_ ;
  assign \new_[69792]_  = A201 & A200;
  assign \new_[69795]_  = ~A265 & ~A203;
  assign \new_[69796]_  = \new_[69795]_  & \new_[69792]_ ;
  assign \new_[69797]_  = \new_[69796]_  & \new_[69789]_ ;
  assign \new_[69801]_  = ~A269 & A267;
  assign \new_[69802]_  = A266 & \new_[69801]_ ;
  assign \new_[69805]_  = ~A299 & A298;
  assign \new_[69808]_  = A301 & A300;
  assign \new_[69809]_  = \new_[69808]_  & \new_[69805]_ ;
  assign \new_[69810]_  = \new_[69809]_  & \new_[69802]_ ;
  assign \new_[69814]_  = ~A199 & ~A168;
  assign \new_[69815]_  = A169 & \new_[69814]_ ;
  assign \new_[69818]_  = A201 & A200;
  assign \new_[69821]_  = ~A265 & ~A203;
  assign \new_[69822]_  = \new_[69821]_  & \new_[69818]_ ;
  assign \new_[69823]_  = \new_[69822]_  & \new_[69815]_ ;
  assign \new_[69827]_  = ~A269 & A267;
  assign \new_[69828]_  = A266 & \new_[69827]_ ;
  assign \new_[69831]_  = ~A299 & A298;
  assign \new_[69834]_  = ~A302 & A300;
  assign \new_[69835]_  = \new_[69834]_  & \new_[69831]_ ;
  assign \new_[69836]_  = \new_[69835]_  & \new_[69828]_ ;
  assign \new_[69840]_  = ~A199 & ~A168;
  assign \new_[69841]_  = A169 & \new_[69840]_ ;
  assign \new_[69844]_  = A201 & A200;
  assign \new_[69847]_  = ~A265 & ~A203;
  assign \new_[69848]_  = \new_[69847]_  & \new_[69844]_ ;
  assign \new_[69849]_  = \new_[69848]_  & \new_[69841]_ ;
  assign \new_[69853]_  = ~A269 & A267;
  assign \new_[69854]_  = A266 & \new_[69853]_ ;
  assign \new_[69857]_  = A299 & ~A298;
  assign \new_[69860]_  = A301 & A300;
  assign \new_[69861]_  = \new_[69860]_  & \new_[69857]_ ;
  assign \new_[69862]_  = \new_[69861]_  & \new_[69854]_ ;
  assign \new_[69866]_  = ~A199 & ~A168;
  assign \new_[69867]_  = A169 & \new_[69866]_ ;
  assign \new_[69870]_  = A201 & A200;
  assign \new_[69873]_  = ~A265 & ~A203;
  assign \new_[69874]_  = \new_[69873]_  & \new_[69870]_ ;
  assign \new_[69875]_  = \new_[69874]_  & \new_[69867]_ ;
  assign \new_[69879]_  = ~A269 & A267;
  assign \new_[69880]_  = A266 & \new_[69879]_ ;
  assign \new_[69883]_  = A299 & ~A298;
  assign \new_[69886]_  = ~A302 & A300;
  assign \new_[69887]_  = \new_[69886]_  & \new_[69883]_ ;
  assign \new_[69888]_  = \new_[69887]_  & \new_[69880]_ ;
  assign \new_[69892]_  = ~A199 & ~A168;
  assign \new_[69893]_  = A169 & \new_[69892]_ ;
  assign \new_[69896]_  = A201 & A200;
  assign \new_[69899]_  = A265 & ~A203;
  assign \new_[69900]_  = \new_[69899]_  & \new_[69896]_ ;
  assign \new_[69901]_  = \new_[69900]_  & \new_[69893]_ ;
  assign \new_[69905]_  = A268 & A267;
  assign \new_[69906]_  = ~A266 & \new_[69905]_ ;
  assign \new_[69909]_  = ~A299 & A298;
  assign \new_[69912]_  = A301 & A300;
  assign \new_[69913]_  = \new_[69912]_  & \new_[69909]_ ;
  assign \new_[69914]_  = \new_[69913]_  & \new_[69906]_ ;
  assign \new_[69918]_  = ~A199 & ~A168;
  assign \new_[69919]_  = A169 & \new_[69918]_ ;
  assign \new_[69922]_  = A201 & A200;
  assign \new_[69925]_  = A265 & ~A203;
  assign \new_[69926]_  = \new_[69925]_  & \new_[69922]_ ;
  assign \new_[69927]_  = \new_[69926]_  & \new_[69919]_ ;
  assign \new_[69931]_  = A268 & A267;
  assign \new_[69932]_  = ~A266 & \new_[69931]_ ;
  assign \new_[69935]_  = ~A299 & A298;
  assign \new_[69938]_  = ~A302 & A300;
  assign \new_[69939]_  = \new_[69938]_  & \new_[69935]_ ;
  assign \new_[69940]_  = \new_[69939]_  & \new_[69932]_ ;
  assign \new_[69944]_  = ~A199 & ~A168;
  assign \new_[69945]_  = A169 & \new_[69944]_ ;
  assign \new_[69948]_  = A201 & A200;
  assign \new_[69951]_  = A265 & ~A203;
  assign \new_[69952]_  = \new_[69951]_  & \new_[69948]_ ;
  assign \new_[69953]_  = \new_[69952]_  & \new_[69945]_ ;
  assign \new_[69957]_  = A268 & A267;
  assign \new_[69958]_  = ~A266 & \new_[69957]_ ;
  assign \new_[69961]_  = A299 & ~A298;
  assign \new_[69964]_  = A301 & A300;
  assign \new_[69965]_  = \new_[69964]_  & \new_[69961]_ ;
  assign \new_[69966]_  = \new_[69965]_  & \new_[69958]_ ;
  assign \new_[69970]_  = ~A199 & ~A168;
  assign \new_[69971]_  = A169 & \new_[69970]_ ;
  assign \new_[69974]_  = A201 & A200;
  assign \new_[69977]_  = A265 & ~A203;
  assign \new_[69978]_  = \new_[69977]_  & \new_[69974]_ ;
  assign \new_[69979]_  = \new_[69978]_  & \new_[69971]_ ;
  assign \new_[69983]_  = A268 & A267;
  assign \new_[69984]_  = ~A266 & \new_[69983]_ ;
  assign \new_[69987]_  = A299 & ~A298;
  assign \new_[69990]_  = ~A302 & A300;
  assign \new_[69991]_  = \new_[69990]_  & \new_[69987]_ ;
  assign \new_[69992]_  = \new_[69991]_  & \new_[69984]_ ;
  assign \new_[69996]_  = ~A199 & ~A168;
  assign \new_[69997]_  = A169 & \new_[69996]_ ;
  assign \new_[70000]_  = A201 & A200;
  assign \new_[70003]_  = A265 & ~A203;
  assign \new_[70004]_  = \new_[70003]_  & \new_[70000]_ ;
  assign \new_[70005]_  = \new_[70004]_  & \new_[69997]_ ;
  assign \new_[70009]_  = ~A269 & A267;
  assign \new_[70010]_  = ~A266 & \new_[70009]_ ;
  assign \new_[70013]_  = ~A299 & A298;
  assign \new_[70016]_  = A301 & A300;
  assign \new_[70017]_  = \new_[70016]_  & \new_[70013]_ ;
  assign \new_[70018]_  = \new_[70017]_  & \new_[70010]_ ;
  assign \new_[70022]_  = ~A199 & ~A168;
  assign \new_[70023]_  = A169 & \new_[70022]_ ;
  assign \new_[70026]_  = A201 & A200;
  assign \new_[70029]_  = A265 & ~A203;
  assign \new_[70030]_  = \new_[70029]_  & \new_[70026]_ ;
  assign \new_[70031]_  = \new_[70030]_  & \new_[70023]_ ;
  assign \new_[70035]_  = ~A269 & A267;
  assign \new_[70036]_  = ~A266 & \new_[70035]_ ;
  assign \new_[70039]_  = ~A299 & A298;
  assign \new_[70042]_  = ~A302 & A300;
  assign \new_[70043]_  = \new_[70042]_  & \new_[70039]_ ;
  assign \new_[70044]_  = \new_[70043]_  & \new_[70036]_ ;
  assign \new_[70048]_  = ~A199 & ~A168;
  assign \new_[70049]_  = A169 & \new_[70048]_ ;
  assign \new_[70052]_  = A201 & A200;
  assign \new_[70055]_  = A265 & ~A203;
  assign \new_[70056]_  = \new_[70055]_  & \new_[70052]_ ;
  assign \new_[70057]_  = \new_[70056]_  & \new_[70049]_ ;
  assign \new_[70061]_  = ~A269 & A267;
  assign \new_[70062]_  = ~A266 & \new_[70061]_ ;
  assign \new_[70065]_  = A299 & ~A298;
  assign \new_[70068]_  = A301 & A300;
  assign \new_[70069]_  = \new_[70068]_  & \new_[70065]_ ;
  assign \new_[70070]_  = \new_[70069]_  & \new_[70062]_ ;
  assign \new_[70074]_  = ~A199 & ~A168;
  assign \new_[70075]_  = A169 & \new_[70074]_ ;
  assign \new_[70078]_  = A201 & A200;
  assign \new_[70081]_  = A265 & ~A203;
  assign \new_[70082]_  = \new_[70081]_  & \new_[70078]_ ;
  assign \new_[70083]_  = \new_[70082]_  & \new_[70075]_ ;
  assign \new_[70087]_  = ~A269 & A267;
  assign \new_[70088]_  = ~A266 & \new_[70087]_ ;
  assign \new_[70091]_  = A299 & ~A298;
  assign \new_[70094]_  = ~A302 & A300;
  assign \new_[70095]_  = \new_[70094]_  & \new_[70091]_ ;
  assign \new_[70096]_  = \new_[70095]_  & \new_[70088]_ ;
  assign \new_[70100]_  = A199 & ~A168;
  assign \new_[70101]_  = A169 & \new_[70100]_ ;
  assign \new_[70104]_  = A201 & ~A200;
  assign \new_[70107]_  = ~A265 & A202;
  assign \new_[70108]_  = \new_[70107]_  & \new_[70104]_ ;
  assign \new_[70109]_  = \new_[70108]_  & \new_[70101]_ ;
  assign \new_[70113]_  = A268 & A267;
  assign \new_[70114]_  = A266 & \new_[70113]_ ;
  assign \new_[70117]_  = ~A299 & A298;
  assign \new_[70120]_  = A301 & A300;
  assign \new_[70121]_  = \new_[70120]_  & \new_[70117]_ ;
  assign \new_[70122]_  = \new_[70121]_  & \new_[70114]_ ;
  assign \new_[70126]_  = A199 & ~A168;
  assign \new_[70127]_  = A169 & \new_[70126]_ ;
  assign \new_[70130]_  = A201 & ~A200;
  assign \new_[70133]_  = ~A265 & A202;
  assign \new_[70134]_  = \new_[70133]_  & \new_[70130]_ ;
  assign \new_[70135]_  = \new_[70134]_  & \new_[70127]_ ;
  assign \new_[70139]_  = A268 & A267;
  assign \new_[70140]_  = A266 & \new_[70139]_ ;
  assign \new_[70143]_  = ~A299 & A298;
  assign \new_[70146]_  = ~A302 & A300;
  assign \new_[70147]_  = \new_[70146]_  & \new_[70143]_ ;
  assign \new_[70148]_  = \new_[70147]_  & \new_[70140]_ ;
  assign \new_[70152]_  = A199 & ~A168;
  assign \new_[70153]_  = A169 & \new_[70152]_ ;
  assign \new_[70156]_  = A201 & ~A200;
  assign \new_[70159]_  = ~A265 & A202;
  assign \new_[70160]_  = \new_[70159]_  & \new_[70156]_ ;
  assign \new_[70161]_  = \new_[70160]_  & \new_[70153]_ ;
  assign \new_[70165]_  = A268 & A267;
  assign \new_[70166]_  = A266 & \new_[70165]_ ;
  assign \new_[70169]_  = A299 & ~A298;
  assign \new_[70172]_  = A301 & A300;
  assign \new_[70173]_  = \new_[70172]_  & \new_[70169]_ ;
  assign \new_[70174]_  = \new_[70173]_  & \new_[70166]_ ;
  assign \new_[70178]_  = A199 & ~A168;
  assign \new_[70179]_  = A169 & \new_[70178]_ ;
  assign \new_[70182]_  = A201 & ~A200;
  assign \new_[70185]_  = ~A265 & A202;
  assign \new_[70186]_  = \new_[70185]_  & \new_[70182]_ ;
  assign \new_[70187]_  = \new_[70186]_  & \new_[70179]_ ;
  assign \new_[70191]_  = A268 & A267;
  assign \new_[70192]_  = A266 & \new_[70191]_ ;
  assign \new_[70195]_  = A299 & ~A298;
  assign \new_[70198]_  = ~A302 & A300;
  assign \new_[70199]_  = \new_[70198]_  & \new_[70195]_ ;
  assign \new_[70200]_  = \new_[70199]_  & \new_[70192]_ ;
  assign \new_[70204]_  = A199 & ~A168;
  assign \new_[70205]_  = A169 & \new_[70204]_ ;
  assign \new_[70208]_  = A201 & ~A200;
  assign \new_[70211]_  = ~A265 & A202;
  assign \new_[70212]_  = \new_[70211]_  & \new_[70208]_ ;
  assign \new_[70213]_  = \new_[70212]_  & \new_[70205]_ ;
  assign \new_[70217]_  = ~A269 & A267;
  assign \new_[70218]_  = A266 & \new_[70217]_ ;
  assign \new_[70221]_  = ~A299 & A298;
  assign \new_[70224]_  = A301 & A300;
  assign \new_[70225]_  = \new_[70224]_  & \new_[70221]_ ;
  assign \new_[70226]_  = \new_[70225]_  & \new_[70218]_ ;
  assign \new_[70230]_  = A199 & ~A168;
  assign \new_[70231]_  = A169 & \new_[70230]_ ;
  assign \new_[70234]_  = A201 & ~A200;
  assign \new_[70237]_  = ~A265 & A202;
  assign \new_[70238]_  = \new_[70237]_  & \new_[70234]_ ;
  assign \new_[70239]_  = \new_[70238]_  & \new_[70231]_ ;
  assign \new_[70243]_  = ~A269 & A267;
  assign \new_[70244]_  = A266 & \new_[70243]_ ;
  assign \new_[70247]_  = ~A299 & A298;
  assign \new_[70250]_  = ~A302 & A300;
  assign \new_[70251]_  = \new_[70250]_  & \new_[70247]_ ;
  assign \new_[70252]_  = \new_[70251]_  & \new_[70244]_ ;
  assign \new_[70256]_  = A199 & ~A168;
  assign \new_[70257]_  = A169 & \new_[70256]_ ;
  assign \new_[70260]_  = A201 & ~A200;
  assign \new_[70263]_  = ~A265 & A202;
  assign \new_[70264]_  = \new_[70263]_  & \new_[70260]_ ;
  assign \new_[70265]_  = \new_[70264]_  & \new_[70257]_ ;
  assign \new_[70269]_  = ~A269 & A267;
  assign \new_[70270]_  = A266 & \new_[70269]_ ;
  assign \new_[70273]_  = A299 & ~A298;
  assign \new_[70276]_  = A301 & A300;
  assign \new_[70277]_  = \new_[70276]_  & \new_[70273]_ ;
  assign \new_[70278]_  = \new_[70277]_  & \new_[70270]_ ;
  assign \new_[70282]_  = A199 & ~A168;
  assign \new_[70283]_  = A169 & \new_[70282]_ ;
  assign \new_[70286]_  = A201 & ~A200;
  assign \new_[70289]_  = ~A265 & A202;
  assign \new_[70290]_  = \new_[70289]_  & \new_[70286]_ ;
  assign \new_[70291]_  = \new_[70290]_  & \new_[70283]_ ;
  assign \new_[70295]_  = ~A269 & A267;
  assign \new_[70296]_  = A266 & \new_[70295]_ ;
  assign \new_[70299]_  = A299 & ~A298;
  assign \new_[70302]_  = ~A302 & A300;
  assign \new_[70303]_  = \new_[70302]_  & \new_[70299]_ ;
  assign \new_[70304]_  = \new_[70303]_  & \new_[70296]_ ;
  assign \new_[70308]_  = A199 & ~A168;
  assign \new_[70309]_  = A169 & \new_[70308]_ ;
  assign \new_[70312]_  = A201 & ~A200;
  assign \new_[70315]_  = A265 & A202;
  assign \new_[70316]_  = \new_[70315]_  & \new_[70312]_ ;
  assign \new_[70317]_  = \new_[70316]_  & \new_[70309]_ ;
  assign \new_[70321]_  = A268 & A267;
  assign \new_[70322]_  = ~A266 & \new_[70321]_ ;
  assign \new_[70325]_  = ~A299 & A298;
  assign \new_[70328]_  = A301 & A300;
  assign \new_[70329]_  = \new_[70328]_  & \new_[70325]_ ;
  assign \new_[70330]_  = \new_[70329]_  & \new_[70322]_ ;
  assign \new_[70334]_  = A199 & ~A168;
  assign \new_[70335]_  = A169 & \new_[70334]_ ;
  assign \new_[70338]_  = A201 & ~A200;
  assign \new_[70341]_  = A265 & A202;
  assign \new_[70342]_  = \new_[70341]_  & \new_[70338]_ ;
  assign \new_[70343]_  = \new_[70342]_  & \new_[70335]_ ;
  assign \new_[70347]_  = A268 & A267;
  assign \new_[70348]_  = ~A266 & \new_[70347]_ ;
  assign \new_[70351]_  = ~A299 & A298;
  assign \new_[70354]_  = ~A302 & A300;
  assign \new_[70355]_  = \new_[70354]_  & \new_[70351]_ ;
  assign \new_[70356]_  = \new_[70355]_  & \new_[70348]_ ;
  assign \new_[70360]_  = A199 & ~A168;
  assign \new_[70361]_  = A169 & \new_[70360]_ ;
  assign \new_[70364]_  = A201 & ~A200;
  assign \new_[70367]_  = A265 & A202;
  assign \new_[70368]_  = \new_[70367]_  & \new_[70364]_ ;
  assign \new_[70369]_  = \new_[70368]_  & \new_[70361]_ ;
  assign \new_[70373]_  = A268 & A267;
  assign \new_[70374]_  = ~A266 & \new_[70373]_ ;
  assign \new_[70377]_  = A299 & ~A298;
  assign \new_[70380]_  = A301 & A300;
  assign \new_[70381]_  = \new_[70380]_  & \new_[70377]_ ;
  assign \new_[70382]_  = \new_[70381]_  & \new_[70374]_ ;
  assign \new_[70386]_  = A199 & ~A168;
  assign \new_[70387]_  = A169 & \new_[70386]_ ;
  assign \new_[70390]_  = A201 & ~A200;
  assign \new_[70393]_  = A265 & A202;
  assign \new_[70394]_  = \new_[70393]_  & \new_[70390]_ ;
  assign \new_[70395]_  = \new_[70394]_  & \new_[70387]_ ;
  assign \new_[70399]_  = A268 & A267;
  assign \new_[70400]_  = ~A266 & \new_[70399]_ ;
  assign \new_[70403]_  = A299 & ~A298;
  assign \new_[70406]_  = ~A302 & A300;
  assign \new_[70407]_  = \new_[70406]_  & \new_[70403]_ ;
  assign \new_[70408]_  = \new_[70407]_  & \new_[70400]_ ;
  assign \new_[70412]_  = A199 & ~A168;
  assign \new_[70413]_  = A169 & \new_[70412]_ ;
  assign \new_[70416]_  = A201 & ~A200;
  assign \new_[70419]_  = A265 & A202;
  assign \new_[70420]_  = \new_[70419]_  & \new_[70416]_ ;
  assign \new_[70421]_  = \new_[70420]_  & \new_[70413]_ ;
  assign \new_[70425]_  = ~A269 & A267;
  assign \new_[70426]_  = ~A266 & \new_[70425]_ ;
  assign \new_[70429]_  = ~A299 & A298;
  assign \new_[70432]_  = A301 & A300;
  assign \new_[70433]_  = \new_[70432]_  & \new_[70429]_ ;
  assign \new_[70434]_  = \new_[70433]_  & \new_[70426]_ ;
  assign \new_[70438]_  = A199 & ~A168;
  assign \new_[70439]_  = A169 & \new_[70438]_ ;
  assign \new_[70442]_  = A201 & ~A200;
  assign \new_[70445]_  = A265 & A202;
  assign \new_[70446]_  = \new_[70445]_  & \new_[70442]_ ;
  assign \new_[70447]_  = \new_[70446]_  & \new_[70439]_ ;
  assign \new_[70451]_  = ~A269 & A267;
  assign \new_[70452]_  = ~A266 & \new_[70451]_ ;
  assign \new_[70455]_  = ~A299 & A298;
  assign \new_[70458]_  = ~A302 & A300;
  assign \new_[70459]_  = \new_[70458]_  & \new_[70455]_ ;
  assign \new_[70460]_  = \new_[70459]_  & \new_[70452]_ ;
  assign \new_[70464]_  = A199 & ~A168;
  assign \new_[70465]_  = A169 & \new_[70464]_ ;
  assign \new_[70468]_  = A201 & ~A200;
  assign \new_[70471]_  = A265 & A202;
  assign \new_[70472]_  = \new_[70471]_  & \new_[70468]_ ;
  assign \new_[70473]_  = \new_[70472]_  & \new_[70465]_ ;
  assign \new_[70477]_  = ~A269 & A267;
  assign \new_[70478]_  = ~A266 & \new_[70477]_ ;
  assign \new_[70481]_  = A299 & ~A298;
  assign \new_[70484]_  = A301 & A300;
  assign \new_[70485]_  = \new_[70484]_  & \new_[70481]_ ;
  assign \new_[70486]_  = \new_[70485]_  & \new_[70478]_ ;
  assign \new_[70490]_  = A199 & ~A168;
  assign \new_[70491]_  = A169 & \new_[70490]_ ;
  assign \new_[70494]_  = A201 & ~A200;
  assign \new_[70497]_  = A265 & A202;
  assign \new_[70498]_  = \new_[70497]_  & \new_[70494]_ ;
  assign \new_[70499]_  = \new_[70498]_  & \new_[70491]_ ;
  assign \new_[70503]_  = ~A269 & A267;
  assign \new_[70504]_  = ~A266 & \new_[70503]_ ;
  assign \new_[70507]_  = A299 & ~A298;
  assign \new_[70510]_  = ~A302 & A300;
  assign \new_[70511]_  = \new_[70510]_  & \new_[70507]_ ;
  assign \new_[70512]_  = \new_[70511]_  & \new_[70504]_ ;
  assign \new_[70516]_  = A199 & ~A168;
  assign \new_[70517]_  = A169 & \new_[70516]_ ;
  assign \new_[70520]_  = A201 & ~A200;
  assign \new_[70523]_  = ~A265 & ~A203;
  assign \new_[70524]_  = \new_[70523]_  & \new_[70520]_ ;
  assign \new_[70525]_  = \new_[70524]_  & \new_[70517]_ ;
  assign \new_[70529]_  = A268 & A267;
  assign \new_[70530]_  = A266 & \new_[70529]_ ;
  assign \new_[70533]_  = ~A299 & A298;
  assign \new_[70536]_  = A301 & A300;
  assign \new_[70537]_  = \new_[70536]_  & \new_[70533]_ ;
  assign \new_[70538]_  = \new_[70537]_  & \new_[70530]_ ;
  assign \new_[70542]_  = A199 & ~A168;
  assign \new_[70543]_  = A169 & \new_[70542]_ ;
  assign \new_[70546]_  = A201 & ~A200;
  assign \new_[70549]_  = ~A265 & ~A203;
  assign \new_[70550]_  = \new_[70549]_  & \new_[70546]_ ;
  assign \new_[70551]_  = \new_[70550]_  & \new_[70543]_ ;
  assign \new_[70555]_  = A268 & A267;
  assign \new_[70556]_  = A266 & \new_[70555]_ ;
  assign \new_[70559]_  = ~A299 & A298;
  assign \new_[70562]_  = ~A302 & A300;
  assign \new_[70563]_  = \new_[70562]_  & \new_[70559]_ ;
  assign \new_[70564]_  = \new_[70563]_  & \new_[70556]_ ;
  assign \new_[70568]_  = A199 & ~A168;
  assign \new_[70569]_  = A169 & \new_[70568]_ ;
  assign \new_[70572]_  = A201 & ~A200;
  assign \new_[70575]_  = ~A265 & ~A203;
  assign \new_[70576]_  = \new_[70575]_  & \new_[70572]_ ;
  assign \new_[70577]_  = \new_[70576]_  & \new_[70569]_ ;
  assign \new_[70581]_  = A268 & A267;
  assign \new_[70582]_  = A266 & \new_[70581]_ ;
  assign \new_[70585]_  = A299 & ~A298;
  assign \new_[70588]_  = A301 & A300;
  assign \new_[70589]_  = \new_[70588]_  & \new_[70585]_ ;
  assign \new_[70590]_  = \new_[70589]_  & \new_[70582]_ ;
  assign \new_[70594]_  = A199 & ~A168;
  assign \new_[70595]_  = A169 & \new_[70594]_ ;
  assign \new_[70598]_  = A201 & ~A200;
  assign \new_[70601]_  = ~A265 & ~A203;
  assign \new_[70602]_  = \new_[70601]_  & \new_[70598]_ ;
  assign \new_[70603]_  = \new_[70602]_  & \new_[70595]_ ;
  assign \new_[70607]_  = A268 & A267;
  assign \new_[70608]_  = A266 & \new_[70607]_ ;
  assign \new_[70611]_  = A299 & ~A298;
  assign \new_[70614]_  = ~A302 & A300;
  assign \new_[70615]_  = \new_[70614]_  & \new_[70611]_ ;
  assign \new_[70616]_  = \new_[70615]_  & \new_[70608]_ ;
  assign \new_[70620]_  = A199 & ~A168;
  assign \new_[70621]_  = A169 & \new_[70620]_ ;
  assign \new_[70624]_  = A201 & ~A200;
  assign \new_[70627]_  = ~A265 & ~A203;
  assign \new_[70628]_  = \new_[70627]_  & \new_[70624]_ ;
  assign \new_[70629]_  = \new_[70628]_  & \new_[70621]_ ;
  assign \new_[70633]_  = ~A269 & A267;
  assign \new_[70634]_  = A266 & \new_[70633]_ ;
  assign \new_[70637]_  = ~A299 & A298;
  assign \new_[70640]_  = A301 & A300;
  assign \new_[70641]_  = \new_[70640]_  & \new_[70637]_ ;
  assign \new_[70642]_  = \new_[70641]_  & \new_[70634]_ ;
  assign \new_[70646]_  = A199 & ~A168;
  assign \new_[70647]_  = A169 & \new_[70646]_ ;
  assign \new_[70650]_  = A201 & ~A200;
  assign \new_[70653]_  = ~A265 & ~A203;
  assign \new_[70654]_  = \new_[70653]_  & \new_[70650]_ ;
  assign \new_[70655]_  = \new_[70654]_  & \new_[70647]_ ;
  assign \new_[70659]_  = ~A269 & A267;
  assign \new_[70660]_  = A266 & \new_[70659]_ ;
  assign \new_[70663]_  = ~A299 & A298;
  assign \new_[70666]_  = ~A302 & A300;
  assign \new_[70667]_  = \new_[70666]_  & \new_[70663]_ ;
  assign \new_[70668]_  = \new_[70667]_  & \new_[70660]_ ;
  assign \new_[70672]_  = A199 & ~A168;
  assign \new_[70673]_  = A169 & \new_[70672]_ ;
  assign \new_[70676]_  = A201 & ~A200;
  assign \new_[70679]_  = ~A265 & ~A203;
  assign \new_[70680]_  = \new_[70679]_  & \new_[70676]_ ;
  assign \new_[70681]_  = \new_[70680]_  & \new_[70673]_ ;
  assign \new_[70685]_  = ~A269 & A267;
  assign \new_[70686]_  = A266 & \new_[70685]_ ;
  assign \new_[70689]_  = A299 & ~A298;
  assign \new_[70692]_  = A301 & A300;
  assign \new_[70693]_  = \new_[70692]_  & \new_[70689]_ ;
  assign \new_[70694]_  = \new_[70693]_  & \new_[70686]_ ;
  assign \new_[70698]_  = A199 & ~A168;
  assign \new_[70699]_  = A169 & \new_[70698]_ ;
  assign \new_[70702]_  = A201 & ~A200;
  assign \new_[70705]_  = ~A265 & ~A203;
  assign \new_[70706]_  = \new_[70705]_  & \new_[70702]_ ;
  assign \new_[70707]_  = \new_[70706]_  & \new_[70699]_ ;
  assign \new_[70711]_  = ~A269 & A267;
  assign \new_[70712]_  = A266 & \new_[70711]_ ;
  assign \new_[70715]_  = A299 & ~A298;
  assign \new_[70718]_  = ~A302 & A300;
  assign \new_[70719]_  = \new_[70718]_  & \new_[70715]_ ;
  assign \new_[70720]_  = \new_[70719]_  & \new_[70712]_ ;
  assign \new_[70724]_  = A199 & ~A168;
  assign \new_[70725]_  = A169 & \new_[70724]_ ;
  assign \new_[70728]_  = A201 & ~A200;
  assign \new_[70731]_  = A265 & ~A203;
  assign \new_[70732]_  = \new_[70731]_  & \new_[70728]_ ;
  assign \new_[70733]_  = \new_[70732]_  & \new_[70725]_ ;
  assign \new_[70737]_  = A268 & A267;
  assign \new_[70738]_  = ~A266 & \new_[70737]_ ;
  assign \new_[70741]_  = ~A299 & A298;
  assign \new_[70744]_  = A301 & A300;
  assign \new_[70745]_  = \new_[70744]_  & \new_[70741]_ ;
  assign \new_[70746]_  = \new_[70745]_  & \new_[70738]_ ;
  assign \new_[70750]_  = A199 & ~A168;
  assign \new_[70751]_  = A169 & \new_[70750]_ ;
  assign \new_[70754]_  = A201 & ~A200;
  assign \new_[70757]_  = A265 & ~A203;
  assign \new_[70758]_  = \new_[70757]_  & \new_[70754]_ ;
  assign \new_[70759]_  = \new_[70758]_  & \new_[70751]_ ;
  assign \new_[70763]_  = A268 & A267;
  assign \new_[70764]_  = ~A266 & \new_[70763]_ ;
  assign \new_[70767]_  = ~A299 & A298;
  assign \new_[70770]_  = ~A302 & A300;
  assign \new_[70771]_  = \new_[70770]_  & \new_[70767]_ ;
  assign \new_[70772]_  = \new_[70771]_  & \new_[70764]_ ;
  assign \new_[70776]_  = A199 & ~A168;
  assign \new_[70777]_  = A169 & \new_[70776]_ ;
  assign \new_[70780]_  = A201 & ~A200;
  assign \new_[70783]_  = A265 & ~A203;
  assign \new_[70784]_  = \new_[70783]_  & \new_[70780]_ ;
  assign \new_[70785]_  = \new_[70784]_  & \new_[70777]_ ;
  assign \new_[70789]_  = A268 & A267;
  assign \new_[70790]_  = ~A266 & \new_[70789]_ ;
  assign \new_[70793]_  = A299 & ~A298;
  assign \new_[70796]_  = A301 & A300;
  assign \new_[70797]_  = \new_[70796]_  & \new_[70793]_ ;
  assign \new_[70798]_  = \new_[70797]_  & \new_[70790]_ ;
  assign \new_[70802]_  = A199 & ~A168;
  assign \new_[70803]_  = A169 & \new_[70802]_ ;
  assign \new_[70806]_  = A201 & ~A200;
  assign \new_[70809]_  = A265 & ~A203;
  assign \new_[70810]_  = \new_[70809]_  & \new_[70806]_ ;
  assign \new_[70811]_  = \new_[70810]_  & \new_[70803]_ ;
  assign \new_[70815]_  = A268 & A267;
  assign \new_[70816]_  = ~A266 & \new_[70815]_ ;
  assign \new_[70819]_  = A299 & ~A298;
  assign \new_[70822]_  = ~A302 & A300;
  assign \new_[70823]_  = \new_[70822]_  & \new_[70819]_ ;
  assign \new_[70824]_  = \new_[70823]_  & \new_[70816]_ ;
  assign \new_[70828]_  = A199 & ~A168;
  assign \new_[70829]_  = A169 & \new_[70828]_ ;
  assign \new_[70832]_  = A201 & ~A200;
  assign \new_[70835]_  = A265 & ~A203;
  assign \new_[70836]_  = \new_[70835]_  & \new_[70832]_ ;
  assign \new_[70837]_  = \new_[70836]_  & \new_[70829]_ ;
  assign \new_[70841]_  = ~A269 & A267;
  assign \new_[70842]_  = ~A266 & \new_[70841]_ ;
  assign \new_[70845]_  = ~A299 & A298;
  assign \new_[70848]_  = A301 & A300;
  assign \new_[70849]_  = \new_[70848]_  & \new_[70845]_ ;
  assign \new_[70850]_  = \new_[70849]_  & \new_[70842]_ ;
  assign \new_[70854]_  = A199 & ~A168;
  assign \new_[70855]_  = A169 & \new_[70854]_ ;
  assign \new_[70858]_  = A201 & ~A200;
  assign \new_[70861]_  = A265 & ~A203;
  assign \new_[70862]_  = \new_[70861]_  & \new_[70858]_ ;
  assign \new_[70863]_  = \new_[70862]_  & \new_[70855]_ ;
  assign \new_[70867]_  = ~A269 & A267;
  assign \new_[70868]_  = ~A266 & \new_[70867]_ ;
  assign \new_[70871]_  = ~A299 & A298;
  assign \new_[70874]_  = ~A302 & A300;
  assign \new_[70875]_  = \new_[70874]_  & \new_[70871]_ ;
  assign \new_[70876]_  = \new_[70875]_  & \new_[70868]_ ;
  assign \new_[70880]_  = A199 & ~A168;
  assign \new_[70881]_  = A169 & \new_[70880]_ ;
  assign \new_[70884]_  = A201 & ~A200;
  assign \new_[70887]_  = A265 & ~A203;
  assign \new_[70888]_  = \new_[70887]_  & \new_[70884]_ ;
  assign \new_[70889]_  = \new_[70888]_  & \new_[70881]_ ;
  assign \new_[70893]_  = ~A269 & A267;
  assign \new_[70894]_  = ~A266 & \new_[70893]_ ;
  assign \new_[70897]_  = A299 & ~A298;
  assign \new_[70900]_  = A301 & A300;
  assign \new_[70901]_  = \new_[70900]_  & \new_[70897]_ ;
  assign \new_[70902]_  = \new_[70901]_  & \new_[70894]_ ;
  assign \new_[70906]_  = A199 & ~A168;
  assign \new_[70907]_  = A169 & \new_[70906]_ ;
  assign \new_[70910]_  = A201 & ~A200;
  assign \new_[70913]_  = A265 & ~A203;
  assign \new_[70914]_  = \new_[70913]_  & \new_[70910]_ ;
  assign \new_[70915]_  = \new_[70914]_  & \new_[70907]_ ;
  assign \new_[70919]_  = ~A269 & A267;
  assign \new_[70920]_  = ~A266 & \new_[70919]_ ;
  assign \new_[70923]_  = A299 & ~A298;
  assign \new_[70926]_  = ~A302 & A300;
  assign \new_[70927]_  = \new_[70926]_  & \new_[70923]_ ;
  assign \new_[70928]_  = \new_[70927]_  & \new_[70920]_ ;
  assign \new_[70932]_  = A168 & ~A169;
  assign \new_[70933]_  = ~A170 & \new_[70932]_ ;
  assign \new_[70936]_  = A200 & ~A199;
  assign \new_[70939]_  = ~A202 & ~A201;
  assign \new_[70940]_  = \new_[70939]_  & \new_[70936]_ ;
  assign \new_[70941]_  = \new_[70940]_  & \new_[70933]_ ;
  assign \new_[70945]_  = ~A268 & A267;
  assign \new_[70946]_  = A203 & \new_[70945]_ ;
  assign \new_[70949]_  = A300 & A269;
  assign \new_[70952]_  = A302 & ~A301;
  assign \new_[70953]_  = \new_[70952]_  & \new_[70949]_ ;
  assign \new_[70954]_  = \new_[70953]_  & \new_[70946]_ ;
  assign \new_[70958]_  = A168 & ~A169;
  assign \new_[70959]_  = ~A170 & \new_[70958]_ ;
  assign \new_[70962]_  = ~A200 & A199;
  assign \new_[70965]_  = ~A202 & ~A201;
  assign \new_[70966]_  = \new_[70965]_  & \new_[70962]_ ;
  assign \new_[70967]_  = \new_[70966]_  & \new_[70959]_ ;
  assign \new_[70971]_  = ~A268 & A267;
  assign \new_[70972]_  = A203 & \new_[70971]_ ;
  assign \new_[70975]_  = A300 & A269;
  assign \new_[70978]_  = A302 & ~A301;
  assign \new_[70979]_  = \new_[70978]_  & \new_[70975]_ ;
  assign \new_[70980]_  = \new_[70979]_  & \new_[70972]_ ;
  assign \new_[70984]_  = ~A168 & ~A169;
  assign \new_[70985]_  = ~A170 & \new_[70984]_ ;
  assign \new_[70988]_  = ~A166 & A167;
  assign \new_[70991]_  = ~A202 & A201;
  assign \new_[70992]_  = \new_[70991]_  & \new_[70988]_ ;
  assign \new_[70993]_  = \new_[70992]_  & \new_[70985]_ ;
  assign \new_[70997]_  = A268 & ~A267;
  assign \new_[70998]_  = A203 & \new_[70997]_ ;
  assign \new_[71001]_  = ~A299 & A298;
  assign \new_[71004]_  = A301 & A300;
  assign \new_[71005]_  = \new_[71004]_  & \new_[71001]_ ;
  assign \new_[71006]_  = \new_[71005]_  & \new_[70998]_ ;
  assign \new_[71010]_  = ~A168 & ~A169;
  assign \new_[71011]_  = ~A170 & \new_[71010]_ ;
  assign \new_[71014]_  = ~A166 & A167;
  assign \new_[71017]_  = ~A202 & A201;
  assign \new_[71018]_  = \new_[71017]_  & \new_[71014]_ ;
  assign \new_[71019]_  = \new_[71018]_  & \new_[71011]_ ;
  assign \new_[71023]_  = A268 & ~A267;
  assign \new_[71024]_  = A203 & \new_[71023]_ ;
  assign \new_[71027]_  = ~A299 & A298;
  assign \new_[71030]_  = ~A302 & A300;
  assign \new_[71031]_  = \new_[71030]_  & \new_[71027]_ ;
  assign \new_[71032]_  = \new_[71031]_  & \new_[71024]_ ;
  assign \new_[71036]_  = ~A168 & ~A169;
  assign \new_[71037]_  = ~A170 & \new_[71036]_ ;
  assign \new_[71040]_  = ~A166 & A167;
  assign \new_[71043]_  = ~A202 & A201;
  assign \new_[71044]_  = \new_[71043]_  & \new_[71040]_ ;
  assign \new_[71045]_  = \new_[71044]_  & \new_[71037]_ ;
  assign \new_[71049]_  = A268 & ~A267;
  assign \new_[71050]_  = A203 & \new_[71049]_ ;
  assign \new_[71053]_  = A299 & ~A298;
  assign \new_[71056]_  = A301 & A300;
  assign \new_[71057]_  = \new_[71056]_  & \new_[71053]_ ;
  assign \new_[71058]_  = \new_[71057]_  & \new_[71050]_ ;
  assign \new_[71062]_  = ~A168 & ~A169;
  assign \new_[71063]_  = ~A170 & \new_[71062]_ ;
  assign \new_[71066]_  = ~A166 & A167;
  assign \new_[71069]_  = ~A202 & A201;
  assign \new_[71070]_  = \new_[71069]_  & \new_[71066]_ ;
  assign \new_[71071]_  = \new_[71070]_  & \new_[71063]_ ;
  assign \new_[71075]_  = A268 & ~A267;
  assign \new_[71076]_  = A203 & \new_[71075]_ ;
  assign \new_[71079]_  = A299 & ~A298;
  assign \new_[71082]_  = ~A302 & A300;
  assign \new_[71083]_  = \new_[71082]_  & \new_[71079]_ ;
  assign \new_[71084]_  = \new_[71083]_  & \new_[71076]_ ;
  assign \new_[71088]_  = ~A168 & ~A169;
  assign \new_[71089]_  = ~A170 & \new_[71088]_ ;
  assign \new_[71092]_  = ~A166 & A167;
  assign \new_[71095]_  = ~A202 & A201;
  assign \new_[71096]_  = \new_[71095]_  & \new_[71092]_ ;
  assign \new_[71097]_  = \new_[71096]_  & \new_[71089]_ ;
  assign \new_[71101]_  = ~A269 & ~A267;
  assign \new_[71102]_  = A203 & \new_[71101]_ ;
  assign \new_[71105]_  = ~A299 & A298;
  assign \new_[71108]_  = A301 & A300;
  assign \new_[71109]_  = \new_[71108]_  & \new_[71105]_ ;
  assign \new_[71110]_  = \new_[71109]_  & \new_[71102]_ ;
  assign \new_[71114]_  = ~A168 & ~A169;
  assign \new_[71115]_  = ~A170 & \new_[71114]_ ;
  assign \new_[71118]_  = ~A166 & A167;
  assign \new_[71121]_  = ~A202 & A201;
  assign \new_[71122]_  = \new_[71121]_  & \new_[71118]_ ;
  assign \new_[71123]_  = \new_[71122]_  & \new_[71115]_ ;
  assign \new_[71127]_  = ~A269 & ~A267;
  assign \new_[71128]_  = A203 & \new_[71127]_ ;
  assign \new_[71131]_  = ~A299 & A298;
  assign \new_[71134]_  = ~A302 & A300;
  assign \new_[71135]_  = \new_[71134]_  & \new_[71131]_ ;
  assign \new_[71136]_  = \new_[71135]_  & \new_[71128]_ ;
  assign \new_[71140]_  = ~A168 & ~A169;
  assign \new_[71141]_  = ~A170 & \new_[71140]_ ;
  assign \new_[71144]_  = ~A166 & A167;
  assign \new_[71147]_  = ~A202 & A201;
  assign \new_[71148]_  = \new_[71147]_  & \new_[71144]_ ;
  assign \new_[71149]_  = \new_[71148]_  & \new_[71141]_ ;
  assign \new_[71153]_  = ~A269 & ~A267;
  assign \new_[71154]_  = A203 & \new_[71153]_ ;
  assign \new_[71157]_  = A299 & ~A298;
  assign \new_[71160]_  = A301 & A300;
  assign \new_[71161]_  = \new_[71160]_  & \new_[71157]_ ;
  assign \new_[71162]_  = \new_[71161]_  & \new_[71154]_ ;
  assign \new_[71166]_  = ~A168 & ~A169;
  assign \new_[71167]_  = ~A170 & \new_[71166]_ ;
  assign \new_[71170]_  = ~A166 & A167;
  assign \new_[71173]_  = ~A202 & A201;
  assign \new_[71174]_  = \new_[71173]_  & \new_[71170]_ ;
  assign \new_[71175]_  = \new_[71174]_  & \new_[71167]_ ;
  assign \new_[71179]_  = ~A269 & ~A267;
  assign \new_[71180]_  = A203 & \new_[71179]_ ;
  assign \new_[71183]_  = A299 & ~A298;
  assign \new_[71186]_  = ~A302 & A300;
  assign \new_[71187]_  = \new_[71186]_  & \new_[71183]_ ;
  assign \new_[71188]_  = \new_[71187]_  & \new_[71180]_ ;
  assign \new_[71192]_  = ~A168 & ~A169;
  assign \new_[71193]_  = ~A170 & \new_[71192]_ ;
  assign \new_[71196]_  = ~A166 & A167;
  assign \new_[71199]_  = ~A202 & A201;
  assign \new_[71200]_  = \new_[71199]_  & \new_[71196]_ ;
  assign \new_[71201]_  = \new_[71200]_  & \new_[71193]_ ;
  assign \new_[71205]_  = A266 & A265;
  assign \new_[71206]_  = A203 & \new_[71205]_ ;
  assign \new_[71209]_  = ~A299 & A298;
  assign \new_[71212]_  = A301 & A300;
  assign \new_[71213]_  = \new_[71212]_  & \new_[71209]_ ;
  assign \new_[71214]_  = \new_[71213]_  & \new_[71206]_ ;
  assign \new_[71218]_  = ~A168 & ~A169;
  assign \new_[71219]_  = ~A170 & \new_[71218]_ ;
  assign \new_[71222]_  = ~A166 & A167;
  assign \new_[71225]_  = ~A202 & A201;
  assign \new_[71226]_  = \new_[71225]_  & \new_[71222]_ ;
  assign \new_[71227]_  = \new_[71226]_  & \new_[71219]_ ;
  assign \new_[71231]_  = A266 & A265;
  assign \new_[71232]_  = A203 & \new_[71231]_ ;
  assign \new_[71235]_  = ~A299 & A298;
  assign \new_[71238]_  = ~A302 & A300;
  assign \new_[71239]_  = \new_[71238]_  & \new_[71235]_ ;
  assign \new_[71240]_  = \new_[71239]_  & \new_[71232]_ ;
  assign \new_[71244]_  = ~A168 & ~A169;
  assign \new_[71245]_  = ~A170 & \new_[71244]_ ;
  assign \new_[71248]_  = ~A166 & A167;
  assign \new_[71251]_  = ~A202 & A201;
  assign \new_[71252]_  = \new_[71251]_  & \new_[71248]_ ;
  assign \new_[71253]_  = \new_[71252]_  & \new_[71245]_ ;
  assign \new_[71257]_  = A266 & A265;
  assign \new_[71258]_  = A203 & \new_[71257]_ ;
  assign \new_[71261]_  = A299 & ~A298;
  assign \new_[71264]_  = A301 & A300;
  assign \new_[71265]_  = \new_[71264]_  & \new_[71261]_ ;
  assign \new_[71266]_  = \new_[71265]_  & \new_[71258]_ ;
  assign \new_[71270]_  = ~A168 & ~A169;
  assign \new_[71271]_  = ~A170 & \new_[71270]_ ;
  assign \new_[71274]_  = ~A166 & A167;
  assign \new_[71277]_  = ~A202 & A201;
  assign \new_[71278]_  = \new_[71277]_  & \new_[71274]_ ;
  assign \new_[71279]_  = \new_[71278]_  & \new_[71271]_ ;
  assign \new_[71283]_  = A266 & A265;
  assign \new_[71284]_  = A203 & \new_[71283]_ ;
  assign \new_[71287]_  = A299 & ~A298;
  assign \new_[71290]_  = ~A302 & A300;
  assign \new_[71291]_  = \new_[71290]_  & \new_[71287]_ ;
  assign \new_[71292]_  = \new_[71291]_  & \new_[71284]_ ;
  assign \new_[71296]_  = ~A168 & ~A169;
  assign \new_[71297]_  = ~A170 & \new_[71296]_ ;
  assign \new_[71300]_  = ~A166 & A167;
  assign \new_[71303]_  = ~A202 & A201;
  assign \new_[71304]_  = \new_[71303]_  & \new_[71300]_ ;
  assign \new_[71305]_  = \new_[71304]_  & \new_[71297]_ ;
  assign \new_[71309]_  = A266 & ~A265;
  assign \new_[71310]_  = A203 & \new_[71309]_ ;
  assign \new_[71313]_  = A268 & A267;
  assign \new_[71316]_  = A301 & ~A300;
  assign \new_[71317]_  = \new_[71316]_  & \new_[71313]_ ;
  assign \new_[71318]_  = \new_[71317]_  & \new_[71310]_ ;
  assign \new_[71322]_  = ~A168 & ~A169;
  assign \new_[71323]_  = ~A170 & \new_[71322]_ ;
  assign \new_[71326]_  = ~A166 & A167;
  assign \new_[71329]_  = ~A202 & A201;
  assign \new_[71330]_  = \new_[71329]_  & \new_[71326]_ ;
  assign \new_[71331]_  = \new_[71330]_  & \new_[71323]_ ;
  assign \new_[71335]_  = A266 & ~A265;
  assign \new_[71336]_  = A203 & \new_[71335]_ ;
  assign \new_[71339]_  = A268 & A267;
  assign \new_[71342]_  = ~A302 & ~A300;
  assign \new_[71343]_  = \new_[71342]_  & \new_[71339]_ ;
  assign \new_[71344]_  = \new_[71343]_  & \new_[71336]_ ;
  assign \new_[71348]_  = ~A168 & ~A169;
  assign \new_[71349]_  = ~A170 & \new_[71348]_ ;
  assign \new_[71352]_  = ~A166 & A167;
  assign \new_[71355]_  = ~A202 & A201;
  assign \new_[71356]_  = \new_[71355]_  & \new_[71352]_ ;
  assign \new_[71357]_  = \new_[71356]_  & \new_[71349]_ ;
  assign \new_[71361]_  = A266 & ~A265;
  assign \new_[71362]_  = A203 & \new_[71361]_ ;
  assign \new_[71365]_  = A268 & A267;
  assign \new_[71368]_  = A299 & A298;
  assign \new_[71369]_  = \new_[71368]_  & \new_[71365]_ ;
  assign \new_[71370]_  = \new_[71369]_  & \new_[71362]_ ;
  assign \new_[71374]_  = ~A168 & ~A169;
  assign \new_[71375]_  = ~A170 & \new_[71374]_ ;
  assign \new_[71378]_  = ~A166 & A167;
  assign \new_[71381]_  = ~A202 & A201;
  assign \new_[71382]_  = \new_[71381]_  & \new_[71378]_ ;
  assign \new_[71383]_  = \new_[71382]_  & \new_[71375]_ ;
  assign \new_[71387]_  = A266 & ~A265;
  assign \new_[71388]_  = A203 & \new_[71387]_ ;
  assign \new_[71391]_  = A268 & A267;
  assign \new_[71394]_  = ~A299 & ~A298;
  assign \new_[71395]_  = \new_[71394]_  & \new_[71391]_ ;
  assign \new_[71396]_  = \new_[71395]_  & \new_[71388]_ ;
  assign \new_[71400]_  = ~A168 & ~A169;
  assign \new_[71401]_  = ~A170 & \new_[71400]_ ;
  assign \new_[71404]_  = ~A166 & A167;
  assign \new_[71407]_  = ~A202 & A201;
  assign \new_[71408]_  = \new_[71407]_  & \new_[71404]_ ;
  assign \new_[71409]_  = \new_[71408]_  & \new_[71401]_ ;
  assign \new_[71413]_  = A266 & ~A265;
  assign \new_[71414]_  = A203 & \new_[71413]_ ;
  assign \new_[71417]_  = ~A269 & A267;
  assign \new_[71420]_  = A301 & ~A300;
  assign \new_[71421]_  = \new_[71420]_  & \new_[71417]_ ;
  assign \new_[71422]_  = \new_[71421]_  & \new_[71414]_ ;
  assign \new_[71426]_  = ~A168 & ~A169;
  assign \new_[71427]_  = ~A170 & \new_[71426]_ ;
  assign \new_[71430]_  = ~A166 & A167;
  assign \new_[71433]_  = ~A202 & A201;
  assign \new_[71434]_  = \new_[71433]_  & \new_[71430]_ ;
  assign \new_[71435]_  = \new_[71434]_  & \new_[71427]_ ;
  assign \new_[71439]_  = A266 & ~A265;
  assign \new_[71440]_  = A203 & \new_[71439]_ ;
  assign \new_[71443]_  = ~A269 & A267;
  assign \new_[71446]_  = ~A302 & ~A300;
  assign \new_[71447]_  = \new_[71446]_  & \new_[71443]_ ;
  assign \new_[71448]_  = \new_[71447]_  & \new_[71440]_ ;
  assign \new_[71452]_  = ~A168 & ~A169;
  assign \new_[71453]_  = ~A170 & \new_[71452]_ ;
  assign \new_[71456]_  = ~A166 & A167;
  assign \new_[71459]_  = ~A202 & A201;
  assign \new_[71460]_  = \new_[71459]_  & \new_[71456]_ ;
  assign \new_[71461]_  = \new_[71460]_  & \new_[71453]_ ;
  assign \new_[71465]_  = A266 & ~A265;
  assign \new_[71466]_  = A203 & \new_[71465]_ ;
  assign \new_[71469]_  = ~A269 & A267;
  assign \new_[71472]_  = A299 & A298;
  assign \new_[71473]_  = \new_[71472]_  & \new_[71469]_ ;
  assign \new_[71474]_  = \new_[71473]_  & \new_[71466]_ ;
  assign \new_[71478]_  = ~A168 & ~A169;
  assign \new_[71479]_  = ~A170 & \new_[71478]_ ;
  assign \new_[71482]_  = ~A166 & A167;
  assign \new_[71485]_  = ~A202 & A201;
  assign \new_[71486]_  = \new_[71485]_  & \new_[71482]_ ;
  assign \new_[71487]_  = \new_[71486]_  & \new_[71479]_ ;
  assign \new_[71491]_  = A266 & ~A265;
  assign \new_[71492]_  = A203 & \new_[71491]_ ;
  assign \new_[71495]_  = ~A269 & A267;
  assign \new_[71498]_  = ~A299 & ~A298;
  assign \new_[71499]_  = \new_[71498]_  & \new_[71495]_ ;
  assign \new_[71500]_  = \new_[71499]_  & \new_[71492]_ ;
  assign \new_[71504]_  = ~A168 & ~A169;
  assign \new_[71505]_  = ~A170 & \new_[71504]_ ;
  assign \new_[71508]_  = ~A166 & A167;
  assign \new_[71511]_  = ~A202 & A201;
  assign \new_[71512]_  = \new_[71511]_  & \new_[71508]_ ;
  assign \new_[71513]_  = \new_[71512]_  & \new_[71505]_ ;
  assign \new_[71517]_  = ~A266 & A265;
  assign \new_[71518]_  = A203 & \new_[71517]_ ;
  assign \new_[71521]_  = A268 & A267;
  assign \new_[71524]_  = A301 & ~A300;
  assign \new_[71525]_  = \new_[71524]_  & \new_[71521]_ ;
  assign \new_[71526]_  = \new_[71525]_  & \new_[71518]_ ;
  assign \new_[71530]_  = ~A168 & ~A169;
  assign \new_[71531]_  = ~A170 & \new_[71530]_ ;
  assign \new_[71534]_  = ~A166 & A167;
  assign \new_[71537]_  = ~A202 & A201;
  assign \new_[71538]_  = \new_[71537]_  & \new_[71534]_ ;
  assign \new_[71539]_  = \new_[71538]_  & \new_[71531]_ ;
  assign \new_[71543]_  = ~A266 & A265;
  assign \new_[71544]_  = A203 & \new_[71543]_ ;
  assign \new_[71547]_  = A268 & A267;
  assign \new_[71550]_  = ~A302 & ~A300;
  assign \new_[71551]_  = \new_[71550]_  & \new_[71547]_ ;
  assign \new_[71552]_  = \new_[71551]_  & \new_[71544]_ ;
  assign \new_[71556]_  = ~A168 & ~A169;
  assign \new_[71557]_  = ~A170 & \new_[71556]_ ;
  assign \new_[71560]_  = ~A166 & A167;
  assign \new_[71563]_  = ~A202 & A201;
  assign \new_[71564]_  = \new_[71563]_  & \new_[71560]_ ;
  assign \new_[71565]_  = \new_[71564]_  & \new_[71557]_ ;
  assign \new_[71569]_  = ~A266 & A265;
  assign \new_[71570]_  = A203 & \new_[71569]_ ;
  assign \new_[71573]_  = A268 & A267;
  assign \new_[71576]_  = A299 & A298;
  assign \new_[71577]_  = \new_[71576]_  & \new_[71573]_ ;
  assign \new_[71578]_  = \new_[71577]_  & \new_[71570]_ ;
  assign \new_[71582]_  = ~A168 & ~A169;
  assign \new_[71583]_  = ~A170 & \new_[71582]_ ;
  assign \new_[71586]_  = ~A166 & A167;
  assign \new_[71589]_  = ~A202 & A201;
  assign \new_[71590]_  = \new_[71589]_  & \new_[71586]_ ;
  assign \new_[71591]_  = \new_[71590]_  & \new_[71583]_ ;
  assign \new_[71595]_  = ~A266 & A265;
  assign \new_[71596]_  = A203 & \new_[71595]_ ;
  assign \new_[71599]_  = A268 & A267;
  assign \new_[71602]_  = ~A299 & ~A298;
  assign \new_[71603]_  = \new_[71602]_  & \new_[71599]_ ;
  assign \new_[71604]_  = \new_[71603]_  & \new_[71596]_ ;
  assign \new_[71608]_  = ~A168 & ~A169;
  assign \new_[71609]_  = ~A170 & \new_[71608]_ ;
  assign \new_[71612]_  = ~A166 & A167;
  assign \new_[71615]_  = ~A202 & A201;
  assign \new_[71616]_  = \new_[71615]_  & \new_[71612]_ ;
  assign \new_[71617]_  = \new_[71616]_  & \new_[71609]_ ;
  assign \new_[71621]_  = ~A266 & A265;
  assign \new_[71622]_  = A203 & \new_[71621]_ ;
  assign \new_[71625]_  = ~A269 & A267;
  assign \new_[71628]_  = A301 & ~A300;
  assign \new_[71629]_  = \new_[71628]_  & \new_[71625]_ ;
  assign \new_[71630]_  = \new_[71629]_  & \new_[71622]_ ;
  assign \new_[71634]_  = ~A168 & ~A169;
  assign \new_[71635]_  = ~A170 & \new_[71634]_ ;
  assign \new_[71638]_  = ~A166 & A167;
  assign \new_[71641]_  = ~A202 & A201;
  assign \new_[71642]_  = \new_[71641]_  & \new_[71638]_ ;
  assign \new_[71643]_  = \new_[71642]_  & \new_[71635]_ ;
  assign \new_[71647]_  = ~A266 & A265;
  assign \new_[71648]_  = A203 & \new_[71647]_ ;
  assign \new_[71651]_  = ~A269 & A267;
  assign \new_[71654]_  = ~A302 & ~A300;
  assign \new_[71655]_  = \new_[71654]_  & \new_[71651]_ ;
  assign \new_[71656]_  = \new_[71655]_  & \new_[71648]_ ;
  assign \new_[71660]_  = ~A168 & ~A169;
  assign \new_[71661]_  = ~A170 & \new_[71660]_ ;
  assign \new_[71664]_  = ~A166 & A167;
  assign \new_[71667]_  = ~A202 & A201;
  assign \new_[71668]_  = \new_[71667]_  & \new_[71664]_ ;
  assign \new_[71669]_  = \new_[71668]_  & \new_[71661]_ ;
  assign \new_[71673]_  = ~A266 & A265;
  assign \new_[71674]_  = A203 & \new_[71673]_ ;
  assign \new_[71677]_  = ~A269 & A267;
  assign \new_[71680]_  = A299 & A298;
  assign \new_[71681]_  = \new_[71680]_  & \new_[71677]_ ;
  assign \new_[71682]_  = \new_[71681]_  & \new_[71674]_ ;
  assign \new_[71686]_  = ~A168 & ~A169;
  assign \new_[71687]_  = ~A170 & \new_[71686]_ ;
  assign \new_[71690]_  = ~A166 & A167;
  assign \new_[71693]_  = ~A202 & A201;
  assign \new_[71694]_  = \new_[71693]_  & \new_[71690]_ ;
  assign \new_[71695]_  = \new_[71694]_  & \new_[71687]_ ;
  assign \new_[71699]_  = ~A266 & A265;
  assign \new_[71700]_  = A203 & \new_[71699]_ ;
  assign \new_[71703]_  = ~A269 & A267;
  assign \new_[71706]_  = ~A299 & ~A298;
  assign \new_[71707]_  = \new_[71706]_  & \new_[71703]_ ;
  assign \new_[71708]_  = \new_[71707]_  & \new_[71700]_ ;
  assign \new_[71712]_  = ~A168 & ~A169;
  assign \new_[71713]_  = ~A170 & \new_[71712]_ ;
  assign \new_[71716]_  = ~A166 & A167;
  assign \new_[71719]_  = ~A202 & A201;
  assign \new_[71720]_  = \new_[71719]_  & \new_[71716]_ ;
  assign \new_[71721]_  = \new_[71720]_  & \new_[71713]_ ;
  assign \new_[71725]_  = ~A266 & ~A265;
  assign \new_[71726]_  = A203 & \new_[71725]_ ;
  assign \new_[71729]_  = ~A299 & A298;
  assign \new_[71732]_  = A301 & A300;
  assign \new_[71733]_  = \new_[71732]_  & \new_[71729]_ ;
  assign \new_[71734]_  = \new_[71733]_  & \new_[71726]_ ;
  assign \new_[71738]_  = ~A168 & ~A169;
  assign \new_[71739]_  = ~A170 & \new_[71738]_ ;
  assign \new_[71742]_  = ~A166 & A167;
  assign \new_[71745]_  = ~A202 & A201;
  assign \new_[71746]_  = \new_[71745]_  & \new_[71742]_ ;
  assign \new_[71747]_  = \new_[71746]_  & \new_[71739]_ ;
  assign \new_[71751]_  = ~A266 & ~A265;
  assign \new_[71752]_  = A203 & \new_[71751]_ ;
  assign \new_[71755]_  = ~A299 & A298;
  assign \new_[71758]_  = ~A302 & A300;
  assign \new_[71759]_  = \new_[71758]_  & \new_[71755]_ ;
  assign \new_[71760]_  = \new_[71759]_  & \new_[71752]_ ;
  assign \new_[71764]_  = ~A168 & ~A169;
  assign \new_[71765]_  = ~A170 & \new_[71764]_ ;
  assign \new_[71768]_  = ~A166 & A167;
  assign \new_[71771]_  = ~A202 & A201;
  assign \new_[71772]_  = \new_[71771]_  & \new_[71768]_ ;
  assign \new_[71773]_  = \new_[71772]_  & \new_[71765]_ ;
  assign \new_[71777]_  = ~A266 & ~A265;
  assign \new_[71778]_  = A203 & \new_[71777]_ ;
  assign \new_[71781]_  = A299 & ~A298;
  assign \new_[71784]_  = A301 & A300;
  assign \new_[71785]_  = \new_[71784]_  & \new_[71781]_ ;
  assign \new_[71786]_  = \new_[71785]_  & \new_[71778]_ ;
  assign \new_[71790]_  = ~A168 & ~A169;
  assign \new_[71791]_  = ~A170 & \new_[71790]_ ;
  assign \new_[71794]_  = ~A166 & A167;
  assign \new_[71797]_  = ~A202 & A201;
  assign \new_[71798]_  = \new_[71797]_  & \new_[71794]_ ;
  assign \new_[71799]_  = \new_[71798]_  & \new_[71791]_ ;
  assign \new_[71803]_  = ~A266 & ~A265;
  assign \new_[71804]_  = A203 & \new_[71803]_ ;
  assign \new_[71807]_  = A299 & ~A298;
  assign \new_[71810]_  = ~A302 & A300;
  assign \new_[71811]_  = \new_[71810]_  & \new_[71807]_ ;
  assign \new_[71812]_  = \new_[71811]_  & \new_[71804]_ ;
  assign \new_[71816]_  = ~A168 & ~A169;
  assign \new_[71817]_  = ~A170 & \new_[71816]_ ;
  assign \new_[71820]_  = ~A166 & A167;
  assign \new_[71823]_  = A202 & ~A201;
  assign \new_[71824]_  = \new_[71823]_  & \new_[71820]_ ;
  assign \new_[71825]_  = \new_[71824]_  & \new_[71817]_ ;
  assign \new_[71829]_  = A269 & ~A268;
  assign \new_[71830]_  = A267 & \new_[71829]_ ;
  assign \new_[71833]_  = ~A299 & A298;
  assign \new_[71836]_  = A301 & A300;
  assign \new_[71837]_  = \new_[71836]_  & \new_[71833]_ ;
  assign \new_[71838]_  = \new_[71837]_  & \new_[71830]_ ;
  assign \new_[71842]_  = ~A168 & ~A169;
  assign \new_[71843]_  = ~A170 & \new_[71842]_ ;
  assign \new_[71846]_  = ~A166 & A167;
  assign \new_[71849]_  = A202 & ~A201;
  assign \new_[71850]_  = \new_[71849]_  & \new_[71846]_ ;
  assign \new_[71851]_  = \new_[71850]_  & \new_[71843]_ ;
  assign \new_[71855]_  = A269 & ~A268;
  assign \new_[71856]_  = A267 & \new_[71855]_ ;
  assign \new_[71859]_  = ~A299 & A298;
  assign \new_[71862]_  = ~A302 & A300;
  assign \new_[71863]_  = \new_[71862]_  & \new_[71859]_ ;
  assign \new_[71864]_  = \new_[71863]_  & \new_[71856]_ ;
  assign \new_[71868]_  = ~A168 & ~A169;
  assign \new_[71869]_  = ~A170 & \new_[71868]_ ;
  assign \new_[71872]_  = ~A166 & A167;
  assign \new_[71875]_  = A202 & ~A201;
  assign \new_[71876]_  = \new_[71875]_  & \new_[71872]_ ;
  assign \new_[71877]_  = \new_[71876]_  & \new_[71869]_ ;
  assign \new_[71881]_  = A269 & ~A268;
  assign \new_[71882]_  = A267 & \new_[71881]_ ;
  assign \new_[71885]_  = A299 & ~A298;
  assign \new_[71888]_  = A301 & A300;
  assign \new_[71889]_  = \new_[71888]_  & \new_[71885]_ ;
  assign \new_[71890]_  = \new_[71889]_  & \new_[71882]_ ;
  assign \new_[71894]_  = ~A168 & ~A169;
  assign \new_[71895]_  = ~A170 & \new_[71894]_ ;
  assign \new_[71898]_  = ~A166 & A167;
  assign \new_[71901]_  = A202 & ~A201;
  assign \new_[71902]_  = \new_[71901]_  & \new_[71898]_ ;
  assign \new_[71903]_  = \new_[71902]_  & \new_[71895]_ ;
  assign \new_[71907]_  = A269 & ~A268;
  assign \new_[71908]_  = A267 & \new_[71907]_ ;
  assign \new_[71911]_  = A299 & ~A298;
  assign \new_[71914]_  = ~A302 & A300;
  assign \new_[71915]_  = \new_[71914]_  & \new_[71911]_ ;
  assign \new_[71916]_  = \new_[71915]_  & \new_[71908]_ ;
  assign \new_[71920]_  = ~A168 & ~A169;
  assign \new_[71921]_  = ~A170 & \new_[71920]_ ;
  assign \new_[71924]_  = ~A166 & A167;
  assign \new_[71927]_  = A202 & ~A201;
  assign \new_[71928]_  = \new_[71927]_  & \new_[71924]_ ;
  assign \new_[71929]_  = \new_[71928]_  & \new_[71921]_ ;
  assign \new_[71933]_  = A298 & A268;
  assign \new_[71934]_  = ~A267 & \new_[71933]_ ;
  assign \new_[71937]_  = ~A300 & ~A299;
  assign \new_[71940]_  = A302 & ~A301;
  assign \new_[71941]_  = \new_[71940]_  & \new_[71937]_ ;
  assign \new_[71942]_  = \new_[71941]_  & \new_[71934]_ ;
  assign \new_[71946]_  = ~A168 & ~A169;
  assign \new_[71947]_  = ~A170 & \new_[71946]_ ;
  assign \new_[71950]_  = ~A166 & A167;
  assign \new_[71953]_  = A202 & ~A201;
  assign \new_[71954]_  = \new_[71953]_  & \new_[71950]_ ;
  assign \new_[71955]_  = \new_[71954]_  & \new_[71947]_ ;
  assign \new_[71959]_  = ~A298 & A268;
  assign \new_[71960]_  = ~A267 & \new_[71959]_ ;
  assign \new_[71963]_  = ~A300 & A299;
  assign \new_[71966]_  = A302 & ~A301;
  assign \new_[71967]_  = \new_[71966]_  & \new_[71963]_ ;
  assign \new_[71968]_  = \new_[71967]_  & \new_[71960]_ ;
  assign \new_[71972]_  = ~A168 & ~A169;
  assign \new_[71973]_  = ~A170 & \new_[71972]_ ;
  assign \new_[71976]_  = ~A166 & A167;
  assign \new_[71979]_  = A202 & ~A201;
  assign \new_[71980]_  = \new_[71979]_  & \new_[71976]_ ;
  assign \new_[71981]_  = \new_[71980]_  & \new_[71973]_ ;
  assign \new_[71985]_  = A298 & ~A269;
  assign \new_[71986]_  = ~A267 & \new_[71985]_ ;
  assign \new_[71989]_  = ~A300 & ~A299;
  assign \new_[71992]_  = A302 & ~A301;
  assign \new_[71993]_  = \new_[71992]_  & \new_[71989]_ ;
  assign \new_[71994]_  = \new_[71993]_  & \new_[71986]_ ;
  assign \new_[71998]_  = ~A168 & ~A169;
  assign \new_[71999]_  = ~A170 & \new_[71998]_ ;
  assign \new_[72002]_  = ~A166 & A167;
  assign \new_[72005]_  = A202 & ~A201;
  assign \new_[72006]_  = \new_[72005]_  & \new_[72002]_ ;
  assign \new_[72007]_  = \new_[72006]_  & \new_[71999]_ ;
  assign \new_[72011]_  = ~A298 & ~A269;
  assign \new_[72012]_  = ~A267 & \new_[72011]_ ;
  assign \new_[72015]_  = ~A300 & A299;
  assign \new_[72018]_  = A302 & ~A301;
  assign \new_[72019]_  = \new_[72018]_  & \new_[72015]_ ;
  assign \new_[72020]_  = \new_[72019]_  & \new_[72012]_ ;
  assign \new_[72024]_  = ~A168 & ~A169;
  assign \new_[72025]_  = ~A170 & \new_[72024]_ ;
  assign \new_[72028]_  = ~A166 & A167;
  assign \new_[72031]_  = A202 & ~A201;
  assign \new_[72032]_  = \new_[72031]_  & \new_[72028]_ ;
  assign \new_[72033]_  = \new_[72032]_  & \new_[72025]_ ;
  assign \new_[72037]_  = A298 & A266;
  assign \new_[72038]_  = A265 & \new_[72037]_ ;
  assign \new_[72041]_  = ~A300 & ~A299;
  assign \new_[72044]_  = A302 & ~A301;
  assign \new_[72045]_  = \new_[72044]_  & \new_[72041]_ ;
  assign \new_[72046]_  = \new_[72045]_  & \new_[72038]_ ;
  assign \new_[72050]_  = ~A168 & ~A169;
  assign \new_[72051]_  = ~A170 & \new_[72050]_ ;
  assign \new_[72054]_  = ~A166 & A167;
  assign \new_[72057]_  = A202 & ~A201;
  assign \new_[72058]_  = \new_[72057]_  & \new_[72054]_ ;
  assign \new_[72059]_  = \new_[72058]_  & \new_[72051]_ ;
  assign \new_[72063]_  = ~A298 & A266;
  assign \new_[72064]_  = A265 & \new_[72063]_ ;
  assign \new_[72067]_  = ~A300 & A299;
  assign \new_[72070]_  = A302 & ~A301;
  assign \new_[72071]_  = \new_[72070]_  & \new_[72067]_ ;
  assign \new_[72072]_  = \new_[72071]_  & \new_[72064]_ ;
  assign \new_[72076]_  = ~A168 & ~A169;
  assign \new_[72077]_  = ~A170 & \new_[72076]_ ;
  assign \new_[72080]_  = ~A166 & A167;
  assign \new_[72083]_  = A202 & ~A201;
  assign \new_[72084]_  = \new_[72083]_  & \new_[72080]_ ;
  assign \new_[72085]_  = \new_[72084]_  & \new_[72077]_ ;
  assign \new_[72089]_  = A267 & A266;
  assign \new_[72090]_  = ~A265 & \new_[72089]_ ;
  assign \new_[72093]_  = A300 & A268;
  assign \new_[72096]_  = A302 & ~A301;
  assign \new_[72097]_  = \new_[72096]_  & \new_[72093]_ ;
  assign \new_[72098]_  = \new_[72097]_  & \new_[72090]_ ;
  assign \new_[72102]_  = ~A168 & ~A169;
  assign \new_[72103]_  = ~A170 & \new_[72102]_ ;
  assign \new_[72106]_  = ~A166 & A167;
  assign \new_[72109]_  = A202 & ~A201;
  assign \new_[72110]_  = \new_[72109]_  & \new_[72106]_ ;
  assign \new_[72111]_  = \new_[72110]_  & \new_[72103]_ ;
  assign \new_[72115]_  = A267 & A266;
  assign \new_[72116]_  = ~A265 & \new_[72115]_ ;
  assign \new_[72119]_  = A300 & ~A269;
  assign \new_[72122]_  = A302 & ~A301;
  assign \new_[72123]_  = \new_[72122]_  & \new_[72119]_ ;
  assign \new_[72124]_  = \new_[72123]_  & \new_[72116]_ ;
  assign \new_[72128]_  = ~A168 & ~A169;
  assign \new_[72129]_  = ~A170 & \new_[72128]_ ;
  assign \new_[72132]_  = ~A166 & A167;
  assign \new_[72135]_  = A202 & ~A201;
  assign \new_[72136]_  = \new_[72135]_  & \new_[72132]_ ;
  assign \new_[72137]_  = \new_[72136]_  & \new_[72129]_ ;
  assign \new_[72141]_  = ~A267 & A266;
  assign \new_[72142]_  = ~A265 & \new_[72141]_ ;
  assign \new_[72145]_  = A269 & ~A268;
  assign \new_[72148]_  = A301 & ~A300;
  assign \new_[72149]_  = \new_[72148]_  & \new_[72145]_ ;
  assign \new_[72150]_  = \new_[72149]_  & \new_[72142]_ ;
  assign \new_[72154]_  = ~A168 & ~A169;
  assign \new_[72155]_  = ~A170 & \new_[72154]_ ;
  assign \new_[72158]_  = ~A166 & A167;
  assign \new_[72161]_  = A202 & ~A201;
  assign \new_[72162]_  = \new_[72161]_  & \new_[72158]_ ;
  assign \new_[72163]_  = \new_[72162]_  & \new_[72155]_ ;
  assign \new_[72167]_  = ~A267 & A266;
  assign \new_[72168]_  = ~A265 & \new_[72167]_ ;
  assign \new_[72171]_  = A269 & ~A268;
  assign \new_[72174]_  = ~A302 & ~A300;
  assign \new_[72175]_  = \new_[72174]_  & \new_[72171]_ ;
  assign \new_[72176]_  = \new_[72175]_  & \new_[72168]_ ;
  assign \new_[72180]_  = ~A168 & ~A169;
  assign \new_[72181]_  = ~A170 & \new_[72180]_ ;
  assign \new_[72184]_  = ~A166 & A167;
  assign \new_[72187]_  = A202 & ~A201;
  assign \new_[72188]_  = \new_[72187]_  & \new_[72184]_ ;
  assign \new_[72189]_  = \new_[72188]_  & \new_[72181]_ ;
  assign \new_[72193]_  = ~A267 & A266;
  assign \new_[72194]_  = ~A265 & \new_[72193]_ ;
  assign \new_[72197]_  = A269 & ~A268;
  assign \new_[72200]_  = A299 & A298;
  assign \new_[72201]_  = \new_[72200]_  & \new_[72197]_ ;
  assign \new_[72202]_  = \new_[72201]_  & \new_[72194]_ ;
  assign \new_[72206]_  = ~A168 & ~A169;
  assign \new_[72207]_  = ~A170 & \new_[72206]_ ;
  assign \new_[72210]_  = ~A166 & A167;
  assign \new_[72213]_  = A202 & ~A201;
  assign \new_[72214]_  = \new_[72213]_  & \new_[72210]_ ;
  assign \new_[72215]_  = \new_[72214]_  & \new_[72207]_ ;
  assign \new_[72219]_  = ~A267 & A266;
  assign \new_[72220]_  = ~A265 & \new_[72219]_ ;
  assign \new_[72223]_  = A269 & ~A268;
  assign \new_[72226]_  = ~A299 & ~A298;
  assign \new_[72227]_  = \new_[72226]_  & \new_[72223]_ ;
  assign \new_[72228]_  = \new_[72227]_  & \new_[72220]_ ;
  assign \new_[72232]_  = ~A168 & ~A169;
  assign \new_[72233]_  = ~A170 & \new_[72232]_ ;
  assign \new_[72236]_  = ~A166 & A167;
  assign \new_[72239]_  = A202 & ~A201;
  assign \new_[72240]_  = \new_[72239]_  & \new_[72236]_ ;
  assign \new_[72241]_  = \new_[72240]_  & \new_[72233]_ ;
  assign \new_[72245]_  = A267 & ~A266;
  assign \new_[72246]_  = A265 & \new_[72245]_ ;
  assign \new_[72249]_  = A300 & A268;
  assign \new_[72252]_  = A302 & ~A301;
  assign \new_[72253]_  = \new_[72252]_  & \new_[72249]_ ;
  assign \new_[72254]_  = \new_[72253]_  & \new_[72246]_ ;
  assign \new_[72258]_  = ~A168 & ~A169;
  assign \new_[72259]_  = ~A170 & \new_[72258]_ ;
  assign \new_[72262]_  = ~A166 & A167;
  assign \new_[72265]_  = A202 & ~A201;
  assign \new_[72266]_  = \new_[72265]_  & \new_[72262]_ ;
  assign \new_[72267]_  = \new_[72266]_  & \new_[72259]_ ;
  assign \new_[72271]_  = A267 & ~A266;
  assign \new_[72272]_  = A265 & \new_[72271]_ ;
  assign \new_[72275]_  = A300 & ~A269;
  assign \new_[72278]_  = A302 & ~A301;
  assign \new_[72279]_  = \new_[72278]_  & \new_[72275]_ ;
  assign \new_[72280]_  = \new_[72279]_  & \new_[72272]_ ;
  assign \new_[72284]_  = ~A168 & ~A169;
  assign \new_[72285]_  = ~A170 & \new_[72284]_ ;
  assign \new_[72288]_  = ~A166 & A167;
  assign \new_[72291]_  = A202 & ~A201;
  assign \new_[72292]_  = \new_[72291]_  & \new_[72288]_ ;
  assign \new_[72293]_  = \new_[72292]_  & \new_[72285]_ ;
  assign \new_[72297]_  = ~A267 & ~A266;
  assign \new_[72298]_  = A265 & \new_[72297]_ ;
  assign \new_[72301]_  = A269 & ~A268;
  assign \new_[72304]_  = A301 & ~A300;
  assign \new_[72305]_  = \new_[72304]_  & \new_[72301]_ ;
  assign \new_[72306]_  = \new_[72305]_  & \new_[72298]_ ;
  assign \new_[72310]_  = ~A168 & ~A169;
  assign \new_[72311]_  = ~A170 & \new_[72310]_ ;
  assign \new_[72314]_  = ~A166 & A167;
  assign \new_[72317]_  = A202 & ~A201;
  assign \new_[72318]_  = \new_[72317]_  & \new_[72314]_ ;
  assign \new_[72319]_  = \new_[72318]_  & \new_[72311]_ ;
  assign \new_[72323]_  = ~A267 & ~A266;
  assign \new_[72324]_  = A265 & \new_[72323]_ ;
  assign \new_[72327]_  = A269 & ~A268;
  assign \new_[72330]_  = ~A302 & ~A300;
  assign \new_[72331]_  = \new_[72330]_  & \new_[72327]_ ;
  assign \new_[72332]_  = \new_[72331]_  & \new_[72324]_ ;
  assign \new_[72336]_  = ~A168 & ~A169;
  assign \new_[72337]_  = ~A170 & \new_[72336]_ ;
  assign \new_[72340]_  = ~A166 & A167;
  assign \new_[72343]_  = A202 & ~A201;
  assign \new_[72344]_  = \new_[72343]_  & \new_[72340]_ ;
  assign \new_[72345]_  = \new_[72344]_  & \new_[72337]_ ;
  assign \new_[72349]_  = ~A267 & ~A266;
  assign \new_[72350]_  = A265 & \new_[72349]_ ;
  assign \new_[72353]_  = A269 & ~A268;
  assign \new_[72356]_  = A299 & A298;
  assign \new_[72357]_  = \new_[72356]_  & \new_[72353]_ ;
  assign \new_[72358]_  = \new_[72357]_  & \new_[72350]_ ;
  assign \new_[72362]_  = ~A168 & ~A169;
  assign \new_[72363]_  = ~A170 & \new_[72362]_ ;
  assign \new_[72366]_  = ~A166 & A167;
  assign \new_[72369]_  = A202 & ~A201;
  assign \new_[72370]_  = \new_[72369]_  & \new_[72366]_ ;
  assign \new_[72371]_  = \new_[72370]_  & \new_[72363]_ ;
  assign \new_[72375]_  = ~A267 & ~A266;
  assign \new_[72376]_  = A265 & \new_[72375]_ ;
  assign \new_[72379]_  = A269 & ~A268;
  assign \new_[72382]_  = ~A299 & ~A298;
  assign \new_[72383]_  = \new_[72382]_  & \new_[72379]_ ;
  assign \new_[72384]_  = \new_[72383]_  & \new_[72376]_ ;
  assign \new_[72388]_  = ~A168 & ~A169;
  assign \new_[72389]_  = ~A170 & \new_[72388]_ ;
  assign \new_[72392]_  = ~A166 & A167;
  assign \new_[72395]_  = A202 & ~A201;
  assign \new_[72396]_  = \new_[72395]_  & \new_[72392]_ ;
  assign \new_[72397]_  = \new_[72396]_  & \new_[72389]_ ;
  assign \new_[72401]_  = A298 & ~A266;
  assign \new_[72402]_  = ~A265 & \new_[72401]_ ;
  assign \new_[72405]_  = ~A300 & ~A299;
  assign \new_[72408]_  = A302 & ~A301;
  assign \new_[72409]_  = \new_[72408]_  & \new_[72405]_ ;
  assign \new_[72410]_  = \new_[72409]_  & \new_[72402]_ ;
  assign \new_[72414]_  = ~A168 & ~A169;
  assign \new_[72415]_  = ~A170 & \new_[72414]_ ;
  assign \new_[72418]_  = ~A166 & A167;
  assign \new_[72421]_  = A202 & ~A201;
  assign \new_[72422]_  = \new_[72421]_  & \new_[72418]_ ;
  assign \new_[72423]_  = \new_[72422]_  & \new_[72415]_ ;
  assign \new_[72427]_  = ~A298 & ~A266;
  assign \new_[72428]_  = ~A265 & \new_[72427]_ ;
  assign \new_[72431]_  = ~A300 & A299;
  assign \new_[72434]_  = A302 & ~A301;
  assign \new_[72435]_  = \new_[72434]_  & \new_[72431]_ ;
  assign \new_[72436]_  = \new_[72435]_  & \new_[72428]_ ;
  assign \new_[72440]_  = ~A168 & ~A169;
  assign \new_[72441]_  = ~A170 & \new_[72440]_ ;
  assign \new_[72444]_  = ~A166 & A167;
  assign \new_[72447]_  = ~A203 & ~A201;
  assign \new_[72448]_  = \new_[72447]_  & \new_[72444]_ ;
  assign \new_[72449]_  = \new_[72448]_  & \new_[72441]_ ;
  assign \new_[72453]_  = A269 & ~A268;
  assign \new_[72454]_  = A267 & \new_[72453]_ ;
  assign \new_[72457]_  = ~A299 & A298;
  assign \new_[72460]_  = A301 & A300;
  assign \new_[72461]_  = \new_[72460]_  & \new_[72457]_ ;
  assign \new_[72462]_  = \new_[72461]_  & \new_[72454]_ ;
  assign \new_[72466]_  = ~A168 & ~A169;
  assign \new_[72467]_  = ~A170 & \new_[72466]_ ;
  assign \new_[72470]_  = ~A166 & A167;
  assign \new_[72473]_  = ~A203 & ~A201;
  assign \new_[72474]_  = \new_[72473]_  & \new_[72470]_ ;
  assign \new_[72475]_  = \new_[72474]_  & \new_[72467]_ ;
  assign \new_[72479]_  = A269 & ~A268;
  assign \new_[72480]_  = A267 & \new_[72479]_ ;
  assign \new_[72483]_  = ~A299 & A298;
  assign \new_[72486]_  = ~A302 & A300;
  assign \new_[72487]_  = \new_[72486]_  & \new_[72483]_ ;
  assign \new_[72488]_  = \new_[72487]_  & \new_[72480]_ ;
  assign \new_[72492]_  = ~A168 & ~A169;
  assign \new_[72493]_  = ~A170 & \new_[72492]_ ;
  assign \new_[72496]_  = ~A166 & A167;
  assign \new_[72499]_  = ~A203 & ~A201;
  assign \new_[72500]_  = \new_[72499]_  & \new_[72496]_ ;
  assign \new_[72501]_  = \new_[72500]_  & \new_[72493]_ ;
  assign \new_[72505]_  = A269 & ~A268;
  assign \new_[72506]_  = A267 & \new_[72505]_ ;
  assign \new_[72509]_  = A299 & ~A298;
  assign \new_[72512]_  = A301 & A300;
  assign \new_[72513]_  = \new_[72512]_  & \new_[72509]_ ;
  assign \new_[72514]_  = \new_[72513]_  & \new_[72506]_ ;
  assign \new_[72518]_  = ~A168 & ~A169;
  assign \new_[72519]_  = ~A170 & \new_[72518]_ ;
  assign \new_[72522]_  = ~A166 & A167;
  assign \new_[72525]_  = ~A203 & ~A201;
  assign \new_[72526]_  = \new_[72525]_  & \new_[72522]_ ;
  assign \new_[72527]_  = \new_[72526]_  & \new_[72519]_ ;
  assign \new_[72531]_  = A269 & ~A268;
  assign \new_[72532]_  = A267 & \new_[72531]_ ;
  assign \new_[72535]_  = A299 & ~A298;
  assign \new_[72538]_  = ~A302 & A300;
  assign \new_[72539]_  = \new_[72538]_  & \new_[72535]_ ;
  assign \new_[72540]_  = \new_[72539]_  & \new_[72532]_ ;
  assign \new_[72544]_  = ~A168 & ~A169;
  assign \new_[72545]_  = ~A170 & \new_[72544]_ ;
  assign \new_[72548]_  = ~A166 & A167;
  assign \new_[72551]_  = ~A203 & ~A201;
  assign \new_[72552]_  = \new_[72551]_  & \new_[72548]_ ;
  assign \new_[72553]_  = \new_[72552]_  & \new_[72545]_ ;
  assign \new_[72557]_  = A298 & A268;
  assign \new_[72558]_  = ~A267 & \new_[72557]_ ;
  assign \new_[72561]_  = ~A300 & ~A299;
  assign \new_[72564]_  = A302 & ~A301;
  assign \new_[72565]_  = \new_[72564]_  & \new_[72561]_ ;
  assign \new_[72566]_  = \new_[72565]_  & \new_[72558]_ ;
  assign \new_[72570]_  = ~A168 & ~A169;
  assign \new_[72571]_  = ~A170 & \new_[72570]_ ;
  assign \new_[72574]_  = ~A166 & A167;
  assign \new_[72577]_  = ~A203 & ~A201;
  assign \new_[72578]_  = \new_[72577]_  & \new_[72574]_ ;
  assign \new_[72579]_  = \new_[72578]_  & \new_[72571]_ ;
  assign \new_[72583]_  = ~A298 & A268;
  assign \new_[72584]_  = ~A267 & \new_[72583]_ ;
  assign \new_[72587]_  = ~A300 & A299;
  assign \new_[72590]_  = A302 & ~A301;
  assign \new_[72591]_  = \new_[72590]_  & \new_[72587]_ ;
  assign \new_[72592]_  = \new_[72591]_  & \new_[72584]_ ;
  assign \new_[72596]_  = ~A168 & ~A169;
  assign \new_[72597]_  = ~A170 & \new_[72596]_ ;
  assign \new_[72600]_  = ~A166 & A167;
  assign \new_[72603]_  = ~A203 & ~A201;
  assign \new_[72604]_  = \new_[72603]_  & \new_[72600]_ ;
  assign \new_[72605]_  = \new_[72604]_  & \new_[72597]_ ;
  assign \new_[72609]_  = A298 & ~A269;
  assign \new_[72610]_  = ~A267 & \new_[72609]_ ;
  assign \new_[72613]_  = ~A300 & ~A299;
  assign \new_[72616]_  = A302 & ~A301;
  assign \new_[72617]_  = \new_[72616]_  & \new_[72613]_ ;
  assign \new_[72618]_  = \new_[72617]_  & \new_[72610]_ ;
  assign \new_[72622]_  = ~A168 & ~A169;
  assign \new_[72623]_  = ~A170 & \new_[72622]_ ;
  assign \new_[72626]_  = ~A166 & A167;
  assign \new_[72629]_  = ~A203 & ~A201;
  assign \new_[72630]_  = \new_[72629]_  & \new_[72626]_ ;
  assign \new_[72631]_  = \new_[72630]_  & \new_[72623]_ ;
  assign \new_[72635]_  = ~A298 & ~A269;
  assign \new_[72636]_  = ~A267 & \new_[72635]_ ;
  assign \new_[72639]_  = ~A300 & A299;
  assign \new_[72642]_  = A302 & ~A301;
  assign \new_[72643]_  = \new_[72642]_  & \new_[72639]_ ;
  assign \new_[72644]_  = \new_[72643]_  & \new_[72636]_ ;
  assign \new_[72648]_  = ~A168 & ~A169;
  assign \new_[72649]_  = ~A170 & \new_[72648]_ ;
  assign \new_[72652]_  = ~A166 & A167;
  assign \new_[72655]_  = ~A203 & ~A201;
  assign \new_[72656]_  = \new_[72655]_  & \new_[72652]_ ;
  assign \new_[72657]_  = \new_[72656]_  & \new_[72649]_ ;
  assign \new_[72661]_  = A298 & A266;
  assign \new_[72662]_  = A265 & \new_[72661]_ ;
  assign \new_[72665]_  = ~A300 & ~A299;
  assign \new_[72668]_  = A302 & ~A301;
  assign \new_[72669]_  = \new_[72668]_  & \new_[72665]_ ;
  assign \new_[72670]_  = \new_[72669]_  & \new_[72662]_ ;
  assign \new_[72674]_  = ~A168 & ~A169;
  assign \new_[72675]_  = ~A170 & \new_[72674]_ ;
  assign \new_[72678]_  = ~A166 & A167;
  assign \new_[72681]_  = ~A203 & ~A201;
  assign \new_[72682]_  = \new_[72681]_  & \new_[72678]_ ;
  assign \new_[72683]_  = \new_[72682]_  & \new_[72675]_ ;
  assign \new_[72687]_  = ~A298 & A266;
  assign \new_[72688]_  = A265 & \new_[72687]_ ;
  assign \new_[72691]_  = ~A300 & A299;
  assign \new_[72694]_  = A302 & ~A301;
  assign \new_[72695]_  = \new_[72694]_  & \new_[72691]_ ;
  assign \new_[72696]_  = \new_[72695]_  & \new_[72688]_ ;
  assign \new_[72700]_  = ~A168 & ~A169;
  assign \new_[72701]_  = ~A170 & \new_[72700]_ ;
  assign \new_[72704]_  = ~A166 & A167;
  assign \new_[72707]_  = ~A203 & ~A201;
  assign \new_[72708]_  = \new_[72707]_  & \new_[72704]_ ;
  assign \new_[72709]_  = \new_[72708]_  & \new_[72701]_ ;
  assign \new_[72713]_  = A267 & A266;
  assign \new_[72714]_  = ~A265 & \new_[72713]_ ;
  assign \new_[72717]_  = A300 & A268;
  assign \new_[72720]_  = A302 & ~A301;
  assign \new_[72721]_  = \new_[72720]_  & \new_[72717]_ ;
  assign \new_[72722]_  = \new_[72721]_  & \new_[72714]_ ;
  assign \new_[72726]_  = ~A168 & ~A169;
  assign \new_[72727]_  = ~A170 & \new_[72726]_ ;
  assign \new_[72730]_  = ~A166 & A167;
  assign \new_[72733]_  = ~A203 & ~A201;
  assign \new_[72734]_  = \new_[72733]_  & \new_[72730]_ ;
  assign \new_[72735]_  = \new_[72734]_  & \new_[72727]_ ;
  assign \new_[72739]_  = A267 & A266;
  assign \new_[72740]_  = ~A265 & \new_[72739]_ ;
  assign \new_[72743]_  = A300 & ~A269;
  assign \new_[72746]_  = A302 & ~A301;
  assign \new_[72747]_  = \new_[72746]_  & \new_[72743]_ ;
  assign \new_[72748]_  = \new_[72747]_  & \new_[72740]_ ;
  assign \new_[72752]_  = ~A168 & ~A169;
  assign \new_[72753]_  = ~A170 & \new_[72752]_ ;
  assign \new_[72756]_  = ~A166 & A167;
  assign \new_[72759]_  = ~A203 & ~A201;
  assign \new_[72760]_  = \new_[72759]_  & \new_[72756]_ ;
  assign \new_[72761]_  = \new_[72760]_  & \new_[72753]_ ;
  assign \new_[72765]_  = ~A267 & A266;
  assign \new_[72766]_  = ~A265 & \new_[72765]_ ;
  assign \new_[72769]_  = A269 & ~A268;
  assign \new_[72772]_  = A301 & ~A300;
  assign \new_[72773]_  = \new_[72772]_  & \new_[72769]_ ;
  assign \new_[72774]_  = \new_[72773]_  & \new_[72766]_ ;
  assign \new_[72778]_  = ~A168 & ~A169;
  assign \new_[72779]_  = ~A170 & \new_[72778]_ ;
  assign \new_[72782]_  = ~A166 & A167;
  assign \new_[72785]_  = ~A203 & ~A201;
  assign \new_[72786]_  = \new_[72785]_  & \new_[72782]_ ;
  assign \new_[72787]_  = \new_[72786]_  & \new_[72779]_ ;
  assign \new_[72791]_  = ~A267 & A266;
  assign \new_[72792]_  = ~A265 & \new_[72791]_ ;
  assign \new_[72795]_  = A269 & ~A268;
  assign \new_[72798]_  = ~A302 & ~A300;
  assign \new_[72799]_  = \new_[72798]_  & \new_[72795]_ ;
  assign \new_[72800]_  = \new_[72799]_  & \new_[72792]_ ;
  assign \new_[72804]_  = ~A168 & ~A169;
  assign \new_[72805]_  = ~A170 & \new_[72804]_ ;
  assign \new_[72808]_  = ~A166 & A167;
  assign \new_[72811]_  = ~A203 & ~A201;
  assign \new_[72812]_  = \new_[72811]_  & \new_[72808]_ ;
  assign \new_[72813]_  = \new_[72812]_  & \new_[72805]_ ;
  assign \new_[72817]_  = ~A267 & A266;
  assign \new_[72818]_  = ~A265 & \new_[72817]_ ;
  assign \new_[72821]_  = A269 & ~A268;
  assign \new_[72824]_  = A299 & A298;
  assign \new_[72825]_  = \new_[72824]_  & \new_[72821]_ ;
  assign \new_[72826]_  = \new_[72825]_  & \new_[72818]_ ;
  assign \new_[72830]_  = ~A168 & ~A169;
  assign \new_[72831]_  = ~A170 & \new_[72830]_ ;
  assign \new_[72834]_  = ~A166 & A167;
  assign \new_[72837]_  = ~A203 & ~A201;
  assign \new_[72838]_  = \new_[72837]_  & \new_[72834]_ ;
  assign \new_[72839]_  = \new_[72838]_  & \new_[72831]_ ;
  assign \new_[72843]_  = ~A267 & A266;
  assign \new_[72844]_  = ~A265 & \new_[72843]_ ;
  assign \new_[72847]_  = A269 & ~A268;
  assign \new_[72850]_  = ~A299 & ~A298;
  assign \new_[72851]_  = \new_[72850]_  & \new_[72847]_ ;
  assign \new_[72852]_  = \new_[72851]_  & \new_[72844]_ ;
  assign \new_[72856]_  = ~A168 & ~A169;
  assign \new_[72857]_  = ~A170 & \new_[72856]_ ;
  assign \new_[72860]_  = ~A166 & A167;
  assign \new_[72863]_  = ~A203 & ~A201;
  assign \new_[72864]_  = \new_[72863]_  & \new_[72860]_ ;
  assign \new_[72865]_  = \new_[72864]_  & \new_[72857]_ ;
  assign \new_[72869]_  = A267 & ~A266;
  assign \new_[72870]_  = A265 & \new_[72869]_ ;
  assign \new_[72873]_  = A300 & A268;
  assign \new_[72876]_  = A302 & ~A301;
  assign \new_[72877]_  = \new_[72876]_  & \new_[72873]_ ;
  assign \new_[72878]_  = \new_[72877]_  & \new_[72870]_ ;
  assign \new_[72882]_  = ~A168 & ~A169;
  assign \new_[72883]_  = ~A170 & \new_[72882]_ ;
  assign \new_[72886]_  = ~A166 & A167;
  assign \new_[72889]_  = ~A203 & ~A201;
  assign \new_[72890]_  = \new_[72889]_  & \new_[72886]_ ;
  assign \new_[72891]_  = \new_[72890]_  & \new_[72883]_ ;
  assign \new_[72895]_  = A267 & ~A266;
  assign \new_[72896]_  = A265 & \new_[72895]_ ;
  assign \new_[72899]_  = A300 & ~A269;
  assign \new_[72902]_  = A302 & ~A301;
  assign \new_[72903]_  = \new_[72902]_  & \new_[72899]_ ;
  assign \new_[72904]_  = \new_[72903]_  & \new_[72896]_ ;
  assign \new_[72908]_  = ~A168 & ~A169;
  assign \new_[72909]_  = ~A170 & \new_[72908]_ ;
  assign \new_[72912]_  = ~A166 & A167;
  assign \new_[72915]_  = ~A203 & ~A201;
  assign \new_[72916]_  = \new_[72915]_  & \new_[72912]_ ;
  assign \new_[72917]_  = \new_[72916]_  & \new_[72909]_ ;
  assign \new_[72921]_  = ~A267 & ~A266;
  assign \new_[72922]_  = A265 & \new_[72921]_ ;
  assign \new_[72925]_  = A269 & ~A268;
  assign \new_[72928]_  = A301 & ~A300;
  assign \new_[72929]_  = \new_[72928]_  & \new_[72925]_ ;
  assign \new_[72930]_  = \new_[72929]_  & \new_[72922]_ ;
  assign \new_[72934]_  = ~A168 & ~A169;
  assign \new_[72935]_  = ~A170 & \new_[72934]_ ;
  assign \new_[72938]_  = ~A166 & A167;
  assign \new_[72941]_  = ~A203 & ~A201;
  assign \new_[72942]_  = \new_[72941]_  & \new_[72938]_ ;
  assign \new_[72943]_  = \new_[72942]_  & \new_[72935]_ ;
  assign \new_[72947]_  = ~A267 & ~A266;
  assign \new_[72948]_  = A265 & \new_[72947]_ ;
  assign \new_[72951]_  = A269 & ~A268;
  assign \new_[72954]_  = ~A302 & ~A300;
  assign \new_[72955]_  = \new_[72954]_  & \new_[72951]_ ;
  assign \new_[72956]_  = \new_[72955]_  & \new_[72948]_ ;
  assign \new_[72960]_  = ~A168 & ~A169;
  assign \new_[72961]_  = ~A170 & \new_[72960]_ ;
  assign \new_[72964]_  = ~A166 & A167;
  assign \new_[72967]_  = ~A203 & ~A201;
  assign \new_[72968]_  = \new_[72967]_  & \new_[72964]_ ;
  assign \new_[72969]_  = \new_[72968]_  & \new_[72961]_ ;
  assign \new_[72973]_  = ~A267 & ~A266;
  assign \new_[72974]_  = A265 & \new_[72973]_ ;
  assign \new_[72977]_  = A269 & ~A268;
  assign \new_[72980]_  = A299 & A298;
  assign \new_[72981]_  = \new_[72980]_  & \new_[72977]_ ;
  assign \new_[72982]_  = \new_[72981]_  & \new_[72974]_ ;
  assign \new_[72986]_  = ~A168 & ~A169;
  assign \new_[72987]_  = ~A170 & \new_[72986]_ ;
  assign \new_[72990]_  = ~A166 & A167;
  assign \new_[72993]_  = ~A203 & ~A201;
  assign \new_[72994]_  = \new_[72993]_  & \new_[72990]_ ;
  assign \new_[72995]_  = \new_[72994]_  & \new_[72987]_ ;
  assign \new_[72999]_  = ~A267 & ~A266;
  assign \new_[73000]_  = A265 & \new_[72999]_ ;
  assign \new_[73003]_  = A269 & ~A268;
  assign \new_[73006]_  = ~A299 & ~A298;
  assign \new_[73007]_  = \new_[73006]_  & \new_[73003]_ ;
  assign \new_[73008]_  = \new_[73007]_  & \new_[73000]_ ;
  assign \new_[73012]_  = ~A168 & ~A169;
  assign \new_[73013]_  = ~A170 & \new_[73012]_ ;
  assign \new_[73016]_  = ~A166 & A167;
  assign \new_[73019]_  = ~A203 & ~A201;
  assign \new_[73020]_  = \new_[73019]_  & \new_[73016]_ ;
  assign \new_[73021]_  = \new_[73020]_  & \new_[73013]_ ;
  assign \new_[73025]_  = A298 & ~A266;
  assign \new_[73026]_  = ~A265 & \new_[73025]_ ;
  assign \new_[73029]_  = ~A300 & ~A299;
  assign \new_[73032]_  = A302 & ~A301;
  assign \new_[73033]_  = \new_[73032]_  & \new_[73029]_ ;
  assign \new_[73034]_  = \new_[73033]_  & \new_[73026]_ ;
  assign \new_[73038]_  = ~A168 & ~A169;
  assign \new_[73039]_  = ~A170 & \new_[73038]_ ;
  assign \new_[73042]_  = ~A166 & A167;
  assign \new_[73045]_  = ~A203 & ~A201;
  assign \new_[73046]_  = \new_[73045]_  & \new_[73042]_ ;
  assign \new_[73047]_  = \new_[73046]_  & \new_[73039]_ ;
  assign \new_[73051]_  = ~A298 & ~A266;
  assign \new_[73052]_  = ~A265 & \new_[73051]_ ;
  assign \new_[73055]_  = ~A300 & A299;
  assign \new_[73058]_  = A302 & ~A301;
  assign \new_[73059]_  = \new_[73058]_  & \new_[73055]_ ;
  assign \new_[73060]_  = \new_[73059]_  & \new_[73052]_ ;
  assign \new_[73064]_  = ~A168 & ~A169;
  assign \new_[73065]_  = ~A170 & \new_[73064]_ ;
  assign \new_[73068]_  = ~A166 & A167;
  assign \new_[73071]_  = A200 & A199;
  assign \new_[73072]_  = \new_[73071]_  & \new_[73068]_ ;
  assign \new_[73073]_  = \new_[73072]_  & \new_[73065]_ ;
  assign \new_[73077]_  = A269 & ~A268;
  assign \new_[73078]_  = A267 & \new_[73077]_ ;
  assign \new_[73081]_  = ~A299 & A298;
  assign \new_[73084]_  = A301 & A300;
  assign \new_[73085]_  = \new_[73084]_  & \new_[73081]_ ;
  assign \new_[73086]_  = \new_[73085]_  & \new_[73078]_ ;
  assign \new_[73090]_  = ~A168 & ~A169;
  assign \new_[73091]_  = ~A170 & \new_[73090]_ ;
  assign \new_[73094]_  = ~A166 & A167;
  assign \new_[73097]_  = A200 & A199;
  assign \new_[73098]_  = \new_[73097]_  & \new_[73094]_ ;
  assign \new_[73099]_  = \new_[73098]_  & \new_[73091]_ ;
  assign \new_[73103]_  = A269 & ~A268;
  assign \new_[73104]_  = A267 & \new_[73103]_ ;
  assign \new_[73107]_  = ~A299 & A298;
  assign \new_[73110]_  = ~A302 & A300;
  assign \new_[73111]_  = \new_[73110]_  & \new_[73107]_ ;
  assign \new_[73112]_  = \new_[73111]_  & \new_[73104]_ ;
  assign \new_[73116]_  = ~A168 & ~A169;
  assign \new_[73117]_  = ~A170 & \new_[73116]_ ;
  assign \new_[73120]_  = ~A166 & A167;
  assign \new_[73123]_  = A200 & A199;
  assign \new_[73124]_  = \new_[73123]_  & \new_[73120]_ ;
  assign \new_[73125]_  = \new_[73124]_  & \new_[73117]_ ;
  assign \new_[73129]_  = A269 & ~A268;
  assign \new_[73130]_  = A267 & \new_[73129]_ ;
  assign \new_[73133]_  = A299 & ~A298;
  assign \new_[73136]_  = A301 & A300;
  assign \new_[73137]_  = \new_[73136]_  & \new_[73133]_ ;
  assign \new_[73138]_  = \new_[73137]_  & \new_[73130]_ ;
  assign \new_[73142]_  = ~A168 & ~A169;
  assign \new_[73143]_  = ~A170 & \new_[73142]_ ;
  assign \new_[73146]_  = ~A166 & A167;
  assign \new_[73149]_  = A200 & A199;
  assign \new_[73150]_  = \new_[73149]_  & \new_[73146]_ ;
  assign \new_[73151]_  = \new_[73150]_  & \new_[73143]_ ;
  assign \new_[73155]_  = A269 & ~A268;
  assign \new_[73156]_  = A267 & \new_[73155]_ ;
  assign \new_[73159]_  = A299 & ~A298;
  assign \new_[73162]_  = ~A302 & A300;
  assign \new_[73163]_  = \new_[73162]_  & \new_[73159]_ ;
  assign \new_[73164]_  = \new_[73163]_  & \new_[73156]_ ;
  assign \new_[73168]_  = ~A168 & ~A169;
  assign \new_[73169]_  = ~A170 & \new_[73168]_ ;
  assign \new_[73172]_  = ~A166 & A167;
  assign \new_[73175]_  = A200 & A199;
  assign \new_[73176]_  = \new_[73175]_  & \new_[73172]_ ;
  assign \new_[73177]_  = \new_[73176]_  & \new_[73169]_ ;
  assign \new_[73181]_  = A298 & A268;
  assign \new_[73182]_  = ~A267 & \new_[73181]_ ;
  assign \new_[73185]_  = ~A300 & ~A299;
  assign \new_[73188]_  = A302 & ~A301;
  assign \new_[73189]_  = \new_[73188]_  & \new_[73185]_ ;
  assign \new_[73190]_  = \new_[73189]_  & \new_[73182]_ ;
  assign \new_[73194]_  = ~A168 & ~A169;
  assign \new_[73195]_  = ~A170 & \new_[73194]_ ;
  assign \new_[73198]_  = ~A166 & A167;
  assign \new_[73201]_  = A200 & A199;
  assign \new_[73202]_  = \new_[73201]_  & \new_[73198]_ ;
  assign \new_[73203]_  = \new_[73202]_  & \new_[73195]_ ;
  assign \new_[73207]_  = ~A298 & A268;
  assign \new_[73208]_  = ~A267 & \new_[73207]_ ;
  assign \new_[73211]_  = ~A300 & A299;
  assign \new_[73214]_  = A302 & ~A301;
  assign \new_[73215]_  = \new_[73214]_  & \new_[73211]_ ;
  assign \new_[73216]_  = \new_[73215]_  & \new_[73208]_ ;
  assign \new_[73220]_  = ~A168 & ~A169;
  assign \new_[73221]_  = ~A170 & \new_[73220]_ ;
  assign \new_[73224]_  = ~A166 & A167;
  assign \new_[73227]_  = A200 & A199;
  assign \new_[73228]_  = \new_[73227]_  & \new_[73224]_ ;
  assign \new_[73229]_  = \new_[73228]_  & \new_[73221]_ ;
  assign \new_[73233]_  = A298 & ~A269;
  assign \new_[73234]_  = ~A267 & \new_[73233]_ ;
  assign \new_[73237]_  = ~A300 & ~A299;
  assign \new_[73240]_  = A302 & ~A301;
  assign \new_[73241]_  = \new_[73240]_  & \new_[73237]_ ;
  assign \new_[73242]_  = \new_[73241]_  & \new_[73234]_ ;
  assign \new_[73246]_  = ~A168 & ~A169;
  assign \new_[73247]_  = ~A170 & \new_[73246]_ ;
  assign \new_[73250]_  = ~A166 & A167;
  assign \new_[73253]_  = A200 & A199;
  assign \new_[73254]_  = \new_[73253]_  & \new_[73250]_ ;
  assign \new_[73255]_  = \new_[73254]_  & \new_[73247]_ ;
  assign \new_[73259]_  = ~A298 & ~A269;
  assign \new_[73260]_  = ~A267 & \new_[73259]_ ;
  assign \new_[73263]_  = ~A300 & A299;
  assign \new_[73266]_  = A302 & ~A301;
  assign \new_[73267]_  = \new_[73266]_  & \new_[73263]_ ;
  assign \new_[73268]_  = \new_[73267]_  & \new_[73260]_ ;
  assign \new_[73272]_  = ~A168 & ~A169;
  assign \new_[73273]_  = ~A170 & \new_[73272]_ ;
  assign \new_[73276]_  = ~A166 & A167;
  assign \new_[73279]_  = A200 & A199;
  assign \new_[73280]_  = \new_[73279]_  & \new_[73276]_ ;
  assign \new_[73281]_  = \new_[73280]_  & \new_[73273]_ ;
  assign \new_[73285]_  = A298 & A266;
  assign \new_[73286]_  = A265 & \new_[73285]_ ;
  assign \new_[73289]_  = ~A300 & ~A299;
  assign \new_[73292]_  = A302 & ~A301;
  assign \new_[73293]_  = \new_[73292]_  & \new_[73289]_ ;
  assign \new_[73294]_  = \new_[73293]_  & \new_[73286]_ ;
  assign \new_[73298]_  = ~A168 & ~A169;
  assign \new_[73299]_  = ~A170 & \new_[73298]_ ;
  assign \new_[73302]_  = ~A166 & A167;
  assign \new_[73305]_  = A200 & A199;
  assign \new_[73306]_  = \new_[73305]_  & \new_[73302]_ ;
  assign \new_[73307]_  = \new_[73306]_  & \new_[73299]_ ;
  assign \new_[73311]_  = ~A298 & A266;
  assign \new_[73312]_  = A265 & \new_[73311]_ ;
  assign \new_[73315]_  = ~A300 & A299;
  assign \new_[73318]_  = A302 & ~A301;
  assign \new_[73319]_  = \new_[73318]_  & \new_[73315]_ ;
  assign \new_[73320]_  = \new_[73319]_  & \new_[73312]_ ;
  assign \new_[73324]_  = ~A168 & ~A169;
  assign \new_[73325]_  = ~A170 & \new_[73324]_ ;
  assign \new_[73328]_  = ~A166 & A167;
  assign \new_[73331]_  = A200 & A199;
  assign \new_[73332]_  = \new_[73331]_  & \new_[73328]_ ;
  assign \new_[73333]_  = \new_[73332]_  & \new_[73325]_ ;
  assign \new_[73337]_  = A267 & A266;
  assign \new_[73338]_  = ~A265 & \new_[73337]_ ;
  assign \new_[73341]_  = A300 & A268;
  assign \new_[73344]_  = A302 & ~A301;
  assign \new_[73345]_  = \new_[73344]_  & \new_[73341]_ ;
  assign \new_[73346]_  = \new_[73345]_  & \new_[73338]_ ;
  assign \new_[73350]_  = ~A168 & ~A169;
  assign \new_[73351]_  = ~A170 & \new_[73350]_ ;
  assign \new_[73354]_  = ~A166 & A167;
  assign \new_[73357]_  = A200 & A199;
  assign \new_[73358]_  = \new_[73357]_  & \new_[73354]_ ;
  assign \new_[73359]_  = \new_[73358]_  & \new_[73351]_ ;
  assign \new_[73363]_  = A267 & A266;
  assign \new_[73364]_  = ~A265 & \new_[73363]_ ;
  assign \new_[73367]_  = A300 & ~A269;
  assign \new_[73370]_  = A302 & ~A301;
  assign \new_[73371]_  = \new_[73370]_  & \new_[73367]_ ;
  assign \new_[73372]_  = \new_[73371]_  & \new_[73364]_ ;
  assign \new_[73376]_  = ~A168 & ~A169;
  assign \new_[73377]_  = ~A170 & \new_[73376]_ ;
  assign \new_[73380]_  = ~A166 & A167;
  assign \new_[73383]_  = A200 & A199;
  assign \new_[73384]_  = \new_[73383]_  & \new_[73380]_ ;
  assign \new_[73385]_  = \new_[73384]_  & \new_[73377]_ ;
  assign \new_[73389]_  = ~A267 & A266;
  assign \new_[73390]_  = ~A265 & \new_[73389]_ ;
  assign \new_[73393]_  = A269 & ~A268;
  assign \new_[73396]_  = A301 & ~A300;
  assign \new_[73397]_  = \new_[73396]_  & \new_[73393]_ ;
  assign \new_[73398]_  = \new_[73397]_  & \new_[73390]_ ;
  assign \new_[73402]_  = ~A168 & ~A169;
  assign \new_[73403]_  = ~A170 & \new_[73402]_ ;
  assign \new_[73406]_  = ~A166 & A167;
  assign \new_[73409]_  = A200 & A199;
  assign \new_[73410]_  = \new_[73409]_  & \new_[73406]_ ;
  assign \new_[73411]_  = \new_[73410]_  & \new_[73403]_ ;
  assign \new_[73415]_  = ~A267 & A266;
  assign \new_[73416]_  = ~A265 & \new_[73415]_ ;
  assign \new_[73419]_  = A269 & ~A268;
  assign \new_[73422]_  = ~A302 & ~A300;
  assign \new_[73423]_  = \new_[73422]_  & \new_[73419]_ ;
  assign \new_[73424]_  = \new_[73423]_  & \new_[73416]_ ;
  assign \new_[73428]_  = ~A168 & ~A169;
  assign \new_[73429]_  = ~A170 & \new_[73428]_ ;
  assign \new_[73432]_  = ~A166 & A167;
  assign \new_[73435]_  = A200 & A199;
  assign \new_[73436]_  = \new_[73435]_  & \new_[73432]_ ;
  assign \new_[73437]_  = \new_[73436]_  & \new_[73429]_ ;
  assign \new_[73441]_  = ~A267 & A266;
  assign \new_[73442]_  = ~A265 & \new_[73441]_ ;
  assign \new_[73445]_  = A269 & ~A268;
  assign \new_[73448]_  = A299 & A298;
  assign \new_[73449]_  = \new_[73448]_  & \new_[73445]_ ;
  assign \new_[73450]_  = \new_[73449]_  & \new_[73442]_ ;
  assign \new_[73454]_  = ~A168 & ~A169;
  assign \new_[73455]_  = ~A170 & \new_[73454]_ ;
  assign \new_[73458]_  = ~A166 & A167;
  assign \new_[73461]_  = A200 & A199;
  assign \new_[73462]_  = \new_[73461]_  & \new_[73458]_ ;
  assign \new_[73463]_  = \new_[73462]_  & \new_[73455]_ ;
  assign \new_[73467]_  = ~A267 & A266;
  assign \new_[73468]_  = ~A265 & \new_[73467]_ ;
  assign \new_[73471]_  = A269 & ~A268;
  assign \new_[73474]_  = ~A299 & ~A298;
  assign \new_[73475]_  = \new_[73474]_  & \new_[73471]_ ;
  assign \new_[73476]_  = \new_[73475]_  & \new_[73468]_ ;
  assign \new_[73480]_  = ~A168 & ~A169;
  assign \new_[73481]_  = ~A170 & \new_[73480]_ ;
  assign \new_[73484]_  = ~A166 & A167;
  assign \new_[73487]_  = A200 & A199;
  assign \new_[73488]_  = \new_[73487]_  & \new_[73484]_ ;
  assign \new_[73489]_  = \new_[73488]_  & \new_[73481]_ ;
  assign \new_[73493]_  = A267 & ~A266;
  assign \new_[73494]_  = A265 & \new_[73493]_ ;
  assign \new_[73497]_  = A300 & A268;
  assign \new_[73500]_  = A302 & ~A301;
  assign \new_[73501]_  = \new_[73500]_  & \new_[73497]_ ;
  assign \new_[73502]_  = \new_[73501]_  & \new_[73494]_ ;
  assign \new_[73506]_  = ~A168 & ~A169;
  assign \new_[73507]_  = ~A170 & \new_[73506]_ ;
  assign \new_[73510]_  = ~A166 & A167;
  assign \new_[73513]_  = A200 & A199;
  assign \new_[73514]_  = \new_[73513]_  & \new_[73510]_ ;
  assign \new_[73515]_  = \new_[73514]_  & \new_[73507]_ ;
  assign \new_[73519]_  = A267 & ~A266;
  assign \new_[73520]_  = A265 & \new_[73519]_ ;
  assign \new_[73523]_  = A300 & ~A269;
  assign \new_[73526]_  = A302 & ~A301;
  assign \new_[73527]_  = \new_[73526]_  & \new_[73523]_ ;
  assign \new_[73528]_  = \new_[73527]_  & \new_[73520]_ ;
  assign \new_[73532]_  = ~A168 & ~A169;
  assign \new_[73533]_  = ~A170 & \new_[73532]_ ;
  assign \new_[73536]_  = ~A166 & A167;
  assign \new_[73539]_  = A200 & A199;
  assign \new_[73540]_  = \new_[73539]_  & \new_[73536]_ ;
  assign \new_[73541]_  = \new_[73540]_  & \new_[73533]_ ;
  assign \new_[73545]_  = ~A267 & ~A266;
  assign \new_[73546]_  = A265 & \new_[73545]_ ;
  assign \new_[73549]_  = A269 & ~A268;
  assign \new_[73552]_  = A301 & ~A300;
  assign \new_[73553]_  = \new_[73552]_  & \new_[73549]_ ;
  assign \new_[73554]_  = \new_[73553]_  & \new_[73546]_ ;
  assign \new_[73558]_  = ~A168 & ~A169;
  assign \new_[73559]_  = ~A170 & \new_[73558]_ ;
  assign \new_[73562]_  = ~A166 & A167;
  assign \new_[73565]_  = A200 & A199;
  assign \new_[73566]_  = \new_[73565]_  & \new_[73562]_ ;
  assign \new_[73567]_  = \new_[73566]_  & \new_[73559]_ ;
  assign \new_[73571]_  = ~A267 & ~A266;
  assign \new_[73572]_  = A265 & \new_[73571]_ ;
  assign \new_[73575]_  = A269 & ~A268;
  assign \new_[73578]_  = ~A302 & ~A300;
  assign \new_[73579]_  = \new_[73578]_  & \new_[73575]_ ;
  assign \new_[73580]_  = \new_[73579]_  & \new_[73572]_ ;
  assign \new_[73584]_  = ~A168 & ~A169;
  assign \new_[73585]_  = ~A170 & \new_[73584]_ ;
  assign \new_[73588]_  = ~A166 & A167;
  assign \new_[73591]_  = A200 & A199;
  assign \new_[73592]_  = \new_[73591]_  & \new_[73588]_ ;
  assign \new_[73593]_  = \new_[73592]_  & \new_[73585]_ ;
  assign \new_[73597]_  = ~A267 & ~A266;
  assign \new_[73598]_  = A265 & \new_[73597]_ ;
  assign \new_[73601]_  = A269 & ~A268;
  assign \new_[73604]_  = A299 & A298;
  assign \new_[73605]_  = \new_[73604]_  & \new_[73601]_ ;
  assign \new_[73606]_  = \new_[73605]_  & \new_[73598]_ ;
  assign \new_[73610]_  = ~A168 & ~A169;
  assign \new_[73611]_  = ~A170 & \new_[73610]_ ;
  assign \new_[73614]_  = ~A166 & A167;
  assign \new_[73617]_  = A200 & A199;
  assign \new_[73618]_  = \new_[73617]_  & \new_[73614]_ ;
  assign \new_[73619]_  = \new_[73618]_  & \new_[73611]_ ;
  assign \new_[73623]_  = ~A267 & ~A266;
  assign \new_[73624]_  = A265 & \new_[73623]_ ;
  assign \new_[73627]_  = A269 & ~A268;
  assign \new_[73630]_  = ~A299 & ~A298;
  assign \new_[73631]_  = \new_[73630]_  & \new_[73627]_ ;
  assign \new_[73632]_  = \new_[73631]_  & \new_[73624]_ ;
  assign \new_[73636]_  = ~A168 & ~A169;
  assign \new_[73637]_  = ~A170 & \new_[73636]_ ;
  assign \new_[73640]_  = ~A166 & A167;
  assign \new_[73643]_  = A200 & A199;
  assign \new_[73644]_  = \new_[73643]_  & \new_[73640]_ ;
  assign \new_[73645]_  = \new_[73644]_  & \new_[73637]_ ;
  assign \new_[73649]_  = A298 & ~A266;
  assign \new_[73650]_  = ~A265 & \new_[73649]_ ;
  assign \new_[73653]_  = ~A300 & ~A299;
  assign \new_[73656]_  = A302 & ~A301;
  assign \new_[73657]_  = \new_[73656]_  & \new_[73653]_ ;
  assign \new_[73658]_  = \new_[73657]_  & \new_[73650]_ ;
  assign \new_[73662]_  = ~A168 & ~A169;
  assign \new_[73663]_  = ~A170 & \new_[73662]_ ;
  assign \new_[73666]_  = ~A166 & A167;
  assign \new_[73669]_  = A200 & A199;
  assign \new_[73670]_  = \new_[73669]_  & \new_[73666]_ ;
  assign \new_[73671]_  = \new_[73670]_  & \new_[73663]_ ;
  assign \new_[73675]_  = ~A298 & ~A266;
  assign \new_[73676]_  = ~A265 & \new_[73675]_ ;
  assign \new_[73679]_  = ~A300 & A299;
  assign \new_[73682]_  = A302 & ~A301;
  assign \new_[73683]_  = \new_[73682]_  & \new_[73679]_ ;
  assign \new_[73684]_  = \new_[73683]_  & \new_[73676]_ ;
  assign \new_[73688]_  = ~A168 & ~A169;
  assign \new_[73689]_  = ~A170 & \new_[73688]_ ;
  assign \new_[73692]_  = ~A166 & A167;
  assign \new_[73695]_  = ~A200 & ~A199;
  assign \new_[73696]_  = \new_[73695]_  & \new_[73692]_ ;
  assign \new_[73697]_  = \new_[73696]_  & \new_[73689]_ ;
  assign \new_[73701]_  = A269 & ~A268;
  assign \new_[73702]_  = A267 & \new_[73701]_ ;
  assign \new_[73705]_  = ~A299 & A298;
  assign \new_[73708]_  = A301 & A300;
  assign \new_[73709]_  = \new_[73708]_  & \new_[73705]_ ;
  assign \new_[73710]_  = \new_[73709]_  & \new_[73702]_ ;
  assign \new_[73714]_  = ~A168 & ~A169;
  assign \new_[73715]_  = ~A170 & \new_[73714]_ ;
  assign \new_[73718]_  = ~A166 & A167;
  assign \new_[73721]_  = ~A200 & ~A199;
  assign \new_[73722]_  = \new_[73721]_  & \new_[73718]_ ;
  assign \new_[73723]_  = \new_[73722]_  & \new_[73715]_ ;
  assign \new_[73727]_  = A269 & ~A268;
  assign \new_[73728]_  = A267 & \new_[73727]_ ;
  assign \new_[73731]_  = ~A299 & A298;
  assign \new_[73734]_  = ~A302 & A300;
  assign \new_[73735]_  = \new_[73734]_  & \new_[73731]_ ;
  assign \new_[73736]_  = \new_[73735]_  & \new_[73728]_ ;
  assign \new_[73740]_  = ~A168 & ~A169;
  assign \new_[73741]_  = ~A170 & \new_[73740]_ ;
  assign \new_[73744]_  = ~A166 & A167;
  assign \new_[73747]_  = ~A200 & ~A199;
  assign \new_[73748]_  = \new_[73747]_  & \new_[73744]_ ;
  assign \new_[73749]_  = \new_[73748]_  & \new_[73741]_ ;
  assign \new_[73753]_  = A269 & ~A268;
  assign \new_[73754]_  = A267 & \new_[73753]_ ;
  assign \new_[73757]_  = A299 & ~A298;
  assign \new_[73760]_  = A301 & A300;
  assign \new_[73761]_  = \new_[73760]_  & \new_[73757]_ ;
  assign \new_[73762]_  = \new_[73761]_  & \new_[73754]_ ;
  assign \new_[73766]_  = ~A168 & ~A169;
  assign \new_[73767]_  = ~A170 & \new_[73766]_ ;
  assign \new_[73770]_  = ~A166 & A167;
  assign \new_[73773]_  = ~A200 & ~A199;
  assign \new_[73774]_  = \new_[73773]_  & \new_[73770]_ ;
  assign \new_[73775]_  = \new_[73774]_  & \new_[73767]_ ;
  assign \new_[73779]_  = A269 & ~A268;
  assign \new_[73780]_  = A267 & \new_[73779]_ ;
  assign \new_[73783]_  = A299 & ~A298;
  assign \new_[73786]_  = ~A302 & A300;
  assign \new_[73787]_  = \new_[73786]_  & \new_[73783]_ ;
  assign \new_[73788]_  = \new_[73787]_  & \new_[73780]_ ;
  assign \new_[73792]_  = ~A168 & ~A169;
  assign \new_[73793]_  = ~A170 & \new_[73792]_ ;
  assign \new_[73796]_  = ~A166 & A167;
  assign \new_[73799]_  = ~A200 & ~A199;
  assign \new_[73800]_  = \new_[73799]_  & \new_[73796]_ ;
  assign \new_[73801]_  = \new_[73800]_  & \new_[73793]_ ;
  assign \new_[73805]_  = A298 & A268;
  assign \new_[73806]_  = ~A267 & \new_[73805]_ ;
  assign \new_[73809]_  = ~A300 & ~A299;
  assign \new_[73812]_  = A302 & ~A301;
  assign \new_[73813]_  = \new_[73812]_  & \new_[73809]_ ;
  assign \new_[73814]_  = \new_[73813]_  & \new_[73806]_ ;
  assign \new_[73818]_  = ~A168 & ~A169;
  assign \new_[73819]_  = ~A170 & \new_[73818]_ ;
  assign \new_[73822]_  = ~A166 & A167;
  assign \new_[73825]_  = ~A200 & ~A199;
  assign \new_[73826]_  = \new_[73825]_  & \new_[73822]_ ;
  assign \new_[73827]_  = \new_[73826]_  & \new_[73819]_ ;
  assign \new_[73831]_  = ~A298 & A268;
  assign \new_[73832]_  = ~A267 & \new_[73831]_ ;
  assign \new_[73835]_  = ~A300 & A299;
  assign \new_[73838]_  = A302 & ~A301;
  assign \new_[73839]_  = \new_[73838]_  & \new_[73835]_ ;
  assign \new_[73840]_  = \new_[73839]_  & \new_[73832]_ ;
  assign \new_[73844]_  = ~A168 & ~A169;
  assign \new_[73845]_  = ~A170 & \new_[73844]_ ;
  assign \new_[73848]_  = ~A166 & A167;
  assign \new_[73851]_  = ~A200 & ~A199;
  assign \new_[73852]_  = \new_[73851]_  & \new_[73848]_ ;
  assign \new_[73853]_  = \new_[73852]_  & \new_[73845]_ ;
  assign \new_[73857]_  = A298 & ~A269;
  assign \new_[73858]_  = ~A267 & \new_[73857]_ ;
  assign \new_[73861]_  = ~A300 & ~A299;
  assign \new_[73864]_  = A302 & ~A301;
  assign \new_[73865]_  = \new_[73864]_  & \new_[73861]_ ;
  assign \new_[73866]_  = \new_[73865]_  & \new_[73858]_ ;
  assign \new_[73870]_  = ~A168 & ~A169;
  assign \new_[73871]_  = ~A170 & \new_[73870]_ ;
  assign \new_[73874]_  = ~A166 & A167;
  assign \new_[73877]_  = ~A200 & ~A199;
  assign \new_[73878]_  = \new_[73877]_  & \new_[73874]_ ;
  assign \new_[73879]_  = \new_[73878]_  & \new_[73871]_ ;
  assign \new_[73883]_  = ~A298 & ~A269;
  assign \new_[73884]_  = ~A267 & \new_[73883]_ ;
  assign \new_[73887]_  = ~A300 & A299;
  assign \new_[73890]_  = A302 & ~A301;
  assign \new_[73891]_  = \new_[73890]_  & \new_[73887]_ ;
  assign \new_[73892]_  = \new_[73891]_  & \new_[73884]_ ;
  assign \new_[73896]_  = ~A168 & ~A169;
  assign \new_[73897]_  = ~A170 & \new_[73896]_ ;
  assign \new_[73900]_  = ~A166 & A167;
  assign \new_[73903]_  = ~A200 & ~A199;
  assign \new_[73904]_  = \new_[73903]_  & \new_[73900]_ ;
  assign \new_[73905]_  = \new_[73904]_  & \new_[73897]_ ;
  assign \new_[73909]_  = A298 & A266;
  assign \new_[73910]_  = A265 & \new_[73909]_ ;
  assign \new_[73913]_  = ~A300 & ~A299;
  assign \new_[73916]_  = A302 & ~A301;
  assign \new_[73917]_  = \new_[73916]_  & \new_[73913]_ ;
  assign \new_[73918]_  = \new_[73917]_  & \new_[73910]_ ;
  assign \new_[73922]_  = ~A168 & ~A169;
  assign \new_[73923]_  = ~A170 & \new_[73922]_ ;
  assign \new_[73926]_  = ~A166 & A167;
  assign \new_[73929]_  = ~A200 & ~A199;
  assign \new_[73930]_  = \new_[73929]_  & \new_[73926]_ ;
  assign \new_[73931]_  = \new_[73930]_  & \new_[73923]_ ;
  assign \new_[73935]_  = ~A298 & A266;
  assign \new_[73936]_  = A265 & \new_[73935]_ ;
  assign \new_[73939]_  = ~A300 & A299;
  assign \new_[73942]_  = A302 & ~A301;
  assign \new_[73943]_  = \new_[73942]_  & \new_[73939]_ ;
  assign \new_[73944]_  = \new_[73943]_  & \new_[73936]_ ;
  assign \new_[73948]_  = ~A168 & ~A169;
  assign \new_[73949]_  = ~A170 & \new_[73948]_ ;
  assign \new_[73952]_  = ~A166 & A167;
  assign \new_[73955]_  = ~A200 & ~A199;
  assign \new_[73956]_  = \new_[73955]_  & \new_[73952]_ ;
  assign \new_[73957]_  = \new_[73956]_  & \new_[73949]_ ;
  assign \new_[73961]_  = A267 & A266;
  assign \new_[73962]_  = ~A265 & \new_[73961]_ ;
  assign \new_[73965]_  = A300 & A268;
  assign \new_[73968]_  = A302 & ~A301;
  assign \new_[73969]_  = \new_[73968]_  & \new_[73965]_ ;
  assign \new_[73970]_  = \new_[73969]_  & \new_[73962]_ ;
  assign \new_[73974]_  = ~A168 & ~A169;
  assign \new_[73975]_  = ~A170 & \new_[73974]_ ;
  assign \new_[73978]_  = ~A166 & A167;
  assign \new_[73981]_  = ~A200 & ~A199;
  assign \new_[73982]_  = \new_[73981]_  & \new_[73978]_ ;
  assign \new_[73983]_  = \new_[73982]_  & \new_[73975]_ ;
  assign \new_[73987]_  = A267 & A266;
  assign \new_[73988]_  = ~A265 & \new_[73987]_ ;
  assign \new_[73991]_  = A300 & ~A269;
  assign \new_[73994]_  = A302 & ~A301;
  assign \new_[73995]_  = \new_[73994]_  & \new_[73991]_ ;
  assign \new_[73996]_  = \new_[73995]_  & \new_[73988]_ ;
  assign \new_[74000]_  = ~A168 & ~A169;
  assign \new_[74001]_  = ~A170 & \new_[74000]_ ;
  assign \new_[74004]_  = ~A166 & A167;
  assign \new_[74007]_  = ~A200 & ~A199;
  assign \new_[74008]_  = \new_[74007]_  & \new_[74004]_ ;
  assign \new_[74009]_  = \new_[74008]_  & \new_[74001]_ ;
  assign \new_[74013]_  = ~A267 & A266;
  assign \new_[74014]_  = ~A265 & \new_[74013]_ ;
  assign \new_[74017]_  = A269 & ~A268;
  assign \new_[74020]_  = A301 & ~A300;
  assign \new_[74021]_  = \new_[74020]_  & \new_[74017]_ ;
  assign \new_[74022]_  = \new_[74021]_  & \new_[74014]_ ;
  assign \new_[74026]_  = ~A168 & ~A169;
  assign \new_[74027]_  = ~A170 & \new_[74026]_ ;
  assign \new_[74030]_  = ~A166 & A167;
  assign \new_[74033]_  = ~A200 & ~A199;
  assign \new_[74034]_  = \new_[74033]_  & \new_[74030]_ ;
  assign \new_[74035]_  = \new_[74034]_  & \new_[74027]_ ;
  assign \new_[74039]_  = ~A267 & A266;
  assign \new_[74040]_  = ~A265 & \new_[74039]_ ;
  assign \new_[74043]_  = A269 & ~A268;
  assign \new_[74046]_  = ~A302 & ~A300;
  assign \new_[74047]_  = \new_[74046]_  & \new_[74043]_ ;
  assign \new_[74048]_  = \new_[74047]_  & \new_[74040]_ ;
  assign \new_[74052]_  = ~A168 & ~A169;
  assign \new_[74053]_  = ~A170 & \new_[74052]_ ;
  assign \new_[74056]_  = ~A166 & A167;
  assign \new_[74059]_  = ~A200 & ~A199;
  assign \new_[74060]_  = \new_[74059]_  & \new_[74056]_ ;
  assign \new_[74061]_  = \new_[74060]_  & \new_[74053]_ ;
  assign \new_[74065]_  = ~A267 & A266;
  assign \new_[74066]_  = ~A265 & \new_[74065]_ ;
  assign \new_[74069]_  = A269 & ~A268;
  assign \new_[74072]_  = A299 & A298;
  assign \new_[74073]_  = \new_[74072]_  & \new_[74069]_ ;
  assign \new_[74074]_  = \new_[74073]_  & \new_[74066]_ ;
  assign \new_[74078]_  = ~A168 & ~A169;
  assign \new_[74079]_  = ~A170 & \new_[74078]_ ;
  assign \new_[74082]_  = ~A166 & A167;
  assign \new_[74085]_  = ~A200 & ~A199;
  assign \new_[74086]_  = \new_[74085]_  & \new_[74082]_ ;
  assign \new_[74087]_  = \new_[74086]_  & \new_[74079]_ ;
  assign \new_[74091]_  = ~A267 & A266;
  assign \new_[74092]_  = ~A265 & \new_[74091]_ ;
  assign \new_[74095]_  = A269 & ~A268;
  assign \new_[74098]_  = ~A299 & ~A298;
  assign \new_[74099]_  = \new_[74098]_  & \new_[74095]_ ;
  assign \new_[74100]_  = \new_[74099]_  & \new_[74092]_ ;
  assign \new_[74104]_  = ~A168 & ~A169;
  assign \new_[74105]_  = ~A170 & \new_[74104]_ ;
  assign \new_[74108]_  = ~A166 & A167;
  assign \new_[74111]_  = ~A200 & ~A199;
  assign \new_[74112]_  = \new_[74111]_  & \new_[74108]_ ;
  assign \new_[74113]_  = \new_[74112]_  & \new_[74105]_ ;
  assign \new_[74117]_  = A267 & ~A266;
  assign \new_[74118]_  = A265 & \new_[74117]_ ;
  assign \new_[74121]_  = A300 & A268;
  assign \new_[74124]_  = A302 & ~A301;
  assign \new_[74125]_  = \new_[74124]_  & \new_[74121]_ ;
  assign \new_[74126]_  = \new_[74125]_  & \new_[74118]_ ;
  assign \new_[74130]_  = ~A168 & ~A169;
  assign \new_[74131]_  = ~A170 & \new_[74130]_ ;
  assign \new_[74134]_  = ~A166 & A167;
  assign \new_[74137]_  = ~A200 & ~A199;
  assign \new_[74138]_  = \new_[74137]_  & \new_[74134]_ ;
  assign \new_[74139]_  = \new_[74138]_  & \new_[74131]_ ;
  assign \new_[74143]_  = A267 & ~A266;
  assign \new_[74144]_  = A265 & \new_[74143]_ ;
  assign \new_[74147]_  = A300 & ~A269;
  assign \new_[74150]_  = A302 & ~A301;
  assign \new_[74151]_  = \new_[74150]_  & \new_[74147]_ ;
  assign \new_[74152]_  = \new_[74151]_  & \new_[74144]_ ;
  assign \new_[74156]_  = ~A168 & ~A169;
  assign \new_[74157]_  = ~A170 & \new_[74156]_ ;
  assign \new_[74160]_  = ~A166 & A167;
  assign \new_[74163]_  = ~A200 & ~A199;
  assign \new_[74164]_  = \new_[74163]_  & \new_[74160]_ ;
  assign \new_[74165]_  = \new_[74164]_  & \new_[74157]_ ;
  assign \new_[74169]_  = ~A267 & ~A266;
  assign \new_[74170]_  = A265 & \new_[74169]_ ;
  assign \new_[74173]_  = A269 & ~A268;
  assign \new_[74176]_  = A301 & ~A300;
  assign \new_[74177]_  = \new_[74176]_  & \new_[74173]_ ;
  assign \new_[74178]_  = \new_[74177]_  & \new_[74170]_ ;
  assign \new_[74182]_  = ~A168 & ~A169;
  assign \new_[74183]_  = ~A170 & \new_[74182]_ ;
  assign \new_[74186]_  = ~A166 & A167;
  assign \new_[74189]_  = ~A200 & ~A199;
  assign \new_[74190]_  = \new_[74189]_  & \new_[74186]_ ;
  assign \new_[74191]_  = \new_[74190]_  & \new_[74183]_ ;
  assign \new_[74195]_  = ~A267 & ~A266;
  assign \new_[74196]_  = A265 & \new_[74195]_ ;
  assign \new_[74199]_  = A269 & ~A268;
  assign \new_[74202]_  = ~A302 & ~A300;
  assign \new_[74203]_  = \new_[74202]_  & \new_[74199]_ ;
  assign \new_[74204]_  = \new_[74203]_  & \new_[74196]_ ;
  assign \new_[74208]_  = ~A168 & ~A169;
  assign \new_[74209]_  = ~A170 & \new_[74208]_ ;
  assign \new_[74212]_  = ~A166 & A167;
  assign \new_[74215]_  = ~A200 & ~A199;
  assign \new_[74216]_  = \new_[74215]_  & \new_[74212]_ ;
  assign \new_[74217]_  = \new_[74216]_  & \new_[74209]_ ;
  assign \new_[74221]_  = ~A267 & ~A266;
  assign \new_[74222]_  = A265 & \new_[74221]_ ;
  assign \new_[74225]_  = A269 & ~A268;
  assign \new_[74228]_  = A299 & A298;
  assign \new_[74229]_  = \new_[74228]_  & \new_[74225]_ ;
  assign \new_[74230]_  = \new_[74229]_  & \new_[74222]_ ;
  assign \new_[74234]_  = ~A168 & ~A169;
  assign \new_[74235]_  = ~A170 & \new_[74234]_ ;
  assign \new_[74238]_  = ~A166 & A167;
  assign \new_[74241]_  = ~A200 & ~A199;
  assign \new_[74242]_  = \new_[74241]_  & \new_[74238]_ ;
  assign \new_[74243]_  = \new_[74242]_  & \new_[74235]_ ;
  assign \new_[74247]_  = ~A267 & ~A266;
  assign \new_[74248]_  = A265 & \new_[74247]_ ;
  assign \new_[74251]_  = A269 & ~A268;
  assign \new_[74254]_  = ~A299 & ~A298;
  assign \new_[74255]_  = \new_[74254]_  & \new_[74251]_ ;
  assign \new_[74256]_  = \new_[74255]_  & \new_[74248]_ ;
  assign \new_[74260]_  = ~A168 & ~A169;
  assign \new_[74261]_  = ~A170 & \new_[74260]_ ;
  assign \new_[74264]_  = ~A166 & A167;
  assign \new_[74267]_  = ~A200 & ~A199;
  assign \new_[74268]_  = \new_[74267]_  & \new_[74264]_ ;
  assign \new_[74269]_  = \new_[74268]_  & \new_[74261]_ ;
  assign \new_[74273]_  = A298 & ~A266;
  assign \new_[74274]_  = ~A265 & \new_[74273]_ ;
  assign \new_[74277]_  = ~A300 & ~A299;
  assign \new_[74280]_  = A302 & ~A301;
  assign \new_[74281]_  = \new_[74280]_  & \new_[74277]_ ;
  assign \new_[74282]_  = \new_[74281]_  & \new_[74274]_ ;
  assign \new_[74286]_  = ~A168 & ~A169;
  assign \new_[74287]_  = ~A170 & \new_[74286]_ ;
  assign \new_[74290]_  = ~A166 & A167;
  assign \new_[74293]_  = ~A200 & ~A199;
  assign \new_[74294]_  = \new_[74293]_  & \new_[74290]_ ;
  assign \new_[74295]_  = \new_[74294]_  & \new_[74287]_ ;
  assign \new_[74299]_  = ~A298 & ~A266;
  assign \new_[74300]_  = ~A265 & \new_[74299]_ ;
  assign \new_[74303]_  = ~A300 & A299;
  assign \new_[74306]_  = A302 & ~A301;
  assign \new_[74307]_  = \new_[74306]_  & \new_[74303]_ ;
  assign \new_[74308]_  = \new_[74307]_  & \new_[74300]_ ;
  assign \new_[74312]_  = ~A168 & ~A169;
  assign \new_[74313]_  = ~A170 & \new_[74312]_ ;
  assign \new_[74316]_  = A166 & ~A167;
  assign \new_[74319]_  = ~A202 & A201;
  assign \new_[74320]_  = \new_[74319]_  & \new_[74316]_ ;
  assign \new_[74321]_  = \new_[74320]_  & \new_[74313]_ ;
  assign \new_[74325]_  = A268 & ~A267;
  assign \new_[74326]_  = A203 & \new_[74325]_ ;
  assign \new_[74329]_  = ~A299 & A298;
  assign \new_[74332]_  = A301 & A300;
  assign \new_[74333]_  = \new_[74332]_  & \new_[74329]_ ;
  assign \new_[74334]_  = \new_[74333]_  & \new_[74326]_ ;
  assign \new_[74338]_  = ~A168 & ~A169;
  assign \new_[74339]_  = ~A170 & \new_[74338]_ ;
  assign \new_[74342]_  = A166 & ~A167;
  assign \new_[74345]_  = ~A202 & A201;
  assign \new_[74346]_  = \new_[74345]_  & \new_[74342]_ ;
  assign \new_[74347]_  = \new_[74346]_  & \new_[74339]_ ;
  assign \new_[74351]_  = A268 & ~A267;
  assign \new_[74352]_  = A203 & \new_[74351]_ ;
  assign \new_[74355]_  = ~A299 & A298;
  assign \new_[74358]_  = ~A302 & A300;
  assign \new_[74359]_  = \new_[74358]_  & \new_[74355]_ ;
  assign \new_[74360]_  = \new_[74359]_  & \new_[74352]_ ;
  assign \new_[74364]_  = ~A168 & ~A169;
  assign \new_[74365]_  = ~A170 & \new_[74364]_ ;
  assign \new_[74368]_  = A166 & ~A167;
  assign \new_[74371]_  = ~A202 & A201;
  assign \new_[74372]_  = \new_[74371]_  & \new_[74368]_ ;
  assign \new_[74373]_  = \new_[74372]_  & \new_[74365]_ ;
  assign \new_[74377]_  = A268 & ~A267;
  assign \new_[74378]_  = A203 & \new_[74377]_ ;
  assign \new_[74381]_  = A299 & ~A298;
  assign \new_[74384]_  = A301 & A300;
  assign \new_[74385]_  = \new_[74384]_  & \new_[74381]_ ;
  assign \new_[74386]_  = \new_[74385]_  & \new_[74378]_ ;
  assign \new_[74390]_  = ~A168 & ~A169;
  assign \new_[74391]_  = ~A170 & \new_[74390]_ ;
  assign \new_[74394]_  = A166 & ~A167;
  assign \new_[74397]_  = ~A202 & A201;
  assign \new_[74398]_  = \new_[74397]_  & \new_[74394]_ ;
  assign \new_[74399]_  = \new_[74398]_  & \new_[74391]_ ;
  assign \new_[74403]_  = A268 & ~A267;
  assign \new_[74404]_  = A203 & \new_[74403]_ ;
  assign \new_[74407]_  = A299 & ~A298;
  assign \new_[74410]_  = ~A302 & A300;
  assign \new_[74411]_  = \new_[74410]_  & \new_[74407]_ ;
  assign \new_[74412]_  = \new_[74411]_  & \new_[74404]_ ;
  assign \new_[74416]_  = ~A168 & ~A169;
  assign \new_[74417]_  = ~A170 & \new_[74416]_ ;
  assign \new_[74420]_  = A166 & ~A167;
  assign \new_[74423]_  = ~A202 & A201;
  assign \new_[74424]_  = \new_[74423]_  & \new_[74420]_ ;
  assign \new_[74425]_  = \new_[74424]_  & \new_[74417]_ ;
  assign \new_[74429]_  = ~A269 & ~A267;
  assign \new_[74430]_  = A203 & \new_[74429]_ ;
  assign \new_[74433]_  = ~A299 & A298;
  assign \new_[74436]_  = A301 & A300;
  assign \new_[74437]_  = \new_[74436]_  & \new_[74433]_ ;
  assign \new_[74438]_  = \new_[74437]_  & \new_[74430]_ ;
  assign \new_[74442]_  = ~A168 & ~A169;
  assign \new_[74443]_  = ~A170 & \new_[74442]_ ;
  assign \new_[74446]_  = A166 & ~A167;
  assign \new_[74449]_  = ~A202 & A201;
  assign \new_[74450]_  = \new_[74449]_  & \new_[74446]_ ;
  assign \new_[74451]_  = \new_[74450]_  & \new_[74443]_ ;
  assign \new_[74455]_  = ~A269 & ~A267;
  assign \new_[74456]_  = A203 & \new_[74455]_ ;
  assign \new_[74459]_  = ~A299 & A298;
  assign \new_[74462]_  = ~A302 & A300;
  assign \new_[74463]_  = \new_[74462]_  & \new_[74459]_ ;
  assign \new_[74464]_  = \new_[74463]_  & \new_[74456]_ ;
  assign \new_[74468]_  = ~A168 & ~A169;
  assign \new_[74469]_  = ~A170 & \new_[74468]_ ;
  assign \new_[74472]_  = A166 & ~A167;
  assign \new_[74475]_  = ~A202 & A201;
  assign \new_[74476]_  = \new_[74475]_  & \new_[74472]_ ;
  assign \new_[74477]_  = \new_[74476]_  & \new_[74469]_ ;
  assign \new_[74481]_  = ~A269 & ~A267;
  assign \new_[74482]_  = A203 & \new_[74481]_ ;
  assign \new_[74485]_  = A299 & ~A298;
  assign \new_[74488]_  = A301 & A300;
  assign \new_[74489]_  = \new_[74488]_  & \new_[74485]_ ;
  assign \new_[74490]_  = \new_[74489]_  & \new_[74482]_ ;
  assign \new_[74494]_  = ~A168 & ~A169;
  assign \new_[74495]_  = ~A170 & \new_[74494]_ ;
  assign \new_[74498]_  = A166 & ~A167;
  assign \new_[74501]_  = ~A202 & A201;
  assign \new_[74502]_  = \new_[74501]_  & \new_[74498]_ ;
  assign \new_[74503]_  = \new_[74502]_  & \new_[74495]_ ;
  assign \new_[74507]_  = ~A269 & ~A267;
  assign \new_[74508]_  = A203 & \new_[74507]_ ;
  assign \new_[74511]_  = A299 & ~A298;
  assign \new_[74514]_  = ~A302 & A300;
  assign \new_[74515]_  = \new_[74514]_  & \new_[74511]_ ;
  assign \new_[74516]_  = \new_[74515]_  & \new_[74508]_ ;
  assign \new_[74520]_  = ~A168 & ~A169;
  assign \new_[74521]_  = ~A170 & \new_[74520]_ ;
  assign \new_[74524]_  = A166 & ~A167;
  assign \new_[74527]_  = ~A202 & A201;
  assign \new_[74528]_  = \new_[74527]_  & \new_[74524]_ ;
  assign \new_[74529]_  = \new_[74528]_  & \new_[74521]_ ;
  assign \new_[74533]_  = A266 & A265;
  assign \new_[74534]_  = A203 & \new_[74533]_ ;
  assign \new_[74537]_  = ~A299 & A298;
  assign \new_[74540]_  = A301 & A300;
  assign \new_[74541]_  = \new_[74540]_  & \new_[74537]_ ;
  assign \new_[74542]_  = \new_[74541]_  & \new_[74534]_ ;
  assign \new_[74546]_  = ~A168 & ~A169;
  assign \new_[74547]_  = ~A170 & \new_[74546]_ ;
  assign \new_[74550]_  = A166 & ~A167;
  assign \new_[74553]_  = ~A202 & A201;
  assign \new_[74554]_  = \new_[74553]_  & \new_[74550]_ ;
  assign \new_[74555]_  = \new_[74554]_  & \new_[74547]_ ;
  assign \new_[74559]_  = A266 & A265;
  assign \new_[74560]_  = A203 & \new_[74559]_ ;
  assign \new_[74563]_  = ~A299 & A298;
  assign \new_[74566]_  = ~A302 & A300;
  assign \new_[74567]_  = \new_[74566]_  & \new_[74563]_ ;
  assign \new_[74568]_  = \new_[74567]_  & \new_[74560]_ ;
  assign \new_[74572]_  = ~A168 & ~A169;
  assign \new_[74573]_  = ~A170 & \new_[74572]_ ;
  assign \new_[74576]_  = A166 & ~A167;
  assign \new_[74579]_  = ~A202 & A201;
  assign \new_[74580]_  = \new_[74579]_  & \new_[74576]_ ;
  assign \new_[74581]_  = \new_[74580]_  & \new_[74573]_ ;
  assign \new_[74585]_  = A266 & A265;
  assign \new_[74586]_  = A203 & \new_[74585]_ ;
  assign \new_[74589]_  = A299 & ~A298;
  assign \new_[74592]_  = A301 & A300;
  assign \new_[74593]_  = \new_[74592]_  & \new_[74589]_ ;
  assign \new_[74594]_  = \new_[74593]_  & \new_[74586]_ ;
  assign \new_[74598]_  = ~A168 & ~A169;
  assign \new_[74599]_  = ~A170 & \new_[74598]_ ;
  assign \new_[74602]_  = A166 & ~A167;
  assign \new_[74605]_  = ~A202 & A201;
  assign \new_[74606]_  = \new_[74605]_  & \new_[74602]_ ;
  assign \new_[74607]_  = \new_[74606]_  & \new_[74599]_ ;
  assign \new_[74611]_  = A266 & A265;
  assign \new_[74612]_  = A203 & \new_[74611]_ ;
  assign \new_[74615]_  = A299 & ~A298;
  assign \new_[74618]_  = ~A302 & A300;
  assign \new_[74619]_  = \new_[74618]_  & \new_[74615]_ ;
  assign \new_[74620]_  = \new_[74619]_  & \new_[74612]_ ;
  assign \new_[74624]_  = ~A168 & ~A169;
  assign \new_[74625]_  = ~A170 & \new_[74624]_ ;
  assign \new_[74628]_  = A166 & ~A167;
  assign \new_[74631]_  = ~A202 & A201;
  assign \new_[74632]_  = \new_[74631]_  & \new_[74628]_ ;
  assign \new_[74633]_  = \new_[74632]_  & \new_[74625]_ ;
  assign \new_[74637]_  = A266 & ~A265;
  assign \new_[74638]_  = A203 & \new_[74637]_ ;
  assign \new_[74641]_  = A268 & A267;
  assign \new_[74644]_  = A301 & ~A300;
  assign \new_[74645]_  = \new_[74644]_  & \new_[74641]_ ;
  assign \new_[74646]_  = \new_[74645]_  & \new_[74638]_ ;
  assign \new_[74650]_  = ~A168 & ~A169;
  assign \new_[74651]_  = ~A170 & \new_[74650]_ ;
  assign \new_[74654]_  = A166 & ~A167;
  assign \new_[74657]_  = ~A202 & A201;
  assign \new_[74658]_  = \new_[74657]_  & \new_[74654]_ ;
  assign \new_[74659]_  = \new_[74658]_  & \new_[74651]_ ;
  assign \new_[74663]_  = A266 & ~A265;
  assign \new_[74664]_  = A203 & \new_[74663]_ ;
  assign \new_[74667]_  = A268 & A267;
  assign \new_[74670]_  = ~A302 & ~A300;
  assign \new_[74671]_  = \new_[74670]_  & \new_[74667]_ ;
  assign \new_[74672]_  = \new_[74671]_  & \new_[74664]_ ;
  assign \new_[74676]_  = ~A168 & ~A169;
  assign \new_[74677]_  = ~A170 & \new_[74676]_ ;
  assign \new_[74680]_  = A166 & ~A167;
  assign \new_[74683]_  = ~A202 & A201;
  assign \new_[74684]_  = \new_[74683]_  & \new_[74680]_ ;
  assign \new_[74685]_  = \new_[74684]_  & \new_[74677]_ ;
  assign \new_[74689]_  = A266 & ~A265;
  assign \new_[74690]_  = A203 & \new_[74689]_ ;
  assign \new_[74693]_  = A268 & A267;
  assign \new_[74696]_  = A299 & A298;
  assign \new_[74697]_  = \new_[74696]_  & \new_[74693]_ ;
  assign \new_[74698]_  = \new_[74697]_  & \new_[74690]_ ;
  assign \new_[74702]_  = ~A168 & ~A169;
  assign \new_[74703]_  = ~A170 & \new_[74702]_ ;
  assign \new_[74706]_  = A166 & ~A167;
  assign \new_[74709]_  = ~A202 & A201;
  assign \new_[74710]_  = \new_[74709]_  & \new_[74706]_ ;
  assign \new_[74711]_  = \new_[74710]_  & \new_[74703]_ ;
  assign \new_[74715]_  = A266 & ~A265;
  assign \new_[74716]_  = A203 & \new_[74715]_ ;
  assign \new_[74719]_  = A268 & A267;
  assign \new_[74722]_  = ~A299 & ~A298;
  assign \new_[74723]_  = \new_[74722]_  & \new_[74719]_ ;
  assign \new_[74724]_  = \new_[74723]_  & \new_[74716]_ ;
  assign \new_[74728]_  = ~A168 & ~A169;
  assign \new_[74729]_  = ~A170 & \new_[74728]_ ;
  assign \new_[74732]_  = A166 & ~A167;
  assign \new_[74735]_  = ~A202 & A201;
  assign \new_[74736]_  = \new_[74735]_  & \new_[74732]_ ;
  assign \new_[74737]_  = \new_[74736]_  & \new_[74729]_ ;
  assign \new_[74741]_  = A266 & ~A265;
  assign \new_[74742]_  = A203 & \new_[74741]_ ;
  assign \new_[74745]_  = ~A269 & A267;
  assign \new_[74748]_  = A301 & ~A300;
  assign \new_[74749]_  = \new_[74748]_  & \new_[74745]_ ;
  assign \new_[74750]_  = \new_[74749]_  & \new_[74742]_ ;
  assign \new_[74754]_  = ~A168 & ~A169;
  assign \new_[74755]_  = ~A170 & \new_[74754]_ ;
  assign \new_[74758]_  = A166 & ~A167;
  assign \new_[74761]_  = ~A202 & A201;
  assign \new_[74762]_  = \new_[74761]_  & \new_[74758]_ ;
  assign \new_[74763]_  = \new_[74762]_  & \new_[74755]_ ;
  assign \new_[74767]_  = A266 & ~A265;
  assign \new_[74768]_  = A203 & \new_[74767]_ ;
  assign \new_[74771]_  = ~A269 & A267;
  assign \new_[74774]_  = ~A302 & ~A300;
  assign \new_[74775]_  = \new_[74774]_  & \new_[74771]_ ;
  assign \new_[74776]_  = \new_[74775]_  & \new_[74768]_ ;
  assign \new_[74780]_  = ~A168 & ~A169;
  assign \new_[74781]_  = ~A170 & \new_[74780]_ ;
  assign \new_[74784]_  = A166 & ~A167;
  assign \new_[74787]_  = ~A202 & A201;
  assign \new_[74788]_  = \new_[74787]_  & \new_[74784]_ ;
  assign \new_[74789]_  = \new_[74788]_  & \new_[74781]_ ;
  assign \new_[74793]_  = A266 & ~A265;
  assign \new_[74794]_  = A203 & \new_[74793]_ ;
  assign \new_[74797]_  = ~A269 & A267;
  assign \new_[74800]_  = A299 & A298;
  assign \new_[74801]_  = \new_[74800]_  & \new_[74797]_ ;
  assign \new_[74802]_  = \new_[74801]_  & \new_[74794]_ ;
  assign \new_[74806]_  = ~A168 & ~A169;
  assign \new_[74807]_  = ~A170 & \new_[74806]_ ;
  assign \new_[74810]_  = A166 & ~A167;
  assign \new_[74813]_  = ~A202 & A201;
  assign \new_[74814]_  = \new_[74813]_  & \new_[74810]_ ;
  assign \new_[74815]_  = \new_[74814]_  & \new_[74807]_ ;
  assign \new_[74819]_  = A266 & ~A265;
  assign \new_[74820]_  = A203 & \new_[74819]_ ;
  assign \new_[74823]_  = ~A269 & A267;
  assign \new_[74826]_  = ~A299 & ~A298;
  assign \new_[74827]_  = \new_[74826]_  & \new_[74823]_ ;
  assign \new_[74828]_  = \new_[74827]_  & \new_[74820]_ ;
  assign \new_[74832]_  = ~A168 & ~A169;
  assign \new_[74833]_  = ~A170 & \new_[74832]_ ;
  assign \new_[74836]_  = A166 & ~A167;
  assign \new_[74839]_  = ~A202 & A201;
  assign \new_[74840]_  = \new_[74839]_  & \new_[74836]_ ;
  assign \new_[74841]_  = \new_[74840]_  & \new_[74833]_ ;
  assign \new_[74845]_  = ~A266 & A265;
  assign \new_[74846]_  = A203 & \new_[74845]_ ;
  assign \new_[74849]_  = A268 & A267;
  assign \new_[74852]_  = A301 & ~A300;
  assign \new_[74853]_  = \new_[74852]_  & \new_[74849]_ ;
  assign \new_[74854]_  = \new_[74853]_  & \new_[74846]_ ;
  assign \new_[74858]_  = ~A168 & ~A169;
  assign \new_[74859]_  = ~A170 & \new_[74858]_ ;
  assign \new_[74862]_  = A166 & ~A167;
  assign \new_[74865]_  = ~A202 & A201;
  assign \new_[74866]_  = \new_[74865]_  & \new_[74862]_ ;
  assign \new_[74867]_  = \new_[74866]_  & \new_[74859]_ ;
  assign \new_[74871]_  = ~A266 & A265;
  assign \new_[74872]_  = A203 & \new_[74871]_ ;
  assign \new_[74875]_  = A268 & A267;
  assign \new_[74878]_  = ~A302 & ~A300;
  assign \new_[74879]_  = \new_[74878]_  & \new_[74875]_ ;
  assign \new_[74880]_  = \new_[74879]_  & \new_[74872]_ ;
  assign \new_[74884]_  = ~A168 & ~A169;
  assign \new_[74885]_  = ~A170 & \new_[74884]_ ;
  assign \new_[74888]_  = A166 & ~A167;
  assign \new_[74891]_  = ~A202 & A201;
  assign \new_[74892]_  = \new_[74891]_  & \new_[74888]_ ;
  assign \new_[74893]_  = \new_[74892]_  & \new_[74885]_ ;
  assign \new_[74897]_  = ~A266 & A265;
  assign \new_[74898]_  = A203 & \new_[74897]_ ;
  assign \new_[74901]_  = A268 & A267;
  assign \new_[74904]_  = A299 & A298;
  assign \new_[74905]_  = \new_[74904]_  & \new_[74901]_ ;
  assign \new_[74906]_  = \new_[74905]_  & \new_[74898]_ ;
  assign \new_[74910]_  = ~A168 & ~A169;
  assign \new_[74911]_  = ~A170 & \new_[74910]_ ;
  assign \new_[74914]_  = A166 & ~A167;
  assign \new_[74917]_  = ~A202 & A201;
  assign \new_[74918]_  = \new_[74917]_  & \new_[74914]_ ;
  assign \new_[74919]_  = \new_[74918]_  & \new_[74911]_ ;
  assign \new_[74923]_  = ~A266 & A265;
  assign \new_[74924]_  = A203 & \new_[74923]_ ;
  assign \new_[74927]_  = A268 & A267;
  assign \new_[74930]_  = ~A299 & ~A298;
  assign \new_[74931]_  = \new_[74930]_  & \new_[74927]_ ;
  assign \new_[74932]_  = \new_[74931]_  & \new_[74924]_ ;
  assign \new_[74936]_  = ~A168 & ~A169;
  assign \new_[74937]_  = ~A170 & \new_[74936]_ ;
  assign \new_[74940]_  = A166 & ~A167;
  assign \new_[74943]_  = ~A202 & A201;
  assign \new_[74944]_  = \new_[74943]_  & \new_[74940]_ ;
  assign \new_[74945]_  = \new_[74944]_  & \new_[74937]_ ;
  assign \new_[74949]_  = ~A266 & A265;
  assign \new_[74950]_  = A203 & \new_[74949]_ ;
  assign \new_[74953]_  = ~A269 & A267;
  assign \new_[74956]_  = A301 & ~A300;
  assign \new_[74957]_  = \new_[74956]_  & \new_[74953]_ ;
  assign \new_[74958]_  = \new_[74957]_  & \new_[74950]_ ;
  assign \new_[74962]_  = ~A168 & ~A169;
  assign \new_[74963]_  = ~A170 & \new_[74962]_ ;
  assign \new_[74966]_  = A166 & ~A167;
  assign \new_[74969]_  = ~A202 & A201;
  assign \new_[74970]_  = \new_[74969]_  & \new_[74966]_ ;
  assign \new_[74971]_  = \new_[74970]_  & \new_[74963]_ ;
  assign \new_[74975]_  = ~A266 & A265;
  assign \new_[74976]_  = A203 & \new_[74975]_ ;
  assign \new_[74979]_  = ~A269 & A267;
  assign \new_[74982]_  = ~A302 & ~A300;
  assign \new_[74983]_  = \new_[74982]_  & \new_[74979]_ ;
  assign \new_[74984]_  = \new_[74983]_  & \new_[74976]_ ;
  assign \new_[74988]_  = ~A168 & ~A169;
  assign \new_[74989]_  = ~A170 & \new_[74988]_ ;
  assign \new_[74992]_  = A166 & ~A167;
  assign \new_[74995]_  = ~A202 & A201;
  assign \new_[74996]_  = \new_[74995]_  & \new_[74992]_ ;
  assign \new_[74997]_  = \new_[74996]_  & \new_[74989]_ ;
  assign \new_[75001]_  = ~A266 & A265;
  assign \new_[75002]_  = A203 & \new_[75001]_ ;
  assign \new_[75005]_  = ~A269 & A267;
  assign \new_[75008]_  = A299 & A298;
  assign \new_[75009]_  = \new_[75008]_  & \new_[75005]_ ;
  assign \new_[75010]_  = \new_[75009]_  & \new_[75002]_ ;
  assign \new_[75014]_  = ~A168 & ~A169;
  assign \new_[75015]_  = ~A170 & \new_[75014]_ ;
  assign \new_[75018]_  = A166 & ~A167;
  assign \new_[75021]_  = ~A202 & A201;
  assign \new_[75022]_  = \new_[75021]_  & \new_[75018]_ ;
  assign \new_[75023]_  = \new_[75022]_  & \new_[75015]_ ;
  assign \new_[75027]_  = ~A266 & A265;
  assign \new_[75028]_  = A203 & \new_[75027]_ ;
  assign \new_[75031]_  = ~A269 & A267;
  assign \new_[75034]_  = ~A299 & ~A298;
  assign \new_[75035]_  = \new_[75034]_  & \new_[75031]_ ;
  assign \new_[75036]_  = \new_[75035]_  & \new_[75028]_ ;
  assign \new_[75040]_  = ~A168 & ~A169;
  assign \new_[75041]_  = ~A170 & \new_[75040]_ ;
  assign \new_[75044]_  = A166 & ~A167;
  assign \new_[75047]_  = ~A202 & A201;
  assign \new_[75048]_  = \new_[75047]_  & \new_[75044]_ ;
  assign \new_[75049]_  = \new_[75048]_  & \new_[75041]_ ;
  assign \new_[75053]_  = ~A266 & ~A265;
  assign \new_[75054]_  = A203 & \new_[75053]_ ;
  assign \new_[75057]_  = ~A299 & A298;
  assign \new_[75060]_  = A301 & A300;
  assign \new_[75061]_  = \new_[75060]_  & \new_[75057]_ ;
  assign \new_[75062]_  = \new_[75061]_  & \new_[75054]_ ;
  assign \new_[75066]_  = ~A168 & ~A169;
  assign \new_[75067]_  = ~A170 & \new_[75066]_ ;
  assign \new_[75070]_  = A166 & ~A167;
  assign \new_[75073]_  = ~A202 & A201;
  assign \new_[75074]_  = \new_[75073]_  & \new_[75070]_ ;
  assign \new_[75075]_  = \new_[75074]_  & \new_[75067]_ ;
  assign \new_[75079]_  = ~A266 & ~A265;
  assign \new_[75080]_  = A203 & \new_[75079]_ ;
  assign \new_[75083]_  = ~A299 & A298;
  assign \new_[75086]_  = ~A302 & A300;
  assign \new_[75087]_  = \new_[75086]_  & \new_[75083]_ ;
  assign \new_[75088]_  = \new_[75087]_  & \new_[75080]_ ;
  assign \new_[75092]_  = ~A168 & ~A169;
  assign \new_[75093]_  = ~A170 & \new_[75092]_ ;
  assign \new_[75096]_  = A166 & ~A167;
  assign \new_[75099]_  = ~A202 & A201;
  assign \new_[75100]_  = \new_[75099]_  & \new_[75096]_ ;
  assign \new_[75101]_  = \new_[75100]_  & \new_[75093]_ ;
  assign \new_[75105]_  = ~A266 & ~A265;
  assign \new_[75106]_  = A203 & \new_[75105]_ ;
  assign \new_[75109]_  = A299 & ~A298;
  assign \new_[75112]_  = A301 & A300;
  assign \new_[75113]_  = \new_[75112]_  & \new_[75109]_ ;
  assign \new_[75114]_  = \new_[75113]_  & \new_[75106]_ ;
  assign \new_[75118]_  = ~A168 & ~A169;
  assign \new_[75119]_  = ~A170 & \new_[75118]_ ;
  assign \new_[75122]_  = A166 & ~A167;
  assign \new_[75125]_  = ~A202 & A201;
  assign \new_[75126]_  = \new_[75125]_  & \new_[75122]_ ;
  assign \new_[75127]_  = \new_[75126]_  & \new_[75119]_ ;
  assign \new_[75131]_  = ~A266 & ~A265;
  assign \new_[75132]_  = A203 & \new_[75131]_ ;
  assign \new_[75135]_  = A299 & ~A298;
  assign \new_[75138]_  = ~A302 & A300;
  assign \new_[75139]_  = \new_[75138]_  & \new_[75135]_ ;
  assign \new_[75140]_  = \new_[75139]_  & \new_[75132]_ ;
  assign \new_[75144]_  = ~A168 & ~A169;
  assign \new_[75145]_  = ~A170 & \new_[75144]_ ;
  assign \new_[75148]_  = A166 & ~A167;
  assign \new_[75151]_  = A202 & ~A201;
  assign \new_[75152]_  = \new_[75151]_  & \new_[75148]_ ;
  assign \new_[75153]_  = \new_[75152]_  & \new_[75145]_ ;
  assign \new_[75157]_  = A269 & ~A268;
  assign \new_[75158]_  = A267 & \new_[75157]_ ;
  assign \new_[75161]_  = ~A299 & A298;
  assign \new_[75164]_  = A301 & A300;
  assign \new_[75165]_  = \new_[75164]_  & \new_[75161]_ ;
  assign \new_[75166]_  = \new_[75165]_  & \new_[75158]_ ;
  assign \new_[75170]_  = ~A168 & ~A169;
  assign \new_[75171]_  = ~A170 & \new_[75170]_ ;
  assign \new_[75174]_  = A166 & ~A167;
  assign \new_[75177]_  = A202 & ~A201;
  assign \new_[75178]_  = \new_[75177]_  & \new_[75174]_ ;
  assign \new_[75179]_  = \new_[75178]_  & \new_[75171]_ ;
  assign \new_[75183]_  = A269 & ~A268;
  assign \new_[75184]_  = A267 & \new_[75183]_ ;
  assign \new_[75187]_  = ~A299 & A298;
  assign \new_[75190]_  = ~A302 & A300;
  assign \new_[75191]_  = \new_[75190]_  & \new_[75187]_ ;
  assign \new_[75192]_  = \new_[75191]_  & \new_[75184]_ ;
  assign \new_[75196]_  = ~A168 & ~A169;
  assign \new_[75197]_  = ~A170 & \new_[75196]_ ;
  assign \new_[75200]_  = A166 & ~A167;
  assign \new_[75203]_  = A202 & ~A201;
  assign \new_[75204]_  = \new_[75203]_  & \new_[75200]_ ;
  assign \new_[75205]_  = \new_[75204]_  & \new_[75197]_ ;
  assign \new_[75209]_  = A269 & ~A268;
  assign \new_[75210]_  = A267 & \new_[75209]_ ;
  assign \new_[75213]_  = A299 & ~A298;
  assign \new_[75216]_  = A301 & A300;
  assign \new_[75217]_  = \new_[75216]_  & \new_[75213]_ ;
  assign \new_[75218]_  = \new_[75217]_  & \new_[75210]_ ;
  assign \new_[75222]_  = ~A168 & ~A169;
  assign \new_[75223]_  = ~A170 & \new_[75222]_ ;
  assign \new_[75226]_  = A166 & ~A167;
  assign \new_[75229]_  = A202 & ~A201;
  assign \new_[75230]_  = \new_[75229]_  & \new_[75226]_ ;
  assign \new_[75231]_  = \new_[75230]_  & \new_[75223]_ ;
  assign \new_[75235]_  = A269 & ~A268;
  assign \new_[75236]_  = A267 & \new_[75235]_ ;
  assign \new_[75239]_  = A299 & ~A298;
  assign \new_[75242]_  = ~A302 & A300;
  assign \new_[75243]_  = \new_[75242]_  & \new_[75239]_ ;
  assign \new_[75244]_  = \new_[75243]_  & \new_[75236]_ ;
  assign \new_[75248]_  = ~A168 & ~A169;
  assign \new_[75249]_  = ~A170 & \new_[75248]_ ;
  assign \new_[75252]_  = A166 & ~A167;
  assign \new_[75255]_  = A202 & ~A201;
  assign \new_[75256]_  = \new_[75255]_  & \new_[75252]_ ;
  assign \new_[75257]_  = \new_[75256]_  & \new_[75249]_ ;
  assign \new_[75261]_  = A298 & A268;
  assign \new_[75262]_  = ~A267 & \new_[75261]_ ;
  assign \new_[75265]_  = ~A300 & ~A299;
  assign \new_[75268]_  = A302 & ~A301;
  assign \new_[75269]_  = \new_[75268]_  & \new_[75265]_ ;
  assign \new_[75270]_  = \new_[75269]_  & \new_[75262]_ ;
  assign \new_[75274]_  = ~A168 & ~A169;
  assign \new_[75275]_  = ~A170 & \new_[75274]_ ;
  assign \new_[75278]_  = A166 & ~A167;
  assign \new_[75281]_  = A202 & ~A201;
  assign \new_[75282]_  = \new_[75281]_  & \new_[75278]_ ;
  assign \new_[75283]_  = \new_[75282]_  & \new_[75275]_ ;
  assign \new_[75287]_  = ~A298 & A268;
  assign \new_[75288]_  = ~A267 & \new_[75287]_ ;
  assign \new_[75291]_  = ~A300 & A299;
  assign \new_[75294]_  = A302 & ~A301;
  assign \new_[75295]_  = \new_[75294]_  & \new_[75291]_ ;
  assign \new_[75296]_  = \new_[75295]_  & \new_[75288]_ ;
  assign \new_[75300]_  = ~A168 & ~A169;
  assign \new_[75301]_  = ~A170 & \new_[75300]_ ;
  assign \new_[75304]_  = A166 & ~A167;
  assign \new_[75307]_  = A202 & ~A201;
  assign \new_[75308]_  = \new_[75307]_  & \new_[75304]_ ;
  assign \new_[75309]_  = \new_[75308]_  & \new_[75301]_ ;
  assign \new_[75313]_  = A298 & ~A269;
  assign \new_[75314]_  = ~A267 & \new_[75313]_ ;
  assign \new_[75317]_  = ~A300 & ~A299;
  assign \new_[75320]_  = A302 & ~A301;
  assign \new_[75321]_  = \new_[75320]_  & \new_[75317]_ ;
  assign \new_[75322]_  = \new_[75321]_  & \new_[75314]_ ;
  assign \new_[75326]_  = ~A168 & ~A169;
  assign \new_[75327]_  = ~A170 & \new_[75326]_ ;
  assign \new_[75330]_  = A166 & ~A167;
  assign \new_[75333]_  = A202 & ~A201;
  assign \new_[75334]_  = \new_[75333]_  & \new_[75330]_ ;
  assign \new_[75335]_  = \new_[75334]_  & \new_[75327]_ ;
  assign \new_[75339]_  = ~A298 & ~A269;
  assign \new_[75340]_  = ~A267 & \new_[75339]_ ;
  assign \new_[75343]_  = ~A300 & A299;
  assign \new_[75346]_  = A302 & ~A301;
  assign \new_[75347]_  = \new_[75346]_  & \new_[75343]_ ;
  assign \new_[75348]_  = \new_[75347]_  & \new_[75340]_ ;
  assign \new_[75352]_  = ~A168 & ~A169;
  assign \new_[75353]_  = ~A170 & \new_[75352]_ ;
  assign \new_[75356]_  = A166 & ~A167;
  assign \new_[75359]_  = A202 & ~A201;
  assign \new_[75360]_  = \new_[75359]_  & \new_[75356]_ ;
  assign \new_[75361]_  = \new_[75360]_  & \new_[75353]_ ;
  assign \new_[75365]_  = A298 & A266;
  assign \new_[75366]_  = A265 & \new_[75365]_ ;
  assign \new_[75369]_  = ~A300 & ~A299;
  assign \new_[75372]_  = A302 & ~A301;
  assign \new_[75373]_  = \new_[75372]_  & \new_[75369]_ ;
  assign \new_[75374]_  = \new_[75373]_  & \new_[75366]_ ;
  assign \new_[75378]_  = ~A168 & ~A169;
  assign \new_[75379]_  = ~A170 & \new_[75378]_ ;
  assign \new_[75382]_  = A166 & ~A167;
  assign \new_[75385]_  = A202 & ~A201;
  assign \new_[75386]_  = \new_[75385]_  & \new_[75382]_ ;
  assign \new_[75387]_  = \new_[75386]_  & \new_[75379]_ ;
  assign \new_[75391]_  = ~A298 & A266;
  assign \new_[75392]_  = A265 & \new_[75391]_ ;
  assign \new_[75395]_  = ~A300 & A299;
  assign \new_[75398]_  = A302 & ~A301;
  assign \new_[75399]_  = \new_[75398]_  & \new_[75395]_ ;
  assign \new_[75400]_  = \new_[75399]_  & \new_[75392]_ ;
  assign \new_[75404]_  = ~A168 & ~A169;
  assign \new_[75405]_  = ~A170 & \new_[75404]_ ;
  assign \new_[75408]_  = A166 & ~A167;
  assign \new_[75411]_  = A202 & ~A201;
  assign \new_[75412]_  = \new_[75411]_  & \new_[75408]_ ;
  assign \new_[75413]_  = \new_[75412]_  & \new_[75405]_ ;
  assign \new_[75417]_  = A267 & A266;
  assign \new_[75418]_  = ~A265 & \new_[75417]_ ;
  assign \new_[75421]_  = A300 & A268;
  assign \new_[75424]_  = A302 & ~A301;
  assign \new_[75425]_  = \new_[75424]_  & \new_[75421]_ ;
  assign \new_[75426]_  = \new_[75425]_  & \new_[75418]_ ;
  assign \new_[75430]_  = ~A168 & ~A169;
  assign \new_[75431]_  = ~A170 & \new_[75430]_ ;
  assign \new_[75434]_  = A166 & ~A167;
  assign \new_[75437]_  = A202 & ~A201;
  assign \new_[75438]_  = \new_[75437]_  & \new_[75434]_ ;
  assign \new_[75439]_  = \new_[75438]_  & \new_[75431]_ ;
  assign \new_[75443]_  = A267 & A266;
  assign \new_[75444]_  = ~A265 & \new_[75443]_ ;
  assign \new_[75447]_  = A300 & ~A269;
  assign \new_[75450]_  = A302 & ~A301;
  assign \new_[75451]_  = \new_[75450]_  & \new_[75447]_ ;
  assign \new_[75452]_  = \new_[75451]_  & \new_[75444]_ ;
  assign \new_[75456]_  = ~A168 & ~A169;
  assign \new_[75457]_  = ~A170 & \new_[75456]_ ;
  assign \new_[75460]_  = A166 & ~A167;
  assign \new_[75463]_  = A202 & ~A201;
  assign \new_[75464]_  = \new_[75463]_  & \new_[75460]_ ;
  assign \new_[75465]_  = \new_[75464]_  & \new_[75457]_ ;
  assign \new_[75469]_  = ~A267 & A266;
  assign \new_[75470]_  = ~A265 & \new_[75469]_ ;
  assign \new_[75473]_  = A269 & ~A268;
  assign \new_[75476]_  = A301 & ~A300;
  assign \new_[75477]_  = \new_[75476]_  & \new_[75473]_ ;
  assign \new_[75478]_  = \new_[75477]_  & \new_[75470]_ ;
  assign \new_[75482]_  = ~A168 & ~A169;
  assign \new_[75483]_  = ~A170 & \new_[75482]_ ;
  assign \new_[75486]_  = A166 & ~A167;
  assign \new_[75489]_  = A202 & ~A201;
  assign \new_[75490]_  = \new_[75489]_  & \new_[75486]_ ;
  assign \new_[75491]_  = \new_[75490]_  & \new_[75483]_ ;
  assign \new_[75495]_  = ~A267 & A266;
  assign \new_[75496]_  = ~A265 & \new_[75495]_ ;
  assign \new_[75499]_  = A269 & ~A268;
  assign \new_[75502]_  = ~A302 & ~A300;
  assign \new_[75503]_  = \new_[75502]_  & \new_[75499]_ ;
  assign \new_[75504]_  = \new_[75503]_  & \new_[75496]_ ;
  assign \new_[75508]_  = ~A168 & ~A169;
  assign \new_[75509]_  = ~A170 & \new_[75508]_ ;
  assign \new_[75512]_  = A166 & ~A167;
  assign \new_[75515]_  = A202 & ~A201;
  assign \new_[75516]_  = \new_[75515]_  & \new_[75512]_ ;
  assign \new_[75517]_  = \new_[75516]_  & \new_[75509]_ ;
  assign \new_[75521]_  = ~A267 & A266;
  assign \new_[75522]_  = ~A265 & \new_[75521]_ ;
  assign \new_[75525]_  = A269 & ~A268;
  assign \new_[75528]_  = A299 & A298;
  assign \new_[75529]_  = \new_[75528]_  & \new_[75525]_ ;
  assign \new_[75530]_  = \new_[75529]_  & \new_[75522]_ ;
  assign \new_[75534]_  = ~A168 & ~A169;
  assign \new_[75535]_  = ~A170 & \new_[75534]_ ;
  assign \new_[75538]_  = A166 & ~A167;
  assign \new_[75541]_  = A202 & ~A201;
  assign \new_[75542]_  = \new_[75541]_  & \new_[75538]_ ;
  assign \new_[75543]_  = \new_[75542]_  & \new_[75535]_ ;
  assign \new_[75547]_  = ~A267 & A266;
  assign \new_[75548]_  = ~A265 & \new_[75547]_ ;
  assign \new_[75551]_  = A269 & ~A268;
  assign \new_[75554]_  = ~A299 & ~A298;
  assign \new_[75555]_  = \new_[75554]_  & \new_[75551]_ ;
  assign \new_[75556]_  = \new_[75555]_  & \new_[75548]_ ;
  assign \new_[75560]_  = ~A168 & ~A169;
  assign \new_[75561]_  = ~A170 & \new_[75560]_ ;
  assign \new_[75564]_  = A166 & ~A167;
  assign \new_[75567]_  = A202 & ~A201;
  assign \new_[75568]_  = \new_[75567]_  & \new_[75564]_ ;
  assign \new_[75569]_  = \new_[75568]_  & \new_[75561]_ ;
  assign \new_[75573]_  = A267 & ~A266;
  assign \new_[75574]_  = A265 & \new_[75573]_ ;
  assign \new_[75577]_  = A300 & A268;
  assign \new_[75580]_  = A302 & ~A301;
  assign \new_[75581]_  = \new_[75580]_  & \new_[75577]_ ;
  assign \new_[75582]_  = \new_[75581]_  & \new_[75574]_ ;
  assign \new_[75586]_  = ~A168 & ~A169;
  assign \new_[75587]_  = ~A170 & \new_[75586]_ ;
  assign \new_[75590]_  = A166 & ~A167;
  assign \new_[75593]_  = A202 & ~A201;
  assign \new_[75594]_  = \new_[75593]_  & \new_[75590]_ ;
  assign \new_[75595]_  = \new_[75594]_  & \new_[75587]_ ;
  assign \new_[75599]_  = A267 & ~A266;
  assign \new_[75600]_  = A265 & \new_[75599]_ ;
  assign \new_[75603]_  = A300 & ~A269;
  assign \new_[75606]_  = A302 & ~A301;
  assign \new_[75607]_  = \new_[75606]_  & \new_[75603]_ ;
  assign \new_[75608]_  = \new_[75607]_  & \new_[75600]_ ;
  assign \new_[75612]_  = ~A168 & ~A169;
  assign \new_[75613]_  = ~A170 & \new_[75612]_ ;
  assign \new_[75616]_  = A166 & ~A167;
  assign \new_[75619]_  = A202 & ~A201;
  assign \new_[75620]_  = \new_[75619]_  & \new_[75616]_ ;
  assign \new_[75621]_  = \new_[75620]_  & \new_[75613]_ ;
  assign \new_[75625]_  = ~A267 & ~A266;
  assign \new_[75626]_  = A265 & \new_[75625]_ ;
  assign \new_[75629]_  = A269 & ~A268;
  assign \new_[75632]_  = A301 & ~A300;
  assign \new_[75633]_  = \new_[75632]_  & \new_[75629]_ ;
  assign \new_[75634]_  = \new_[75633]_  & \new_[75626]_ ;
  assign \new_[75638]_  = ~A168 & ~A169;
  assign \new_[75639]_  = ~A170 & \new_[75638]_ ;
  assign \new_[75642]_  = A166 & ~A167;
  assign \new_[75645]_  = A202 & ~A201;
  assign \new_[75646]_  = \new_[75645]_  & \new_[75642]_ ;
  assign \new_[75647]_  = \new_[75646]_  & \new_[75639]_ ;
  assign \new_[75651]_  = ~A267 & ~A266;
  assign \new_[75652]_  = A265 & \new_[75651]_ ;
  assign \new_[75655]_  = A269 & ~A268;
  assign \new_[75658]_  = ~A302 & ~A300;
  assign \new_[75659]_  = \new_[75658]_  & \new_[75655]_ ;
  assign \new_[75660]_  = \new_[75659]_  & \new_[75652]_ ;
  assign \new_[75664]_  = ~A168 & ~A169;
  assign \new_[75665]_  = ~A170 & \new_[75664]_ ;
  assign \new_[75668]_  = A166 & ~A167;
  assign \new_[75671]_  = A202 & ~A201;
  assign \new_[75672]_  = \new_[75671]_  & \new_[75668]_ ;
  assign \new_[75673]_  = \new_[75672]_  & \new_[75665]_ ;
  assign \new_[75677]_  = ~A267 & ~A266;
  assign \new_[75678]_  = A265 & \new_[75677]_ ;
  assign \new_[75681]_  = A269 & ~A268;
  assign \new_[75684]_  = A299 & A298;
  assign \new_[75685]_  = \new_[75684]_  & \new_[75681]_ ;
  assign \new_[75686]_  = \new_[75685]_  & \new_[75678]_ ;
  assign \new_[75690]_  = ~A168 & ~A169;
  assign \new_[75691]_  = ~A170 & \new_[75690]_ ;
  assign \new_[75694]_  = A166 & ~A167;
  assign \new_[75697]_  = A202 & ~A201;
  assign \new_[75698]_  = \new_[75697]_  & \new_[75694]_ ;
  assign \new_[75699]_  = \new_[75698]_  & \new_[75691]_ ;
  assign \new_[75703]_  = ~A267 & ~A266;
  assign \new_[75704]_  = A265 & \new_[75703]_ ;
  assign \new_[75707]_  = A269 & ~A268;
  assign \new_[75710]_  = ~A299 & ~A298;
  assign \new_[75711]_  = \new_[75710]_  & \new_[75707]_ ;
  assign \new_[75712]_  = \new_[75711]_  & \new_[75704]_ ;
  assign \new_[75716]_  = ~A168 & ~A169;
  assign \new_[75717]_  = ~A170 & \new_[75716]_ ;
  assign \new_[75720]_  = A166 & ~A167;
  assign \new_[75723]_  = A202 & ~A201;
  assign \new_[75724]_  = \new_[75723]_  & \new_[75720]_ ;
  assign \new_[75725]_  = \new_[75724]_  & \new_[75717]_ ;
  assign \new_[75729]_  = A298 & ~A266;
  assign \new_[75730]_  = ~A265 & \new_[75729]_ ;
  assign \new_[75733]_  = ~A300 & ~A299;
  assign \new_[75736]_  = A302 & ~A301;
  assign \new_[75737]_  = \new_[75736]_  & \new_[75733]_ ;
  assign \new_[75738]_  = \new_[75737]_  & \new_[75730]_ ;
  assign \new_[75742]_  = ~A168 & ~A169;
  assign \new_[75743]_  = ~A170 & \new_[75742]_ ;
  assign \new_[75746]_  = A166 & ~A167;
  assign \new_[75749]_  = A202 & ~A201;
  assign \new_[75750]_  = \new_[75749]_  & \new_[75746]_ ;
  assign \new_[75751]_  = \new_[75750]_  & \new_[75743]_ ;
  assign \new_[75755]_  = ~A298 & ~A266;
  assign \new_[75756]_  = ~A265 & \new_[75755]_ ;
  assign \new_[75759]_  = ~A300 & A299;
  assign \new_[75762]_  = A302 & ~A301;
  assign \new_[75763]_  = \new_[75762]_  & \new_[75759]_ ;
  assign \new_[75764]_  = \new_[75763]_  & \new_[75756]_ ;
  assign \new_[75768]_  = ~A168 & ~A169;
  assign \new_[75769]_  = ~A170 & \new_[75768]_ ;
  assign \new_[75772]_  = A166 & ~A167;
  assign \new_[75775]_  = ~A203 & ~A201;
  assign \new_[75776]_  = \new_[75775]_  & \new_[75772]_ ;
  assign \new_[75777]_  = \new_[75776]_  & \new_[75769]_ ;
  assign \new_[75781]_  = A269 & ~A268;
  assign \new_[75782]_  = A267 & \new_[75781]_ ;
  assign \new_[75785]_  = ~A299 & A298;
  assign \new_[75788]_  = A301 & A300;
  assign \new_[75789]_  = \new_[75788]_  & \new_[75785]_ ;
  assign \new_[75790]_  = \new_[75789]_  & \new_[75782]_ ;
  assign \new_[75794]_  = ~A168 & ~A169;
  assign \new_[75795]_  = ~A170 & \new_[75794]_ ;
  assign \new_[75798]_  = A166 & ~A167;
  assign \new_[75801]_  = ~A203 & ~A201;
  assign \new_[75802]_  = \new_[75801]_  & \new_[75798]_ ;
  assign \new_[75803]_  = \new_[75802]_  & \new_[75795]_ ;
  assign \new_[75807]_  = A269 & ~A268;
  assign \new_[75808]_  = A267 & \new_[75807]_ ;
  assign \new_[75811]_  = ~A299 & A298;
  assign \new_[75814]_  = ~A302 & A300;
  assign \new_[75815]_  = \new_[75814]_  & \new_[75811]_ ;
  assign \new_[75816]_  = \new_[75815]_  & \new_[75808]_ ;
  assign \new_[75820]_  = ~A168 & ~A169;
  assign \new_[75821]_  = ~A170 & \new_[75820]_ ;
  assign \new_[75824]_  = A166 & ~A167;
  assign \new_[75827]_  = ~A203 & ~A201;
  assign \new_[75828]_  = \new_[75827]_  & \new_[75824]_ ;
  assign \new_[75829]_  = \new_[75828]_  & \new_[75821]_ ;
  assign \new_[75833]_  = A269 & ~A268;
  assign \new_[75834]_  = A267 & \new_[75833]_ ;
  assign \new_[75837]_  = A299 & ~A298;
  assign \new_[75840]_  = A301 & A300;
  assign \new_[75841]_  = \new_[75840]_  & \new_[75837]_ ;
  assign \new_[75842]_  = \new_[75841]_  & \new_[75834]_ ;
  assign \new_[75846]_  = ~A168 & ~A169;
  assign \new_[75847]_  = ~A170 & \new_[75846]_ ;
  assign \new_[75850]_  = A166 & ~A167;
  assign \new_[75853]_  = ~A203 & ~A201;
  assign \new_[75854]_  = \new_[75853]_  & \new_[75850]_ ;
  assign \new_[75855]_  = \new_[75854]_  & \new_[75847]_ ;
  assign \new_[75859]_  = A269 & ~A268;
  assign \new_[75860]_  = A267 & \new_[75859]_ ;
  assign \new_[75863]_  = A299 & ~A298;
  assign \new_[75866]_  = ~A302 & A300;
  assign \new_[75867]_  = \new_[75866]_  & \new_[75863]_ ;
  assign \new_[75868]_  = \new_[75867]_  & \new_[75860]_ ;
  assign \new_[75872]_  = ~A168 & ~A169;
  assign \new_[75873]_  = ~A170 & \new_[75872]_ ;
  assign \new_[75876]_  = A166 & ~A167;
  assign \new_[75879]_  = ~A203 & ~A201;
  assign \new_[75880]_  = \new_[75879]_  & \new_[75876]_ ;
  assign \new_[75881]_  = \new_[75880]_  & \new_[75873]_ ;
  assign \new_[75885]_  = A298 & A268;
  assign \new_[75886]_  = ~A267 & \new_[75885]_ ;
  assign \new_[75889]_  = ~A300 & ~A299;
  assign \new_[75892]_  = A302 & ~A301;
  assign \new_[75893]_  = \new_[75892]_  & \new_[75889]_ ;
  assign \new_[75894]_  = \new_[75893]_  & \new_[75886]_ ;
  assign \new_[75898]_  = ~A168 & ~A169;
  assign \new_[75899]_  = ~A170 & \new_[75898]_ ;
  assign \new_[75902]_  = A166 & ~A167;
  assign \new_[75905]_  = ~A203 & ~A201;
  assign \new_[75906]_  = \new_[75905]_  & \new_[75902]_ ;
  assign \new_[75907]_  = \new_[75906]_  & \new_[75899]_ ;
  assign \new_[75911]_  = ~A298 & A268;
  assign \new_[75912]_  = ~A267 & \new_[75911]_ ;
  assign \new_[75915]_  = ~A300 & A299;
  assign \new_[75918]_  = A302 & ~A301;
  assign \new_[75919]_  = \new_[75918]_  & \new_[75915]_ ;
  assign \new_[75920]_  = \new_[75919]_  & \new_[75912]_ ;
  assign \new_[75924]_  = ~A168 & ~A169;
  assign \new_[75925]_  = ~A170 & \new_[75924]_ ;
  assign \new_[75928]_  = A166 & ~A167;
  assign \new_[75931]_  = ~A203 & ~A201;
  assign \new_[75932]_  = \new_[75931]_  & \new_[75928]_ ;
  assign \new_[75933]_  = \new_[75932]_  & \new_[75925]_ ;
  assign \new_[75937]_  = A298 & ~A269;
  assign \new_[75938]_  = ~A267 & \new_[75937]_ ;
  assign \new_[75941]_  = ~A300 & ~A299;
  assign \new_[75944]_  = A302 & ~A301;
  assign \new_[75945]_  = \new_[75944]_  & \new_[75941]_ ;
  assign \new_[75946]_  = \new_[75945]_  & \new_[75938]_ ;
  assign \new_[75950]_  = ~A168 & ~A169;
  assign \new_[75951]_  = ~A170 & \new_[75950]_ ;
  assign \new_[75954]_  = A166 & ~A167;
  assign \new_[75957]_  = ~A203 & ~A201;
  assign \new_[75958]_  = \new_[75957]_  & \new_[75954]_ ;
  assign \new_[75959]_  = \new_[75958]_  & \new_[75951]_ ;
  assign \new_[75963]_  = ~A298 & ~A269;
  assign \new_[75964]_  = ~A267 & \new_[75963]_ ;
  assign \new_[75967]_  = ~A300 & A299;
  assign \new_[75970]_  = A302 & ~A301;
  assign \new_[75971]_  = \new_[75970]_  & \new_[75967]_ ;
  assign \new_[75972]_  = \new_[75971]_  & \new_[75964]_ ;
  assign \new_[75976]_  = ~A168 & ~A169;
  assign \new_[75977]_  = ~A170 & \new_[75976]_ ;
  assign \new_[75980]_  = A166 & ~A167;
  assign \new_[75983]_  = ~A203 & ~A201;
  assign \new_[75984]_  = \new_[75983]_  & \new_[75980]_ ;
  assign \new_[75985]_  = \new_[75984]_  & \new_[75977]_ ;
  assign \new_[75989]_  = A298 & A266;
  assign \new_[75990]_  = A265 & \new_[75989]_ ;
  assign \new_[75993]_  = ~A300 & ~A299;
  assign \new_[75996]_  = A302 & ~A301;
  assign \new_[75997]_  = \new_[75996]_  & \new_[75993]_ ;
  assign \new_[75998]_  = \new_[75997]_  & \new_[75990]_ ;
  assign \new_[76002]_  = ~A168 & ~A169;
  assign \new_[76003]_  = ~A170 & \new_[76002]_ ;
  assign \new_[76006]_  = A166 & ~A167;
  assign \new_[76009]_  = ~A203 & ~A201;
  assign \new_[76010]_  = \new_[76009]_  & \new_[76006]_ ;
  assign \new_[76011]_  = \new_[76010]_  & \new_[76003]_ ;
  assign \new_[76015]_  = ~A298 & A266;
  assign \new_[76016]_  = A265 & \new_[76015]_ ;
  assign \new_[76019]_  = ~A300 & A299;
  assign \new_[76022]_  = A302 & ~A301;
  assign \new_[76023]_  = \new_[76022]_  & \new_[76019]_ ;
  assign \new_[76024]_  = \new_[76023]_  & \new_[76016]_ ;
  assign \new_[76028]_  = ~A168 & ~A169;
  assign \new_[76029]_  = ~A170 & \new_[76028]_ ;
  assign \new_[76032]_  = A166 & ~A167;
  assign \new_[76035]_  = ~A203 & ~A201;
  assign \new_[76036]_  = \new_[76035]_  & \new_[76032]_ ;
  assign \new_[76037]_  = \new_[76036]_  & \new_[76029]_ ;
  assign \new_[76041]_  = A267 & A266;
  assign \new_[76042]_  = ~A265 & \new_[76041]_ ;
  assign \new_[76045]_  = A300 & A268;
  assign \new_[76048]_  = A302 & ~A301;
  assign \new_[76049]_  = \new_[76048]_  & \new_[76045]_ ;
  assign \new_[76050]_  = \new_[76049]_  & \new_[76042]_ ;
  assign \new_[76054]_  = ~A168 & ~A169;
  assign \new_[76055]_  = ~A170 & \new_[76054]_ ;
  assign \new_[76058]_  = A166 & ~A167;
  assign \new_[76061]_  = ~A203 & ~A201;
  assign \new_[76062]_  = \new_[76061]_  & \new_[76058]_ ;
  assign \new_[76063]_  = \new_[76062]_  & \new_[76055]_ ;
  assign \new_[76067]_  = A267 & A266;
  assign \new_[76068]_  = ~A265 & \new_[76067]_ ;
  assign \new_[76071]_  = A300 & ~A269;
  assign \new_[76074]_  = A302 & ~A301;
  assign \new_[76075]_  = \new_[76074]_  & \new_[76071]_ ;
  assign \new_[76076]_  = \new_[76075]_  & \new_[76068]_ ;
  assign \new_[76080]_  = ~A168 & ~A169;
  assign \new_[76081]_  = ~A170 & \new_[76080]_ ;
  assign \new_[76084]_  = A166 & ~A167;
  assign \new_[76087]_  = ~A203 & ~A201;
  assign \new_[76088]_  = \new_[76087]_  & \new_[76084]_ ;
  assign \new_[76089]_  = \new_[76088]_  & \new_[76081]_ ;
  assign \new_[76093]_  = ~A267 & A266;
  assign \new_[76094]_  = ~A265 & \new_[76093]_ ;
  assign \new_[76097]_  = A269 & ~A268;
  assign \new_[76100]_  = A301 & ~A300;
  assign \new_[76101]_  = \new_[76100]_  & \new_[76097]_ ;
  assign \new_[76102]_  = \new_[76101]_  & \new_[76094]_ ;
  assign \new_[76106]_  = ~A168 & ~A169;
  assign \new_[76107]_  = ~A170 & \new_[76106]_ ;
  assign \new_[76110]_  = A166 & ~A167;
  assign \new_[76113]_  = ~A203 & ~A201;
  assign \new_[76114]_  = \new_[76113]_  & \new_[76110]_ ;
  assign \new_[76115]_  = \new_[76114]_  & \new_[76107]_ ;
  assign \new_[76119]_  = ~A267 & A266;
  assign \new_[76120]_  = ~A265 & \new_[76119]_ ;
  assign \new_[76123]_  = A269 & ~A268;
  assign \new_[76126]_  = ~A302 & ~A300;
  assign \new_[76127]_  = \new_[76126]_  & \new_[76123]_ ;
  assign \new_[76128]_  = \new_[76127]_  & \new_[76120]_ ;
  assign \new_[76132]_  = ~A168 & ~A169;
  assign \new_[76133]_  = ~A170 & \new_[76132]_ ;
  assign \new_[76136]_  = A166 & ~A167;
  assign \new_[76139]_  = ~A203 & ~A201;
  assign \new_[76140]_  = \new_[76139]_  & \new_[76136]_ ;
  assign \new_[76141]_  = \new_[76140]_  & \new_[76133]_ ;
  assign \new_[76145]_  = ~A267 & A266;
  assign \new_[76146]_  = ~A265 & \new_[76145]_ ;
  assign \new_[76149]_  = A269 & ~A268;
  assign \new_[76152]_  = A299 & A298;
  assign \new_[76153]_  = \new_[76152]_  & \new_[76149]_ ;
  assign \new_[76154]_  = \new_[76153]_  & \new_[76146]_ ;
  assign \new_[76158]_  = ~A168 & ~A169;
  assign \new_[76159]_  = ~A170 & \new_[76158]_ ;
  assign \new_[76162]_  = A166 & ~A167;
  assign \new_[76165]_  = ~A203 & ~A201;
  assign \new_[76166]_  = \new_[76165]_  & \new_[76162]_ ;
  assign \new_[76167]_  = \new_[76166]_  & \new_[76159]_ ;
  assign \new_[76171]_  = ~A267 & A266;
  assign \new_[76172]_  = ~A265 & \new_[76171]_ ;
  assign \new_[76175]_  = A269 & ~A268;
  assign \new_[76178]_  = ~A299 & ~A298;
  assign \new_[76179]_  = \new_[76178]_  & \new_[76175]_ ;
  assign \new_[76180]_  = \new_[76179]_  & \new_[76172]_ ;
  assign \new_[76184]_  = ~A168 & ~A169;
  assign \new_[76185]_  = ~A170 & \new_[76184]_ ;
  assign \new_[76188]_  = A166 & ~A167;
  assign \new_[76191]_  = ~A203 & ~A201;
  assign \new_[76192]_  = \new_[76191]_  & \new_[76188]_ ;
  assign \new_[76193]_  = \new_[76192]_  & \new_[76185]_ ;
  assign \new_[76197]_  = A267 & ~A266;
  assign \new_[76198]_  = A265 & \new_[76197]_ ;
  assign \new_[76201]_  = A300 & A268;
  assign \new_[76204]_  = A302 & ~A301;
  assign \new_[76205]_  = \new_[76204]_  & \new_[76201]_ ;
  assign \new_[76206]_  = \new_[76205]_  & \new_[76198]_ ;
  assign \new_[76210]_  = ~A168 & ~A169;
  assign \new_[76211]_  = ~A170 & \new_[76210]_ ;
  assign \new_[76214]_  = A166 & ~A167;
  assign \new_[76217]_  = ~A203 & ~A201;
  assign \new_[76218]_  = \new_[76217]_  & \new_[76214]_ ;
  assign \new_[76219]_  = \new_[76218]_  & \new_[76211]_ ;
  assign \new_[76223]_  = A267 & ~A266;
  assign \new_[76224]_  = A265 & \new_[76223]_ ;
  assign \new_[76227]_  = A300 & ~A269;
  assign \new_[76230]_  = A302 & ~A301;
  assign \new_[76231]_  = \new_[76230]_  & \new_[76227]_ ;
  assign \new_[76232]_  = \new_[76231]_  & \new_[76224]_ ;
  assign \new_[76236]_  = ~A168 & ~A169;
  assign \new_[76237]_  = ~A170 & \new_[76236]_ ;
  assign \new_[76240]_  = A166 & ~A167;
  assign \new_[76243]_  = ~A203 & ~A201;
  assign \new_[76244]_  = \new_[76243]_  & \new_[76240]_ ;
  assign \new_[76245]_  = \new_[76244]_  & \new_[76237]_ ;
  assign \new_[76249]_  = ~A267 & ~A266;
  assign \new_[76250]_  = A265 & \new_[76249]_ ;
  assign \new_[76253]_  = A269 & ~A268;
  assign \new_[76256]_  = A301 & ~A300;
  assign \new_[76257]_  = \new_[76256]_  & \new_[76253]_ ;
  assign \new_[76258]_  = \new_[76257]_  & \new_[76250]_ ;
  assign \new_[76262]_  = ~A168 & ~A169;
  assign \new_[76263]_  = ~A170 & \new_[76262]_ ;
  assign \new_[76266]_  = A166 & ~A167;
  assign \new_[76269]_  = ~A203 & ~A201;
  assign \new_[76270]_  = \new_[76269]_  & \new_[76266]_ ;
  assign \new_[76271]_  = \new_[76270]_  & \new_[76263]_ ;
  assign \new_[76275]_  = ~A267 & ~A266;
  assign \new_[76276]_  = A265 & \new_[76275]_ ;
  assign \new_[76279]_  = A269 & ~A268;
  assign \new_[76282]_  = ~A302 & ~A300;
  assign \new_[76283]_  = \new_[76282]_  & \new_[76279]_ ;
  assign \new_[76284]_  = \new_[76283]_  & \new_[76276]_ ;
  assign \new_[76288]_  = ~A168 & ~A169;
  assign \new_[76289]_  = ~A170 & \new_[76288]_ ;
  assign \new_[76292]_  = A166 & ~A167;
  assign \new_[76295]_  = ~A203 & ~A201;
  assign \new_[76296]_  = \new_[76295]_  & \new_[76292]_ ;
  assign \new_[76297]_  = \new_[76296]_  & \new_[76289]_ ;
  assign \new_[76301]_  = ~A267 & ~A266;
  assign \new_[76302]_  = A265 & \new_[76301]_ ;
  assign \new_[76305]_  = A269 & ~A268;
  assign \new_[76308]_  = A299 & A298;
  assign \new_[76309]_  = \new_[76308]_  & \new_[76305]_ ;
  assign \new_[76310]_  = \new_[76309]_  & \new_[76302]_ ;
  assign \new_[76314]_  = ~A168 & ~A169;
  assign \new_[76315]_  = ~A170 & \new_[76314]_ ;
  assign \new_[76318]_  = A166 & ~A167;
  assign \new_[76321]_  = ~A203 & ~A201;
  assign \new_[76322]_  = \new_[76321]_  & \new_[76318]_ ;
  assign \new_[76323]_  = \new_[76322]_  & \new_[76315]_ ;
  assign \new_[76327]_  = ~A267 & ~A266;
  assign \new_[76328]_  = A265 & \new_[76327]_ ;
  assign \new_[76331]_  = A269 & ~A268;
  assign \new_[76334]_  = ~A299 & ~A298;
  assign \new_[76335]_  = \new_[76334]_  & \new_[76331]_ ;
  assign \new_[76336]_  = \new_[76335]_  & \new_[76328]_ ;
  assign \new_[76340]_  = ~A168 & ~A169;
  assign \new_[76341]_  = ~A170 & \new_[76340]_ ;
  assign \new_[76344]_  = A166 & ~A167;
  assign \new_[76347]_  = ~A203 & ~A201;
  assign \new_[76348]_  = \new_[76347]_  & \new_[76344]_ ;
  assign \new_[76349]_  = \new_[76348]_  & \new_[76341]_ ;
  assign \new_[76353]_  = A298 & ~A266;
  assign \new_[76354]_  = ~A265 & \new_[76353]_ ;
  assign \new_[76357]_  = ~A300 & ~A299;
  assign \new_[76360]_  = A302 & ~A301;
  assign \new_[76361]_  = \new_[76360]_  & \new_[76357]_ ;
  assign \new_[76362]_  = \new_[76361]_  & \new_[76354]_ ;
  assign \new_[76366]_  = ~A168 & ~A169;
  assign \new_[76367]_  = ~A170 & \new_[76366]_ ;
  assign \new_[76370]_  = A166 & ~A167;
  assign \new_[76373]_  = ~A203 & ~A201;
  assign \new_[76374]_  = \new_[76373]_  & \new_[76370]_ ;
  assign \new_[76375]_  = \new_[76374]_  & \new_[76367]_ ;
  assign \new_[76379]_  = ~A298 & ~A266;
  assign \new_[76380]_  = ~A265 & \new_[76379]_ ;
  assign \new_[76383]_  = ~A300 & A299;
  assign \new_[76386]_  = A302 & ~A301;
  assign \new_[76387]_  = \new_[76386]_  & \new_[76383]_ ;
  assign \new_[76388]_  = \new_[76387]_  & \new_[76380]_ ;
  assign \new_[76392]_  = ~A168 & ~A169;
  assign \new_[76393]_  = ~A170 & \new_[76392]_ ;
  assign \new_[76396]_  = A166 & ~A167;
  assign \new_[76399]_  = A200 & A199;
  assign \new_[76400]_  = \new_[76399]_  & \new_[76396]_ ;
  assign \new_[76401]_  = \new_[76400]_  & \new_[76393]_ ;
  assign \new_[76405]_  = A269 & ~A268;
  assign \new_[76406]_  = A267 & \new_[76405]_ ;
  assign \new_[76409]_  = ~A299 & A298;
  assign \new_[76412]_  = A301 & A300;
  assign \new_[76413]_  = \new_[76412]_  & \new_[76409]_ ;
  assign \new_[76414]_  = \new_[76413]_  & \new_[76406]_ ;
  assign \new_[76418]_  = ~A168 & ~A169;
  assign \new_[76419]_  = ~A170 & \new_[76418]_ ;
  assign \new_[76422]_  = A166 & ~A167;
  assign \new_[76425]_  = A200 & A199;
  assign \new_[76426]_  = \new_[76425]_  & \new_[76422]_ ;
  assign \new_[76427]_  = \new_[76426]_  & \new_[76419]_ ;
  assign \new_[76431]_  = A269 & ~A268;
  assign \new_[76432]_  = A267 & \new_[76431]_ ;
  assign \new_[76435]_  = ~A299 & A298;
  assign \new_[76438]_  = ~A302 & A300;
  assign \new_[76439]_  = \new_[76438]_  & \new_[76435]_ ;
  assign \new_[76440]_  = \new_[76439]_  & \new_[76432]_ ;
  assign \new_[76444]_  = ~A168 & ~A169;
  assign \new_[76445]_  = ~A170 & \new_[76444]_ ;
  assign \new_[76448]_  = A166 & ~A167;
  assign \new_[76451]_  = A200 & A199;
  assign \new_[76452]_  = \new_[76451]_  & \new_[76448]_ ;
  assign \new_[76453]_  = \new_[76452]_  & \new_[76445]_ ;
  assign \new_[76457]_  = A269 & ~A268;
  assign \new_[76458]_  = A267 & \new_[76457]_ ;
  assign \new_[76461]_  = A299 & ~A298;
  assign \new_[76464]_  = A301 & A300;
  assign \new_[76465]_  = \new_[76464]_  & \new_[76461]_ ;
  assign \new_[76466]_  = \new_[76465]_  & \new_[76458]_ ;
  assign \new_[76470]_  = ~A168 & ~A169;
  assign \new_[76471]_  = ~A170 & \new_[76470]_ ;
  assign \new_[76474]_  = A166 & ~A167;
  assign \new_[76477]_  = A200 & A199;
  assign \new_[76478]_  = \new_[76477]_  & \new_[76474]_ ;
  assign \new_[76479]_  = \new_[76478]_  & \new_[76471]_ ;
  assign \new_[76483]_  = A269 & ~A268;
  assign \new_[76484]_  = A267 & \new_[76483]_ ;
  assign \new_[76487]_  = A299 & ~A298;
  assign \new_[76490]_  = ~A302 & A300;
  assign \new_[76491]_  = \new_[76490]_  & \new_[76487]_ ;
  assign \new_[76492]_  = \new_[76491]_  & \new_[76484]_ ;
  assign \new_[76496]_  = ~A168 & ~A169;
  assign \new_[76497]_  = ~A170 & \new_[76496]_ ;
  assign \new_[76500]_  = A166 & ~A167;
  assign \new_[76503]_  = A200 & A199;
  assign \new_[76504]_  = \new_[76503]_  & \new_[76500]_ ;
  assign \new_[76505]_  = \new_[76504]_  & \new_[76497]_ ;
  assign \new_[76509]_  = A298 & A268;
  assign \new_[76510]_  = ~A267 & \new_[76509]_ ;
  assign \new_[76513]_  = ~A300 & ~A299;
  assign \new_[76516]_  = A302 & ~A301;
  assign \new_[76517]_  = \new_[76516]_  & \new_[76513]_ ;
  assign \new_[76518]_  = \new_[76517]_  & \new_[76510]_ ;
  assign \new_[76522]_  = ~A168 & ~A169;
  assign \new_[76523]_  = ~A170 & \new_[76522]_ ;
  assign \new_[76526]_  = A166 & ~A167;
  assign \new_[76529]_  = A200 & A199;
  assign \new_[76530]_  = \new_[76529]_  & \new_[76526]_ ;
  assign \new_[76531]_  = \new_[76530]_  & \new_[76523]_ ;
  assign \new_[76535]_  = ~A298 & A268;
  assign \new_[76536]_  = ~A267 & \new_[76535]_ ;
  assign \new_[76539]_  = ~A300 & A299;
  assign \new_[76542]_  = A302 & ~A301;
  assign \new_[76543]_  = \new_[76542]_  & \new_[76539]_ ;
  assign \new_[76544]_  = \new_[76543]_  & \new_[76536]_ ;
  assign \new_[76548]_  = ~A168 & ~A169;
  assign \new_[76549]_  = ~A170 & \new_[76548]_ ;
  assign \new_[76552]_  = A166 & ~A167;
  assign \new_[76555]_  = A200 & A199;
  assign \new_[76556]_  = \new_[76555]_  & \new_[76552]_ ;
  assign \new_[76557]_  = \new_[76556]_  & \new_[76549]_ ;
  assign \new_[76561]_  = A298 & ~A269;
  assign \new_[76562]_  = ~A267 & \new_[76561]_ ;
  assign \new_[76565]_  = ~A300 & ~A299;
  assign \new_[76568]_  = A302 & ~A301;
  assign \new_[76569]_  = \new_[76568]_  & \new_[76565]_ ;
  assign \new_[76570]_  = \new_[76569]_  & \new_[76562]_ ;
  assign \new_[76574]_  = ~A168 & ~A169;
  assign \new_[76575]_  = ~A170 & \new_[76574]_ ;
  assign \new_[76578]_  = A166 & ~A167;
  assign \new_[76581]_  = A200 & A199;
  assign \new_[76582]_  = \new_[76581]_  & \new_[76578]_ ;
  assign \new_[76583]_  = \new_[76582]_  & \new_[76575]_ ;
  assign \new_[76587]_  = ~A298 & ~A269;
  assign \new_[76588]_  = ~A267 & \new_[76587]_ ;
  assign \new_[76591]_  = ~A300 & A299;
  assign \new_[76594]_  = A302 & ~A301;
  assign \new_[76595]_  = \new_[76594]_  & \new_[76591]_ ;
  assign \new_[76596]_  = \new_[76595]_  & \new_[76588]_ ;
  assign \new_[76600]_  = ~A168 & ~A169;
  assign \new_[76601]_  = ~A170 & \new_[76600]_ ;
  assign \new_[76604]_  = A166 & ~A167;
  assign \new_[76607]_  = A200 & A199;
  assign \new_[76608]_  = \new_[76607]_  & \new_[76604]_ ;
  assign \new_[76609]_  = \new_[76608]_  & \new_[76601]_ ;
  assign \new_[76613]_  = A298 & A266;
  assign \new_[76614]_  = A265 & \new_[76613]_ ;
  assign \new_[76617]_  = ~A300 & ~A299;
  assign \new_[76620]_  = A302 & ~A301;
  assign \new_[76621]_  = \new_[76620]_  & \new_[76617]_ ;
  assign \new_[76622]_  = \new_[76621]_  & \new_[76614]_ ;
  assign \new_[76626]_  = ~A168 & ~A169;
  assign \new_[76627]_  = ~A170 & \new_[76626]_ ;
  assign \new_[76630]_  = A166 & ~A167;
  assign \new_[76633]_  = A200 & A199;
  assign \new_[76634]_  = \new_[76633]_  & \new_[76630]_ ;
  assign \new_[76635]_  = \new_[76634]_  & \new_[76627]_ ;
  assign \new_[76639]_  = ~A298 & A266;
  assign \new_[76640]_  = A265 & \new_[76639]_ ;
  assign \new_[76643]_  = ~A300 & A299;
  assign \new_[76646]_  = A302 & ~A301;
  assign \new_[76647]_  = \new_[76646]_  & \new_[76643]_ ;
  assign \new_[76648]_  = \new_[76647]_  & \new_[76640]_ ;
  assign \new_[76652]_  = ~A168 & ~A169;
  assign \new_[76653]_  = ~A170 & \new_[76652]_ ;
  assign \new_[76656]_  = A166 & ~A167;
  assign \new_[76659]_  = A200 & A199;
  assign \new_[76660]_  = \new_[76659]_  & \new_[76656]_ ;
  assign \new_[76661]_  = \new_[76660]_  & \new_[76653]_ ;
  assign \new_[76665]_  = A267 & A266;
  assign \new_[76666]_  = ~A265 & \new_[76665]_ ;
  assign \new_[76669]_  = A300 & A268;
  assign \new_[76672]_  = A302 & ~A301;
  assign \new_[76673]_  = \new_[76672]_  & \new_[76669]_ ;
  assign \new_[76674]_  = \new_[76673]_  & \new_[76666]_ ;
  assign \new_[76678]_  = ~A168 & ~A169;
  assign \new_[76679]_  = ~A170 & \new_[76678]_ ;
  assign \new_[76682]_  = A166 & ~A167;
  assign \new_[76685]_  = A200 & A199;
  assign \new_[76686]_  = \new_[76685]_  & \new_[76682]_ ;
  assign \new_[76687]_  = \new_[76686]_  & \new_[76679]_ ;
  assign \new_[76691]_  = A267 & A266;
  assign \new_[76692]_  = ~A265 & \new_[76691]_ ;
  assign \new_[76695]_  = A300 & ~A269;
  assign \new_[76698]_  = A302 & ~A301;
  assign \new_[76699]_  = \new_[76698]_  & \new_[76695]_ ;
  assign \new_[76700]_  = \new_[76699]_  & \new_[76692]_ ;
  assign \new_[76704]_  = ~A168 & ~A169;
  assign \new_[76705]_  = ~A170 & \new_[76704]_ ;
  assign \new_[76708]_  = A166 & ~A167;
  assign \new_[76711]_  = A200 & A199;
  assign \new_[76712]_  = \new_[76711]_  & \new_[76708]_ ;
  assign \new_[76713]_  = \new_[76712]_  & \new_[76705]_ ;
  assign \new_[76717]_  = ~A267 & A266;
  assign \new_[76718]_  = ~A265 & \new_[76717]_ ;
  assign \new_[76721]_  = A269 & ~A268;
  assign \new_[76724]_  = A301 & ~A300;
  assign \new_[76725]_  = \new_[76724]_  & \new_[76721]_ ;
  assign \new_[76726]_  = \new_[76725]_  & \new_[76718]_ ;
  assign \new_[76730]_  = ~A168 & ~A169;
  assign \new_[76731]_  = ~A170 & \new_[76730]_ ;
  assign \new_[76734]_  = A166 & ~A167;
  assign \new_[76737]_  = A200 & A199;
  assign \new_[76738]_  = \new_[76737]_  & \new_[76734]_ ;
  assign \new_[76739]_  = \new_[76738]_  & \new_[76731]_ ;
  assign \new_[76743]_  = ~A267 & A266;
  assign \new_[76744]_  = ~A265 & \new_[76743]_ ;
  assign \new_[76747]_  = A269 & ~A268;
  assign \new_[76750]_  = ~A302 & ~A300;
  assign \new_[76751]_  = \new_[76750]_  & \new_[76747]_ ;
  assign \new_[76752]_  = \new_[76751]_  & \new_[76744]_ ;
  assign \new_[76756]_  = ~A168 & ~A169;
  assign \new_[76757]_  = ~A170 & \new_[76756]_ ;
  assign \new_[76760]_  = A166 & ~A167;
  assign \new_[76763]_  = A200 & A199;
  assign \new_[76764]_  = \new_[76763]_  & \new_[76760]_ ;
  assign \new_[76765]_  = \new_[76764]_  & \new_[76757]_ ;
  assign \new_[76769]_  = ~A267 & A266;
  assign \new_[76770]_  = ~A265 & \new_[76769]_ ;
  assign \new_[76773]_  = A269 & ~A268;
  assign \new_[76776]_  = A299 & A298;
  assign \new_[76777]_  = \new_[76776]_  & \new_[76773]_ ;
  assign \new_[76778]_  = \new_[76777]_  & \new_[76770]_ ;
  assign \new_[76782]_  = ~A168 & ~A169;
  assign \new_[76783]_  = ~A170 & \new_[76782]_ ;
  assign \new_[76786]_  = A166 & ~A167;
  assign \new_[76789]_  = A200 & A199;
  assign \new_[76790]_  = \new_[76789]_  & \new_[76786]_ ;
  assign \new_[76791]_  = \new_[76790]_  & \new_[76783]_ ;
  assign \new_[76795]_  = ~A267 & A266;
  assign \new_[76796]_  = ~A265 & \new_[76795]_ ;
  assign \new_[76799]_  = A269 & ~A268;
  assign \new_[76802]_  = ~A299 & ~A298;
  assign \new_[76803]_  = \new_[76802]_  & \new_[76799]_ ;
  assign \new_[76804]_  = \new_[76803]_  & \new_[76796]_ ;
  assign \new_[76808]_  = ~A168 & ~A169;
  assign \new_[76809]_  = ~A170 & \new_[76808]_ ;
  assign \new_[76812]_  = A166 & ~A167;
  assign \new_[76815]_  = A200 & A199;
  assign \new_[76816]_  = \new_[76815]_  & \new_[76812]_ ;
  assign \new_[76817]_  = \new_[76816]_  & \new_[76809]_ ;
  assign \new_[76821]_  = A267 & ~A266;
  assign \new_[76822]_  = A265 & \new_[76821]_ ;
  assign \new_[76825]_  = A300 & A268;
  assign \new_[76828]_  = A302 & ~A301;
  assign \new_[76829]_  = \new_[76828]_  & \new_[76825]_ ;
  assign \new_[76830]_  = \new_[76829]_  & \new_[76822]_ ;
  assign \new_[76834]_  = ~A168 & ~A169;
  assign \new_[76835]_  = ~A170 & \new_[76834]_ ;
  assign \new_[76838]_  = A166 & ~A167;
  assign \new_[76841]_  = A200 & A199;
  assign \new_[76842]_  = \new_[76841]_  & \new_[76838]_ ;
  assign \new_[76843]_  = \new_[76842]_  & \new_[76835]_ ;
  assign \new_[76847]_  = A267 & ~A266;
  assign \new_[76848]_  = A265 & \new_[76847]_ ;
  assign \new_[76851]_  = A300 & ~A269;
  assign \new_[76854]_  = A302 & ~A301;
  assign \new_[76855]_  = \new_[76854]_  & \new_[76851]_ ;
  assign \new_[76856]_  = \new_[76855]_  & \new_[76848]_ ;
  assign \new_[76860]_  = ~A168 & ~A169;
  assign \new_[76861]_  = ~A170 & \new_[76860]_ ;
  assign \new_[76864]_  = A166 & ~A167;
  assign \new_[76867]_  = A200 & A199;
  assign \new_[76868]_  = \new_[76867]_  & \new_[76864]_ ;
  assign \new_[76869]_  = \new_[76868]_  & \new_[76861]_ ;
  assign \new_[76873]_  = ~A267 & ~A266;
  assign \new_[76874]_  = A265 & \new_[76873]_ ;
  assign \new_[76877]_  = A269 & ~A268;
  assign \new_[76880]_  = A301 & ~A300;
  assign \new_[76881]_  = \new_[76880]_  & \new_[76877]_ ;
  assign \new_[76882]_  = \new_[76881]_  & \new_[76874]_ ;
  assign \new_[76886]_  = ~A168 & ~A169;
  assign \new_[76887]_  = ~A170 & \new_[76886]_ ;
  assign \new_[76890]_  = A166 & ~A167;
  assign \new_[76893]_  = A200 & A199;
  assign \new_[76894]_  = \new_[76893]_  & \new_[76890]_ ;
  assign \new_[76895]_  = \new_[76894]_  & \new_[76887]_ ;
  assign \new_[76899]_  = ~A267 & ~A266;
  assign \new_[76900]_  = A265 & \new_[76899]_ ;
  assign \new_[76903]_  = A269 & ~A268;
  assign \new_[76906]_  = ~A302 & ~A300;
  assign \new_[76907]_  = \new_[76906]_  & \new_[76903]_ ;
  assign \new_[76908]_  = \new_[76907]_  & \new_[76900]_ ;
  assign \new_[76912]_  = ~A168 & ~A169;
  assign \new_[76913]_  = ~A170 & \new_[76912]_ ;
  assign \new_[76916]_  = A166 & ~A167;
  assign \new_[76919]_  = A200 & A199;
  assign \new_[76920]_  = \new_[76919]_  & \new_[76916]_ ;
  assign \new_[76921]_  = \new_[76920]_  & \new_[76913]_ ;
  assign \new_[76925]_  = ~A267 & ~A266;
  assign \new_[76926]_  = A265 & \new_[76925]_ ;
  assign \new_[76929]_  = A269 & ~A268;
  assign \new_[76932]_  = A299 & A298;
  assign \new_[76933]_  = \new_[76932]_  & \new_[76929]_ ;
  assign \new_[76934]_  = \new_[76933]_  & \new_[76926]_ ;
  assign \new_[76938]_  = ~A168 & ~A169;
  assign \new_[76939]_  = ~A170 & \new_[76938]_ ;
  assign \new_[76942]_  = A166 & ~A167;
  assign \new_[76945]_  = A200 & A199;
  assign \new_[76946]_  = \new_[76945]_  & \new_[76942]_ ;
  assign \new_[76947]_  = \new_[76946]_  & \new_[76939]_ ;
  assign \new_[76951]_  = ~A267 & ~A266;
  assign \new_[76952]_  = A265 & \new_[76951]_ ;
  assign \new_[76955]_  = A269 & ~A268;
  assign \new_[76958]_  = ~A299 & ~A298;
  assign \new_[76959]_  = \new_[76958]_  & \new_[76955]_ ;
  assign \new_[76960]_  = \new_[76959]_  & \new_[76952]_ ;
  assign \new_[76964]_  = ~A168 & ~A169;
  assign \new_[76965]_  = ~A170 & \new_[76964]_ ;
  assign \new_[76968]_  = A166 & ~A167;
  assign \new_[76971]_  = A200 & A199;
  assign \new_[76972]_  = \new_[76971]_  & \new_[76968]_ ;
  assign \new_[76973]_  = \new_[76972]_  & \new_[76965]_ ;
  assign \new_[76977]_  = A298 & ~A266;
  assign \new_[76978]_  = ~A265 & \new_[76977]_ ;
  assign \new_[76981]_  = ~A300 & ~A299;
  assign \new_[76984]_  = A302 & ~A301;
  assign \new_[76985]_  = \new_[76984]_  & \new_[76981]_ ;
  assign \new_[76986]_  = \new_[76985]_  & \new_[76978]_ ;
  assign \new_[76990]_  = ~A168 & ~A169;
  assign \new_[76991]_  = ~A170 & \new_[76990]_ ;
  assign \new_[76994]_  = A166 & ~A167;
  assign \new_[76997]_  = A200 & A199;
  assign \new_[76998]_  = \new_[76997]_  & \new_[76994]_ ;
  assign \new_[76999]_  = \new_[76998]_  & \new_[76991]_ ;
  assign \new_[77003]_  = ~A298 & ~A266;
  assign \new_[77004]_  = ~A265 & \new_[77003]_ ;
  assign \new_[77007]_  = ~A300 & A299;
  assign \new_[77010]_  = A302 & ~A301;
  assign \new_[77011]_  = \new_[77010]_  & \new_[77007]_ ;
  assign \new_[77012]_  = \new_[77011]_  & \new_[77004]_ ;
  assign \new_[77016]_  = ~A168 & ~A169;
  assign \new_[77017]_  = ~A170 & \new_[77016]_ ;
  assign \new_[77020]_  = A166 & ~A167;
  assign \new_[77023]_  = ~A200 & ~A199;
  assign \new_[77024]_  = \new_[77023]_  & \new_[77020]_ ;
  assign \new_[77025]_  = \new_[77024]_  & \new_[77017]_ ;
  assign \new_[77029]_  = A269 & ~A268;
  assign \new_[77030]_  = A267 & \new_[77029]_ ;
  assign \new_[77033]_  = ~A299 & A298;
  assign \new_[77036]_  = A301 & A300;
  assign \new_[77037]_  = \new_[77036]_  & \new_[77033]_ ;
  assign \new_[77038]_  = \new_[77037]_  & \new_[77030]_ ;
  assign \new_[77042]_  = ~A168 & ~A169;
  assign \new_[77043]_  = ~A170 & \new_[77042]_ ;
  assign \new_[77046]_  = A166 & ~A167;
  assign \new_[77049]_  = ~A200 & ~A199;
  assign \new_[77050]_  = \new_[77049]_  & \new_[77046]_ ;
  assign \new_[77051]_  = \new_[77050]_  & \new_[77043]_ ;
  assign \new_[77055]_  = A269 & ~A268;
  assign \new_[77056]_  = A267 & \new_[77055]_ ;
  assign \new_[77059]_  = ~A299 & A298;
  assign \new_[77062]_  = ~A302 & A300;
  assign \new_[77063]_  = \new_[77062]_  & \new_[77059]_ ;
  assign \new_[77064]_  = \new_[77063]_  & \new_[77056]_ ;
  assign \new_[77068]_  = ~A168 & ~A169;
  assign \new_[77069]_  = ~A170 & \new_[77068]_ ;
  assign \new_[77072]_  = A166 & ~A167;
  assign \new_[77075]_  = ~A200 & ~A199;
  assign \new_[77076]_  = \new_[77075]_  & \new_[77072]_ ;
  assign \new_[77077]_  = \new_[77076]_  & \new_[77069]_ ;
  assign \new_[77081]_  = A269 & ~A268;
  assign \new_[77082]_  = A267 & \new_[77081]_ ;
  assign \new_[77085]_  = A299 & ~A298;
  assign \new_[77088]_  = A301 & A300;
  assign \new_[77089]_  = \new_[77088]_  & \new_[77085]_ ;
  assign \new_[77090]_  = \new_[77089]_  & \new_[77082]_ ;
  assign \new_[77094]_  = ~A168 & ~A169;
  assign \new_[77095]_  = ~A170 & \new_[77094]_ ;
  assign \new_[77098]_  = A166 & ~A167;
  assign \new_[77101]_  = ~A200 & ~A199;
  assign \new_[77102]_  = \new_[77101]_  & \new_[77098]_ ;
  assign \new_[77103]_  = \new_[77102]_  & \new_[77095]_ ;
  assign \new_[77107]_  = A269 & ~A268;
  assign \new_[77108]_  = A267 & \new_[77107]_ ;
  assign \new_[77111]_  = A299 & ~A298;
  assign \new_[77114]_  = ~A302 & A300;
  assign \new_[77115]_  = \new_[77114]_  & \new_[77111]_ ;
  assign \new_[77116]_  = \new_[77115]_  & \new_[77108]_ ;
  assign \new_[77120]_  = ~A168 & ~A169;
  assign \new_[77121]_  = ~A170 & \new_[77120]_ ;
  assign \new_[77124]_  = A166 & ~A167;
  assign \new_[77127]_  = ~A200 & ~A199;
  assign \new_[77128]_  = \new_[77127]_  & \new_[77124]_ ;
  assign \new_[77129]_  = \new_[77128]_  & \new_[77121]_ ;
  assign \new_[77133]_  = A298 & A268;
  assign \new_[77134]_  = ~A267 & \new_[77133]_ ;
  assign \new_[77137]_  = ~A300 & ~A299;
  assign \new_[77140]_  = A302 & ~A301;
  assign \new_[77141]_  = \new_[77140]_  & \new_[77137]_ ;
  assign \new_[77142]_  = \new_[77141]_  & \new_[77134]_ ;
  assign \new_[77146]_  = ~A168 & ~A169;
  assign \new_[77147]_  = ~A170 & \new_[77146]_ ;
  assign \new_[77150]_  = A166 & ~A167;
  assign \new_[77153]_  = ~A200 & ~A199;
  assign \new_[77154]_  = \new_[77153]_  & \new_[77150]_ ;
  assign \new_[77155]_  = \new_[77154]_  & \new_[77147]_ ;
  assign \new_[77159]_  = ~A298 & A268;
  assign \new_[77160]_  = ~A267 & \new_[77159]_ ;
  assign \new_[77163]_  = ~A300 & A299;
  assign \new_[77166]_  = A302 & ~A301;
  assign \new_[77167]_  = \new_[77166]_  & \new_[77163]_ ;
  assign \new_[77168]_  = \new_[77167]_  & \new_[77160]_ ;
  assign \new_[77172]_  = ~A168 & ~A169;
  assign \new_[77173]_  = ~A170 & \new_[77172]_ ;
  assign \new_[77176]_  = A166 & ~A167;
  assign \new_[77179]_  = ~A200 & ~A199;
  assign \new_[77180]_  = \new_[77179]_  & \new_[77176]_ ;
  assign \new_[77181]_  = \new_[77180]_  & \new_[77173]_ ;
  assign \new_[77185]_  = A298 & ~A269;
  assign \new_[77186]_  = ~A267 & \new_[77185]_ ;
  assign \new_[77189]_  = ~A300 & ~A299;
  assign \new_[77192]_  = A302 & ~A301;
  assign \new_[77193]_  = \new_[77192]_  & \new_[77189]_ ;
  assign \new_[77194]_  = \new_[77193]_  & \new_[77186]_ ;
  assign \new_[77198]_  = ~A168 & ~A169;
  assign \new_[77199]_  = ~A170 & \new_[77198]_ ;
  assign \new_[77202]_  = A166 & ~A167;
  assign \new_[77205]_  = ~A200 & ~A199;
  assign \new_[77206]_  = \new_[77205]_  & \new_[77202]_ ;
  assign \new_[77207]_  = \new_[77206]_  & \new_[77199]_ ;
  assign \new_[77211]_  = ~A298 & ~A269;
  assign \new_[77212]_  = ~A267 & \new_[77211]_ ;
  assign \new_[77215]_  = ~A300 & A299;
  assign \new_[77218]_  = A302 & ~A301;
  assign \new_[77219]_  = \new_[77218]_  & \new_[77215]_ ;
  assign \new_[77220]_  = \new_[77219]_  & \new_[77212]_ ;
  assign \new_[77224]_  = ~A168 & ~A169;
  assign \new_[77225]_  = ~A170 & \new_[77224]_ ;
  assign \new_[77228]_  = A166 & ~A167;
  assign \new_[77231]_  = ~A200 & ~A199;
  assign \new_[77232]_  = \new_[77231]_  & \new_[77228]_ ;
  assign \new_[77233]_  = \new_[77232]_  & \new_[77225]_ ;
  assign \new_[77237]_  = A298 & A266;
  assign \new_[77238]_  = A265 & \new_[77237]_ ;
  assign \new_[77241]_  = ~A300 & ~A299;
  assign \new_[77244]_  = A302 & ~A301;
  assign \new_[77245]_  = \new_[77244]_  & \new_[77241]_ ;
  assign \new_[77246]_  = \new_[77245]_  & \new_[77238]_ ;
  assign \new_[77250]_  = ~A168 & ~A169;
  assign \new_[77251]_  = ~A170 & \new_[77250]_ ;
  assign \new_[77254]_  = A166 & ~A167;
  assign \new_[77257]_  = ~A200 & ~A199;
  assign \new_[77258]_  = \new_[77257]_  & \new_[77254]_ ;
  assign \new_[77259]_  = \new_[77258]_  & \new_[77251]_ ;
  assign \new_[77263]_  = ~A298 & A266;
  assign \new_[77264]_  = A265 & \new_[77263]_ ;
  assign \new_[77267]_  = ~A300 & A299;
  assign \new_[77270]_  = A302 & ~A301;
  assign \new_[77271]_  = \new_[77270]_  & \new_[77267]_ ;
  assign \new_[77272]_  = \new_[77271]_  & \new_[77264]_ ;
  assign \new_[77276]_  = ~A168 & ~A169;
  assign \new_[77277]_  = ~A170 & \new_[77276]_ ;
  assign \new_[77280]_  = A166 & ~A167;
  assign \new_[77283]_  = ~A200 & ~A199;
  assign \new_[77284]_  = \new_[77283]_  & \new_[77280]_ ;
  assign \new_[77285]_  = \new_[77284]_  & \new_[77277]_ ;
  assign \new_[77289]_  = A267 & A266;
  assign \new_[77290]_  = ~A265 & \new_[77289]_ ;
  assign \new_[77293]_  = A300 & A268;
  assign \new_[77296]_  = A302 & ~A301;
  assign \new_[77297]_  = \new_[77296]_  & \new_[77293]_ ;
  assign \new_[77298]_  = \new_[77297]_  & \new_[77290]_ ;
  assign \new_[77302]_  = ~A168 & ~A169;
  assign \new_[77303]_  = ~A170 & \new_[77302]_ ;
  assign \new_[77306]_  = A166 & ~A167;
  assign \new_[77309]_  = ~A200 & ~A199;
  assign \new_[77310]_  = \new_[77309]_  & \new_[77306]_ ;
  assign \new_[77311]_  = \new_[77310]_  & \new_[77303]_ ;
  assign \new_[77315]_  = A267 & A266;
  assign \new_[77316]_  = ~A265 & \new_[77315]_ ;
  assign \new_[77319]_  = A300 & ~A269;
  assign \new_[77322]_  = A302 & ~A301;
  assign \new_[77323]_  = \new_[77322]_  & \new_[77319]_ ;
  assign \new_[77324]_  = \new_[77323]_  & \new_[77316]_ ;
  assign \new_[77328]_  = ~A168 & ~A169;
  assign \new_[77329]_  = ~A170 & \new_[77328]_ ;
  assign \new_[77332]_  = A166 & ~A167;
  assign \new_[77335]_  = ~A200 & ~A199;
  assign \new_[77336]_  = \new_[77335]_  & \new_[77332]_ ;
  assign \new_[77337]_  = \new_[77336]_  & \new_[77329]_ ;
  assign \new_[77341]_  = ~A267 & A266;
  assign \new_[77342]_  = ~A265 & \new_[77341]_ ;
  assign \new_[77345]_  = A269 & ~A268;
  assign \new_[77348]_  = A301 & ~A300;
  assign \new_[77349]_  = \new_[77348]_  & \new_[77345]_ ;
  assign \new_[77350]_  = \new_[77349]_  & \new_[77342]_ ;
  assign \new_[77354]_  = ~A168 & ~A169;
  assign \new_[77355]_  = ~A170 & \new_[77354]_ ;
  assign \new_[77358]_  = A166 & ~A167;
  assign \new_[77361]_  = ~A200 & ~A199;
  assign \new_[77362]_  = \new_[77361]_  & \new_[77358]_ ;
  assign \new_[77363]_  = \new_[77362]_  & \new_[77355]_ ;
  assign \new_[77367]_  = ~A267 & A266;
  assign \new_[77368]_  = ~A265 & \new_[77367]_ ;
  assign \new_[77371]_  = A269 & ~A268;
  assign \new_[77374]_  = ~A302 & ~A300;
  assign \new_[77375]_  = \new_[77374]_  & \new_[77371]_ ;
  assign \new_[77376]_  = \new_[77375]_  & \new_[77368]_ ;
  assign \new_[77380]_  = ~A168 & ~A169;
  assign \new_[77381]_  = ~A170 & \new_[77380]_ ;
  assign \new_[77384]_  = A166 & ~A167;
  assign \new_[77387]_  = ~A200 & ~A199;
  assign \new_[77388]_  = \new_[77387]_  & \new_[77384]_ ;
  assign \new_[77389]_  = \new_[77388]_  & \new_[77381]_ ;
  assign \new_[77393]_  = ~A267 & A266;
  assign \new_[77394]_  = ~A265 & \new_[77393]_ ;
  assign \new_[77397]_  = A269 & ~A268;
  assign \new_[77400]_  = A299 & A298;
  assign \new_[77401]_  = \new_[77400]_  & \new_[77397]_ ;
  assign \new_[77402]_  = \new_[77401]_  & \new_[77394]_ ;
  assign \new_[77406]_  = ~A168 & ~A169;
  assign \new_[77407]_  = ~A170 & \new_[77406]_ ;
  assign \new_[77410]_  = A166 & ~A167;
  assign \new_[77413]_  = ~A200 & ~A199;
  assign \new_[77414]_  = \new_[77413]_  & \new_[77410]_ ;
  assign \new_[77415]_  = \new_[77414]_  & \new_[77407]_ ;
  assign \new_[77419]_  = ~A267 & A266;
  assign \new_[77420]_  = ~A265 & \new_[77419]_ ;
  assign \new_[77423]_  = A269 & ~A268;
  assign \new_[77426]_  = ~A299 & ~A298;
  assign \new_[77427]_  = \new_[77426]_  & \new_[77423]_ ;
  assign \new_[77428]_  = \new_[77427]_  & \new_[77420]_ ;
  assign \new_[77432]_  = ~A168 & ~A169;
  assign \new_[77433]_  = ~A170 & \new_[77432]_ ;
  assign \new_[77436]_  = A166 & ~A167;
  assign \new_[77439]_  = ~A200 & ~A199;
  assign \new_[77440]_  = \new_[77439]_  & \new_[77436]_ ;
  assign \new_[77441]_  = \new_[77440]_  & \new_[77433]_ ;
  assign \new_[77445]_  = A267 & ~A266;
  assign \new_[77446]_  = A265 & \new_[77445]_ ;
  assign \new_[77449]_  = A300 & A268;
  assign \new_[77452]_  = A302 & ~A301;
  assign \new_[77453]_  = \new_[77452]_  & \new_[77449]_ ;
  assign \new_[77454]_  = \new_[77453]_  & \new_[77446]_ ;
  assign \new_[77458]_  = ~A168 & ~A169;
  assign \new_[77459]_  = ~A170 & \new_[77458]_ ;
  assign \new_[77462]_  = A166 & ~A167;
  assign \new_[77465]_  = ~A200 & ~A199;
  assign \new_[77466]_  = \new_[77465]_  & \new_[77462]_ ;
  assign \new_[77467]_  = \new_[77466]_  & \new_[77459]_ ;
  assign \new_[77471]_  = A267 & ~A266;
  assign \new_[77472]_  = A265 & \new_[77471]_ ;
  assign \new_[77475]_  = A300 & ~A269;
  assign \new_[77478]_  = A302 & ~A301;
  assign \new_[77479]_  = \new_[77478]_  & \new_[77475]_ ;
  assign \new_[77480]_  = \new_[77479]_  & \new_[77472]_ ;
  assign \new_[77484]_  = ~A168 & ~A169;
  assign \new_[77485]_  = ~A170 & \new_[77484]_ ;
  assign \new_[77488]_  = A166 & ~A167;
  assign \new_[77491]_  = ~A200 & ~A199;
  assign \new_[77492]_  = \new_[77491]_  & \new_[77488]_ ;
  assign \new_[77493]_  = \new_[77492]_  & \new_[77485]_ ;
  assign \new_[77497]_  = ~A267 & ~A266;
  assign \new_[77498]_  = A265 & \new_[77497]_ ;
  assign \new_[77501]_  = A269 & ~A268;
  assign \new_[77504]_  = A301 & ~A300;
  assign \new_[77505]_  = \new_[77504]_  & \new_[77501]_ ;
  assign \new_[77506]_  = \new_[77505]_  & \new_[77498]_ ;
  assign \new_[77510]_  = ~A168 & ~A169;
  assign \new_[77511]_  = ~A170 & \new_[77510]_ ;
  assign \new_[77514]_  = A166 & ~A167;
  assign \new_[77517]_  = ~A200 & ~A199;
  assign \new_[77518]_  = \new_[77517]_  & \new_[77514]_ ;
  assign \new_[77519]_  = \new_[77518]_  & \new_[77511]_ ;
  assign \new_[77523]_  = ~A267 & ~A266;
  assign \new_[77524]_  = A265 & \new_[77523]_ ;
  assign \new_[77527]_  = A269 & ~A268;
  assign \new_[77530]_  = ~A302 & ~A300;
  assign \new_[77531]_  = \new_[77530]_  & \new_[77527]_ ;
  assign \new_[77532]_  = \new_[77531]_  & \new_[77524]_ ;
  assign \new_[77536]_  = ~A168 & ~A169;
  assign \new_[77537]_  = ~A170 & \new_[77536]_ ;
  assign \new_[77540]_  = A166 & ~A167;
  assign \new_[77543]_  = ~A200 & ~A199;
  assign \new_[77544]_  = \new_[77543]_  & \new_[77540]_ ;
  assign \new_[77545]_  = \new_[77544]_  & \new_[77537]_ ;
  assign \new_[77549]_  = ~A267 & ~A266;
  assign \new_[77550]_  = A265 & \new_[77549]_ ;
  assign \new_[77553]_  = A269 & ~A268;
  assign \new_[77556]_  = A299 & A298;
  assign \new_[77557]_  = \new_[77556]_  & \new_[77553]_ ;
  assign \new_[77558]_  = \new_[77557]_  & \new_[77550]_ ;
  assign \new_[77562]_  = ~A168 & ~A169;
  assign \new_[77563]_  = ~A170 & \new_[77562]_ ;
  assign \new_[77566]_  = A166 & ~A167;
  assign \new_[77569]_  = ~A200 & ~A199;
  assign \new_[77570]_  = \new_[77569]_  & \new_[77566]_ ;
  assign \new_[77571]_  = \new_[77570]_  & \new_[77563]_ ;
  assign \new_[77575]_  = ~A267 & ~A266;
  assign \new_[77576]_  = A265 & \new_[77575]_ ;
  assign \new_[77579]_  = A269 & ~A268;
  assign \new_[77582]_  = ~A299 & ~A298;
  assign \new_[77583]_  = \new_[77582]_  & \new_[77579]_ ;
  assign \new_[77584]_  = \new_[77583]_  & \new_[77576]_ ;
  assign \new_[77588]_  = ~A168 & ~A169;
  assign \new_[77589]_  = ~A170 & \new_[77588]_ ;
  assign \new_[77592]_  = A166 & ~A167;
  assign \new_[77595]_  = ~A200 & ~A199;
  assign \new_[77596]_  = \new_[77595]_  & \new_[77592]_ ;
  assign \new_[77597]_  = \new_[77596]_  & \new_[77589]_ ;
  assign \new_[77601]_  = A298 & ~A266;
  assign \new_[77602]_  = ~A265 & \new_[77601]_ ;
  assign \new_[77605]_  = ~A300 & ~A299;
  assign \new_[77608]_  = A302 & ~A301;
  assign \new_[77609]_  = \new_[77608]_  & \new_[77605]_ ;
  assign \new_[77610]_  = \new_[77609]_  & \new_[77602]_ ;
  assign \new_[77614]_  = ~A168 & ~A169;
  assign \new_[77615]_  = ~A170 & \new_[77614]_ ;
  assign \new_[77618]_  = A166 & ~A167;
  assign \new_[77621]_  = ~A200 & ~A199;
  assign \new_[77622]_  = \new_[77621]_  & \new_[77618]_ ;
  assign \new_[77623]_  = \new_[77622]_  & \new_[77615]_ ;
  assign \new_[77627]_  = ~A298 & ~A266;
  assign \new_[77628]_  = ~A265 & \new_[77627]_ ;
  assign \new_[77631]_  = ~A300 & A299;
  assign \new_[77634]_  = A302 & ~A301;
  assign \new_[77635]_  = \new_[77634]_  & \new_[77631]_ ;
  assign \new_[77636]_  = \new_[77635]_  & \new_[77628]_ ;
  assign \new_[77640]_  = ~A199 & A166;
  assign \new_[77641]_  = A167 & \new_[77640]_ ;
  assign \new_[77644]_  = A201 & A200;
  assign \new_[77647]_  = ~A265 & A202;
  assign \new_[77648]_  = \new_[77647]_  & \new_[77644]_ ;
  assign \new_[77649]_  = \new_[77648]_  & \new_[77641]_ ;
  assign \new_[77652]_  = A267 & A266;
  assign \new_[77655]_  = A298 & A268;
  assign \new_[77656]_  = \new_[77655]_  & \new_[77652]_ ;
  assign \new_[77659]_  = ~A300 & ~A299;
  assign \new_[77662]_  = A302 & ~A301;
  assign \new_[77663]_  = \new_[77662]_  & \new_[77659]_ ;
  assign \new_[77664]_  = \new_[77663]_  & \new_[77656]_ ;
  assign \new_[77668]_  = ~A199 & A166;
  assign \new_[77669]_  = A167 & \new_[77668]_ ;
  assign \new_[77672]_  = A201 & A200;
  assign \new_[77675]_  = ~A265 & A202;
  assign \new_[77676]_  = \new_[77675]_  & \new_[77672]_ ;
  assign \new_[77677]_  = \new_[77676]_  & \new_[77669]_ ;
  assign \new_[77680]_  = A267 & A266;
  assign \new_[77683]_  = ~A298 & A268;
  assign \new_[77684]_  = \new_[77683]_  & \new_[77680]_ ;
  assign \new_[77687]_  = ~A300 & A299;
  assign \new_[77690]_  = A302 & ~A301;
  assign \new_[77691]_  = \new_[77690]_  & \new_[77687]_ ;
  assign \new_[77692]_  = \new_[77691]_  & \new_[77684]_ ;
  assign \new_[77696]_  = ~A199 & A166;
  assign \new_[77697]_  = A167 & \new_[77696]_ ;
  assign \new_[77700]_  = A201 & A200;
  assign \new_[77703]_  = ~A265 & A202;
  assign \new_[77704]_  = \new_[77703]_  & \new_[77700]_ ;
  assign \new_[77705]_  = \new_[77704]_  & \new_[77697]_ ;
  assign \new_[77708]_  = A267 & A266;
  assign \new_[77711]_  = A298 & ~A269;
  assign \new_[77712]_  = \new_[77711]_  & \new_[77708]_ ;
  assign \new_[77715]_  = ~A300 & ~A299;
  assign \new_[77718]_  = A302 & ~A301;
  assign \new_[77719]_  = \new_[77718]_  & \new_[77715]_ ;
  assign \new_[77720]_  = \new_[77719]_  & \new_[77712]_ ;
  assign \new_[77724]_  = ~A199 & A166;
  assign \new_[77725]_  = A167 & \new_[77724]_ ;
  assign \new_[77728]_  = A201 & A200;
  assign \new_[77731]_  = ~A265 & A202;
  assign \new_[77732]_  = \new_[77731]_  & \new_[77728]_ ;
  assign \new_[77733]_  = \new_[77732]_  & \new_[77725]_ ;
  assign \new_[77736]_  = A267 & A266;
  assign \new_[77739]_  = ~A298 & ~A269;
  assign \new_[77740]_  = \new_[77739]_  & \new_[77736]_ ;
  assign \new_[77743]_  = ~A300 & A299;
  assign \new_[77746]_  = A302 & ~A301;
  assign \new_[77747]_  = \new_[77746]_  & \new_[77743]_ ;
  assign \new_[77748]_  = \new_[77747]_  & \new_[77740]_ ;
  assign \new_[77752]_  = ~A199 & A166;
  assign \new_[77753]_  = A167 & \new_[77752]_ ;
  assign \new_[77756]_  = A201 & A200;
  assign \new_[77759]_  = ~A265 & A202;
  assign \new_[77760]_  = \new_[77759]_  & \new_[77756]_ ;
  assign \new_[77761]_  = \new_[77760]_  & \new_[77753]_ ;
  assign \new_[77764]_  = ~A267 & A266;
  assign \new_[77767]_  = A269 & ~A268;
  assign \new_[77768]_  = \new_[77767]_  & \new_[77764]_ ;
  assign \new_[77771]_  = ~A299 & A298;
  assign \new_[77774]_  = A301 & A300;
  assign \new_[77775]_  = \new_[77774]_  & \new_[77771]_ ;
  assign \new_[77776]_  = \new_[77775]_  & \new_[77768]_ ;
  assign \new_[77780]_  = ~A199 & A166;
  assign \new_[77781]_  = A167 & \new_[77780]_ ;
  assign \new_[77784]_  = A201 & A200;
  assign \new_[77787]_  = ~A265 & A202;
  assign \new_[77788]_  = \new_[77787]_  & \new_[77784]_ ;
  assign \new_[77789]_  = \new_[77788]_  & \new_[77781]_ ;
  assign \new_[77792]_  = ~A267 & A266;
  assign \new_[77795]_  = A269 & ~A268;
  assign \new_[77796]_  = \new_[77795]_  & \new_[77792]_ ;
  assign \new_[77799]_  = ~A299 & A298;
  assign \new_[77802]_  = ~A302 & A300;
  assign \new_[77803]_  = \new_[77802]_  & \new_[77799]_ ;
  assign \new_[77804]_  = \new_[77803]_  & \new_[77796]_ ;
  assign \new_[77808]_  = ~A199 & A166;
  assign \new_[77809]_  = A167 & \new_[77808]_ ;
  assign \new_[77812]_  = A201 & A200;
  assign \new_[77815]_  = ~A265 & A202;
  assign \new_[77816]_  = \new_[77815]_  & \new_[77812]_ ;
  assign \new_[77817]_  = \new_[77816]_  & \new_[77809]_ ;
  assign \new_[77820]_  = ~A267 & A266;
  assign \new_[77823]_  = A269 & ~A268;
  assign \new_[77824]_  = \new_[77823]_  & \new_[77820]_ ;
  assign \new_[77827]_  = A299 & ~A298;
  assign \new_[77830]_  = A301 & A300;
  assign \new_[77831]_  = \new_[77830]_  & \new_[77827]_ ;
  assign \new_[77832]_  = \new_[77831]_  & \new_[77824]_ ;
  assign \new_[77836]_  = ~A199 & A166;
  assign \new_[77837]_  = A167 & \new_[77836]_ ;
  assign \new_[77840]_  = A201 & A200;
  assign \new_[77843]_  = ~A265 & A202;
  assign \new_[77844]_  = \new_[77843]_  & \new_[77840]_ ;
  assign \new_[77845]_  = \new_[77844]_  & \new_[77837]_ ;
  assign \new_[77848]_  = ~A267 & A266;
  assign \new_[77851]_  = A269 & ~A268;
  assign \new_[77852]_  = \new_[77851]_  & \new_[77848]_ ;
  assign \new_[77855]_  = A299 & ~A298;
  assign \new_[77858]_  = ~A302 & A300;
  assign \new_[77859]_  = \new_[77858]_  & \new_[77855]_ ;
  assign \new_[77860]_  = \new_[77859]_  & \new_[77852]_ ;
  assign \new_[77864]_  = ~A199 & A166;
  assign \new_[77865]_  = A167 & \new_[77864]_ ;
  assign \new_[77868]_  = A201 & A200;
  assign \new_[77871]_  = A265 & A202;
  assign \new_[77872]_  = \new_[77871]_  & \new_[77868]_ ;
  assign \new_[77873]_  = \new_[77872]_  & \new_[77865]_ ;
  assign \new_[77876]_  = A267 & ~A266;
  assign \new_[77879]_  = A298 & A268;
  assign \new_[77880]_  = \new_[77879]_  & \new_[77876]_ ;
  assign \new_[77883]_  = ~A300 & ~A299;
  assign \new_[77886]_  = A302 & ~A301;
  assign \new_[77887]_  = \new_[77886]_  & \new_[77883]_ ;
  assign \new_[77888]_  = \new_[77887]_  & \new_[77880]_ ;
  assign \new_[77892]_  = ~A199 & A166;
  assign \new_[77893]_  = A167 & \new_[77892]_ ;
  assign \new_[77896]_  = A201 & A200;
  assign \new_[77899]_  = A265 & A202;
  assign \new_[77900]_  = \new_[77899]_  & \new_[77896]_ ;
  assign \new_[77901]_  = \new_[77900]_  & \new_[77893]_ ;
  assign \new_[77904]_  = A267 & ~A266;
  assign \new_[77907]_  = ~A298 & A268;
  assign \new_[77908]_  = \new_[77907]_  & \new_[77904]_ ;
  assign \new_[77911]_  = ~A300 & A299;
  assign \new_[77914]_  = A302 & ~A301;
  assign \new_[77915]_  = \new_[77914]_  & \new_[77911]_ ;
  assign \new_[77916]_  = \new_[77915]_  & \new_[77908]_ ;
  assign \new_[77920]_  = ~A199 & A166;
  assign \new_[77921]_  = A167 & \new_[77920]_ ;
  assign \new_[77924]_  = A201 & A200;
  assign \new_[77927]_  = A265 & A202;
  assign \new_[77928]_  = \new_[77927]_  & \new_[77924]_ ;
  assign \new_[77929]_  = \new_[77928]_  & \new_[77921]_ ;
  assign \new_[77932]_  = A267 & ~A266;
  assign \new_[77935]_  = A298 & ~A269;
  assign \new_[77936]_  = \new_[77935]_  & \new_[77932]_ ;
  assign \new_[77939]_  = ~A300 & ~A299;
  assign \new_[77942]_  = A302 & ~A301;
  assign \new_[77943]_  = \new_[77942]_  & \new_[77939]_ ;
  assign \new_[77944]_  = \new_[77943]_  & \new_[77936]_ ;
  assign \new_[77948]_  = ~A199 & A166;
  assign \new_[77949]_  = A167 & \new_[77948]_ ;
  assign \new_[77952]_  = A201 & A200;
  assign \new_[77955]_  = A265 & A202;
  assign \new_[77956]_  = \new_[77955]_  & \new_[77952]_ ;
  assign \new_[77957]_  = \new_[77956]_  & \new_[77949]_ ;
  assign \new_[77960]_  = A267 & ~A266;
  assign \new_[77963]_  = ~A298 & ~A269;
  assign \new_[77964]_  = \new_[77963]_  & \new_[77960]_ ;
  assign \new_[77967]_  = ~A300 & A299;
  assign \new_[77970]_  = A302 & ~A301;
  assign \new_[77971]_  = \new_[77970]_  & \new_[77967]_ ;
  assign \new_[77972]_  = \new_[77971]_  & \new_[77964]_ ;
  assign \new_[77976]_  = ~A199 & A166;
  assign \new_[77977]_  = A167 & \new_[77976]_ ;
  assign \new_[77980]_  = A201 & A200;
  assign \new_[77983]_  = A265 & A202;
  assign \new_[77984]_  = \new_[77983]_  & \new_[77980]_ ;
  assign \new_[77985]_  = \new_[77984]_  & \new_[77977]_ ;
  assign \new_[77988]_  = ~A267 & ~A266;
  assign \new_[77991]_  = A269 & ~A268;
  assign \new_[77992]_  = \new_[77991]_  & \new_[77988]_ ;
  assign \new_[77995]_  = ~A299 & A298;
  assign \new_[77998]_  = A301 & A300;
  assign \new_[77999]_  = \new_[77998]_  & \new_[77995]_ ;
  assign \new_[78000]_  = \new_[77999]_  & \new_[77992]_ ;
  assign \new_[78004]_  = ~A199 & A166;
  assign \new_[78005]_  = A167 & \new_[78004]_ ;
  assign \new_[78008]_  = A201 & A200;
  assign \new_[78011]_  = A265 & A202;
  assign \new_[78012]_  = \new_[78011]_  & \new_[78008]_ ;
  assign \new_[78013]_  = \new_[78012]_  & \new_[78005]_ ;
  assign \new_[78016]_  = ~A267 & ~A266;
  assign \new_[78019]_  = A269 & ~A268;
  assign \new_[78020]_  = \new_[78019]_  & \new_[78016]_ ;
  assign \new_[78023]_  = ~A299 & A298;
  assign \new_[78026]_  = ~A302 & A300;
  assign \new_[78027]_  = \new_[78026]_  & \new_[78023]_ ;
  assign \new_[78028]_  = \new_[78027]_  & \new_[78020]_ ;
  assign \new_[78032]_  = ~A199 & A166;
  assign \new_[78033]_  = A167 & \new_[78032]_ ;
  assign \new_[78036]_  = A201 & A200;
  assign \new_[78039]_  = A265 & A202;
  assign \new_[78040]_  = \new_[78039]_  & \new_[78036]_ ;
  assign \new_[78041]_  = \new_[78040]_  & \new_[78033]_ ;
  assign \new_[78044]_  = ~A267 & ~A266;
  assign \new_[78047]_  = A269 & ~A268;
  assign \new_[78048]_  = \new_[78047]_  & \new_[78044]_ ;
  assign \new_[78051]_  = A299 & ~A298;
  assign \new_[78054]_  = A301 & A300;
  assign \new_[78055]_  = \new_[78054]_  & \new_[78051]_ ;
  assign \new_[78056]_  = \new_[78055]_  & \new_[78048]_ ;
  assign \new_[78060]_  = ~A199 & A166;
  assign \new_[78061]_  = A167 & \new_[78060]_ ;
  assign \new_[78064]_  = A201 & A200;
  assign \new_[78067]_  = A265 & A202;
  assign \new_[78068]_  = \new_[78067]_  & \new_[78064]_ ;
  assign \new_[78069]_  = \new_[78068]_  & \new_[78061]_ ;
  assign \new_[78072]_  = ~A267 & ~A266;
  assign \new_[78075]_  = A269 & ~A268;
  assign \new_[78076]_  = \new_[78075]_  & \new_[78072]_ ;
  assign \new_[78079]_  = A299 & ~A298;
  assign \new_[78082]_  = ~A302 & A300;
  assign \new_[78083]_  = \new_[78082]_  & \new_[78079]_ ;
  assign \new_[78084]_  = \new_[78083]_  & \new_[78076]_ ;
  assign \new_[78088]_  = ~A199 & A166;
  assign \new_[78089]_  = A167 & \new_[78088]_ ;
  assign \new_[78092]_  = A201 & A200;
  assign \new_[78095]_  = ~A265 & ~A203;
  assign \new_[78096]_  = \new_[78095]_  & \new_[78092]_ ;
  assign \new_[78097]_  = \new_[78096]_  & \new_[78089]_ ;
  assign \new_[78100]_  = A267 & A266;
  assign \new_[78103]_  = A298 & A268;
  assign \new_[78104]_  = \new_[78103]_  & \new_[78100]_ ;
  assign \new_[78107]_  = ~A300 & ~A299;
  assign \new_[78110]_  = A302 & ~A301;
  assign \new_[78111]_  = \new_[78110]_  & \new_[78107]_ ;
  assign \new_[78112]_  = \new_[78111]_  & \new_[78104]_ ;
  assign \new_[78116]_  = ~A199 & A166;
  assign \new_[78117]_  = A167 & \new_[78116]_ ;
  assign \new_[78120]_  = A201 & A200;
  assign \new_[78123]_  = ~A265 & ~A203;
  assign \new_[78124]_  = \new_[78123]_  & \new_[78120]_ ;
  assign \new_[78125]_  = \new_[78124]_  & \new_[78117]_ ;
  assign \new_[78128]_  = A267 & A266;
  assign \new_[78131]_  = ~A298 & A268;
  assign \new_[78132]_  = \new_[78131]_  & \new_[78128]_ ;
  assign \new_[78135]_  = ~A300 & A299;
  assign \new_[78138]_  = A302 & ~A301;
  assign \new_[78139]_  = \new_[78138]_  & \new_[78135]_ ;
  assign \new_[78140]_  = \new_[78139]_  & \new_[78132]_ ;
  assign \new_[78144]_  = ~A199 & A166;
  assign \new_[78145]_  = A167 & \new_[78144]_ ;
  assign \new_[78148]_  = A201 & A200;
  assign \new_[78151]_  = ~A265 & ~A203;
  assign \new_[78152]_  = \new_[78151]_  & \new_[78148]_ ;
  assign \new_[78153]_  = \new_[78152]_  & \new_[78145]_ ;
  assign \new_[78156]_  = A267 & A266;
  assign \new_[78159]_  = A298 & ~A269;
  assign \new_[78160]_  = \new_[78159]_  & \new_[78156]_ ;
  assign \new_[78163]_  = ~A300 & ~A299;
  assign \new_[78166]_  = A302 & ~A301;
  assign \new_[78167]_  = \new_[78166]_  & \new_[78163]_ ;
  assign \new_[78168]_  = \new_[78167]_  & \new_[78160]_ ;
  assign \new_[78172]_  = ~A199 & A166;
  assign \new_[78173]_  = A167 & \new_[78172]_ ;
  assign \new_[78176]_  = A201 & A200;
  assign \new_[78179]_  = ~A265 & ~A203;
  assign \new_[78180]_  = \new_[78179]_  & \new_[78176]_ ;
  assign \new_[78181]_  = \new_[78180]_  & \new_[78173]_ ;
  assign \new_[78184]_  = A267 & A266;
  assign \new_[78187]_  = ~A298 & ~A269;
  assign \new_[78188]_  = \new_[78187]_  & \new_[78184]_ ;
  assign \new_[78191]_  = ~A300 & A299;
  assign \new_[78194]_  = A302 & ~A301;
  assign \new_[78195]_  = \new_[78194]_  & \new_[78191]_ ;
  assign \new_[78196]_  = \new_[78195]_  & \new_[78188]_ ;
  assign \new_[78200]_  = ~A199 & A166;
  assign \new_[78201]_  = A167 & \new_[78200]_ ;
  assign \new_[78204]_  = A201 & A200;
  assign \new_[78207]_  = ~A265 & ~A203;
  assign \new_[78208]_  = \new_[78207]_  & \new_[78204]_ ;
  assign \new_[78209]_  = \new_[78208]_  & \new_[78201]_ ;
  assign \new_[78212]_  = ~A267 & A266;
  assign \new_[78215]_  = A269 & ~A268;
  assign \new_[78216]_  = \new_[78215]_  & \new_[78212]_ ;
  assign \new_[78219]_  = ~A299 & A298;
  assign \new_[78222]_  = A301 & A300;
  assign \new_[78223]_  = \new_[78222]_  & \new_[78219]_ ;
  assign \new_[78224]_  = \new_[78223]_  & \new_[78216]_ ;
  assign \new_[78228]_  = ~A199 & A166;
  assign \new_[78229]_  = A167 & \new_[78228]_ ;
  assign \new_[78232]_  = A201 & A200;
  assign \new_[78235]_  = ~A265 & ~A203;
  assign \new_[78236]_  = \new_[78235]_  & \new_[78232]_ ;
  assign \new_[78237]_  = \new_[78236]_  & \new_[78229]_ ;
  assign \new_[78240]_  = ~A267 & A266;
  assign \new_[78243]_  = A269 & ~A268;
  assign \new_[78244]_  = \new_[78243]_  & \new_[78240]_ ;
  assign \new_[78247]_  = ~A299 & A298;
  assign \new_[78250]_  = ~A302 & A300;
  assign \new_[78251]_  = \new_[78250]_  & \new_[78247]_ ;
  assign \new_[78252]_  = \new_[78251]_  & \new_[78244]_ ;
  assign \new_[78256]_  = ~A199 & A166;
  assign \new_[78257]_  = A167 & \new_[78256]_ ;
  assign \new_[78260]_  = A201 & A200;
  assign \new_[78263]_  = ~A265 & ~A203;
  assign \new_[78264]_  = \new_[78263]_  & \new_[78260]_ ;
  assign \new_[78265]_  = \new_[78264]_  & \new_[78257]_ ;
  assign \new_[78268]_  = ~A267 & A266;
  assign \new_[78271]_  = A269 & ~A268;
  assign \new_[78272]_  = \new_[78271]_  & \new_[78268]_ ;
  assign \new_[78275]_  = A299 & ~A298;
  assign \new_[78278]_  = A301 & A300;
  assign \new_[78279]_  = \new_[78278]_  & \new_[78275]_ ;
  assign \new_[78280]_  = \new_[78279]_  & \new_[78272]_ ;
  assign \new_[78284]_  = ~A199 & A166;
  assign \new_[78285]_  = A167 & \new_[78284]_ ;
  assign \new_[78288]_  = A201 & A200;
  assign \new_[78291]_  = ~A265 & ~A203;
  assign \new_[78292]_  = \new_[78291]_  & \new_[78288]_ ;
  assign \new_[78293]_  = \new_[78292]_  & \new_[78285]_ ;
  assign \new_[78296]_  = ~A267 & A266;
  assign \new_[78299]_  = A269 & ~A268;
  assign \new_[78300]_  = \new_[78299]_  & \new_[78296]_ ;
  assign \new_[78303]_  = A299 & ~A298;
  assign \new_[78306]_  = ~A302 & A300;
  assign \new_[78307]_  = \new_[78306]_  & \new_[78303]_ ;
  assign \new_[78308]_  = \new_[78307]_  & \new_[78300]_ ;
  assign \new_[78312]_  = ~A199 & A166;
  assign \new_[78313]_  = A167 & \new_[78312]_ ;
  assign \new_[78316]_  = A201 & A200;
  assign \new_[78319]_  = A265 & ~A203;
  assign \new_[78320]_  = \new_[78319]_  & \new_[78316]_ ;
  assign \new_[78321]_  = \new_[78320]_  & \new_[78313]_ ;
  assign \new_[78324]_  = A267 & ~A266;
  assign \new_[78327]_  = A298 & A268;
  assign \new_[78328]_  = \new_[78327]_  & \new_[78324]_ ;
  assign \new_[78331]_  = ~A300 & ~A299;
  assign \new_[78334]_  = A302 & ~A301;
  assign \new_[78335]_  = \new_[78334]_  & \new_[78331]_ ;
  assign \new_[78336]_  = \new_[78335]_  & \new_[78328]_ ;
  assign \new_[78340]_  = ~A199 & A166;
  assign \new_[78341]_  = A167 & \new_[78340]_ ;
  assign \new_[78344]_  = A201 & A200;
  assign \new_[78347]_  = A265 & ~A203;
  assign \new_[78348]_  = \new_[78347]_  & \new_[78344]_ ;
  assign \new_[78349]_  = \new_[78348]_  & \new_[78341]_ ;
  assign \new_[78352]_  = A267 & ~A266;
  assign \new_[78355]_  = ~A298 & A268;
  assign \new_[78356]_  = \new_[78355]_  & \new_[78352]_ ;
  assign \new_[78359]_  = ~A300 & A299;
  assign \new_[78362]_  = A302 & ~A301;
  assign \new_[78363]_  = \new_[78362]_  & \new_[78359]_ ;
  assign \new_[78364]_  = \new_[78363]_  & \new_[78356]_ ;
  assign \new_[78368]_  = ~A199 & A166;
  assign \new_[78369]_  = A167 & \new_[78368]_ ;
  assign \new_[78372]_  = A201 & A200;
  assign \new_[78375]_  = A265 & ~A203;
  assign \new_[78376]_  = \new_[78375]_  & \new_[78372]_ ;
  assign \new_[78377]_  = \new_[78376]_  & \new_[78369]_ ;
  assign \new_[78380]_  = A267 & ~A266;
  assign \new_[78383]_  = A298 & ~A269;
  assign \new_[78384]_  = \new_[78383]_  & \new_[78380]_ ;
  assign \new_[78387]_  = ~A300 & ~A299;
  assign \new_[78390]_  = A302 & ~A301;
  assign \new_[78391]_  = \new_[78390]_  & \new_[78387]_ ;
  assign \new_[78392]_  = \new_[78391]_  & \new_[78384]_ ;
  assign \new_[78396]_  = ~A199 & A166;
  assign \new_[78397]_  = A167 & \new_[78396]_ ;
  assign \new_[78400]_  = A201 & A200;
  assign \new_[78403]_  = A265 & ~A203;
  assign \new_[78404]_  = \new_[78403]_  & \new_[78400]_ ;
  assign \new_[78405]_  = \new_[78404]_  & \new_[78397]_ ;
  assign \new_[78408]_  = A267 & ~A266;
  assign \new_[78411]_  = ~A298 & ~A269;
  assign \new_[78412]_  = \new_[78411]_  & \new_[78408]_ ;
  assign \new_[78415]_  = ~A300 & A299;
  assign \new_[78418]_  = A302 & ~A301;
  assign \new_[78419]_  = \new_[78418]_  & \new_[78415]_ ;
  assign \new_[78420]_  = \new_[78419]_  & \new_[78412]_ ;
  assign \new_[78424]_  = ~A199 & A166;
  assign \new_[78425]_  = A167 & \new_[78424]_ ;
  assign \new_[78428]_  = A201 & A200;
  assign \new_[78431]_  = A265 & ~A203;
  assign \new_[78432]_  = \new_[78431]_  & \new_[78428]_ ;
  assign \new_[78433]_  = \new_[78432]_  & \new_[78425]_ ;
  assign \new_[78436]_  = ~A267 & ~A266;
  assign \new_[78439]_  = A269 & ~A268;
  assign \new_[78440]_  = \new_[78439]_  & \new_[78436]_ ;
  assign \new_[78443]_  = ~A299 & A298;
  assign \new_[78446]_  = A301 & A300;
  assign \new_[78447]_  = \new_[78446]_  & \new_[78443]_ ;
  assign \new_[78448]_  = \new_[78447]_  & \new_[78440]_ ;
  assign \new_[78452]_  = ~A199 & A166;
  assign \new_[78453]_  = A167 & \new_[78452]_ ;
  assign \new_[78456]_  = A201 & A200;
  assign \new_[78459]_  = A265 & ~A203;
  assign \new_[78460]_  = \new_[78459]_  & \new_[78456]_ ;
  assign \new_[78461]_  = \new_[78460]_  & \new_[78453]_ ;
  assign \new_[78464]_  = ~A267 & ~A266;
  assign \new_[78467]_  = A269 & ~A268;
  assign \new_[78468]_  = \new_[78467]_  & \new_[78464]_ ;
  assign \new_[78471]_  = ~A299 & A298;
  assign \new_[78474]_  = ~A302 & A300;
  assign \new_[78475]_  = \new_[78474]_  & \new_[78471]_ ;
  assign \new_[78476]_  = \new_[78475]_  & \new_[78468]_ ;
  assign \new_[78480]_  = ~A199 & A166;
  assign \new_[78481]_  = A167 & \new_[78480]_ ;
  assign \new_[78484]_  = A201 & A200;
  assign \new_[78487]_  = A265 & ~A203;
  assign \new_[78488]_  = \new_[78487]_  & \new_[78484]_ ;
  assign \new_[78489]_  = \new_[78488]_  & \new_[78481]_ ;
  assign \new_[78492]_  = ~A267 & ~A266;
  assign \new_[78495]_  = A269 & ~A268;
  assign \new_[78496]_  = \new_[78495]_  & \new_[78492]_ ;
  assign \new_[78499]_  = A299 & ~A298;
  assign \new_[78502]_  = A301 & A300;
  assign \new_[78503]_  = \new_[78502]_  & \new_[78499]_ ;
  assign \new_[78504]_  = \new_[78503]_  & \new_[78496]_ ;
  assign \new_[78508]_  = ~A199 & A166;
  assign \new_[78509]_  = A167 & \new_[78508]_ ;
  assign \new_[78512]_  = A201 & A200;
  assign \new_[78515]_  = A265 & ~A203;
  assign \new_[78516]_  = \new_[78515]_  & \new_[78512]_ ;
  assign \new_[78517]_  = \new_[78516]_  & \new_[78509]_ ;
  assign \new_[78520]_  = ~A267 & ~A266;
  assign \new_[78523]_  = A269 & ~A268;
  assign \new_[78524]_  = \new_[78523]_  & \new_[78520]_ ;
  assign \new_[78527]_  = A299 & ~A298;
  assign \new_[78530]_  = ~A302 & A300;
  assign \new_[78531]_  = \new_[78530]_  & \new_[78527]_ ;
  assign \new_[78532]_  = \new_[78531]_  & \new_[78524]_ ;
  assign \new_[78536]_  = ~A199 & A166;
  assign \new_[78537]_  = A167 & \new_[78536]_ ;
  assign \new_[78540]_  = ~A201 & A200;
  assign \new_[78543]_  = A203 & ~A202;
  assign \new_[78544]_  = \new_[78543]_  & \new_[78540]_ ;
  assign \new_[78545]_  = \new_[78544]_  & \new_[78537]_ ;
  assign \new_[78548]_  = A266 & ~A265;
  assign \new_[78551]_  = A268 & A267;
  assign \new_[78552]_  = \new_[78551]_  & \new_[78548]_ ;
  assign \new_[78555]_  = ~A299 & A298;
  assign \new_[78558]_  = A301 & A300;
  assign \new_[78559]_  = \new_[78558]_  & \new_[78555]_ ;
  assign \new_[78560]_  = \new_[78559]_  & \new_[78552]_ ;
  assign \new_[78564]_  = ~A199 & A166;
  assign \new_[78565]_  = A167 & \new_[78564]_ ;
  assign \new_[78568]_  = ~A201 & A200;
  assign \new_[78571]_  = A203 & ~A202;
  assign \new_[78572]_  = \new_[78571]_  & \new_[78568]_ ;
  assign \new_[78573]_  = \new_[78572]_  & \new_[78565]_ ;
  assign \new_[78576]_  = A266 & ~A265;
  assign \new_[78579]_  = A268 & A267;
  assign \new_[78580]_  = \new_[78579]_  & \new_[78576]_ ;
  assign \new_[78583]_  = ~A299 & A298;
  assign \new_[78586]_  = ~A302 & A300;
  assign \new_[78587]_  = \new_[78586]_  & \new_[78583]_ ;
  assign \new_[78588]_  = \new_[78587]_  & \new_[78580]_ ;
  assign \new_[78592]_  = ~A199 & A166;
  assign \new_[78593]_  = A167 & \new_[78592]_ ;
  assign \new_[78596]_  = ~A201 & A200;
  assign \new_[78599]_  = A203 & ~A202;
  assign \new_[78600]_  = \new_[78599]_  & \new_[78596]_ ;
  assign \new_[78601]_  = \new_[78600]_  & \new_[78593]_ ;
  assign \new_[78604]_  = A266 & ~A265;
  assign \new_[78607]_  = A268 & A267;
  assign \new_[78608]_  = \new_[78607]_  & \new_[78604]_ ;
  assign \new_[78611]_  = A299 & ~A298;
  assign \new_[78614]_  = A301 & A300;
  assign \new_[78615]_  = \new_[78614]_  & \new_[78611]_ ;
  assign \new_[78616]_  = \new_[78615]_  & \new_[78608]_ ;
  assign \new_[78620]_  = ~A199 & A166;
  assign \new_[78621]_  = A167 & \new_[78620]_ ;
  assign \new_[78624]_  = ~A201 & A200;
  assign \new_[78627]_  = A203 & ~A202;
  assign \new_[78628]_  = \new_[78627]_  & \new_[78624]_ ;
  assign \new_[78629]_  = \new_[78628]_  & \new_[78621]_ ;
  assign \new_[78632]_  = A266 & ~A265;
  assign \new_[78635]_  = A268 & A267;
  assign \new_[78636]_  = \new_[78635]_  & \new_[78632]_ ;
  assign \new_[78639]_  = A299 & ~A298;
  assign \new_[78642]_  = ~A302 & A300;
  assign \new_[78643]_  = \new_[78642]_  & \new_[78639]_ ;
  assign \new_[78644]_  = \new_[78643]_  & \new_[78636]_ ;
  assign \new_[78648]_  = ~A199 & A166;
  assign \new_[78649]_  = A167 & \new_[78648]_ ;
  assign \new_[78652]_  = ~A201 & A200;
  assign \new_[78655]_  = A203 & ~A202;
  assign \new_[78656]_  = \new_[78655]_  & \new_[78652]_ ;
  assign \new_[78657]_  = \new_[78656]_  & \new_[78649]_ ;
  assign \new_[78660]_  = A266 & ~A265;
  assign \new_[78663]_  = ~A269 & A267;
  assign \new_[78664]_  = \new_[78663]_  & \new_[78660]_ ;
  assign \new_[78667]_  = ~A299 & A298;
  assign \new_[78670]_  = A301 & A300;
  assign \new_[78671]_  = \new_[78670]_  & \new_[78667]_ ;
  assign \new_[78672]_  = \new_[78671]_  & \new_[78664]_ ;
  assign \new_[78676]_  = ~A199 & A166;
  assign \new_[78677]_  = A167 & \new_[78676]_ ;
  assign \new_[78680]_  = ~A201 & A200;
  assign \new_[78683]_  = A203 & ~A202;
  assign \new_[78684]_  = \new_[78683]_  & \new_[78680]_ ;
  assign \new_[78685]_  = \new_[78684]_  & \new_[78677]_ ;
  assign \new_[78688]_  = A266 & ~A265;
  assign \new_[78691]_  = ~A269 & A267;
  assign \new_[78692]_  = \new_[78691]_  & \new_[78688]_ ;
  assign \new_[78695]_  = ~A299 & A298;
  assign \new_[78698]_  = ~A302 & A300;
  assign \new_[78699]_  = \new_[78698]_  & \new_[78695]_ ;
  assign \new_[78700]_  = \new_[78699]_  & \new_[78692]_ ;
  assign \new_[78704]_  = ~A199 & A166;
  assign \new_[78705]_  = A167 & \new_[78704]_ ;
  assign \new_[78708]_  = ~A201 & A200;
  assign \new_[78711]_  = A203 & ~A202;
  assign \new_[78712]_  = \new_[78711]_  & \new_[78708]_ ;
  assign \new_[78713]_  = \new_[78712]_  & \new_[78705]_ ;
  assign \new_[78716]_  = A266 & ~A265;
  assign \new_[78719]_  = ~A269 & A267;
  assign \new_[78720]_  = \new_[78719]_  & \new_[78716]_ ;
  assign \new_[78723]_  = A299 & ~A298;
  assign \new_[78726]_  = A301 & A300;
  assign \new_[78727]_  = \new_[78726]_  & \new_[78723]_ ;
  assign \new_[78728]_  = \new_[78727]_  & \new_[78720]_ ;
  assign \new_[78732]_  = ~A199 & A166;
  assign \new_[78733]_  = A167 & \new_[78732]_ ;
  assign \new_[78736]_  = ~A201 & A200;
  assign \new_[78739]_  = A203 & ~A202;
  assign \new_[78740]_  = \new_[78739]_  & \new_[78736]_ ;
  assign \new_[78741]_  = \new_[78740]_  & \new_[78733]_ ;
  assign \new_[78744]_  = A266 & ~A265;
  assign \new_[78747]_  = ~A269 & A267;
  assign \new_[78748]_  = \new_[78747]_  & \new_[78744]_ ;
  assign \new_[78751]_  = A299 & ~A298;
  assign \new_[78754]_  = ~A302 & A300;
  assign \new_[78755]_  = \new_[78754]_  & \new_[78751]_ ;
  assign \new_[78756]_  = \new_[78755]_  & \new_[78748]_ ;
  assign \new_[78760]_  = ~A199 & A166;
  assign \new_[78761]_  = A167 & \new_[78760]_ ;
  assign \new_[78764]_  = ~A201 & A200;
  assign \new_[78767]_  = A203 & ~A202;
  assign \new_[78768]_  = \new_[78767]_  & \new_[78764]_ ;
  assign \new_[78769]_  = \new_[78768]_  & \new_[78761]_ ;
  assign \new_[78772]_  = ~A266 & A265;
  assign \new_[78775]_  = A268 & A267;
  assign \new_[78776]_  = \new_[78775]_  & \new_[78772]_ ;
  assign \new_[78779]_  = ~A299 & A298;
  assign \new_[78782]_  = A301 & A300;
  assign \new_[78783]_  = \new_[78782]_  & \new_[78779]_ ;
  assign \new_[78784]_  = \new_[78783]_  & \new_[78776]_ ;
  assign \new_[78788]_  = ~A199 & A166;
  assign \new_[78789]_  = A167 & \new_[78788]_ ;
  assign \new_[78792]_  = ~A201 & A200;
  assign \new_[78795]_  = A203 & ~A202;
  assign \new_[78796]_  = \new_[78795]_  & \new_[78792]_ ;
  assign \new_[78797]_  = \new_[78796]_  & \new_[78789]_ ;
  assign \new_[78800]_  = ~A266 & A265;
  assign \new_[78803]_  = A268 & A267;
  assign \new_[78804]_  = \new_[78803]_  & \new_[78800]_ ;
  assign \new_[78807]_  = ~A299 & A298;
  assign \new_[78810]_  = ~A302 & A300;
  assign \new_[78811]_  = \new_[78810]_  & \new_[78807]_ ;
  assign \new_[78812]_  = \new_[78811]_  & \new_[78804]_ ;
  assign \new_[78816]_  = ~A199 & A166;
  assign \new_[78817]_  = A167 & \new_[78816]_ ;
  assign \new_[78820]_  = ~A201 & A200;
  assign \new_[78823]_  = A203 & ~A202;
  assign \new_[78824]_  = \new_[78823]_  & \new_[78820]_ ;
  assign \new_[78825]_  = \new_[78824]_  & \new_[78817]_ ;
  assign \new_[78828]_  = ~A266 & A265;
  assign \new_[78831]_  = A268 & A267;
  assign \new_[78832]_  = \new_[78831]_  & \new_[78828]_ ;
  assign \new_[78835]_  = A299 & ~A298;
  assign \new_[78838]_  = A301 & A300;
  assign \new_[78839]_  = \new_[78838]_  & \new_[78835]_ ;
  assign \new_[78840]_  = \new_[78839]_  & \new_[78832]_ ;
  assign \new_[78844]_  = ~A199 & A166;
  assign \new_[78845]_  = A167 & \new_[78844]_ ;
  assign \new_[78848]_  = ~A201 & A200;
  assign \new_[78851]_  = A203 & ~A202;
  assign \new_[78852]_  = \new_[78851]_  & \new_[78848]_ ;
  assign \new_[78853]_  = \new_[78852]_  & \new_[78845]_ ;
  assign \new_[78856]_  = ~A266 & A265;
  assign \new_[78859]_  = A268 & A267;
  assign \new_[78860]_  = \new_[78859]_  & \new_[78856]_ ;
  assign \new_[78863]_  = A299 & ~A298;
  assign \new_[78866]_  = ~A302 & A300;
  assign \new_[78867]_  = \new_[78866]_  & \new_[78863]_ ;
  assign \new_[78868]_  = \new_[78867]_  & \new_[78860]_ ;
  assign \new_[78872]_  = ~A199 & A166;
  assign \new_[78873]_  = A167 & \new_[78872]_ ;
  assign \new_[78876]_  = ~A201 & A200;
  assign \new_[78879]_  = A203 & ~A202;
  assign \new_[78880]_  = \new_[78879]_  & \new_[78876]_ ;
  assign \new_[78881]_  = \new_[78880]_  & \new_[78873]_ ;
  assign \new_[78884]_  = ~A266 & A265;
  assign \new_[78887]_  = ~A269 & A267;
  assign \new_[78888]_  = \new_[78887]_  & \new_[78884]_ ;
  assign \new_[78891]_  = ~A299 & A298;
  assign \new_[78894]_  = A301 & A300;
  assign \new_[78895]_  = \new_[78894]_  & \new_[78891]_ ;
  assign \new_[78896]_  = \new_[78895]_  & \new_[78888]_ ;
  assign \new_[78900]_  = ~A199 & A166;
  assign \new_[78901]_  = A167 & \new_[78900]_ ;
  assign \new_[78904]_  = ~A201 & A200;
  assign \new_[78907]_  = A203 & ~A202;
  assign \new_[78908]_  = \new_[78907]_  & \new_[78904]_ ;
  assign \new_[78909]_  = \new_[78908]_  & \new_[78901]_ ;
  assign \new_[78912]_  = ~A266 & A265;
  assign \new_[78915]_  = ~A269 & A267;
  assign \new_[78916]_  = \new_[78915]_  & \new_[78912]_ ;
  assign \new_[78919]_  = ~A299 & A298;
  assign \new_[78922]_  = ~A302 & A300;
  assign \new_[78923]_  = \new_[78922]_  & \new_[78919]_ ;
  assign \new_[78924]_  = \new_[78923]_  & \new_[78916]_ ;
  assign \new_[78928]_  = ~A199 & A166;
  assign \new_[78929]_  = A167 & \new_[78928]_ ;
  assign \new_[78932]_  = ~A201 & A200;
  assign \new_[78935]_  = A203 & ~A202;
  assign \new_[78936]_  = \new_[78935]_  & \new_[78932]_ ;
  assign \new_[78937]_  = \new_[78936]_  & \new_[78929]_ ;
  assign \new_[78940]_  = ~A266 & A265;
  assign \new_[78943]_  = ~A269 & A267;
  assign \new_[78944]_  = \new_[78943]_  & \new_[78940]_ ;
  assign \new_[78947]_  = A299 & ~A298;
  assign \new_[78950]_  = A301 & A300;
  assign \new_[78951]_  = \new_[78950]_  & \new_[78947]_ ;
  assign \new_[78952]_  = \new_[78951]_  & \new_[78944]_ ;
  assign \new_[78956]_  = ~A199 & A166;
  assign \new_[78957]_  = A167 & \new_[78956]_ ;
  assign \new_[78960]_  = ~A201 & A200;
  assign \new_[78963]_  = A203 & ~A202;
  assign \new_[78964]_  = \new_[78963]_  & \new_[78960]_ ;
  assign \new_[78965]_  = \new_[78964]_  & \new_[78957]_ ;
  assign \new_[78968]_  = ~A266 & A265;
  assign \new_[78971]_  = ~A269 & A267;
  assign \new_[78972]_  = \new_[78971]_  & \new_[78968]_ ;
  assign \new_[78975]_  = A299 & ~A298;
  assign \new_[78978]_  = ~A302 & A300;
  assign \new_[78979]_  = \new_[78978]_  & \new_[78975]_ ;
  assign \new_[78980]_  = \new_[78979]_  & \new_[78972]_ ;
  assign \new_[78984]_  = A199 & A166;
  assign \new_[78985]_  = A167 & \new_[78984]_ ;
  assign \new_[78988]_  = A201 & ~A200;
  assign \new_[78991]_  = ~A265 & A202;
  assign \new_[78992]_  = \new_[78991]_  & \new_[78988]_ ;
  assign \new_[78993]_  = \new_[78992]_  & \new_[78985]_ ;
  assign \new_[78996]_  = A267 & A266;
  assign \new_[78999]_  = A298 & A268;
  assign \new_[79000]_  = \new_[78999]_  & \new_[78996]_ ;
  assign \new_[79003]_  = ~A300 & ~A299;
  assign \new_[79006]_  = A302 & ~A301;
  assign \new_[79007]_  = \new_[79006]_  & \new_[79003]_ ;
  assign \new_[79008]_  = \new_[79007]_  & \new_[79000]_ ;
  assign \new_[79012]_  = A199 & A166;
  assign \new_[79013]_  = A167 & \new_[79012]_ ;
  assign \new_[79016]_  = A201 & ~A200;
  assign \new_[79019]_  = ~A265 & A202;
  assign \new_[79020]_  = \new_[79019]_  & \new_[79016]_ ;
  assign \new_[79021]_  = \new_[79020]_  & \new_[79013]_ ;
  assign \new_[79024]_  = A267 & A266;
  assign \new_[79027]_  = ~A298 & A268;
  assign \new_[79028]_  = \new_[79027]_  & \new_[79024]_ ;
  assign \new_[79031]_  = ~A300 & A299;
  assign \new_[79034]_  = A302 & ~A301;
  assign \new_[79035]_  = \new_[79034]_  & \new_[79031]_ ;
  assign \new_[79036]_  = \new_[79035]_  & \new_[79028]_ ;
  assign \new_[79040]_  = A199 & A166;
  assign \new_[79041]_  = A167 & \new_[79040]_ ;
  assign \new_[79044]_  = A201 & ~A200;
  assign \new_[79047]_  = ~A265 & A202;
  assign \new_[79048]_  = \new_[79047]_  & \new_[79044]_ ;
  assign \new_[79049]_  = \new_[79048]_  & \new_[79041]_ ;
  assign \new_[79052]_  = A267 & A266;
  assign \new_[79055]_  = A298 & ~A269;
  assign \new_[79056]_  = \new_[79055]_  & \new_[79052]_ ;
  assign \new_[79059]_  = ~A300 & ~A299;
  assign \new_[79062]_  = A302 & ~A301;
  assign \new_[79063]_  = \new_[79062]_  & \new_[79059]_ ;
  assign \new_[79064]_  = \new_[79063]_  & \new_[79056]_ ;
  assign \new_[79068]_  = A199 & A166;
  assign \new_[79069]_  = A167 & \new_[79068]_ ;
  assign \new_[79072]_  = A201 & ~A200;
  assign \new_[79075]_  = ~A265 & A202;
  assign \new_[79076]_  = \new_[79075]_  & \new_[79072]_ ;
  assign \new_[79077]_  = \new_[79076]_  & \new_[79069]_ ;
  assign \new_[79080]_  = A267 & A266;
  assign \new_[79083]_  = ~A298 & ~A269;
  assign \new_[79084]_  = \new_[79083]_  & \new_[79080]_ ;
  assign \new_[79087]_  = ~A300 & A299;
  assign \new_[79090]_  = A302 & ~A301;
  assign \new_[79091]_  = \new_[79090]_  & \new_[79087]_ ;
  assign \new_[79092]_  = \new_[79091]_  & \new_[79084]_ ;
  assign \new_[79096]_  = A199 & A166;
  assign \new_[79097]_  = A167 & \new_[79096]_ ;
  assign \new_[79100]_  = A201 & ~A200;
  assign \new_[79103]_  = ~A265 & A202;
  assign \new_[79104]_  = \new_[79103]_  & \new_[79100]_ ;
  assign \new_[79105]_  = \new_[79104]_  & \new_[79097]_ ;
  assign \new_[79108]_  = ~A267 & A266;
  assign \new_[79111]_  = A269 & ~A268;
  assign \new_[79112]_  = \new_[79111]_  & \new_[79108]_ ;
  assign \new_[79115]_  = ~A299 & A298;
  assign \new_[79118]_  = A301 & A300;
  assign \new_[79119]_  = \new_[79118]_  & \new_[79115]_ ;
  assign \new_[79120]_  = \new_[79119]_  & \new_[79112]_ ;
  assign \new_[79124]_  = A199 & A166;
  assign \new_[79125]_  = A167 & \new_[79124]_ ;
  assign \new_[79128]_  = A201 & ~A200;
  assign \new_[79131]_  = ~A265 & A202;
  assign \new_[79132]_  = \new_[79131]_  & \new_[79128]_ ;
  assign \new_[79133]_  = \new_[79132]_  & \new_[79125]_ ;
  assign \new_[79136]_  = ~A267 & A266;
  assign \new_[79139]_  = A269 & ~A268;
  assign \new_[79140]_  = \new_[79139]_  & \new_[79136]_ ;
  assign \new_[79143]_  = ~A299 & A298;
  assign \new_[79146]_  = ~A302 & A300;
  assign \new_[79147]_  = \new_[79146]_  & \new_[79143]_ ;
  assign \new_[79148]_  = \new_[79147]_  & \new_[79140]_ ;
  assign \new_[79152]_  = A199 & A166;
  assign \new_[79153]_  = A167 & \new_[79152]_ ;
  assign \new_[79156]_  = A201 & ~A200;
  assign \new_[79159]_  = ~A265 & A202;
  assign \new_[79160]_  = \new_[79159]_  & \new_[79156]_ ;
  assign \new_[79161]_  = \new_[79160]_  & \new_[79153]_ ;
  assign \new_[79164]_  = ~A267 & A266;
  assign \new_[79167]_  = A269 & ~A268;
  assign \new_[79168]_  = \new_[79167]_  & \new_[79164]_ ;
  assign \new_[79171]_  = A299 & ~A298;
  assign \new_[79174]_  = A301 & A300;
  assign \new_[79175]_  = \new_[79174]_  & \new_[79171]_ ;
  assign \new_[79176]_  = \new_[79175]_  & \new_[79168]_ ;
  assign \new_[79180]_  = A199 & A166;
  assign \new_[79181]_  = A167 & \new_[79180]_ ;
  assign \new_[79184]_  = A201 & ~A200;
  assign \new_[79187]_  = ~A265 & A202;
  assign \new_[79188]_  = \new_[79187]_  & \new_[79184]_ ;
  assign \new_[79189]_  = \new_[79188]_  & \new_[79181]_ ;
  assign \new_[79192]_  = ~A267 & A266;
  assign \new_[79195]_  = A269 & ~A268;
  assign \new_[79196]_  = \new_[79195]_  & \new_[79192]_ ;
  assign \new_[79199]_  = A299 & ~A298;
  assign \new_[79202]_  = ~A302 & A300;
  assign \new_[79203]_  = \new_[79202]_  & \new_[79199]_ ;
  assign \new_[79204]_  = \new_[79203]_  & \new_[79196]_ ;
  assign \new_[79208]_  = A199 & A166;
  assign \new_[79209]_  = A167 & \new_[79208]_ ;
  assign \new_[79212]_  = A201 & ~A200;
  assign \new_[79215]_  = A265 & A202;
  assign \new_[79216]_  = \new_[79215]_  & \new_[79212]_ ;
  assign \new_[79217]_  = \new_[79216]_  & \new_[79209]_ ;
  assign \new_[79220]_  = A267 & ~A266;
  assign \new_[79223]_  = A298 & A268;
  assign \new_[79224]_  = \new_[79223]_  & \new_[79220]_ ;
  assign \new_[79227]_  = ~A300 & ~A299;
  assign \new_[79230]_  = A302 & ~A301;
  assign \new_[79231]_  = \new_[79230]_  & \new_[79227]_ ;
  assign \new_[79232]_  = \new_[79231]_  & \new_[79224]_ ;
  assign \new_[79236]_  = A199 & A166;
  assign \new_[79237]_  = A167 & \new_[79236]_ ;
  assign \new_[79240]_  = A201 & ~A200;
  assign \new_[79243]_  = A265 & A202;
  assign \new_[79244]_  = \new_[79243]_  & \new_[79240]_ ;
  assign \new_[79245]_  = \new_[79244]_  & \new_[79237]_ ;
  assign \new_[79248]_  = A267 & ~A266;
  assign \new_[79251]_  = ~A298 & A268;
  assign \new_[79252]_  = \new_[79251]_  & \new_[79248]_ ;
  assign \new_[79255]_  = ~A300 & A299;
  assign \new_[79258]_  = A302 & ~A301;
  assign \new_[79259]_  = \new_[79258]_  & \new_[79255]_ ;
  assign \new_[79260]_  = \new_[79259]_  & \new_[79252]_ ;
  assign \new_[79264]_  = A199 & A166;
  assign \new_[79265]_  = A167 & \new_[79264]_ ;
  assign \new_[79268]_  = A201 & ~A200;
  assign \new_[79271]_  = A265 & A202;
  assign \new_[79272]_  = \new_[79271]_  & \new_[79268]_ ;
  assign \new_[79273]_  = \new_[79272]_  & \new_[79265]_ ;
  assign \new_[79276]_  = A267 & ~A266;
  assign \new_[79279]_  = A298 & ~A269;
  assign \new_[79280]_  = \new_[79279]_  & \new_[79276]_ ;
  assign \new_[79283]_  = ~A300 & ~A299;
  assign \new_[79286]_  = A302 & ~A301;
  assign \new_[79287]_  = \new_[79286]_  & \new_[79283]_ ;
  assign \new_[79288]_  = \new_[79287]_  & \new_[79280]_ ;
  assign \new_[79292]_  = A199 & A166;
  assign \new_[79293]_  = A167 & \new_[79292]_ ;
  assign \new_[79296]_  = A201 & ~A200;
  assign \new_[79299]_  = A265 & A202;
  assign \new_[79300]_  = \new_[79299]_  & \new_[79296]_ ;
  assign \new_[79301]_  = \new_[79300]_  & \new_[79293]_ ;
  assign \new_[79304]_  = A267 & ~A266;
  assign \new_[79307]_  = ~A298 & ~A269;
  assign \new_[79308]_  = \new_[79307]_  & \new_[79304]_ ;
  assign \new_[79311]_  = ~A300 & A299;
  assign \new_[79314]_  = A302 & ~A301;
  assign \new_[79315]_  = \new_[79314]_  & \new_[79311]_ ;
  assign \new_[79316]_  = \new_[79315]_  & \new_[79308]_ ;
  assign \new_[79320]_  = A199 & A166;
  assign \new_[79321]_  = A167 & \new_[79320]_ ;
  assign \new_[79324]_  = A201 & ~A200;
  assign \new_[79327]_  = A265 & A202;
  assign \new_[79328]_  = \new_[79327]_  & \new_[79324]_ ;
  assign \new_[79329]_  = \new_[79328]_  & \new_[79321]_ ;
  assign \new_[79332]_  = ~A267 & ~A266;
  assign \new_[79335]_  = A269 & ~A268;
  assign \new_[79336]_  = \new_[79335]_  & \new_[79332]_ ;
  assign \new_[79339]_  = ~A299 & A298;
  assign \new_[79342]_  = A301 & A300;
  assign \new_[79343]_  = \new_[79342]_  & \new_[79339]_ ;
  assign \new_[79344]_  = \new_[79343]_  & \new_[79336]_ ;
  assign \new_[79348]_  = A199 & A166;
  assign \new_[79349]_  = A167 & \new_[79348]_ ;
  assign \new_[79352]_  = A201 & ~A200;
  assign \new_[79355]_  = A265 & A202;
  assign \new_[79356]_  = \new_[79355]_  & \new_[79352]_ ;
  assign \new_[79357]_  = \new_[79356]_  & \new_[79349]_ ;
  assign \new_[79360]_  = ~A267 & ~A266;
  assign \new_[79363]_  = A269 & ~A268;
  assign \new_[79364]_  = \new_[79363]_  & \new_[79360]_ ;
  assign \new_[79367]_  = ~A299 & A298;
  assign \new_[79370]_  = ~A302 & A300;
  assign \new_[79371]_  = \new_[79370]_  & \new_[79367]_ ;
  assign \new_[79372]_  = \new_[79371]_  & \new_[79364]_ ;
  assign \new_[79376]_  = A199 & A166;
  assign \new_[79377]_  = A167 & \new_[79376]_ ;
  assign \new_[79380]_  = A201 & ~A200;
  assign \new_[79383]_  = A265 & A202;
  assign \new_[79384]_  = \new_[79383]_  & \new_[79380]_ ;
  assign \new_[79385]_  = \new_[79384]_  & \new_[79377]_ ;
  assign \new_[79388]_  = ~A267 & ~A266;
  assign \new_[79391]_  = A269 & ~A268;
  assign \new_[79392]_  = \new_[79391]_  & \new_[79388]_ ;
  assign \new_[79395]_  = A299 & ~A298;
  assign \new_[79398]_  = A301 & A300;
  assign \new_[79399]_  = \new_[79398]_  & \new_[79395]_ ;
  assign \new_[79400]_  = \new_[79399]_  & \new_[79392]_ ;
  assign \new_[79404]_  = A199 & A166;
  assign \new_[79405]_  = A167 & \new_[79404]_ ;
  assign \new_[79408]_  = A201 & ~A200;
  assign \new_[79411]_  = A265 & A202;
  assign \new_[79412]_  = \new_[79411]_  & \new_[79408]_ ;
  assign \new_[79413]_  = \new_[79412]_  & \new_[79405]_ ;
  assign \new_[79416]_  = ~A267 & ~A266;
  assign \new_[79419]_  = A269 & ~A268;
  assign \new_[79420]_  = \new_[79419]_  & \new_[79416]_ ;
  assign \new_[79423]_  = A299 & ~A298;
  assign \new_[79426]_  = ~A302 & A300;
  assign \new_[79427]_  = \new_[79426]_  & \new_[79423]_ ;
  assign \new_[79428]_  = \new_[79427]_  & \new_[79420]_ ;
  assign \new_[79432]_  = A199 & A166;
  assign \new_[79433]_  = A167 & \new_[79432]_ ;
  assign \new_[79436]_  = A201 & ~A200;
  assign \new_[79439]_  = ~A265 & ~A203;
  assign \new_[79440]_  = \new_[79439]_  & \new_[79436]_ ;
  assign \new_[79441]_  = \new_[79440]_  & \new_[79433]_ ;
  assign \new_[79444]_  = A267 & A266;
  assign \new_[79447]_  = A298 & A268;
  assign \new_[79448]_  = \new_[79447]_  & \new_[79444]_ ;
  assign \new_[79451]_  = ~A300 & ~A299;
  assign \new_[79454]_  = A302 & ~A301;
  assign \new_[79455]_  = \new_[79454]_  & \new_[79451]_ ;
  assign \new_[79456]_  = \new_[79455]_  & \new_[79448]_ ;
  assign \new_[79460]_  = A199 & A166;
  assign \new_[79461]_  = A167 & \new_[79460]_ ;
  assign \new_[79464]_  = A201 & ~A200;
  assign \new_[79467]_  = ~A265 & ~A203;
  assign \new_[79468]_  = \new_[79467]_  & \new_[79464]_ ;
  assign \new_[79469]_  = \new_[79468]_  & \new_[79461]_ ;
  assign \new_[79472]_  = A267 & A266;
  assign \new_[79475]_  = ~A298 & A268;
  assign \new_[79476]_  = \new_[79475]_  & \new_[79472]_ ;
  assign \new_[79479]_  = ~A300 & A299;
  assign \new_[79482]_  = A302 & ~A301;
  assign \new_[79483]_  = \new_[79482]_  & \new_[79479]_ ;
  assign \new_[79484]_  = \new_[79483]_  & \new_[79476]_ ;
  assign \new_[79488]_  = A199 & A166;
  assign \new_[79489]_  = A167 & \new_[79488]_ ;
  assign \new_[79492]_  = A201 & ~A200;
  assign \new_[79495]_  = ~A265 & ~A203;
  assign \new_[79496]_  = \new_[79495]_  & \new_[79492]_ ;
  assign \new_[79497]_  = \new_[79496]_  & \new_[79489]_ ;
  assign \new_[79500]_  = A267 & A266;
  assign \new_[79503]_  = A298 & ~A269;
  assign \new_[79504]_  = \new_[79503]_  & \new_[79500]_ ;
  assign \new_[79507]_  = ~A300 & ~A299;
  assign \new_[79510]_  = A302 & ~A301;
  assign \new_[79511]_  = \new_[79510]_  & \new_[79507]_ ;
  assign \new_[79512]_  = \new_[79511]_  & \new_[79504]_ ;
  assign \new_[79516]_  = A199 & A166;
  assign \new_[79517]_  = A167 & \new_[79516]_ ;
  assign \new_[79520]_  = A201 & ~A200;
  assign \new_[79523]_  = ~A265 & ~A203;
  assign \new_[79524]_  = \new_[79523]_  & \new_[79520]_ ;
  assign \new_[79525]_  = \new_[79524]_  & \new_[79517]_ ;
  assign \new_[79528]_  = A267 & A266;
  assign \new_[79531]_  = ~A298 & ~A269;
  assign \new_[79532]_  = \new_[79531]_  & \new_[79528]_ ;
  assign \new_[79535]_  = ~A300 & A299;
  assign \new_[79538]_  = A302 & ~A301;
  assign \new_[79539]_  = \new_[79538]_  & \new_[79535]_ ;
  assign \new_[79540]_  = \new_[79539]_  & \new_[79532]_ ;
  assign \new_[79544]_  = A199 & A166;
  assign \new_[79545]_  = A167 & \new_[79544]_ ;
  assign \new_[79548]_  = A201 & ~A200;
  assign \new_[79551]_  = ~A265 & ~A203;
  assign \new_[79552]_  = \new_[79551]_  & \new_[79548]_ ;
  assign \new_[79553]_  = \new_[79552]_  & \new_[79545]_ ;
  assign \new_[79556]_  = ~A267 & A266;
  assign \new_[79559]_  = A269 & ~A268;
  assign \new_[79560]_  = \new_[79559]_  & \new_[79556]_ ;
  assign \new_[79563]_  = ~A299 & A298;
  assign \new_[79566]_  = A301 & A300;
  assign \new_[79567]_  = \new_[79566]_  & \new_[79563]_ ;
  assign \new_[79568]_  = \new_[79567]_  & \new_[79560]_ ;
  assign \new_[79572]_  = A199 & A166;
  assign \new_[79573]_  = A167 & \new_[79572]_ ;
  assign \new_[79576]_  = A201 & ~A200;
  assign \new_[79579]_  = ~A265 & ~A203;
  assign \new_[79580]_  = \new_[79579]_  & \new_[79576]_ ;
  assign \new_[79581]_  = \new_[79580]_  & \new_[79573]_ ;
  assign \new_[79584]_  = ~A267 & A266;
  assign \new_[79587]_  = A269 & ~A268;
  assign \new_[79588]_  = \new_[79587]_  & \new_[79584]_ ;
  assign \new_[79591]_  = ~A299 & A298;
  assign \new_[79594]_  = ~A302 & A300;
  assign \new_[79595]_  = \new_[79594]_  & \new_[79591]_ ;
  assign \new_[79596]_  = \new_[79595]_  & \new_[79588]_ ;
  assign \new_[79600]_  = A199 & A166;
  assign \new_[79601]_  = A167 & \new_[79600]_ ;
  assign \new_[79604]_  = A201 & ~A200;
  assign \new_[79607]_  = ~A265 & ~A203;
  assign \new_[79608]_  = \new_[79607]_  & \new_[79604]_ ;
  assign \new_[79609]_  = \new_[79608]_  & \new_[79601]_ ;
  assign \new_[79612]_  = ~A267 & A266;
  assign \new_[79615]_  = A269 & ~A268;
  assign \new_[79616]_  = \new_[79615]_  & \new_[79612]_ ;
  assign \new_[79619]_  = A299 & ~A298;
  assign \new_[79622]_  = A301 & A300;
  assign \new_[79623]_  = \new_[79622]_  & \new_[79619]_ ;
  assign \new_[79624]_  = \new_[79623]_  & \new_[79616]_ ;
  assign \new_[79628]_  = A199 & A166;
  assign \new_[79629]_  = A167 & \new_[79628]_ ;
  assign \new_[79632]_  = A201 & ~A200;
  assign \new_[79635]_  = ~A265 & ~A203;
  assign \new_[79636]_  = \new_[79635]_  & \new_[79632]_ ;
  assign \new_[79637]_  = \new_[79636]_  & \new_[79629]_ ;
  assign \new_[79640]_  = ~A267 & A266;
  assign \new_[79643]_  = A269 & ~A268;
  assign \new_[79644]_  = \new_[79643]_  & \new_[79640]_ ;
  assign \new_[79647]_  = A299 & ~A298;
  assign \new_[79650]_  = ~A302 & A300;
  assign \new_[79651]_  = \new_[79650]_  & \new_[79647]_ ;
  assign \new_[79652]_  = \new_[79651]_  & \new_[79644]_ ;
  assign \new_[79656]_  = A199 & A166;
  assign \new_[79657]_  = A167 & \new_[79656]_ ;
  assign \new_[79660]_  = A201 & ~A200;
  assign \new_[79663]_  = A265 & ~A203;
  assign \new_[79664]_  = \new_[79663]_  & \new_[79660]_ ;
  assign \new_[79665]_  = \new_[79664]_  & \new_[79657]_ ;
  assign \new_[79668]_  = A267 & ~A266;
  assign \new_[79671]_  = A298 & A268;
  assign \new_[79672]_  = \new_[79671]_  & \new_[79668]_ ;
  assign \new_[79675]_  = ~A300 & ~A299;
  assign \new_[79678]_  = A302 & ~A301;
  assign \new_[79679]_  = \new_[79678]_  & \new_[79675]_ ;
  assign \new_[79680]_  = \new_[79679]_  & \new_[79672]_ ;
  assign \new_[79684]_  = A199 & A166;
  assign \new_[79685]_  = A167 & \new_[79684]_ ;
  assign \new_[79688]_  = A201 & ~A200;
  assign \new_[79691]_  = A265 & ~A203;
  assign \new_[79692]_  = \new_[79691]_  & \new_[79688]_ ;
  assign \new_[79693]_  = \new_[79692]_  & \new_[79685]_ ;
  assign \new_[79696]_  = A267 & ~A266;
  assign \new_[79699]_  = ~A298 & A268;
  assign \new_[79700]_  = \new_[79699]_  & \new_[79696]_ ;
  assign \new_[79703]_  = ~A300 & A299;
  assign \new_[79706]_  = A302 & ~A301;
  assign \new_[79707]_  = \new_[79706]_  & \new_[79703]_ ;
  assign \new_[79708]_  = \new_[79707]_  & \new_[79700]_ ;
  assign \new_[79712]_  = A199 & A166;
  assign \new_[79713]_  = A167 & \new_[79712]_ ;
  assign \new_[79716]_  = A201 & ~A200;
  assign \new_[79719]_  = A265 & ~A203;
  assign \new_[79720]_  = \new_[79719]_  & \new_[79716]_ ;
  assign \new_[79721]_  = \new_[79720]_  & \new_[79713]_ ;
  assign \new_[79724]_  = A267 & ~A266;
  assign \new_[79727]_  = A298 & ~A269;
  assign \new_[79728]_  = \new_[79727]_  & \new_[79724]_ ;
  assign \new_[79731]_  = ~A300 & ~A299;
  assign \new_[79734]_  = A302 & ~A301;
  assign \new_[79735]_  = \new_[79734]_  & \new_[79731]_ ;
  assign \new_[79736]_  = \new_[79735]_  & \new_[79728]_ ;
  assign \new_[79740]_  = A199 & A166;
  assign \new_[79741]_  = A167 & \new_[79740]_ ;
  assign \new_[79744]_  = A201 & ~A200;
  assign \new_[79747]_  = A265 & ~A203;
  assign \new_[79748]_  = \new_[79747]_  & \new_[79744]_ ;
  assign \new_[79749]_  = \new_[79748]_  & \new_[79741]_ ;
  assign \new_[79752]_  = A267 & ~A266;
  assign \new_[79755]_  = ~A298 & ~A269;
  assign \new_[79756]_  = \new_[79755]_  & \new_[79752]_ ;
  assign \new_[79759]_  = ~A300 & A299;
  assign \new_[79762]_  = A302 & ~A301;
  assign \new_[79763]_  = \new_[79762]_  & \new_[79759]_ ;
  assign \new_[79764]_  = \new_[79763]_  & \new_[79756]_ ;
  assign \new_[79768]_  = A199 & A166;
  assign \new_[79769]_  = A167 & \new_[79768]_ ;
  assign \new_[79772]_  = A201 & ~A200;
  assign \new_[79775]_  = A265 & ~A203;
  assign \new_[79776]_  = \new_[79775]_  & \new_[79772]_ ;
  assign \new_[79777]_  = \new_[79776]_  & \new_[79769]_ ;
  assign \new_[79780]_  = ~A267 & ~A266;
  assign \new_[79783]_  = A269 & ~A268;
  assign \new_[79784]_  = \new_[79783]_  & \new_[79780]_ ;
  assign \new_[79787]_  = ~A299 & A298;
  assign \new_[79790]_  = A301 & A300;
  assign \new_[79791]_  = \new_[79790]_  & \new_[79787]_ ;
  assign \new_[79792]_  = \new_[79791]_  & \new_[79784]_ ;
  assign \new_[79796]_  = A199 & A166;
  assign \new_[79797]_  = A167 & \new_[79796]_ ;
  assign \new_[79800]_  = A201 & ~A200;
  assign \new_[79803]_  = A265 & ~A203;
  assign \new_[79804]_  = \new_[79803]_  & \new_[79800]_ ;
  assign \new_[79805]_  = \new_[79804]_  & \new_[79797]_ ;
  assign \new_[79808]_  = ~A267 & ~A266;
  assign \new_[79811]_  = A269 & ~A268;
  assign \new_[79812]_  = \new_[79811]_  & \new_[79808]_ ;
  assign \new_[79815]_  = ~A299 & A298;
  assign \new_[79818]_  = ~A302 & A300;
  assign \new_[79819]_  = \new_[79818]_  & \new_[79815]_ ;
  assign \new_[79820]_  = \new_[79819]_  & \new_[79812]_ ;
  assign \new_[79824]_  = A199 & A166;
  assign \new_[79825]_  = A167 & \new_[79824]_ ;
  assign \new_[79828]_  = A201 & ~A200;
  assign \new_[79831]_  = A265 & ~A203;
  assign \new_[79832]_  = \new_[79831]_  & \new_[79828]_ ;
  assign \new_[79833]_  = \new_[79832]_  & \new_[79825]_ ;
  assign \new_[79836]_  = ~A267 & ~A266;
  assign \new_[79839]_  = A269 & ~A268;
  assign \new_[79840]_  = \new_[79839]_  & \new_[79836]_ ;
  assign \new_[79843]_  = A299 & ~A298;
  assign \new_[79846]_  = A301 & A300;
  assign \new_[79847]_  = \new_[79846]_  & \new_[79843]_ ;
  assign \new_[79848]_  = \new_[79847]_  & \new_[79840]_ ;
  assign \new_[79852]_  = A199 & A166;
  assign \new_[79853]_  = A167 & \new_[79852]_ ;
  assign \new_[79856]_  = A201 & ~A200;
  assign \new_[79859]_  = A265 & ~A203;
  assign \new_[79860]_  = \new_[79859]_  & \new_[79856]_ ;
  assign \new_[79861]_  = \new_[79860]_  & \new_[79853]_ ;
  assign \new_[79864]_  = ~A267 & ~A266;
  assign \new_[79867]_  = A269 & ~A268;
  assign \new_[79868]_  = \new_[79867]_  & \new_[79864]_ ;
  assign \new_[79871]_  = A299 & ~A298;
  assign \new_[79874]_  = ~A302 & A300;
  assign \new_[79875]_  = \new_[79874]_  & \new_[79871]_ ;
  assign \new_[79876]_  = \new_[79875]_  & \new_[79868]_ ;
  assign \new_[79880]_  = A199 & A166;
  assign \new_[79881]_  = A167 & \new_[79880]_ ;
  assign \new_[79884]_  = ~A201 & ~A200;
  assign \new_[79887]_  = A203 & ~A202;
  assign \new_[79888]_  = \new_[79887]_  & \new_[79884]_ ;
  assign \new_[79889]_  = \new_[79888]_  & \new_[79881]_ ;
  assign \new_[79892]_  = A266 & ~A265;
  assign \new_[79895]_  = A268 & A267;
  assign \new_[79896]_  = \new_[79895]_  & \new_[79892]_ ;
  assign \new_[79899]_  = ~A299 & A298;
  assign \new_[79902]_  = A301 & A300;
  assign \new_[79903]_  = \new_[79902]_  & \new_[79899]_ ;
  assign \new_[79904]_  = \new_[79903]_  & \new_[79896]_ ;
  assign \new_[79908]_  = A199 & A166;
  assign \new_[79909]_  = A167 & \new_[79908]_ ;
  assign \new_[79912]_  = ~A201 & ~A200;
  assign \new_[79915]_  = A203 & ~A202;
  assign \new_[79916]_  = \new_[79915]_  & \new_[79912]_ ;
  assign \new_[79917]_  = \new_[79916]_  & \new_[79909]_ ;
  assign \new_[79920]_  = A266 & ~A265;
  assign \new_[79923]_  = A268 & A267;
  assign \new_[79924]_  = \new_[79923]_  & \new_[79920]_ ;
  assign \new_[79927]_  = ~A299 & A298;
  assign \new_[79930]_  = ~A302 & A300;
  assign \new_[79931]_  = \new_[79930]_  & \new_[79927]_ ;
  assign \new_[79932]_  = \new_[79931]_  & \new_[79924]_ ;
  assign \new_[79936]_  = A199 & A166;
  assign \new_[79937]_  = A167 & \new_[79936]_ ;
  assign \new_[79940]_  = ~A201 & ~A200;
  assign \new_[79943]_  = A203 & ~A202;
  assign \new_[79944]_  = \new_[79943]_  & \new_[79940]_ ;
  assign \new_[79945]_  = \new_[79944]_  & \new_[79937]_ ;
  assign \new_[79948]_  = A266 & ~A265;
  assign \new_[79951]_  = A268 & A267;
  assign \new_[79952]_  = \new_[79951]_  & \new_[79948]_ ;
  assign \new_[79955]_  = A299 & ~A298;
  assign \new_[79958]_  = A301 & A300;
  assign \new_[79959]_  = \new_[79958]_  & \new_[79955]_ ;
  assign \new_[79960]_  = \new_[79959]_  & \new_[79952]_ ;
  assign \new_[79964]_  = A199 & A166;
  assign \new_[79965]_  = A167 & \new_[79964]_ ;
  assign \new_[79968]_  = ~A201 & ~A200;
  assign \new_[79971]_  = A203 & ~A202;
  assign \new_[79972]_  = \new_[79971]_  & \new_[79968]_ ;
  assign \new_[79973]_  = \new_[79972]_  & \new_[79965]_ ;
  assign \new_[79976]_  = A266 & ~A265;
  assign \new_[79979]_  = A268 & A267;
  assign \new_[79980]_  = \new_[79979]_  & \new_[79976]_ ;
  assign \new_[79983]_  = A299 & ~A298;
  assign \new_[79986]_  = ~A302 & A300;
  assign \new_[79987]_  = \new_[79986]_  & \new_[79983]_ ;
  assign \new_[79988]_  = \new_[79987]_  & \new_[79980]_ ;
  assign \new_[79992]_  = A199 & A166;
  assign \new_[79993]_  = A167 & \new_[79992]_ ;
  assign \new_[79996]_  = ~A201 & ~A200;
  assign \new_[79999]_  = A203 & ~A202;
  assign \new_[80000]_  = \new_[79999]_  & \new_[79996]_ ;
  assign \new_[80001]_  = \new_[80000]_  & \new_[79993]_ ;
  assign \new_[80004]_  = A266 & ~A265;
  assign \new_[80007]_  = ~A269 & A267;
  assign \new_[80008]_  = \new_[80007]_  & \new_[80004]_ ;
  assign \new_[80011]_  = ~A299 & A298;
  assign \new_[80014]_  = A301 & A300;
  assign \new_[80015]_  = \new_[80014]_  & \new_[80011]_ ;
  assign \new_[80016]_  = \new_[80015]_  & \new_[80008]_ ;
  assign \new_[80020]_  = A199 & A166;
  assign \new_[80021]_  = A167 & \new_[80020]_ ;
  assign \new_[80024]_  = ~A201 & ~A200;
  assign \new_[80027]_  = A203 & ~A202;
  assign \new_[80028]_  = \new_[80027]_  & \new_[80024]_ ;
  assign \new_[80029]_  = \new_[80028]_  & \new_[80021]_ ;
  assign \new_[80032]_  = A266 & ~A265;
  assign \new_[80035]_  = ~A269 & A267;
  assign \new_[80036]_  = \new_[80035]_  & \new_[80032]_ ;
  assign \new_[80039]_  = ~A299 & A298;
  assign \new_[80042]_  = ~A302 & A300;
  assign \new_[80043]_  = \new_[80042]_  & \new_[80039]_ ;
  assign \new_[80044]_  = \new_[80043]_  & \new_[80036]_ ;
  assign \new_[80048]_  = A199 & A166;
  assign \new_[80049]_  = A167 & \new_[80048]_ ;
  assign \new_[80052]_  = ~A201 & ~A200;
  assign \new_[80055]_  = A203 & ~A202;
  assign \new_[80056]_  = \new_[80055]_  & \new_[80052]_ ;
  assign \new_[80057]_  = \new_[80056]_  & \new_[80049]_ ;
  assign \new_[80060]_  = A266 & ~A265;
  assign \new_[80063]_  = ~A269 & A267;
  assign \new_[80064]_  = \new_[80063]_  & \new_[80060]_ ;
  assign \new_[80067]_  = A299 & ~A298;
  assign \new_[80070]_  = A301 & A300;
  assign \new_[80071]_  = \new_[80070]_  & \new_[80067]_ ;
  assign \new_[80072]_  = \new_[80071]_  & \new_[80064]_ ;
  assign \new_[80076]_  = A199 & A166;
  assign \new_[80077]_  = A167 & \new_[80076]_ ;
  assign \new_[80080]_  = ~A201 & ~A200;
  assign \new_[80083]_  = A203 & ~A202;
  assign \new_[80084]_  = \new_[80083]_  & \new_[80080]_ ;
  assign \new_[80085]_  = \new_[80084]_  & \new_[80077]_ ;
  assign \new_[80088]_  = A266 & ~A265;
  assign \new_[80091]_  = ~A269 & A267;
  assign \new_[80092]_  = \new_[80091]_  & \new_[80088]_ ;
  assign \new_[80095]_  = A299 & ~A298;
  assign \new_[80098]_  = ~A302 & A300;
  assign \new_[80099]_  = \new_[80098]_  & \new_[80095]_ ;
  assign \new_[80100]_  = \new_[80099]_  & \new_[80092]_ ;
  assign \new_[80104]_  = A199 & A166;
  assign \new_[80105]_  = A167 & \new_[80104]_ ;
  assign \new_[80108]_  = ~A201 & ~A200;
  assign \new_[80111]_  = A203 & ~A202;
  assign \new_[80112]_  = \new_[80111]_  & \new_[80108]_ ;
  assign \new_[80113]_  = \new_[80112]_  & \new_[80105]_ ;
  assign \new_[80116]_  = ~A266 & A265;
  assign \new_[80119]_  = A268 & A267;
  assign \new_[80120]_  = \new_[80119]_  & \new_[80116]_ ;
  assign \new_[80123]_  = ~A299 & A298;
  assign \new_[80126]_  = A301 & A300;
  assign \new_[80127]_  = \new_[80126]_  & \new_[80123]_ ;
  assign \new_[80128]_  = \new_[80127]_  & \new_[80120]_ ;
  assign \new_[80132]_  = A199 & A166;
  assign \new_[80133]_  = A167 & \new_[80132]_ ;
  assign \new_[80136]_  = ~A201 & ~A200;
  assign \new_[80139]_  = A203 & ~A202;
  assign \new_[80140]_  = \new_[80139]_  & \new_[80136]_ ;
  assign \new_[80141]_  = \new_[80140]_  & \new_[80133]_ ;
  assign \new_[80144]_  = ~A266 & A265;
  assign \new_[80147]_  = A268 & A267;
  assign \new_[80148]_  = \new_[80147]_  & \new_[80144]_ ;
  assign \new_[80151]_  = ~A299 & A298;
  assign \new_[80154]_  = ~A302 & A300;
  assign \new_[80155]_  = \new_[80154]_  & \new_[80151]_ ;
  assign \new_[80156]_  = \new_[80155]_  & \new_[80148]_ ;
  assign \new_[80160]_  = A199 & A166;
  assign \new_[80161]_  = A167 & \new_[80160]_ ;
  assign \new_[80164]_  = ~A201 & ~A200;
  assign \new_[80167]_  = A203 & ~A202;
  assign \new_[80168]_  = \new_[80167]_  & \new_[80164]_ ;
  assign \new_[80169]_  = \new_[80168]_  & \new_[80161]_ ;
  assign \new_[80172]_  = ~A266 & A265;
  assign \new_[80175]_  = A268 & A267;
  assign \new_[80176]_  = \new_[80175]_  & \new_[80172]_ ;
  assign \new_[80179]_  = A299 & ~A298;
  assign \new_[80182]_  = A301 & A300;
  assign \new_[80183]_  = \new_[80182]_  & \new_[80179]_ ;
  assign \new_[80184]_  = \new_[80183]_  & \new_[80176]_ ;
  assign \new_[80188]_  = A199 & A166;
  assign \new_[80189]_  = A167 & \new_[80188]_ ;
  assign \new_[80192]_  = ~A201 & ~A200;
  assign \new_[80195]_  = A203 & ~A202;
  assign \new_[80196]_  = \new_[80195]_  & \new_[80192]_ ;
  assign \new_[80197]_  = \new_[80196]_  & \new_[80189]_ ;
  assign \new_[80200]_  = ~A266 & A265;
  assign \new_[80203]_  = A268 & A267;
  assign \new_[80204]_  = \new_[80203]_  & \new_[80200]_ ;
  assign \new_[80207]_  = A299 & ~A298;
  assign \new_[80210]_  = ~A302 & A300;
  assign \new_[80211]_  = \new_[80210]_  & \new_[80207]_ ;
  assign \new_[80212]_  = \new_[80211]_  & \new_[80204]_ ;
  assign \new_[80216]_  = A199 & A166;
  assign \new_[80217]_  = A167 & \new_[80216]_ ;
  assign \new_[80220]_  = ~A201 & ~A200;
  assign \new_[80223]_  = A203 & ~A202;
  assign \new_[80224]_  = \new_[80223]_  & \new_[80220]_ ;
  assign \new_[80225]_  = \new_[80224]_  & \new_[80217]_ ;
  assign \new_[80228]_  = ~A266 & A265;
  assign \new_[80231]_  = ~A269 & A267;
  assign \new_[80232]_  = \new_[80231]_  & \new_[80228]_ ;
  assign \new_[80235]_  = ~A299 & A298;
  assign \new_[80238]_  = A301 & A300;
  assign \new_[80239]_  = \new_[80238]_  & \new_[80235]_ ;
  assign \new_[80240]_  = \new_[80239]_  & \new_[80232]_ ;
  assign \new_[80244]_  = A199 & A166;
  assign \new_[80245]_  = A167 & \new_[80244]_ ;
  assign \new_[80248]_  = ~A201 & ~A200;
  assign \new_[80251]_  = A203 & ~A202;
  assign \new_[80252]_  = \new_[80251]_  & \new_[80248]_ ;
  assign \new_[80253]_  = \new_[80252]_  & \new_[80245]_ ;
  assign \new_[80256]_  = ~A266 & A265;
  assign \new_[80259]_  = ~A269 & A267;
  assign \new_[80260]_  = \new_[80259]_  & \new_[80256]_ ;
  assign \new_[80263]_  = ~A299 & A298;
  assign \new_[80266]_  = ~A302 & A300;
  assign \new_[80267]_  = \new_[80266]_  & \new_[80263]_ ;
  assign \new_[80268]_  = \new_[80267]_  & \new_[80260]_ ;
  assign \new_[80272]_  = A199 & A166;
  assign \new_[80273]_  = A167 & \new_[80272]_ ;
  assign \new_[80276]_  = ~A201 & ~A200;
  assign \new_[80279]_  = A203 & ~A202;
  assign \new_[80280]_  = \new_[80279]_  & \new_[80276]_ ;
  assign \new_[80281]_  = \new_[80280]_  & \new_[80273]_ ;
  assign \new_[80284]_  = ~A266 & A265;
  assign \new_[80287]_  = ~A269 & A267;
  assign \new_[80288]_  = \new_[80287]_  & \new_[80284]_ ;
  assign \new_[80291]_  = A299 & ~A298;
  assign \new_[80294]_  = A301 & A300;
  assign \new_[80295]_  = \new_[80294]_  & \new_[80291]_ ;
  assign \new_[80296]_  = \new_[80295]_  & \new_[80288]_ ;
  assign \new_[80300]_  = A199 & A166;
  assign \new_[80301]_  = A167 & \new_[80300]_ ;
  assign \new_[80304]_  = ~A201 & ~A200;
  assign \new_[80307]_  = A203 & ~A202;
  assign \new_[80308]_  = \new_[80307]_  & \new_[80304]_ ;
  assign \new_[80309]_  = \new_[80308]_  & \new_[80301]_ ;
  assign \new_[80312]_  = ~A266 & A265;
  assign \new_[80315]_  = ~A269 & A267;
  assign \new_[80316]_  = \new_[80315]_  & \new_[80312]_ ;
  assign \new_[80319]_  = A299 & ~A298;
  assign \new_[80322]_  = ~A302 & A300;
  assign \new_[80323]_  = \new_[80322]_  & \new_[80319]_ ;
  assign \new_[80324]_  = \new_[80323]_  & \new_[80316]_ ;
  assign \new_[80328]_  = ~A199 & ~A166;
  assign \new_[80329]_  = ~A167 & \new_[80328]_ ;
  assign \new_[80332]_  = A201 & A200;
  assign \new_[80335]_  = ~A265 & A202;
  assign \new_[80336]_  = \new_[80335]_  & \new_[80332]_ ;
  assign \new_[80337]_  = \new_[80336]_  & \new_[80329]_ ;
  assign \new_[80340]_  = A267 & A266;
  assign \new_[80343]_  = A298 & A268;
  assign \new_[80344]_  = \new_[80343]_  & \new_[80340]_ ;
  assign \new_[80347]_  = ~A300 & ~A299;
  assign \new_[80350]_  = A302 & ~A301;
  assign \new_[80351]_  = \new_[80350]_  & \new_[80347]_ ;
  assign \new_[80352]_  = \new_[80351]_  & \new_[80344]_ ;
  assign \new_[80356]_  = ~A199 & ~A166;
  assign \new_[80357]_  = ~A167 & \new_[80356]_ ;
  assign \new_[80360]_  = A201 & A200;
  assign \new_[80363]_  = ~A265 & A202;
  assign \new_[80364]_  = \new_[80363]_  & \new_[80360]_ ;
  assign \new_[80365]_  = \new_[80364]_  & \new_[80357]_ ;
  assign \new_[80368]_  = A267 & A266;
  assign \new_[80371]_  = ~A298 & A268;
  assign \new_[80372]_  = \new_[80371]_  & \new_[80368]_ ;
  assign \new_[80375]_  = ~A300 & A299;
  assign \new_[80378]_  = A302 & ~A301;
  assign \new_[80379]_  = \new_[80378]_  & \new_[80375]_ ;
  assign \new_[80380]_  = \new_[80379]_  & \new_[80372]_ ;
  assign \new_[80384]_  = ~A199 & ~A166;
  assign \new_[80385]_  = ~A167 & \new_[80384]_ ;
  assign \new_[80388]_  = A201 & A200;
  assign \new_[80391]_  = ~A265 & A202;
  assign \new_[80392]_  = \new_[80391]_  & \new_[80388]_ ;
  assign \new_[80393]_  = \new_[80392]_  & \new_[80385]_ ;
  assign \new_[80396]_  = A267 & A266;
  assign \new_[80399]_  = A298 & ~A269;
  assign \new_[80400]_  = \new_[80399]_  & \new_[80396]_ ;
  assign \new_[80403]_  = ~A300 & ~A299;
  assign \new_[80406]_  = A302 & ~A301;
  assign \new_[80407]_  = \new_[80406]_  & \new_[80403]_ ;
  assign \new_[80408]_  = \new_[80407]_  & \new_[80400]_ ;
  assign \new_[80412]_  = ~A199 & ~A166;
  assign \new_[80413]_  = ~A167 & \new_[80412]_ ;
  assign \new_[80416]_  = A201 & A200;
  assign \new_[80419]_  = ~A265 & A202;
  assign \new_[80420]_  = \new_[80419]_  & \new_[80416]_ ;
  assign \new_[80421]_  = \new_[80420]_  & \new_[80413]_ ;
  assign \new_[80424]_  = A267 & A266;
  assign \new_[80427]_  = ~A298 & ~A269;
  assign \new_[80428]_  = \new_[80427]_  & \new_[80424]_ ;
  assign \new_[80431]_  = ~A300 & A299;
  assign \new_[80434]_  = A302 & ~A301;
  assign \new_[80435]_  = \new_[80434]_  & \new_[80431]_ ;
  assign \new_[80436]_  = \new_[80435]_  & \new_[80428]_ ;
  assign \new_[80440]_  = ~A199 & ~A166;
  assign \new_[80441]_  = ~A167 & \new_[80440]_ ;
  assign \new_[80444]_  = A201 & A200;
  assign \new_[80447]_  = ~A265 & A202;
  assign \new_[80448]_  = \new_[80447]_  & \new_[80444]_ ;
  assign \new_[80449]_  = \new_[80448]_  & \new_[80441]_ ;
  assign \new_[80452]_  = ~A267 & A266;
  assign \new_[80455]_  = A269 & ~A268;
  assign \new_[80456]_  = \new_[80455]_  & \new_[80452]_ ;
  assign \new_[80459]_  = ~A299 & A298;
  assign \new_[80462]_  = A301 & A300;
  assign \new_[80463]_  = \new_[80462]_  & \new_[80459]_ ;
  assign \new_[80464]_  = \new_[80463]_  & \new_[80456]_ ;
  assign \new_[80468]_  = ~A199 & ~A166;
  assign \new_[80469]_  = ~A167 & \new_[80468]_ ;
  assign \new_[80472]_  = A201 & A200;
  assign \new_[80475]_  = ~A265 & A202;
  assign \new_[80476]_  = \new_[80475]_  & \new_[80472]_ ;
  assign \new_[80477]_  = \new_[80476]_  & \new_[80469]_ ;
  assign \new_[80480]_  = ~A267 & A266;
  assign \new_[80483]_  = A269 & ~A268;
  assign \new_[80484]_  = \new_[80483]_  & \new_[80480]_ ;
  assign \new_[80487]_  = ~A299 & A298;
  assign \new_[80490]_  = ~A302 & A300;
  assign \new_[80491]_  = \new_[80490]_  & \new_[80487]_ ;
  assign \new_[80492]_  = \new_[80491]_  & \new_[80484]_ ;
  assign \new_[80496]_  = ~A199 & ~A166;
  assign \new_[80497]_  = ~A167 & \new_[80496]_ ;
  assign \new_[80500]_  = A201 & A200;
  assign \new_[80503]_  = ~A265 & A202;
  assign \new_[80504]_  = \new_[80503]_  & \new_[80500]_ ;
  assign \new_[80505]_  = \new_[80504]_  & \new_[80497]_ ;
  assign \new_[80508]_  = ~A267 & A266;
  assign \new_[80511]_  = A269 & ~A268;
  assign \new_[80512]_  = \new_[80511]_  & \new_[80508]_ ;
  assign \new_[80515]_  = A299 & ~A298;
  assign \new_[80518]_  = A301 & A300;
  assign \new_[80519]_  = \new_[80518]_  & \new_[80515]_ ;
  assign \new_[80520]_  = \new_[80519]_  & \new_[80512]_ ;
  assign \new_[80524]_  = ~A199 & ~A166;
  assign \new_[80525]_  = ~A167 & \new_[80524]_ ;
  assign \new_[80528]_  = A201 & A200;
  assign \new_[80531]_  = ~A265 & A202;
  assign \new_[80532]_  = \new_[80531]_  & \new_[80528]_ ;
  assign \new_[80533]_  = \new_[80532]_  & \new_[80525]_ ;
  assign \new_[80536]_  = ~A267 & A266;
  assign \new_[80539]_  = A269 & ~A268;
  assign \new_[80540]_  = \new_[80539]_  & \new_[80536]_ ;
  assign \new_[80543]_  = A299 & ~A298;
  assign \new_[80546]_  = ~A302 & A300;
  assign \new_[80547]_  = \new_[80546]_  & \new_[80543]_ ;
  assign \new_[80548]_  = \new_[80547]_  & \new_[80540]_ ;
  assign \new_[80552]_  = ~A199 & ~A166;
  assign \new_[80553]_  = ~A167 & \new_[80552]_ ;
  assign \new_[80556]_  = A201 & A200;
  assign \new_[80559]_  = A265 & A202;
  assign \new_[80560]_  = \new_[80559]_  & \new_[80556]_ ;
  assign \new_[80561]_  = \new_[80560]_  & \new_[80553]_ ;
  assign \new_[80564]_  = A267 & ~A266;
  assign \new_[80567]_  = A298 & A268;
  assign \new_[80568]_  = \new_[80567]_  & \new_[80564]_ ;
  assign \new_[80571]_  = ~A300 & ~A299;
  assign \new_[80574]_  = A302 & ~A301;
  assign \new_[80575]_  = \new_[80574]_  & \new_[80571]_ ;
  assign \new_[80576]_  = \new_[80575]_  & \new_[80568]_ ;
  assign \new_[80580]_  = ~A199 & ~A166;
  assign \new_[80581]_  = ~A167 & \new_[80580]_ ;
  assign \new_[80584]_  = A201 & A200;
  assign \new_[80587]_  = A265 & A202;
  assign \new_[80588]_  = \new_[80587]_  & \new_[80584]_ ;
  assign \new_[80589]_  = \new_[80588]_  & \new_[80581]_ ;
  assign \new_[80592]_  = A267 & ~A266;
  assign \new_[80595]_  = ~A298 & A268;
  assign \new_[80596]_  = \new_[80595]_  & \new_[80592]_ ;
  assign \new_[80599]_  = ~A300 & A299;
  assign \new_[80602]_  = A302 & ~A301;
  assign \new_[80603]_  = \new_[80602]_  & \new_[80599]_ ;
  assign \new_[80604]_  = \new_[80603]_  & \new_[80596]_ ;
  assign \new_[80608]_  = ~A199 & ~A166;
  assign \new_[80609]_  = ~A167 & \new_[80608]_ ;
  assign \new_[80612]_  = A201 & A200;
  assign \new_[80615]_  = A265 & A202;
  assign \new_[80616]_  = \new_[80615]_  & \new_[80612]_ ;
  assign \new_[80617]_  = \new_[80616]_  & \new_[80609]_ ;
  assign \new_[80620]_  = A267 & ~A266;
  assign \new_[80623]_  = A298 & ~A269;
  assign \new_[80624]_  = \new_[80623]_  & \new_[80620]_ ;
  assign \new_[80627]_  = ~A300 & ~A299;
  assign \new_[80630]_  = A302 & ~A301;
  assign \new_[80631]_  = \new_[80630]_  & \new_[80627]_ ;
  assign \new_[80632]_  = \new_[80631]_  & \new_[80624]_ ;
  assign \new_[80636]_  = ~A199 & ~A166;
  assign \new_[80637]_  = ~A167 & \new_[80636]_ ;
  assign \new_[80640]_  = A201 & A200;
  assign \new_[80643]_  = A265 & A202;
  assign \new_[80644]_  = \new_[80643]_  & \new_[80640]_ ;
  assign \new_[80645]_  = \new_[80644]_  & \new_[80637]_ ;
  assign \new_[80648]_  = A267 & ~A266;
  assign \new_[80651]_  = ~A298 & ~A269;
  assign \new_[80652]_  = \new_[80651]_  & \new_[80648]_ ;
  assign \new_[80655]_  = ~A300 & A299;
  assign \new_[80658]_  = A302 & ~A301;
  assign \new_[80659]_  = \new_[80658]_  & \new_[80655]_ ;
  assign \new_[80660]_  = \new_[80659]_  & \new_[80652]_ ;
  assign \new_[80664]_  = ~A199 & ~A166;
  assign \new_[80665]_  = ~A167 & \new_[80664]_ ;
  assign \new_[80668]_  = A201 & A200;
  assign \new_[80671]_  = A265 & A202;
  assign \new_[80672]_  = \new_[80671]_  & \new_[80668]_ ;
  assign \new_[80673]_  = \new_[80672]_  & \new_[80665]_ ;
  assign \new_[80676]_  = ~A267 & ~A266;
  assign \new_[80679]_  = A269 & ~A268;
  assign \new_[80680]_  = \new_[80679]_  & \new_[80676]_ ;
  assign \new_[80683]_  = ~A299 & A298;
  assign \new_[80686]_  = A301 & A300;
  assign \new_[80687]_  = \new_[80686]_  & \new_[80683]_ ;
  assign \new_[80688]_  = \new_[80687]_  & \new_[80680]_ ;
  assign \new_[80692]_  = ~A199 & ~A166;
  assign \new_[80693]_  = ~A167 & \new_[80692]_ ;
  assign \new_[80696]_  = A201 & A200;
  assign \new_[80699]_  = A265 & A202;
  assign \new_[80700]_  = \new_[80699]_  & \new_[80696]_ ;
  assign \new_[80701]_  = \new_[80700]_  & \new_[80693]_ ;
  assign \new_[80704]_  = ~A267 & ~A266;
  assign \new_[80707]_  = A269 & ~A268;
  assign \new_[80708]_  = \new_[80707]_  & \new_[80704]_ ;
  assign \new_[80711]_  = ~A299 & A298;
  assign \new_[80714]_  = ~A302 & A300;
  assign \new_[80715]_  = \new_[80714]_  & \new_[80711]_ ;
  assign \new_[80716]_  = \new_[80715]_  & \new_[80708]_ ;
  assign \new_[80720]_  = ~A199 & ~A166;
  assign \new_[80721]_  = ~A167 & \new_[80720]_ ;
  assign \new_[80724]_  = A201 & A200;
  assign \new_[80727]_  = A265 & A202;
  assign \new_[80728]_  = \new_[80727]_  & \new_[80724]_ ;
  assign \new_[80729]_  = \new_[80728]_  & \new_[80721]_ ;
  assign \new_[80732]_  = ~A267 & ~A266;
  assign \new_[80735]_  = A269 & ~A268;
  assign \new_[80736]_  = \new_[80735]_  & \new_[80732]_ ;
  assign \new_[80739]_  = A299 & ~A298;
  assign \new_[80742]_  = A301 & A300;
  assign \new_[80743]_  = \new_[80742]_  & \new_[80739]_ ;
  assign \new_[80744]_  = \new_[80743]_  & \new_[80736]_ ;
  assign \new_[80748]_  = ~A199 & ~A166;
  assign \new_[80749]_  = ~A167 & \new_[80748]_ ;
  assign \new_[80752]_  = A201 & A200;
  assign \new_[80755]_  = A265 & A202;
  assign \new_[80756]_  = \new_[80755]_  & \new_[80752]_ ;
  assign \new_[80757]_  = \new_[80756]_  & \new_[80749]_ ;
  assign \new_[80760]_  = ~A267 & ~A266;
  assign \new_[80763]_  = A269 & ~A268;
  assign \new_[80764]_  = \new_[80763]_  & \new_[80760]_ ;
  assign \new_[80767]_  = A299 & ~A298;
  assign \new_[80770]_  = ~A302 & A300;
  assign \new_[80771]_  = \new_[80770]_  & \new_[80767]_ ;
  assign \new_[80772]_  = \new_[80771]_  & \new_[80764]_ ;
  assign \new_[80776]_  = ~A199 & ~A166;
  assign \new_[80777]_  = ~A167 & \new_[80776]_ ;
  assign \new_[80780]_  = A201 & A200;
  assign \new_[80783]_  = ~A265 & ~A203;
  assign \new_[80784]_  = \new_[80783]_  & \new_[80780]_ ;
  assign \new_[80785]_  = \new_[80784]_  & \new_[80777]_ ;
  assign \new_[80788]_  = A267 & A266;
  assign \new_[80791]_  = A298 & A268;
  assign \new_[80792]_  = \new_[80791]_  & \new_[80788]_ ;
  assign \new_[80795]_  = ~A300 & ~A299;
  assign \new_[80798]_  = A302 & ~A301;
  assign \new_[80799]_  = \new_[80798]_  & \new_[80795]_ ;
  assign \new_[80800]_  = \new_[80799]_  & \new_[80792]_ ;
  assign \new_[80804]_  = ~A199 & ~A166;
  assign \new_[80805]_  = ~A167 & \new_[80804]_ ;
  assign \new_[80808]_  = A201 & A200;
  assign \new_[80811]_  = ~A265 & ~A203;
  assign \new_[80812]_  = \new_[80811]_  & \new_[80808]_ ;
  assign \new_[80813]_  = \new_[80812]_  & \new_[80805]_ ;
  assign \new_[80816]_  = A267 & A266;
  assign \new_[80819]_  = ~A298 & A268;
  assign \new_[80820]_  = \new_[80819]_  & \new_[80816]_ ;
  assign \new_[80823]_  = ~A300 & A299;
  assign \new_[80826]_  = A302 & ~A301;
  assign \new_[80827]_  = \new_[80826]_  & \new_[80823]_ ;
  assign \new_[80828]_  = \new_[80827]_  & \new_[80820]_ ;
  assign \new_[80832]_  = ~A199 & ~A166;
  assign \new_[80833]_  = ~A167 & \new_[80832]_ ;
  assign \new_[80836]_  = A201 & A200;
  assign \new_[80839]_  = ~A265 & ~A203;
  assign \new_[80840]_  = \new_[80839]_  & \new_[80836]_ ;
  assign \new_[80841]_  = \new_[80840]_  & \new_[80833]_ ;
  assign \new_[80844]_  = A267 & A266;
  assign \new_[80847]_  = A298 & ~A269;
  assign \new_[80848]_  = \new_[80847]_  & \new_[80844]_ ;
  assign \new_[80851]_  = ~A300 & ~A299;
  assign \new_[80854]_  = A302 & ~A301;
  assign \new_[80855]_  = \new_[80854]_  & \new_[80851]_ ;
  assign \new_[80856]_  = \new_[80855]_  & \new_[80848]_ ;
  assign \new_[80860]_  = ~A199 & ~A166;
  assign \new_[80861]_  = ~A167 & \new_[80860]_ ;
  assign \new_[80864]_  = A201 & A200;
  assign \new_[80867]_  = ~A265 & ~A203;
  assign \new_[80868]_  = \new_[80867]_  & \new_[80864]_ ;
  assign \new_[80869]_  = \new_[80868]_  & \new_[80861]_ ;
  assign \new_[80872]_  = A267 & A266;
  assign \new_[80875]_  = ~A298 & ~A269;
  assign \new_[80876]_  = \new_[80875]_  & \new_[80872]_ ;
  assign \new_[80879]_  = ~A300 & A299;
  assign \new_[80882]_  = A302 & ~A301;
  assign \new_[80883]_  = \new_[80882]_  & \new_[80879]_ ;
  assign \new_[80884]_  = \new_[80883]_  & \new_[80876]_ ;
  assign \new_[80888]_  = ~A199 & ~A166;
  assign \new_[80889]_  = ~A167 & \new_[80888]_ ;
  assign \new_[80892]_  = A201 & A200;
  assign \new_[80895]_  = ~A265 & ~A203;
  assign \new_[80896]_  = \new_[80895]_  & \new_[80892]_ ;
  assign \new_[80897]_  = \new_[80896]_  & \new_[80889]_ ;
  assign \new_[80900]_  = ~A267 & A266;
  assign \new_[80903]_  = A269 & ~A268;
  assign \new_[80904]_  = \new_[80903]_  & \new_[80900]_ ;
  assign \new_[80907]_  = ~A299 & A298;
  assign \new_[80910]_  = A301 & A300;
  assign \new_[80911]_  = \new_[80910]_  & \new_[80907]_ ;
  assign \new_[80912]_  = \new_[80911]_  & \new_[80904]_ ;
  assign \new_[80916]_  = ~A199 & ~A166;
  assign \new_[80917]_  = ~A167 & \new_[80916]_ ;
  assign \new_[80920]_  = A201 & A200;
  assign \new_[80923]_  = ~A265 & ~A203;
  assign \new_[80924]_  = \new_[80923]_  & \new_[80920]_ ;
  assign \new_[80925]_  = \new_[80924]_  & \new_[80917]_ ;
  assign \new_[80928]_  = ~A267 & A266;
  assign \new_[80931]_  = A269 & ~A268;
  assign \new_[80932]_  = \new_[80931]_  & \new_[80928]_ ;
  assign \new_[80935]_  = ~A299 & A298;
  assign \new_[80938]_  = ~A302 & A300;
  assign \new_[80939]_  = \new_[80938]_  & \new_[80935]_ ;
  assign \new_[80940]_  = \new_[80939]_  & \new_[80932]_ ;
  assign \new_[80944]_  = ~A199 & ~A166;
  assign \new_[80945]_  = ~A167 & \new_[80944]_ ;
  assign \new_[80948]_  = A201 & A200;
  assign \new_[80951]_  = ~A265 & ~A203;
  assign \new_[80952]_  = \new_[80951]_  & \new_[80948]_ ;
  assign \new_[80953]_  = \new_[80952]_  & \new_[80945]_ ;
  assign \new_[80956]_  = ~A267 & A266;
  assign \new_[80959]_  = A269 & ~A268;
  assign \new_[80960]_  = \new_[80959]_  & \new_[80956]_ ;
  assign \new_[80963]_  = A299 & ~A298;
  assign \new_[80966]_  = A301 & A300;
  assign \new_[80967]_  = \new_[80966]_  & \new_[80963]_ ;
  assign \new_[80968]_  = \new_[80967]_  & \new_[80960]_ ;
  assign \new_[80972]_  = ~A199 & ~A166;
  assign \new_[80973]_  = ~A167 & \new_[80972]_ ;
  assign \new_[80976]_  = A201 & A200;
  assign \new_[80979]_  = ~A265 & ~A203;
  assign \new_[80980]_  = \new_[80979]_  & \new_[80976]_ ;
  assign \new_[80981]_  = \new_[80980]_  & \new_[80973]_ ;
  assign \new_[80984]_  = ~A267 & A266;
  assign \new_[80987]_  = A269 & ~A268;
  assign \new_[80988]_  = \new_[80987]_  & \new_[80984]_ ;
  assign \new_[80991]_  = A299 & ~A298;
  assign \new_[80994]_  = ~A302 & A300;
  assign \new_[80995]_  = \new_[80994]_  & \new_[80991]_ ;
  assign \new_[80996]_  = \new_[80995]_  & \new_[80988]_ ;
  assign \new_[81000]_  = ~A199 & ~A166;
  assign \new_[81001]_  = ~A167 & \new_[81000]_ ;
  assign \new_[81004]_  = A201 & A200;
  assign \new_[81007]_  = A265 & ~A203;
  assign \new_[81008]_  = \new_[81007]_  & \new_[81004]_ ;
  assign \new_[81009]_  = \new_[81008]_  & \new_[81001]_ ;
  assign \new_[81012]_  = A267 & ~A266;
  assign \new_[81015]_  = A298 & A268;
  assign \new_[81016]_  = \new_[81015]_  & \new_[81012]_ ;
  assign \new_[81019]_  = ~A300 & ~A299;
  assign \new_[81022]_  = A302 & ~A301;
  assign \new_[81023]_  = \new_[81022]_  & \new_[81019]_ ;
  assign \new_[81024]_  = \new_[81023]_  & \new_[81016]_ ;
  assign \new_[81028]_  = ~A199 & ~A166;
  assign \new_[81029]_  = ~A167 & \new_[81028]_ ;
  assign \new_[81032]_  = A201 & A200;
  assign \new_[81035]_  = A265 & ~A203;
  assign \new_[81036]_  = \new_[81035]_  & \new_[81032]_ ;
  assign \new_[81037]_  = \new_[81036]_  & \new_[81029]_ ;
  assign \new_[81040]_  = A267 & ~A266;
  assign \new_[81043]_  = ~A298 & A268;
  assign \new_[81044]_  = \new_[81043]_  & \new_[81040]_ ;
  assign \new_[81047]_  = ~A300 & A299;
  assign \new_[81050]_  = A302 & ~A301;
  assign \new_[81051]_  = \new_[81050]_  & \new_[81047]_ ;
  assign \new_[81052]_  = \new_[81051]_  & \new_[81044]_ ;
  assign \new_[81056]_  = ~A199 & ~A166;
  assign \new_[81057]_  = ~A167 & \new_[81056]_ ;
  assign \new_[81060]_  = A201 & A200;
  assign \new_[81063]_  = A265 & ~A203;
  assign \new_[81064]_  = \new_[81063]_  & \new_[81060]_ ;
  assign \new_[81065]_  = \new_[81064]_  & \new_[81057]_ ;
  assign \new_[81068]_  = A267 & ~A266;
  assign \new_[81071]_  = A298 & ~A269;
  assign \new_[81072]_  = \new_[81071]_  & \new_[81068]_ ;
  assign \new_[81075]_  = ~A300 & ~A299;
  assign \new_[81078]_  = A302 & ~A301;
  assign \new_[81079]_  = \new_[81078]_  & \new_[81075]_ ;
  assign \new_[81080]_  = \new_[81079]_  & \new_[81072]_ ;
  assign \new_[81084]_  = ~A199 & ~A166;
  assign \new_[81085]_  = ~A167 & \new_[81084]_ ;
  assign \new_[81088]_  = A201 & A200;
  assign \new_[81091]_  = A265 & ~A203;
  assign \new_[81092]_  = \new_[81091]_  & \new_[81088]_ ;
  assign \new_[81093]_  = \new_[81092]_  & \new_[81085]_ ;
  assign \new_[81096]_  = A267 & ~A266;
  assign \new_[81099]_  = ~A298 & ~A269;
  assign \new_[81100]_  = \new_[81099]_  & \new_[81096]_ ;
  assign \new_[81103]_  = ~A300 & A299;
  assign \new_[81106]_  = A302 & ~A301;
  assign \new_[81107]_  = \new_[81106]_  & \new_[81103]_ ;
  assign \new_[81108]_  = \new_[81107]_  & \new_[81100]_ ;
  assign \new_[81112]_  = ~A199 & ~A166;
  assign \new_[81113]_  = ~A167 & \new_[81112]_ ;
  assign \new_[81116]_  = A201 & A200;
  assign \new_[81119]_  = A265 & ~A203;
  assign \new_[81120]_  = \new_[81119]_  & \new_[81116]_ ;
  assign \new_[81121]_  = \new_[81120]_  & \new_[81113]_ ;
  assign \new_[81124]_  = ~A267 & ~A266;
  assign \new_[81127]_  = A269 & ~A268;
  assign \new_[81128]_  = \new_[81127]_  & \new_[81124]_ ;
  assign \new_[81131]_  = ~A299 & A298;
  assign \new_[81134]_  = A301 & A300;
  assign \new_[81135]_  = \new_[81134]_  & \new_[81131]_ ;
  assign \new_[81136]_  = \new_[81135]_  & \new_[81128]_ ;
  assign \new_[81140]_  = ~A199 & ~A166;
  assign \new_[81141]_  = ~A167 & \new_[81140]_ ;
  assign \new_[81144]_  = A201 & A200;
  assign \new_[81147]_  = A265 & ~A203;
  assign \new_[81148]_  = \new_[81147]_  & \new_[81144]_ ;
  assign \new_[81149]_  = \new_[81148]_  & \new_[81141]_ ;
  assign \new_[81152]_  = ~A267 & ~A266;
  assign \new_[81155]_  = A269 & ~A268;
  assign \new_[81156]_  = \new_[81155]_  & \new_[81152]_ ;
  assign \new_[81159]_  = ~A299 & A298;
  assign \new_[81162]_  = ~A302 & A300;
  assign \new_[81163]_  = \new_[81162]_  & \new_[81159]_ ;
  assign \new_[81164]_  = \new_[81163]_  & \new_[81156]_ ;
  assign \new_[81168]_  = ~A199 & ~A166;
  assign \new_[81169]_  = ~A167 & \new_[81168]_ ;
  assign \new_[81172]_  = A201 & A200;
  assign \new_[81175]_  = A265 & ~A203;
  assign \new_[81176]_  = \new_[81175]_  & \new_[81172]_ ;
  assign \new_[81177]_  = \new_[81176]_  & \new_[81169]_ ;
  assign \new_[81180]_  = ~A267 & ~A266;
  assign \new_[81183]_  = A269 & ~A268;
  assign \new_[81184]_  = \new_[81183]_  & \new_[81180]_ ;
  assign \new_[81187]_  = A299 & ~A298;
  assign \new_[81190]_  = A301 & A300;
  assign \new_[81191]_  = \new_[81190]_  & \new_[81187]_ ;
  assign \new_[81192]_  = \new_[81191]_  & \new_[81184]_ ;
  assign \new_[81196]_  = ~A199 & ~A166;
  assign \new_[81197]_  = ~A167 & \new_[81196]_ ;
  assign \new_[81200]_  = A201 & A200;
  assign \new_[81203]_  = A265 & ~A203;
  assign \new_[81204]_  = \new_[81203]_  & \new_[81200]_ ;
  assign \new_[81205]_  = \new_[81204]_  & \new_[81197]_ ;
  assign \new_[81208]_  = ~A267 & ~A266;
  assign \new_[81211]_  = A269 & ~A268;
  assign \new_[81212]_  = \new_[81211]_  & \new_[81208]_ ;
  assign \new_[81215]_  = A299 & ~A298;
  assign \new_[81218]_  = ~A302 & A300;
  assign \new_[81219]_  = \new_[81218]_  & \new_[81215]_ ;
  assign \new_[81220]_  = \new_[81219]_  & \new_[81212]_ ;
  assign \new_[81224]_  = ~A199 & ~A166;
  assign \new_[81225]_  = ~A167 & \new_[81224]_ ;
  assign \new_[81228]_  = ~A201 & A200;
  assign \new_[81231]_  = A203 & ~A202;
  assign \new_[81232]_  = \new_[81231]_  & \new_[81228]_ ;
  assign \new_[81233]_  = \new_[81232]_  & \new_[81225]_ ;
  assign \new_[81236]_  = A266 & ~A265;
  assign \new_[81239]_  = A268 & A267;
  assign \new_[81240]_  = \new_[81239]_  & \new_[81236]_ ;
  assign \new_[81243]_  = ~A299 & A298;
  assign \new_[81246]_  = A301 & A300;
  assign \new_[81247]_  = \new_[81246]_  & \new_[81243]_ ;
  assign \new_[81248]_  = \new_[81247]_  & \new_[81240]_ ;
  assign \new_[81252]_  = ~A199 & ~A166;
  assign \new_[81253]_  = ~A167 & \new_[81252]_ ;
  assign \new_[81256]_  = ~A201 & A200;
  assign \new_[81259]_  = A203 & ~A202;
  assign \new_[81260]_  = \new_[81259]_  & \new_[81256]_ ;
  assign \new_[81261]_  = \new_[81260]_  & \new_[81253]_ ;
  assign \new_[81264]_  = A266 & ~A265;
  assign \new_[81267]_  = A268 & A267;
  assign \new_[81268]_  = \new_[81267]_  & \new_[81264]_ ;
  assign \new_[81271]_  = ~A299 & A298;
  assign \new_[81274]_  = ~A302 & A300;
  assign \new_[81275]_  = \new_[81274]_  & \new_[81271]_ ;
  assign \new_[81276]_  = \new_[81275]_  & \new_[81268]_ ;
  assign \new_[81280]_  = ~A199 & ~A166;
  assign \new_[81281]_  = ~A167 & \new_[81280]_ ;
  assign \new_[81284]_  = ~A201 & A200;
  assign \new_[81287]_  = A203 & ~A202;
  assign \new_[81288]_  = \new_[81287]_  & \new_[81284]_ ;
  assign \new_[81289]_  = \new_[81288]_  & \new_[81281]_ ;
  assign \new_[81292]_  = A266 & ~A265;
  assign \new_[81295]_  = A268 & A267;
  assign \new_[81296]_  = \new_[81295]_  & \new_[81292]_ ;
  assign \new_[81299]_  = A299 & ~A298;
  assign \new_[81302]_  = A301 & A300;
  assign \new_[81303]_  = \new_[81302]_  & \new_[81299]_ ;
  assign \new_[81304]_  = \new_[81303]_  & \new_[81296]_ ;
  assign \new_[81308]_  = ~A199 & ~A166;
  assign \new_[81309]_  = ~A167 & \new_[81308]_ ;
  assign \new_[81312]_  = ~A201 & A200;
  assign \new_[81315]_  = A203 & ~A202;
  assign \new_[81316]_  = \new_[81315]_  & \new_[81312]_ ;
  assign \new_[81317]_  = \new_[81316]_  & \new_[81309]_ ;
  assign \new_[81320]_  = A266 & ~A265;
  assign \new_[81323]_  = A268 & A267;
  assign \new_[81324]_  = \new_[81323]_  & \new_[81320]_ ;
  assign \new_[81327]_  = A299 & ~A298;
  assign \new_[81330]_  = ~A302 & A300;
  assign \new_[81331]_  = \new_[81330]_  & \new_[81327]_ ;
  assign \new_[81332]_  = \new_[81331]_  & \new_[81324]_ ;
  assign \new_[81336]_  = ~A199 & ~A166;
  assign \new_[81337]_  = ~A167 & \new_[81336]_ ;
  assign \new_[81340]_  = ~A201 & A200;
  assign \new_[81343]_  = A203 & ~A202;
  assign \new_[81344]_  = \new_[81343]_  & \new_[81340]_ ;
  assign \new_[81345]_  = \new_[81344]_  & \new_[81337]_ ;
  assign \new_[81348]_  = A266 & ~A265;
  assign \new_[81351]_  = ~A269 & A267;
  assign \new_[81352]_  = \new_[81351]_  & \new_[81348]_ ;
  assign \new_[81355]_  = ~A299 & A298;
  assign \new_[81358]_  = A301 & A300;
  assign \new_[81359]_  = \new_[81358]_  & \new_[81355]_ ;
  assign \new_[81360]_  = \new_[81359]_  & \new_[81352]_ ;
  assign \new_[81364]_  = ~A199 & ~A166;
  assign \new_[81365]_  = ~A167 & \new_[81364]_ ;
  assign \new_[81368]_  = ~A201 & A200;
  assign \new_[81371]_  = A203 & ~A202;
  assign \new_[81372]_  = \new_[81371]_  & \new_[81368]_ ;
  assign \new_[81373]_  = \new_[81372]_  & \new_[81365]_ ;
  assign \new_[81376]_  = A266 & ~A265;
  assign \new_[81379]_  = ~A269 & A267;
  assign \new_[81380]_  = \new_[81379]_  & \new_[81376]_ ;
  assign \new_[81383]_  = ~A299 & A298;
  assign \new_[81386]_  = ~A302 & A300;
  assign \new_[81387]_  = \new_[81386]_  & \new_[81383]_ ;
  assign \new_[81388]_  = \new_[81387]_  & \new_[81380]_ ;
  assign \new_[81392]_  = ~A199 & ~A166;
  assign \new_[81393]_  = ~A167 & \new_[81392]_ ;
  assign \new_[81396]_  = ~A201 & A200;
  assign \new_[81399]_  = A203 & ~A202;
  assign \new_[81400]_  = \new_[81399]_  & \new_[81396]_ ;
  assign \new_[81401]_  = \new_[81400]_  & \new_[81393]_ ;
  assign \new_[81404]_  = A266 & ~A265;
  assign \new_[81407]_  = ~A269 & A267;
  assign \new_[81408]_  = \new_[81407]_  & \new_[81404]_ ;
  assign \new_[81411]_  = A299 & ~A298;
  assign \new_[81414]_  = A301 & A300;
  assign \new_[81415]_  = \new_[81414]_  & \new_[81411]_ ;
  assign \new_[81416]_  = \new_[81415]_  & \new_[81408]_ ;
  assign \new_[81420]_  = ~A199 & ~A166;
  assign \new_[81421]_  = ~A167 & \new_[81420]_ ;
  assign \new_[81424]_  = ~A201 & A200;
  assign \new_[81427]_  = A203 & ~A202;
  assign \new_[81428]_  = \new_[81427]_  & \new_[81424]_ ;
  assign \new_[81429]_  = \new_[81428]_  & \new_[81421]_ ;
  assign \new_[81432]_  = A266 & ~A265;
  assign \new_[81435]_  = ~A269 & A267;
  assign \new_[81436]_  = \new_[81435]_  & \new_[81432]_ ;
  assign \new_[81439]_  = A299 & ~A298;
  assign \new_[81442]_  = ~A302 & A300;
  assign \new_[81443]_  = \new_[81442]_  & \new_[81439]_ ;
  assign \new_[81444]_  = \new_[81443]_  & \new_[81436]_ ;
  assign \new_[81448]_  = ~A199 & ~A166;
  assign \new_[81449]_  = ~A167 & \new_[81448]_ ;
  assign \new_[81452]_  = ~A201 & A200;
  assign \new_[81455]_  = A203 & ~A202;
  assign \new_[81456]_  = \new_[81455]_  & \new_[81452]_ ;
  assign \new_[81457]_  = \new_[81456]_  & \new_[81449]_ ;
  assign \new_[81460]_  = ~A266 & A265;
  assign \new_[81463]_  = A268 & A267;
  assign \new_[81464]_  = \new_[81463]_  & \new_[81460]_ ;
  assign \new_[81467]_  = ~A299 & A298;
  assign \new_[81470]_  = A301 & A300;
  assign \new_[81471]_  = \new_[81470]_  & \new_[81467]_ ;
  assign \new_[81472]_  = \new_[81471]_  & \new_[81464]_ ;
  assign \new_[81476]_  = ~A199 & ~A166;
  assign \new_[81477]_  = ~A167 & \new_[81476]_ ;
  assign \new_[81480]_  = ~A201 & A200;
  assign \new_[81483]_  = A203 & ~A202;
  assign \new_[81484]_  = \new_[81483]_  & \new_[81480]_ ;
  assign \new_[81485]_  = \new_[81484]_  & \new_[81477]_ ;
  assign \new_[81488]_  = ~A266 & A265;
  assign \new_[81491]_  = A268 & A267;
  assign \new_[81492]_  = \new_[81491]_  & \new_[81488]_ ;
  assign \new_[81495]_  = ~A299 & A298;
  assign \new_[81498]_  = ~A302 & A300;
  assign \new_[81499]_  = \new_[81498]_  & \new_[81495]_ ;
  assign \new_[81500]_  = \new_[81499]_  & \new_[81492]_ ;
  assign \new_[81504]_  = ~A199 & ~A166;
  assign \new_[81505]_  = ~A167 & \new_[81504]_ ;
  assign \new_[81508]_  = ~A201 & A200;
  assign \new_[81511]_  = A203 & ~A202;
  assign \new_[81512]_  = \new_[81511]_  & \new_[81508]_ ;
  assign \new_[81513]_  = \new_[81512]_  & \new_[81505]_ ;
  assign \new_[81516]_  = ~A266 & A265;
  assign \new_[81519]_  = A268 & A267;
  assign \new_[81520]_  = \new_[81519]_  & \new_[81516]_ ;
  assign \new_[81523]_  = A299 & ~A298;
  assign \new_[81526]_  = A301 & A300;
  assign \new_[81527]_  = \new_[81526]_  & \new_[81523]_ ;
  assign \new_[81528]_  = \new_[81527]_  & \new_[81520]_ ;
  assign \new_[81532]_  = ~A199 & ~A166;
  assign \new_[81533]_  = ~A167 & \new_[81532]_ ;
  assign \new_[81536]_  = ~A201 & A200;
  assign \new_[81539]_  = A203 & ~A202;
  assign \new_[81540]_  = \new_[81539]_  & \new_[81536]_ ;
  assign \new_[81541]_  = \new_[81540]_  & \new_[81533]_ ;
  assign \new_[81544]_  = ~A266 & A265;
  assign \new_[81547]_  = A268 & A267;
  assign \new_[81548]_  = \new_[81547]_  & \new_[81544]_ ;
  assign \new_[81551]_  = A299 & ~A298;
  assign \new_[81554]_  = ~A302 & A300;
  assign \new_[81555]_  = \new_[81554]_  & \new_[81551]_ ;
  assign \new_[81556]_  = \new_[81555]_  & \new_[81548]_ ;
  assign \new_[81560]_  = ~A199 & ~A166;
  assign \new_[81561]_  = ~A167 & \new_[81560]_ ;
  assign \new_[81564]_  = ~A201 & A200;
  assign \new_[81567]_  = A203 & ~A202;
  assign \new_[81568]_  = \new_[81567]_  & \new_[81564]_ ;
  assign \new_[81569]_  = \new_[81568]_  & \new_[81561]_ ;
  assign \new_[81572]_  = ~A266 & A265;
  assign \new_[81575]_  = ~A269 & A267;
  assign \new_[81576]_  = \new_[81575]_  & \new_[81572]_ ;
  assign \new_[81579]_  = ~A299 & A298;
  assign \new_[81582]_  = A301 & A300;
  assign \new_[81583]_  = \new_[81582]_  & \new_[81579]_ ;
  assign \new_[81584]_  = \new_[81583]_  & \new_[81576]_ ;
  assign \new_[81588]_  = ~A199 & ~A166;
  assign \new_[81589]_  = ~A167 & \new_[81588]_ ;
  assign \new_[81592]_  = ~A201 & A200;
  assign \new_[81595]_  = A203 & ~A202;
  assign \new_[81596]_  = \new_[81595]_  & \new_[81592]_ ;
  assign \new_[81597]_  = \new_[81596]_  & \new_[81589]_ ;
  assign \new_[81600]_  = ~A266 & A265;
  assign \new_[81603]_  = ~A269 & A267;
  assign \new_[81604]_  = \new_[81603]_  & \new_[81600]_ ;
  assign \new_[81607]_  = ~A299 & A298;
  assign \new_[81610]_  = ~A302 & A300;
  assign \new_[81611]_  = \new_[81610]_  & \new_[81607]_ ;
  assign \new_[81612]_  = \new_[81611]_  & \new_[81604]_ ;
  assign \new_[81616]_  = ~A199 & ~A166;
  assign \new_[81617]_  = ~A167 & \new_[81616]_ ;
  assign \new_[81620]_  = ~A201 & A200;
  assign \new_[81623]_  = A203 & ~A202;
  assign \new_[81624]_  = \new_[81623]_  & \new_[81620]_ ;
  assign \new_[81625]_  = \new_[81624]_  & \new_[81617]_ ;
  assign \new_[81628]_  = ~A266 & A265;
  assign \new_[81631]_  = ~A269 & A267;
  assign \new_[81632]_  = \new_[81631]_  & \new_[81628]_ ;
  assign \new_[81635]_  = A299 & ~A298;
  assign \new_[81638]_  = A301 & A300;
  assign \new_[81639]_  = \new_[81638]_  & \new_[81635]_ ;
  assign \new_[81640]_  = \new_[81639]_  & \new_[81632]_ ;
  assign \new_[81644]_  = ~A199 & ~A166;
  assign \new_[81645]_  = ~A167 & \new_[81644]_ ;
  assign \new_[81648]_  = ~A201 & A200;
  assign \new_[81651]_  = A203 & ~A202;
  assign \new_[81652]_  = \new_[81651]_  & \new_[81648]_ ;
  assign \new_[81653]_  = \new_[81652]_  & \new_[81645]_ ;
  assign \new_[81656]_  = ~A266 & A265;
  assign \new_[81659]_  = ~A269 & A267;
  assign \new_[81660]_  = \new_[81659]_  & \new_[81656]_ ;
  assign \new_[81663]_  = A299 & ~A298;
  assign \new_[81666]_  = ~A302 & A300;
  assign \new_[81667]_  = \new_[81666]_  & \new_[81663]_ ;
  assign \new_[81668]_  = \new_[81667]_  & \new_[81660]_ ;
  assign \new_[81672]_  = A199 & ~A166;
  assign \new_[81673]_  = ~A167 & \new_[81672]_ ;
  assign \new_[81676]_  = A201 & ~A200;
  assign \new_[81679]_  = ~A265 & A202;
  assign \new_[81680]_  = \new_[81679]_  & \new_[81676]_ ;
  assign \new_[81681]_  = \new_[81680]_  & \new_[81673]_ ;
  assign \new_[81684]_  = A267 & A266;
  assign \new_[81687]_  = A298 & A268;
  assign \new_[81688]_  = \new_[81687]_  & \new_[81684]_ ;
  assign \new_[81691]_  = ~A300 & ~A299;
  assign \new_[81694]_  = A302 & ~A301;
  assign \new_[81695]_  = \new_[81694]_  & \new_[81691]_ ;
  assign \new_[81696]_  = \new_[81695]_  & \new_[81688]_ ;
  assign \new_[81700]_  = A199 & ~A166;
  assign \new_[81701]_  = ~A167 & \new_[81700]_ ;
  assign \new_[81704]_  = A201 & ~A200;
  assign \new_[81707]_  = ~A265 & A202;
  assign \new_[81708]_  = \new_[81707]_  & \new_[81704]_ ;
  assign \new_[81709]_  = \new_[81708]_  & \new_[81701]_ ;
  assign \new_[81712]_  = A267 & A266;
  assign \new_[81715]_  = ~A298 & A268;
  assign \new_[81716]_  = \new_[81715]_  & \new_[81712]_ ;
  assign \new_[81719]_  = ~A300 & A299;
  assign \new_[81722]_  = A302 & ~A301;
  assign \new_[81723]_  = \new_[81722]_  & \new_[81719]_ ;
  assign \new_[81724]_  = \new_[81723]_  & \new_[81716]_ ;
  assign \new_[81728]_  = A199 & ~A166;
  assign \new_[81729]_  = ~A167 & \new_[81728]_ ;
  assign \new_[81732]_  = A201 & ~A200;
  assign \new_[81735]_  = ~A265 & A202;
  assign \new_[81736]_  = \new_[81735]_  & \new_[81732]_ ;
  assign \new_[81737]_  = \new_[81736]_  & \new_[81729]_ ;
  assign \new_[81740]_  = A267 & A266;
  assign \new_[81743]_  = A298 & ~A269;
  assign \new_[81744]_  = \new_[81743]_  & \new_[81740]_ ;
  assign \new_[81747]_  = ~A300 & ~A299;
  assign \new_[81750]_  = A302 & ~A301;
  assign \new_[81751]_  = \new_[81750]_  & \new_[81747]_ ;
  assign \new_[81752]_  = \new_[81751]_  & \new_[81744]_ ;
  assign \new_[81756]_  = A199 & ~A166;
  assign \new_[81757]_  = ~A167 & \new_[81756]_ ;
  assign \new_[81760]_  = A201 & ~A200;
  assign \new_[81763]_  = ~A265 & A202;
  assign \new_[81764]_  = \new_[81763]_  & \new_[81760]_ ;
  assign \new_[81765]_  = \new_[81764]_  & \new_[81757]_ ;
  assign \new_[81768]_  = A267 & A266;
  assign \new_[81771]_  = ~A298 & ~A269;
  assign \new_[81772]_  = \new_[81771]_  & \new_[81768]_ ;
  assign \new_[81775]_  = ~A300 & A299;
  assign \new_[81778]_  = A302 & ~A301;
  assign \new_[81779]_  = \new_[81778]_  & \new_[81775]_ ;
  assign \new_[81780]_  = \new_[81779]_  & \new_[81772]_ ;
  assign \new_[81784]_  = A199 & ~A166;
  assign \new_[81785]_  = ~A167 & \new_[81784]_ ;
  assign \new_[81788]_  = A201 & ~A200;
  assign \new_[81791]_  = ~A265 & A202;
  assign \new_[81792]_  = \new_[81791]_  & \new_[81788]_ ;
  assign \new_[81793]_  = \new_[81792]_  & \new_[81785]_ ;
  assign \new_[81796]_  = ~A267 & A266;
  assign \new_[81799]_  = A269 & ~A268;
  assign \new_[81800]_  = \new_[81799]_  & \new_[81796]_ ;
  assign \new_[81803]_  = ~A299 & A298;
  assign \new_[81806]_  = A301 & A300;
  assign \new_[81807]_  = \new_[81806]_  & \new_[81803]_ ;
  assign \new_[81808]_  = \new_[81807]_  & \new_[81800]_ ;
  assign \new_[81812]_  = A199 & ~A166;
  assign \new_[81813]_  = ~A167 & \new_[81812]_ ;
  assign \new_[81816]_  = A201 & ~A200;
  assign \new_[81819]_  = ~A265 & A202;
  assign \new_[81820]_  = \new_[81819]_  & \new_[81816]_ ;
  assign \new_[81821]_  = \new_[81820]_  & \new_[81813]_ ;
  assign \new_[81824]_  = ~A267 & A266;
  assign \new_[81827]_  = A269 & ~A268;
  assign \new_[81828]_  = \new_[81827]_  & \new_[81824]_ ;
  assign \new_[81831]_  = ~A299 & A298;
  assign \new_[81834]_  = ~A302 & A300;
  assign \new_[81835]_  = \new_[81834]_  & \new_[81831]_ ;
  assign \new_[81836]_  = \new_[81835]_  & \new_[81828]_ ;
  assign \new_[81840]_  = A199 & ~A166;
  assign \new_[81841]_  = ~A167 & \new_[81840]_ ;
  assign \new_[81844]_  = A201 & ~A200;
  assign \new_[81847]_  = ~A265 & A202;
  assign \new_[81848]_  = \new_[81847]_  & \new_[81844]_ ;
  assign \new_[81849]_  = \new_[81848]_  & \new_[81841]_ ;
  assign \new_[81852]_  = ~A267 & A266;
  assign \new_[81855]_  = A269 & ~A268;
  assign \new_[81856]_  = \new_[81855]_  & \new_[81852]_ ;
  assign \new_[81859]_  = A299 & ~A298;
  assign \new_[81862]_  = A301 & A300;
  assign \new_[81863]_  = \new_[81862]_  & \new_[81859]_ ;
  assign \new_[81864]_  = \new_[81863]_  & \new_[81856]_ ;
  assign \new_[81868]_  = A199 & ~A166;
  assign \new_[81869]_  = ~A167 & \new_[81868]_ ;
  assign \new_[81872]_  = A201 & ~A200;
  assign \new_[81875]_  = ~A265 & A202;
  assign \new_[81876]_  = \new_[81875]_  & \new_[81872]_ ;
  assign \new_[81877]_  = \new_[81876]_  & \new_[81869]_ ;
  assign \new_[81880]_  = ~A267 & A266;
  assign \new_[81883]_  = A269 & ~A268;
  assign \new_[81884]_  = \new_[81883]_  & \new_[81880]_ ;
  assign \new_[81887]_  = A299 & ~A298;
  assign \new_[81890]_  = ~A302 & A300;
  assign \new_[81891]_  = \new_[81890]_  & \new_[81887]_ ;
  assign \new_[81892]_  = \new_[81891]_  & \new_[81884]_ ;
  assign \new_[81896]_  = A199 & ~A166;
  assign \new_[81897]_  = ~A167 & \new_[81896]_ ;
  assign \new_[81900]_  = A201 & ~A200;
  assign \new_[81903]_  = A265 & A202;
  assign \new_[81904]_  = \new_[81903]_  & \new_[81900]_ ;
  assign \new_[81905]_  = \new_[81904]_  & \new_[81897]_ ;
  assign \new_[81908]_  = A267 & ~A266;
  assign \new_[81911]_  = A298 & A268;
  assign \new_[81912]_  = \new_[81911]_  & \new_[81908]_ ;
  assign \new_[81915]_  = ~A300 & ~A299;
  assign \new_[81918]_  = A302 & ~A301;
  assign \new_[81919]_  = \new_[81918]_  & \new_[81915]_ ;
  assign \new_[81920]_  = \new_[81919]_  & \new_[81912]_ ;
  assign \new_[81924]_  = A199 & ~A166;
  assign \new_[81925]_  = ~A167 & \new_[81924]_ ;
  assign \new_[81928]_  = A201 & ~A200;
  assign \new_[81931]_  = A265 & A202;
  assign \new_[81932]_  = \new_[81931]_  & \new_[81928]_ ;
  assign \new_[81933]_  = \new_[81932]_  & \new_[81925]_ ;
  assign \new_[81936]_  = A267 & ~A266;
  assign \new_[81939]_  = ~A298 & A268;
  assign \new_[81940]_  = \new_[81939]_  & \new_[81936]_ ;
  assign \new_[81943]_  = ~A300 & A299;
  assign \new_[81946]_  = A302 & ~A301;
  assign \new_[81947]_  = \new_[81946]_  & \new_[81943]_ ;
  assign \new_[81948]_  = \new_[81947]_  & \new_[81940]_ ;
  assign \new_[81952]_  = A199 & ~A166;
  assign \new_[81953]_  = ~A167 & \new_[81952]_ ;
  assign \new_[81956]_  = A201 & ~A200;
  assign \new_[81959]_  = A265 & A202;
  assign \new_[81960]_  = \new_[81959]_  & \new_[81956]_ ;
  assign \new_[81961]_  = \new_[81960]_  & \new_[81953]_ ;
  assign \new_[81964]_  = A267 & ~A266;
  assign \new_[81967]_  = A298 & ~A269;
  assign \new_[81968]_  = \new_[81967]_  & \new_[81964]_ ;
  assign \new_[81971]_  = ~A300 & ~A299;
  assign \new_[81974]_  = A302 & ~A301;
  assign \new_[81975]_  = \new_[81974]_  & \new_[81971]_ ;
  assign \new_[81976]_  = \new_[81975]_  & \new_[81968]_ ;
  assign \new_[81980]_  = A199 & ~A166;
  assign \new_[81981]_  = ~A167 & \new_[81980]_ ;
  assign \new_[81984]_  = A201 & ~A200;
  assign \new_[81987]_  = A265 & A202;
  assign \new_[81988]_  = \new_[81987]_  & \new_[81984]_ ;
  assign \new_[81989]_  = \new_[81988]_  & \new_[81981]_ ;
  assign \new_[81992]_  = A267 & ~A266;
  assign \new_[81995]_  = ~A298 & ~A269;
  assign \new_[81996]_  = \new_[81995]_  & \new_[81992]_ ;
  assign \new_[81999]_  = ~A300 & A299;
  assign \new_[82002]_  = A302 & ~A301;
  assign \new_[82003]_  = \new_[82002]_  & \new_[81999]_ ;
  assign \new_[82004]_  = \new_[82003]_  & \new_[81996]_ ;
  assign \new_[82008]_  = A199 & ~A166;
  assign \new_[82009]_  = ~A167 & \new_[82008]_ ;
  assign \new_[82012]_  = A201 & ~A200;
  assign \new_[82015]_  = A265 & A202;
  assign \new_[82016]_  = \new_[82015]_  & \new_[82012]_ ;
  assign \new_[82017]_  = \new_[82016]_  & \new_[82009]_ ;
  assign \new_[82020]_  = ~A267 & ~A266;
  assign \new_[82023]_  = A269 & ~A268;
  assign \new_[82024]_  = \new_[82023]_  & \new_[82020]_ ;
  assign \new_[82027]_  = ~A299 & A298;
  assign \new_[82030]_  = A301 & A300;
  assign \new_[82031]_  = \new_[82030]_  & \new_[82027]_ ;
  assign \new_[82032]_  = \new_[82031]_  & \new_[82024]_ ;
  assign \new_[82036]_  = A199 & ~A166;
  assign \new_[82037]_  = ~A167 & \new_[82036]_ ;
  assign \new_[82040]_  = A201 & ~A200;
  assign \new_[82043]_  = A265 & A202;
  assign \new_[82044]_  = \new_[82043]_  & \new_[82040]_ ;
  assign \new_[82045]_  = \new_[82044]_  & \new_[82037]_ ;
  assign \new_[82048]_  = ~A267 & ~A266;
  assign \new_[82051]_  = A269 & ~A268;
  assign \new_[82052]_  = \new_[82051]_  & \new_[82048]_ ;
  assign \new_[82055]_  = ~A299 & A298;
  assign \new_[82058]_  = ~A302 & A300;
  assign \new_[82059]_  = \new_[82058]_  & \new_[82055]_ ;
  assign \new_[82060]_  = \new_[82059]_  & \new_[82052]_ ;
  assign \new_[82064]_  = A199 & ~A166;
  assign \new_[82065]_  = ~A167 & \new_[82064]_ ;
  assign \new_[82068]_  = A201 & ~A200;
  assign \new_[82071]_  = A265 & A202;
  assign \new_[82072]_  = \new_[82071]_  & \new_[82068]_ ;
  assign \new_[82073]_  = \new_[82072]_  & \new_[82065]_ ;
  assign \new_[82076]_  = ~A267 & ~A266;
  assign \new_[82079]_  = A269 & ~A268;
  assign \new_[82080]_  = \new_[82079]_  & \new_[82076]_ ;
  assign \new_[82083]_  = A299 & ~A298;
  assign \new_[82086]_  = A301 & A300;
  assign \new_[82087]_  = \new_[82086]_  & \new_[82083]_ ;
  assign \new_[82088]_  = \new_[82087]_  & \new_[82080]_ ;
  assign \new_[82092]_  = A199 & ~A166;
  assign \new_[82093]_  = ~A167 & \new_[82092]_ ;
  assign \new_[82096]_  = A201 & ~A200;
  assign \new_[82099]_  = A265 & A202;
  assign \new_[82100]_  = \new_[82099]_  & \new_[82096]_ ;
  assign \new_[82101]_  = \new_[82100]_  & \new_[82093]_ ;
  assign \new_[82104]_  = ~A267 & ~A266;
  assign \new_[82107]_  = A269 & ~A268;
  assign \new_[82108]_  = \new_[82107]_  & \new_[82104]_ ;
  assign \new_[82111]_  = A299 & ~A298;
  assign \new_[82114]_  = ~A302 & A300;
  assign \new_[82115]_  = \new_[82114]_  & \new_[82111]_ ;
  assign \new_[82116]_  = \new_[82115]_  & \new_[82108]_ ;
  assign \new_[82120]_  = A199 & ~A166;
  assign \new_[82121]_  = ~A167 & \new_[82120]_ ;
  assign \new_[82124]_  = A201 & ~A200;
  assign \new_[82127]_  = ~A265 & ~A203;
  assign \new_[82128]_  = \new_[82127]_  & \new_[82124]_ ;
  assign \new_[82129]_  = \new_[82128]_  & \new_[82121]_ ;
  assign \new_[82132]_  = A267 & A266;
  assign \new_[82135]_  = A298 & A268;
  assign \new_[82136]_  = \new_[82135]_  & \new_[82132]_ ;
  assign \new_[82139]_  = ~A300 & ~A299;
  assign \new_[82142]_  = A302 & ~A301;
  assign \new_[82143]_  = \new_[82142]_  & \new_[82139]_ ;
  assign \new_[82144]_  = \new_[82143]_  & \new_[82136]_ ;
  assign \new_[82148]_  = A199 & ~A166;
  assign \new_[82149]_  = ~A167 & \new_[82148]_ ;
  assign \new_[82152]_  = A201 & ~A200;
  assign \new_[82155]_  = ~A265 & ~A203;
  assign \new_[82156]_  = \new_[82155]_  & \new_[82152]_ ;
  assign \new_[82157]_  = \new_[82156]_  & \new_[82149]_ ;
  assign \new_[82160]_  = A267 & A266;
  assign \new_[82163]_  = ~A298 & A268;
  assign \new_[82164]_  = \new_[82163]_  & \new_[82160]_ ;
  assign \new_[82167]_  = ~A300 & A299;
  assign \new_[82170]_  = A302 & ~A301;
  assign \new_[82171]_  = \new_[82170]_  & \new_[82167]_ ;
  assign \new_[82172]_  = \new_[82171]_  & \new_[82164]_ ;
  assign \new_[82176]_  = A199 & ~A166;
  assign \new_[82177]_  = ~A167 & \new_[82176]_ ;
  assign \new_[82180]_  = A201 & ~A200;
  assign \new_[82183]_  = ~A265 & ~A203;
  assign \new_[82184]_  = \new_[82183]_  & \new_[82180]_ ;
  assign \new_[82185]_  = \new_[82184]_  & \new_[82177]_ ;
  assign \new_[82188]_  = A267 & A266;
  assign \new_[82191]_  = A298 & ~A269;
  assign \new_[82192]_  = \new_[82191]_  & \new_[82188]_ ;
  assign \new_[82195]_  = ~A300 & ~A299;
  assign \new_[82198]_  = A302 & ~A301;
  assign \new_[82199]_  = \new_[82198]_  & \new_[82195]_ ;
  assign \new_[82200]_  = \new_[82199]_  & \new_[82192]_ ;
  assign \new_[82204]_  = A199 & ~A166;
  assign \new_[82205]_  = ~A167 & \new_[82204]_ ;
  assign \new_[82208]_  = A201 & ~A200;
  assign \new_[82211]_  = ~A265 & ~A203;
  assign \new_[82212]_  = \new_[82211]_  & \new_[82208]_ ;
  assign \new_[82213]_  = \new_[82212]_  & \new_[82205]_ ;
  assign \new_[82216]_  = A267 & A266;
  assign \new_[82219]_  = ~A298 & ~A269;
  assign \new_[82220]_  = \new_[82219]_  & \new_[82216]_ ;
  assign \new_[82223]_  = ~A300 & A299;
  assign \new_[82226]_  = A302 & ~A301;
  assign \new_[82227]_  = \new_[82226]_  & \new_[82223]_ ;
  assign \new_[82228]_  = \new_[82227]_  & \new_[82220]_ ;
  assign \new_[82232]_  = A199 & ~A166;
  assign \new_[82233]_  = ~A167 & \new_[82232]_ ;
  assign \new_[82236]_  = A201 & ~A200;
  assign \new_[82239]_  = ~A265 & ~A203;
  assign \new_[82240]_  = \new_[82239]_  & \new_[82236]_ ;
  assign \new_[82241]_  = \new_[82240]_  & \new_[82233]_ ;
  assign \new_[82244]_  = ~A267 & A266;
  assign \new_[82247]_  = A269 & ~A268;
  assign \new_[82248]_  = \new_[82247]_  & \new_[82244]_ ;
  assign \new_[82251]_  = ~A299 & A298;
  assign \new_[82254]_  = A301 & A300;
  assign \new_[82255]_  = \new_[82254]_  & \new_[82251]_ ;
  assign \new_[82256]_  = \new_[82255]_  & \new_[82248]_ ;
  assign \new_[82260]_  = A199 & ~A166;
  assign \new_[82261]_  = ~A167 & \new_[82260]_ ;
  assign \new_[82264]_  = A201 & ~A200;
  assign \new_[82267]_  = ~A265 & ~A203;
  assign \new_[82268]_  = \new_[82267]_  & \new_[82264]_ ;
  assign \new_[82269]_  = \new_[82268]_  & \new_[82261]_ ;
  assign \new_[82272]_  = ~A267 & A266;
  assign \new_[82275]_  = A269 & ~A268;
  assign \new_[82276]_  = \new_[82275]_  & \new_[82272]_ ;
  assign \new_[82279]_  = ~A299 & A298;
  assign \new_[82282]_  = ~A302 & A300;
  assign \new_[82283]_  = \new_[82282]_  & \new_[82279]_ ;
  assign \new_[82284]_  = \new_[82283]_  & \new_[82276]_ ;
  assign \new_[82288]_  = A199 & ~A166;
  assign \new_[82289]_  = ~A167 & \new_[82288]_ ;
  assign \new_[82292]_  = A201 & ~A200;
  assign \new_[82295]_  = ~A265 & ~A203;
  assign \new_[82296]_  = \new_[82295]_  & \new_[82292]_ ;
  assign \new_[82297]_  = \new_[82296]_  & \new_[82289]_ ;
  assign \new_[82300]_  = ~A267 & A266;
  assign \new_[82303]_  = A269 & ~A268;
  assign \new_[82304]_  = \new_[82303]_  & \new_[82300]_ ;
  assign \new_[82307]_  = A299 & ~A298;
  assign \new_[82310]_  = A301 & A300;
  assign \new_[82311]_  = \new_[82310]_  & \new_[82307]_ ;
  assign \new_[82312]_  = \new_[82311]_  & \new_[82304]_ ;
  assign \new_[82316]_  = A199 & ~A166;
  assign \new_[82317]_  = ~A167 & \new_[82316]_ ;
  assign \new_[82320]_  = A201 & ~A200;
  assign \new_[82323]_  = ~A265 & ~A203;
  assign \new_[82324]_  = \new_[82323]_  & \new_[82320]_ ;
  assign \new_[82325]_  = \new_[82324]_  & \new_[82317]_ ;
  assign \new_[82328]_  = ~A267 & A266;
  assign \new_[82331]_  = A269 & ~A268;
  assign \new_[82332]_  = \new_[82331]_  & \new_[82328]_ ;
  assign \new_[82335]_  = A299 & ~A298;
  assign \new_[82338]_  = ~A302 & A300;
  assign \new_[82339]_  = \new_[82338]_  & \new_[82335]_ ;
  assign \new_[82340]_  = \new_[82339]_  & \new_[82332]_ ;
  assign \new_[82344]_  = A199 & ~A166;
  assign \new_[82345]_  = ~A167 & \new_[82344]_ ;
  assign \new_[82348]_  = A201 & ~A200;
  assign \new_[82351]_  = A265 & ~A203;
  assign \new_[82352]_  = \new_[82351]_  & \new_[82348]_ ;
  assign \new_[82353]_  = \new_[82352]_  & \new_[82345]_ ;
  assign \new_[82356]_  = A267 & ~A266;
  assign \new_[82359]_  = A298 & A268;
  assign \new_[82360]_  = \new_[82359]_  & \new_[82356]_ ;
  assign \new_[82363]_  = ~A300 & ~A299;
  assign \new_[82366]_  = A302 & ~A301;
  assign \new_[82367]_  = \new_[82366]_  & \new_[82363]_ ;
  assign \new_[82368]_  = \new_[82367]_  & \new_[82360]_ ;
  assign \new_[82372]_  = A199 & ~A166;
  assign \new_[82373]_  = ~A167 & \new_[82372]_ ;
  assign \new_[82376]_  = A201 & ~A200;
  assign \new_[82379]_  = A265 & ~A203;
  assign \new_[82380]_  = \new_[82379]_  & \new_[82376]_ ;
  assign \new_[82381]_  = \new_[82380]_  & \new_[82373]_ ;
  assign \new_[82384]_  = A267 & ~A266;
  assign \new_[82387]_  = ~A298 & A268;
  assign \new_[82388]_  = \new_[82387]_  & \new_[82384]_ ;
  assign \new_[82391]_  = ~A300 & A299;
  assign \new_[82394]_  = A302 & ~A301;
  assign \new_[82395]_  = \new_[82394]_  & \new_[82391]_ ;
  assign \new_[82396]_  = \new_[82395]_  & \new_[82388]_ ;
  assign \new_[82400]_  = A199 & ~A166;
  assign \new_[82401]_  = ~A167 & \new_[82400]_ ;
  assign \new_[82404]_  = A201 & ~A200;
  assign \new_[82407]_  = A265 & ~A203;
  assign \new_[82408]_  = \new_[82407]_  & \new_[82404]_ ;
  assign \new_[82409]_  = \new_[82408]_  & \new_[82401]_ ;
  assign \new_[82412]_  = A267 & ~A266;
  assign \new_[82415]_  = A298 & ~A269;
  assign \new_[82416]_  = \new_[82415]_  & \new_[82412]_ ;
  assign \new_[82419]_  = ~A300 & ~A299;
  assign \new_[82422]_  = A302 & ~A301;
  assign \new_[82423]_  = \new_[82422]_  & \new_[82419]_ ;
  assign \new_[82424]_  = \new_[82423]_  & \new_[82416]_ ;
  assign \new_[82428]_  = A199 & ~A166;
  assign \new_[82429]_  = ~A167 & \new_[82428]_ ;
  assign \new_[82432]_  = A201 & ~A200;
  assign \new_[82435]_  = A265 & ~A203;
  assign \new_[82436]_  = \new_[82435]_  & \new_[82432]_ ;
  assign \new_[82437]_  = \new_[82436]_  & \new_[82429]_ ;
  assign \new_[82440]_  = A267 & ~A266;
  assign \new_[82443]_  = ~A298 & ~A269;
  assign \new_[82444]_  = \new_[82443]_  & \new_[82440]_ ;
  assign \new_[82447]_  = ~A300 & A299;
  assign \new_[82450]_  = A302 & ~A301;
  assign \new_[82451]_  = \new_[82450]_  & \new_[82447]_ ;
  assign \new_[82452]_  = \new_[82451]_  & \new_[82444]_ ;
  assign \new_[82456]_  = A199 & ~A166;
  assign \new_[82457]_  = ~A167 & \new_[82456]_ ;
  assign \new_[82460]_  = A201 & ~A200;
  assign \new_[82463]_  = A265 & ~A203;
  assign \new_[82464]_  = \new_[82463]_  & \new_[82460]_ ;
  assign \new_[82465]_  = \new_[82464]_  & \new_[82457]_ ;
  assign \new_[82468]_  = ~A267 & ~A266;
  assign \new_[82471]_  = A269 & ~A268;
  assign \new_[82472]_  = \new_[82471]_  & \new_[82468]_ ;
  assign \new_[82475]_  = ~A299 & A298;
  assign \new_[82478]_  = A301 & A300;
  assign \new_[82479]_  = \new_[82478]_  & \new_[82475]_ ;
  assign \new_[82480]_  = \new_[82479]_  & \new_[82472]_ ;
  assign \new_[82484]_  = A199 & ~A166;
  assign \new_[82485]_  = ~A167 & \new_[82484]_ ;
  assign \new_[82488]_  = A201 & ~A200;
  assign \new_[82491]_  = A265 & ~A203;
  assign \new_[82492]_  = \new_[82491]_  & \new_[82488]_ ;
  assign \new_[82493]_  = \new_[82492]_  & \new_[82485]_ ;
  assign \new_[82496]_  = ~A267 & ~A266;
  assign \new_[82499]_  = A269 & ~A268;
  assign \new_[82500]_  = \new_[82499]_  & \new_[82496]_ ;
  assign \new_[82503]_  = ~A299 & A298;
  assign \new_[82506]_  = ~A302 & A300;
  assign \new_[82507]_  = \new_[82506]_  & \new_[82503]_ ;
  assign \new_[82508]_  = \new_[82507]_  & \new_[82500]_ ;
  assign \new_[82512]_  = A199 & ~A166;
  assign \new_[82513]_  = ~A167 & \new_[82512]_ ;
  assign \new_[82516]_  = A201 & ~A200;
  assign \new_[82519]_  = A265 & ~A203;
  assign \new_[82520]_  = \new_[82519]_  & \new_[82516]_ ;
  assign \new_[82521]_  = \new_[82520]_  & \new_[82513]_ ;
  assign \new_[82524]_  = ~A267 & ~A266;
  assign \new_[82527]_  = A269 & ~A268;
  assign \new_[82528]_  = \new_[82527]_  & \new_[82524]_ ;
  assign \new_[82531]_  = A299 & ~A298;
  assign \new_[82534]_  = A301 & A300;
  assign \new_[82535]_  = \new_[82534]_  & \new_[82531]_ ;
  assign \new_[82536]_  = \new_[82535]_  & \new_[82528]_ ;
  assign \new_[82540]_  = A199 & ~A166;
  assign \new_[82541]_  = ~A167 & \new_[82540]_ ;
  assign \new_[82544]_  = A201 & ~A200;
  assign \new_[82547]_  = A265 & ~A203;
  assign \new_[82548]_  = \new_[82547]_  & \new_[82544]_ ;
  assign \new_[82549]_  = \new_[82548]_  & \new_[82541]_ ;
  assign \new_[82552]_  = ~A267 & ~A266;
  assign \new_[82555]_  = A269 & ~A268;
  assign \new_[82556]_  = \new_[82555]_  & \new_[82552]_ ;
  assign \new_[82559]_  = A299 & ~A298;
  assign \new_[82562]_  = ~A302 & A300;
  assign \new_[82563]_  = \new_[82562]_  & \new_[82559]_ ;
  assign \new_[82564]_  = \new_[82563]_  & \new_[82556]_ ;
  assign \new_[82568]_  = A199 & ~A166;
  assign \new_[82569]_  = ~A167 & \new_[82568]_ ;
  assign \new_[82572]_  = ~A201 & ~A200;
  assign \new_[82575]_  = A203 & ~A202;
  assign \new_[82576]_  = \new_[82575]_  & \new_[82572]_ ;
  assign \new_[82577]_  = \new_[82576]_  & \new_[82569]_ ;
  assign \new_[82580]_  = A266 & ~A265;
  assign \new_[82583]_  = A268 & A267;
  assign \new_[82584]_  = \new_[82583]_  & \new_[82580]_ ;
  assign \new_[82587]_  = ~A299 & A298;
  assign \new_[82590]_  = A301 & A300;
  assign \new_[82591]_  = \new_[82590]_  & \new_[82587]_ ;
  assign \new_[82592]_  = \new_[82591]_  & \new_[82584]_ ;
  assign \new_[82596]_  = A199 & ~A166;
  assign \new_[82597]_  = ~A167 & \new_[82596]_ ;
  assign \new_[82600]_  = ~A201 & ~A200;
  assign \new_[82603]_  = A203 & ~A202;
  assign \new_[82604]_  = \new_[82603]_  & \new_[82600]_ ;
  assign \new_[82605]_  = \new_[82604]_  & \new_[82597]_ ;
  assign \new_[82608]_  = A266 & ~A265;
  assign \new_[82611]_  = A268 & A267;
  assign \new_[82612]_  = \new_[82611]_  & \new_[82608]_ ;
  assign \new_[82615]_  = ~A299 & A298;
  assign \new_[82618]_  = ~A302 & A300;
  assign \new_[82619]_  = \new_[82618]_  & \new_[82615]_ ;
  assign \new_[82620]_  = \new_[82619]_  & \new_[82612]_ ;
  assign \new_[82624]_  = A199 & ~A166;
  assign \new_[82625]_  = ~A167 & \new_[82624]_ ;
  assign \new_[82628]_  = ~A201 & ~A200;
  assign \new_[82631]_  = A203 & ~A202;
  assign \new_[82632]_  = \new_[82631]_  & \new_[82628]_ ;
  assign \new_[82633]_  = \new_[82632]_  & \new_[82625]_ ;
  assign \new_[82636]_  = A266 & ~A265;
  assign \new_[82639]_  = A268 & A267;
  assign \new_[82640]_  = \new_[82639]_  & \new_[82636]_ ;
  assign \new_[82643]_  = A299 & ~A298;
  assign \new_[82646]_  = A301 & A300;
  assign \new_[82647]_  = \new_[82646]_  & \new_[82643]_ ;
  assign \new_[82648]_  = \new_[82647]_  & \new_[82640]_ ;
  assign \new_[82652]_  = A199 & ~A166;
  assign \new_[82653]_  = ~A167 & \new_[82652]_ ;
  assign \new_[82656]_  = ~A201 & ~A200;
  assign \new_[82659]_  = A203 & ~A202;
  assign \new_[82660]_  = \new_[82659]_  & \new_[82656]_ ;
  assign \new_[82661]_  = \new_[82660]_  & \new_[82653]_ ;
  assign \new_[82664]_  = A266 & ~A265;
  assign \new_[82667]_  = A268 & A267;
  assign \new_[82668]_  = \new_[82667]_  & \new_[82664]_ ;
  assign \new_[82671]_  = A299 & ~A298;
  assign \new_[82674]_  = ~A302 & A300;
  assign \new_[82675]_  = \new_[82674]_  & \new_[82671]_ ;
  assign \new_[82676]_  = \new_[82675]_  & \new_[82668]_ ;
  assign \new_[82680]_  = A199 & ~A166;
  assign \new_[82681]_  = ~A167 & \new_[82680]_ ;
  assign \new_[82684]_  = ~A201 & ~A200;
  assign \new_[82687]_  = A203 & ~A202;
  assign \new_[82688]_  = \new_[82687]_  & \new_[82684]_ ;
  assign \new_[82689]_  = \new_[82688]_  & \new_[82681]_ ;
  assign \new_[82692]_  = A266 & ~A265;
  assign \new_[82695]_  = ~A269 & A267;
  assign \new_[82696]_  = \new_[82695]_  & \new_[82692]_ ;
  assign \new_[82699]_  = ~A299 & A298;
  assign \new_[82702]_  = A301 & A300;
  assign \new_[82703]_  = \new_[82702]_  & \new_[82699]_ ;
  assign \new_[82704]_  = \new_[82703]_  & \new_[82696]_ ;
  assign \new_[82708]_  = A199 & ~A166;
  assign \new_[82709]_  = ~A167 & \new_[82708]_ ;
  assign \new_[82712]_  = ~A201 & ~A200;
  assign \new_[82715]_  = A203 & ~A202;
  assign \new_[82716]_  = \new_[82715]_  & \new_[82712]_ ;
  assign \new_[82717]_  = \new_[82716]_  & \new_[82709]_ ;
  assign \new_[82720]_  = A266 & ~A265;
  assign \new_[82723]_  = ~A269 & A267;
  assign \new_[82724]_  = \new_[82723]_  & \new_[82720]_ ;
  assign \new_[82727]_  = ~A299 & A298;
  assign \new_[82730]_  = ~A302 & A300;
  assign \new_[82731]_  = \new_[82730]_  & \new_[82727]_ ;
  assign \new_[82732]_  = \new_[82731]_  & \new_[82724]_ ;
  assign \new_[82736]_  = A199 & ~A166;
  assign \new_[82737]_  = ~A167 & \new_[82736]_ ;
  assign \new_[82740]_  = ~A201 & ~A200;
  assign \new_[82743]_  = A203 & ~A202;
  assign \new_[82744]_  = \new_[82743]_  & \new_[82740]_ ;
  assign \new_[82745]_  = \new_[82744]_  & \new_[82737]_ ;
  assign \new_[82748]_  = A266 & ~A265;
  assign \new_[82751]_  = ~A269 & A267;
  assign \new_[82752]_  = \new_[82751]_  & \new_[82748]_ ;
  assign \new_[82755]_  = A299 & ~A298;
  assign \new_[82758]_  = A301 & A300;
  assign \new_[82759]_  = \new_[82758]_  & \new_[82755]_ ;
  assign \new_[82760]_  = \new_[82759]_  & \new_[82752]_ ;
  assign \new_[82764]_  = A199 & ~A166;
  assign \new_[82765]_  = ~A167 & \new_[82764]_ ;
  assign \new_[82768]_  = ~A201 & ~A200;
  assign \new_[82771]_  = A203 & ~A202;
  assign \new_[82772]_  = \new_[82771]_  & \new_[82768]_ ;
  assign \new_[82773]_  = \new_[82772]_  & \new_[82765]_ ;
  assign \new_[82776]_  = A266 & ~A265;
  assign \new_[82779]_  = ~A269 & A267;
  assign \new_[82780]_  = \new_[82779]_  & \new_[82776]_ ;
  assign \new_[82783]_  = A299 & ~A298;
  assign \new_[82786]_  = ~A302 & A300;
  assign \new_[82787]_  = \new_[82786]_  & \new_[82783]_ ;
  assign \new_[82788]_  = \new_[82787]_  & \new_[82780]_ ;
  assign \new_[82792]_  = A199 & ~A166;
  assign \new_[82793]_  = ~A167 & \new_[82792]_ ;
  assign \new_[82796]_  = ~A201 & ~A200;
  assign \new_[82799]_  = A203 & ~A202;
  assign \new_[82800]_  = \new_[82799]_  & \new_[82796]_ ;
  assign \new_[82801]_  = \new_[82800]_  & \new_[82793]_ ;
  assign \new_[82804]_  = ~A266 & A265;
  assign \new_[82807]_  = A268 & A267;
  assign \new_[82808]_  = \new_[82807]_  & \new_[82804]_ ;
  assign \new_[82811]_  = ~A299 & A298;
  assign \new_[82814]_  = A301 & A300;
  assign \new_[82815]_  = \new_[82814]_  & \new_[82811]_ ;
  assign \new_[82816]_  = \new_[82815]_  & \new_[82808]_ ;
  assign \new_[82820]_  = A199 & ~A166;
  assign \new_[82821]_  = ~A167 & \new_[82820]_ ;
  assign \new_[82824]_  = ~A201 & ~A200;
  assign \new_[82827]_  = A203 & ~A202;
  assign \new_[82828]_  = \new_[82827]_  & \new_[82824]_ ;
  assign \new_[82829]_  = \new_[82828]_  & \new_[82821]_ ;
  assign \new_[82832]_  = ~A266 & A265;
  assign \new_[82835]_  = A268 & A267;
  assign \new_[82836]_  = \new_[82835]_  & \new_[82832]_ ;
  assign \new_[82839]_  = ~A299 & A298;
  assign \new_[82842]_  = ~A302 & A300;
  assign \new_[82843]_  = \new_[82842]_  & \new_[82839]_ ;
  assign \new_[82844]_  = \new_[82843]_  & \new_[82836]_ ;
  assign \new_[82848]_  = A199 & ~A166;
  assign \new_[82849]_  = ~A167 & \new_[82848]_ ;
  assign \new_[82852]_  = ~A201 & ~A200;
  assign \new_[82855]_  = A203 & ~A202;
  assign \new_[82856]_  = \new_[82855]_  & \new_[82852]_ ;
  assign \new_[82857]_  = \new_[82856]_  & \new_[82849]_ ;
  assign \new_[82860]_  = ~A266 & A265;
  assign \new_[82863]_  = A268 & A267;
  assign \new_[82864]_  = \new_[82863]_  & \new_[82860]_ ;
  assign \new_[82867]_  = A299 & ~A298;
  assign \new_[82870]_  = A301 & A300;
  assign \new_[82871]_  = \new_[82870]_  & \new_[82867]_ ;
  assign \new_[82872]_  = \new_[82871]_  & \new_[82864]_ ;
  assign \new_[82876]_  = A199 & ~A166;
  assign \new_[82877]_  = ~A167 & \new_[82876]_ ;
  assign \new_[82880]_  = ~A201 & ~A200;
  assign \new_[82883]_  = A203 & ~A202;
  assign \new_[82884]_  = \new_[82883]_  & \new_[82880]_ ;
  assign \new_[82885]_  = \new_[82884]_  & \new_[82877]_ ;
  assign \new_[82888]_  = ~A266 & A265;
  assign \new_[82891]_  = A268 & A267;
  assign \new_[82892]_  = \new_[82891]_  & \new_[82888]_ ;
  assign \new_[82895]_  = A299 & ~A298;
  assign \new_[82898]_  = ~A302 & A300;
  assign \new_[82899]_  = \new_[82898]_  & \new_[82895]_ ;
  assign \new_[82900]_  = \new_[82899]_  & \new_[82892]_ ;
  assign \new_[82904]_  = A199 & ~A166;
  assign \new_[82905]_  = ~A167 & \new_[82904]_ ;
  assign \new_[82908]_  = ~A201 & ~A200;
  assign \new_[82911]_  = A203 & ~A202;
  assign \new_[82912]_  = \new_[82911]_  & \new_[82908]_ ;
  assign \new_[82913]_  = \new_[82912]_  & \new_[82905]_ ;
  assign \new_[82916]_  = ~A266 & A265;
  assign \new_[82919]_  = ~A269 & A267;
  assign \new_[82920]_  = \new_[82919]_  & \new_[82916]_ ;
  assign \new_[82923]_  = ~A299 & A298;
  assign \new_[82926]_  = A301 & A300;
  assign \new_[82927]_  = \new_[82926]_  & \new_[82923]_ ;
  assign \new_[82928]_  = \new_[82927]_  & \new_[82920]_ ;
  assign \new_[82932]_  = A199 & ~A166;
  assign \new_[82933]_  = ~A167 & \new_[82932]_ ;
  assign \new_[82936]_  = ~A201 & ~A200;
  assign \new_[82939]_  = A203 & ~A202;
  assign \new_[82940]_  = \new_[82939]_  & \new_[82936]_ ;
  assign \new_[82941]_  = \new_[82940]_  & \new_[82933]_ ;
  assign \new_[82944]_  = ~A266 & A265;
  assign \new_[82947]_  = ~A269 & A267;
  assign \new_[82948]_  = \new_[82947]_  & \new_[82944]_ ;
  assign \new_[82951]_  = ~A299 & A298;
  assign \new_[82954]_  = ~A302 & A300;
  assign \new_[82955]_  = \new_[82954]_  & \new_[82951]_ ;
  assign \new_[82956]_  = \new_[82955]_  & \new_[82948]_ ;
  assign \new_[82960]_  = A199 & ~A166;
  assign \new_[82961]_  = ~A167 & \new_[82960]_ ;
  assign \new_[82964]_  = ~A201 & ~A200;
  assign \new_[82967]_  = A203 & ~A202;
  assign \new_[82968]_  = \new_[82967]_  & \new_[82964]_ ;
  assign \new_[82969]_  = \new_[82968]_  & \new_[82961]_ ;
  assign \new_[82972]_  = ~A266 & A265;
  assign \new_[82975]_  = ~A269 & A267;
  assign \new_[82976]_  = \new_[82975]_  & \new_[82972]_ ;
  assign \new_[82979]_  = A299 & ~A298;
  assign \new_[82982]_  = A301 & A300;
  assign \new_[82983]_  = \new_[82982]_  & \new_[82979]_ ;
  assign \new_[82984]_  = \new_[82983]_  & \new_[82976]_ ;
  assign \new_[82988]_  = A199 & ~A166;
  assign \new_[82989]_  = ~A167 & \new_[82988]_ ;
  assign \new_[82992]_  = ~A201 & ~A200;
  assign \new_[82995]_  = A203 & ~A202;
  assign \new_[82996]_  = \new_[82995]_  & \new_[82992]_ ;
  assign \new_[82997]_  = \new_[82996]_  & \new_[82989]_ ;
  assign \new_[83000]_  = ~A266 & A265;
  assign \new_[83003]_  = ~A269 & A267;
  assign \new_[83004]_  = \new_[83003]_  & \new_[83000]_ ;
  assign \new_[83007]_  = A299 & ~A298;
  assign \new_[83010]_  = ~A302 & A300;
  assign \new_[83011]_  = \new_[83010]_  & \new_[83007]_ ;
  assign \new_[83012]_  = \new_[83011]_  & \new_[83004]_ ;
  assign \new_[83016]_  = A167 & A168;
  assign \new_[83017]_  = A170 & \new_[83016]_ ;
  assign \new_[83020]_  = A201 & ~A166;
  assign \new_[83023]_  = A203 & ~A202;
  assign \new_[83024]_  = \new_[83023]_  & \new_[83020]_ ;
  assign \new_[83025]_  = \new_[83024]_  & \new_[83017]_ ;
  assign \new_[83028]_  = ~A268 & A267;
  assign \new_[83031]_  = A298 & A269;
  assign \new_[83032]_  = \new_[83031]_  & \new_[83028]_ ;
  assign \new_[83035]_  = ~A300 & ~A299;
  assign \new_[83038]_  = A302 & ~A301;
  assign \new_[83039]_  = \new_[83038]_  & \new_[83035]_ ;
  assign \new_[83040]_  = \new_[83039]_  & \new_[83032]_ ;
  assign \new_[83044]_  = A167 & A168;
  assign \new_[83045]_  = A170 & \new_[83044]_ ;
  assign \new_[83048]_  = A201 & ~A166;
  assign \new_[83051]_  = A203 & ~A202;
  assign \new_[83052]_  = \new_[83051]_  & \new_[83048]_ ;
  assign \new_[83053]_  = \new_[83052]_  & \new_[83045]_ ;
  assign \new_[83056]_  = ~A268 & A267;
  assign \new_[83059]_  = ~A298 & A269;
  assign \new_[83060]_  = \new_[83059]_  & \new_[83056]_ ;
  assign \new_[83063]_  = ~A300 & A299;
  assign \new_[83066]_  = A302 & ~A301;
  assign \new_[83067]_  = \new_[83066]_  & \new_[83063]_ ;
  assign \new_[83068]_  = \new_[83067]_  & \new_[83060]_ ;
  assign \new_[83072]_  = A167 & A168;
  assign \new_[83073]_  = A170 & \new_[83072]_ ;
  assign \new_[83076]_  = A201 & ~A166;
  assign \new_[83079]_  = A203 & ~A202;
  assign \new_[83080]_  = \new_[83079]_  & \new_[83076]_ ;
  assign \new_[83081]_  = \new_[83080]_  & \new_[83073]_ ;
  assign \new_[83084]_  = A266 & ~A265;
  assign \new_[83087]_  = ~A268 & ~A267;
  assign \new_[83088]_  = \new_[83087]_  & \new_[83084]_ ;
  assign \new_[83091]_  = A300 & A269;
  assign \new_[83094]_  = A302 & ~A301;
  assign \new_[83095]_  = \new_[83094]_  & \new_[83091]_ ;
  assign \new_[83096]_  = \new_[83095]_  & \new_[83088]_ ;
  assign \new_[83100]_  = A167 & A168;
  assign \new_[83101]_  = A170 & \new_[83100]_ ;
  assign \new_[83104]_  = A201 & ~A166;
  assign \new_[83107]_  = A203 & ~A202;
  assign \new_[83108]_  = \new_[83107]_  & \new_[83104]_ ;
  assign \new_[83109]_  = \new_[83108]_  & \new_[83101]_ ;
  assign \new_[83112]_  = ~A266 & A265;
  assign \new_[83115]_  = ~A268 & ~A267;
  assign \new_[83116]_  = \new_[83115]_  & \new_[83112]_ ;
  assign \new_[83119]_  = A300 & A269;
  assign \new_[83122]_  = A302 & ~A301;
  assign \new_[83123]_  = \new_[83122]_  & \new_[83119]_ ;
  assign \new_[83124]_  = \new_[83123]_  & \new_[83116]_ ;
  assign \new_[83128]_  = ~A167 & A168;
  assign \new_[83129]_  = A170 & \new_[83128]_ ;
  assign \new_[83132]_  = A201 & A166;
  assign \new_[83135]_  = A203 & ~A202;
  assign \new_[83136]_  = \new_[83135]_  & \new_[83132]_ ;
  assign \new_[83137]_  = \new_[83136]_  & \new_[83129]_ ;
  assign \new_[83140]_  = ~A268 & A267;
  assign \new_[83143]_  = A298 & A269;
  assign \new_[83144]_  = \new_[83143]_  & \new_[83140]_ ;
  assign \new_[83147]_  = ~A300 & ~A299;
  assign \new_[83150]_  = A302 & ~A301;
  assign \new_[83151]_  = \new_[83150]_  & \new_[83147]_ ;
  assign \new_[83152]_  = \new_[83151]_  & \new_[83144]_ ;
  assign \new_[83156]_  = ~A167 & A168;
  assign \new_[83157]_  = A170 & \new_[83156]_ ;
  assign \new_[83160]_  = A201 & A166;
  assign \new_[83163]_  = A203 & ~A202;
  assign \new_[83164]_  = \new_[83163]_  & \new_[83160]_ ;
  assign \new_[83165]_  = \new_[83164]_  & \new_[83157]_ ;
  assign \new_[83168]_  = ~A268 & A267;
  assign \new_[83171]_  = ~A298 & A269;
  assign \new_[83172]_  = \new_[83171]_  & \new_[83168]_ ;
  assign \new_[83175]_  = ~A300 & A299;
  assign \new_[83178]_  = A302 & ~A301;
  assign \new_[83179]_  = \new_[83178]_  & \new_[83175]_ ;
  assign \new_[83180]_  = \new_[83179]_  & \new_[83172]_ ;
  assign \new_[83184]_  = ~A167 & A168;
  assign \new_[83185]_  = A170 & \new_[83184]_ ;
  assign \new_[83188]_  = A201 & A166;
  assign \new_[83191]_  = A203 & ~A202;
  assign \new_[83192]_  = \new_[83191]_  & \new_[83188]_ ;
  assign \new_[83193]_  = \new_[83192]_  & \new_[83185]_ ;
  assign \new_[83196]_  = A266 & ~A265;
  assign \new_[83199]_  = ~A268 & ~A267;
  assign \new_[83200]_  = \new_[83199]_  & \new_[83196]_ ;
  assign \new_[83203]_  = A300 & A269;
  assign \new_[83206]_  = A302 & ~A301;
  assign \new_[83207]_  = \new_[83206]_  & \new_[83203]_ ;
  assign \new_[83208]_  = \new_[83207]_  & \new_[83200]_ ;
  assign \new_[83212]_  = ~A167 & A168;
  assign \new_[83213]_  = A170 & \new_[83212]_ ;
  assign \new_[83216]_  = A201 & A166;
  assign \new_[83219]_  = A203 & ~A202;
  assign \new_[83220]_  = \new_[83219]_  & \new_[83216]_ ;
  assign \new_[83221]_  = \new_[83220]_  & \new_[83213]_ ;
  assign \new_[83224]_  = ~A266 & A265;
  assign \new_[83227]_  = ~A268 & ~A267;
  assign \new_[83228]_  = \new_[83227]_  & \new_[83224]_ ;
  assign \new_[83231]_  = A300 & A269;
  assign \new_[83234]_  = A302 & ~A301;
  assign \new_[83235]_  = \new_[83234]_  & \new_[83231]_ ;
  assign \new_[83236]_  = \new_[83235]_  & \new_[83228]_ ;
  assign \new_[83240]_  = ~A199 & ~A168;
  assign \new_[83241]_  = A170 & \new_[83240]_ ;
  assign \new_[83244]_  = A201 & A200;
  assign \new_[83247]_  = ~A265 & A202;
  assign \new_[83248]_  = \new_[83247]_  & \new_[83244]_ ;
  assign \new_[83249]_  = \new_[83248]_  & \new_[83241]_ ;
  assign \new_[83252]_  = A267 & A266;
  assign \new_[83255]_  = A298 & A268;
  assign \new_[83256]_  = \new_[83255]_  & \new_[83252]_ ;
  assign \new_[83259]_  = ~A300 & ~A299;
  assign \new_[83262]_  = A302 & ~A301;
  assign \new_[83263]_  = \new_[83262]_  & \new_[83259]_ ;
  assign \new_[83264]_  = \new_[83263]_  & \new_[83256]_ ;
  assign \new_[83268]_  = ~A199 & ~A168;
  assign \new_[83269]_  = A170 & \new_[83268]_ ;
  assign \new_[83272]_  = A201 & A200;
  assign \new_[83275]_  = ~A265 & A202;
  assign \new_[83276]_  = \new_[83275]_  & \new_[83272]_ ;
  assign \new_[83277]_  = \new_[83276]_  & \new_[83269]_ ;
  assign \new_[83280]_  = A267 & A266;
  assign \new_[83283]_  = ~A298 & A268;
  assign \new_[83284]_  = \new_[83283]_  & \new_[83280]_ ;
  assign \new_[83287]_  = ~A300 & A299;
  assign \new_[83290]_  = A302 & ~A301;
  assign \new_[83291]_  = \new_[83290]_  & \new_[83287]_ ;
  assign \new_[83292]_  = \new_[83291]_  & \new_[83284]_ ;
  assign \new_[83296]_  = ~A199 & ~A168;
  assign \new_[83297]_  = A170 & \new_[83296]_ ;
  assign \new_[83300]_  = A201 & A200;
  assign \new_[83303]_  = ~A265 & A202;
  assign \new_[83304]_  = \new_[83303]_  & \new_[83300]_ ;
  assign \new_[83305]_  = \new_[83304]_  & \new_[83297]_ ;
  assign \new_[83308]_  = A267 & A266;
  assign \new_[83311]_  = A298 & ~A269;
  assign \new_[83312]_  = \new_[83311]_  & \new_[83308]_ ;
  assign \new_[83315]_  = ~A300 & ~A299;
  assign \new_[83318]_  = A302 & ~A301;
  assign \new_[83319]_  = \new_[83318]_  & \new_[83315]_ ;
  assign \new_[83320]_  = \new_[83319]_  & \new_[83312]_ ;
  assign \new_[83324]_  = ~A199 & ~A168;
  assign \new_[83325]_  = A170 & \new_[83324]_ ;
  assign \new_[83328]_  = A201 & A200;
  assign \new_[83331]_  = ~A265 & A202;
  assign \new_[83332]_  = \new_[83331]_  & \new_[83328]_ ;
  assign \new_[83333]_  = \new_[83332]_  & \new_[83325]_ ;
  assign \new_[83336]_  = A267 & A266;
  assign \new_[83339]_  = ~A298 & ~A269;
  assign \new_[83340]_  = \new_[83339]_  & \new_[83336]_ ;
  assign \new_[83343]_  = ~A300 & A299;
  assign \new_[83346]_  = A302 & ~A301;
  assign \new_[83347]_  = \new_[83346]_  & \new_[83343]_ ;
  assign \new_[83348]_  = \new_[83347]_  & \new_[83340]_ ;
  assign \new_[83352]_  = ~A199 & ~A168;
  assign \new_[83353]_  = A170 & \new_[83352]_ ;
  assign \new_[83356]_  = A201 & A200;
  assign \new_[83359]_  = ~A265 & A202;
  assign \new_[83360]_  = \new_[83359]_  & \new_[83356]_ ;
  assign \new_[83361]_  = \new_[83360]_  & \new_[83353]_ ;
  assign \new_[83364]_  = ~A267 & A266;
  assign \new_[83367]_  = A269 & ~A268;
  assign \new_[83368]_  = \new_[83367]_  & \new_[83364]_ ;
  assign \new_[83371]_  = ~A299 & A298;
  assign \new_[83374]_  = A301 & A300;
  assign \new_[83375]_  = \new_[83374]_  & \new_[83371]_ ;
  assign \new_[83376]_  = \new_[83375]_  & \new_[83368]_ ;
  assign \new_[83380]_  = ~A199 & ~A168;
  assign \new_[83381]_  = A170 & \new_[83380]_ ;
  assign \new_[83384]_  = A201 & A200;
  assign \new_[83387]_  = ~A265 & A202;
  assign \new_[83388]_  = \new_[83387]_  & \new_[83384]_ ;
  assign \new_[83389]_  = \new_[83388]_  & \new_[83381]_ ;
  assign \new_[83392]_  = ~A267 & A266;
  assign \new_[83395]_  = A269 & ~A268;
  assign \new_[83396]_  = \new_[83395]_  & \new_[83392]_ ;
  assign \new_[83399]_  = ~A299 & A298;
  assign \new_[83402]_  = ~A302 & A300;
  assign \new_[83403]_  = \new_[83402]_  & \new_[83399]_ ;
  assign \new_[83404]_  = \new_[83403]_  & \new_[83396]_ ;
  assign \new_[83408]_  = ~A199 & ~A168;
  assign \new_[83409]_  = A170 & \new_[83408]_ ;
  assign \new_[83412]_  = A201 & A200;
  assign \new_[83415]_  = ~A265 & A202;
  assign \new_[83416]_  = \new_[83415]_  & \new_[83412]_ ;
  assign \new_[83417]_  = \new_[83416]_  & \new_[83409]_ ;
  assign \new_[83420]_  = ~A267 & A266;
  assign \new_[83423]_  = A269 & ~A268;
  assign \new_[83424]_  = \new_[83423]_  & \new_[83420]_ ;
  assign \new_[83427]_  = A299 & ~A298;
  assign \new_[83430]_  = A301 & A300;
  assign \new_[83431]_  = \new_[83430]_  & \new_[83427]_ ;
  assign \new_[83432]_  = \new_[83431]_  & \new_[83424]_ ;
  assign \new_[83436]_  = ~A199 & ~A168;
  assign \new_[83437]_  = A170 & \new_[83436]_ ;
  assign \new_[83440]_  = A201 & A200;
  assign \new_[83443]_  = ~A265 & A202;
  assign \new_[83444]_  = \new_[83443]_  & \new_[83440]_ ;
  assign \new_[83445]_  = \new_[83444]_  & \new_[83437]_ ;
  assign \new_[83448]_  = ~A267 & A266;
  assign \new_[83451]_  = A269 & ~A268;
  assign \new_[83452]_  = \new_[83451]_  & \new_[83448]_ ;
  assign \new_[83455]_  = A299 & ~A298;
  assign \new_[83458]_  = ~A302 & A300;
  assign \new_[83459]_  = \new_[83458]_  & \new_[83455]_ ;
  assign \new_[83460]_  = \new_[83459]_  & \new_[83452]_ ;
  assign \new_[83464]_  = ~A199 & ~A168;
  assign \new_[83465]_  = A170 & \new_[83464]_ ;
  assign \new_[83468]_  = A201 & A200;
  assign \new_[83471]_  = A265 & A202;
  assign \new_[83472]_  = \new_[83471]_  & \new_[83468]_ ;
  assign \new_[83473]_  = \new_[83472]_  & \new_[83465]_ ;
  assign \new_[83476]_  = A267 & ~A266;
  assign \new_[83479]_  = A298 & A268;
  assign \new_[83480]_  = \new_[83479]_  & \new_[83476]_ ;
  assign \new_[83483]_  = ~A300 & ~A299;
  assign \new_[83486]_  = A302 & ~A301;
  assign \new_[83487]_  = \new_[83486]_  & \new_[83483]_ ;
  assign \new_[83488]_  = \new_[83487]_  & \new_[83480]_ ;
  assign \new_[83492]_  = ~A199 & ~A168;
  assign \new_[83493]_  = A170 & \new_[83492]_ ;
  assign \new_[83496]_  = A201 & A200;
  assign \new_[83499]_  = A265 & A202;
  assign \new_[83500]_  = \new_[83499]_  & \new_[83496]_ ;
  assign \new_[83501]_  = \new_[83500]_  & \new_[83493]_ ;
  assign \new_[83504]_  = A267 & ~A266;
  assign \new_[83507]_  = ~A298 & A268;
  assign \new_[83508]_  = \new_[83507]_  & \new_[83504]_ ;
  assign \new_[83511]_  = ~A300 & A299;
  assign \new_[83514]_  = A302 & ~A301;
  assign \new_[83515]_  = \new_[83514]_  & \new_[83511]_ ;
  assign \new_[83516]_  = \new_[83515]_  & \new_[83508]_ ;
  assign \new_[83520]_  = ~A199 & ~A168;
  assign \new_[83521]_  = A170 & \new_[83520]_ ;
  assign \new_[83524]_  = A201 & A200;
  assign \new_[83527]_  = A265 & A202;
  assign \new_[83528]_  = \new_[83527]_  & \new_[83524]_ ;
  assign \new_[83529]_  = \new_[83528]_  & \new_[83521]_ ;
  assign \new_[83532]_  = A267 & ~A266;
  assign \new_[83535]_  = A298 & ~A269;
  assign \new_[83536]_  = \new_[83535]_  & \new_[83532]_ ;
  assign \new_[83539]_  = ~A300 & ~A299;
  assign \new_[83542]_  = A302 & ~A301;
  assign \new_[83543]_  = \new_[83542]_  & \new_[83539]_ ;
  assign \new_[83544]_  = \new_[83543]_  & \new_[83536]_ ;
  assign \new_[83548]_  = ~A199 & ~A168;
  assign \new_[83549]_  = A170 & \new_[83548]_ ;
  assign \new_[83552]_  = A201 & A200;
  assign \new_[83555]_  = A265 & A202;
  assign \new_[83556]_  = \new_[83555]_  & \new_[83552]_ ;
  assign \new_[83557]_  = \new_[83556]_  & \new_[83549]_ ;
  assign \new_[83560]_  = A267 & ~A266;
  assign \new_[83563]_  = ~A298 & ~A269;
  assign \new_[83564]_  = \new_[83563]_  & \new_[83560]_ ;
  assign \new_[83567]_  = ~A300 & A299;
  assign \new_[83570]_  = A302 & ~A301;
  assign \new_[83571]_  = \new_[83570]_  & \new_[83567]_ ;
  assign \new_[83572]_  = \new_[83571]_  & \new_[83564]_ ;
  assign \new_[83576]_  = ~A199 & ~A168;
  assign \new_[83577]_  = A170 & \new_[83576]_ ;
  assign \new_[83580]_  = A201 & A200;
  assign \new_[83583]_  = A265 & A202;
  assign \new_[83584]_  = \new_[83583]_  & \new_[83580]_ ;
  assign \new_[83585]_  = \new_[83584]_  & \new_[83577]_ ;
  assign \new_[83588]_  = ~A267 & ~A266;
  assign \new_[83591]_  = A269 & ~A268;
  assign \new_[83592]_  = \new_[83591]_  & \new_[83588]_ ;
  assign \new_[83595]_  = ~A299 & A298;
  assign \new_[83598]_  = A301 & A300;
  assign \new_[83599]_  = \new_[83598]_  & \new_[83595]_ ;
  assign \new_[83600]_  = \new_[83599]_  & \new_[83592]_ ;
  assign \new_[83604]_  = ~A199 & ~A168;
  assign \new_[83605]_  = A170 & \new_[83604]_ ;
  assign \new_[83608]_  = A201 & A200;
  assign \new_[83611]_  = A265 & A202;
  assign \new_[83612]_  = \new_[83611]_  & \new_[83608]_ ;
  assign \new_[83613]_  = \new_[83612]_  & \new_[83605]_ ;
  assign \new_[83616]_  = ~A267 & ~A266;
  assign \new_[83619]_  = A269 & ~A268;
  assign \new_[83620]_  = \new_[83619]_  & \new_[83616]_ ;
  assign \new_[83623]_  = ~A299 & A298;
  assign \new_[83626]_  = ~A302 & A300;
  assign \new_[83627]_  = \new_[83626]_  & \new_[83623]_ ;
  assign \new_[83628]_  = \new_[83627]_  & \new_[83620]_ ;
  assign \new_[83632]_  = ~A199 & ~A168;
  assign \new_[83633]_  = A170 & \new_[83632]_ ;
  assign \new_[83636]_  = A201 & A200;
  assign \new_[83639]_  = A265 & A202;
  assign \new_[83640]_  = \new_[83639]_  & \new_[83636]_ ;
  assign \new_[83641]_  = \new_[83640]_  & \new_[83633]_ ;
  assign \new_[83644]_  = ~A267 & ~A266;
  assign \new_[83647]_  = A269 & ~A268;
  assign \new_[83648]_  = \new_[83647]_  & \new_[83644]_ ;
  assign \new_[83651]_  = A299 & ~A298;
  assign \new_[83654]_  = A301 & A300;
  assign \new_[83655]_  = \new_[83654]_  & \new_[83651]_ ;
  assign \new_[83656]_  = \new_[83655]_  & \new_[83648]_ ;
  assign \new_[83660]_  = ~A199 & ~A168;
  assign \new_[83661]_  = A170 & \new_[83660]_ ;
  assign \new_[83664]_  = A201 & A200;
  assign \new_[83667]_  = A265 & A202;
  assign \new_[83668]_  = \new_[83667]_  & \new_[83664]_ ;
  assign \new_[83669]_  = \new_[83668]_  & \new_[83661]_ ;
  assign \new_[83672]_  = ~A267 & ~A266;
  assign \new_[83675]_  = A269 & ~A268;
  assign \new_[83676]_  = \new_[83675]_  & \new_[83672]_ ;
  assign \new_[83679]_  = A299 & ~A298;
  assign \new_[83682]_  = ~A302 & A300;
  assign \new_[83683]_  = \new_[83682]_  & \new_[83679]_ ;
  assign \new_[83684]_  = \new_[83683]_  & \new_[83676]_ ;
  assign \new_[83688]_  = ~A199 & ~A168;
  assign \new_[83689]_  = A170 & \new_[83688]_ ;
  assign \new_[83692]_  = A201 & A200;
  assign \new_[83695]_  = ~A265 & ~A203;
  assign \new_[83696]_  = \new_[83695]_  & \new_[83692]_ ;
  assign \new_[83697]_  = \new_[83696]_  & \new_[83689]_ ;
  assign \new_[83700]_  = A267 & A266;
  assign \new_[83703]_  = A298 & A268;
  assign \new_[83704]_  = \new_[83703]_  & \new_[83700]_ ;
  assign \new_[83707]_  = ~A300 & ~A299;
  assign \new_[83710]_  = A302 & ~A301;
  assign \new_[83711]_  = \new_[83710]_  & \new_[83707]_ ;
  assign \new_[83712]_  = \new_[83711]_  & \new_[83704]_ ;
  assign \new_[83716]_  = ~A199 & ~A168;
  assign \new_[83717]_  = A170 & \new_[83716]_ ;
  assign \new_[83720]_  = A201 & A200;
  assign \new_[83723]_  = ~A265 & ~A203;
  assign \new_[83724]_  = \new_[83723]_  & \new_[83720]_ ;
  assign \new_[83725]_  = \new_[83724]_  & \new_[83717]_ ;
  assign \new_[83728]_  = A267 & A266;
  assign \new_[83731]_  = ~A298 & A268;
  assign \new_[83732]_  = \new_[83731]_  & \new_[83728]_ ;
  assign \new_[83735]_  = ~A300 & A299;
  assign \new_[83738]_  = A302 & ~A301;
  assign \new_[83739]_  = \new_[83738]_  & \new_[83735]_ ;
  assign \new_[83740]_  = \new_[83739]_  & \new_[83732]_ ;
  assign \new_[83744]_  = ~A199 & ~A168;
  assign \new_[83745]_  = A170 & \new_[83744]_ ;
  assign \new_[83748]_  = A201 & A200;
  assign \new_[83751]_  = ~A265 & ~A203;
  assign \new_[83752]_  = \new_[83751]_  & \new_[83748]_ ;
  assign \new_[83753]_  = \new_[83752]_  & \new_[83745]_ ;
  assign \new_[83756]_  = A267 & A266;
  assign \new_[83759]_  = A298 & ~A269;
  assign \new_[83760]_  = \new_[83759]_  & \new_[83756]_ ;
  assign \new_[83763]_  = ~A300 & ~A299;
  assign \new_[83766]_  = A302 & ~A301;
  assign \new_[83767]_  = \new_[83766]_  & \new_[83763]_ ;
  assign \new_[83768]_  = \new_[83767]_  & \new_[83760]_ ;
  assign \new_[83772]_  = ~A199 & ~A168;
  assign \new_[83773]_  = A170 & \new_[83772]_ ;
  assign \new_[83776]_  = A201 & A200;
  assign \new_[83779]_  = ~A265 & ~A203;
  assign \new_[83780]_  = \new_[83779]_  & \new_[83776]_ ;
  assign \new_[83781]_  = \new_[83780]_  & \new_[83773]_ ;
  assign \new_[83784]_  = A267 & A266;
  assign \new_[83787]_  = ~A298 & ~A269;
  assign \new_[83788]_  = \new_[83787]_  & \new_[83784]_ ;
  assign \new_[83791]_  = ~A300 & A299;
  assign \new_[83794]_  = A302 & ~A301;
  assign \new_[83795]_  = \new_[83794]_  & \new_[83791]_ ;
  assign \new_[83796]_  = \new_[83795]_  & \new_[83788]_ ;
  assign \new_[83800]_  = ~A199 & ~A168;
  assign \new_[83801]_  = A170 & \new_[83800]_ ;
  assign \new_[83804]_  = A201 & A200;
  assign \new_[83807]_  = ~A265 & ~A203;
  assign \new_[83808]_  = \new_[83807]_  & \new_[83804]_ ;
  assign \new_[83809]_  = \new_[83808]_  & \new_[83801]_ ;
  assign \new_[83812]_  = ~A267 & A266;
  assign \new_[83815]_  = A269 & ~A268;
  assign \new_[83816]_  = \new_[83815]_  & \new_[83812]_ ;
  assign \new_[83819]_  = ~A299 & A298;
  assign \new_[83822]_  = A301 & A300;
  assign \new_[83823]_  = \new_[83822]_  & \new_[83819]_ ;
  assign \new_[83824]_  = \new_[83823]_  & \new_[83816]_ ;
  assign \new_[83828]_  = ~A199 & ~A168;
  assign \new_[83829]_  = A170 & \new_[83828]_ ;
  assign \new_[83832]_  = A201 & A200;
  assign \new_[83835]_  = ~A265 & ~A203;
  assign \new_[83836]_  = \new_[83835]_  & \new_[83832]_ ;
  assign \new_[83837]_  = \new_[83836]_  & \new_[83829]_ ;
  assign \new_[83840]_  = ~A267 & A266;
  assign \new_[83843]_  = A269 & ~A268;
  assign \new_[83844]_  = \new_[83843]_  & \new_[83840]_ ;
  assign \new_[83847]_  = ~A299 & A298;
  assign \new_[83850]_  = ~A302 & A300;
  assign \new_[83851]_  = \new_[83850]_  & \new_[83847]_ ;
  assign \new_[83852]_  = \new_[83851]_  & \new_[83844]_ ;
  assign \new_[83856]_  = ~A199 & ~A168;
  assign \new_[83857]_  = A170 & \new_[83856]_ ;
  assign \new_[83860]_  = A201 & A200;
  assign \new_[83863]_  = ~A265 & ~A203;
  assign \new_[83864]_  = \new_[83863]_  & \new_[83860]_ ;
  assign \new_[83865]_  = \new_[83864]_  & \new_[83857]_ ;
  assign \new_[83868]_  = ~A267 & A266;
  assign \new_[83871]_  = A269 & ~A268;
  assign \new_[83872]_  = \new_[83871]_  & \new_[83868]_ ;
  assign \new_[83875]_  = A299 & ~A298;
  assign \new_[83878]_  = A301 & A300;
  assign \new_[83879]_  = \new_[83878]_  & \new_[83875]_ ;
  assign \new_[83880]_  = \new_[83879]_  & \new_[83872]_ ;
  assign \new_[83884]_  = ~A199 & ~A168;
  assign \new_[83885]_  = A170 & \new_[83884]_ ;
  assign \new_[83888]_  = A201 & A200;
  assign \new_[83891]_  = ~A265 & ~A203;
  assign \new_[83892]_  = \new_[83891]_  & \new_[83888]_ ;
  assign \new_[83893]_  = \new_[83892]_  & \new_[83885]_ ;
  assign \new_[83896]_  = ~A267 & A266;
  assign \new_[83899]_  = A269 & ~A268;
  assign \new_[83900]_  = \new_[83899]_  & \new_[83896]_ ;
  assign \new_[83903]_  = A299 & ~A298;
  assign \new_[83906]_  = ~A302 & A300;
  assign \new_[83907]_  = \new_[83906]_  & \new_[83903]_ ;
  assign \new_[83908]_  = \new_[83907]_  & \new_[83900]_ ;
  assign \new_[83912]_  = ~A199 & ~A168;
  assign \new_[83913]_  = A170 & \new_[83912]_ ;
  assign \new_[83916]_  = A201 & A200;
  assign \new_[83919]_  = A265 & ~A203;
  assign \new_[83920]_  = \new_[83919]_  & \new_[83916]_ ;
  assign \new_[83921]_  = \new_[83920]_  & \new_[83913]_ ;
  assign \new_[83924]_  = A267 & ~A266;
  assign \new_[83927]_  = A298 & A268;
  assign \new_[83928]_  = \new_[83927]_  & \new_[83924]_ ;
  assign \new_[83931]_  = ~A300 & ~A299;
  assign \new_[83934]_  = A302 & ~A301;
  assign \new_[83935]_  = \new_[83934]_  & \new_[83931]_ ;
  assign \new_[83936]_  = \new_[83935]_  & \new_[83928]_ ;
  assign \new_[83940]_  = ~A199 & ~A168;
  assign \new_[83941]_  = A170 & \new_[83940]_ ;
  assign \new_[83944]_  = A201 & A200;
  assign \new_[83947]_  = A265 & ~A203;
  assign \new_[83948]_  = \new_[83947]_  & \new_[83944]_ ;
  assign \new_[83949]_  = \new_[83948]_  & \new_[83941]_ ;
  assign \new_[83952]_  = A267 & ~A266;
  assign \new_[83955]_  = ~A298 & A268;
  assign \new_[83956]_  = \new_[83955]_  & \new_[83952]_ ;
  assign \new_[83959]_  = ~A300 & A299;
  assign \new_[83962]_  = A302 & ~A301;
  assign \new_[83963]_  = \new_[83962]_  & \new_[83959]_ ;
  assign \new_[83964]_  = \new_[83963]_  & \new_[83956]_ ;
  assign \new_[83968]_  = ~A199 & ~A168;
  assign \new_[83969]_  = A170 & \new_[83968]_ ;
  assign \new_[83972]_  = A201 & A200;
  assign \new_[83975]_  = A265 & ~A203;
  assign \new_[83976]_  = \new_[83975]_  & \new_[83972]_ ;
  assign \new_[83977]_  = \new_[83976]_  & \new_[83969]_ ;
  assign \new_[83980]_  = A267 & ~A266;
  assign \new_[83983]_  = A298 & ~A269;
  assign \new_[83984]_  = \new_[83983]_  & \new_[83980]_ ;
  assign \new_[83987]_  = ~A300 & ~A299;
  assign \new_[83990]_  = A302 & ~A301;
  assign \new_[83991]_  = \new_[83990]_  & \new_[83987]_ ;
  assign \new_[83992]_  = \new_[83991]_  & \new_[83984]_ ;
  assign \new_[83996]_  = ~A199 & ~A168;
  assign \new_[83997]_  = A170 & \new_[83996]_ ;
  assign \new_[84000]_  = A201 & A200;
  assign \new_[84003]_  = A265 & ~A203;
  assign \new_[84004]_  = \new_[84003]_  & \new_[84000]_ ;
  assign \new_[84005]_  = \new_[84004]_  & \new_[83997]_ ;
  assign \new_[84008]_  = A267 & ~A266;
  assign \new_[84011]_  = ~A298 & ~A269;
  assign \new_[84012]_  = \new_[84011]_  & \new_[84008]_ ;
  assign \new_[84015]_  = ~A300 & A299;
  assign \new_[84018]_  = A302 & ~A301;
  assign \new_[84019]_  = \new_[84018]_  & \new_[84015]_ ;
  assign \new_[84020]_  = \new_[84019]_  & \new_[84012]_ ;
  assign \new_[84024]_  = ~A199 & ~A168;
  assign \new_[84025]_  = A170 & \new_[84024]_ ;
  assign \new_[84028]_  = A201 & A200;
  assign \new_[84031]_  = A265 & ~A203;
  assign \new_[84032]_  = \new_[84031]_  & \new_[84028]_ ;
  assign \new_[84033]_  = \new_[84032]_  & \new_[84025]_ ;
  assign \new_[84036]_  = ~A267 & ~A266;
  assign \new_[84039]_  = A269 & ~A268;
  assign \new_[84040]_  = \new_[84039]_  & \new_[84036]_ ;
  assign \new_[84043]_  = ~A299 & A298;
  assign \new_[84046]_  = A301 & A300;
  assign \new_[84047]_  = \new_[84046]_  & \new_[84043]_ ;
  assign \new_[84048]_  = \new_[84047]_  & \new_[84040]_ ;
  assign \new_[84052]_  = ~A199 & ~A168;
  assign \new_[84053]_  = A170 & \new_[84052]_ ;
  assign \new_[84056]_  = A201 & A200;
  assign \new_[84059]_  = A265 & ~A203;
  assign \new_[84060]_  = \new_[84059]_  & \new_[84056]_ ;
  assign \new_[84061]_  = \new_[84060]_  & \new_[84053]_ ;
  assign \new_[84064]_  = ~A267 & ~A266;
  assign \new_[84067]_  = A269 & ~A268;
  assign \new_[84068]_  = \new_[84067]_  & \new_[84064]_ ;
  assign \new_[84071]_  = ~A299 & A298;
  assign \new_[84074]_  = ~A302 & A300;
  assign \new_[84075]_  = \new_[84074]_  & \new_[84071]_ ;
  assign \new_[84076]_  = \new_[84075]_  & \new_[84068]_ ;
  assign \new_[84080]_  = ~A199 & ~A168;
  assign \new_[84081]_  = A170 & \new_[84080]_ ;
  assign \new_[84084]_  = A201 & A200;
  assign \new_[84087]_  = A265 & ~A203;
  assign \new_[84088]_  = \new_[84087]_  & \new_[84084]_ ;
  assign \new_[84089]_  = \new_[84088]_  & \new_[84081]_ ;
  assign \new_[84092]_  = ~A267 & ~A266;
  assign \new_[84095]_  = A269 & ~A268;
  assign \new_[84096]_  = \new_[84095]_  & \new_[84092]_ ;
  assign \new_[84099]_  = A299 & ~A298;
  assign \new_[84102]_  = A301 & A300;
  assign \new_[84103]_  = \new_[84102]_  & \new_[84099]_ ;
  assign \new_[84104]_  = \new_[84103]_  & \new_[84096]_ ;
  assign \new_[84108]_  = ~A199 & ~A168;
  assign \new_[84109]_  = A170 & \new_[84108]_ ;
  assign \new_[84112]_  = A201 & A200;
  assign \new_[84115]_  = A265 & ~A203;
  assign \new_[84116]_  = \new_[84115]_  & \new_[84112]_ ;
  assign \new_[84117]_  = \new_[84116]_  & \new_[84109]_ ;
  assign \new_[84120]_  = ~A267 & ~A266;
  assign \new_[84123]_  = A269 & ~A268;
  assign \new_[84124]_  = \new_[84123]_  & \new_[84120]_ ;
  assign \new_[84127]_  = A299 & ~A298;
  assign \new_[84130]_  = ~A302 & A300;
  assign \new_[84131]_  = \new_[84130]_  & \new_[84127]_ ;
  assign \new_[84132]_  = \new_[84131]_  & \new_[84124]_ ;
  assign \new_[84136]_  = ~A199 & ~A168;
  assign \new_[84137]_  = A170 & \new_[84136]_ ;
  assign \new_[84140]_  = ~A201 & A200;
  assign \new_[84143]_  = A203 & ~A202;
  assign \new_[84144]_  = \new_[84143]_  & \new_[84140]_ ;
  assign \new_[84145]_  = \new_[84144]_  & \new_[84137]_ ;
  assign \new_[84148]_  = A266 & ~A265;
  assign \new_[84151]_  = A268 & A267;
  assign \new_[84152]_  = \new_[84151]_  & \new_[84148]_ ;
  assign \new_[84155]_  = ~A299 & A298;
  assign \new_[84158]_  = A301 & A300;
  assign \new_[84159]_  = \new_[84158]_  & \new_[84155]_ ;
  assign \new_[84160]_  = \new_[84159]_  & \new_[84152]_ ;
  assign \new_[84164]_  = ~A199 & ~A168;
  assign \new_[84165]_  = A170 & \new_[84164]_ ;
  assign \new_[84168]_  = ~A201 & A200;
  assign \new_[84171]_  = A203 & ~A202;
  assign \new_[84172]_  = \new_[84171]_  & \new_[84168]_ ;
  assign \new_[84173]_  = \new_[84172]_  & \new_[84165]_ ;
  assign \new_[84176]_  = A266 & ~A265;
  assign \new_[84179]_  = A268 & A267;
  assign \new_[84180]_  = \new_[84179]_  & \new_[84176]_ ;
  assign \new_[84183]_  = ~A299 & A298;
  assign \new_[84186]_  = ~A302 & A300;
  assign \new_[84187]_  = \new_[84186]_  & \new_[84183]_ ;
  assign \new_[84188]_  = \new_[84187]_  & \new_[84180]_ ;
  assign \new_[84192]_  = ~A199 & ~A168;
  assign \new_[84193]_  = A170 & \new_[84192]_ ;
  assign \new_[84196]_  = ~A201 & A200;
  assign \new_[84199]_  = A203 & ~A202;
  assign \new_[84200]_  = \new_[84199]_  & \new_[84196]_ ;
  assign \new_[84201]_  = \new_[84200]_  & \new_[84193]_ ;
  assign \new_[84204]_  = A266 & ~A265;
  assign \new_[84207]_  = A268 & A267;
  assign \new_[84208]_  = \new_[84207]_  & \new_[84204]_ ;
  assign \new_[84211]_  = A299 & ~A298;
  assign \new_[84214]_  = A301 & A300;
  assign \new_[84215]_  = \new_[84214]_  & \new_[84211]_ ;
  assign \new_[84216]_  = \new_[84215]_  & \new_[84208]_ ;
  assign \new_[84220]_  = ~A199 & ~A168;
  assign \new_[84221]_  = A170 & \new_[84220]_ ;
  assign \new_[84224]_  = ~A201 & A200;
  assign \new_[84227]_  = A203 & ~A202;
  assign \new_[84228]_  = \new_[84227]_  & \new_[84224]_ ;
  assign \new_[84229]_  = \new_[84228]_  & \new_[84221]_ ;
  assign \new_[84232]_  = A266 & ~A265;
  assign \new_[84235]_  = A268 & A267;
  assign \new_[84236]_  = \new_[84235]_  & \new_[84232]_ ;
  assign \new_[84239]_  = A299 & ~A298;
  assign \new_[84242]_  = ~A302 & A300;
  assign \new_[84243]_  = \new_[84242]_  & \new_[84239]_ ;
  assign \new_[84244]_  = \new_[84243]_  & \new_[84236]_ ;
  assign \new_[84248]_  = ~A199 & ~A168;
  assign \new_[84249]_  = A170 & \new_[84248]_ ;
  assign \new_[84252]_  = ~A201 & A200;
  assign \new_[84255]_  = A203 & ~A202;
  assign \new_[84256]_  = \new_[84255]_  & \new_[84252]_ ;
  assign \new_[84257]_  = \new_[84256]_  & \new_[84249]_ ;
  assign \new_[84260]_  = A266 & ~A265;
  assign \new_[84263]_  = ~A269 & A267;
  assign \new_[84264]_  = \new_[84263]_  & \new_[84260]_ ;
  assign \new_[84267]_  = ~A299 & A298;
  assign \new_[84270]_  = A301 & A300;
  assign \new_[84271]_  = \new_[84270]_  & \new_[84267]_ ;
  assign \new_[84272]_  = \new_[84271]_  & \new_[84264]_ ;
  assign \new_[84276]_  = ~A199 & ~A168;
  assign \new_[84277]_  = A170 & \new_[84276]_ ;
  assign \new_[84280]_  = ~A201 & A200;
  assign \new_[84283]_  = A203 & ~A202;
  assign \new_[84284]_  = \new_[84283]_  & \new_[84280]_ ;
  assign \new_[84285]_  = \new_[84284]_  & \new_[84277]_ ;
  assign \new_[84288]_  = A266 & ~A265;
  assign \new_[84291]_  = ~A269 & A267;
  assign \new_[84292]_  = \new_[84291]_  & \new_[84288]_ ;
  assign \new_[84295]_  = ~A299 & A298;
  assign \new_[84298]_  = ~A302 & A300;
  assign \new_[84299]_  = \new_[84298]_  & \new_[84295]_ ;
  assign \new_[84300]_  = \new_[84299]_  & \new_[84292]_ ;
  assign \new_[84304]_  = ~A199 & ~A168;
  assign \new_[84305]_  = A170 & \new_[84304]_ ;
  assign \new_[84308]_  = ~A201 & A200;
  assign \new_[84311]_  = A203 & ~A202;
  assign \new_[84312]_  = \new_[84311]_  & \new_[84308]_ ;
  assign \new_[84313]_  = \new_[84312]_  & \new_[84305]_ ;
  assign \new_[84316]_  = A266 & ~A265;
  assign \new_[84319]_  = ~A269 & A267;
  assign \new_[84320]_  = \new_[84319]_  & \new_[84316]_ ;
  assign \new_[84323]_  = A299 & ~A298;
  assign \new_[84326]_  = A301 & A300;
  assign \new_[84327]_  = \new_[84326]_  & \new_[84323]_ ;
  assign \new_[84328]_  = \new_[84327]_  & \new_[84320]_ ;
  assign \new_[84332]_  = ~A199 & ~A168;
  assign \new_[84333]_  = A170 & \new_[84332]_ ;
  assign \new_[84336]_  = ~A201 & A200;
  assign \new_[84339]_  = A203 & ~A202;
  assign \new_[84340]_  = \new_[84339]_  & \new_[84336]_ ;
  assign \new_[84341]_  = \new_[84340]_  & \new_[84333]_ ;
  assign \new_[84344]_  = A266 & ~A265;
  assign \new_[84347]_  = ~A269 & A267;
  assign \new_[84348]_  = \new_[84347]_  & \new_[84344]_ ;
  assign \new_[84351]_  = A299 & ~A298;
  assign \new_[84354]_  = ~A302 & A300;
  assign \new_[84355]_  = \new_[84354]_  & \new_[84351]_ ;
  assign \new_[84356]_  = \new_[84355]_  & \new_[84348]_ ;
  assign \new_[84360]_  = ~A199 & ~A168;
  assign \new_[84361]_  = A170 & \new_[84360]_ ;
  assign \new_[84364]_  = ~A201 & A200;
  assign \new_[84367]_  = A203 & ~A202;
  assign \new_[84368]_  = \new_[84367]_  & \new_[84364]_ ;
  assign \new_[84369]_  = \new_[84368]_  & \new_[84361]_ ;
  assign \new_[84372]_  = ~A266 & A265;
  assign \new_[84375]_  = A268 & A267;
  assign \new_[84376]_  = \new_[84375]_  & \new_[84372]_ ;
  assign \new_[84379]_  = ~A299 & A298;
  assign \new_[84382]_  = A301 & A300;
  assign \new_[84383]_  = \new_[84382]_  & \new_[84379]_ ;
  assign \new_[84384]_  = \new_[84383]_  & \new_[84376]_ ;
  assign \new_[84388]_  = ~A199 & ~A168;
  assign \new_[84389]_  = A170 & \new_[84388]_ ;
  assign \new_[84392]_  = ~A201 & A200;
  assign \new_[84395]_  = A203 & ~A202;
  assign \new_[84396]_  = \new_[84395]_  & \new_[84392]_ ;
  assign \new_[84397]_  = \new_[84396]_  & \new_[84389]_ ;
  assign \new_[84400]_  = ~A266 & A265;
  assign \new_[84403]_  = A268 & A267;
  assign \new_[84404]_  = \new_[84403]_  & \new_[84400]_ ;
  assign \new_[84407]_  = ~A299 & A298;
  assign \new_[84410]_  = ~A302 & A300;
  assign \new_[84411]_  = \new_[84410]_  & \new_[84407]_ ;
  assign \new_[84412]_  = \new_[84411]_  & \new_[84404]_ ;
  assign \new_[84416]_  = ~A199 & ~A168;
  assign \new_[84417]_  = A170 & \new_[84416]_ ;
  assign \new_[84420]_  = ~A201 & A200;
  assign \new_[84423]_  = A203 & ~A202;
  assign \new_[84424]_  = \new_[84423]_  & \new_[84420]_ ;
  assign \new_[84425]_  = \new_[84424]_  & \new_[84417]_ ;
  assign \new_[84428]_  = ~A266 & A265;
  assign \new_[84431]_  = A268 & A267;
  assign \new_[84432]_  = \new_[84431]_  & \new_[84428]_ ;
  assign \new_[84435]_  = A299 & ~A298;
  assign \new_[84438]_  = A301 & A300;
  assign \new_[84439]_  = \new_[84438]_  & \new_[84435]_ ;
  assign \new_[84440]_  = \new_[84439]_  & \new_[84432]_ ;
  assign \new_[84444]_  = ~A199 & ~A168;
  assign \new_[84445]_  = A170 & \new_[84444]_ ;
  assign \new_[84448]_  = ~A201 & A200;
  assign \new_[84451]_  = A203 & ~A202;
  assign \new_[84452]_  = \new_[84451]_  & \new_[84448]_ ;
  assign \new_[84453]_  = \new_[84452]_  & \new_[84445]_ ;
  assign \new_[84456]_  = ~A266 & A265;
  assign \new_[84459]_  = A268 & A267;
  assign \new_[84460]_  = \new_[84459]_  & \new_[84456]_ ;
  assign \new_[84463]_  = A299 & ~A298;
  assign \new_[84466]_  = ~A302 & A300;
  assign \new_[84467]_  = \new_[84466]_  & \new_[84463]_ ;
  assign \new_[84468]_  = \new_[84467]_  & \new_[84460]_ ;
  assign \new_[84472]_  = ~A199 & ~A168;
  assign \new_[84473]_  = A170 & \new_[84472]_ ;
  assign \new_[84476]_  = ~A201 & A200;
  assign \new_[84479]_  = A203 & ~A202;
  assign \new_[84480]_  = \new_[84479]_  & \new_[84476]_ ;
  assign \new_[84481]_  = \new_[84480]_  & \new_[84473]_ ;
  assign \new_[84484]_  = ~A266 & A265;
  assign \new_[84487]_  = ~A269 & A267;
  assign \new_[84488]_  = \new_[84487]_  & \new_[84484]_ ;
  assign \new_[84491]_  = ~A299 & A298;
  assign \new_[84494]_  = A301 & A300;
  assign \new_[84495]_  = \new_[84494]_  & \new_[84491]_ ;
  assign \new_[84496]_  = \new_[84495]_  & \new_[84488]_ ;
  assign \new_[84500]_  = ~A199 & ~A168;
  assign \new_[84501]_  = A170 & \new_[84500]_ ;
  assign \new_[84504]_  = ~A201 & A200;
  assign \new_[84507]_  = A203 & ~A202;
  assign \new_[84508]_  = \new_[84507]_  & \new_[84504]_ ;
  assign \new_[84509]_  = \new_[84508]_  & \new_[84501]_ ;
  assign \new_[84512]_  = ~A266 & A265;
  assign \new_[84515]_  = ~A269 & A267;
  assign \new_[84516]_  = \new_[84515]_  & \new_[84512]_ ;
  assign \new_[84519]_  = ~A299 & A298;
  assign \new_[84522]_  = ~A302 & A300;
  assign \new_[84523]_  = \new_[84522]_  & \new_[84519]_ ;
  assign \new_[84524]_  = \new_[84523]_  & \new_[84516]_ ;
  assign \new_[84528]_  = ~A199 & ~A168;
  assign \new_[84529]_  = A170 & \new_[84528]_ ;
  assign \new_[84532]_  = ~A201 & A200;
  assign \new_[84535]_  = A203 & ~A202;
  assign \new_[84536]_  = \new_[84535]_  & \new_[84532]_ ;
  assign \new_[84537]_  = \new_[84536]_  & \new_[84529]_ ;
  assign \new_[84540]_  = ~A266 & A265;
  assign \new_[84543]_  = ~A269 & A267;
  assign \new_[84544]_  = \new_[84543]_  & \new_[84540]_ ;
  assign \new_[84547]_  = A299 & ~A298;
  assign \new_[84550]_  = A301 & A300;
  assign \new_[84551]_  = \new_[84550]_  & \new_[84547]_ ;
  assign \new_[84552]_  = \new_[84551]_  & \new_[84544]_ ;
  assign \new_[84556]_  = ~A199 & ~A168;
  assign \new_[84557]_  = A170 & \new_[84556]_ ;
  assign \new_[84560]_  = ~A201 & A200;
  assign \new_[84563]_  = A203 & ~A202;
  assign \new_[84564]_  = \new_[84563]_  & \new_[84560]_ ;
  assign \new_[84565]_  = \new_[84564]_  & \new_[84557]_ ;
  assign \new_[84568]_  = ~A266 & A265;
  assign \new_[84571]_  = ~A269 & A267;
  assign \new_[84572]_  = \new_[84571]_  & \new_[84568]_ ;
  assign \new_[84575]_  = A299 & ~A298;
  assign \new_[84578]_  = ~A302 & A300;
  assign \new_[84579]_  = \new_[84578]_  & \new_[84575]_ ;
  assign \new_[84580]_  = \new_[84579]_  & \new_[84572]_ ;
  assign \new_[84584]_  = A199 & ~A168;
  assign \new_[84585]_  = A170 & \new_[84584]_ ;
  assign \new_[84588]_  = A201 & ~A200;
  assign \new_[84591]_  = ~A265 & A202;
  assign \new_[84592]_  = \new_[84591]_  & \new_[84588]_ ;
  assign \new_[84593]_  = \new_[84592]_  & \new_[84585]_ ;
  assign \new_[84596]_  = A267 & A266;
  assign \new_[84599]_  = A298 & A268;
  assign \new_[84600]_  = \new_[84599]_  & \new_[84596]_ ;
  assign \new_[84603]_  = ~A300 & ~A299;
  assign \new_[84606]_  = A302 & ~A301;
  assign \new_[84607]_  = \new_[84606]_  & \new_[84603]_ ;
  assign \new_[84608]_  = \new_[84607]_  & \new_[84600]_ ;
  assign \new_[84612]_  = A199 & ~A168;
  assign \new_[84613]_  = A170 & \new_[84612]_ ;
  assign \new_[84616]_  = A201 & ~A200;
  assign \new_[84619]_  = ~A265 & A202;
  assign \new_[84620]_  = \new_[84619]_  & \new_[84616]_ ;
  assign \new_[84621]_  = \new_[84620]_  & \new_[84613]_ ;
  assign \new_[84624]_  = A267 & A266;
  assign \new_[84627]_  = ~A298 & A268;
  assign \new_[84628]_  = \new_[84627]_  & \new_[84624]_ ;
  assign \new_[84631]_  = ~A300 & A299;
  assign \new_[84634]_  = A302 & ~A301;
  assign \new_[84635]_  = \new_[84634]_  & \new_[84631]_ ;
  assign \new_[84636]_  = \new_[84635]_  & \new_[84628]_ ;
  assign \new_[84640]_  = A199 & ~A168;
  assign \new_[84641]_  = A170 & \new_[84640]_ ;
  assign \new_[84644]_  = A201 & ~A200;
  assign \new_[84647]_  = ~A265 & A202;
  assign \new_[84648]_  = \new_[84647]_  & \new_[84644]_ ;
  assign \new_[84649]_  = \new_[84648]_  & \new_[84641]_ ;
  assign \new_[84652]_  = A267 & A266;
  assign \new_[84655]_  = A298 & ~A269;
  assign \new_[84656]_  = \new_[84655]_  & \new_[84652]_ ;
  assign \new_[84659]_  = ~A300 & ~A299;
  assign \new_[84662]_  = A302 & ~A301;
  assign \new_[84663]_  = \new_[84662]_  & \new_[84659]_ ;
  assign \new_[84664]_  = \new_[84663]_  & \new_[84656]_ ;
  assign \new_[84668]_  = A199 & ~A168;
  assign \new_[84669]_  = A170 & \new_[84668]_ ;
  assign \new_[84672]_  = A201 & ~A200;
  assign \new_[84675]_  = ~A265 & A202;
  assign \new_[84676]_  = \new_[84675]_  & \new_[84672]_ ;
  assign \new_[84677]_  = \new_[84676]_  & \new_[84669]_ ;
  assign \new_[84680]_  = A267 & A266;
  assign \new_[84683]_  = ~A298 & ~A269;
  assign \new_[84684]_  = \new_[84683]_  & \new_[84680]_ ;
  assign \new_[84687]_  = ~A300 & A299;
  assign \new_[84690]_  = A302 & ~A301;
  assign \new_[84691]_  = \new_[84690]_  & \new_[84687]_ ;
  assign \new_[84692]_  = \new_[84691]_  & \new_[84684]_ ;
  assign \new_[84696]_  = A199 & ~A168;
  assign \new_[84697]_  = A170 & \new_[84696]_ ;
  assign \new_[84700]_  = A201 & ~A200;
  assign \new_[84703]_  = ~A265 & A202;
  assign \new_[84704]_  = \new_[84703]_  & \new_[84700]_ ;
  assign \new_[84705]_  = \new_[84704]_  & \new_[84697]_ ;
  assign \new_[84708]_  = ~A267 & A266;
  assign \new_[84711]_  = A269 & ~A268;
  assign \new_[84712]_  = \new_[84711]_  & \new_[84708]_ ;
  assign \new_[84715]_  = ~A299 & A298;
  assign \new_[84718]_  = A301 & A300;
  assign \new_[84719]_  = \new_[84718]_  & \new_[84715]_ ;
  assign \new_[84720]_  = \new_[84719]_  & \new_[84712]_ ;
  assign \new_[84724]_  = A199 & ~A168;
  assign \new_[84725]_  = A170 & \new_[84724]_ ;
  assign \new_[84728]_  = A201 & ~A200;
  assign \new_[84731]_  = ~A265 & A202;
  assign \new_[84732]_  = \new_[84731]_  & \new_[84728]_ ;
  assign \new_[84733]_  = \new_[84732]_  & \new_[84725]_ ;
  assign \new_[84736]_  = ~A267 & A266;
  assign \new_[84739]_  = A269 & ~A268;
  assign \new_[84740]_  = \new_[84739]_  & \new_[84736]_ ;
  assign \new_[84743]_  = ~A299 & A298;
  assign \new_[84746]_  = ~A302 & A300;
  assign \new_[84747]_  = \new_[84746]_  & \new_[84743]_ ;
  assign \new_[84748]_  = \new_[84747]_  & \new_[84740]_ ;
  assign \new_[84752]_  = A199 & ~A168;
  assign \new_[84753]_  = A170 & \new_[84752]_ ;
  assign \new_[84756]_  = A201 & ~A200;
  assign \new_[84759]_  = ~A265 & A202;
  assign \new_[84760]_  = \new_[84759]_  & \new_[84756]_ ;
  assign \new_[84761]_  = \new_[84760]_  & \new_[84753]_ ;
  assign \new_[84764]_  = ~A267 & A266;
  assign \new_[84767]_  = A269 & ~A268;
  assign \new_[84768]_  = \new_[84767]_  & \new_[84764]_ ;
  assign \new_[84771]_  = A299 & ~A298;
  assign \new_[84774]_  = A301 & A300;
  assign \new_[84775]_  = \new_[84774]_  & \new_[84771]_ ;
  assign \new_[84776]_  = \new_[84775]_  & \new_[84768]_ ;
  assign \new_[84780]_  = A199 & ~A168;
  assign \new_[84781]_  = A170 & \new_[84780]_ ;
  assign \new_[84784]_  = A201 & ~A200;
  assign \new_[84787]_  = ~A265 & A202;
  assign \new_[84788]_  = \new_[84787]_  & \new_[84784]_ ;
  assign \new_[84789]_  = \new_[84788]_  & \new_[84781]_ ;
  assign \new_[84792]_  = ~A267 & A266;
  assign \new_[84795]_  = A269 & ~A268;
  assign \new_[84796]_  = \new_[84795]_  & \new_[84792]_ ;
  assign \new_[84799]_  = A299 & ~A298;
  assign \new_[84802]_  = ~A302 & A300;
  assign \new_[84803]_  = \new_[84802]_  & \new_[84799]_ ;
  assign \new_[84804]_  = \new_[84803]_  & \new_[84796]_ ;
  assign \new_[84808]_  = A199 & ~A168;
  assign \new_[84809]_  = A170 & \new_[84808]_ ;
  assign \new_[84812]_  = A201 & ~A200;
  assign \new_[84815]_  = A265 & A202;
  assign \new_[84816]_  = \new_[84815]_  & \new_[84812]_ ;
  assign \new_[84817]_  = \new_[84816]_  & \new_[84809]_ ;
  assign \new_[84820]_  = A267 & ~A266;
  assign \new_[84823]_  = A298 & A268;
  assign \new_[84824]_  = \new_[84823]_  & \new_[84820]_ ;
  assign \new_[84827]_  = ~A300 & ~A299;
  assign \new_[84830]_  = A302 & ~A301;
  assign \new_[84831]_  = \new_[84830]_  & \new_[84827]_ ;
  assign \new_[84832]_  = \new_[84831]_  & \new_[84824]_ ;
  assign \new_[84836]_  = A199 & ~A168;
  assign \new_[84837]_  = A170 & \new_[84836]_ ;
  assign \new_[84840]_  = A201 & ~A200;
  assign \new_[84843]_  = A265 & A202;
  assign \new_[84844]_  = \new_[84843]_  & \new_[84840]_ ;
  assign \new_[84845]_  = \new_[84844]_  & \new_[84837]_ ;
  assign \new_[84848]_  = A267 & ~A266;
  assign \new_[84851]_  = ~A298 & A268;
  assign \new_[84852]_  = \new_[84851]_  & \new_[84848]_ ;
  assign \new_[84855]_  = ~A300 & A299;
  assign \new_[84858]_  = A302 & ~A301;
  assign \new_[84859]_  = \new_[84858]_  & \new_[84855]_ ;
  assign \new_[84860]_  = \new_[84859]_  & \new_[84852]_ ;
  assign \new_[84864]_  = A199 & ~A168;
  assign \new_[84865]_  = A170 & \new_[84864]_ ;
  assign \new_[84868]_  = A201 & ~A200;
  assign \new_[84871]_  = A265 & A202;
  assign \new_[84872]_  = \new_[84871]_  & \new_[84868]_ ;
  assign \new_[84873]_  = \new_[84872]_  & \new_[84865]_ ;
  assign \new_[84876]_  = A267 & ~A266;
  assign \new_[84879]_  = A298 & ~A269;
  assign \new_[84880]_  = \new_[84879]_  & \new_[84876]_ ;
  assign \new_[84883]_  = ~A300 & ~A299;
  assign \new_[84886]_  = A302 & ~A301;
  assign \new_[84887]_  = \new_[84886]_  & \new_[84883]_ ;
  assign \new_[84888]_  = \new_[84887]_  & \new_[84880]_ ;
  assign \new_[84892]_  = A199 & ~A168;
  assign \new_[84893]_  = A170 & \new_[84892]_ ;
  assign \new_[84896]_  = A201 & ~A200;
  assign \new_[84899]_  = A265 & A202;
  assign \new_[84900]_  = \new_[84899]_  & \new_[84896]_ ;
  assign \new_[84901]_  = \new_[84900]_  & \new_[84893]_ ;
  assign \new_[84904]_  = A267 & ~A266;
  assign \new_[84907]_  = ~A298 & ~A269;
  assign \new_[84908]_  = \new_[84907]_  & \new_[84904]_ ;
  assign \new_[84911]_  = ~A300 & A299;
  assign \new_[84914]_  = A302 & ~A301;
  assign \new_[84915]_  = \new_[84914]_  & \new_[84911]_ ;
  assign \new_[84916]_  = \new_[84915]_  & \new_[84908]_ ;
  assign \new_[84920]_  = A199 & ~A168;
  assign \new_[84921]_  = A170 & \new_[84920]_ ;
  assign \new_[84924]_  = A201 & ~A200;
  assign \new_[84927]_  = A265 & A202;
  assign \new_[84928]_  = \new_[84927]_  & \new_[84924]_ ;
  assign \new_[84929]_  = \new_[84928]_  & \new_[84921]_ ;
  assign \new_[84932]_  = ~A267 & ~A266;
  assign \new_[84935]_  = A269 & ~A268;
  assign \new_[84936]_  = \new_[84935]_  & \new_[84932]_ ;
  assign \new_[84939]_  = ~A299 & A298;
  assign \new_[84942]_  = A301 & A300;
  assign \new_[84943]_  = \new_[84942]_  & \new_[84939]_ ;
  assign \new_[84944]_  = \new_[84943]_  & \new_[84936]_ ;
  assign \new_[84948]_  = A199 & ~A168;
  assign \new_[84949]_  = A170 & \new_[84948]_ ;
  assign \new_[84952]_  = A201 & ~A200;
  assign \new_[84955]_  = A265 & A202;
  assign \new_[84956]_  = \new_[84955]_  & \new_[84952]_ ;
  assign \new_[84957]_  = \new_[84956]_  & \new_[84949]_ ;
  assign \new_[84960]_  = ~A267 & ~A266;
  assign \new_[84963]_  = A269 & ~A268;
  assign \new_[84964]_  = \new_[84963]_  & \new_[84960]_ ;
  assign \new_[84967]_  = ~A299 & A298;
  assign \new_[84970]_  = ~A302 & A300;
  assign \new_[84971]_  = \new_[84970]_  & \new_[84967]_ ;
  assign \new_[84972]_  = \new_[84971]_  & \new_[84964]_ ;
  assign \new_[84976]_  = A199 & ~A168;
  assign \new_[84977]_  = A170 & \new_[84976]_ ;
  assign \new_[84980]_  = A201 & ~A200;
  assign \new_[84983]_  = A265 & A202;
  assign \new_[84984]_  = \new_[84983]_  & \new_[84980]_ ;
  assign \new_[84985]_  = \new_[84984]_  & \new_[84977]_ ;
  assign \new_[84988]_  = ~A267 & ~A266;
  assign \new_[84991]_  = A269 & ~A268;
  assign \new_[84992]_  = \new_[84991]_  & \new_[84988]_ ;
  assign \new_[84995]_  = A299 & ~A298;
  assign \new_[84998]_  = A301 & A300;
  assign \new_[84999]_  = \new_[84998]_  & \new_[84995]_ ;
  assign \new_[85000]_  = \new_[84999]_  & \new_[84992]_ ;
  assign \new_[85004]_  = A199 & ~A168;
  assign \new_[85005]_  = A170 & \new_[85004]_ ;
  assign \new_[85008]_  = A201 & ~A200;
  assign \new_[85011]_  = A265 & A202;
  assign \new_[85012]_  = \new_[85011]_  & \new_[85008]_ ;
  assign \new_[85013]_  = \new_[85012]_  & \new_[85005]_ ;
  assign \new_[85016]_  = ~A267 & ~A266;
  assign \new_[85019]_  = A269 & ~A268;
  assign \new_[85020]_  = \new_[85019]_  & \new_[85016]_ ;
  assign \new_[85023]_  = A299 & ~A298;
  assign \new_[85026]_  = ~A302 & A300;
  assign \new_[85027]_  = \new_[85026]_  & \new_[85023]_ ;
  assign \new_[85028]_  = \new_[85027]_  & \new_[85020]_ ;
  assign \new_[85032]_  = A199 & ~A168;
  assign \new_[85033]_  = A170 & \new_[85032]_ ;
  assign \new_[85036]_  = A201 & ~A200;
  assign \new_[85039]_  = ~A265 & ~A203;
  assign \new_[85040]_  = \new_[85039]_  & \new_[85036]_ ;
  assign \new_[85041]_  = \new_[85040]_  & \new_[85033]_ ;
  assign \new_[85044]_  = A267 & A266;
  assign \new_[85047]_  = A298 & A268;
  assign \new_[85048]_  = \new_[85047]_  & \new_[85044]_ ;
  assign \new_[85051]_  = ~A300 & ~A299;
  assign \new_[85054]_  = A302 & ~A301;
  assign \new_[85055]_  = \new_[85054]_  & \new_[85051]_ ;
  assign \new_[85056]_  = \new_[85055]_  & \new_[85048]_ ;
  assign \new_[85060]_  = A199 & ~A168;
  assign \new_[85061]_  = A170 & \new_[85060]_ ;
  assign \new_[85064]_  = A201 & ~A200;
  assign \new_[85067]_  = ~A265 & ~A203;
  assign \new_[85068]_  = \new_[85067]_  & \new_[85064]_ ;
  assign \new_[85069]_  = \new_[85068]_  & \new_[85061]_ ;
  assign \new_[85072]_  = A267 & A266;
  assign \new_[85075]_  = ~A298 & A268;
  assign \new_[85076]_  = \new_[85075]_  & \new_[85072]_ ;
  assign \new_[85079]_  = ~A300 & A299;
  assign \new_[85082]_  = A302 & ~A301;
  assign \new_[85083]_  = \new_[85082]_  & \new_[85079]_ ;
  assign \new_[85084]_  = \new_[85083]_  & \new_[85076]_ ;
  assign \new_[85088]_  = A199 & ~A168;
  assign \new_[85089]_  = A170 & \new_[85088]_ ;
  assign \new_[85092]_  = A201 & ~A200;
  assign \new_[85095]_  = ~A265 & ~A203;
  assign \new_[85096]_  = \new_[85095]_  & \new_[85092]_ ;
  assign \new_[85097]_  = \new_[85096]_  & \new_[85089]_ ;
  assign \new_[85100]_  = A267 & A266;
  assign \new_[85103]_  = A298 & ~A269;
  assign \new_[85104]_  = \new_[85103]_  & \new_[85100]_ ;
  assign \new_[85107]_  = ~A300 & ~A299;
  assign \new_[85110]_  = A302 & ~A301;
  assign \new_[85111]_  = \new_[85110]_  & \new_[85107]_ ;
  assign \new_[85112]_  = \new_[85111]_  & \new_[85104]_ ;
  assign \new_[85116]_  = A199 & ~A168;
  assign \new_[85117]_  = A170 & \new_[85116]_ ;
  assign \new_[85120]_  = A201 & ~A200;
  assign \new_[85123]_  = ~A265 & ~A203;
  assign \new_[85124]_  = \new_[85123]_  & \new_[85120]_ ;
  assign \new_[85125]_  = \new_[85124]_  & \new_[85117]_ ;
  assign \new_[85128]_  = A267 & A266;
  assign \new_[85131]_  = ~A298 & ~A269;
  assign \new_[85132]_  = \new_[85131]_  & \new_[85128]_ ;
  assign \new_[85135]_  = ~A300 & A299;
  assign \new_[85138]_  = A302 & ~A301;
  assign \new_[85139]_  = \new_[85138]_  & \new_[85135]_ ;
  assign \new_[85140]_  = \new_[85139]_  & \new_[85132]_ ;
  assign \new_[85144]_  = A199 & ~A168;
  assign \new_[85145]_  = A170 & \new_[85144]_ ;
  assign \new_[85148]_  = A201 & ~A200;
  assign \new_[85151]_  = ~A265 & ~A203;
  assign \new_[85152]_  = \new_[85151]_  & \new_[85148]_ ;
  assign \new_[85153]_  = \new_[85152]_  & \new_[85145]_ ;
  assign \new_[85156]_  = ~A267 & A266;
  assign \new_[85159]_  = A269 & ~A268;
  assign \new_[85160]_  = \new_[85159]_  & \new_[85156]_ ;
  assign \new_[85163]_  = ~A299 & A298;
  assign \new_[85166]_  = A301 & A300;
  assign \new_[85167]_  = \new_[85166]_  & \new_[85163]_ ;
  assign \new_[85168]_  = \new_[85167]_  & \new_[85160]_ ;
  assign \new_[85172]_  = A199 & ~A168;
  assign \new_[85173]_  = A170 & \new_[85172]_ ;
  assign \new_[85176]_  = A201 & ~A200;
  assign \new_[85179]_  = ~A265 & ~A203;
  assign \new_[85180]_  = \new_[85179]_  & \new_[85176]_ ;
  assign \new_[85181]_  = \new_[85180]_  & \new_[85173]_ ;
  assign \new_[85184]_  = ~A267 & A266;
  assign \new_[85187]_  = A269 & ~A268;
  assign \new_[85188]_  = \new_[85187]_  & \new_[85184]_ ;
  assign \new_[85191]_  = ~A299 & A298;
  assign \new_[85194]_  = ~A302 & A300;
  assign \new_[85195]_  = \new_[85194]_  & \new_[85191]_ ;
  assign \new_[85196]_  = \new_[85195]_  & \new_[85188]_ ;
  assign \new_[85200]_  = A199 & ~A168;
  assign \new_[85201]_  = A170 & \new_[85200]_ ;
  assign \new_[85204]_  = A201 & ~A200;
  assign \new_[85207]_  = ~A265 & ~A203;
  assign \new_[85208]_  = \new_[85207]_  & \new_[85204]_ ;
  assign \new_[85209]_  = \new_[85208]_  & \new_[85201]_ ;
  assign \new_[85212]_  = ~A267 & A266;
  assign \new_[85215]_  = A269 & ~A268;
  assign \new_[85216]_  = \new_[85215]_  & \new_[85212]_ ;
  assign \new_[85219]_  = A299 & ~A298;
  assign \new_[85222]_  = A301 & A300;
  assign \new_[85223]_  = \new_[85222]_  & \new_[85219]_ ;
  assign \new_[85224]_  = \new_[85223]_  & \new_[85216]_ ;
  assign \new_[85228]_  = A199 & ~A168;
  assign \new_[85229]_  = A170 & \new_[85228]_ ;
  assign \new_[85232]_  = A201 & ~A200;
  assign \new_[85235]_  = ~A265 & ~A203;
  assign \new_[85236]_  = \new_[85235]_  & \new_[85232]_ ;
  assign \new_[85237]_  = \new_[85236]_  & \new_[85229]_ ;
  assign \new_[85240]_  = ~A267 & A266;
  assign \new_[85243]_  = A269 & ~A268;
  assign \new_[85244]_  = \new_[85243]_  & \new_[85240]_ ;
  assign \new_[85247]_  = A299 & ~A298;
  assign \new_[85250]_  = ~A302 & A300;
  assign \new_[85251]_  = \new_[85250]_  & \new_[85247]_ ;
  assign \new_[85252]_  = \new_[85251]_  & \new_[85244]_ ;
  assign \new_[85256]_  = A199 & ~A168;
  assign \new_[85257]_  = A170 & \new_[85256]_ ;
  assign \new_[85260]_  = A201 & ~A200;
  assign \new_[85263]_  = A265 & ~A203;
  assign \new_[85264]_  = \new_[85263]_  & \new_[85260]_ ;
  assign \new_[85265]_  = \new_[85264]_  & \new_[85257]_ ;
  assign \new_[85268]_  = A267 & ~A266;
  assign \new_[85271]_  = A298 & A268;
  assign \new_[85272]_  = \new_[85271]_  & \new_[85268]_ ;
  assign \new_[85275]_  = ~A300 & ~A299;
  assign \new_[85278]_  = A302 & ~A301;
  assign \new_[85279]_  = \new_[85278]_  & \new_[85275]_ ;
  assign \new_[85280]_  = \new_[85279]_  & \new_[85272]_ ;
  assign \new_[85284]_  = A199 & ~A168;
  assign \new_[85285]_  = A170 & \new_[85284]_ ;
  assign \new_[85288]_  = A201 & ~A200;
  assign \new_[85291]_  = A265 & ~A203;
  assign \new_[85292]_  = \new_[85291]_  & \new_[85288]_ ;
  assign \new_[85293]_  = \new_[85292]_  & \new_[85285]_ ;
  assign \new_[85296]_  = A267 & ~A266;
  assign \new_[85299]_  = ~A298 & A268;
  assign \new_[85300]_  = \new_[85299]_  & \new_[85296]_ ;
  assign \new_[85303]_  = ~A300 & A299;
  assign \new_[85306]_  = A302 & ~A301;
  assign \new_[85307]_  = \new_[85306]_  & \new_[85303]_ ;
  assign \new_[85308]_  = \new_[85307]_  & \new_[85300]_ ;
  assign \new_[85312]_  = A199 & ~A168;
  assign \new_[85313]_  = A170 & \new_[85312]_ ;
  assign \new_[85316]_  = A201 & ~A200;
  assign \new_[85319]_  = A265 & ~A203;
  assign \new_[85320]_  = \new_[85319]_  & \new_[85316]_ ;
  assign \new_[85321]_  = \new_[85320]_  & \new_[85313]_ ;
  assign \new_[85324]_  = A267 & ~A266;
  assign \new_[85327]_  = A298 & ~A269;
  assign \new_[85328]_  = \new_[85327]_  & \new_[85324]_ ;
  assign \new_[85331]_  = ~A300 & ~A299;
  assign \new_[85334]_  = A302 & ~A301;
  assign \new_[85335]_  = \new_[85334]_  & \new_[85331]_ ;
  assign \new_[85336]_  = \new_[85335]_  & \new_[85328]_ ;
  assign \new_[85340]_  = A199 & ~A168;
  assign \new_[85341]_  = A170 & \new_[85340]_ ;
  assign \new_[85344]_  = A201 & ~A200;
  assign \new_[85347]_  = A265 & ~A203;
  assign \new_[85348]_  = \new_[85347]_  & \new_[85344]_ ;
  assign \new_[85349]_  = \new_[85348]_  & \new_[85341]_ ;
  assign \new_[85352]_  = A267 & ~A266;
  assign \new_[85355]_  = ~A298 & ~A269;
  assign \new_[85356]_  = \new_[85355]_  & \new_[85352]_ ;
  assign \new_[85359]_  = ~A300 & A299;
  assign \new_[85362]_  = A302 & ~A301;
  assign \new_[85363]_  = \new_[85362]_  & \new_[85359]_ ;
  assign \new_[85364]_  = \new_[85363]_  & \new_[85356]_ ;
  assign \new_[85368]_  = A199 & ~A168;
  assign \new_[85369]_  = A170 & \new_[85368]_ ;
  assign \new_[85372]_  = A201 & ~A200;
  assign \new_[85375]_  = A265 & ~A203;
  assign \new_[85376]_  = \new_[85375]_  & \new_[85372]_ ;
  assign \new_[85377]_  = \new_[85376]_  & \new_[85369]_ ;
  assign \new_[85380]_  = ~A267 & ~A266;
  assign \new_[85383]_  = A269 & ~A268;
  assign \new_[85384]_  = \new_[85383]_  & \new_[85380]_ ;
  assign \new_[85387]_  = ~A299 & A298;
  assign \new_[85390]_  = A301 & A300;
  assign \new_[85391]_  = \new_[85390]_  & \new_[85387]_ ;
  assign \new_[85392]_  = \new_[85391]_  & \new_[85384]_ ;
  assign \new_[85396]_  = A199 & ~A168;
  assign \new_[85397]_  = A170 & \new_[85396]_ ;
  assign \new_[85400]_  = A201 & ~A200;
  assign \new_[85403]_  = A265 & ~A203;
  assign \new_[85404]_  = \new_[85403]_  & \new_[85400]_ ;
  assign \new_[85405]_  = \new_[85404]_  & \new_[85397]_ ;
  assign \new_[85408]_  = ~A267 & ~A266;
  assign \new_[85411]_  = A269 & ~A268;
  assign \new_[85412]_  = \new_[85411]_  & \new_[85408]_ ;
  assign \new_[85415]_  = ~A299 & A298;
  assign \new_[85418]_  = ~A302 & A300;
  assign \new_[85419]_  = \new_[85418]_  & \new_[85415]_ ;
  assign \new_[85420]_  = \new_[85419]_  & \new_[85412]_ ;
  assign \new_[85424]_  = A199 & ~A168;
  assign \new_[85425]_  = A170 & \new_[85424]_ ;
  assign \new_[85428]_  = A201 & ~A200;
  assign \new_[85431]_  = A265 & ~A203;
  assign \new_[85432]_  = \new_[85431]_  & \new_[85428]_ ;
  assign \new_[85433]_  = \new_[85432]_  & \new_[85425]_ ;
  assign \new_[85436]_  = ~A267 & ~A266;
  assign \new_[85439]_  = A269 & ~A268;
  assign \new_[85440]_  = \new_[85439]_  & \new_[85436]_ ;
  assign \new_[85443]_  = A299 & ~A298;
  assign \new_[85446]_  = A301 & A300;
  assign \new_[85447]_  = \new_[85446]_  & \new_[85443]_ ;
  assign \new_[85448]_  = \new_[85447]_  & \new_[85440]_ ;
  assign \new_[85452]_  = A199 & ~A168;
  assign \new_[85453]_  = A170 & \new_[85452]_ ;
  assign \new_[85456]_  = A201 & ~A200;
  assign \new_[85459]_  = A265 & ~A203;
  assign \new_[85460]_  = \new_[85459]_  & \new_[85456]_ ;
  assign \new_[85461]_  = \new_[85460]_  & \new_[85453]_ ;
  assign \new_[85464]_  = ~A267 & ~A266;
  assign \new_[85467]_  = A269 & ~A268;
  assign \new_[85468]_  = \new_[85467]_  & \new_[85464]_ ;
  assign \new_[85471]_  = A299 & ~A298;
  assign \new_[85474]_  = ~A302 & A300;
  assign \new_[85475]_  = \new_[85474]_  & \new_[85471]_ ;
  assign \new_[85476]_  = \new_[85475]_  & \new_[85468]_ ;
  assign \new_[85480]_  = A199 & ~A168;
  assign \new_[85481]_  = A170 & \new_[85480]_ ;
  assign \new_[85484]_  = ~A201 & ~A200;
  assign \new_[85487]_  = A203 & ~A202;
  assign \new_[85488]_  = \new_[85487]_  & \new_[85484]_ ;
  assign \new_[85489]_  = \new_[85488]_  & \new_[85481]_ ;
  assign \new_[85492]_  = A266 & ~A265;
  assign \new_[85495]_  = A268 & A267;
  assign \new_[85496]_  = \new_[85495]_  & \new_[85492]_ ;
  assign \new_[85499]_  = ~A299 & A298;
  assign \new_[85502]_  = A301 & A300;
  assign \new_[85503]_  = \new_[85502]_  & \new_[85499]_ ;
  assign \new_[85504]_  = \new_[85503]_  & \new_[85496]_ ;
  assign \new_[85508]_  = A199 & ~A168;
  assign \new_[85509]_  = A170 & \new_[85508]_ ;
  assign \new_[85512]_  = ~A201 & ~A200;
  assign \new_[85515]_  = A203 & ~A202;
  assign \new_[85516]_  = \new_[85515]_  & \new_[85512]_ ;
  assign \new_[85517]_  = \new_[85516]_  & \new_[85509]_ ;
  assign \new_[85520]_  = A266 & ~A265;
  assign \new_[85523]_  = A268 & A267;
  assign \new_[85524]_  = \new_[85523]_  & \new_[85520]_ ;
  assign \new_[85527]_  = ~A299 & A298;
  assign \new_[85530]_  = ~A302 & A300;
  assign \new_[85531]_  = \new_[85530]_  & \new_[85527]_ ;
  assign \new_[85532]_  = \new_[85531]_  & \new_[85524]_ ;
  assign \new_[85536]_  = A199 & ~A168;
  assign \new_[85537]_  = A170 & \new_[85536]_ ;
  assign \new_[85540]_  = ~A201 & ~A200;
  assign \new_[85543]_  = A203 & ~A202;
  assign \new_[85544]_  = \new_[85543]_  & \new_[85540]_ ;
  assign \new_[85545]_  = \new_[85544]_  & \new_[85537]_ ;
  assign \new_[85548]_  = A266 & ~A265;
  assign \new_[85551]_  = A268 & A267;
  assign \new_[85552]_  = \new_[85551]_  & \new_[85548]_ ;
  assign \new_[85555]_  = A299 & ~A298;
  assign \new_[85558]_  = A301 & A300;
  assign \new_[85559]_  = \new_[85558]_  & \new_[85555]_ ;
  assign \new_[85560]_  = \new_[85559]_  & \new_[85552]_ ;
  assign \new_[85564]_  = A199 & ~A168;
  assign \new_[85565]_  = A170 & \new_[85564]_ ;
  assign \new_[85568]_  = ~A201 & ~A200;
  assign \new_[85571]_  = A203 & ~A202;
  assign \new_[85572]_  = \new_[85571]_  & \new_[85568]_ ;
  assign \new_[85573]_  = \new_[85572]_  & \new_[85565]_ ;
  assign \new_[85576]_  = A266 & ~A265;
  assign \new_[85579]_  = A268 & A267;
  assign \new_[85580]_  = \new_[85579]_  & \new_[85576]_ ;
  assign \new_[85583]_  = A299 & ~A298;
  assign \new_[85586]_  = ~A302 & A300;
  assign \new_[85587]_  = \new_[85586]_  & \new_[85583]_ ;
  assign \new_[85588]_  = \new_[85587]_  & \new_[85580]_ ;
  assign \new_[85592]_  = A199 & ~A168;
  assign \new_[85593]_  = A170 & \new_[85592]_ ;
  assign \new_[85596]_  = ~A201 & ~A200;
  assign \new_[85599]_  = A203 & ~A202;
  assign \new_[85600]_  = \new_[85599]_  & \new_[85596]_ ;
  assign \new_[85601]_  = \new_[85600]_  & \new_[85593]_ ;
  assign \new_[85604]_  = A266 & ~A265;
  assign \new_[85607]_  = ~A269 & A267;
  assign \new_[85608]_  = \new_[85607]_  & \new_[85604]_ ;
  assign \new_[85611]_  = ~A299 & A298;
  assign \new_[85614]_  = A301 & A300;
  assign \new_[85615]_  = \new_[85614]_  & \new_[85611]_ ;
  assign \new_[85616]_  = \new_[85615]_  & \new_[85608]_ ;
  assign \new_[85620]_  = A199 & ~A168;
  assign \new_[85621]_  = A170 & \new_[85620]_ ;
  assign \new_[85624]_  = ~A201 & ~A200;
  assign \new_[85627]_  = A203 & ~A202;
  assign \new_[85628]_  = \new_[85627]_  & \new_[85624]_ ;
  assign \new_[85629]_  = \new_[85628]_  & \new_[85621]_ ;
  assign \new_[85632]_  = A266 & ~A265;
  assign \new_[85635]_  = ~A269 & A267;
  assign \new_[85636]_  = \new_[85635]_  & \new_[85632]_ ;
  assign \new_[85639]_  = ~A299 & A298;
  assign \new_[85642]_  = ~A302 & A300;
  assign \new_[85643]_  = \new_[85642]_  & \new_[85639]_ ;
  assign \new_[85644]_  = \new_[85643]_  & \new_[85636]_ ;
  assign \new_[85648]_  = A199 & ~A168;
  assign \new_[85649]_  = A170 & \new_[85648]_ ;
  assign \new_[85652]_  = ~A201 & ~A200;
  assign \new_[85655]_  = A203 & ~A202;
  assign \new_[85656]_  = \new_[85655]_  & \new_[85652]_ ;
  assign \new_[85657]_  = \new_[85656]_  & \new_[85649]_ ;
  assign \new_[85660]_  = A266 & ~A265;
  assign \new_[85663]_  = ~A269 & A267;
  assign \new_[85664]_  = \new_[85663]_  & \new_[85660]_ ;
  assign \new_[85667]_  = A299 & ~A298;
  assign \new_[85670]_  = A301 & A300;
  assign \new_[85671]_  = \new_[85670]_  & \new_[85667]_ ;
  assign \new_[85672]_  = \new_[85671]_  & \new_[85664]_ ;
  assign \new_[85676]_  = A199 & ~A168;
  assign \new_[85677]_  = A170 & \new_[85676]_ ;
  assign \new_[85680]_  = ~A201 & ~A200;
  assign \new_[85683]_  = A203 & ~A202;
  assign \new_[85684]_  = \new_[85683]_  & \new_[85680]_ ;
  assign \new_[85685]_  = \new_[85684]_  & \new_[85677]_ ;
  assign \new_[85688]_  = A266 & ~A265;
  assign \new_[85691]_  = ~A269 & A267;
  assign \new_[85692]_  = \new_[85691]_  & \new_[85688]_ ;
  assign \new_[85695]_  = A299 & ~A298;
  assign \new_[85698]_  = ~A302 & A300;
  assign \new_[85699]_  = \new_[85698]_  & \new_[85695]_ ;
  assign \new_[85700]_  = \new_[85699]_  & \new_[85692]_ ;
  assign \new_[85704]_  = A199 & ~A168;
  assign \new_[85705]_  = A170 & \new_[85704]_ ;
  assign \new_[85708]_  = ~A201 & ~A200;
  assign \new_[85711]_  = A203 & ~A202;
  assign \new_[85712]_  = \new_[85711]_  & \new_[85708]_ ;
  assign \new_[85713]_  = \new_[85712]_  & \new_[85705]_ ;
  assign \new_[85716]_  = ~A266 & A265;
  assign \new_[85719]_  = A268 & A267;
  assign \new_[85720]_  = \new_[85719]_  & \new_[85716]_ ;
  assign \new_[85723]_  = ~A299 & A298;
  assign \new_[85726]_  = A301 & A300;
  assign \new_[85727]_  = \new_[85726]_  & \new_[85723]_ ;
  assign \new_[85728]_  = \new_[85727]_  & \new_[85720]_ ;
  assign \new_[85732]_  = A199 & ~A168;
  assign \new_[85733]_  = A170 & \new_[85732]_ ;
  assign \new_[85736]_  = ~A201 & ~A200;
  assign \new_[85739]_  = A203 & ~A202;
  assign \new_[85740]_  = \new_[85739]_  & \new_[85736]_ ;
  assign \new_[85741]_  = \new_[85740]_  & \new_[85733]_ ;
  assign \new_[85744]_  = ~A266 & A265;
  assign \new_[85747]_  = A268 & A267;
  assign \new_[85748]_  = \new_[85747]_  & \new_[85744]_ ;
  assign \new_[85751]_  = ~A299 & A298;
  assign \new_[85754]_  = ~A302 & A300;
  assign \new_[85755]_  = \new_[85754]_  & \new_[85751]_ ;
  assign \new_[85756]_  = \new_[85755]_  & \new_[85748]_ ;
  assign \new_[85760]_  = A199 & ~A168;
  assign \new_[85761]_  = A170 & \new_[85760]_ ;
  assign \new_[85764]_  = ~A201 & ~A200;
  assign \new_[85767]_  = A203 & ~A202;
  assign \new_[85768]_  = \new_[85767]_  & \new_[85764]_ ;
  assign \new_[85769]_  = \new_[85768]_  & \new_[85761]_ ;
  assign \new_[85772]_  = ~A266 & A265;
  assign \new_[85775]_  = A268 & A267;
  assign \new_[85776]_  = \new_[85775]_  & \new_[85772]_ ;
  assign \new_[85779]_  = A299 & ~A298;
  assign \new_[85782]_  = A301 & A300;
  assign \new_[85783]_  = \new_[85782]_  & \new_[85779]_ ;
  assign \new_[85784]_  = \new_[85783]_  & \new_[85776]_ ;
  assign \new_[85788]_  = A199 & ~A168;
  assign \new_[85789]_  = A170 & \new_[85788]_ ;
  assign \new_[85792]_  = ~A201 & ~A200;
  assign \new_[85795]_  = A203 & ~A202;
  assign \new_[85796]_  = \new_[85795]_  & \new_[85792]_ ;
  assign \new_[85797]_  = \new_[85796]_  & \new_[85789]_ ;
  assign \new_[85800]_  = ~A266 & A265;
  assign \new_[85803]_  = A268 & A267;
  assign \new_[85804]_  = \new_[85803]_  & \new_[85800]_ ;
  assign \new_[85807]_  = A299 & ~A298;
  assign \new_[85810]_  = ~A302 & A300;
  assign \new_[85811]_  = \new_[85810]_  & \new_[85807]_ ;
  assign \new_[85812]_  = \new_[85811]_  & \new_[85804]_ ;
  assign \new_[85816]_  = A199 & ~A168;
  assign \new_[85817]_  = A170 & \new_[85816]_ ;
  assign \new_[85820]_  = ~A201 & ~A200;
  assign \new_[85823]_  = A203 & ~A202;
  assign \new_[85824]_  = \new_[85823]_  & \new_[85820]_ ;
  assign \new_[85825]_  = \new_[85824]_  & \new_[85817]_ ;
  assign \new_[85828]_  = ~A266 & A265;
  assign \new_[85831]_  = ~A269 & A267;
  assign \new_[85832]_  = \new_[85831]_  & \new_[85828]_ ;
  assign \new_[85835]_  = ~A299 & A298;
  assign \new_[85838]_  = A301 & A300;
  assign \new_[85839]_  = \new_[85838]_  & \new_[85835]_ ;
  assign \new_[85840]_  = \new_[85839]_  & \new_[85832]_ ;
  assign \new_[85844]_  = A199 & ~A168;
  assign \new_[85845]_  = A170 & \new_[85844]_ ;
  assign \new_[85848]_  = ~A201 & ~A200;
  assign \new_[85851]_  = A203 & ~A202;
  assign \new_[85852]_  = \new_[85851]_  & \new_[85848]_ ;
  assign \new_[85853]_  = \new_[85852]_  & \new_[85845]_ ;
  assign \new_[85856]_  = ~A266 & A265;
  assign \new_[85859]_  = ~A269 & A267;
  assign \new_[85860]_  = \new_[85859]_  & \new_[85856]_ ;
  assign \new_[85863]_  = ~A299 & A298;
  assign \new_[85866]_  = ~A302 & A300;
  assign \new_[85867]_  = \new_[85866]_  & \new_[85863]_ ;
  assign \new_[85868]_  = \new_[85867]_  & \new_[85860]_ ;
  assign \new_[85872]_  = A199 & ~A168;
  assign \new_[85873]_  = A170 & \new_[85872]_ ;
  assign \new_[85876]_  = ~A201 & ~A200;
  assign \new_[85879]_  = A203 & ~A202;
  assign \new_[85880]_  = \new_[85879]_  & \new_[85876]_ ;
  assign \new_[85881]_  = \new_[85880]_  & \new_[85873]_ ;
  assign \new_[85884]_  = ~A266 & A265;
  assign \new_[85887]_  = ~A269 & A267;
  assign \new_[85888]_  = \new_[85887]_  & \new_[85884]_ ;
  assign \new_[85891]_  = A299 & ~A298;
  assign \new_[85894]_  = A301 & A300;
  assign \new_[85895]_  = \new_[85894]_  & \new_[85891]_ ;
  assign \new_[85896]_  = \new_[85895]_  & \new_[85888]_ ;
  assign \new_[85900]_  = A199 & ~A168;
  assign \new_[85901]_  = A170 & \new_[85900]_ ;
  assign \new_[85904]_  = ~A201 & ~A200;
  assign \new_[85907]_  = A203 & ~A202;
  assign \new_[85908]_  = \new_[85907]_  & \new_[85904]_ ;
  assign \new_[85909]_  = \new_[85908]_  & \new_[85901]_ ;
  assign \new_[85912]_  = ~A266 & A265;
  assign \new_[85915]_  = ~A269 & A267;
  assign \new_[85916]_  = \new_[85915]_  & \new_[85912]_ ;
  assign \new_[85919]_  = A299 & ~A298;
  assign \new_[85922]_  = ~A302 & A300;
  assign \new_[85923]_  = \new_[85922]_  & \new_[85919]_ ;
  assign \new_[85924]_  = \new_[85923]_  & \new_[85916]_ ;
  assign \new_[85928]_  = A167 & A168;
  assign \new_[85929]_  = A169 & \new_[85928]_ ;
  assign \new_[85932]_  = A201 & ~A166;
  assign \new_[85935]_  = A203 & ~A202;
  assign \new_[85936]_  = \new_[85935]_  & \new_[85932]_ ;
  assign \new_[85937]_  = \new_[85936]_  & \new_[85929]_ ;
  assign \new_[85940]_  = ~A268 & A267;
  assign \new_[85943]_  = A298 & A269;
  assign \new_[85944]_  = \new_[85943]_  & \new_[85940]_ ;
  assign \new_[85947]_  = ~A300 & ~A299;
  assign \new_[85950]_  = A302 & ~A301;
  assign \new_[85951]_  = \new_[85950]_  & \new_[85947]_ ;
  assign \new_[85952]_  = \new_[85951]_  & \new_[85944]_ ;
  assign \new_[85956]_  = A167 & A168;
  assign \new_[85957]_  = A169 & \new_[85956]_ ;
  assign \new_[85960]_  = A201 & ~A166;
  assign \new_[85963]_  = A203 & ~A202;
  assign \new_[85964]_  = \new_[85963]_  & \new_[85960]_ ;
  assign \new_[85965]_  = \new_[85964]_  & \new_[85957]_ ;
  assign \new_[85968]_  = ~A268 & A267;
  assign \new_[85971]_  = ~A298 & A269;
  assign \new_[85972]_  = \new_[85971]_  & \new_[85968]_ ;
  assign \new_[85975]_  = ~A300 & A299;
  assign \new_[85978]_  = A302 & ~A301;
  assign \new_[85979]_  = \new_[85978]_  & \new_[85975]_ ;
  assign \new_[85980]_  = \new_[85979]_  & \new_[85972]_ ;
  assign \new_[85984]_  = A167 & A168;
  assign \new_[85985]_  = A169 & \new_[85984]_ ;
  assign \new_[85988]_  = A201 & ~A166;
  assign \new_[85991]_  = A203 & ~A202;
  assign \new_[85992]_  = \new_[85991]_  & \new_[85988]_ ;
  assign \new_[85993]_  = \new_[85992]_  & \new_[85985]_ ;
  assign \new_[85996]_  = A266 & ~A265;
  assign \new_[85999]_  = ~A268 & ~A267;
  assign \new_[86000]_  = \new_[85999]_  & \new_[85996]_ ;
  assign \new_[86003]_  = A300 & A269;
  assign \new_[86006]_  = A302 & ~A301;
  assign \new_[86007]_  = \new_[86006]_  & \new_[86003]_ ;
  assign \new_[86008]_  = \new_[86007]_  & \new_[86000]_ ;
  assign \new_[86012]_  = A167 & A168;
  assign \new_[86013]_  = A169 & \new_[86012]_ ;
  assign \new_[86016]_  = A201 & ~A166;
  assign \new_[86019]_  = A203 & ~A202;
  assign \new_[86020]_  = \new_[86019]_  & \new_[86016]_ ;
  assign \new_[86021]_  = \new_[86020]_  & \new_[86013]_ ;
  assign \new_[86024]_  = ~A266 & A265;
  assign \new_[86027]_  = ~A268 & ~A267;
  assign \new_[86028]_  = \new_[86027]_  & \new_[86024]_ ;
  assign \new_[86031]_  = A300 & A269;
  assign \new_[86034]_  = A302 & ~A301;
  assign \new_[86035]_  = \new_[86034]_  & \new_[86031]_ ;
  assign \new_[86036]_  = \new_[86035]_  & \new_[86028]_ ;
  assign \new_[86040]_  = ~A167 & A168;
  assign \new_[86041]_  = A169 & \new_[86040]_ ;
  assign \new_[86044]_  = A201 & A166;
  assign \new_[86047]_  = A203 & ~A202;
  assign \new_[86048]_  = \new_[86047]_  & \new_[86044]_ ;
  assign \new_[86049]_  = \new_[86048]_  & \new_[86041]_ ;
  assign \new_[86052]_  = ~A268 & A267;
  assign \new_[86055]_  = A298 & A269;
  assign \new_[86056]_  = \new_[86055]_  & \new_[86052]_ ;
  assign \new_[86059]_  = ~A300 & ~A299;
  assign \new_[86062]_  = A302 & ~A301;
  assign \new_[86063]_  = \new_[86062]_  & \new_[86059]_ ;
  assign \new_[86064]_  = \new_[86063]_  & \new_[86056]_ ;
  assign \new_[86068]_  = ~A167 & A168;
  assign \new_[86069]_  = A169 & \new_[86068]_ ;
  assign \new_[86072]_  = A201 & A166;
  assign \new_[86075]_  = A203 & ~A202;
  assign \new_[86076]_  = \new_[86075]_  & \new_[86072]_ ;
  assign \new_[86077]_  = \new_[86076]_  & \new_[86069]_ ;
  assign \new_[86080]_  = ~A268 & A267;
  assign \new_[86083]_  = ~A298 & A269;
  assign \new_[86084]_  = \new_[86083]_  & \new_[86080]_ ;
  assign \new_[86087]_  = ~A300 & A299;
  assign \new_[86090]_  = A302 & ~A301;
  assign \new_[86091]_  = \new_[86090]_  & \new_[86087]_ ;
  assign \new_[86092]_  = \new_[86091]_  & \new_[86084]_ ;
  assign \new_[86096]_  = ~A167 & A168;
  assign \new_[86097]_  = A169 & \new_[86096]_ ;
  assign \new_[86100]_  = A201 & A166;
  assign \new_[86103]_  = A203 & ~A202;
  assign \new_[86104]_  = \new_[86103]_  & \new_[86100]_ ;
  assign \new_[86105]_  = \new_[86104]_  & \new_[86097]_ ;
  assign \new_[86108]_  = A266 & ~A265;
  assign \new_[86111]_  = ~A268 & ~A267;
  assign \new_[86112]_  = \new_[86111]_  & \new_[86108]_ ;
  assign \new_[86115]_  = A300 & A269;
  assign \new_[86118]_  = A302 & ~A301;
  assign \new_[86119]_  = \new_[86118]_  & \new_[86115]_ ;
  assign \new_[86120]_  = \new_[86119]_  & \new_[86112]_ ;
  assign \new_[86124]_  = ~A167 & A168;
  assign \new_[86125]_  = A169 & \new_[86124]_ ;
  assign \new_[86128]_  = A201 & A166;
  assign \new_[86131]_  = A203 & ~A202;
  assign \new_[86132]_  = \new_[86131]_  & \new_[86128]_ ;
  assign \new_[86133]_  = \new_[86132]_  & \new_[86125]_ ;
  assign \new_[86136]_  = ~A266 & A265;
  assign \new_[86139]_  = ~A268 & ~A267;
  assign \new_[86140]_  = \new_[86139]_  & \new_[86136]_ ;
  assign \new_[86143]_  = A300 & A269;
  assign \new_[86146]_  = A302 & ~A301;
  assign \new_[86147]_  = \new_[86146]_  & \new_[86143]_ ;
  assign \new_[86148]_  = \new_[86147]_  & \new_[86140]_ ;
  assign \new_[86152]_  = ~A199 & ~A168;
  assign \new_[86153]_  = A169 & \new_[86152]_ ;
  assign \new_[86156]_  = A201 & A200;
  assign \new_[86159]_  = ~A265 & A202;
  assign \new_[86160]_  = \new_[86159]_  & \new_[86156]_ ;
  assign \new_[86161]_  = \new_[86160]_  & \new_[86153]_ ;
  assign \new_[86164]_  = A267 & A266;
  assign \new_[86167]_  = A298 & A268;
  assign \new_[86168]_  = \new_[86167]_  & \new_[86164]_ ;
  assign \new_[86171]_  = ~A300 & ~A299;
  assign \new_[86174]_  = A302 & ~A301;
  assign \new_[86175]_  = \new_[86174]_  & \new_[86171]_ ;
  assign \new_[86176]_  = \new_[86175]_  & \new_[86168]_ ;
  assign \new_[86180]_  = ~A199 & ~A168;
  assign \new_[86181]_  = A169 & \new_[86180]_ ;
  assign \new_[86184]_  = A201 & A200;
  assign \new_[86187]_  = ~A265 & A202;
  assign \new_[86188]_  = \new_[86187]_  & \new_[86184]_ ;
  assign \new_[86189]_  = \new_[86188]_  & \new_[86181]_ ;
  assign \new_[86192]_  = A267 & A266;
  assign \new_[86195]_  = ~A298 & A268;
  assign \new_[86196]_  = \new_[86195]_  & \new_[86192]_ ;
  assign \new_[86199]_  = ~A300 & A299;
  assign \new_[86202]_  = A302 & ~A301;
  assign \new_[86203]_  = \new_[86202]_  & \new_[86199]_ ;
  assign \new_[86204]_  = \new_[86203]_  & \new_[86196]_ ;
  assign \new_[86208]_  = ~A199 & ~A168;
  assign \new_[86209]_  = A169 & \new_[86208]_ ;
  assign \new_[86212]_  = A201 & A200;
  assign \new_[86215]_  = ~A265 & A202;
  assign \new_[86216]_  = \new_[86215]_  & \new_[86212]_ ;
  assign \new_[86217]_  = \new_[86216]_  & \new_[86209]_ ;
  assign \new_[86220]_  = A267 & A266;
  assign \new_[86223]_  = A298 & ~A269;
  assign \new_[86224]_  = \new_[86223]_  & \new_[86220]_ ;
  assign \new_[86227]_  = ~A300 & ~A299;
  assign \new_[86230]_  = A302 & ~A301;
  assign \new_[86231]_  = \new_[86230]_  & \new_[86227]_ ;
  assign \new_[86232]_  = \new_[86231]_  & \new_[86224]_ ;
  assign \new_[86236]_  = ~A199 & ~A168;
  assign \new_[86237]_  = A169 & \new_[86236]_ ;
  assign \new_[86240]_  = A201 & A200;
  assign \new_[86243]_  = ~A265 & A202;
  assign \new_[86244]_  = \new_[86243]_  & \new_[86240]_ ;
  assign \new_[86245]_  = \new_[86244]_  & \new_[86237]_ ;
  assign \new_[86248]_  = A267 & A266;
  assign \new_[86251]_  = ~A298 & ~A269;
  assign \new_[86252]_  = \new_[86251]_  & \new_[86248]_ ;
  assign \new_[86255]_  = ~A300 & A299;
  assign \new_[86258]_  = A302 & ~A301;
  assign \new_[86259]_  = \new_[86258]_  & \new_[86255]_ ;
  assign \new_[86260]_  = \new_[86259]_  & \new_[86252]_ ;
  assign \new_[86264]_  = ~A199 & ~A168;
  assign \new_[86265]_  = A169 & \new_[86264]_ ;
  assign \new_[86268]_  = A201 & A200;
  assign \new_[86271]_  = ~A265 & A202;
  assign \new_[86272]_  = \new_[86271]_  & \new_[86268]_ ;
  assign \new_[86273]_  = \new_[86272]_  & \new_[86265]_ ;
  assign \new_[86276]_  = ~A267 & A266;
  assign \new_[86279]_  = A269 & ~A268;
  assign \new_[86280]_  = \new_[86279]_  & \new_[86276]_ ;
  assign \new_[86283]_  = ~A299 & A298;
  assign \new_[86286]_  = A301 & A300;
  assign \new_[86287]_  = \new_[86286]_  & \new_[86283]_ ;
  assign \new_[86288]_  = \new_[86287]_  & \new_[86280]_ ;
  assign \new_[86292]_  = ~A199 & ~A168;
  assign \new_[86293]_  = A169 & \new_[86292]_ ;
  assign \new_[86296]_  = A201 & A200;
  assign \new_[86299]_  = ~A265 & A202;
  assign \new_[86300]_  = \new_[86299]_  & \new_[86296]_ ;
  assign \new_[86301]_  = \new_[86300]_  & \new_[86293]_ ;
  assign \new_[86304]_  = ~A267 & A266;
  assign \new_[86307]_  = A269 & ~A268;
  assign \new_[86308]_  = \new_[86307]_  & \new_[86304]_ ;
  assign \new_[86311]_  = ~A299 & A298;
  assign \new_[86314]_  = ~A302 & A300;
  assign \new_[86315]_  = \new_[86314]_  & \new_[86311]_ ;
  assign \new_[86316]_  = \new_[86315]_  & \new_[86308]_ ;
  assign \new_[86320]_  = ~A199 & ~A168;
  assign \new_[86321]_  = A169 & \new_[86320]_ ;
  assign \new_[86324]_  = A201 & A200;
  assign \new_[86327]_  = ~A265 & A202;
  assign \new_[86328]_  = \new_[86327]_  & \new_[86324]_ ;
  assign \new_[86329]_  = \new_[86328]_  & \new_[86321]_ ;
  assign \new_[86332]_  = ~A267 & A266;
  assign \new_[86335]_  = A269 & ~A268;
  assign \new_[86336]_  = \new_[86335]_  & \new_[86332]_ ;
  assign \new_[86339]_  = A299 & ~A298;
  assign \new_[86342]_  = A301 & A300;
  assign \new_[86343]_  = \new_[86342]_  & \new_[86339]_ ;
  assign \new_[86344]_  = \new_[86343]_  & \new_[86336]_ ;
  assign \new_[86348]_  = ~A199 & ~A168;
  assign \new_[86349]_  = A169 & \new_[86348]_ ;
  assign \new_[86352]_  = A201 & A200;
  assign \new_[86355]_  = ~A265 & A202;
  assign \new_[86356]_  = \new_[86355]_  & \new_[86352]_ ;
  assign \new_[86357]_  = \new_[86356]_  & \new_[86349]_ ;
  assign \new_[86360]_  = ~A267 & A266;
  assign \new_[86363]_  = A269 & ~A268;
  assign \new_[86364]_  = \new_[86363]_  & \new_[86360]_ ;
  assign \new_[86367]_  = A299 & ~A298;
  assign \new_[86370]_  = ~A302 & A300;
  assign \new_[86371]_  = \new_[86370]_  & \new_[86367]_ ;
  assign \new_[86372]_  = \new_[86371]_  & \new_[86364]_ ;
  assign \new_[86376]_  = ~A199 & ~A168;
  assign \new_[86377]_  = A169 & \new_[86376]_ ;
  assign \new_[86380]_  = A201 & A200;
  assign \new_[86383]_  = A265 & A202;
  assign \new_[86384]_  = \new_[86383]_  & \new_[86380]_ ;
  assign \new_[86385]_  = \new_[86384]_  & \new_[86377]_ ;
  assign \new_[86388]_  = A267 & ~A266;
  assign \new_[86391]_  = A298 & A268;
  assign \new_[86392]_  = \new_[86391]_  & \new_[86388]_ ;
  assign \new_[86395]_  = ~A300 & ~A299;
  assign \new_[86398]_  = A302 & ~A301;
  assign \new_[86399]_  = \new_[86398]_  & \new_[86395]_ ;
  assign \new_[86400]_  = \new_[86399]_  & \new_[86392]_ ;
  assign \new_[86404]_  = ~A199 & ~A168;
  assign \new_[86405]_  = A169 & \new_[86404]_ ;
  assign \new_[86408]_  = A201 & A200;
  assign \new_[86411]_  = A265 & A202;
  assign \new_[86412]_  = \new_[86411]_  & \new_[86408]_ ;
  assign \new_[86413]_  = \new_[86412]_  & \new_[86405]_ ;
  assign \new_[86416]_  = A267 & ~A266;
  assign \new_[86419]_  = ~A298 & A268;
  assign \new_[86420]_  = \new_[86419]_  & \new_[86416]_ ;
  assign \new_[86423]_  = ~A300 & A299;
  assign \new_[86426]_  = A302 & ~A301;
  assign \new_[86427]_  = \new_[86426]_  & \new_[86423]_ ;
  assign \new_[86428]_  = \new_[86427]_  & \new_[86420]_ ;
  assign \new_[86432]_  = ~A199 & ~A168;
  assign \new_[86433]_  = A169 & \new_[86432]_ ;
  assign \new_[86436]_  = A201 & A200;
  assign \new_[86439]_  = A265 & A202;
  assign \new_[86440]_  = \new_[86439]_  & \new_[86436]_ ;
  assign \new_[86441]_  = \new_[86440]_  & \new_[86433]_ ;
  assign \new_[86444]_  = A267 & ~A266;
  assign \new_[86447]_  = A298 & ~A269;
  assign \new_[86448]_  = \new_[86447]_  & \new_[86444]_ ;
  assign \new_[86451]_  = ~A300 & ~A299;
  assign \new_[86454]_  = A302 & ~A301;
  assign \new_[86455]_  = \new_[86454]_  & \new_[86451]_ ;
  assign \new_[86456]_  = \new_[86455]_  & \new_[86448]_ ;
  assign \new_[86460]_  = ~A199 & ~A168;
  assign \new_[86461]_  = A169 & \new_[86460]_ ;
  assign \new_[86464]_  = A201 & A200;
  assign \new_[86467]_  = A265 & A202;
  assign \new_[86468]_  = \new_[86467]_  & \new_[86464]_ ;
  assign \new_[86469]_  = \new_[86468]_  & \new_[86461]_ ;
  assign \new_[86472]_  = A267 & ~A266;
  assign \new_[86475]_  = ~A298 & ~A269;
  assign \new_[86476]_  = \new_[86475]_  & \new_[86472]_ ;
  assign \new_[86479]_  = ~A300 & A299;
  assign \new_[86482]_  = A302 & ~A301;
  assign \new_[86483]_  = \new_[86482]_  & \new_[86479]_ ;
  assign \new_[86484]_  = \new_[86483]_  & \new_[86476]_ ;
  assign \new_[86488]_  = ~A199 & ~A168;
  assign \new_[86489]_  = A169 & \new_[86488]_ ;
  assign \new_[86492]_  = A201 & A200;
  assign \new_[86495]_  = A265 & A202;
  assign \new_[86496]_  = \new_[86495]_  & \new_[86492]_ ;
  assign \new_[86497]_  = \new_[86496]_  & \new_[86489]_ ;
  assign \new_[86500]_  = ~A267 & ~A266;
  assign \new_[86503]_  = A269 & ~A268;
  assign \new_[86504]_  = \new_[86503]_  & \new_[86500]_ ;
  assign \new_[86507]_  = ~A299 & A298;
  assign \new_[86510]_  = A301 & A300;
  assign \new_[86511]_  = \new_[86510]_  & \new_[86507]_ ;
  assign \new_[86512]_  = \new_[86511]_  & \new_[86504]_ ;
  assign \new_[86516]_  = ~A199 & ~A168;
  assign \new_[86517]_  = A169 & \new_[86516]_ ;
  assign \new_[86520]_  = A201 & A200;
  assign \new_[86523]_  = A265 & A202;
  assign \new_[86524]_  = \new_[86523]_  & \new_[86520]_ ;
  assign \new_[86525]_  = \new_[86524]_  & \new_[86517]_ ;
  assign \new_[86528]_  = ~A267 & ~A266;
  assign \new_[86531]_  = A269 & ~A268;
  assign \new_[86532]_  = \new_[86531]_  & \new_[86528]_ ;
  assign \new_[86535]_  = ~A299 & A298;
  assign \new_[86538]_  = ~A302 & A300;
  assign \new_[86539]_  = \new_[86538]_  & \new_[86535]_ ;
  assign \new_[86540]_  = \new_[86539]_  & \new_[86532]_ ;
  assign \new_[86544]_  = ~A199 & ~A168;
  assign \new_[86545]_  = A169 & \new_[86544]_ ;
  assign \new_[86548]_  = A201 & A200;
  assign \new_[86551]_  = A265 & A202;
  assign \new_[86552]_  = \new_[86551]_  & \new_[86548]_ ;
  assign \new_[86553]_  = \new_[86552]_  & \new_[86545]_ ;
  assign \new_[86556]_  = ~A267 & ~A266;
  assign \new_[86559]_  = A269 & ~A268;
  assign \new_[86560]_  = \new_[86559]_  & \new_[86556]_ ;
  assign \new_[86563]_  = A299 & ~A298;
  assign \new_[86566]_  = A301 & A300;
  assign \new_[86567]_  = \new_[86566]_  & \new_[86563]_ ;
  assign \new_[86568]_  = \new_[86567]_  & \new_[86560]_ ;
  assign \new_[86572]_  = ~A199 & ~A168;
  assign \new_[86573]_  = A169 & \new_[86572]_ ;
  assign \new_[86576]_  = A201 & A200;
  assign \new_[86579]_  = A265 & A202;
  assign \new_[86580]_  = \new_[86579]_  & \new_[86576]_ ;
  assign \new_[86581]_  = \new_[86580]_  & \new_[86573]_ ;
  assign \new_[86584]_  = ~A267 & ~A266;
  assign \new_[86587]_  = A269 & ~A268;
  assign \new_[86588]_  = \new_[86587]_  & \new_[86584]_ ;
  assign \new_[86591]_  = A299 & ~A298;
  assign \new_[86594]_  = ~A302 & A300;
  assign \new_[86595]_  = \new_[86594]_  & \new_[86591]_ ;
  assign \new_[86596]_  = \new_[86595]_  & \new_[86588]_ ;
  assign \new_[86600]_  = ~A199 & ~A168;
  assign \new_[86601]_  = A169 & \new_[86600]_ ;
  assign \new_[86604]_  = A201 & A200;
  assign \new_[86607]_  = ~A265 & ~A203;
  assign \new_[86608]_  = \new_[86607]_  & \new_[86604]_ ;
  assign \new_[86609]_  = \new_[86608]_  & \new_[86601]_ ;
  assign \new_[86612]_  = A267 & A266;
  assign \new_[86615]_  = A298 & A268;
  assign \new_[86616]_  = \new_[86615]_  & \new_[86612]_ ;
  assign \new_[86619]_  = ~A300 & ~A299;
  assign \new_[86622]_  = A302 & ~A301;
  assign \new_[86623]_  = \new_[86622]_  & \new_[86619]_ ;
  assign \new_[86624]_  = \new_[86623]_  & \new_[86616]_ ;
  assign \new_[86628]_  = ~A199 & ~A168;
  assign \new_[86629]_  = A169 & \new_[86628]_ ;
  assign \new_[86632]_  = A201 & A200;
  assign \new_[86635]_  = ~A265 & ~A203;
  assign \new_[86636]_  = \new_[86635]_  & \new_[86632]_ ;
  assign \new_[86637]_  = \new_[86636]_  & \new_[86629]_ ;
  assign \new_[86640]_  = A267 & A266;
  assign \new_[86643]_  = ~A298 & A268;
  assign \new_[86644]_  = \new_[86643]_  & \new_[86640]_ ;
  assign \new_[86647]_  = ~A300 & A299;
  assign \new_[86650]_  = A302 & ~A301;
  assign \new_[86651]_  = \new_[86650]_  & \new_[86647]_ ;
  assign \new_[86652]_  = \new_[86651]_  & \new_[86644]_ ;
  assign \new_[86656]_  = ~A199 & ~A168;
  assign \new_[86657]_  = A169 & \new_[86656]_ ;
  assign \new_[86660]_  = A201 & A200;
  assign \new_[86663]_  = ~A265 & ~A203;
  assign \new_[86664]_  = \new_[86663]_  & \new_[86660]_ ;
  assign \new_[86665]_  = \new_[86664]_  & \new_[86657]_ ;
  assign \new_[86668]_  = A267 & A266;
  assign \new_[86671]_  = A298 & ~A269;
  assign \new_[86672]_  = \new_[86671]_  & \new_[86668]_ ;
  assign \new_[86675]_  = ~A300 & ~A299;
  assign \new_[86678]_  = A302 & ~A301;
  assign \new_[86679]_  = \new_[86678]_  & \new_[86675]_ ;
  assign \new_[86680]_  = \new_[86679]_  & \new_[86672]_ ;
  assign \new_[86684]_  = ~A199 & ~A168;
  assign \new_[86685]_  = A169 & \new_[86684]_ ;
  assign \new_[86688]_  = A201 & A200;
  assign \new_[86691]_  = ~A265 & ~A203;
  assign \new_[86692]_  = \new_[86691]_  & \new_[86688]_ ;
  assign \new_[86693]_  = \new_[86692]_  & \new_[86685]_ ;
  assign \new_[86696]_  = A267 & A266;
  assign \new_[86699]_  = ~A298 & ~A269;
  assign \new_[86700]_  = \new_[86699]_  & \new_[86696]_ ;
  assign \new_[86703]_  = ~A300 & A299;
  assign \new_[86706]_  = A302 & ~A301;
  assign \new_[86707]_  = \new_[86706]_  & \new_[86703]_ ;
  assign \new_[86708]_  = \new_[86707]_  & \new_[86700]_ ;
  assign \new_[86712]_  = ~A199 & ~A168;
  assign \new_[86713]_  = A169 & \new_[86712]_ ;
  assign \new_[86716]_  = A201 & A200;
  assign \new_[86719]_  = ~A265 & ~A203;
  assign \new_[86720]_  = \new_[86719]_  & \new_[86716]_ ;
  assign \new_[86721]_  = \new_[86720]_  & \new_[86713]_ ;
  assign \new_[86724]_  = ~A267 & A266;
  assign \new_[86727]_  = A269 & ~A268;
  assign \new_[86728]_  = \new_[86727]_  & \new_[86724]_ ;
  assign \new_[86731]_  = ~A299 & A298;
  assign \new_[86734]_  = A301 & A300;
  assign \new_[86735]_  = \new_[86734]_  & \new_[86731]_ ;
  assign \new_[86736]_  = \new_[86735]_  & \new_[86728]_ ;
  assign \new_[86740]_  = ~A199 & ~A168;
  assign \new_[86741]_  = A169 & \new_[86740]_ ;
  assign \new_[86744]_  = A201 & A200;
  assign \new_[86747]_  = ~A265 & ~A203;
  assign \new_[86748]_  = \new_[86747]_  & \new_[86744]_ ;
  assign \new_[86749]_  = \new_[86748]_  & \new_[86741]_ ;
  assign \new_[86752]_  = ~A267 & A266;
  assign \new_[86755]_  = A269 & ~A268;
  assign \new_[86756]_  = \new_[86755]_  & \new_[86752]_ ;
  assign \new_[86759]_  = ~A299 & A298;
  assign \new_[86762]_  = ~A302 & A300;
  assign \new_[86763]_  = \new_[86762]_  & \new_[86759]_ ;
  assign \new_[86764]_  = \new_[86763]_  & \new_[86756]_ ;
  assign \new_[86768]_  = ~A199 & ~A168;
  assign \new_[86769]_  = A169 & \new_[86768]_ ;
  assign \new_[86772]_  = A201 & A200;
  assign \new_[86775]_  = ~A265 & ~A203;
  assign \new_[86776]_  = \new_[86775]_  & \new_[86772]_ ;
  assign \new_[86777]_  = \new_[86776]_  & \new_[86769]_ ;
  assign \new_[86780]_  = ~A267 & A266;
  assign \new_[86783]_  = A269 & ~A268;
  assign \new_[86784]_  = \new_[86783]_  & \new_[86780]_ ;
  assign \new_[86787]_  = A299 & ~A298;
  assign \new_[86790]_  = A301 & A300;
  assign \new_[86791]_  = \new_[86790]_  & \new_[86787]_ ;
  assign \new_[86792]_  = \new_[86791]_  & \new_[86784]_ ;
  assign \new_[86796]_  = ~A199 & ~A168;
  assign \new_[86797]_  = A169 & \new_[86796]_ ;
  assign \new_[86800]_  = A201 & A200;
  assign \new_[86803]_  = ~A265 & ~A203;
  assign \new_[86804]_  = \new_[86803]_  & \new_[86800]_ ;
  assign \new_[86805]_  = \new_[86804]_  & \new_[86797]_ ;
  assign \new_[86808]_  = ~A267 & A266;
  assign \new_[86811]_  = A269 & ~A268;
  assign \new_[86812]_  = \new_[86811]_  & \new_[86808]_ ;
  assign \new_[86815]_  = A299 & ~A298;
  assign \new_[86818]_  = ~A302 & A300;
  assign \new_[86819]_  = \new_[86818]_  & \new_[86815]_ ;
  assign \new_[86820]_  = \new_[86819]_  & \new_[86812]_ ;
  assign \new_[86824]_  = ~A199 & ~A168;
  assign \new_[86825]_  = A169 & \new_[86824]_ ;
  assign \new_[86828]_  = A201 & A200;
  assign \new_[86831]_  = A265 & ~A203;
  assign \new_[86832]_  = \new_[86831]_  & \new_[86828]_ ;
  assign \new_[86833]_  = \new_[86832]_  & \new_[86825]_ ;
  assign \new_[86836]_  = A267 & ~A266;
  assign \new_[86839]_  = A298 & A268;
  assign \new_[86840]_  = \new_[86839]_  & \new_[86836]_ ;
  assign \new_[86843]_  = ~A300 & ~A299;
  assign \new_[86846]_  = A302 & ~A301;
  assign \new_[86847]_  = \new_[86846]_  & \new_[86843]_ ;
  assign \new_[86848]_  = \new_[86847]_  & \new_[86840]_ ;
  assign \new_[86852]_  = ~A199 & ~A168;
  assign \new_[86853]_  = A169 & \new_[86852]_ ;
  assign \new_[86856]_  = A201 & A200;
  assign \new_[86859]_  = A265 & ~A203;
  assign \new_[86860]_  = \new_[86859]_  & \new_[86856]_ ;
  assign \new_[86861]_  = \new_[86860]_  & \new_[86853]_ ;
  assign \new_[86864]_  = A267 & ~A266;
  assign \new_[86867]_  = ~A298 & A268;
  assign \new_[86868]_  = \new_[86867]_  & \new_[86864]_ ;
  assign \new_[86871]_  = ~A300 & A299;
  assign \new_[86874]_  = A302 & ~A301;
  assign \new_[86875]_  = \new_[86874]_  & \new_[86871]_ ;
  assign \new_[86876]_  = \new_[86875]_  & \new_[86868]_ ;
  assign \new_[86880]_  = ~A199 & ~A168;
  assign \new_[86881]_  = A169 & \new_[86880]_ ;
  assign \new_[86884]_  = A201 & A200;
  assign \new_[86887]_  = A265 & ~A203;
  assign \new_[86888]_  = \new_[86887]_  & \new_[86884]_ ;
  assign \new_[86889]_  = \new_[86888]_  & \new_[86881]_ ;
  assign \new_[86892]_  = A267 & ~A266;
  assign \new_[86895]_  = A298 & ~A269;
  assign \new_[86896]_  = \new_[86895]_  & \new_[86892]_ ;
  assign \new_[86899]_  = ~A300 & ~A299;
  assign \new_[86902]_  = A302 & ~A301;
  assign \new_[86903]_  = \new_[86902]_  & \new_[86899]_ ;
  assign \new_[86904]_  = \new_[86903]_  & \new_[86896]_ ;
  assign \new_[86908]_  = ~A199 & ~A168;
  assign \new_[86909]_  = A169 & \new_[86908]_ ;
  assign \new_[86912]_  = A201 & A200;
  assign \new_[86915]_  = A265 & ~A203;
  assign \new_[86916]_  = \new_[86915]_  & \new_[86912]_ ;
  assign \new_[86917]_  = \new_[86916]_  & \new_[86909]_ ;
  assign \new_[86920]_  = A267 & ~A266;
  assign \new_[86923]_  = ~A298 & ~A269;
  assign \new_[86924]_  = \new_[86923]_  & \new_[86920]_ ;
  assign \new_[86927]_  = ~A300 & A299;
  assign \new_[86930]_  = A302 & ~A301;
  assign \new_[86931]_  = \new_[86930]_  & \new_[86927]_ ;
  assign \new_[86932]_  = \new_[86931]_  & \new_[86924]_ ;
  assign \new_[86936]_  = ~A199 & ~A168;
  assign \new_[86937]_  = A169 & \new_[86936]_ ;
  assign \new_[86940]_  = A201 & A200;
  assign \new_[86943]_  = A265 & ~A203;
  assign \new_[86944]_  = \new_[86943]_  & \new_[86940]_ ;
  assign \new_[86945]_  = \new_[86944]_  & \new_[86937]_ ;
  assign \new_[86948]_  = ~A267 & ~A266;
  assign \new_[86951]_  = A269 & ~A268;
  assign \new_[86952]_  = \new_[86951]_  & \new_[86948]_ ;
  assign \new_[86955]_  = ~A299 & A298;
  assign \new_[86958]_  = A301 & A300;
  assign \new_[86959]_  = \new_[86958]_  & \new_[86955]_ ;
  assign \new_[86960]_  = \new_[86959]_  & \new_[86952]_ ;
  assign \new_[86964]_  = ~A199 & ~A168;
  assign \new_[86965]_  = A169 & \new_[86964]_ ;
  assign \new_[86968]_  = A201 & A200;
  assign \new_[86971]_  = A265 & ~A203;
  assign \new_[86972]_  = \new_[86971]_  & \new_[86968]_ ;
  assign \new_[86973]_  = \new_[86972]_  & \new_[86965]_ ;
  assign \new_[86976]_  = ~A267 & ~A266;
  assign \new_[86979]_  = A269 & ~A268;
  assign \new_[86980]_  = \new_[86979]_  & \new_[86976]_ ;
  assign \new_[86983]_  = ~A299 & A298;
  assign \new_[86986]_  = ~A302 & A300;
  assign \new_[86987]_  = \new_[86986]_  & \new_[86983]_ ;
  assign \new_[86988]_  = \new_[86987]_  & \new_[86980]_ ;
  assign \new_[86992]_  = ~A199 & ~A168;
  assign \new_[86993]_  = A169 & \new_[86992]_ ;
  assign \new_[86996]_  = A201 & A200;
  assign \new_[86999]_  = A265 & ~A203;
  assign \new_[87000]_  = \new_[86999]_  & \new_[86996]_ ;
  assign \new_[87001]_  = \new_[87000]_  & \new_[86993]_ ;
  assign \new_[87004]_  = ~A267 & ~A266;
  assign \new_[87007]_  = A269 & ~A268;
  assign \new_[87008]_  = \new_[87007]_  & \new_[87004]_ ;
  assign \new_[87011]_  = A299 & ~A298;
  assign \new_[87014]_  = A301 & A300;
  assign \new_[87015]_  = \new_[87014]_  & \new_[87011]_ ;
  assign \new_[87016]_  = \new_[87015]_  & \new_[87008]_ ;
  assign \new_[87020]_  = ~A199 & ~A168;
  assign \new_[87021]_  = A169 & \new_[87020]_ ;
  assign \new_[87024]_  = A201 & A200;
  assign \new_[87027]_  = A265 & ~A203;
  assign \new_[87028]_  = \new_[87027]_  & \new_[87024]_ ;
  assign \new_[87029]_  = \new_[87028]_  & \new_[87021]_ ;
  assign \new_[87032]_  = ~A267 & ~A266;
  assign \new_[87035]_  = A269 & ~A268;
  assign \new_[87036]_  = \new_[87035]_  & \new_[87032]_ ;
  assign \new_[87039]_  = A299 & ~A298;
  assign \new_[87042]_  = ~A302 & A300;
  assign \new_[87043]_  = \new_[87042]_  & \new_[87039]_ ;
  assign \new_[87044]_  = \new_[87043]_  & \new_[87036]_ ;
  assign \new_[87048]_  = ~A199 & ~A168;
  assign \new_[87049]_  = A169 & \new_[87048]_ ;
  assign \new_[87052]_  = ~A201 & A200;
  assign \new_[87055]_  = A203 & ~A202;
  assign \new_[87056]_  = \new_[87055]_  & \new_[87052]_ ;
  assign \new_[87057]_  = \new_[87056]_  & \new_[87049]_ ;
  assign \new_[87060]_  = A266 & ~A265;
  assign \new_[87063]_  = A268 & A267;
  assign \new_[87064]_  = \new_[87063]_  & \new_[87060]_ ;
  assign \new_[87067]_  = ~A299 & A298;
  assign \new_[87070]_  = A301 & A300;
  assign \new_[87071]_  = \new_[87070]_  & \new_[87067]_ ;
  assign \new_[87072]_  = \new_[87071]_  & \new_[87064]_ ;
  assign \new_[87076]_  = ~A199 & ~A168;
  assign \new_[87077]_  = A169 & \new_[87076]_ ;
  assign \new_[87080]_  = ~A201 & A200;
  assign \new_[87083]_  = A203 & ~A202;
  assign \new_[87084]_  = \new_[87083]_  & \new_[87080]_ ;
  assign \new_[87085]_  = \new_[87084]_  & \new_[87077]_ ;
  assign \new_[87088]_  = A266 & ~A265;
  assign \new_[87091]_  = A268 & A267;
  assign \new_[87092]_  = \new_[87091]_  & \new_[87088]_ ;
  assign \new_[87095]_  = ~A299 & A298;
  assign \new_[87098]_  = ~A302 & A300;
  assign \new_[87099]_  = \new_[87098]_  & \new_[87095]_ ;
  assign \new_[87100]_  = \new_[87099]_  & \new_[87092]_ ;
  assign \new_[87104]_  = ~A199 & ~A168;
  assign \new_[87105]_  = A169 & \new_[87104]_ ;
  assign \new_[87108]_  = ~A201 & A200;
  assign \new_[87111]_  = A203 & ~A202;
  assign \new_[87112]_  = \new_[87111]_  & \new_[87108]_ ;
  assign \new_[87113]_  = \new_[87112]_  & \new_[87105]_ ;
  assign \new_[87116]_  = A266 & ~A265;
  assign \new_[87119]_  = A268 & A267;
  assign \new_[87120]_  = \new_[87119]_  & \new_[87116]_ ;
  assign \new_[87123]_  = A299 & ~A298;
  assign \new_[87126]_  = A301 & A300;
  assign \new_[87127]_  = \new_[87126]_  & \new_[87123]_ ;
  assign \new_[87128]_  = \new_[87127]_  & \new_[87120]_ ;
  assign \new_[87132]_  = ~A199 & ~A168;
  assign \new_[87133]_  = A169 & \new_[87132]_ ;
  assign \new_[87136]_  = ~A201 & A200;
  assign \new_[87139]_  = A203 & ~A202;
  assign \new_[87140]_  = \new_[87139]_  & \new_[87136]_ ;
  assign \new_[87141]_  = \new_[87140]_  & \new_[87133]_ ;
  assign \new_[87144]_  = A266 & ~A265;
  assign \new_[87147]_  = A268 & A267;
  assign \new_[87148]_  = \new_[87147]_  & \new_[87144]_ ;
  assign \new_[87151]_  = A299 & ~A298;
  assign \new_[87154]_  = ~A302 & A300;
  assign \new_[87155]_  = \new_[87154]_  & \new_[87151]_ ;
  assign \new_[87156]_  = \new_[87155]_  & \new_[87148]_ ;
  assign \new_[87160]_  = ~A199 & ~A168;
  assign \new_[87161]_  = A169 & \new_[87160]_ ;
  assign \new_[87164]_  = ~A201 & A200;
  assign \new_[87167]_  = A203 & ~A202;
  assign \new_[87168]_  = \new_[87167]_  & \new_[87164]_ ;
  assign \new_[87169]_  = \new_[87168]_  & \new_[87161]_ ;
  assign \new_[87172]_  = A266 & ~A265;
  assign \new_[87175]_  = ~A269 & A267;
  assign \new_[87176]_  = \new_[87175]_  & \new_[87172]_ ;
  assign \new_[87179]_  = ~A299 & A298;
  assign \new_[87182]_  = A301 & A300;
  assign \new_[87183]_  = \new_[87182]_  & \new_[87179]_ ;
  assign \new_[87184]_  = \new_[87183]_  & \new_[87176]_ ;
  assign \new_[87188]_  = ~A199 & ~A168;
  assign \new_[87189]_  = A169 & \new_[87188]_ ;
  assign \new_[87192]_  = ~A201 & A200;
  assign \new_[87195]_  = A203 & ~A202;
  assign \new_[87196]_  = \new_[87195]_  & \new_[87192]_ ;
  assign \new_[87197]_  = \new_[87196]_  & \new_[87189]_ ;
  assign \new_[87200]_  = A266 & ~A265;
  assign \new_[87203]_  = ~A269 & A267;
  assign \new_[87204]_  = \new_[87203]_  & \new_[87200]_ ;
  assign \new_[87207]_  = ~A299 & A298;
  assign \new_[87210]_  = ~A302 & A300;
  assign \new_[87211]_  = \new_[87210]_  & \new_[87207]_ ;
  assign \new_[87212]_  = \new_[87211]_  & \new_[87204]_ ;
  assign \new_[87216]_  = ~A199 & ~A168;
  assign \new_[87217]_  = A169 & \new_[87216]_ ;
  assign \new_[87220]_  = ~A201 & A200;
  assign \new_[87223]_  = A203 & ~A202;
  assign \new_[87224]_  = \new_[87223]_  & \new_[87220]_ ;
  assign \new_[87225]_  = \new_[87224]_  & \new_[87217]_ ;
  assign \new_[87228]_  = A266 & ~A265;
  assign \new_[87231]_  = ~A269 & A267;
  assign \new_[87232]_  = \new_[87231]_  & \new_[87228]_ ;
  assign \new_[87235]_  = A299 & ~A298;
  assign \new_[87238]_  = A301 & A300;
  assign \new_[87239]_  = \new_[87238]_  & \new_[87235]_ ;
  assign \new_[87240]_  = \new_[87239]_  & \new_[87232]_ ;
  assign \new_[87244]_  = ~A199 & ~A168;
  assign \new_[87245]_  = A169 & \new_[87244]_ ;
  assign \new_[87248]_  = ~A201 & A200;
  assign \new_[87251]_  = A203 & ~A202;
  assign \new_[87252]_  = \new_[87251]_  & \new_[87248]_ ;
  assign \new_[87253]_  = \new_[87252]_  & \new_[87245]_ ;
  assign \new_[87256]_  = A266 & ~A265;
  assign \new_[87259]_  = ~A269 & A267;
  assign \new_[87260]_  = \new_[87259]_  & \new_[87256]_ ;
  assign \new_[87263]_  = A299 & ~A298;
  assign \new_[87266]_  = ~A302 & A300;
  assign \new_[87267]_  = \new_[87266]_  & \new_[87263]_ ;
  assign \new_[87268]_  = \new_[87267]_  & \new_[87260]_ ;
  assign \new_[87272]_  = ~A199 & ~A168;
  assign \new_[87273]_  = A169 & \new_[87272]_ ;
  assign \new_[87276]_  = ~A201 & A200;
  assign \new_[87279]_  = A203 & ~A202;
  assign \new_[87280]_  = \new_[87279]_  & \new_[87276]_ ;
  assign \new_[87281]_  = \new_[87280]_  & \new_[87273]_ ;
  assign \new_[87284]_  = ~A266 & A265;
  assign \new_[87287]_  = A268 & A267;
  assign \new_[87288]_  = \new_[87287]_  & \new_[87284]_ ;
  assign \new_[87291]_  = ~A299 & A298;
  assign \new_[87294]_  = A301 & A300;
  assign \new_[87295]_  = \new_[87294]_  & \new_[87291]_ ;
  assign \new_[87296]_  = \new_[87295]_  & \new_[87288]_ ;
  assign \new_[87300]_  = ~A199 & ~A168;
  assign \new_[87301]_  = A169 & \new_[87300]_ ;
  assign \new_[87304]_  = ~A201 & A200;
  assign \new_[87307]_  = A203 & ~A202;
  assign \new_[87308]_  = \new_[87307]_  & \new_[87304]_ ;
  assign \new_[87309]_  = \new_[87308]_  & \new_[87301]_ ;
  assign \new_[87312]_  = ~A266 & A265;
  assign \new_[87315]_  = A268 & A267;
  assign \new_[87316]_  = \new_[87315]_  & \new_[87312]_ ;
  assign \new_[87319]_  = ~A299 & A298;
  assign \new_[87322]_  = ~A302 & A300;
  assign \new_[87323]_  = \new_[87322]_  & \new_[87319]_ ;
  assign \new_[87324]_  = \new_[87323]_  & \new_[87316]_ ;
  assign \new_[87328]_  = ~A199 & ~A168;
  assign \new_[87329]_  = A169 & \new_[87328]_ ;
  assign \new_[87332]_  = ~A201 & A200;
  assign \new_[87335]_  = A203 & ~A202;
  assign \new_[87336]_  = \new_[87335]_  & \new_[87332]_ ;
  assign \new_[87337]_  = \new_[87336]_  & \new_[87329]_ ;
  assign \new_[87340]_  = ~A266 & A265;
  assign \new_[87343]_  = A268 & A267;
  assign \new_[87344]_  = \new_[87343]_  & \new_[87340]_ ;
  assign \new_[87347]_  = A299 & ~A298;
  assign \new_[87350]_  = A301 & A300;
  assign \new_[87351]_  = \new_[87350]_  & \new_[87347]_ ;
  assign \new_[87352]_  = \new_[87351]_  & \new_[87344]_ ;
  assign \new_[87356]_  = ~A199 & ~A168;
  assign \new_[87357]_  = A169 & \new_[87356]_ ;
  assign \new_[87360]_  = ~A201 & A200;
  assign \new_[87363]_  = A203 & ~A202;
  assign \new_[87364]_  = \new_[87363]_  & \new_[87360]_ ;
  assign \new_[87365]_  = \new_[87364]_  & \new_[87357]_ ;
  assign \new_[87368]_  = ~A266 & A265;
  assign \new_[87371]_  = A268 & A267;
  assign \new_[87372]_  = \new_[87371]_  & \new_[87368]_ ;
  assign \new_[87375]_  = A299 & ~A298;
  assign \new_[87378]_  = ~A302 & A300;
  assign \new_[87379]_  = \new_[87378]_  & \new_[87375]_ ;
  assign \new_[87380]_  = \new_[87379]_  & \new_[87372]_ ;
  assign \new_[87384]_  = ~A199 & ~A168;
  assign \new_[87385]_  = A169 & \new_[87384]_ ;
  assign \new_[87388]_  = ~A201 & A200;
  assign \new_[87391]_  = A203 & ~A202;
  assign \new_[87392]_  = \new_[87391]_  & \new_[87388]_ ;
  assign \new_[87393]_  = \new_[87392]_  & \new_[87385]_ ;
  assign \new_[87396]_  = ~A266 & A265;
  assign \new_[87399]_  = ~A269 & A267;
  assign \new_[87400]_  = \new_[87399]_  & \new_[87396]_ ;
  assign \new_[87403]_  = ~A299 & A298;
  assign \new_[87406]_  = A301 & A300;
  assign \new_[87407]_  = \new_[87406]_  & \new_[87403]_ ;
  assign \new_[87408]_  = \new_[87407]_  & \new_[87400]_ ;
  assign \new_[87412]_  = ~A199 & ~A168;
  assign \new_[87413]_  = A169 & \new_[87412]_ ;
  assign \new_[87416]_  = ~A201 & A200;
  assign \new_[87419]_  = A203 & ~A202;
  assign \new_[87420]_  = \new_[87419]_  & \new_[87416]_ ;
  assign \new_[87421]_  = \new_[87420]_  & \new_[87413]_ ;
  assign \new_[87424]_  = ~A266 & A265;
  assign \new_[87427]_  = ~A269 & A267;
  assign \new_[87428]_  = \new_[87427]_  & \new_[87424]_ ;
  assign \new_[87431]_  = ~A299 & A298;
  assign \new_[87434]_  = ~A302 & A300;
  assign \new_[87435]_  = \new_[87434]_  & \new_[87431]_ ;
  assign \new_[87436]_  = \new_[87435]_  & \new_[87428]_ ;
  assign \new_[87440]_  = ~A199 & ~A168;
  assign \new_[87441]_  = A169 & \new_[87440]_ ;
  assign \new_[87444]_  = ~A201 & A200;
  assign \new_[87447]_  = A203 & ~A202;
  assign \new_[87448]_  = \new_[87447]_  & \new_[87444]_ ;
  assign \new_[87449]_  = \new_[87448]_  & \new_[87441]_ ;
  assign \new_[87452]_  = ~A266 & A265;
  assign \new_[87455]_  = ~A269 & A267;
  assign \new_[87456]_  = \new_[87455]_  & \new_[87452]_ ;
  assign \new_[87459]_  = A299 & ~A298;
  assign \new_[87462]_  = A301 & A300;
  assign \new_[87463]_  = \new_[87462]_  & \new_[87459]_ ;
  assign \new_[87464]_  = \new_[87463]_  & \new_[87456]_ ;
  assign \new_[87468]_  = ~A199 & ~A168;
  assign \new_[87469]_  = A169 & \new_[87468]_ ;
  assign \new_[87472]_  = ~A201 & A200;
  assign \new_[87475]_  = A203 & ~A202;
  assign \new_[87476]_  = \new_[87475]_  & \new_[87472]_ ;
  assign \new_[87477]_  = \new_[87476]_  & \new_[87469]_ ;
  assign \new_[87480]_  = ~A266 & A265;
  assign \new_[87483]_  = ~A269 & A267;
  assign \new_[87484]_  = \new_[87483]_  & \new_[87480]_ ;
  assign \new_[87487]_  = A299 & ~A298;
  assign \new_[87490]_  = ~A302 & A300;
  assign \new_[87491]_  = \new_[87490]_  & \new_[87487]_ ;
  assign \new_[87492]_  = \new_[87491]_  & \new_[87484]_ ;
  assign \new_[87496]_  = A199 & ~A168;
  assign \new_[87497]_  = A169 & \new_[87496]_ ;
  assign \new_[87500]_  = A201 & ~A200;
  assign \new_[87503]_  = ~A265 & A202;
  assign \new_[87504]_  = \new_[87503]_  & \new_[87500]_ ;
  assign \new_[87505]_  = \new_[87504]_  & \new_[87497]_ ;
  assign \new_[87508]_  = A267 & A266;
  assign \new_[87511]_  = A298 & A268;
  assign \new_[87512]_  = \new_[87511]_  & \new_[87508]_ ;
  assign \new_[87515]_  = ~A300 & ~A299;
  assign \new_[87518]_  = A302 & ~A301;
  assign \new_[87519]_  = \new_[87518]_  & \new_[87515]_ ;
  assign \new_[87520]_  = \new_[87519]_  & \new_[87512]_ ;
  assign \new_[87524]_  = A199 & ~A168;
  assign \new_[87525]_  = A169 & \new_[87524]_ ;
  assign \new_[87528]_  = A201 & ~A200;
  assign \new_[87531]_  = ~A265 & A202;
  assign \new_[87532]_  = \new_[87531]_  & \new_[87528]_ ;
  assign \new_[87533]_  = \new_[87532]_  & \new_[87525]_ ;
  assign \new_[87536]_  = A267 & A266;
  assign \new_[87539]_  = ~A298 & A268;
  assign \new_[87540]_  = \new_[87539]_  & \new_[87536]_ ;
  assign \new_[87543]_  = ~A300 & A299;
  assign \new_[87546]_  = A302 & ~A301;
  assign \new_[87547]_  = \new_[87546]_  & \new_[87543]_ ;
  assign \new_[87548]_  = \new_[87547]_  & \new_[87540]_ ;
  assign \new_[87552]_  = A199 & ~A168;
  assign \new_[87553]_  = A169 & \new_[87552]_ ;
  assign \new_[87556]_  = A201 & ~A200;
  assign \new_[87559]_  = ~A265 & A202;
  assign \new_[87560]_  = \new_[87559]_  & \new_[87556]_ ;
  assign \new_[87561]_  = \new_[87560]_  & \new_[87553]_ ;
  assign \new_[87564]_  = A267 & A266;
  assign \new_[87567]_  = A298 & ~A269;
  assign \new_[87568]_  = \new_[87567]_  & \new_[87564]_ ;
  assign \new_[87571]_  = ~A300 & ~A299;
  assign \new_[87574]_  = A302 & ~A301;
  assign \new_[87575]_  = \new_[87574]_  & \new_[87571]_ ;
  assign \new_[87576]_  = \new_[87575]_  & \new_[87568]_ ;
  assign \new_[87580]_  = A199 & ~A168;
  assign \new_[87581]_  = A169 & \new_[87580]_ ;
  assign \new_[87584]_  = A201 & ~A200;
  assign \new_[87587]_  = ~A265 & A202;
  assign \new_[87588]_  = \new_[87587]_  & \new_[87584]_ ;
  assign \new_[87589]_  = \new_[87588]_  & \new_[87581]_ ;
  assign \new_[87592]_  = A267 & A266;
  assign \new_[87595]_  = ~A298 & ~A269;
  assign \new_[87596]_  = \new_[87595]_  & \new_[87592]_ ;
  assign \new_[87599]_  = ~A300 & A299;
  assign \new_[87602]_  = A302 & ~A301;
  assign \new_[87603]_  = \new_[87602]_  & \new_[87599]_ ;
  assign \new_[87604]_  = \new_[87603]_  & \new_[87596]_ ;
  assign \new_[87608]_  = A199 & ~A168;
  assign \new_[87609]_  = A169 & \new_[87608]_ ;
  assign \new_[87612]_  = A201 & ~A200;
  assign \new_[87615]_  = ~A265 & A202;
  assign \new_[87616]_  = \new_[87615]_  & \new_[87612]_ ;
  assign \new_[87617]_  = \new_[87616]_  & \new_[87609]_ ;
  assign \new_[87620]_  = ~A267 & A266;
  assign \new_[87623]_  = A269 & ~A268;
  assign \new_[87624]_  = \new_[87623]_  & \new_[87620]_ ;
  assign \new_[87627]_  = ~A299 & A298;
  assign \new_[87630]_  = A301 & A300;
  assign \new_[87631]_  = \new_[87630]_  & \new_[87627]_ ;
  assign \new_[87632]_  = \new_[87631]_  & \new_[87624]_ ;
  assign \new_[87636]_  = A199 & ~A168;
  assign \new_[87637]_  = A169 & \new_[87636]_ ;
  assign \new_[87640]_  = A201 & ~A200;
  assign \new_[87643]_  = ~A265 & A202;
  assign \new_[87644]_  = \new_[87643]_  & \new_[87640]_ ;
  assign \new_[87645]_  = \new_[87644]_  & \new_[87637]_ ;
  assign \new_[87648]_  = ~A267 & A266;
  assign \new_[87651]_  = A269 & ~A268;
  assign \new_[87652]_  = \new_[87651]_  & \new_[87648]_ ;
  assign \new_[87655]_  = ~A299 & A298;
  assign \new_[87658]_  = ~A302 & A300;
  assign \new_[87659]_  = \new_[87658]_  & \new_[87655]_ ;
  assign \new_[87660]_  = \new_[87659]_  & \new_[87652]_ ;
  assign \new_[87664]_  = A199 & ~A168;
  assign \new_[87665]_  = A169 & \new_[87664]_ ;
  assign \new_[87668]_  = A201 & ~A200;
  assign \new_[87671]_  = ~A265 & A202;
  assign \new_[87672]_  = \new_[87671]_  & \new_[87668]_ ;
  assign \new_[87673]_  = \new_[87672]_  & \new_[87665]_ ;
  assign \new_[87676]_  = ~A267 & A266;
  assign \new_[87679]_  = A269 & ~A268;
  assign \new_[87680]_  = \new_[87679]_  & \new_[87676]_ ;
  assign \new_[87683]_  = A299 & ~A298;
  assign \new_[87686]_  = A301 & A300;
  assign \new_[87687]_  = \new_[87686]_  & \new_[87683]_ ;
  assign \new_[87688]_  = \new_[87687]_  & \new_[87680]_ ;
  assign \new_[87692]_  = A199 & ~A168;
  assign \new_[87693]_  = A169 & \new_[87692]_ ;
  assign \new_[87696]_  = A201 & ~A200;
  assign \new_[87699]_  = ~A265 & A202;
  assign \new_[87700]_  = \new_[87699]_  & \new_[87696]_ ;
  assign \new_[87701]_  = \new_[87700]_  & \new_[87693]_ ;
  assign \new_[87704]_  = ~A267 & A266;
  assign \new_[87707]_  = A269 & ~A268;
  assign \new_[87708]_  = \new_[87707]_  & \new_[87704]_ ;
  assign \new_[87711]_  = A299 & ~A298;
  assign \new_[87714]_  = ~A302 & A300;
  assign \new_[87715]_  = \new_[87714]_  & \new_[87711]_ ;
  assign \new_[87716]_  = \new_[87715]_  & \new_[87708]_ ;
  assign \new_[87720]_  = A199 & ~A168;
  assign \new_[87721]_  = A169 & \new_[87720]_ ;
  assign \new_[87724]_  = A201 & ~A200;
  assign \new_[87727]_  = A265 & A202;
  assign \new_[87728]_  = \new_[87727]_  & \new_[87724]_ ;
  assign \new_[87729]_  = \new_[87728]_  & \new_[87721]_ ;
  assign \new_[87732]_  = A267 & ~A266;
  assign \new_[87735]_  = A298 & A268;
  assign \new_[87736]_  = \new_[87735]_  & \new_[87732]_ ;
  assign \new_[87739]_  = ~A300 & ~A299;
  assign \new_[87742]_  = A302 & ~A301;
  assign \new_[87743]_  = \new_[87742]_  & \new_[87739]_ ;
  assign \new_[87744]_  = \new_[87743]_  & \new_[87736]_ ;
  assign \new_[87748]_  = A199 & ~A168;
  assign \new_[87749]_  = A169 & \new_[87748]_ ;
  assign \new_[87752]_  = A201 & ~A200;
  assign \new_[87755]_  = A265 & A202;
  assign \new_[87756]_  = \new_[87755]_  & \new_[87752]_ ;
  assign \new_[87757]_  = \new_[87756]_  & \new_[87749]_ ;
  assign \new_[87760]_  = A267 & ~A266;
  assign \new_[87763]_  = ~A298 & A268;
  assign \new_[87764]_  = \new_[87763]_  & \new_[87760]_ ;
  assign \new_[87767]_  = ~A300 & A299;
  assign \new_[87770]_  = A302 & ~A301;
  assign \new_[87771]_  = \new_[87770]_  & \new_[87767]_ ;
  assign \new_[87772]_  = \new_[87771]_  & \new_[87764]_ ;
  assign \new_[87776]_  = A199 & ~A168;
  assign \new_[87777]_  = A169 & \new_[87776]_ ;
  assign \new_[87780]_  = A201 & ~A200;
  assign \new_[87783]_  = A265 & A202;
  assign \new_[87784]_  = \new_[87783]_  & \new_[87780]_ ;
  assign \new_[87785]_  = \new_[87784]_  & \new_[87777]_ ;
  assign \new_[87788]_  = A267 & ~A266;
  assign \new_[87791]_  = A298 & ~A269;
  assign \new_[87792]_  = \new_[87791]_  & \new_[87788]_ ;
  assign \new_[87795]_  = ~A300 & ~A299;
  assign \new_[87798]_  = A302 & ~A301;
  assign \new_[87799]_  = \new_[87798]_  & \new_[87795]_ ;
  assign \new_[87800]_  = \new_[87799]_  & \new_[87792]_ ;
  assign \new_[87804]_  = A199 & ~A168;
  assign \new_[87805]_  = A169 & \new_[87804]_ ;
  assign \new_[87808]_  = A201 & ~A200;
  assign \new_[87811]_  = A265 & A202;
  assign \new_[87812]_  = \new_[87811]_  & \new_[87808]_ ;
  assign \new_[87813]_  = \new_[87812]_  & \new_[87805]_ ;
  assign \new_[87816]_  = A267 & ~A266;
  assign \new_[87819]_  = ~A298 & ~A269;
  assign \new_[87820]_  = \new_[87819]_  & \new_[87816]_ ;
  assign \new_[87823]_  = ~A300 & A299;
  assign \new_[87826]_  = A302 & ~A301;
  assign \new_[87827]_  = \new_[87826]_  & \new_[87823]_ ;
  assign \new_[87828]_  = \new_[87827]_  & \new_[87820]_ ;
  assign \new_[87832]_  = A199 & ~A168;
  assign \new_[87833]_  = A169 & \new_[87832]_ ;
  assign \new_[87836]_  = A201 & ~A200;
  assign \new_[87839]_  = A265 & A202;
  assign \new_[87840]_  = \new_[87839]_  & \new_[87836]_ ;
  assign \new_[87841]_  = \new_[87840]_  & \new_[87833]_ ;
  assign \new_[87844]_  = ~A267 & ~A266;
  assign \new_[87847]_  = A269 & ~A268;
  assign \new_[87848]_  = \new_[87847]_  & \new_[87844]_ ;
  assign \new_[87851]_  = ~A299 & A298;
  assign \new_[87854]_  = A301 & A300;
  assign \new_[87855]_  = \new_[87854]_  & \new_[87851]_ ;
  assign \new_[87856]_  = \new_[87855]_  & \new_[87848]_ ;
  assign \new_[87860]_  = A199 & ~A168;
  assign \new_[87861]_  = A169 & \new_[87860]_ ;
  assign \new_[87864]_  = A201 & ~A200;
  assign \new_[87867]_  = A265 & A202;
  assign \new_[87868]_  = \new_[87867]_  & \new_[87864]_ ;
  assign \new_[87869]_  = \new_[87868]_  & \new_[87861]_ ;
  assign \new_[87872]_  = ~A267 & ~A266;
  assign \new_[87875]_  = A269 & ~A268;
  assign \new_[87876]_  = \new_[87875]_  & \new_[87872]_ ;
  assign \new_[87879]_  = ~A299 & A298;
  assign \new_[87882]_  = ~A302 & A300;
  assign \new_[87883]_  = \new_[87882]_  & \new_[87879]_ ;
  assign \new_[87884]_  = \new_[87883]_  & \new_[87876]_ ;
  assign \new_[87888]_  = A199 & ~A168;
  assign \new_[87889]_  = A169 & \new_[87888]_ ;
  assign \new_[87892]_  = A201 & ~A200;
  assign \new_[87895]_  = A265 & A202;
  assign \new_[87896]_  = \new_[87895]_  & \new_[87892]_ ;
  assign \new_[87897]_  = \new_[87896]_  & \new_[87889]_ ;
  assign \new_[87900]_  = ~A267 & ~A266;
  assign \new_[87903]_  = A269 & ~A268;
  assign \new_[87904]_  = \new_[87903]_  & \new_[87900]_ ;
  assign \new_[87907]_  = A299 & ~A298;
  assign \new_[87910]_  = A301 & A300;
  assign \new_[87911]_  = \new_[87910]_  & \new_[87907]_ ;
  assign \new_[87912]_  = \new_[87911]_  & \new_[87904]_ ;
  assign \new_[87916]_  = A199 & ~A168;
  assign \new_[87917]_  = A169 & \new_[87916]_ ;
  assign \new_[87920]_  = A201 & ~A200;
  assign \new_[87923]_  = A265 & A202;
  assign \new_[87924]_  = \new_[87923]_  & \new_[87920]_ ;
  assign \new_[87925]_  = \new_[87924]_  & \new_[87917]_ ;
  assign \new_[87928]_  = ~A267 & ~A266;
  assign \new_[87931]_  = A269 & ~A268;
  assign \new_[87932]_  = \new_[87931]_  & \new_[87928]_ ;
  assign \new_[87935]_  = A299 & ~A298;
  assign \new_[87938]_  = ~A302 & A300;
  assign \new_[87939]_  = \new_[87938]_  & \new_[87935]_ ;
  assign \new_[87940]_  = \new_[87939]_  & \new_[87932]_ ;
  assign \new_[87944]_  = A199 & ~A168;
  assign \new_[87945]_  = A169 & \new_[87944]_ ;
  assign \new_[87948]_  = A201 & ~A200;
  assign \new_[87951]_  = ~A265 & ~A203;
  assign \new_[87952]_  = \new_[87951]_  & \new_[87948]_ ;
  assign \new_[87953]_  = \new_[87952]_  & \new_[87945]_ ;
  assign \new_[87956]_  = A267 & A266;
  assign \new_[87959]_  = A298 & A268;
  assign \new_[87960]_  = \new_[87959]_  & \new_[87956]_ ;
  assign \new_[87963]_  = ~A300 & ~A299;
  assign \new_[87966]_  = A302 & ~A301;
  assign \new_[87967]_  = \new_[87966]_  & \new_[87963]_ ;
  assign \new_[87968]_  = \new_[87967]_  & \new_[87960]_ ;
  assign \new_[87972]_  = A199 & ~A168;
  assign \new_[87973]_  = A169 & \new_[87972]_ ;
  assign \new_[87976]_  = A201 & ~A200;
  assign \new_[87979]_  = ~A265 & ~A203;
  assign \new_[87980]_  = \new_[87979]_  & \new_[87976]_ ;
  assign \new_[87981]_  = \new_[87980]_  & \new_[87973]_ ;
  assign \new_[87984]_  = A267 & A266;
  assign \new_[87987]_  = ~A298 & A268;
  assign \new_[87988]_  = \new_[87987]_  & \new_[87984]_ ;
  assign \new_[87991]_  = ~A300 & A299;
  assign \new_[87994]_  = A302 & ~A301;
  assign \new_[87995]_  = \new_[87994]_  & \new_[87991]_ ;
  assign \new_[87996]_  = \new_[87995]_  & \new_[87988]_ ;
  assign \new_[88000]_  = A199 & ~A168;
  assign \new_[88001]_  = A169 & \new_[88000]_ ;
  assign \new_[88004]_  = A201 & ~A200;
  assign \new_[88007]_  = ~A265 & ~A203;
  assign \new_[88008]_  = \new_[88007]_  & \new_[88004]_ ;
  assign \new_[88009]_  = \new_[88008]_  & \new_[88001]_ ;
  assign \new_[88012]_  = A267 & A266;
  assign \new_[88015]_  = A298 & ~A269;
  assign \new_[88016]_  = \new_[88015]_  & \new_[88012]_ ;
  assign \new_[88019]_  = ~A300 & ~A299;
  assign \new_[88022]_  = A302 & ~A301;
  assign \new_[88023]_  = \new_[88022]_  & \new_[88019]_ ;
  assign \new_[88024]_  = \new_[88023]_  & \new_[88016]_ ;
  assign \new_[88028]_  = A199 & ~A168;
  assign \new_[88029]_  = A169 & \new_[88028]_ ;
  assign \new_[88032]_  = A201 & ~A200;
  assign \new_[88035]_  = ~A265 & ~A203;
  assign \new_[88036]_  = \new_[88035]_  & \new_[88032]_ ;
  assign \new_[88037]_  = \new_[88036]_  & \new_[88029]_ ;
  assign \new_[88040]_  = A267 & A266;
  assign \new_[88043]_  = ~A298 & ~A269;
  assign \new_[88044]_  = \new_[88043]_  & \new_[88040]_ ;
  assign \new_[88047]_  = ~A300 & A299;
  assign \new_[88050]_  = A302 & ~A301;
  assign \new_[88051]_  = \new_[88050]_  & \new_[88047]_ ;
  assign \new_[88052]_  = \new_[88051]_  & \new_[88044]_ ;
  assign \new_[88056]_  = A199 & ~A168;
  assign \new_[88057]_  = A169 & \new_[88056]_ ;
  assign \new_[88060]_  = A201 & ~A200;
  assign \new_[88063]_  = ~A265 & ~A203;
  assign \new_[88064]_  = \new_[88063]_  & \new_[88060]_ ;
  assign \new_[88065]_  = \new_[88064]_  & \new_[88057]_ ;
  assign \new_[88068]_  = ~A267 & A266;
  assign \new_[88071]_  = A269 & ~A268;
  assign \new_[88072]_  = \new_[88071]_  & \new_[88068]_ ;
  assign \new_[88075]_  = ~A299 & A298;
  assign \new_[88078]_  = A301 & A300;
  assign \new_[88079]_  = \new_[88078]_  & \new_[88075]_ ;
  assign \new_[88080]_  = \new_[88079]_  & \new_[88072]_ ;
  assign \new_[88084]_  = A199 & ~A168;
  assign \new_[88085]_  = A169 & \new_[88084]_ ;
  assign \new_[88088]_  = A201 & ~A200;
  assign \new_[88091]_  = ~A265 & ~A203;
  assign \new_[88092]_  = \new_[88091]_  & \new_[88088]_ ;
  assign \new_[88093]_  = \new_[88092]_  & \new_[88085]_ ;
  assign \new_[88096]_  = ~A267 & A266;
  assign \new_[88099]_  = A269 & ~A268;
  assign \new_[88100]_  = \new_[88099]_  & \new_[88096]_ ;
  assign \new_[88103]_  = ~A299 & A298;
  assign \new_[88106]_  = ~A302 & A300;
  assign \new_[88107]_  = \new_[88106]_  & \new_[88103]_ ;
  assign \new_[88108]_  = \new_[88107]_  & \new_[88100]_ ;
  assign \new_[88112]_  = A199 & ~A168;
  assign \new_[88113]_  = A169 & \new_[88112]_ ;
  assign \new_[88116]_  = A201 & ~A200;
  assign \new_[88119]_  = ~A265 & ~A203;
  assign \new_[88120]_  = \new_[88119]_  & \new_[88116]_ ;
  assign \new_[88121]_  = \new_[88120]_  & \new_[88113]_ ;
  assign \new_[88124]_  = ~A267 & A266;
  assign \new_[88127]_  = A269 & ~A268;
  assign \new_[88128]_  = \new_[88127]_  & \new_[88124]_ ;
  assign \new_[88131]_  = A299 & ~A298;
  assign \new_[88134]_  = A301 & A300;
  assign \new_[88135]_  = \new_[88134]_  & \new_[88131]_ ;
  assign \new_[88136]_  = \new_[88135]_  & \new_[88128]_ ;
  assign \new_[88140]_  = A199 & ~A168;
  assign \new_[88141]_  = A169 & \new_[88140]_ ;
  assign \new_[88144]_  = A201 & ~A200;
  assign \new_[88147]_  = ~A265 & ~A203;
  assign \new_[88148]_  = \new_[88147]_  & \new_[88144]_ ;
  assign \new_[88149]_  = \new_[88148]_  & \new_[88141]_ ;
  assign \new_[88152]_  = ~A267 & A266;
  assign \new_[88155]_  = A269 & ~A268;
  assign \new_[88156]_  = \new_[88155]_  & \new_[88152]_ ;
  assign \new_[88159]_  = A299 & ~A298;
  assign \new_[88162]_  = ~A302 & A300;
  assign \new_[88163]_  = \new_[88162]_  & \new_[88159]_ ;
  assign \new_[88164]_  = \new_[88163]_  & \new_[88156]_ ;
  assign \new_[88168]_  = A199 & ~A168;
  assign \new_[88169]_  = A169 & \new_[88168]_ ;
  assign \new_[88172]_  = A201 & ~A200;
  assign \new_[88175]_  = A265 & ~A203;
  assign \new_[88176]_  = \new_[88175]_  & \new_[88172]_ ;
  assign \new_[88177]_  = \new_[88176]_  & \new_[88169]_ ;
  assign \new_[88180]_  = A267 & ~A266;
  assign \new_[88183]_  = A298 & A268;
  assign \new_[88184]_  = \new_[88183]_  & \new_[88180]_ ;
  assign \new_[88187]_  = ~A300 & ~A299;
  assign \new_[88190]_  = A302 & ~A301;
  assign \new_[88191]_  = \new_[88190]_  & \new_[88187]_ ;
  assign \new_[88192]_  = \new_[88191]_  & \new_[88184]_ ;
  assign \new_[88196]_  = A199 & ~A168;
  assign \new_[88197]_  = A169 & \new_[88196]_ ;
  assign \new_[88200]_  = A201 & ~A200;
  assign \new_[88203]_  = A265 & ~A203;
  assign \new_[88204]_  = \new_[88203]_  & \new_[88200]_ ;
  assign \new_[88205]_  = \new_[88204]_  & \new_[88197]_ ;
  assign \new_[88208]_  = A267 & ~A266;
  assign \new_[88211]_  = ~A298 & A268;
  assign \new_[88212]_  = \new_[88211]_  & \new_[88208]_ ;
  assign \new_[88215]_  = ~A300 & A299;
  assign \new_[88218]_  = A302 & ~A301;
  assign \new_[88219]_  = \new_[88218]_  & \new_[88215]_ ;
  assign \new_[88220]_  = \new_[88219]_  & \new_[88212]_ ;
  assign \new_[88224]_  = A199 & ~A168;
  assign \new_[88225]_  = A169 & \new_[88224]_ ;
  assign \new_[88228]_  = A201 & ~A200;
  assign \new_[88231]_  = A265 & ~A203;
  assign \new_[88232]_  = \new_[88231]_  & \new_[88228]_ ;
  assign \new_[88233]_  = \new_[88232]_  & \new_[88225]_ ;
  assign \new_[88236]_  = A267 & ~A266;
  assign \new_[88239]_  = A298 & ~A269;
  assign \new_[88240]_  = \new_[88239]_  & \new_[88236]_ ;
  assign \new_[88243]_  = ~A300 & ~A299;
  assign \new_[88246]_  = A302 & ~A301;
  assign \new_[88247]_  = \new_[88246]_  & \new_[88243]_ ;
  assign \new_[88248]_  = \new_[88247]_  & \new_[88240]_ ;
  assign \new_[88252]_  = A199 & ~A168;
  assign \new_[88253]_  = A169 & \new_[88252]_ ;
  assign \new_[88256]_  = A201 & ~A200;
  assign \new_[88259]_  = A265 & ~A203;
  assign \new_[88260]_  = \new_[88259]_  & \new_[88256]_ ;
  assign \new_[88261]_  = \new_[88260]_  & \new_[88253]_ ;
  assign \new_[88264]_  = A267 & ~A266;
  assign \new_[88267]_  = ~A298 & ~A269;
  assign \new_[88268]_  = \new_[88267]_  & \new_[88264]_ ;
  assign \new_[88271]_  = ~A300 & A299;
  assign \new_[88274]_  = A302 & ~A301;
  assign \new_[88275]_  = \new_[88274]_  & \new_[88271]_ ;
  assign \new_[88276]_  = \new_[88275]_  & \new_[88268]_ ;
  assign \new_[88280]_  = A199 & ~A168;
  assign \new_[88281]_  = A169 & \new_[88280]_ ;
  assign \new_[88284]_  = A201 & ~A200;
  assign \new_[88287]_  = A265 & ~A203;
  assign \new_[88288]_  = \new_[88287]_  & \new_[88284]_ ;
  assign \new_[88289]_  = \new_[88288]_  & \new_[88281]_ ;
  assign \new_[88292]_  = ~A267 & ~A266;
  assign \new_[88295]_  = A269 & ~A268;
  assign \new_[88296]_  = \new_[88295]_  & \new_[88292]_ ;
  assign \new_[88299]_  = ~A299 & A298;
  assign \new_[88302]_  = A301 & A300;
  assign \new_[88303]_  = \new_[88302]_  & \new_[88299]_ ;
  assign \new_[88304]_  = \new_[88303]_  & \new_[88296]_ ;
  assign \new_[88308]_  = A199 & ~A168;
  assign \new_[88309]_  = A169 & \new_[88308]_ ;
  assign \new_[88312]_  = A201 & ~A200;
  assign \new_[88315]_  = A265 & ~A203;
  assign \new_[88316]_  = \new_[88315]_  & \new_[88312]_ ;
  assign \new_[88317]_  = \new_[88316]_  & \new_[88309]_ ;
  assign \new_[88320]_  = ~A267 & ~A266;
  assign \new_[88323]_  = A269 & ~A268;
  assign \new_[88324]_  = \new_[88323]_  & \new_[88320]_ ;
  assign \new_[88327]_  = ~A299 & A298;
  assign \new_[88330]_  = ~A302 & A300;
  assign \new_[88331]_  = \new_[88330]_  & \new_[88327]_ ;
  assign \new_[88332]_  = \new_[88331]_  & \new_[88324]_ ;
  assign \new_[88336]_  = A199 & ~A168;
  assign \new_[88337]_  = A169 & \new_[88336]_ ;
  assign \new_[88340]_  = A201 & ~A200;
  assign \new_[88343]_  = A265 & ~A203;
  assign \new_[88344]_  = \new_[88343]_  & \new_[88340]_ ;
  assign \new_[88345]_  = \new_[88344]_  & \new_[88337]_ ;
  assign \new_[88348]_  = ~A267 & ~A266;
  assign \new_[88351]_  = A269 & ~A268;
  assign \new_[88352]_  = \new_[88351]_  & \new_[88348]_ ;
  assign \new_[88355]_  = A299 & ~A298;
  assign \new_[88358]_  = A301 & A300;
  assign \new_[88359]_  = \new_[88358]_  & \new_[88355]_ ;
  assign \new_[88360]_  = \new_[88359]_  & \new_[88352]_ ;
  assign \new_[88364]_  = A199 & ~A168;
  assign \new_[88365]_  = A169 & \new_[88364]_ ;
  assign \new_[88368]_  = A201 & ~A200;
  assign \new_[88371]_  = A265 & ~A203;
  assign \new_[88372]_  = \new_[88371]_  & \new_[88368]_ ;
  assign \new_[88373]_  = \new_[88372]_  & \new_[88365]_ ;
  assign \new_[88376]_  = ~A267 & ~A266;
  assign \new_[88379]_  = A269 & ~A268;
  assign \new_[88380]_  = \new_[88379]_  & \new_[88376]_ ;
  assign \new_[88383]_  = A299 & ~A298;
  assign \new_[88386]_  = ~A302 & A300;
  assign \new_[88387]_  = \new_[88386]_  & \new_[88383]_ ;
  assign \new_[88388]_  = \new_[88387]_  & \new_[88380]_ ;
  assign \new_[88392]_  = A199 & ~A168;
  assign \new_[88393]_  = A169 & \new_[88392]_ ;
  assign \new_[88396]_  = ~A201 & ~A200;
  assign \new_[88399]_  = A203 & ~A202;
  assign \new_[88400]_  = \new_[88399]_  & \new_[88396]_ ;
  assign \new_[88401]_  = \new_[88400]_  & \new_[88393]_ ;
  assign \new_[88404]_  = A266 & ~A265;
  assign \new_[88407]_  = A268 & A267;
  assign \new_[88408]_  = \new_[88407]_  & \new_[88404]_ ;
  assign \new_[88411]_  = ~A299 & A298;
  assign \new_[88414]_  = A301 & A300;
  assign \new_[88415]_  = \new_[88414]_  & \new_[88411]_ ;
  assign \new_[88416]_  = \new_[88415]_  & \new_[88408]_ ;
  assign \new_[88420]_  = A199 & ~A168;
  assign \new_[88421]_  = A169 & \new_[88420]_ ;
  assign \new_[88424]_  = ~A201 & ~A200;
  assign \new_[88427]_  = A203 & ~A202;
  assign \new_[88428]_  = \new_[88427]_  & \new_[88424]_ ;
  assign \new_[88429]_  = \new_[88428]_  & \new_[88421]_ ;
  assign \new_[88432]_  = A266 & ~A265;
  assign \new_[88435]_  = A268 & A267;
  assign \new_[88436]_  = \new_[88435]_  & \new_[88432]_ ;
  assign \new_[88439]_  = ~A299 & A298;
  assign \new_[88442]_  = ~A302 & A300;
  assign \new_[88443]_  = \new_[88442]_  & \new_[88439]_ ;
  assign \new_[88444]_  = \new_[88443]_  & \new_[88436]_ ;
  assign \new_[88448]_  = A199 & ~A168;
  assign \new_[88449]_  = A169 & \new_[88448]_ ;
  assign \new_[88452]_  = ~A201 & ~A200;
  assign \new_[88455]_  = A203 & ~A202;
  assign \new_[88456]_  = \new_[88455]_  & \new_[88452]_ ;
  assign \new_[88457]_  = \new_[88456]_  & \new_[88449]_ ;
  assign \new_[88460]_  = A266 & ~A265;
  assign \new_[88463]_  = A268 & A267;
  assign \new_[88464]_  = \new_[88463]_  & \new_[88460]_ ;
  assign \new_[88467]_  = A299 & ~A298;
  assign \new_[88470]_  = A301 & A300;
  assign \new_[88471]_  = \new_[88470]_  & \new_[88467]_ ;
  assign \new_[88472]_  = \new_[88471]_  & \new_[88464]_ ;
  assign \new_[88476]_  = A199 & ~A168;
  assign \new_[88477]_  = A169 & \new_[88476]_ ;
  assign \new_[88480]_  = ~A201 & ~A200;
  assign \new_[88483]_  = A203 & ~A202;
  assign \new_[88484]_  = \new_[88483]_  & \new_[88480]_ ;
  assign \new_[88485]_  = \new_[88484]_  & \new_[88477]_ ;
  assign \new_[88488]_  = A266 & ~A265;
  assign \new_[88491]_  = A268 & A267;
  assign \new_[88492]_  = \new_[88491]_  & \new_[88488]_ ;
  assign \new_[88495]_  = A299 & ~A298;
  assign \new_[88498]_  = ~A302 & A300;
  assign \new_[88499]_  = \new_[88498]_  & \new_[88495]_ ;
  assign \new_[88500]_  = \new_[88499]_  & \new_[88492]_ ;
  assign \new_[88504]_  = A199 & ~A168;
  assign \new_[88505]_  = A169 & \new_[88504]_ ;
  assign \new_[88508]_  = ~A201 & ~A200;
  assign \new_[88511]_  = A203 & ~A202;
  assign \new_[88512]_  = \new_[88511]_  & \new_[88508]_ ;
  assign \new_[88513]_  = \new_[88512]_  & \new_[88505]_ ;
  assign \new_[88516]_  = A266 & ~A265;
  assign \new_[88519]_  = ~A269 & A267;
  assign \new_[88520]_  = \new_[88519]_  & \new_[88516]_ ;
  assign \new_[88523]_  = ~A299 & A298;
  assign \new_[88526]_  = A301 & A300;
  assign \new_[88527]_  = \new_[88526]_  & \new_[88523]_ ;
  assign \new_[88528]_  = \new_[88527]_  & \new_[88520]_ ;
  assign \new_[88532]_  = A199 & ~A168;
  assign \new_[88533]_  = A169 & \new_[88532]_ ;
  assign \new_[88536]_  = ~A201 & ~A200;
  assign \new_[88539]_  = A203 & ~A202;
  assign \new_[88540]_  = \new_[88539]_  & \new_[88536]_ ;
  assign \new_[88541]_  = \new_[88540]_  & \new_[88533]_ ;
  assign \new_[88544]_  = A266 & ~A265;
  assign \new_[88547]_  = ~A269 & A267;
  assign \new_[88548]_  = \new_[88547]_  & \new_[88544]_ ;
  assign \new_[88551]_  = ~A299 & A298;
  assign \new_[88554]_  = ~A302 & A300;
  assign \new_[88555]_  = \new_[88554]_  & \new_[88551]_ ;
  assign \new_[88556]_  = \new_[88555]_  & \new_[88548]_ ;
  assign \new_[88560]_  = A199 & ~A168;
  assign \new_[88561]_  = A169 & \new_[88560]_ ;
  assign \new_[88564]_  = ~A201 & ~A200;
  assign \new_[88567]_  = A203 & ~A202;
  assign \new_[88568]_  = \new_[88567]_  & \new_[88564]_ ;
  assign \new_[88569]_  = \new_[88568]_  & \new_[88561]_ ;
  assign \new_[88572]_  = A266 & ~A265;
  assign \new_[88575]_  = ~A269 & A267;
  assign \new_[88576]_  = \new_[88575]_  & \new_[88572]_ ;
  assign \new_[88579]_  = A299 & ~A298;
  assign \new_[88582]_  = A301 & A300;
  assign \new_[88583]_  = \new_[88582]_  & \new_[88579]_ ;
  assign \new_[88584]_  = \new_[88583]_  & \new_[88576]_ ;
  assign \new_[88588]_  = A199 & ~A168;
  assign \new_[88589]_  = A169 & \new_[88588]_ ;
  assign \new_[88592]_  = ~A201 & ~A200;
  assign \new_[88595]_  = A203 & ~A202;
  assign \new_[88596]_  = \new_[88595]_  & \new_[88592]_ ;
  assign \new_[88597]_  = \new_[88596]_  & \new_[88589]_ ;
  assign \new_[88600]_  = A266 & ~A265;
  assign \new_[88603]_  = ~A269 & A267;
  assign \new_[88604]_  = \new_[88603]_  & \new_[88600]_ ;
  assign \new_[88607]_  = A299 & ~A298;
  assign \new_[88610]_  = ~A302 & A300;
  assign \new_[88611]_  = \new_[88610]_  & \new_[88607]_ ;
  assign \new_[88612]_  = \new_[88611]_  & \new_[88604]_ ;
  assign \new_[88616]_  = A199 & ~A168;
  assign \new_[88617]_  = A169 & \new_[88616]_ ;
  assign \new_[88620]_  = ~A201 & ~A200;
  assign \new_[88623]_  = A203 & ~A202;
  assign \new_[88624]_  = \new_[88623]_  & \new_[88620]_ ;
  assign \new_[88625]_  = \new_[88624]_  & \new_[88617]_ ;
  assign \new_[88628]_  = ~A266 & A265;
  assign \new_[88631]_  = A268 & A267;
  assign \new_[88632]_  = \new_[88631]_  & \new_[88628]_ ;
  assign \new_[88635]_  = ~A299 & A298;
  assign \new_[88638]_  = A301 & A300;
  assign \new_[88639]_  = \new_[88638]_  & \new_[88635]_ ;
  assign \new_[88640]_  = \new_[88639]_  & \new_[88632]_ ;
  assign \new_[88644]_  = A199 & ~A168;
  assign \new_[88645]_  = A169 & \new_[88644]_ ;
  assign \new_[88648]_  = ~A201 & ~A200;
  assign \new_[88651]_  = A203 & ~A202;
  assign \new_[88652]_  = \new_[88651]_  & \new_[88648]_ ;
  assign \new_[88653]_  = \new_[88652]_  & \new_[88645]_ ;
  assign \new_[88656]_  = ~A266 & A265;
  assign \new_[88659]_  = A268 & A267;
  assign \new_[88660]_  = \new_[88659]_  & \new_[88656]_ ;
  assign \new_[88663]_  = ~A299 & A298;
  assign \new_[88666]_  = ~A302 & A300;
  assign \new_[88667]_  = \new_[88666]_  & \new_[88663]_ ;
  assign \new_[88668]_  = \new_[88667]_  & \new_[88660]_ ;
  assign \new_[88672]_  = A199 & ~A168;
  assign \new_[88673]_  = A169 & \new_[88672]_ ;
  assign \new_[88676]_  = ~A201 & ~A200;
  assign \new_[88679]_  = A203 & ~A202;
  assign \new_[88680]_  = \new_[88679]_  & \new_[88676]_ ;
  assign \new_[88681]_  = \new_[88680]_  & \new_[88673]_ ;
  assign \new_[88684]_  = ~A266 & A265;
  assign \new_[88687]_  = A268 & A267;
  assign \new_[88688]_  = \new_[88687]_  & \new_[88684]_ ;
  assign \new_[88691]_  = A299 & ~A298;
  assign \new_[88694]_  = A301 & A300;
  assign \new_[88695]_  = \new_[88694]_  & \new_[88691]_ ;
  assign \new_[88696]_  = \new_[88695]_  & \new_[88688]_ ;
  assign \new_[88700]_  = A199 & ~A168;
  assign \new_[88701]_  = A169 & \new_[88700]_ ;
  assign \new_[88704]_  = ~A201 & ~A200;
  assign \new_[88707]_  = A203 & ~A202;
  assign \new_[88708]_  = \new_[88707]_  & \new_[88704]_ ;
  assign \new_[88709]_  = \new_[88708]_  & \new_[88701]_ ;
  assign \new_[88712]_  = ~A266 & A265;
  assign \new_[88715]_  = A268 & A267;
  assign \new_[88716]_  = \new_[88715]_  & \new_[88712]_ ;
  assign \new_[88719]_  = A299 & ~A298;
  assign \new_[88722]_  = ~A302 & A300;
  assign \new_[88723]_  = \new_[88722]_  & \new_[88719]_ ;
  assign \new_[88724]_  = \new_[88723]_  & \new_[88716]_ ;
  assign \new_[88728]_  = A199 & ~A168;
  assign \new_[88729]_  = A169 & \new_[88728]_ ;
  assign \new_[88732]_  = ~A201 & ~A200;
  assign \new_[88735]_  = A203 & ~A202;
  assign \new_[88736]_  = \new_[88735]_  & \new_[88732]_ ;
  assign \new_[88737]_  = \new_[88736]_  & \new_[88729]_ ;
  assign \new_[88740]_  = ~A266 & A265;
  assign \new_[88743]_  = ~A269 & A267;
  assign \new_[88744]_  = \new_[88743]_  & \new_[88740]_ ;
  assign \new_[88747]_  = ~A299 & A298;
  assign \new_[88750]_  = A301 & A300;
  assign \new_[88751]_  = \new_[88750]_  & \new_[88747]_ ;
  assign \new_[88752]_  = \new_[88751]_  & \new_[88744]_ ;
  assign \new_[88756]_  = A199 & ~A168;
  assign \new_[88757]_  = A169 & \new_[88756]_ ;
  assign \new_[88760]_  = ~A201 & ~A200;
  assign \new_[88763]_  = A203 & ~A202;
  assign \new_[88764]_  = \new_[88763]_  & \new_[88760]_ ;
  assign \new_[88765]_  = \new_[88764]_  & \new_[88757]_ ;
  assign \new_[88768]_  = ~A266 & A265;
  assign \new_[88771]_  = ~A269 & A267;
  assign \new_[88772]_  = \new_[88771]_  & \new_[88768]_ ;
  assign \new_[88775]_  = ~A299 & A298;
  assign \new_[88778]_  = ~A302 & A300;
  assign \new_[88779]_  = \new_[88778]_  & \new_[88775]_ ;
  assign \new_[88780]_  = \new_[88779]_  & \new_[88772]_ ;
  assign \new_[88784]_  = A199 & ~A168;
  assign \new_[88785]_  = A169 & \new_[88784]_ ;
  assign \new_[88788]_  = ~A201 & ~A200;
  assign \new_[88791]_  = A203 & ~A202;
  assign \new_[88792]_  = \new_[88791]_  & \new_[88788]_ ;
  assign \new_[88793]_  = \new_[88792]_  & \new_[88785]_ ;
  assign \new_[88796]_  = ~A266 & A265;
  assign \new_[88799]_  = ~A269 & A267;
  assign \new_[88800]_  = \new_[88799]_  & \new_[88796]_ ;
  assign \new_[88803]_  = A299 & ~A298;
  assign \new_[88806]_  = A301 & A300;
  assign \new_[88807]_  = \new_[88806]_  & \new_[88803]_ ;
  assign \new_[88808]_  = \new_[88807]_  & \new_[88800]_ ;
  assign \new_[88812]_  = A199 & ~A168;
  assign \new_[88813]_  = A169 & \new_[88812]_ ;
  assign \new_[88816]_  = ~A201 & ~A200;
  assign \new_[88819]_  = A203 & ~A202;
  assign \new_[88820]_  = \new_[88819]_  & \new_[88816]_ ;
  assign \new_[88821]_  = \new_[88820]_  & \new_[88813]_ ;
  assign \new_[88824]_  = ~A266 & A265;
  assign \new_[88827]_  = ~A269 & A267;
  assign \new_[88828]_  = \new_[88827]_  & \new_[88824]_ ;
  assign \new_[88831]_  = A299 & ~A298;
  assign \new_[88834]_  = ~A302 & A300;
  assign \new_[88835]_  = \new_[88834]_  & \new_[88831]_ ;
  assign \new_[88836]_  = \new_[88835]_  & \new_[88828]_ ;
  assign \new_[88840]_  = A168 & ~A169;
  assign \new_[88841]_  = ~A170 & \new_[88840]_ ;
  assign \new_[88844]_  = A200 & ~A199;
  assign \new_[88847]_  = A202 & A201;
  assign \new_[88848]_  = \new_[88847]_  & \new_[88844]_ ;
  assign \new_[88849]_  = \new_[88848]_  & \new_[88841]_ ;
  assign \new_[88852]_  = A266 & ~A265;
  assign \new_[88855]_  = A268 & A267;
  assign \new_[88856]_  = \new_[88855]_  & \new_[88852]_ ;
  assign \new_[88859]_  = ~A299 & A298;
  assign \new_[88862]_  = A301 & A300;
  assign \new_[88863]_  = \new_[88862]_  & \new_[88859]_ ;
  assign \new_[88864]_  = \new_[88863]_  & \new_[88856]_ ;
  assign \new_[88868]_  = A168 & ~A169;
  assign \new_[88869]_  = ~A170 & \new_[88868]_ ;
  assign \new_[88872]_  = A200 & ~A199;
  assign \new_[88875]_  = A202 & A201;
  assign \new_[88876]_  = \new_[88875]_  & \new_[88872]_ ;
  assign \new_[88877]_  = \new_[88876]_  & \new_[88869]_ ;
  assign \new_[88880]_  = A266 & ~A265;
  assign \new_[88883]_  = A268 & A267;
  assign \new_[88884]_  = \new_[88883]_  & \new_[88880]_ ;
  assign \new_[88887]_  = ~A299 & A298;
  assign \new_[88890]_  = ~A302 & A300;
  assign \new_[88891]_  = \new_[88890]_  & \new_[88887]_ ;
  assign \new_[88892]_  = \new_[88891]_  & \new_[88884]_ ;
  assign \new_[88896]_  = A168 & ~A169;
  assign \new_[88897]_  = ~A170 & \new_[88896]_ ;
  assign \new_[88900]_  = A200 & ~A199;
  assign \new_[88903]_  = A202 & A201;
  assign \new_[88904]_  = \new_[88903]_  & \new_[88900]_ ;
  assign \new_[88905]_  = \new_[88904]_  & \new_[88897]_ ;
  assign \new_[88908]_  = A266 & ~A265;
  assign \new_[88911]_  = A268 & A267;
  assign \new_[88912]_  = \new_[88911]_  & \new_[88908]_ ;
  assign \new_[88915]_  = A299 & ~A298;
  assign \new_[88918]_  = A301 & A300;
  assign \new_[88919]_  = \new_[88918]_  & \new_[88915]_ ;
  assign \new_[88920]_  = \new_[88919]_  & \new_[88912]_ ;
  assign \new_[88924]_  = A168 & ~A169;
  assign \new_[88925]_  = ~A170 & \new_[88924]_ ;
  assign \new_[88928]_  = A200 & ~A199;
  assign \new_[88931]_  = A202 & A201;
  assign \new_[88932]_  = \new_[88931]_  & \new_[88928]_ ;
  assign \new_[88933]_  = \new_[88932]_  & \new_[88925]_ ;
  assign \new_[88936]_  = A266 & ~A265;
  assign \new_[88939]_  = A268 & A267;
  assign \new_[88940]_  = \new_[88939]_  & \new_[88936]_ ;
  assign \new_[88943]_  = A299 & ~A298;
  assign \new_[88946]_  = ~A302 & A300;
  assign \new_[88947]_  = \new_[88946]_  & \new_[88943]_ ;
  assign \new_[88948]_  = \new_[88947]_  & \new_[88940]_ ;
  assign \new_[88952]_  = A168 & ~A169;
  assign \new_[88953]_  = ~A170 & \new_[88952]_ ;
  assign \new_[88956]_  = A200 & ~A199;
  assign \new_[88959]_  = A202 & A201;
  assign \new_[88960]_  = \new_[88959]_  & \new_[88956]_ ;
  assign \new_[88961]_  = \new_[88960]_  & \new_[88953]_ ;
  assign \new_[88964]_  = A266 & ~A265;
  assign \new_[88967]_  = ~A269 & A267;
  assign \new_[88968]_  = \new_[88967]_  & \new_[88964]_ ;
  assign \new_[88971]_  = ~A299 & A298;
  assign \new_[88974]_  = A301 & A300;
  assign \new_[88975]_  = \new_[88974]_  & \new_[88971]_ ;
  assign \new_[88976]_  = \new_[88975]_  & \new_[88968]_ ;
  assign \new_[88980]_  = A168 & ~A169;
  assign \new_[88981]_  = ~A170 & \new_[88980]_ ;
  assign \new_[88984]_  = A200 & ~A199;
  assign \new_[88987]_  = A202 & A201;
  assign \new_[88988]_  = \new_[88987]_  & \new_[88984]_ ;
  assign \new_[88989]_  = \new_[88988]_  & \new_[88981]_ ;
  assign \new_[88992]_  = A266 & ~A265;
  assign \new_[88995]_  = ~A269 & A267;
  assign \new_[88996]_  = \new_[88995]_  & \new_[88992]_ ;
  assign \new_[88999]_  = ~A299 & A298;
  assign \new_[89002]_  = ~A302 & A300;
  assign \new_[89003]_  = \new_[89002]_  & \new_[88999]_ ;
  assign \new_[89004]_  = \new_[89003]_  & \new_[88996]_ ;
  assign \new_[89008]_  = A168 & ~A169;
  assign \new_[89009]_  = ~A170 & \new_[89008]_ ;
  assign \new_[89012]_  = A200 & ~A199;
  assign \new_[89015]_  = A202 & A201;
  assign \new_[89016]_  = \new_[89015]_  & \new_[89012]_ ;
  assign \new_[89017]_  = \new_[89016]_  & \new_[89009]_ ;
  assign \new_[89020]_  = A266 & ~A265;
  assign \new_[89023]_  = ~A269 & A267;
  assign \new_[89024]_  = \new_[89023]_  & \new_[89020]_ ;
  assign \new_[89027]_  = A299 & ~A298;
  assign \new_[89030]_  = A301 & A300;
  assign \new_[89031]_  = \new_[89030]_  & \new_[89027]_ ;
  assign \new_[89032]_  = \new_[89031]_  & \new_[89024]_ ;
  assign \new_[89036]_  = A168 & ~A169;
  assign \new_[89037]_  = ~A170 & \new_[89036]_ ;
  assign \new_[89040]_  = A200 & ~A199;
  assign \new_[89043]_  = A202 & A201;
  assign \new_[89044]_  = \new_[89043]_  & \new_[89040]_ ;
  assign \new_[89045]_  = \new_[89044]_  & \new_[89037]_ ;
  assign \new_[89048]_  = A266 & ~A265;
  assign \new_[89051]_  = ~A269 & A267;
  assign \new_[89052]_  = \new_[89051]_  & \new_[89048]_ ;
  assign \new_[89055]_  = A299 & ~A298;
  assign \new_[89058]_  = ~A302 & A300;
  assign \new_[89059]_  = \new_[89058]_  & \new_[89055]_ ;
  assign \new_[89060]_  = \new_[89059]_  & \new_[89052]_ ;
  assign \new_[89064]_  = A168 & ~A169;
  assign \new_[89065]_  = ~A170 & \new_[89064]_ ;
  assign \new_[89068]_  = A200 & ~A199;
  assign \new_[89071]_  = A202 & A201;
  assign \new_[89072]_  = \new_[89071]_  & \new_[89068]_ ;
  assign \new_[89073]_  = \new_[89072]_  & \new_[89065]_ ;
  assign \new_[89076]_  = ~A266 & A265;
  assign \new_[89079]_  = A268 & A267;
  assign \new_[89080]_  = \new_[89079]_  & \new_[89076]_ ;
  assign \new_[89083]_  = ~A299 & A298;
  assign \new_[89086]_  = A301 & A300;
  assign \new_[89087]_  = \new_[89086]_  & \new_[89083]_ ;
  assign \new_[89088]_  = \new_[89087]_  & \new_[89080]_ ;
  assign \new_[89092]_  = A168 & ~A169;
  assign \new_[89093]_  = ~A170 & \new_[89092]_ ;
  assign \new_[89096]_  = A200 & ~A199;
  assign \new_[89099]_  = A202 & A201;
  assign \new_[89100]_  = \new_[89099]_  & \new_[89096]_ ;
  assign \new_[89101]_  = \new_[89100]_  & \new_[89093]_ ;
  assign \new_[89104]_  = ~A266 & A265;
  assign \new_[89107]_  = A268 & A267;
  assign \new_[89108]_  = \new_[89107]_  & \new_[89104]_ ;
  assign \new_[89111]_  = ~A299 & A298;
  assign \new_[89114]_  = ~A302 & A300;
  assign \new_[89115]_  = \new_[89114]_  & \new_[89111]_ ;
  assign \new_[89116]_  = \new_[89115]_  & \new_[89108]_ ;
  assign \new_[89120]_  = A168 & ~A169;
  assign \new_[89121]_  = ~A170 & \new_[89120]_ ;
  assign \new_[89124]_  = A200 & ~A199;
  assign \new_[89127]_  = A202 & A201;
  assign \new_[89128]_  = \new_[89127]_  & \new_[89124]_ ;
  assign \new_[89129]_  = \new_[89128]_  & \new_[89121]_ ;
  assign \new_[89132]_  = ~A266 & A265;
  assign \new_[89135]_  = A268 & A267;
  assign \new_[89136]_  = \new_[89135]_  & \new_[89132]_ ;
  assign \new_[89139]_  = A299 & ~A298;
  assign \new_[89142]_  = A301 & A300;
  assign \new_[89143]_  = \new_[89142]_  & \new_[89139]_ ;
  assign \new_[89144]_  = \new_[89143]_  & \new_[89136]_ ;
  assign \new_[89148]_  = A168 & ~A169;
  assign \new_[89149]_  = ~A170 & \new_[89148]_ ;
  assign \new_[89152]_  = A200 & ~A199;
  assign \new_[89155]_  = A202 & A201;
  assign \new_[89156]_  = \new_[89155]_  & \new_[89152]_ ;
  assign \new_[89157]_  = \new_[89156]_  & \new_[89149]_ ;
  assign \new_[89160]_  = ~A266 & A265;
  assign \new_[89163]_  = A268 & A267;
  assign \new_[89164]_  = \new_[89163]_  & \new_[89160]_ ;
  assign \new_[89167]_  = A299 & ~A298;
  assign \new_[89170]_  = ~A302 & A300;
  assign \new_[89171]_  = \new_[89170]_  & \new_[89167]_ ;
  assign \new_[89172]_  = \new_[89171]_  & \new_[89164]_ ;
  assign \new_[89176]_  = A168 & ~A169;
  assign \new_[89177]_  = ~A170 & \new_[89176]_ ;
  assign \new_[89180]_  = A200 & ~A199;
  assign \new_[89183]_  = A202 & A201;
  assign \new_[89184]_  = \new_[89183]_  & \new_[89180]_ ;
  assign \new_[89185]_  = \new_[89184]_  & \new_[89177]_ ;
  assign \new_[89188]_  = ~A266 & A265;
  assign \new_[89191]_  = ~A269 & A267;
  assign \new_[89192]_  = \new_[89191]_  & \new_[89188]_ ;
  assign \new_[89195]_  = ~A299 & A298;
  assign \new_[89198]_  = A301 & A300;
  assign \new_[89199]_  = \new_[89198]_  & \new_[89195]_ ;
  assign \new_[89200]_  = \new_[89199]_  & \new_[89192]_ ;
  assign \new_[89204]_  = A168 & ~A169;
  assign \new_[89205]_  = ~A170 & \new_[89204]_ ;
  assign \new_[89208]_  = A200 & ~A199;
  assign \new_[89211]_  = A202 & A201;
  assign \new_[89212]_  = \new_[89211]_  & \new_[89208]_ ;
  assign \new_[89213]_  = \new_[89212]_  & \new_[89205]_ ;
  assign \new_[89216]_  = ~A266 & A265;
  assign \new_[89219]_  = ~A269 & A267;
  assign \new_[89220]_  = \new_[89219]_  & \new_[89216]_ ;
  assign \new_[89223]_  = ~A299 & A298;
  assign \new_[89226]_  = ~A302 & A300;
  assign \new_[89227]_  = \new_[89226]_  & \new_[89223]_ ;
  assign \new_[89228]_  = \new_[89227]_  & \new_[89220]_ ;
  assign \new_[89232]_  = A168 & ~A169;
  assign \new_[89233]_  = ~A170 & \new_[89232]_ ;
  assign \new_[89236]_  = A200 & ~A199;
  assign \new_[89239]_  = A202 & A201;
  assign \new_[89240]_  = \new_[89239]_  & \new_[89236]_ ;
  assign \new_[89241]_  = \new_[89240]_  & \new_[89233]_ ;
  assign \new_[89244]_  = ~A266 & A265;
  assign \new_[89247]_  = ~A269 & A267;
  assign \new_[89248]_  = \new_[89247]_  & \new_[89244]_ ;
  assign \new_[89251]_  = A299 & ~A298;
  assign \new_[89254]_  = A301 & A300;
  assign \new_[89255]_  = \new_[89254]_  & \new_[89251]_ ;
  assign \new_[89256]_  = \new_[89255]_  & \new_[89248]_ ;
  assign \new_[89260]_  = A168 & ~A169;
  assign \new_[89261]_  = ~A170 & \new_[89260]_ ;
  assign \new_[89264]_  = A200 & ~A199;
  assign \new_[89267]_  = A202 & A201;
  assign \new_[89268]_  = \new_[89267]_  & \new_[89264]_ ;
  assign \new_[89269]_  = \new_[89268]_  & \new_[89261]_ ;
  assign \new_[89272]_  = ~A266 & A265;
  assign \new_[89275]_  = ~A269 & A267;
  assign \new_[89276]_  = \new_[89275]_  & \new_[89272]_ ;
  assign \new_[89279]_  = A299 & ~A298;
  assign \new_[89282]_  = ~A302 & A300;
  assign \new_[89283]_  = \new_[89282]_  & \new_[89279]_ ;
  assign \new_[89284]_  = \new_[89283]_  & \new_[89276]_ ;
  assign \new_[89288]_  = A168 & ~A169;
  assign \new_[89289]_  = ~A170 & \new_[89288]_ ;
  assign \new_[89292]_  = A200 & ~A199;
  assign \new_[89295]_  = ~A203 & A201;
  assign \new_[89296]_  = \new_[89295]_  & \new_[89292]_ ;
  assign \new_[89297]_  = \new_[89296]_  & \new_[89289]_ ;
  assign \new_[89300]_  = A266 & ~A265;
  assign \new_[89303]_  = A268 & A267;
  assign \new_[89304]_  = \new_[89303]_  & \new_[89300]_ ;
  assign \new_[89307]_  = ~A299 & A298;
  assign \new_[89310]_  = A301 & A300;
  assign \new_[89311]_  = \new_[89310]_  & \new_[89307]_ ;
  assign \new_[89312]_  = \new_[89311]_  & \new_[89304]_ ;
  assign \new_[89316]_  = A168 & ~A169;
  assign \new_[89317]_  = ~A170 & \new_[89316]_ ;
  assign \new_[89320]_  = A200 & ~A199;
  assign \new_[89323]_  = ~A203 & A201;
  assign \new_[89324]_  = \new_[89323]_  & \new_[89320]_ ;
  assign \new_[89325]_  = \new_[89324]_  & \new_[89317]_ ;
  assign \new_[89328]_  = A266 & ~A265;
  assign \new_[89331]_  = A268 & A267;
  assign \new_[89332]_  = \new_[89331]_  & \new_[89328]_ ;
  assign \new_[89335]_  = ~A299 & A298;
  assign \new_[89338]_  = ~A302 & A300;
  assign \new_[89339]_  = \new_[89338]_  & \new_[89335]_ ;
  assign \new_[89340]_  = \new_[89339]_  & \new_[89332]_ ;
  assign \new_[89344]_  = A168 & ~A169;
  assign \new_[89345]_  = ~A170 & \new_[89344]_ ;
  assign \new_[89348]_  = A200 & ~A199;
  assign \new_[89351]_  = ~A203 & A201;
  assign \new_[89352]_  = \new_[89351]_  & \new_[89348]_ ;
  assign \new_[89353]_  = \new_[89352]_  & \new_[89345]_ ;
  assign \new_[89356]_  = A266 & ~A265;
  assign \new_[89359]_  = A268 & A267;
  assign \new_[89360]_  = \new_[89359]_  & \new_[89356]_ ;
  assign \new_[89363]_  = A299 & ~A298;
  assign \new_[89366]_  = A301 & A300;
  assign \new_[89367]_  = \new_[89366]_  & \new_[89363]_ ;
  assign \new_[89368]_  = \new_[89367]_  & \new_[89360]_ ;
  assign \new_[89372]_  = A168 & ~A169;
  assign \new_[89373]_  = ~A170 & \new_[89372]_ ;
  assign \new_[89376]_  = A200 & ~A199;
  assign \new_[89379]_  = ~A203 & A201;
  assign \new_[89380]_  = \new_[89379]_  & \new_[89376]_ ;
  assign \new_[89381]_  = \new_[89380]_  & \new_[89373]_ ;
  assign \new_[89384]_  = A266 & ~A265;
  assign \new_[89387]_  = A268 & A267;
  assign \new_[89388]_  = \new_[89387]_  & \new_[89384]_ ;
  assign \new_[89391]_  = A299 & ~A298;
  assign \new_[89394]_  = ~A302 & A300;
  assign \new_[89395]_  = \new_[89394]_  & \new_[89391]_ ;
  assign \new_[89396]_  = \new_[89395]_  & \new_[89388]_ ;
  assign \new_[89400]_  = A168 & ~A169;
  assign \new_[89401]_  = ~A170 & \new_[89400]_ ;
  assign \new_[89404]_  = A200 & ~A199;
  assign \new_[89407]_  = ~A203 & A201;
  assign \new_[89408]_  = \new_[89407]_  & \new_[89404]_ ;
  assign \new_[89409]_  = \new_[89408]_  & \new_[89401]_ ;
  assign \new_[89412]_  = A266 & ~A265;
  assign \new_[89415]_  = ~A269 & A267;
  assign \new_[89416]_  = \new_[89415]_  & \new_[89412]_ ;
  assign \new_[89419]_  = ~A299 & A298;
  assign \new_[89422]_  = A301 & A300;
  assign \new_[89423]_  = \new_[89422]_  & \new_[89419]_ ;
  assign \new_[89424]_  = \new_[89423]_  & \new_[89416]_ ;
  assign \new_[89428]_  = A168 & ~A169;
  assign \new_[89429]_  = ~A170 & \new_[89428]_ ;
  assign \new_[89432]_  = A200 & ~A199;
  assign \new_[89435]_  = ~A203 & A201;
  assign \new_[89436]_  = \new_[89435]_  & \new_[89432]_ ;
  assign \new_[89437]_  = \new_[89436]_  & \new_[89429]_ ;
  assign \new_[89440]_  = A266 & ~A265;
  assign \new_[89443]_  = ~A269 & A267;
  assign \new_[89444]_  = \new_[89443]_  & \new_[89440]_ ;
  assign \new_[89447]_  = ~A299 & A298;
  assign \new_[89450]_  = ~A302 & A300;
  assign \new_[89451]_  = \new_[89450]_  & \new_[89447]_ ;
  assign \new_[89452]_  = \new_[89451]_  & \new_[89444]_ ;
  assign \new_[89456]_  = A168 & ~A169;
  assign \new_[89457]_  = ~A170 & \new_[89456]_ ;
  assign \new_[89460]_  = A200 & ~A199;
  assign \new_[89463]_  = ~A203 & A201;
  assign \new_[89464]_  = \new_[89463]_  & \new_[89460]_ ;
  assign \new_[89465]_  = \new_[89464]_  & \new_[89457]_ ;
  assign \new_[89468]_  = A266 & ~A265;
  assign \new_[89471]_  = ~A269 & A267;
  assign \new_[89472]_  = \new_[89471]_  & \new_[89468]_ ;
  assign \new_[89475]_  = A299 & ~A298;
  assign \new_[89478]_  = A301 & A300;
  assign \new_[89479]_  = \new_[89478]_  & \new_[89475]_ ;
  assign \new_[89480]_  = \new_[89479]_  & \new_[89472]_ ;
  assign \new_[89484]_  = A168 & ~A169;
  assign \new_[89485]_  = ~A170 & \new_[89484]_ ;
  assign \new_[89488]_  = A200 & ~A199;
  assign \new_[89491]_  = ~A203 & A201;
  assign \new_[89492]_  = \new_[89491]_  & \new_[89488]_ ;
  assign \new_[89493]_  = \new_[89492]_  & \new_[89485]_ ;
  assign \new_[89496]_  = A266 & ~A265;
  assign \new_[89499]_  = ~A269 & A267;
  assign \new_[89500]_  = \new_[89499]_  & \new_[89496]_ ;
  assign \new_[89503]_  = A299 & ~A298;
  assign \new_[89506]_  = ~A302 & A300;
  assign \new_[89507]_  = \new_[89506]_  & \new_[89503]_ ;
  assign \new_[89508]_  = \new_[89507]_  & \new_[89500]_ ;
  assign \new_[89512]_  = A168 & ~A169;
  assign \new_[89513]_  = ~A170 & \new_[89512]_ ;
  assign \new_[89516]_  = A200 & ~A199;
  assign \new_[89519]_  = ~A203 & A201;
  assign \new_[89520]_  = \new_[89519]_  & \new_[89516]_ ;
  assign \new_[89521]_  = \new_[89520]_  & \new_[89513]_ ;
  assign \new_[89524]_  = ~A266 & A265;
  assign \new_[89527]_  = A268 & A267;
  assign \new_[89528]_  = \new_[89527]_  & \new_[89524]_ ;
  assign \new_[89531]_  = ~A299 & A298;
  assign \new_[89534]_  = A301 & A300;
  assign \new_[89535]_  = \new_[89534]_  & \new_[89531]_ ;
  assign \new_[89536]_  = \new_[89535]_  & \new_[89528]_ ;
  assign \new_[89540]_  = A168 & ~A169;
  assign \new_[89541]_  = ~A170 & \new_[89540]_ ;
  assign \new_[89544]_  = A200 & ~A199;
  assign \new_[89547]_  = ~A203 & A201;
  assign \new_[89548]_  = \new_[89547]_  & \new_[89544]_ ;
  assign \new_[89549]_  = \new_[89548]_  & \new_[89541]_ ;
  assign \new_[89552]_  = ~A266 & A265;
  assign \new_[89555]_  = A268 & A267;
  assign \new_[89556]_  = \new_[89555]_  & \new_[89552]_ ;
  assign \new_[89559]_  = ~A299 & A298;
  assign \new_[89562]_  = ~A302 & A300;
  assign \new_[89563]_  = \new_[89562]_  & \new_[89559]_ ;
  assign \new_[89564]_  = \new_[89563]_  & \new_[89556]_ ;
  assign \new_[89568]_  = A168 & ~A169;
  assign \new_[89569]_  = ~A170 & \new_[89568]_ ;
  assign \new_[89572]_  = A200 & ~A199;
  assign \new_[89575]_  = ~A203 & A201;
  assign \new_[89576]_  = \new_[89575]_  & \new_[89572]_ ;
  assign \new_[89577]_  = \new_[89576]_  & \new_[89569]_ ;
  assign \new_[89580]_  = ~A266 & A265;
  assign \new_[89583]_  = A268 & A267;
  assign \new_[89584]_  = \new_[89583]_  & \new_[89580]_ ;
  assign \new_[89587]_  = A299 & ~A298;
  assign \new_[89590]_  = A301 & A300;
  assign \new_[89591]_  = \new_[89590]_  & \new_[89587]_ ;
  assign \new_[89592]_  = \new_[89591]_  & \new_[89584]_ ;
  assign \new_[89596]_  = A168 & ~A169;
  assign \new_[89597]_  = ~A170 & \new_[89596]_ ;
  assign \new_[89600]_  = A200 & ~A199;
  assign \new_[89603]_  = ~A203 & A201;
  assign \new_[89604]_  = \new_[89603]_  & \new_[89600]_ ;
  assign \new_[89605]_  = \new_[89604]_  & \new_[89597]_ ;
  assign \new_[89608]_  = ~A266 & A265;
  assign \new_[89611]_  = A268 & A267;
  assign \new_[89612]_  = \new_[89611]_  & \new_[89608]_ ;
  assign \new_[89615]_  = A299 & ~A298;
  assign \new_[89618]_  = ~A302 & A300;
  assign \new_[89619]_  = \new_[89618]_  & \new_[89615]_ ;
  assign \new_[89620]_  = \new_[89619]_  & \new_[89612]_ ;
  assign \new_[89624]_  = A168 & ~A169;
  assign \new_[89625]_  = ~A170 & \new_[89624]_ ;
  assign \new_[89628]_  = A200 & ~A199;
  assign \new_[89631]_  = ~A203 & A201;
  assign \new_[89632]_  = \new_[89631]_  & \new_[89628]_ ;
  assign \new_[89633]_  = \new_[89632]_  & \new_[89625]_ ;
  assign \new_[89636]_  = ~A266 & A265;
  assign \new_[89639]_  = ~A269 & A267;
  assign \new_[89640]_  = \new_[89639]_  & \new_[89636]_ ;
  assign \new_[89643]_  = ~A299 & A298;
  assign \new_[89646]_  = A301 & A300;
  assign \new_[89647]_  = \new_[89646]_  & \new_[89643]_ ;
  assign \new_[89648]_  = \new_[89647]_  & \new_[89640]_ ;
  assign \new_[89652]_  = A168 & ~A169;
  assign \new_[89653]_  = ~A170 & \new_[89652]_ ;
  assign \new_[89656]_  = A200 & ~A199;
  assign \new_[89659]_  = ~A203 & A201;
  assign \new_[89660]_  = \new_[89659]_  & \new_[89656]_ ;
  assign \new_[89661]_  = \new_[89660]_  & \new_[89653]_ ;
  assign \new_[89664]_  = ~A266 & A265;
  assign \new_[89667]_  = ~A269 & A267;
  assign \new_[89668]_  = \new_[89667]_  & \new_[89664]_ ;
  assign \new_[89671]_  = ~A299 & A298;
  assign \new_[89674]_  = ~A302 & A300;
  assign \new_[89675]_  = \new_[89674]_  & \new_[89671]_ ;
  assign \new_[89676]_  = \new_[89675]_  & \new_[89668]_ ;
  assign \new_[89680]_  = A168 & ~A169;
  assign \new_[89681]_  = ~A170 & \new_[89680]_ ;
  assign \new_[89684]_  = A200 & ~A199;
  assign \new_[89687]_  = ~A203 & A201;
  assign \new_[89688]_  = \new_[89687]_  & \new_[89684]_ ;
  assign \new_[89689]_  = \new_[89688]_  & \new_[89681]_ ;
  assign \new_[89692]_  = ~A266 & A265;
  assign \new_[89695]_  = ~A269 & A267;
  assign \new_[89696]_  = \new_[89695]_  & \new_[89692]_ ;
  assign \new_[89699]_  = A299 & ~A298;
  assign \new_[89702]_  = A301 & A300;
  assign \new_[89703]_  = \new_[89702]_  & \new_[89699]_ ;
  assign \new_[89704]_  = \new_[89703]_  & \new_[89696]_ ;
  assign \new_[89708]_  = A168 & ~A169;
  assign \new_[89709]_  = ~A170 & \new_[89708]_ ;
  assign \new_[89712]_  = A200 & ~A199;
  assign \new_[89715]_  = ~A203 & A201;
  assign \new_[89716]_  = \new_[89715]_  & \new_[89712]_ ;
  assign \new_[89717]_  = \new_[89716]_  & \new_[89709]_ ;
  assign \new_[89720]_  = ~A266 & A265;
  assign \new_[89723]_  = ~A269 & A267;
  assign \new_[89724]_  = \new_[89723]_  & \new_[89720]_ ;
  assign \new_[89727]_  = A299 & ~A298;
  assign \new_[89730]_  = ~A302 & A300;
  assign \new_[89731]_  = \new_[89730]_  & \new_[89727]_ ;
  assign \new_[89732]_  = \new_[89731]_  & \new_[89724]_ ;
  assign \new_[89736]_  = A168 & ~A169;
  assign \new_[89737]_  = ~A170 & \new_[89736]_ ;
  assign \new_[89740]_  = ~A200 & A199;
  assign \new_[89743]_  = A202 & A201;
  assign \new_[89744]_  = \new_[89743]_  & \new_[89740]_ ;
  assign \new_[89745]_  = \new_[89744]_  & \new_[89737]_ ;
  assign \new_[89748]_  = A266 & ~A265;
  assign \new_[89751]_  = A268 & A267;
  assign \new_[89752]_  = \new_[89751]_  & \new_[89748]_ ;
  assign \new_[89755]_  = ~A299 & A298;
  assign \new_[89758]_  = A301 & A300;
  assign \new_[89759]_  = \new_[89758]_  & \new_[89755]_ ;
  assign \new_[89760]_  = \new_[89759]_  & \new_[89752]_ ;
  assign \new_[89764]_  = A168 & ~A169;
  assign \new_[89765]_  = ~A170 & \new_[89764]_ ;
  assign \new_[89768]_  = ~A200 & A199;
  assign \new_[89771]_  = A202 & A201;
  assign \new_[89772]_  = \new_[89771]_  & \new_[89768]_ ;
  assign \new_[89773]_  = \new_[89772]_  & \new_[89765]_ ;
  assign \new_[89776]_  = A266 & ~A265;
  assign \new_[89779]_  = A268 & A267;
  assign \new_[89780]_  = \new_[89779]_  & \new_[89776]_ ;
  assign \new_[89783]_  = ~A299 & A298;
  assign \new_[89786]_  = ~A302 & A300;
  assign \new_[89787]_  = \new_[89786]_  & \new_[89783]_ ;
  assign \new_[89788]_  = \new_[89787]_  & \new_[89780]_ ;
  assign \new_[89792]_  = A168 & ~A169;
  assign \new_[89793]_  = ~A170 & \new_[89792]_ ;
  assign \new_[89796]_  = ~A200 & A199;
  assign \new_[89799]_  = A202 & A201;
  assign \new_[89800]_  = \new_[89799]_  & \new_[89796]_ ;
  assign \new_[89801]_  = \new_[89800]_  & \new_[89793]_ ;
  assign \new_[89804]_  = A266 & ~A265;
  assign \new_[89807]_  = A268 & A267;
  assign \new_[89808]_  = \new_[89807]_  & \new_[89804]_ ;
  assign \new_[89811]_  = A299 & ~A298;
  assign \new_[89814]_  = A301 & A300;
  assign \new_[89815]_  = \new_[89814]_  & \new_[89811]_ ;
  assign \new_[89816]_  = \new_[89815]_  & \new_[89808]_ ;
  assign \new_[89820]_  = A168 & ~A169;
  assign \new_[89821]_  = ~A170 & \new_[89820]_ ;
  assign \new_[89824]_  = ~A200 & A199;
  assign \new_[89827]_  = A202 & A201;
  assign \new_[89828]_  = \new_[89827]_  & \new_[89824]_ ;
  assign \new_[89829]_  = \new_[89828]_  & \new_[89821]_ ;
  assign \new_[89832]_  = A266 & ~A265;
  assign \new_[89835]_  = A268 & A267;
  assign \new_[89836]_  = \new_[89835]_  & \new_[89832]_ ;
  assign \new_[89839]_  = A299 & ~A298;
  assign \new_[89842]_  = ~A302 & A300;
  assign \new_[89843]_  = \new_[89842]_  & \new_[89839]_ ;
  assign \new_[89844]_  = \new_[89843]_  & \new_[89836]_ ;
  assign \new_[89848]_  = A168 & ~A169;
  assign \new_[89849]_  = ~A170 & \new_[89848]_ ;
  assign \new_[89852]_  = ~A200 & A199;
  assign \new_[89855]_  = A202 & A201;
  assign \new_[89856]_  = \new_[89855]_  & \new_[89852]_ ;
  assign \new_[89857]_  = \new_[89856]_  & \new_[89849]_ ;
  assign \new_[89860]_  = A266 & ~A265;
  assign \new_[89863]_  = ~A269 & A267;
  assign \new_[89864]_  = \new_[89863]_  & \new_[89860]_ ;
  assign \new_[89867]_  = ~A299 & A298;
  assign \new_[89870]_  = A301 & A300;
  assign \new_[89871]_  = \new_[89870]_  & \new_[89867]_ ;
  assign \new_[89872]_  = \new_[89871]_  & \new_[89864]_ ;
  assign \new_[89876]_  = A168 & ~A169;
  assign \new_[89877]_  = ~A170 & \new_[89876]_ ;
  assign \new_[89880]_  = ~A200 & A199;
  assign \new_[89883]_  = A202 & A201;
  assign \new_[89884]_  = \new_[89883]_  & \new_[89880]_ ;
  assign \new_[89885]_  = \new_[89884]_  & \new_[89877]_ ;
  assign \new_[89888]_  = A266 & ~A265;
  assign \new_[89891]_  = ~A269 & A267;
  assign \new_[89892]_  = \new_[89891]_  & \new_[89888]_ ;
  assign \new_[89895]_  = ~A299 & A298;
  assign \new_[89898]_  = ~A302 & A300;
  assign \new_[89899]_  = \new_[89898]_  & \new_[89895]_ ;
  assign \new_[89900]_  = \new_[89899]_  & \new_[89892]_ ;
  assign \new_[89904]_  = A168 & ~A169;
  assign \new_[89905]_  = ~A170 & \new_[89904]_ ;
  assign \new_[89908]_  = ~A200 & A199;
  assign \new_[89911]_  = A202 & A201;
  assign \new_[89912]_  = \new_[89911]_  & \new_[89908]_ ;
  assign \new_[89913]_  = \new_[89912]_  & \new_[89905]_ ;
  assign \new_[89916]_  = A266 & ~A265;
  assign \new_[89919]_  = ~A269 & A267;
  assign \new_[89920]_  = \new_[89919]_  & \new_[89916]_ ;
  assign \new_[89923]_  = A299 & ~A298;
  assign \new_[89926]_  = A301 & A300;
  assign \new_[89927]_  = \new_[89926]_  & \new_[89923]_ ;
  assign \new_[89928]_  = \new_[89927]_  & \new_[89920]_ ;
  assign \new_[89932]_  = A168 & ~A169;
  assign \new_[89933]_  = ~A170 & \new_[89932]_ ;
  assign \new_[89936]_  = ~A200 & A199;
  assign \new_[89939]_  = A202 & A201;
  assign \new_[89940]_  = \new_[89939]_  & \new_[89936]_ ;
  assign \new_[89941]_  = \new_[89940]_  & \new_[89933]_ ;
  assign \new_[89944]_  = A266 & ~A265;
  assign \new_[89947]_  = ~A269 & A267;
  assign \new_[89948]_  = \new_[89947]_  & \new_[89944]_ ;
  assign \new_[89951]_  = A299 & ~A298;
  assign \new_[89954]_  = ~A302 & A300;
  assign \new_[89955]_  = \new_[89954]_  & \new_[89951]_ ;
  assign \new_[89956]_  = \new_[89955]_  & \new_[89948]_ ;
  assign \new_[89960]_  = A168 & ~A169;
  assign \new_[89961]_  = ~A170 & \new_[89960]_ ;
  assign \new_[89964]_  = ~A200 & A199;
  assign \new_[89967]_  = A202 & A201;
  assign \new_[89968]_  = \new_[89967]_  & \new_[89964]_ ;
  assign \new_[89969]_  = \new_[89968]_  & \new_[89961]_ ;
  assign \new_[89972]_  = ~A266 & A265;
  assign \new_[89975]_  = A268 & A267;
  assign \new_[89976]_  = \new_[89975]_  & \new_[89972]_ ;
  assign \new_[89979]_  = ~A299 & A298;
  assign \new_[89982]_  = A301 & A300;
  assign \new_[89983]_  = \new_[89982]_  & \new_[89979]_ ;
  assign \new_[89984]_  = \new_[89983]_  & \new_[89976]_ ;
  assign \new_[89988]_  = A168 & ~A169;
  assign \new_[89989]_  = ~A170 & \new_[89988]_ ;
  assign \new_[89992]_  = ~A200 & A199;
  assign \new_[89995]_  = A202 & A201;
  assign \new_[89996]_  = \new_[89995]_  & \new_[89992]_ ;
  assign \new_[89997]_  = \new_[89996]_  & \new_[89989]_ ;
  assign \new_[90000]_  = ~A266 & A265;
  assign \new_[90003]_  = A268 & A267;
  assign \new_[90004]_  = \new_[90003]_  & \new_[90000]_ ;
  assign \new_[90007]_  = ~A299 & A298;
  assign \new_[90010]_  = ~A302 & A300;
  assign \new_[90011]_  = \new_[90010]_  & \new_[90007]_ ;
  assign \new_[90012]_  = \new_[90011]_  & \new_[90004]_ ;
  assign \new_[90016]_  = A168 & ~A169;
  assign \new_[90017]_  = ~A170 & \new_[90016]_ ;
  assign \new_[90020]_  = ~A200 & A199;
  assign \new_[90023]_  = A202 & A201;
  assign \new_[90024]_  = \new_[90023]_  & \new_[90020]_ ;
  assign \new_[90025]_  = \new_[90024]_  & \new_[90017]_ ;
  assign \new_[90028]_  = ~A266 & A265;
  assign \new_[90031]_  = A268 & A267;
  assign \new_[90032]_  = \new_[90031]_  & \new_[90028]_ ;
  assign \new_[90035]_  = A299 & ~A298;
  assign \new_[90038]_  = A301 & A300;
  assign \new_[90039]_  = \new_[90038]_  & \new_[90035]_ ;
  assign \new_[90040]_  = \new_[90039]_  & \new_[90032]_ ;
  assign \new_[90044]_  = A168 & ~A169;
  assign \new_[90045]_  = ~A170 & \new_[90044]_ ;
  assign \new_[90048]_  = ~A200 & A199;
  assign \new_[90051]_  = A202 & A201;
  assign \new_[90052]_  = \new_[90051]_  & \new_[90048]_ ;
  assign \new_[90053]_  = \new_[90052]_  & \new_[90045]_ ;
  assign \new_[90056]_  = ~A266 & A265;
  assign \new_[90059]_  = A268 & A267;
  assign \new_[90060]_  = \new_[90059]_  & \new_[90056]_ ;
  assign \new_[90063]_  = A299 & ~A298;
  assign \new_[90066]_  = ~A302 & A300;
  assign \new_[90067]_  = \new_[90066]_  & \new_[90063]_ ;
  assign \new_[90068]_  = \new_[90067]_  & \new_[90060]_ ;
  assign \new_[90072]_  = A168 & ~A169;
  assign \new_[90073]_  = ~A170 & \new_[90072]_ ;
  assign \new_[90076]_  = ~A200 & A199;
  assign \new_[90079]_  = A202 & A201;
  assign \new_[90080]_  = \new_[90079]_  & \new_[90076]_ ;
  assign \new_[90081]_  = \new_[90080]_  & \new_[90073]_ ;
  assign \new_[90084]_  = ~A266 & A265;
  assign \new_[90087]_  = ~A269 & A267;
  assign \new_[90088]_  = \new_[90087]_  & \new_[90084]_ ;
  assign \new_[90091]_  = ~A299 & A298;
  assign \new_[90094]_  = A301 & A300;
  assign \new_[90095]_  = \new_[90094]_  & \new_[90091]_ ;
  assign \new_[90096]_  = \new_[90095]_  & \new_[90088]_ ;
  assign \new_[90100]_  = A168 & ~A169;
  assign \new_[90101]_  = ~A170 & \new_[90100]_ ;
  assign \new_[90104]_  = ~A200 & A199;
  assign \new_[90107]_  = A202 & A201;
  assign \new_[90108]_  = \new_[90107]_  & \new_[90104]_ ;
  assign \new_[90109]_  = \new_[90108]_  & \new_[90101]_ ;
  assign \new_[90112]_  = ~A266 & A265;
  assign \new_[90115]_  = ~A269 & A267;
  assign \new_[90116]_  = \new_[90115]_  & \new_[90112]_ ;
  assign \new_[90119]_  = ~A299 & A298;
  assign \new_[90122]_  = ~A302 & A300;
  assign \new_[90123]_  = \new_[90122]_  & \new_[90119]_ ;
  assign \new_[90124]_  = \new_[90123]_  & \new_[90116]_ ;
  assign \new_[90128]_  = A168 & ~A169;
  assign \new_[90129]_  = ~A170 & \new_[90128]_ ;
  assign \new_[90132]_  = ~A200 & A199;
  assign \new_[90135]_  = A202 & A201;
  assign \new_[90136]_  = \new_[90135]_  & \new_[90132]_ ;
  assign \new_[90137]_  = \new_[90136]_  & \new_[90129]_ ;
  assign \new_[90140]_  = ~A266 & A265;
  assign \new_[90143]_  = ~A269 & A267;
  assign \new_[90144]_  = \new_[90143]_  & \new_[90140]_ ;
  assign \new_[90147]_  = A299 & ~A298;
  assign \new_[90150]_  = A301 & A300;
  assign \new_[90151]_  = \new_[90150]_  & \new_[90147]_ ;
  assign \new_[90152]_  = \new_[90151]_  & \new_[90144]_ ;
  assign \new_[90156]_  = A168 & ~A169;
  assign \new_[90157]_  = ~A170 & \new_[90156]_ ;
  assign \new_[90160]_  = ~A200 & A199;
  assign \new_[90163]_  = A202 & A201;
  assign \new_[90164]_  = \new_[90163]_  & \new_[90160]_ ;
  assign \new_[90165]_  = \new_[90164]_  & \new_[90157]_ ;
  assign \new_[90168]_  = ~A266 & A265;
  assign \new_[90171]_  = ~A269 & A267;
  assign \new_[90172]_  = \new_[90171]_  & \new_[90168]_ ;
  assign \new_[90175]_  = A299 & ~A298;
  assign \new_[90178]_  = ~A302 & A300;
  assign \new_[90179]_  = \new_[90178]_  & \new_[90175]_ ;
  assign \new_[90180]_  = \new_[90179]_  & \new_[90172]_ ;
  assign \new_[90184]_  = A168 & ~A169;
  assign \new_[90185]_  = ~A170 & \new_[90184]_ ;
  assign \new_[90188]_  = ~A200 & A199;
  assign \new_[90191]_  = ~A203 & A201;
  assign \new_[90192]_  = \new_[90191]_  & \new_[90188]_ ;
  assign \new_[90193]_  = \new_[90192]_  & \new_[90185]_ ;
  assign \new_[90196]_  = A266 & ~A265;
  assign \new_[90199]_  = A268 & A267;
  assign \new_[90200]_  = \new_[90199]_  & \new_[90196]_ ;
  assign \new_[90203]_  = ~A299 & A298;
  assign \new_[90206]_  = A301 & A300;
  assign \new_[90207]_  = \new_[90206]_  & \new_[90203]_ ;
  assign \new_[90208]_  = \new_[90207]_  & \new_[90200]_ ;
  assign \new_[90212]_  = A168 & ~A169;
  assign \new_[90213]_  = ~A170 & \new_[90212]_ ;
  assign \new_[90216]_  = ~A200 & A199;
  assign \new_[90219]_  = ~A203 & A201;
  assign \new_[90220]_  = \new_[90219]_  & \new_[90216]_ ;
  assign \new_[90221]_  = \new_[90220]_  & \new_[90213]_ ;
  assign \new_[90224]_  = A266 & ~A265;
  assign \new_[90227]_  = A268 & A267;
  assign \new_[90228]_  = \new_[90227]_  & \new_[90224]_ ;
  assign \new_[90231]_  = ~A299 & A298;
  assign \new_[90234]_  = ~A302 & A300;
  assign \new_[90235]_  = \new_[90234]_  & \new_[90231]_ ;
  assign \new_[90236]_  = \new_[90235]_  & \new_[90228]_ ;
  assign \new_[90240]_  = A168 & ~A169;
  assign \new_[90241]_  = ~A170 & \new_[90240]_ ;
  assign \new_[90244]_  = ~A200 & A199;
  assign \new_[90247]_  = ~A203 & A201;
  assign \new_[90248]_  = \new_[90247]_  & \new_[90244]_ ;
  assign \new_[90249]_  = \new_[90248]_  & \new_[90241]_ ;
  assign \new_[90252]_  = A266 & ~A265;
  assign \new_[90255]_  = A268 & A267;
  assign \new_[90256]_  = \new_[90255]_  & \new_[90252]_ ;
  assign \new_[90259]_  = A299 & ~A298;
  assign \new_[90262]_  = A301 & A300;
  assign \new_[90263]_  = \new_[90262]_  & \new_[90259]_ ;
  assign \new_[90264]_  = \new_[90263]_  & \new_[90256]_ ;
  assign \new_[90268]_  = A168 & ~A169;
  assign \new_[90269]_  = ~A170 & \new_[90268]_ ;
  assign \new_[90272]_  = ~A200 & A199;
  assign \new_[90275]_  = ~A203 & A201;
  assign \new_[90276]_  = \new_[90275]_  & \new_[90272]_ ;
  assign \new_[90277]_  = \new_[90276]_  & \new_[90269]_ ;
  assign \new_[90280]_  = A266 & ~A265;
  assign \new_[90283]_  = A268 & A267;
  assign \new_[90284]_  = \new_[90283]_  & \new_[90280]_ ;
  assign \new_[90287]_  = A299 & ~A298;
  assign \new_[90290]_  = ~A302 & A300;
  assign \new_[90291]_  = \new_[90290]_  & \new_[90287]_ ;
  assign \new_[90292]_  = \new_[90291]_  & \new_[90284]_ ;
  assign \new_[90296]_  = A168 & ~A169;
  assign \new_[90297]_  = ~A170 & \new_[90296]_ ;
  assign \new_[90300]_  = ~A200 & A199;
  assign \new_[90303]_  = ~A203 & A201;
  assign \new_[90304]_  = \new_[90303]_  & \new_[90300]_ ;
  assign \new_[90305]_  = \new_[90304]_  & \new_[90297]_ ;
  assign \new_[90308]_  = A266 & ~A265;
  assign \new_[90311]_  = ~A269 & A267;
  assign \new_[90312]_  = \new_[90311]_  & \new_[90308]_ ;
  assign \new_[90315]_  = ~A299 & A298;
  assign \new_[90318]_  = A301 & A300;
  assign \new_[90319]_  = \new_[90318]_  & \new_[90315]_ ;
  assign \new_[90320]_  = \new_[90319]_  & \new_[90312]_ ;
  assign \new_[90324]_  = A168 & ~A169;
  assign \new_[90325]_  = ~A170 & \new_[90324]_ ;
  assign \new_[90328]_  = ~A200 & A199;
  assign \new_[90331]_  = ~A203 & A201;
  assign \new_[90332]_  = \new_[90331]_  & \new_[90328]_ ;
  assign \new_[90333]_  = \new_[90332]_  & \new_[90325]_ ;
  assign \new_[90336]_  = A266 & ~A265;
  assign \new_[90339]_  = ~A269 & A267;
  assign \new_[90340]_  = \new_[90339]_  & \new_[90336]_ ;
  assign \new_[90343]_  = ~A299 & A298;
  assign \new_[90346]_  = ~A302 & A300;
  assign \new_[90347]_  = \new_[90346]_  & \new_[90343]_ ;
  assign \new_[90348]_  = \new_[90347]_  & \new_[90340]_ ;
  assign \new_[90352]_  = A168 & ~A169;
  assign \new_[90353]_  = ~A170 & \new_[90352]_ ;
  assign \new_[90356]_  = ~A200 & A199;
  assign \new_[90359]_  = ~A203 & A201;
  assign \new_[90360]_  = \new_[90359]_  & \new_[90356]_ ;
  assign \new_[90361]_  = \new_[90360]_  & \new_[90353]_ ;
  assign \new_[90364]_  = A266 & ~A265;
  assign \new_[90367]_  = ~A269 & A267;
  assign \new_[90368]_  = \new_[90367]_  & \new_[90364]_ ;
  assign \new_[90371]_  = A299 & ~A298;
  assign \new_[90374]_  = A301 & A300;
  assign \new_[90375]_  = \new_[90374]_  & \new_[90371]_ ;
  assign \new_[90376]_  = \new_[90375]_  & \new_[90368]_ ;
  assign \new_[90380]_  = A168 & ~A169;
  assign \new_[90381]_  = ~A170 & \new_[90380]_ ;
  assign \new_[90384]_  = ~A200 & A199;
  assign \new_[90387]_  = ~A203 & A201;
  assign \new_[90388]_  = \new_[90387]_  & \new_[90384]_ ;
  assign \new_[90389]_  = \new_[90388]_  & \new_[90381]_ ;
  assign \new_[90392]_  = A266 & ~A265;
  assign \new_[90395]_  = ~A269 & A267;
  assign \new_[90396]_  = \new_[90395]_  & \new_[90392]_ ;
  assign \new_[90399]_  = A299 & ~A298;
  assign \new_[90402]_  = ~A302 & A300;
  assign \new_[90403]_  = \new_[90402]_  & \new_[90399]_ ;
  assign \new_[90404]_  = \new_[90403]_  & \new_[90396]_ ;
  assign \new_[90408]_  = A168 & ~A169;
  assign \new_[90409]_  = ~A170 & \new_[90408]_ ;
  assign \new_[90412]_  = ~A200 & A199;
  assign \new_[90415]_  = ~A203 & A201;
  assign \new_[90416]_  = \new_[90415]_  & \new_[90412]_ ;
  assign \new_[90417]_  = \new_[90416]_  & \new_[90409]_ ;
  assign \new_[90420]_  = ~A266 & A265;
  assign \new_[90423]_  = A268 & A267;
  assign \new_[90424]_  = \new_[90423]_  & \new_[90420]_ ;
  assign \new_[90427]_  = ~A299 & A298;
  assign \new_[90430]_  = A301 & A300;
  assign \new_[90431]_  = \new_[90430]_  & \new_[90427]_ ;
  assign \new_[90432]_  = \new_[90431]_  & \new_[90424]_ ;
  assign \new_[90436]_  = A168 & ~A169;
  assign \new_[90437]_  = ~A170 & \new_[90436]_ ;
  assign \new_[90440]_  = ~A200 & A199;
  assign \new_[90443]_  = ~A203 & A201;
  assign \new_[90444]_  = \new_[90443]_  & \new_[90440]_ ;
  assign \new_[90445]_  = \new_[90444]_  & \new_[90437]_ ;
  assign \new_[90448]_  = ~A266 & A265;
  assign \new_[90451]_  = A268 & A267;
  assign \new_[90452]_  = \new_[90451]_  & \new_[90448]_ ;
  assign \new_[90455]_  = ~A299 & A298;
  assign \new_[90458]_  = ~A302 & A300;
  assign \new_[90459]_  = \new_[90458]_  & \new_[90455]_ ;
  assign \new_[90460]_  = \new_[90459]_  & \new_[90452]_ ;
  assign \new_[90464]_  = A168 & ~A169;
  assign \new_[90465]_  = ~A170 & \new_[90464]_ ;
  assign \new_[90468]_  = ~A200 & A199;
  assign \new_[90471]_  = ~A203 & A201;
  assign \new_[90472]_  = \new_[90471]_  & \new_[90468]_ ;
  assign \new_[90473]_  = \new_[90472]_  & \new_[90465]_ ;
  assign \new_[90476]_  = ~A266 & A265;
  assign \new_[90479]_  = A268 & A267;
  assign \new_[90480]_  = \new_[90479]_  & \new_[90476]_ ;
  assign \new_[90483]_  = A299 & ~A298;
  assign \new_[90486]_  = A301 & A300;
  assign \new_[90487]_  = \new_[90486]_  & \new_[90483]_ ;
  assign \new_[90488]_  = \new_[90487]_  & \new_[90480]_ ;
  assign \new_[90492]_  = A168 & ~A169;
  assign \new_[90493]_  = ~A170 & \new_[90492]_ ;
  assign \new_[90496]_  = ~A200 & A199;
  assign \new_[90499]_  = ~A203 & A201;
  assign \new_[90500]_  = \new_[90499]_  & \new_[90496]_ ;
  assign \new_[90501]_  = \new_[90500]_  & \new_[90493]_ ;
  assign \new_[90504]_  = ~A266 & A265;
  assign \new_[90507]_  = A268 & A267;
  assign \new_[90508]_  = \new_[90507]_  & \new_[90504]_ ;
  assign \new_[90511]_  = A299 & ~A298;
  assign \new_[90514]_  = ~A302 & A300;
  assign \new_[90515]_  = \new_[90514]_  & \new_[90511]_ ;
  assign \new_[90516]_  = \new_[90515]_  & \new_[90508]_ ;
  assign \new_[90520]_  = A168 & ~A169;
  assign \new_[90521]_  = ~A170 & \new_[90520]_ ;
  assign \new_[90524]_  = ~A200 & A199;
  assign \new_[90527]_  = ~A203 & A201;
  assign \new_[90528]_  = \new_[90527]_  & \new_[90524]_ ;
  assign \new_[90529]_  = \new_[90528]_  & \new_[90521]_ ;
  assign \new_[90532]_  = ~A266 & A265;
  assign \new_[90535]_  = ~A269 & A267;
  assign \new_[90536]_  = \new_[90535]_  & \new_[90532]_ ;
  assign \new_[90539]_  = ~A299 & A298;
  assign \new_[90542]_  = A301 & A300;
  assign \new_[90543]_  = \new_[90542]_  & \new_[90539]_ ;
  assign \new_[90544]_  = \new_[90543]_  & \new_[90536]_ ;
  assign \new_[90548]_  = A168 & ~A169;
  assign \new_[90549]_  = ~A170 & \new_[90548]_ ;
  assign \new_[90552]_  = ~A200 & A199;
  assign \new_[90555]_  = ~A203 & A201;
  assign \new_[90556]_  = \new_[90555]_  & \new_[90552]_ ;
  assign \new_[90557]_  = \new_[90556]_  & \new_[90549]_ ;
  assign \new_[90560]_  = ~A266 & A265;
  assign \new_[90563]_  = ~A269 & A267;
  assign \new_[90564]_  = \new_[90563]_  & \new_[90560]_ ;
  assign \new_[90567]_  = ~A299 & A298;
  assign \new_[90570]_  = ~A302 & A300;
  assign \new_[90571]_  = \new_[90570]_  & \new_[90567]_ ;
  assign \new_[90572]_  = \new_[90571]_  & \new_[90564]_ ;
  assign \new_[90576]_  = A168 & ~A169;
  assign \new_[90577]_  = ~A170 & \new_[90576]_ ;
  assign \new_[90580]_  = ~A200 & A199;
  assign \new_[90583]_  = ~A203 & A201;
  assign \new_[90584]_  = \new_[90583]_  & \new_[90580]_ ;
  assign \new_[90585]_  = \new_[90584]_  & \new_[90577]_ ;
  assign \new_[90588]_  = ~A266 & A265;
  assign \new_[90591]_  = ~A269 & A267;
  assign \new_[90592]_  = \new_[90591]_  & \new_[90588]_ ;
  assign \new_[90595]_  = A299 & ~A298;
  assign \new_[90598]_  = A301 & A300;
  assign \new_[90599]_  = \new_[90598]_  & \new_[90595]_ ;
  assign \new_[90600]_  = \new_[90599]_  & \new_[90592]_ ;
  assign \new_[90604]_  = A168 & ~A169;
  assign \new_[90605]_  = ~A170 & \new_[90604]_ ;
  assign \new_[90608]_  = ~A200 & A199;
  assign \new_[90611]_  = ~A203 & A201;
  assign \new_[90612]_  = \new_[90611]_  & \new_[90608]_ ;
  assign \new_[90613]_  = \new_[90612]_  & \new_[90605]_ ;
  assign \new_[90616]_  = ~A266 & A265;
  assign \new_[90619]_  = ~A269 & A267;
  assign \new_[90620]_  = \new_[90619]_  & \new_[90616]_ ;
  assign \new_[90623]_  = A299 & ~A298;
  assign \new_[90626]_  = ~A302 & A300;
  assign \new_[90627]_  = \new_[90626]_  & \new_[90623]_ ;
  assign \new_[90628]_  = \new_[90627]_  & \new_[90620]_ ;
  assign \new_[90632]_  = ~A168 & ~A169;
  assign \new_[90633]_  = ~A170 & \new_[90632]_ ;
  assign \new_[90636]_  = ~A166 & A167;
  assign \new_[90639]_  = ~A202 & A201;
  assign \new_[90640]_  = \new_[90639]_  & \new_[90636]_ ;
  assign \new_[90641]_  = \new_[90640]_  & \new_[90633]_ ;
  assign \new_[90644]_  = A267 & A203;
  assign \new_[90647]_  = A269 & ~A268;
  assign \new_[90648]_  = \new_[90647]_  & \new_[90644]_ ;
  assign \new_[90651]_  = ~A299 & A298;
  assign \new_[90654]_  = A301 & A300;
  assign \new_[90655]_  = \new_[90654]_  & \new_[90651]_ ;
  assign \new_[90656]_  = \new_[90655]_  & \new_[90648]_ ;
  assign \new_[90660]_  = ~A168 & ~A169;
  assign \new_[90661]_  = ~A170 & \new_[90660]_ ;
  assign \new_[90664]_  = ~A166 & A167;
  assign \new_[90667]_  = ~A202 & A201;
  assign \new_[90668]_  = \new_[90667]_  & \new_[90664]_ ;
  assign \new_[90669]_  = \new_[90668]_  & \new_[90661]_ ;
  assign \new_[90672]_  = A267 & A203;
  assign \new_[90675]_  = A269 & ~A268;
  assign \new_[90676]_  = \new_[90675]_  & \new_[90672]_ ;
  assign \new_[90679]_  = ~A299 & A298;
  assign \new_[90682]_  = ~A302 & A300;
  assign \new_[90683]_  = \new_[90682]_  & \new_[90679]_ ;
  assign \new_[90684]_  = \new_[90683]_  & \new_[90676]_ ;
  assign \new_[90688]_  = ~A168 & ~A169;
  assign \new_[90689]_  = ~A170 & \new_[90688]_ ;
  assign \new_[90692]_  = ~A166 & A167;
  assign \new_[90695]_  = ~A202 & A201;
  assign \new_[90696]_  = \new_[90695]_  & \new_[90692]_ ;
  assign \new_[90697]_  = \new_[90696]_  & \new_[90689]_ ;
  assign \new_[90700]_  = A267 & A203;
  assign \new_[90703]_  = A269 & ~A268;
  assign \new_[90704]_  = \new_[90703]_  & \new_[90700]_ ;
  assign \new_[90707]_  = A299 & ~A298;
  assign \new_[90710]_  = A301 & A300;
  assign \new_[90711]_  = \new_[90710]_  & \new_[90707]_ ;
  assign \new_[90712]_  = \new_[90711]_  & \new_[90704]_ ;
  assign \new_[90716]_  = ~A168 & ~A169;
  assign \new_[90717]_  = ~A170 & \new_[90716]_ ;
  assign \new_[90720]_  = ~A166 & A167;
  assign \new_[90723]_  = ~A202 & A201;
  assign \new_[90724]_  = \new_[90723]_  & \new_[90720]_ ;
  assign \new_[90725]_  = \new_[90724]_  & \new_[90717]_ ;
  assign \new_[90728]_  = A267 & A203;
  assign \new_[90731]_  = A269 & ~A268;
  assign \new_[90732]_  = \new_[90731]_  & \new_[90728]_ ;
  assign \new_[90735]_  = A299 & ~A298;
  assign \new_[90738]_  = ~A302 & A300;
  assign \new_[90739]_  = \new_[90738]_  & \new_[90735]_ ;
  assign \new_[90740]_  = \new_[90739]_  & \new_[90732]_ ;
  assign \new_[90744]_  = ~A168 & ~A169;
  assign \new_[90745]_  = ~A170 & \new_[90744]_ ;
  assign \new_[90748]_  = ~A166 & A167;
  assign \new_[90751]_  = ~A202 & A201;
  assign \new_[90752]_  = \new_[90751]_  & \new_[90748]_ ;
  assign \new_[90753]_  = \new_[90752]_  & \new_[90745]_ ;
  assign \new_[90756]_  = ~A267 & A203;
  assign \new_[90759]_  = A298 & A268;
  assign \new_[90760]_  = \new_[90759]_  & \new_[90756]_ ;
  assign \new_[90763]_  = ~A300 & ~A299;
  assign \new_[90766]_  = A302 & ~A301;
  assign \new_[90767]_  = \new_[90766]_  & \new_[90763]_ ;
  assign \new_[90768]_  = \new_[90767]_  & \new_[90760]_ ;
  assign \new_[90772]_  = ~A168 & ~A169;
  assign \new_[90773]_  = ~A170 & \new_[90772]_ ;
  assign \new_[90776]_  = ~A166 & A167;
  assign \new_[90779]_  = ~A202 & A201;
  assign \new_[90780]_  = \new_[90779]_  & \new_[90776]_ ;
  assign \new_[90781]_  = \new_[90780]_  & \new_[90773]_ ;
  assign \new_[90784]_  = ~A267 & A203;
  assign \new_[90787]_  = ~A298 & A268;
  assign \new_[90788]_  = \new_[90787]_  & \new_[90784]_ ;
  assign \new_[90791]_  = ~A300 & A299;
  assign \new_[90794]_  = A302 & ~A301;
  assign \new_[90795]_  = \new_[90794]_  & \new_[90791]_ ;
  assign \new_[90796]_  = \new_[90795]_  & \new_[90788]_ ;
  assign \new_[90800]_  = ~A168 & ~A169;
  assign \new_[90801]_  = ~A170 & \new_[90800]_ ;
  assign \new_[90804]_  = ~A166 & A167;
  assign \new_[90807]_  = ~A202 & A201;
  assign \new_[90808]_  = \new_[90807]_  & \new_[90804]_ ;
  assign \new_[90809]_  = \new_[90808]_  & \new_[90801]_ ;
  assign \new_[90812]_  = ~A267 & A203;
  assign \new_[90815]_  = A298 & ~A269;
  assign \new_[90816]_  = \new_[90815]_  & \new_[90812]_ ;
  assign \new_[90819]_  = ~A300 & ~A299;
  assign \new_[90822]_  = A302 & ~A301;
  assign \new_[90823]_  = \new_[90822]_  & \new_[90819]_ ;
  assign \new_[90824]_  = \new_[90823]_  & \new_[90816]_ ;
  assign \new_[90828]_  = ~A168 & ~A169;
  assign \new_[90829]_  = ~A170 & \new_[90828]_ ;
  assign \new_[90832]_  = ~A166 & A167;
  assign \new_[90835]_  = ~A202 & A201;
  assign \new_[90836]_  = \new_[90835]_  & \new_[90832]_ ;
  assign \new_[90837]_  = \new_[90836]_  & \new_[90829]_ ;
  assign \new_[90840]_  = ~A267 & A203;
  assign \new_[90843]_  = ~A298 & ~A269;
  assign \new_[90844]_  = \new_[90843]_  & \new_[90840]_ ;
  assign \new_[90847]_  = ~A300 & A299;
  assign \new_[90850]_  = A302 & ~A301;
  assign \new_[90851]_  = \new_[90850]_  & \new_[90847]_ ;
  assign \new_[90852]_  = \new_[90851]_  & \new_[90844]_ ;
  assign \new_[90856]_  = ~A168 & ~A169;
  assign \new_[90857]_  = ~A170 & \new_[90856]_ ;
  assign \new_[90860]_  = ~A166 & A167;
  assign \new_[90863]_  = ~A202 & A201;
  assign \new_[90864]_  = \new_[90863]_  & \new_[90860]_ ;
  assign \new_[90865]_  = \new_[90864]_  & \new_[90857]_ ;
  assign \new_[90868]_  = A265 & A203;
  assign \new_[90871]_  = A298 & A266;
  assign \new_[90872]_  = \new_[90871]_  & \new_[90868]_ ;
  assign \new_[90875]_  = ~A300 & ~A299;
  assign \new_[90878]_  = A302 & ~A301;
  assign \new_[90879]_  = \new_[90878]_  & \new_[90875]_ ;
  assign \new_[90880]_  = \new_[90879]_  & \new_[90872]_ ;
  assign \new_[90884]_  = ~A168 & ~A169;
  assign \new_[90885]_  = ~A170 & \new_[90884]_ ;
  assign \new_[90888]_  = ~A166 & A167;
  assign \new_[90891]_  = ~A202 & A201;
  assign \new_[90892]_  = \new_[90891]_  & \new_[90888]_ ;
  assign \new_[90893]_  = \new_[90892]_  & \new_[90885]_ ;
  assign \new_[90896]_  = A265 & A203;
  assign \new_[90899]_  = ~A298 & A266;
  assign \new_[90900]_  = \new_[90899]_  & \new_[90896]_ ;
  assign \new_[90903]_  = ~A300 & A299;
  assign \new_[90906]_  = A302 & ~A301;
  assign \new_[90907]_  = \new_[90906]_  & \new_[90903]_ ;
  assign \new_[90908]_  = \new_[90907]_  & \new_[90900]_ ;
  assign \new_[90912]_  = ~A168 & ~A169;
  assign \new_[90913]_  = ~A170 & \new_[90912]_ ;
  assign \new_[90916]_  = ~A166 & A167;
  assign \new_[90919]_  = ~A202 & A201;
  assign \new_[90920]_  = \new_[90919]_  & \new_[90916]_ ;
  assign \new_[90921]_  = \new_[90920]_  & \new_[90913]_ ;
  assign \new_[90924]_  = ~A265 & A203;
  assign \new_[90927]_  = A267 & A266;
  assign \new_[90928]_  = \new_[90927]_  & \new_[90924]_ ;
  assign \new_[90931]_  = A300 & A268;
  assign \new_[90934]_  = A302 & ~A301;
  assign \new_[90935]_  = \new_[90934]_  & \new_[90931]_ ;
  assign \new_[90936]_  = \new_[90935]_  & \new_[90928]_ ;
  assign \new_[90940]_  = ~A168 & ~A169;
  assign \new_[90941]_  = ~A170 & \new_[90940]_ ;
  assign \new_[90944]_  = ~A166 & A167;
  assign \new_[90947]_  = ~A202 & A201;
  assign \new_[90948]_  = \new_[90947]_  & \new_[90944]_ ;
  assign \new_[90949]_  = \new_[90948]_  & \new_[90941]_ ;
  assign \new_[90952]_  = ~A265 & A203;
  assign \new_[90955]_  = A267 & A266;
  assign \new_[90956]_  = \new_[90955]_  & \new_[90952]_ ;
  assign \new_[90959]_  = A300 & ~A269;
  assign \new_[90962]_  = A302 & ~A301;
  assign \new_[90963]_  = \new_[90962]_  & \new_[90959]_ ;
  assign \new_[90964]_  = \new_[90963]_  & \new_[90956]_ ;
  assign \new_[90968]_  = ~A168 & ~A169;
  assign \new_[90969]_  = ~A170 & \new_[90968]_ ;
  assign \new_[90972]_  = ~A166 & A167;
  assign \new_[90975]_  = ~A202 & A201;
  assign \new_[90976]_  = \new_[90975]_  & \new_[90972]_ ;
  assign \new_[90977]_  = \new_[90976]_  & \new_[90969]_ ;
  assign \new_[90980]_  = ~A265 & A203;
  assign \new_[90983]_  = ~A267 & A266;
  assign \new_[90984]_  = \new_[90983]_  & \new_[90980]_ ;
  assign \new_[90987]_  = A269 & ~A268;
  assign \new_[90990]_  = A301 & ~A300;
  assign \new_[90991]_  = \new_[90990]_  & \new_[90987]_ ;
  assign \new_[90992]_  = \new_[90991]_  & \new_[90984]_ ;
  assign \new_[90996]_  = ~A168 & ~A169;
  assign \new_[90997]_  = ~A170 & \new_[90996]_ ;
  assign \new_[91000]_  = ~A166 & A167;
  assign \new_[91003]_  = ~A202 & A201;
  assign \new_[91004]_  = \new_[91003]_  & \new_[91000]_ ;
  assign \new_[91005]_  = \new_[91004]_  & \new_[90997]_ ;
  assign \new_[91008]_  = ~A265 & A203;
  assign \new_[91011]_  = ~A267 & A266;
  assign \new_[91012]_  = \new_[91011]_  & \new_[91008]_ ;
  assign \new_[91015]_  = A269 & ~A268;
  assign \new_[91018]_  = ~A302 & ~A300;
  assign \new_[91019]_  = \new_[91018]_  & \new_[91015]_ ;
  assign \new_[91020]_  = \new_[91019]_  & \new_[91012]_ ;
  assign \new_[91024]_  = ~A168 & ~A169;
  assign \new_[91025]_  = ~A170 & \new_[91024]_ ;
  assign \new_[91028]_  = ~A166 & A167;
  assign \new_[91031]_  = ~A202 & A201;
  assign \new_[91032]_  = \new_[91031]_  & \new_[91028]_ ;
  assign \new_[91033]_  = \new_[91032]_  & \new_[91025]_ ;
  assign \new_[91036]_  = ~A265 & A203;
  assign \new_[91039]_  = ~A267 & A266;
  assign \new_[91040]_  = \new_[91039]_  & \new_[91036]_ ;
  assign \new_[91043]_  = A269 & ~A268;
  assign \new_[91046]_  = A299 & A298;
  assign \new_[91047]_  = \new_[91046]_  & \new_[91043]_ ;
  assign \new_[91048]_  = \new_[91047]_  & \new_[91040]_ ;
  assign \new_[91052]_  = ~A168 & ~A169;
  assign \new_[91053]_  = ~A170 & \new_[91052]_ ;
  assign \new_[91056]_  = ~A166 & A167;
  assign \new_[91059]_  = ~A202 & A201;
  assign \new_[91060]_  = \new_[91059]_  & \new_[91056]_ ;
  assign \new_[91061]_  = \new_[91060]_  & \new_[91053]_ ;
  assign \new_[91064]_  = ~A265 & A203;
  assign \new_[91067]_  = ~A267 & A266;
  assign \new_[91068]_  = \new_[91067]_  & \new_[91064]_ ;
  assign \new_[91071]_  = A269 & ~A268;
  assign \new_[91074]_  = ~A299 & ~A298;
  assign \new_[91075]_  = \new_[91074]_  & \new_[91071]_ ;
  assign \new_[91076]_  = \new_[91075]_  & \new_[91068]_ ;
  assign \new_[91080]_  = ~A168 & ~A169;
  assign \new_[91081]_  = ~A170 & \new_[91080]_ ;
  assign \new_[91084]_  = ~A166 & A167;
  assign \new_[91087]_  = ~A202 & A201;
  assign \new_[91088]_  = \new_[91087]_  & \new_[91084]_ ;
  assign \new_[91089]_  = \new_[91088]_  & \new_[91081]_ ;
  assign \new_[91092]_  = A265 & A203;
  assign \new_[91095]_  = A267 & ~A266;
  assign \new_[91096]_  = \new_[91095]_  & \new_[91092]_ ;
  assign \new_[91099]_  = A300 & A268;
  assign \new_[91102]_  = A302 & ~A301;
  assign \new_[91103]_  = \new_[91102]_  & \new_[91099]_ ;
  assign \new_[91104]_  = \new_[91103]_  & \new_[91096]_ ;
  assign \new_[91108]_  = ~A168 & ~A169;
  assign \new_[91109]_  = ~A170 & \new_[91108]_ ;
  assign \new_[91112]_  = ~A166 & A167;
  assign \new_[91115]_  = ~A202 & A201;
  assign \new_[91116]_  = \new_[91115]_  & \new_[91112]_ ;
  assign \new_[91117]_  = \new_[91116]_  & \new_[91109]_ ;
  assign \new_[91120]_  = A265 & A203;
  assign \new_[91123]_  = A267 & ~A266;
  assign \new_[91124]_  = \new_[91123]_  & \new_[91120]_ ;
  assign \new_[91127]_  = A300 & ~A269;
  assign \new_[91130]_  = A302 & ~A301;
  assign \new_[91131]_  = \new_[91130]_  & \new_[91127]_ ;
  assign \new_[91132]_  = \new_[91131]_  & \new_[91124]_ ;
  assign \new_[91136]_  = ~A168 & ~A169;
  assign \new_[91137]_  = ~A170 & \new_[91136]_ ;
  assign \new_[91140]_  = ~A166 & A167;
  assign \new_[91143]_  = ~A202 & A201;
  assign \new_[91144]_  = \new_[91143]_  & \new_[91140]_ ;
  assign \new_[91145]_  = \new_[91144]_  & \new_[91137]_ ;
  assign \new_[91148]_  = A265 & A203;
  assign \new_[91151]_  = ~A267 & ~A266;
  assign \new_[91152]_  = \new_[91151]_  & \new_[91148]_ ;
  assign \new_[91155]_  = A269 & ~A268;
  assign \new_[91158]_  = A301 & ~A300;
  assign \new_[91159]_  = \new_[91158]_  & \new_[91155]_ ;
  assign \new_[91160]_  = \new_[91159]_  & \new_[91152]_ ;
  assign \new_[91164]_  = ~A168 & ~A169;
  assign \new_[91165]_  = ~A170 & \new_[91164]_ ;
  assign \new_[91168]_  = ~A166 & A167;
  assign \new_[91171]_  = ~A202 & A201;
  assign \new_[91172]_  = \new_[91171]_  & \new_[91168]_ ;
  assign \new_[91173]_  = \new_[91172]_  & \new_[91165]_ ;
  assign \new_[91176]_  = A265 & A203;
  assign \new_[91179]_  = ~A267 & ~A266;
  assign \new_[91180]_  = \new_[91179]_  & \new_[91176]_ ;
  assign \new_[91183]_  = A269 & ~A268;
  assign \new_[91186]_  = ~A302 & ~A300;
  assign \new_[91187]_  = \new_[91186]_  & \new_[91183]_ ;
  assign \new_[91188]_  = \new_[91187]_  & \new_[91180]_ ;
  assign \new_[91192]_  = ~A168 & ~A169;
  assign \new_[91193]_  = ~A170 & \new_[91192]_ ;
  assign \new_[91196]_  = ~A166 & A167;
  assign \new_[91199]_  = ~A202 & A201;
  assign \new_[91200]_  = \new_[91199]_  & \new_[91196]_ ;
  assign \new_[91201]_  = \new_[91200]_  & \new_[91193]_ ;
  assign \new_[91204]_  = A265 & A203;
  assign \new_[91207]_  = ~A267 & ~A266;
  assign \new_[91208]_  = \new_[91207]_  & \new_[91204]_ ;
  assign \new_[91211]_  = A269 & ~A268;
  assign \new_[91214]_  = A299 & A298;
  assign \new_[91215]_  = \new_[91214]_  & \new_[91211]_ ;
  assign \new_[91216]_  = \new_[91215]_  & \new_[91208]_ ;
  assign \new_[91220]_  = ~A168 & ~A169;
  assign \new_[91221]_  = ~A170 & \new_[91220]_ ;
  assign \new_[91224]_  = ~A166 & A167;
  assign \new_[91227]_  = ~A202 & A201;
  assign \new_[91228]_  = \new_[91227]_  & \new_[91224]_ ;
  assign \new_[91229]_  = \new_[91228]_  & \new_[91221]_ ;
  assign \new_[91232]_  = A265 & A203;
  assign \new_[91235]_  = ~A267 & ~A266;
  assign \new_[91236]_  = \new_[91235]_  & \new_[91232]_ ;
  assign \new_[91239]_  = A269 & ~A268;
  assign \new_[91242]_  = ~A299 & ~A298;
  assign \new_[91243]_  = \new_[91242]_  & \new_[91239]_ ;
  assign \new_[91244]_  = \new_[91243]_  & \new_[91236]_ ;
  assign \new_[91248]_  = ~A168 & ~A169;
  assign \new_[91249]_  = ~A170 & \new_[91248]_ ;
  assign \new_[91252]_  = ~A166 & A167;
  assign \new_[91255]_  = ~A202 & A201;
  assign \new_[91256]_  = \new_[91255]_  & \new_[91252]_ ;
  assign \new_[91257]_  = \new_[91256]_  & \new_[91249]_ ;
  assign \new_[91260]_  = ~A265 & A203;
  assign \new_[91263]_  = A298 & ~A266;
  assign \new_[91264]_  = \new_[91263]_  & \new_[91260]_ ;
  assign \new_[91267]_  = ~A300 & ~A299;
  assign \new_[91270]_  = A302 & ~A301;
  assign \new_[91271]_  = \new_[91270]_  & \new_[91267]_ ;
  assign \new_[91272]_  = \new_[91271]_  & \new_[91264]_ ;
  assign \new_[91276]_  = ~A168 & ~A169;
  assign \new_[91277]_  = ~A170 & \new_[91276]_ ;
  assign \new_[91280]_  = ~A166 & A167;
  assign \new_[91283]_  = ~A202 & A201;
  assign \new_[91284]_  = \new_[91283]_  & \new_[91280]_ ;
  assign \new_[91285]_  = \new_[91284]_  & \new_[91277]_ ;
  assign \new_[91288]_  = ~A265 & A203;
  assign \new_[91291]_  = ~A298 & ~A266;
  assign \new_[91292]_  = \new_[91291]_  & \new_[91288]_ ;
  assign \new_[91295]_  = ~A300 & A299;
  assign \new_[91298]_  = A302 & ~A301;
  assign \new_[91299]_  = \new_[91298]_  & \new_[91295]_ ;
  assign \new_[91300]_  = \new_[91299]_  & \new_[91292]_ ;
  assign \new_[91304]_  = ~A168 & ~A169;
  assign \new_[91305]_  = ~A170 & \new_[91304]_ ;
  assign \new_[91308]_  = ~A166 & A167;
  assign \new_[91311]_  = A202 & ~A201;
  assign \new_[91312]_  = \new_[91311]_  & \new_[91308]_ ;
  assign \new_[91313]_  = \new_[91312]_  & \new_[91305]_ ;
  assign \new_[91316]_  = ~A268 & A267;
  assign \new_[91319]_  = A298 & A269;
  assign \new_[91320]_  = \new_[91319]_  & \new_[91316]_ ;
  assign \new_[91323]_  = ~A300 & ~A299;
  assign \new_[91326]_  = A302 & ~A301;
  assign \new_[91327]_  = \new_[91326]_  & \new_[91323]_ ;
  assign \new_[91328]_  = \new_[91327]_  & \new_[91320]_ ;
  assign \new_[91332]_  = ~A168 & ~A169;
  assign \new_[91333]_  = ~A170 & \new_[91332]_ ;
  assign \new_[91336]_  = ~A166 & A167;
  assign \new_[91339]_  = A202 & ~A201;
  assign \new_[91340]_  = \new_[91339]_  & \new_[91336]_ ;
  assign \new_[91341]_  = \new_[91340]_  & \new_[91333]_ ;
  assign \new_[91344]_  = ~A268 & A267;
  assign \new_[91347]_  = ~A298 & A269;
  assign \new_[91348]_  = \new_[91347]_  & \new_[91344]_ ;
  assign \new_[91351]_  = ~A300 & A299;
  assign \new_[91354]_  = A302 & ~A301;
  assign \new_[91355]_  = \new_[91354]_  & \new_[91351]_ ;
  assign \new_[91356]_  = \new_[91355]_  & \new_[91348]_ ;
  assign \new_[91360]_  = ~A168 & ~A169;
  assign \new_[91361]_  = ~A170 & \new_[91360]_ ;
  assign \new_[91364]_  = ~A166 & A167;
  assign \new_[91367]_  = A202 & ~A201;
  assign \new_[91368]_  = \new_[91367]_  & \new_[91364]_ ;
  assign \new_[91369]_  = \new_[91368]_  & \new_[91361]_ ;
  assign \new_[91372]_  = A266 & ~A265;
  assign \new_[91375]_  = ~A268 & ~A267;
  assign \new_[91376]_  = \new_[91375]_  & \new_[91372]_ ;
  assign \new_[91379]_  = A300 & A269;
  assign \new_[91382]_  = A302 & ~A301;
  assign \new_[91383]_  = \new_[91382]_  & \new_[91379]_ ;
  assign \new_[91384]_  = \new_[91383]_  & \new_[91376]_ ;
  assign \new_[91388]_  = ~A168 & ~A169;
  assign \new_[91389]_  = ~A170 & \new_[91388]_ ;
  assign \new_[91392]_  = ~A166 & A167;
  assign \new_[91395]_  = A202 & ~A201;
  assign \new_[91396]_  = \new_[91395]_  & \new_[91392]_ ;
  assign \new_[91397]_  = \new_[91396]_  & \new_[91389]_ ;
  assign \new_[91400]_  = ~A266 & A265;
  assign \new_[91403]_  = ~A268 & ~A267;
  assign \new_[91404]_  = \new_[91403]_  & \new_[91400]_ ;
  assign \new_[91407]_  = A300 & A269;
  assign \new_[91410]_  = A302 & ~A301;
  assign \new_[91411]_  = \new_[91410]_  & \new_[91407]_ ;
  assign \new_[91412]_  = \new_[91411]_  & \new_[91404]_ ;
  assign \new_[91416]_  = ~A168 & ~A169;
  assign \new_[91417]_  = ~A170 & \new_[91416]_ ;
  assign \new_[91420]_  = ~A166 & A167;
  assign \new_[91423]_  = ~A203 & ~A201;
  assign \new_[91424]_  = \new_[91423]_  & \new_[91420]_ ;
  assign \new_[91425]_  = \new_[91424]_  & \new_[91417]_ ;
  assign \new_[91428]_  = ~A268 & A267;
  assign \new_[91431]_  = A298 & A269;
  assign \new_[91432]_  = \new_[91431]_  & \new_[91428]_ ;
  assign \new_[91435]_  = ~A300 & ~A299;
  assign \new_[91438]_  = A302 & ~A301;
  assign \new_[91439]_  = \new_[91438]_  & \new_[91435]_ ;
  assign \new_[91440]_  = \new_[91439]_  & \new_[91432]_ ;
  assign \new_[91444]_  = ~A168 & ~A169;
  assign \new_[91445]_  = ~A170 & \new_[91444]_ ;
  assign \new_[91448]_  = ~A166 & A167;
  assign \new_[91451]_  = ~A203 & ~A201;
  assign \new_[91452]_  = \new_[91451]_  & \new_[91448]_ ;
  assign \new_[91453]_  = \new_[91452]_  & \new_[91445]_ ;
  assign \new_[91456]_  = ~A268 & A267;
  assign \new_[91459]_  = ~A298 & A269;
  assign \new_[91460]_  = \new_[91459]_  & \new_[91456]_ ;
  assign \new_[91463]_  = ~A300 & A299;
  assign \new_[91466]_  = A302 & ~A301;
  assign \new_[91467]_  = \new_[91466]_  & \new_[91463]_ ;
  assign \new_[91468]_  = \new_[91467]_  & \new_[91460]_ ;
  assign \new_[91472]_  = ~A168 & ~A169;
  assign \new_[91473]_  = ~A170 & \new_[91472]_ ;
  assign \new_[91476]_  = ~A166 & A167;
  assign \new_[91479]_  = ~A203 & ~A201;
  assign \new_[91480]_  = \new_[91479]_  & \new_[91476]_ ;
  assign \new_[91481]_  = \new_[91480]_  & \new_[91473]_ ;
  assign \new_[91484]_  = A266 & ~A265;
  assign \new_[91487]_  = ~A268 & ~A267;
  assign \new_[91488]_  = \new_[91487]_  & \new_[91484]_ ;
  assign \new_[91491]_  = A300 & A269;
  assign \new_[91494]_  = A302 & ~A301;
  assign \new_[91495]_  = \new_[91494]_  & \new_[91491]_ ;
  assign \new_[91496]_  = \new_[91495]_  & \new_[91488]_ ;
  assign \new_[91500]_  = ~A168 & ~A169;
  assign \new_[91501]_  = ~A170 & \new_[91500]_ ;
  assign \new_[91504]_  = ~A166 & A167;
  assign \new_[91507]_  = ~A203 & ~A201;
  assign \new_[91508]_  = \new_[91507]_  & \new_[91504]_ ;
  assign \new_[91509]_  = \new_[91508]_  & \new_[91501]_ ;
  assign \new_[91512]_  = ~A266 & A265;
  assign \new_[91515]_  = ~A268 & ~A267;
  assign \new_[91516]_  = \new_[91515]_  & \new_[91512]_ ;
  assign \new_[91519]_  = A300 & A269;
  assign \new_[91522]_  = A302 & ~A301;
  assign \new_[91523]_  = \new_[91522]_  & \new_[91519]_ ;
  assign \new_[91524]_  = \new_[91523]_  & \new_[91516]_ ;
  assign \new_[91528]_  = ~A168 & ~A169;
  assign \new_[91529]_  = ~A170 & \new_[91528]_ ;
  assign \new_[91532]_  = ~A166 & A167;
  assign \new_[91535]_  = A200 & A199;
  assign \new_[91536]_  = \new_[91535]_  & \new_[91532]_ ;
  assign \new_[91537]_  = \new_[91536]_  & \new_[91529]_ ;
  assign \new_[91540]_  = ~A268 & A267;
  assign \new_[91543]_  = A298 & A269;
  assign \new_[91544]_  = \new_[91543]_  & \new_[91540]_ ;
  assign \new_[91547]_  = ~A300 & ~A299;
  assign \new_[91550]_  = A302 & ~A301;
  assign \new_[91551]_  = \new_[91550]_  & \new_[91547]_ ;
  assign \new_[91552]_  = \new_[91551]_  & \new_[91544]_ ;
  assign \new_[91556]_  = ~A168 & ~A169;
  assign \new_[91557]_  = ~A170 & \new_[91556]_ ;
  assign \new_[91560]_  = ~A166 & A167;
  assign \new_[91563]_  = A200 & A199;
  assign \new_[91564]_  = \new_[91563]_  & \new_[91560]_ ;
  assign \new_[91565]_  = \new_[91564]_  & \new_[91557]_ ;
  assign \new_[91568]_  = ~A268 & A267;
  assign \new_[91571]_  = ~A298 & A269;
  assign \new_[91572]_  = \new_[91571]_  & \new_[91568]_ ;
  assign \new_[91575]_  = ~A300 & A299;
  assign \new_[91578]_  = A302 & ~A301;
  assign \new_[91579]_  = \new_[91578]_  & \new_[91575]_ ;
  assign \new_[91580]_  = \new_[91579]_  & \new_[91572]_ ;
  assign \new_[91584]_  = ~A168 & ~A169;
  assign \new_[91585]_  = ~A170 & \new_[91584]_ ;
  assign \new_[91588]_  = ~A166 & A167;
  assign \new_[91591]_  = A200 & A199;
  assign \new_[91592]_  = \new_[91591]_  & \new_[91588]_ ;
  assign \new_[91593]_  = \new_[91592]_  & \new_[91585]_ ;
  assign \new_[91596]_  = A266 & ~A265;
  assign \new_[91599]_  = ~A268 & ~A267;
  assign \new_[91600]_  = \new_[91599]_  & \new_[91596]_ ;
  assign \new_[91603]_  = A300 & A269;
  assign \new_[91606]_  = A302 & ~A301;
  assign \new_[91607]_  = \new_[91606]_  & \new_[91603]_ ;
  assign \new_[91608]_  = \new_[91607]_  & \new_[91600]_ ;
  assign \new_[91612]_  = ~A168 & ~A169;
  assign \new_[91613]_  = ~A170 & \new_[91612]_ ;
  assign \new_[91616]_  = ~A166 & A167;
  assign \new_[91619]_  = A200 & A199;
  assign \new_[91620]_  = \new_[91619]_  & \new_[91616]_ ;
  assign \new_[91621]_  = \new_[91620]_  & \new_[91613]_ ;
  assign \new_[91624]_  = ~A266 & A265;
  assign \new_[91627]_  = ~A268 & ~A267;
  assign \new_[91628]_  = \new_[91627]_  & \new_[91624]_ ;
  assign \new_[91631]_  = A300 & A269;
  assign \new_[91634]_  = A302 & ~A301;
  assign \new_[91635]_  = \new_[91634]_  & \new_[91631]_ ;
  assign \new_[91636]_  = \new_[91635]_  & \new_[91628]_ ;
  assign \new_[91640]_  = ~A168 & ~A169;
  assign \new_[91641]_  = ~A170 & \new_[91640]_ ;
  assign \new_[91644]_  = ~A166 & A167;
  assign \new_[91647]_  = ~A200 & ~A199;
  assign \new_[91648]_  = \new_[91647]_  & \new_[91644]_ ;
  assign \new_[91649]_  = \new_[91648]_  & \new_[91641]_ ;
  assign \new_[91652]_  = ~A268 & A267;
  assign \new_[91655]_  = A298 & A269;
  assign \new_[91656]_  = \new_[91655]_  & \new_[91652]_ ;
  assign \new_[91659]_  = ~A300 & ~A299;
  assign \new_[91662]_  = A302 & ~A301;
  assign \new_[91663]_  = \new_[91662]_  & \new_[91659]_ ;
  assign \new_[91664]_  = \new_[91663]_  & \new_[91656]_ ;
  assign \new_[91668]_  = ~A168 & ~A169;
  assign \new_[91669]_  = ~A170 & \new_[91668]_ ;
  assign \new_[91672]_  = ~A166 & A167;
  assign \new_[91675]_  = ~A200 & ~A199;
  assign \new_[91676]_  = \new_[91675]_  & \new_[91672]_ ;
  assign \new_[91677]_  = \new_[91676]_  & \new_[91669]_ ;
  assign \new_[91680]_  = ~A268 & A267;
  assign \new_[91683]_  = ~A298 & A269;
  assign \new_[91684]_  = \new_[91683]_  & \new_[91680]_ ;
  assign \new_[91687]_  = ~A300 & A299;
  assign \new_[91690]_  = A302 & ~A301;
  assign \new_[91691]_  = \new_[91690]_  & \new_[91687]_ ;
  assign \new_[91692]_  = \new_[91691]_  & \new_[91684]_ ;
  assign \new_[91696]_  = ~A168 & ~A169;
  assign \new_[91697]_  = ~A170 & \new_[91696]_ ;
  assign \new_[91700]_  = ~A166 & A167;
  assign \new_[91703]_  = ~A200 & ~A199;
  assign \new_[91704]_  = \new_[91703]_  & \new_[91700]_ ;
  assign \new_[91705]_  = \new_[91704]_  & \new_[91697]_ ;
  assign \new_[91708]_  = A266 & ~A265;
  assign \new_[91711]_  = ~A268 & ~A267;
  assign \new_[91712]_  = \new_[91711]_  & \new_[91708]_ ;
  assign \new_[91715]_  = A300 & A269;
  assign \new_[91718]_  = A302 & ~A301;
  assign \new_[91719]_  = \new_[91718]_  & \new_[91715]_ ;
  assign \new_[91720]_  = \new_[91719]_  & \new_[91712]_ ;
  assign \new_[91724]_  = ~A168 & ~A169;
  assign \new_[91725]_  = ~A170 & \new_[91724]_ ;
  assign \new_[91728]_  = ~A166 & A167;
  assign \new_[91731]_  = ~A200 & ~A199;
  assign \new_[91732]_  = \new_[91731]_  & \new_[91728]_ ;
  assign \new_[91733]_  = \new_[91732]_  & \new_[91725]_ ;
  assign \new_[91736]_  = ~A266 & A265;
  assign \new_[91739]_  = ~A268 & ~A267;
  assign \new_[91740]_  = \new_[91739]_  & \new_[91736]_ ;
  assign \new_[91743]_  = A300 & A269;
  assign \new_[91746]_  = A302 & ~A301;
  assign \new_[91747]_  = \new_[91746]_  & \new_[91743]_ ;
  assign \new_[91748]_  = \new_[91747]_  & \new_[91740]_ ;
  assign \new_[91752]_  = ~A168 & ~A169;
  assign \new_[91753]_  = ~A170 & \new_[91752]_ ;
  assign \new_[91756]_  = A166 & ~A167;
  assign \new_[91759]_  = ~A202 & A201;
  assign \new_[91760]_  = \new_[91759]_  & \new_[91756]_ ;
  assign \new_[91761]_  = \new_[91760]_  & \new_[91753]_ ;
  assign \new_[91764]_  = A267 & A203;
  assign \new_[91767]_  = A269 & ~A268;
  assign \new_[91768]_  = \new_[91767]_  & \new_[91764]_ ;
  assign \new_[91771]_  = ~A299 & A298;
  assign \new_[91774]_  = A301 & A300;
  assign \new_[91775]_  = \new_[91774]_  & \new_[91771]_ ;
  assign \new_[91776]_  = \new_[91775]_  & \new_[91768]_ ;
  assign \new_[91780]_  = ~A168 & ~A169;
  assign \new_[91781]_  = ~A170 & \new_[91780]_ ;
  assign \new_[91784]_  = A166 & ~A167;
  assign \new_[91787]_  = ~A202 & A201;
  assign \new_[91788]_  = \new_[91787]_  & \new_[91784]_ ;
  assign \new_[91789]_  = \new_[91788]_  & \new_[91781]_ ;
  assign \new_[91792]_  = A267 & A203;
  assign \new_[91795]_  = A269 & ~A268;
  assign \new_[91796]_  = \new_[91795]_  & \new_[91792]_ ;
  assign \new_[91799]_  = ~A299 & A298;
  assign \new_[91802]_  = ~A302 & A300;
  assign \new_[91803]_  = \new_[91802]_  & \new_[91799]_ ;
  assign \new_[91804]_  = \new_[91803]_  & \new_[91796]_ ;
  assign \new_[91808]_  = ~A168 & ~A169;
  assign \new_[91809]_  = ~A170 & \new_[91808]_ ;
  assign \new_[91812]_  = A166 & ~A167;
  assign \new_[91815]_  = ~A202 & A201;
  assign \new_[91816]_  = \new_[91815]_  & \new_[91812]_ ;
  assign \new_[91817]_  = \new_[91816]_  & \new_[91809]_ ;
  assign \new_[91820]_  = A267 & A203;
  assign \new_[91823]_  = A269 & ~A268;
  assign \new_[91824]_  = \new_[91823]_  & \new_[91820]_ ;
  assign \new_[91827]_  = A299 & ~A298;
  assign \new_[91830]_  = A301 & A300;
  assign \new_[91831]_  = \new_[91830]_  & \new_[91827]_ ;
  assign \new_[91832]_  = \new_[91831]_  & \new_[91824]_ ;
  assign \new_[91836]_  = ~A168 & ~A169;
  assign \new_[91837]_  = ~A170 & \new_[91836]_ ;
  assign \new_[91840]_  = A166 & ~A167;
  assign \new_[91843]_  = ~A202 & A201;
  assign \new_[91844]_  = \new_[91843]_  & \new_[91840]_ ;
  assign \new_[91845]_  = \new_[91844]_  & \new_[91837]_ ;
  assign \new_[91848]_  = A267 & A203;
  assign \new_[91851]_  = A269 & ~A268;
  assign \new_[91852]_  = \new_[91851]_  & \new_[91848]_ ;
  assign \new_[91855]_  = A299 & ~A298;
  assign \new_[91858]_  = ~A302 & A300;
  assign \new_[91859]_  = \new_[91858]_  & \new_[91855]_ ;
  assign \new_[91860]_  = \new_[91859]_  & \new_[91852]_ ;
  assign \new_[91864]_  = ~A168 & ~A169;
  assign \new_[91865]_  = ~A170 & \new_[91864]_ ;
  assign \new_[91868]_  = A166 & ~A167;
  assign \new_[91871]_  = ~A202 & A201;
  assign \new_[91872]_  = \new_[91871]_  & \new_[91868]_ ;
  assign \new_[91873]_  = \new_[91872]_  & \new_[91865]_ ;
  assign \new_[91876]_  = ~A267 & A203;
  assign \new_[91879]_  = A298 & A268;
  assign \new_[91880]_  = \new_[91879]_  & \new_[91876]_ ;
  assign \new_[91883]_  = ~A300 & ~A299;
  assign \new_[91886]_  = A302 & ~A301;
  assign \new_[91887]_  = \new_[91886]_  & \new_[91883]_ ;
  assign \new_[91888]_  = \new_[91887]_  & \new_[91880]_ ;
  assign \new_[91892]_  = ~A168 & ~A169;
  assign \new_[91893]_  = ~A170 & \new_[91892]_ ;
  assign \new_[91896]_  = A166 & ~A167;
  assign \new_[91899]_  = ~A202 & A201;
  assign \new_[91900]_  = \new_[91899]_  & \new_[91896]_ ;
  assign \new_[91901]_  = \new_[91900]_  & \new_[91893]_ ;
  assign \new_[91904]_  = ~A267 & A203;
  assign \new_[91907]_  = ~A298 & A268;
  assign \new_[91908]_  = \new_[91907]_  & \new_[91904]_ ;
  assign \new_[91911]_  = ~A300 & A299;
  assign \new_[91914]_  = A302 & ~A301;
  assign \new_[91915]_  = \new_[91914]_  & \new_[91911]_ ;
  assign \new_[91916]_  = \new_[91915]_  & \new_[91908]_ ;
  assign \new_[91920]_  = ~A168 & ~A169;
  assign \new_[91921]_  = ~A170 & \new_[91920]_ ;
  assign \new_[91924]_  = A166 & ~A167;
  assign \new_[91927]_  = ~A202 & A201;
  assign \new_[91928]_  = \new_[91927]_  & \new_[91924]_ ;
  assign \new_[91929]_  = \new_[91928]_  & \new_[91921]_ ;
  assign \new_[91932]_  = ~A267 & A203;
  assign \new_[91935]_  = A298 & ~A269;
  assign \new_[91936]_  = \new_[91935]_  & \new_[91932]_ ;
  assign \new_[91939]_  = ~A300 & ~A299;
  assign \new_[91942]_  = A302 & ~A301;
  assign \new_[91943]_  = \new_[91942]_  & \new_[91939]_ ;
  assign \new_[91944]_  = \new_[91943]_  & \new_[91936]_ ;
  assign \new_[91948]_  = ~A168 & ~A169;
  assign \new_[91949]_  = ~A170 & \new_[91948]_ ;
  assign \new_[91952]_  = A166 & ~A167;
  assign \new_[91955]_  = ~A202 & A201;
  assign \new_[91956]_  = \new_[91955]_  & \new_[91952]_ ;
  assign \new_[91957]_  = \new_[91956]_  & \new_[91949]_ ;
  assign \new_[91960]_  = ~A267 & A203;
  assign \new_[91963]_  = ~A298 & ~A269;
  assign \new_[91964]_  = \new_[91963]_  & \new_[91960]_ ;
  assign \new_[91967]_  = ~A300 & A299;
  assign \new_[91970]_  = A302 & ~A301;
  assign \new_[91971]_  = \new_[91970]_  & \new_[91967]_ ;
  assign \new_[91972]_  = \new_[91971]_  & \new_[91964]_ ;
  assign \new_[91976]_  = ~A168 & ~A169;
  assign \new_[91977]_  = ~A170 & \new_[91976]_ ;
  assign \new_[91980]_  = A166 & ~A167;
  assign \new_[91983]_  = ~A202 & A201;
  assign \new_[91984]_  = \new_[91983]_  & \new_[91980]_ ;
  assign \new_[91985]_  = \new_[91984]_  & \new_[91977]_ ;
  assign \new_[91988]_  = A265 & A203;
  assign \new_[91991]_  = A298 & A266;
  assign \new_[91992]_  = \new_[91991]_  & \new_[91988]_ ;
  assign \new_[91995]_  = ~A300 & ~A299;
  assign \new_[91998]_  = A302 & ~A301;
  assign \new_[91999]_  = \new_[91998]_  & \new_[91995]_ ;
  assign \new_[92000]_  = \new_[91999]_  & \new_[91992]_ ;
  assign \new_[92004]_  = ~A168 & ~A169;
  assign \new_[92005]_  = ~A170 & \new_[92004]_ ;
  assign \new_[92008]_  = A166 & ~A167;
  assign \new_[92011]_  = ~A202 & A201;
  assign \new_[92012]_  = \new_[92011]_  & \new_[92008]_ ;
  assign \new_[92013]_  = \new_[92012]_  & \new_[92005]_ ;
  assign \new_[92016]_  = A265 & A203;
  assign \new_[92019]_  = ~A298 & A266;
  assign \new_[92020]_  = \new_[92019]_  & \new_[92016]_ ;
  assign \new_[92023]_  = ~A300 & A299;
  assign \new_[92026]_  = A302 & ~A301;
  assign \new_[92027]_  = \new_[92026]_  & \new_[92023]_ ;
  assign \new_[92028]_  = \new_[92027]_  & \new_[92020]_ ;
  assign \new_[92032]_  = ~A168 & ~A169;
  assign \new_[92033]_  = ~A170 & \new_[92032]_ ;
  assign \new_[92036]_  = A166 & ~A167;
  assign \new_[92039]_  = ~A202 & A201;
  assign \new_[92040]_  = \new_[92039]_  & \new_[92036]_ ;
  assign \new_[92041]_  = \new_[92040]_  & \new_[92033]_ ;
  assign \new_[92044]_  = ~A265 & A203;
  assign \new_[92047]_  = A267 & A266;
  assign \new_[92048]_  = \new_[92047]_  & \new_[92044]_ ;
  assign \new_[92051]_  = A300 & A268;
  assign \new_[92054]_  = A302 & ~A301;
  assign \new_[92055]_  = \new_[92054]_  & \new_[92051]_ ;
  assign \new_[92056]_  = \new_[92055]_  & \new_[92048]_ ;
  assign \new_[92060]_  = ~A168 & ~A169;
  assign \new_[92061]_  = ~A170 & \new_[92060]_ ;
  assign \new_[92064]_  = A166 & ~A167;
  assign \new_[92067]_  = ~A202 & A201;
  assign \new_[92068]_  = \new_[92067]_  & \new_[92064]_ ;
  assign \new_[92069]_  = \new_[92068]_  & \new_[92061]_ ;
  assign \new_[92072]_  = ~A265 & A203;
  assign \new_[92075]_  = A267 & A266;
  assign \new_[92076]_  = \new_[92075]_  & \new_[92072]_ ;
  assign \new_[92079]_  = A300 & ~A269;
  assign \new_[92082]_  = A302 & ~A301;
  assign \new_[92083]_  = \new_[92082]_  & \new_[92079]_ ;
  assign \new_[92084]_  = \new_[92083]_  & \new_[92076]_ ;
  assign \new_[92088]_  = ~A168 & ~A169;
  assign \new_[92089]_  = ~A170 & \new_[92088]_ ;
  assign \new_[92092]_  = A166 & ~A167;
  assign \new_[92095]_  = ~A202 & A201;
  assign \new_[92096]_  = \new_[92095]_  & \new_[92092]_ ;
  assign \new_[92097]_  = \new_[92096]_  & \new_[92089]_ ;
  assign \new_[92100]_  = ~A265 & A203;
  assign \new_[92103]_  = ~A267 & A266;
  assign \new_[92104]_  = \new_[92103]_  & \new_[92100]_ ;
  assign \new_[92107]_  = A269 & ~A268;
  assign \new_[92110]_  = A301 & ~A300;
  assign \new_[92111]_  = \new_[92110]_  & \new_[92107]_ ;
  assign \new_[92112]_  = \new_[92111]_  & \new_[92104]_ ;
  assign \new_[92116]_  = ~A168 & ~A169;
  assign \new_[92117]_  = ~A170 & \new_[92116]_ ;
  assign \new_[92120]_  = A166 & ~A167;
  assign \new_[92123]_  = ~A202 & A201;
  assign \new_[92124]_  = \new_[92123]_  & \new_[92120]_ ;
  assign \new_[92125]_  = \new_[92124]_  & \new_[92117]_ ;
  assign \new_[92128]_  = ~A265 & A203;
  assign \new_[92131]_  = ~A267 & A266;
  assign \new_[92132]_  = \new_[92131]_  & \new_[92128]_ ;
  assign \new_[92135]_  = A269 & ~A268;
  assign \new_[92138]_  = ~A302 & ~A300;
  assign \new_[92139]_  = \new_[92138]_  & \new_[92135]_ ;
  assign \new_[92140]_  = \new_[92139]_  & \new_[92132]_ ;
  assign \new_[92144]_  = ~A168 & ~A169;
  assign \new_[92145]_  = ~A170 & \new_[92144]_ ;
  assign \new_[92148]_  = A166 & ~A167;
  assign \new_[92151]_  = ~A202 & A201;
  assign \new_[92152]_  = \new_[92151]_  & \new_[92148]_ ;
  assign \new_[92153]_  = \new_[92152]_  & \new_[92145]_ ;
  assign \new_[92156]_  = ~A265 & A203;
  assign \new_[92159]_  = ~A267 & A266;
  assign \new_[92160]_  = \new_[92159]_  & \new_[92156]_ ;
  assign \new_[92163]_  = A269 & ~A268;
  assign \new_[92166]_  = A299 & A298;
  assign \new_[92167]_  = \new_[92166]_  & \new_[92163]_ ;
  assign \new_[92168]_  = \new_[92167]_  & \new_[92160]_ ;
  assign \new_[92172]_  = ~A168 & ~A169;
  assign \new_[92173]_  = ~A170 & \new_[92172]_ ;
  assign \new_[92176]_  = A166 & ~A167;
  assign \new_[92179]_  = ~A202 & A201;
  assign \new_[92180]_  = \new_[92179]_  & \new_[92176]_ ;
  assign \new_[92181]_  = \new_[92180]_  & \new_[92173]_ ;
  assign \new_[92184]_  = ~A265 & A203;
  assign \new_[92187]_  = ~A267 & A266;
  assign \new_[92188]_  = \new_[92187]_  & \new_[92184]_ ;
  assign \new_[92191]_  = A269 & ~A268;
  assign \new_[92194]_  = ~A299 & ~A298;
  assign \new_[92195]_  = \new_[92194]_  & \new_[92191]_ ;
  assign \new_[92196]_  = \new_[92195]_  & \new_[92188]_ ;
  assign \new_[92200]_  = ~A168 & ~A169;
  assign \new_[92201]_  = ~A170 & \new_[92200]_ ;
  assign \new_[92204]_  = A166 & ~A167;
  assign \new_[92207]_  = ~A202 & A201;
  assign \new_[92208]_  = \new_[92207]_  & \new_[92204]_ ;
  assign \new_[92209]_  = \new_[92208]_  & \new_[92201]_ ;
  assign \new_[92212]_  = A265 & A203;
  assign \new_[92215]_  = A267 & ~A266;
  assign \new_[92216]_  = \new_[92215]_  & \new_[92212]_ ;
  assign \new_[92219]_  = A300 & A268;
  assign \new_[92222]_  = A302 & ~A301;
  assign \new_[92223]_  = \new_[92222]_  & \new_[92219]_ ;
  assign \new_[92224]_  = \new_[92223]_  & \new_[92216]_ ;
  assign \new_[92228]_  = ~A168 & ~A169;
  assign \new_[92229]_  = ~A170 & \new_[92228]_ ;
  assign \new_[92232]_  = A166 & ~A167;
  assign \new_[92235]_  = ~A202 & A201;
  assign \new_[92236]_  = \new_[92235]_  & \new_[92232]_ ;
  assign \new_[92237]_  = \new_[92236]_  & \new_[92229]_ ;
  assign \new_[92240]_  = A265 & A203;
  assign \new_[92243]_  = A267 & ~A266;
  assign \new_[92244]_  = \new_[92243]_  & \new_[92240]_ ;
  assign \new_[92247]_  = A300 & ~A269;
  assign \new_[92250]_  = A302 & ~A301;
  assign \new_[92251]_  = \new_[92250]_  & \new_[92247]_ ;
  assign \new_[92252]_  = \new_[92251]_  & \new_[92244]_ ;
  assign \new_[92256]_  = ~A168 & ~A169;
  assign \new_[92257]_  = ~A170 & \new_[92256]_ ;
  assign \new_[92260]_  = A166 & ~A167;
  assign \new_[92263]_  = ~A202 & A201;
  assign \new_[92264]_  = \new_[92263]_  & \new_[92260]_ ;
  assign \new_[92265]_  = \new_[92264]_  & \new_[92257]_ ;
  assign \new_[92268]_  = A265 & A203;
  assign \new_[92271]_  = ~A267 & ~A266;
  assign \new_[92272]_  = \new_[92271]_  & \new_[92268]_ ;
  assign \new_[92275]_  = A269 & ~A268;
  assign \new_[92278]_  = A301 & ~A300;
  assign \new_[92279]_  = \new_[92278]_  & \new_[92275]_ ;
  assign \new_[92280]_  = \new_[92279]_  & \new_[92272]_ ;
  assign \new_[92284]_  = ~A168 & ~A169;
  assign \new_[92285]_  = ~A170 & \new_[92284]_ ;
  assign \new_[92288]_  = A166 & ~A167;
  assign \new_[92291]_  = ~A202 & A201;
  assign \new_[92292]_  = \new_[92291]_  & \new_[92288]_ ;
  assign \new_[92293]_  = \new_[92292]_  & \new_[92285]_ ;
  assign \new_[92296]_  = A265 & A203;
  assign \new_[92299]_  = ~A267 & ~A266;
  assign \new_[92300]_  = \new_[92299]_  & \new_[92296]_ ;
  assign \new_[92303]_  = A269 & ~A268;
  assign \new_[92306]_  = ~A302 & ~A300;
  assign \new_[92307]_  = \new_[92306]_  & \new_[92303]_ ;
  assign \new_[92308]_  = \new_[92307]_  & \new_[92300]_ ;
  assign \new_[92312]_  = ~A168 & ~A169;
  assign \new_[92313]_  = ~A170 & \new_[92312]_ ;
  assign \new_[92316]_  = A166 & ~A167;
  assign \new_[92319]_  = ~A202 & A201;
  assign \new_[92320]_  = \new_[92319]_  & \new_[92316]_ ;
  assign \new_[92321]_  = \new_[92320]_  & \new_[92313]_ ;
  assign \new_[92324]_  = A265 & A203;
  assign \new_[92327]_  = ~A267 & ~A266;
  assign \new_[92328]_  = \new_[92327]_  & \new_[92324]_ ;
  assign \new_[92331]_  = A269 & ~A268;
  assign \new_[92334]_  = A299 & A298;
  assign \new_[92335]_  = \new_[92334]_  & \new_[92331]_ ;
  assign \new_[92336]_  = \new_[92335]_  & \new_[92328]_ ;
  assign \new_[92340]_  = ~A168 & ~A169;
  assign \new_[92341]_  = ~A170 & \new_[92340]_ ;
  assign \new_[92344]_  = A166 & ~A167;
  assign \new_[92347]_  = ~A202 & A201;
  assign \new_[92348]_  = \new_[92347]_  & \new_[92344]_ ;
  assign \new_[92349]_  = \new_[92348]_  & \new_[92341]_ ;
  assign \new_[92352]_  = A265 & A203;
  assign \new_[92355]_  = ~A267 & ~A266;
  assign \new_[92356]_  = \new_[92355]_  & \new_[92352]_ ;
  assign \new_[92359]_  = A269 & ~A268;
  assign \new_[92362]_  = ~A299 & ~A298;
  assign \new_[92363]_  = \new_[92362]_  & \new_[92359]_ ;
  assign \new_[92364]_  = \new_[92363]_  & \new_[92356]_ ;
  assign \new_[92368]_  = ~A168 & ~A169;
  assign \new_[92369]_  = ~A170 & \new_[92368]_ ;
  assign \new_[92372]_  = A166 & ~A167;
  assign \new_[92375]_  = ~A202 & A201;
  assign \new_[92376]_  = \new_[92375]_  & \new_[92372]_ ;
  assign \new_[92377]_  = \new_[92376]_  & \new_[92369]_ ;
  assign \new_[92380]_  = ~A265 & A203;
  assign \new_[92383]_  = A298 & ~A266;
  assign \new_[92384]_  = \new_[92383]_  & \new_[92380]_ ;
  assign \new_[92387]_  = ~A300 & ~A299;
  assign \new_[92390]_  = A302 & ~A301;
  assign \new_[92391]_  = \new_[92390]_  & \new_[92387]_ ;
  assign \new_[92392]_  = \new_[92391]_  & \new_[92384]_ ;
  assign \new_[92396]_  = ~A168 & ~A169;
  assign \new_[92397]_  = ~A170 & \new_[92396]_ ;
  assign \new_[92400]_  = A166 & ~A167;
  assign \new_[92403]_  = ~A202 & A201;
  assign \new_[92404]_  = \new_[92403]_  & \new_[92400]_ ;
  assign \new_[92405]_  = \new_[92404]_  & \new_[92397]_ ;
  assign \new_[92408]_  = ~A265 & A203;
  assign \new_[92411]_  = ~A298 & ~A266;
  assign \new_[92412]_  = \new_[92411]_  & \new_[92408]_ ;
  assign \new_[92415]_  = ~A300 & A299;
  assign \new_[92418]_  = A302 & ~A301;
  assign \new_[92419]_  = \new_[92418]_  & \new_[92415]_ ;
  assign \new_[92420]_  = \new_[92419]_  & \new_[92412]_ ;
  assign \new_[92424]_  = ~A168 & ~A169;
  assign \new_[92425]_  = ~A170 & \new_[92424]_ ;
  assign \new_[92428]_  = A166 & ~A167;
  assign \new_[92431]_  = A202 & ~A201;
  assign \new_[92432]_  = \new_[92431]_  & \new_[92428]_ ;
  assign \new_[92433]_  = \new_[92432]_  & \new_[92425]_ ;
  assign \new_[92436]_  = ~A268 & A267;
  assign \new_[92439]_  = A298 & A269;
  assign \new_[92440]_  = \new_[92439]_  & \new_[92436]_ ;
  assign \new_[92443]_  = ~A300 & ~A299;
  assign \new_[92446]_  = A302 & ~A301;
  assign \new_[92447]_  = \new_[92446]_  & \new_[92443]_ ;
  assign \new_[92448]_  = \new_[92447]_  & \new_[92440]_ ;
  assign \new_[92452]_  = ~A168 & ~A169;
  assign \new_[92453]_  = ~A170 & \new_[92452]_ ;
  assign \new_[92456]_  = A166 & ~A167;
  assign \new_[92459]_  = A202 & ~A201;
  assign \new_[92460]_  = \new_[92459]_  & \new_[92456]_ ;
  assign \new_[92461]_  = \new_[92460]_  & \new_[92453]_ ;
  assign \new_[92464]_  = ~A268 & A267;
  assign \new_[92467]_  = ~A298 & A269;
  assign \new_[92468]_  = \new_[92467]_  & \new_[92464]_ ;
  assign \new_[92471]_  = ~A300 & A299;
  assign \new_[92474]_  = A302 & ~A301;
  assign \new_[92475]_  = \new_[92474]_  & \new_[92471]_ ;
  assign \new_[92476]_  = \new_[92475]_  & \new_[92468]_ ;
  assign \new_[92480]_  = ~A168 & ~A169;
  assign \new_[92481]_  = ~A170 & \new_[92480]_ ;
  assign \new_[92484]_  = A166 & ~A167;
  assign \new_[92487]_  = A202 & ~A201;
  assign \new_[92488]_  = \new_[92487]_  & \new_[92484]_ ;
  assign \new_[92489]_  = \new_[92488]_  & \new_[92481]_ ;
  assign \new_[92492]_  = A266 & ~A265;
  assign \new_[92495]_  = ~A268 & ~A267;
  assign \new_[92496]_  = \new_[92495]_  & \new_[92492]_ ;
  assign \new_[92499]_  = A300 & A269;
  assign \new_[92502]_  = A302 & ~A301;
  assign \new_[92503]_  = \new_[92502]_  & \new_[92499]_ ;
  assign \new_[92504]_  = \new_[92503]_  & \new_[92496]_ ;
  assign \new_[92508]_  = ~A168 & ~A169;
  assign \new_[92509]_  = ~A170 & \new_[92508]_ ;
  assign \new_[92512]_  = A166 & ~A167;
  assign \new_[92515]_  = A202 & ~A201;
  assign \new_[92516]_  = \new_[92515]_  & \new_[92512]_ ;
  assign \new_[92517]_  = \new_[92516]_  & \new_[92509]_ ;
  assign \new_[92520]_  = ~A266 & A265;
  assign \new_[92523]_  = ~A268 & ~A267;
  assign \new_[92524]_  = \new_[92523]_  & \new_[92520]_ ;
  assign \new_[92527]_  = A300 & A269;
  assign \new_[92530]_  = A302 & ~A301;
  assign \new_[92531]_  = \new_[92530]_  & \new_[92527]_ ;
  assign \new_[92532]_  = \new_[92531]_  & \new_[92524]_ ;
  assign \new_[92536]_  = ~A168 & ~A169;
  assign \new_[92537]_  = ~A170 & \new_[92536]_ ;
  assign \new_[92540]_  = A166 & ~A167;
  assign \new_[92543]_  = ~A203 & ~A201;
  assign \new_[92544]_  = \new_[92543]_  & \new_[92540]_ ;
  assign \new_[92545]_  = \new_[92544]_  & \new_[92537]_ ;
  assign \new_[92548]_  = ~A268 & A267;
  assign \new_[92551]_  = A298 & A269;
  assign \new_[92552]_  = \new_[92551]_  & \new_[92548]_ ;
  assign \new_[92555]_  = ~A300 & ~A299;
  assign \new_[92558]_  = A302 & ~A301;
  assign \new_[92559]_  = \new_[92558]_  & \new_[92555]_ ;
  assign \new_[92560]_  = \new_[92559]_  & \new_[92552]_ ;
  assign \new_[92564]_  = ~A168 & ~A169;
  assign \new_[92565]_  = ~A170 & \new_[92564]_ ;
  assign \new_[92568]_  = A166 & ~A167;
  assign \new_[92571]_  = ~A203 & ~A201;
  assign \new_[92572]_  = \new_[92571]_  & \new_[92568]_ ;
  assign \new_[92573]_  = \new_[92572]_  & \new_[92565]_ ;
  assign \new_[92576]_  = ~A268 & A267;
  assign \new_[92579]_  = ~A298 & A269;
  assign \new_[92580]_  = \new_[92579]_  & \new_[92576]_ ;
  assign \new_[92583]_  = ~A300 & A299;
  assign \new_[92586]_  = A302 & ~A301;
  assign \new_[92587]_  = \new_[92586]_  & \new_[92583]_ ;
  assign \new_[92588]_  = \new_[92587]_  & \new_[92580]_ ;
  assign \new_[92592]_  = ~A168 & ~A169;
  assign \new_[92593]_  = ~A170 & \new_[92592]_ ;
  assign \new_[92596]_  = A166 & ~A167;
  assign \new_[92599]_  = ~A203 & ~A201;
  assign \new_[92600]_  = \new_[92599]_  & \new_[92596]_ ;
  assign \new_[92601]_  = \new_[92600]_  & \new_[92593]_ ;
  assign \new_[92604]_  = A266 & ~A265;
  assign \new_[92607]_  = ~A268 & ~A267;
  assign \new_[92608]_  = \new_[92607]_  & \new_[92604]_ ;
  assign \new_[92611]_  = A300 & A269;
  assign \new_[92614]_  = A302 & ~A301;
  assign \new_[92615]_  = \new_[92614]_  & \new_[92611]_ ;
  assign \new_[92616]_  = \new_[92615]_  & \new_[92608]_ ;
  assign \new_[92620]_  = ~A168 & ~A169;
  assign \new_[92621]_  = ~A170 & \new_[92620]_ ;
  assign \new_[92624]_  = A166 & ~A167;
  assign \new_[92627]_  = ~A203 & ~A201;
  assign \new_[92628]_  = \new_[92627]_  & \new_[92624]_ ;
  assign \new_[92629]_  = \new_[92628]_  & \new_[92621]_ ;
  assign \new_[92632]_  = ~A266 & A265;
  assign \new_[92635]_  = ~A268 & ~A267;
  assign \new_[92636]_  = \new_[92635]_  & \new_[92632]_ ;
  assign \new_[92639]_  = A300 & A269;
  assign \new_[92642]_  = A302 & ~A301;
  assign \new_[92643]_  = \new_[92642]_  & \new_[92639]_ ;
  assign \new_[92644]_  = \new_[92643]_  & \new_[92636]_ ;
  assign \new_[92648]_  = ~A168 & ~A169;
  assign \new_[92649]_  = ~A170 & \new_[92648]_ ;
  assign \new_[92652]_  = A166 & ~A167;
  assign \new_[92655]_  = A200 & A199;
  assign \new_[92656]_  = \new_[92655]_  & \new_[92652]_ ;
  assign \new_[92657]_  = \new_[92656]_  & \new_[92649]_ ;
  assign \new_[92660]_  = ~A268 & A267;
  assign \new_[92663]_  = A298 & A269;
  assign \new_[92664]_  = \new_[92663]_  & \new_[92660]_ ;
  assign \new_[92667]_  = ~A300 & ~A299;
  assign \new_[92670]_  = A302 & ~A301;
  assign \new_[92671]_  = \new_[92670]_  & \new_[92667]_ ;
  assign \new_[92672]_  = \new_[92671]_  & \new_[92664]_ ;
  assign \new_[92676]_  = ~A168 & ~A169;
  assign \new_[92677]_  = ~A170 & \new_[92676]_ ;
  assign \new_[92680]_  = A166 & ~A167;
  assign \new_[92683]_  = A200 & A199;
  assign \new_[92684]_  = \new_[92683]_  & \new_[92680]_ ;
  assign \new_[92685]_  = \new_[92684]_  & \new_[92677]_ ;
  assign \new_[92688]_  = ~A268 & A267;
  assign \new_[92691]_  = ~A298 & A269;
  assign \new_[92692]_  = \new_[92691]_  & \new_[92688]_ ;
  assign \new_[92695]_  = ~A300 & A299;
  assign \new_[92698]_  = A302 & ~A301;
  assign \new_[92699]_  = \new_[92698]_  & \new_[92695]_ ;
  assign \new_[92700]_  = \new_[92699]_  & \new_[92692]_ ;
  assign \new_[92704]_  = ~A168 & ~A169;
  assign \new_[92705]_  = ~A170 & \new_[92704]_ ;
  assign \new_[92708]_  = A166 & ~A167;
  assign \new_[92711]_  = A200 & A199;
  assign \new_[92712]_  = \new_[92711]_  & \new_[92708]_ ;
  assign \new_[92713]_  = \new_[92712]_  & \new_[92705]_ ;
  assign \new_[92716]_  = A266 & ~A265;
  assign \new_[92719]_  = ~A268 & ~A267;
  assign \new_[92720]_  = \new_[92719]_  & \new_[92716]_ ;
  assign \new_[92723]_  = A300 & A269;
  assign \new_[92726]_  = A302 & ~A301;
  assign \new_[92727]_  = \new_[92726]_  & \new_[92723]_ ;
  assign \new_[92728]_  = \new_[92727]_  & \new_[92720]_ ;
  assign \new_[92732]_  = ~A168 & ~A169;
  assign \new_[92733]_  = ~A170 & \new_[92732]_ ;
  assign \new_[92736]_  = A166 & ~A167;
  assign \new_[92739]_  = A200 & A199;
  assign \new_[92740]_  = \new_[92739]_  & \new_[92736]_ ;
  assign \new_[92741]_  = \new_[92740]_  & \new_[92733]_ ;
  assign \new_[92744]_  = ~A266 & A265;
  assign \new_[92747]_  = ~A268 & ~A267;
  assign \new_[92748]_  = \new_[92747]_  & \new_[92744]_ ;
  assign \new_[92751]_  = A300 & A269;
  assign \new_[92754]_  = A302 & ~A301;
  assign \new_[92755]_  = \new_[92754]_  & \new_[92751]_ ;
  assign \new_[92756]_  = \new_[92755]_  & \new_[92748]_ ;
  assign \new_[92760]_  = ~A168 & ~A169;
  assign \new_[92761]_  = ~A170 & \new_[92760]_ ;
  assign \new_[92764]_  = A166 & ~A167;
  assign \new_[92767]_  = ~A200 & ~A199;
  assign \new_[92768]_  = \new_[92767]_  & \new_[92764]_ ;
  assign \new_[92769]_  = \new_[92768]_  & \new_[92761]_ ;
  assign \new_[92772]_  = ~A268 & A267;
  assign \new_[92775]_  = A298 & A269;
  assign \new_[92776]_  = \new_[92775]_  & \new_[92772]_ ;
  assign \new_[92779]_  = ~A300 & ~A299;
  assign \new_[92782]_  = A302 & ~A301;
  assign \new_[92783]_  = \new_[92782]_  & \new_[92779]_ ;
  assign \new_[92784]_  = \new_[92783]_  & \new_[92776]_ ;
  assign \new_[92788]_  = ~A168 & ~A169;
  assign \new_[92789]_  = ~A170 & \new_[92788]_ ;
  assign \new_[92792]_  = A166 & ~A167;
  assign \new_[92795]_  = ~A200 & ~A199;
  assign \new_[92796]_  = \new_[92795]_  & \new_[92792]_ ;
  assign \new_[92797]_  = \new_[92796]_  & \new_[92789]_ ;
  assign \new_[92800]_  = ~A268 & A267;
  assign \new_[92803]_  = ~A298 & A269;
  assign \new_[92804]_  = \new_[92803]_  & \new_[92800]_ ;
  assign \new_[92807]_  = ~A300 & A299;
  assign \new_[92810]_  = A302 & ~A301;
  assign \new_[92811]_  = \new_[92810]_  & \new_[92807]_ ;
  assign \new_[92812]_  = \new_[92811]_  & \new_[92804]_ ;
  assign \new_[92816]_  = ~A168 & ~A169;
  assign \new_[92817]_  = ~A170 & \new_[92816]_ ;
  assign \new_[92820]_  = A166 & ~A167;
  assign \new_[92823]_  = ~A200 & ~A199;
  assign \new_[92824]_  = \new_[92823]_  & \new_[92820]_ ;
  assign \new_[92825]_  = \new_[92824]_  & \new_[92817]_ ;
  assign \new_[92828]_  = A266 & ~A265;
  assign \new_[92831]_  = ~A268 & ~A267;
  assign \new_[92832]_  = \new_[92831]_  & \new_[92828]_ ;
  assign \new_[92835]_  = A300 & A269;
  assign \new_[92838]_  = A302 & ~A301;
  assign \new_[92839]_  = \new_[92838]_  & \new_[92835]_ ;
  assign \new_[92840]_  = \new_[92839]_  & \new_[92832]_ ;
  assign \new_[92844]_  = ~A168 & ~A169;
  assign \new_[92845]_  = ~A170 & \new_[92844]_ ;
  assign \new_[92848]_  = A166 & ~A167;
  assign \new_[92851]_  = ~A200 & ~A199;
  assign \new_[92852]_  = \new_[92851]_  & \new_[92848]_ ;
  assign \new_[92853]_  = \new_[92852]_  & \new_[92845]_ ;
  assign \new_[92856]_  = ~A266 & A265;
  assign \new_[92859]_  = ~A268 & ~A267;
  assign \new_[92860]_  = \new_[92859]_  & \new_[92856]_ ;
  assign \new_[92863]_  = A300 & A269;
  assign \new_[92866]_  = A302 & ~A301;
  assign \new_[92867]_  = \new_[92866]_  & \new_[92863]_ ;
  assign \new_[92868]_  = \new_[92867]_  & \new_[92860]_ ;
  assign \new_[92871]_  = A166 & A167;
  assign \new_[92874]_  = A200 & ~A199;
  assign \new_[92875]_  = \new_[92874]_  & \new_[92871]_ ;
  assign \new_[92878]_  = A202 & A201;
  assign \new_[92881]_  = A266 & ~A265;
  assign \new_[92882]_  = \new_[92881]_  & \new_[92878]_ ;
  assign \new_[92883]_  = \new_[92882]_  & \new_[92875]_ ;
  assign \new_[92886]_  = ~A268 & ~A267;
  assign \new_[92889]_  = A298 & A269;
  assign \new_[92890]_  = \new_[92889]_  & \new_[92886]_ ;
  assign \new_[92893]_  = ~A300 & ~A299;
  assign \new_[92896]_  = A302 & ~A301;
  assign \new_[92897]_  = \new_[92896]_  & \new_[92893]_ ;
  assign \new_[92898]_  = \new_[92897]_  & \new_[92890]_ ;
  assign \new_[92901]_  = A166 & A167;
  assign \new_[92904]_  = A200 & ~A199;
  assign \new_[92905]_  = \new_[92904]_  & \new_[92901]_ ;
  assign \new_[92908]_  = A202 & A201;
  assign \new_[92911]_  = A266 & ~A265;
  assign \new_[92912]_  = \new_[92911]_  & \new_[92908]_ ;
  assign \new_[92913]_  = \new_[92912]_  & \new_[92905]_ ;
  assign \new_[92916]_  = ~A268 & ~A267;
  assign \new_[92919]_  = ~A298 & A269;
  assign \new_[92920]_  = \new_[92919]_  & \new_[92916]_ ;
  assign \new_[92923]_  = ~A300 & A299;
  assign \new_[92926]_  = A302 & ~A301;
  assign \new_[92927]_  = \new_[92926]_  & \new_[92923]_ ;
  assign \new_[92928]_  = \new_[92927]_  & \new_[92920]_ ;
  assign \new_[92931]_  = A166 & A167;
  assign \new_[92934]_  = A200 & ~A199;
  assign \new_[92935]_  = \new_[92934]_  & \new_[92931]_ ;
  assign \new_[92938]_  = A202 & A201;
  assign \new_[92941]_  = ~A266 & A265;
  assign \new_[92942]_  = \new_[92941]_  & \new_[92938]_ ;
  assign \new_[92943]_  = \new_[92942]_  & \new_[92935]_ ;
  assign \new_[92946]_  = ~A268 & ~A267;
  assign \new_[92949]_  = A298 & A269;
  assign \new_[92950]_  = \new_[92949]_  & \new_[92946]_ ;
  assign \new_[92953]_  = ~A300 & ~A299;
  assign \new_[92956]_  = A302 & ~A301;
  assign \new_[92957]_  = \new_[92956]_  & \new_[92953]_ ;
  assign \new_[92958]_  = \new_[92957]_  & \new_[92950]_ ;
  assign \new_[92961]_  = A166 & A167;
  assign \new_[92964]_  = A200 & ~A199;
  assign \new_[92965]_  = \new_[92964]_  & \new_[92961]_ ;
  assign \new_[92968]_  = A202 & A201;
  assign \new_[92971]_  = ~A266 & A265;
  assign \new_[92972]_  = \new_[92971]_  & \new_[92968]_ ;
  assign \new_[92973]_  = \new_[92972]_  & \new_[92965]_ ;
  assign \new_[92976]_  = ~A268 & ~A267;
  assign \new_[92979]_  = ~A298 & A269;
  assign \new_[92980]_  = \new_[92979]_  & \new_[92976]_ ;
  assign \new_[92983]_  = ~A300 & A299;
  assign \new_[92986]_  = A302 & ~A301;
  assign \new_[92987]_  = \new_[92986]_  & \new_[92983]_ ;
  assign \new_[92988]_  = \new_[92987]_  & \new_[92980]_ ;
  assign \new_[92991]_  = A166 & A167;
  assign \new_[92994]_  = A200 & ~A199;
  assign \new_[92995]_  = \new_[92994]_  & \new_[92991]_ ;
  assign \new_[92998]_  = ~A203 & A201;
  assign \new_[93001]_  = A266 & ~A265;
  assign \new_[93002]_  = \new_[93001]_  & \new_[92998]_ ;
  assign \new_[93003]_  = \new_[93002]_  & \new_[92995]_ ;
  assign \new_[93006]_  = ~A268 & ~A267;
  assign \new_[93009]_  = A298 & A269;
  assign \new_[93010]_  = \new_[93009]_  & \new_[93006]_ ;
  assign \new_[93013]_  = ~A300 & ~A299;
  assign \new_[93016]_  = A302 & ~A301;
  assign \new_[93017]_  = \new_[93016]_  & \new_[93013]_ ;
  assign \new_[93018]_  = \new_[93017]_  & \new_[93010]_ ;
  assign \new_[93021]_  = A166 & A167;
  assign \new_[93024]_  = A200 & ~A199;
  assign \new_[93025]_  = \new_[93024]_  & \new_[93021]_ ;
  assign \new_[93028]_  = ~A203 & A201;
  assign \new_[93031]_  = A266 & ~A265;
  assign \new_[93032]_  = \new_[93031]_  & \new_[93028]_ ;
  assign \new_[93033]_  = \new_[93032]_  & \new_[93025]_ ;
  assign \new_[93036]_  = ~A268 & ~A267;
  assign \new_[93039]_  = ~A298 & A269;
  assign \new_[93040]_  = \new_[93039]_  & \new_[93036]_ ;
  assign \new_[93043]_  = ~A300 & A299;
  assign \new_[93046]_  = A302 & ~A301;
  assign \new_[93047]_  = \new_[93046]_  & \new_[93043]_ ;
  assign \new_[93048]_  = \new_[93047]_  & \new_[93040]_ ;
  assign \new_[93051]_  = A166 & A167;
  assign \new_[93054]_  = A200 & ~A199;
  assign \new_[93055]_  = \new_[93054]_  & \new_[93051]_ ;
  assign \new_[93058]_  = ~A203 & A201;
  assign \new_[93061]_  = ~A266 & A265;
  assign \new_[93062]_  = \new_[93061]_  & \new_[93058]_ ;
  assign \new_[93063]_  = \new_[93062]_  & \new_[93055]_ ;
  assign \new_[93066]_  = ~A268 & ~A267;
  assign \new_[93069]_  = A298 & A269;
  assign \new_[93070]_  = \new_[93069]_  & \new_[93066]_ ;
  assign \new_[93073]_  = ~A300 & ~A299;
  assign \new_[93076]_  = A302 & ~A301;
  assign \new_[93077]_  = \new_[93076]_  & \new_[93073]_ ;
  assign \new_[93078]_  = \new_[93077]_  & \new_[93070]_ ;
  assign \new_[93081]_  = A166 & A167;
  assign \new_[93084]_  = A200 & ~A199;
  assign \new_[93085]_  = \new_[93084]_  & \new_[93081]_ ;
  assign \new_[93088]_  = ~A203 & A201;
  assign \new_[93091]_  = ~A266 & A265;
  assign \new_[93092]_  = \new_[93091]_  & \new_[93088]_ ;
  assign \new_[93093]_  = \new_[93092]_  & \new_[93085]_ ;
  assign \new_[93096]_  = ~A268 & ~A267;
  assign \new_[93099]_  = ~A298 & A269;
  assign \new_[93100]_  = \new_[93099]_  & \new_[93096]_ ;
  assign \new_[93103]_  = ~A300 & A299;
  assign \new_[93106]_  = A302 & ~A301;
  assign \new_[93107]_  = \new_[93106]_  & \new_[93103]_ ;
  assign \new_[93108]_  = \new_[93107]_  & \new_[93100]_ ;
  assign \new_[93111]_  = A166 & A167;
  assign \new_[93114]_  = A200 & ~A199;
  assign \new_[93115]_  = \new_[93114]_  & \new_[93111]_ ;
  assign \new_[93118]_  = ~A202 & ~A201;
  assign \new_[93121]_  = ~A265 & A203;
  assign \new_[93122]_  = \new_[93121]_  & \new_[93118]_ ;
  assign \new_[93123]_  = \new_[93122]_  & \new_[93115]_ ;
  assign \new_[93126]_  = A267 & A266;
  assign \new_[93129]_  = A298 & A268;
  assign \new_[93130]_  = \new_[93129]_  & \new_[93126]_ ;
  assign \new_[93133]_  = ~A300 & ~A299;
  assign \new_[93136]_  = A302 & ~A301;
  assign \new_[93137]_  = \new_[93136]_  & \new_[93133]_ ;
  assign \new_[93138]_  = \new_[93137]_  & \new_[93130]_ ;
  assign \new_[93141]_  = A166 & A167;
  assign \new_[93144]_  = A200 & ~A199;
  assign \new_[93145]_  = \new_[93144]_  & \new_[93141]_ ;
  assign \new_[93148]_  = ~A202 & ~A201;
  assign \new_[93151]_  = ~A265 & A203;
  assign \new_[93152]_  = \new_[93151]_  & \new_[93148]_ ;
  assign \new_[93153]_  = \new_[93152]_  & \new_[93145]_ ;
  assign \new_[93156]_  = A267 & A266;
  assign \new_[93159]_  = ~A298 & A268;
  assign \new_[93160]_  = \new_[93159]_  & \new_[93156]_ ;
  assign \new_[93163]_  = ~A300 & A299;
  assign \new_[93166]_  = A302 & ~A301;
  assign \new_[93167]_  = \new_[93166]_  & \new_[93163]_ ;
  assign \new_[93168]_  = \new_[93167]_  & \new_[93160]_ ;
  assign \new_[93171]_  = A166 & A167;
  assign \new_[93174]_  = A200 & ~A199;
  assign \new_[93175]_  = \new_[93174]_  & \new_[93171]_ ;
  assign \new_[93178]_  = ~A202 & ~A201;
  assign \new_[93181]_  = ~A265 & A203;
  assign \new_[93182]_  = \new_[93181]_  & \new_[93178]_ ;
  assign \new_[93183]_  = \new_[93182]_  & \new_[93175]_ ;
  assign \new_[93186]_  = A267 & A266;
  assign \new_[93189]_  = A298 & ~A269;
  assign \new_[93190]_  = \new_[93189]_  & \new_[93186]_ ;
  assign \new_[93193]_  = ~A300 & ~A299;
  assign \new_[93196]_  = A302 & ~A301;
  assign \new_[93197]_  = \new_[93196]_  & \new_[93193]_ ;
  assign \new_[93198]_  = \new_[93197]_  & \new_[93190]_ ;
  assign \new_[93201]_  = A166 & A167;
  assign \new_[93204]_  = A200 & ~A199;
  assign \new_[93205]_  = \new_[93204]_  & \new_[93201]_ ;
  assign \new_[93208]_  = ~A202 & ~A201;
  assign \new_[93211]_  = ~A265 & A203;
  assign \new_[93212]_  = \new_[93211]_  & \new_[93208]_ ;
  assign \new_[93213]_  = \new_[93212]_  & \new_[93205]_ ;
  assign \new_[93216]_  = A267 & A266;
  assign \new_[93219]_  = ~A298 & ~A269;
  assign \new_[93220]_  = \new_[93219]_  & \new_[93216]_ ;
  assign \new_[93223]_  = ~A300 & A299;
  assign \new_[93226]_  = A302 & ~A301;
  assign \new_[93227]_  = \new_[93226]_  & \new_[93223]_ ;
  assign \new_[93228]_  = \new_[93227]_  & \new_[93220]_ ;
  assign \new_[93231]_  = A166 & A167;
  assign \new_[93234]_  = A200 & ~A199;
  assign \new_[93235]_  = \new_[93234]_  & \new_[93231]_ ;
  assign \new_[93238]_  = ~A202 & ~A201;
  assign \new_[93241]_  = ~A265 & A203;
  assign \new_[93242]_  = \new_[93241]_  & \new_[93238]_ ;
  assign \new_[93243]_  = \new_[93242]_  & \new_[93235]_ ;
  assign \new_[93246]_  = ~A267 & A266;
  assign \new_[93249]_  = A269 & ~A268;
  assign \new_[93250]_  = \new_[93249]_  & \new_[93246]_ ;
  assign \new_[93253]_  = ~A299 & A298;
  assign \new_[93256]_  = A301 & A300;
  assign \new_[93257]_  = \new_[93256]_  & \new_[93253]_ ;
  assign \new_[93258]_  = \new_[93257]_  & \new_[93250]_ ;
  assign \new_[93261]_  = A166 & A167;
  assign \new_[93264]_  = A200 & ~A199;
  assign \new_[93265]_  = \new_[93264]_  & \new_[93261]_ ;
  assign \new_[93268]_  = ~A202 & ~A201;
  assign \new_[93271]_  = ~A265 & A203;
  assign \new_[93272]_  = \new_[93271]_  & \new_[93268]_ ;
  assign \new_[93273]_  = \new_[93272]_  & \new_[93265]_ ;
  assign \new_[93276]_  = ~A267 & A266;
  assign \new_[93279]_  = A269 & ~A268;
  assign \new_[93280]_  = \new_[93279]_  & \new_[93276]_ ;
  assign \new_[93283]_  = ~A299 & A298;
  assign \new_[93286]_  = ~A302 & A300;
  assign \new_[93287]_  = \new_[93286]_  & \new_[93283]_ ;
  assign \new_[93288]_  = \new_[93287]_  & \new_[93280]_ ;
  assign \new_[93291]_  = A166 & A167;
  assign \new_[93294]_  = A200 & ~A199;
  assign \new_[93295]_  = \new_[93294]_  & \new_[93291]_ ;
  assign \new_[93298]_  = ~A202 & ~A201;
  assign \new_[93301]_  = ~A265 & A203;
  assign \new_[93302]_  = \new_[93301]_  & \new_[93298]_ ;
  assign \new_[93303]_  = \new_[93302]_  & \new_[93295]_ ;
  assign \new_[93306]_  = ~A267 & A266;
  assign \new_[93309]_  = A269 & ~A268;
  assign \new_[93310]_  = \new_[93309]_  & \new_[93306]_ ;
  assign \new_[93313]_  = A299 & ~A298;
  assign \new_[93316]_  = A301 & A300;
  assign \new_[93317]_  = \new_[93316]_  & \new_[93313]_ ;
  assign \new_[93318]_  = \new_[93317]_  & \new_[93310]_ ;
  assign \new_[93321]_  = A166 & A167;
  assign \new_[93324]_  = A200 & ~A199;
  assign \new_[93325]_  = \new_[93324]_  & \new_[93321]_ ;
  assign \new_[93328]_  = ~A202 & ~A201;
  assign \new_[93331]_  = ~A265 & A203;
  assign \new_[93332]_  = \new_[93331]_  & \new_[93328]_ ;
  assign \new_[93333]_  = \new_[93332]_  & \new_[93325]_ ;
  assign \new_[93336]_  = ~A267 & A266;
  assign \new_[93339]_  = A269 & ~A268;
  assign \new_[93340]_  = \new_[93339]_  & \new_[93336]_ ;
  assign \new_[93343]_  = A299 & ~A298;
  assign \new_[93346]_  = ~A302 & A300;
  assign \new_[93347]_  = \new_[93346]_  & \new_[93343]_ ;
  assign \new_[93348]_  = \new_[93347]_  & \new_[93340]_ ;
  assign \new_[93351]_  = A166 & A167;
  assign \new_[93354]_  = A200 & ~A199;
  assign \new_[93355]_  = \new_[93354]_  & \new_[93351]_ ;
  assign \new_[93358]_  = ~A202 & ~A201;
  assign \new_[93361]_  = A265 & A203;
  assign \new_[93362]_  = \new_[93361]_  & \new_[93358]_ ;
  assign \new_[93363]_  = \new_[93362]_  & \new_[93355]_ ;
  assign \new_[93366]_  = A267 & ~A266;
  assign \new_[93369]_  = A298 & A268;
  assign \new_[93370]_  = \new_[93369]_  & \new_[93366]_ ;
  assign \new_[93373]_  = ~A300 & ~A299;
  assign \new_[93376]_  = A302 & ~A301;
  assign \new_[93377]_  = \new_[93376]_  & \new_[93373]_ ;
  assign \new_[93378]_  = \new_[93377]_  & \new_[93370]_ ;
  assign \new_[93381]_  = A166 & A167;
  assign \new_[93384]_  = A200 & ~A199;
  assign \new_[93385]_  = \new_[93384]_  & \new_[93381]_ ;
  assign \new_[93388]_  = ~A202 & ~A201;
  assign \new_[93391]_  = A265 & A203;
  assign \new_[93392]_  = \new_[93391]_  & \new_[93388]_ ;
  assign \new_[93393]_  = \new_[93392]_  & \new_[93385]_ ;
  assign \new_[93396]_  = A267 & ~A266;
  assign \new_[93399]_  = ~A298 & A268;
  assign \new_[93400]_  = \new_[93399]_  & \new_[93396]_ ;
  assign \new_[93403]_  = ~A300 & A299;
  assign \new_[93406]_  = A302 & ~A301;
  assign \new_[93407]_  = \new_[93406]_  & \new_[93403]_ ;
  assign \new_[93408]_  = \new_[93407]_  & \new_[93400]_ ;
  assign \new_[93411]_  = A166 & A167;
  assign \new_[93414]_  = A200 & ~A199;
  assign \new_[93415]_  = \new_[93414]_  & \new_[93411]_ ;
  assign \new_[93418]_  = ~A202 & ~A201;
  assign \new_[93421]_  = A265 & A203;
  assign \new_[93422]_  = \new_[93421]_  & \new_[93418]_ ;
  assign \new_[93423]_  = \new_[93422]_  & \new_[93415]_ ;
  assign \new_[93426]_  = A267 & ~A266;
  assign \new_[93429]_  = A298 & ~A269;
  assign \new_[93430]_  = \new_[93429]_  & \new_[93426]_ ;
  assign \new_[93433]_  = ~A300 & ~A299;
  assign \new_[93436]_  = A302 & ~A301;
  assign \new_[93437]_  = \new_[93436]_  & \new_[93433]_ ;
  assign \new_[93438]_  = \new_[93437]_  & \new_[93430]_ ;
  assign \new_[93441]_  = A166 & A167;
  assign \new_[93444]_  = A200 & ~A199;
  assign \new_[93445]_  = \new_[93444]_  & \new_[93441]_ ;
  assign \new_[93448]_  = ~A202 & ~A201;
  assign \new_[93451]_  = A265 & A203;
  assign \new_[93452]_  = \new_[93451]_  & \new_[93448]_ ;
  assign \new_[93453]_  = \new_[93452]_  & \new_[93445]_ ;
  assign \new_[93456]_  = A267 & ~A266;
  assign \new_[93459]_  = ~A298 & ~A269;
  assign \new_[93460]_  = \new_[93459]_  & \new_[93456]_ ;
  assign \new_[93463]_  = ~A300 & A299;
  assign \new_[93466]_  = A302 & ~A301;
  assign \new_[93467]_  = \new_[93466]_  & \new_[93463]_ ;
  assign \new_[93468]_  = \new_[93467]_  & \new_[93460]_ ;
  assign \new_[93471]_  = A166 & A167;
  assign \new_[93474]_  = A200 & ~A199;
  assign \new_[93475]_  = \new_[93474]_  & \new_[93471]_ ;
  assign \new_[93478]_  = ~A202 & ~A201;
  assign \new_[93481]_  = A265 & A203;
  assign \new_[93482]_  = \new_[93481]_  & \new_[93478]_ ;
  assign \new_[93483]_  = \new_[93482]_  & \new_[93475]_ ;
  assign \new_[93486]_  = ~A267 & ~A266;
  assign \new_[93489]_  = A269 & ~A268;
  assign \new_[93490]_  = \new_[93489]_  & \new_[93486]_ ;
  assign \new_[93493]_  = ~A299 & A298;
  assign \new_[93496]_  = A301 & A300;
  assign \new_[93497]_  = \new_[93496]_  & \new_[93493]_ ;
  assign \new_[93498]_  = \new_[93497]_  & \new_[93490]_ ;
  assign \new_[93501]_  = A166 & A167;
  assign \new_[93504]_  = A200 & ~A199;
  assign \new_[93505]_  = \new_[93504]_  & \new_[93501]_ ;
  assign \new_[93508]_  = ~A202 & ~A201;
  assign \new_[93511]_  = A265 & A203;
  assign \new_[93512]_  = \new_[93511]_  & \new_[93508]_ ;
  assign \new_[93513]_  = \new_[93512]_  & \new_[93505]_ ;
  assign \new_[93516]_  = ~A267 & ~A266;
  assign \new_[93519]_  = A269 & ~A268;
  assign \new_[93520]_  = \new_[93519]_  & \new_[93516]_ ;
  assign \new_[93523]_  = ~A299 & A298;
  assign \new_[93526]_  = ~A302 & A300;
  assign \new_[93527]_  = \new_[93526]_  & \new_[93523]_ ;
  assign \new_[93528]_  = \new_[93527]_  & \new_[93520]_ ;
  assign \new_[93531]_  = A166 & A167;
  assign \new_[93534]_  = A200 & ~A199;
  assign \new_[93535]_  = \new_[93534]_  & \new_[93531]_ ;
  assign \new_[93538]_  = ~A202 & ~A201;
  assign \new_[93541]_  = A265 & A203;
  assign \new_[93542]_  = \new_[93541]_  & \new_[93538]_ ;
  assign \new_[93543]_  = \new_[93542]_  & \new_[93535]_ ;
  assign \new_[93546]_  = ~A267 & ~A266;
  assign \new_[93549]_  = A269 & ~A268;
  assign \new_[93550]_  = \new_[93549]_  & \new_[93546]_ ;
  assign \new_[93553]_  = A299 & ~A298;
  assign \new_[93556]_  = A301 & A300;
  assign \new_[93557]_  = \new_[93556]_  & \new_[93553]_ ;
  assign \new_[93558]_  = \new_[93557]_  & \new_[93550]_ ;
  assign \new_[93561]_  = A166 & A167;
  assign \new_[93564]_  = A200 & ~A199;
  assign \new_[93565]_  = \new_[93564]_  & \new_[93561]_ ;
  assign \new_[93568]_  = ~A202 & ~A201;
  assign \new_[93571]_  = A265 & A203;
  assign \new_[93572]_  = \new_[93571]_  & \new_[93568]_ ;
  assign \new_[93573]_  = \new_[93572]_  & \new_[93565]_ ;
  assign \new_[93576]_  = ~A267 & ~A266;
  assign \new_[93579]_  = A269 & ~A268;
  assign \new_[93580]_  = \new_[93579]_  & \new_[93576]_ ;
  assign \new_[93583]_  = A299 & ~A298;
  assign \new_[93586]_  = ~A302 & A300;
  assign \new_[93587]_  = \new_[93586]_  & \new_[93583]_ ;
  assign \new_[93588]_  = \new_[93587]_  & \new_[93580]_ ;
  assign \new_[93591]_  = A166 & A167;
  assign \new_[93594]_  = ~A200 & A199;
  assign \new_[93595]_  = \new_[93594]_  & \new_[93591]_ ;
  assign \new_[93598]_  = A202 & A201;
  assign \new_[93601]_  = A266 & ~A265;
  assign \new_[93602]_  = \new_[93601]_  & \new_[93598]_ ;
  assign \new_[93603]_  = \new_[93602]_  & \new_[93595]_ ;
  assign \new_[93606]_  = ~A268 & ~A267;
  assign \new_[93609]_  = A298 & A269;
  assign \new_[93610]_  = \new_[93609]_  & \new_[93606]_ ;
  assign \new_[93613]_  = ~A300 & ~A299;
  assign \new_[93616]_  = A302 & ~A301;
  assign \new_[93617]_  = \new_[93616]_  & \new_[93613]_ ;
  assign \new_[93618]_  = \new_[93617]_  & \new_[93610]_ ;
  assign \new_[93621]_  = A166 & A167;
  assign \new_[93624]_  = ~A200 & A199;
  assign \new_[93625]_  = \new_[93624]_  & \new_[93621]_ ;
  assign \new_[93628]_  = A202 & A201;
  assign \new_[93631]_  = A266 & ~A265;
  assign \new_[93632]_  = \new_[93631]_  & \new_[93628]_ ;
  assign \new_[93633]_  = \new_[93632]_  & \new_[93625]_ ;
  assign \new_[93636]_  = ~A268 & ~A267;
  assign \new_[93639]_  = ~A298 & A269;
  assign \new_[93640]_  = \new_[93639]_  & \new_[93636]_ ;
  assign \new_[93643]_  = ~A300 & A299;
  assign \new_[93646]_  = A302 & ~A301;
  assign \new_[93647]_  = \new_[93646]_  & \new_[93643]_ ;
  assign \new_[93648]_  = \new_[93647]_  & \new_[93640]_ ;
  assign \new_[93651]_  = A166 & A167;
  assign \new_[93654]_  = ~A200 & A199;
  assign \new_[93655]_  = \new_[93654]_  & \new_[93651]_ ;
  assign \new_[93658]_  = A202 & A201;
  assign \new_[93661]_  = ~A266 & A265;
  assign \new_[93662]_  = \new_[93661]_  & \new_[93658]_ ;
  assign \new_[93663]_  = \new_[93662]_  & \new_[93655]_ ;
  assign \new_[93666]_  = ~A268 & ~A267;
  assign \new_[93669]_  = A298 & A269;
  assign \new_[93670]_  = \new_[93669]_  & \new_[93666]_ ;
  assign \new_[93673]_  = ~A300 & ~A299;
  assign \new_[93676]_  = A302 & ~A301;
  assign \new_[93677]_  = \new_[93676]_  & \new_[93673]_ ;
  assign \new_[93678]_  = \new_[93677]_  & \new_[93670]_ ;
  assign \new_[93681]_  = A166 & A167;
  assign \new_[93684]_  = ~A200 & A199;
  assign \new_[93685]_  = \new_[93684]_  & \new_[93681]_ ;
  assign \new_[93688]_  = A202 & A201;
  assign \new_[93691]_  = ~A266 & A265;
  assign \new_[93692]_  = \new_[93691]_  & \new_[93688]_ ;
  assign \new_[93693]_  = \new_[93692]_  & \new_[93685]_ ;
  assign \new_[93696]_  = ~A268 & ~A267;
  assign \new_[93699]_  = ~A298 & A269;
  assign \new_[93700]_  = \new_[93699]_  & \new_[93696]_ ;
  assign \new_[93703]_  = ~A300 & A299;
  assign \new_[93706]_  = A302 & ~A301;
  assign \new_[93707]_  = \new_[93706]_  & \new_[93703]_ ;
  assign \new_[93708]_  = \new_[93707]_  & \new_[93700]_ ;
  assign \new_[93711]_  = A166 & A167;
  assign \new_[93714]_  = ~A200 & A199;
  assign \new_[93715]_  = \new_[93714]_  & \new_[93711]_ ;
  assign \new_[93718]_  = ~A203 & A201;
  assign \new_[93721]_  = A266 & ~A265;
  assign \new_[93722]_  = \new_[93721]_  & \new_[93718]_ ;
  assign \new_[93723]_  = \new_[93722]_  & \new_[93715]_ ;
  assign \new_[93726]_  = ~A268 & ~A267;
  assign \new_[93729]_  = A298 & A269;
  assign \new_[93730]_  = \new_[93729]_  & \new_[93726]_ ;
  assign \new_[93733]_  = ~A300 & ~A299;
  assign \new_[93736]_  = A302 & ~A301;
  assign \new_[93737]_  = \new_[93736]_  & \new_[93733]_ ;
  assign \new_[93738]_  = \new_[93737]_  & \new_[93730]_ ;
  assign \new_[93741]_  = A166 & A167;
  assign \new_[93744]_  = ~A200 & A199;
  assign \new_[93745]_  = \new_[93744]_  & \new_[93741]_ ;
  assign \new_[93748]_  = ~A203 & A201;
  assign \new_[93751]_  = A266 & ~A265;
  assign \new_[93752]_  = \new_[93751]_  & \new_[93748]_ ;
  assign \new_[93753]_  = \new_[93752]_  & \new_[93745]_ ;
  assign \new_[93756]_  = ~A268 & ~A267;
  assign \new_[93759]_  = ~A298 & A269;
  assign \new_[93760]_  = \new_[93759]_  & \new_[93756]_ ;
  assign \new_[93763]_  = ~A300 & A299;
  assign \new_[93766]_  = A302 & ~A301;
  assign \new_[93767]_  = \new_[93766]_  & \new_[93763]_ ;
  assign \new_[93768]_  = \new_[93767]_  & \new_[93760]_ ;
  assign \new_[93771]_  = A166 & A167;
  assign \new_[93774]_  = ~A200 & A199;
  assign \new_[93775]_  = \new_[93774]_  & \new_[93771]_ ;
  assign \new_[93778]_  = ~A203 & A201;
  assign \new_[93781]_  = ~A266 & A265;
  assign \new_[93782]_  = \new_[93781]_  & \new_[93778]_ ;
  assign \new_[93783]_  = \new_[93782]_  & \new_[93775]_ ;
  assign \new_[93786]_  = ~A268 & ~A267;
  assign \new_[93789]_  = A298 & A269;
  assign \new_[93790]_  = \new_[93789]_  & \new_[93786]_ ;
  assign \new_[93793]_  = ~A300 & ~A299;
  assign \new_[93796]_  = A302 & ~A301;
  assign \new_[93797]_  = \new_[93796]_  & \new_[93793]_ ;
  assign \new_[93798]_  = \new_[93797]_  & \new_[93790]_ ;
  assign \new_[93801]_  = A166 & A167;
  assign \new_[93804]_  = ~A200 & A199;
  assign \new_[93805]_  = \new_[93804]_  & \new_[93801]_ ;
  assign \new_[93808]_  = ~A203 & A201;
  assign \new_[93811]_  = ~A266 & A265;
  assign \new_[93812]_  = \new_[93811]_  & \new_[93808]_ ;
  assign \new_[93813]_  = \new_[93812]_  & \new_[93805]_ ;
  assign \new_[93816]_  = ~A268 & ~A267;
  assign \new_[93819]_  = ~A298 & A269;
  assign \new_[93820]_  = \new_[93819]_  & \new_[93816]_ ;
  assign \new_[93823]_  = ~A300 & A299;
  assign \new_[93826]_  = A302 & ~A301;
  assign \new_[93827]_  = \new_[93826]_  & \new_[93823]_ ;
  assign \new_[93828]_  = \new_[93827]_  & \new_[93820]_ ;
  assign \new_[93831]_  = A166 & A167;
  assign \new_[93834]_  = ~A200 & A199;
  assign \new_[93835]_  = \new_[93834]_  & \new_[93831]_ ;
  assign \new_[93838]_  = ~A202 & ~A201;
  assign \new_[93841]_  = ~A265 & A203;
  assign \new_[93842]_  = \new_[93841]_  & \new_[93838]_ ;
  assign \new_[93843]_  = \new_[93842]_  & \new_[93835]_ ;
  assign \new_[93846]_  = A267 & A266;
  assign \new_[93849]_  = A298 & A268;
  assign \new_[93850]_  = \new_[93849]_  & \new_[93846]_ ;
  assign \new_[93853]_  = ~A300 & ~A299;
  assign \new_[93856]_  = A302 & ~A301;
  assign \new_[93857]_  = \new_[93856]_  & \new_[93853]_ ;
  assign \new_[93858]_  = \new_[93857]_  & \new_[93850]_ ;
  assign \new_[93861]_  = A166 & A167;
  assign \new_[93864]_  = ~A200 & A199;
  assign \new_[93865]_  = \new_[93864]_  & \new_[93861]_ ;
  assign \new_[93868]_  = ~A202 & ~A201;
  assign \new_[93871]_  = ~A265 & A203;
  assign \new_[93872]_  = \new_[93871]_  & \new_[93868]_ ;
  assign \new_[93873]_  = \new_[93872]_  & \new_[93865]_ ;
  assign \new_[93876]_  = A267 & A266;
  assign \new_[93879]_  = ~A298 & A268;
  assign \new_[93880]_  = \new_[93879]_  & \new_[93876]_ ;
  assign \new_[93883]_  = ~A300 & A299;
  assign \new_[93886]_  = A302 & ~A301;
  assign \new_[93887]_  = \new_[93886]_  & \new_[93883]_ ;
  assign \new_[93888]_  = \new_[93887]_  & \new_[93880]_ ;
  assign \new_[93891]_  = A166 & A167;
  assign \new_[93894]_  = ~A200 & A199;
  assign \new_[93895]_  = \new_[93894]_  & \new_[93891]_ ;
  assign \new_[93898]_  = ~A202 & ~A201;
  assign \new_[93901]_  = ~A265 & A203;
  assign \new_[93902]_  = \new_[93901]_  & \new_[93898]_ ;
  assign \new_[93903]_  = \new_[93902]_  & \new_[93895]_ ;
  assign \new_[93906]_  = A267 & A266;
  assign \new_[93909]_  = A298 & ~A269;
  assign \new_[93910]_  = \new_[93909]_  & \new_[93906]_ ;
  assign \new_[93913]_  = ~A300 & ~A299;
  assign \new_[93916]_  = A302 & ~A301;
  assign \new_[93917]_  = \new_[93916]_  & \new_[93913]_ ;
  assign \new_[93918]_  = \new_[93917]_  & \new_[93910]_ ;
  assign \new_[93921]_  = A166 & A167;
  assign \new_[93924]_  = ~A200 & A199;
  assign \new_[93925]_  = \new_[93924]_  & \new_[93921]_ ;
  assign \new_[93928]_  = ~A202 & ~A201;
  assign \new_[93931]_  = ~A265 & A203;
  assign \new_[93932]_  = \new_[93931]_  & \new_[93928]_ ;
  assign \new_[93933]_  = \new_[93932]_  & \new_[93925]_ ;
  assign \new_[93936]_  = A267 & A266;
  assign \new_[93939]_  = ~A298 & ~A269;
  assign \new_[93940]_  = \new_[93939]_  & \new_[93936]_ ;
  assign \new_[93943]_  = ~A300 & A299;
  assign \new_[93946]_  = A302 & ~A301;
  assign \new_[93947]_  = \new_[93946]_  & \new_[93943]_ ;
  assign \new_[93948]_  = \new_[93947]_  & \new_[93940]_ ;
  assign \new_[93951]_  = A166 & A167;
  assign \new_[93954]_  = ~A200 & A199;
  assign \new_[93955]_  = \new_[93954]_  & \new_[93951]_ ;
  assign \new_[93958]_  = ~A202 & ~A201;
  assign \new_[93961]_  = ~A265 & A203;
  assign \new_[93962]_  = \new_[93961]_  & \new_[93958]_ ;
  assign \new_[93963]_  = \new_[93962]_  & \new_[93955]_ ;
  assign \new_[93966]_  = ~A267 & A266;
  assign \new_[93969]_  = A269 & ~A268;
  assign \new_[93970]_  = \new_[93969]_  & \new_[93966]_ ;
  assign \new_[93973]_  = ~A299 & A298;
  assign \new_[93976]_  = A301 & A300;
  assign \new_[93977]_  = \new_[93976]_  & \new_[93973]_ ;
  assign \new_[93978]_  = \new_[93977]_  & \new_[93970]_ ;
  assign \new_[93981]_  = A166 & A167;
  assign \new_[93984]_  = ~A200 & A199;
  assign \new_[93985]_  = \new_[93984]_  & \new_[93981]_ ;
  assign \new_[93988]_  = ~A202 & ~A201;
  assign \new_[93991]_  = ~A265 & A203;
  assign \new_[93992]_  = \new_[93991]_  & \new_[93988]_ ;
  assign \new_[93993]_  = \new_[93992]_  & \new_[93985]_ ;
  assign \new_[93996]_  = ~A267 & A266;
  assign \new_[93999]_  = A269 & ~A268;
  assign \new_[94000]_  = \new_[93999]_  & \new_[93996]_ ;
  assign \new_[94003]_  = ~A299 & A298;
  assign \new_[94006]_  = ~A302 & A300;
  assign \new_[94007]_  = \new_[94006]_  & \new_[94003]_ ;
  assign \new_[94008]_  = \new_[94007]_  & \new_[94000]_ ;
  assign \new_[94011]_  = A166 & A167;
  assign \new_[94014]_  = ~A200 & A199;
  assign \new_[94015]_  = \new_[94014]_  & \new_[94011]_ ;
  assign \new_[94018]_  = ~A202 & ~A201;
  assign \new_[94021]_  = ~A265 & A203;
  assign \new_[94022]_  = \new_[94021]_  & \new_[94018]_ ;
  assign \new_[94023]_  = \new_[94022]_  & \new_[94015]_ ;
  assign \new_[94026]_  = ~A267 & A266;
  assign \new_[94029]_  = A269 & ~A268;
  assign \new_[94030]_  = \new_[94029]_  & \new_[94026]_ ;
  assign \new_[94033]_  = A299 & ~A298;
  assign \new_[94036]_  = A301 & A300;
  assign \new_[94037]_  = \new_[94036]_  & \new_[94033]_ ;
  assign \new_[94038]_  = \new_[94037]_  & \new_[94030]_ ;
  assign \new_[94041]_  = A166 & A167;
  assign \new_[94044]_  = ~A200 & A199;
  assign \new_[94045]_  = \new_[94044]_  & \new_[94041]_ ;
  assign \new_[94048]_  = ~A202 & ~A201;
  assign \new_[94051]_  = ~A265 & A203;
  assign \new_[94052]_  = \new_[94051]_  & \new_[94048]_ ;
  assign \new_[94053]_  = \new_[94052]_  & \new_[94045]_ ;
  assign \new_[94056]_  = ~A267 & A266;
  assign \new_[94059]_  = A269 & ~A268;
  assign \new_[94060]_  = \new_[94059]_  & \new_[94056]_ ;
  assign \new_[94063]_  = A299 & ~A298;
  assign \new_[94066]_  = ~A302 & A300;
  assign \new_[94067]_  = \new_[94066]_  & \new_[94063]_ ;
  assign \new_[94068]_  = \new_[94067]_  & \new_[94060]_ ;
  assign \new_[94071]_  = A166 & A167;
  assign \new_[94074]_  = ~A200 & A199;
  assign \new_[94075]_  = \new_[94074]_  & \new_[94071]_ ;
  assign \new_[94078]_  = ~A202 & ~A201;
  assign \new_[94081]_  = A265 & A203;
  assign \new_[94082]_  = \new_[94081]_  & \new_[94078]_ ;
  assign \new_[94083]_  = \new_[94082]_  & \new_[94075]_ ;
  assign \new_[94086]_  = A267 & ~A266;
  assign \new_[94089]_  = A298 & A268;
  assign \new_[94090]_  = \new_[94089]_  & \new_[94086]_ ;
  assign \new_[94093]_  = ~A300 & ~A299;
  assign \new_[94096]_  = A302 & ~A301;
  assign \new_[94097]_  = \new_[94096]_  & \new_[94093]_ ;
  assign \new_[94098]_  = \new_[94097]_  & \new_[94090]_ ;
  assign \new_[94101]_  = A166 & A167;
  assign \new_[94104]_  = ~A200 & A199;
  assign \new_[94105]_  = \new_[94104]_  & \new_[94101]_ ;
  assign \new_[94108]_  = ~A202 & ~A201;
  assign \new_[94111]_  = A265 & A203;
  assign \new_[94112]_  = \new_[94111]_  & \new_[94108]_ ;
  assign \new_[94113]_  = \new_[94112]_  & \new_[94105]_ ;
  assign \new_[94116]_  = A267 & ~A266;
  assign \new_[94119]_  = ~A298 & A268;
  assign \new_[94120]_  = \new_[94119]_  & \new_[94116]_ ;
  assign \new_[94123]_  = ~A300 & A299;
  assign \new_[94126]_  = A302 & ~A301;
  assign \new_[94127]_  = \new_[94126]_  & \new_[94123]_ ;
  assign \new_[94128]_  = \new_[94127]_  & \new_[94120]_ ;
  assign \new_[94131]_  = A166 & A167;
  assign \new_[94134]_  = ~A200 & A199;
  assign \new_[94135]_  = \new_[94134]_  & \new_[94131]_ ;
  assign \new_[94138]_  = ~A202 & ~A201;
  assign \new_[94141]_  = A265 & A203;
  assign \new_[94142]_  = \new_[94141]_  & \new_[94138]_ ;
  assign \new_[94143]_  = \new_[94142]_  & \new_[94135]_ ;
  assign \new_[94146]_  = A267 & ~A266;
  assign \new_[94149]_  = A298 & ~A269;
  assign \new_[94150]_  = \new_[94149]_  & \new_[94146]_ ;
  assign \new_[94153]_  = ~A300 & ~A299;
  assign \new_[94156]_  = A302 & ~A301;
  assign \new_[94157]_  = \new_[94156]_  & \new_[94153]_ ;
  assign \new_[94158]_  = \new_[94157]_  & \new_[94150]_ ;
  assign \new_[94161]_  = A166 & A167;
  assign \new_[94164]_  = ~A200 & A199;
  assign \new_[94165]_  = \new_[94164]_  & \new_[94161]_ ;
  assign \new_[94168]_  = ~A202 & ~A201;
  assign \new_[94171]_  = A265 & A203;
  assign \new_[94172]_  = \new_[94171]_  & \new_[94168]_ ;
  assign \new_[94173]_  = \new_[94172]_  & \new_[94165]_ ;
  assign \new_[94176]_  = A267 & ~A266;
  assign \new_[94179]_  = ~A298 & ~A269;
  assign \new_[94180]_  = \new_[94179]_  & \new_[94176]_ ;
  assign \new_[94183]_  = ~A300 & A299;
  assign \new_[94186]_  = A302 & ~A301;
  assign \new_[94187]_  = \new_[94186]_  & \new_[94183]_ ;
  assign \new_[94188]_  = \new_[94187]_  & \new_[94180]_ ;
  assign \new_[94191]_  = A166 & A167;
  assign \new_[94194]_  = ~A200 & A199;
  assign \new_[94195]_  = \new_[94194]_  & \new_[94191]_ ;
  assign \new_[94198]_  = ~A202 & ~A201;
  assign \new_[94201]_  = A265 & A203;
  assign \new_[94202]_  = \new_[94201]_  & \new_[94198]_ ;
  assign \new_[94203]_  = \new_[94202]_  & \new_[94195]_ ;
  assign \new_[94206]_  = ~A267 & ~A266;
  assign \new_[94209]_  = A269 & ~A268;
  assign \new_[94210]_  = \new_[94209]_  & \new_[94206]_ ;
  assign \new_[94213]_  = ~A299 & A298;
  assign \new_[94216]_  = A301 & A300;
  assign \new_[94217]_  = \new_[94216]_  & \new_[94213]_ ;
  assign \new_[94218]_  = \new_[94217]_  & \new_[94210]_ ;
  assign \new_[94221]_  = A166 & A167;
  assign \new_[94224]_  = ~A200 & A199;
  assign \new_[94225]_  = \new_[94224]_  & \new_[94221]_ ;
  assign \new_[94228]_  = ~A202 & ~A201;
  assign \new_[94231]_  = A265 & A203;
  assign \new_[94232]_  = \new_[94231]_  & \new_[94228]_ ;
  assign \new_[94233]_  = \new_[94232]_  & \new_[94225]_ ;
  assign \new_[94236]_  = ~A267 & ~A266;
  assign \new_[94239]_  = A269 & ~A268;
  assign \new_[94240]_  = \new_[94239]_  & \new_[94236]_ ;
  assign \new_[94243]_  = ~A299 & A298;
  assign \new_[94246]_  = ~A302 & A300;
  assign \new_[94247]_  = \new_[94246]_  & \new_[94243]_ ;
  assign \new_[94248]_  = \new_[94247]_  & \new_[94240]_ ;
  assign \new_[94251]_  = A166 & A167;
  assign \new_[94254]_  = ~A200 & A199;
  assign \new_[94255]_  = \new_[94254]_  & \new_[94251]_ ;
  assign \new_[94258]_  = ~A202 & ~A201;
  assign \new_[94261]_  = A265 & A203;
  assign \new_[94262]_  = \new_[94261]_  & \new_[94258]_ ;
  assign \new_[94263]_  = \new_[94262]_  & \new_[94255]_ ;
  assign \new_[94266]_  = ~A267 & ~A266;
  assign \new_[94269]_  = A269 & ~A268;
  assign \new_[94270]_  = \new_[94269]_  & \new_[94266]_ ;
  assign \new_[94273]_  = A299 & ~A298;
  assign \new_[94276]_  = A301 & A300;
  assign \new_[94277]_  = \new_[94276]_  & \new_[94273]_ ;
  assign \new_[94278]_  = \new_[94277]_  & \new_[94270]_ ;
  assign \new_[94281]_  = A166 & A167;
  assign \new_[94284]_  = ~A200 & A199;
  assign \new_[94285]_  = \new_[94284]_  & \new_[94281]_ ;
  assign \new_[94288]_  = ~A202 & ~A201;
  assign \new_[94291]_  = A265 & A203;
  assign \new_[94292]_  = \new_[94291]_  & \new_[94288]_ ;
  assign \new_[94293]_  = \new_[94292]_  & \new_[94285]_ ;
  assign \new_[94296]_  = ~A267 & ~A266;
  assign \new_[94299]_  = A269 & ~A268;
  assign \new_[94300]_  = \new_[94299]_  & \new_[94296]_ ;
  assign \new_[94303]_  = A299 & ~A298;
  assign \new_[94306]_  = ~A302 & A300;
  assign \new_[94307]_  = \new_[94306]_  & \new_[94303]_ ;
  assign \new_[94308]_  = \new_[94307]_  & \new_[94300]_ ;
  assign \new_[94311]_  = ~A166 & ~A167;
  assign \new_[94314]_  = A200 & ~A199;
  assign \new_[94315]_  = \new_[94314]_  & \new_[94311]_ ;
  assign \new_[94318]_  = A202 & A201;
  assign \new_[94321]_  = A266 & ~A265;
  assign \new_[94322]_  = \new_[94321]_  & \new_[94318]_ ;
  assign \new_[94323]_  = \new_[94322]_  & \new_[94315]_ ;
  assign \new_[94326]_  = ~A268 & ~A267;
  assign \new_[94329]_  = A298 & A269;
  assign \new_[94330]_  = \new_[94329]_  & \new_[94326]_ ;
  assign \new_[94333]_  = ~A300 & ~A299;
  assign \new_[94336]_  = A302 & ~A301;
  assign \new_[94337]_  = \new_[94336]_  & \new_[94333]_ ;
  assign \new_[94338]_  = \new_[94337]_  & \new_[94330]_ ;
  assign \new_[94341]_  = ~A166 & ~A167;
  assign \new_[94344]_  = A200 & ~A199;
  assign \new_[94345]_  = \new_[94344]_  & \new_[94341]_ ;
  assign \new_[94348]_  = A202 & A201;
  assign \new_[94351]_  = A266 & ~A265;
  assign \new_[94352]_  = \new_[94351]_  & \new_[94348]_ ;
  assign \new_[94353]_  = \new_[94352]_  & \new_[94345]_ ;
  assign \new_[94356]_  = ~A268 & ~A267;
  assign \new_[94359]_  = ~A298 & A269;
  assign \new_[94360]_  = \new_[94359]_  & \new_[94356]_ ;
  assign \new_[94363]_  = ~A300 & A299;
  assign \new_[94366]_  = A302 & ~A301;
  assign \new_[94367]_  = \new_[94366]_  & \new_[94363]_ ;
  assign \new_[94368]_  = \new_[94367]_  & \new_[94360]_ ;
  assign \new_[94371]_  = ~A166 & ~A167;
  assign \new_[94374]_  = A200 & ~A199;
  assign \new_[94375]_  = \new_[94374]_  & \new_[94371]_ ;
  assign \new_[94378]_  = A202 & A201;
  assign \new_[94381]_  = ~A266 & A265;
  assign \new_[94382]_  = \new_[94381]_  & \new_[94378]_ ;
  assign \new_[94383]_  = \new_[94382]_  & \new_[94375]_ ;
  assign \new_[94386]_  = ~A268 & ~A267;
  assign \new_[94389]_  = A298 & A269;
  assign \new_[94390]_  = \new_[94389]_  & \new_[94386]_ ;
  assign \new_[94393]_  = ~A300 & ~A299;
  assign \new_[94396]_  = A302 & ~A301;
  assign \new_[94397]_  = \new_[94396]_  & \new_[94393]_ ;
  assign \new_[94398]_  = \new_[94397]_  & \new_[94390]_ ;
  assign \new_[94401]_  = ~A166 & ~A167;
  assign \new_[94404]_  = A200 & ~A199;
  assign \new_[94405]_  = \new_[94404]_  & \new_[94401]_ ;
  assign \new_[94408]_  = A202 & A201;
  assign \new_[94411]_  = ~A266 & A265;
  assign \new_[94412]_  = \new_[94411]_  & \new_[94408]_ ;
  assign \new_[94413]_  = \new_[94412]_  & \new_[94405]_ ;
  assign \new_[94416]_  = ~A268 & ~A267;
  assign \new_[94419]_  = ~A298 & A269;
  assign \new_[94420]_  = \new_[94419]_  & \new_[94416]_ ;
  assign \new_[94423]_  = ~A300 & A299;
  assign \new_[94426]_  = A302 & ~A301;
  assign \new_[94427]_  = \new_[94426]_  & \new_[94423]_ ;
  assign \new_[94428]_  = \new_[94427]_  & \new_[94420]_ ;
  assign \new_[94431]_  = ~A166 & ~A167;
  assign \new_[94434]_  = A200 & ~A199;
  assign \new_[94435]_  = \new_[94434]_  & \new_[94431]_ ;
  assign \new_[94438]_  = ~A203 & A201;
  assign \new_[94441]_  = A266 & ~A265;
  assign \new_[94442]_  = \new_[94441]_  & \new_[94438]_ ;
  assign \new_[94443]_  = \new_[94442]_  & \new_[94435]_ ;
  assign \new_[94446]_  = ~A268 & ~A267;
  assign \new_[94449]_  = A298 & A269;
  assign \new_[94450]_  = \new_[94449]_  & \new_[94446]_ ;
  assign \new_[94453]_  = ~A300 & ~A299;
  assign \new_[94456]_  = A302 & ~A301;
  assign \new_[94457]_  = \new_[94456]_  & \new_[94453]_ ;
  assign \new_[94458]_  = \new_[94457]_  & \new_[94450]_ ;
  assign \new_[94461]_  = ~A166 & ~A167;
  assign \new_[94464]_  = A200 & ~A199;
  assign \new_[94465]_  = \new_[94464]_  & \new_[94461]_ ;
  assign \new_[94468]_  = ~A203 & A201;
  assign \new_[94471]_  = A266 & ~A265;
  assign \new_[94472]_  = \new_[94471]_  & \new_[94468]_ ;
  assign \new_[94473]_  = \new_[94472]_  & \new_[94465]_ ;
  assign \new_[94476]_  = ~A268 & ~A267;
  assign \new_[94479]_  = ~A298 & A269;
  assign \new_[94480]_  = \new_[94479]_  & \new_[94476]_ ;
  assign \new_[94483]_  = ~A300 & A299;
  assign \new_[94486]_  = A302 & ~A301;
  assign \new_[94487]_  = \new_[94486]_  & \new_[94483]_ ;
  assign \new_[94488]_  = \new_[94487]_  & \new_[94480]_ ;
  assign \new_[94491]_  = ~A166 & ~A167;
  assign \new_[94494]_  = A200 & ~A199;
  assign \new_[94495]_  = \new_[94494]_  & \new_[94491]_ ;
  assign \new_[94498]_  = ~A203 & A201;
  assign \new_[94501]_  = ~A266 & A265;
  assign \new_[94502]_  = \new_[94501]_  & \new_[94498]_ ;
  assign \new_[94503]_  = \new_[94502]_  & \new_[94495]_ ;
  assign \new_[94506]_  = ~A268 & ~A267;
  assign \new_[94509]_  = A298 & A269;
  assign \new_[94510]_  = \new_[94509]_  & \new_[94506]_ ;
  assign \new_[94513]_  = ~A300 & ~A299;
  assign \new_[94516]_  = A302 & ~A301;
  assign \new_[94517]_  = \new_[94516]_  & \new_[94513]_ ;
  assign \new_[94518]_  = \new_[94517]_  & \new_[94510]_ ;
  assign \new_[94521]_  = ~A166 & ~A167;
  assign \new_[94524]_  = A200 & ~A199;
  assign \new_[94525]_  = \new_[94524]_  & \new_[94521]_ ;
  assign \new_[94528]_  = ~A203 & A201;
  assign \new_[94531]_  = ~A266 & A265;
  assign \new_[94532]_  = \new_[94531]_  & \new_[94528]_ ;
  assign \new_[94533]_  = \new_[94532]_  & \new_[94525]_ ;
  assign \new_[94536]_  = ~A268 & ~A267;
  assign \new_[94539]_  = ~A298 & A269;
  assign \new_[94540]_  = \new_[94539]_  & \new_[94536]_ ;
  assign \new_[94543]_  = ~A300 & A299;
  assign \new_[94546]_  = A302 & ~A301;
  assign \new_[94547]_  = \new_[94546]_  & \new_[94543]_ ;
  assign \new_[94548]_  = \new_[94547]_  & \new_[94540]_ ;
  assign \new_[94551]_  = ~A166 & ~A167;
  assign \new_[94554]_  = A200 & ~A199;
  assign \new_[94555]_  = \new_[94554]_  & \new_[94551]_ ;
  assign \new_[94558]_  = ~A202 & ~A201;
  assign \new_[94561]_  = ~A265 & A203;
  assign \new_[94562]_  = \new_[94561]_  & \new_[94558]_ ;
  assign \new_[94563]_  = \new_[94562]_  & \new_[94555]_ ;
  assign \new_[94566]_  = A267 & A266;
  assign \new_[94569]_  = A298 & A268;
  assign \new_[94570]_  = \new_[94569]_  & \new_[94566]_ ;
  assign \new_[94573]_  = ~A300 & ~A299;
  assign \new_[94576]_  = A302 & ~A301;
  assign \new_[94577]_  = \new_[94576]_  & \new_[94573]_ ;
  assign \new_[94578]_  = \new_[94577]_  & \new_[94570]_ ;
  assign \new_[94581]_  = ~A166 & ~A167;
  assign \new_[94584]_  = A200 & ~A199;
  assign \new_[94585]_  = \new_[94584]_  & \new_[94581]_ ;
  assign \new_[94588]_  = ~A202 & ~A201;
  assign \new_[94591]_  = ~A265 & A203;
  assign \new_[94592]_  = \new_[94591]_  & \new_[94588]_ ;
  assign \new_[94593]_  = \new_[94592]_  & \new_[94585]_ ;
  assign \new_[94596]_  = A267 & A266;
  assign \new_[94599]_  = ~A298 & A268;
  assign \new_[94600]_  = \new_[94599]_  & \new_[94596]_ ;
  assign \new_[94603]_  = ~A300 & A299;
  assign \new_[94606]_  = A302 & ~A301;
  assign \new_[94607]_  = \new_[94606]_  & \new_[94603]_ ;
  assign \new_[94608]_  = \new_[94607]_  & \new_[94600]_ ;
  assign \new_[94611]_  = ~A166 & ~A167;
  assign \new_[94614]_  = A200 & ~A199;
  assign \new_[94615]_  = \new_[94614]_  & \new_[94611]_ ;
  assign \new_[94618]_  = ~A202 & ~A201;
  assign \new_[94621]_  = ~A265 & A203;
  assign \new_[94622]_  = \new_[94621]_  & \new_[94618]_ ;
  assign \new_[94623]_  = \new_[94622]_  & \new_[94615]_ ;
  assign \new_[94626]_  = A267 & A266;
  assign \new_[94629]_  = A298 & ~A269;
  assign \new_[94630]_  = \new_[94629]_  & \new_[94626]_ ;
  assign \new_[94633]_  = ~A300 & ~A299;
  assign \new_[94636]_  = A302 & ~A301;
  assign \new_[94637]_  = \new_[94636]_  & \new_[94633]_ ;
  assign \new_[94638]_  = \new_[94637]_  & \new_[94630]_ ;
  assign \new_[94641]_  = ~A166 & ~A167;
  assign \new_[94644]_  = A200 & ~A199;
  assign \new_[94645]_  = \new_[94644]_  & \new_[94641]_ ;
  assign \new_[94648]_  = ~A202 & ~A201;
  assign \new_[94651]_  = ~A265 & A203;
  assign \new_[94652]_  = \new_[94651]_  & \new_[94648]_ ;
  assign \new_[94653]_  = \new_[94652]_  & \new_[94645]_ ;
  assign \new_[94656]_  = A267 & A266;
  assign \new_[94659]_  = ~A298 & ~A269;
  assign \new_[94660]_  = \new_[94659]_  & \new_[94656]_ ;
  assign \new_[94663]_  = ~A300 & A299;
  assign \new_[94666]_  = A302 & ~A301;
  assign \new_[94667]_  = \new_[94666]_  & \new_[94663]_ ;
  assign \new_[94668]_  = \new_[94667]_  & \new_[94660]_ ;
  assign \new_[94671]_  = ~A166 & ~A167;
  assign \new_[94674]_  = A200 & ~A199;
  assign \new_[94675]_  = \new_[94674]_  & \new_[94671]_ ;
  assign \new_[94678]_  = ~A202 & ~A201;
  assign \new_[94681]_  = ~A265 & A203;
  assign \new_[94682]_  = \new_[94681]_  & \new_[94678]_ ;
  assign \new_[94683]_  = \new_[94682]_  & \new_[94675]_ ;
  assign \new_[94686]_  = ~A267 & A266;
  assign \new_[94689]_  = A269 & ~A268;
  assign \new_[94690]_  = \new_[94689]_  & \new_[94686]_ ;
  assign \new_[94693]_  = ~A299 & A298;
  assign \new_[94696]_  = A301 & A300;
  assign \new_[94697]_  = \new_[94696]_  & \new_[94693]_ ;
  assign \new_[94698]_  = \new_[94697]_  & \new_[94690]_ ;
  assign \new_[94701]_  = ~A166 & ~A167;
  assign \new_[94704]_  = A200 & ~A199;
  assign \new_[94705]_  = \new_[94704]_  & \new_[94701]_ ;
  assign \new_[94708]_  = ~A202 & ~A201;
  assign \new_[94711]_  = ~A265 & A203;
  assign \new_[94712]_  = \new_[94711]_  & \new_[94708]_ ;
  assign \new_[94713]_  = \new_[94712]_  & \new_[94705]_ ;
  assign \new_[94716]_  = ~A267 & A266;
  assign \new_[94719]_  = A269 & ~A268;
  assign \new_[94720]_  = \new_[94719]_  & \new_[94716]_ ;
  assign \new_[94723]_  = ~A299 & A298;
  assign \new_[94726]_  = ~A302 & A300;
  assign \new_[94727]_  = \new_[94726]_  & \new_[94723]_ ;
  assign \new_[94728]_  = \new_[94727]_  & \new_[94720]_ ;
  assign \new_[94731]_  = ~A166 & ~A167;
  assign \new_[94734]_  = A200 & ~A199;
  assign \new_[94735]_  = \new_[94734]_  & \new_[94731]_ ;
  assign \new_[94738]_  = ~A202 & ~A201;
  assign \new_[94741]_  = ~A265 & A203;
  assign \new_[94742]_  = \new_[94741]_  & \new_[94738]_ ;
  assign \new_[94743]_  = \new_[94742]_  & \new_[94735]_ ;
  assign \new_[94746]_  = ~A267 & A266;
  assign \new_[94749]_  = A269 & ~A268;
  assign \new_[94750]_  = \new_[94749]_  & \new_[94746]_ ;
  assign \new_[94753]_  = A299 & ~A298;
  assign \new_[94756]_  = A301 & A300;
  assign \new_[94757]_  = \new_[94756]_  & \new_[94753]_ ;
  assign \new_[94758]_  = \new_[94757]_  & \new_[94750]_ ;
  assign \new_[94761]_  = ~A166 & ~A167;
  assign \new_[94764]_  = A200 & ~A199;
  assign \new_[94765]_  = \new_[94764]_  & \new_[94761]_ ;
  assign \new_[94768]_  = ~A202 & ~A201;
  assign \new_[94771]_  = ~A265 & A203;
  assign \new_[94772]_  = \new_[94771]_  & \new_[94768]_ ;
  assign \new_[94773]_  = \new_[94772]_  & \new_[94765]_ ;
  assign \new_[94776]_  = ~A267 & A266;
  assign \new_[94779]_  = A269 & ~A268;
  assign \new_[94780]_  = \new_[94779]_  & \new_[94776]_ ;
  assign \new_[94783]_  = A299 & ~A298;
  assign \new_[94786]_  = ~A302 & A300;
  assign \new_[94787]_  = \new_[94786]_  & \new_[94783]_ ;
  assign \new_[94788]_  = \new_[94787]_  & \new_[94780]_ ;
  assign \new_[94791]_  = ~A166 & ~A167;
  assign \new_[94794]_  = A200 & ~A199;
  assign \new_[94795]_  = \new_[94794]_  & \new_[94791]_ ;
  assign \new_[94798]_  = ~A202 & ~A201;
  assign \new_[94801]_  = A265 & A203;
  assign \new_[94802]_  = \new_[94801]_  & \new_[94798]_ ;
  assign \new_[94803]_  = \new_[94802]_  & \new_[94795]_ ;
  assign \new_[94806]_  = A267 & ~A266;
  assign \new_[94809]_  = A298 & A268;
  assign \new_[94810]_  = \new_[94809]_  & \new_[94806]_ ;
  assign \new_[94813]_  = ~A300 & ~A299;
  assign \new_[94816]_  = A302 & ~A301;
  assign \new_[94817]_  = \new_[94816]_  & \new_[94813]_ ;
  assign \new_[94818]_  = \new_[94817]_  & \new_[94810]_ ;
  assign \new_[94821]_  = ~A166 & ~A167;
  assign \new_[94824]_  = A200 & ~A199;
  assign \new_[94825]_  = \new_[94824]_  & \new_[94821]_ ;
  assign \new_[94828]_  = ~A202 & ~A201;
  assign \new_[94831]_  = A265 & A203;
  assign \new_[94832]_  = \new_[94831]_  & \new_[94828]_ ;
  assign \new_[94833]_  = \new_[94832]_  & \new_[94825]_ ;
  assign \new_[94836]_  = A267 & ~A266;
  assign \new_[94839]_  = ~A298 & A268;
  assign \new_[94840]_  = \new_[94839]_  & \new_[94836]_ ;
  assign \new_[94843]_  = ~A300 & A299;
  assign \new_[94846]_  = A302 & ~A301;
  assign \new_[94847]_  = \new_[94846]_  & \new_[94843]_ ;
  assign \new_[94848]_  = \new_[94847]_  & \new_[94840]_ ;
  assign \new_[94851]_  = ~A166 & ~A167;
  assign \new_[94854]_  = A200 & ~A199;
  assign \new_[94855]_  = \new_[94854]_  & \new_[94851]_ ;
  assign \new_[94858]_  = ~A202 & ~A201;
  assign \new_[94861]_  = A265 & A203;
  assign \new_[94862]_  = \new_[94861]_  & \new_[94858]_ ;
  assign \new_[94863]_  = \new_[94862]_  & \new_[94855]_ ;
  assign \new_[94866]_  = A267 & ~A266;
  assign \new_[94869]_  = A298 & ~A269;
  assign \new_[94870]_  = \new_[94869]_  & \new_[94866]_ ;
  assign \new_[94873]_  = ~A300 & ~A299;
  assign \new_[94876]_  = A302 & ~A301;
  assign \new_[94877]_  = \new_[94876]_  & \new_[94873]_ ;
  assign \new_[94878]_  = \new_[94877]_  & \new_[94870]_ ;
  assign \new_[94881]_  = ~A166 & ~A167;
  assign \new_[94884]_  = A200 & ~A199;
  assign \new_[94885]_  = \new_[94884]_  & \new_[94881]_ ;
  assign \new_[94888]_  = ~A202 & ~A201;
  assign \new_[94891]_  = A265 & A203;
  assign \new_[94892]_  = \new_[94891]_  & \new_[94888]_ ;
  assign \new_[94893]_  = \new_[94892]_  & \new_[94885]_ ;
  assign \new_[94896]_  = A267 & ~A266;
  assign \new_[94899]_  = ~A298 & ~A269;
  assign \new_[94900]_  = \new_[94899]_  & \new_[94896]_ ;
  assign \new_[94903]_  = ~A300 & A299;
  assign \new_[94906]_  = A302 & ~A301;
  assign \new_[94907]_  = \new_[94906]_  & \new_[94903]_ ;
  assign \new_[94908]_  = \new_[94907]_  & \new_[94900]_ ;
  assign \new_[94911]_  = ~A166 & ~A167;
  assign \new_[94914]_  = A200 & ~A199;
  assign \new_[94915]_  = \new_[94914]_  & \new_[94911]_ ;
  assign \new_[94918]_  = ~A202 & ~A201;
  assign \new_[94921]_  = A265 & A203;
  assign \new_[94922]_  = \new_[94921]_  & \new_[94918]_ ;
  assign \new_[94923]_  = \new_[94922]_  & \new_[94915]_ ;
  assign \new_[94926]_  = ~A267 & ~A266;
  assign \new_[94929]_  = A269 & ~A268;
  assign \new_[94930]_  = \new_[94929]_  & \new_[94926]_ ;
  assign \new_[94933]_  = ~A299 & A298;
  assign \new_[94936]_  = A301 & A300;
  assign \new_[94937]_  = \new_[94936]_  & \new_[94933]_ ;
  assign \new_[94938]_  = \new_[94937]_  & \new_[94930]_ ;
  assign \new_[94941]_  = ~A166 & ~A167;
  assign \new_[94944]_  = A200 & ~A199;
  assign \new_[94945]_  = \new_[94944]_  & \new_[94941]_ ;
  assign \new_[94948]_  = ~A202 & ~A201;
  assign \new_[94951]_  = A265 & A203;
  assign \new_[94952]_  = \new_[94951]_  & \new_[94948]_ ;
  assign \new_[94953]_  = \new_[94952]_  & \new_[94945]_ ;
  assign \new_[94956]_  = ~A267 & ~A266;
  assign \new_[94959]_  = A269 & ~A268;
  assign \new_[94960]_  = \new_[94959]_  & \new_[94956]_ ;
  assign \new_[94963]_  = ~A299 & A298;
  assign \new_[94966]_  = ~A302 & A300;
  assign \new_[94967]_  = \new_[94966]_  & \new_[94963]_ ;
  assign \new_[94968]_  = \new_[94967]_  & \new_[94960]_ ;
  assign \new_[94971]_  = ~A166 & ~A167;
  assign \new_[94974]_  = A200 & ~A199;
  assign \new_[94975]_  = \new_[94974]_  & \new_[94971]_ ;
  assign \new_[94978]_  = ~A202 & ~A201;
  assign \new_[94981]_  = A265 & A203;
  assign \new_[94982]_  = \new_[94981]_  & \new_[94978]_ ;
  assign \new_[94983]_  = \new_[94982]_  & \new_[94975]_ ;
  assign \new_[94986]_  = ~A267 & ~A266;
  assign \new_[94989]_  = A269 & ~A268;
  assign \new_[94990]_  = \new_[94989]_  & \new_[94986]_ ;
  assign \new_[94993]_  = A299 & ~A298;
  assign \new_[94996]_  = A301 & A300;
  assign \new_[94997]_  = \new_[94996]_  & \new_[94993]_ ;
  assign \new_[94998]_  = \new_[94997]_  & \new_[94990]_ ;
  assign \new_[95001]_  = ~A166 & ~A167;
  assign \new_[95004]_  = A200 & ~A199;
  assign \new_[95005]_  = \new_[95004]_  & \new_[95001]_ ;
  assign \new_[95008]_  = ~A202 & ~A201;
  assign \new_[95011]_  = A265 & A203;
  assign \new_[95012]_  = \new_[95011]_  & \new_[95008]_ ;
  assign \new_[95013]_  = \new_[95012]_  & \new_[95005]_ ;
  assign \new_[95016]_  = ~A267 & ~A266;
  assign \new_[95019]_  = A269 & ~A268;
  assign \new_[95020]_  = \new_[95019]_  & \new_[95016]_ ;
  assign \new_[95023]_  = A299 & ~A298;
  assign \new_[95026]_  = ~A302 & A300;
  assign \new_[95027]_  = \new_[95026]_  & \new_[95023]_ ;
  assign \new_[95028]_  = \new_[95027]_  & \new_[95020]_ ;
  assign \new_[95031]_  = ~A166 & ~A167;
  assign \new_[95034]_  = ~A200 & A199;
  assign \new_[95035]_  = \new_[95034]_  & \new_[95031]_ ;
  assign \new_[95038]_  = A202 & A201;
  assign \new_[95041]_  = A266 & ~A265;
  assign \new_[95042]_  = \new_[95041]_  & \new_[95038]_ ;
  assign \new_[95043]_  = \new_[95042]_  & \new_[95035]_ ;
  assign \new_[95046]_  = ~A268 & ~A267;
  assign \new_[95049]_  = A298 & A269;
  assign \new_[95050]_  = \new_[95049]_  & \new_[95046]_ ;
  assign \new_[95053]_  = ~A300 & ~A299;
  assign \new_[95056]_  = A302 & ~A301;
  assign \new_[95057]_  = \new_[95056]_  & \new_[95053]_ ;
  assign \new_[95058]_  = \new_[95057]_  & \new_[95050]_ ;
  assign \new_[95061]_  = ~A166 & ~A167;
  assign \new_[95064]_  = ~A200 & A199;
  assign \new_[95065]_  = \new_[95064]_  & \new_[95061]_ ;
  assign \new_[95068]_  = A202 & A201;
  assign \new_[95071]_  = A266 & ~A265;
  assign \new_[95072]_  = \new_[95071]_  & \new_[95068]_ ;
  assign \new_[95073]_  = \new_[95072]_  & \new_[95065]_ ;
  assign \new_[95076]_  = ~A268 & ~A267;
  assign \new_[95079]_  = ~A298 & A269;
  assign \new_[95080]_  = \new_[95079]_  & \new_[95076]_ ;
  assign \new_[95083]_  = ~A300 & A299;
  assign \new_[95086]_  = A302 & ~A301;
  assign \new_[95087]_  = \new_[95086]_  & \new_[95083]_ ;
  assign \new_[95088]_  = \new_[95087]_  & \new_[95080]_ ;
  assign \new_[95091]_  = ~A166 & ~A167;
  assign \new_[95094]_  = ~A200 & A199;
  assign \new_[95095]_  = \new_[95094]_  & \new_[95091]_ ;
  assign \new_[95098]_  = A202 & A201;
  assign \new_[95101]_  = ~A266 & A265;
  assign \new_[95102]_  = \new_[95101]_  & \new_[95098]_ ;
  assign \new_[95103]_  = \new_[95102]_  & \new_[95095]_ ;
  assign \new_[95106]_  = ~A268 & ~A267;
  assign \new_[95109]_  = A298 & A269;
  assign \new_[95110]_  = \new_[95109]_  & \new_[95106]_ ;
  assign \new_[95113]_  = ~A300 & ~A299;
  assign \new_[95116]_  = A302 & ~A301;
  assign \new_[95117]_  = \new_[95116]_  & \new_[95113]_ ;
  assign \new_[95118]_  = \new_[95117]_  & \new_[95110]_ ;
  assign \new_[95121]_  = ~A166 & ~A167;
  assign \new_[95124]_  = ~A200 & A199;
  assign \new_[95125]_  = \new_[95124]_  & \new_[95121]_ ;
  assign \new_[95128]_  = A202 & A201;
  assign \new_[95131]_  = ~A266 & A265;
  assign \new_[95132]_  = \new_[95131]_  & \new_[95128]_ ;
  assign \new_[95133]_  = \new_[95132]_  & \new_[95125]_ ;
  assign \new_[95136]_  = ~A268 & ~A267;
  assign \new_[95139]_  = ~A298 & A269;
  assign \new_[95140]_  = \new_[95139]_  & \new_[95136]_ ;
  assign \new_[95143]_  = ~A300 & A299;
  assign \new_[95146]_  = A302 & ~A301;
  assign \new_[95147]_  = \new_[95146]_  & \new_[95143]_ ;
  assign \new_[95148]_  = \new_[95147]_  & \new_[95140]_ ;
  assign \new_[95151]_  = ~A166 & ~A167;
  assign \new_[95154]_  = ~A200 & A199;
  assign \new_[95155]_  = \new_[95154]_  & \new_[95151]_ ;
  assign \new_[95158]_  = ~A203 & A201;
  assign \new_[95161]_  = A266 & ~A265;
  assign \new_[95162]_  = \new_[95161]_  & \new_[95158]_ ;
  assign \new_[95163]_  = \new_[95162]_  & \new_[95155]_ ;
  assign \new_[95166]_  = ~A268 & ~A267;
  assign \new_[95169]_  = A298 & A269;
  assign \new_[95170]_  = \new_[95169]_  & \new_[95166]_ ;
  assign \new_[95173]_  = ~A300 & ~A299;
  assign \new_[95176]_  = A302 & ~A301;
  assign \new_[95177]_  = \new_[95176]_  & \new_[95173]_ ;
  assign \new_[95178]_  = \new_[95177]_  & \new_[95170]_ ;
  assign \new_[95181]_  = ~A166 & ~A167;
  assign \new_[95184]_  = ~A200 & A199;
  assign \new_[95185]_  = \new_[95184]_  & \new_[95181]_ ;
  assign \new_[95188]_  = ~A203 & A201;
  assign \new_[95191]_  = A266 & ~A265;
  assign \new_[95192]_  = \new_[95191]_  & \new_[95188]_ ;
  assign \new_[95193]_  = \new_[95192]_  & \new_[95185]_ ;
  assign \new_[95196]_  = ~A268 & ~A267;
  assign \new_[95199]_  = ~A298 & A269;
  assign \new_[95200]_  = \new_[95199]_  & \new_[95196]_ ;
  assign \new_[95203]_  = ~A300 & A299;
  assign \new_[95206]_  = A302 & ~A301;
  assign \new_[95207]_  = \new_[95206]_  & \new_[95203]_ ;
  assign \new_[95208]_  = \new_[95207]_  & \new_[95200]_ ;
  assign \new_[95211]_  = ~A166 & ~A167;
  assign \new_[95214]_  = ~A200 & A199;
  assign \new_[95215]_  = \new_[95214]_  & \new_[95211]_ ;
  assign \new_[95218]_  = ~A203 & A201;
  assign \new_[95221]_  = ~A266 & A265;
  assign \new_[95222]_  = \new_[95221]_  & \new_[95218]_ ;
  assign \new_[95223]_  = \new_[95222]_  & \new_[95215]_ ;
  assign \new_[95226]_  = ~A268 & ~A267;
  assign \new_[95229]_  = A298 & A269;
  assign \new_[95230]_  = \new_[95229]_  & \new_[95226]_ ;
  assign \new_[95233]_  = ~A300 & ~A299;
  assign \new_[95236]_  = A302 & ~A301;
  assign \new_[95237]_  = \new_[95236]_  & \new_[95233]_ ;
  assign \new_[95238]_  = \new_[95237]_  & \new_[95230]_ ;
  assign \new_[95241]_  = ~A166 & ~A167;
  assign \new_[95244]_  = ~A200 & A199;
  assign \new_[95245]_  = \new_[95244]_  & \new_[95241]_ ;
  assign \new_[95248]_  = ~A203 & A201;
  assign \new_[95251]_  = ~A266 & A265;
  assign \new_[95252]_  = \new_[95251]_  & \new_[95248]_ ;
  assign \new_[95253]_  = \new_[95252]_  & \new_[95245]_ ;
  assign \new_[95256]_  = ~A268 & ~A267;
  assign \new_[95259]_  = ~A298 & A269;
  assign \new_[95260]_  = \new_[95259]_  & \new_[95256]_ ;
  assign \new_[95263]_  = ~A300 & A299;
  assign \new_[95266]_  = A302 & ~A301;
  assign \new_[95267]_  = \new_[95266]_  & \new_[95263]_ ;
  assign \new_[95268]_  = \new_[95267]_  & \new_[95260]_ ;
  assign \new_[95271]_  = ~A166 & ~A167;
  assign \new_[95274]_  = ~A200 & A199;
  assign \new_[95275]_  = \new_[95274]_  & \new_[95271]_ ;
  assign \new_[95278]_  = ~A202 & ~A201;
  assign \new_[95281]_  = ~A265 & A203;
  assign \new_[95282]_  = \new_[95281]_  & \new_[95278]_ ;
  assign \new_[95283]_  = \new_[95282]_  & \new_[95275]_ ;
  assign \new_[95286]_  = A267 & A266;
  assign \new_[95289]_  = A298 & A268;
  assign \new_[95290]_  = \new_[95289]_  & \new_[95286]_ ;
  assign \new_[95293]_  = ~A300 & ~A299;
  assign \new_[95296]_  = A302 & ~A301;
  assign \new_[95297]_  = \new_[95296]_  & \new_[95293]_ ;
  assign \new_[95298]_  = \new_[95297]_  & \new_[95290]_ ;
  assign \new_[95301]_  = ~A166 & ~A167;
  assign \new_[95304]_  = ~A200 & A199;
  assign \new_[95305]_  = \new_[95304]_  & \new_[95301]_ ;
  assign \new_[95308]_  = ~A202 & ~A201;
  assign \new_[95311]_  = ~A265 & A203;
  assign \new_[95312]_  = \new_[95311]_  & \new_[95308]_ ;
  assign \new_[95313]_  = \new_[95312]_  & \new_[95305]_ ;
  assign \new_[95316]_  = A267 & A266;
  assign \new_[95319]_  = ~A298 & A268;
  assign \new_[95320]_  = \new_[95319]_  & \new_[95316]_ ;
  assign \new_[95323]_  = ~A300 & A299;
  assign \new_[95326]_  = A302 & ~A301;
  assign \new_[95327]_  = \new_[95326]_  & \new_[95323]_ ;
  assign \new_[95328]_  = \new_[95327]_  & \new_[95320]_ ;
  assign \new_[95331]_  = ~A166 & ~A167;
  assign \new_[95334]_  = ~A200 & A199;
  assign \new_[95335]_  = \new_[95334]_  & \new_[95331]_ ;
  assign \new_[95338]_  = ~A202 & ~A201;
  assign \new_[95341]_  = ~A265 & A203;
  assign \new_[95342]_  = \new_[95341]_  & \new_[95338]_ ;
  assign \new_[95343]_  = \new_[95342]_  & \new_[95335]_ ;
  assign \new_[95346]_  = A267 & A266;
  assign \new_[95349]_  = A298 & ~A269;
  assign \new_[95350]_  = \new_[95349]_  & \new_[95346]_ ;
  assign \new_[95353]_  = ~A300 & ~A299;
  assign \new_[95356]_  = A302 & ~A301;
  assign \new_[95357]_  = \new_[95356]_  & \new_[95353]_ ;
  assign \new_[95358]_  = \new_[95357]_  & \new_[95350]_ ;
  assign \new_[95361]_  = ~A166 & ~A167;
  assign \new_[95364]_  = ~A200 & A199;
  assign \new_[95365]_  = \new_[95364]_  & \new_[95361]_ ;
  assign \new_[95368]_  = ~A202 & ~A201;
  assign \new_[95371]_  = ~A265 & A203;
  assign \new_[95372]_  = \new_[95371]_  & \new_[95368]_ ;
  assign \new_[95373]_  = \new_[95372]_  & \new_[95365]_ ;
  assign \new_[95376]_  = A267 & A266;
  assign \new_[95379]_  = ~A298 & ~A269;
  assign \new_[95380]_  = \new_[95379]_  & \new_[95376]_ ;
  assign \new_[95383]_  = ~A300 & A299;
  assign \new_[95386]_  = A302 & ~A301;
  assign \new_[95387]_  = \new_[95386]_  & \new_[95383]_ ;
  assign \new_[95388]_  = \new_[95387]_  & \new_[95380]_ ;
  assign \new_[95391]_  = ~A166 & ~A167;
  assign \new_[95394]_  = ~A200 & A199;
  assign \new_[95395]_  = \new_[95394]_  & \new_[95391]_ ;
  assign \new_[95398]_  = ~A202 & ~A201;
  assign \new_[95401]_  = ~A265 & A203;
  assign \new_[95402]_  = \new_[95401]_  & \new_[95398]_ ;
  assign \new_[95403]_  = \new_[95402]_  & \new_[95395]_ ;
  assign \new_[95406]_  = ~A267 & A266;
  assign \new_[95409]_  = A269 & ~A268;
  assign \new_[95410]_  = \new_[95409]_  & \new_[95406]_ ;
  assign \new_[95413]_  = ~A299 & A298;
  assign \new_[95416]_  = A301 & A300;
  assign \new_[95417]_  = \new_[95416]_  & \new_[95413]_ ;
  assign \new_[95418]_  = \new_[95417]_  & \new_[95410]_ ;
  assign \new_[95421]_  = ~A166 & ~A167;
  assign \new_[95424]_  = ~A200 & A199;
  assign \new_[95425]_  = \new_[95424]_  & \new_[95421]_ ;
  assign \new_[95428]_  = ~A202 & ~A201;
  assign \new_[95431]_  = ~A265 & A203;
  assign \new_[95432]_  = \new_[95431]_  & \new_[95428]_ ;
  assign \new_[95433]_  = \new_[95432]_  & \new_[95425]_ ;
  assign \new_[95436]_  = ~A267 & A266;
  assign \new_[95439]_  = A269 & ~A268;
  assign \new_[95440]_  = \new_[95439]_  & \new_[95436]_ ;
  assign \new_[95443]_  = ~A299 & A298;
  assign \new_[95446]_  = ~A302 & A300;
  assign \new_[95447]_  = \new_[95446]_  & \new_[95443]_ ;
  assign \new_[95448]_  = \new_[95447]_  & \new_[95440]_ ;
  assign \new_[95451]_  = ~A166 & ~A167;
  assign \new_[95454]_  = ~A200 & A199;
  assign \new_[95455]_  = \new_[95454]_  & \new_[95451]_ ;
  assign \new_[95458]_  = ~A202 & ~A201;
  assign \new_[95461]_  = ~A265 & A203;
  assign \new_[95462]_  = \new_[95461]_  & \new_[95458]_ ;
  assign \new_[95463]_  = \new_[95462]_  & \new_[95455]_ ;
  assign \new_[95466]_  = ~A267 & A266;
  assign \new_[95469]_  = A269 & ~A268;
  assign \new_[95470]_  = \new_[95469]_  & \new_[95466]_ ;
  assign \new_[95473]_  = A299 & ~A298;
  assign \new_[95476]_  = A301 & A300;
  assign \new_[95477]_  = \new_[95476]_  & \new_[95473]_ ;
  assign \new_[95478]_  = \new_[95477]_  & \new_[95470]_ ;
  assign \new_[95481]_  = ~A166 & ~A167;
  assign \new_[95484]_  = ~A200 & A199;
  assign \new_[95485]_  = \new_[95484]_  & \new_[95481]_ ;
  assign \new_[95488]_  = ~A202 & ~A201;
  assign \new_[95491]_  = ~A265 & A203;
  assign \new_[95492]_  = \new_[95491]_  & \new_[95488]_ ;
  assign \new_[95493]_  = \new_[95492]_  & \new_[95485]_ ;
  assign \new_[95496]_  = ~A267 & A266;
  assign \new_[95499]_  = A269 & ~A268;
  assign \new_[95500]_  = \new_[95499]_  & \new_[95496]_ ;
  assign \new_[95503]_  = A299 & ~A298;
  assign \new_[95506]_  = ~A302 & A300;
  assign \new_[95507]_  = \new_[95506]_  & \new_[95503]_ ;
  assign \new_[95508]_  = \new_[95507]_  & \new_[95500]_ ;
  assign \new_[95511]_  = ~A166 & ~A167;
  assign \new_[95514]_  = ~A200 & A199;
  assign \new_[95515]_  = \new_[95514]_  & \new_[95511]_ ;
  assign \new_[95518]_  = ~A202 & ~A201;
  assign \new_[95521]_  = A265 & A203;
  assign \new_[95522]_  = \new_[95521]_  & \new_[95518]_ ;
  assign \new_[95523]_  = \new_[95522]_  & \new_[95515]_ ;
  assign \new_[95526]_  = A267 & ~A266;
  assign \new_[95529]_  = A298 & A268;
  assign \new_[95530]_  = \new_[95529]_  & \new_[95526]_ ;
  assign \new_[95533]_  = ~A300 & ~A299;
  assign \new_[95536]_  = A302 & ~A301;
  assign \new_[95537]_  = \new_[95536]_  & \new_[95533]_ ;
  assign \new_[95538]_  = \new_[95537]_  & \new_[95530]_ ;
  assign \new_[95541]_  = ~A166 & ~A167;
  assign \new_[95544]_  = ~A200 & A199;
  assign \new_[95545]_  = \new_[95544]_  & \new_[95541]_ ;
  assign \new_[95548]_  = ~A202 & ~A201;
  assign \new_[95551]_  = A265 & A203;
  assign \new_[95552]_  = \new_[95551]_  & \new_[95548]_ ;
  assign \new_[95553]_  = \new_[95552]_  & \new_[95545]_ ;
  assign \new_[95556]_  = A267 & ~A266;
  assign \new_[95559]_  = ~A298 & A268;
  assign \new_[95560]_  = \new_[95559]_  & \new_[95556]_ ;
  assign \new_[95563]_  = ~A300 & A299;
  assign \new_[95566]_  = A302 & ~A301;
  assign \new_[95567]_  = \new_[95566]_  & \new_[95563]_ ;
  assign \new_[95568]_  = \new_[95567]_  & \new_[95560]_ ;
  assign \new_[95571]_  = ~A166 & ~A167;
  assign \new_[95574]_  = ~A200 & A199;
  assign \new_[95575]_  = \new_[95574]_  & \new_[95571]_ ;
  assign \new_[95578]_  = ~A202 & ~A201;
  assign \new_[95581]_  = A265 & A203;
  assign \new_[95582]_  = \new_[95581]_  & \new_[95578]_ ;
  assign \new_[95583]_  = \new_[95582]_  & \new_[95575]_ ;
  assign \new_[95586]_  = A267 & ~A266;
  assign \new_[95589]_  = A298 & ~A269;
  assign \new_[95590]_  = \new_[95589]_  & \new_[95586]_ ;
  assign \new_[95593]_  = ~A300 & ~A299;
  assign \new_[95596]_  = A302 & ~A301;
  assign \new_[95597]_  = \new_[95596]_  & \new_[95593]_ ;
  assign \new_[95598]_  = \new_[95597]_  & \new_[95590]_ ;
  assign \new_[95601]_  = ~A166 & ~A167;
  assign \new_[95604]_  = ~A200 & A199;
  assign \new_[95605]_  = \new_[95604]_  & \new_[95601]_ ;
  assign \new_[95608]_  = ~A202 & ~A201;
  assign \new_[95611]_  = A265 & A203;
  assign \new_[95612]_  = \new_[95611]_  & \new_[95608]_ ;
  assign \new_[95613]_  = \new_[95612]_  & \new_[95605]_ ;
  assign \new_[95616]_  = A267 & ~A266;
  assign \new_[95619]_  = ~A298 & ~A269;
  assign \new_[95620]_  = \new_[95619]_  & \new_[95616]_ ;
  assign \new_[95623]_  = ~A300 & A299;
  assign \new_[95626]_  = A302 & ~A301;
  assign \new_[95627]_  = \new_[95626]_  & \new_[95623]_ ;
  assign \new_[95628]_  = \new_[95627]_  & \new_[95620]_ ;
  assign \new_[95631]_  = ~A166 & ~A167;
  assign \new_[95634]_  = ~A200 & A199;
  assign \new_[95635]_  = \new_[95634]_  & \new_[95631]_ ;
  assign \new_[95638]_  = ~A202 & ~A201;
  assign \new_[95641]_  = A265 & A203;
  assign \new_[95642]_  = \new_[95641]_  & \new_[95638]_ ;
  assign \new_[95643]_  = \new_[95642]_  & \new_[95635]_ ;
  assign \new_[95646]_  = ~A267 & ~A266;
  assign \new_[95649]_  = A269 & ~A268;
  assign \new_[95650]_  = \new_[95649]_  & \new_[95646]_ ;
  assign \new_[95653]_  = ~A299 & A298;
  assign \new_[95656]_  = A301 & A300;
  assign \new_[95657]_  = \new_[95656]_  & \new_[95653]_ ;
  assign \new_[95658]_  = \new_[95657]_  & \new_[95650]_ ;
  assign \new_[95661]_  = ~A166 & ~A167;
  assign \new_[95664]_  = ~A200 & A199;
  assign \new_[95665]_  = \new_[95664]_  & \new_[95661]_ ;
  assign \new_[95668]_  = ~A202 & ~A201;
  assign \new_[95671]_  = A265 & A203;
  assign \new_[95672]_  = \new_[95671]_  & \new_[95668]_ ;
  assign \new_[95673]_  = \new_[95672]_  & \new_[95665]_ ;
  assign \new_[95676]_  = ~A267 & ~A266;
  assign \new_[95679]_  = A269 & ~A268;
  assign \new_[95680]_  = \new_[95679]_  & \new_[95676]_ ;
  assign \new_[95683]_  = ~A299 & A298;
  assign \new_[95686]_  = ~A302 & A300;
  assign \new_[95687]_  = \new_[95686]_  & \new_[95683]_ ;
  assign \new_[95688]_  = \new_[95687]_  & \new_[95680]_ ;
  assign \new_[95691]_  = ~A166 & ~A167;
  assign \new_[95694]_  = ~A200 & A199;
  assign \new_[95695]_  = \new_[95694]_  & \new_[95691]_ ;
  assign \new_[95698]_  = ~A202 & ~A201;
  assign \new_[95701]_  = A265 & A203;
  assign \new_[95702]_  = \new_[95701]_  & \new_[95698]_ ;
  assign \new_[95703]_  = \new_[95702]_  & \new_[95695]_ ;
  assign \new_[95706]_  = ~A267 & ~A266;
  assign \new_[95709]_  = A269 & ~A268;
  assign \new_[95710]_  = \new_[95709]_  & \new_[95706]_ ;
  assign \new_[95713]_  = A299 & ~A298;
  assign \new_[95716]_  = A301 & A300;
  assign \new_[95717]_  = \new_[95716]_  & \new_[95713]_ ;
  assign \new_[95718]_  = \new_[95717]_  & \new_[95710]_ ;
  assign \new_[95721]_  = ~A166 & ~A167;
  assign \new_[95724]_  = ~A200 & A199;
  assign \new_[95725]_  = \new_[95724]_  & \new_[95721]_ ;
  assign \new_[95728]_  = ~A202 & ~A201;
  assign \new_[95731]_  = A265 & A203;
  assign \new_[95732]_  = \new_[95731]_  & \new_[95728]_ ;
  assign \new_[95733]_  = \new_[95732]_  & \new_[95725]_ ;
  assign \new_[95736]_  = ~A267 & ~A266;
  assign \new_[95739]_  = A269 & ~A268;
  assign \new_[95740]_  = \new_[95739]_  & \new_[95736]_ ;
  assign \new_[95743]_  = A299 & ~A298;
  assign \new_[95746]_  = ~A302 & A300;
  assign \new_[95747]_  = \new_[95746]_  & \new_[95743]_ ;
  assign \new_[95748]_  = \new_[95747]_  & \new_[95740]_ ;
  assign \new_[95751]_  = ~A168 & A170;
  assign \new_[95754]_  = A200 & ~A199;
  assign \new_[95755]_  = \new_[95754]_  & \new_[95751]_ ;
  assign \new_[95758]_  = A202 & A201;
  assign \new_[95761]_  = A266 & ~A265;
  assign \new_[95762]_  = \new_[95761]_  & \new_[95758]_ ;
  assign \new_[95763]_  = \new_[95762]_  & \new_[95755]_ ;
  assign \new_[95766]_  = ~A268 & ~A267;
  assign \new_[95769]_  = A298 & A269;
  assign \new_[95770]_  = \new_[95769]_  & \new_[95766]_ ;
  assign \new_[95773]_  = ~A300 & ~A299;
  assign \new_[95776]_  = A302 & ~A301;
  assign \new_[95777]_  = \new_[95776]_  & \new_[95773]_ ;
  assign \new_[95778]_  = \new_[95777]_  & \new_[95770]_ ;
  assign \new_[95781]_  = ~A168 & A170;
  assign \new_[95784]_  = A200 & ~A199;
  assign \new_[95785]_  = \new_[95784]_  & \new_[95781]_ ;
  assign \new_[95788]_  = A202 & A201;
  assign \new_[95791]_  = A266 & ~A265;
  assign \new_[95792]_  = \new_[95791]_  & \new_[95788]_ ;
  assign \new_[95793]_  = \new_[95792]_  & \new_[95785]_ ;
  assign \new_[95796]_  = ~A268 & ~A267;
  assign \new_[95799]_  = ~A298 & A269;
  assign \new_[95800]_  = \new_[95799]_  & \new_[95796]_ ;
  assign \new_[95803]_  = ~A300 & A299;
  assign \new_[95806]_  = A302 & ~A301;
  assign \new_[95807]_  = \new_[95806]_  & \new_[95803]_ ;
  assign \new_[95808]_  = \new_[95807]_  & \new_[95800]_ ;
  assign \new_[95811]_  = ~A168 & A170;
  assign \new_[95814]_  = A200 & ~A199;
  assign \new_[95815]_  = \new_[95814]_  & \new_[95811]_ ;
  assign \new_[95818]_  = A202 & A201;
  assign \new_[95821]_  = ~A266 & A265;
  assign \new_[95822]_  = \new_[95821]_  & \new_[95818]_ ;
  assign \new_[95823]_  = \new_[95822]_  & \new_[95815]_ ;
  assign \new_[95826]_  = ~A268 & ~A267;
  assign \new_[95829]_  = A298 & A269;
  assign \new_[95830]_  = \new_[95829]_  & \new_[95826]_ ;
  assign \new_[95833]_  = ~A300 & ~A299;
  assign \new_[95836]_  = A302 & ~A301;
  assign \new_[95837]_  = \new_[95836]_  & \new_[95833]_ ;
  assign \new_[95838]_  = \new_[95837]_  & \new_[95830]_ ;
  assign \new_[95841]_  = ~A168 & A170;
  assign \new_[95844]_  = A200 & ~A199;
  assign \new_[95845]_  = \new_[95844]_  & \new_[95841]_ ;
  assign \new_[95848]_  = A202 & A201;
  assign \new_[95851]_  = ~A266 & A265;
  assign \new_[95852]_  = \new_[95851]_  & \new_[95848]_ ;
  assign \new_[95853]_  = \new_[95852]_  & \new_[95845]_ ;
  assign \new_[95856]_  = ~A268 & ~A267;
  assign \new_[95859]_  = ~A298 & A269;
  assign \new_[95860]_  = \new_[95859]_  & \new_[95856]_ ;
  assign \new_[95863]_  = ~A300 & A299;
  assign \new_[95866]_  = A302 & ~A301;
  assign \new_[95867]_  = \new_[95866]_  & \new_[95863]_ ;
  assign \new_[95868]_  = \new_[95867]_  & \new_[95860]_ ;
  assign \new_[95871]_  = ~A168 & A170;
  assign \new_[95874]_  = A200 & ~A199;
  assign \new_[95875]_  = \new_[95874]_  & \new_[95871]_ ;
  assign \new_[95878]_  = ~A203 & A201;
  assign \new_[95881]_  = A266 & ~A265;
  assign \new_[95882]_  = \new_[95881]_  & \new_[95878]_ ;
  assign \new_[95883]_  = \new_[95882]_  & \new_[95875]_ ;
  assign \new_[95886]_  = ~A268 & ~A267;
  assign \new_[95889]_  = A298 & A269;
  assign \new_[95890]_  = \new_[95889]_  & \new_[95886]_ ;
  assign \new_[95893]_  = ~A300 & ~A299;
  assign \new_[95896]_  = A302 & ~A301;
  assign \new_[95897]_  = \new_[95896]_  & \new_[95893]_ ;
  assign \new_[95898]_  = \new_[95897]_  & \new_[95890]_ ;
  assign \new_[95901]_  = ~A168 & A170;
  assign \new_[95904]_  = A200 & ~A199;
  assign \new_[95905]_  = \new_[95904]_  & \new_[95901]_ ;
  assign \new_[95908]_  = ~A203 & A201;
  assign \new_[95911]_  = A266 & ~A265;
  assign \new_[95912]_  = \new_[95911]_  & \new_[95908]_ ;
  assign \new_[95913]_  = \new_[95912]_  & \new_[95905]_ ;
  assign \new_[95916]_  = ~A268 & ~A267;
  assign \new_[95919]_  = ~A298 & A269;
  assign \new_[95920]_  = \new_[95919]_  & \new_[95916]_ ;
  assign \new_[95923]_  = ~A300 & A299;
  assign \new_[95926]_  = A302 & ~A301;
  assign \new_[95927]_  = \new_[95926]_  & \new_[95923]_ ;
  assign \new_[95928]_  = \new_[95927]_  & \new_[95920]_ ;
  assign \new_[95931]_  = ~A168 & A170;
  assign \new_[95934]_  = A200 & ~A199;
  assign \new_[95935]_  = \new_[95934]_  & \new_[95931]_ ;
  assign \new_[95938]_  = ~A203 & A201;
  assign \new_[95941]_  = ~A266 & A265;
  assign \new_[95942]_  = \new_[95941]_  & \new_[95938]_ ;
  assign \new_[95943]_  = \new_[95942]_  & \new_[95935]_ ;
  assign \new_[95946]_  = ~A268 & ~A267;
  assign \new_[95949]_  = A298 & A269;
  assign \new_[95950]_  = \new_[95949]_  & \new_[95946]_ ;
  assign \new_[95953]_  = ~A300 & ~A299;
  assign \new_[95956]_  = A302 & ~A301;
  assign \new_[95957]_  = \new_[95956]_  & \new_[95953]_ ;
  assign \new_[95958]_  = \new_[95957]_  & \new_[95950]_ ;
  assign \new_[95961]_  = ~A168 & A170;
  assign \new_[95964]_  = A200 & ~A199;
  assign \new_[95965]_  = \new_[95964]_  & \new_[95961]_ ;
  assign \new_[95968]_  = ~A203 & A201;
  assign \new_[95971]_  = ~A266 & A265;
  assign \new_[95972]_  = \new_[95971]_  & \new_[95968]_ ;
  assign \new_[95973]_  = \new_[95972]_  & \new_[95965]_ ;
  assign \new_[95976]_  = ~A268 & ~A267;
  assign \new_[95979]_  = ~A298 & A269;
  assign \new_[95980]_  = \new_[95979]_  & \new_[95976]_ ;
  assign \new_[95983]_  = ~A300 & A299;
  assign \new_[95986]_  = A302 & ~A301;
  assign \new_[95987]_  = \new_[95986]_  & \new_[95983]_ ;
  assign \new_[95988]_  = \new_[95987]_  & \new_[95980]_ ;
  assign \new_[95991]_  = ~A168 & A170;
  assign \new_[95994]_  = A200 & ~A199;
  assign \new_[95995]_  = \new_[95994]_  & \new_[95991]_ ;
  assign \new_[95998]_  = ~A202 & ~A201;
  assign \new_[96001]_  = ~A265 & A203;
  assign \new_[96002]_  = \new_[96001]_  & \new_[95998]_ ;
  assign \new_[96003]_  = \new_[96002]_  & \new_[95995]_ ;
  assign \new_[96006]_  = A267 & A266;
  assign \new_[96009]_  = A298 & A268;
  assign \new_[96010]_  = \new_[96009]_  & \new_[96006]_ ;
  assign \new_[96013]_  = ~A300 & ~A299;
  assign \new_[96016]_  = A302 & ~A301;
  assign \new_[96017]_  = \new_[96016]_  & \new_[96013]_ ;
  assign \new_[96018]_  = \new_[96017]_  & \new_[96010]_ ;
  assign \new_[96021]_  = ~A168 & A170;
  assign \new_[96024]_  = A200 & ~A199;
  assign \new_[96025]_  = \new_[96024]_  & \new_[96021]_ ;
  assign \new_[96028]_  = ~A202 & ~A201;
  assign \new_[96031]_  = ~A265 & A203;
  assign \new_[96032]_  = \new_[96031]_  & \new_[96028]_ ;
  assign \new_[96033]_  = \new_[96032]_  & \new_[96025]_ ;
  assign \new_[96036]_  = A267 & A266;
  assign \new_[96039]_  = ~A298 & A268;
  assign \new_[96040]_  = \new_[96039]_  & \new_[96036]_ ;
  assign \new_[96043]_  = ~A300 & A299;
  assign \new_[96046]_  = A302 & ~A301;
  assign \new_[96047]_  = \new_[96046]_  & \new_[96043]_ ;
  assign \new_[96048]_  = \new_[96047]_  & \new_[96040]_ ;
  assign \new_[96051]_  = ~A168 & A170;
  assign \new_[96054]_  = A200 & ~A199;
  assign \new_[96055]_  = \new_[96054]_  & \new_[96051]_ ;
  assign \new_[96058]_  = ~A202 & ~A201;
  assign \new_[96061]_  = ~A265 & A203;
  assign \new_[96062]_  = \new_[96061]_  & \new_[96058]_ ;
  assign \new_[96063]_  = \new_[96062]_  & \new_[96055]_ ;
  assign \new_[96066]_  = A267 & A266;
  assign \new_[96069]_  = A298 & ~A269;
  assign \new_[96070]_  = \new_[96069]_  & \new_[96066]_ ;
  assign \new_[96073]_  = ~A300 & ~A299;
  assign \new_[96076]_  = A302 & ~A301;
  assign \new_[96077]_  = \new_[96076]_  & \new_[96073]_ ;
  assign \new_[96078]_  = \new_[96077]_  & \new_[96070]_ ;
  assign \new_[96081]_  = ~A168 & A170;
  assign \new_[96084]_  = A200 & ~A199;
  assign \new_[96085]_  = \new_[96084]_  & \new_[96081]_ ;
  assign \new_[96088]_  = ~A202 & ~A201;
  assign \new_[96091]_  = ~A265 & A203;
  assign \new_[96092]_  = \new_[96091]_  & \new_[96088]_ ;
  assign \new_[96093]_  = \new_[96092]_  & \new_[96085]_ ;
  assign \new_[96096]_  = A267 & A266;
  assign \new_[96099]_  = ~A298 & ~A269;
  assign \new_[96100]_  = \new_[96099]_  & \new_[96096]_ ;
  assign \new_[96103]_  = ~A300 & A299;
  assign \new_[96106]_  = A302 & ~A301;
  assign \new_[96107]_  = \new_[96106]_  & \new_[96103]_ ;
  assign \new_[96108]_  = \new_[96107]_  & \new_[96100]_ ;
  assign \new_[96111]_  = ~A168 & A170;
  assign \new_[96114]_  = A200 & ~A199;
  assign \new_[96115]_  = \new_[96114]_  & \new_[96111]_ ;
  assign \new_[96118]_  = ~A202 & ~A201;
  assign \new_[96121]_  = ~A265 & A203;
  assign \new_[96122]_  = \new_[96121]_  & \new_[96118]_ ;
  assign \new_[96123]_  = \new_[96122]_  & \new_[96115]_ ;
  assign \new_[96126]_  = ~A267 & A266;
  assign \new_[96129]_  = A269 & ~A268;
  assign \new_[96130]_  = \new_[96129]_  & \new_[96126]_ ;
  assign \new_[96133]_  = ~A299 & A298;
  assign \new_[96136]_  = A301 & A300;
  assign \new_[96137]_  = \new_[96136]_  & \new_[96133]_ ;
  assign \new_[96138]_  = \new_[96137]_  & \new_[96130]_ ;
  assign \new_[96141]_  = ~A168 & A170;
  assign \new_[96144]_  = A200 & ~A199;
  assign \new_[96145]_  = \new_[96144]_  & \new_[96141]_ ;
  assign \new_[96148]_  = ~A202 & ~A201;
  assign \new_[96151]_  = ~A265 & A203;
  assign \new_[96152]_  = \new_[96151]_  & \new_[96148]_ ;
  assign \new_[96153]_  = \new_[96152]_  & \new_[96145]_ ;
  assign \new_[96156]_  = ~A267 & A266;
  assign \new_[96159]_  = A269 & ~A268;
  assign \new_[96160]_  = \new_[96159]_  & \new_[96156]_ ;
  assign \new_[96163]_  = ~A299 & A298;
  assign \new_[96166]_  = ~A302 & A300;
  assign \new_[96167]_  = \new_[96166]_  & \new_[96163]_ ;
  assign \new_[96168]_  = \new_[96167]_  & \new_[96160]_ ;
  assign \new_[96171]_  = ~A168 & A170;
  assign \new_[96174]_  = A200 & ~A199;
  assign \new_[96175]_  = \new_[96174]_  & \new_[96171]_ ;
  assign \new_[96178]_  = ~A202 & ~A201;
  assign \new_[96181]_  = ~A265 & A203;
  assign \new_[96182]_  = \new_[96181]_  & \new_[96178]_ ;
  assign \new_[96183]_  = \new_[96182]_  & \new_[96175]_ ;
  assign \new_[96186]_  = ~A267 & A266;
  assign \new_[96189]_  = A269 & ~A268;
  assign \new_[96190]_  = \new_[96189]_  & \new_[96186]_ ;
  assign \new_[96193]_  = A299 & ~A298;
  assign \new_[96196]_  = A301 & A300;
  assign \new_[96197]_  = \new_[96196]_  & \new_[96193]_ ;
  assign \new_[96198]_  = \new_[96197]_  & \new_[96190]_ ;
  assign \new_[96201]_  = ~A168 & A170;
  assign \new_[96204]_  = A200 & ~A199;
  assign \new_[96205]_  = \new_[96204]_  & \new_[96201]_ ;
  assign \new_[96208]_  = ~A202 & ~A201;
  assign \new_[96211]_  = ~A265 & A203;
  assign \new_[96212]_  = \new_[96211]_  & \new_[96208]_ ;
  assign \new_[96213]_  = \new_[96212]_  & \new_[96205]_ ;
  assign \new_[96216]_  = ~A267 & A266;
  assign \new_[96219]_  = A269 & ~A268;
  assign \new_[96220]_  = \new_[96219]_  & \new_[96216]_ ;
  assign \new_[96223]_  = A299 & ~A298;
  assign \new_[96226]_  = ~A302 & A300;
  assign \new_[96227]_  = \new_[96226]_  & \new_[96223]_ ;
  assign \new_[96228]_  = \new_[96227]_  & \new_[96220]_ ;
  assign \new_[96231]_  = ~A168 & A170;
  assign \new_[96234]_  = A200 & ~A199;
  assign \new_[96235]_  = \new_[96234]_  & \new_[96231]_ ;
  assign \new_[96238]_  = ~A202 & ~A201;
  assign \new_[96241]_  = A265 & A203;
  assign \new_[96242]_  = \new_[96241]_  & \new_[96238]_ ;
  assign \new_[96243]_  = \new_[96242]_  & \new_[96235]_ ;
  assign \new_[96246]_  = A267 & ~A266;
  assign \new_[96249]_  = A298 & A268;
  assign \new_[96250]_  = \new_[96249]_  & \new_[96246]_ ;
  assign \new_[96253]_  = ~A300 & ~A299;
  assign \new_[96256]_  = A302 & ~A301;
  assign \new_[96257]_  = \new_[96256]_  & \new_[96253]_ ;
  assign \new_[96258]_  = \new_[96257]_  & \new_[96250]_ ;
  assign \new_[96261]_  = ~A168 & A170;
  assign \new_[96264]_  = A200 & ~A199;
  assign \new_[96265]_  = \new_[96264]_  & \new_[96261]_ ;
  assign \new_[96268]_  = ~A202 & ~A201;
  assign \new_[96271]_  = A265 & A203;
  assign \new_[96272]_  = \new_[96271]_  & \new_[96268]_ ;
  assign \new_[96273]_  = \new_[96272]_  & \new_[96265]_ ;
  assign \new_[96276]_  = A267 & ~A266;
  assign \new_[96279]_  = ~A298 & A268;
  assign \new_[96280]_  = \new_[96279]_  & \new_[96276]_ ;
  assign \new_[96283]_  = ~A300 & A299;
  assign \new_[96286]_  = A302 & ~A301;
  assign \new_[96287]_  = \new_[96286]_  & \new_[96283]_ ;
  assign \new_[96288]_  = \new_[96287]_  & \new_[96280]_ ;
  assign \new_[96291]_  = ~A168 & A170;
  assign \new_[96294]_  = A200 & ~A199;
  assign \new_[96295]_  = \new_[96294]_  & \new_[96291]_ ;
  assign \new_[96298]_  = ~A202 & ~A201;
  assign \new_[96301]_  = A265 & A203;
  assign \new_[96302]_  = \new_[96301]_  & \new_[96298]_ ;
  assign \new_[96303]_  = \new_[96302]_  & \new_[96295]_ ;
  assign \new_[96306]_  = A267 & ~A266;
  assign \new_[96309]_  = A298 & ~A269;
  assign \new_[96310]_  = \new_[96309]_  & \new_[96306]_ ;
  assign \new_[96313]_  = ~A300 & ~A299;
  assign \new_[96316]_  = A302 & ~A301;
  assign \new_[96317]_  = \new_[96316]_  & \new_[96313]_ ;
  assign \new_[96318]_  = \new_[96317]_  & \new_[96310]_ ;
  assign \new_[96321]_  = ~A168 & A170;
  assign \new_[96324]_  = A200 & ~A199;
  assign \new_[96325]_  = \new_[96324]_  & \new_[96321]_ ;
  assign \new_[96328]_  = ~A202 & ~A201;
  assign \new_[96331]_  = A265 & A203;
  assign \new_[96332]_  = \new_[96331]_  & \new_[96328]_ ;
  assign \new_[96333]_  = \new_[96332]_  & \new_[96325]_ ;
  assign \new_[96336]_  = A267 & ~A266;
  assign \new_[96339]_  = ~A298 & ~A269;
  assign \new_[96340]_  = \new_[96339]_  & \new_[96336]_ ;
  assign \new_[96343]_  = ~A300 & A299;
  assign \new_[96346]_  = A302 & ~A301;
  assign \new_[96347]_  = \new_[96346]_  & \new_[96343]_ ;
  assign \new_[96348]_  = \new_[96347]_  & \new_[96340]_ ;
  assign \new_[96351]_  = ~A168 & A170;
  assign \new_[96354]_  = A200 & ~A199;
  assign \new_[96355]_  = \new_[96354]_  & \new_[96351]_ ;
  assign \new_[96358]_  = ~A202 & ~A201;
  assign \new_[96361]_  = A265 & A203;
  assign \new_[96362]_  = \new_[96361]_  & \new_[96358]_ ;
  assign \new_[96363]_  = \new_[96362]_  & \new_[96355]_ ;
  assign \new_[96366]_  = ~A267 & ~A266;
  assign \new_[96369]_  = A269 & ~A268;
  assign \new_[96370]_  = \new_[96369]_  & \new_[96366]_ ;
  assign \new_[96373]_  = ~A299 & A298;
  assign \new_[96376]_  = A301 & A300;
  assign \new_[96377]_  = \new_[96376]_  & \new_[96373]_ ;
  assign \new_[96378]_  = \new_[96377]_  & \new_[96370]_ ;
  assign \new_[96381]_  = ~A168 & A170;
  assign \new_[96384]_  = A200 & ~A199;
  assign \new_[96385]_  = \new_[96384]_  & \new_[96381]_ ;
  assign \new_[96388]_  = ~A202 & ~A201;
  assign \new_[96391]_  = A265 & A203;
  assign \new_[96392]_  = \new_[96391]_  & \new_[96388]_ ;
  assign \new_[96393]_  = \new_[96392]_  & \new_[96385]_ ;
  assign \new_[96396]_  = ~A267 & ~A266;
  assign \new_[96399]_  = A269 & ~A268;
  assign \new_[96400]_  = \new_[96399]_  & \new_[96396]_ ;
  assign \new_[96403]_  = ~A299 & A298;
  assign \new_[96406]_  = ~A302 & A300;
  assign \new_[96407]_  = \new_[96406]_  & \new_[96403]_ ;
  assign \new_[96408]_  = \new_[96407]_  & \new_[96400]_ ;
  assign \new_[96411]_  = ~A168 & A170;
  assign \new_[96414]_  = A200 & ~A199;
  assign \new_[96415]_  = \new_[96414]_  & \new_[96411]_ ;
  assign \new_[96418]_  = ~A202 & ~A201;
  assign \new_[96421]_  = A265 & A203;
  assign \new_[96422]_  = \new_[96421]_  & \new_[96418]_ ;
  assign \new_[96423]_  = \new_[96422]_  & \new_[96415]_ ;
  assign \new_[96426]_  = ~A267 & ~A266;
  assign \new_[96429]_  = A269 & ~A268;
  assign \new_[96430]_  = \new_[96429]_  & \new_[96426]_ ;
  assign \new_[96433]_  = A299 & ~A298;
  assign \new_[96436]_  = A301 & A300;
  assign \new_[96437]_  = \new_[96436]_  & \new_[96433]_ ;
  assign \new_[96438]_  = \new_[96437]_  & \new_[96430]_ ;
  assign \new_[96441]_  = ~A168 & A170;
  assign \new_[96444]_  = A200 & ~A199;
  assign \new_[96445]_  = \new_[96444]_  & \new_[96441]_ ;
  assign \new_[96448]_  = ~A202 & ~A201;
  assign \new_[96451]_  = A265 & A203;
  assign \new_[96452]_  = \new_[96451]_  & \new_[96448]_ ;
  assign \new_[96453]_  = \new_[96452]_  & \new_[96445]_ ;
  assign \new_[96456]_  = ~A267 & ~A266;
  assign \new_[96459]_  = A269 & ~A268;
  assign \new_[96460]_  = \new_[96459]_  & \new_[96456]_ ;
  assign \new_[96463]_  = A299 & ~A298;
  assign \new_[96466]_  = ~A302 & A300;
  assign \new_[96467]_  = \new_[96466]_  & \new_[96463]_ ;
  assign \new_[96468]_  = \new_[96467]_  & \new_[96460]_ ;
  assign \new_[96471]_  = ~A168 & A170;
  assign \new_[96474]_  = ~A200 & A199;
  assign \new_[96475]_  = \new_[96474]_  & \new_[96471]_ ;
  assign \new_[96478]_  = A202 & A201;
  assign \new_[96481]_  = A266 & ~A265;
  assign \new_[96482]_  = \new_[96481]_  & \new_[96478]_ ;
  assign \new_[96483]_  = \new_[96482]_  & \new_[96475]_ ;
  assign \new_[96486]_  = ~A268 & ~A267;
  assign \new_[96489]_  = A298 & A269;
  assign \new_[96490]_  = \new_[96489]_  & \new_[96486]_ ;
  assign \new_[96493]_  = ~A300 & ~A299;
  assign \new_[96496]_  = A302 & ~A301;
  assign \new_[96497]_  = \new_[96496]_  & \new_[96493]_ ;
  assign \new_[96498]_  = \new_[96497]_  & \new_[96490]_ ;
  assign \new_[96501]_  = ~A168 & A170;
  assign \new_[96504]_  = ~A200 & A199;
  assign \new_[96505]_  = \new_[96504]_  & \new_[96501]_ ;
  assign \new_[96508]_  = A202 & A201;
  assign \new_[96511]_  = A266 & ~A265;
  assign \new_[96512]_  = \new_[96511]_  & \new_[96508]_ ;
  assign \new_[96513]_  = \new_[96512]_  & \new_[96505]_ ;
  assign \new_[96516]_  = ~A268 & ~A267;
  assign \new_[96519]_  = ~A298 & A269;
  assign \new_[96520]_  = \new_[96519]_  & \new_[96516]_ ;
  assign \new_[96523]_  = ~A300 & A299;
  assign \new_[96526]_  = A302 & ~A301;
  assign \new_[96527]_  = \new_[96526]_  & \new_[96523]_ ;
  assign \new_[96528]_  = \new_[96527]_  & \new_[96520]_ ;
  assign \new_[96531]_  = ~A168 & A170;
  assign \new_[96534]_  = ~A200 & A199;
  assign \new_[96535]_  = \new_[96534]_  & \new_[96531]_ ;
  assign \new_[96538]_  = A202 & A201;
  assign \new_[96541]_  = ~A266 & A265;
  assign \new_[96542]_  = \new_[96541]_  & \new_[96538]_ ;
  assign \new_[96543]_  = \new_[96542]_  & \new_[96535]_ ;
  assign \new_[96546]_  = ~A268 & ~A267;
  assign \new_[96549]_  = A298 & A269;
  assign \new_[96550]_  = \new_[96549]_  & \new_[96546]_ ;
  assign \new_[96553]_  = ~A300 & ~A299;
  assign \new_[96556]_  = A302 & ~A301;
  assign \new_[96557]_  = \new_[96556]_  & \new_[96553]_ ;
  assign \new_[96558]_  = \new_[96557]_  & \new_[96550]_ ;
  assign \new_[96561]_  = ~A168 & A170;
  assign \new_[96564]_  = ~A200 & A199;
  assign \new_[96565]_  = \new_[96564]_  & \new_[96561]_ ;
  assign \new_[96568]_  = A202 & A201;
  assign \new_[96571]_  = ~A266 & A265;
  assign \new_[96572]_  = \new_[96571]_  & \new_[96568]_ ;
  assign \new_[96573]_  = \new_[96572]_  & \new_[96565]_ ;
  assign \new_[96576]_  = ~A268 & ~A267;
  assign \new_[96579]_  = ~A298 & A269;
  assign \new_[96580]_  = \new_[96579]_  & \new_[96576]_ ;
  assign \new_[96583]_  = ~A300 & A299;
  assign \new_[96586]_  = A302 & ~A301;
  assign \new_[96587]_  = \new_[96586]_  & \new_[96583]_ ;
  assign \new_[96588]_  = \new_[96587]_  & \new_[96580]_ ;
  assign \new_[96591]_  = ~A168 & A170;
  assign \new_[96594]_  = ~A200 & A199;
  assign \new_[96595]_  = \new_[96594]_  & \new_[96591]_ ;
  assign \new_[96598]_  = ~A203 & A201;
  assign \new_[96601]_  = A266 & ~A265;
  assign \new_[96602]_  = \new_[96601]_  & \new_[96598]_ ;
  assign \new_[96603]_  = \new_[96602]_  & \new_[96595]_ ;
  assign \new_[96606]_  = ~A268 & ~A267;
  assign \new_[96609]_  = A298 & A269;
  assign \new_[96610]_  = \new_[96609]_  & \new_[96606]_ ;
  assign \new_[96613]_  = ~A300 & ~A299;
  assign \new_[96616]_  = A302 & ~A301;
  assign \new_[96617]_  = \new_[96616]_  & \new_[96613]_ ;
  assign \new_[96618]_  = \new_[96617]_  & \new_[96610]_ ;
  assign \new_[96621]_  = ~A168 & A170;
  assign \new_[96624]_  = ~A200 & A199;
  assign \new_[96625]_  = \new_[96624]_  & \new_[96621]_ ;
  assign \new_[96628]_  = ~A203 & A201;
  assign \new_[96631]_  = A266 & ~A265;
  assign \new_[96632]_  = \new_[96631]_  & \new_[96628]_ ;
  assign \new_[96633]_  = \new_[96632]_  & \new_[96625]_ ;
  assign \new_[96636]_  = ~A268 & ~A267;
  assign \new_[96639]_  = ~A298 & A269;
  assign \new_[96640]_  = \new_[96639]_  & \new_[96636]_ ;
  assign \new_[96643]_  = ~A300 & A299;
  assign \new_[96646]_  = A302 & ~A301;
  assign \new_[96647]_  = \new_[96646]_  & \new_[96643]_ ;
  assign \new_[96648]_  = \new_[96647]_  & \new_[96640]_ ;
  assign \new_[96651]_  = ~A168 & A170;
  assign \new_[96654]_  = ~A200 & A199;
  assign \new_[96655]_  = \new_[96654]_  & \new_[96651]_ ;
  assign \new_[96658]_  = ~A203 & A201;
  assign \new_[96661]_  = ~A266 & A265;
  assign \new_[96662]_  = \new_[96661]_  & \new_[96658]_ ;
  assign \new_[96663]_  = \new_[96662]_  & \new_[96655]_ ;
  assign \new_[96666]_  = ~A268 & ~A267;
  assign \new_[96669]_  = A298 & A269;
  assign \new_[96670]_  = \new_[96669]_  & \new_[96666]_ ;
  assign \new_[96673]_  = ~A300 & ~A299;
  assign \new_[96676]_  = A302 & ~A301;
  assign \new_[96677]_  = \new_[96676]_  & \new_[96673]_ ;
  assign \new_[96678]_  = \new_[96677]_  & \new_[96670]_ ;
  assign \new_[96681]_  = ~A168 & A170;
  assign \new_[96684]_  = ~A200 & A199;
  assign \new_[96685]_  = \new_[96684]_  & \new_[96681]_ ;
  assign \new_[96688]_  = ~A203 & A201;
  assign \new_[96691]_  = ~A266 & A265;
  assign \new_[96692]_  = \new_[96691]_  & \new_[96688]_ ;
  assign \new_[96693]_  = \new_[96692]_  & \new_[96685]_ ;
  assign \new_[96696]_  = ~A268 & ~A267;
  assign \new_[96699]_  = ~A298 & A269;
  assign \new_[96700]_  = \new_[96699]_  & \new_[96696]_ ;
  assign \new_[96703]_  = ~A300 & A299;
  assign \new_[96706]_  = A302 & ~A301;
  assign \new_[96707]_  = \new_[96706]_  & \new_[96703]_ ;
  assign \new_[96708]_  = \new_[96707]_  & \new_[96700]_ ;
  assign \new_[96711]_  = ~A168 & A170;
  assign \new_[96714]_  = ~A200 & A199;
  assign \new_[96715]_  = \new_[96714]_  & \new_[96711]_ ;
  assign \new_[96718]_  = ~A202 & ~A201;
  assign \new_[96721]_  = ~A265 & A203;
  assign \new_[96722]_  = \new_[96721]_  & \new_[96718]_ ;
  assign \new_[96723]_  = \new_[96722]_  & \new_[96715]_ ;
  assign \new_[96726]_  = A267 & A266;
  assign \new_[96729]_  = A298 & A268;
  assign \new_[96730]_  = \new_[96729]_  & \new_[96726]_ ;
  assign \new_[96733]_  = ~A300 & ~A299;
  assign \new_[96736]_  = A302 & ~A301;
  assign \new_[96737]_  = \new_[96736]_  & \new_[96733]_ ;
  assign \new_[96738]_  = \new_[96737]_  & \new_[96730]_ ;
  assign \new_[96741]_  = ~A168 & A170;
  assign \new_[96744]_  = ~A200 & A199;
  assign \new_[96745]_  = \new_[96744]_  & \new_[96741]_ ;
  assign \new_[96748]_  = ~A202 & ~A201;
  assign \new_[96751]_  = ~A265 & A203;
  assign \new_[96752]_  = \new_[96751]_  & \new_[96748]_ ;
  assign \new_[96753]_  = \new_[96752]_  & \new_[96745]_ ;
  assign \new_[96756]_  = A267 & A266;
  assign \new_[96759]_  = ~A298 & A268;
  assign \new_[96760]_  = \new_[96759]_  & \new_[96756]_ ;
  assign \new_[96763]_  = ~A300 & A299;
  assign \new_[96766]_  = A302 & ~A301;
  assign \new_[96767]_  = \new_[96766]_  & \new_[96763]_ ;
  assign \new_[96768]_  = \new_[96767]_  & \new_[96760]_ ;
  assign \new_[96771]_  = ~A168 & A170;
  assign \new_[96774]_  = ~A200 & A199;
  assign \new_[96775]_  = \new_[96774]_  & \new_[96771]_ ;
  assign \new_[96778]_  = ~A202 & ~A201;
  assign \new_[96781]_  = ~A265 & A203;
  assign \new_[96782]_  = \new_[96781]_  & \new_[96778]_ ;
  assign \new_[96783]_  = \new_[96782]_  & \new_[96775]_ ;
  assign \new_[96786]_  = A267 & A266;
  assign \new_[96789]_  = A298 & ~A269;
  assign \new_[96790]_  = \new_[96789]_  & \new_[96786]_ ;
  assign \new_[96793]_  = ~A300 & ~A299;
  assign \new_[96796]_  = A302 & ~A301;
  assign \new_[96797]_  = \new_[96796]_  & \new_[96793]_ ;
  assign \new_[96798]_  = \new_[96797]_  & \new_[96790]_ ;
  assign \new_[96801]_  = ~A168 & A170;
  assign \new_[96804]_  = ~A200 & A199;
  assign \new_[96805]_  = \new_[96804]_  & \new_[96801]_ ;
  assign \new_[96808]_  = ~A202 & ~A201;
  assign \new_[96811]_  = ~A265 & A203;
  assign \new_[96812]_  = \new_[96811]_  & \new_[96808]_ ;
  assign \new_[96813]_  = \new_[96812]_  & \new_[96805]_ ;
  assign \new_[96816]_  = A267 & A266;
  assign \new_[96819]_  = ~A298 & ~A269;
  assign \new_[96820]_  = \new_[96819]_  & \new_[96816]_ ;
  assign \new_[96823]_  = ~A300 & A299;
  assign \new_[96826]_  = A302 & ~A301;
  assign \new_[96827]_  = \new_[96826]_  & \new_[96823]_ ;
  assign \new_[96828]_  = \new_[96827]_  & \new_[96820]_ ;
  assign \new_[96831]_  = ~A168 & A170;
  assign \new_[96834]_  = ~A200 & A199;
  assign \new_[96835]_  = \new_[96834]_  & \new_[96831]_ ;
  assign \new_[96838]_  = ~A202 & ~A201;
  assign \new_[96841]_  = ~A265 & A203;
  assign \new_[96842]_  = \new_[96841]_  & \new_[96838]_ ;
  assign \new_[96843]_  = \new_[96842]_  & \new_[96835]_ ;
  assign \new_[96846]_  = ~A267 & A266;
  assign \new_[96849]_  = A269 & ~A268;
  assign \new_[96850]_  = \new_[96849]_  & \new_[96846]_ ;
  assign \new_[96853]_  = ~A299 & A298;
  assign \new_[96856]_  = A301 & A300;
  assign \new_[96857]_  = \new_[96856]_  & \new_[96853]_ ;
  assign \new_[96858]_  = \new_[96857]_  & \new_[96850]_ ;
  assign \new_[96861]_  = ~A168 & A170;
  assign \new_[96864]_  = ~A200 & A199;
  assign \new_[96865]_  = \new_[96864]_  & \new_[96861]_ ;
  assign \new_[96868]_  = ~A202 & ~A201;
  assign \new_[96871]_  = ~A265 & A203;
  assign \new_[96872]_  = \new_[96871]_  & \new_[96868]_ ;
  assign \new_[96873]_  = \new_[96872]_  & \new_[96865]_ ;
  assign \new_[96876]_  = ~A267 & A266;
  assign \new_[96879]_  = A269 & ~A268;
  assign \new_[96880]_  = \new_[96879]_  & \new_[96876]_ ;
  assign \new_[96883]_  = ~A299 & A298;
  assign \new_[96886]_  = ~A302 & A300;
  assign \new_[96887]_  = \new_[96886]_  & \new_[96883]_ ;
  assign \new_[96888]_  = \new_[96887]_  & \new_[96880]_ ;
  assign \new_[96891]_  = ~A168 & A170;
  assign \new_[96894]_  = ~A200 & A199;
  assign \new_[96895]_  = \new_[96894]_  & \new_[96891]_ ;
  assign \new_[96898]_  = ~A202 & ~A201;
  assign \new_[96901]_  = ~A265 & A203;
  assign \new_[96902]_  = \new_[96901]_  & \new_[96898]_ ;
  assign \new_[96903]_  = \new_[96902]_  & \new_[96895]_ ;
  assign \new_[96906]_  = ~A267 & A266;
  assign \new_[96909]_  = A269 & ~A268;
  assign \new_[96910]_  = \new_[96909]_  & \new_[96906]_ ;
  assign \new_[96913]_  = A299 & ~A298;
  assign \new_[96916]_  = A301 & A300;
  assign \new_[96917]_  = \new_[96916]_  & \new_[96913]_ ;
  assign \new_[96918]_  = \new_[96917]_  & \new_[96910]_ ;
  assign \new_[96921]_  = ~A168 & A170;
  assign \new_[96924]_  = ~A200 & A199;
  assign \new_[96925]_  = \new_[96924]_  & \new_[96921]_ ;
  assign \new_[96928]_  = ~A202 & ~A201;
  assign \new_[96931]_  = ~A265 & A203;
  assign \new_[96932]_  = \new_[96931]_  & \new_[96928]_ ;
  assign \new_[96933]_  = \new_[96932]_  & \new_[96925]_ ;
  assign \new_[96936]_  = ~A267 & A266;
  assign \new_[96939]_  = A269 & ~A268;
  assign \new_[96940]_  = \new_[96939]_  & \new_[96936]_ ;
  assign \new_[96943]_  = A299 & ~A298;
  assign \new_[96946]_  = ~A302 & A300;
  assign \new_[96947]_  = \new_[96946]_  & \new_[96943]_ ;
  assign \new_[96948]_  = \new_[96947]_  & \new_[96940]_ ;
  assign \new_[96951]_  = ~A168 & A170;
  assign \new_[96954]_  = ~A200 & A199;
  assign \new_[96955]_  = \new_[96954]_  & \new_[96951]_ ;
  assign \new_[96958]_  = ~A202 & ~A201;
  assign \new_[96961]_  = A265 & A203;
  assign \new_[96962]_  = \new_[96961]_  & \new_[96958]_ ;
  assign \new_[96963]_  = \new_[96962]_  & \new_[96955]_ ;
  assign \new_[96966]_  = A267 & ~A266;
  assign \new_[96969]_  = A298 & A268;
  assign \new_[96970]_  = \new_[96969]_  & \new_[96966]_ ;
  assign \new_[96973]_  = ~A300 & ~A299;
  assign \new_[96976]_  = A302 & ~A301;
  assign \new_[96977]_  = \new_[96976]_  & \new_[96973]_ ;
  assign \new_[96978]_  = \new_[96977]_  & \new_[96970]_ ;
  assign \new_[96981]_  = ~A168 & A170;
  assign \new_[96984]_  = ~A200 & A199;
  assign \new_[96985]_  = \new_[96984]_  & \new_[96981]_ ;
  assign \new_[96988]_  = ~A202 & ~A201;
  assign \new_[96991]_  = A265 & A203;
  assign \new_[96992]_  = \new_[96991]_  & \new_[96988]_ ;
  assign \new_[96993]_  = \new_[96992]_  & \new_[96985]_ ;
  assign \new_[96996]_  = A267 & ~A266;
  assign \new_[96999]_  = ~A298 & A268;
  assign \new_[97000]_  = \new_[96999]_  & \new_[96996]_ ;
  assign \new_[97003]_  = ~A300 & A299;
  assign \new_[97006]_  = A302 & ~A301;
  assign \new_[97007]_  = \new_[97006]_  & \new_[97003]_ ;
  assign \new_[97008]_  = \new_[97007]_  & \new_[97000]_ ;
  assign \new_[97011]_  = ~A168 & A170;
  assign \new_[97014]_  = ~A200 & A199;
  assign \new_[97015]_  = \new_[97014]_  & \new_[97011]_ ;
  assign \new_[97018]_  = ~A202 & ~A201;
  assign \new_[97021]_  = A265 & A203;
  assign \new_[97022]_  = \new_[97021]_  & \new_[97018]_ ;
  assign \new_[97023]_  = \new_[97022]_  & \new_[97015]_ ;
  assign \new_[97026]_  = A267 & ~A266;
  assign \new_[97029]_  = A298 & ~A269;
  assign \new_[97030]_  = \new_[97029]_  & \new_[97026]_ ;
  assign \new_[97033]_  = ~A300 & ~A299;
  assign \new_[97036]_  = A302 & ~A301;
  assign \new_[97037]_  = \new_[97036]_  & \new_[97033]_ ;
  assign \new_[97038]_  = \new_[97037]_  & \new_[97030]_ ;
  assign \new_[97041]_  = ~A168 & A170;
  assign \new_[97044]_  = ~A200 & A199;
  assign \new_[97045]_  = \new_[97044]_  & \new_[97041]_ ;
  assign \new_[97048]_  = ~A202 & ~A201;
  assign \new_[97051]_  = A265 & A203;
  assign \new_[97052]_  = \new_[97051]_  & \new_[97048]_ ;
  assign \new_[97053]_  = \new_[97052]_  & \new_[97045]_ ;
  assign \new_[97056]_  = A267 & ~A266;
  assign \new_[97059]_  = ~A298 & ~A269;
  assign \new_[97060]_  = \new_[97059]_  & \new_[97056]_ ;
  assign \new_[97063]_  = ~A300 & A299;
  assign \new_[97066]_  = A302 & ~A301;
  assign \new_[97067]_  = \new_[97066]_  & \new_[97063]_ ;
  assign \new_[97068]_  = \new_[97067]_  & \new_[97060]_ ;
  assign \new_[97071]_  = ~A168 & A170;
  assign \new_[97074]_  = ~A200 & A199;
  assign \new_[97075]_  = \new_[97074]_  & \new_[97071]_ ;
  assign \new_[97078]_  = ~A202 & ~A201;
  assign \new_[97081]_  = A265 & A203;
  assign \new_[97082]_  = \new_[97081]_  & \new_[97078]_ ;
  assign \new_[97083]_  = \new_[97082]_  & \new_[97075]_ ;
  assign \new_[97086]_  = ~A267 & ~A266;
  assign \new_[97089]_  = A269 & ~A268;
  assign \new_[97090]_  = \new_[97089]_  & \new_[97086]_ ;
  assign \new_[97093]_  = ~A299 & A298;
  assign \new_[97096]_  = A301 & A300;
  assign \new_[97097]_  = \new_[97096]_  & \new_[97093]_ ;
  assign \new_[97098]_  = \new_[97097]_  & \new_[97090]_ ;
  assign \new_[97101]_  = ~A168 & A170;
  assign \new_[97104]_  = ~A200 & A199;
  assign \new_[97105]_  = \new_[97104]_  & \new_[97101]_ ;
  assign \new_[97108]_  = ~A202 & ~A201;
  assign \new_[97111]_  = A265 & A203;
  assign \new_[97112]_  = \new_[97111]_  & \new_[97108]_ ;
  assign \new_[97113]_  = \new_[97112]_  & \new_[97105]_ ;
  assign \new_[97116]_  = ~A267 & ~A266;
  assign \new_[97119]_  = A269 & ~A268;
  assign \new_[97120]_  = \new_[97119]_  & \new_[97116]_ ;
  assign \new_[97123]_  = ~A299 & A298;
  assign \new_[97126]_  = ~A302 & A300;
  assign \new_[97127]_  = \new_[97126]_  & \new_[97123]_ ;
  assign \new_[97128]_  = \new_[97127]_  & \new_[97120]_ ;
  assign \new_[97131]_  = ~A168 & A170;
  assign \new_[97134]_  = ~A200 & A199;
  assign \new_[97135]_  = \new_[97134]_  & \new_[97131]_ ;
  assign \new_[97138]_  = ~A202 & ~A201;
  assign \new_[97141]_  = A265 & A203;
  assign \new_[97142]_  = \new_[97141]_  & \new_[97138]_ ;
  assign \new_[97143]_  = \new_[97142]_  & \new_[97135]_ ;
  assign \new_[97146]_  = ~A267 & ~A266;
  assign \new_[97149]_  = A269 & ~A268;
  assign \new_[97150]_  = \new_[97149]_  & \new_[97146]_ ;
  assign \new_[97153]_  = A299 & ~A298;
  assign \new_[97156]_  = A301 & A300;
  assign \new_[97157]_  = \new_[97156]_  & \new_[97153]_ ;
  assign \new_[97158]_  = \new_[97157]_  & \new_[97150]_ ;
  assign \new_[97161]_  = ~A168 & A170;
  assign \new_[97164]_  = ~A200 & A199;
  assign \new_[97165]_  = \new_[97164]_  & \new_[97161]_ ;
  assign \new_[97168]_  = ~A202 & ~A201;
  assign \new_[97171]_  = A265 & A203;
  assign \new_[97172]_  = \new_[97171]_  & \new_[97168]_ ;
  assign \new_[97173]_  = \new_[97172]_  & \new_[97165]_ ;
  assign \new_[97176]_  = ~A267 & ~A266;
  assign \new_[97179]_  = A269 & ~A268;
  assign \new_[97180]_  = \new_[97179]_  & \new_[97176]_ ;
  assign \new_[97183]_  = A299 & ~A298;
  assign \new_[97186]_  = ~A302 & A300;
  assign \new_[97187]_  = \new_[97186]_  & \new_[97183]_ ;
  assign \new_[97188]_  = \new_[97187]_  & \new_[97180]_ ;
  assign \new_[97191]_  = ~A168 & A169;
  assign \new_[97194]_  = A200 & ~A199;
  assign \new_[97195]_  = \new_[97194]_  & \new_[97191]_ ;
  assign \new_[97198]_  = A202 & A201;
  assign \new_[97201]_  = A266 & ~A265;
  assign \new_[97202]_  = \new_[97201]_  & \new_[97198]_ ;
  assign \new_[97203]_  = \new_[97202]_  & \new_[97195]_ ;
  assign \new_[97206]_  = ~A268 & ~A267;
  assign \new_[97209]_  = A298 & A269;
  assign \new_[97210]_  = \new_[97209]_  & \new_[97206]_ ;
  assign \new_[97213]_  = ~A300 & ~A299;
  assign \new_[97216]_  = A302 & ~A301;
  assign \new_[97217]_  = \new_[97216]_  & \new_[97213]_ ;
  assign \new_[97218]_  = \new_[97217]_  & \new_[97210]_ ;
  assign \new_[97221]_  = ~A168 & A169;
  assign \new_[97224]_  = A200 & ~A199;
  assign \new_[97225]_  = \new_[97224]_  & \new_[97221]_ ;
  assign \new_[97228]_  = A202 & A201;
  assign \new_[97231]_  = A266 & ~A265;
  assign \new_[97232]_  = \new_[97231]_  & \new_[97228]_ ;
  assign \new_[97233]_  = \new_[97232]_  & \new_[97225]_ ;
  assign \new_[97236]_  = ~A268 & ~A267;
  assign \new_[97239]_  = ~A298 & A269;
  assign \new_[97240]_  = \new_[97239]_  & \new_[97236]_ ;
  assign \new_[97243]_  = ~A300 & A299;
  assign \new_[97246]_  = A302 & ~A301;
  assign \new_[97247]_  = \new_[97246]_  & \new_[97243]_ ;
  assign \new_[97248]_  = \new_[97247]_  & \new_[97240]_ ;
  assign \new_[97251]_  = ~A168 & A169;
  assign \new_[97254]_  = A200 & ~A199;
  assign \new_[97255]_  = \new_[97254]_  & \new_[97251]_ ;
  assign \new_[97258]_  = A202 & A201;
  assign \new_[97261]_  = ~A266 & A265;
  assign \new_[97262]_  = \new_[97261]_  & \new_[97258]_ ;
  assign \new_[97263]_  = \new_[97262]_  & \new_[97255]_ ;
  assign \new_[97266]_  = ~A268 & ~A267;
  assign \new_[97269]_  = A298 & A269;
  assign \new_[97270]_  = \new_[97269]_  & \new_[97266]_ ;
  assign \new_[97273]_  = ~A300 & ~A299;
  assign \new_[97276]_  = A302 & ~A301;
  assign \new_[97277]_  = \new_[97276]_  & \new_[97273]_ ;
  assign \new_[97278]_  = \new_[97277]_  & \new_[97270]_ ;
  assign \new_[97281]_  = ~A168 & A169;
  assign \new_[97284]_  = A200 & ~A199;
  assign \new_[97285]_  = \new_[97284]_  & \new_[97281]_ ;
  assign \new_[97288]_  = A202 & A201;
  assign \new_[97291]_  = ~A266 & A265;
  assign \new_[97292]_  = \new_[97291]_  & \new_[97288]_ ;
  assign \new_[97293]_  = \new_[97292]_  & \new_[97285]_ ;
  assign \new_[97296]_  = ~A268 & ~A267;
  assign \new_[97299]_  = ~A298 & A269;
  assign \new_[97300]_  = \new_[97299]_  & \new_[97296]_ ;
  assign \new_[97303]_  = ~A300 & A299;
  assign \new_[97306]_  = A302 & ~A301;
  assign \new_[97307]_  = \new_[97306]_  & \new_[97303]_ ;
  assign \new_[97308]_  = \new_[97307]_  & \new_[97300]_ ;
  assign \new_[97311]_  = ~A168 & A169;
  assign \new_[97314]_  = A200 & ~A199;
  assign \new_[97315]_  = \new_[97314]_  & \new_[97311]_ ;
  assign \new_[97318]_  = ~A203 & A201;
  assign \new_[97321]_  = A266 & ~A265;
  assign \new_[97322]_  = \new_[97321]_  & \new_[97318]_ ;
  assign \new_[97323]_  = \new_[97322]_  & \new_[97315]_ ;
  assign \new_[97326]_  = ~A268 & ~A267;
  assign \new_[97329]_  = A298 & A269;
  assign \new_[97330]_  = \new_[97329]_  & \new_[97326]_ ;
  assign \new_[97333]_  = ~A300 & ~A299;
  assign \new_[97336]_  = A302 & ~A301;
  assign \new_[97337]_  = \new_[97336]_  & \new_[97333]_ ;
  assign \new_[97338]_  = \new_[97337]_  & \new_[97330]_ ;
  assign \new_[97341]_  = ~A168 & A169;
  assign \new_[97344]_  = A200 & ~A199;
  assign \new_[97345]_  = \new_[97344]_  & \new_[97341]_ ;
  assign \new_[97348]_  = ~A203 & A201;
  assign \new_[97351]_  = A266 & ~A265;
  assign \new_[97352]_  = \new_[97351]_  & \new_[97348]_ ;
  assign \new_[97353]_  = \new_[97352]_  & \new_[97345]_ ;
  assign \new_[97356]_  = ~A268 & ~A267;
  assign \new_[97359]_  = ~A298 & A269;
  assign \new_[97360]_  = \new_[97359]_  & \new_[97356]_ ;
  assign \new_[97363]_  = ~A300 & A299;
  assign \new_[97366]_  = A302 & ~A301;
  assign \new_[97367]_  = \new_[97366]_  & \new_[97363]_ ;
  assign \new_[97368]_  = \new_[97367]_  & \new_[97360]_ ;
  assign \new_[97371]_  = ~A168 & A169;
  assign \new_[97374]_  = A200 & ~A199;
  assign \new_[97375]_  = \new_[97374]_  & \new_[97371]_ ;
  assign \new_[97378]_  = ~A203 & A201;
  assign \new_[97381]_  = ~A266 & A265;
  assign \new_[97382]_  = \new_[97381]_  & \new_[97378]_ ;
  assign \new_[97383]_  = \new_[97382]_  & \new_[97375]_ ;
  assign \new_[97386]_  = ~A268 & ~A267;
  assign \new_[97389]_  = A298 & A269;
  assign \new_[97390]_  = \new_[97389]_  & \new_[97386]_ ;
  assign \new_[97393]_  = ~A300 & ~A299;
  assign \new_[97396]_  = A302 & ~A301;
  assign \new_[97397]_  = \new_[97396]_  & \new_[97393]_ ;
  assign \new_[97398]_  = \new_[97397]_  & \new_[97390]_ ;
  assign \new_[97401]_  = ~A168 & A169;
  assign \new_[97404]_  = A200 & ~A199;
  assign \new_[97405]_  = \new_[97404]_  & \new_[97401]_ ;
  assign \new_[97408]_  = ~A203 & A201;
  assign \new_[97411]_  = ~A266 & A265;
  assign \new_[97412]_  = \new_[97411]_  & \new_[97408]_ ;
  assign \new_[97413]_  = \new_[97412]_  & \new_[97405]_ ;
  assign \new_[97416]_  = ~A268 & ~A267;
  assign \new_[97419]_  = ~A298 & A269;
  assign \new_[97420]_  = \new_[97419]_  & \new_[97416]_ ;
  assign \new_[97423]_  = ~A300 & A299;
  assign \new_[97426]_  = A302 & ~A301;
  assign \new_[97427]_  = \new_[97426]_  & \new_[97423]_ ;
  assign \new_[97428]_  = \new_[97427]_  & \new_[97420]_ ;
  assign \new_[97431]_  = ~A168 & A169;
  assign \new_[97434]_  = A200 & ~A199;
  assign \new_[97435]_  = \new_[97434]_  & \new_[97431]_ ;
  assign \new_[97438]_  = ~A202 & ~A201;
  assign \new_[97441]_  = ~A265 & A203;
  assign \new_[97442]_  = \new_[97441]_  & \new_[97438]_ ;
  assign \new_[97443]_  = \new_[97442]_  & \new_[97435]_ ;
  assign \new_[97446]_  = A267 & A266;
  assign \new_[97449]_  = A298 & A268;
  assign \new_[97450]_  = \new_[97449]_  & \new_[97446]_ ;
  assign \new_[97453]_  = ~A300 & ~A299;
  assign \new_[97456]_  = A302 & ~A301;
  assign \new_[97457]_  = \new_[97456]_  & \new_[97453]_ ;
  assign \new_[97458]_  = \new_[97457]_  & \new_[97450]_ ;
  assign \new_[97461]_  = ~A168 & A169;
  assign \new_[97464]_  = A200 & ~A199;
  assign \new_[97465]_  = \new_[97464]_  & \new_[97461]_ ;
  assign \new_[97468]_  = ~A202 & ~A201;
  assign \new_[97471]_  = ~A265 & A203;
  assign \new_[97472]_  = \new_[97471]_  & \new_[97468]_ ;
  assign \new_[97473]_  = \new_[97472]_  & \new_[97465]_ ;
  assign \new_[97476]_  = A267 & A266;
  assign \new_[97479]_  = ~A298 & A268;
  assign \new_[97480]_  = \new_[97479]_  & \new_[97476]_ ;
  assign \new_[97483]_  = ~A300 & A299;
  assign \new_[97486]_  = A302 & ~A301;
  assign \new_[97487]_  = \new_[97486]_  & \new_[97483]_ ;
  assign \new_[97488]_  = \new_[97487]_  & \new_[97480]_ ;
  assign \new_[97491]_  = ~A168 & A169;
  assign \new_[97494]_  = A200 & ~A199;
  assign \new_[97495]_  = \new_[97494]_  & \new_[97491]_ ;
  assign \new_[97498]_  = ~A202 & ~A201;
  assign \new_[97501]_  = ~A265 & A203;
  assign \new_[97502]_  = \new_[97501]_  & \new_[97498]_ ;
  assign \new_[97503]_  = \new_[97502]_  & \new_[97495]_ ;
  assign \new_[97506]_  = A267 & A266;
  assign \new_[97509]_  = A298 & ~A269;
  assign \new_[97510]_  = \new_[97509]_  & \new_[97506]_ ;
  assign \new_[97513]_  = ~A300 & ~A299;
  assign \new_[97516]_  = A302 & ~A301;
  assign \new_[97517]_  = \new_[97516]_  & \new_[97513]_ ;
  assign \new_[97518]_  = \new_[97517]_  & \new_[97510]_ ;
  assign \new_[97521]_  = ~A168 & A169;
  assign \new_[97524]_  = A200 & ~A199;
  assign \new_[97525]_  = \new_[97524]_  & \new_[97521]_ ;
  assign \new_[97528]_  = ~A202 & ~A201;
  assign \new_[97531]_  = ~A265 & A203;
  assign \new_[97532]_  = \new_[97531]_  & \new_[97528]_ ;
  assign \new_[97533]_  = \new_[97532]_  & \new_[97525]_ ;
  assign \new_[97536]_  = A267 & A266;
  assign \new_[97539]_  = ~A298 & ~A269;
  assign \new_[97540]_  = \new_[97539]_  & \new_[97536]_ ;
  assign \new_[97543]_  = ~A300 & A299;
  assign \new_[97546]_  = A302 & ~A301;
  assign \new_[97547]_  = \new_[97546]_  & \new_[97543]_ ;
  assign \new_[97548]_  = \new_[97547]_  & \new_[97540]_ ;
  assign \new_[97551]_  = ~A168 & A169;
  assign \new_[97554]_  = A200 & ~A199;
  assign \new_[97555]_  = \new_[97554]_  & \new_[97551]_ ;
  assign \new_[97558]_  = ~A202 & ~A201;
  assign \new_[97561]_  = ~A265 & A203;
  assign \new_[97562]_  = \new_[97561]_  & \new_[97558]_ ;
  assign \new_[97563]_  = \new_[97562]_  & \new_[97555]_ ;
  assign \new_[97566]_  = ~A267 & A266;
  assign \new_[97569]_  = A269 & ~A268;
  assign \new_[97570]_  = \new_[97569]_  & \new_[97566]_ ;
  assign \new_[97573]_  = ~A299 & A298;
  assign \new_[97576]_  = A301 & A300;
  assign \new_[97577]_  = \new_[97576]_  & \new_[97573]_ ;
  assign \new_[97578]_  = \new_[97577]_  & \new_[97570]_ ;
  assign \new_[97581]_  = ~A168 & A169;
  assign \new_[97584]_  = A200 & ~A199;
  assign \new_[97585]_  = \new_[97584]_  & \new_[97581]_ ;
  assign \new_[97588]_  = ~A202 & ~A201;
  assign \new_[97591]_  = ~A265 & A203;
  assign \new_[97592]_  = \new_[97591]_  & \new_[97588]_ ;
  assign \new_[97593]_  = \new_[97592]_  & \new_[97585]_ ;
  assign \new_[97596]_  = ~A267 & A266;
  assign \new_[97599]_  = A269 & ~A268;
  assign \new_[97600]_  = \new_[97599]_  & \new_[97596]_ ;
  assign \new_[97603]_  = ~A299 & A298;
  assign \new_[97606]_  = ~A302 & A300;
  assign \new_[97607]_  = \new_[97606]_  & \new_[97603]_ ;
  assign \new_[97608]_  = \new_[97607]_  & \new_[97600]_ ;
  assign \new_[97611]_  = ~A168 & A169;
  assign \new_[97614]_  = A200 & ~A199;
  assign \new_[97615]_  = \new_[97614]_  & \new_[97611]_ ;
  assign \new_[97618]_  = ~A202 & ~A201;
  assign \new_[97621]_  = ~A265 & A203;
  assign \new_[97622]_  = \new_[97621]_  & \new_[97618]_ ;
  assign \new_[97623]_  = \new_[97622]_  & \new_[97615]_ ;
  assign \new_[97626]_  = ~A267 & A266;
  assign \new_[97629]_  = A269 & ~A268;
  assign \new_[97630]_  = \new_[97629]_  & \new_[97626]_ ;
  assign \new_[97633]_  = A299 & ~A298;
  assign \new_[97636]_  = A301 & A300;
  assign \new_[97637]_  = \new_[97636]_  & \new_[97633]_ ;
  assign \new_[97638]_  = \new_[97637]_  & \new_[97630]_ ;
  assign \new_[97641]_  = ~A168 & A169;
  assign \new_[97644]_  = A200 & ~A199;
  assign \new_[97645]_  = \new_[97644]_  & \new_[97641]_ ;
  assign \new_[97648]_  = ~A202 & ~A201;
  assign \new_[97651]_  = ~A265 & A203;
  assign \new_[97652]_  = \new_[97651]_  & \new_[97648]_ ;
  assign \new_[97653]_  = \new_[97652]_  & \new_[97645]_ ;
  assign \new_[97656]_  = ~A267 & A266;
  assign \new_[97659]_  = A269 & ~A268;
  assign \new_[97660]_  = \new_[97659]_  & \new_[97656]_ ;
  assign \new_[97663]_  = A299 & ~A298;
  assign \new_[97666]_  = ~A302 & A300;
  assign \new_[97667]_  = \new_[97666]_  & \new_[97663]_ ;
  assign \new_[97668]_  = \new_[97667]_  & \new_[97660]_ ;
  assign \new_[97671]_  = ~A168 & A169;
  assign \new_[97674]_  = A200 & ~A199;
  assign \new_[97675]_  = \new_[97674]_  & \new_[97671]_ ;
  assign \new_[97678]_  = ~A202 & ~A201;
  assign \new_[97681]_  = A265 & A203;
  assign \new_[97682]_  = \new_[97681]_  & \new_[97678]_ ;
  assign \new_[97683]_  = \new_[97682]_  & \new_[97675]_ ;
  assign \new_[97686]_  = A267 & ~A266;
  assign \new_[97689]_  = A298 & A268;
  assign \new_[97690]_  = \new_[97689]_  & \new_[97686]_ ;
  assign \new_[97693]_  = ~A300 & ~A299;
  assign \new_[97696]_  = A302 & ~A301;
  assign \new_[97697]_  = \new_[97696]_  & \new_[97693]_ ;
  assign \new_[97698]_  = \new_[97697]_  & \new_[97690]_ ;
  assign \new_[97701]_  = ~A168 & A169;
  assign \new_[97704]_  = A200 & ~A199;
  assign \new_[97705]_  = \new_[97704]_  & \new_[97701]_ ;
  assign \new_[97708]_  = ~A202 & ~A201;
  assign \new_[97711]_  = A265 & A203;
  assign \new_[97712]_  = \new_[97711]_  & \new_[97708]_ ;
  assign \new_[97713]_  = \new_[97712]_  & \new_[97705]_ ;
  assign \new_[97716]_  = A267 & ~A266;
  assign \new_[97719]_  = ~A298 & A268;
  assign \new_[97720]_  = \new_[97719]_  & \new_[97716]_ ;
  assign \new_[97723]_  = ~A300 & A299;
  assign \new_[97726]_  = A302 & ~A301;
  assign \new_[97727]_  = \new_[97726]_  & \new_[97723]_ ;
  assign \new_[97728]_  = \new_[97727]_  & \new_[97720]_ ;
  assign \new_[97731]_  = ~A168 & A169;
  assign \new_[97734]_  = A200 & ~A199;
  assign \new_[97735]_  = \new_[97734]_  & \new_[97731]_ ;
  assign \new_[97738]_  = ~A202 & ~A201;
  assign \new_[97741]_  = A265 & A203;
  assign \new_[97742]_  = \new_[97741]_  & \new_[97738]_ ;
  assign \new_[97743]_  = \new_[97742]_  & \new_[97735]_ ;
  assign \new_[97746]_  = A267 & ~A266;
  assign \new_[97749]_  = A298 & ~A269;
  assign \new_[97750]_  = \new_[97749]_  & \new_[97746]_ ;
  assign \new_[97753]_  = ~A300 & ~A299;
  assign \new_[97756]_  = A302 & ~A301;
  assign \new_[97757]_  = \new_[97756]_  & \new_[97753]_ ;
  assign \new_[97758]_  = \new_[97757]_  & \new_[97750]_ ;
  assign \new_[97761]_  = ~A168 & A169;
  assign \new_[97764]_  = A200 & ~A199;
  assign \new_[97765]_  = \new_[97764]_  & \new_[97761]_ ;
  assign \new_[97768]_  = ~A202 & ~A201;
  assign \new_[97771]_  = A265 & A203;
  assign \new_[97772]_  = \new_[97771]_  & \new_[97768]_ ;
  assign \new_[97773]_  = \new_[97772]_  & \new_[97765]_ ;
  assign \new_[97776]_  = A267 & ~A266;
  assign \new_[97779]_  = ~A298 & ~A269;
  assign \new_[97780]_  = \new_[97779]_  & \new_[97776]_ ;
  assign \new_[97783]_  = ~A300 & A299;
  assign \new_[97786]_  = A302 & ~A301;
  assign \new_[97787]_  = \new_[97786]_  & \new_[97783]_ ;
  assign \new_[97788]_  = \new_[97787]_  & \new_[97780]_ ;
  assign \new_[97791]_  = ~A168 & A169;
  assign \new_[97794]_  = A200 & ~A199;
  assign \new_[97795]_  = \new_[97794]_  & \new_[97791]_ ;
  assign \new_[97798]_  = ~A202 & ~A201;
  assign \new_[97801]_  = A265 & A203;
  assign \new_[97802]_  = \new_[97801]_  & \new_[97798]_ ;
  assign \new_[97803]_  = \new_[97802]_  & \new_[97795]_ ;
  assign \new_[97806]_  = ~A267 & ~A266;
  assign \new_[97809]_  = A269 & ~A268;
  assign \new_[97810]_  = \new_[97809]_  & \new_[97806]_ ;
  assign \new_[97813]_  = ~A299 & A298;
  assign \new_[97816]_  = A301 & A300;
  assign \new_[97817]_  = \new_[97816]_  & \new_[97813]_ ;
  assign \new_[97818]_  = \new_[97817]_  & \new_[97810]_ ;
  assign \new_[97821]_  = ~A168 & A169;
  assign \new_[97824]_  = A200 & ~A199;
  assign \new_[97825]_  = \new_[97824]_  & \new_[97821]_ ;
  assign \new_[97828]_  = ~A202 & ~A201;
  assign \new_[97831]_  = A265 & A203;
  assign \new_[97832]_  = \new_[97831]_  & \new_[97828]_ ;
  assign \new_[97833]_  = \new_[97832]_  & \new_[97825]_ ;
  assign \new_[97836]_  = ~A267 & ~A266;
  assign \new_[97839]_  = A269 & ~A268;
  assign \new_[97840]_  = \new_[97839]_  & \new_[97836]_ ;
  assign \new_[97843]_  = ~A299 & A298;
  assign \new_[97846]_  = ~A302 & A300;
  assign \new_[97847]_  = \new_[97846]_  & \new_[97843]_ ;
  assign \new_[97848]_  = \new_[97847]_  & \new_[97840]_ ;
  assign \new_[97851]_  = ~A168 & A169;
  assign \new_[97854]_  = A200 & ~A199;
  assign \new_[97855]_  = \new_[97854]_  & \new_[97851]_ ;
  assign \new_[97858]_  = ~A202 & ~A201;
  assign \new_[97861]_  = A265 & A203;
  assign \new_[97862]_  = \new_[97861]_  & \new_[97858]_ ;
  assign \new_[97863]_  = \new_[97862]_  & \new_[97855]_ ;
  assign \new_[97866]_  = ~A267 & ~A266;
  assign \new_[97869]_  = A269 & ~A268;
  assign \new_[97870]_  = \new_[97869]_  & \new_[97866]_ ;
  assign \new_[97873]_  = A299 & ~A298;
  assign \new_[97876]_  = A301 & A300;
  assign \new_[97877]_  = \new_[97876]_  & \new_[97873]_ ;
  assign \new_[97878]_  = \new_[97877]_  & \new_[97870]_ ;
  assign \new_[97881]_  = ~A168 & A169;
  assign \new_[97884]_  = A200 & ~A199;
  assign \new_[97885]_  = \new_[97884]_  & \new_[97881]_ ;
  assign \new_[97888]_  = ~A202 & ~A201;
  assign \new_[97891]_  = A265 & A203;
  assign \new_[97892]_  = \new_[97891]_  & \new_[97888]_ ;
  assign \new_[97893]_  = \new_[97892]_  & \new_[97885]_ ;
  assign \new_[97896]_  = ~A267 & ~A266;
  assign \new_[97899]_  = A269 & ~A268;
  assign \new_[97900]_  = \new_[97899]_  & \new_[97896]_ ;
  assign \new_[97903]_  = A299 & ~A298;
  assign \new_[97906]_  = ~A302 & A300;
  assign \new_[97907]_  = \new_[97906]_  & \new_[97903]_ ;
  assign \new_[97908]_  = \new_[97907]_  & \new_[97900]_ ;
  assign \new_[97911]_  = ~A168 & A169;
  assign \new_[97914]_  = ~A200 & A199;
  assign \new_[97915]_  = \new_[97914]_  & \new_[97911]_ ;
  assign \new_[97918]_  = A202 & A201;
  assign \new_[97921]_  = A266 & ~A265;
  assign \new_[97922]_  = \new_[97921]_  & \new_[97918]_ ;
  assign \new_[97923]_  = \new_[97922]_  & \new_[97915]_ ;
  assign \new_[97926]_  = ~A268 & ~A267;
  assign \new_[97929]_  = A298 & A269;
  assign \new_[97930]_  = \new_[97929]_  & \new_[97926]_ ;
  assign \new_[97933]_  = ~A300 & ~A299;
  assign \new_[97936]_  = A302 & ~A301;
  assign \new_[97937]_  = \new_[97936]_  & \new_[97933]_ ;
  assign \new_[97938]_  = \new_[97937]_  & \new_[97930]_ ;
  assign \new_[97941]_  = ~A168 & A169;
  assign \new_[97944]_  = ~A200 & A199;
  assign \new_[97945]_  = \new_[97944]_  & \new_[97941]_ ;
  assign \new_[97948]_  = A202 & A201;
  assign \new_[97951]_  = A266 & ~A265;
  assign \new_[97952]_  = \new_[97951]_  & \new_[97948]_ ;
  assign \new_[97953]_  = \new_[97952]_  & \new_[97945]_ ;
  assign \new_[97956]_  = ~A268 & ~A267;
  assign \new_[97959]_  = ~A298 & A269;
  assign \new_[97960]_  = \new_[97959]_  & \new_[97956]_ ;
  assign \new_[97963]_  = ~A300 & A299;
  assign \new_[97966]_  = A302 & ~A301;
  assign \new_[97967]_  = \new_[97966]_  & \new_[97963]_ ;
  assign \new_[97968]_  = \new_[97967]_  & \new_[97960]_ ;
  assign \new_[97971]_  = ~A168 & A169;
  assign \new_[97974]_  = ~A200 & A199;
  assign \new_[97975]_  = \new_[97974]_  & \new_[97971]_ ;
  assign \new_[97978]_  = A202 & A201;
  assign \new_[97981]_  = ~A266 & A265;
  assign \new_[97982]_  = \new_[97981]_  & \new_[97978]_ ;
  assign \new_[97983]_  = \new_[97982]_  & \new_[97975]_ ;
  assign \new_[97986]_  = ~A268 & ~A267;
  assign \new_[97989]_  = A298 & A269;
  assign \new_[97990]_  = \new_[97989]_  & \new_[97986]_ ;
  assign \new_[97993]_  = ~A300 & ~A299;
  assign \new_[97996]_  = A302 & ~A301;
  assign \new_[97997]_  = \new_[97996]_  & \new_[97993]_ ;
  assign \new_[97998]_  = \new_[97997]_  & \new_[97990]_ ;
  assign \new_[98001]_  = ~A168 & A169;
  assign \new_[98004]_  = ~A200 & A199;
  assign \new_[98005]_  = \new_[98004]_  & \new_[98001]_ ;
  assign \new_[98008]_  = A202 & A201;
  assign \new_[98011]_  = ~A266 & A265;
  assign \new_[98012]_  = \new_[98011]_  & \new_[98008]_ ;
  assign \new_[98013]_  = \new_[98012]_  & \new_[98005]_ ;
  assign \new_[98016]_  = ~A268 & ~A267;
  assign \new_[98019]_  = ~A298 & A269;
  assign \new_[98020]_  = \new_[98019]_  & \new_[98016]_ ;
  assign \new_[98023]_  = ~A300 & A299;
  assign \new_[98026]_  = A302 & ~A301;
  assign \new_[98027]_  = \new_[98026]_  & \new_[98023]_ ;
  assign \new_[98028]_  = \new_[98027]_  & \new_[98020]_ ;
  assign \new_[98031]_  = ~A168 & A169;
  assign \new_[98034]_  = ~A200 & A199;
  assign \new_[98035]_  = \new_[98034]_  & \new_[98031]_ ;
  assign \new_[98038]_  = ~A203 & A201;
  assign \new_[98041]_  = A266 & ~A265;
  assign \new_[98042]_  = \new_[98041]_  & \new_[98038]_ ;
  assign \new_[98043]_  = \new_[98042]_  & \new_[98035]_ ;
  assign \new_[98046]_  = ~A268 & ~A267;
  assign \new_[98049]_  = A298 & A269;
  assign \new_[98050]_  = \new_[98049]_  & \new_[98046]_ ;
  assign \new_[98053]_  = ~A300 & ~A299;
  assign \new_[98056]_  = A302 & ~A301;
  assign \new_[98057]_  = \new_[98056]_  & \new_[98053]_ ;
  assign \new_[98058]_  = \new_[98057]_  & \new_[98050]_ ;
  assign \new_[98061]_  = ~A168 & A169;
  assign \new_[98064]_  = ~A200 & A199;
  assign \new_[98065]_  = \new_[98064]_  & \new_[98061]_ ;
  assign \new_[98068]_  = ~A203 & A201;
  assign \new_[98071]_  = A266 & ~A265;
  assign \new_[98072]_  = \new_[98071]_  & \new_[98068]_ ;
  assign \new_[98073]_  = \new_[98072]_  & \new_[98065]_ ;
  assign \new_[98076]_  = ~A268 & ~A267;
  assign \new_[98079]_  = ~A298 & A269;
  assign \new_[98080]_  = \new_[98079]_  & \new_[98076]_ ;
  assign \new_[98083]_  = ~A300 & A299;
  assign \new_[98086]_  = A302 & ~A301;
  assign \new_[98087]_  = \new_[98086]_  & \new_[98083]_ ;
  assign \new_[98088]_  = \new_[98087]_  & \new_[98080]_ ;
  assign \new_[98091]_  = ~A168 & A169;
  assign \new_[98094]_  = ~A200 & A199;
  assign \new_[98095]_  = \new_[98094]_  & \new_[98091]_ ;
  assign \new_[98098]_  = ~A203 & A201;
  assign \new_[98101]_  = ~A266 & A265;
  assign \new_[98102]_  = \new_[98101]_  & \new_[98098]_ ;
  assign \new_[98103]_  = \new_[98102]_  & \new_[98095]_ ;
  assign \new_[98106]_  = ~A268 & ~A267;
  assign \new_[98109]_  = A298 & A269;
  assign \new_[98110]_  = \new_[98109]_  & \new_[98106]_ ;
  assign \new_[98113]_  = ~A300 & ~A299;
  assign \new_[98116]_  = A302 & ~A301;
  assign \new_[98117]_  = \new_[98116]_  & \new_[98113]_ ;
  assign \new_[98118]_  = \new_[98117]_  & \new_[98110]_ ;
  assign \new_[98121]_  = ~A168 & A169;
  assign \new_[98124]_  = ~A200 & A199;
  assign \new_[98125]_  = \new_[98124]_  & \new_[98121]_ ;
  assign \new_[98128]_  = ~A203 & A201;
  assign \new_[98131]_  = ~A266 & A265;
  assign \new_[98132]_  = \new_[98131]_  & \new_[98128]_ ;
  assign \new_[98133]_  = \new_[98132]_  & \new_[98125]_ ;
  assign \new_[98136]_  = ~A268 & ~A267;
  assign \new_[98139]_  = ~A298 & A269;
  assign \new_[98140]_  = \new_[98139]_  & \new_[98136]_ ;
  assign \new_[98143]_  = ~A300 & A299;
  assign \new_[98146]_  = A302 & ~A301;
  assign \new_[98147]_  = \new_[98146]_  & \new_[98143]_ ;
  assign \new_[98148]_  = \new_[98147]_  & \new_[98140]_ ;
  assign \new_[98151]_  = ~A168 & A169;
  assign \new_[98154]_  = ~A200 & A199;
  assign \new_[98155]_  = \new_[98154]_  & \new_[98151]_ ;
  assign \new_[98158]_  = ~A202 & ~A201;
  assign \new_[98161]_  = ~A265 & A203;
  assign \new_[98162]_  = \new_[98161]_  & \new_[98158]_ ;
  assign \new_[98163]_  = \new_[98162]_  & \new_[98155]_ ;
  assign \new_[98166]_  = A267 & A266;
  assign \new_[98169]_  = A298 & A268;
  assign \new_[98170]_  = \new_[98169]_  & \new_[98166]_ ;
  assign \new_[98173]_  = ~A300 & ~A299;
  assign \new_[98176]_  = A302 & ~A301;
  assign \new_[98177]_  = \new_[98176]_  & \new_[98173]_ ;
  assign \new_[98178]_  = \new_[98177]_  & \new_[98170]_ ;
  assign \new_[98181]_  = ~A168 & A169;
  assign \new_[98184]_  = ~A200 & A199;
  assign \new_[98185]_  = \new_[98184]_  & \new_[98181]_ ;
  assign \new_[98188]_  = ~A202 & ~A201;
  assign \new_[98191]_  = ~A265 & A203;
  assign \new_[98192]_  = \new_[98191]_  & \new_[98188]_ ;
  assign \new_[98193]_  = \new_[98192]_  & \new_[98185]_ ;
  assign \new_[98196]_  = A267 & A266;
  assign \new_[98199]_  = ~A298 & A268;
  assign \new_[98200]_  = \new_[98199]_  & \new_[98196]_ ;
  assign \new_[98203]_  = ~A300 & A299;
  assign \new_[98206]_  = A302 & ~A301;
  assign \new_[98207]_  = \new_[98206]_  & \new_[98203]_ ;
  assign \new_[98208]_  = \new_[98207]_  & \new_[98200]_ ;
  assign \new_[98211]_  = ~A168 & A169;
  assign \new_[98214]_  = ~A200 & A199;
  assign \new_[98215]_  = \new_[98214]_  & \new_[98211]_ ;
  assign \new_[98218]_  = ~A202 & ~A201;
  assign \new_[98221]_  = ~A265 & A203;
  assign \new_[98222]_  = \new_[98221]_  & \new_[98218]_ ;
  assign \new_[98223]_  = \new_[98222]_  & \new_[98215]_ ;
  assign \new_[98226]_  = A267 & A266;
  assign \new_[98229]_  = A298 & ~A269;
  assign \new_[98230]_  = \new_[98229]_  & \new_[98226]_ ;
  assign \new_[98233]_  = ~A300 & ~A299;
  assign \new_[98236]_  = A302 & ~A301;
  assign \new_[98237]_  = \new_[98236]_  & \new_[98233]_ ;
  assign \new_[98238]_  = \new_[98237]_  & \new_[98230]_ ;
  assign \new_[98241]_  = ~A168 & A169;
  assign \new_[98244]_  = ~A200 & A199;
  assign \new_[98245]_  = \new_[98244]_  & \new_[98241]_ ;
  assign \new_[98248]_  = ~A202 & ~A201;
  assign \new_[98251]_  = ~A265 & A203;
  assign \new_[98252]_  = \new_[98251]_  & \new_[98248]_ ;
  assign \new_[98253]_  = \new_[98252]_  & \new_[98245]_ ;
  assign \new_[98256]_  = A267 & A266;
  assign \new_[98259]_  = ~A298 & ~A269;
  assign \new_[98260]_  = \new_[98259]_  & \new_[98256]_ ;
  assign \new_[98263]_  = ~A300 & A299;
  assign \new_[98266]_  = A302 & ~A301;
  assign \new_[98267]_  = \new_[98266]_  & \new_[98263]_ ;
  assign \new_[98268]_  = \new_[98267]_  & \new_[98260]_ ;
  assign \new_[98271]_  = ~A168 & A169;
  assign \new_[98274]_  = ~A200 & A199;
  assign \new_[98275]_  = \new_[98274]_  & \new_[98271]_ ;
  assign \new_[98278]_  = ~A202 & ~A201;
  assign \new_[98281]_  = ~A265 & A203;
  assign \new_[98282]_  = \new_[98281]_  & \new_[98278]_ ;
  assign \new_[98283]_  = \new_[98282]_  & \new_[98275]_ ;
  assign \new_[98286]_  = ~A267 & A266;
  assign \new_[98289]_  = A269 & ~A268;
  assign \new_[98290]_  = \new_[98289]_  & \new_[98286]_ ;
  assign \new_[98293]_  = ~A299 & A298;
  assign \new_[98296]_  = A301 & A300;
  assign \new_[98297]_  = \new_[98296]_  & \new_[98293]_ ;
  assign \new_[98298]_  = \new_[98297]_  & \new_[98290]_ ;
  assign \new_[98301]_  = ~A168 & A169;
  assign \new_[98304]_  = ~A200 & A199;
  assign \new_[98305]_  = \new_[98304]_  & \new_[98301]_ ;
  assign \new_[98308]_  = ~A202 & ~A201;
  assign \new_[98311]_  = ~A265 & A203;
  assign \new_[98312]_  = \new_[98311]_  & \new_[98308]_ ;
  assign \new_[98313]_  = \new_[98312]_  & \new_[98305]_ ;
  assign \new_[98316]_  = ~A267 & A266;
  assign \new_[98319]_  = A269 & ~A268;
  assign \new_[98320]_  = \new_[98319]_  & \new_[98316]_ ;
  assign \new_[98323]_  = ~A299 & A298;
  assign \new_[98326]_  = ~A302 & A300;
  assign \new_[98327]_  = \new_[98326]_  & \new_[98323]_ ;
  assign \new_[98328]_  = \new_[98327]_  & \new_[98320]_ ;
  assign \new_[98331]_  = ~A168 & A169;
  assign \new_[98334]_  = ~A200 & A199;
  assign \new_[98335]_  = \new_[98334]_  & \new_[98331]_ ;
  assign \new_[98338]_  = ~A202 & ~A201;
  assign \new_[98341]_  = ~A265 & A203;
  assign \new_[98342]_  = \new_[98341]_  & \new_[98338]_ ;
  assign \new_[98343]_  = \new_[98342]_  & \new_[98335]_ ;
  assign \new_[98346]_  = ~A267 & A266;
  assign \new_[98349]_  = A269 & ~A268;
  assign \new_[98350]_  = \new_[98349]_  & \new_[98346]_ ;
  assign \new_[98353]_  = A299 & ~A298;
  assign \new_[98356]_  = A301 & A300;
  assign \new_[98357]_  = \new_[98356]_  & \new_[98353]_ ;
  assign \new_[98358]_  = \new_[98357]_  & \new_[98350]_ ;
  assign \new_[98361]_  = ~A168 & A169;
  assign \new_[98364]_  = ~A200 & A199;
  assign \new_[98365]_  = \new_[98364]_  & \new_[98361]_ ;
  assign \new_[98368]_  = ~A202 & ~A201;
  assign \new_[98371]_  = ~A265 & A203;
  assign \new_[98372]_  = \new_[98371]_  & \new_[98368]_ ;
  assign \new_[98373]_  = \new_[98372]_  & \new_[98365]_ ;
  assign \new_[98376]_  = ~A267 & A266;
  assign \new_[98379]_  = A269 & ~A268;
  assign \new_[98380]_  = \new_[98379]_  & \new_[98376]_ ;
  assign \new_[98383]_  = A299 & ~A298;
  assign \new_[98386]_  = ~A302 & A300;
  assign \new_[98387]_  = \new_[98386]_  & \new_[98383]_ ;
  assign \new_[98388]_  = \new_[98387]_  & \new_[98380]_ ;
  assign \new_[98391]_  = ~A168 & A169;
  assign \new_[98394]_  = ~A200 & A199;
  assign \new_[98395]_  = \new_[98394]_  & \new_[98391]_ ;
  assign \new_[98398]_  = ~A202 & ~A201;
  assign \new_[98401]_  = A265 & A203;
  assign \new_[98402]_  = \new_[98401]_  & \new_[98398]_ ;
  assign \new_[98403]_  = \new_[98402]_  & \new_[98395]_ ;
  assign \new_[98406]_  = A267 & ~A266;
  assign \new_[98409]_  = A298 & A268;
  assign \new_[98410]_  = \new_[98409]_  & \new_[98406]_ ;
  assign \new_[98413]_  = ~A300 & ~A299;
  assign \new_[98416]_  = A302 & ~A301;
  assign \new_[98417]_  = \new_[98416]_  & \new_[98413]_ ;
  assign \new_[98418]_  = \new_[98417]_  & \new_[98410]_ ;
  assign \new_[98421]_  = ~A168 & A169;
  assign \new_[98424]_  = ~A200 & A199;
  assign \new_[98425]_  = \new_[98424]_  & \new_[98421]_ ;
  assign \new_[98428]_  = ~A202 & ~A201;
  assign \new_[98431]_  = A265 & A203;
  assign \new_[98432]_  = \new_[98431]_  & \new_[98428]_ ;
  assign \new_[98433]_  = \new_[98432]_  & \new_[98425]_ ;
  assign \new_[98436]_  = A267 & ~A266;
  assign \new_[98439]_  = ~A298 & A268;
  assign \new_[98440]_  = \new_[98439]_  & \new_[98436]_ ;
  assign \new_[98443]_  = ~A300 & A299;
  assign \new_[98446]_  = A302 & ~A301;
  assign \new_[98447]_  = \new_[98446]_  & \new_[98443]_ ;
  assign \new_[98448]_  = \new_[98447]_  & \new_[98440]_ ;
  assign \new_[98451]_  = ~A168 & A169;
  assign \new_[98454]_  = ~A200 & A199;
  assign \new_[98455]_  = \new_[98454]_  & \new_[98451]_ ;
  assign \new_[98458]_  = ~A202 & ~A201;
  assign \new_[98461]_  = A265 & A203;
  assign \new_[98462]_  = \new_[98461]_  & \new_[98458]_ ;
  assign \new_[98463]_  = \new_[98462]_  & \new_[98455]_ ;
  assign \new_[98466]_  = A267 & ~A266;
  assign \new_[98469]_  = A298 & ~A269;
  assign \new_[98470]_  = \new_[98469]_  & \new_[98466]_ ;
  assign \new_[98473]_  = ~A300 & ~A299;
  assign \new_[98476]_  = A302 & ~A301;
  assign \new_[98477]_  = \new_[98476]_  & \new_[98473]_ ;
  assign \new_[98478]_  = \new_[98477]_  & \new_[98470]_ ;
  assign \new_[98481]_  = ~A168 & A169;
  assign \new_[98484]_  = ~A200 & A199;
  assign \new_[98485]_  = \new_[98484]_  & \new_[98481]_ ;
  assign \new_[98488]_  = ~A202 & ~A201;
  assign \new_[98491]_  = A265 & A203;
  assign \new_[98492]_  = \new_[98491]_  & \new_[98488]_ ;
  assign \new_[98493]_  = \new_[98492]_  & \new_[98485]_ ;
  assign \new_[98496]_  = A267 & ~A266;
  assign \new_[98499]_  = ~A298 & ~A269;
  assign \new_[98500]_  = \new_[98499]_  & \new_[98496]_ ;
  assign \new_[98503]_  = ~A300 & A299;
  assign \new_[98506]_  = A302 & ~A301;
  assign \new_[98507]_  = \new_[98506]_  & \new_[98503]_ ;
  assign \new_[98508]_  = \new_[98507]_  & \new_[98500]_ ;
  assign \new_[98511]_  = ~A168 & A169;
  assign \new_[98514]_  = ~A200 & A199;
  assign \new_[98515]_  = \new_[98514]_  & \new_[98511]_ ;
  assign \new_[98518]_  = ~A202 & ~A201;
  assign \new_[98521]_  = A265 & A203;
  assign \new_[98522]_  = \new_[98521]_  & \new_[98518]_ ;
  assign \new_[98523]_  = \new_[98522]_  & \new_[98515]_ ;
  assign \new_[98526]_  = ~A267 & ~A266;
  assign \new_[98529]_  = A269 & ~A268;
  assign \new_[98530]_  = \new_[98529]_  & \new_[98526]_ ;
  assign \new_[98533]_  = ~A299 & A298;
  assign \new_[98536]_  = A301 & A300;
  assign \new_[98537]_  = \new_[98536]_  & \new_[98533]_ ;
  assign \new_[98538]_  = \new_[98537]_  & \new_[98530]_ ;
  assign \new_[98541]_  = ~A168 & A169;
  assign \new_[98544]_  = ~A200 & A199;
  assign \new_[98545]_  = \new_[98544]_  & \new_[98541]_ ;
  assign \new_[98548]_  = ~A202 & ~A201;
  assign \new_[98551]_  = A265 & A203;
  assign \new_[98552]_  = \new_[98551]_  & \new_[98548]_ ;
  assign \new_[98553]_  = \new_[98552]_  & \new_[98545]_ ;
  assign \new_[98556]_  = ~A267 & ~A266;
  assign \new_[98559]_  = A269 & ~A268;
  assign \new_[98560]_  = \new_[98559]_  & \new_[98556]_ ;
  assign \new_[98563]_  = ~A299 & A298;
  assign \new_[98566]_  = ~A302 & A300;
  assign \new_[98567]_  = \new_[98566]_  & \new_[98563]_ ;
  assign \new_[98568]_  = \new_[98567]_  & \new_[98560]_ ;
  assign \new_[98571]_  = ~A168 & A169;
  assign \new_[98574]_  = ~A200 & A199;
  assign \new_[98575]_  = \new_[98574]_  & \new_[98571]_ ;
  assign \new_[98578]_  = ~A202 & ~A201;
  assign \new_[98581]_  = A265 & A203;
  assign \new_[98582]_  = \new_[98581]_  & \new_[98578]_ ;
  assign \new_[98583]_  = \new_[98582]_  & \new_[98575]_ ;
  assign \new_[98586]_  = ~A267 & ~A266;
  assign \new_[98589]_  = A269 & ~A268;
  assign \new_[98590]_  = \new_[98589]_  & \new_[98586]_ ;
  assign \new_[98593]_  = A299 & ~A298;
  assign \new_[98596]_  = A301 & A300;
  assign \new_[98597]_  = \new_[98596]_  & \new_[98593]_ ;
  assign \new_[98598]_  = \new_[98597]_  & \new_[98590]_ ;
  assign \new_[98601]_  = ~A168 & A169;
  assign \new_[98604]_  = ~A200 & A199;
  assign \new_[98605]_  = \new_[98604]_  & \new_[98601]_ ;
  assign \new_[98608]_  = ~A202 & ~A201;
  assign \new_[98611]_  = A265 & A203;
  assign \new_[98612]_  = \new_[98611]_  & \new_[98608]_ ;
  assign \new_[98613]_  = \new_[98612]_  & \new_[98605]_ ;
  assign \new_[98616]_  = ~A267 & ~A266;
  assign \new_[98619]_  = A269 & ~A268;
  assign \new_[98620]_  = \new_[98619]_  & \new_[98616]_ ;
  assign \new_[98623]_  = A299 & ~A298;
  assign \new_[98626]_  = ~A302 & A300;
  assign \new_[98627]_  = \new_[98626]_  & \new_[98623]_ ;
  assign \new_[98628]_  = \new_[98627]_  & \new_[98620]_ ;
  assign \new_[98631]_  = ~A169 & ~A170;
  assign \new_[98634]_  = ~A199 & A168;
  assign \new_[98635]_  = \new_[98634]_  & \new_[98631]_ ;
  assign \new_[98638]_  = A201 & A200;
  assign \new_[98641]_  = ~A265 & A202;
  assign \new_[98642]_  = \new_[98641]_  & \new_[98638]_ ;
  assign \new_[98643]_  = \new_[98642]_  & \new_[98635]_ ;
  assign \new_[98646]_  = A267 & A266;
  assign \new_[98649]_  = A298 & A268;
  assign \new_[98650]_  = \new_[98649]_  & \new_[98646]_ ;
  assign \new_[98653]_  = ~A300 & ~A299;
  assign \new_[98656]_  = A302 & ~A301;
  assign \new_[98657]_  = \new_[98656]_  & \new_[98653]_ ;
  assign \new_[98658]_  = \new_[98657]_  & \new_[98650]_ ;
  assign \new_[98661]_  = ~A169 & ~A170;
  assign \new_[98664]_  = ~A199 & A168;
  assign \new_[98665]_  = \new_[98664]_  & \new_[98661]_ ;
  assign \new_[98668]_  = A201 & A200;
  assign \new_[98671]_  = ~A265 & A202;
  assign \new_[98672]_  = \new_[98671]_  & \new_[98668]_ ;
  assign \new_[98673]_  = \new_[98672]_  & \new_[98665]_ ;
  assign \new_[98676]_  = A267 & A266;
  assign \new_[98679]_  = ~A298 & A268;
  assign \new_[98680]_  = \new_[98679]_  & \new_[98676]_ ;
  assign \new_[98683]_  = ~A300 & A299;
  assign \new_[98686]_  = A302 & ~A301;
  assign \new_[98687]_  = \new_[98686]_  & \new_[98683]_ ;
  assign \new_[98688]_  = \new_[98687]_  & \new_[98680]_ ;
  assign \new_[98691]_  = ~A169 & ~A170;
  assign \new_[98694]_  = ~A199 & A168;
  assign \new_[98695]_  = \new_[98694]_  & \new_[98691]_ ;
  assign \new_[98698]_  = A201 & A200;
  assign \new_[98701]_  = ~A265 & A202;
  assign \new_[98702]_  = \new_[98701]_  & \new_[98698]_ ;
  assign \new_[98703]_  = \new_[98702]_  & \new_[98695]_ ;
  assign \new_[98706]_  = A267 & A266;
  assign \new_[98709]_  = A298 & ~A269;
  assign \new_[98710]_  = \new_[98709]_  & \new_[98706]_ ;
  assign \new_[98713]_  = ~A300 & ~A299;
  assign \new_[98716]_  = A302 & ~A301;
  assign \new_[98717]_  = \new_[98716]_  & \new_[98713]_ ;
  assign \new_[98718]_  = \new_[98717]_  & \new_[98710]_ ;
  assign \new_[98721]_  = ~A169 & ~A170;
  assign \new_[98724]_  = ~A199 & A168;
  assign \new_[98725]_  = \new_[98724]_  & \new_[98721]_ ;
  assign \new_[98728]_  = A201 & A200;
  assign \new_[98731]_  = ~A265 & A202;
  assign \new_[98732]_  = \new_[98731]_  & \new_[98728]_ ;
  assign \new_[98733]_  = \new_[98732]_  & \new_[98725]_ ;
  assign \new_[98736]_  = A267 & A266;
  assign \new_[98739]_  = ~A298 & ~A269;
  assign \new_[98740]_  = \new_[98739]_  & \new_[98736]_ ;
  assign \new_[98743]_  = ~A300 & A299;
  assign \new_[98746]_  = A302 & ~A301;
  assign \new_[98747]_  = \new_[98746]_  & \new_[98743]_ ;
  assign \new_[98748]_  = \new_[98747]_  & \new_[98740]_ ;
  assign \new_[98751]_  = ~A169 & ~A170;
  assign \new_[98754]_  = ~A199 & A168;
  assign \new_[98755]_  = \new_[98754]_  & \new_[98751]_ ;
  assign \new_[98758]_  = A201 & A200;
  assign \new_[98761]_  = ~A265 & A202;
  assign \new_[98762]_  = \new_[98761]_  & \new_[98758]_ ;
  assign \new_[98763]_  = \new_[98762]_  & \new_[98755]_ ;
  assign \new_[98766]_  = ~A267 & A266;
  assign \new_[98769]_  = A269 & ~A268;
  assign \new_[98770]_  = \new_[98769]_  & \new_[98766]_ ;
  assign \new_[98773]_  = ~A299 & A298;
  assign \new_[98776]_  = A301 & A300;
  assign \new_[98777]_  = \new_[98776]_  & \new_[98773]_ ;
  assign \new_[98778]_  = \new_[98777]_  & \new_[98770]_ ;
  assign \new_[98781]_  = ~A169 & ~A170;
  assign \new_[98784]_  = ~A199 & A168;
  assign \new_[98785]_  = \new_[98784]_  & \new_[98781]_ ;
  assign \new_[98788]_  = A201 & A200;
  assign \new_[98791]_  = ~A265 & A202;
  assign \new_[98792]_  = \new_[98791]_  & \new_[98788]_ ;
  assign \new_[98793]_  = \new_[98792]_  & \new_[98785]_ ;
  assign \new_[98796]_  = ~A267 & A266;
  assign \new_[98799]_  = A269 & ~A268;
  assign \new_[98800]_  = \new_[98799]_  & \new_[98796]_ ;
  assign \new_[98803]_  = ~A299 & A298;
  assign \new_[98806]_  = ~A302 & A300;
  assign \new_[98807]_  = \new_[98806]_  & \new_[98803]_ ;
  assign \new_[98808]_  = \new_[98807]_  & \new_[98800]_ ;
  assign \new_[98811]_  = ~A169 & ~A170;
  assign \new_[98814]_  = ~A199 & A168;
  assign \new_[98815]_  = \new_[98814]_  & \new_[98811]_ ;
  assign \new_[98818]_  = A201 & A200;
  assign \new_[98821]_  = ~A265 & A202;
  assign \new_[98822]_  = \new_[98821]_  & \new_[98818]_ ;
  assign \new_[98823]_  = \new_[98822]_  & \new_[98815]_ ;
  assign \new_[98826]_  = ~A267 & A266;
  assign \new_[98829]_  = A269 & ~A268;
  assign \new_[98830]_  = \new_[98829]_  & \new_[98826]_ ;
  assign \new_[98833]_  = A299 & ~A298;
  assign \new_[98836]_  = A301 & A300;
  assign \new_[98837]_  = \new_[98836]_  & \new_[98833]_ ;
  assign \new_[98838]_  = \new_[98837]_  & \new_[98830]_ ;
  assign \new_[98841]_  = ~A169 & ~A170;
  assign \new_[98844]_  = ~A199 & A168;
  assign \new_[98845]_  = \new_[98844]_  & \new_[98841]_ ;
  assign \new_[98848]_  = A201 & A200;
  assign \new_[98851]_  = ~A265 & A202;
  assign \new_[98852]_  = \new_[98851]_  & \new_[98848]_ ;
  assign \new_[98853]_  = \new_[98852]_  & \new_[98845]_ ;
  assign \new_[98856]_  = ~A267 & A266;
  assign \new_[98859]_  = A269 & ~A268;
  assign \new_[98860]_  = \new_[98859]_  & \new_[98856]_ ;
  assign \new_[98863]_  = A299 & ~A298;
  assign \new_[98866]_  = ~A302 & A300;
  assign \new_[98867]_  = \new_[98866]_  & \new_[98863]_ ;
  assign \new_[98868]_  = \new_[98867]_  & \new_[98860]_ ;
  assign \new_[98871]_  = ~A169 & ~A170;
  assign \new_[98874]_  = ~A199 & A168;
  assign \new_[98875]_  = \new_[98874]_  & \new_[98871]_ ;
  assign \new_[98878]_  = A201 & A200;
  assign \new_[98881]_  = A265 & A202;
  assign \new_[98882]_  = \new_[98881]_  & \new_[98878]_ ;
  assign \new_[98883]_  = \new_[98882]_  & \new_[98875]_ ;
  assign \new_[98886]_  = A267 & ~A266;
  assign \new_[98889]_  = A298 & A268;
  assign \new_[98890]_  = \new_[98889]_  & \new_[98886]_ ;
  assign \new_[98893]_  = ~A300 & ~A299;
  assign \new_[98896]_  = A302 & ~A301;
  assign \new_[98897]_  = \new_[98896]_  & \new_[98893]_ ;
  assign \new_[98898]_  = \new_[98897]_  & \new_[98890]_ ;
  assign \new_[98901]_  = ~A169 & ~A170;
  assign \new_[98904]_  = ~A199 & A168;
  assign \new_[98905]_  = \new_[98904]_  & \new_[98901]_ ;
  assign \new_[98908]_  = A201 & A200;
  assign \new_[98911]_  = A265 & A202;
  assign \new_[98912]_  = \new_[98911]_  & \new_[98908]_ ;
  assign \new_[98913]_  = \new_[98912]_  & \new_[98905]_ ;
  assign \new_[98916]_  = A267 & ~A266;
  assign \new_[98919]_  = ~A298 & A268;
  assign \new_[98920]_  = \new_[98919]_  & \new_[98916]_ ;
  assign \new_[98923]_  = ~A300 & A299;
  assign \new_[98926]_  = A302 & ~A301;
  assign \new_[98927]_  = \new_[98926]_  & \new_[98923]_ ;
  assign \new_[98928]_  = \new_[98927]_  & \new_[98920]_ ;
  assign \new_[98931]_  = ~A169 & ~A170;
  assign \new_[98934]_  = ~A199 & A168;
  assign \new_[98935]_  = \new_[98934]_  & \new_[98931]_ ;
  assign \new_[98938]_  = A201 & A200;
  assign \new_[98941]_  = A265 & A202;
  assign \new_[98942]_  = \new_[98941]_  & \new_[98938]_ ;
  assign \new_[98943]_  = \new_[98942]_  & \new_[98935]_ ;
  assign \new_[98946]_  = A267 & ~A266;
  assign \new_[98949]_  = A298 & ~A269;
  assign \new_[98950]_  = \new_[98949]_  & \new_[98946]_ ;
  assign \new_[98953]_  = ~A300 & ~A299;
  assign \new_[98956]_  = A302 & ~A301;
  assign \new_[98957]_  = \new_[98956]_  & \new_[98953]_ ;
  assign \new_[98958]_  = \new_[98957]_  & \new_[98950]_ ;
  assign \new_[98961]_  = ~A169 & ~A170;
  assign \new_[98964]_  = ~A199 & A168;
  assign \new_[98965]_  = \new_[98964]_  & \new_[98961]_ ;
  assign \new_[98968]_  = A201 & A200;
  assign \new_[98971]_  = A265 & A202;
  assign \new_[98972]_  = \new_[98971]_  & \new_[98968]_ ;
  assign \new_[98973]_  = \new_[98972]_  & \new_[98965]_ ;
  assign \new_[98976]_  = A267 & ~A266;
  assign \new_[98979]_  = ~A298 & ~A269;
  assign \new_[98980]_  = \new_[98979]_  & \new_[98976]_ ;
  assign \new_[98983]_  = ~A300 & A299;
  assign \new_[98986]_  = A302 & ~A301;
  assign \new_[98987]_  = \new_[98986]_  & \new_[98983]_ ;
  assign \new_[98988]_  = \new_[98987]_  & \new_[98980]_ ;
  assign \new_[98991]_  = ~A169 & ~A170;
  assign \new_[98994]_  = ~A199 & A168;
  assign \new_[98995]_  = \new_[98994]_  & \new_[98991]_ ;
  assign \new_[98998]_  = A201 & A200;
  assign \new_[99001]_  = A265 & A202;
  assign \new_[99002]_  = \new_[99001]_  & \new_[98998]_ ;
  assign \new_[99003]_  = \new_[99002]_  & \new_[98995]_ ;
  assign \new_[99006]_  = ~A267 & ~A266;
  assign \new_[99009]_  = A269 & ~A268;
  assign \new_[99010]_  = \new_[99009]_  & \new_[99006]_ ;
  assign \new_[99013]_  = ~A299 & A298;
  assign \new_[99016]_  = A301 & A300;
  assign \new_[99017]_  = \new_[99016]_  & \new_[99013]_ ;
  assign \new_[99018]_  = \new_[99017]_  & \new_[99010]_ ;
  assign \new_[99021]_  = ~A169 & ~A170;
  assign \new_[99024]_  = ~A199 & A168;
  assign \new_[99025]_  = \new_[99024]_  & \new_[99021]_ ;
  assign \new_[99028]_  = A201 & A200;
  assign \new_[99031]_  = A265 & A202;
  assign \new_[99032]_  = \new_[99031]_  & \new_[99028]_ ;
  assign \new_[99033]_  = \new_[99032]_  & \new_[99025]_ ;
  assign \new_[99036]_  = ~A267 & ~A266;
  assign \new_[99039]_  = A269 & ~A268;
  assign \new_[99040]_  = \new_[99039]_  & \new_[99036]_ ;
  assign \new_[99043]_  = ~A299 & A298;
  assign \new_[99046]_  = ~A302 & A300;
  assign \new_[99047]_  = \new_[99046]_  & \new_[99043]_ ;
  assign \new_[99048]_  = \new_[99047]_  & \new_[99040]_ ;
  assign \new_[99051]_  = ~A169 & ~A170;
  assign \new_[99054]_  = ~A199 & A168;
  assign \new_[99055]_  = \new_[99054]_  & \new_[99051]_ ;
  assign \new_[99058]_  = A201 & A200;
  assign \new_[99061]_  = A265 & A202;
  assign \new_[99062]_  = \new_[99061]_  & \new_[99058]_ ;
  assign \new_[99063]_  = \new_[99062]_  & \new_[99055]_ ;
  assign \new_[99066]_  = ~A267 & ~A266;
  assign \new_[99069]_  = A269 & ~A268;
  assign \new_[99070]_  = \new_[99069]_  & \new_[99066]_ ;
  assign \new_[99073]_  = A299 & ~A298;
  assign \new_[99076]_  = A301 & A300;
  assign \new_[99077]_  = \new_[99076]_  & \new_[99073]_ ;
  assign \new_[99078]_  = \new_[99077]_  & \new_[99070]_ ;
  assign \new_[99081]_  = ~A169 & ~A170;
  assign \new_[99084]_  = ~A199 & A168;
  assign \new_[99085]_  = \new_[99084]_  & \new_[99081]_ ;
  assign \new_[99088]_  = A201 & A200;
  assign \new_[99091]_  = A265 & A202;
  assign \new_[99092]_  = \new_[99091]_  & \new_[99088]_ ;
  assign \new_[99093]_  = \new_[99092]_  & \new_[99085]_ ;
  assign \new_[99096]_  = ~A267 & ~A266;
  assign \new_[99099]_  = A269 & ~A268;
  assign \new_[99100]_  = \new_[99099]_  & \new_[99096]_ ;
  assign \new_[99103]_  = A299 & ~A298;
  assign \new_[99106]_  = ~A302 & A300;
  assign \new_[99107]_  = \new_[99106]_  & \new_[99103]_ ;
  assign \new_[99108]_  = \new_[99107]_  & \new_[99100]_ ;
  assign \new_[99111]_  = ~A169 & ~A170;
  assign \new_[99114]_  = ~A199 & A168;
  assign \new_[99115]_  = \new_[99114]_  & \new_[99111]_ ;
  assign \new_[99118]_  = A201 & A200;
  assign \new_[99121]_  = ~A265 & ~A203;
  assign \new_[99122]_  = \new_[99121]_  & \new_[99118]_ ;
  assign \new_[99123]_  = \new_[99122]_  & \new_[99115]_ ;
  assign \new_[99126]_  = A267 & A266;
  assign \new_[99129]_  = A298 & A268;
  assign \new_[99130]_  = \new_[99129]_  & \new_[99126]_ ;
  assign \new_[99133]_  = ~A300 & ~A299;
  assign \new_[99136]_  = A302 & ~A301;
  assign \new_[99137]_  = \new_[99136]_  & \new_[99133]_ ;
  assign \new_[99138]_  = \new_[99137]_  & \new_[99130]_ ;
  assign \new_[99141]_  = ~A169 & ~A170;
  assign \new_[99144]_  = ~A199 & A168;
  assign \new_[99145]_  = \new_[99144]_  & \new_[99141]_ ;
  assign \new_[99148]_  = A201 & A200;
  assign \new_[99151]_  = ~A265 & ~A203;
  assign \new_[99152]_  = \new_[99151]_  & \new_[99148]_ ;
  assign \new_[99153]_  = \new_[99152]_  & \new_[99145]_ ;
  assign \new_[99156]_  = A267 & A266;
  assign \new_[99159]_  = ~A298 & A268;
  assign \new_[99160]_  = \new_[99159]_  & \new_[99156]_ ;
  assign \new_[99163]_  = ~A300 & A299;
  assign \new_[99166]_  = A302 & ~A301;
  assign \new_[99167]_  = \new_[99166]_  & \new_[99163]_ ;
  assign \new_[99168]_  = \new_[99167]_  & \new_[99160]_ ;
  assign \new_[99171]_  = ~A169 & ~A170;
  assign \new_[99174]_  = ~A199 & A168;
  assign \new_[99175]_  = \new_[99174]_  & \new_[99171]_ ;
  assign \new_[99178]_  = A201 & A200;
  assign \new_[99181]_  = ~A265 & ~A203;
  assign \new_[99182]_  = \new_[99181]_  & \new_[99178]_ ;
  assign \new_[99183]_  = \new_[99182]_  & \new_[99175]_ ;
  assign \new_[99186]_  = A267 & A266;
  assign \new_[99189]_  = A298 & ~A269;
  assign \new_[99190]_  = \new_[99189]_  & \new_[99186]_ ;
  assign \new_[99193]_  = ~A300 & ~A299;
  assign \new_[99196]_  = A302 & ~A301;
  assign \new_[99197]_  = \new_[99196]_  & \new_[99193]_ ;
  assign \new_[99198]_  = \new_[99197]_  & \new_[99190]_ ;
  assign \new_[99201]_  = ~A169 & ~A170;
  assign \new_[99204]_  = ~A199 & A168;
  assign \new_[99205]_  = \new_[99204]_  & \new_[99201]_ ;
  assign \new_[99208]_  = A201 & A200;
  assign \new_[99211]_  = ~A265 & ~A203;
  assign \new_[99212]_  = \new_[99211]_  & \new_[99208]_ ;
  assign \new_[99213]_  = \new_[99212]_  & \new_[99205]_ ;
  assign \new_[99216]_  = A267 & A266;
  assign \new_[99219]_  = ~A298 & ~A269;
  assign \new_[99220]_  = \new_[99219]_  & \new_[99216]_ ;
  assign \new_[99223]_  = ~A300 & A299;
  assign \new_[99226]_  = A302 & ~A301;
  assign \new_[99227]_  = \new_[99226]_  & \new_[99223]_ ;
  assign \new_[99228]_  = \new_[99227]_  & \new_[99220]_ ;
  assign \new_[99231]_  = ~A169 & ~A170;
  assign \new_[99234]_  = ~A199 & A168;
  assign \new_[99235]_  = \new_[99234]_  & \new_[99231]_ ;
  assign \new_[99238]_  = A201 & A200;
  assign \new_[99241]_  = ~A265 & ~A203;
  assign \new_[99242]_  = \new_[99241]_  & \new_[99238]_ ;
  assign \new_[99243]_  = \new_[99242]_  & \new_[99235]_ ;
  assign \new_[99246]_  = ~A267 & A266;
  assign \new_[99249]_  = A269 & ~A268;
  assign \new_[99250]_  = \new_[99249]_  & \new_[99246]_ ;
  assign \new_[99253]_  = ~A299 & A298;
  assign \new_[99256]_  = A301 & A300;
  assign \new_[99257]_  = \new_[99256]_  & \new_[99253]_ ;
  assign \new_[99258]_  = \new_[99257]_  & \new_[99250]_ ;
  assign \new_[99261]_  = ~A169 & ~A170;
  assign \new_[99264]_  = ~A199 & A168;
  assign \new_[99265]_  = \new_[99264]_  & \new_[99261]_ ;
  assign \new_[99268]_  = A201 & A200;
  assign \new_[99271]_  = ~A265 & ~A203;
  assign \new_[99272]_  = \new_[99271]_  & \new_[99268]_ ;
  assign \new_[99273]_  = \new_[99272]_  & \new_[99265]_ ;
  assign \new_[99276]_  = ~A267 & A266;
  assign \new_[99279]_  = A269 & ~A268;
  assign \new_[99280]_  = \new_[99279]_  & \new_[99276]_ ;
  assign \new_[99283]_  = ~A299 & A298;
  assign \new_[99286]_  = ~A302 & A300;
  assign \new_[99287]_  = \new_[99286]_  & \new_[99283]_ ;
  assign \new_[99288]_  = \new_[99287]_  & \new_[99280]_ ;
  assign \new_[99291]_  = ~A169 & ~A170;
  assign \new_[99294]_  = ~A199 & A168;
  assign \new_[99295]_  = \new_[99294]_  & \new_[99291]_ ;
  assign \new_[99298]_  = A201 & A200;
  assign \new_[99301]_  = ~A265 & ~A203;
  assign \new_[99302]_  = \new_[99301]_  & \new_[99298]_ ;
  assign \new_[99303]_  = \new_[99302]_  & \new_[99295]_ ;
  assign \new_[99306]_  = ~A267 & A266;
  assign \new_[99309]_  = A269 & ~A268;
  assign \new_[99310]_  = \new_[99309]_  & \new_[99306]_ ;
  assign \new_[99313]_  = A299 & ~A298;
  assign \new_[99316]_  = A301 & A300;
  assign \new_[99317]_  = \new_[99316]_  & \new_[99313]_ ;
  assign \new_[99318]_  = \new_[99317]_  & \new_[99310]_ ;
  assign \new_[99321]_  = ~A169 & ~A170;
  assign \new_[99324]_  = ~A199 & A168;
  assign \new_[99325]_  = \new_[99324]_  & \new_[99321]_ ;
  assign \new_[99328]_  = A201 & A200;
  assign \new_[99331]_  = ~A265 & ~A203;
  assign \new_[99332]_  = \new_[99331]_  & \new_[99328]_ ;
  assign \new_[99333]_  = \new_[99332]_  & \new_[99325]_ ;
  assign \new_[99336]_  = ~A267 & A266;
  assign \new_[99339]_  = A269 & ~A268;
  assign \new_[99340]_  = \new_[99339]_  & \new_[99336]_ ;
  assign \new_[99343]_  = A299 & ~A298;
  assign \new_[99346]_  = ~A302 & A300;
  assign \new_[99347]_  = \new_[99346]_  & \new_[99343]_ ;
  assign \new_[99348]_  = \new_[99347]_  & \new_[99340]_ ;
  assign \new_[99351]_  = ~A169 & ~A170;
  assign \new_[99354]_  = ~A199 & A168;
  assign \new_[99355]_  = \new_[99354]_  & \new_[99351]_ ;
  assign \new_[99358]_  = A201 & A200;
  assign \new_[99361]_  = A265 & ~A203;
  assign \new_[99362]_  = \new_[99361]_  & \new_[99358]_ ;
  assign \new_[99363]_  = \new_[99362]_  & \new_[99355]_ ;
  assign \new_[99366]_  = A267 & ~A266;
  assign \new_[99369]_  = A298 & A268;
  assign \new_[99370]_  = \new_[99369]_  & \new_[99366]_ ;
  assign \new_[99373]_  = ~A300 & ~A299;
  assign \new_[99376]_  = A302 & ~A301;
  assign \new_[99377]_  = \new_[99376]_  & \new_[99373]_ ;
  assign \new_[99378]_  = \new_[99377]_  & \new_[99370]_ ;
  assign \new_[99381]_  = ~A169 & ~A170;
  assign \new_[99384]_  = ~A199 & A168;
  assign \new_[99385]_  = \new_[99384]_  & \new_[99381]_ ;
  assign \new_[99388]_  = A201 & A200;
  assign \new_[99391]_  = A265 & ~A203;
  assign \new_[99392]_  = \new_[99391]_  & \new_[99388]_ ;
  assign \new_[99393]_  = \new_[99392]_  & \new_[99385]_ ;
  assign \new_[99396]_  = A267 & ~A266;
  assign \new_[99399]_  = ~A298 & A268;
  assign \new_[99400]_  = \new_[99399]_  & \new_[99396]_ ;
  assign \new_[99403]_  = ~A300 & A299;
  assign \new_[99406]_  = A302 & ~A301;
  assign \new_[99407]_  = \new_[99406]_  & \new_[99403]_ ;
  assign \new_[99408]_  = \new_[99407]_  & \new_[99400]_ ;
  assign \new_[99411]_  = ~A169 & ~A170;
  assign \new_[99414]_  = ~A199 & A168;
  assign \new_[99415]_  = \new_[99414]_  & \new_[99411]_ ;
  assign \new_[99418]_  = A201 & A200;
  assign \new_[99421]_  = A265 & ~A203;
  assign \new_[99422]_  = \new_[99421]_  & \new_[99418]_ ;
  assign \new_[99423]_  = \new_[99422]_  & \new_[99415]_ ;
  assign \new_[99426]_  = A267 & ~A266;
  assign \new_[99429]_  = A298 & ~A269;
  assign \new_[99430]_  = \new_[99429]_  & \new_[99426]_ ;
  assign \new_[99433]_  = ~A300 & ~A299;
  assign \new_[99436]_  = A302 & ~A301;
  assign \new_[99437]_  = \new_[99436]_  & \new_[99433]_ ;
  assign \new_[99438]_  = \new_[99437]_  & \new_[99430]_ ;
  assign \new_[99441]_  = ~A169 & ~A170;
  assign \new_[99444]_  = ~A199 & A168;
  assign \new_[99445]_  = \new_[99444]_  & \new_[99441]_ ;
  assign \new_[99448]_  = A201 & A200;
  assign \new_[99451]_  = A265 & ~A203;
  assign \new_[99452]_  = \new_[99451]_  & \new_[99448]_ ;
  assign \new_[99453]_  = \new_[99452]_  & \new_[99445]_ ;
  assign \new_[99456]_  = A267 & ~A266;
  assign \new_[99459]_  = ~A298 & ~A269;
  assign \new_[99460]_  = \new_[99459]_  & \new_[99456]_ ;
  assign \new_[99463]_  = ~A300 & A299;
  assign \new_[99466]_  = A302 & ~A301;
  assign \new_[99467]_  = \new_[99466]_  & \new_[99463]_ ;
  assign \new_[99468]_  = \new_[99467]_  & \new_[99460]_ ;
  assign \new_[99471]_  = ~A169 & ~A170;
  assign \new_[99474]_  = ~A199 & A168;
  assign \new_[99475]_  = \new_[99474]_  & \new_[99471]_ ;
  assign \new_[99478]_  = A201 & A200;
  assign \new_[99481]_  = A265 & ~A203;
  assign \new_[99482]_  = \new_[99481]_  & \new_[99478]_ ;
  assign \new_[99483]_  = \new_[99482]_  & \new_[99475]_ ;
  assign \new_[99486]_  = ~A267 & ~A266;
  assign \new_[99489]_  = A269 & ~A268;
  assign \new_[99490]_  = \new_[99489]_  & \new_[99486]_ ;
  assign \new_[99493]_  = ~A299 & A298;
  assign \new_[99496]_  = A301 & A300;
  assign \new_[99497]_  = \new_[99496]_  & \new_[99493]_ ;
  assign \new_[99498]_  = \new_[99497]_  & \new_[99490]_ ;
  assign \new_[99501]_  = ~A169 & ~A170;
  assign \new_[99504]_  = ~A199 & A168;
  assign \new_[99505]_  = \new_[99504]_  & \new_[99501]_ ;
  assign \new_[99508]_  = A201 & A200;
  assign \new_[99511]_  = A265 & ~A203;
  assign \new_[99512]_  = \new_[99511]_  & \new_[99508]_ ;
  assign \new_[99513]_  = \new_[99512]_  & \new_[99505]_ ;
  assign \new_[99516]_  = ~A267 & ~A266;
  assign \new_[99519]_  = A269 & ~A268;
  assign \new_[99520]_  = \new_[99519]_  & \new_[99516]_ ;
  assign \new_[99523]_  = ~A299 & A298;
  assign \new_[99526]_  = ~A302 & A300;
  assign \new_[99527]_  = \new_[99526]_  & \new_[99523]_ ;
  assign \new_[99528]_  = \new_[99527]_  & \new_[99520]_ ;
  assign \new_[99531]_  = ~A169 & ~A170;
  assign \new_[99534]_  = ~A199 & A168;
  assign \new_[99535]_  = \new_[99534]_  & \new_[99531]_ ;
  assign \new_[99538]_  = A201 & A200;
  assign \new_[99541]_  = A265 & ~A203;
  assign \new_[99542]_  = \new_[99541]_  & \new_[99538]_ ;
  assign \new_[99543]_  = \new_[99542]_  & \new_[99535]_ ;
  assign \new_[99546]_  = ~A267 & ~A266;
  assign \new_[99549]_  = A269 & ~A268;
  assign \new_[99550]_  = \new_[99549]_  & \new_[99546]_ ;
  assign \new_[99553]_  = A299 & ~A298;
  assign \new_[99556]_  = A301 & A300;
  assign \new_[99557]_  = \new_[99556]_  & \new_[99553]_ ;
  assign \new_[99558]_  = \new_[99557]_  & \new_[99550]_ ;
  assign \new_[99561]_  = ~A169 & ~A170;
  assign \new_[99564]_  = ~A199 & A168;
  assign \new_[99565]_  = \new_[99564]_  & \new_[99561]_ ;
  assign \new_[99568]_  = A201 & A200;
  assign \new_[99571]_  = A265 & ~A203;
  assign \new_[99572]_  = \new_[99571]_  & \new_[99568]_ ;
  assign \new_[99573]_  = \new_[99572]_  & \new_[99565]_ ;
  assign \new_[99576]_  = ~A267 & ~A266;
  assign \new_[99579]_  = A269 & ~A268;
  assign \new_[99580]_  = \new_[99579]_  & \new_[99576]_ ;
  assign \new_[99583]_  = A299 & ~A298;
  assign \new_[99586]_  = ~A302 & A300;
  assign \new_[99587]_  = \new_[99586]_  & \new_[99583]_ ;
  assign \new_[99588]_  = \new_[99587]_  & \new_[99580]_ ;
  assign \new_[99591]_  = ~A169 & ~A170;
  assign \new_[99594]_  = ~A199 & A168;
  assign \new_[99595]_  = \new_[99594]_  & \new_[99591]_ ;
  assign \new_[99598]_  = ~A201 & A200;
  assign \new_[99601]_  = A203 & ~A202;
  assign \new_[99602]_  = \new_[99601]_  & \new_[99598]_ ;
  assign \new_[99603]_  = \new_[99602]_  & \new_[99595]_ ;
  assign \new_[99606]_  = A266 & ~A265;
  assign \new_[99609]_  = A268 & A267;
  assign \new_[99610]_  = \new_[99609]_  & \new_[99606]_ ;
  assign \new_[99613]_  = ~A299 & A298;
  assign \new_[99616]_  = A301 & A300;
  assign \new_[99617]_  = \new_[99616]_  & \new_[99613]_ ;
  assign \new_[99618]_  = \new_[99617]_  & \new_[99610]_ ;
  assign \new_[99621]_  = ~A169 & ~A170;
  assign \new_[99624]_  = ~A199 & A168;
  assign \new_[99625]_  = \new_[99624]_  & \new_[99621]_ ;
  assign \new_[99628]_  = ~A201 & A200;
  assign \new_[99631]_  = A203 & ~A202;
  assign \new_[99632]_  = \new_[99631]_  & \new_[99628]_ ;
  assign \new_[99633]_  = \new_[99632]_  & \new_[99625]_ ;
  assign \new_[99636]_  = A266 & ~A265;
  assign \new_[99639]_  = A268 & A267;
  assign \new_[99640]_  = \new_[99639]_  & \new_[99636]_ ;
  assign \new_[99643]_  = ~A299 & A298;
  assign \new_[99646]_  = ~A302 & A300;
  assign \new_[99647]_  = \new_[99646]_  & \new_[99643]_ ;
  assign \new_[99648]_  = \new_[99647]_  & \new_[99640]_ ;
  assign \new_[99651]_  = ~A169 & ~A170;
  assign \new_[99654]_  = ~A199 & A168;
  assign \new_[99655]_  = \new_[99654]_  & \new_[99651]_ ;
  assign \new_[99658]_  = ~A201 & A200;
  assign \new_[99661]_  = A203 & ~A202;
  assign \new_[99662]_  = \new_[99661]_  & \new_[99658]_ ;
  assign \new_[99663]_  = \new_[99662]_  & \new_[99655]_ ;
  assign \new_[99666]_  = A266 & ~A265;
  assign \new_[99669]_  = A268 & A267;
  assign \new_[99670]_  = \new_[99669]_  & \new_[99666]_ ;
  assign \new_[99673]_  = A299 & ~A298;
  assign \new_[99676]_  = A301 & A300;
  assign \new_[99677]_  = \new_[99676]_  & \new_[99673]_ ;
  assign \new_[99678]_  = \new_[99677]_  & \new_[99670]_ ;
  assign \new_[99681]_  = ~A169 & ~A170;
  assign \new_[99684]_  = ~A199 & A168;
  assign \new_[99685]_  = \new_[99684]_  & \new_[99681]_ ;
  assign \new_[99688]_  = ~A201 & A200;
  assign \new_[99691]_  = A203 & ~A202;
  assign \new_[99692]_  = \new_[99691]_  & \new_[99688]_ ;
  assign \new_[99693]_  = \new_[99692]_  & \new_[99685]_ ;
  assign \new_[99696]_  = A266 & ~A265;
  assign \new_[99699]_  = A268 & A267;
  assign \new_[99700]_  = \new_[99699]_  & \new_[99696]_ ;
  assign \new_[99703]_  = A299 & ~A298;
  assign \new_[99706]_  = ~A302 & A300;
  assign \new_[99707]_  = \new_[99706]_  & \new_[99703]_ ;
  assign \new_[99708]_  = \new_[99707]_  & \new_[99700]_ ;
  assign \new_[99711]_  = ~A169 & ~A170;
  assign \new_[99714]_  = ~A199 & A168;
  assign \new_[99715]_  = \new_[99714]_  & \new_[99711]_ ;
  assign \new_[99718]_  = ~A201 & A200;
  assign \new_[99721]_  = A203 & ~A202;
  assign \new_[99722]_  = \new_[99721]_  & \new_[99718]_ ;
  assign \new_[99723]_  = \new_[99722]_  & \new_[99715]_ ;
  assign \new_[99726]_  = A266 & ~A265;
  assign \new_[99729]_  = ~A269 & A267;
  assign \new_[99730]_  = \new_[99729]_  & \new_[99726]_ ;
  assign \new_[99733]_  = ~A299 & A298;
  assign \new_[99736]_  = A301 & A300;
  assign \new_[99737]_  = \new_[99736]_  & \new_[99733]_ ;
  assign \new_[99738]_  = \new_[99737]_  & \new_[99730]_ ;
  assign \new_[99741]_  = ~A169 & ~A170;
  assign \new_[99744]_  = ~A199 & A168;
  assign \new_[99745]_  = \new_[99744]_  & \new_[99741]_ ;
  assign \new_[99748]_  = ~A201 & A200;
  assign \new_[99751]_  = A203 & ~A202;
  assign \new_[99752]_  = \new_[99751]_  & \new_[99748]_ ;
  assign \new_[99753]_  = \new_[99752]_  & \new_[99745]_ ;
  assign \new_[99756]_  = A266 & ~A265;
  assign \new_[99759]_  = ~A269 & A267;
  assign \new_[99760]_  = \new_[99759]_  & \new_[99756]_ ;
  assign \new_[99763]_  = ~A299 & A298;
  assign \new_[99766]_  = ~A302 & A300;
  assign \new_[99767]_  = \new_[99766]_  & \new_[99763]_ ;
  assign \new_[99768]_  = \new_[99767]_  & \new_[99760]_ ;
  assign \new_[99771]_  = ~A169 & ~A170;
  assign \new_[99774]_  = ~A199 & A168;
  assign \new_[99775]_  = \new_[99774]_  & \new_[99771]_ ;
  assign \new_[99778]_  = ~A201 & A200;
  assign \new_[99781]_  = A203 & ~A202;
  assign \new_[99782]_  = \new_[99781]_  & \new_[99778]_ ;
  assign \new_[99783]_  = \new_[99782]_  & \new_[99775]_ ;
  assign \new_[99786]_  = A266 & ~A265;
  assign \new_[99789]_  = ~A269 & A267;
  assign \new_[99790]_  = \new_[99789]_  & \new_[99786]_ ;
  assign \new_[99793]_  = A299 & ~A298;
  assign \new_[99796]_  = A301 & A300;
  assign \new_[99797]_  = \new_[99796]_  & \new_[99793]_ ;
  assign \new_[99798]_  = \new_[99797]_  & \new_[99790]_ ;
  assign \new_[99801]_  = ~A169 & ~A170;
  assign \new_[99804]_  = ~A199 & A168;
  assign \new_[99805]_  = \new_[99804]_  & \new_[99801]_ ;
  assign \new_[99808]_  = ~A201 & A200;
  assign \new_[99811]_  = A203 & ~A202;
  assign \new_[99812]_  = \new_[99811]_  & \new_[99808]_ ;
  assign \new_[99813]_  = \new_[99812]_  & \new_[99805]_ ;
  assign \new_[99816]_  = A266 & ~A265;
  assign \new_[99819]_  = ~A269 & A267;
  assign \new_[99820]_  = \new_[99819]_  & \new_[99816]_ ;
  assign \new_[99823]_  = A299 & ~A298;
  assign \new_[99826]_  = ~A302 & A300;
  assign \new_[99827]_  = \new_[99826]_  & \new_[99823]_ ;
  assign \new_[99828]_  = \new_[99827]_  & \new_[99820]_ ;
  assign \new_[99831]_  = ~A169 & ~A170;
  assign \new_[99834]_  = ~A199 & A168;
  assign \new_[99835]_  = \new_[99834]_  & \new_[99831]_ ;
  assign \new_[99838]_  = ~A201 & A200;
  assign \new_[99841]_  = A203 & ~A202;
  assign \new_[99842]_  = \new_[99841]_  & \new_[99838]_ ;
  assign \new_[99843]_  = \new_[99842]_  & \new_[99835]_ ;
  assign \new_[99846]_  = ~A266 & A265;
  assign \new_[99849]_  = A268 & A267;
  assign \new_[99850]_  = \new_[99849]_  & \new_[99846]_ ;
  assign \new_[99853]_  = ~A299 & A298;
  assign \new_[99856]_  = A301 & A300;
  assign \new_[99857]_  = \new_[99856]_  & \new_[99853]_ ;
  assign \new_[99858]_  = \new_[99857]_  & \new_[99850]_ ;
  assign \new_[99861]_  = ~A169 & ~A170;
  assign \new_[99864]_  = ~A199 & A168;
  assign \new_[99865]_  = \new_[99864]_  & \new_[99861]_ ;
  assign \new_[99868]_  = ~A201 & A200;
  assign \new_[99871]_  = A203 & ~A202;
  assign \new_[99872]_  = \new_[99871]_  & \new_[99868]_ ;
  assign \new_[99873]_  = \new_[99872]_  & \new_[99865]_ ;
  assign \new_[99876]_  = ~A266 & A265;
  assign \new_[99879]_  = A268 & A267;
  assign \new_[99880]_  = \new_[99879]_  & \new_[99876]_ ;
  assign \new_[99883]_  = ~A299 & A298;
  assign \new_[99886]_  = ~A302 & A300;
  assign \new_[99887]_  = \new_[99886]_  & \new_[99883]_ ;
  assign \new_[99888]_  = \new_[99887]_  & \new_[99880]_ ;
  assign \new_[99891]_  = ~A169 & ~A170;
  assign \new_[99894]_  = ~A199 & A168;
  assign \new_[99895]_  = \new_[99894]_  & \new_[99891]_ ;
  assign \new_[99898]_  = ~A201 & A200;
  assign \new_[99901]_  = A203 & ~A202;
  assign \new_[99902]_  = \new_[99901]_  & \new_[99898]_ ;
  assign \new_[99903]_  = \new_[99902]_  & \new_[99895]_ ;
  assign \new_[99906]_  = ~A266 & A265;
  assign \new_[99909]_  = A268 & A267;
  assign \new_[99910]_  = \new_[99909]_  & \new_[99906]_ ;
  assign \new_[99913]_  = A299 & ~A298;
  assign \new_[99916]_  = A301 & A300;
  assign \new_[99917]_  = \new_[99916]_  & \new_[99913]_ ;
  assign \new_[99918]_  = \new_[99917]_  & \new_[99910]_ ;
  assign \new_[99921]_  = ~A169 & ~A170;
  assign \new_[99924]_  = ~A199 & A168;
  assign \new_[99925]_  = \new_[99924]_  & \new_[99921]_ ;
  assign \new_[99928]_  = ~A201 & A200;
  assign \new_[99931]_  = A203 & ~A202;
  assign \new_[99932]_  = \new_[99931]_  & \new_[99928]_ ;
  assign \new_[99933]_  = \new_[99932]_  & \new_[99925]_ ;
  assign \new_[99936]_  = ~A266 & A265;
  assign \new_[99939]_  = A268 & A267;
  assign \new_[99940]_  = \new_[99939]_  & \new_[99936]_ ;
  assign \new_[99943]_  = A299 & ~A298;
  assign \new_[99946]_  = ~A302 & A300;
  assign \new_[99947]_  = \new_[99946]_  & \new_[99943]_ ;
  assign \new_[99948]_  = \new_[99947]_  & \new_[99940]_ ;
  assign \new_[99951]_  = ~A169 & ~A170;
  assign \new_[99954]_  = ~A199 & A168;
  assign \new_[99955]_  = \new_[99954]_  & \new_[99951]_ ;
  assign \new_[99958]_  = ~A201 & A200;
  assign \new_[99961]_  = A203 & ~A202;
  assign \new_[99962]_  = \new_[99961]_  & \new_[99958]_ ;
  assign \new_[99963]_  = \new_[99962]_  & \new_[99955]_ ;
  assign \new_[99966]_  = ~A266 & A265;
  assign \new_[99969]_  = ~A269 & A267;
  assign \new_[99970]_  = \new_[99969]_  & \new_[99966]_ ;
  assign \new_[99973]_  = ~A299 & A298;
  assign \new_[99976]_  = A301 & A300;
  assign \new_[99977]_  = \new_[99976]_  & \new_[99973]_ ;
  assign \new_[99978]_  = \new_[99977]_  & \new_[99970]_ ;
  assign \new_[99981]_  = ~A169 & ~A170;
  assign \new_[99984]_  = ~A199 & A168;
  assign \new_[99985]_  = \new_[99984]_  & \new_[99981]_ ;
  assign \new_[99988]_  = ~A201 & A200;
  assign \new_[99991]_  = A203 & ~A202;
  assign \new_[99992]_  = \new_[99991]_  & \new_[99988]_ ;
  assign \new_[99993]_  = \new_[99992]_  & \new_[99985]_ ;
  assign \new_[99996]_  = ~A266 & A265;
  assign \new_[99999]_  = ~A269 & A267;
  assign \new_[100000]_  = \new_[99999]_  & \new_[99996]_ ;
  assign \new_[100003]_  = ~A299 & A298;
  assign \new_[100006]_  = ~A302 & A300;
  assign \new_[100007]_  = \new_[100006]_  & \new_[100003]_ ;
  assign \new_[100008]_  = \new_[100007]_  & \new_[100000]_ ;
  assign \new_[100011]_  = ~A169 & ~A170;
  assign \new_[100014]_  = ~A199 & A168;
  assign \new_[100015]_  = \new_[100014]_  & \new_[100011]_ ;
  assign \new_[100018]_  = ~A201 & A200;
  assign \new_[100021]_  = A203 & ~A202;
  assign \new_[100022]_  = \new_[100021]_  & \new_[100018]_ ;
  assign \new_[100023]_  = \new_[100022]_  & \new_[100015]_ ;
  assign \new_[100026]_  = ~A266 & A265;
  assign \new_[100029]_  = ~A269 & A267;
  assign \new_[100030]_  = \new_[100029]_  & \new_[100026]_ ;
  assign \new_[100033]_  = A299 & ~A298;
  assign \new_[100036]_  = A301 & A300;
  assign \new_[100037]_  = \new_[100036]_  & \new_[100033]_ ;
  assign \new_[100038]_  = \new_[100037]_  & \new_[100030]_ ;
  assign \new_[100041]_  = ~A169 & ~A170;
  assign \new_[100044]_  = ~A199 & A168;
  assign \new_[100045]_  = \new_[100044]_  & \new_[100041]_ ;
  assign \new_[100048]_  = ~A201 & A200;
  assign \new_[100051]_  = A203 & ~A202;
  assign \new_[100052]_  = \new_[100051]_  & \new_[100048]_ ;
  assign \new_[100053]_  = \new_[100052]_  & \new_[100045]_ ;
  assign \new_[100056]_  = ~A266 & A265;
  assign \new_[100059]_  = ~A269 & A267;
  assign \new_[100060]_  = \new_[100059]_  & \new_[100056]_ ;
  assign \new_[100063]_  = A299 & ~A298;
  assign \new_[100066]_  = ~A302 & A300;
  assign \new_[100067]_  = \new_[100066]_  & \new_[100063]_ ;
  assign \new_[100068]_  = \new_[100067]_  & \new_[100060]_ ;
  assign \new_[100071]_  = ~A169 & ~A170;
  assign \new_[100074]_  = A199 & A168;
  assign \new_[100075]_  = \new_[100074]_  & \new_[100071]_ ;
  assign \new_[100078]_  = A201 & ~A200;
  assign \new_[100081]_  = ~A265 & A202;
  assign \new_[100082]_  = \new_[100081]_  & \new_[100078]_ ;
  assign \new_[100083]_  = \new_[100082]_  & \new_[100075]_ ;
  assign \new_[100086]_  = A267 & A266;
  assign \new_[100089]_  = A298 & A268;
  assign \new_[100090]_  = \new_[100089]_  & \new_[100086]_ ;
  assign \new_[100093]_  = ~A300 & ~A299;
  assign \new_[100096]_  = A302 & ~A301;
  assign \new_[100097]_  = \new_[100096]_  & \new_[100093]_ ;
  assign \new_[100098]_  = \new_[100097]_  & \new_[100090]_ ;
  assign \new_[100101]_  = ~A169 & ~A170;
  assign \new_[100104]_  = A199 & A168;
  assign \new_[100105]_  = \new_[100104]_  & \new_[100101]_ ;
  assign \new_[100108]_  = A201 & ~A200;
  assign \new_[100111]_  = ~A265 & A202;
  assign \new_[100112]_  = \new_[100111]_  & \new_[100108]_ ;
  assign \new_[100113]_  = \new_[100112]_  & \new_[100105]_ ;
  assign \new_[100116]_  = A267 & A266;
  assign \new_[100119]_  = ~A298 & A268;
  assign \new_[100120]_  = \new_[100119]_  & \new_[100116]_ ;
  assign \new_[100123]_  = ~A300 & A299;
  assign \new_[100126]_  = A302 & ~A301;
  assign \new_[100127]_  = \new_[100126]_  & \new_[100123]_ ;
  assign \new_[100128]_  = \new_[100127]_  & \new_[100120]_ ;
  assign \new_[100131]_  = ~A169 & ~A170;
  assign \new_[100134]_  = A199 & A168;
  assign \new_[100135]_  = \new_[100134]_  & \new_[100131]_ ;
  assign \new_[100138]_  = A201 & ~A200;
  assign \new_[100141]_  = ~A265 & A202;
  assign \new_[100142]_  = \new_[100141]_  & \new_[100138]_ ;
  assign \new_[100143]_  = \new_[100142]_  & \new_[100135]_ ;
  assign \new_[100146]_  = A267 & A266;
  assign \new_[100149]_  = A298 & ~A269;
  assign \new_[100150]_  = \new_[100149]_  & \new_[100146]_ ;
  assign \new_[100153]_  = ~A300 & ~A299;
  assign \new_[100156]_  = A302 & ~A301;
  assign \new_[100157]_  = \new_[100156]_  & \new_[100153]_ ;
  assign \new_[100158]_  = \new_[100157]_  & \new_[100150]_ ;
  assign \new_[100161]_  = ~A169 & ~A170;
  assign \new_[100164]_  = A199 & A168;
  assign \new_[100165]_  = \new_[100164]_  & \new_[100161]_ ;
  assign \new_[100168]_  = A201 & ~A200;
  assign \new_[100171]_  = ~A265 & A202;
  assign \new_[100172]_  = \new_[100171]_  & \new_[100168]_ ;
  assign \new_[100173]_  = \new_[100172]_  & \new_[100165]_ ;
  assign \new_[100176]_  = A267 & A266;
  assign \new_[100179]_  = ~A298 & ~A269;
  assign \new_[100180]_  = \new_[100179]_  & \new_[100176]_ ;
  assign \new_[100183]_  = ~A300 & A299;
  assign \new_[100186]_  = A302 & ~A301;
  assign \new_[100187]_  = \new_[100186]_  & \new_[100183]_ ;
  assign \new_[100188]_  = \new_[100187]_  & \new_[100180]_ ;
  assign \new_[100191]_  = ~A169 & ~A170;
  assign \new_[100194]_  = A199 & A168;
  assign \new_[100195]_  = \new_[100194]_  & \new_[100191]_ ;
  assign \new_[100198]_  = A201 & ~A200;
  assign \new_[100201]_  = ~A265 & A202;
  assign \new_[100202]_  = \new_[100201]_  & \new_[100198]_ ;
  assign \new_[100203]_  = \new_[100202]_  & \new_[100195]_ ;
  assign \new_[100206]_  = ~A267 & A266;
  assign \new_[100209]_  = A269 & ~A268;
  assign \new_[100210]_  = \new_[100209]_  & \new_[100206]_ ;
  assign \new_[100213]_  = ~A299 & A298;
  assign \new_[100216]_  = A301 & A300;
  assign \new_[100217]_  = \new_[100216]_  & \new_[100213]_ ;
  assign \new_[100218]_  = \new_[100217]_  & \new_[100210]_ ;
  assign \new_[100221]_  = ~A169 & ~A170;
  assign \new_[100224]_  = A199 & A168;
  assign \new_[100225]_  = \new_[100224]_  & \new_[100221]_ ;
  assign \new_[100228]_  = A201 & ~A200;
  assign \new_[100231]_  = ~A265 & A202;
  assign \new_[100232]_  = \new_[100231]_  & \new_[100228]_ ;
  assign \new_[100233]_  = \new_[100232]_  & \new_[100225]_ ;
  assign \new_[100236]_  = ~A267 & A266;
  assign \new_[100239]_  = A269 & ~A268;
  assign \new_[100240]_  = \new_[100239]_  & \new_[100236]_ ;
  assign \new_[100243]_  = ~A299 & A298;
  assign \new_[100246]_  = ~A302 & A300;
  assign \new_[100247]_  = \new_[100246]_  & \new_[100243]_ ;
  assign \new_[100248]_  = \new_[100247]_  & \new_[100240]_ ;
  assign \new_[100251]_  = ~A169 & ~A170;
  assign \new_[100254]_  = A199 & A168;
  assign \new_[100255]_  = \new_[100254]_  & \new_[100251]_ ;
  assign \new_[100258]_  = A201 & ~A200;
  assign \new_[100261]_  = ~A265 & A202;
  assign \new_[100262]_  = \new_[100261]_  & \new_[100258]_ ;
  assign \new_[100263]_  = \new_[100262]_  & \new_[100255]_ ;
  assign \new_[100266]_  = ~A267 & A266;
  assign \new_[100269]_  = A269 & ~A268;
  assign \new_[100270]_  = \new_[100269]_  & \new_[100266]_ ;
  assign \new_[100273]_  = A299 & ~A298;
  assign \new_[100276]_  = A301 & A300;
  assign \new_[100277]_  = \new_[100276]_  & \new_[100273]_ ;
  assign \new_[100278]_  = \new_[100277]_  & \new_[100270]_ ;
  assign \new_[100281]_  = ~A169 & ~A170;
  assign \new_[100284]_  = A199 & A168;
  assign \new_[100285]_  = \new_[100284]_  & \new_[100281]_ ;
  assign \new_[100288]_  = A201 & ~A200;
  assign \new_[100291]_  = ~A265 & A202;
  assign \new_[100292]_  = \new_[100291]_  & \new_[100288]_ ;
  assign \new_[100293]_  = \new_[100292]_  & \new_[100285]_ ;
  assign \new_[100296]_  = ~A267 & A266;
  assign \new_[100299]_  = A269 & ~A268;
  assign \new_[100300]_  = \new_[100299]_  & \new_[100296]_ ;
  assign \new_[100303]_  = A299 & ~A298;
  assign \new_[100306]_  = ~A302 & A300;
  assign \new_[100307]_  = \new_[100306]_  & \new_[100303]_ ;
  assign \new_[100308]_  = \new_[100307]_  & \new_[100300]_ ;
  assign \new_[100311]_  = ~A169 & ~A170;
  assign \new_[100314]_  = A199 & A168;
  assign \new_[100315]_  = \new_[100314]_  & \new_[100311]_ ;
  assign \new_[100318]_  = A201 & ~A200;
  assign \new_[100321]_  = A265 & A202;
  assign \new_[100322]_  = \new_[100321]_  & \new_[100318]_ ;
  assign \new_[100323]_  = \new_[100322]_  & \new_[100315]_ ;
  assign \new_[100326]_  = A267 & ~A266;
  assign \new_[100329]_  = A298 & A268;
  assign \new_[100330]_  = \new_[100329]_  & \new_[100326]_ ;
  assign \new_[100333]_  = ~A300 & ~A299;
  assign \new_[100336]_  = A302 & ~A301;
  assign \new_[100337]_  = \new_[100336]_  & \new_[100333]_ ;
  assign \new_[100338]_  = \new_[100337]_  & \new_[100330]_ ;
  assign \new_[100341]_  = ~A169 & ~A170;
  assign \new_[100344]_  = A199 & A168;
  assign \new_[100345]_  = \new_[100344]_  & \new_[100341]_ ;
  assign \new_[100348]_  = A201 & ~A200;
  assign \new_[100351]_  = A265 & A202;
  assign \new_[100352]_  = \new_[100351]_  & \new_[100348]_ ;
  assign \new_[100353]_  = \new_[100352]_  & \new_[100345]_ ;
  assign \new_[100356]_  = A267 & ~A266;
  assign \new_[100359]_  = ~A298 & A268;
  assign \new_[100360]_  = \new_[100359]_  & \new_[100356]_ ;
  assign \new_[100363]_  = ~A300 & A299;
  assign \new_[100366]_  = A302 & ~A301;
  assign \new_[100367]_  = \new_[100366]_  & \new_[100363]_ ;
  assign \new_[100368]_  = \new_[100367]_  & \new_[100360]_ ;
  assign \new_[100371]_  = ~A169 & ~A170;
  assign \new_[100374]_  = A199 & A168;
  assign \new_[100375]_  = \new_[100374]_  & \new_[100371]_ ;
  assign \new_[100378]_  = A201 & ~A200;
  assign \new_[100381]_  = A265 & A202;
  assign \new_[100382]_  = \new_[100381]_  & \new_[100378]_ ;
  assign \new_[100383]_  = \new_[100382]_  & \new_[100375]_ ;
  assign \new_[100386]_  = A267 & ~A266;
  assign \new_[100389]_  = A298 & ~A269;
  assign \new_[100390]_  = \new_[100389]_  & \new_[100386]_ ;
  assign \new_[100393]_  = ~A300 & ~A299;
  assign \new_[100396]_  = A302 & ~A301;
  assign \new_[100397]_  = \new_[100396]_  & \new_[100393]_ ;
  assign \new_[100398]_  = \new_[100397]_  & \new_[100390]_ ;
  assign \new_[100401]_  = ~A169 & ~A170;
  assign \new_[100404]_  = A199 & A168;
  assign \new_[100405]_  = \new_[100404]_  & \new_[100401]_ ;
  assign \new_[100408]_  = A201 & ~A200;
  assign \new_[100411]_  = A265 & A202;
  assign \new_[100412]_  = \new_[100411]_  & \new_[100408]_ ;
  assign \new_[100413]_  = \new_[100412]_  & \new_[100405]_ ;
  assign \new_[100416]_  = A267 & ~A266;
  assign \new_[100419]_  = ~A298 & ~A269;
  assign \new_[100420]_  = \new_[100419]_  & \new_[100416]_ ;
  assign \new_[100423]_  = ~A300 & A299;
  assign \new_[100426]_  = A302 & ~A301;
  assign \new_[100427]_  = \new_[100426]_  & \new_[100423]_ ;
  assign \new_[100428]_  = \new_[100427]_  & \new_[100420]_ ;
  assign \new_[100431]_  = ~A169 & ~A170;
  assign \new_[100434]_  = A199 & A168;
  assign \new_[100435]_  = \new_[100434]_  & \new_[100431]_ ;
  assign \new_[100438]_  = A201 & ~A200;
  assign \new_[100441]_  = A265 & A202;
  assign \new_[100442]_  = \new_[100441]_  & \new_[100438]_ ;
  assign \new_[100443]_  = \new_[100442]_  & \new_[100435]_ ;
  assign \new_[100446]_  = ~A267 & ~A266;
  assign \new_[100449]_  = A269 & ~A268;
  assign \new_[100450]_  = \new_[100449]_  & \new_[100446]_ ;
  assign \new_[100453]_  = ~A299 & A298;
  assign \new_[100456]_  = A301 & A300;
  assign \new_[100457]_  = \new_[100456]_  & \new_[100453]_ ;
  assign \new_[100458]_  = \new_[100457]_  & \new_[100450]_ ;
  assign \new_[100461]_  = ~A169 & ~A170;
  assign \new_[100464]_  = A199 & A168;
  assign \new_[100465]_  = \new_[100464]_  & \new_[100461]_ ;
  assign \new_[100468]_  = A201 & ~A200;
  assign \new_[100471]_  = A265 & A202;
  assign \new_[100472]_  = \new_[100471]_  & \new_[100468]_ ;
  assign \new_[100473]_  = \new_[100472]_  & \new_[100465]_ ;
  assign \new_[100476]_  = ~A267 & ~A266;
  assign \new_[100479]_  = A269 & ~A268;
  assign \new_[100480]_  = \new_[100479]_  & \new_[100476]_ ;
  assign \new_[100483]_  = ~A299 & A298;
  assign \new_[100486]_  = ~A302 & A300;
  assign \new_[100487]_  = \new_[100486]_  & \new_[100483]_ ;
  assign \new_[100488]_  = \new_[100487]_  & \new_[100480]_ ;
  assign \new_[100491]_  = ~A169 & ~A170;
  assign \new_[100494]_  = A199 & A168;
  assign \new_[100495]_  = \new_[100494]_  & \new_[100491]_ ;
  assign \new_[100498]_  = A201 & ~A200;
  assign \new_[100501]_  = A265 & A202;
  assign \new_[100502]_  = \new_[100501]_  & \new_[100498]_ ;
  assign \new_[100503]_  = \new_[100502]_  & \new_[100495]_ ;
  assign \new_[100506]_  = ~A267 & ~A266;
  assign \new_[100509]_  = A269 & ~A268;
  assign \new_[100510]_  = \new_[100509]_  & \new_[100506]_ ;
  assign \new_[100513]_  = A299 & ~A298;
  assign \new_[100516]_  = A301 & A300;
  assign \new_[100517]_  = \new_[100516]_  & \new_[100513]_ ;
  assign \new_[100518]_  = \new_[100517]_  & \new_[100510]_ ;
  assign \new_[100521]_  = ~A169 & ~A170;
  assign \new_[100524]_  = A199 & A168;
  assign \new_[100525]_  = \new_[100524]_  & \new_[100521]_ ;
  assign \new_[100528]_  = A201 & ~A200;
  assign \new_[100531]_  = A265 & A202;
  assign \new_[100532]_  = \new_[100531]_  & \new_[100528]_ ;
  assign \new_[100533]_  = \new_[100532]_  & \new_[100525]_ ;
  assign \new_[100536]_  = ~A267 & ~A266;
  assign \new_[100539]_  = A269 & ~A268;
  assign \new_[100540]_  = \new_[100539]_  & \new_[100536]_ ;
  assign \new_[100543]_  = A299 & ~A298;
  assign \new_[100546]_  = ~A302 & A300;
  assign \new_[100547]_  = \new_[100546]_  & \new_[100543]_ ;
  assign \new_[100548]_  = \new_[100547]_  & \new_[100540]_ ;
  assign \new_[100551]_  = ~A169 & ~A170;
  assign \new_[100554]_  = A199 & A168;
  assign \new_[100555]_  = \new_[100554]_  & \new_[100551]_ ;
  assign \new_[100558]_  = A201 & ~A200;
  assign \new_[100561]_  = ~A265 & ~A203;
  assign \new_[100562]_  = \new_[100561]_  & \new_[100558]_ ;
  assign \new_[100563]_  = \new_[100562]_  & \new_[100555]_ ;
  assign \new_[100566]_  = A267 & A266;
  assign \new_[100569]_  = A298 & A268;
  assign \new_[100570]_  = \new_[100569]_  & \new_[100566]_ ;
  assign \new_[100573]_  = ~A300 & ~A299;
  assign \new_[100576]_  = A302 & ~A301;
  assign \new_[100577]_  = \new_[100576]_  & \new_[100573]_ ;
  assign \new_[100578]_  = \new_[100577]_  & \new_[100570]_ ;
  assign \new_[100581]_  = ~A169 & ~A170;
  assign \new_[100584]_  = A199 & A168;
  assign \new_[100585]_  = \new_[100584]_  & \new_[100581]_ ;
  assign \new_[100588]_  = A201 & ~A200;
  assign \new_[100591]_  = ~A265 & ~A203;
  assign \new_[100592]_  = \new_[100591]_  & \new_[100588]_ ;
  assign \new_[100593]_  = \new_[100592]_  & \new_[100585]_ ;
  assign \new_[100596]_  = A267 & A266;
  assign \new_[100599]_  = ~A298 & A268;
  assign \new_[100600]_  = \new_[100599]_  & \new_[100596]_ ;
  assign \new_[100603]_  = ~A300 & A299;
  assign \new_[100606]_  = A302 & ~A301;
  assign \new_[100607]_  = \new_[100606]_  & \new_[100603]_ ;
  assign \new_[100608]_  = \new_[100607]_  & \new_[100600]_ ;
  assign \new_[100611]_  = ~A169 & ~A170;
  assign \new_[100614]_  = A199 & A168;
  assign \new_[100615]_  = \new_[100614]_  & \new_[100611]_ ;
  assign \new_[100618]_  = A201 & ~A200;
  assign \new_[100621]_  = ~A265 & ~A203;
  assign \new_[100622]_  = \new_[100621]_  & \new_[100618]_ ;
  assign \new_[100623]_  = \new_[100622]_  & \new_[100615]_ ;
  assign \new_[100626]_  = A267 & A266;
  assign \new_[100629]_  = A298 & ~A269;
  assign \new_[100630]_  = \new_[100629]_  & \new_[100626]_ ;
  assign \new_[100633]_  = ~A300 & ~A299;
  assign \new_[100636]_  = A302 & ~A301;
  assign \new_[100637]_  = \new_[100636]_  & \new_[100633]_ ;
  assign \new_[100638]_  = \new_[100637]_  & \new_[100630]_ ;
  assign \new_[100641]_  = ~A169 & ~A170;
  assign \new_[100644]_  = A199 & A168;
  assign \new_[100645]_  = \new_[100644]_  & \new_[100641]_ ;
  assign \new_[100648]_  = A201 & ~A200;
  assign \new_[100651]_  = ~A265 & ~A203;
  assign \new_[100652]_  = \new_[100651]_  & \new_[100648]_ ;
  assign \new_[100653]_  = \new_[100652]_  & \new_[100645]_ ;
  assign \new_[100656]_  = A267 & A266;
  assign \new_[100659]_  = ~A298 & ~A269;
  assign \new_[100660]_  = \new_[100659]_  & \new_[100656]_ ;
  assign \new_[100663]_  = ~A300 & A299;
  assign \new_[100666]_  = A302 & ~A301;
  assign \new_[100667]_  = \new_[100666]_  & \new_[100663]_ ;
  assign \new_[100668]_  = \new_[100667]_  & \new_[100660]_ ;
  assign \new_[100671]_  = ~A169 & ~A170;
  assign \new_[100674]_  = A199 & A168;
  assign \new_[100675]_  = \new_[100674]_  & \new_[100671]_ ;
  assign \new_[100678]_  = A201 & ~A200;
  assign \new_[100681]_  = ~A265 & ~A203;
  assign \new_[100682]_  = \new_[100681]_  & \new_[100678]_ ;
  assign \new_[100683]_  = \new_[100682]_  & \new_[100675]_ ;
  assign \new_[100686]_  = ~A267 & A266;
  assign \new_[100689]_  = A269 & ~A268;
  assign \new_[100690]_  = \new_[100689]_  & \new_[100686]_ ;
  assign \new_[100693]_  = ~A299 & A298;
  assign \new_[100696]_  = A301 & A300;
  assign \new_[100697]_  = \new_[100696]_  & \new_[100693]_ ;
  assign \new_[100698]_  = \new_[100697]_  & \new_[100690]_ ;
  assign \new_[100701]_  = ~A169 & ~A170;
  assign \new_[100704]_  = A199 & A168;
  assign \new_[100705]_  = \new_[100704]_  & \new_[100701]_ ;
  assign \new_[100708]_  = A201 & ~A200;
  assign \new_[100711]_  = ~A265 & ~A203;
  assign \new_[100712]_  = \new_[100711]_  & \new_[100708]_ ;
  assign \new_[100713]_  = \new_[100712]_  & \new_[100705]_ ;
  assign \new_[100716]_  = ~A267 & A266;
  assign \new_[100719]_  = A269 & ~A268;
  assign \new_[100720]_  = \new_[100719]_  & \new_[100716]_ ;
  assign \new_[100723]_  = ~A299 & A298;
  assign \new_[100726]_  = ~A302 & A300;
  assign \new_[100727]_  = \new_[100726]_  & \new_[100723]_ ;
  assign \new_[100728]_  = \new_[100727]_  & \new_[100720]_ ;
  assign \new_[100731]_  = ~A169 & ~A170;
  assign \new_[100734]_  = A199 & A168;
  assign \new_[100735]_  = \new_[100734]_  & \new_[100731]_ ;
  assign \new_[100738]_  = A201 & ~A200;
  assign \new_[100741]_  = ~A265 & ~A203;
  assign \new_[100742]_  = \new_[100741]_  & \new_[100738]_ ;
  assign \new_[100743]_  = \new_[100742]_  & \new_[100735]_ ;
  assign \new_[100746]_  = ~A267 & A266;
  assign \new_[100749]_  = A269 & ~A268;
  assign \new_[100750]_  = \new_[100749]_  & \new_[100746]_ ;
  assign \new_[100753]_  = A299 & ~A298;
  assign \new_[100756]_  = A301 & A300;
  assign \new_[100757]_  = \new_[100756]_  & \new_[100753]_ ;
  assign \new_[100758]_  = \new_[100757]_  & \new_[100750]_ ;
  assign \new_[100761]_  = ~A169 & ~A170;
  assign \new_[100764]_  = A199 & A168;
  assign \new_[100765]_  = \new_[100764]_  & \new_[100761]_ ;
  assign \new_[100768]_  = A201 & ~A200;
  assign \new_[100771]_  = ~A265 & ~A203;
  assign \new_[100772]_  = \new_[100771]_  & \new_[100768]_ ;
  assign \new_[100773]_  = \new_[100772]_  & \new_[100765]_ ;
  assign \new_[100776]_  = ~A267 & A266;
  assign \new_[100779]_  = A269 & ~A268;
  assign \new_[100780]_  = \new_[100779]_  & \new_[100776]_ ;
  assign \new_[100783]_  = A299 & ~A298;
  assign \new_[100786]_  = ~A302 & A300;
  assign \new_[100787]_  = \new_[100786]_  & \new_[100783]_ ;
  assign \new_[100788]_  = \new_[100787]_  & \new_[100780]_ ;
  assign \new_[100791]_  = ~A169 & ~A170;
  assign \new_[100794]_  = A199 & A168;
  assign \new_[100795]_  = \new_[100794]_  & \new_[100791]_ ;
  assign \new_[100798]_  = A201 & ~A200;
  assign \new_[100801]_  = A265 & ~A203;
  assign \new_[100802]_  = \new_[100801]_  & \new_[100798]_ ;
  assign \new_[100803]_  = \new_[100802]_  & \new_[100795]_ ;
  assign \new_[100806]_  = A267 & ~A266;
  assign \new_[100809]_  = A298 & A268;
  assign \new_[100810]_  = \new_[100809]_  & \new_[100806]_ ;
  assign \new_[100813]_  = ~A300 & ~A299;
  assign \new_[100816]_  = A302 & ~A301;
  assign \new_[100817]_  = \new_[100816]_  & \new_[100813]_ ;
  assign \new_[100818]_  = \new_[100817]_  & \new_[100810]_ ;
  assign \new_[100821]_  = ~A169 & ~A170;
  assign \new_[100824]_  = A199 & A168;
  assign \new_[100825]_  = \new_[100824]_  & \new_[100821]_ ;
  assign \new_[100828]_  = A201 & ~A200;
  assign \new_[100831]_  = A265 & ~A203;
  assign \new_[100832]_  = \new_[100831]_  & \new_[100828]_ ;
  assign \new_[100833]_  = \new_[100832]_  & \new_[100825]_ ;
  assign \new_[100836]_  = A267 & ~A266;
  assign \new_[100839]_  = ~A298 & A268;
  assign \new_[100840]_  = \new_[100839]_  & \new_[100836]_ ;
  assign \new_[100843]_  = ~A300 & A299;
  assign \new_[100846]_  = A302 & ~A301;
  assign \new_[100847]_  = \new_[100846]_  & \new_[100843]_ ;
  assign \new_[100848]_  = \new_[100847]_  & \new_[100840]_ ;
  assign \new_[100851]_  = ~A169 & ~A170;
  assign \new_[100854]_  = A199 & A168;
  assign \new_[100855]_  = \new_[100854]_  & \new_[100851]_ ;
  assign \new_[100858]_  = A201 & ~A200;
  assign \new_[100861]_  = A265 & ~A203;
  assign \new_[100862]_  = \new_[100861]_  & \new_[100858]_ ;
  assign \new_[100863]_  = \new_[100862]_  & \new_[100855]_ ;
  assign \new_[100866]_  = A267 & ~A266;
  assign \new_[100869]_  = A298 & ~A269;
  assign \new_[100870]_  = \new_[100869]_  & \new_[100866]_ ;
  assign \new_[100873]_  = ~A300 & ~A299;
  assign \new_[100876]_  = A302 & ~A301;
  assign \new_[100877]_  = \new_[100876]_  & \new_[100873]_ ;
  assign \new_[100878]_  = \new_[100877]_  & \new_[100870]_ ;
  assign \new_[100881]_  = ~A169 & ~A170;
  assign \new_[100884]_  = A199 & A168;
  assign \new_[100885]_  = \new_[100884]_  & \new_[100881]_ ;
  assign \new_[100888]_  = A201 & ~A200;
  assign \new_[100891]_  = A265 & ~A203;
  assign \new_[100892]_  = \new_[100891]_  & \new_[100888]_ ;
  assign \new_[100893]_  = \new_[100892]_  & \new_[100885]_ ;
  assign \new_[100896]_  = A267 & ~A266;
  assign \new_[100899]_  = ~A298 & ~A269;
  assign \new_[100900]_  = \new_[100899]_  & \new_[100896]_ ;
  assign \new_[100903]_  = ~A300 & A299;
  assign \new_[100906]_  = A302 & ~A301;
  assign \new_[100907]_  = \new_[100906]_  & \new_[100903]_ ;
  assign \new_[100908]_  = \new_[100907]_  & \new_[100900]_ ;
  assign \new_[100911]_  = ~A169 & ~A170;
  assign \new_[100914]_  = A199 & A168;
  assign \new_[100915]_  = \new_[100914]_  & \new_[100911]_ ;
  assign \new_[100918]_  = A201 & ~A200;
  assign \new_[100921]_  = A265 & ~A203;
  assign \new_[100922]_  = \new_[100921]_  & \new_[100918]_ ;
  assign \new_[100923]_  = \new_[100922]_  & \new_[100915]_ ;
  assign \new_[100926]_  = ~A267 & ~A266;
  assign \new_[100929]_  = A269 & ~A268;
  assign \new_[100930]_  = \new_[100929]_  & \new_[100926]_ ;
  assign \new_[100933]_  = ~A299 & A298;
  assign \new_[100936]_  = A301 & A300;
  assign \new_[100937]_  = \new_[100936]_  & \new_[100933]_ ;
  assign \new_[100938]_  = \new_[100937]_  & \new_[100930]_ ;
  assign \new_[100941]_  = ~A169 & ~A170;
  assign \new_[100944]_  = A199 & A168;
  assign \new_[100945]_  = \new_[100944]_  & \new_[100941]_ ;
  assign \new_[100948]_  = A201 & ~A200;
  assign \new_[100951]_  = A265 & ~A203;
  assign \new_[100952]_  = \new_[100951]_  & \new_[100948]_ ;
  assign \new_[100953]_  = \new_[100952]_  & \new_[100945]_ ;
  assign \new_[100956]_  = ~A267 & ~A266;
  assign \new_[100959]_  = A269 & ~A268;
  assign \new_[100960]_  = \new_[100959]_  & \new_[100956]_ ;
  assign \new_[100963]_  = ~A299 & A298;
  assign \new_[100966]_  = ~A302 & A300;
  assign \new_[100967]_  = \new_[100966]_  & \new_[100963]_ ;
  assign \new_[100968]_  = \new_[100967]_  & \new_[100960]_ ;
  assign \new_[100971]_  = ~A169 & ~A170;
  assign \new_[100974]_  = A199 & A168;
  assign \new_[100975]_  = \new_[100974]_  & \new_[100971]_ ;
  assign \new_[100978]_  = A201 & ~A200;
  assign \new_[100981]_  = A265 & ~A203;
  assign \new_[100982]_  = \new_[100981]_  & \new_[100978]_ ;
  assign \new_[100983]_  = \new_[100982]_  & \new_[100975]_ ;
  assign \new_[100986]_  = ~A267 & ~A266;
  assign \new_[100989]_  = A269 & ~A268;
  assign \new_[100990]_  = \new_[100989]_  & \new_[100986]_ ;
  assign \new_[100993]_  = A299 & ~A298;
  assign \new_[100996]_  = A301 & A300;
  assign \new_[100997]_  = \new_[100996]_  & \new_[100993]_ ;
  assign \new_[100998]_  = \new_[100997]_  & \new_[100990]_ ;
  assign \new_[101001]_  = ~A169 & ~A170;
  assign \new_[101004]_  = A199 & A168;
  assign \new_[101005]_  = \new_[101004]_  & \new_[101001]_ ;
  assign \new_[101008]_  = A201 & ~A200;
  assign \new_[101011]_  = A265 & ~A203;
  assign \new_[101012]_  = \new_[101011]_  & \new_[101008]_ ;
  assign \new_[101013]_  = \new_[101012]_  & \new_[101005]_ ;
  assign \new_[101016]_  = ~A267 & ~A266;
  assign \new_[101019]_  = A269 & ~A268;
  assign \new_[101020]_  = \new_[101019]_  & \new_[101016]_ ;
  assign \new_[101023]_  = A299 & ~A298;
  assign \new_[101026]_  = ~A302 & A300;
  assign \new_[101027]_  = \new_[101026]_  & \new_[101023]_ ;
  assign \new_[101028]_  = \new_[101027]_  & \new_[101020]_ ;
  assign \new_[101031]_  = ~A169 & ~A170;
  assign \new_[101034]_  = A199 & A168;
  assign \new_[101035]_  = \new_[101034]_  & \new_[101031]_ ;
  assign \new_[101038]_  = ~A201 & ~A200;
  assign \new_[101041]_  = A203 & ~A202;
  assign \new_[101042]_  = \new_[101041]_  & \new_[101038]_ ;
  assign \new_[101043]_  = \new_[101042]_  & \new_[101035]_ ;
  assign \new_[101046]_  = A266 & ~A265;
  assign \new_[101049]_  = A268 & A267;
  assign \new_[101050]_  = \new_[101049]_  & \new_[101046]_ ;
  assign \new_[101053]_  = ~A299 & A298;
  assign \new_[101056]_  = A301 & A300;
  assign \new_[101057]_  = \new_[101056]_  & \new_[101053]_ ;
  assign \new_[101058]_  = \new_[101057]_  & \new_[101050]_ ;
  assign \new_[101061]_  = ~A169 & ~A170;
  assign \new_[101064]_  = A199 & A168;
  assign \new_[101065]_  = \new_[101064]_  & \new_[101061]_ ;
  assign \new_[101068]_  = ~A201 & ~A200;
  assign \new_[101071]_  = A203 & ~A202;
  assign \new_[101072]_  = \new_[101071]_  & \new_[101068]_ ;
  assign \new_[101073]_  = \new_[101072]_  & \new_[101065]_ ;
  assign \new_[101076]_  = A266 & ~A265;
  assign \new_[101079]_  = A268 & A267;
  assign \new_[101080]_  = \new_[101079]_  & \new_[101076]_ ;
  assign \new_[101083]_  = ~A299 & A298;
  assign \new_[101086]_  = ~A302 & A300;
  assign \new_[101087]_  = \new_[101086]_  & \new_[101083]_ ;
  assign \new_[101088]_  = \new_[101087]_  & \new_[101080]_ ;
  assign \new_[101091]_  = ~A169 & ~A170;
  assign \new_[101094]_  = A199 & A168;
  assign \new_[101095]_  = \new_[101094]_  & \new_[101091]_ ;
  assign \new_[101098]_  = ~A201 & ~A200;
  assign \new_[101101]_  = A203 & ~A202;
  assign \new_[101102]_  = \new_[101101]_  & \new_[101098]_ ;
  assign \new_[101103]_  = \new_[101102]_  & \new_[101095]_ ;
  assign \new_[101106]_  = A266 & ~A265;
  assign \new_[101109]_  = A268 & A267;
  assign \new_[101110]_  = \new_[101109]_  & \new_[101106]_ ;
  assign \new_[101113]_  = A299 & ~A298;
  assign \new_[101116]_  = A301 & A300;
  assign \new_[101117]_  = \new_[101116]_  & \new_[101113]_ ;
  assign \new_[101118]_  = \new_[101117]_  & \new_[101110]_ ;
  assign \new_[101121]_  = ~A169 & ~A170;
  assign \new_[101124]_  = A199 & A168;
  assign \new_[101125]_  = \new_[101124]_  & \new_[101121]_ ;
  assign \new_[101128]_  = ~A201 & ~A200;
  assign \new_[101131]_  = A203 & ~A202;
  assign \new_[101132]_  = \new_[101131]_  & \new_[101128]_ ;
  assign \new_[101133]_  = \new_[101132]_  & \new_[101125]_ ;
  assign \new_[101136]_  = A266 & ~A265;
  assign \new_[101139]_  = A268 & A267;
  assign \new_[101140]_  = \new_[101139]_  & \new_[101136]_ ;
  assign \new_[101143]_  = A299 & ~A298;
  assign \new_[101146]_  = ~A302 & A300;
  assign \new_[101147]_  = \new_[101146]_  & \new_[101143]_ ;
  assign \new_[101148]_  = \new_[101147]_  & \new_[101140]_ ;
  assign \new_[101151]_  = ~A169 & ~A170;
  assign \new_[101154]_  = A199 & A168;
  assign \new_[101155]_  = \new_[101154]_  & \new_[101151]_ ;
  assign \new_[101158]_  = ~A201 & ~A200;
  assign \new_[101161]_  = A203 & ~A202;
  assign \new_[101162]_  = \new_[101161]_  & \new_[101158]_ ;
  assign \new_[101163]_  = \new_[101162]_  & \new_[101155]_ ;
  assign \new_[101166]_  = A266 & ~A265;
  assign \new_[101169]_  = ~A269 & A267;
  assign \new_[101170]_  = \new_[101169]_  & \new_[101166]_ ;
  assign \new_[101173]_  = ~A299 & A298;
  assign \new_[101176]_  = A301 & A300;
  assign \new_[101177]_  = \new_[101176]_  & \new_[101173]_ ;
  assign \new_[101178]_  = \new_[101177]_  & \new_[101170]_ ;
  assign \new_[101181]_  = ~A169 & ~A170;
  assign \new_[101184]_  = A199 & A168;
  assign \new_[101185]_  = \new_[101184]_  & \new_[101181]_ ;
  assign \new_[101188]_  = ~A201 & ~A200;
  assign \new_[101191]_  = A203 & ~A202;
  assign \new_[101192]_  = \new_[101191]_  & \new_[101188]_ ;
  assign \new_[101193]_  = \new_[101192]_  & \new_[101185]_ ;
  assign \new_[101196]_  = A266 & ~A265;
  assign \new_[101199]_  = ~A269 & A267;
  assign \new_[101200]_  = \new_[101199]_  & \new_[101196]_ ;
  assign \new_[101203]_  = ~A299 & A298;
  assign \new_[101206]_  = ~A302 & A300;
  assign \new_[101207]_  = \new_[101206]_  & \new_[101203]_ ;
  assign \new_[101208]_  = \new_[101207]_  & \new_[101200]_ ;
  assign \new_[101211]_  = ~A169 & ~A170;
  assign \new_[101214]_  = A199 & A168;
  assign \new_[101215]_  = \new_[101214]_  & \new_[101211]_ ;
  assign \new_[101218]_  = ~A201 & ~A200;
  assign \new_[101221]_  = A203 & ~A202;
  assign \new_[101222]_  = \new_[101221]_  & \new_[101218]_ ;
  assign \new_[101223]_  = \new_[101222]_  & \new_[101215]_ ;
  assign \new_[101226]_  = A266 & ~A265;
  assign \new_[101229]_  = ~A269 & A267;
  assign \new_[101230]_  = \new_[101229]_  & \new_[101226]_ ;
  assign \new_[101233]_  = A299 & ~A298;
  assign \new_[101236]_  = A301 & A300;
  assign \new_[101237]_  = \new_[101236]_  & \new_[101233]_ ;
  assign \new_[101238]_  = \new_[101237]_  & \new_[101230]_ ;
  assign \new_[101241]_  = ~A169 & ~A170;
  assign \new_[101244]_  = A199 & A168;
  assign \new_[101245]_  = \new_[101244]_  & \new_[101241]_ ;
  assign \new_[101248]_  = ~A201 & ~A200;
  assign \new_[101251]_  = A203 & ~A202;
  assign \new_[101252]_  = \new_[101251]_  & \new_[101248]_ ;
  assign \new_[101253]_  = \new_[101252]_  & \new_[101245]_ ;
  assign \new_[101256]_  = A266 & ~A265;
  assign \new_[101259]_  = ~A269 & A267;
  assign \new_[101260]_  = \new_[101259]_  & \new_[101256]_ ;
  assign \new_[101263]_  = A299 & ~A298;
  assign \new_[101266]_  = ~A302 & A300;
  assign \new_[101267]_  = \new_[101266]_  & \new_[101263]_ ;
  assign \new_[101268]_  = \new_[101267]_  & \new_[101260]_ ;
  assign \new_[101271]_  = ~A169 & ~A170;
  assign \new_[101274]_  = A199 & A168;
  assign \new_[101275]_  = \new_[101274]_  & \new_[101271]_ ;
  assign \new_[101278]_  = ~A201 & ~A200;
  assign \new_[101281]_  = A203 & ~A202;
  assign \new_[101282]_  = \new_[101281]_  & \new_[101278]_ ;
  assign \new_[101283]_  = \new_[101282]_  & \new_[101275]_ ;
  assign \new_[101286]_  = ~A266 & A265;
  assign \new_[101289]_  = A268 & A267;
  assign \new_[101290]_  = \new_[101289]_  & \new_[101286]_ ;
  assign \new_[101293]_  = ~A299 & A298;
  assign \new_[101296]_  = A301 & A300;
  assign \new_[101297]_  = \new_[101296]_  & \new_[101293]_ ;
  assign \new_[101298]_  = \new_[101297]_  & \new_[101290]_ ;
  assign \new_[101301]_  = ~A169 & ~A170;
  assign \new_[101304]_  = A199 & A168;
  assign \new_[101305]_  = \new_[101304]_  & \new_[101301]_ ;
  assign \new_[101308]_  = ~A201 & ~A200;
  assign \new_[101311]_  = A203 & ~A202;
  assign \new_[101312]_  = \new_[101311]_  & \new_[101308]_ ;
  assign \new_[101313]_  = \new_[101312]_  & \new_[101305]_ ;
  assign \new_[101316]_  = ~A266 & A265;
  assign \new_[101319]_  = A268 & A267;
  assign \new_[101320]_  = \new_[101319]_  & \new_[101316]_ ;
  assign \new_[101323]_  = ~A299 & A298;
  assign \new_[101326]_  = ~A302 & A300;
  assign \new_[101327]_  = \new_[101326]_  & \new_[101323]_ ;
  assign \new_[101328]_  = \new_[101327]_  & \new_[101320]_ ;
  assign \new_[101331]_  = ~A169 & ~A170;
  assign \new_[101334]_  = A199 & A168;
  assign \new_[101335]_  = \new_[101334]_  & \new_[101331]_ ;
  assign \new_[101338]_  = ~A201 & ~A200;
  assign \new_[101341]_  = A203 & ~A202;
  assign \new_[101342]_  = \new_[101341]_  & \new_[101338]_ ;
  assign \new_[101343]_  = \new_[101342]_  & \new_[101335]_ ;
  assign \new_[101346]_  = ~A266 & A265;
  assign \new_[101349]_  = A268 & A267;
  assign \new_[101350]_  = \new_[101349]_  & \new_[101346]_ ;
  assign \new_[101353]_  = A299 & ~A298;
  assign \new_[101356]_  = A301 & A300;
  assign \new_[101357]_  = \new_[101356]_  & \new_[101353]_ ;
  assign \new_[101358]_  = \new_[101357]_  & \new_[101350]_ ;
  assign \new_[101361]_  = ~A169 & ~A170;
  assign \new_[101364]_  = A199 & A168;
  assign \new_[101365]_  = \new_[101364]_  & \new_[101361]_ ;
  assign \new_[101368]_  = ~A201 & ~A200;
  assign \new_[101371]_  = A203 & ~A202;
  assign \new_[101372]_  = \new_[101371]_  & \new_[101368]_ ;
  assign \new_[101373]_  = \new_[101372]_  & \new_[101365]_ ;
  assign \new_[101376]_  = ~A266 & A265;
  assign \new_[101379]_  = A268 & A267;
  assign \new_[101380]_  = \new_[101379]_  & \new_[101376]_ ;
  assign \new_[101383]_  = A299 & ~A298;
  assign \new_[101386]_  = ~A302 & A300;
  assign \new_[101387]_  = \new_[101386]_  & \new_[101383]_ ;
  assign \new_[101388]_  = \new_[101387]_  & \new_[101380]_ ;
  assign \new_[101391]_  = ~A169 & ~A170;
  assign \new_[101394]_  = A199 & A168;
  assign \new_[101395]_  = \new_[101394]_  & \new_[101391]_ ;
  assign \new_[101398]_  = ~A201 & ~A200;
  assign \new_[101401]_  = A203 & ~A202;
  assign \new_[101402]_  = \new_[101401]_  & \new_[101398]_ ;
  assign \new_[101403]_  = \new_[101402]_  & \new_[101395]_ ;
  assign \new_[101406]_  = ~A266 & A265;
  assign \new_[101409]_  = ~A269 & A267;
  assign \new_[101410]_  = \new_[101409]_  & \new_[101406]_ ;
  assign \new_[101413]_  = ~A299 & A298;
  assign \new_[101416]_  = A301 & A300;
  assign \new_[101417]_  = \new_[101416]_  & \new_[101413]_ ;
  assign \new_[101418]_  = \new_[101417]_  & \new_[101410]_ ;
  assign \new_[101421]_  = ~A169 & ~A170;
  assign \new_[101424]_  = A199 & A168;
  assign \new_[101425]_  = \new_[101424]_  & \new_[101421]_ ;
  assign \new_[101428]_  = ~A201 & ~A200;
  assign \new_[101431]_  = A203 & ~A202;
  assign \new_[101432]_  = \new_[101431]_  & \new_[101428]_ ;
  assign \new_[101433]_  = \new_[101432]_  & \new_[101425]_ ;
  assign \new_[101436]_  = ~A266 & A265;
  assign \new_[101439]_  = ~A269 & A267;
  assign \new_[101440]_  = \new_[101439]_  & \new_[101436]_ ;
  assign \new_[101443]_  = ~A299 & A298;
  assign \new_[101446]_  = ~A302 & A300;
  assign \new_[101447]_  = \new_[101446]_  & \new_[101443]_ ;
  assign \new_[101448]_  = \new_[101447]_  & \new_[101440]_ ;
  assign \new_[101451]_  = ~A169 & ~A170;
  assign \new_[101454]_  = A199 & A168;
  assign \new_[101455]_  = \new_[101454]_  & \new_[101451]_ ;
  assign \new_[101458]_  = ~A201 & ~A200;
  assign \new_[101461]_  = A203 & ~A202;
  assign \new_[101462]_  = \new_[101461]_  & \new_[101458]_ ;
  assign \new_[101463]_  = \new_[101462]_  & \new_[101455]_ ;
  assign \new_[101466]_  = ~A266 & A265;
  assign \new_[101469]_  = ~A269 & A267;
  assign \new_[101470]_  = \new_[101469]_  & \new_[101466]_ ;
  assign \new_[101473]_  = A299 & ~A298;
  assign \new_[101476]_  = A301 & A300;
  assign \new_[101477]_  = \new_[101476]_  & \new_[101473]_ ;
  assign \new_[101478]_  = \new_[101477]_  & \new_[101470]_ ;
  assign \new_[101481]_  = ~A169 & ~A170;
  assign \new_[101484]_  = A199 & A168;
  assign \new_[101485]_  = \new_[101484]_  & \new_[101481]_ ;
  assign \new_[101488]_  = ~A201 & ~A200;
  assign \new_[101491]_  = A203 & ~A202;
  assign \new_[101492]_  = \new_[101491]_  & \new_[101488]_ ;
  assign \new_[101493]_  = \new_[101492]_  & \new_[101485]_ ;
  assign \new_[101496]_  = ~A266 & A265;
  assign \new_[101499]_  = ~A269 & A267;
  assign \new_[101500]_  = \new_[101499]_  & \new_[101496]_ ;
  assign \new_[101503]_  = A299 & ~A298;
  assign \new_[101506]_  = ~A302 & A300;
  assign \new_[101507]_  = \new_[101506]_  & \new_[101503]_ ;
  assign \new_[101508]_  = \new_[101507]_  & \new_[101500]_ ;
  assign \new_[101511]_  = ~A169 & ~A170;
  assign \new_[101514]_  = A167 & ~A168;
  assign \new_[101515]_  = \new_[101514]_  & \new_[101511]_ ;
  assign \new_[101518]_  = A201 & ~A166;
  assign \new_[101521]_  = A203 & ~A202;
  assign \new_[101522]_  = \new_[101521]_  & \new_[101518]_ ;
  assign \new_[101523]_  = \new_[101522]_  & \new_[101515]_ ;
  assign \new_[101526]_  = ~A268 & A267;
  assign \new_[101529]_  = A298 & A269;
  assign \new_[101530]_  = \new_[101529]_  & \new_[101526]_ ;
  assign \new_[101533]_  = ~A300 & ~A299;
  assign \new_[101536]_  = A302 & ~A301;
  assign \new_[101537]_  = \new_[101536]_  & \new_[101533]_ ;
  assign \new_[101538]_  = \new_[101537]_  & \new_[101530]_ ;
  assign \new_[101541]_  = ~A169 & ~A170;
  assign \new_[101544]_  = A167 & ~A168;
  assign \new_[101545]_  = \new_[101544]_  & \new_[101541]_ ;
  assign \new_[101548]_  = A201 & ~A166;
  assign \new_[101551]_  = A203 & ~A202;
  assign \new_[101552]_  = \new_[101551]_  & \new_[101548]_ ;
  assign \new_[101553]_  = \new_[101552]_  & \new_[101545]_ ;
  assign \new_[101556]_  = ~A268 & A267;
  assign \new_[101559]_  = ~A298 & A269;
  assign \new_[101560]_  = \new_[101559]_  & \new_[101556]_ ;
  assign \new_[101563]_  = ~A300 & A299;
  assign \new_[101566]_  = A302 & ~A301;
  assign \new_[101567]_  = \new_[101566]_  & \new_[101563]_ ;
  assign \new_[101568]_  = \new_[101567]_  & \new_[101560]_ ;
  assign \new_[101571]_  = ~A169 & ~A170;
  assign \new_[101574]_  = A167 & ~A168;
  assign \new_[101575]_  = \new_[101574]_  & \new_[101571]_ ;
  assign \new_[101578]_  = A201 & ~A166;
  assign \new_[101581]_  = A203 & ~A202;
  assign \new_[101582]_  = \new_[101581]_  & \new_[101578]_ ;
  assign \new_[101583]_  = \new_[101582]_  & \new_[101575]_ ;
  assign \new_[101586]_  = A266 & ~A265;
  assign \new_[101589]_  = ~A268 & ~A267;
  assign \new_[101590]_  = \new_[101589]_  & \new_[101586]_ ;
  assign \new_[101593]_  = A300 & A269;
  assign \new_[101596]_  = A302 & ~A301;
  assign \new_[101597]_  = \new_[101596]_  & \new_[101593]_ ;
  assign \new_[101598]_  = \new_[101597]_  & \new_[101590]_ ;
  assign \new_[101601]_  = ~A169 & ~A170;
  assign \new_[101604]_  = A167 & ~A168;
  assign \new_[101605]_  = \new_[101604]_  & \new_[101601]_ ;
  assign \new_[101608]_  = A201 & ~A166;
  assign \new_[101611]_  = A203 & ~A202;
  assign \new_[101612]_  = \new_[101611]_  & \new_[101608]_ ;
  assign \new_[101613]_  = \new_[101612]_  & \new_[101605]_ ;
  assign \new_[101616]_  = ~A266 & A265;
  assign \new_[101619]_  = ~A268 & ~A267;
  assign \new_[101620]_  = \new_[101619]_  & \new_[101616]_ ;
  assign \new_[101623]_  = A300 & A269;
  assign \new_[101626]_  = A302 & ~A301;
  assign \new_[101627]_  = \new_[101626]_  & \new_[101623]_ ;
  assign \new_[101628]_  = \new_[101627]_  & \new_[101620]_ ;
  assign \new_[101631]_  = ~A169 & ~A170;
  assign \new_[101634]_  = ~A167 & ~A168;
  assign \new_[101635]_  = \new_[101634]_  & \new_[101631]_ ;
  assign \new_[101638]_  = A201 & A166;
  assign \new_[101641]_  = A203 & ~A202;
  assign \new_[101642]_  = \new_[101641]_  & \new_[101638]_ ;
  assign \new_[101643]_  = \new_[101642]_  & \new_[101635]_ ;
  assign \new_[101646]_  = ~A268 & A267;
  assign \new_[101649]_  = A298 & A269;
  assign \new_[101650]_  = \new_[101649]_  & \new_[101646]_ ;
  assign \new_[101653]_  = ~A300 & ~A299;
  assign \new_[101656]_  = A302 & ~A301;
  assign \new_[101657]_  = \new_[101656]_  & \new_[101653]_ ;
  assign \new_[101658]_  = \new_[101657]_  & \new_[101650]_ ;
  assign \new_[101661]_  = ~A169 & ~A170;
  assign \new_[101664]_  = ~A167 & ~A168;
  assign \new_[101665]_  = \new_[101664]_  & \new_[101661]_ ;
  assign \new_[101668]_  = A201 & A166;
  assign \new_[101671]_  = A203 & ~A202;
  assign \new_[101672]_  = \new_[101671]_  & \new_[101668]_ ;
  assign \new_[101673]_  = \new_[101672]_  & \new_[101665]_ ;
  assign \new_[101676]_  = ~A268 & A267;
  assign \new_[101679]_  = ~A298 & A269;
  assign \new_[101680]_  = \new_[101679]_  & \new_[101676]_ ;
  assign \new_[101683]_  = ~A300 & A299;
  assign \new_[101686]_  = A302 & ~A301;
  assign \new_[101687]_  = \new_[101686]_  & \new_[101683]_ ;
  assign \new_[101688]_  = \new_[101687]_  & \new_[101680]_ ;
  assign \new_[101691]_  = ~A169 & ~A170;
  assign \new_[101694]_  = ~A167 & ~A168;
  assign \new_[101695]_  = \new_[101694]_  & \new_[101691]_ ;
  assign \new_[101698]_  = A201 & A166;
  assign \new_[101701]_  = A203 & ~A202;
  assign \new_[101702]_  = \new_[101701]_  & \new_[101698]_ ;
  assign \new_[101703]_  = \new_[101702]_  & \new_[101695]_ ;
  assign \new_[101706]_  = A266 & ~A265;
  assign \new_[101709]_  = ~A268 & ~A267;
  assign \new_[101710]_  = \new_[101709]_  & \new_[101706]_ ;
  assign \new_[101713]_  = A300 & A269;
  assign \new_[101716]_  = A302 & ~A301;
  assign \new_[101717]_  = \new_[101716]_  & \new_[101713]_ ;
  assign \new_[101718]_  = \new_[101717]_  & \new_[101710]_ ;
  assign \new_[101721]_  = ~A169 & ~A170;
  assign \new_[101724]_  = ~A167 & ~A168;
  assign \new_[101725]_  = \new_[101724]_  & \new_[101721]_ ;
  assign \new_[101728]_  = A201 & A166;
  assign \new_[101731]_  = A203 & ~A202;
  assign \new_[101732]_  = \new_[101731]_  & \new_[101728]_ ;
  assign \new_[101733]_  = \new_[101732]_  & \new_[101725]_ ;
  assign \new_[101736]_  = ~A266 & A265;
  assign \new_[101739]_  = ~A268 & ~A267;
  assign \new_[101740]_  = \new_[101739]_  & \new_[101736]_ ;
  assign \new_[101743]_  = A300 & A269;
  assign \new_[101746]_  = A302 & ~A301;
  assign \new_[101747]_  = \new_[101746]_  & \new_[101743]_ ;
  assign \new_[101748]_  = \new_[101747]_  & \new_[101740]_ ;
  assign \new_[101751]_  = A166 & A167;
  assign \new_[101754]_  = A200 & ~A199;
  assign \new_[101755]_  = \new_[101754]_  & \new_[101751]_ ;
  assign \new_[101758]_  = ~A202 & ~A201;
  assign \new_[101761]_  = ~A265 & A203;
  assign \new_[101762]_  = \new_[101761]_  & \new_[101758]_ ;
  assign \new_[101763]_  = \new_[101762]_  & \new_[101755]_ ;
  assign \new_[101766]_  = ~A267 & A266;
  assign \new_[101769]_  = A269 & ~A268;
  assign \new_[101770]_  = \new_[101769]_  & \new_[101766]_ ;
  assign \new_[101773]_  = ~A299 & A298;
  assign \new_[101777]_  = A302 & ~A301;
  assign \new_[101778]_  = ~A300 & \new_[101777]_ ;
  assign \new_[101779]_  = \new_[101778]_  & \new_[101773]_ ;
  assign \new_[101780]_  = \new_[101779]_  & \new_[101770]_ ;
  assign \new_[101783]_  = A166 & A167;
  assign \new_[101786]_  = A200 & ~A199;
  assign \new_[101787]_  = \new_[101786]_  & \new_[101783]_ ;
  assign \new_[101790]_  = ~A202 & ~A201;
  assign \new_[101793]_  = ~A265 & A203;
  assign \new_[101794]_  = \new_[101793]_  & \new_[101790]_ ;
  assign \new_[101795]_  = \new_[101794]_  & \new_[101787]_ ;
  assign \new_[101798]_  = ~A267 & A266;
  assign \new_[101801]_  = A269 & ~A268;
  assign \new_[101802]_  = \new_[101801]_  & \new_[101798]_ ;
  assign \new_[101805]_  = A299 & ~A298;
  assign \new_[101809]_  = A302 & ~A301;
  assign \new_[101810]_  = ~A300 & \new_[101809]_ ;
  assign \new_[101811]_  = \new_[101810]_  & \new_[101805]_ ;
  assign \new_[101812]_  = \new_[101811]_  & \new_[101802]_ ;
  assign \new_[101815]_  = A166 & A167;
  assign \new_[101818]_  = A200 & ~A199;
  assign \new_[101819]_  = \new_[101818]_  & \new_[101815]_ ;
  assign \new_[101822]_  = ~A202 & ~A201;
  assign \new_[101825]_  = A265 & A203;
  assign \new_[101826]_  = \new_[101825]_  & \new_[101822]_ ;
  assign \new_[101827]_  = \new_[101826]_  & \new_[101819]_ ;
  assign \new_[101830]_  = ~A267 & ~A266;
  assign \new_[101833]_  = A269 & ~A268;
  assign \new_[101834]_  = \new_[101833]_  & \new_[101830]_ ;
  assign \new_[101837]_  = ~A299 & A298;
  assign \new_[101841]_  = A302 & ~A301;
  assign \new_[101842]_  = ~A300 & \new_[101841]_ ;
  assign \new_[101843]_  = \new_[101842]_  & \new_[101837]_ ;
  assign \new_[101844]_  = \new_[101843]_  & \new_[101834]_ ;
  assign \new_[101847]_  = A166 & A167;
  assign \new_[101850]_  = A200 & ~A199;
  assign \new_[101851]_  = \new_[101850]_  & \new_[101847]_ ;
  assign \new_[101854]_  = ~A202 & ~A201;
  assign \new_[101857]_  = A265 & A203;
  assign \new_[101858]_  = \new_[101857]_  & \new_[101854]_ ;
  assign \new_[101859]_  = \new_[101858]_  & \new_[101851]_ ;
  assign \new_[101862]_  = ~A267 & ~A266;
  assign \new_[101865]_  = A269 & ~A268;
  assign \new_[101866]_  = \new_[101865]_  & \new_[101862]_ ;
  assign \new_[101869]_  = A299 & ~A298;
  assign \new_[101873]_  = A302 & ~A301;
  assign \new_[101874]_  = ~A300 & \new_[101873]_ ;
  assign \new_[101875]_  = \new_[101874]_  & \new_[101869]_ ;
  assign \new_[101876]_  = \new_[101875]_  & \new_[101866]_ ;
  assign \new_[101879]_  = A166 & A167;
  assign \new_[101882]_  = ~A200 & A199;
  assign \new_[101883]_  = \new_[101882]_  & \new_[101879]_ ;
  assign \new_[101886]_  = ~A202 & ~A201;
  assign \new_[101889]_  = ~A265 & A203;
  assign \new_[101890]_  = \new_[101889]_  & \new_[101886]_ ;
  assign \new_[101891]_  = \new_[101890]_  & \new_[101883]_ ;
  assign \new_[101894]_  = ~A267 & A266;
  assign \new_[101897]_  = A269 & ~A268;
  assign \new_[101898]_  = \new_[101897]_  & \new_[101894]_ ;
  assign \new_[101901]_  = ~A299 & A298;
  assign \new_[101905]_  = A302 & ~A301;
  assign \new_[101906]_  = ~A300 & \new_[101905]_ ;
  assign \new_[101907]_  = \new_[101906]_  & \new_[101901]_ ;
  assign \new_[101908]_  = \new_[101907]_  & \new_[101898]_ ;
  assign \new_[101911]_  = A166 & A167;
  assign \new_[101914]_  = ~A200 & A199;
  assign \new_[101915]_  = \new_[101914]_  & \new_[101911]_ ;
  assign \new_[101918]_  = ~A202 & ~A201;
  assign \new_[101921]_  = ~A265 & A203;
  assign \new_[101922]_  = \new_[101921]_  & \new_[101918]_ ;
  assign \new_[101923]_  = \new_[101922]_  & \new_[101915]_ ;
  assign \new_[101926]_  = ~A267 & A266;
  assign \new_[101929]_  = A269 & ~A268;
  assign \new_[101930]_  = \new_[101929]_  & \new_[101926]_ ;
  assign \new_[101933]_  = A299 & ~A298;
  assign \new_[101937]_  = A302 & ~A301;
  assign \new_[101938]_  = ~A300 & \new_[101937]_ ;
  assign \new_[101939]_  = \new_[101938]_  & \new_[101933]_ ;
  assign \new_[101940]_  = \new_[101939]_  & \new_[101930]_ ;
  assign \new_[101943]_  = A166 & A167;
  assign \new_[101946]_  = ~A200 & A199;
  assign \new_[101947]_  = \new_[101946]_  & \new_[101943]_ ;
  assign \new_[101950]_  = ~A202 & ~A201;
  assign \new_[101953]_  = A265 & A203;
  assign \new_[101954]_  = \new_[101953]_  & \new_[101950]_ ;
  assign \new_[101955]_  = \new_[101954]_  & \new_[101947]_ ;
  assign \new_[101958]_  = ~A267 & ~A266;
  assign \new_[101961]_  = A269 & ~A268;
  assign \new_[101962]_  = \new_[101961]_  & \new_[101958]_ ;
  assign \new_[101965]_  = ~A299 & A298;
  assign \new_[101969]_  = A302 & ~A301;
  assign \new_[101970]_  = ~A300 & \new_[101969]_ ;
  assign \new_[101971]_  = \new_[101970]_  & \new_[101965]_ ;
  assign \new_[101972]_  = \new_[101971]_  & \new_[101962]_ ;
  assign \new_[101975]_  = A166 & A167;
  assign \new_[101978]_  = ~A200 & A199;
  assign \new_[101979]_  = \new_[101978]_  & \new_[101975]_ ;
  assign \new_[101982]_  = ~A202 & ~A201;
  assign \new_[101985]_  = A265 & A203;
  assign \new_[101986]_  = \new_[101985]_  & \new_[101982]_ ;
  assign \new_[101987]_  = \new_[101986]_  & \new_[101979]_ ;
  assign \new_[101990]_  = ~A267 & ~A266;
  assign \new_[101993]_  = A269 & ~A268;
  assign \new_[101994]_  = \new_[101993]_  & \new_[101990]_ ;
  assign \new_[101997]_  = A299 & ~A298;
  assign \new_[102001]_  = A302 & ~A301;
  assign \new_[102002]_  = ~A300 & \new_[102001]_ ;
  assign \new_[102003]_  = \new_[102002]_  & \new_[101997]_ ;
  assign \new_[102004]_  = \new_[102003]_  & \new_[101994]_ ;
  assign \new_[102007]_  = ~A166 & ~A167;
  assign \new_[102010]_  = A200 & ~A199;
  assign \new_[102011]_  = \new_[102010]_  & \new_[102007]_ ;
  assign \new_[102014]_  = ~A202 & ~A201;
  assign \new_[102017]_  = ~A265 & A203;
  assign \new_[102018]_  = \new_[102017]_  & \new_[102014]_ ;
  assign \new_[102019]_  = \new_[102018]_  & \new_[102011]_ ;
  assign \new_[102022]_  = ~A267 & A266;
  assign \new_[102025]_  = A269 & ~A268;
  assign \new_[102026]_  = \new_[102025]_  & \new_[102022]_ ;
  assign \new_[102029]_  = ~A299 & A298;
  assign \new_[102033]_  = A302 & ~A301;
  assign \new_[102034]_  = ~A300 & \new_[102033]_ ;
  assign \new_[102035]_  = \new_[102034]_  & \new_[102029]_ ;
  assign \new_[102036]_  = \new_[102035]_  & \new_[102026]_ ;
  assign \new_[102039]_  = ~A166 & ~A167;
  assign \new_[102042]_  = A200 & ~A199;
  assign \new_[102043]_  = \new_[102042]_  & \new_[102039]_ ;
  assign \new_[102046]_  = ~A202 & ~A201;
  assign \new_[102049]_  = ~A265 & A203;
  assign \new_[102050]_  = \new_[102049]_  & \new_[102046]_ ;
  assign \new_[102051]_  = \new_[102050]_  & \new_[102043]_ ;
  assign \new_[102054]_  = ~A267 & A266;
  assign \new_[102057]_  = A269 & ~A268;
  assign \new_[102058]_  = \new_[102057]_  & \new_[102054]_ ;
  assign \new_[102061]_  = A299 & ~A298;
  assign \new_[102065]_  = A302 & ~A301;
  assign \new_[102066]_  = ~A300 & \new_[102065]_ ;
  assign \new_[102067]_  = \new_[102066]_  & \new_[102061]_ ;
  assign \new_[102068]_  = \new_[102067]_  & \new_[102058]_ ;
  assign \new_[102071]_  = ~A166 & ~A167;
  assign \new_[102074]_  = A200 & ~A199;
  assign \new_[102075]_  = \new_[102074]_  & \new_[102071]_ ;
  assign \new_[102078]_  = ~A202 & ~A201;
  assign \new_[102081]_  = A265 & A203;
  assign \new_[102082]_  = \new_[102081]_  & \new_[102078]_ ;
  assign \new_[102083]_  = \new_[102082]_  & \new_[102075]_ ;
  assign \new_[102086]_  = ~A267 & ~A266;
  assign \new_[102089]_  = A269 & ~A268;
  assign \new_[102090]_  = \new_[102089]_  & \new_[102086]_ ;
  assign \new_[102093]_  = ~A299 & A298;
  assign \new_[102097]_  = A302 & ~A301;
  assign \new_[102098]_  = ~A300 & \new_[102097]_ ;
  assign \new_[102099]_  = \new_[102098]_  & \new_[102093]_ ;
  assign \new_[102100]_  = \new_[102099]_  & \new_[102090]_ ;
  assign \new_[102103]_  = ~A166 & ~A167;
  assign \new_[102106]_  = A200 & ~A199;
  assign \new_[102107]_  = \new_[102106]_  & \new_[102103]_ ;
  assign \new_[102110]_  = ~A202 & ~A201;
  assign \new_[102113]_  = A265 & A203;
  assign \new_[102114]_  = \new_[102113]_  & \new_[102110]_ ;
  assign \new_[102115]_  = \new_[102114]_  & \new_[102107]_ ;
  assign \new_[102118]_  = ~A267 & ~A266;
  assign \new_[102121]_  = A269 & ~A268;
  assign \new_[102122]_  = \new_[102121]_  & \new_[102118]_ ;
  assign \new_[102125]_  = A299 & ~A298;
  assign \new_[102129]_  = A302 & ~A301;
  assign \new_[102130]_  = ~A300 & \new_[102129]_ ;
  assign \new_[102131]_  = \new_[102130]_  & \new_[102125]_ ;
  assign \new_[102132]_  = \new_[102131]_  & \new_[102122]_ ;
  assign \new_[102135]_  = ~A166 & ~A167;
  assign \new_[102138]_  = ~A200 & A199;
  assign \new_[102139]_  = \new_[102138]_  & \new_[102135]_ ;
  assign \new_[102142]_  = ~A202 & ~A201;
  assign \new_[102145]_  = ~A265 & A203;
  assign \new_[102146]_  = \new_[102145]_  & \new_[102142]_ ;
  assign \new_[102147]_  = \new_[102146]_  & \new_[102139]_ ;
  assign \new_[102150]_  = ~A267 & A266;
  assign \new_[102153]_  = A269 & ~A268;
  assign \new_[102154]_  = \new_[102153]_  & \new_[102150]_ ;
  assign \new_[102157]_  = ~A299 & A298;
  assign \new_[102161]_  = A302 & ~A301;
  assign \new_[102162]_  = ~A300 & \new_[102161]_ ;
  assign \new_[102163]_  = \new_[102162]_  & \new_[102157]_ ;
  assign \new_[102164]_  = \new_[102163]_  & \new_[102154]_ ;
  assign \new_[102167]_  = ~A166 & ~A167;
  assign \new_[102170]_  = ~A200 & A199;
  assign \new_[102171]_  = \new_[102170]_  & \new_[102167]_ ;
  assign \new_[102174]_  = ~A202 & ~A201;
  assign \new_[102177]_  = ~A265 & A203;
  assign \new_[102178]_  = \new_[102177]_  & \new_[102174]_ ;
  assign \new_[102179]_  = \new_[102178]_  & \new_[102171]_ ;
  assign \new_[102182]_  = ~A267 & A266;
  assign \new_[102185]_  = A269 & ~A268;
  assign \new_[102186]_  = \new_[102185]_  & \new_[102182]_ ;
  assign \new_[102189]_  = A299 & ~A298;
  assign \new_[102193]_  = A302 & ~A301;
  assign \new_[102194]_  = ~A300 & \new_[102193]_ ;
  assign \new_[102195]_  = \new_[102194]_  & \new_[102189]_ ;
  assign \new_[102196]_  = \new_[102195]_  & \new_[102186]_ ;
  assign \new_[102199]_  = ~A166 & ~A167;
  assign \new_[102202]_  = ~A200 & A199;
  assign \new_[102203]_  = \new_[102202]_  & \new_[102199]_ ;
  assign \new_[102206]_  = ~A202 & ~A201;
  assign \new_[102209]_  = A265 & A203;
  assign \new_[102210]_  = \new_[102209]_  & \new_[102206]_ ;
  assign \new_[102211]_  = \new_[102210]_  & \new_[102203]_ ;
  assign \new_[102214]_  = ~A267 & ~A266;
  assign \new_[102217]_  = A269 & ~A268;
  assign \new_[102218]_  = \new_[102217]_  & \new_[102214]_ ;
  assign \new_[102221]_  = ~A299 & A298;
  assign \new_[102225]_  = A302 & ~A301;
  assign \new_[102226]_  = ~A300 & \new_[102225]_ ;
  assign \new_[102227]_  = \new_[102226]_  & \new_[102221]_ ;
  assign \new_[102228]_  = \new_[102227]_  & \new_[102218]_ ;
  assign \new_[102231]_  = ~A166 & ~A167;
  assign \new_[102234]_  = ~A200 & A199;
  assign \new_[102235]_  = \new_[102234]_  & \new_[102231]_ ;
  assign \new_[102238]_  = ~A202 & ~A201;
  assign \new_[102241]_  = A265 & A203;
  assign \new_[102242]_  = \new_[102241]_  & \new_[102238]_ ;
  assign \new_[102243]_  = \new_[102242]_  & \new_[102235]_ ;
  assign \new_[102246]_  = ~A267 & ~A266;
  assign \new_[102249]_  = A269 & ~A268;
  assign \new_[102250]_  = \new_[102249]_  & \new_[102246]_ ;
  assign \new_[102253]_  = A299 & ~A298;
  assign \new_[102257]_  = A302 & ~A301;
  assign \new_[102258]_  = ~A300 & \new_[102257]_ ;
  assign \new_[102259]_  = \new_[102258]_  & \new_[102253]_ ;
  assign \new_[102260]_  = \new_[102259]_  & \new_[102250]_ ;
  assign \new_[102263]_  = ~A168 & A170;
  assign \new_[102266]_  = A200 & ~A199;
  assign \new_[102267]_  = \new_[102266]_  & \new_[102263]_ ;
  assign \new_[102270]_  = ~A202 & ~A201;
  assign \new_[102273]_  = ~A265 & A203;
  assign \new_[102274]_  = \new_[102273]_  & \new_[102270]_ ;
  assign \new_[102275]_  = \new_[102274]_  & \new_[102267]_ ;
  assign \new_[102278]_  = ~A267 & A266;
  assign \new_[102281]_  = A269 & ~A268;
  assign \new_[102282]_  = \new_[102281]_  & \new_[102278]_ ;
  assign \new_[102285]_  = ~A299 & A298;
  assign \new_[102289]_  = A302 & ~A301;
  assign \new_[102290]_  = ~A300 & \new_[102289]_ ;
  assign \new_[102291]_  = \new_[102290]_  & \new_[102285]_ ;
  assign \new_[102292]_  = \new_[102291]_  & \new_[102282]_ ;
  assign \new_[102295]_  = ~A168 & A170;
  assign \new_[102298]_  = A200 & ~A199;
  assign \new_[102299]_  = \new_[102298]_  & \new_[102295]_ ;
  assign \new_[102302]_  = ~A202 & ~A201;
  assign \new_[102305]_  = ~A265 & A203;
  assign \new_[102306]_  = \new_[102305]_  & \new_[102302]_ ;
  assign \new_[102307]_  = \new_[102306]_  & \new_[102299]_ ;
  assign \new_[102310]_  = ~A267 & A266;
  assign \new_[102313]_  = A269 & ~A268;
  assign \new_[102314]_  = \new_[102313]_  & \new_[102310]_ ;
  assign \new_[102317]_  = A299 & ~A298;
  assign \new_[102321]_  = A302 & ~A301;
  assign \new_[102322]_  = ~A300 & \new_[102321]_ ;
  assign \new_[102323]_  = \new_[102322]_  & \new_[102317]_ ;
  assign \new_[102324]_  = \new_[102323]_  & \new_[102314]_ ;
  assign \new_[102327]_  = ~A168 & A170;
  assign \new_[102330]_  = A200 & ~A199;
  assign \new_[102331]_  = \new_[102330]_  & \new_[102327]_ ;
  assign \new_[102334]_  = ~A202 & ~A201;
  assign \new_[102337]_  = A265 & A203;
  assign \new_[102338]_  = \new_[102337]_  & \new_[102334]_ ;
  assign \new_[102339]_  = \new_[102338]_  & \new_[102331]_ ;
  assign \new_[102342]_  = ~A267 & ~A266;
  assign \new_[102345]_  = A269 & ~A268;
  assign \new_[102346]_  = \new_[102345]_  & \new_[102342]_ ;
  assign \new_[102349]_  = ~A299 & A298;
  assign \new_[102353]_  = A302 & ~A301;
  assign \new_[102354]_  = ~A300 & \new_[102353]_ ;
  assign \new_[102355]_  = \new_[102354]_  & \new_[102349]_ ;
  assign \new_[102356]_  = \new_[102355]_  & \new_[102346]_ ;
  assign \new_[102359]_  = ~A168 & A170;
  assign \new_[102362]_  = A200 & ~A199;
  assign \new_[102363]_  = \new_[102362]_  & \new_[102359]_ ;
  assign \new_[102366]_  = ~A202 & ~A201;
  assign \new_[102369]_  = A265 & A203;
  assign \new_[102370]_  = \new_[102369]_  & \new_[102366]_ ;
  assign \new_[102371]_  = \new_[102370]_  & \new_[102363]_ ;
  assign \new_[102374]_  = ~A267 & ~A266;
  assign \new_[102377]_  = A269 & ~A268;
  assign \new_[102378]_  = \new_[102377]_  & \new_[102374]_ ;
  assign \new_[102381]_  = A299 & ~A298;
  assign \new_[102385]_  = A302 & ~A301;
  assign \new_[102386]_  = ~A300 & \new_[102385]_ ;
  assign \new_[102387]_  = \new_[102386]_  & \new_[102381]_ ;
  assign \new_[102388]_  = \new_[102387]_  & \new_[102378]_ ;
  assign \new_[102391]_  = ~A168 & A170;
  assign \new_[102394]_  = ~A200 & A199;
  assign \new_[102395]_  = \new_[102394]_  & \new_[102391]_ ;
  assign \new_[102398]_  = ~A202 & ~A201;
  assign \new_[102401]_  = ~A265 & A203;
  assign \new_[102402]_  = \new_[102401]_  & \new_[102398]_ ;
  assign \new_[102403]_  = \new_[102402]_  & \new_[102395]_ ;
  assign \new_[102406]_  = ~A267 & A266;
  assign \new_[102409]_  = A269 & ~A268;
  assign \new_[102410]_  = \new_[102409]_  & \new_[102406]_ ;
  assign \new_[102413]_  = ~A299 & A298;
  assign \new_[102417]_  = A302 & ~A301;
  assign \new_[102418]_  = ~A300 & \new_[102417]_ ;
  assign \new_[102419]_  = \new_[102418]_  & \new_[102413]_ ;
  assign \new_[102420]_  = \new_[102419]_  & \new_[102410]_ ;
  assign \new_[102423]_  = ~A168 & A170;
  assign \new_[102426]_  = ~A200 & A199;
  assign \new_[102427]_  = \new_[102426]_  & \new_[102423]_ ;
  assign \new_[102430]_  = ~A202 & ~A201;
  assign \new_[102433]_  = ~A265 & A203;
  assign \new_[102434]_  = \new_[102433]_  & \new_[102430]_ ;
  assign \new_[102435]_  = \new_[102434]_  & \new_[102427]_ ;
  assign \new_[102438]_  = ~A267 & A266;
  assign \new_[102441]_  = A269 & ~A268;
  assign \new_[102442]_  = \new_[102441]_  & \new_[102438]_ ;
  assign \new_[102445]_  = A299 & ~A298;
  assign \new_[102449]_  = A302 & ~A301;
  assign \new_[102450]_  = ~A300 & \new_[102449]_ ;
  assign \new_[102451]_  = \new_[102450]_  & \new_[102445]_ ;
  assign \new_[102452]_  = \new_[102451]_  & \new_[102442]_ ;
  assign \new_[102455]_  = ~A168 & A170;
  assign \new_[102458]_  = ~A200 & A199;
  assign \new_[102459]_  = \new_[102458]_  & \new_[102455]_ ;
  assign \new_[102462]_  = ~A202 & ~A201;
  assign \new_[102465]_  = A265 & A203;
  assign \new_[102466]_  = \new_[102465]_  & \new_[102462]_ ;
  assign \new_[102467]_  = \new_[102466]_  & \new_[102459]_ ;
  assign \new_[102470]_  = ~A267 & ~A266;
  assign \new_[102473]_  = A269 & ~A268;
  assign \new_[102474]_  = \new_[102473]_  & \new_[102470]_ ;
  assign \new_[102477]_  = ~A299 & A298;
  assign \new_[102481]_  = A302 & ~A301;
  assign \new_[102482]_  = ~A300 & \new_[102481]_ ;
  assign \new_[102483]_  = \new_[102482]_  & \new_[102477]_ ;
  assign \new_[102484]_  = \new_[102483]_  & \new_[102474]_ ;
  assign \new_[102487]_  = ~A168 & A170;
  assign \new_[102490]_  = ~A200 & A199;
  assign \new_[102491]_  = \new_[102490]_  & \new_[102487]_ ;
  assign \new_[102494]_  = ~A202 & ~A201;
  assign \new_[102497]_  = A265 & A203;
  assign \new_[102498]_  = \new_[102497]_  & \new_[102494]_ ;
  assign \new_[102499]_  = \new_[102498]_  & \new_[102491]_ ;
  assign \new_[102502]_  = ~A267 & ~A266;
  assign \new_[102505]_  = A269 & ~A268;
  assign \new_[102506]_  = \new_[102505]_  & \new_[102502]_ ;
  assign \new_[102509]_  = A299 & ~A298;
  assign \new_[102513]_  = A302 & ~A301;
  assign \new_[102514]_  = ~A300 & \new_[102513]_ ;
  assign \new_[102515]_  = \new_[102514]_  & \new_[102509]_ ;
  assign \new_[102516]_  = \new_[102515]_  & \new_[102506]_ ;
  assign \new_[102519]_  = ~A168 & A169;
  assign \new_[102522]_  = A200 & ~A199;
  assign \new_[102523]_  = \new_[102522]_  & \new_[102519]_ ;
  assign \new_[102526]_  = ~A202 & ~A201;
  assign \new_[102529]_  = ~A265 & A203;
  assign \new_[102530]_  = \new_[102529]_  & \new_[102526]_ ;
  assign \new_[102531]_  = \new_[102530]_  & \new_[102523]_ ;
  assign \new_[102534]_  = ~A267 & A266;
  assign \new_[102537]_  = A269 & ~A268;
  assign \new_[102538]_  = \new_[102537]_  & \new_[102534]_ ;
  assign \new_[102541]_  = ~A299 & A298;
  assign \new_[102545]_  = A302 & ~A301;
  assign \new_[102546]_  = ~A300 & \new_[102545]_ ;
  assign \new_[102547]_  = \new_[102546]_  & \new_[102541]_ ;
  assign \new_[102548]_  = \new_[102547]_  & \new_[102538]_ ;
  assign \new_[102551]_  = ~A168 & A169;
  assign \new_[102554]_  = A200 & ~A199;
  assign \new_[102555]_  = \new_[102554]_  & \new_[102551]_ ;
  assign \new_[102558]_  = ~A202 & ~A201;
  assign \new_[102561]_  = ~A265 & A203;
  assign \new_[102562]_  = \new_[102561]_  & \new_[102558]_ ;
  assign \new_[102563]_  = \new_[102562]_  & \new_[102555]_ ;
  assign \new_[102566]_  = ~A267 & A266;
  assign \new_[102569]_  = A269 & ~A268;
  assign \new_[102570]_  = \new_[102569]_  & \new_[102566]_ ;
  assign \new_[102573]_  = A299 & ~A298;
  assign \new_[102577]_  = A302 & ~A301;
  assign \new_[102578]_  = ~A300 & \new_[102577]_ ;
  assign \new_[102579]_  = \new_[102578]_  & \new_[102573]_ ;
  assign \new_[102580]_  = \new_[102579]_  & \new_[102570]_ ;
  assign \new_[102583]_  = ~A168 & A169;
  assign \new_[102586]_  = A200 & ~A199;
  assign \new_[102587]_  = \new_[102586]_  & \new_[102583]_ ;
  assign \new_[102590]_  = ~A202 & ~A201;
  assign \new_[102593]_  = A265 & A203;
  assign \new_[102594]_  = \new_[102593]_  & \new_[102590]_ ;
  assign \new_[102595]_  = \new_[102594]_  & \new_[102587]_ ;
  assign \new_[102598]_  = ~A267 & ~A266;
  assign \new_[102601]_  = A269 & ~A268;
  assign \new_[102602]_  = \new_[102601]_  & \new_[102598]_ ;
  assign \new_[102605]_  = ~A299 & A298;
  assign \new_[102609]_  = A302 & ~A301;
  assign \new_[102610]_  = ~A300 & \new_[102609]_ ;
  assign \new_[102611]_  = \new_[102610]_  & \new_[102605]_ ;
  assign \new_[102612]_  = \new_[102611]_  & \new_[102602]_ ;
  assign \new_[102615]_  = ~A168 & A169;
  assign \new_[102618]_  = A200 & ~A199;
  assign \new_[102619]_  = \new_[102618]_  & \new_[102615]_ ;
  assign \new_[102622]_  = ~A202 & ~A201;
  assign \new_[102625]_  = A265 & A203;
  assign \new_[102626]_  = \new_[102625]_  & \new_[102622]_ ;
  assign \new_[102627]_  = \new_[102626]_  & \new_[102619]_ ;
  assign \new_[102630]_  = ~A267 & ~A266;
  assign \new_[102633]_  = A269 & ~A268;
  assign \new_[102634]_  = \new_[102633]_  & \new_[102630]_ ;
  assign \new_[102637]_  = A299 & ~A298;
  assign \new_[102641]_  = A302 & ~A301;
  assign \new_[102642]_  = ~A300 & \new_[102641]_ ;
  assign \new_[102643]_  = \new_[102642]_  & \new_[102637]_ ;
  assign \new_[102644]_  = \new_[102643]_  & \new_[102634]_ ;
  assign \new_[102647]_  = ~A168 & A169;
  assign \new_[102650]_  = ~A200 & A199;
  assign \new_[102651]_  = \new_[102650]_  & \new_[102647]_ ;
  assign \new_[102654]_  = ~A202 & ~A201;
  assign \new_[102657]_  = ~A265 & A203;
  assign \new_[102658]_  = \new_[102657]_  & \new_[102654]_ ;
  assign \new_[102659]_  = \new_[102658]_  & \new_[102651]_ ;
  assign \new_[102662]_  = ~A267 & A266;
  assign \new_[102665]_  = A269 & ~A268;
  assign \new_[102666]_  = \new_[102665]_  & \new_[102662]_ ;
  assign \new_[102669]_  = ~A299 & A298;
  assign \new_[102673]_  = A302 & ~A301;
  assign \new_[102674]_  = ~A300 & \new_[102673]_ ;
  assign \new_[102675]_  = \new_[102674]_  & \new_[102669]_ ;
  assign \new_[102676]_  = \new_[102675]_  & \new_[102666]_ ;
  assign \new_[102679]_  = ~A168 & A169;
  assign \new_[102682]_  = ~A200 & A199;
  assign \new_[102683]_  = \new_[102682]_  & \new_[102679]_ ;
  assign \new_[102686]_  = ~A202 & ~A201;
  assign \new_[102689]_  = ~A265 & A203;
  assign \new_[102690]_  = \new_[102689]_  & \new_[102686]_ ;
  assign \new_[102691]_  = \new_[102690]_  & \new_[102683]_ ;
  assign \new_[102694]_  = ~A267 & A266;
  assign \new_[102697]_  = A269 & ~A268;
  assign \new_[102698]_  = \new_[102697]_  & \new_[102694]_ ;
  assign \new_[102701]_  = A299 & ~A298;
  assign \new_[102705]_  = A302 & ~A301;
  assign \new_[102706]_  = ~A300 & \new_[102705]_ ;
  assign \new_[102707]_  = \new_[102706]_  & \new_[102701]_ ;
  assign \new_[102708]_  = \new_[102707]_  & \new_[102698]_ ;
  assign \new_[102711]_  = ~A168 & A169;
  assign \new_[102714]_  = ~A200 & A199;
  assign \new_[102715]_  = \new_[102714]_  & \new_[102711]_ ;
  assign \new_[102718]_  = ~A202 & ~A201;
  assign \new_[102721]_  = A265 & A203;
  assign \new_[102722]_  = \new_[102721]_  & \new_[102718]_ ;
  assign \new_[102723]_  = \new_[102722]_  & \new_[102715]_ ;
  assign \new_[102726]_  = ~A267 & ~A266;
  assign \new_[102729]_  = A269 & ~A268;
  assign \new_[102730]_  = \new_[102729]_  & \new_[102726]_ ;
  assign \new_[102733]_  = ~A299 & A298;
  assign \new_[102737]_  = A302 & ~A301;
  assign \new_[102738]_  = ~A300 & \new_[102737]_ ;
  assign \new_[102739]_  = \new_[102738]_  & \new_[102733]_ ;
  assign \new_[102740]_  = \new_[102739]_  & \new_[102730]_ ;
  assign \new_[102743]_  = ~A168 & A169;
  assign \new_[102746]_  = ~A200 & A199;
  assign \new_[102747]_  = \new_[102746]_  & \new_[102743]_ ;
  assign \new_[102750]_  = ~A202 & ~A201;
  assign \new_[102753]_  = A265 & A203;
  assign \new_[102754]_  = \new_[102753]_  & \new_[102750]_ ;
  assign \new_[102755]_  = \new_[102754]_  & \new_[102747]_ ;
  assign \new_[102758]_  = ~A267 & ~A266;
  assign \new_[102761]_  = A269 & ~A268;
  assign \new_[102762]_  = \new_[102761]_  & \new_[102758]_ ;
  assign \new_[102765]_  = A299 & ~A298;
  assign \new_[102769]_  = A302 & ~A301;
  assign \new_[102770]_  = ~A300 & \new_[102769]_ ;
  assign \new_[102771]_  = \new_[102770]_  & \new_[102765]_ ;
  assign \new_[102772]_  = \new_[102771]_  & \new_[102762]_ ;
  assign \new_[102775]_  = ~A169 & ~A170;
  assign \new_[102778]_  = ~A199 & A168;
  assign \new_[102779]_  = \new_[102778]_  & \new_[102775]_ ;
  assign \new_[102782]_  = A201 & A200;
  assign \new_[102785]_  = ~A265 & A202;
  assign \new_[102786]_  = \new_[102785]_  & \new_[102782]_ ;
  assign \new_[102787]_  = \new_[102786]_  & \new_[102779]_ ;
  assign \new_[102790]_  = ~A267 & A266;
  assign \new_[102793]_  = A269 & ~A268;
  assign \new_[102794]_  = \new_[102793]_  & \new_[102790]_ ;
  assign \new_[102797]_  = ~A299 & A298;
  assign \new_[102801]_  = A302 & ~A301;
  assign \new_[102802]_  = ~A300 & \new_[102801]_ ;
  assign \new_[102803]_  = \new_[102802]_  & \new_[102797]_ ;
  assign \new_[102804]_  = \new_[102803]_  & \new_[102794]_ ;
  assign \new_[102807]_  = ~A169 & ~A170;
  assign \new_[102810]_  = ~A199 & A168;
  assign \new_[102811]_  = \new_[102810]_  & \new_[102807]_ ;
  assign \new_[102814]_  = A201 & A200;
  assign \new_[102817]_  = ~A265 & A202;
  assign \new_[102818]_  = \new_[102817]_  & \new_[102814]_ ;
  assign \new_[102819]_  = \new_[102818]_  & \new_[102811]_ ;
  assign \new_[102822]_  = ~A267 & A266;
  assign \new_[102825]_  = A269 & ~A268;
  assign \new_[102826]_  = \new_[102825]_  & \new_[102822]_ ;
  assign \new_[102829]_  = A299 & ~A298;
  assign \new_[102833]_  = A302 & ~A301;
  assign \new_[102834]_  = ~A300 & \new_[102833]_ ;
  assign \new_[102835]_  = \new_[102834]_  & \new_[102829]_ ;
  assign \new_[102836]_  = \new_[102835]_  & \new_[102826]_ ;
  assign \new_[102839]_  = ~A169 & ~A170;
  assign \new_[102842]_  = ~A199 & A168;
  assign \new_[102843]_  = \new_[102842]_  & \new_[102839]_ ;
  assign \new_[102846]_  = A201 & A200;
  assign \new_[102849]_  = A265 & A202;
  assign \new_[102850]_  = \new_[102849]_  & \new_[102846]_ ;
  assign \new_[102851]_  = \new_[102850]_  & \new_[102843]_ ;
  assign \new_[102854]_  = ~A267 & ~A266;
  assign \new_[102857]_  = A269 & ~A268;
  assign \new_[102858]_  = \new_[102857]_  & \new_[102854]_ ;
  assign \new_[102861]_  = ~A299 & A298;
  assign \new_[102865]_  = A302 & ~A301;
  assign \new_[102866]_  = ~A300 & \new_[102865]_ ;
  assign \new_[102867]_  = \new_[102866]_  & \new_[102861]_ ;
  assign \new_[102868]_  = \new_[102867]_  & \new_[102858]_ ;
  assign \new_[102871]_  = ~A169 & ~A170;
  assign \new_[102874]_  = ~A199 & A168;
  assign \new_[102875]_  = \new_[102874]_  & \new_[102871]_ ;
  assign \new_[102878]_  = A201 & A200;
  assign \new_[102881]_  = A265 & A202;
  assign \new_[102882]_  = \new_[102881]_  & \new_[102878]_ ;
  assign \new_[102883]_  = \new_[102882]_  & \new_[102875]_ ;
  assign \new_[102886]_  = ~A267 & ~A266;
  assign \new_[102889]_  = A269 & ~A268;
  assign \new_[102890]_  = \new_[102889]_  & \new_[102886]_ ;
  assign \new_[102893]_  = A299 & ~A298;
  assign \new_[102897]_  = A302 & ~A301;
  assign \new_[102898]_  = ~A300 & \new_[102897]_ ;
  assign \new_[102899]_  = \new_[102898]_  & \new_[102893]_ ;
  assign \new_[102900]_  = \new_[102899]_  & \new_[102890]_ ;
  assign \new_[102903]_  = ~A169 & ~A170;
  assign \new_[102906]_  = ~A199 & A168;
  assign \new_[102907]_  = \new_[102906]_  & \new_[102903]_ ;
  assign \new_[102910]_  = A201 & A200;
  assign \new_[102913]_  = ~A265 & ~A203;
  assign \new_[102914]_  = \new_[102913]_  & \new_[102910]_ ;
  assign \new_[102915]_  = \new_[102914]_  & \new_[102907]_ ;
  assign \new_[102918]_  = ~A267 & A266;
  assign \new_[102921]_  = A269 & ~A268;
  assign \new_[102922]_  = \new_[102921]_  & \new_[102918]_ ;
  assign \new_[102925]_  = ~A299 & A298;
  assign \new_[102929]_  = A302 & ~A301;
  assign \new_[102930]_  = ~A300 & \new_[102929]_ ;
  assign \new_[102931]_  = \new_[102930]_  & \new_[102925]_ ;
  assign \new_[102932]_  = \new_[102931]_  & \new_[102922]_ ;
  assign \new_[102935]_  = ~A169 & ~A170;
  assign \new_[102938]_  = ~A199 & A168;
  assign \new_[102939]_  = \new_[102938]_  & \new_[102935]_ ;
  assign \new_[102942]_  = A201 & A200;
  assign \new_[102945]_  = ~A265 & ~A203;
  assign \new_[102946]_  = \new_[102945]_  & \new_[102942]_ ;
  assign \new_[102947]_  = \new_[102946]_  & \new_[102939]_ ;
  assign \new_[102950]_  = ~A267 & A266;
  assign \new_[102953]_  = A269 & ~A268;
  assign \new_[102954]_  = \new_[102953]_  & \new_[102950]_ ;
  assign \new_[102957]_  = A299 & ~A298;
  assign \new_[102961]_  = A302 & ~A301;
  assign \new_[102962]_  = ~A300 & \new_[102961]_ ;
  assign \new_[102963]_  = \new_[102962]_  & \new_[102957]_ ;
  assign \new_[102964]_  = \new_[102963]_  & \new_[102954]_ ;
  assign \new_[102967]_  = ~A169 & ~A170;
  assign \new_[102970]_  = ~A199 & A168;
  assign \new_[102971]_  = \new_[102970]_  & \new_[102967]_ ;
  assign \new_[102974]_  = A201 & A200;
  assign \new_[102977]_  = A265 & ~A203;
  assign \new_[102978]_  = \new_[102977]_  & \new_[102974]_ ;
  assign \new_[102979]_  = \new_[102978]_  & \new_[102971]_ ;
  assign \new_[102982]_  = ~A267 & ~A266;
  assign \new_[102985]_  = A269 & ~A268;
  assign \new_[102986]_  = \new_[102985]_  & \new_[102982]_ ;
  assign \new_[102989]_  = ~A299 & A298;
  assign \new_[102993]_  = A302 & ~A301;
  assign \new_[102994]_  = ~A300 & \new_[102993]_ ;
  assign \new_[102995]_  = \new_[102994]_  & \new_[102989]_ ;
  assign \new_[102996]_  = \new_[102995]_  & \new_[102986]_ ;
  assign \new_[102999]_  = ~A169 & ~A170;
  assign \new_[103002]_  = ~A199 & A168;
  assign \new_[103003]_  = \new_[103002]_  & \new_[102999]_ ;
  assign \new_[103006]_  = A201 & A200;
  assign \new_[103009]_  = A265 & ~A203;
  assign \new_[103010]_  = \new_[103009]_  & \new_[103006]_ ;
  assign \new_[103011]_  = \new_[103010]_  & \new_[103003]_ ;
  assign \new_[103014]_  = ~A267 & ~A266;
  assign \new_[103017]_  = A269 & ~A268;
  assign \new_[103018]_  = \new_[103017]_  & \new_[103014]_ ;
  assign \new_[103021]_  = A299 & ~A298;
  assign \new_[103025]_  = A302 & ~A301;
  assign \new_[103026]_  = ~A300 & \new_[103025]_ ;
  assign \new_[103027]_  = \new_[103026]_  & \new_[103021]_ ;
  assign \new_[103028]_  = \new_[103027]_  & \new_[103018]_ ;
  assign \new_[103031]_  = ~A169 & ~A170;
  assign \new_[103034]_  = ~A199 & A168;
  assign \new_[103035]_  = \new_[103034]_  & \new_[103031]_ ;
  assign \new_[103038]_  = ~A201 & A200;
  assign \new_[103041]_  = A203 & ~A202;
  assign \new_[103042]_  = \new_[103041]_  & \new_[103038]_ ;
  assign \new_[103043]_  = \new_[103042]_  & \new_[103035]_ ;
  assign \new_[103046]_  = A266 & ~A265;
  assign \new_[103049]_  = A268 & A267;
  assign \new_[103050]_  = \new_[103049]_  & \new_[103046]_ ;
  assign \new_[103053]_  = ~A299 & A298;
  assign \new_[103057]_  = A302 & ~A301;
  assign \new_[103058]_  = ~A300 & \new_[103057]_ ;
  assign \new_[103059]_  = \new_[103058]_  & \new_[103053]_ ;
  assign \new_[103060]_  = \new_[103059]_  & \new_[103050]_ ;
  assign \new_[103063]_  = ~A169 & ~A170;
  assign \new_[103066]_  = ~A199 & A168;
  assign \new_[103067]_  = \new_[103066]_  & \new_[103063]_ ;
  assign \new_[103070]_  = ~A201 & A200;
  assign \new_[103073]_  = A203 & ~A202;
  assign \new_[103074]_  = \new_[103073]_  & \new_[103070]_ ;
  assign \new_[103075]_  = \new_[103074]_  & \new_[103067]_ ;
  assign \new_[103078]_  = A266 & ~A265;
  assign \new_[103081]_  = A268 & A267;
  assign \new_[103082]_  = \new_[103081]_  & \new_[103078]_ ;
  assign \new_[103085]_  = A299 & ~A298;
  assign \new_[103089]_  = A302 & ~A301;
  assign \new_[103090]_  = ~A300 & \new_[103089]_ ;
  assign \new_[103091]_  = \new_[103090]_  & \new_[103085]_ ;
  assign \new_[103092]_  = \new_[103091]_  & \new_[103082]_ ;
  assign \new_[103095]_  = ~A169 & ~A170;
  assign \new_[103098]_  = ~A199 & A168;
  assign \new_[103099]_  = \new_[103098]_  & \new_[103095]_ ;
  assign \new_[103102]_  = ~A201 & A200;
  assign \new_[103105]_  = A203 & ~A202;
  assign \new_[103106]_  = \new_[103105]_  & \new_[103102]_ ;
  assign \new_[103107]_  = \new_[103106]_  & \new_[103099]_ ;
  assign \new_[103110]_  = A266 & ~A265;
  assign \new_[103113]_  = ~A269 & A267;
  assign \new_[103114]_  = \new_[103113]_  & \new_[103110]_ ;
  assign \new_[103117]_  = ~A299 & A298;
  assign \new_[103121]_  = A302 & ~A301;
  assign \new_[103122]_  = ~A300 & \new_[103121]_ ;
  assign \new_[103123]_  = \new_[103122]_  & \new_[103117]_ ;
  assign \new_[103124]_  = \new_[103123]_  & \new_[103114]_ ;
  assign \new_[103127]_  = ~A169 & ~A170;
  assign \new_[103130]_  = ~A199 & A168;
  assign \new_[103131]_  = \new_[103130]_  & \new_[103127]_ ;
  assign \new_[103134]_  = ~A201 & A200;
  assign \new_[103137]_  = A203 & ~A202;
  assign \new_[103138]_  = \new_[103137]_  & \new_[103134]_ ;
  assign \new_[103139]_  = \new_[103138]_  & \new_[103131]_ ;
  assign \new_[103142]_  = A266 & ~A265;
  assign \new_[103145]_  = ~A269 & A267;
  assign \new_[103146]_  = \new_[103145]_  & \new_[103142]_ ;
  assign \new_[103149]_  = A299 & ~A298;
  assign \new_[103153]_  = A302 & ~A301;
  assign \new_[103154]_  = ~A300 & \new_[103153]_ ;
  assign \new_[103155]_  = \new_[103154]_  & \new_[103149]_ ;
  assign \new_[103156]_  = \new_[103155]_  & \new_[103146]_ ;
  assign \new_[103159]_  = ~A169 & ~A170;
  assign \new_[103162]_  = ~A199 & A168;
  assign \new_[103163]_  = \new_[103162]_  & \new_[103159]_ ;
  assign \new_[103166]_  = ~A201 & A200;
  assign \new_[103169]_  = A203 & ~A202;
  assign \new_[103170]_  = \new_[103169]_  & \new_[103166]_ ;
  assign \new_[103171]_  = \new_[103170]_  & \new_[103163]_ ;
  assign \new_[103174]_  = A266 & ~A265;
  assign \new_[103177]_  = ~A268 & ~A267;
  assign \new_[103178]_  = \new_[103177]_  & \new_[103174]_ ;
  assign \new_[103181]_  = A298 & A269;
  assign \new_[103185]_  = A301 & A300;
  assign \new_[103186]_  = ~A299 & \new_[103185]_ ;
  assign \new_[103187]_  = \new_[103186]_  & \new_[103181]_ ;
  assign \new_[103188]_  = \new_[103187]_  & \new_[103178]_ ;
  assign \new_[103191]_  = ~A169 & ~A170;
  assign \new_[103194]_  = ~A199 & A168;
  assign \new_[103195]_  = \new_[103194]_  & \new_[103191]_ ;
  assign \new_[103198]_  = ~A201 & A200;
  assign \new_[103201]_  = A203 & ~A202;
  assign \new_[103202]_  = \new_[103201]_  & \new_[103198]_ ;
  assign \new_[103203]_  = \new_[103202]_  & \new_[103195]_ ;
  assign \new_[103206]_  = A266 & ~A265;
  assign \new_[103209]_  = ~A268 & ~A267;
  assign \new_[103210]_  = \new_[103209]_  & \new_[103206]_ ;
  assign \new_[103213]_  = A298 & A269;
  assign \new_[103217]_  = ~A302 & A300;
  assign \new_[103218]_  = ~A299 & \new_[103217]_ ;
  assign \new_[103219]_  = \new_[103218]_  & \new_[103213]_ ;
  assign \new_[103220]_  = \new_[103219]_  & \new_[103210]_ ;
  assign \new_[103223]_  = ~A169 & ~A170;
  assign \new_[103226]_  = ~A199 & A168;
  assign \new_[103227]_  = \new_[103226]_  & \new_[103223]_ ;
  assign \new_[103230]_  = ~A201 & A200;
  assign \new_[103233]_  = A203 & ~A202;
  assign \new_[103234]_  = \new_[103233]_  & \new_[103230]_ ;
  assign \new_[103235]_  = \new_[103234]_  & \new_[103227]_ ;
  assign \new_[103238]_  = A266 & ~A265;
  assign \new_[103241]_  = ~A268 & ~A267;
  assign \new_[103242]_  = \new_[103241]_  & \new_[103238]_ ;
  assign \new_[103245]_  = ~A298 & A269;
  assign \new_[103249]_  = A301 & A300;
  assign \new_[103250]_  = A299 & \new_[103249]_ ;
  assign \new_[103251]_  = \new_[103250]_  & \new_[103245]_ ;
  assign \new_[103252]_  = \new_[103251]_  & \new_[103242]_ ;
  assign \new_[103255]_  = ~A169 & ~A170;
  assign \new_[103258]_  = ~A199 & A168;
  assign \new_[103259]_  = \new_[103258]_  & \new_[103255]_ ;
  assign \new_[103262]_  = ~A201 & A200;
  assign \new_[103265]_  = A203 & ~A202;
  assign \new_[103266]_  = \new_[103265]_  & \new_[103262]_ ;
  assign \new_[103267]_  = \new_[103266]_  & \new_[103259]_ ;
  assign \new_[103270]_  = A266 & ~A265;
  assign \new_[103273]_  = ~A268 & ~A267;
  assign \new_[103274]_  = \new_[103273]_  & \new_[103270]_ ;
  assign \new_[103277]_  = ~A298 & A269;
  assign \new_[103281]_  = ~A302 & A300;
  assign \new_[103282]_  = A299 & \new_[103281]_ ;
  assign \new_[103283]_  = \new_[103282]_  & \new_[103277]_ ;
  assign \new_[103284]_  = \new_[103283]_  & \new_[103274]_ ;
  assign \new_[103287]_  = ~A169 & ~A170;
  assign \new_[103290]_  = ~A199 & A168;
  assign \new_[103291]_  = \new_[103290]_  & \new_[103287]_ ;
  assign \new_[103294]_  = ~A201 & A200;
  assign \new_[103297]_  = A203 & ~A202;
  assign \new_[103298]_  = \new_[103297]_  & \new_[103294]_ ;
  assign \new_[103299]_  = \new_[103298]_  & \new_[103291]_ ;
  assign \new_[103302]_  = ~A266 & A265;
  assign \new_[103305]_  = A268 & A267;
  assign \new_[103306]_  = \new_[103305]_  & \new_[103302]_ ;
  assign \new_[103309]_  = ~A299 & A298;
  assign \new_[103313]_  = A302 & ~A301;
  assign \new_[103314]_  = ~A300 & \new_[103313]_ ;
  assign \new_[103315]_  = \new_[103314]_  & \new_[103309]_ ;
  assign \new_[103316]_  = \new_[103315]_  & \new_[103306]_ ;
  assign \new_[103319]_  = ~A169 & ~A170;
  assign \new_[103322]_  = ~A199 & A168;
  assign \new_[103323]_  = \new_[103322]_  & \new_[103319]_ ;
  assign \new_[103326]_  = ~A201 & A200;
  assign \new_[103329]_  = A203 & ~A202;
  assign \new_[103330]_  = \new_[103329]_  & \new_[103326]_ ;
  assign \new_[103331]_  = \new_[103330]_  & \new_[103323]_ ;
  assign \new_[103334]_  = ~A266 & A265;
  assign \new_[103337]_  = A268 & A267;
  assign \new_[103338]_  = \new_[103337]_  & \new_[103334]_ ;
  assign \new_[103341]_  = A299 & ~A298;
  assign \new_[103345]_  = A302 & ~A301;
  assign \new_[103346]_  = ~A300 & \new_[103345]_ ;
  assign \new_[103347]_  = \new_[103346]_  & \new_[103341]_ ;
  assign \new_[103348]_  = \new_[103347]_  & \new_[103338]_ ;
  assign \new_[103351]_  = ~A169 & ~A170;
  assign \new_[103354]_  = ~A199 & A168;
  assign \new_[103355]_  = \new_[103354]_  & \new_[103351]_ ;
  assign \new_[103358]_  = ~A201 & A200;
  assign \new_[103361]_  = A203 & ~A202;
  assign \new_[103362]_  = \new_[103361]_  & \new_[103358]_ ;
  assign \new_[103363]_  = \new_[103362]_  & \new_[103355]_ ;
  assign \new_[103366]_  = ~A266 & A265;
  assign \new_[103369]_  = ~A269 & A267;
  assign \new_[103370]_  = \new_[103369]_  & \new_[103366]_ ;
  assign \new_[103373]_  = ~A299 & A298;
  assign \new_[103377]_  = A302 & ~A301;
  assign \new_[103378]_  = ~A300 & \new_[103377]_ ;
  assign \new_[103379]_  = \new_[103378]_  & \new_[103373]_ ;
  assign \new_[103380]_  = \new_[103379]_  & \new_[103370]_ ;
  assign \new_[103383]_  = ~A169 & ~A170;
  assign \new_[103386]_  = ~A199 & A168;
  assign \new_[103387]_  = \new_[103386]_  & \new_[103383]_ ;
  assign \new_[103390]_  = ~A201 & A200;
  assign \new_[103393]_  = A203 & ~A202;
  assign \new_[103394]_  = \new_[103393]_  & \new_[103390]_ ;
  assign \new_[103395]_  = \new_[103394]_  & \new_[103387]_ ;
  assign \new_[103398]_  = ~A266 & A265;
  assign \new_[103401]_  = ~A269 & A267;
  assign \new_[103402]_  = \new_[103401]_  & \new_[103398]_ ;
  assign \new_[103405]_  = A299 & ~A298;
  assign \new_[103409]_  = A302 & ~A301;
  assign \new_[103410]_  = ~A300 & \new_[103409]_ ;
  assign \new_[103411]_  = \new_[103410]_  & \new_[103405]_ ;
  assign \new_[103412]_  = \new_[103411]_  & \new_[103402]_ ;
  assign \new_[103415]_  = ~A169 & ~A170;
  assign \new_[103418]_  = ~A199 & A168;
  assign \new_[103419]_  = \new_[103418]_  & \new_[103415]_ ;
  assign \new_[103422]_  = ~A201 & A200;
  assign \new_[103425]_  = A203 & ~A202;
  assign \new_[103426]_  = \new_[103425]_  & \new_[103422]_ ;
  assign \new_[103427]_  = \new_[103426]_  & \new_[103419]_ ;
  assign \new_[103430]_  = ~A266 & A265;
  assign \new_[103433]_  = ~A268 & ~A267;
  assign \new_[103434]_  = \new_[103433]_  & \new_[103430]_ ;
  assign \new_[103437]_  = A298 & A269;
  assign \new_[103441]_  = A301 & A300;
  assign \new_[103442]_  = ~A299 & \new_[103441]_ ;
  assign \new_[103443]_  = \new_[103442]_  & \new_[103437]_ ;
  assign \new_[103444]_  = \new_[103443]_  & \new_[103434]_ ;
  assign \new_[103447]_  = ~A169 & ~A170;
  assign \new_[103450]_  = ~A199 & A168;
  assign \new_[103451]_  = \new_[103450]_  & \new_[103447]_ ;
  assign \new_[103454]_  = ~A201 & A200;
  assign \new_[103457]_  = A203 & ~A202;
  assign \new_[103458]_  = \new_[103457]_  & \new_[103454]_ ;
  assign \new_[103459]_  = \new_[103458]_  & \new_[103451]_ ;
  assign \new_[103462]_  = ~A266 & A265;
  assign \new_[103465]_  = ~A268 & ~A267;
  assign \new_[103466]_  = \new_[103465]_  & \new_[103462]_ ;
  assign \new_[103469]_  = A298 & A269;
  assign \new_[103473]_  = ~A302 & A300;
  assign \new_[103474]_  = ~A299 & \new_[103473]_ ;
  assign \new_[103475]_  = \new_[103474]_  & \new_[103469]_ ;
  assign \new_[103476]_  = \new_[103475]_  & \new_[103466]_ ;
  assign \new_[103479]_  = ~A169 & ~A170;
  assign \new_[103482]_  = ~A199 & A168;
  assign \new_[103483]_  = \new_[103482]_  & \new_[103479]_ ;
  assign \new_[103486]_  = ~A201 & A200;
  assign \new_[103489]_  = A203 & ~A202;
  assign \new_[103490]_  = \new_[103489]_  & \new_[103486]_ ;
  assign \new_[103491]_  = \new_[103490]_  & \new_[103483]_ ;
  assign \new_[103494]_  = ~A266 & A265;
  assign \new_[103497]_  = ~A268 & ~A267;
  assign \new_[103498]_  = \new_[103497]_  & \new_[103494]_ ;
  assign \new_[103501]_  = ~A298 & A269;
  assign \new_[103505]_  = A301 & A300;
  assign \new_[103506]_  = A299 & \new_[103505]_ ;
  assign \new_[103507]_  = \new_[103506]_  & \new_[103501]_ ;
  assign \new_[103508]_  = \new_[103507]_  & \new_[103498]_ ;
  assign \new_[103511]_  = ~A169 & ~A170;
  assign \new_[103514]_  = ~A199 & A168;
  assign \new_[103515]_  = \new_[103514]_  & \new_[103511]_ ;
  assign \new_[103518]_  = ~A201 & A200;
  assign \new_[103521]_  = A203 & ~A202;
  assign \new_[103522]_  = \new_[103521]_  & \new_[103518]_ ;
  assign \new_[103523]_  = \new_[103522]_  & \new_[103515]_ ;
  assign \new_[103526]_  = ~A266 & A265;
  assign \new_[103529]_  = ~A268 & ~A267;
  assign \new_[103530]_  = \new_[103529]_  & \new_[103526]_ ;
  assign \new_[103533]_  = ~A298 & A269;
  assign \new_[103537]_  = ~A302 & A300;
  assign \new_[103538]_  = A299 & \new_[103537]_ ;
  assign \new_[103539]_  = \new_[103538]_  & \new_[103533]_ ;
  assign \new_[103540]_  = \new_[103539]_  & \new_[103530]_ ;
  assign \new_[103543]_  = ~A169 & ~A170;
  assign \new_[103546]_  = A199 & A168;
  assign \new_[103547]_  = \new_[103546]_  & \new_[103543]_ ;
  assign \new_[103550]_  = A201 & ~A200;
  assign \new_[103553]_  = ~A265 & A202;
  assign \new_[103554]_  = \new_[103553]_  & \new_[103550]_ ;
  assign \new_[103555]_  = \new_[103554]_  & \new_[103547]_ ;
  assign \new_[103558]_  = ~A267 & A266;
  assign \new_[103561]_  = A269 & ~A268;
  assign \new_[103562]_  = \new_[103561]_  & \new_[103558]_ ;
  assign \new_[103565]_  = ~A299 & A298;
  assign \new_[103569]_  = A302 & ~A301;
  assign \new_[103570]_  = ~A300 & \new_[103569]_ ;
  assign \new_[103571]_  = \new_[103570]_  & \new_[103565]_ ;
  assign \new_[103572]_  = \new_[103571]_  & \new_[103562]_ ;
  assign \new_[103575]_  = ~A169 & ~A170;
  assign \new_[103578]_  = A199 & A168;
  assign \new_[103579]_  = \new_[103578]_  & \new_[103575]_ ;
  assign \new_[103582]_  = A201 & ~A200;
  assign \new_[103585]_  = ~A265 & A202;
  assign \new_[103586]_  = \new_[103585]_  & \new_[103582]_ ;
  assign \new_[103587]_  = \new_[103586]_  & \new_[103579]_ ;
  assign \new_[103590]_  = ~A267 & A266;
  assign \new_[103593]_  = A269 & ~A268;
  assign \new_[103594]_  = \new_[103593]_  & \new_[103590]_ ;
  assign \new_[103597]_  = A299 & ~A298;
  assign \new_[103601]_  = A302 & ~A301;
  assign \new_[103602]_  = ~A300 & \new_[103601]_ ;
  assign \new_[103603]_  = \new_[103602]_  & \new_[103597]_ ;
  assign \new_[103604]_  = \new_[103603]_  & \new_[103594]_ ;
  assign \new_[103607]_  = ~A169 & ~A170;
  assign \new_[103610]_  = A199 & A168;
  assign \new_[103611]_  = \new_[103610]_  & \new_[103607]_ ;
  assign \new_[103614]_  = A201 & ~A200;
  assign \new_[103617]_  = A265 & A202;
  assign \new_[103618]_  = \new_[103617]_  & \new_[103614]_ ;
  assign \new_[103619]_  = \new_[103618]_  & \new_[103611]_ ;
  assign \new_[103622]_  = ~A267 & ~A266;
  assign \new_[103625]_  = A269 & ~A268;
  assign \new_[103626]_  = \new_[103625]_  & \new_[103622]_ ;
  assign \new_[103629]_  = ~A299 & A298;
  assign \new_[103633]_  = A302 & ~A301;
  assign \new_[103634]_  = ~A300 & \new_[103633]_ ;
  assign \new_[103635]_  = \new_[103634]_  & \new_[103629]_ ;
  assign \new_[103636]_  = \new_[103635]_  & \new_[103626]_ ;
  assign \new_[103639]_  = ~A169 & ~A170;
  assign \new_[103642]_  = A199 & A168;
  assign \new_[103643]_  = \new_[103642]_  & \new_[103639]_ ;
  assign \new_[103646]_  = A201 & ~A200;
  assign \new_[103649]_  = A265 & A202;
  assign \new_[103650]_  = \new_[103649]_  & \new_[103646]_ ;
  assign \new_[103651]_  = \new_[103650]_  & \new_[103643]_ ;
  assign \new_[103654]_  = ~A267 & ~A266;
  assign \new_[103657]_  = A269 & ~A268;
  assign \new_[103658]_  = \new_[103657]_  & \new_[103654]_ ;
  assign \new_[103661]_  = A299 & ~A298;
  assign \new_[103665]_  = A302 & ~A301;
  assign \new_[103666]_  = ~A300 & \new_[103665]_ ;
  assign \new_[103667]_  = \new_[103666]_  & \new_[103661]_ ;
  assign \new_[103668]_  = \new_[103667]_  & \new_[103658]_ ;
  assign \new_[103671]_  = ~A169 & ~A170;
  assign \new_[103674]_  = A199 & A168;
  assign \new_[103675]_  = \new_[103674]_  & \new_[103671]_ ;
  assign \new_[103678]_  = A201 & ~A200;
  assign \new_[103681]_  = ~A265 & ~A203;
  assign \new_[103682]_  = \new_[103681]_  & \new_[103678]_ ;
  assign \new_[103683]_  = \new_[103682]_  & \new_[103675]_ ;
  assign \new_[103686]_  = ~A267 & A266;
  assign \new_[103689]_  = A269 & ~A268;
  assign \new_[103690]_  = \new_[103689]_  & \new_[103686]_ ;
  assign \new_[103693]_  = ~A299 & A298;
  assign \new_[103697]_  = A302 & ~A301;
  assign \new_[103698]_  = ~A300 & \new_[103697]_ ;
  assign \new_[103699]_  = \new_[103698]_  & \new_[103693]_ ;
  assign \new_[103700]_  = \new_[103699]_  & \new_[103690]_ ;
  assign \new_[103703]_  = ~A169 & ~A170;
  assign \new_[103706]_  = A199 & A168;
  assign \new_[103707]_  = \new_[103706]_  & \new_[103703]_ ;
  assign \new_[103710]_  = A201 & ~A200;
  assign \new_[103713]_  = ~A265 & ~A203;
  assign \new_[103714]_  = \new_[103713]_  & \new_[103710]_ ;
  assign \new_[103715]_  = \new_[103714]_  & \new_[103707]_ ;
  assign \new_[103718]_  = ~A267 & A266;
  assign \new_[103721]_  = A269 & ~A268;
  assign \new_[103722]_  = \new_[103721]_  & \new_[103718]_ ;
  assign \new_[103725]_  = A299 & ~A298;
  assign \new_[103729]_  = A302 & ~A301;
  assign \new_[103730]_  = ~A300 & \new_[103729]_ ;
  assign \new_[103731]_  = \new_[103730]_  & \new_[103725]_ ;
  assign \new_[103732]_  = \new_[103731]_  & \new_[103722]_ ;
  assign \new_[103735]_  = ~A169 & ~A170;
  assign \new_[103738]_  = A199 & A168;
  assign \new_[103739]_  = \new_[103738]_  & \new_[103735]_ ;
  assign \new_[103742]_  = A201 & ~A200;
  assign \new_[103745]_  = A265 & ~A203;
  assign \new_[103746]_  = \new_[103745]_  & \new_[103742]_ ;
  assign \new_[103747]_  = \new_[103746]_  & \new_[103739]_ ;
  assign \new_[103750]_  = ~A267 & ~A266;
  assign \new_[103753]_  = A269 & ~A268;
  assign \new_[103754]_  = \new_[103753]_  & \new_[103750]_ ;
  assign \new_[103757]_  = ~A299 & A298;
  assign \new_[103761]_  = A302 & ~A301;
  assign \new_[103762]_  = ~A300 & \new_[103761]_ ;
  assign \new_[103763]_  = \new_[103762]_  & \new_[103757]_ ;
  assign \new_[103764]_  = \new_[103763]_  & \new_[103754]_ ;
  assign \new_[103767]_  = ~A169 & ~A170;
  assign \new_[103770]_  = A199 & A168;
  assign \new_[103771]_  = \new_[103770]_  & \new_[103767]_ ;
  assign \new_[103774]_  = A201 & ~A200;
  assign \new_[103777]_  = A265 & ~A203;
  assign \new_[103778]_  = \new_[103777]_  & \new_[103774]_ ;
  assign \new_[103779]_  = \new_[103778]_  & \new_[103771]_ ;
  assign \new_[103782]_  = ~A267 & ~A266;
  assign \new_[103785]_  = A269 & ~A268;
  assign \new_[103786]_  = \new_[103785]_  & \new_[103782]_ ;
  assign \new_[103789]_  = A299 & ~A298;
  assign \new_[103793]_  = A302 & ~A301;
  assign \new_[103794]_  = ~A300 & \new_[103793]_ ;
  assign \new_[103795]_  = \new_[103794]_  & \new_[103789]_ ;
  assign \new_[103796]_  = \new_[103795]_  & \new_[103786]_ ;
  assign \new_[103799]_  = ~A169 & ~A170;
  assign \new_[103802]_  = A199 & A168;
  assign \new_[103803]_  = \new_[103802]_  & \new_[103799]_ ;
  assign \new_[103806]_  = ~A201 & ~A200;
  assign \new_[103809]_  = A203 & ~A202;
  assign \new_[103810]_  = \new_[103809]_  & \new_[103806]_ ;
  assign \new_[103811]_  = \new_[103810]_  & \new_[103803]_ ;
  assign \new_[103814]_  = A266 & ~A265;
  assign \new_[103817]_  = A268 & A267;
  assign \new_[103818]_  = \new_[103817]_  & \new_[103814]_ ;
  assign \new_[103821]_  = ~A299 & A298;
  assign \new_[103825]_  = A302 & ~A301;
  assign \new_[103826]_  = ~A300 & \new_[103825]_ ;
  assign \new_[103827]_  = \new_[103826]_  & \new_[103821]_ ;
  assign \new_[103828]_  = \new_[103827]_  & \new_[103818]_ ;
  assign \new_[103831]_  = ~A169 & ~A170;
  assign \new_[103834]_  = A199 & A168;
  assign \new_[103835]_  = \new_[103834]_  & \new_[103831]_ ;
  assign \new_[103838]_  = ~A201 & ~A200;
  assign \new_[103841]_  = A203 & ~A202;
  assign \new_[103842]_  = \new_[103841]_  & \new_[103838]_ ;
  assign \new_[103843]_  = \new_[103842]_  & \new_[103835]_ ;
  assign \new_[103846]_  = A266 & ~A265;
  assign \new_[103849]_  = A268 & A267;
  assign \new_[103850]_  = \new_[103849]_  & \new_[103846]_ ;
  assign \new_[103853]_  = A299 & ~A298;
  assign \new_[103857]_  = A302 & ~A301;
  assign \new_[103858]_  = ~A300 & \new_[103857]_ ;
  assign \new_[103859]_  = \new_[103858]_  & \new_[103853]_ ;
  assign \new_[103860]_  = \new_[103859]_  & \new_[103850]_ ;
  assign \new_[103863]_  = ~A169 & ~A170;
  assign \new_[103866]_  = A199 & A168;
  assign \new_[103867]_  = \new_[103866]_  & \new_[103863]_ ;
  assign \new_[103870]_  = ~A201 & ~A200;
  assign \new_[103873]_  = A203 & ~A202;
  assign \new_[103874]_  = \new_[103873]_  & \new_[103870]_ ;
  assign \new_[103875]_  = \new_[103874]_  & \new_[103867]_ ;
  assign \new_[103878]_  = A266 & ~A265;
  assign \new_[103881]_  = ~A269 & A267;
  assign \new_[103882]_  = \new_[103881]_  & \new_[103878]_ ;
  assign \new_[103885]_  = ~A299 & A298;
  assign \new_[103889]_  = A302 & ~A301;
  assign \new_[103890]_  = ~A300 & \new_[103889]_ ;
  assign \new_[103891]_  = \new_[103890]_  & \new_[103885]_ ;
  assign \new_[103892]_  = \new_[103891]_  & \new_[103882]_ ;
  assign \new_[103895]_  = ~A169 & ~A170;
  assign \new_[103898]_  = A199 & A168;
  assign \new_[103899]_  = \new_[103898]_  & \new_[103895]_ ;
  assign \new_[103902]_  = ~A201 & ~A200;
  assign \new_[103905]_  = A203 & ~A202;
  assign \new_[103906]_  = \new_[103905]_  & \new_[103902]_ ;
  assign \new_[103907]_  = \new_[103906]_  & \new_[103899]_ ;
  assign \new_[103910]_  = A266 & ~A265;
  assign \new_[103913]_  = ~A269 & A267;
  assign \new_[103914]_  = \new_[103913]_  & \new_[103910]_ ;
  assign \new_[103917]_  = A299 & ~A298;
  assign \new_[103921]_  = A302 & ~A301;
  assign \new_[103922]_  = ~A300 & \new_[103921]_ ;
  assign \new_[103923]_  = \new_[103922]_  & \new_[103917]_ ;
  assign \new_[103924]_  = \new_[103923]_  & \new_[103914]_ ;
  assign \new_[103927]_  = ~A169 & ~A170;
  assign \new_[103930]_  = A199 & A168;
  assign \new_[103931]_  = \new_[103930]_  & \new_[103927]_ ;
  assign \new_[103934]_  = ~A201 & ~A200;
  assign \new_[103937]_  = A203 & ~A202;
  assign \new_[103938]_  = \new_[103937]_  & \new_[103934]_ ;
  assign \new_[103939]_  = \new_[103938]_  & \new_[103931]_ ;
  assign \new_[103942]_  = A266 & ~A265;
  assign \new_[103945]_  = ~A268 & ~A267;
  assign \new_[103946]_  = \new_[103945]_  & \new_[103942]_ ;
  assign \new_[103949]_  = A298 & A269;
  assign \new_[103953]_  = A301 & A300;
  assign \new_[103954]_  = ~A299 & \new_[103953]_ ;
  assign \new_[103955]_  = \new_[103954]_  & \new_[103949]_ ;
  assign \new_[103956]_  = \new_[103955]_  & \new_[103946]_ ;
  assign \new_[103959]_  = ~A169 & ~A170;
  assign \new_[103962]_  = A199 & A168;
  assign \new_[103963]_  = \new_[103962]_  & \new_[103959]_ ;
  assign \new_[103966]_  = ~A201 & ~A200;
  assign \new_[103969]_  = A203 & ~A202;
  assign \new_[103970]_  = \new_[103969]_  & \new_[103966]_ ;
  assign \new_[103971]_  = \new_[103970]_  & \new_[103963]_ ;
  assign \new_[103974]_  = A266 & ~A265;
  assign \new_[103977]_  = ~A268 & ~A267;
  assign \new_[103978]_  = \new_[103977]_  & \new_[103974]_ ;
  assign \new_[103981]_  = A298 & A269;
  assign \new_[103985]_  = ~A302 & A300;
  assign \new_[103986]_  = ~A299 & \new_[103985]_ ;
  assign \new_[103987]_  = \new_[103986]_  & \new_[103981]_ ;
  assign \new_[103988]_  = \new_[103987]_  & \new_[103978]_ ;
  assign \new_[103991]_  = ~A169 & ~A170;
  assign \new_[103994]_  = A199 & A168;
  assign \new_[103995]_  = \new_[103994]_  & \new_[103991]_ ;
  assign \new_[103998]_  = ~A201 & ~A200;
  assign \new_[104001]_  = A203 & ~A202;
  assign \new_[104002]_  = \new_[104001]_  & \new_[103998]_ ;
  assign \new_[104003]_  = \new_[104002]_  & \new_[103995]_ ;
  assign \new_[104006]_  = A266 & ~A265;
  assign \new_[104009]_  = ~A268 & ~A267;
  assign \new_[104010]_  = \new_[104009]_  & \new_[104006]_ ;
  assign \new_[104013]_  = ~A298 & A269;
  assign \new_[104017]_  = A301 & A300;
  assign \new_[104018]_  = A299 & \new_[104017]_ ;
  assign \new_[104019]_  = \new_[104018]_  & \new_[104013]_ ;
  assign \new_[104020]_  = \new_[104019]_  & \new_[104010]_ ;
  assign \new_[104023]_  = ~A169 & ~A170;
  assign \new_[104026]_  = A199 & A168;
  assign \new_[104027]_  = \new_[104026]_  & \new_[104023]_ ;
  assign \new_[104030]_  = ~A201 & ~A200;
  assign \new_[104033]_  = A203 & ~A202;
  assign \new_[104034]_  = \new_[104033]_  & \new_[104030]_ ;
  assign \new_[104035]_  = \new_[104034]_  & \new_[104027]_ ;
  assign \new_[104038]_  = A266 & ~A265;
  assign \new_[104041]_  = ~A268 & ~A267;
  assign \new_[104042]_  = \new_[104041]_  & \new_[104038]_ ;
  assign \new_[104045]_  = ~A298 & A269;
  assign \new_[104049]_  = ~A302 & A300;
  assign \new_[104050]_  = A299 & \new_[104049]_ ;
  assign \new_[104051]_  = \new_[104050]_  & \new_[104045]_ ;
  assign \new_[104052]_  = \new_[104051]_  & \new_[104042]_ ;
  assign \new_[104055]_  = ~A169 & ~A170;
  assign \new_[104058]_  = A199 & A168;
  assign \new_[104059]_  = \new_[104058]_  & \new_[104055]_ ;
  assign \new_[104062]_  = ~A201 & ~A200;
  assign \new_[104065]_  = A203 & ~A202;
  assign \new_[104066]_  = \new_[104065]_  & \new_[104062]_ ;
  assign \new_[104067]_  = \new_[104066]_  & \new_[104059]_ ;
  assign \new_[104070]_  = ~A266 & A265;
  assign \new_[104073]_  = A268 & A267;
  assign \new_[104074]_  = \new_[104073]_  & \new_[104070]_ ;
  assign \new_[104077]_  = ~A299 & A298;
  assign \new_[104081]_  = A302 & ~A301;
  assign \new_[104082]_  = ~A300 & \new_[104081]_ ;
  assign \new_[104083]_  = \new_[104082]_  & \new_[104077]_ ;
  assign \new_[104084]_  = \new_[104083]_  & \new_[104074]_ ;
  assign \new_[104087]_  = ~A169 & ~A170;
  assign \new_[104090]_  = A199 & A168;
  assign \new_[104091]_  = \new_[104090]_  & \new_[104087]_ ;
  assign \new_[104094]_  = ~A201 & ~A200;
  assign \new_[104097]_  = A203 & ~A202;
  assign \new_[104098]_  = \new_[104097]_  & \new_[104094]_ ;
  assign \new_[104099]_  = \new_[104098]_  & \new_[104091]_ ;
  assign \new_[104102]_  = ~A266 & A265;
  assign \new_[104105]_  = A268 & A267;
  assign \new_[104106]_  = \new_[104105]_  & \new_[104102]_ ;
  assign \new_[104109]_  = A299 & ~A298;
  assign \new_[104113]_  = A302 & ~A301;
  assign \new_[104114]_  = ~A300 & \new_[104113]_ ;
  assign \new_[104115]_  = \new_[104114]_  & \new_[104109]_ ;
  assign \new_[104116]_  = \new_[104115]_  & \new_[104106]_ ;
  assign \new_[104119]_  = ~A169 & ~A170;
  assign \new_[104122]_  = A199 & A168;
  assign \new_[104123]_  = \new_[104122]_  & \new_[104119]_ ;
  assign \new_[104126]_  = ~A201 & ~A200;
  assign \new_[104129]_  = A203 & ~A202;
  assign \new_[104130]_  = \new_[104129]_  & \new_[104126]_ ;
  assign \new_[104131]_  = \new_[104130]_  & \new_[104123]_ ;
  assign \new_[104134]_  = ~A266 & A265;
  assign \new_[104137]_  = ~A269 & A267;
  assign \new_[104138]_  = \new_[104137]_  & \new_[104134]_ ;
  assign \new_[104141]_  = ~A299 & A298;
  assign \new_[104145]_  = A302 & ~A301;
  assign \new_[104146]_  = ~A300 & \new_[104145]_ ;
  assign \new_[104147]_  = \new_[104146]_  & \new_[104141]_ ;
  assign \new_[104148]_  = \new_[104147]_  & \new_[104138]_ ;
  assign \new_[104151]_  = ~A169 & ~A170;
  assign \new_[104154]_  = A199 & A168;
  assign \new_[104155]_  = \new_[104154]_  & \new_[104151]_ ;
  assign \new_[104158]_  = ~A201 & ~A200;
  assign \new_[104161]_  = A203 & ~A202;
  assign \new_[104162]_  = \new_[104161]_  & \new_[104158]_ ;
  assign \new_[104163]_  = \new_[104162]_  & \new_[104155]_ ;
  assign \new_[104166]_  = ~A266 & A265;
  assign \new_[104169]_  = ~A269 & A267;
  assign \new_[104170]_  = \new_[104169]_  & \new_[104166]_ ;
  assign \new_[104173]_  = A299 & ~A298;
  assign \new_[104177]_  = A302 & ~A301;
  assign \new_[104178]_  = ~A300 & \new_[104177]_ ;
  assign \new_[104179]_  = \new_[104178]_  & \new_[104173]_ ;
  assign \new_[104180]_  = \new_[104179]_  & \new_[104170]_ ;
  assign \new_[104183]_  = ~A169 & ~A170;
  assign \new_[104186]_  = A199 & A168;
  assign \new_[104187]_  = \new_[104186]_  & \new_[104183]_ ;
  assign \new_[104190]_  = ~A201 & ~A200;
  assign \new_[104193]_  = A203 & ~A202;
  assign \new_[104194]_  = \new_[104193]_  & \new_[104190]_ ;
  assign \new_[104195]_  = \new_[104194]_  & \new_[104187]_ ;
  assign \new_[104198]_  = ~A266 & A265;
  assign \new_[104201]_  = ~A268 & ~A267;
  assign \new_[104202]_  = \new_[104201]_  & \new_[104198]_ ;
  assign \new_[104205]_  = A298 & A269;
  assign \new_[104209]_  = A301 & A300;
  assign \new_[104210]_  = ~A299 & \new_[104209]_ ;
  assign \new_[104211]_  = \new_[104210]_  & \new_[104205]_ ;
  assign \new_[104212]_  = \new_[104211]_  & \new_[104202]_ ;
  assign \new_[104215]_  = ~A169 & ~A170;
  assign \new_[104218]_  = A199 & A168;
  assign \new_[104219]_  = \new_[104218]_  & \new_[104215]_ ;
  assign \new_[104222]_  = ~A201 & ~A200;
  assign \new_[104225]_  = A203 & ~A202;
  assign \new_[104226]_  = \new_[104225]_  & \new_[104222]_ ;
  assign \new_[104227]_  = \new_[104226]_  & \new_[104219]_ ;
  assign \new_[104230]_  = ~A266 & A265;
  assign \new_[104233]_  = ~A268 & ~A267;
  assign \new_[104234]_  = \new_[104233]_  & \new_[104230]_ ;
  assign \new_[104237]_  = A298 & A269;
  assign \new_[104241]_  = ~A302 & A300;
  assign \new_[104242]_  = ~A299 & \new_[104241]_ ;
  assign \new_[104243]_  = \new_[104242]_  & \new_[104237]_ ;
  assign \new_[104244]_  = \new_[104243]_  & \new_[104234]_ ;
  assign \new_[104247]_  = ~A169 & ~A170;
  assign \new_[104250]_  = A199 & A168;
  assign \new_[104251]_  = \new_[104250]_  & \new_[104247]_ ;
  assign \new_[104254]_  = ~A201 & ~A200;
  assign \new_[104257]_  = A203 & ~A202;
  assign \new_[104258]_  = \new_[104257]_  & \new_[104254]_ ;
  assign \new_[104259]_  = \new_[104258]_  & \new_[104251]_ ;
  assign \new_[104262]_  = ~A266 & A265;
  assign \new_[104265]_  = ~A268 & ~A267;
  assign \new_[104266]_  = \new_[104265]_  & \new_[104262]_ ;
  assign \new_[104269]_  = ~A298 & A269;
  assign \new_[104273]_  = A301 & A300;
  assign \new_[104274]_  = A299 & \new_[104273]_ ;
  assign \new_[104275]_  = \new_[104274]_  & \new_[104269]_ ;
  assign \new_[104276]_  = \new_[104275]_  & \new_[104266]_ ;
  assign \new_[104279]_  = ~A169 & ~A170;
  assign \new_[104282]_  = A199 & A168;
  assign \new_[104283]_  = \new_[104282]_  & \new_[104279]_ ;
  assign \new_[104286]_  = ~A201 & ~A200;
  assign \new_[104289]_  = A203 & ~A202;
  assign \new_[104290]_  = \new_[104289]_  & \new_[104286]_ ;
  assign \new_[104291]_  = \new_[104290]_  & \new_[104283]_ ;
  assign \new_[104294]_  = ~A266 & A265;
  assign \new_[104297]_  = ~A268 & ~A267;
  assign \new_[104298]_  = \new_[104297]_  & \new_[104294]_ ;
  assign \new_[104301]_  = ~A298 & A269;
  assign \new_[104305]_  = ~A302 & A300;
  assign \new_[104306]_  = A299 & \new_[104305]_ ;
  assign \new_[104307]_  = \new_[104306]_  & \new_[104301]_ ;
  assign \new_[104308]_  = \new_[104307]_  & \new_[104298]_ ;
  assign \new_[104311]_  = ~A169 & ~A170;
  assign \new_[104314]_  = ~A199 & A168;
  assign \new_[104315]_  = \new_[104314]_  & \new_[104311]_ ;
  assign \new_[104318]_  = ~A201 & A200;
  assign \new_[104322]_  = ~A265 & A203;
  assign \new_[104323]_  = ~A202 & \new_[104322]_ ;
  assign \new_[104324]_  = \new_[104323]_  & \new_[104318]_ ;
  assign \new_[104325]_  = \new_[104324]_  & \new_[104315]_ ;
  assign \new_[104328]_  = ~A267 & A266;
  assign \new_[104331]_  = A269 & ~A268;
  assign \new_[104332]_  = \new_[104331]_  & \new_[104328]_ ;
  assign \new_[104335]_  = ~A299 & A298;
  assign \new_[104339]_  = A302 & ~A301;
  assign \new_[104340]_  = ~A300 & \new_[104339]_ ;
  assign \new_[104341]_  = \new_[104340]_  & \new_[104335]_ ;
  assign \new_[104342]_  = \new_[104341]_  & \new_[104332]_ ;
  assign \new_[104345]_  = ~A169 & ~A170;
  assign \new_[104348]_  = ~A199 & A168;
  assign \new_[104349]_  = \new_[104348]_  & \new_[104345]_ ;
  assign \new_[104352]_  = ~A201 & A200;
  assign \new_[104356]_  = ~A265 & A203;
  assign \new_[104357]_  = ~A202 & \new_[104356]_ ;
  assign \new_[104358]_  = \new_[104357]_  & \new_[104352]_ ;
  assign \new_[104359]_  = \new_[104358]_  & \new_[104349]_ ;
  assign \new_[104362]_  = ~A267 & A266;
  assign \new_[104365]_  = A269 & ~A268;
  assign \new_[104366]_  = \new_[104365]_  & \new_[104362]_ ;
  assign \new_[104369]_  = A299 & ~A298;
  assign \new_[104373]_  = A302 & ~A301;
  assign \new_[104374]_  = ~A300 & \new_[104373]_ ;
  assign \new_[104375]_  = \new_[104374]_  & \new_[104369]_ ;
  assign \new_[104376]_  = \new_[104375]_  & \new_[104366]_ ;
  assign \new_[104379]_  = ~A169 & ~A170;
  assign \new_[104382]_  = ~A199 & A168;
  assign \new_[104383]_  = \new_[104382]_  & \new_[104379]_ ;
  assign \new_[104386]_  = ~A201 & A200;
  assign \new_[104390]_  = A265 & A203;
  assign \new_[104391]_  = ~A202 & \new_[104390]_ ;
  assign \new_[104392]_  = \new_[104391]_  & \new_[104386]_ ;
  assign \new_[104393]_  = \new_[104392]_  & \new_[104383]_ ;
  assign \new_[104396]_  = ~A267 & ~A266;
  assign \new_[104399]_  = A269 & ~A268;
  assign \new_[104400]_  = \new_[104399]_  & \new_[104396]_ ;
  assign \new_[104403]_  = ~A299 & A298;
  assign \new_[104407]_  = A302 & ~A301;
  assign \new_[104408]_  = ~A300 & \new_[104407]_ ;
  assign \new_[104409]_  = \new_[104408]_  & \new_[104403]_ ;
  assign \new_[104410]_  = \new_[104409]_  & \new_[104400]_ ;
  assign \new_[104413]_  = ~A169 & ~A170;
  assign \new_[104416]_  = ~A199 & A168;
  assign \new_[104417]_  = \new_[104416]_  & \new_[104413]_ ;
  assign \new_[104420]_  = ~A201 & A200;
  assign \new_[104424]_  = A265 & A203;
  assign \new_[104425]_  = ~A202 & \new_[104424]_ ;
  assign \new_[104426]_  = \new_[104425]_  & \new_[104420]_ ;
  assign \new_[104427]_  = \new_[104426]_  & \new_[104417]_ ;
  assign \new_[104430]_  = ~A267 & ~A266;
  assign \new_[104433]_  = A269 & ~A268;
  assign \new_[104434]_  = \new_[104433]_  & \new_[104430]_ ;
  assign \new_[104437]_  = A299 & ~A298;
  assign \new_[104441]_  = A302 & ~A301;
  assign \new_[104442]_  = ~A300 & \new_[104441]_ ;
  assign \new_[104443]_  = \new_[104442]_  & \new_[104437]_ ;
  assign \new_[104444]_  = \new_[104443]_  & \new_[104434]_ ;
  assign \new_[104447]_  = ~A169 & ~A170;
  assign \new_[104450]_  = A199 & A168;
  assign \new_[104451]_  = \new_[104450]_  & \new_[104447]_ ;
  assign \new_[104454]_  = ~A201 & ~A200;
  assign \new_[104458]_  = ~A265 & A203;
  assign \new_[104459]_  = ~A202 & \new_[104458]_ ;
  assign \new_[104460]_  = \new_[104459]_  & \new_[104454]_ ;
  assign \new_[104461]_  = \new_[104460]_  & \new_[104451]_ ;
  assign \new_[104464]_  = ~A267 & A266;
  assign \new_[104467]_  = A269 & ~A268;
  assign \new_[104468]_  = \new_[104467]_  & \new_[104464]_ ;
  assign \new_[104471]_  = ~A299 & A298;
  assign \new_[104475]_  = A302 & ~A301;
  assign \new_[104476]_  = ~A300 & \new_[104475]_ ;
  assign \new_[104477]_  = \new_[104476]_  & \new_[104471]_ ;
  assign \new_[104478]_  = \new_[104477]_  & \new_[104468]_ ;
  assign \new_[104481]_  = ~A169 & ~A170;
  assign \new_[104484]_  = A199 & A168;
  assign \new_[104485]_  = \new_[104484]_  & \new_[104481]_ ;
  assign \new_[104488]_  = ~A201 & ~A200;
  assign \new_[104492]_  = ~A265 & A203;
  assign \new_[104493]_  = ~A202 & \new_[104492]_ ;
  assign \new_[104494]_  = \new_[104493]_  & \new_[104488]_ ;
  assign \new_[104495]_  = \new_[104494]_  & \new_[104485]_ ;
  assign \new_[104498]_  = ~A267 & A266;
  assign \new_[104501]_  = A269 & ~A268;
  assign \new_[104502]_  = \new_[104501]_  & \new_[104498]_ ;
  assign \new_[104505]_  = A299 & ~A298;
  assign \new_[104509]_  = A302 & ~A301;
  assign \new_[104510]_  = ~A300 & \new_[104509]_ ;
  assign \new_[104511]_  = \new_[104510]_  & \new_[104505]_ ;
  assign \new_[104512]_  = \new_[104511]_  & \new_[104502]_ ;
  assign \new_[104515]_  = ~A169 & ~A170;
  assign \new_[104518]_  = A199 & A168;
  assign \new_[104519]_  = \new_[104518]_  & \new_[104515]_ ;
  assign \new_[104522]_  = ~A201 & ~A200;
  assign \new_[104526]_  = A265 & A203;
  assign \new_[104527]_  = ~A202 & \new_[104526]_ ;
  assign \new_[104528]_  = \new_[104527]_  & \new_[104522]_ ;
  assign \new_[104529]_  = \new_[104528]_  & \new_[104519]_ ;
  assign \new_[104532]_  = ~A267 & ~A266;
  assign \new_[104535]_  = A269 & ~A268;
  assign \new_[104536]_  = \new_[104535]_  & \new_[104532]_ ;
  assign \new_[104539]_  = ~A299 & A298;
  assign \new_[104543]_  = A302 & ~A301;
  assign \new_[104544]_  = ~A300 & \new_[104543]_ ;
  assign \new_[104545]_  = \new_[104544]_  & \new_[104539]_ ;
  assign \new_[104546]_  = \new_[104545]_  & \new_[104536]_ ;
  assign \new_[104549]_  = ~A169 & ~A170;
  assign \new_[104552]_  = A199 & A168;
  assign \new_[104553]_  = \new_[104552]_  & \new_[104549]_ ;
  assign \new_[104556]_  = ~A201 & ~A200;
  assign \new_[104560]_  = A265 & A203;
  assign \new_[104561]_  = ~A202 & \new_[104560]_ ;
  assign \new_[104562]_  = \new_[104561]_  & \new_[104556]_ ;
  assign \new_[104563]_  = \new_[104562]_  & \new_[104553]_ ;
  assign \new_[104566]_  = ~A267 & ~A266;
  assign \new_[104569]_  = A269 & ~A268;
  assign \new_[104570]_  = \new_[104569]_  & \new_[104566]_ ;
  assign \new_[104573]_  = A299 & ~A298;
  assign \new_[104577]_  = A302 & ~A301;
  assign \new_[104578]_  = ~A300 & \new_[104577]_ ;
  assign \new_[104579]_  = \new_[104578]_  & \new_[104573]_ ;
  assign \new_[104580]_  = \new_[104579]_  & \new_[104570]_ ;
endmodule


