module top ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, a0, q, b0, r, c0, s,
    d0, t, e0, u, f0, v, g0, w, h0, x, i0, y, j0, z, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, c1, b1, e1, d1, g1, f1,
    i1, h1, j1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, a0, q, b0, r,
    c0, s, d0, t, e0, u, f0, v, g0, w, h0, x, i0, y, j0, z, k0, l0, m0, n0,
    o0;
  output p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, c1, b1, e1, d1, g1,
    f1, i1, h1, j1;
  wire new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n78_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n105_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n120_, new_n121_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n171_, new_n172_, new_n174_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_;
  assign new_n63_ = c0 & j0;
  assign new_n64_ = ~l0 & ~new_n63_;
  assign new_n65_ = b0 & ~new_n64_;
  assign new_n66_ = ~n0 & ~new_n65_;
  assign new_n67_ = c0 & ~k0;
  assign new_n68_ = ~j0 & ~k0;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = ~e & new_n69_;
  assign new_n71_ = ~e & k;
  assign new_n72_ = ~new_n70_ & ~new_n71_;
  assign new_n73_ = ~b0 & ~new_n71_;
  assign new_n74_ = ~new_n72_ & ~new_n73_;
  assign new_n75_ = o0 & new_n74_;
  assign new_n76_ = ~new_n65_ & ~new_n75_;
  assign b1 = new_n66_ | new_n76_;
  assign new_n78_ = ~p & ~b1;
  assign p0 = ~q | new_n78_;
  assign new_n80_ = e & j0;
  assign new_n81_ = b0 & ~c0;
  assign new_n82_ = new_n80_ & new_n81_;
  assign new_n83_ = ~e0 & ~g0;
  assign new_n84_ = e & ~new_n83_;
  assign new_n85_ = b0 & k0;
  assign new_n86_ = e & new_n85_;
  assign new_n87_ = ~new_n82_ & ~new_n84_;
  assign q0 = ~new_n86_ & new_n87_;
  assign new_n89_ = ~c0 & j0;
  assign new_n90_ = b0 & new_n89_;
  assign new_n91_ = i & new_n89_;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign new_n93_ = e & new_n92_;
  assign new_n94_ = i & d0;
  assign new_n95_ = ~c & ~new_n94_;
  assign new_n96_ = ~new_n93_ & ~new_n95_;
  assign x0 = n0 & o0;
  assign r0 = ~new_n96_ | ~x0;
  assign new_n99_ = ~b0 & ~l0;
  assign new_n100_ = b0 & ~new_n63_;
  assign new_n101_ = ~new_n64_ & ~new_n99_;
  assign new_n102_ = ~new_n100_ & new_n101_;
  assign s0 = ~v | ~new_n102_;
  assign t0 = v | ~new_n102_;
  assign new_n105_ = b0 & c0;
  assign v0 = ~l0 & ~new_n105_;
  assign new_n107_ = ~p & r;
  assign new_n108_ = ~f0 & ~h0;
  assign new_n109_ = ~new_n107_ & new_n108_;
  assign new_n110_ = o & ~new_n109_;
  assign new_n111_ = d & ~new_n110_;
  assign new_n112_ = ~m0 & new_n111_;
  assign new_n113_ = ~a & o;
  assign new_n114_ = o & z;
  assign new_n115_ = ~a & ~z;
  assign new_n116_ = ~new_n113_ & ~new_n114_;
  assign new_n117_ = ~new_n115_ & new_n116_;
  assign new_n118_ = new_n111_ & new_n117_;
  assign w0 = new_n112_ | new_n118_;
  assign new_n120_ = a0 & i0;
  assign new_n121_ = b0 & new_n120_;
  assign y0 = l & new_n121_;
  assign new_n123_ = o0 & ~new_n83_;
  assign new_n124_ = o0 & new_n69_;
  assign new_n125_ = b0 & new_n124_;
  assign new_n126_ = ~new_n123_ & ~new_n125_;
  assign new_n127_ = n0 & ~new_n126_;
  assign new_n128_ = ~e & f;
  assign new_n129_ = new_n127_ & new_n128_;
  assign new_n130_ = h & b0;
  assign new_n131_ = new_n70_ & new_n130_;
  assign new_n132_ = ~n0 & new_n131_;
  assign new_n133_ = ~o0 & new_n131_;
  assign new_n134_ = ~new_n132_ & ~new_n133_;
  assign new_n135_ = g & l0;
  assign new_n136_ = b0 & new_n135_;
  assign new_n137_ = ~new_n129_ & new_n134_;
  assign z0 = new_n136_ | ~new_n137_;
  assign new_n139_ = o0 & new_n94_;
  assign new_n140_ = b0 & j0;
  assign new_n141_ = ~e & ~c0;
  assign new_n142_ = new_n140_ & new_n141_;
  assign new_n143_ = i & ~c0;
  assign new_n144_ = j0 & new_n143_;
  assign new_n145_ = ~b0 & new_n144_;
  assign new_n146_ = ~j & ~e0;
  assign new_n147_ = ~new_n142_ & ~new_n145_;
  assign new_n148_ = new_n146_ & new_n147_;
  assign new_n149_ = ~new_n139_ & new_n148_;
  assign new_n150_ = ~n0 & new_n148_;
  assign h1 = ~new_n149_ & ~new_n150_;
  assign new_n152_ = ~e & o0;
  assign new_n153_ = j0 & k0;
  assign new_n154_ = c0 & ~new_n153_;
  assign new_n155_ = new_n83_ & new_n154_;
  assign new_n156_ = ~b0 & new_n83_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = new_n152_ & new_n157_;
  assign new_n159_ = ~n & new_n158_;
  assign new_n160_ = ~j0 & ~l0;
  assign new_n161_ = ~c0 & ~l0;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign new_n163_ = ~s & u;
  assign new_n164_ = ~t & new_n163_;
  assign new_n165_ = new_n162_ & new_n164_;
  assign new_n166_ = b0 & new_n165_;
  assign new_n167_ = ~new_n159_ & ~new_n166_;
  assign new_n168_ = ~n0 & ~new_n166_;
  assign c1 = ~new_n167_ & ~new_n168_;
  assign e1 = m & new_n121_;
  assign new_n171_ = w & ~y;
  assign new_n172_ = b & x;
  assign g1 = new_n171_ & new_n172_;
  assign new_n174_ = b & w;
  assign f1 = ~x & new_n174_;
  assign new_n176_ = i & j0;
  assign new_n177_ = ~c0 & new_n176_;
  assign new_n178_ = ~e0 & ~new_n140_;
  assign new_n179_ = ~j & ~new_n177_;
  assign new_n180_ = new_n178_ & new_n179_;
  assign new_n181_ = ~new_n139_ & new_n180_;
  assign new_n182_ = ~n0 & new_n180_;
  assign j1 = new_n181_ | new_n182_;
  assign u0 = ~v0;
  assign a1 = ~h1;
  assign d1 = ~c1;
  assign i1 = a1;
endmodule

