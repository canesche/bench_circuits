module MultiplierB_16 ( clock, 
    \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    50  );
  input  clock;
  input  \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18;
  output 50;
  reg 2, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48;
  wire new_n109_, new_n110_, new_n111_, new_n112_, new_n113_1_, new_n114_,
    new_n117_, new_n118_1_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_1_, new_n129_,
    new_n131_, new_n132_, new_n133_1_, new_n134_, new_n135_, new_n136_,
    new_n138_1_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_1_,
    new_n145_, new_n146_, new_n147_, new_n148_1_, new_n149_, new_n150_,
    new_n152_, new_n153_1_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_1_, new_n164_,
    new_n166_, new_n167_, new_n168_1_, new_n169_, new_n170_, new_n171_,
    new_n173_1_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_1_,
    new_n180_, new_n181_, new_n182_, new_n183_1_, new_n184_, new_n185_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n285_, new_n286_, new_n287_, new_n288_, n38,
    n43, n48, n53, n58, n63, n68, n73, n78, n83, n88, n93, n98, n103, n108,
    n113, n118, n123, n128, n133, n138, n143, n148, n153, n158, n163, n168,
    n173, n178, n183;
  assign new_n109_ = \1  & 3;
  assign new_n110_ = ~20 & 34;
  assign new_n111_ = 20 & ~34;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign new_n113_1_ = new_n109_ & new_n112_;
  assign new_n114_ = ~new_n109_ & ~new_n112_;
  assign 50 = new_n113_1_ | new_n114_;
  assign n38 = \1  & 18;
  assign new_n117_ = \1  & 4;
  assign new_n118_1_ = ~21 & 35;
  assign new_n119_ = 21 & ~35;
  assign new_n120_ = ~new_n118_1_ & ~new_n119_;
  assign new_n121_ = new_n117_ & new_n120_;
  assign new_n122_ = ~new_n117_ & ~new_n120_;
  assign n43 = new_n121_ | new_n122_;
  assign new_n124_ = \1  & 5;
  assign new_n125_ = ~22 & 36;
  assign new_n126_ = 22 & ~36;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_1_ = new_n124_ & new_n127_;
  assign new_n129_ = ~new_n124_ & ~new_n127_;
  assign n48 = new_n128_1_ | new_n129_;
  assign new_n131_ = \1  & 6;
  assign new_n132_ = ~23 & 37;
  assign new_n133_1_ = 23 & ~37;
  assign new_n134_ = ~new_n132_ & ~new_n133_1_;
  assign new_n135_ = new_n131_ & new_n134_;
  assign new_n136_ = ~new_n131_ & ~new_n134_;
  assign n53 = new_n135_ | new_n136_;
  assign new_n138_1_ = \1  & 7;
  assign new_n139_ = ~24 & 38;
  assign new_n140_ = 24 & ~38;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = new_n138_1_ & new_n141_;
  assign new_n143_1_ = ~new_n138_1_ & ~new_n141_;
  assign n58 = new_n142_ | new_n143_1_;
  assign new_n145_ = \1  & 8;
  assign new_n146_ = ~25 & 39;
  assign new_n147_ = 25 & ~39;
  assign new_n148_1_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = new_n145_ & new_n148_1_;
  assign new_n150_ = ~new_n145_ & ~new_n148_1_;
  assign n63 = new_n149_ | new_n150_;
  assign new_n152_ = \1  & 9;
  assign new_n153_1_ = ~26 & 40;
  assign new_n154_ = 26 & ~40;
  assign new_n155_ = ~new_n153_1_ & ~new_n154_;
  assign new_n156_ = new_n152_ & new_n155_;
  assign new_n157_ = ~new_n152_ & ~new_n155_;
  assign n68 = new_n156_ | new_n157_;
  assign new_n159_ = \1  & 10;
  assign new_n160_ = ~27 & 41;
  assign new_n161_ = 27 & ~41;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign new_n163_1_ = new_n159_ & new_n162_;
  assign new_n164_ = ~new_n159_ & ~new_n162_;
  assign n73 = new_n163_1_ | new_n164_;
  assign new_n166_ = \1  & 11;
  assign new_n167_ = ~28 & 42;
  assign new_n168_1_ = 28 & ~42;
  assign new_n169_ = ~new_n167_ & ~new_n168_1_;
  assign new_n170_ = new_n166_ & new_n169_;
  assign new_n171_ = ~new_n166_ & ~new_n169_;
  assign n78 = new_n170_ | new_n171_;
  assign new_n173_1_ = \1  & 12;
  assign new_n174_ = ~29 & 43;
  assign new_n175_ = 29 & ~43;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = new_n173_1_ & new_n176_;
  assign new_n178_1_ = ~new_n173_1_ & ~new_n176_;
  assign n83 = new_n177_ | new_n178_1_;
  assign new_n180_ = \1  & 13;
  assign new_n181_ = ~30 & 44;
  assign new_n182_ = 30 & ~44;
  assign new_n183_1_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = new_n180_ & new_n183_1_;
  assign new_n185_ = ~new_n180_ & ~new_n183_1_;
  assign n88 = new_n184_ | new_n185_;
  assign new_n187_ = \1  & 14;
  assign new_n188_ = ~31 & 45;
  assign new_n189_ = 31 & ~45;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = new_n187_ & new_n190_;
  assign new_n192_ = ~new_n187_ & ~new_n190_;
  assign n93 = new_n191_ | new_n192_;
  assign new_n194_ = \1  & 15;
  assign new_n195_ = ~32 & 46;
  assign new_n196_ = 32 & ~46;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = new_n194_ & new_n197_;
  assign new_n199_ = ~new_n194_ & ~new_n197_;
  assign n98 = new_n198_ | new_n199_;
  assign new_n201_ = \1  & 16;
  assign new_n202_ = ~33 & 47;
  assign new_n203_ = 33 & ~47;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = new_n201_ & new_n204_;
  assign new_n206_ = ~new_n201_ & ~new_n204_;
  assign n103 = new_n205_ | new_n206_;
  assign new_n208_ = \1  & 17;
  assign new_n209_ = ~2 & 48;
  assign new_n210_ = 2 & ~48;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = new_n208_ & new_n211_;
  assign new_n213_ = ~new_n208_ & ~new_n211_;
  assign n108 = new_n212_ | new_n213_;
  assign new_n215_ = 20 & 34;
  assign new_n216_ = 20 & new_n109_;
  assign new_n217_ = 34 & new_n109_;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign n113 = new_n215_ | ~new_n218_;
  assign new_n220_ = 21 & 35;
  assign new_n221_ = 21 & new_n117_;
  assign new_n222_ = 35 & new_n117_;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign n118 = new_n220_ | ~new_n223_;
  assign new_n225_ = 22 & 36;
  assign new_n226_ = 22 & new_n124_;
  assign new_n227_ = 36 & new_n124_;
  assign new_n228_ = ~new_n226_ & ~new_n227_;
  assign n123 = new_n225_ | ~new_n228_;
  assign new_n230_ = 23 & 37;
  assign new_n231_ = 23 & new_n131_;
  assign new_n232_ = 37 & new_n131_;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign n128 = new_n230_ | ~new_n233_;
  assign new_n235_ = 24 & 38;
  assign new_n236_ = 24 & new_n138_1_;
  assign new_n237_ = 38 & new_n138_1_;
  assign new_n238_ = ~new_n236_ & ~new_n237_;
  assign n133 = new_n235_ | ~new_n238_;
  assign new_n240_ = 25 & 39;
  assign new_n241_ = 25 & new_n145_;
  assign new_n242_ = 39 & new_n145_;
  assign new_n243_ = ~new_n241_ & ~new_n242_;
  assign n138 = new_n240_ | ~new_n243_;
  assign new_n245_ = 26 & 40;
  assign new_n246_ = 26 & new_n152_;
  assign new_n247_ = 40 & new_n152_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign n143 = new_n245_ | ~new_n248_;
  assign new_n250_ = 27 & 41;
  assign new_n251_ = 27 & new_n159_;
  assign new_n252_ = 41 & new_n159_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign n148 = new_n250_ | ~new_n253_;
  assign new_n255_ = 28 & 42;
  assign new_n256_ = 28 & new_n166_;
  assign new_n257_ = 42 & new_n166_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign n153 = new_n255_ | ~new_n258_;
  assign new_n260_ = 29 & 43;
  assign new_n261_ = 29 & new_n173_1_;
  assign new_n262_ = 43 & new_n173_1_;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign n158 = new_n260_ | ~new_n263_;
  assign new_n265_ = 30 & 44;
  assign new_n266_ = 30 & new_n180_;
  assign new_n267_ = 44 & new_n180_;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign n163 = new_n265_ | ~new_n268_;
  assign new_n270_ = 31 & 45;
  assign new_n271_ = 31 & new_n187_;
  assign new_n272_ = 45 & new_n187_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign n168 = new_n270_ | ~new_n273_;
  assign new_n275_ = 32 & 46;
  assign new_n276_ = 32 & new_n194_;
  assign new_n277_ = 46 & new_n194_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign n173 = new_n275_ | ~new_n278_;
  assign new_n280_ = 33 & 47;
  assign new_n281_ = 33 & new_n201_;
  assign new_n282_ = 47 & new_n201_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign n178 = new_n280_ | ~new_n283_;
  assign new_n285_ = 2 & 48;
  assign new_n286_ = 2 & new_n208_;
  assign new_n287_ = 48 & new_n208_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign n183 = new_n285_ | ~new_n288_;
  always @ (posedge clock) begin
    2 <= n38;
    20 <= n43;
    21 <= n48;
    22 <= n53;
    23 <= n58;
    24 <= n63;
    25 <= n68;
    26 <= n73;
    27 <= n78;
    28 <= n83;
    29 <= n88;
    30 <= n93;
    31 <= n98;
    32 <= n103;
    33 <= n108;
    34 <= n113;
    35 <= n118;
    36 <= n123;
    37 <= n128;
    38 <= n133;
    39 <= n138;
    40 <= n143;
    41 <= n148;
    42 <= n153;
    43 <= n158;
    44 <= n163;
    45 <= n168;
    46 <= n173;
    47 <= n178;
    48 <= n183;
  end
  initial begin
    2 <= 1'b0;
    20 <= 1'b0;
    21 <= 1'b0;
    22 <= 1'b0;
    23 <= 1'b0;
    24 <= 1'b0;
    25 <= 1'b0;
    26 <= 1'b0;
    27 <= 1'b0;
    28 <= 1'b0;
    29 <= 1'b0;
    30 <= 1'b0;
    31 <= 1'b0;
    32 <= 1'b0;
    33 <= 1'b0;
    34 <= 1'b0;
    35 <= 1'b0;
    36 <= 1'b0;
    37 <= 1'b0;
    38 <= 1'b0;
    39 <= 1'b0;
    40 <= 1'b0;
    41 <= 1'b0;
    42 <= 1'b0;
    43 <= 1'b0;
    44 <= 1'b0;
    45 <= 1'b0;
    46 <= 1'b0;
    47 <= 1'b0;
    48 <= 1'b0;
  end
endmodule

