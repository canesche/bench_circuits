module rot ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1,
    i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1,
    a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2,
    s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3,
    k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4,
    c4, d4, e4,
    f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4,
    x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5,
    p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6,
    h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6,
    z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7,
    r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1,
    g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1,
    y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2,
    q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3,
    i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3,
    a4, b4, c4, d4, e4;
  output f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4,
    w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5,
    o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6,
    g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6,
    y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7,
    q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8;
  wire new_n243_, new_n244_, new_n245_, new_n247_, new_n248_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n283_,
    new_n284_, new_n285_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n369_, new_n370_, new_n371_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n402_, new_n403_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n441_, new_n442_,
    new_n443_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n459_, new_n462_, new_n463_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n476_, new_n478_, new_n479_, new_n481_, new_n483_,
    new_n484_, new_n486_, new_n488_, new_n490_, new_n491_, new_n493_,
    new_n495_, new_n496_, new_n497_, new_n499_, new_n501_, new_n502_,
    new_n503_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n583_,
    new_n584_, new_n585_, new_n587_, new_n588_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n613_, new_n614_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n645_, new_n646_, new_n647_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n704_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n782_, new_n783_, new_n786_, new_n787_, new_n789_, new_n791_;
  assign new_n243_ = x & ~y;
  assign new_n244_ = e0 & ~new_n243_;
  assign new_n245_ = j1 & new_n243_;
  assign f4 = new_n244_ | new_n245_;
  assign new_n247_ = p0 & ~y1;
  assign new_n248_ = k1 & y1;
  assign g4 = new_n247_ | new_n248_;
  assign new_n250_ = x1 & m2;
  assign new_n251_ = y1 & new_n250_;
  assign new_n252_ = ~u & s0;
  assign new_n253_ = ~h0 & ~s0;
  assign new_n254_ = ~new_n252_ & ~new_n253_;
  assign new_n255_ = ~k & d0;
  assign new_n256_ = ~m & ~d0;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = x2 & ~new_n257_;
  assign new_n259_ = ~w2 & new_n258_;
  assign new_n260_ = ~h & u3;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = ~new_n254_ & ~new_n261_;
  assign new_n263_ = u2 & new_n262_;
  assign new_n264_ = ~i & u3;
  assign new_n265_ = g & ~new_n264_;
  assign new_n266_ = ~j & d0;
  assign new_n267_ = ~l & ~d0;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = new_n265_ & new_n268_;
  assign new_n270_ = ~new_n263_ & new_n269_;
  assign new_n271_ = x2 & ~new_n251_;
  assign new_n272_ = x2 & ~new_n270_;
  assign new_n273_ = w2 & ~new_n272_;
  assign d8 = new_n271_ | new_n273_;
  assign h4 = v2 | d8;
  assign new_n276_ = u & s0;
  assign new_n277_ = ~t & new_n276_;
  assign new_n278_ = h0 & ~s0;
  assign new_n279_ = ~g0 & new_n278_;
  assign new_n280_ = ~new_n277_ & ~new_n279_;
  assign new_n281_ = u2 & ~new_n280_;
  assign i4 = d8 | new_n281_;
  assign new_n283_ = ~new_n276_ & ~new_n278_;
  assign new_n284_ = u2 & ~new_n283_;
  assign new_n285_ = c2 & d8;
  assign j4 = new_n284_ | new_n285_;
  assign new_n287_ = p2 & q2;
  assign new_n288_ = m2 & ~new_n287_;
  assign new_n289_ = ~y1 & new_n288_;
  assign new_n290_ = x1 & new_n289_;
  assign new_n291_ = r0 & new_n290_;
  assign new_n292_ = ~x1 & y1;
  assign new_n293_ = m2 & new_n292_;
  assign new_n294_ = d1 & e1;
  assign new_n295_ = c1 & new_n294_;
  assign new_n296_ = n & ~new_n295_;
  assign new_n297_ = new_n293_ & ~new_n296_;
  assign new_n298_ = ~w1 & new_n251_;
  assign new_n299_ = ~new_n291_ & ~new_n298_;
  assign n4 = new_n297_ | ~new_n299_;
  assign o4 = w1 & new_n251_;
  assign new_n302_ = b2 & ~d8;
  assign new_n303_ = ~s1 & new_n302_;
  assign new_n304_ = s0 & ~new_n303_;
  assign new_n305_ = ~r1 & s1;
  assign new_n306_ = new_n302_ & new_n305_;
  assign new_n307_ = n1 & ~new_n306_;
  assign new_n308_ = f2 & ~h2;
  assign new_n309_ = ~f2 & h2;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~g2 & ~new_n310_;
  assign new_n312_ = ~f2 & ~h2;
  assign new_n313_ = r1 & ~s1;
  assign new_n314_ = ~new_n305_ & ~new_n313_;
  assign new_n315_ = l2 & new_n311_;
  assign new_n316_ = ~z1 & ~new_n315_;
  assign new_n317_ = ~new_n314_ & ~new_n316_;
  assign new_n318_ = ~new_n312_ & new_n317_;
  assign new_n319_ = o2 & new_n318_;
  assign new_n320_ = ~p1 & new_n319_;
  assign new_n321_ = r1 & new_n320_;
  assign new_n322_ = v1 & b2;
  assign new_n323_ = ~d8 & new_n322_;
  assign new_n324_ = ~i3 & m3;
  assign new_n325_ = h3 & new_n324_;
  assign new_n326_ = ~e3 & ~new_n325_;
  assign new_n327_ = ~new_n323_ & ~new_n326_;
  assign new_n328_ = i3 & m3;
  assign new_n329_ = ~h3 & new_n328_;
  assign new_n330_ = ~f3 & ~new_n329_;
  assign new_n331_ = ~new_n323_ & ~new_n330_;
  assign new_n332_ = ~new_n327_ & ~new_n331_;
  assign new_n333_ = g3 & ~new_n323_;
  assign new_n334_ = ~new_n321_ & new_n333_;
  assign new_n335_ = ~new_n332_ & new_n334_;
  assign new_n336_ = ~s & ~l3;
  assign new_n337_ = ~new_n304_ & ~new_n336_;
  assign new_n338_ = u2 & ~new_n337_;
  assign new_n339_ = y3 & ~new_n307_;
  assign new_n340_ = v2 & ~new_n339_;
  assign new_n341_ = y2 & ~new_n321_;
  assign new_n342_ = ~new_n332_ & new_n335_;
  assign new_n343_ = new_n341_ & new_n342_;
  assign new_n344_ = ~new_n340_ & ~new_n343_;
  assign new_n345_ = ~new_n338_ & new_n344_;
  assign new_n346_ = ~z3 & ~new_n345_;
  assign new_n347_ = ~d8 & new_n346_;
  assign new_n348_ = new_n251_ & new_n270_;
  assign new_n349_ = x2 & ~new_n348_;
  assign new_n350_ = w2 & ~new_n349_;
  assign new_n351_ = ~new_n347_ & ~new_n350_;
  assign new_n352_ = a & f0;
  assign new_n353_ = ~j4 & new_n320_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = r2 & new_n354_;
  assign new_n356_ = new_n351_ & ~new_n355_;
  assign new_n357_ = ~t1 & t2;
  assign new_n358_ = f2 & h2;
  assign new_n359_ = ~g2 & l2;
  assign new_n360_ = ~z1 & ~new_n359_;
  assign new_n361_ = ~new_n358_ & ~new_n360_;
  assign new_n362_ = g2 & l2;
  assign new_n363_ = z1 & ~new_n362_;
  assign new_n364_ = ~new_n312_ & ~new_n363_;
  assign new_n365_ = ~new_n361_ & new_n364_;
  assign new_n366_ = ~new_n357_ & ~new_n365_;
  assign new_n367_ = ~new_n356_ & new_n366_;
  assign p4 = ~a & new_n367_;
  assign new_n369_ = ~a & ~t1;
  assign new_n370_ = new_n312_ & new_n369_;
  assign new_n371_ = ~a1 & ~new_n370_;
  assign q4 = t2 & ~new_n371_;
  assign new_n373_ = a & ~h2;
  assign new_n374_ = ~r1 & ~s1;
  assign new_n375_ = ~q1 & new_n374_;
  assign new_n376_ = new_n373_ & new_n375_;
  assign new_n377_ = ~o & h2;
  assign new_n378_ = ~p & ~q;
  assign new_n379_ = new_n377_ & new_n378_;
  assign new_n380_ = ~new_n376_ & ~new_n379_;
  assign new_n381_ = ~o0 & new_n380_;
  assign new_n382_ = ~l2 & ~new_n381_;
  assign new_n383_ = ~f1 & ~g1;
  assign new_n384_ = ~h1 & g2;
  assign new_n385_ = new_n383_ & new_n384_;
  assign new_n386_ = ~q1 & ~r1;
  assign new_n387_ = ~s1 & ~g2;
  assign new_n388_ = new_n386_ & new_n387_;
  assign new_n389_ = ~new_n385_ & ~new_n388_;
  assign new_n390_ = ~o0 & ~new_n379_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = g2 & ~new_n385_;
  assign new_n393_ = ~s1 & ~new_n392_;
  assign new_n394_ = ~r1 & new_n393_;
  assign new_n395_ = ~q1 & new_n394_;
  assign new_n396_ = ~h2 & new_n395_;
  assign new_n397_ = ~new_n391_ & ~new_n396_;
  assign new_n398_ = a & ~new_n397_;
  assign new_n399_ = ~new_n311_ & new_n391_;
  assign new_n400_ = ~new_n398_ & ~new_n399_;
  assign r4 = new_n382_ | ~new_n400_;
  assign new_n402_ = j4 & new_n320_;
  assign new_n403_ = ~f0 & ~new_n402_;
  assign s4 = ~a & ~new_n403_;
  assign new_n405_ = ~new_n351_ & ~new_n355_;
  assign new_n406_ = e & f;
  assign new_n407_ = d & new_n406_;
  assign new_n408_ = ~r1 & ~new_n407_;
  assign new_n409_ = n & s1;
  assign new_n410_ = new_n408_ & new_n409_;
  assign new_n411_ = a & ~new_n410_;
  assign new_n412_ = ~n2 & ~o2;
  assign new_n413_ = new_n411_ & ~new_n412_;
  assign new_n414_ = ~n2 & new_n413_;
  assign new_n415_ = n2 & ~new_n413_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~new_n405_ & ~new_n416_;
  assign new_n418_ = v & s0;
  assign new_n419_ = i0 & ~s0;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = ~h4 & new_n420_;
  assign new_n422_ = ~i4 & ~new_n421_;
  assign new_n423_ = ~h4 & i4;
  assign new_n424_ = y2 & ~new_n332_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign new_n426_ = ~new_n422_ & new_n425_;
  assign new_n427_ = new_n405_ & ~new_n426_;
  assign t4 = new_n417_ | new_n427_;
  assign new_n429_ = o2 & ~new_n414_;
  assign new_n430_ = ~o2 & new_n413_;
  assign new_n431_ = ~n2 & new_n430_;
  assign new_n432_ = ~new_n429_ & ~new_n431_;
  assign new_n433_ = ~new_n405_ & ~new_n432_;
  assign new_n434_ = h4 & ~i4;
  assign new_n435_ = new_n327_ & new_n331_;
  assign new_n436_ = y2 & new_n435_;
  assign new_n437_ = ~new_n423_ & ~new_n436_;
  assign new_n438_ = ~new_n434_ & new_n437_;
  assign new_n439_ = new_n405_ & ~new_n438_;
  assign u4 = new_n433_ | new_n439_;
  assign new_n441_ = ~r2 & new_n351_;
  assign new_n442_ = new_n411_ & new_n412_;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign v4 = new_n354_ & new_n443_;
  assign new_n445_ = d2 & new_n405_;
  assign new_n446_ = b & ~new_n411_;
  assign new_n447_ = ~b & new_n411_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = ~new_n405_ & ~new_n448_;
  assign w4 = new_n445_ | new_n449_;
  assign new_n451_ = e2 & new_n405_;
  assign new_n452_ = b & new_n411_;
  assign new_n453_ = c & ~new_n452_;
  assign new_n454_ = ~c & new_n411_;
  assign new_n455_ = b & new_n454_;
  assign new_n456_ = ~new_n453_ & ~new_n455_;
  assign new_n457_ = ~new_n405_ & ~new_n456_;
  assign x4 = new_n451_ | new_n457_;
  assign new_n459_ = v0 & ~x3;
  assign y4 = a | new_n459_;
  assign z4 = v0 & b4;
  assign new_n462_ = ~c1 & d1;
  assign new_n463_ = c1 & ~d1;
  assign b5 = new_n462_ | new_n463_;
  assign new_n465_ = c1 & d1;
  assign new_n466_ = e1 & ~new_n465_;
  assign new_n467_ = d1 & ~e1;
  assign new_n468_ = c1 & new_n467_;
  assign c5 = new_n466_ | new_n468_;
  assign new_n470_ = n & ~p;
  assign new_n471_ = q & new_n470_;
  assign new_n472_ = ~d1 & ~e1;
  assign new_n473_ = ~c1 & new_n472_;
  assign new_n474_ = new_n471_ & ~new_n473_;
  assign d5 = l2 & ~new_n474_;
  assign new_n476_ = new_n471_ & ~new_n472_;
  assign e5 = l2 & ~new_n476_;
  assign new_n478_ = ~c1 & ~e1;
  assign new_n479_ = new_n471_ & ~new_n478_;
  assign f5 = l2 & ~new_n479_;
  assign new_n481_ = e1 & new_n471_;
  assign g5 = l2 & ~new_n481_;
  assign new_n483_ = ~c1 & ~d1;
  assign new_n484_ = new_n471_ & ~new_n483_;
  assign h5 = l2 & ~new_n484_;
  assign new_n486_ = d1 & new_n471_;
  assign i5 = l2 & ~new_n486_;
  assign new_n488_ = c1 & new_n471_;
  assign j5 = l2 & ~new_n488_;
  assign new_n490_ = n & c1;
  assign new_n491_ = d1 & new_n490_;
  assign l5 = e1 & new_n491_;
  assign new_n493_ = ~b1 & ~new_n305_;
  assign m5 = ~new_n407_ & ~new_n493_;
  assign new_n495_ = ~f2 & g2;
  assign new_n496_ = h2 & ~l2;
  assign new_n497_ = new_n495_ & new_n496_;
  assign n5 = a | new_n497_;
  assign new_n499_ = ~l2 & ~new_n495_;
  assign o5 = h2 & new_n499_;
  assign new_n501_ = ~h2 & ~l2;
  assign new_n502_ = ~f2 & ~g2;
  assign new_n503_ = ~new_n496_ & ~new_n502_;
  assign p5 = new_n501_ | new_n503_;
  assign new_n505_ = o & ~p;
  assign new_n506_ = ~q & new_n505_;
  assign new_n507_ = ~z2 & ~a3;
  assign new_n508_ = ~b3 & ~d3;
  assign new_n509_ = o0 & l2;
  assign new_n510_ = b3 & new_n509_;
  assign new_n511_ = ~new_n508_ & ~new_n510_;
  assign new_n512_ = ~c3 & ~new_n511_;
  assign new_n513_ = d3 & new_n509_;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = a3 & new_n321_;
  assign new_n516_ = ~z2 & new_n515_;
  assign new_n517_ = ~new_n514_ & ~new_n516_;
  assign new_n518_ = new_n507_ & new_n517_;
  assign new_n519_ = m3 & ~new_n321_;
  assign new_n520_ = h3 & i3;
  assign new_n521_ = ~new_n519_ & ~new_n520_;
  assign new_n522_ = new_n507_ & ~new_n521_;
  assign new_n523_ = ~new_n518_ & new_n522_;
  assign new_n524_ = w0 & z0;
  assign new_n525_ = ~x0 & y0;
  assign new_n526_ = x0 & ~y0;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = ~z0 & ~new_n527_;
  assign new_n529_ = ~w0 & new_n528_;
  assign new_n530_ = ~new_n524_ & ~new_n529_;
  assign new_n531_ = ~x0 & ~z0;
  assign new_n532_ = x0 & z0;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = ~w0 & ~y0;
  assign new_n535_ = w0 & y0;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = ~new_n533_ & ~new_n536_;
  assign new_n538_ = u1 & new_n537_;
  assign new_n539_ = new_n530_ & ~new_n538_;
  assign new_n540_ = j2 & ~new_n539_;
  assign new_n541_ = ~h3 & i3;
  assign new_n542_ = h3 & ~i3;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = ~n3 & ~o3;
  assign new_n545_ = ~t3 & new_n544_;
  assign new_n546_ = a2 & ~new_n545_;
  assign new_n547_ = g0 & t0;
  assign new_n548_ = ~l2 & new_n547_;
  assign new_n549_ = new_n538_ & new_n548_;
  assign new_n550_ = ~z3 & ~d8;
  assign new_n551_ = ~new_n254_ & ~new_n550_;
  assign new_n552_ = new_n506_ & ~new_n530_;
  assign new_n553_ = l2 & new_n552_;
  assign new_n554_ = new_n540_ & ~new_n553_;
  assign new_n555_ = ~h0 & new_n507_;
  assign new_n556_ = ~new_n355_ & ~new_n555_;
  assign new_n557_ = u2 & new_n556_;
  assign new_n558_ = t0 & ~new_n557_;
  assign new_n559_ = ~l3 & new_n558_;
  assign new_n560_ = ~new_n549_ & ~new_n559_;
  assign new_n561_ = new_n546_ & ~new_n560_;
  assign new_n562_ = ~new_n523_ & ~new_n543_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = ~new_n554_ & new_n563_;
  assign new_n565_ = ~new_n551_ & new_n564_;
  assign new_n566_ = k0 & l0;
  assign new_n567_ = m0 & new_n566_;
  assign new_n568_ = ~new_n540_ & new_n567_;
  assign new_n569_ = ~h0 & t0;
  assign new_n570_ = n3 & new_n569_;
  assign new_n571_ = ~j0 & ~new_n546_;
  assign new_n572_ = new_n568_ & ~new_n570_;
  assign new_n573_ = new_n565_ & new_n572_;
  assign q5 = ~new_n571_ & ~new_n573_;
  assign new_n575_ = ~g0 & h0;
  assign new_n576_ = t0 & new_n575_;
  assign new_n577_ = ~l3 & new_n576_;
  assign new_n578_ = new_n546_ & ~new_n570_;
  assign new_n579_ = ~j0 & ~new_n578_;
  assign new_n580_ = new_n568_ & ~new_n579_;
  assign new_n581_ = new_n565_ & ~new_n577_;
  assign r5 = new_n580_ & new_n581_;
  assign new_n583_ = j2 & new_n530_;
  assign new_n584_ = ~new_n538_ & new_n583_;
  assign new_n585_ = ~o3 & new_n546_;
  assign s5 = new_n584_ | new_n585_;
  assign new_n587_ = new_n546_ & new_n555_;
  assign new_n588_ = k0 & ~new_n587_;
  assign t5 = l2 | new_n588_;
  assign new_n590_ = u2 & ~new_n355_;
  assign new_n591_ = new_n546_ & ~new_n590_;
  assign new_n592_ = s0 & new_n591_;
  assign new_n593_ = l0 & ~new_n592_;
  assign u5 = ~new_n316_ | new_n593_;
  assign new_n595_ = ~o & ~new_n541_;
  assign new_n596_ = ~p2 & ~new_n595_;
  assign new_n597_ = l2 & ~new_n596_;
  assign new_n598_ = ~q & new_n597_;
  assign new_n599_ = p & new_n598_;
  assign new_n600_ = ~y1 & m2;
  assign new_n601_ = ~w1 & x1;
  assign new_n602_ = new_n600_ & new_n601_;
  assign new_n603_ = ~m0 & ~new_n602_;
  assign new_n604_ = ~new_n599_ & new_n603_;
  assign v5 = ~new_n577_ & ~new_n604_;
  assign w5 = n3 & new_n580_;
  assign new_n607_ = l2 & new_n506_;
  assign new_n608_ = k2 & ~new_n607_;
  assign x5 = new_n549_ | new_n608_;
  assign new_n610_ = t0 & l3;
  assign new_n611_ = g0 & new_n610_;
  assign y5 = new_n540_ | new_n611_;
  assign new_n613_ = ~i2 & ~k2;
  assign new_n614_ = ~d8 & ~new_n570_;
  assign z5 = ~new_n613_ | ~new_n614_;
  assign new_n616_ = ~x & y;
  assign new_n617_ = n0 & ~new_n616_;
  assign new_n618_ = e0 & new_n616_;
  assign a6 = new_n617_ | new_n618_;
  assign new_n620_ = ~m1 & ~q2;
  assign new_n621_ = ~r0 & new_n620_;
  assign b6 = m2 & ~new_n621_;
  assign new_n623_ = w1 & x1;
  assign new_n624_ = ~y1 & new_n623_;
  assign c6 = m2 & new_n624_;
  assign new_n626_ = ~p2 & q2;
  assign new_n627_ = p2 & ~q2;
  assign e6 = new_n626_ | new_n627_;
  assign new_n629_ = ~p2 & ~q2;
  assign new_n630_ = ~r0 & new_n629_;
  assign f6 = m2 & ~new_n630_;
  assign new_n632_ = p & ~m2;
  assign new_n633_ = new_n287_ & new_n632_;
  assign new_n634_ = ~new_n291_ & ~new_n633_;
  assign new_n635_ = ~p0 & ~new_n634_;
  assign new_n636_ = v3 & new_n634_;
  assign g6 = new_n635_ | new_n636_;
  assign new_n638_ = w3 & new_n634_;
  assign new_n639_ = p0 & ~q0;
  assign new_n640_ = ~p0 & q0;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n634_ & ~new_n641_;
  assign h6 = new_n638_ | new_n642_;
  assign i6 = l3 & new_n580_;
  assign new_n645_ = l2 & new_n287_;
  assign new_n646_ = ~new_n321_ & ~new_n645_;
  assign new_n647_ = r0 & new_n646_;
  assign j6 = new_n577_ | new_n647_;
  assign k6 = ~m0 & ~k2;
  assign new_n650_ = m0 & ~p2;
  assign new_n651_ = m2 & ~new_n541_;
  assign new_n652_ = new_n650_ & ~new_n651_;
  assign l6 = ~k2 & ~new_n652_;
  assign new_n654_ = ~new_n518_ & new_n569_;
  assign new_n655_ = new_n507_ & new_n654_;
  assign new_n656_ = h3 & new_n523_;
  assign new_n657_ = ~new_n577_ & ~new_n656_;
  assign m6 = new_n655_ | ~new_n657_;
  assign new_n659_ = i3 & new_n523_;
  assign new_n660_ = ~i3 & ~new_n523_;
  assign new_n661_ = h3 & new_n660_;
  assign new_n662_ = ~new_n659_ & ~new_n661_;
  assign n6 = new_n655_ | ~new_n662_;
  assign new_n664_ = new_n507_ & ~new_n518_;
  assign new_n665_ = ~new_n321_ & ~new_n543_;
  assign new_n666_ = m3 & new_n665_;
  assign new_n667_ = ~new_n655_ & ~new_n666_;
  assign new_n668_ = ~new_n520_ & new_n667_;
  assign new_n669_ = ~new_n664_ & ~new_n668_;
  assign new_n670_ = new_n518_ & ~new_n669_;
  assign new_n671_ = new_n543_ & ~new_n670_;
  assign new_n672_ = ~new_n518_ & ~new_n669_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign new_n674_ = z2 & ~new_n673_;
  assign new_n675_ = ~new_n254_ & new_n669_;
  assign o6 = new_n674_ | new_n675_;
  assign new_n677_ = ~z2 & new_n321_;
  assign new_n678_ = ~new_n283_ & ~new_n670_;
  assign new_n679_ = ~new_n672_ & ~new_n678_;
  assign new_n680_ = ~new_n677_ & ~new_n679_;
  assign new_n681_ = a3 & new_n680_;
  assign new_n682_ = ~u & new_n418_;
  assign new_n683_ = ~h0 & new_n419_;
  assign new_n684_ = ~new_n682_ & ~new_n683_;
  assign new_n685_ = new_n543_ & new_n684_;
  assign new_n686_ = new_n669_ & ~new_n685_;
  assign p6 = new_n681_ | new_n686_;
  assign new_n688_ = ~b3 & ~c3;
  assign new_n689_ = o0 & ~new_n688_;
  assign new_n690_ = z2 & new_n518_;
  assign new_n691_ = ~new_n518_ & ~new_n689_;
  assign new_n692_ = b3 & new_n691_;
  assign q6 = new_n690_ | new_n692_;
  assign new_n694_ = ~b3 & new_n321_;
  assign new_n695_ = ~new_n518_ & ~new_n694_;
  assign new_n696_ = ~new_n689_ & new_n695_;
  assign new_n697_ = c3 & new_n696_;
  assign new_n698_ = a3 & new_n518_;
  assign r6 = new_n697_ | new_n698_;
  assign new_n700_ = c3 & new_n689_;
  assign new_n701_ = ~o0 & ~new_n518_;
  assign new_n702_ = d3 & new_n701_;
  assign s6 = new_n700_ | new_n702_;
  assign new_n704_ = ~k2 & new_n607_;
  assign t6 = new_n584_ | new_n704_;
  assign u6 = ~new_n538_ & new_n547_;
  assign v6 = ~y0 & ~z0;
  assign x6 = ~w0 & ~x0;
  assign new_n709_ = q & l2;
  assign new_n710_ = p2 & new_n709_;
  assign new_n711_ = q2 & new_n710_;
  assign new_n712_ = s1 & new_n320_;
  assign new_n713_ = o1 & ~y3;
  assign new_n714_ = ~m1 & ~new_n713_;
  assign new_n715_ = ~new_n712_ & ~new_n714_;
  assign c7 = ~new_n711_ & new_n715_;
  assign new_n717_ = ~i1 & ~new_n713_;
  assign new_n718_ = m1 & ~new_n712_;
  assign new_n719_ = new_n629_ & new_n709_;
  assign new_n720_ = ~new_n718_ & new_n719_;
  assign new_n721_ = ~new_n717_ & ~new_n720_;
  assign d7 = ~new_n711_ & new_n721_;
  assign new_n723_ = i1 & e4;
  assign new_n724_ = z3 & ~new_n336_;
  assign new_n725_ = y3 & new_n724_;
  assign e7 = new_n723_ & new_n725_;
  assign new_n727_ = ~m1 & new_n629_;
  assign f7 = m2 & ~new_n727_;
  assign new_n729_ = ~new_n287_ & new_n293_;
  assign new_n730_ = q & ~m2;
  assign new_n731_ = new_n287_ & new_n730_;
  assign new_n732_ = ~new_n729_ & ~new_n731_;
  assign new_n733_ = ~k1 & ~new_n732_;
  assign new_n734_ = q3 & new_n732_;
  assign g7 = new_n733_ | new_n734_;
  assign new_n736_ = r3 & new_n732_;
  assign new_n737_ = k1 & ~l1;
  assign new_n738_ = ~k1 & l1;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = ~new_n732_ & ~new_n739_;
  assign h7 = new_n736_ | new_n740_;
  assign i7 = y3 & new_n723_;
  assign j7 = ~m1 & ~d8;
  assign k7 = i1 | new_n293_;
  assign new_n745_ = s & ~l3;
  assign new_n746_ = u2 & new_n405_;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign l7 = new_n335_ | ~new_n747_;
  assign new_n749_ = ~new_n307_ & ~new_n545_;
  assign m7 = ~new_n335_ & new_n749_;
  assign n7 = ~new_n307_ & new_n335_;
  assign new_n752_ = ~new_n335_ & new_n545_;
  assign o7 = new_n307_ | new_n752_;
  assign new_n754_ = v2 & new_n355_;
  assign new_n755_ = new_n307_ & ~new_n754_;
  assign new_n756_ = ~new_n580_ & ~new_n723_;
  assign new_n757_ = ~new_n338_ & ~new_n756_;
  assign new_n758_ = ~new_n335_ & new_n757_;
  assign new_n759_ = ~new_n321_ & ~new_n332_;
  assign new_n760_ = y2 & new_n759_;
  assign new_n761_ = new_n335_ & ~new_n760_;
  assign new_n762_ = ~new_n758_ & ~new_n761_;
  assign new_n763_ = ~new_n340_ & ~new_n762_;
  assign new_n764_ = ~new_n335_ & ~new_n723_;
  assign new_n765_ = ~new_n580_ & new_n764_;
  assign new_n766_ = ~new_n355_ & ~new_n765_;
  assign new_n767_ = ~new_n763_ & ~new_n766_;
  assign new_n768_ = ~new_n755_ & new_n767_;
  assign new_n769_ = a4 & ~new_n768_;
  assign p7 = ~d8 & new_n769_;
  assign new_n771_ = new_n251_ & ~new_n270_;
  assign new_n772_ = ~d4 & ~new_n771_;
  assign new_n773_ = ~d8 & new_n772_;
  assign q7 = ~s1 & ~new_n773_;
  assign new_n775_ = s1 & ~new_n773_;
  assign r7 = ~r1 & new_n775_;
  assign new_n777_ = u0 & s2;
  assign new_n778_ = ~k3 & p3;
  assign new_n779_ = r & ~new_n778_;
  assign x7 = new_n777_ | new_n779_;
  assign y7 = j3 & p3;
  assign new_n782_ = k & ~d0;
  assign new_n783_ = m & d0;
  assign z7 = new_n782_ | new_n783_;
  assign a8 = c4 | new_n771_;
  assign new_n786_ = ~w2 & x2;
  assign new_n787_ = new_n251_ & new_n786_;
  assign b8 = new_n270_ & new_n787_;
  assign new_n789_ = w2 & ~new_n251_;
  assign c8 = ~a4 | new_n789_;
  assign new_n791_ = x2 & ~d8;
  assign h8 = ~w2 & ~new_n791_;
  assign l4 = ~o3;
  assign d6 = ~p2;
  assign k4 = s3;
  assign m4 = t3;
  assign a5 = m2;
  assign k5 = l2;
  assign w6 = y0;
  assign y6 = w0;
  assign z6 = v6;
  assign a7 = y0;
  assign b7 = z0;
  assign s7 = w;
  assign t7 = z;
  assign u7 = a0;
  assign v7 = b0;
  assign w7 = c0;
  assign e8 = x6;
  assign f8 = w0;
  assign g8 = x0;
endmodule

