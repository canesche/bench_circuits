module top ( 
    pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps, pd0, pe1,
    pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0, pl0, pm1,
    pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1, pr2, pa,
    pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1, pv2, pt1,
    pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1, py0, pz0,
    pk, pz1, pl, pm, pn, po,
    pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4  );
  input  pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps,
    pd0, pe1, pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0,
    pw, ph0, pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0,
    pl0, pm1, pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1,
    pr2, pa, pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1,
    pv2, pt1, pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1,
    py0, pz0, pk, pz1, pl, pm, pn, po;
  output pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4;
  wire new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n408_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n442_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n464_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n489_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n513_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_;
  assign new_n166_ = ~ph0 & pt2;
  assign new_n167_ = ph0 & ~pt2;
  assign new_n168_ = ~pq2 & ~pi;
  assign new_n169_ = ~new_n166_ & ~new_n167_;
  assign new_n170_ = ~new_n168_ & new_n169_;
  assign new_n171_ = pn2 & ~pp2;
  assign new_n172_ = ~po2 & pr2;
  assign new_n173_ = new_n171_ & new_n172_;
  assign new_n174_ = pe1 & new_n170_;
  assign new_n175_ = new_n173_ & new_n174_;
  assign new_n176_ = ~pi0 & new_n175_;
  assign new_n177_ = pe1 & ~new_n168_;
  assign new_n178_ = pn2 & ~po2;
  assign new_n179_ = new_n177_ & new_n178_;
  assign new_n180_ = pr2 & new_n179_;
  assign new_n181_ = ~pp2 & new_n180_;
  assign new_n182_ = ps2 & ~new_n181_;
  assign new_n183_ = ~pi0 & new_n182_;
  assign pc3 = new_n176_ | new_n183_;
  assign new_n185_ = po2 & ~pq2;
  assign new_n186_ = ~pp2 & new_n185_;
  assign new_n187_ = ~pr2 & new_n186_;
  assign new_n188_ = ~pc1 & pk1;
  assign new_n189_ = ~new_n187_ & new_n188_;
  assign new_n190_ = ~pp2 & ~pq2;
  assign new_n191_ = ~pr2 & new_n190_;
  assign new_n192_ = ~pn2 & new_n191_;
  assign new_n193_ = pe1 & po2;
  assign new_n194_ = new_n192_ & new_n193_;
  assign new_n195_ = ~pc1 & new_n194_;
  assign new_n196_ = pn2 & new_n195_;
  assign new_n197_ = ~pe1 & new_n188_;
  assign new_n198_ = pt0 & new_n188_;
  assign new_n199_ = pn2 & new_n188_;
  assign new_n200_ = ~new_n187_ & new_n195_;
  assign new_n201_ = ~pe1 & new_n195_;
  assign new_n202_ = pt0 & new_n195_;
  assign new_n203_ = ~new_n189_ & ~new_n196_;
  assign new_n204_ = ~new_n197_ & ~new_n198_;
  assign new_n205_ = new_n203_ & new_n204_;
  assign new_n206_ = ~new_n201_ & ~new_n202_;
  assign new_n207_ = ~new_n199_ & ~new_n200_;
  assign new_n208_ = new_n206_ & new_n207_;
  assign pd4 = ~new_n205_ | ~new_n208_;
  assign new_n210_ = pb & ~pu0;
  assign new_n211_ = ~pk2 & ~pl2;
  assign new_n212_ = ~pk2 & pm2;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~pc1 & new_n213_;
  assign new_n215_ = new_n210_ & new_n214_;
  assign new_n216_ = ~pk2 & new_n215_;
  assign new_n217_ = ~pl2 & new_n215_;
  assign new_n218_ = pu2 & new_n214_;
  assign new_n219_ = ~pk2 & new_n218_;
  assign new_n220_ = ~pl2 & new_n218_;
  assign new_n221_ = pl2 & new_n214_;
  assign new_n222_ = ~pk2 & new_n221_;
  assign new_n223_ = ~pu2 & ~new_n210_;
  assign new_n224_ = new_n214_ & new_n223_;
  assign new_n225_ = new_n210_ & new_n224_;
  assign new_n226_ = pl2 & new_n224_;
  assign new_n227_ = pu2 & new_n224_;
  assign new_n228_ = ~new_n216_ & ~new_n217_;
  assign new_n229_ = ~new_n219_ & ~new_n220_;
  assign new_n230_ = new_n228_ & new_n229_;
  assign new_n231_ = ~new_n226_ & ~new_n227_;
  assign new_n232_ = ~new_n222_ & ~new_n225_;
  assign new_n233_ = new_n231_ & new_n232_;
  assign pe5 = ~new_n230_ | ~new_n233_;
  assign new_n235_ = pk2 & pu2;
  assign new_n236_ = pk2 & pb;
  assign new_n237_ = ~pu0 & new_n236_;
  assign new_n238_ = ~new_n235_ & ~new_n237_;
  assign new_n239_ = ~pc1 & new_n238_;
  assign new_n240_ = pk2 & new_n239_;
  assign new_n241_ = new_n210_ & new_n239_;
  assign new_n242_ = pu2 & new_n239_;
  assign new_n243_ = ~new_n240_ & ~new_n241_;
  assign pd5 = new_n242_ | ~new_n243_;
  assign new_n245_ = ~po2 & ~pq2;
  assign new_n246_ = ~pr2 & ~pp2;
  assign new_n247_ = new_n245_ & new_n246_;
  assign new_n248_ = pe1 & new_n247_;
  assign new_n249_ = pn2 & new_n248_;
  assign new_n250_ = ~pc1 & new_n249_;
  assign new_n251_ = ~pc1 & pl1;
  assign pe4 = new_n250_ | new_n251_;
  assign new_n253_ = pg0 & pv2;
  assign new_n254_ = ~pi0 & ~new_n253_;
  assign new_n255_ = pl2 & pm2;
  assign new_n256_ = ~ph & new_n255_;
  assign new_n257_ = ~pk2 & ~pg;
  assign new_n258_ = new_n256_ & new_n257_;
  assign new_n259_ = new_n254_ & new_n258_;
  assign new_n260_ = pm1 & new_n254_;
  assign pf4 = new_n259_ | new_n260_;
  assign new_n262_ = pn2 & pm2;
  assign new_n263_ = pl2 & new_n262_;
  assign new_n264_ = ~pk2 & new_n263_;
  assign new_n265_ = pe1 & pn2;
  assign new_n266_ = pd1 & pn2;
  assign new_n267_ = ~new_n264_ & ~new_n265_;
  assign new_n268_ = ~pc1 & ~new_n266_;
  assign new_n269_ = new_n267_ & new_n268_;
  assign new_n270_ = ~pk2 & pl2;
  assign new_n271_ = pm2 & new_n270_;
  assign new_n272_ = new_n269_ & new_n271_;
  assign new_n273_ = pe1 & new_n269_;
  assign new_n274_ = pd1 & new_n269_;
  assign new_n275_ = pn2 & new_n269_;
  assign new_n276_ = ~new_n272_ & ~new_n273_;
  assign new_n277_ = ~new_n274_ & ~new_n275_;
  assign pg5 = ~new_n276_ | ~new_n277_;
  assign new_n279_ = ~pl2 & ~pm2;
  assign new_n280_ = ~pk2 & ~pm2;
  assign new_n281_ = ~new_n270_ & ~new_n279_;
  assign new_n282_ = ~pc1 & ~new_n280_;
  assign new_n283_ = new_n281_ & new_n282_;
  assign new_n284_ = new_n210_ & new_n283_;
  assign new_n285_ = ~pl2 & new_n284_;
  assign new_n286_ = ~pm2 & new_n284_;
  assign new_n287_ = pu2 & new_n283_;
  assign new_n288_ = ~pl2 & new_n287_;
  assign new_n289_ = ~pm2 & new_n287_;
  assign new_n290_ = pm2 & new_n283_;
  assign new_n291_ = ~pl2 & new_n290_;
  assign new_n292_ = new_n223_ & new_n283_;
  assign new_n293_ = new_n210_ & new_n292_;
  assign new_n294_ = pm2 & new_n292_;
  assign new_n295_ = pu2 & new_n292_;
  assign new_n296_ = ~new_n285_ & ~new_n286_;
  assign new_n297_ = ~new_n288_ & ~new_n289_;
  assign new_n298_ = new_n296_ & new_n297_;
  assign new_n299_ = ~new_n294_ & ~new_n295_;
  assign new_n300_ = ~new_n291_ & ~new_n293_;
  assign new_n301_ = new_n299_ & new_n300_;
  assign pf5 = ~new_n298_ | ~new_n301_;
  assign new_n303_ = pg0 & pm1;
  assign new_n304_ = pv2 & new_n303_;
  assign new_n305_ = ph & new_n304_;
  assign new_n306_ = ~ph0 & new_n304_;
  assign new_n307_ = pg & new_n304_;
  assign new_n308_ = ~new_n305_ & ~new_n306_;
  assign new_n309_ = ~new_n307_ & new_n308_;
  assign new_n310_ = pe1 & ~po1;
  assign new_n311_ = ~pm0 & new_n309_;
  assign new_n312_ = new_n310_ & new_n311_;
  assign new_n313_ = ~pi0 & new_n312_;
  assign new_n314_ = pm1 & pv2;
  assign new_n315_ = pg0 & new_n314_;
  assign new_n316_ = pi & new_n315_;
  assign new_n317_ = ~pi0 & new_n316_;
  assign new_n318_ = ph & new_n303_;
  assign new_n319_ = pv2 & new_n318_;
  assign new_n320_ = ~ph0 & new_n315_;
  assign new_n321_ = pg & new_n303_;
  assign new_n322_ = pv2 & new_n321_;
  assign new_n323_ = pe1 & ~pm0;
  assign new_n324_ = ~new_n319_ & ~new_n320_;
  assign new_n325_ = ~new_n322_ & ~new_n323_;
  assign new_n326_ = new_n324_ & new_n325_;
  assign new_n327_ = pn1 & new_n326_;
  assign new_n328_ = ~pi0 & new_n327_;
  assign new_n329_ = ~new_n313_ & ~new_n317_;
  assign pg4 = new_n328_ | ~new_n329_;
  assign new_n331_ = ~pg & ~pi;
  assign new_n332_ = ~ph & new_n331_;
  assign new_n333_ = ph0 & new_n332_;
  assign new_n334_ = ~pi0 & pm1;
  assign new_n335_ = pv2 & new_n334_;
  assign new_n336_ = pc0 & ~new_n333_;
  assign new_n337_ = new_n335_ & new_n336_;
  assign new_n338_ = pg0 & new_n337_;
  assign new_n339_ = pe1 & pi2;
  assign new_n340_ = pi & new_n304_;
  assign new_n341_ = ~new_n307_ & ~new_n340_;
  assign new_n342_ = new_n308_ & new_n341_;
  assign new_n343_ = ~pm0 & new_n339_;
  assign new_n344_ = new_n342_ & new_n343_;
  assign new_n345_ = ~pi0 & new_n344_;
  assign new_n346_ = pm1 & ~new_n333_;
  assign new_n347_ = pg0 & new_n346_;
  assign new_n348_ = pv2 & new_n347_;
  assign new_n349_ = ~new_n323_ & ~new_n348_;
  assign new_n350_ = ph2 & new_n349_;
  assign new_n351_ = ~pi0 & new_n350_;
  assign new_n352_ = ~new_n338_ & ~new_n345_;
  assign pa5 = new_n351_ | ~new_n352_;
  assign new_n354_ = ~pn0 & ~new_n191_;
  assign new_n355_ = ~pn2 & ~pn0;
  assign new_n356_ = ~pe1 & ~pn0;
  assign new_n357_ = po2 & ~pn0;
  assign new_n358_ = ~new_n354_ & ~new_n355_;
  assign new_n359_ = ~new_n356_ & ~new_n357_;
  assign new_n360_ = new_n358_ & new_n359_;
  assign new_n361_ = ~pi0 & new_n360_;
  assign pg3 = ~pc1 & new_n361_;
  assign new_n363_ = ~pc1 & ph1;
  assign new_n364_ = ~new_n187_ & new_n363_;
  assign new_n365_ = ~pe1 & new_n363_;
  assign new_n366_ = pq0 & new_n363_;
  assign new_n367_ = pn2 & new_n363_;
  assign new_n368_ = pq0 & new_n195_;
  assign new_n369_ = ~new_n196_ & ~new_n364_;
  assign new_n370_ = ~new_n365_ & ~new_n366_;
  assign new_n371_ = new_n369_ & new_n370_;
  assign new_n372_ = ~new_n201_ & ~new_n368_;
  assign new_n373_ = ~new_n200_ & ~new_n367_;
  assign new_n374_ = new_n372_ & new_n373_;
  assign pa4 = ~new_n371_ | ~new_n374_;
  assign new_n376_ = ~ph0 & pm1;
  assign new_n377_ = pm1 & ph;
  assign new_n378_ = pm1 & pi;
  assign new_n379_ = pm1 & pg;
  assign new_n380_ = ~new_n376_ & ~new_n377_;
  assign new_n381_ = ~new_n378_ & ~new_n379_;
  assign new_n382_ = new_n380_ & new_n381_;
  assign new_n383_ = pg0 & new_n382_;
  assign new_n384_ = pv2 & new_n383_;
  assign new_n385_ = ~pi0 & new_n253_;
  assign new_n386_ = ~pi0 & ~pm0;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign pf3 = new_n384_ | new_n387_;
  assign new_n389_ = ~pc1 & pi1;
  assign new_n390_ = ~new_n187_ & new_n389_;
  assign new_n391_ = ~pe1 & new_n389_;
  assign new_n392_ = pr0 & new_n389_;
  assign new_n393_ = pn2 & new_n389_;
  assign new_n394_ = pr0 & new_n195_;
  assign new_n395_ = ~new_n196_ & ~new_n390_;
  assign new_n396_ = ~new_n391_ & ~new_n392_;
  assign new_n397_ = new_n395_ & new_n396_;
  assign new_n398_ = ~new_n201_ & ~new_n394_;
  assign new_n399_ = ~new_n200_ & ~new_n393_;
  assign new_n400_ = new_n398_ & new_n399_;
  assign pb4 = ~new_n397_ | ~new_n400_;
  assign new_n402_ = pe0 & ~new_n333_;
  assign new_n403_ = new_n335_ & new_n402_;
  assign new_n404_ = pg0 & new_n403_;
  assign new_n405_ = ~pi0 & new_n349_;
  assign new_n406_ = pj2 & new_n405_;
  assign pc5 = new_n404_ | new_n406_;
  assign new_n408_ = ~pc1 & pl0;
  assign pe3 = new_n250_ | new_n408_;
  assign new_n410_ = pd0 & ~new_n333_;
  assign new_n411_ = new_n335_ & new_n410_;
  assign new_n412_ = pg0 & new_n411_;
  assign new_n413_ = pe1 & pj2;
  assign new_n414_ = ~pm0 & new_n413_;
  assign new_n415_ = new_n342_ & new_n414_;
  assign new_n416_ = ~pi0 & new_n415_;
  assign new_n417_ = pi2 & new_n349_;
  assign new_n418_ = ~pi0 & new_n417_;
  assign new_n419_ = ~new_n412_ & ~new_n416_;
  assign pb5 = new_n418_ | ~new_n419_;
  assign new_n421_ = ~pc1 & pj1;
  assign new_n422_ = ~new_n187_ & new_n421_;
  assign new_n423_ = ~pe1 & new_n421_;
  assign new_n424_ = ps0 & new_n421_;
  assign new_n425_ = pn2 & new_n421_;
  assign new_n426_ = ps0 & new_n195_;
  assign new_n427_ = ~new_n196_ & ~new_n422_;
  assign new_n428_ = ~new_n423_ & ~new_n424_;
  assign new_n429_ = new_n427_ & new_n428_;
  assign new_n430_ = ~new_n201_ & ~new_n426_;
  assign new_n431_ = ~new_n200_ & ~new_n425_;
  assign new_n432_ = new_n430_ & new_n431_;
  assign pc4 = ~new_n429_ | ~new_n432_;
  assign new_n434_ = ~pc1 & new_n382_;
  assign new_n435_ = pg0 & new_n434_;
  assign new_n436_ = pv2 & new_n435_;
  assign new_n437_ = ~pf0 & ~pk0;
  assign new_n438_ = ~pk0 & ~pv2;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_ = ~pc1 & new_n439_;
  assign pd3 = new_n436_ | new_n440_;
  assign new_n442_ = ~pi0 & pr0;
  assign pk3 = ~pc1 & new_n442_;
  assign new_n444_ = pn & ~new_n333_;
  assign new_n445_ = new_n335_ & new_n444_;
  assign new_n446_ = pg0 & new_n445_;
  assign new_n447_ = pe1 & pt1;
  assign new_n448_ = ~pm0 & new_n447_;
  assign new_n449_ = new_n342_ & new_n448_;
  assign new_n450_ = ~pi0 & new_n449_;
  assign new_n451_ = ps1 & new_n349_;
  assign new_n452_ = ~pi0 & new_n451_;
  assign new_n453_ = ~new_n446_ & ~new_n450_;
  assign pl4 = new_n452_ | ~new_n453_;
  assign new_n455_ = ~ps2 & pt2;
  assign new_n456_ = ~pc1 & new_n455_;
  assign new_n457_ = pl1 & ~pt2;
  assign new_n458_ = ps2 & new_n457_;
  assign new_n459_ = ~pc1 & new_n458_;
  assign new_n460_ = ~pl1 & pt2;
  assign new_n461_ = ~pc1 & new_n460_;
  assign new_n462_ = ~new_n456_ & ~new_n459_;
  assign pm5 = new_n461_ | ~new_n462_;
  assign new_n464_ = ~pi0 & pq0;
  assign pj3 = ~pc1 & new_n464_;
  assign new_n466_ = ~pm0 & pn1;
  assign new_n467_ = pe1 & new_n466_;
  assign new_n468_ = ~pi0 & new_n467_;
  assign new_n469_ = pb1 & ~pe1;
  assign new_n470_ = ~pi0 & new_n469_;
  assign new_n471_ = pb1 & pn1;
  assign new_n472_ = ~pi0 & new_n471_;
  assign new_n473_ = pb1 & pm0;
  assign new_n474_ = ~pi0 & new_n473_;
  assign new_n475_ = ~new_n468_ & ~new_n470_;
  assign new_n476_ = ~new_n472_ & ~new_n474_;
  assign pl5 = ~new_n475_ | ~new_n476_;
  assign new_n478_ = po & ~new_n333_;
  assign new_n479_ = new_n335_ & new_n478_;
  assign new_n480_ = pg0 & new_n479_;
  assign new_n481_ = pe1 & pu1;
  assign new_n482_ = ~pm0 & new_n481_;
  assign new_n483_ = new_n342_ & new_n482_;
  assign new_n484_ = ~pi0 & new_n483_;
  assign new_n485_ = pt1 & new_n349_;
  assign new_n486_ = ~pi0 & new_n485_;
  assign new_n487_ = ~new_n480_ & ~new_n484_;
  assign pm4 = new_n486_ | ~new_n487_;
  assign new_n489_ = ~pi0 & pp0;
  assign pi3 = ~pc1 & new_n489_;
  assign new_n491_ = pp & ~new_n333_;
  assign new_n492_ = new_n335_ & new_n491_;
  assign new_n493_ = pg0 & new_n492_;
  assign new_n494_ = pe1 & pv1;
  assign new_n495_ = ~pm0 & new_n494_;
  assign new_n496_ = new_n342_ & new_n495_;
  assign new_n497_ = ~pi0 & new_n496_;
  assign new_n498_ = pu1 & new_n349_;
  assign new_n499_ = ~pi0 & new_n498_;
  assign new_n500_ = ~new_n493_ & ~new_n497_;
  assign pn4 = new_n499_ | ~new_n500_;
  assign new_n502_ = pv2 & new_n254_;
  assign new_n503_ = ~pf0 & new_n502_;
  assign new_n504_ = pr2 & ~pp2;
  assign new_n505_ = ~po2 & new_n504_;
  assign new_n506_ = pq2 & new_n505_;
  assign new_n507_ = pi & new_n505_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = pn2 & ~new_n508_;
  assign new_n510_ = pe1 & new_n509_;
  assign new_n511_ = new_n254_ & new_n510_;
  assign po5 = new_n503_ | new_n511_;
  assign new_n513_ = ~pi0 & po0;
  assign ph3 = ~pc1 & new_n513_;
  assign new_n515_ = ~pb & ~pu2;
  assign new_n516_ = pu0 & ~pu2;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = ~pi0 & new_n517_;
  assign new_n519_ = new_n210_ & new_n518_;
  assign new_n520_ = ~pl2 & new_n518_;
  assign new_n521_ = pk2 & new_n518_;
  assign new_n522_ = ~pm2 & new_n518_;
  assign new_n523_ = ~new_n519_ & ~new_n520_;
  assign new_n524_ = ~new_n521_ & ~new_n522_;
  assign pn5 = ~new_n523_ | ~new_n524_;
  assign new_n526_ = pq & ~new_n333_;
  assign new_n527_ = new_n335_ & new_n526_;
  assign new_n528_ = pg0 & new_n527_;
  assign new_n529_ = pe1 & pw1;
  assign new_n530_ = ~pm0 & new_n529_;
  assign new_n531_ = new_n342_ & new_n530_;
  assign new_n532_ = ~pi0 & new_n531_;
  assign new_n533_ = pv1 & new_n349_;
  assign new_n534_ = ~pi0 & new_n533_;
  assign new_n535_ = ~new_n528_ & ~new_n532_;
  assign po4 = new_n534_ | ~new_n535_;
  assign new_n537_ = ~pm0 & pp1;
  assign new_n538_ = pe1 & new_n537_;
  assign new_n539_ = ~pi0 & new_n538_;
  assign new_n540_ = ~pe1 & ~po1;
  assign new_n541_ = ~pi0 & new_n540_;
  assign new_n542_ = ~po1 & pp1;
  assign new_n543_ = ~pi0 & new_n542_;
  assign new_n544_ = pm0 & ~po1;
  assign new_n545_ = ~pi0 & new_n544_;
  assign new_n546_ = ~new_n539_ & ~new_n541_;
  assign new_n547_ = ~new_n543_ & ~new_n545_;
  assign new_n548_ = new_n546_ & new_n547_;
  assign ph4 = new_n348_ | new_n548_;
  assign new_n550_ = ~pn2 & ~pp2;
  assign new_n551_ = ~po2 & ~pp2;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~pc1 & new_n552_;
  assign new_n554_ = pe1 & new_n553_;
  assign new_n555_ = ~po2 & new_n554_;
  assign new_n556_ = ~pp2 & new_n554_;
  assign new_n557_ = pp2 & new_n553_;
  assign new_n558_ = ~po2 & new_n557_;
  assign new_n559_ = ~pn2 & new_n554_;
  assign new_n560_ = ~pn2 & new_n557_;
  assign new_n561_ = ~pk2 & new_n255_;
  assign new_n562_ = ~pd1 & ~new_n561_;
  assign new_n563_ = ~pe1 & new_n562_;
  assign new_n564_ = new_n553_ & new_n563_;
  assign new_n565_ = pe1 & new_n564_;
  assign new_n566_ = pd1 & new_n564_;
  assign new_n567_ = new_n271_ & new_n564_;
  assign new_n568_ = new_n271_ & new_n553_;
  assign new_n569_ = ~pp2 & new_n568_;
  assign new_n570_ = pp2 & new_n564_;
  assign new_n571_ = ~po2 & new_n568_;
  assign new_n572_ = pd1 & new_n553_;
  assign new_n573_ = ~pp2 & new_n572_;
  assign new_n574_ = ~pn2 & new_n568_;
  assign new_n575_ = ~pn2 & new_n572_;
  assign new_n576_ = ~po2 & new_n572_;
  assign new_n577_ = ~new_n555_ & ~new_n556_;
  assign new_n578_ = ~new_n558_ & ~new_n559_;
  assign new_n579_ = new_n577_ & new_n578_;
  assign new_n580_ = ~new_n566_ & ~new_n567_;
  assign new_n581_ = ~new_n560_ & ~new_n565_;
  assign new_n582_ = new_n580_ & new_n581_;
  assign new_n583_ = new_n579_ & new_n582_;
  assign new_n584_ = ~new_n574_ & ~new_n575_;
  assign new_n585_ = ~new_n576_ & new_n584_;
  assign new_n586_ = ~new_n571_ & ~new_n573_;
  assign new_n587_ = ~new_n569_ & ~new_n570_;
  assign new_n588_ = new_n586_ & new_n587_;
  assign new_n589_ = new_n585_ & new_n588_;
  assign pi5 = ~new_n583_ | ~new_n589_;
  assign po3 = ~pi0 & pa;
  assign new_n592_ = ~pn2 & ~po2;
  assign new_n593_ = ~pc1 & ~new_n592_;
  assign new_n594_ = pd1 & new_n593_;
  assign new_n595_ = ~pn2 & new_n594_;
  assign new_n596_ = ~po2 & new_n594_;
  assign new_n597_ = pe1 & new_n593_;
  assign new_n598_ = ~pn2 & new_n597_;
  assign new_n599_ = ~po2 & new_n597_;
  assign new_n600_ = po2 & new_n593_;
  assign new_n601_ = ~pn2 & new_n600_;
  assign new_n602_ = new_n563_ & new_n593_;
  assign new_n603_ = new_n271_ & new_n602_;
  assign new_n604_ = pd1 & new_n602_;
  assign new_n605_ = po2 & new_n602_;
  assign new_n606_ = pe1 & new_n602_;
  assign new_n607_ = new_n271_ & new_n593_;
  assign new_n608_ = ~pn2 & new_n607_;
  assign new_n609_ = ~po2 & new_n607_;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign new_n611_ = ~new_n604_ & ~new_n605_;
  assign new_n612_ = ~new_n606_ & new_n611_;
  assign new_n613_ = new_n610_ & new_n612_;
  assign new_n614_ = ~new_n595_ & ~new_n596_;
  assign new_n615_ = ~new_n598_ & new_n614_;
  assign new_n616_ = ~new_n599_ & ~new_n601_;
  assign new_n617_ = ~new_n603_ & new_n616_;
  assign new_n618_ = new_n615_ & new_n617_;
  assign ph5 = ~new_n613_ | ~new_n618_;
  assign new_n620_ = ~new_n333_ & new_n335_;
  assign new_n621_ = pk & new_n620_;
  assign new_n622_ = pg0 & new_n621_;
  assign new_n623_ = pe1 & pq1;
  assign new_n624_ = ~pm0 & new_n342_;
  assign new_n625_ = new_n623_ & new_n624_;
  assign new_n626_ = ~pi0 & new_n625_;
  assign new_n627_ = pp1 & new_n349_;
  assign new_n628_ = ~pi0 & new_n627_;
  assign new_n629_ = ~new_n622_ & ~new_n626_;
  assign pi4 = new_n628_ | ~new_n629_;
  assign pn3 = ~pi0 & pb;
  assign new_n632_ = pl & ~new_n333_;
  assign new_n633_ = new_n335_ & new_n632_;
  assign new_n634_ = pg0 & new_n633_;
  assign new_n635_ = pe1 & pr1;
  assign new_n636_ = ~pm0 & new_n635_;
  assign new_n637_ = new_n342_ & new_n636_;
  assign new_n638_ = ~pi0 & new_n637_;
  assign new_n639_ = pq1 & new_n349_;
  assign new_n640_ = ~pi0 & new_n639_;
  assign new_n641_ = ~new_n634_ & ~new_n638_;
  assign pj4 = new_n640_ | ~new_n641_;
  assign new_n643_ = pp2 & pq2;
  assign new_n644_ = pr2 & new_n643_;
  assign new_n645_ = ~pc1 & ~new_n644_;
  assign new_n646_ = pr2 & new_n645_;
  assign new_n647_ = pn2 & pp2;
  assign new_n648_ = po2 & pq2;
  assign new_n649_ = new_n647_ & new_n648_;
  assign new_n650_ = ~pc1 & pe1;
  assign new_n651_ = new_n649_ & new_n650_;
  assign new_n652_ = ~pn2 & new_n651_;
  assign new_n653_ = ~pc1 & pr2;
  assign new_n654_ = ~po2 & new_n653_;
  assign new_n655_ = ~pc1 & new_n563_;
  assign new_n656_ = pr2 & new_n655_;
  assign new_n657_ = ~pn2 & new_n653_;
  assign new_n658_ = new_n649_ & new_n655_;
  assign new_n659_ = new_n271_ & new_n658_;
  assign new_n660_ = new_n645_ & new_n649_;
  assign new_n661_ = pe1 & new_n660_;
  assign new_n662_ = pd1 & new_n660_;
  assign new_n663_ = new_n271_ & new_n660_;
  assign new_n664_ = pe1 & new_n658_;
  assign new_n665_ = pd1 & new_n658_;
  assign new_n666_ = ~pc1 & new_n271_;
  assign new_n667_ = new_n649_ & new_n666_;
  assign new_n668_ = ~po2 & new_n667_;
  assign new_n669_ = ~pc1 & pd1;
  assign new_n670_ = new_n649_ & new_n669_;
  assign new_n671_ = ~po2 & new_n670_;
  assign new_n672_ = ~pn2 & new_n667_;
  assign new_n673_ = ~po2 & new_n651_;
  assign new_n674_ = ~pn2 & new_n670_;
  assign new_n675_ = ~new_n646_ & ~new_n652_;
  assign new_n676_ = ~new_n654_ & ~new_n656_;
  assign new_n677_ = new_n675_ & new_n676_;
  assign new_n678_ = ~new_n661_ & ~new_n662_;
  assign new_n679_ = ~new_n657_ & ~new_n659_;
  assign new_n680_ = new_n678_ & new_n679_;
  assign new_n681_ = new_n677_ & new_n680_;
  assign new_n682_ = ~new_n665_ & ~new_n668_;
  assign new_n683_ = ~new_n663_ & ~new_n664_;
  assign new_n684_ = new_n682_ & new_n683_;
  assign new_n685_ = ~new_n671_ & ~new_n672_;
  assign new_n686_ = ~new_n673_ & ~new_n674_;
  assign new_n687_ = new_n685_ & new_n686_;
  assign new_n688_ = new_n684_ & new_n687_;
  assign pk5 = ~new_n681_ | ~new_n688_;
  assign new_n690_ = ~pi0 & pt0;
  assign pm3 = ~pc1 & new_n690_;
  assign new_n692_ = ~pn2 & ~pq2;
  assign new_n693_ = ~new_n190_ & ~new_n692_;
  assign new_n694_ = ~pc1 & ~new_n245_;
  assign new_n695_ = new_n693_ & new_n694_;
  assign new_n696_ = pq2 & new_n695_;
  assign new_n697_ = new_n563_ & new_n696_;
  assign new_n698_ = pe1 & new_n695_;
  assign new_n699_ = ~po2 & new_n698_;
  assign new_n700_ = ~pn2 & new_n696_;
  assign new_n701_ = ~new_n643_ & new_n696_;
  assign new_n702_ = ~po2 & new_n696_;
  assign new_n703_ = new_n271_ & new_n695_;
  assign new_n704_ = ~po2 & new_n703_;
  assign new_n705_ = ~pn2 & new_n703_;
  assign new_n706_ = ~new_n643_ & new_n703_;
  assign new_n707_ = new_n563_ & new_n703_;
  assign new_n708_ = pd1 & new_n695_;
  assign new_n709_ = ~new_n643_ & new_n708_;
  assign new_n710_ = new_n563_ & new_n708_;
  assign new_n711_ = ~pn2 & new_n708_;
  assign new_n712_ = new_n563_ & new_n698_;
  assign new_n713_ = ~po2 & new_n708_;
  assign new_n714_ = ~pn2 & new_n698_;
  assign new_n715_ = ~new_n643_ & new_n698_;
  assign new_n716_ = ~new_n697_ & ~new_n699_;
  assign new_n717_ = ~new_n700_ & ~new_n701_;
  assign new_n718_ = new_n716_ & new_n717_;
  assign new_n719_ = ~new_n705_ & ~new_n706_;
  assign new_n720_ = ~new_n702_ & ~new_n704_;
  assign new_n721_ = new_n719_ & new_n720_;
  assign new_n722_ = new_n718_ & new_n721_;
  assign new_n723_ = ~new_n710_ & ~new_n711_;
  assign new_n724_ = ~new_n707_ & ~new_n709_;
  assign new_n725_ = new_n723_ & new_n724_;
  assign new_n726_ = ~new_n712_ & ~new_n713_;
  assign new_n727_ = ~new_n714_ & ~new_n715_;
  assign new_n728_ = new_n726_ & new_n727_;
  assign new_n729_ = new_n725_ & new_n728_;
  assign pj5 = ~new_n722_ | ~new_n729_;
  assign new_n731_ = pm & ~new_n333_;
  assign new_n732_ = new_n335_ & new_n731_;
  assign new_n733_ = pg0 & new_n732_;
  assign new_n734_ = pe1 & ps1;
  assign new_n735_ = ~pm0 & new_n734_;
  assign new_n736_ = new_n342_ & new_n735_;
  assign new_n737_ = ~pi0 & new_n736_;
  assign new_n738_ = pr1 & new_n349_;
  assign new_n739_ = ~pi0 & new_n738_;
  assign new_n740_ = ~new_n733_ & ~new_n737_;
  assign pk4 = new_n739_ | ~new_n740_;
  assign new_n742_ = ~pi0 & ps0;
  assign pl3 = ~pc1 & new_n742_;
  assign ps3 = ~pi0 & py0;
  assign new_n745_ = pv & ~new_n333_;
  assign new_n746_ = new_n335_ & new_n745_;
  assign new_n747_ = pg0 & new_n746_;
  assign new_n748_ = pb2 & pe1;
  assign new_n749_ = ~pm0 & new_n748_;
  assign new_n750_ = new_n342_ & new_n749_;
  assign new_n751_ = ~pi0 & new_n750_;
  assign new_n752_ = pa2 & new_n349_;
  assign new_n753_ = ~pi0 & new_n752_;
  assign new_n754_ = ~new_n747_ & ~new_n751_;
  assign pt4 = new_n753_ | ~new_n754_;
  assign pr3 = ~pi0 & px0;
  assign new_n757_ = pw & ~new_n333_;
  assign new_n758_ = new_n335_ & new_n757_;
  assign new_n759_ = pg0 & new_n758_;
  assign new_n760_ = pc2 & pe1;
  assign new_n761_ = ~pm0 & new_n760_;
  assign new_n762_ = new_n342_ & new_n761_;
  assign new_n763_ = ~pi0 & new_n762_;
  assign new_n764_ = pb2 & new_n349_;
  assign new_n765_ = ~pi0 & new_n764_;
  assign new_n766_ = ~new_n759_ & ~new_n763_;
  assign pu4 = new_n765_ | ~new_n766_;
  assign pq3 = ~pi0 & pw0;
  assign new_n769_ = px & ~new_n333_;
  assign new_n770_ = new_n335_ & new_n769_;
  assign new_n771_ = pg0 & new_n770_;
  assign new_n772_ = pe1 & pd2;
  assign new_n773_ = ~pm0 & new_n772_;
  assign new_n774_ = new_n342_ & new_n773_;
  assign new_n775_ = ~pi0 & new_n774_;
  assign new_n776_ = pc2 & new_n349_;
  assign new_n777_ = ~pi0 & new_n776_;
  assign new_n778_ = ~new_n771_ & ~new_n775_;
  assign pv4 = new_n777_ | ~new_n778_;
  assign pp3 = ~pi0 & pv0;
  assign new_n781_ = py & ~new_n333_;
  assign new_n782_ = new_n335_ & new_n781_;
  assign new_n783_ = pg0 & new_n782_;
  assign new_n784_ = pe1 & pe2;
  assign new_n785_ = ~pm0 & new_n784_;
  assign new_n786_ = new_n342_ & new_n785_;
  assign new_n787_ = ~pi0 & new_n786_;
  assign new_n788_ = pd2 & new_n349_;
  assign new_n789_ = ~pi0 & new_n788_;
  assign new_n790_ = ~new_n783_ & ~new_n787_;
  assign pw4 = new_n789_ | ~new_n790_;
  assign new_n792_ = pr & ~new_n333_;
  assign new_n793_ = new_n335_ & new_n792_;
  assign new_n794_ = pg0 & new_n793_;
  assign new_n795_ = pe1 & px1;
  assign new_n796_ = ~pm0 & new_n795_;
  assign new_n797_ = new_n342_ & new_n796_;
  assign new_n798_ = ~pi0 & new_n797_;
  assign new_n799_ = pw1 & new_n349_;
  assign new_n800_ = ~pi0 & new_n799_;
  assign new_n801_ = ~new_n794_ & ~new_n798_;
  assign pp4 = new_n800_ | ~new_n801_;
  assign new_n803_ = ph0 & ~ph;
  assign new_n804_ = ~pi & new_n803_;
  assign new_n805_ = ~pg & new_n804_;
  assign new_n806_ = ~pg0 & ~new_n805_;
  assign new_n807_ = pi0 & ~pm1;
  assign new_n808_ = new_n806_ & new_n807_;
  assign pw3 = pv2 & new_n808_;
  assign new_n810_ = ps & ~new_n333_;
  assign new_n811_ = new_n335_ & new_n810_;
  assign new_n812_ = pg0 & new_n811_;
  assign new_n813_ = pe1 & py1;
  assign new_n814_ = ~pm0 & new_n813_;
  assign new_n815_ = new_n342_ & new_n814_;
  assign new_n816_ = ~pi0 & new_n815_;
  assign new_n817_ = px1 & new_n349_;
  assign new_n818_ = ~pi0 & new_n817_;
  assign new_n819_ = ~new_n812_ & ~new_n816_;
  assign pq4 = new_n818_ | ~new_n819_;
  assign new_n821_ = pr2 & new_n551_;
  assign new_n822_ = new_n177_ & new_n821_;
  assign new_n823_ = pn2 & new_n822_;
  assign new_n824_ = ~pi0 & ~pv2;
  assign new_n825_ = ~pf0 & ~pi0;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = ~new_n384_ & ~new_n823_;
  assign pv3 = new_n826_ | ~new_n827_;
  assign new_n829_ = pt & ~new_n333_;
  assign new_n830_ = new_n335_ & new_n829_;
  assign new_n831_ = pg0 & new_n830_;
  assign new_n832_ = pe1 & pz1;
  assign new_n833_ = ~pm0 & new_n832_;
  assign new_n834_ = new_n342_ & new_n833_;
  assign new_n835_ = ~pi0 & new_n834_;
  assign new_n836_ = py1 & new_n349_;
  assign new_n837_ = ~pi0 & new_n836_;
  assign new_n838_ = ~new_n831_ & ~new_n835_;
  assign pr4 = new_n837_ | ~new_n838_;
  assign pu3 = pa1 & ~pi0;
  assign new_n841_ = pu & ~new_n333_;
  assign new_n842_ = new_n335_ & new_n841_;
  assign new_n843_ = pg0 & new_n842_;
  assign new_n844_ = pa2 & pe1;
  assign new_n845_ = ~pm0 & new_n844_;
  assign new_n846_ = new_n342_ & new_n845_;
  assign new_n847_ = ~pi0 & new_n846_;
  assign new_n848_ = pz1 & new_n349_;
  assign new_n849_ = ~pi0 & new_n848_;
  assign new_n850_ = ~new_n843_ & ~new_n847_;
  assign ps4 = new_n849_ | ~new_n850_;
  assign pt3 = ~pi0 & pz0;
  assign new_n853_ = ~pc1 & pg1;
  assign new_n854_ = ~new_n187_ & new_n853_;
  assign new_n855_ = ~pe1 & new_n853_;
  assign new_n856_ = pp0 & new_n853_;
  assign new_n857_ = pn2 & new_n853_;
  assign new_n858_ = pp0 & new_n195_;
  assign new_n859_ = ~new_n196_ & ~new_n854_;
  assign new_n860_ = ~new_n855_ & ~new_n856_;
  assign new_n861_ = new_n859_ & new_n860_;
  assign new_n862_ = ~new_n201_ & ~new_n858_;
  assign new_n863_ = ~new_n200_ & ~new_n857_;
  assign new_n864_ = new_n862_ & new_n863_;
  assign pz3 = ~new_n861_ | ~new_n864_;
  assign new_n866_ = ~pc1 & pf1;
  assign new_n867_ = ~new_n187_ & new_n866_;
  assign new_n868_ = ~pe1 & new_n866_;
  assign new_n869_ = po0 & new_n866_;
  assign new_n870_ = pn2 & new_n866_;
  assign new_n871_ = po0 & new_n195_;
  assign new_n872_ = ~new_n196_ & ~new_n867_;
  assign new_n873_ = ~new_n868_ & ~new_n869_;
  assign new_n874_ = new_n872_ & new_n873_;
  assign new_n875_ = ~new_n201_ & ~new_n871_;
  assign new_n876_ = ~new_n200_ & ~new_n870_;
  assign new_n877_ = new_n875_ & new_n876_;
  assign py3 = ~new_n874_ | ~new_n877_;
  assign new_n879_ = pl2 & new_n212_;
  assign new_n880_ = ~pc1 & new_n879_;
  assign new_n881_ = ~new_n669_ & ~new_n880_;
  assign px3 = new_n650_ | ~new_n881_;
  assign new_n883_ = pz & ~new_n333_;
  assign new_n884_ = new_n335_ & new_n883_;
  assign new_n885_ = pg0 & new_n884_;
  assign new_n886_ = pe1 & pf2;
  assign new_n887_ = ~pm0 & new_n886_;
  assign new_n888_ = new_n342_ & new_n887_;
  assign new_n889_ = ~pi0 & new_n888_;
  assign new_n890_ = pe2 & new_n349_;
  assign new_n891_ = ~pi0 & new_n890_;
  assign new_n892_ = ~new_n885_ & ~new_n889_;
  assign px4 = new_n891_ | ~new_n892_;
  assign new_n894_ = pa0 & ~new_n333_;
  assign new_n895_ = new_n335_ & new_n894_;
  assign new_n896_ = pg0 & new_n895_;
  assign new_n897_ = pe1 & pg2;
  assign new_n898_ = ~pm0 & new_n897_;
  assign new_n899_ = new_n342_ & new_n898_;
  assign new_n900_ = ~pi0 & new_n899_;
  assign new_n901_ = pf2 & new_n349_;
  assign new_n902_ = ~pi0 & new_n901_;
  assign new_n903_ = ~new_n896_ & ~new_n900_;
  assign py4 = new_n902_ | ~new_n903_;
  assign new_n905_ = pb0 & ~new_n333_;
  assign new_n906_ = new_n335_ & new_n905_;
  assign new_n907_ = pg0 & new_n906_;
  assign new_n908_ = pe1 & ph2;
  assign new_n909_ = ~pm0 & new_n908_;
  assign new_n910_ = new_n342_ & new_n909_;
  assign new_n911_ = ~pi0 & new_n910_;
  assign new_n912_ = pg2 & new_n349_;
  assign new_n913_ = ~pi0 & new_n912_;
  assign new_n914_ = ~new_n907_ & ~new_n911_;
  assign pz4 = new_n913_ | ~new_n914_;
  assign pb3 = ~pk1;
  assign pa3 = ~pj1;
  assign pw2 = ~pf1;
  assign pz2 = ~pi1;
  assign px2 = ~pg1;
  assign py2 = ~ph1;
endmodule

