// Benchmark "top" written by ABC on Thu Oct  8 22:52:00 2020

module top ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3122_, new_n3123_, new_n3125_, new_n3126_, new_n3128_, new_n3129_,
    new_n3131_, new_n3132_, new_n3134_, new_n3135_, new_n3137_, new_n3138_,
    new_n3140_, new_n3141_, new_n3143_, new_n3144_, new_n3146_, new_n3147_,
    new_n3149_, new_n3150_, new_n3152_, new_n3153_, new_n3155_, new_n3156_,
    new_n3158_, new_n3159_, new_n3161_, new_n3162_, new_n3164_, new_n3165_,
    new_n3167_, new_n3168_, new_n3170_, new_n3171_, new_n3173_, new_n3174_,
    new_n3176_, new_n3177_, new_n3179_, new_n3180_, new_n3182_, new_n3183_,
    new_n3185_, new_n3186_, new_n3188_, new_n3189_, new_n3191_, new_n3192_,
    new_n3194_, new_n3195_, new_n3197_, new_n3198_, new_n3200_, new_n3201_,
    new_n3203_, new_n3204_, new_n3206_, new_n3207_, new_n3209_, new_n3210_,
    new_n3212_, new_n3213_, new_n3215_, new_n3216_, new_n3218_, new_n3219_,
    new_n3221_, new_n3222_, new_n3224_, new_n3225_, new_n3227_, new_n3228_,
    new_n3230_, new_n3231_, new_n3233_, new_n3234_, new_n3236_, new_n3237_,
    new_n3239_, new_n3240_, new_n3242_, new_n3243_, new_n3245_, new_n3246_,
    new_n3248_, new_n3249_, new_n3251_, new_n3252_, new_n3254_, new_n3255_,
    new_n3257_, new_n3258_, new_n3260_, new_n3261_, new_n3263_, new_n3264_,
    new_n3266_, new_n3267_, new_n3269_, new_n3270_, new_n3272_, new_n3273_,
    new_n3275_, new_n3276_, new_n3278_, new_n3279_, new_n3281_, new_n3282_,
    new_n3284_, new_n3285_, new_n3287_, new_n3288_, new_n3290_, new_n3291_,
    new_n3293_, new_n3294_, new_n3296_, new_n3297_, new_n3299_, new_n3300_,
    new_n3302_, new_n3303_, new_n3305_, new_n3306_, new_n3308_, new_n3309_,
    new_n3311_, new_n3312_, new_n3314_, new_n3315_, new_n3317_, new_n3318_,
    new_n3320_, new_n3321_, new_n3323_, new_n3324_, new_n3326_, new_n3327_,
    new_n3329_, new_n3330_, new_n3332_, new_n3333_, new_n3335_, new_n3336_,
    new_n3338_, new_n3339_, new_n3341_, new_n3342_, new_n3344_, new_n3345_,
    new_n3347_, new_n3348_, new_n3350_, new_n3351_, new_n3353_, new_n3354_,
    new_n3356_, new_n3357_, new_n3359_, new_n3360_, new_n3362_, new_n3363_,
    new_n3365_, new_n3366_, new_n3368_, new_n3369_, new_n3371_, new_n3372_,
    new_n3374_, new_n3375_, new_n3377_, new_n3378_, new_n3380_, new_n3381_,
    new_n3383_, new_n3384_, new_n3386_, new_n3387_, new_n3389_, new_n3390_,
    new_n3392_, new_n3393_, new_n3395_, new_n3396_, new_n3398_, new_n3399_,
    new_n3401_, new_n3402_, new_n3404_, new_n3405_, new_n3407_, new_n3408_,
    new_n3410_, new_n3411_, new_n3413_, new_n3414_, new_n3416_, new_n3417_,
    new_n3419_, new_n3420_, new_n3422_, new_n3423_, new_n3425_, new_n3426_,
    new_n3428_, new_n3429_, new_n3431_, new_n3432_, new_n3434_, new_n3435_,
    new_n3437_, new_n3438_, new_n3440_, new_n3441_, new_n3443_, new_n3444_,
    new_n3446_, new_n3447_, new_n3449_, new_n3450_, new_n3452_, new_n3453_,
    new_n3455_, new_n3456_, new_n3458_, new_n3459_, new_n3461_, new_n3462_,
    new_n3464_, new_n3465_, new_n3467_, new_n3468_, new_n3470_, new_n3471_,
    new_n3473_, new_n3474_, new_n3476_, new_n3477_, new_n3479_, new_n3480_,
    new_n3482_, new_n3483_, new_n3485_, new_n3486_, new_n3488_, new_n3489_,
    new_n3491_, new_n3492_, new_n3494_, new_n3495_, new_n3497_, new_n3498_,
    new_n3500_, new_n3501_, new_n3503_, new_n3505_, new_n3506_;
  assign new_n643_ = \in2[119]  & ~\in3[119] ;
  assign new_n644_ = ~\in2[119]  & \in3[119] ;
  assign new_n645_ = ~\in2[118]  & \in3[118] ;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = ~\in2[117]  & \in3[117] ;
  assign new_n648_ = \in2[116]  & ~\in3[116] ;
  assign new_n649_ = ~new_n647_ & new_n648_;
  assign new_n650_ = \in2[117]  & ~\in3[117] ;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = new_n646_ & ~new_n651_;
  assign new_n653_ = ~\in3[118]  & ~new_n644_;
  assign new_n654_ = \in2[118]  & new_n653_;
  assign new_n655_ = ~\in2[112]  & \in3[112] ;
  assign new_n656_ = ~\in2[115]  & \in3[115] ;
  assign new_n657_ = ~\in2[114]  & \in3[114] ;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = ~\in2[113]  & \in3[113] ;
  assign new_n660_ = \in2[111]  & ~\in3[111] ;
  assign new_n661_ = ~\in2[111]  & \in3[111] ;
  assign new_n662_ = ~\in2[110]  & \in3[110] ;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign new_n664_ = ~\in2[109]  & \in3[109] ;
  assign new_n665_ = \in2[108]  & ~\in3[108] ;
  assign new_n666_ = ~new_n664_ & new_n665_;
  assign new_n667_ = \in2[109]  & ~\in3[109] ;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = new_n663_ & ~new_n668_;
  assign new_n670_ = ~\in3[110]  & ~new_n661_;
  assign new_n671_ = \in2[110]  & new_n670_;
  assign new_n672_ = \in2[103]  & ~\in3[103] ;
  assign new_n673_ = ~\in2[103]  & \in3[103] ;
  assign new_n674_ = ~\in2[102]  & \in3[102] ;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~\in2[101]  & \in3[101] ;
  assign new_n677_ = \in2[100]  & ~\in3[100] ;
  assign new_n678_ = ~new_n676_ & new_n677_;
  assign new_n679_ = \in2[101]  & ~\in3[101] ;
  assign new_n680_ = ~new_n678_ & ~new_n679_;
  assign new_n681_ = new_n675_ & ~new_n680_;
  assign new_n682_ = ~\in3[102]  & ~new_n673_;
  assign new_n683_ = \in2[102]  & new_n682_;
  assign new_n684_ = ~\in2[96]  & \in3[96] ;
  assign new_n685_ = ~\in2[99]  & \in3[99] ;
  assign new_n686_ = ~\in2[98]  & \in3[98] ;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign new_n688_ = ~\in2[97]  & \in3[97] ;
  assign new_n689_ = \in2[95]  & ~\in3[95] ;
  assign new_n690_ = ~\in2[95]  & \in3[95] ;
  assign new_n691_ = ~\in2[94]  & \in3[94] ;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = ~\in2[93]  & \in3[93] ;
  assign new_n694_ = \in2[92]  & ~\in3[92] ;
  assign new_n695_ = ~new_n693_ & new_n694_;
  assign new_n696_ = \in2[93]  & ~\in3[93] ;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = new_n692_ & ~new_n697_;
  assign new_n699_ = ~\in3[94]  & ~new_n690_;
  assign new_n700_ = \in2[94]  & new_n699_;
  assign new_n701_ = \in2[87]  & ~\in3[87] ;
  assign new_n702_ = ~\in2[87]  & \in3[87] ;
  assign new_n703_ = ~\in2[86]  & \in3[86] ;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = ~\in2[85]  & \in3[85] ;
  assign new_n706_ = \in2[84]  & ~\in3[84] ;
  assign new_n707_ = ~new_n705_ & new_n706_;
  assign new_n708_ = \in2[85]  & ~\in3[85] ;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = new_n704_ & ~new_n709_;
  assign new_n711_ = ~\in3[86]  & ~new_n702_;
  assign new_n712_ = \in2[86]  & new_n711_;
  assign new_n713_ = ~\in2[80]  & \in3[80] ;
  assign new_n714_ = ~\in2[83]  & \in3[83] ;
  assign new_n715_ = ~\in2[82]  & \in3[82] ;
  assign new_n716_ = ~new_n714_ & ~new_n715_;
  assign new_n717_ = ~\in2[81]  & \in3[81] ;
  assign new_n718_ = \in2[79]  & ~\in3[79] ;
  assign new_n719_ = ~\in2[79]  & \in3[79] ;
  assign new_n720_ = ~\in2[78]  & \in3[78] ;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = ~\in2[77]  & \in3[77] ;
  assign new_n723_ = \in2[76]  & ~\in3[76] ;
  assign new_n724_ = ~new_n722_ & new_n723_;
  assign new_n725_ = \in2[77]  & ~\in3[77] ;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = new_n721_ & ~new_n726_;
  assign new_n728_ = ~\in3[78]  & ~new_n719_;
  assign new_n729_ = \in2[78]  & new_n728_;
  assign new_n730_ = \in2[71]  & ~\in3[71] ;
  assign new_n731_ = ~\in2[71]  & \in3[71] ;
  assign new_n732_ = ~\in2[70]  & \in3[70] ;
  assign new_n733_ = ~new_n731_ & ~new_n732_;
  assign new_n734_ = ~\in2[69]  & \in3[69] ;
  assign new_n735_ = \in2[68]  & ~\in3[68] ;
  assign new_n736_ = ~new_n734_ & new_n735_;
  assign new_n737_ = \in2[69]  & ~\in3[69] ;
  assign new_n738_ = ~new_n736_ & ~new_n737_;
  assign new_n739_ = new_n733_ & ~new_n738_;
  assign new_n740_ = ~\in3[70]  & ~new_n731_;
  assign new_n741_ = \in2[70]  & new_n740_;
  assign new_n742_ = ~\in2[67]  & \in3[67] ;
  assign new_n743_ = ~\in2[66]  & \in3[66] ;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = ~\in2[65]  & \in3[65] ;
  assign new_n746_ = \in2[63]  & ~\in3[63] ;
  assign new_n747_ = ~\in2[63]  & \in3[63] ;
  assign new_n748_ = ~\in2[62]  & \in3[62] ;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign new_n750_ = ~\in2[60]  & \in3[60] ;
  assign new_n751_ = ~\in2[61]  & \in3[61] ;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = new_n749_ & new_n752_;
  assign new_n754_ = \in2[59]  & ~\in3[59] ;
  assign new_n755_ = ~\in2[59]  & \in3[59] ;
  assign new_n756_ = ~\in2[58]  & \in3[58] ;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = ~\in2[57]  & \in3[57] ;
  assign new_n759_ = \in2[56]  & ~\in3[56] ;
  assign new_n760_ = ~new_n758_ & new_n759_;
  assign new_n761_ = \in2[57]  & ~\in3[57] ;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = \in2[58]  & ~\in3[58] ;
  assign new_n764_ = new_n762_ & ~new_n763_;
  assign new_n765_ = new_n757_ & ~new_n764_;
  assign new_n766_ = ~new_n754_ & ~new_n765_;
  assign new_n767_ = new_n753_ & ~new_n766_;
  assign new_n768_ = \in2[60]  & ~\in3[60] ;
  assign new_n769_ = ~new_n751_ & new_n768_;
  assign new_n770_ = \in2[61]  & ~\in3[61] ;
  assign new_n771_ = ~new_n769_ & ~new_n770_;
  assign new_n772_ = new_n749_ & ~new_n771_;
  assign new_n773_ = ~\in3[62]  & ~new_n747_;
  assign new_n774_ = \in2[62]  & new_n773_;
  assign new_n775_ = \in2[47]  & ~\in3[47] ;
  assign new_n776_ = ~\in2[47]  & \in3[47] ;
  assign new_n777_ = ~\in2[46]  & \in3[46] ;
  assign new_n778_ = ~new_n776_ & ~new_n777_;
  assign new_n779_ = ~\in2[44]  & \in3[44] ;
  assign new_n780_ = ~\in2[45]  & \in3[45] ;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = new_n778_ & new_n781_;
  assign new_n783_ = \in2[43]  & ~\in3[43] ;
  assign new_n784_ = ~\in2[43]  & \in3[43] ;
  assign new_n785_ = ~\in2[42]  & \in3[42] ;
  assign new_n786_ = ~new_n784_ & ~new_n785_;
  assign new_n787_ = ~\in2[41]  & \in3[41] ;
  assign new_n788_ = \in2[40]  & ~\in3[40] ;
  assign new_n789_ = ~new_n787_ & new_n788_;
  assign new_n790_ = \in2[41]  & ~\in3[41] ;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = \in2[42]  & ~\in3[42] ;
  assign new_n793_ = new_n791_ & ~new_n792_;
  assign new_n794_ = new_n786_ & ~new_n793_;
  assign new_n795_ = ~new_n783_ & ~new_n794_;
  assign new_n796_ = new_n782_ & ~new_n795_;
  assign new_n797_ = \in2[44]  & ~\in3[44] ;
  assign new_n798_ = ~new_n780_ & new_n797_;
  assign new_n799_ = \in2[45]  & ~\in3[45] ;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = new_n778_ & ~new_n800_;
  assign new_n802_ = ~\in3[46]  & ~new_n776_;
  assign new_n803_ = \in2[46]  & new_n802_;
  assign new_n804_ = ~\in2[32]  & \in3[32] ;
  assign new_n805_ = ~\in2[31]  & \in3[31] ;
  assign new_n806_ = ~\in2[30]  & \in3[30] ;
  assign new_n807_ = ~\in2[29]  & \in3[29] ;
  assign new_n808_ = ~\in2[28]  & \in3[28] ;
  assign new_n809_ = ~\in2[27]  & \in3[27] ;
  assign new_n810_ = ~\in2[26]  & \in3[26] ;
  assign new_n811_ = ~\in2[23]  & \in3[23] ;
  assign new_n812_ = ~\in2[22]  & \in3[22] ;
  assign new_n813_ = ~\in2[21]  & \in3[21] ;
  assign new_n814_ = ~\in2[20]  & \in3[20] ;
  assign new_n815_ = ~\in2[19]  & \in3[19] ;
  assign new_n816_ = ~\in2[18]  & \in3[18] ;
  assign new_n817_ = ~\in2[15]  & \in3[15] ;
  assign new_n818_ = ~\in2[14]  & \in3[14] ;
  assign new_n819_ = ~\in2[13]  & \in3[13] ;
  assign new_n820_ = ~\in2[12]  & \in3[12] ;
  assign new_n821_ = ~\in2[11]  & \in3[11] ;
  assign new_n822_ = ~\in2[10]  & \in3[10] ;
  assign new_n823_ = ~\in2[7]  & \in3[7] ;
  assign new_n824_ = ~\in2[6]  & \in3[6] ;
  assign new_n825_ = ~\in2[3]  & \in3[3] ;
  assign new_n826_ = \in2[0]  & ~\in3[0] ;
  assign new_n827_ = \in2[1]  & new_n826_;
  assign new_n828_ = \in3[1]  & ~new_n827_;
  assign new_n829_ = ~\in2[2]  & \in3[2] ;
  assign new_n830_ = ~\in2[1]  & ~new_n826_;
  assign new_n831_ = ~new_n829_ & ~new_n830_;
  assign new_n832_ = ~new_n828_ & new_n831_;
  assign new_n833_ = \in2[2]  & ~\in3[2] ;
  assign new_n834_ = ~new_n832_ & ~new_n833_;
  assign new_n835_ = ~new_n825_ & ~new_n834_;
  assign new_n836_ = \in2[3]  & ~\in3[3] ;
  assign new_n837_ = ~new_n835_ & ~new_n836_;
  assign new_n838_ = ~\in2[4]  & new_n837_;
  assign new_n839_ = ~\in3[4]  & ~new_n838_;
  assign new_n840_ = \in2[4]  & ~new_n837_;
  assign new_n841_ = ~new_n839_ & ~new_n840_;
  assign new_n842_ = ~\in2[5]  & new_n841_;
  assign new_n843_ = ~\in3[5]  & ~new_n842_;
  assign new_n844_ = \in2[5]  & ~new_n841_;
  assign new_n845_ = ~new_n843_ & ~new_n844_;
  assign new_n846_ = ~new_n824_ & ~new_n845_;
  assign new_n847_ = \in2[6]  & ~\in3[6] ;
  assign new_n848_ = ~new_n846_ & ~new_n847_;
  assign new_n849_ = ~new_n823_ & ~new_n848_;
  assign new_n850_ = \in2[7]  & ~\in3[7] ;
  assign new_n851_ = ~new_n849_ & ~new_n850_;
  assign new_n852_ = ~\in2[8]  & new_n851_;
  assign new_n853_ = ~\in3[8]  & ~new_n852_;
  assign new_n854_ = \in2[8]  & ~new_n851_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign new_n856_ = ~\in2[9]  & new_n855_;
  assign new_n857_ = ~\in3[9]  & ~new_n856_;
  assign new_n858_ = \in2[9]  & ~new_n855_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~new_n822_ & ~new_n859_;
  assign new_n861_ = \in2[10]  & ~\in3[10] ;
  assign new_n862_ = ~new_n860_ & ~new_n861_;
  assign new_n863_ = ~new_n821_ & ~new_n862_;
  assign new_n864_ = \in2[11]  & ~\in3[11] ;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = ~new_n820_ & ~new_n865_;
  assign new_n867_ = \in2[12]  & ~\in3[12] ;
  assign new_n868_ = ~new_n866_ & ~new_n867_;
  assign new_n869_ = ~new_n819_ & ~new_n868_;
  assign new_n870_ = \in2[13]  & ~\in3[13] ;
  assign new_n871_ = ~new_n869_ & ~new_n870_;
  assign new_n872_ = ~new_n818_ & ~new_n871_;
  assign new_n873_ = \in2[14]  & ~\in3[14] ;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = ~new_n817_ & ~new_n874_;
  assign new_n876_ = \in2[15]  & ~\in3[15] ;
  assign new_n877_ = ~new_n875_ & ~new_n876_;
  assign new_n878_ = ~\in2[16]  & new_n877_;
  assign new_n879_ = ~\in3[16]  & ~new_n878_;
  assign new_n880_ = \in2[16]  & ~new_n877_;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = ~\in2[17]  & new_n881_;
  assign new_n883_ = ~\in3[17]  & ~new_n882_;
  assign new_n884_ = \in2[17]  & ~new_n881_;
  assign new_n885_ = ~new_n883_ & ~new_n884_;
  assign new_n886_ = ~new_n816_ & ~new_n885_;
  assign new_n887_ = \in2[18]  & ~\in3[18] ;
  assign new_n888_ = ~new_n886_ & ~new_n887_;
  assign new_n889_ = ~new_n815_ & ~new_n888_;
  assign new_n890_ = \in2[19]  & ~\in3[19] ;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = ~new_n814_ & ~new_n891_;
  assign new_n893_ = \in2[20]  & ~\in3[20] ;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = ~new_n813_ & ~new_n894_;
  assign new_n896_ = \in2[21]  & ~\in3[21] ;
  assign new_n897_ = ~new_n895_ & ~new_n896_;
  assign new_n898_ = ~new_n812_ & ~new_n897_;
  assign new_n899_ = \in2[22]  & ~\in3[22] ;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~new_n811_ & ~new_n900_;
  assign new_n902_ = \in2[23]  & ~\in3[23] ;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = ~\in2[24]  & new_n903_;
  assign new_n905_ = ~\in3[24]  & ~new_n904_;
  assign new_n906_ = \in2[24]  & ~new_n903_;
  assign new_n907_ = ~new_n905_ & ~new_n906_;
  assign new_n908_ = ~\in2[25]  & new_n907_;
  assign new_n909_ = ~\in3[25]  & ~new_n908_;
  assign new_n910_ = \in2[25]  & ~new_n907_;
  assign new_n911_ = ~new_n909_ & ~new_n910_;
  assign new_n912_ = ~new_n810_ & ~new_n911_;
  assign new_n913_ = \in2[26]  & ~\in3[26] ;
  assign new_n914_ = ~new_n912_ & ~new_n913_;
  assign new_n915_ = ~new_n809_ & ~new_n914_;
  assign new_n916_ = \in2[27]  & ~\in3[27] ;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = ~new_n808_ & ~new_n917_;
  assign new_n919_ = \in2[28]  & ~\in3[28] ;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~new_n807_ & ~new_n920_;
  assign new_n922_ = \in2[29]  & ~\in3[29] ;
  assign new_n923_ = ~new_n921_ & ~new_n922_;
  assign new_n924_ = ~new_n806_ & ~new_n923_;
  assign new_n925_ = \in2[30]  & ~\in3[30] ;
  assign new_n926_ = ~new_n924_ & ~new_n925_;
  assign new_n927_ = ~new_n805_ & ~new_n926_;
  assign new_n928_ = \in2[31]  & ~\in3[31] ;
  assign new_n929_ = ~new_n927_ & ~new_n928_;
  assign new_n930_ = ~\in2[39]  & \in3[39] ;
  assign new_n931_ = ~\in2[38]  & \in3[38] ;
  assign new_n932_ = ~new_n930_ & ~new_n931_;
  assign new_n933_ = ~\in2[36]  & \in3[36] ;
  assign new_n934_ = ~\in2[37]  & \in3[37] ;
  assign new_n935_ = ~new_n933_ & ~new_n934_;
  assign new_n936_ = new_n932_ & new_n935_;
  assign new_n937_ = ~\in2[33]  & \in3[33] ;
  assign new_n938_ = ~\in2[35]  & \in3[35] ;
  assign new_n939_ = ~\in2[34]  & \in3[34] ;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = ~new_n937_ & new_n940_;
  assign new_n942_ = new_n936_ & new_n941_;
  assign new_n943_ = ~new_n929_ & new_n942_;
  assign new_n944_ = ~new_n804_ & new_n943_;
  assign new_n945_ = \in2[39]  & ~\in3[39] ;
  assign new_n946_ = \in2[36]  & ~\in3[36] ;
  assign new_n947_ = ~new_n934_ & new_n946_;
  assign new_n948_ = \in2[37]  & ~\in3[37] ;
  assign new_n949_ = ~new_n947_ & ~new_n948_;
  assign new_n950_ = new_n932_ & ~new_n949_;
  assign new_n951_ = ~\in3[38]  & ~new_n930_;
  assign new_n952_ = \in2[38]  & new_n951_;
  assign new_n953_ = \in2[35]  & ~\in3[35] ;
  assign new_n954_ = ~\in3[32]  & ~new_n937_;
  assign new_n955_ = \in2[32]  & new_n954_;
  assign new_n956_ = \in2[33]  & ~\in3[33] ;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = \in2[34]  & ~\in3[34] ;
  assign new_n959_ = new_n957_ & ~new_n958_;
  assign new_n960_ = new_n940_ & ~new_n959_;
  assign new_n961_ = ~new_n953_ & ~new_n960_;
  assign new_n962_ = new_n936_ & ~new_n961_;
  assign new_n963_ = ~new_n952_ & ~new_n962_;
  assign new_n964_ = ~new_n950_ & new_n963_;
  assign new_n965_ = ~new_n945_ & new_n964_;
  assign new_n966_ = ~new_n944_ & new_n965_;
  assign new_n967_ = ~\in2[40]  & \in3[40] ;
  assign new_n968_ = ~new_n787_ & ~new_n967_;
  assign new_n969_ = new_n786_ & new_n968_;
  assign new_n970_ = new_n782_ & new_n969_;
  assign new_n971_ = ~new_n966_ & new_n970_;
  assign new_n972_ = ~new_n803_ & ~new_n971_;
  assign new_n973_ = ~new_n801_ & new_n972_;
  assign new_n974_ = ~new_n796_ & new_n973_;
  assign new_n975_ = ~new_n775_ & new_n974_;
  assign new_n976_ = ~\in2[48]  & \in3[48] ;
  assign new_n977_ = ~\in2[55]  & \in3[55] ;
  assign new_n978_ = ~\in2[54]  & \in3[54] ;
  assign new_n979_ = ~new_n977_ & ~new_n978_;
  assign new_n980_ = ~\in2[53]  & \in3[53] ;
  assign new_n981_ = ~\in2[52]  & \in3[52] ;
  assign new_n982_ = ~new_n980_ & ~new_n981_;
  assign new_n983_ = new_n979_ & new_n982_;
  assign new_n984_ = ~\in2[49]  & \in3[49] ;
  assign new_n985_ = ~\in2[51]  & \in3[51] ;
  assign new_n986_ = ~\in2[50]  & \in3[50] ;
  assign new_n987_ = ~new_n985_ & ~new_n986_;
  assign new_n988_ = ~new_n984_ & new_n987_;
  assign new_n989_ = new_n983_ & new_n988_;
  assign new_n990_ = ~new_n976_ & new_n989_;
  assign new_n991_ = ~new_n975_ & new_n990_;
  assign new_n992_ = \in2[55]  & ~\in3[55] ;
  assign new_n993_ = \in2[51]  & ~\in3[51] ;
  assign new_n994_ = ~\in3[48]  & ~new_n984_;
  assign new_n995_ = \in2[48]  & new_n994_;
  assign new_n996_ = \in2[49]  & ~\in3[49] ;
  assign new_n997_ = ~new_n995_ & ~new_n996_;
  assign new_n998_ = \in2[50]  & ~\in3[50] ;
  assign new_n999_ = new_n997_ & ~new_n998_;
  assign new_n1000_ = new_n987_ & ~new_n999_;
  assign new_n1001_ = ~new_n993_ & ~new_n1000_;
  assign new_n1002_ = new_n983_ & ~new_n1001_;
  assign new_n1003_ = \in2[52]  & ~\in3[52] ;
  assign new_n1004_ = ~new_n980_ & new_n1003_;
  assign new_n1005_ = \in2[53]  & ~\in3[53] ;
  assign new_n1006_ = ~new_n1004_ & ~new_n1005_;
  assign new_n1007_ = \in2[54]  & ~\in3[54] ;
  assign new_n1008_ = new_n1006_ & ~new_n1007_;
  assign new_n1009_ = new_n979_ & ~new_n1008_;
  assign new_n1010_ = ~new_n1002_ & ~new_n1009_;
  assign new_n1011_ = ~new_n992_ & new_n1010_;
  assign new_n1012_ = ~new_n991_ & new_n1011_;
  assign new_n1013_ = ~\in2[56]  & \in3[56] ;
  assign new_n1014_ = ~new_n758_ & ~new_n1013_;
  assign new_n1015_ = new_n753_ & new_n1014_;
  assign new_n1016_ = new_n757_ & new_n1015_;
  assign new_n1017_ = ~new_n1012_ & new_n1016_;
  assign new_n1018_ = ~new_n774_ & ~new_n1017_;
  assign new_n1019_ = ~new_n772_ & new_n1018_;
  assign new_n1020_ = ~new_n767_ & new_n1019_;
  assign new_n1021_ = ~new_n746_ & new_n1020_;
  assign new_n1022_ = ~\in2[64]  & \in3[64] ;
  assign new_n1023_ = ~new_n1021_ & ~new_n1022_;
  assign new_n1024_ = ~new_n745_ & new_n1023_;
  assign new_n1025_ = new_n744_ & new_n1024_;
  assign new_n1026_ = \in2[67]  & ~\in3[67] ;
  assign new_n1027_ = \in2[64]  & ~\in3[64] ;
  assign new_n1028_ = ~new_n745_ & new_n1027_;
  assign new_n1029_ = \in2[65]  & ~\in3[65] ;
  assign new_n1030_ = ~new_n1028_ & ~new_n1029_;
  assign new_n1031_ = \in2[66]  & ~\in3[66] ;
  assign new_n1032_ = new_n1030_ & ~new_n1031_;
  assign new_n1033_ = new_n744_ & ~new_n1032_;
  assign new_n1034_ = ~new_n1026_ & ~new_n1033_;
  assign new_n1035_ = ~new_n1025_ & new_n1034_;
  assign new_n1036_ = ~\in2[68]  & \in3[68] ;
  assign new_n1037_ = ~new_n734_ & ~new_n1036_;
  assign new_n1038_ = new_n733_ & new_n1037_;
  assign new_n1039_ = ~new_n1035_ & new_n1038_;
  assign new_n1040_ = ~new_n741_ & ~new_n1039_;
  assign new_n1041_ = ~new_n739_ & new_n1040_;
  assign new_n1042_ = ~new_n730_ & new_n1041_;
  assign new_n1043_ = ~\in2[75]  & \in3[75] ;
  assign new_n1044_ = ~\in2[74]  & \in3[74] ;
  assign new_n1045_ = ~new_n1043_ & ~new_n1044_;
  assign new_n1046_ = ~\in2[73]  & \in3[73] ;
  assign new_n1047_ = ~\in2[72]  & \in3[72] ;
  assign new_n1048_ = ~new_n1046_ & ~new_n1047_;
  assign new_n1049_ = new_n1045_ & new_n1048_;
  assign new_n1050_ = ~new_n1042_ & new_n1049_;
  assign new_n1051_ = \in2[75]  & ~\in3[75] ;
  assign new_n1052_ = \in2[72]  & ~\in3[72] ;
  assign new_n1053_ = ~new_n1046_ & new_n1052_;
  assign new_n1054_ = \in2[73]  & ~\in3[73] ;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = \in2[74]  & ~\in3[74] ;
  assign new_n1057_ = new_n1055_ & ~new_n1056_;
  assign new_n1058_ = new_n1045_ & ~new_n1057_;
  assign new_n1059_ = ~new_n1051_ & ~new_n1058_;
  assign new_n1060_ = ~new_n1050_ & new_n1059_;
  assign new_n1061_ = ~\in2[76]  & \in3[76] ;
  assign new_n1062_ = ~new_n722_ & ~new_n1061_;
  assign new_n1063_ = new_n721_ & new_n1062_;
  assign new_n1064_ = ~new_n1060_ & new_n1063_;
  assign new_n1065_ = ~new_n729_ & ~new_n1064_;
  assign new_n1066_ = ~new_n727_ & new_n1065_;
  assign new_n1067_ = ~new_n718_ & new_n1066_;
  assign new_n1068_ = ~new_n717_ & ~new_n1067_;
  assign new_n1069_ = new_n716_ & new_n1068_;
  assign new_n1070_ = ~new_n713_ & new_n1069_;
  assign new_n1071_ = \in2[83]  & ~\in3[83] ;
  assign new_n1072_ = ~\in3[80]  & ~new_n717_;
  assign new_n1073_ = \in2[80]  & new_n1072_;
  assign new_n1074_ = \in2[81]  & ~\in3[81] ;
  assign new_n1075_ = ~new_n1073_ & ~new_n1074_;
  assign new_n1076_ = \in2[82]  & ~\in3[82] ;
  assign new_n1077_ = new_n1075_ & ~new_n1076_;
  assign new_n1078_ = new_n716_ & ~new_n1077_;
  assign new_n1079_ = ~new_n1071_ & ~new_n1078_;
  assign new_n1080_ = ~new_n1070_ & new_n1079_;
  assign new_n1081_ = ~\in2[84]  & \in3[84] ;
  assign new_n1082_ = ~new_n705_ & ~new_n1081_;
  assign new_n1083_ = new_n704_ & new_n1082_;
  assign new_n1084_ = ~new_n1080_ & new_n1083_;
  assign new_n1085_ = ~new_n712_ & ~new_n1084_;
  assign new_n1086_ = ~new_n710_ & new_n1085_;
  assign new_n1087_ = ~new_n701_ & new_n1086_;
  assign new_n1088_ = ~\in2[91]  & \in3[91] ;
  assign new_n1089_ = ~\in2[90]  & \in3[90] ;
  assign new_n1090_ = ~new_n1088_ & ~new_n1089_;
  assign new_n1091_ = ~\in2[89]  & \in3[89] ;
  assign new_n1092_ = ~\in2[88]  & \in3[88] ;
  assign new_n1093_ = ~new_n1091_ & ~new_n1092_;
  assign new_n1094_ = new_n1090_ & new_n1093_;
  assign new_n1095_ = ~new_n1087_ & new_n1094_;
  assign new_n1096_ = \in2[91]  & ~\in3[91] ;
  assign new_n1097_ = \in2[88]  & ~\in3[88] ;
  assign new_n1098_ = ~new_n1091_ & new_n1097_;
  assign new_n1099_ = \in2[89]  & ~\in3[89] ;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = \in2[90]  & ~\in3[90] ;
  assign new_n1102_ = new_n1100_ & ~new_n1101_;
  assign new_n1103_ = new_n1090_ & ~new_n1102_;
  assign new_n1104_ = ~new_n1096_ & ~new_n1103_;
  assign new_n1105_ = ~new_n1095_ & new_n1104_;
  assign new_n1106_ = ~\in2[92]  & \in3[92] ;
  assign new_n1107_ = ~new_n693_ & ~new_n1106_;
  assign new_n1108_ = new_n692_ & new_n1107_;
  assign new_n1109_ = ~new_n1105_ & new_n1108_;
  assign new_n1110_ = ~new_n700_ & ~new_n1109_;
  assign new_n1111_ = ~new_n698_ & new_n1110_;
  assign new_n1112_ = ~new_n689_ & new_n1111_;
  assign new_n1113_ = ~new_n688_ & ~new_n1112_;
  assign new_n1114_ = new_n687_ & new_n1113_;
  assign new_n1115_ = ~new_n684_ & new_n1114_;
  assign new_n1116_ = \in2[99]  & ~\in3[99] ;
  assign new_n1117_ = ~\in3[96]  & ~new_n688_;
  assign new_n1118_ = \in2[96]  & new_n1117_;
  assign new_n1119_ = \in2[97]  & ~\in3[97] ;
  assign new_n1120_ = ~new_n1118_ & ~new_n1119_;
  assign new_n1121_ = \in2[98]  & ~\in3[98] ;
  assign new_n1122_ = new_n1120_ & ~new_n1121_;
  assign new_n1123_ = new_n687_ & ~new_n1122_;
  assign new_n1124_ = ~new_n1116_ & ~new_n1123_;
  assign new_n1125_ = ~new_n1115_ & new_n1124_;
  assign new_n1126_ = ~\in2[100]  & \in3[100] ;
  assign new_n1127_ = ~new_n676_ & ~new_n1126_;
  assign new_n1128_ = new_n675_ & new_n1127_;
  assign new_n1129_ = ~new_n1125_ & new_n1128_;
  assign new_n1130_ = ~new_n683_ & ~new_n1129_;
  assign new_n1131_ = ~new_n681_ & new_n1130_;
  assign new_n1132_ = ~new_n672_ & new_n1131_;
  assign new_n1133_ = ~\in2[107]  & \in3[107] ;
  assign new_n1134_ = ~\in2[106]  & \in3[106] ;
  assign new_n1135_ = ~new_n1133_ & ~new_n1134_;
  assign new_n1136_ = ~\in2[105]  & \in3[105] ;
  assign new_n1137_ = ~\in2[104]  & \in3[104] ;
  assign new_n1138_ = ~new_n1136_ & ~new_n1137_;
  assign new_n1139_ = new_n1135_ & new_n1138_;
  assign new_n1140_ = ~new_n1132_ & new_n1139_;
  assign new_n1141_ = \in2[107]  & ~\in3[107] ;
  assign new_n1142_ = \in2[104]  & ~\in3[104] ;
  assign new_n1143_ = ~new_n1136_ & new_n1142_;
  assign new_n1144_ = \in2[105]  & ~\in3[105] ;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = \in2[106]  & ~\in3[106] ;
  assign new_n1147_ = new_n1145_ & ~new_n1146_;
  assign new_n1148_ = new_n1135_ & ~new_n1147_;
  assign new_n1149_ = ~new_n1141_ & ~new_n1148_;
  assign new_n1150_ = ~new_n1140_ & new_n1149_;
  assign new_n1151_ = ~\in2[108]  & \in3[108] ;
  assign new_n1152_ = ~new_n664_ & ~new_n1151_;
  assign new_n1153_ = new_n663_ & new_n1152_;
  assign new_n1154_ = ~new_n1150_ & new_n1153_;
  assign new_n1155_ = ~new_n671_ & ~new_n1154_;
  assign new_n1156_ = ~new_n669_ & new_n1155_;
  assign new_n1157_ = ~new_n660_ & new_n1156_;
  assign new_n1158_ = ~new_n659_ & ~new_n1157_;
  assign new_n1159_ = new_n658_ & new_n1158_;
  assign new_n1160_ = ~new_n655_ & new_n1159_;
  assign new_n1161_ = \in2[115]  & ~\in3[115] ;
  assign new_n1162_ = ~\in3[112]  & ~new_n659_;
  assign new_n1163_ = \in2[112]  & new_n1162_;
  assign new_n1164_ = \in2[113]  & ~\in3[113] ;
  assign new_n1165_ = ~new_n1163_ & ~new_n1164_;
  assign new_n1166_ = \in2[114]  & ~\in3[114] ;
  assign new_n1167_ = new_n1165_ & ~new_n1166_;
  assign new_n1168_ = new_n658_ & ~new_n1167_;
  assign new_n1169_ = ~new_n1161_ & ~new_n1168_;
  assign new_n1170_ = ~new_n1160_ & new_n1169_;
  assign new_n1171_ = ~\in2[116]  & \in3[116] ;
  assign new_n1172_ = ~new_n647_ & ~new_n1171_;
  assign new_n1173_ = new_n646_ & new_n1172_;
  assign new_n1174_ = ~new_n1170_ & new_n1173_;
  assign new_n1175_ = ~new_n654_ & ~new_n1174_;
  assign new_n1176_ = ~new_n652_ & new_n1175_;
  assign new_n1177_ = ~new_n643_ & new_n1176_;
  assign new_n1178_ = ~\in2[123]  & \in3[123] ;
  assign new_n1179_ = ~\in2[122]  & \in3[122] ;
  assign new_n1180_ = ~new_n1178_ & ~new_n1179_;
  assign new_n1181_ = ~\in2[121]  & \in3[121] ;
  assign new_n1182_ = ~\in2[120]  & \in3[120] ;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_ = new_n1180_ & new_n1183_;
  assign new_n1185_ = ~new_n1177_ & new_n1184_;
  assign new_n1186_ = \in2[123]  & ~\in3[123] ;
  assign new_n1187_ = \in2[120]  & ~\in3[120] ;
  assign new_n1188_ = ~new_n1181_ & new_n1187_;
  assign new_n1189_ = \in2[121]  & ~\in3[121] ;
  assign new_n1190_ = ~new_n1188_ & ~new_n1189_;
  assign new_n1191_ = \in2[122]  & ~\in3[122] ;
  assign new_n1192_ = new_n1190_ & ~new_n1191_;
  assign new_n1193_ = new_n1180_ & ~new_n1192_;
  assign new_n1194_ = ~new_n1186_ & ~new_n1193_;
  assign new_n1195_ = ~new_n1185_ & new_n1194_;
  assign new_n1196_ = ~\in2[124]  & \in3[124] ;
  assign new_n1197_ = \in2[127]  & ~\in3[127] ;
  assign new_n1198_ = ~\in2[126]  & \in3[126] ;
  assign new_n1199_ = ~\in2[125]  & \in3[125] ;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = ~new_n1197_ & new_n1200_;
  assign new_n1202_ = ~new_n1196_ & new_n1201_;
  assign new_n1203_ = ~new_n1195_ & new_n1202_;
  assign new_n1204_ = \in2[124]  & ~\in3[124] ;
  assign new_n1205_ = \in2[125]  & ~\in3[125] ;
  assign new_n1206_ = ~new_n1204_ & ~new_n1205_;
  assign new_n1207_ = new_n1200_ & ~new_n1206_;
  assign new_n1208_ = \in2[126]  & ~\in3[126] ;
  assign new_n1209_ = ~new_n1207_ & ~new_n1208_;
  assign new_n1210_ = ~new_n1197_ & ~new_n1209_;
  assign new_n1211_ = ~new_n1203_ & ~new_n1210_;
  assign new_n1212_ = ~\in3[127]  & new_n1211_;
  assign new_n1213_ = \in2[127]  & ~new_n1212_;
  assign new_n1214_ = \in0[119]  & ~\in1[119] ;
  assign new_n1215_ = ~\in0[119]  & \in1[119] ;
  assign new_n1216_ = ~\in0[118]  & \in1[118] ;
  assign new_n1217_ = ~new_n1215_ & ~new_n1216_;
  assign new_n1218_ = ~\in0[117]  & \in1[117] ;
  assign new_n1219_ = \in0[116]  & ~\in1[116] ;
  assign new_n1220_ = ~new_n1218_ & new_n1219_;
  assign new_n1221_ = \in0[117]  & ~\in1[117] ;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = new_n1217_ & ~new_n1222_;
  assign new_n1224_ = ~\in1[118]  & ~new_n1215_;
  assign new_n1225_ = \in0[118]  & new_n1224_;
  assign new_n1226_ = ~\in0[112]  & \in1[112] ;
  assign new_n1227_ = ~\in0[115]  & \in1[115] ;
  assign new_n1228_ = ~\in0[114]  & \in1[114] ;
  assign new_n1229_ = ~new_n1227_ & ~new_n1228_;
  assign new_n1230_ = ~\in0[113]  & \in1[113] ;
  assign new_n1231_ = \in0[111]  & ~\in1[111] ;
  assign new_n1232_ = ~\in0[111]  & \in1[111] ;
  assign new_n1233_ = ~\in0[110]  & \in1[110] ;
  assign new_n1234_ = ~new_n1232_ & ~new_n1233_;
  assign new_n1235_ = ~\in0[109]  & \in1[109] ;
  assign new_n1236_ = \in0[108]  & ~\in1[108] ;
  assign new_n1237_ = ~new_n1235_ & new_n1236_;
  assign new_n1238_ = \in0[109]  & ~\in1[109] ;
  assign new_n1239_ = ~new_n1237_ & ~new_n1238_;
  assign new_n1240_ = new_n1234_ & ~new_n1239_;
  assign new_n1241_ = ~\in1[110]  & ~new_n1232_;
  assign new_n1242_ = \in0[110]  & new_n1241_;
  assign new_n1243_ = \in0[103]  & ~\in1[103] ;
  assign new_n1244_ = ~\in0[103]  & \in1[103] ;
  assign new_n1245_ = ~\in0[102]  & \in1[102] ;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = ~\in0[101]  & \in1[101] ;
  assign new_n1248_ = \in0[100]  & ~\in1[100] ;
  assign new_n1249_ = ~new_n1247_ & new_n1248_;
  assign new_n1250_ = \in0[101]  & ~\in1[101] ;
  assign new_n1251_ = ~new_n1249_ & ~new_n1250_;
  assign new_n1252_ = new_n1246_ & ~new_n1251_;
  assign new_n1253_ = ~\in1[102]  & ~new_n1244_;
  assign new_n1254_ = \in0[102]  & new_n1253_;
  assign new_n1255_ = ~\in0[96]  & \in1[96] ;
  assign new_n1256_ = ~\in0[99]  & \in1[99] ;
  assign new_n1257_ = ~\in0[98]  & \in1[98] ;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = ~\in0[97]  & \in1[97] ;
  assign new_n1260_ = \in0[95]  & ~\in1[95] ;
  assign new_n1261_ = ~\in0[95]  & \in1[95] ;
  assign new_n1262_ = ~\in0[94]  & \in1[94] ;
  assign new_n1263_ = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = ~\in0[93]  & \in1[93] ;
  assign new_n1265_ = \in0[92]  & ~\in1[92] ;
  assign new_n1266_ = ~new_n1264_ & new_n1265_;
  assign new_n1267_ = \in0[93]  & ~\in1[93] ;
  assign new_n1268_ = ~new_n1266_ & ~new_n1267_;
  assign new_n1269_ = new_n1263_ & ~new_n1268_;
  assign new_n1270_ = ~\in1[94]  & ~new_n1261_;
  assign new_n1271_ = \in0[94]  & new_n1270_;
  assign new_n1272_ = \in0[87]  & ~\in1[87] ;
  assign new_n1273_ = ~\in0[87]  & \in1[87] ;
  assign new_n1274_ = ~\in0[86]  & \in1[86] ;
  assign new_n1275_ = ~new_n1273_ & ~new_n1274_;
  assign new_n1276_ = ~\in0[85]  & \in1[85] ;
  assign new_n1277_ = \in0[84]  & ~\in1[84] ;
  assign new_n1278_ = ~new_n1276_ & new_n1277_;
  assign new_n1279_ = \in0[85]  & ~\in1[85] ;
  assign new_n1280_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = new_n1275_ & ~new_n1280_;
  assign new_n1282_ = ~\in1[86]  & ~new_n1273_;
  assign new_n1283_ = \in0[86]  & new_n1282_;
  assign new_n1284_ = ~\in0[80]  & \in1[80] ;
  assign new_n1285_ = ~\in0[83]  & \in1[83] ;
  assign new_n1286_ = ~\in0[82]  & \in1[82] ;
  assign new_n1287_ = ~new_n1285_ & ~new_n1286_;
  assign new_n1288_ = ~\in0[81]  & \in1[81] ;
  assign new_n1289_ = \in0[79]  & ~\in1[79] ;
  assign new_n1290_ = ~\in0[79]  & \in1[79] ;
  assign new_n1291_ = ~\in0[78]  & \in1[78] ;
  assign new_n1292_ = ~new_n1290_ & ~new_n1291_;
  assign new_n1293_ = ~\in0[77]  & \in1[77] ;
  assign new_n1294_ = \in0[76]  & ~\in1[76] ;
  assign new_n1295_ = ~new_n1293_ & new_n1294_;
  assign new_n1296_ = \in0[77]  & ~\in1[77] ;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = new_n1292_ & ~new_n1297_;
  assign new_n1299_ = ~\in1[78]  & ~new_n1290_;
  assign new_n1300_ = \in0[78]  & new_n1299_;
  assign new_n1301_ = \in0[71]  & ~\in1[71] ;
  assign new_n1302_ = ~\in0[71]  & \in1[71] ;
  assign new_n1303_ = ~\in0[70]  & \in1[70] ;
  assign new_n1304_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = ~\in0[69]  & \in1[69] ;
  assign new_n1306_ = \in0[68]  & ~\in1[68] ;
  assign new_n1307_ = ~new_n1305_ & new_n1306_;
  assign new_n1308_ = \in0[69]  & ~\in1[69] ;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_ = new_n1304_ & ~new_n1309_;
  assign new_n1311_ = ~\in1[70]  & ~new_n1302_;
  assign new_n1312_ = \in0[70]  & new_n1311_;
  assign new_n1313_ = ~\in0[67]  & \in1[67] ;
  assign new_n1314_ = ~\in0[66]  & \in1[66] ;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1316_ = ~\in0[65]  & \in1[65] ;
  assign new_n1317_ = \in0[63]  & ~\in1[63] ;
  assign new_n1318_ = ~\in0[63]  & \in1[63] ;
  assign new_n1319_ = ~\in0[62]  & \in1[62] ;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = ~\in0[60]  & \in1[60] ;
  assign new_n1322_ = ~\in0[61]  & \in1[61] ;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign new_n1324_ = new_n1320_ & new_n1323_;
  assign new_n1325_ = \in0[59]  & ~\in1[59] ;
  assign new_n1326_ = ~\in0[59]  & \in1[59] ;
  assign new_n1327_ = ~\in0[58]  & \in1[58] ;
  assign new_n1328_ = ~new_n1326_ & ~new_n1327_;
  assign new_n1329_ = ~\in0[57]  & \in1[57] ;
  assign new_n1330_ = \in0[56]  & ~\in1[56] ;
  assign new_n1331_ = ~new_n1329_ & new_n1330_;
  assign new_n1332_ = \in0[57]  & ~\in1[57] ;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = \in0[58]  & ~\in1[58] ;
  assign new_n1335_ = new_n1333_ & ~new_n1334_;
  assign new_n1336_ = new_n1328_ & ~new_n1335_;
  assign new_n1337_ = ~new_n1325_ & ~new_n1336_;
  assign new_n1338_ = new_n1324_ & ~new_n1337_;
  assign new_n1339_ = \in0[60]  & ~\in1[60] ;
  assign new_n1340_ = ~new_n1322_ & new_n1339_;
  assign new_n1341_ = \in0[61]  & ~\in1[61] ;
  assign new_n1342_ = ~new_n1340_ & ~new_n1341_;
  assign new_n1343_ = new_n1320_ & ~new_n1342_;
  assign new_n1344_ = ~\in1[62]  & ~new_n1318_;
  assign new_n1345_ = \in0[62]  & new_n1344_;
  assign new_n1346_ = \in0[47]  & ~\in1[47] ;
  assign new_n1347_ = ~\in0[47]  & \in1[47] ;
  assign new_n1348_ = ~\in0[46]  & \in1[46] ;
  assign new_n1349_ = ~new_n1347_ & ~new_n1348_;
  assign new_n1350_ = ~\in0[44]  & \in1[44] ;
  assign new_n1351_ = ~\in0[45]  & \in1[45] ;
  assign new_n1352_ = ~new_n1350_ & ~new_n1351_;
  assign new_n1353_ = new_n1349_ & new_n1352_;
  assign new_n1354_ = \in0[43]  & ~\in1[43] ;
  assign new_n1355_ = ~\in0[43]  & \in1[43] ;
  assign new_n1356_ = ~\in0[42]  & \in1[42] ;
  assign new_n1357_ = ~new_n1355_ & ~new_n1356_;
  assign new_n1358_ = ~\in0[41]  & \in1[41] ;
  assign new_n1359_ = \in0[40]  & ~\in1[40] ;
  assign new_n1360_ = ~new_n1358_ & new_n1359_;
  assign new_n1361_ = \in0[41]  & ~\in1[41] ;
  assign new_n1362_ = ~new_n1360_ & ~new_n1361_;
  assign new_n1363_ = \in0[42]  & ~\in1[42] ;
  assign new_n1364_ = new_n1362_ & ~new_n1363_;
  assign new_n1365_ = new_n1357_ & ~new_n1364_;
  assign new_n1366_ = ~new_n1354_ & ~new_n1365_;
  assign new_n1367_ = new_n1353_ & ~new_n1366_;
  assign new_n1368_ = \in0[44]  & ~\in1[44] ;
  assign new_n1369_ = ~new_n1351_ & new_n1368_;
  assign new_n1370_ = \in0[45]  & ~\in1[45] ;
  assign new_n1371_ = ~new_n1369_ & ~new_n1370_;
  assign new_n1372_ = new_n1349_ & ~new_n1371_;
  assign new_n1373_ = ~\in1[46]  & ~new_n1347_;
  assign new_n1374_ = \in0[46]  & new_n1373_;
  assign new_n1375_ = ~\in0[32]  & \in1[32] ;
  assign new_n1376_ = ~\in0[31]  & \in1[31] ;
  assign new_n1377_ = ~\in0[30]  & \in1[30] ;
  assign new_n1378_ = ~\in0[29]  & \in1[29] ;
  assign new_n1379_ = ~\in0[28]  & \in1[28] ;
  assign new_n1380_ = ~\in0[27]  & \in1[27] ;
  assign new_n1381_ = ~\in0[26]  & \in1[26] ;
  assign new_n1382_ = ~\in0[23]  & \in1[23] ;
  assign new_n1383_ = ~\in0[22]  & \in1[22] ;
  assign new_n1384_ = ~\in0[21]  & \in1[21] ;
  assign new_n1385_ = ~\in0[20]  & \in1[20] ;
  assign new_n1386_ = ~\in0[19]  & \in1[19] ;
  assign new_n1387_ = ~\in0[18]  & \in1[18] ;
  assign new_n1388_ = ~\in0[15]  & \in1[15] ;
  assign new_n1389_ = ~\in0[14]  & \in1[14] ;
  assign new_n1390_ = ~\in0[13]  & \in1[13] ;
  assign new_n1391_ = ~\in0[12]  & \in1[12] ;
  assign new_n1392_ = ~\in0[11]  & \in1[11] ;
  assign new_n1393_ = ~\in0[10]  & \in1[10] ;
  assign new_n1394_ = ~\in0[7]  & \in1[7] ;
  assign new_n1395_ = ~\in0[6]  & \in1[6] ;
  assign new_n1396_ = ~\in0[3]  & \in1[3] ;
  assign new_n1397_ = \in0[0]  & ~\in1[0] ;
  assign new_n1398_ = \in0[1]  & ~\in1[1] ;
  assign new_n1399_ = ~new_n1397_ & ~new_n1398_;
  assign new_n1400_ = ~\in0[2]  & \in1[2] ;
  assign new_n1401_ = ~\in0[1]  & \in1[1] ;
  assign new_n1402_ = ~new_n1400_ & ~new_n1401_;
  assign new_n1403_ = ~new_n1399_ & new_n1402_;
  assign new_n1404_ = \in0[2]  & ~\in1[2] ;
  assign new_n1405_ = ~new_n1403_ & ~new_n1404_;
  assign new_n1406_ = ~new_n1396_ & ~new_n1405_;
  assign new_n1407_ = \in0[3]  & ~\in1[3] ;
  assign new_n1408_ = ~new_n1406_ & ~new_n1407_;
  assign new_n1409_ = ~\in0[4]  & new_n1408_;
  assign new_n1410_ = ~\in1[4]  & ~new_n1409_;
  assign new_n1411_ = \in0[4]  & ~new_n1408_;
  assign new_n1412_ = ~new_n1410_ & ~new_n1411_;
  assign new_n1413_ = ~\in0[5]  & new_n1412_;
  assign new_n1414_ = ~\in1[5]  & ~new_n1413_;
  assign new_n1415_ = \in0[5]  & ~new_n1412_;
  assign new_n1416_ = ~new_n1414_ & ~new_n1415_;
  assign new_n1417_ = ~new_n1395_ & ~new_n1416_;
  assign new_n1418_ = \in0[6]  & ~\in1[6] ;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_ = ~new_n1394_ & ~new_n1419_;
  assign new_n1421_ = \in0[7]  & ~\in1[7] ;
  assign new_n1422_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = ~\in0[8]  & new_n1422_;
  assign new_n1424_ = ~\in1[8]  & ~new_n1423_;
  assign new_n1425_ = \in0[8]  & ~new_n1422_;
  assign new_n1426_ = ~new_n1424_ & ~new_n1425_;
  assign new_n1427_ = ~\in0[9]  & new_n1426_;
  assign new_n1428_ = ~\in1[9]  & ~new_n1427_;
  assign new_n1429_ = \in0[9]  & ~new_n1426_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n1393_ & ~new_n1430_;
  assign new_n1432_ = \in0[10]  & ~\in1[10] ;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = ~new_n1392_ & ~new_n1433_;
  assign new_n1435_ = \in0[11]  & ~\in1[11] ;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = ~new_n1391_ & ~new_n1436_;
  assign new_n1438_ = \in0[12]  & ~\in1[12] ;
  assign new_n1439_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1440_ = ~new_n1390_ & ~new_n1439_;
  assign new_n1441_ = \in0[13]  & ~\in1[13] ;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1443_ = ~new_n1389_ & ~new_n1442_;
  assign new_n1444_ = \in0[14]  & ~\in1[14] ;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = ~new_n1388_ & ~new_n1445_;
  assign new_n1447_ = \in0[15]  & ~\in1[15] ;
  assign new_n1448_ = ~new_n1446_ & ~new_n1447_;
  assign new_n1449_ = ~\in0[16]  & new_n1448_;
  assign new_n1450_ = ~\in1[16]  & ~new_n1449_;
  assign new_n1451_ = \in0[16]  & ~new_n1448_;
  assign new_n1452_ = ~new_n1450_ & ~new_n1451_;
  assign new_n1453_ = ~\in0[17]  & new_n1452_;
  assign new_n1454_ = ~\in1[17]  & ~new_n1453_;
  assign new_n1455_ = \in0[17]  & ~new_n1452_;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1457_ = ~new_n1387_ & ~new_n1456_;
  assign new_n1458_ = \in0[18]  & ~\in1[18] ;
  assign new_n1459_ = ~new_n1457_ & ~new_n1458_;
  assign new_n1460_ = ~new_n1386_ & ~new_n1459_;
  assign new_n1461_ = \in0[19]  & ~\in1[19] ;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = ~new_n1385_ & ~new_n1462_;
  assign new_n1464_ = \in0[20]  & ~\in1[20] ;
  assign new_n1465_ = ~new_n1463_ & ~new_n1464_;
  assign new_n1466_ = ~new_n1384_ & ~new_n1465_;
  assign new_n1467_ = \in0[21]  & ~\in1[21] ;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = ~new_n1383_ & ~new_n1468_;
  assign new_n1470_ = \in0[22]  & ~\in1[22] ;
  assign new_n1471_ = ~new_n1469_ & ~new_n1470_;
  assign new_n1472_ = ~new_n1382_ & ~new_n1471_;
  assign new_n1473_ = \in0[23]  & ~\in1[23] ;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = ~\in0[24]  & new_n1474_;
  assign new_n1476_ = ~\in1[24]  & ~new_n1475_;
  assign new_n1477_ = \in0[24]  & ~new_n1474_;
  assign new_n1478_ = ~new_n1476_ & ~new_n1477_;
  assign new_n1479_ = ~\in0[25]  & new_n1478_;
  assign new_n1480_ = ~\in1[25]  & ~new_n1479_;
  assign new_n1481_ = \in0[25]  & ~new_n1478_;
  assign new_n1482_ = ~new_n1480_ & ~new_n1481_;
  assign new_n1483_ = ~new_n1381_ & ~new_n1482_;
  assign new_n1484_ = \in0[26]  & ~\in1[26] ;
  assign new_n1485_ = ~new_n1483_ & ~new_n1484_;
  assign new_n1486_ = ~new_n1380_ & ~new_n1485_;
  assign new_n1487_ = \in0[27]  & ~\in1[27] ;
  assign new_n1488_ = ~new_n1486_ & ~new_n1487_;
  assign new_n1489_ = ~new_n1379_ & ~new_n1488_;
  assign new_n1490_ = \in0[28]  & ~\in1[28] ;
  assign new_n1491_ = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = ~new_n1378_ & ~new_n1491_;
  assign new_n1493_ = \in0[29]  & ~\in1[29] ;
  assign new_n1494_ = ~new_n1492_ & ~new_n1493_;
  assign new_n1495_ = ~new_n1377_ & ~new_n1494_;
  assign new_n1496_ = \in0[30]  & ~\in1[30] ;
  assign new_n1497_ = ~new_n1495_ & ~new_n1496_;
  assign new_n1498_ = ~new_n1376_ & ~new_n1497_;
  assign new_n1499_ = \in0[31]  & ~\in1[31] ;
  assign new_n1500_ = ~new_n1498_ & ~new_n1499_;
  assign new_n1501_ = ~\in0[39]  & \in1[39] ;
  assign new_n1502_ = ~\in0[38]  & \in1[38] ;
  assign new_n1503_ = ~new_n1501_ & ~new_n1502_;
  assign new_n1504_ = ~\in0[36]  & \in1[36] ;
  assign new_n1505_ = ~\in0[37]  & \in1[37] ;
  assign new_n1506_ = ~new_n1504_ & ~new_n1505_;
  assign new_n1507_ = new_n1503_ & new_n1506_;
  assign new_n1508_ = ~\in0[33]  & \in1[33] ;
  assign new_n1509_ = ~\in0[35]  & \in1[35] ;
  assign new_n1510_ = ~\in0[34]  & \in1[34] ;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = ~new_n1508_ & new_n1511_;
  assign new_n1513_ = new_n1507_ & new_n1512_;
  assign new_n1514_ = ~new_n1500_ & new_n1513_;
  assign new_n1515_ = ~new_n1375_ & new_n1514_;
  assign new_n1516_ = \in0[39]  & ~\in1[39] ;
  assign new_n1517_ = \in0[36]  & ~\in1[36] ;
  assign new_n1518_ = ~new_n1505_ & new_n1517_;
  assign new_n1519_ = \in0[37]  & ~\in1[37] ;
  assign new_n1520_ = ~new_n1518_ & ~new_n1519_;
  assign new_n1521_ = new_n1503_ & ~new_n1520_;
  assign new_n1522_ = ~\in1[38]  & ~new_n1501_;
  assign new_n1523_ = \in0[38]  & new_n1522_;
  assign new_n1524_ = \in0[35]  & ~\in1[35] ;
  assign new_n1525_ = ~\in1[32]  & ~new_n1508_;
  assign new_n1526_ = \in0[32]  & new_n1525_;
  assign new_n1527_ = \in0[33]  & ~\in1[33] ;
  assign new_n1528_ = ~new_n1526_ & ~new_n1527_;
  assign new_n1529_ = \in0[34]  & ~\in1[34] ;
  assign new_n1530_ = new_n1528_ & ~new_n1529_;
  assign new_n1531_ = new_n1511_ & ~new_n1530_;
  assign new_n1532_ = ~new_n1524_ & ~new_n1531_;
  assign new_n1533_ = new_n1507_ & ~new_n1532_;
  assign new_n1534_ = ~new_n1523_ & ~new_n1533_;
  assign new_n1535_ = ~new_n1521_ & new_n1534_;
  assign new_n1536_ = ~new_n1516_ & new_n1535_;
  assign new_n1537_ = ~new_n1515_ & new_n1536_;
  assign new_n1538_ = ~\in0[40]  & \in1[40] ;
  assign new_n1539_ = ~new_n1358_ & ~new_n1538_;
  assign new_n1540_ = new_n1357_ & new_n1539_;
  assign new_n1541_ = new_n1353_ & new_n1540_;
  assign new_n1542_ = ~new_n1537_ & new_n1541_;
  assign new_n1543_ = ~new_n1374_ & ~new_n1542_;
  assign new_n1544_ = ~new_n1372_ & new_n1543_;
  assign new_n1545_ = ~new_n1367_ & new_n1544_;
  assign new_n1546_ = ~new_n1346_ & new_n1545_;
  assign new_n1547_ = ~\in0[48]  & \in1[48] ;
  assign new_n1548_ = ~\in0[55]  & \in1[55] ;
  assign new_n1549_ = ~\in0[54]  & \in1[54] ;
  assign new_n1550_ = ~new_n1548_ & ~new_n1549_;
  assign new_n1551_ = ~\in0[53]  & \in1[53] ;
  assign new_n1552_ = ~\in0[52]  & \in1[52] ;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_ = new_n1550_ & new_n1553_;
  assign new_n1555_ = ~\in0[49]  & \in1[49] ;
  assign new_n1556_ = ~\in0[51]  & \in1[51] ;
  assign new_n1557_ = ~\in0[50]  & \in1[50] ;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = ~new_n1555_ & new_n1558_;
  assign new_n1560_ = new_n1554_ & new_n1559_;
  assign new_n1561_ = ~new_n1547_ & new_n1560_;
  assign new_n1562_ = ~new_n1546_ & new_n1561_;
  assign new_n1563_ = \in0[55]  & ~\in1[55] ;
  assign new_n1564_ = \in0[51]  & ~\in1[51] ;
  assign new_n1565_ = ~\in1[48]  & ~new_n1555_;
  assign new_n1566_ = \in0[48]  & new_n1565_;
  assign new_n1567_ = \in0[49]  & ~\in1[49] ;
  assign new_n1568_ = ~new_n1566_ & ~new_n1567_;
  assign new_n1569_ = \in0[50]  & ~\in1[50] ;
  assign new_n1570_ = new_n1568_ & ~new_n1569_;
  assign new_n1571_ = new_n1558_ & ~new_n1570_;
  assign new_n1572_ = ~new_n1564_ & ~new_n1571_;
  assign new_n1573_ = new_n1554_ & ~new_n1572_;
  assign new_n1574_ = \in0[52]  & ~\in1[52] ;
  assign new_n1575_ = ~new_n1551_ & new_n1574_;
  assign new_n1576_ = \in0[53]  & ~\in1[53] ;
  assign new_n1577_ = ~new_n1575_ & ~new_n1576_;
  assign new_n1578_ = \in0[54]  & ~\in1[54] ;
  assign new_n1579_ = new_n1577_ & ~new_n1578_;
  assign new_n1580_ = new_n1550_ & ~new_n1579_;
  assign new_n1581_ = ~new_n1573_ & ~new_n1580_;
  assign new_n1582_ = ~new_n1563_ & new_n1581_;
  assign new_n1583_ = ~new_n1562_ & new_n1582_;
  assign new_n1584_ = ~\in0[56]  & \in1[56] ;
  assign new_n1585_ = ~new_n1329_ & ~new_n1584_;
  assign new_n1586_ = new_n1324_ & new_n1585_;
  assign new_n1587_ = new_n1328_ & new_n1586_;
  assign new_n1588_ = ~new_n1583_ & new_n1587_;
  assign new_n1589_ = ~new_n1345_ & ~new_n1588_;
  assign new_n1590_ = ~new_n1343_ & new_n1589_;
  assign new_n1591_ = ~new_n1338_ & new_n1590_;
  assign new_n1592_ = ~new_n1317_ & new_n1591_;
  assign new_n1593_ = ~\in0[64]  & \in1[64] ;
  assign new_n1594_ = ~new_n1592_ & ~new_n1593_;
  assign new_n1595_ = ~new_n1316_ & new_n1594_;
  assign new_n1596_ = new_n1315_ & new_n1595_;
  assign new_n1597_ = \in0[67]  & ~\in1[67] ;
  assign new_n1598_ = \in0[64]  & ~\in1[64] ;
  assign new_n1599_ = ~new_n1316_ & new_n1598_;
  assign new_n1600_ = \in0[65]  & ~\in1[65] ;
  assign new_n1601_ = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = \in0[66]  & ~\in1[66] ;
  assign new_n1603_ = new_n1601_ & ~new_n1602_;
  assign new_n1604_ = new_n1315_ & ~new_n1603_;
  assign new_n1605_ = ~new_n1597_ & ~new_n1604_;
  assign new_n1606_ = ~new_n1596_ & new_n1605_;
  assign new_n1607_ = ~\in0[68]  & \in1[68] ;
  assign new_n1608_ = ~new_n1305_ & ~new_n1607_;
  assign new_n1609_ = new_n1304_ & new_n1608_;
  assign new_n1610_ = ~new_n1606_ & new_n1609_;
  assign new_n1611_ = ~new_n1312_ & ~new_n1610_;
  assign new_n1612_ = ~new_n1310_ & new_n1611_;
  assign new_n1613_ = ~new_n1301_ & new_n1612_;
  assign new_n1614_ = ~\in0[75]  & \in1[75] ;
  assign new_n1615_ = ~\in0[74]  & \in1[74] ;
  assign new_n1616_ = ~new_n1614_ & ~new_n1615_;
  assign new_n1617_ = ~\in0[73]  & \in1[73] ;
  assign new_n1618_ = ~\in0[72]  & \in1[72] ;
  assign new_n1619_ = ~new_n1617_ & ~new_n1618_;
  assign new_n1620_ = new_n1616_ & new_n1619_;
  assign new_n1621_ = ~new_n1613_ & new_n1620_;
  assign new_n1622_ = \in0[75]  & ~\in1[75] ;
  assign new_n1623_ = \in0[72]  & ~\in1[72] ;
  assign new_n1624_ = ~new_n1617_ & new_n1623_;
  assign new_n1625_ = \in0[73]  & ~\in1[73] ;
  assign new_n1626_ = ~new_n1624_ & ~new_n1625_;
  assign new_n1627_ = \in0[74]  & ~\in1[74] ;
  assign new_n1628_ = new_n1626_ & ~new_n1627_;
  assign new_n1629_ = new_n1616_ & ~new_n1628_;
  assign new_n1630_ = ~new_n1622_ & ~new_n1629_;
  assign new_n1631_ = ~new_n1621_ & new_n1630_;
  assign new_n1632_ = ~\in0[76]  & \in1[76] ;
  assign new_n1633_ = ~new_n1293_ & ~new_n1632_;
  assign new_n1634_ = new_n1292_ & new_n1633_;
  assign new_n1635_ = ~new_n1631_ & new_n1634_;
  assign new_n1636_ = ~new_n1300_ & ~new_n1635_;
  assign new_n1637_ = ~new_n1298_ & new_n1636_;
  assign new_n1638_ = ~new_n1289_ & new_n1637_;
  assign new_n1639_ = ~new_n1288_ & ~new_n1638_;
  assign new_n1640_ = new_n1287_ & new_n1639_;
  assign new_n1641_ = ~new_n1284_ & new_n1640_;
  assign new_n1642_ = \in0[83]  & ~\in1[83] ;
  assign new_n1643_ = ~\in1[80]  & ~new_n1288_;
  assign new_n1644_ = \in0[80]  & new_n1643_;
  assign new_n1645_ = \in0[81]  & ~\in1[81] ;
  assign new_n1646_ = ~new_n1644_ & ~new_n1645_;
  assign new_n1647_ = \in0[82]  & ~\in1[82] ;
  assign new_n1648_ = new_n1646_ & ~new_n1647_;
  assign new_n1649_ = new_n1287_ & ~new_n1648_;
  assign new_n1650_ = ~new_n1642_ & ~new_n1649_;
  assign new_n1651_ = ~new_n1641_ & new_n1650_;
  assign new_n1652_ = ~\in0[84]  & \in1[84] ;
  assign new_n1653_ = ~new_n1276_ & ~new_n1652_;
  assign new_n1654_ = new_n1275_ & new_n1653_;
  assign new_n1655_ = ~new_n1651_ & new_n1654_;
  assign new_n1656_ = ~new_n1283_ & ~new_n1655_;
  assign new_n1657_ = ~new_n1281_ & new_n1656_;
  assign new_n1658_ = ~new_n1272_ & new_n1657_;
  assign new_n1659_ = ~\in0[91]  & \in1[91] ;
  assign new_n1660_ = ~\in0[90]  & \in1[90] ;
  assign new_n1661_ = ~new_n1659_ & ~new_n1660_;
  assign new_n1662_ = ~\in0[89]  & \in1[89] ;
  assign new_n1663_ = ~\in0[88]  & \in1[88] ;
  assign new_n1664_ = ~new_n1662_ & ~new_n1663_;
  assign new_n1665_ = new_n1661_ & new_n1664_;
  assign new_n1666_ = ~new_n1658_ & new_n1665_;
  assign new_n1667_ = \in0[91]  & ~\in1[91] ;
  assign new_n1668_ = \in0[88]  & ~\in1[88] ;
  assign new_n1669_ = ~new_n1662_ & new_n1668_;
  assign new_n1670_ = \in0[89]  & ~\in1[89] ;
  assign new_n1671_ = ~new_n1669_ & ~new_n1670_;
  assign new_n1672_ = \in0[90]  & ~\in1[90] ;
  assign new_n1673_ = new_n1671_ & ~new_n1672_;
  assign new_n1674_ = new_n1661_ & ~new_n1673_;
  assign new_n1675_ = ~new_n1667_ & ~new_n1674_;
  assign new_n1676_ = ~new_n1666_ & new_n1675_;
  assign new_n1677_ = ~\in0[92]  & \in1[92] ;
  assign new_n1678_ = ~new_n1264_ & ~new_n1677_;
  assign new_n1679_ = new_n1263_ & new_n1678_;
  assign new_n1680_ = ~new_n1676_ & new_n1679_;
  assign new_n1681_ = ~new_n1271_ & ~new_n1680_;
  assign new_n1682_ = ~new_n1269_ & new_n1681_;
  assign new_n1683_ = ~new_n1260_ & new_n1682_;
  assign new_n1684_ = ~new_n1259_ & ~new_n1683_;
  assign new_n1685_ = new_n1258_ & new_n1684_;
  assign new_n1686_ = ~new_n1255_ & new_n1685_;
  assign new_n1687_ = \in0[99]  & ~\in1[99] ;
  assign new_n1688_ = ~\in1[96]  & ~new_n1259_;
  assign new_n1689_ = \in0[96]  & new_n1688_;
  assign new_n1690_ = \in0[97]  & ~\in1[97] ;
  assign new_n1691_ = ~new_n1689_ & ~new_n1690_;
  assign new_n1692_ = \in0[98]  & ~\in1[98] ;
  assign new_n1693_ = new_n1691_ & ~new_n1692_;
  assign new_n1694_ = new_n1258_ & ~new_n1693_;
  assign new_n1695_ = ~new_n1687_ & ~new_n1694_;
  assign new_n1696_ = ~new_n1686_ & new_n1695_;
  assign new_n1697_ = ~\in0[100]  & \in1[100] ;
  assign new_n1698_ = ~new_n1247_ & ~new_n1697_;
  assign new_n1699_ = new_n1246_ & new_n1698_;
  assign new_n1700_ = ~new_n1696_ & new_n1699_;
  assign new_n1701_ = ~new_n1254_ & ~new_n1700_;
  assign new_n1702_ = ~new_n1252_ & new_n1701_;
  assign new_n1703_ = ~new_n1243_ & new_n1702_;
  assign new_n1704_ = ~\in0[107]  & \in1[107] ;
  assign new_n1705_ = ~\in0[106]  & \in1[106] ;
  assign new_n1706_ = ~new_n1704_ & ~new_n1705_;
  assign new_n1707_ = ~\in0[105]  & \in1[105] ;
  assign new_n1708_ = ~\in0[104]  & \in1[104] ;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_ = new_n1706_ & new_n1709_;
  assign new_n1711_ = ~new_n1703_ & new_n1710_;
  assign new_n1712_ = \in0[107]  & ~\in1[107] ;
  assign new_n1713_ = \in0[104]  & ~\in1[104] ;
  assign new_n1714_ = ~new_n1707_ & new_n1713_;
  assign new_n1715_ = \in0[105]  & ~\in1[105] ;
  assign new_n1716_ = ~new_n1714_ & ~new_n1715_;
  assign new_n1717_ = \in0[106]  & ~\in1[106] ;
  assign new_n1718_ = new_n1716_ & ~new_n1717_;
  assign new_n1719_ = new_n1706_ & ~new_n1718_;
  assign new_n1720_ = ~new_n1712_ & ~new_n1719_;
  assign new_n1721_ = ~new_n1711_ & new_n1720_;
  assign new_n1722_ = ~\in0[108]  & \in1[108] ;
  assign new_n1723_ = ~new_n1235_ & ~new_n1722_;
  assign new_n1724_ = new_n1234_ & new_n1723_;
  assign new_n1725_ = ~new_n1721_ & new_n1724_;
  assign new_n1726_ = ~new_n1242_ & ~new_n1725_;
  assign new_n1727_ = ~new_n1240_ & new_n1726_;
  assign new_n1728_ = ~new_n1231_ & new_n1727_;
  assign new_n1729_ = ~new_n1230_ & ~new_n1728_;
  assign new_n1730_ = new_n1229_ & new_n1729_;
  assign new_n1731_ = ~new_n1226_ & new_n1730_;
  assign new_n1732_ = \in0[115]  & ~\in1[115] ;
  assign new_n1733_ = ~\in1[112]  & ~new_n1230_;
  assign new_n1734_ = \in0[112]  & new_n1733_;
  assign new_n1735_ = \in0[113]  & ~\in1[113] ;
  assign new_n1736_ = ~new_n1734_ & ~new_n1735_;
  assign new_n1737_ = \in0[114]  & ~\in1[114] ;
  assign new_n1738_ = new_n1736_ & ~new_n1737_;
  assign new_n1739_ = new_n1229_ & ~new_n1738_;
  assign new_n1740_ = ~new_n1732_ & ~new_n1739_;
  assign new_n1741_ = ~new_n1731_ & new_n1740_;
  assign new_n1742_ = ~\in0[116]  & \in1[116] ;
  assign new_n1743_ = ~new_n1218_ & ~new_n1742_;
  assign new_n1744_ = new_n1217_ & new_n1743_;
  assign new_n1745_ = ~new_n1741_ & new_n1744_;
  assign new_n1746_ = ~new_n1225_ & ~new_n1745_;
  assign new_n1747_ = ~new_n1223_ & new_n1746_;
  assign new_n1748_ = ~new_n1214_ & new_n1747_;
  assign new_n1749_ = ~\in0[123]  & \in1[123] ;
  assign new_n1750_ = ~\in0[122]  & \in1[122] ;
  assign new_n1751_ = ~new_n1749_ & ~new_n1750_;
  assign new_n1752_ = ~\in0[121]  & \in1[121] ;
  assign new_n1753_ = ~\in0[120]  & \in1[120] ;
  assign new_n1754_ = ~new_n1752_ & ~new_n1753_;
  assign new_n1755_ = new_n1751_ & new_n1754_;
  assign new_n1756_ = ~new_n1748_ & new_n1755_;
  assign new_n1757_ = \in0[123]  & ~\in1[123] ;
  assign new_n1758_ = \in0[120]  & ~\in1[120] ;
  assign new_n1759_ = ~new_n1752_ & new_n1758_;
  assign new_n1760_ = \in0[121]  & ~\in1[121] ;
  assign new_n1761_ = ~new_n1759_ & ~new_n1760_;
  assign new_n1762_ = \in0[122]  & ~\in1[122] ;
  assign new_n1763_ = new_n1761_ & ~new_n1762_;
  assign new_n1764_ = new_n1751_ & ~new_n1763_;
  assign new_n1765_ = ~new_n1757_ & ~new_n1764_;
  assign new_n1766_ = ~new_n1756_ & new_n1765_;
  assign new_n1767_ = ~\in0[124]  & \in1[124] ;
  assign new_n1768_ = \in0[127]  & ~\in1[127] ;
  assign new_n1769_ = ~\in0[126]  & \in1[126] ;
  assign new_n1770_ = ~\in0[125]  & \in1[125] ;
  assign new_n1771_ = ~new_n1769_ & ~new_n1770_;
  assign new_n1772_ = ~new_n1768_ & new_n1771_;
  assign new_n1773_ = ~new_n1767_ & new_n1772_;
  assign new_n1774_ = ~new_n1766_ & new_n1773_;
  assign new_n1775_ = \in0[124]  & ~\in1[124] ;
  assign new_n1776_ = \in0[125]  & ~\in1[125] ;
  assign new_n1777_ = ~new_n1775_ & ~new_n1776_;
  assign new_n1778_ = new_n1771_ & ~new_n1777_;
  assign new_n1779_ = \in0[126]  & ~\in1[126] ;
  assign new_n1780_ = ~new_n1778_ & ~new_n1779_;
  assign new_n1781_ = ~new_n1768_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1774_ & ~new_n1781_;
  assign new_n1783_ = ~\in1[127]  & new_n1782_;
  assign new_n1784_ = \in0[127]  & ~new_n1783_;
  assign new_n1785_ = new_n1213_ & ~new_n1784_;
  assign new_n1786_ = ~\in0[127]  & \in1[127] ;
  assign new_n1787_ = new_n1782_ & ~new_n1786_;
  assign new_n1788_ = \in1[119]  & new_n1787_;
  assign new_n1789_ = \in0[119]  & ~new_n1787_;
  assign new_n1790_ = ~new_n1788_ & ~new_n1789_;
  assign new_n1791_ = ~\in2[127]  & \in3[127] ;
  assign new_n1792_ = new_n1211_ & ~new_n1791_;
  assign new_n1793_ = \in3[119]  & new_n1792_;
  assign new_n1794_ = \in2[119]  & ~new_n1792_;
  assign new_n1795_ = ~new_n1793_ & ~new_n1794_;
  assign new_n1796_ = ~new_n1790_ & new_n1795_;
  assign new_n1797_ = new_n1790_ & ~new_n1795_;
  assign new_n1798_ = \in3[118]  & new_n1792_;
  assign new_n1799_ = \in2[118]  & ~new_n1792_;
  assign new_n1800_ = ~new_n1798_ & ~new_n1799_;
  assign new_n1801_ = \in1[118]  & new_n1787_;
  assign new_n1802_ = \in0[118]  & ~new_n1787_;
  assign new_n1803_ = ~new_n1801_ & ~new_n1802_;
  assign new_n1804_ = ~new_n1800_ & new_n1803_;
  assign new_n1805_ = ~new_n1797_ & ~new_n1804_;
  assign new_n1806_ = \in1[116]  & new_n1787_;
  assign new_n1807_ = \in0[116]  & ~new_n1787_;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_ = \in1[117]  & new_n1787_;
  assign new_n1810_ = \in0[117]  & ~new_n1787_;
  assign new_n1811_ = ~new_n1809_ & ~new_n1810_;
  assign new_n1812_ = \in3[117]  & new_n1792_;
  assign new_n1813_ = \in2[117]  & ~new_n1792_;
  assign new_n1814_ = ~new_n1812_ & ~new_n1813_;
  assign new_n1815_ = new_n1811_ & ~new_n1814_;
  assign new_n1816_ = \in3[116]  & new_n1792_;
  assign new_n1817_ = \in2[116]  & ~new_n1792_;
  assign new_n1818_ = ~new_n1816_ & ~new_n1817_;
  assign new_n1819_ = ~new_n1815_ & new_n1818_;
  assign new_n1820_ = ~new_n1808_ & new_n1819_;
  assign new_n1821_ = ~new_n1811_ & new_n1814_;
  assign new_n1822_ = ~new_n1820_ & ~new_n1821_;
  assign new_n1823_ = new_n1805_ & ~new_n1822_;
  assign new_n1824_ = new_n1800_ & ~new_n1803_;
  assign new_n1825_ = ~new_n1797_ & new_n1824_;
  assign new_n1826_ = \in3[112]  & new_n1792_;
  assign new_n1827_ = \in2[112]  & ~new_n1792_;
  assign new_n1828_ = ~new_n1826_ & ~new_n1827_;
  assign new_n1829_ = \in1[112]  & new_n1787_;
  assign new_n1830_ = \in0[112]  & ~new_n1787_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = ~new_n1828_ & new_n1831_;
  assign new_n1833_ = \in1[115]  & new_n1787_;
  assign new_n1834_ = \in0[115]  & ~new_n1787_;
  assign new_n1835_ = ~new_n1833_ & ~new_n1834_;
  assign new_n1836_ = \in3[115]  & new_n1792_;
  assign new_n1837_ = \in2[115]  & ~new_n1792_;
  assign new_n1838_ = ~new_n1836_ & ~new_n1837_;
  assign new_n1839_ = new_n1835_ & ~new_n1838_;
  assign new_n1840_ = \in3[114]  & new_n1792_;
  assign new_n1841_ = \in2[114]  & ~new_n1792_;
  assign new_n1842_ = ~new_n1840_ & ~new_n1841_;
  assign new_n1843_ = \in1[114]  & new_n1787_;
  assign new_n1844_ = \in0[114]  & ~new_n1787_;
  assign new_n1845_ = ~new_n1843_ & ~new_n1844_;
  assign new_n1846_ = ~new_n1842_ & new_n1845_;
  assign new_n1847_ = ~new_n1839_ & ~new_n1846_;
  assign new_n1848_ = \in1[113]  & new_n1787_;
  assign new_n1849_ = \in0[113]  & ~new_n1787_;
  assign new_n1850_ = ~new_n1848_ & ~new_n1849_;
  assign new_n1851_ = \in3[113]  & new_n1792_;
  assign new_n1852_ = \in2[113]  & ~new_n1792_;
  assign new_n1853_ = ~new_n1851_ & ~new_n1852_;
  assign new_n1854_ = new_n1850_ & ~new_n1853_;
  assign new_n1855_ = \in1[111]  & new_n1787_;
  assign new_n1856_ = \in0[111]  & ~new_n1787_;
  assign new_n1857_ = ~new_n1855_ & ~new_n1856_;
  assign new_n1858_ = \in3[111]  & new_n1792_;
  assign new_n1859_ = \in2[111]  & ~new_n1792_;
  assign new_n1860_ = ~new_n1858_ & ~new_n1859_;
  assign new_n1861_ = ~new_n1857_ & new_n1860_;
  assign new_n1862_ = new_n1857_ & ~new_n1860_;
  assign new_n1863_ = \in3[110]  & new_n1792_;
  assign new_n1864_ = \in2[110]  & ~new_n1792_;
  assign new_n1865_ = ~new_n1863_ & ~new_n1864_;
  assign new_n1866_ = \in1[110]  & new_n1787_;
  assign new_n1867_ = \in0[110]  & ~new_n1787_;
  assign new_n1868_ = ~new_n1866_ & ~new_n1867_;
  assign new_n1869_ = ~new_n1865_ & new_n1868_;
  assign new_n1870_ = ~new_n1862_ & ~new_n1869_;
  assign new_n1871_ = \in1[109]  & new_n1787_;
  assign new_n1872_ = \in0[109]  & ~new_n1787_;
  assign new_n1873_ = ~new_n1871_ & ~new_n1872_;
  assign new_n1874_ = \in3[109]  & new_n1792_;
  assign new_n1875_ = \in2[109]  & ~new_n1792_;
  assign new_n1876_ = ~new_n1874_ & ~new_n1875_;
  assign new_n1877_ = new_n1873_ & ~new_n1876_;
  assign new_n1878_ = \in1[108]  & new_n1787_;
  assign new_n1879_ = \in0[108]  & ~new_n1787_;
  assign new_n1880_ = ~new_n1878_ & ~new_n1879_;
  assign new_n1881_ = \in3[108]  & new_n1792_;
  assign new_n1882_ = \in2[108]  & ~new_n1792_;
  assign new_n1883_ = ~new_n1881_ & ~new_n1882_;
  assign new_n1884_ = ~new_n1880_ & new_n1883_;
  assign new_n1885_ = ~new_n1877_ & new_n1884_;
  assign new_n1886_ = ~new_n1873_ & new_n1876_;
  assign new_n1887_ = ~new_n1885_ & ~new_n1886_;
  assign new_n1888_ = new_n1870_ & ~new_n1887_;
  assign new_n1889_ = new_n1865_ & ~new_n1868_;
  assign new_n1890_ = ~new_n1862_ & new_n1889_;
  assign new_n1891_ = \in1[103]  & new_n1787_;
  assign new_n1892_ = \in0[103]  & ~new_n1787_;
  assign new_n1893_ = ~new_n1891_ & ~new_n1892_;
  assign new_n1894_ = \in3[103]  & new_n1792_;
  assign new_n1895_ = \in2[103]  & ~new_n1792_;
  assign new_n1896_ = ~new_n1894_ & ~new_n1895_;
  assign new_n1897_ = ~new_n1893_ & new_n1896_;
  assign new_n1898_ = new_n1893_ & ~new_n1896_;
  assign new_n1899_ = \in3[102]  & new_n1792_;
  assign new_n1900_ = \in2[102]  & ~new_n1792_;
  assign new_n1901_ = ~new_n1899_ & ~new_n1900_;
  assign new_n1902_ = \in1[102]  & new_n1787_;
  assign new_n1903_ = \in0[102]  & ~new_n1787_;
  assign new_n1904_ = ~new_n1902_ & ~new_n1903_;
  assign new_n1905_ = ~new_n1901_ & new_n1904_;
  assign new_n1906_ = ~new_n1898_ & ~new_n1905_;
  assign new_n1907_ = \in1[101]  & new_n1787_;
  assign new_n1908_ = \in0[101]  & ~new_n1787_;
  assign new_n1909_ = ~new_n1907_ & ~new_n1908_;
  assign new_n1910_ = \in3[101]  & new_n1792_;
  assign new_n1911_ = \in2[101]  & ~new_n1792_;
  assign new_n1912_ = ~new_n1910_ & ~new_n1911_;
  assign new_n1913_ = new_n1909_ & ~new_n1912_;
  assign new_n1914_ = \in1[100]  & new_n1787_;
  assign new_n1915_ = \in0[100]  & ~new_n1787_;
  assign new_n1916_ = ~new_n1914_ & ~new_n1915_;
  assign new_n1917_ = \in3[100]  & new_n1792_;
  assign new_n1918_ = \in2[100]  & ~new_n1792_;
  assign new_n1919_ = ~new_n1917_ & ~new_n1918_;
  assign new_n1920_ = ~new_n1916_ & new_n1919_;
  assign new_n1921_ = ~new_n1913_ & new_n1920_;
  assign new_n1922_ = ~new_n1909_ & new_n1912_;
  assign new_n1923_ = ~new_n1921_ & ~new_n1922_;
  assign new_n1924_ = new_n1906_ & ~new_n1923_;
  assign new_n1925_ = new_n1901_ & ~new_n1904_;
  assign new_n1926_ = ~new_n1898_ & new_n1925_;
  assign new_n1927_ = \in3[96]  & new_n1792_;
  assign new_n1928_ = \in2[96]  & ~new_n1792_;
  assign new_n1929_ = ~new_n1927_ & ~new_n1928_;
  assign new_n1930_ = \in1[96]  & new_n1787_;
  assign new_n1931_ = \in0[96]  & ~new_n1787_;
  assign new_n1932_ = ~new_n1930_ & ~new_n1931_;
  assign new_n1933_ = ~new_n1929_ & new_n1932_;
  assign new_n1934_ = \in1[99]  & new_n1787_;
  assign new_n1935_ = \in0[99]  & ~new_n1787_;
  assign new_n1936_ = ~new_n1934_ & ~new_n1935_;
  assign new_n1937_ = \in3[99]  & new_n1792_;
  assign new_n1938_ = \in2[99]  & ~new_n1792_;
  assign new_n1939_ = ~new_n1937_ & ~new_n1938_;
  assign new_n1940_ = new_n1936_ & ~new_n1939_;
  assign new_n1941_ = \in3[98]  & new_n1792_;
  assign new_n1942_ = \in2[98]  & ~new_n1792_;
  assign new_n1943_ = ~new_n1941_ & ~new_n1942_;
  assign new_n1944_ = \in1[98]  & new_n1787_;
  assign new_n1945_ = \in0[98]  & ~new_n1787_;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = ~new_n1943_ & new_n1946_;
  assign new_n1948_ = ~new_n1940_ & ~new_n1947_;
  assign new_n1949_ = \in1[97]  & new_n1787_;
  assign new_n1950_ = \in0[97]  & ~new_n1787_;
  assign new_n1951_ = ~new_n1949_ & ~new_n1950_;
  assign new_n1952_ = \in3[97]  & new_n1792_;
  assign new_n1953_ = \in2[97]  & ~new_n1792_;
  assign new_n1954_ = ~new_n1952_ & ~new_n1953_;
  assign new_n1955_ = new_n1951_ & ~new_n1954_;
  assign new_n1956_ = \in1[95]  & new_n1787_;
  assign new_n1957_ = \in0[95]  & ~new_n1787_;
  assign new_n1958_ = ~new_n1956_ & ~new_n1957_;
  assign new_n1959_ = \in3[95]  & new_n1792_;
  assign new_n1960_ = \in2[95]  & ~new_n1792_;
  assign new_n1961_ = ~new_n1959_ & ~new_n1960_;
  assign new_n1962_ = ~new_n1958_ & new_n1961_;
  assign new_n1963_ = new_n1958_ & ~new_n1961_;
  assign new_n1964_ = \in3[94]  & new_n1792_;
  assign new_n1965_ = \in2[94]  & ~new_n1792_;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = \in1[94]  & new_n1787_;
  assign new_n1968_ = \in0[94]  & ~new_n1787_;
  assign new_n1969_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1970_ = ~new_n1966_ & new_n1969_;
  assign new_n1971_ = ~new_n1963_ & ~new_n1970_;
  assign new_n1972_ = \in1[93]  & new_n1787_;
  assign new_n1973_ = \in0[93]  & ~new_n1787_;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1975_ = \in3[93]  & new_n1792_;
  assign new_n1976_ = \in2[93]  & ~new_n1792_;
  assign new_n1977_ = ~new_n1975_ & ~new_n1976_;
  assign new_n1978_ = new_n1974_ & ~new_n1977_;
  assign new_n1979_ = \in1[92]  & new_n1787_;
  assign new_n1980_ = \in0[92]  & ~new_n1787_;
  assign new_n1981_ = ~new_n1979_ & ~new_n1980_;
  assign new_n1982_ = \in3[92]  & new_n1792_;
  assign new_n1983_ = \in2[92]  & ~new_n1792_;
  assign new_n1984_ = ~new_n1982_ & ~new_n1983_;
  assign new_n1985_ = ~new_n1981_ & new_n1984_;
  assign new_n1986_ = ~new_n1978_ & new_n1985_;
  assign new_n1987_ = ~new_n1974_ & new_n1977_;
  assign new_n1988_ = ~new_n1986_ & ~new_n1987_;
  assign new_n1989_ = new_n1971_ & ~new_n1988_;
  assign new_n1990_ = new_n1966_ & ~new_n1969_;
  assign new_n1991_ = ~new_n1963_ & new_n1990_;
  assign new_n1992_ = \in1[87]  & new_n1787_;
  assign new_n1993_ = \in0[87]  & ~new_n1787_;
  assign new_n1994_ = ~new_n1992_ & ~new_n1993_;
  assign new_n1995_ = \in3[87]  & new_n1792_;
  assign new_n1996_ = \in2[87]  & ~new_n1792_;
  assign new_n1997_ = ~new_n1995_ & ~new_n1996_;
  assign new_n1998_ = ~new_n1994_ & new_n1997_;
  assign new_n1999_ = new_n1994_ & ~new_n1997_;
  assign new_n2000_ = \in3[86]  & new_n1792_;
  assign new_n2001_ = \in2[86]  & ~new_n1792_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = \in1[86]  & new_n1787_;
  assign new_n2004_ = \in0[86]  & ~new_n1787_;
  assign new_n2005_ = ~new_n2003_ & ~new_n2004_;
  assign new_n2006_ = ~new_n2002_ & new_n2005_;
  assign new_n2007_ = ~new_n1999_ & ~new_n2006_;
  assign new_n2008_ = \in1[85]  & new_n1787_;
  assign new_n2009_ = \in0[85]  & ~new_n1787_;
  assign new_n2010_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2011_ = \in3[85]  & new_n1792_;
  assign new_n2012_ = \in2[85]  & ~new_n1792_;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = new_n2010_ & ~new_n2013_;
  assign new_n2015_ = \in1[84]  & new_n1787_;
  assign new_n2016_ = \in0[84]  & ~new_n1787_;
  assign new_n2017_ = ~new_n2015_ & ~new_n2016_;
  assign new_n2018_ = \in3[84]  & new_n1792_;
  assign new_n2019_ = \in2[84]  & ~new_n1792_;
  assign new_n2020_ = ~new_n2018_ & ~new_n2019_;
  assign new_n2021_ = ~new_n2017_ & new_n2020_;
  assign new_n2022_ = ~new_n2014_ & new_n2021_;
  assign new_n2023_ = ~new_n2010_ & new_n2013_;
  assign new_n2024_ = ~new_n2022_ & ~new_n2023_;
  assign new_n2025_ = new_n2007_ & ~new_n2024_;
  assign new_n2026_ = new_n2002_ & ~new_n2005_;
  assign new_n2027_ = ~new_n1999_ & new_n2026_;
  assign new_n2028_ = \in3[80]  & new_n1792_;
  assign new_n2029_ = \in2[80]  & ~new_n1792_;
  assign new_n2030_ = ~new_n2028_ & ~new_n2029_;
  assign new_n2031_ = \in1[80]  & new_n1787_;
  assign new_n2032_ = \in0[80]  & ~new_n1787_;
  assign new_n2033_ = ~new_n2031_ & ~new_n2032_;
  assign new_n2034_ = ~new_n2030_ & new_n2033_;
  assign new_n2035_ = \in1[83]  & new_n1787_;
  assign new_n2036_ = \in0[83]  & ~new_n1787_;
  assign new_n2037_ = ~new_n2035_ & ~new_n2036_;
  assign new_n2038_ = \in3[83]  & new_n1792_;
  assign new_n2039_ = \in2[83]  & ~new_n1792_;
  assign new_n2040_ = ~new_n2038_ & ~new_n2039_;
  assign new_n2041_ = new_n2037_ & ~new_n2040_;
  assign new_n2042_ = \in3[82]  & new_n1792_;
  assign new_n2043_ = \in2[82]  & ~new_n1792_;
  assign new_n2044_ = ~new_n2042_ & ~new_n2043_;
  assign new_n2045_ = \in1[82]  & new_n1787_;
  assign new_n2046_ = \in0[82]  & ~new_n1787_;
  assign new_n2047_ = ~new_n2045_ & ~new_n2046_;
  assign new_n2048_ = ~new_n2044_ & new_n2047_;
  assign new_n2049_ = ~new_n2041_ & ~new_n2048_;
  assign new_n2050_ = \in1[81]  & new_n1787_;
  assign new_n2051_ = \in0[81]  & ~new_n1787_;
  assign new_n2052_ = ~new_n2050_ & ~new_n2051_;
  assign new_n2053_ = \in3[81]  & new_n1792_;
  assign new_n2054_ = \in2[81]  & ~new_n1792_;
  assign new_n2055_ = ~new_n2053_ & ~new_n2054_;
  assign new_n2056_ = new_n2052_ & ~new_n2055_;
  assign new_n2057_ = \in1[79]  & new_n1787_;
  assign new_n2058_ = \in0[79]  & ~new_n1787_;
  assign new_n2059_ = ~new_n2057_ & ~new_n2058_;
  assign new_n2060_ = \in3[79]  & new_n1792_;
  assign new_n2061_ = \in2[79]  & ~new_n1792_;
  assign new_n2062_ = ~new_n2060_ & ~new_n2061_;
  assign new_n2063_ = ~new_n2059_ & new_n2062_;
  assign new_n2064_ = new_n2059_ & ~new_n2062_;
  assign new_n2065_ = \in3[78]  & new_n1792_;
  assign new_n2066_ = \in2[78]  & ~new_n1792_;
  assign new_n2067_ = ~new_n2065_ & ~new_n2066_;
  assign new_n2068_ = \in1[78]  & new_n1787_;
  assign new_n2069_ = \in0[78]  & ~new_n1787_;
  assign new_n2070_ = ~new_n2068_ & ~new_n2069_;
  assign new_n2071_ = ~new_n2067_ & new_n2070_;
  assign new_n2072_ = ~new_n2064_ & ~new_n2071_;
  assign new_n2073_ = \in1[77]  & new_n1787_;
  assign new_n2074_ = \in0[77]  & ~new_n1787_;
  assign new_n2075_ = ~new_n2073_ & ~new_n2074_;
  assign new_n2076_ = \in3[77]  & new_n1792_;
  assign new_n2077_ = \in2[77]  & ~new_n1792_;
  assign new_n2078_ = ~new_n2076_ & ~new_n2077_;
  assign new_n2079_ = new_n2075_ & ~new_n2078_;
  assign new_n2080_ = \in1[76]  & new_n1787_;
  assign new_n2081_ = \in0[76]  & ~new_n1787_;
  assign new_n2082_ = ~new_n2080_ & ~new_n2081_;
  assign new_n2083_ = \in3[76]  & new_n1792_;
  assign new_n2084_ = \in2[76]  & ~new_n1792_;
  assign new_n2085_ = ~new_n2083_ & ~new_n2084_;
  assign new_n2086_ = ~new_n2082_ & new_n2085_;
  assign new_n2087_ = ~new_n2079_ & new_n2086_;
  assign new_n2088_ = ~new_n2075_ & new_n2078_;
  assign new_n2089_ = ~new_n2087_ & ~new_n2088_;
  assign new_n2090_ = new_n2072_ & ~new_n2089_;
  assign new_n2091_ = new_n2067_ & ~new_n2070_;
  assign new_n2092_ = ~new_n2064_ & new_n2091_;
  assign new_n2093_ = \in1[71]  & new_n1787_;
  assign new_n2094_ = \in0[71]  & ~new_n1787_;
  assign new_n2095_ = ~new_n2093_ & ~new_n2094_;
  assign new_n2096_ = \in3[71]  & new_n1792_;
  assign new_n2097_ = \in2[71]  & ~new_n1792_;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = ~new_n2095_ & new_n2098_;
  assign new_n2100_ = new_n2095_ & ~new_n2098_;
  assign new_n2101_ = \in3[70]  & new_n1792_;
  assign new_n2102_ = \in2[70]  & ~new_n1792_;
  assign new_n2103_ = ~new_n2101_ & ~new_n2102_;
  assign new_n2104_ = \in1[70]  & new_n1787_;
  assign new_n2105_ = \in0[70]  & ~new_n1787_;
  assign new_n2106_ = ~new_n2104_ & ~new_n2105_;
  assign new_n2107_ = ~new_n2103_ & new_n2106_;
  assign new_n2108_ = ~new_n2100_ & ~new_n2107_;
  assign new_n2109_ = \in1[69]  & new_n1787_;
  assign new_n2110_ = \in0[69]  & ~new_n1787_;
  assign new_n2111_ = ~new_n2109_ & ~new_n2110_;
  assign new_n2112_ = \in3[69]  & new_n1792_;
  assign new_n2113_ = \in2[69]  & ~new_n1792_;
  assign new_n2114_ = ~new_n2112_ & ~new_n2113_;
  assign new_n2115_ = new_n2111_ & ~new_n2114_;
  assign new_n2116_ = \in1[68]  & new_n1787_;
  assign new_n2117_ = \in0[68]  & ~new_n1787_;
  assign new_n2118_ = ~new_n2116_ & ~new_n2117_;
  assign new_n2119_ = \in3[68]  & new_n1792_;
  assign new_n2120_ = \in2[68]  & ~new_n1792_;
  assign new_n2121_ = ~new_n2119_ & ~new_n2120_;
  assign new_n2122_ = ~new_n2118_ & new_n2121_;
  assign new_n2123_ = ~new_n2115_ & new_n2122_;
  assign new_n2124_ = ~new_n2111_ & new_n2114_;
  assign new_n2125_ = ~new_n2123_ & ~new_n2124_;
  assign new_n2126_ = new_n2108_ & ~new_n2125_;
  assign new_n2127_ = new_n2103_ & ~new_n2106_;
  assign new_n2128_ = ~new_n2100_ & new_n2127_;
  assign new_n2129_ = \in1[67]  & new_n1787_;
  assign new_n2130_ = \in0[67]  & ~new_n1787_;
  assign new_n2131_ = ~new_n2129_ & ~new_n2130_;
  assign new_n2132_ = \in3[67]  & new_n1792_;
  assign new_n2133_ = \in2[67]  & ~new_n1792_;
  assign new_n2134_ = ~new_n2132_ & ~new_n2133_;
  assign new_n2135_ = new_n2131_ & ~new_n2134_;
  assign new_n2136_ = \in3[66]  & new_n1792_;
  assign new_n2137_ = \in2[66]  & ~new_n1792_;
  assign new_n2138_ = ~new_n2136_ & ~new_n2137_;
  assign new_n2139_ = \in1[66]  & new_n1787_;
  assign new_n2140_ = \in0[66]  & ~new_n1787_;
  assign new_n2141_ = ~new_n2139_ & ~new_n2140_;
  assign new_n2142_ = ~new_n2138_ & new_n2141_;
  assign new_n2143_ = ~new_n2135_ & ~new_n2142_;
  assign new_n2144_ = \in3[64]  & new_n1792_;
  assign new_n2145_ = \in2[64]  & ~new_n1792_;
  assign new_n2146_ = ~new_n2144_ & ~new_n2145_;
  assign new_n2147_ = \in1[64]  & new_n1787_;
  assign new_n2148_ = \in0[64]  & ~new_n1787_;
  assign new_n2149_ = ~new_n2147_ & ~new_n2148_;
  assign new_n2150_ = ~new_n2146_ & new_n2149_;
  assign new_n2151_ = \in1[65]  & new_n1787_;
  assign new_n2152_ = \in0[65]  & ~new_n1787_;
  assign new_n2153_ = ~new_n2151_ & ~new_n2152_;
  assign new_n2154_ = \in3[65]  & new_n1792_;
  assign new_n2155_ = \in2[65]  & ~new_n1792_;
  assign new_n2156_ = ~new_n2154_ & ~new_n2155_;
  assign new_n2157_ = new_n2153_ & ~new_n2156_;
  assign new_n2158_ = \in1[63]  & new_n1787_;
  assign new_n2159_ = \in0[63]  & ~new_n1787_;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = \in3[63]  & new_n1792_;
  assign new_n2162_ = \in2[63]  & ~new_n1792_;
  assign new_n2163_ = ~new_n2161_ & ~new_n2162_;
  assign new_n2164_ = ~new_n2160_ & new_n2163_;
  assign new_n2165_ = new_n2160_ & ~new_n2163_;
  assign new_n2166_ = \in3[62]  & new_n1792_;
  assign new_n2167_ = \in2[62]  & ~new_n1792_;
  assign new_n2168_ = ~new_n2166_ & ~new_n2167_;
  assign new_n2169_ = \in1[62]  & new_n1787_;
  assign new_n2170_ = \in0[62]  & ~new_n1787_;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = ~new_n2168_ & new_n2171_;
  assign new_n2173_ = ~new_n2165_ & ~new_n2172_;
  assign new_n2174_ = \in1[60]  & new_n1787_;
  assign new_n2175_ = \in0[60]  & ~new_n1787_;
  assign new_n2176_ = ~new_n2174_ & ~new_n2175_;
  assign new_n2177_ = \in3[60]  & new_n1792_;
  assign new_n2178_ = \in2[60]  & ~new_n1792_;
  assign new_n2179_ = ~new_n2177_ & ~new_n2178_;
  assign new_n2180_ = new_n2176_ & ~new_n2179_;
  assign new_n2181_ = \in1[61]  & new_n1787_;
  assign new_n2182_ = \in0[61]  & ~new_n1787_;
  assign new_n2183_ = ~new_n2181_ & ~new_n2182_;
  assign new_n2184_ = \in3[61]  & new_n1792_;
  assign new_n2185_ = \in2[61]  & ~new_n1792_;
  assign new_n2186_ = ~new_n2184_ & ~new_n2185_;
  assign new_n2187_ = new_n2183_ & ~new_n2186_;
  assign new_n2188_ = ~new_n2180_ & ~new_n2187_;
  assign new_n2189_ = new_n2173_ & new_n2188_;
  assign new_n2190_ = \in1[59]  & new_n1787_;
  assign new_n2191_ = \in0[59]  & ~new_n1787_;
  assign new_n2192_ = ~new_n2190_ & ~new_n2191_;
  assign new_n2193_ = \in3[59]  & new_n1792_;
  assign new_n2194_ = \in2[59]  & ~new_n1792_;
  assign new_n2195_ = ~new_n2193_ & ~new_n2194_;
  assign new_n2196_ = ~new_n2192_ & new_n2195_;
  assign new_n2197_ = new_n2192_ & ~new_n2195_;
  assign new_n2198_ = \in1[58]  & new_n1787_;
  assign new_n2199_ = \in0[58]  & ~new_n1787_;
  assign new_n2200_ = ~new_n2198_ & ~new_n2199_;
  assign new_n2201_ = \in3[58]  & new_n1792_;
  assign new_n2202_ = \in2[58]  & ~new_n1792_;
  assign new_n2203_ = ~new_n2201_ & ~new_n2202_;
  assign new_n2204_ = new_n2200_ & ~new_n2203_;
  assign new_n2205_ = ~new_n2197_ & ~new_n2204_;
  assign new_n2206_ = \in1[57]  & new_n1787_;
  assign new_n2207_ = \in0[57]  & ~new_n1787_;
  assign new_n2208_ = ~new_n2206_ & ~new_n2207_;
  assign new_n2209_ = \in3[57]  & new_n1792_;
  assign new_n2210_ = \in2[57]  & ~new_n1792_;
  assign new_n2211_ = ~new_n2209_ & ~new_n2210_;
  assign new_n2212_ = new_n2208_ & ~new_n2211_;
  assign new_n2213_ = \in1[56]  & new_n1787_;
  assign new_n2214_ = \in0[56]  & ~new_n1787_;
  assign new_n2215_ = ~new_n2213_ & ~new_n2214_;
  assign new_n2216_ = \in3[56]  & new_n1792_;
  assign new_n2217_ = \in2[56]  & ~new_n1792_;
  assign new_n2218_ = ~new_n2216_ & ~new_n2217_;
  assign new_n2219_ = ~new_n2215_ & new_n2218_;
  assign new_n2220_ = ~new_n2212_ & new_n2219_;
  assign new_n2221_ = ~new_n2208_ & new_n2211_;
  assign new_n2222_ = ~new_n2220_ & ~new_n2221_;
  assign new_n2223_ = ~new_n2200_ & new_n2203_;
  assign new_n2224_ = new_n2222_ & ~new_n2223_;
  assign new_n2225_ = new_n2205_ & ~new_n2224_;
  assign new_n2226_ = ~new_n2196_ & ~new_n2225_;
  assign new_n2227_ = new_n2189_ & ~new_n2226_;
  assign new_n2228_ = ~new_n2176_ & new_n2179_;
  assign new_n2229_ = ~new_n2187_ & new_n2228_;
  assign new_n2230_ = ~new_n2183_ & new_n2186_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = new_n2173_ & ~new_n2231_;
  assign new_n2233_ = new_n2168_ & ~new_n2171_;
  assign new_n2234_ = ~new_n2165_ & new_n2233_;
  assign new_n2235_ = \in1[47]  & new_n1787_;
  assign new_n2236_ = \in0[47]  & ~new_n1787_;
  assign new_n2237_ = ~new_n2235_ & ~new_n2236_;
  assign new_n2238_ = \in3[47]  & new_n1792_;
  assign new_n2239_ = \in2[47]  & ~new_n1792_;
  assign new_n2240_ = ~new_n2238_ & ~new_n2239_;
  assign new_n2241_ = ~new_n2237_ & new_n2240_;
  assign new_n2242_ = new_n2237_ & ~new_n2240_;
  assign new_n2243_ = \in3[46]  & new_n1792_;
  assign new_n2244_ = \in2[46]  & ~new_n1792_;
  assign new_n2245_ = ~new_n2243_ & ~new_n2244_;
  assign new_n2246_ = \in1[46]  & new_n1787_;
  assign new_n2247_ = \in0[46]  & ~new_n1787_;
  assign new_n2248_ = ~new_n2246_ & ~new_n2247_;
  assign new_n2249_ = ~new_n2245_ & new_n2248_;
  assign new_n2250_ = ~new_n2242_ & ~new_n2249_;
  assign new_n2251_ = \in1[44]  & new_n1787_;
  assign new_n2252_ = \in0[44]  & ~new_n1787_;
  assign new_n2253_ = ~new_n2251_ & ~new_n2252_;
  assign new_n2254_ = \in3[44]  & new_n1792_;
  assign new_n2255_ = \in2[44]  & ~new_n1792_;
  assign new_n2256_ = ~new_n2254_ & ~new_n2255_;
  assign new_n2257_ = new_n2253_ & ~new_n2256_;
  assign new_n2258_ = \in1[45]  & new_n1787_;
  assign new_n2259_ = \in0[45]  & ~new_n1787_;
  assign new_n2260_ = ~new_n2258_ & ~new_n2259_;
  assign new_n2261_ = \in3[45]  & new_n1792_;
  assign new_n2262_ = \in2[45]  & ~new_n1792_;
  assign new_n2263_ = ~new_n2261_ & ~new_n2262_;
  assign new_n2264_ = new_n2260_ & ~new_n2263_;
  assign new_n2265_ = ~new_n2257_ & ~new_n2264_;
  assign new_n2266_ = new_n2250_ & new_n2265_;
  assign new_n2267_ = \in1[43]  & new_n1787_;
  assign new_n2268_ = \in0[43]  & ~new_n1787_;
  assign new_n2269_ = ~new_n2267_ & ~new_n2268_;
  assign new_n2270_ = \in3[43]  & new_n1792_;
  assign new_n2271_ = \in2[43]  & ~new_n1792_;
  assign new_n2272_ = ~new_n2270_ & ~new_n2271_;
  assign new_n2273_ = ~new_n2269_ & new_n2272_;
  assign new_n2274_ = new_n2269_ & ~new_n2272_;
  assign new_n2275_ = \in1[42]  & new_n1787_;
  assign new_n2276_ = \in0[42]  & ~new_n1787_;
  assign new_n2277_ = ~new_n2275_ & ~new_n2276_;
  assign new_n2278_ = \in3[42]  & new_n1792_;
  assign new_n2279_ = \in2[42]  & ~new_n1792_;
  assign new_n2280_ = ~new_n2278_ & ~new_n2279_;
  assign new_n2281_ = new_n2277_ & ~new_n2280_;
  assign new_n2282_ = ~new_n2274_ & ~new_n2281_;
  assign new_n2283_ = \in1[41]  & new_n1787_;
  assign new_n2284_ = \in0[41]  & ~new_n1787_;
  assign new_n2285_ = ~new_n2283_ & ~new_n2284_;
  assign new_n2286_ = \in3[41]  & new_n1792_;
  assign new_n2287_ = \in2[41]  & ~new_n1792_;
  assign new_n2288_ = ~new_n2286_ & ~new_n2287_;
  assign new_n2289_ = new_n2285_ & ~new_n2288_;
  assign new_n2290_ = \in1[40]  & new_n1787_;
  assign new_n2291_ = \in0[40]  & ~new_n1787_;
  assign new_n2292_ = ~new_n2290_ & ~new_n2291_;
  assign new_n2293_ = \in3[40]  & new_n1792_;
  assign new_n2294_ = \in2[40]  & ~new_n1792_;
  assign new_n2295_ = ~new_n2293_ & ~new_n2294_;
  assign new_n2296_ = ~new_n2292_ & new_n2295_;
  assign new_n2297_ = ~new_n2289_ & new_n2296_;
  assign new_n2298_ = ~new_n2285_ & new_n2288_;
  assign new_n2299_ = ~new_n2297_ & ~new_n2298_;
  assign new_n2300_ = ~new_n2277_ & new_n2280_;
  assign new_n2301_ = new_n2299_ & ~new_n2300_;
  assign new_n2302_ = new_n2282_ & ~new_n2301_;
  assign new_n2303_ = ~new_n2273_ & ~new_n2302_;
  assign new_n2304_ = new_n2266_ & ~new_n2303_;
  assign new_n2305_ = ~new_n2253_ & new_n2256_;
  assign new_n2306_ = ~new_n2264_ & new_n2305_;
  assign new_n2307_ = ~new_n2260_ & new_n2263_;
  assign new_n2308_ = ~new_n2306_ & ~new_n2307_;
  assign new_n2309_ = new_n2250_ & ~new_n2308_;
  assign new_n2310_ = new_n2245_ & ~new_n2248_;
  assign new_n2311_ = ~new_n2242_ & new_n2310_;
  assign new_n2312_ = \in3[32]  & new_n1792_;
  assign new_n2313_ = \in2[32]  & ~new_n1792_;
  assign new_n2314_ = ~new_n2312_ & ~new_n2313_;
  assign new_n2315_ = \in1[32]  & new_n1787_;
  assign new_n2316_ = \in0[32]  & ~new_n1787_;
  assign new_n2317_ = ~new_n2315_ & ~new_n2316_;
  assign new_n2318_ = ~new_n2314_ & new_n2317_;
  assign new_n2319_ = \in1[31]  & new_n1787_;
  assign new_n2320_ = \in0[31]  & ~new_n1787_;
  assign new_n2321_ = ~new_n2319_ & ~new_n2320_;
  assign new_n2322_ = \in3[31]  & new_n1792_;
  assign new_n2323_ = \in2[31]  & ~new_n1792_;
  assign new_n2324_ = ~new_n2322_ & ~new_n2323_;
  assign new_n2325_ = new_n2321_ & ~new_n2324_;
  assign new_n2326_ = \in1[30]  & new_n1787_;
  assign new_n2327_ = \in0[30]  & ~new_n1787_;
  assign new_n2328_ = ~new_n2326_ & ~new_n2327_;
  assign new_n2329_ = \in3[30]  & new_n1792_;
  assign new_n2330_ = \in2[30]  & ~new_n1792_;
  assign new_n2331_ = ~new_n2329_ & ~new_n2330_;
  assign new_n2332_ = new_n2328_ & ~new_n2331_;
  assign new_n2333_ = \in1[29]  & new_n1787_;
  assign new_n2334_ = \in0[29]  & ~new_n1787_;
  assign new_n2335_ = ~new_n2333_ & ~new_n2334_;
  assign new_n2336_ = \in3[29]  & new_n1792_;
  assign new_n2337_ = \in2[29]  & ~new_n1792_;
  assign new_n2338_ = ~new_n2336_ & ~new_n2337_;
  assign new_n2339_ = new_n2335_ & ~new_n2338_;
  assign new_n2340_ = \in1[28]  & new_n1787_;
  assign new_n2341_ = \in0[28]  & ~new_n1787_;
  assign new_n2342_ = ~new_n2340_ & ~new_n2341_;
  assign new_n2343_ = \in3[28]  & new_n1792_;
  assign new_n2344_ = \in2[28]  & ~new_n1792_;
  assign new_n2345_ = ~new_n2343_ & ~new_n2344_;
  assign new_n2346_ = new_n2342_ & ~new_n2345_;
  assign new_n2347_ = \in1[27]  & new_n1787_;
  assign new_n2348_ = \in0[27]  & ~new_n1787_;
  assign new_n2349_ = ~new_n2347_ & ~new_n2348_;
  assign new_n2350_ = \in3[27]  & new_n1792_;
  assign new_n2351_ = \in2[27]  & ~new_n1792_;
  assign new_n2352_ = ~new_n2350_ & ~new_n2351_;
  assign new_n2353_ = new_n2349_ & ~new_n2352_;
  assign new_n2354_ = \in1[26]  & new_n1787_;
  assign new_n2355_ = \in0[26]  & ~new_n1787_;
  assign new_n2356_ = ~new_n2354_ & ~new_n2355_;
  assign new_n2357_ = \in3[26]  & new_n1792_;
  assign new_n2358_ = \in2[26]  & ~new_n1792_;
  assign new_n2359_ = ~new_n2357_ & ~new_n2358_;
  assign new_n2360_ = new_n2356_ & ~new_n2359_;
  assign new_n2361_ = \in3[25]  & new_n1792_;
  assign new_n2362_ = \in2[25]  & ~new_n1792_;
  assign new_n2363_ = ~new_n2361_ & ~new_n2362_;
  assign new_n2364_ = \in3[24]  & new_n1792_;
  assign new_n2365_ = \in2[24]  & ~new_n1792_;
  assign new_n2366_ = ~new_n2364_ & ~new_n2365_;
  assign new_n2367_ = \in1[23]  & new_n1787_;
  assign new_n2368_ = \in0[23]  & ~new_n1787_;
  assign new_n2369_ = ~new_n2367_ & ~new_n2368_;
  assign new_n2370_ = \in3[23]  & new_n1792_;
  assign new_n2371_ = \in2[23]  & ~new_n1792_;
  assign new_n2372_ = ~new_n2370_ & ~new_n2371_;
  assign new_n2373_ = new_n2369_ & ~new_n2372_;
  assign new_n2374_ = \in1[22]  & new_n1787_;
  assign new_n2375_ = \in0[22]  & ~new_n1787_;
  assign new_n2376_ = ~new_n2374_ & ~new_n2375_;
  assign new_n2377_ = \in3[22]  & new_n1792_;
  assign new_n2378_ = \in2[22]  & ~new_n1792_;
  assign new_n2379_ = ~new_n2377_ & ~new_n2378_;
  assign new_n2380_ = new_n2376_ & ~new_n2379_;
  assign new_n2381_ = \in1[21]  & new_n1787_;
  assign new_n2382_ = \in0[21]  & ~new_n1787_;
  assign new_n2383_ = ~new_n2381_ & ~new_n2382_;
  assign new_n2384_ = \in3[21]  & new_n1792_;
  assign new_n2385_ = \in2[21]  & ~new_n1792_;
  assign new_n2386_ = ~new_n2384_ & ~new_n2385_;
  assign new_n2387_ = new_n2383_ & ~new_n2386_;
  assign new_n2388_ = \in1[20]  & new_n1787_;
  assign new_n2389_ = \in0[20]  & ~new_n1787_;
  assign new_n2390_ = ~new_n2388_ & ~new_n2389_;
  assign new_n2391_ = \in3[20]  & new_n1792_;
  assign new_n2392_ = \in2[20]  & ~new_n1792_;
  assign new_n2393_ = ~new_n2391_ & ~new_n2392_;
  assign new_n2394_ = new_n2390_ & ~new_n2393_;
  assign new_n2395_ = \in1[19]  & new_n1787_;
  assign new_n2396_ = \in0[19]  & ~new_n1787_;
  assign new_n2397_ = ~new_n2395_ & ~new_n2396_;
  assign new_n2398_ = \in3[19]  & new_n1792_;
  assign new_n2399_ = \in2[19]  & ~new_n1792_;
  assign new_n2400_ = ~new_n2398_ & ~new_n2399_;
  assign new_n2401_ = new_n2397_ & ~new_n2400_;
  assign new_n2402_ = \in1[18]  & new_n1787_;
  assign new_n2403_ = \in0[18]  & ~new_n1787_;
  assign new_n2404_ = ~new_n2402_ & ~new_n2403_;
  assign new_n2405_ = \in3[18]  & new_n1792_;
  assign new_n2406_ = \in2[18]  & ~new_n1792_;
  assign new_n2407_ = ~new_n2405_ & ~new_n2406_;
  assign new_n2408_ = new_n2404_ & ~new_n2407_;
  assign new_n2409_ = \in3[17]  & new_n1792_;
  assign new_n2410_ = \in2[17]  & ~new_n1792_;
  assign new_n2411_ = ~new_n2409_ & ~new_n2410_;
  assign new_n2412_ = \in3[16]  & new_n1792_;
  assign new_n2413_ = \in2[16]  & ~new_n1792_;
  assign new_n2414_ = ~new_n2412_ & ~new_n2413_;
  assign new_n2415_ = \in1[15]  & new_n1787_;
  assign new_n2416_ = \in0[15]  & ~new_n1787_;
  assign new_n2417_ = ~new_n2415_ & ~new_n2416_;
  assign new_n2418_ = \in3[15]  & new_n1792_;
  assign new_n2419_ = \in2[15]  & ~new_n1792_;
  assign new_n2420_ = ~new_n2418_ & ~new_n2419_;
  assign new_n2421_ = new_n2417_ & ~new_n2420_;
  assign new_n2422_ = \in1[14]  & new_n1787_;
  assign new_n2423_ = \in0[14]  & ~new_n1787_;
  assign new_n2424_ = ~new_n2422_ & ~new_n2423_;
  assign new_n2425_ = \in3[14]  & new_n1792_;
  assign new_n2426_ = \in2[14]  & ~new_n1792_;
  assign new_n2427_ = ~new_n2425_ & ~new_n2426_;
  assign new_n2428_ = new_n2424_ & ~new_n2427_;
  assign new_n2429_ = \in1[13]  & new_n1787_;
  assign new_n2430_ = \in0[13]  & ~new_n1787_;
  assign new_n2431_ = ~new_n2429_ & ~new_n2430_;
  assign new_n2432_ = \in3[13]  & new_n1792_;
  assign new_n2433_ = \in2[13]  & ~new_n1792_;
  assign new_n2434_ = ~new_n2432_ & ~new_n2433_;
  assign new_n2435_ = new_n2431_ & ~new_n2434_;
  assign new_n2436_ = \in1[12]  & new_n1787_;
  assign new_n2437_ = \in0[12]  & ~new_n1787_;
  assign new_n2438_ = ~new_n2436_ & ~new_n2437_;
  assign new_n2439_ = \in3[12]  & new_n1792_;
  assign new_n2440_ = \in2[12]  & ~new_n1792_;
  assign new_n2441_ = ~new_n2439_ & ~new_n2440_;
  assign new_n2442_ = new_n2438_ & ~new_n2441_;
  assign new_n2443_ = \in1[11]  & new_n1787_;
  assign new_n2444_ = \in0[11]  & ~new_n1787_;
  assign new_n2445_ = ~new_n2443_ & ~new_n2444_;
  assign new_n2446_ = \in3[11]  & new_n1792_;
  assign new_n2447_ = \in2[11]  & ~new_n1792_;
  assign new_n2448_ = ~new_n2446_ & ~new_n2447_;
  assign new_n2449_ = new_n2445_ & ~new_n2448_;
  assign new_n2450_ = \in1[10]  & new_n1787_;
  assign new_n2451_ = \in0[10]  & ~new_n1787_;
  assign new_n2452_ = ~new_n2450_ & ~new_n2451_;
  assign new_n2453_ = \in3[10]  & new_n1792_;
  assign new_n2454_ = \in2[10]  & ~new_n1792_;
  assign new_n2455_ = ~new_n2453_ & ~new_n2454_;
  assign new_n2456_ = new_n2452_ & ~new_n2455_;
  assign new_n2457_ = \in3[9]  & new_n1792_;
  assign new_n2458_ = \in2[9]  & ~new_n1792_;
  assign new_n2459_ = ~new_n2457_ & ~new_n2458_;
  assign new_n2460_ = \in3[8]  & new_n1792_;
  assign new_n2461_ = \in2[8]  & ~new_n1792_;
  assign new_n2462_ = ~new_n2460_ & ~new_n2461_;
  assign new_n2463_ = \in1[7]  & new_n1787_;
  assign new_n2464_ = \in0[7]  & ~new_n1787_;
  assign new_n2465_ = ~new_n2463_ & ~new_n2464_;
  assign new_n2466_ = \in3[7]  & new_n1792_;
  assign new_n2467_ = \in2[7]  & ~new_n1792_;
  assign new_n2468_ = ~new_n2466_ & ~new_n2467_;
  assign new_n2469_ = new_n2465_ & ~new_n2468_;
  assign new_n2470_ = \in3[6]  & new_n1792_;
  assign new_n2471_ = \in2[6]  & ~new_n1792_;
  assign new_n2472_ = ~new_n2470_ & ~new_n2471_;
  assign new_n2473_ = \in1[6]  & new_n1787_;
  assign new_n2474_ = \in0[6]  & ~new_n1787_;
  assign new_n2475_ = ~new_n2473_ & ~new_n2474_;
  assign new_n2476_ = \in3[5]  & new_n1792_;
  assign new_n2477_ = \in2[5]  & ~new_n1792_;
  assign new_n2478_ = ~new_n2476_ & ~new_n2477_;
  assign new_n2479_ = \in1[5]  & new_n1787_;
  assign new_n2480_ = \in0[5]  & ~new_n1787_;
  assign new_n2481_ = ~new_n2479_ & ~new_n2480_;
  assign new_n2482_ = \in3[4]  & new_n1792_;
  assign new_n2483_ = \in2[4]  & ~new_n1792_;
  assign new_n2484_ = ~new_n2482_ & ~new_n2483_;
  assign new_n2485_ = \in1[4]  & new_n1787_;
  assign new_n2486_ = \in0[4]  & ~new_n1787_;
  assign new_n2487_ = ~new_n2485_ & ~new_n2486_;
  assign new_n2488_ = \in1[3]  & new_n1787_;
  assign new_n2489_ = \in0[3]  & ~new_n1787_;
  assign new_n2490_ = ~new_n2488_ & ~new_n2489_;
  assign new_n2491_ = \in3[3]  & new_n1792_;
  assign new_n2492_ = \in2[3]  & ~new_n1792_;
  assign new_n2493_ = ~new_n2491_ & ~new_n2492_;
  assign new_n2494_ = new_n2490_ & ~new_n2493_;
  assign new_n2495_ = \in3[1]  & new_n1792_;
  assign new_n2496_ = \in2[1]  & ~new_n1792_;
  assign new_n2497_ = ~new_n2495_ & ~new_n2496_;
  assign new_n2498_ = \in1[0]  & new_n1787_;
  assign new_n2499_ = \in0[0]  & ~new_n1787_;
  assign new_n2500_ = ~new_n2498_ & ~new_n2499_;
  assign new_n2501_ = \in3[0]  & new_n1792_;
  assign new_n2502_ = \in2[0]  & ~new_n1792_;
  assign new_n2503_ = ~new_n2501_ & ~new_n2502_;
  assign new_n2504_ = ~new_n2500_ & new_n2503_;
  assign new_n2505_ = new_n2497_ & new_n2504_;
  assign new_n2506_ = \in1[1]  & new_n1787_;
  assign new_n2507_ = \in0[1]  & ~new_n1787_;
  assign new_n2508_ = ~new_n2506_ & ~new_n2507_;
  assign new_n2509_ = ~new_n2505_ & new_n2508_;
  assign new_n2510_ = \in1[2]  & new_n1787_;
  assign new_n2511_ = \in0[2]  & ~new_n1787_;
  assign new_n2512_ = ~new_n2510_ & ~new_n2511_;
  assign new_n2513_ = \in3[2]  & new_n1792_;
  assign new_n2514_ = \in2[2]  & ~new_n1792_;
  assign new_n2515_ = ~new_n2513_ & ~new_n2514_;
  assign new_n2516_ = new_n2512_ & ~new_n2515_;
  assign new_n2517_ = ~new_n2497_ & ~new_n2504_;
  assign new_n2518_ = ~new_n2516_ & ~new_n2517_;
  assign new_n2519_ = ~new_n2509_ & new_n2518_;
  assign new_n2520_ = ~new_n2512_ & new_n2515_;
  assign new_n2521_ = ~new_n2519_ & ~new_n2520_;
  assign new_n2522_ = ~new_n2494_ & ~new_n2521_;
  assign new_n2523_ = ~new_n2490_ & new_n2493_;
  assign new_n2524_ = ~new_n2522_ & ~new_n2523_;
  assign new_n2525_ = new_n2487_ & new_n2524_;
  assign new_n2526_ = new_n2484_ & ~new_n2525_;
  assign new_n2527_ = ~new_n2487_ & ~new_n2524_;
  assign new_n2528_ = ~new_n2526_ & ~new_n2527_;
  assign new_n2529_ = new_n2481_ & new_n2528_;
  assign new_n2530_ = new_n2478_ & ~new_n2529_;
  assign new_n2531_ = ~new_n2481_ & ~new_n2528_;
  assign new_n2532_ = ~new_n2530_ & ~new_n2531_;
  assign new_n2533_ = new_n2475_ & new_n2532_;
  assign new_n2534_ = new_n2472_ & ~new_n2533_;
  assign new_n2535_ = ~new_n2475_ & ~new_n2532_;
  assign new_n2536_ = ~new_n2534_ & ~new_n2535_;
  assign new_n2537_ = ~new_n2469_ & ~new_n2536_;
  assign new_n2538_ = ~new_n2465_ & new_n2468_;
  assign new_n2539_ = ~new_n2537_ & ~new_n2538_;
  assign new_n2540_ = \in1[8]  & new_n1787_;
  assign new_n2541_ = \in0[8]  & ~new_n1787_;
  assign new_n2542_ = ~new_n2540_ & ~new_n2541_;
  assign new_n2543_ = new_n2539_ & new_n2542_;
  assign new_n2544_ = new_n2462_ & ~new_n2543_;
  assign new_n2545_ = ~new_n2539_ & ~new_n2542_;
  assign new_n2546_ = ~new_n2544_ & ~new_n2545_;
  assign new_n2547_ = \in1[9]  & new_n1787_;
  assign new_n2548_ = \in0[9]  & ~new_n1787_;
  assign new_n2549_ = ~new_n2547_ & ~new_n2548_;
  assign new_n2550_ = new_n2546_ & new_n2549_;
  assign new_n2551_ = new_n2459_ & ~new_n2550_;
  assign new_n2552_ = ~new_n2546_ & ~new_n2549_;
  assign new_n2553_ = ~new_n2551_ & ~new_n2552_;
  assign new_n2554_ = ~new_n2456_ & ~new_n2553_;
  assign new_n2555_ = ~new_n2452_ & new_n2455_;
  assign new_n2556_ = ~new_n2554_ & ~new_n2555_;
  assign new_n2557_ = ~new_n2449_ & ~new_n2556_;
  assign new_n2558_ = ~new_n2445_ & new_n2448_;
  assign new_n2559_ = ~new_n2557_ & ~new_n2558_;
  assign new_n2560_ = ~new_n2442_ & ~new_n2559_;
  assign new_n2561_ = ~new_n2438_ & new_n2441_;
  assign new_n2562_ = ~new_n2560_ & ~new_n2561_;
  assign new_n2563_ = ~new_n2435_ & ~new_n2562_;
  assign new_n2564_ = ~new_n2431_ & new_n2434_;
  assign new_n2565_ = ~new_n2563_ & ~new_n2564_;
  assign new_n2566_ = ~new_n2428_ & ~new_n2565_;
  assign new_n2567_ = ~new_n2424_ & new_n2427_;
  assign new_n2568_ = ~new_n2566_ & ~new_n2567_;
  assign new_n2569_ = ~new_n2421_ & ~new_n2568_;
  assign new_n2570_ = ~new_n2417_ & new_n2420_;
  assign new_n2571_ = ~new_n2569_ & ~new_n2570_;
  assign new_n2572_ = \in1[16]  & new_n1787_;
  assign new_n2573_ = \in0[16]  & ~new_n1787_;
  assign new_n2574_ = ~new_n2572_ & ~new_n2573_;
  assign new_n2575_ = new_n2571_ & new_n2574_;
  assign new_n2576_ = new_n2414_ & ~new_n2575_;
  assign new_n2577_ = ~new_n2571_ & ~new_n2574_;
  assign new_n2578_ = ~new_n2576_ & ~new_n2577_;
  assign new_n2579_ = \in1[17]  & new_n1787_;
  assign new_n2580_ = \in0[17]  & ~new_n1787_;
  assign new_n2581_ = ~new_n2579_ & ~new_n2580_;
  assign new_n2582_ = new_n2578_ & new_n2581_;
  assign new_n2583_ = new_n2411_ & ~new_n2582_;
  assign new_n2584_ = ~new_n2578_ & ~new_n2581_;
  assign new_n2585_ = ~new_n2583_ & ~new_n2584_;
  assign new_n2586_ = ~new_n2408_ & ~new_n2585_;
  assign new_n2587_ = ~new_n2404_ & new_n2407_;
  assign new_n2588_ = ~new_n2586_ & ~new_n2587_;
  assign new_n2589_ = ~new_n2401_ & ~new_n2588_;
  assign new_n2590_ = ~new_n2397_ & new_n2400_;
  assign new_n2591_ = ~new_n2589_ & ~new_n2590_;
  assign new_n2592_ = ~new_n2394_ & ~new_n2591_;
  assign new_n2593_ = ~new_n2390_ & new_n2393_;
  assign new_n2594_ = ~new_n2592_ & ~new_n2593_;
  assign new_n2595_ = ~new_n2387_ & ~new_n2594_;
  assign new_n2596_ = ~new_n2383_ & new_n2386_;
  assign new_n2597_ = ~new_n2595_ & ~new_n2596_;
  assign new_n2598_ = ~new_n2380_ & ~new_n2597_;
  assign new_n2599_ = ~new_n2376_ & new_n2379_;
  assign new_n2600_ = ~new_n2598_ & ~new_n2599_;
  assign new_n2601_ = ~new_n2373_ & ~new_n2600_;
  assign new_n2602_ = ~new_n2369_ & new_n2372_;
  assign new_n2603_ = ~new_n2601_ & ~new_n2602_;
  assign new_n2604_ = \in1[24]  & new_n1787_;
  assign new_n2605_ = \in0[24]  & ~new_n1787_;
  assign new_n2606_ = ~new_n2604_ & ~new_n2605_;
  assign new_n2607_ = new_n2603_ & new_n2606_;
  assign new_n2608_ = new_n2366_ & ~new_n2607_;
  assign new_n2609_ = ~new_n2603_ & ~new_n2606_;
  assign new_n2610_ = ~new_n2608_ & ~new_n2609_;
  assign new_n2611_ = \in1[25]  & new_n1787_;
  assign new_n2612_ = \in0[25]  & ~new_n1787_;
  assign new_n2613_ = ~new_n2611_ & ~new_n2612_;
  assign new_n2614_ = new_n2610_ & new_n2613_;
  assign new_n2615_ = new_n2363_ & ~new_n2614_;
  assign new_n2616_ = ~new_n2610_ & ~new_n2613_;
  assign new_n2617_ = ~new_n2615_ & ~new_n2616_;
  assign new_n2618_ = ~new_n2360_ & ~new_n2617_;
  assign new_n2619_ = ~new_n2356_ & new_n2359_;
  assign new_n2620_ = ~new_n2618_ & ~new_n2619_;
  assign new_n2621_ = ~new_n2353_ & ~new_n2620_;
  assign new_n2622_ = ~new_n2349_ & new_n2352_;
  assign new_n2623_ = ~new_n2621_ & ~new_n2622_;
  assign new_n2624_ = ~new_n2346_ & ~new_n2623_;
  assign new_n2625_ = ~new_n2342_ & new_n2345_;
  assign new_n2626_ = ~new_n2624_ & ~new_n2625_;
  assign new_n2627_ = ~new_n2339_ & ~new_n2626_;
  assign new_n2628_ = ~new_n2335_ & new_n2338_;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = ~new_n2332_ & ~new_n2629_;
  assign new_n2631_ = ~new_n2328_ & new_n2331_;
  assign new_n2632_ = ~new_n2630_ & ~new_n2631_;
  assign new_n2633_ = ~new_n2325_ & ~new_n2632_;
  assign new_n2634_ = ~new_n2321_ & new_n2324_;
  assign new_n2635_ = ~new_n2633_ & ~new_n2634_;
  assign new_n2636_ = \in1[39]  & new_n1787_;
  assign new_n2637_ = \in0[39]  & ~new_n1787_;
  assign new_n2638_ = ~new_n2636_ & ~new_n2637_;
  assign new_n2639_ = \in3[39]  & new_n1792_;
  assign new_n2640_ = \in2[39]  & ~new_n1792_;
  assign new_n2641_ = ~new_n2639_ & ~new_n2640_;
  assign new_n2642_ = new_n2638_ & ~new_n2641_;
  assign new_n2643_ = \in3[38]  & new_n1792_;
  assign new_n2644_ = \in2[38]  & ~new_n1792_;
  assign new_n2645_ = ~new_n2643_ & ~new_n2644_;
  assign new_n2646_ = \in1[38]  & new_n1787_;
  assign new_n2647_ = \in0[38]  & ~new_n1787_;
  assign new_n2648_ = ~new_n2646_ & ~new_n2647_;
  assign new_n2649_ = ~new_n2645_ & new_n2648_;
  assign new_n2650_ = ~new_n2642_ & ~new_n2649_;
  assign new_n2651_ = \in1[36]  & new_n1787_;
  assign new_n2652_ = \in0[36]  & ~new_n1787_;
  assign new_n2653_ = ~new_n2651_ & ~new_n2652_;
  assign new_n2654_ = \in3[36]  & new_n1792_;
  assign new_n2655_ = \in2[36]  & ~new_n1792_;
  assign new_n2656_ = ~new_n2654_ & ~new_n2655_;
  assign new_n2657_ = new_n2653_ & ~new_n2656_;
  assign new_n2658_ = \in1[37]  & new_n1787_;
  assign new_n2659_ = \in0[37]  & ~new_n1787_;
  assign new_n2660_ = ~new_n2658_ & ~new_n2659_;
  assign new_n2661_ = \in3[37]  & new_n1792_;
  assign new_n2662_ = \in2[37]  & ~new_n1792_;
  assign new_n2663_ = ~new_n2661_ & ~new_n2662_;
  assign new_n2664_ = new_n2660_ & ~new_n2663_;
  assign new_n2665_ = ~new_n2657_ & ~new_n2664_;
  assign new_n2666_ = new_n2650_ & new_n2665_;
  assign new_n2667_ = \in1[33]  & new_n1787_;
  assign new_n2668_ = \in0[33]  & ~new_n1787_;
  assign new_n2669_ = ~new_n2667_ & ~new_n2668_;
  assign new_n2670_ = \in3[33]  & new_n1792_;
  assign new_n2671_ = \in2[33]  & ~new_n1792_;
  assign new_n2672_ = ~new_n2670_ & ~new_n2671_;
  assign new_n2673_ = new_n2669_ & ~new_n2672_;
  assign new_n2674_ = \in1[35]  & new_n1787_;
  assign new_n2675_ = \in0[35]  & ~new_n1787_;
  assign new_n2676_ = ~new_n2674_ & ~new_n2675_;
  assign new_n2677_ = \in3[35]  & new_n1792_;
  assign new_n2678_ = \in2[35]  & ~new_n1792_;
  assign new_n2679_ = ~new_n2677_ & ~new_n2678_;
  assign new_n2680_ = new_n2676_ & ~new_n2679_;
  assign new_n2681_ = \in3[34]  & new_n1792_;
  assign new_n2682_ = \in2[34]  & ~new_n1792_;
  assign new_n2683_ = ~new_n2681_ & ~new_n2682_;
  assign new_n2684_ = \in1[34]  & new_n1787_;
  assign new_n2685_ = \in0[34]  & ~new_n1787_;
  assign new_n2686_ = ~new_n2684_ & ~new_n2685_;
  assign new_n2687_ = ~new_n2683_ & new_n2686_;
  assign new_n2688_ = ~new_n2680_ & ~new_n2687_;
  assign new_n2689_ = ~new_n2673_ & new_n2688_;
  assign new_n2690_ = new_n2666_ & new_n2689_;
  assign new_n2691_ = ~new_n2635_ & new_n2690_;
  assign new_n2692_ = ~new_n2318_ & new_n2691_;
  assign new_n2693_ = ~new_n2638_ & new_n2641_;
  assign new_n2694_ = ~new_n2653_ & new_n2656_;
  assign new_n2695_ = ~new_n2664_ & new_n2694_;
  assign new_n2696_ = ~new_n2660_ & new_n2663_;
  assign new_n2697_ = ~new_n2695_ & ~new_n2696_;
  assign new_n2698_ = new_n2650_ & ~new_n2697_;
  assign new_n2699_ = ~new_n2642_ & new_n2645_;
  assign new_n2700_ = ~new_n2648_ & new_n2699_;
  assign new_n2701_ = ~new_n2676_ & new_n2679_;
  assign new_n2702_ = ~new_n2680_ & new_n2683_;
  assign new_n2703_ = ~new_n2686_ & new_n2702_;
  assign new_n2704_ = new_n2314_ & ~new_n2317_;
  assign new_n2705_ = ~new_n2669_ & new_n2672_;
  assign new_n2706_ = ~new_n2704_ & ~new_n2705_;
  assign new_n2707_ = new_n2689_ & ~new_n2706_;
  assign new_n2708_ = ~new_n2703_ & ~new_n2707_;
  assign new_n2709_ = ~new_n2701_ & new_n2708_;
  assign new_n2710_ = new_n2666_ & ~new_n2709_;
  assign new_n2711_ = ~new_n2700_ & ~new_n2710_;
  assign new_n2712_ = ~new_n2698_ & new_n2711_;
  assign new_n2713_ = ~new_n2693_ & new_n2712_;
  assign new_n2714_ = ~new_n2692_ & new_n2713_;
  assign new_n2715_ = new_n2292_ & ~new_n2295_;
  assign new_n2716_ = ~new_n2289_ & ~new_n2715_;
  assign new_n2717_ = new_n2282_ & new_n2716_;
  assign new_n2718_ = new_n2266_ & new_n2717_;
  assign new_n2719_ = ~new_n2714_ & new_n2718_;
  assign new_n2720_ = ~new_n2311_ & ~new_n2719_;
  assign new_n2721_ = ~new_n2309_ & new_n2720_;
  assign new_n2722_ = ~new_n2304_ & new_n2721_;
  assign new_n2723_ = ~new_n2241_ & new_n2722_;
  assign new_n2724_ = \in3[48]  & new_n1792_;
  assign new_n2725_ = \in2[48]  & ~new_n1792_;
  assign new_n2726_ = ~new_n2724_ & ~new_n2725_;
  assign new_n2727_ = \in1[48]  & new_n1787_;
  assign new_n2728_ = \in0[48]  & ~new_n1787_;
  assign new_n2729_ = ~new_n2727_ & ~new_n2728_;
  assign new_n2730_ = ~new_n2726_ & new_n2729_;
  assign new_n2731_ = \in1[55]  & new_n1787_;
  assign new_n2732_ = \in0[55]  & ~new_n1787_;
  assign new_n2733_ = ~new_n2731_ & ~new_n2732_;
  assign new_n2734_ = \in3[55]  & new_n1792_;
  assign new_n2735_ = \in2[55]  & ~new_n1792_;
  assign new_n2736_ = ~new_n2734_ & ~new_n2735_;
  assign new_n2737_ = new_n2733_ & ~new_n2736_;
  assign new_n2738_ = \in3[54]  & new_n1792_;
  assign new_n2739_ = \in2[54]  & ~new_n1792_;
  assign new_n2740_ = ~new_n2738_ & ~new_n2739_;
  assign new_n2741_ = \in1[54]  & new_n1787_;
  assign new_n2742_ = \in0[54]  & ~new_n1787_;
  assign new_n2743_ = ~new_n2741_ & ~new_n2742_;
  assign new_n2744_ = ~new_n2740_ & new_n2743_;
  assign new_n2745_ = ~new_n2737_ & ~new_n2744_;
  assign new_n2746_ = \in1[53]  & new_n1787_;
  assign new_n2747_ = \in0[53]  & ~new_n1787_;
  assign new_n2748_ = ~new_n2746_ & ~new_n2747_;
  assign new_n2749_ = \in3[53]  & new_n1792_;
  assign new_n2750_ = \in2[53]  & ~new_n1792_;
  assign new_n2751_ = ~new_n2749_ & ~new_n2750_;
  assign new_n2752_ = new_n2748_ & ~new_n2751_;
  assign new_n2753_ = \in3[52]  & new_n1792_;
  assign new_n2754_ = \in2[52]  & ~new_n1792_;
  assign new_n2755_ = ~new_n2753_ & ~new_n2754_;
  assign new_n2756_ = \in1[52]  & new_n1787_;
  assign new_n2757_ = \in0[52]  & ~new_n1787_;
  assign new_n2758_ = ~new_n2756_ & ~new_n2757_;
  assign new_n2759_ = ~new_n2755_ & new_n2758_;
  assign new_n2760_ = ~new_n2752_ & ~new_n2759_;
  assign new_n2761_ = new_n2745_ & new_n2760_;
  assign new_n2762_ = \in1[49]  & new_n1787_;
  assign new_n2763_ = \in0[49]  & ~new_n1787_;
  assign new_n2764_ = ~new_n2762_ & ~new_n2763_;
  assign new_n2765_ = \in3[49]  & new_n1792_;
  assign new_n2766_ = \in2[49]  & ~new_n1792_;
  assign new_n2767_ = ~new_n2765_ & ~new_n2766_;
  assign new_n2768_ = new_n2764_ & ~new_n2767_;
  assign new_n2769_ = \in1[51]  & new_n1787_;
  assign new_n2770_ = \in0[51]  & ~new_n1787_;
  assign new_n2771_ = ~new_n2769_ & ~new_n2770_;
  assign new_n2772_ = \in3[51]  & new_n1792_;
  assign new_n2773_ = \in2[51]  & ~new_n1792_;
  assign new_n2774_ = ~new_n2772_ & ~new_n2773_;
  assign new_n2775_ = new_n2771_ & ~new_n2774_;
  assign new_n2776_ = \in3[50]  & new_n1792_;
  assign new_n2777_ = \in2[50]  & ~new_n1792_;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = \in1[50]  & new_n1787_;
  assign new_n2780_ = \in0[50]  & ~new_n1787_;
  assign new_n2781_ = ~new_n2779_ & ~new_n2780_;
  assign new_n2782_ = ~new_n2778_ & new_n2781_;
  assign new_n2783_ = ~new_n2775_ & ~new_n2782_;
  assign new_n2784_ = ~new_n2768_ & new_n2783_;
  assign new_n2785_ = new_n2761_ & new_n2784_;
  assign new_n2786_ = ~new_n2730_ & new_n2785_;
  assign new_n2787_ = ~new_n2723_ & new_n2786_;
  assign new_n2788_ = ~new_n2733_ & new_n2736_;
  assign new_n2789_ = ~new_n2771_ & new_n2774_;
  assign new_n2790_ = ~new_n2775_ & new_n2778_;
  assign new_n2791_ = ~new_n2781_ & new_n2790_;
  assign new_n2792_ = new_n2726_ & ~new_n2729_;
  assign new_n2793_ = ~new_n2764_ & new_n2767_;
  assign new_n2794_ = ~new_n2792_ & ~new_n2793_;
  assign new_n2795_ = new_n2784_ & ~new_n2794_;
  assign new_n2796_ = ~new_n2791_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2789_ & new_n2796_;
  assign new_n2798_ = new_n2761_ & ~new_n2797_;
  assign new_n2799_ = new_n2755_ & ~new_n2758_;
  assign new_n2800_ = ~new_n2752_ & new_n2799_;
  assign new_n2801_ = ~new_n2748_ & new_n2751_;
  assign new_n2802_ = ~new_n2800_ & ~new_n2801_;
  assign new_n2803_ = new_n2740_ & ~new_n2743_;
  assign new_n2804_ = new_n2802_ & ~new_n2803_;
  assign new_n2805_ = new_n2745_ & ~new_n2804_;
  assign new_n2806_ = ~new_n2798_ & ~new_n2805_;
  assign new_n2807_ = ~new_n2788_ & new_n2806_;
  assign new_n2808_ = ~new_n2787_ & new_n2807_;
  assign new_n2809_ = new_n2215_ & ~new_n2218_;
  assign new_n2810_ = ~new_n2212_ & ~new_n2809_;
  assign new_n2811_ = new_n2189_ & new_n2810_;
  assign new_n2812_ = new_n2205_ & new_n2811_;
  assign new_n2813_ = ~new_n2808_ & new_n2812_;
  assign new_n2814_ = ~new_n2234_ & ~new_n2813_;
  assign new_n2815_ = ~new_n2232_ & new_n2814_;
  assign new_n2816_ = ~new_n2227_ & new_n2815_;
  assign new_n2817_ = ~new_n2164_ & new_n2816_;
  assign new_n2818_ = ~new_n2157_ & ~new_n2817_;
  assign new_n2819_ = ~new_n2150_ & new_n2818_;
  assign new_n2820_ = new_n2143_ & new_n2819_;
  assign new_n2821_ = ~new_n2131_ & new_n2134_;
  assign new_n2822_ = new_n2146_ & ~new_n2157_;
  assign new_n2823_ = ~new_n2149_ & new_n2822_;
  assign new_n2824_ = ~new_n2153_ & new_n2156_;
  assign new_n2825_ = ~new_n2823_ & ~new_n2824_;
  assign new_n2826_ = new_n2138_ & ~new_n2141_;
  assign new_n2827_ = new_n2825_ & ~new_n2826_;
  assign new_n2828_ = new_n2143_ & ~new_n2827_;
  assign new_n2829_ = ~new_n2821_ & ~new_n2828_;
  assign new_n2830_ = ~new_n2820_ & new_n2829_;
  assign new_n2831_ = new_n2118_ & ~new_n2121_;
  assign new_n2832_ = ~new_n2115_ & ~new_n2831_;
  assign new_n2833_ = new_n2108_ & new_n2832_;
  assign new_n2834_ = ~new_n2830_ & new_n2833_;
  assign new_n2835_ = ~new_n2128_ & ~new_n2834_;
  assign new_n2836_ = ~new_n2126_ & new_n2835_;
  assign new_n2837_ = ~new_n2099_ & new_n2836_;
  assign new_n2838_ = \in1[75]  & new_n1787_;
  assign new_n2839_ = \in0[75]  & ~new_n1787_;
  assign new_n2840_ = ~new_n2838_ & ~new_n2839_;
  assign new_n2841_ = \in3[75]  & new_n1792_;
  assign new_n2842_ = \in2[75]  & ~new_n1792_;
  assign new_n2843_ = ~new_n2841_ & ~new_n2842_;
  assign new_n2844_ = new_n2840_ & ~new_n2843_;
  assign new_n2845_ = \in3[74]  & new_n1792_;
  assign new_n2846_ = \in2[74]  & ~new_n1792_;
  assign new_n2847_ = ~new_n2845_ & ~new_n2846_;
  assign new_n2848_ = \in1[74]  & new_n1787_;
  assign new_n2849_ = \in0[74]  & ~new_n1787_;
  assign new_n2850_ = ~new_n2848_ & ~new_n2849_;
  assign new_n2851_ = ~new_n2847_ & new_n2850_;
  assign new_n2852_ = ~new_n2844_ & ~new_n2851_;
  assign new_n2853_ = \in1[73]  & new_n1787_;
  assign new_n2854_ = \in0[73]  & ~new_n1787_;
  assign new_n2855_ = ~new_n2853_ & ~new_n2854_;
  assign new_n2856_ = \in3[73]  & new_n1792_;
  assign new_n2857_ = \in2[73]  & ~new_n1792_;
  assign new_n2858_ = ~new_n2856_ & ~new_n2857_;
  assign new_n2859_ = new_n2855_ & ~new_n2858_;
  assign new_n2860_ = \in3[72]  & new_n1792_;
  assign new_n2861_ = \in2[72]  & ~new_n1792_;
  assign new_n2862_ = ~new_n2860_ & ~new_n2861_;
  assign new_n2863_ = \in1[72]  & new_n1787_;
  assign new_n2864_ = \in0[72]  & ~new_n1787_;
  assign new_n2865_ = ~new_n2863_ & ~new_n2864_;
  assign new_n2866_ = ~new_n2862_ & new_n2865_;
  assign new_n2867_ = ~new_n2859_ & ~new_n2866_;
  assign new_n2868_ = new_n2852_ & new_n2867_;
  assign new_n2869_ = ~new_n2837_ & new_n2868_;
  assign new_n2870_ = ~new_n2840_ & new_n2843_;
  assign new_n2871_ = new_n2862_ & ~new_n2865_;
  assign new_n2872_ = ~new_n2859_ & new_n2871_;
  assign new_n2873_ = ~new_n2855_ & new_n2858_;
  assign new_n2874_ = ~new_n2872_ & ~new_n2873_;
  assign new_n2875_ = new_n2847_ & ~new_n2850_;
  assign new_n2876_ = new_n2874_ & ~new_n2875_;
  assign new_n2877_ = new_n2852_ & ~new_n2876_;
  assign new_n2878_ = ~new_n2870_ & ~new_n2877_;
  assign new_n2879_ = ~new_n2869_ & new_n2878_;
  assign new_n2880_ = new_n2082_ & ~new_n2085_;
  assign new_n2881_ = ~new_n2079_ & ~new_n2880_;
  assign new_n2882_ = new_n2072_ & new_n2881_;
  assign new_n2883_ = ~new_n2879_ & new_n2882_;
  assign new_n2884_ = ~new_n2092_ & ~new_n2883_;
  assign new_n2885_ = ~new_n2090_ & new_n2884_;
  assign new_n2886_ = ~new_n2063_ & new_n2885_;
  assign new_n2887_ = ~new_n2056_ & ~new_n2886_;
  assign new_n2888_ = new_n2049_ & new_n2887_;
  assign new_n2889_ = ~new_n2034_ & new_n2888_;
  assign new_n2890_ = ~new_n2037_ & new_n2040_;
  assign new_n2891_ = new_n2030_ & ~new_n2056_;
  assign new_n2892_ = ~new_n2033_ & new_n2891_;
  assign new_n2893_ = ~new_n2052_ & new_n2055_;
  assign new_n2894_ = ~new_n2892_ & ~new_n2893_;
  assign new_n2895_ = new_n2044_ & ~new_n2047_;
  assign new_n2896_ = new_n2894_ & ~new_n2895_;
  assign new_n2897_ = new_n2049_ & ~new_n2896_;
  assign new_n2898_ = ~new_n2890_ & ~new_n2897_;
  assign new_n2899_ = ~new_n2889_ & new_n2898_;
  assign new_n2900_ = new_n2017_ & ~new_n2020_;
  assign new_n2901_ = ~new_n2014_ & ~new_n2900_;
  assign new_n2902_ = new_n2007_ & new_n2901_;
  assign new_n2903_ = ~new_n2899_ & new_n2902_;
  assign new_n2904_ = ~new_n2027_ & ~new_n2903_;
  assign new_n2905_ = ~new_n2025_ & new_n2904_;
  assign new_n2906_ = ~new_n1998_ & new_n2905_;
  assign new_n2907_ = \in1[91]  & new_n1787_;
  assign new_n2908_ = \in0[91]  & ~new_n1787_;
  assign new_n2909_ = ~new_n2907_ & ~new_n2908_;
  assign new_n2910_ = \in3[91]  & new_n1792_;
  assign new_n2911_ = \in2[91]  & ~new_n1792_;
  assign new_n2912_ = ~new_n2910_ & ~new_n2911_;
  assign new_n2913_ = new_n2909_ & ~new_n2912_;
  assign new_n2914_ = \in3[90]  & new_n1792_;
  assign new_n2915_ = \in2[90]  & ~new_n1792_;
  assign new_n2916_ = ~new_n2914_ & ~new_n2915_;
  assign new_n2917_ = \in1[90]  & new_n1787_;
  assign new_n2918_ = \in0[90]  & ~new_n1787_;
  assign new_n2919_ = ~new_n2917_ & ~new_n2918_;
  assign new_n2920_ = ~new_n2916_ & new_n2919_;
  assign new_n2921_ = ~new_n2913_ & ~new_n2920_;
  assign new_n2922_ = \in1[89]  & new_n1787_;
  assign new_n2923_ = \in0[89]  & ~new_n1787_;
  assign new_n2924_ = ~new_n2922_ & ~new_n2923_;
  assign new_n2925_ = \in3[89]  & new_n1792_;
  assign new_n2926_ = \in2[89]  & ~new_n1792_;
  assign new_n2927_ = ~new_n2925_ & ~new_n2926_;
  assign new_n2928_ = new_n2924_ & ~new_n2927_;
  assign new_n2929_ = \in3[88]  & new_n1792_;
  assign new_n2930_ = \in2[88]  & ~new_n1792_;
  assign new_n2931_ = ~new_n2929_ & ~new_n2930_;
  assign new_n2932_ = \in1[88]  & new_n1787_;
  assign new_n2933_ = \in0[88]  & ~new_n1787_;
  assign new_n2934_ = ~new_n2932_ & ~new_n2933_;
  assign new_n2935_ = ~new_n2931_ & new_n2934_;
  assign new_n2936_ = ~new_n2928_ & ~new_n2935_;
  assign new_n2937_ = new_n2921_ & new_n2936_;
  assign new_n2938_ = ~new_n2906_ & new_n2937_;
  assign new_n2939_ = ~new_n2909_ & new_n2912_;
  assign new_n2940_ = new_n2931_ & ~new_n2934_;
  assign new_n2941_ = ~new_n2928_ & new_n2940_;
  assign new_n2942_ = ~new_n2924_ & new_n2927_;
  assign new_n2943_ = ~new_n2941_ & ~new_n2942_;
  assign new_n2944_ = new_n2916_ & ~new_n2919_;
  assign new_n2945_ = new_n2943_ & ~new_n2944_;
  assign new_n2946_ = new_n2921_ & ~new_n2945_;
  assign new_n2947_ = ~new_n2939_ & ~new_n2946_;
  assign new_n2948_ = ~new_n2938_ & new_n2947_;
  assign new_n2949_ = new_n1981_ & ~new_n1984_;
  assign new_n2950_ = ~new_n1978_ & ~new_n2949_;
  assign new_n2951_ = new_n1971_ & new_n2950_;
  assign new_n2952_ = ~new_n2948_ & new_n2951_;
  assign new_n2953_ = ~new_n1991_ & ~new_n2952_;
  assign new_n2954_ = ~new_n1989_ & new_n2953_;
  assign new_n2955_ = ~new_n1962_ & new_n2954_;
  assign new_n2956_ = ~new_n1955_ & ~new_n2955_;
  assign new_n2957_ = new_n1948_ & new_n2956_;
  assign new_n2958_ = ~new_n1933_ & new_n2957_;
  assign new_n2959_ = ~new_n1936_ & new_n1939_;
  assign new_n2960_ = new_n1929_ & ~new_n1955_;
  assign new_n2961_ = ~new_n1932_ & new_n2960_;
  assign new_n2962_ = ~new_n1951_ & new_n1954_;
  assign new_n2963_ = ~new_n2961_ & ~new_n2962_;
  assign new_n2964_ = new_n1943_ & ~new_n1946_;
  assign new_n2965_ = new_n2963_ & ~new_n2964_;
  assign new_n2966_ = new_n1948_ & ~new_n2965_;
  assign new_n2967_ = ~new_n2959_ & ~new_n2966_;
  assign new_n2968_ = ~new_n2958_ & new_n2967_;
  assign new_n2969_ = new_n1916_ & ~new_n1919_;
  assign new_n2970_ = ~new_n1913_ & ~new_n2969_;
  assign new_n2971_ = new_n1906_ & new_n2970_;
  assign new_n2972_ = ~new_n2968_ & new_n2971_;
  assign new_n2973_ = ~new_n1926_ & ~new_n2972_;
  assign new_n2974_ = ~new_n1924_ & new_n2973_;
  assign new_n2975_ = ~new_n1897_ & new_n2974_;
  assign new_n2976_ = \in1[107]  & new_n1787_;
  assign new_n2977_ = \in0[107]  & ~new_n1787_;
  assign new_n2978_ = ~new_n2976_ & ~new_n2977_;
  assign new_n2979_ = \in3[107]  & new_n1792_;
  assign new_n2980_ = \in2[107]  & ~new_n1792_;
  assign new_n2981_ = ~new_n2979_ & ~new_n2980_;
  assign new_n2982_ = new_n2978_ & ~new_n2981_;
  assign new_n2983_ = \in3[106]  & new_n1792_;
  assign new_n2984_ = \in2[106]  & ~new_n1792_;
  assign new_n2985_ = ~new_n2983_ & ~new_n2984_;
  assign new_n2986_ = \in1[106]  & new_n1787_;
  assign new_n2987_ = \in0[106]  & ~new_n1787_;
  assign new_n2988_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2989_ = ~new_n2985_ & new_n2988_;
  assign new_n2990_ = ~new_n2982_ & ~new_n2989_;
  assign new_n2991_ = \in1[105]  & new_n1787_;
  assign new_n2992_ = \in0[105]  & ~new_n1787_;
  assign new_n2993_ = ~new_n2991_ & ~new_n2992_;
  assign new_n2994_ = \in3[105]  & new_n1792_;
  assign new_n2995_ = \in2[105]  & ~new_n1792_;
  assign new_n2996_ = ~new_n2994_ & ~new_n2995_;
  assign new_n2997_ = new_n2993_ & ~new_n2996_;
  assign new_n2998_ = \in3[104]  & new_n1792_;
  assign new_n2999_ = \in2[104]  & ~new_n1792_;
  assign new_n3000_ = ~new_n2998_ & ~new_n2999_;
  assign new_n3001_ = \in1[104]  & new_n1787_;
  assign new_n3002_ = \in0[104]  & ~new_n1787_;
  assign new_n3003_ = ~new_n3001_ & ~new_n3002_;
  assign new_n3004_ = ~new_n3000_ & new_n3003_;
  assign new_n3005_ = ~new_n2997_ & ~new_n3004_;
  assign new_n3006_ = new_n2990_ & new_n3005_;
  assign new_n3007_ = ~new_n2975_ & new_n3006_;
  assign new_n3008_ = ~new_n2978_ & new_n2981_;
  assign new_n3009_ = new_n3000_ & ~new_n3003_;
  assign new_n3010_ = ~new_n2997_ & new_n3009_;
  assign new_n3011_ = ~new_n2993_ & new_n2996_;
  assign new_n3012_ = ~new_n3010_ & ~new_n3011_;
  assign new_n3013_ = new_n2985_ & ~new_n2988_;
  assign new_n3014_ = new_n3012_ & ~new_n3013_;
  assign new_n3015_ = new_n2990_ & ~new_n3014_;
  assign new_n3016_ = ~new_n3008_ & ~new_n3015_;
  assign new_n3017_ = ~new_n3007_ & new_n3016_;
  assign new_n3018_ = new_n1880_ & ~new_n1883_;
  assign new_n3019_ = ~new_n1877_ & ~new_n3018_;
  assign new_n3020_ = new_n1870_ & new_n3019_;
  assign new_n3021_ = ~new_n3017_ & new_n3020_;
  assign new_n3022_ = ~new_n1890_ & ~new_n3021_;
  assign new_n3023_ = ~new_n1888_ & new_n3022_;
  assign new_n3024_ = ~new_n1861_ & new_n3023_;
  assign new_n3025_ = ~new_n1854_ & ~new_n3024_;
  assign new_n3026_ = new_n1847_ & new_n3025_;
  assign new_n3027_ = ~new_n1832_ & new_n3026_;
  assign new_n3028_ = ~new_n1835_ & new_n1838_;
  assign new_n3029_ = new_n1828_ & ~new_n1854_;
  assign new_n3030_ = ~new_n1831_ & new_n3029_;
  assign new_n3031_ = ~new_n1850_ & new_n1853_;
  assign new_n3032_ = ~new_n3030_ & ~new_n3031_;
  assign new_n3033_ = new_n1842_ & ~new_n1845_;
  assign new_n3034_ = new_n3032_ & ~new_n3033_;
  assign new_n3035_ = new_n1847_ & ~new_n3034_;
  assign new_n3036_ = ~new_n3028_ & ~new_n3035_;
  assign new_n3037_ = ~new_n3027_ & new_n3036_;
  assign new_n3038_ = new_n1808_ & ~new_n1818_;
  assign new_n3039_ = ~new_n1815_ & ~new_n3038_;
  assign new_n3040_ = new_n1805_ & new_n3039_;
  assign new_n3041_ = ~new_n3037_ & new_n3040_;
  assign new_n3042_ = ~new_n1825_ & ~new_n3041_;
  assign new_n3043_ = ~new_n1823_ & new_n3042_;
  assign new_n3044_ = ~new_n1796_ & new_n3043_;
  assign new_n3045_ = \in1[123]  & new_n1787_;
  assign new_n3046_ = \in0[123]  & ~new_n1787_;
  assign new_n3047_ = ~new_n3045_ & ~new_n3046_;
  assign new_n3048_ = \in3[123]  & new_n1792_;
  assign new_n3049_ = \in2[123]  & ~new_n1792_;
  assign new_n3050_ = ~new_n3048_ & ~new_n3049_;
  assign new_n3051_ = new_n3047_ & ~new_n3050_;
  assign new_n3052_ = \in3[122]  & new_n1792_;
  assign new_n3053_ = \in2[122]  & ~new_n1792_;
  assign new_n3054_ = ~new_n3052_ & ~new_n3053_;
  assign new_n3055_ = \in1[122]  & new_n1787_;
  assign new_n3056_ = \in0[122]  & ~new_n1787_;
  assign new_n3057_ = ~new_n3055_ & ~new_n3056_;
  assign new_n3058_ = ~new_n3054_ & new_n3057_;
  assign new_n3059_ = ~new_n3051_ & ~new_n3058_;
  assign new_n3060_ = \in1[121]  & new_n1787_;
  assign new_n3061_ = \in0[121]  & ~new_n1787_;
  assign new_n3062_ = ~new_n3060_ & ~new_n3061_;
  assign new_n3063_ = \in3[121]  & new_n1792_;
  assign new_n3064_ = \in2[121]  & ~new_n1792_;
  assign new_n3065_ = ~new_n3063_ & ~new_n3064_;
  assign new_n3066_ = new_n3062_ & ~new_n3065_;
  assign new_n3067_ = \in3[120]  & new_n1792_;
  assign new_n3068_ = \in2[120]  & ~new_n1792_;
  assign new_n3069_ = ~new_n3067_ & ~new_n3068_;
  assign new_n3070_ = \in1[120]  & new_n1787_;
  assign new_n3071_ = \in0[120]  & ~new_n1787_;
  assign new_n3072_ = ~new_n3070_ & ~new_n3071_;
  assign new_n3073_ = ~new_n3069_ & new_n3072_;
  assign new_n3074_ = ~new_n3066_ & ~new_n3073_;
  assign new_n3075_ = new_n3059_ & new_n3074_;
  assign new_n3076_ = ~new_n3044_ & new_n3075_;
  assign new_n3077_ = ~new_n3047_ & new_n3050_;
  assign new_n3078_ = ~new_n3066_ & new_n3069_;
  assign new_n3079_ = ~new_n3072_ & new_n3078_;
  assign new_n3080_ = ~new_n3062_ & new_n3065_;
  assign new_n3081_ = ~new_n3079_ & ~new_n3080_;
  assign new_n3082_ = new_n3054_ & ~new_n3057_;
  assign new_n3083_ = new_n3081_ & ~new_n3082_;
  assign new_n3084_ = new_n3059_ & ~new_n3083_;
  assign new_n3085_ = ~new_n3077_ & ~new_n3084_;
  assign new_n3086_ = ~new_n3076_ & new_n3085_;
  assign new_n3087_ = \in1[124]  & new_n1787_;
  assign new_n3088_ = \in0[124]  & ~new_n1787_;
  assign new_n3089_ = ~new_n3087_ & ~new_n3088_;
  assign new_n3090_ = \in3[124]  & new_n1792_;
  assign new_n3091_ = \in2[124]  & ~new_n1792_;
  assign new_n3092_ = ~new_n3090_ & ~new_n3091_;
  assign new_n3093_ = new_n3089_ & ~new_n3092_;
  assign new_n3094_ = ~new_n1213_ & new_n1784_;
  assign new_n3095_ = \in1[126]  & new_n1787_;
  assign new_n3096_ = \in0[126]  & ~new_n1787_;
  assign new_n3097_ = ~new_n3095_ & ~new_n3096_;
  assign new_n3098_ = \in3[126]  & new_n1792_;
  assign new_n3099_ = \in2[126]  & ~new_n1792_;
  assign new_n3100_ = ~new_n3098_ & ~new_n3099_;
  assign new_n3101_ = new_n3097_ & ~new_n3100_;
  assign new_n3102_ = \in1[125]  & new_n1787_;
  assign new_n3103_ = \in0[125]  & ~new_n1787_;
  assign new_n3104_ = ~new_n3102_ & ~new_n3103_;
  assign new_n3105_ = \in3[125]  & new_n1792_;
  assign new_n3106_ = \in2[125]  & ~new_n1792_;
  assign new_n3107_ = ~new_n3105_ & ~new_n3106_;
  assign new_n3108_ = new_n3104_ & ~new_n3107_;
  assign new_n3109_ = ~new_n3101_ & ~new_n3108_;
  assign new_n3110_ = ~new_n3094_ & new_n3109_;
  assign new_n3111_ = ~new_n3093_ & new_n3110_;
  assign new_n3112_ = ~new_n3086_ & new_n3111_;
  assign new_n3113_ = ~new_n3089_ & new_n3092_;
  assign new_n3114_ = ~new_n3104_ & new_n3107_;
  assign new_n3115_ = ~new_n3113_ & ~new_n3114_;
  assign new_n3116_ = new_n3109_ & ~new_n3115_;
  assign new_n3117_ = ~new_n3097_ & new_n3100_;
  assign new_n3118_ = ~new_n3116_ & ~new_n3117_;
  assign new_n3119_ = ~new_n3094_ & ~new_n3118_;
  assign new_n3120_ = ~new_n3112_ & ~new_n3119_;
  assign \address[1]  = ~new_n1785_ & new_n3120_;
  assign new_n3122_ = ~new_n2503_ & \address[1] ;
  assign new_n3123_ = ~new_n2500_ & ~\address[1] ;
  assign \result[0]  = new_n3122_ | new_n3123_;
  assign new_n3125_ = ~new_n2497_ & \address[1] ;
  assign new_n3126_ = ~new_n2508_ & ~\address[1] ;
  assign \result[1]  = new_n3125_ | new_n3126_;
  assign new_n3128_ = ~new_n2515_ & \address[1] ;
  assign new_n3129_ = ~new_n2512_ & ~\address[1] ;
  assign \result[2]  = new_n3128_ | new_n3129_;
  assign new_n3131_ = ~new_n2493_ & \address[1] ;
  assign new_n3132_ = ~new_n2490_ & ~\address[1] ;
  assign \result[3]  = new_n3131_ | new_n3132_;
  assign new_n3134_ = ~new_n2484_ & \address[1] ;
  assign new_n3135_ = ~new_n2487_ & ~\address[1] ;
  assign \result[4]  = new_n3134_ | new_n3135_;
  assign new_n3137_ = ~new_n2478_ & \address[1] ;
  assign new_n3138_ = ~new_n2481_ & ~\address[1] ;
  assign \result[5]  = new_n3137_ | new_n3138_;
  assign new_n3140_ = ~new_n2472_ & \address[1] ;
  assign new_n3141_ = ~new_n2475_ & ~\address[1] ;
  assign \result[6]  = new_n3140_ | new_n3141_;
  assign new_n3143_ = ~new_n2468_ & \address[1] ;
  assign new_n3144_ = ~new_n2465_ & ~\address[1] ;
  assign \result[7]  = new_n3143_ | new_n3144_;
  assign new_n3146_ = ~new_n2462_ & \address[1] ;
  assign new_n3147_ = ~new_n2542_ & ~\address[1] ;
  assign \result[8]  = new_n3146_ | new_n3147_;
  assign new_n3149_ = ~new_n2459_ & \address[1] ;
  assign new_n3150_ = ~new_n2549_ & ~\address[1] ;
  assign \result[9]  = new_n3149_ | new_n3150_;
  assign new_n3152_ = ~new_n2455_ & \address[1] ;
  assign new_n3153_ = ~new_n2452_ & ~\address[1] ;
  assign \result[10]  = new_n3152_ | new_n3153_;
  assign new_n3155_ = ~new_n2448_ & \address[1] ;
  assign new_n3156_ = ~new_n2445_ & ~\address[1] ;
  assign \result[11]  = new_n3155_ | new_n3156_;
  assign new_n3158_ = ~new_n2441_ & \address[1] ;
  assign new_n3159_ = ~new_n2438_ & ~\address[1] ;
  assign \result[12]  = new_n3158_ | new_n3159_;
  assign new_n3161_ = ~new_n2434_ & \address[1] ;
  assign new_n3162_ = ~new_n2431_ & ~\address[1] ;
  assign \result[13]  = new_n3161_ | new_n3162_;
  assign new_n3164_ = ~new_n2427_ & \address[1] ;
  assign new_n3165_ = ~new_n2424_ & ~\address[1] ;
  assign \result[14]  = new_n3164_ | new_n3165_;
  assign new_n3167_ = ~new_n2420_ & \address[1] ;
  assign new_n3168_ = ~new_n2417_ & ~\address[1] ;
  assign \result[15]  = new_n3167_ | new_n3168_;
  assign new_n3170_ = ~new_n2414_ & \address[1] ;
  assign new_n3171_ = ~new_n2574_ & ~\address[1] ;
  assign \result[16]  = new_n3170_ | new_n3171_;
  assign new_n3173_ = ~new_n2411_ & \address[1] ;
  assign new_n3174_ = ~new_n2581_ & ~\address[1] ;
  assign \result[17]  = new_n3173_ | new_n3174_;
  assign new_n3176_ = ~new_n2407_ & \address[1] ;
  assign new_n3177_ = ~new_n2404_ & ~\address[1] ;
  assign \result[18]  = new_n3176_ | new_n3177_;
  assign new_n3179_ = ~new_n2400_ & \address[1] ;
  assign new_n3180_ = ~new_n2397_ & ~\address[1] ;
  assign \result[19]  = new_n3179_ | new_n3180_;
  assign new_n3182_ = ~new_n2393_ & \address[1] ;
  assign new_n3183_ = ~new_n2390_ & ~\address[1] ;
  assign \result[20]  = new_n3182_ | new_n3183_;
  assign new_n3185_ = ~new_n2386_ & \address[1] ;
  assign new_n3186_ = ~new_n2383_ & ~\address[1] ;
  assign \result[21]  = new_n3185_ | new_n3186_;
  assign new_n3188_ = ~new_n2379_ & \address[1] ;
  assign new_n3189_ = ~new_n2376_ & ~\address[1] ;
  assign \result[22]  = new_n3188_ | new_n3189_;
  assign new_n3191_ = ~new_n2372_ & \address[1] ;
  assign new_n3192_ = ~new_n2369_ & ~\address[1] ;
  assign \result[23]  = new_n3191_ | new_n3192_;
  assign new_n3194_ = ~new_n2366_ & \address[1] ;
  assign new_n3195_ = ~new_n2606_ & ~\address[1] ;
  assign \result[24]  = new_n3194_ | new_n3195_;
  assign new_n3197_ = ~new_n2363_ & \address[1] ;
  assign new_n3198_ = ~new_n2613_ & ~\address[1] ;
  assign \result[25]  = new_n3197_ | new_n3198_;
  assign new_n3200_ = ~new_n2359_ & \address[1] ;
  assign new_n3201_ = ~new_n2356_ & ~\address[1] ;
  assign \result[26]  = new_n3200_ | new_n3201_;
  assign new_n3203_ = ~new_n2352_ & \address[1] ;
  assign new_n3204_ = ~new_n2349_ & ~\address[1] ;
  assign \result[27]  = new_n3203_ | new_n3204_;
  assign new_n3206_ = ~new_n2345_ & \address[1] ;
  assign new_n3207_ = ~new_n2342_ & ~\address[1] ;
  assign \result[28]  = new_n3206_ | new_n3207_;
  assign new_n3209_ = ~new_n2338_ & \address[1] ;
  assign new_n3210_ = ~new_n2335_ & ~\address[1] ;
  assign \result[29]  = new_n3209_ | new_n3210_;
  assign new_n3212_ = ~new_n2331_ & \address[1] ;
  assign new_n3213_ = ~new_n2328_ & ~\address[1] ;
  assign \result[30]  = new_n3212_ | new_n3213_;
  assign new_n3215_ = ~new_n2324_ & \address[1] ;
  assign new_n3216_ = ~new_n2321_ & ~\address[1] ;
  assign \result[31]  = new_n3215_ | new_n3216_;
  assign new_n3218_ = ~new_n2314_ & \address[1] ;
  assign new_n3219_ = ~new_n2317_ & ~\address[1] ;
  assign \result[32]  = new_n3218_ | new_n3219_;
  assign new_n3221_ = ~new_n2672_ & \address[1] ;
  assign new_n3222_ = ~new_n2669_ & ~\address[1] ;
  assign \result[33]  = new_n3221_ | new_n3222_;
  assign new_n3224_ = ~new_n2683_ & \address[1] ;
  assign new_n3225_ = ~new_n2686_ & ~\address[1] ;
  assign \result[34]  = new_n3224_ | new_n3225_;
  assign new_n3227_ = ~new_n2679_ & \address[1] ;
  assign new_n3228_ = ~new_n2676_ & ~\address[1] ;
  assign \result[35]  = new_n3227_ | new_n3228_;
  assign new_n3230_ = ~new_n2656_ & \address[1] ;
  assign new_n3231_ = ~new_n2653_ & ~\address[1] ;
  assign \result[36]  = new_n3230_ | new_n3231_;
  assign new_n3233_ = ~new_n2663_ & \address[1] ;
  assign new_n3234_ = ~new_n2660_ & ~\address[1] ;
  assign \result[37]  = new_n3233_ | new_n3234_;
  assign new_n3236_ = ~new_n2645_ & \address[1] ;
  assign new_n3237_ = ~new_n2648_ & ~\address[1] ;
  assign \result[38]  = new_n3236_ | new_n3237_;
  assign new_n3239_ = ~new_n2641_ & \address[1] ;
  assign new_n3240_ = ~new_n2638_ & ~\address[1] ;
  assign \result[39]  = new_n3239_ | new_n3240_;
  assign new_n3242_ = ~new_n2295_ & \address[1] ;
  assign new_n3243_ = ~new_n2292_ & ~\address[1] ;
  assign \result[40]  = new_n3242_ | new_n3243_;
  assign new_n3245_ = ~new_n2288_ & \address[1] ;
  assign new_n3246_ = ~new_n2285_ & ~\address[1] ;
  assign \result[41]  = new_n3245_ | new_n3246_;
  assign new_n3248_ = ~new_n2280_ & \address[1] ;
  assign new_n3249_ = ~new_n2277_ & ~\address[1] ;
  assign \result[42]  = new_n3248_ | new_n3249_;
  assign new_n3251_ = ~new_n2272_ & \address[1] ;
  assign new_n3252_ = ~new_n2269_ & ~\address[1] ;
  assign \result[43]  = new_n3251_ | new_n3252_;
  assign new_n3254_ = ~new_n2256_ & \address[1] ;
  assign new_n3255_ = ~new_n2253_ & ~\address[1] ;
  assign \result[44]  = new_n3254_ | new_n3255_;
  assign new_n3257_ = ~new_n2263_ & \address[1] ;
  assign new_n3258_ = ~new_n2260_ & ~\address[1] ;
  assign \result[45]  = new_n3257_ | new_n3258_;
  assign new_n3260_ = ~new_n2245_ & \address[1] ;
  assign new_n3261_ = ~new_n2248_ & ~\address[1] ;
  assign \result[46]  = new_n3260_ | new_n3261_;
  assign new_n3263_ = ~new_n2240_ & \address[1] ;
  assign new_n3264_ = ~new_n2237_ & ~\address[1] ;
  assign \result[47]  = new_n3263_ | new_n3264_;
  assign new_n3266_ = ~new_n2726_ & \address[1] ;
  assign new_n3267_ = ~new_n2729_ & ~\address[1] ;
  assign \result[48]  = new_n3266_ | new_n3267_;
  assign new_n3269_ = ~new_n2767_ & \address[1] ;
  assign new_n3270_ = ~new_n2764_ & ~\address[1] ;
  assign \result[49]  = new_n3269_ | new_n3270_;
  assign new_n3272_ = ~new_n2778_ & \address[1] ;
  assign new_n3273_ = ~new_n2781_ & ~\address[1] ;
  assign \result[50]  = new_n3272_ | new_n3273_;
  assign new_n3275_ = ~new_n2774_ & \address[1] ;
  assign new_n3276_ = ~new_n2771_ & ~\address[1] ;
  assign \result[51]  = new_n3275_ | new_n3276_;
  assign new_n3278_ = ~new_n2755_ & \address[1] ;
  assign new_n3279_ = ~new_n2758_ & ~\address[1] ;
  assign \result[52]  = new_n3278_ | new_n3279_;
  assign new_n3281_ = ~new_n2751_ & \address[1] ;
  assign new_n3282_ = ~new_n2748_ & ~\address[1] ;
  assign \result[53]  = new_n3281_ | new_n3282_;
  assign new_n3284_ = ~new_n2740_ & \address[1] ;
  assign new_n3285_ = ~new_n2743_ & ~\address[1] ;
  assign \result[54]  = new_n3284_ | new_n3285_;
  assign new_n3287_ = ~new_n2736_ & \address[1] ;
  assign new_n3288_ = ~new_n2733_ & ~\address[1] ;
  assign \result[55]  = new_n3287_ | new_n3288_;
  assign new_n3290_ = ~new_n2218_ & \address[1] ;
  assign new_n3291_ = ~new_n2215_ & ~\address[1] ;
  assign \result[56]  = new_n3290_ | new_n3291_;
  assign new_n3293_ = ~new_n2211_ & \address[1] ;
  assign new_n3294_ = ~new_n2208_ & ~\address[1] ;
  assign \result[57]  = new_n3293_ | new_n3294_;
  assign new_n3296_ = ~new_n2203_ & \address[1] ;
  assign new_n3297_ = ~new_n2200_ & ~\address[1] ;
  assign \result[58]  = new_n3296_ | new_n3297_;
  assign new_n3299_ = ~new_n2195_ & \address[1] ;
  assign new_n3300_ = ~new_n2192_ & ~\address[1] ;
  assign \result[59]  = new_n3299_ | new_n3300_;
  assign new_n3302_ = ~new_n2179_ & \address[1] ;
  assign new_n3303_ = ~new_n2176_ & ~\address[1] ;
  assign \result[60]  = new_n3302_ | new_n3303_;
  assign new_n3305_ = ~new_n2186_ & \address[1] ;
  assign new_n3306_ = ~new_n2183_ & ~\address[1] ;
  assign \result[61]  = new_n3305_ | new_n3306_;
  assign new_n3308_ = ~new_n2168_ & \address[1] ;
  assign new_n3309_ = ~new_n2171_ & ~\address[1] ;
  assign \result[62]  = new_n3308_ | new_n3309_;
  assign new_n3311_ = ~new_n2163_ & \address[1] ;
  assign new_n3312_ = ~new_n2160_ & ~\address[1] ;
  assign \result[63]  = new_n3311_ | new_n3312_;
  assign new_n3314_ = ~new_n2146_ & \address[1] ;
  assign new_n3315_ = ~new_n2149_ & ~\address[1] ;
  assign \result[64]  = new_n3314_ | new_n3315_;
  assign new_n3317_ = ~new_n2156_ & \address[1] ;
  assign new_n3318_ = ~new_n2153_ & ~\address[1] ;
  assign \result[65]  = new_n3317_ | new_n3318_;
  assign new_n3320_ = ~new_n2138_ & \address[1] ;
  assign new_n3321_ = ~new_n2141_ & ~\address[1] ;
  assign \result[66]  = new_n3320_ | new_n3321_;
  assign new_n3323_ = ~new_n2134_ & \address[1] ;
  assign new_n3324_ = ~new_n2131_ & ~\address[1] ;
  assign \result[67]  = new_n3323_ | new_n3324_;
  assign new_n3326_ = ~new_n2121_ & \address[1] ;
  assign new_n3327_ = ~new_n2118_ & ~\address[1] ;
  assign \result[68]  = new_n3326_ | new_n3327_;
  assign new_n3329_ = ~new_n2114_ & \address[1] ;
  assign new_n3330_ = ~new_n2111_ & ~\address[1] ;
  assign \result[69]  = new_n3329_ | new_n3330_;
  assign new_n3332_ = ~new_n2103_ & \address[1] ;
  assign new_n3333_ = ~new_n2106_ & ~\address[1] ;
  assign \result[70]  = new_n3332_ | new_n3333_;
  assign new_n3335_ = ~new_n2098_ & \address[1] ;
  assign new_n3336_ = ~new_n2095_ & ~\address[1] ;
  assign \result[71]  = new_n3335_ | new_n3336_;
  assign new_n3338_ = ~new_n2862_ & \address[1] ;
  assign new_n3339_ = ~new_n2865_ & ~\address[1] ;
  assign \result[72]  = new_n3338_ | new_n3339_;
  assign new_n3341_ = ~new_n2858_ & \address[1] ;
  assign new_n3342_ = ~new_n2855_ & ~\address[1] ;
  assign \result[73]  = new_n3341_ | new_n3342_;
  assign new_n3344_ = ~new_n2847_ & \address[1] ;
  assign new_n3345_ = ~new_n2850_ & ~\address[1] ;
  assign \result[74]  = new_n3344_ | new_n3345_;
  assign new_n3347_ = ~new_n2843_ & \address[1] ;
  assign new_n3348_ = ~new_n2840_ & ~\address[1] ;
  assign \result[75]  = new_n3347_ | new_n3348_;
  assign new_n3350_ = ~new_n2085_ & \address[1] ;
  assign new_n3351_ = ~new_n2082_ & ~\address[1] ;
  assign \result[76]  = new_n3350_ | new_n3351_;
  assign new_n3353_ = ~new_n2078_ & \address[1] ;
  assign new_n3354_ = ~new_n2075_ & ~\address[1] ;
  assign \result[77]  = new_n3353_ | new_n3354_;
  assign new_n3356_ = ~new_n2067_ & \address[1] ;
  assign new_n3357_ = ~new_n2070_ & ~\address[1] ;
  assign \result[78]  = new_n3356_ | new_n3357_;
  assign new_n3359_ = ~new_n2062_ & \address[1] ;
  assign new_n3360_ = ~new_n2059_ & ~\address[1] ;
  assign \result[79]  = new_n3359_ | new_n3360_;
  assign new_n3362_ = ~new_n2030_ & \address[1] ;
  assign new_n3363_ = ~new_n2033_ & ~\address[1] ;
  assign \result[80]  = new_n3362_ | new_n3363_;
  assign new_n3365_ = ~new_n2055_ & \address[1] ;
  assign new_n3366_ = ~new_n2052_ & ~\address[1] ;
  assign \result[81]  = new_n3365_ | new_n3366_;
  assign new_n3368_ = ~new_n2044_ & \address[1] ;
  assign new_n3369_ = ~new_n2047_ & ~\address[1] ;
  assign \result[82]  = new_n3368_ | new_n3369_;
  assign new_n3371_ = ~new_n2040_ & \address[1] ;
  assign new_n3372_ = ~new_n2037_ & ~\address[1] ;
  assign \result[83]  = new_n3371_ | new_n3372_;
  assign new_n3374_ = ~new_n2020_ & \address[1] ;
  assign new_n3375_ = ~new_n2017_ & ~\address[1] ;
  assign \result[84]  = new_n3374_ | new_n3375_;
  assign new_n3377_ = ~new_n2013_ & \address[1] ;
  assign new_n3378_ = ~new_n2010_ & ~\address[1] ;
  assign \result[85]  = new_n3377_ | new_n3378_;
  assign new_n3380_ = ~new_n2002_ & \address[1] ;
  assign new_n3381_ = ~new_n2005_ & ~\address[1] ;
  assign \result[86]  = new_n3380_ | new_n3381_;
  assign new_n3383_ = ~new_n1997_ & \address[1] ;
  assign new_n3384_ = ~new_n1994_ & ~\address[1] ;
  assign \result[87]  = new_n3383_ | new_n3384_;
  assign new_n3386_ = ~new_n2931_ & \address[1] ;
  assign new_n3387_ = ~new_n2934_ & ~\address[1] ;
  assign \result[88]  = new_n3386_ | new_n3387_;
  assign new_n3389_ = ~new_n2927_ & \address[1] ;
  assign new_n3390_ = ~new_n2924_ & ~\address[1] ;
  assign \result[89]  = new_n3389_ | new_n3390_;
  assign new_n3392_ = ~new_n2916_ & \address[1] ;
  assign new_n3393_ = ~new_n2919_ & ~\address[1] ;
  assign \result[90]  = new_n3392_ | new_n3393_;
  assign new_n3395_ = ~new_n2912_ & \address[1] ;
  assign new_n3396_ = ~new_n2909_ & ~\address[1] ;
  assign \result[91]  = new_n3395_ | new_n3396_;
  assign new_n3398_ = ~new_n1984_ & \address[1] ;
  assign new_n3399_ = ~new_n1981_ & ~\address[1] ;
  assign \result[92]  = new_n3398_ | new_n3399_;
  assign new_n3401_ = ~new_n1977_ & \address[1] ;
  assign new_n3402_ = ~new_n1974_ & ~\address[1] ;
  assign \result[93]  = new_n3401_ | new_n3402_;
  assign new_n3404_ = ~new_n1966_ & \address[1] ;
  assign new_n3405_ = ~new_n1969_ & ~\address[1] ;
  assign \result[94]  = new_n3404_ | new_n3405_;
  assign new_n3407_ = ~new_n1961_ & \address[1] ;
  assign new_n3408_ = ~new_n1958_ & ~\address[1] ;
  assign \result[95]  = new_n3407_ | new_n3408_;
  assign new_n3410_ = ~new_n1929_ & \address[1] ;
  assign new_n3411_ = ~new_n1932_ & ~\address[1] ;
  assign \result[96]  = new_n3410_ | new_n3411_;
  assign new_n3413_ = ~new_n1954_ & \address[1] ;
  assign new_n3414_ = ~new_n1951_ & ~\address[1] ;
  assign \result[97]  = new_n3413_ | new_n3414_;
  assign new_n3416_ = ~new_n1943_ & \address[1] ;
  assign new_n3417_ = ~new_n1946_ & ~\address[1] ;
  assign \result[98]  = new_n3416_ | new_n3417_;
  assign new_n3419_ = ~new_n1939_ & \address[1] ;
  assign new_n3420_ = ~new_n1936_ & ~\address[1] ;
  assign \result[99]  = new_n3419_ | new_n3420_;
  assign new_n3422_ = ~new_n1919_ & \address[1] ;
  assign new_n3423_ = ~new_n1916_ & ~\address[1] ;
  assign \result[100]  = new_n3422_ | new_n3423_;
  assign new_n3425_ = ~new_n1912_ & \address[1] ;
  assign new_n3426_ = ~new_n1909_ & ~\address[1] ;
  assign \result[101]  = new_n3425_ | new_n3426_;
  assign new_n3428_ = ~new_n1901_ & \address[1] ;
  assign new_n3429_ = ~new_n1904_ & ~\address[1] ;
  assign \result[102]  = new_n3428_ | new_n3429_;
  assign new_n3431_ = ~new_n1896_ & \address[1] ;
  assign new_n3432_ = ~new_n1893_ & ~\address[1] ;
  assign \result[103]  = new_n3431_ | new_n3432_;
  assign new_n3434_ = ~new_n3000_ & \address[1] ;
  assign new_n3435_ = ~new_n3003_ & ~\address[1] ;
  assign \result[104]  = new_n3434_ | new_n3435_;
  assign new_n3437_ = ~new_n2996_ & \address[1] ;
  assign new_n3438_ = ~new_n2993_ & ~\address[1] ;
  assign \result[105]  = new_n3437_ | new_n3438_;
  assign new_n3440_ = ~new_n2985_ & \address[1] ;
  assign new_n3441_ = ~new_n2988_ & ~\address[1] ;
  assign \result[106]  = new_n3440_ | new_n3441_;
  assign new_n3443_ = ~new_n2981_ & \address[1] ;
  assign new_n3444_ = ~new_n2978_ & ~\address[1] ;
  assign \result[107]  = new_n3443_ | new_n3444_;
  assign new_n3446_ = ~new_n1883_ & \address[1] ;
  assign new_n3447_ = ~new_n1880_ & ~\address[1] ;
  assign \result[108]  = new_n3446_ | new_n3447_;
  assign new_n3449_ = ~new_n1876_ & \address[1] ;
  assign new_n3450_ = ~new_n1873_ & ~\address[1] ;
  assign \result[109]  = new_n3449_ | new_n3450_;
  assign new_n3452_ = ~new_n1865_ & \address[1] ;
  assign new_n3453_ = ~new_n1868_ & ~\address[1] ;
  assign \result[110]  = new_n3452_ | new_n3453_;
  assign new_n3455_ = ~new_n1860_ & \address[1] ;
  assign new_n3456_ = ~new_n1857_ & ~\address[1] ;
  assign \result[111]  = new_n3455_ | new_n3456_;
  assign new_n3458_ = ~new_n1828_ & \address[1] ;
  assign new_n3459_ = ~new_n1831_ & ~\address[1] ;
  assign \result[112]  = new_n3458_ | new_n3459_;
  assign new_n3461_ = ~new_n1853_ & \address[1] ;
  assign new_n3462_ = ~new_n1850_ & ~\address[1] ;
  assign \result[113]  = new_n3461_ | new_n3462_;
  assign new_n3464_ = ~new_n1842_ & \address[1] ;
  assign new_n3465_ = ~new_n1845_ & ~\address[1] ;
  assign \result[114]  = new_n3464_ | new_n3465_;
  assign new_n3467_ = ~new_n1838_ & \address[1] ;
  assign new_n3468_ = ~new_n1835_ & ~\address[1] ;
  assign \result[115]  = new_n3467_ | new_n3468_;
  assign new_n3470_ = ~new_n1818_ & \address[1] ;
  assign new_n3471_ = ~new_n1808_ & ~\address[1] ;
  assign \result[116]  = new_n3470_ | new_n3471_;
  assign new_n3473_ = ~new_n1814_ & \address[1] ;
  assign new_n3474_ = ~new_n1811_ & ~\address[1] ;
  assign \result[117]  = new_n3473_ | new_n3474_;
  assign new_n3476_ = ~new_n1800_ & \address[1] ;
  assign new_n3477_ = ~new_n1803_ & ~\address[1] ;
  assign \result[118]  = new_n3476_ | new_n3477_;
  assign new_n3479_ = ~new_n1795_ & \address[1] ;
  assign new_n3480_ = ~new_n1790_ & ~\address[1] ;
  assign \result[119]  = new_n3479_ | new_n3480_;
  assign new_n3482_ = ~new_n3069_ & \address[1] ;
  assign new_n3483_ = ~new_n3072_ & ~\address[1] ;
  assign \result[120]  = new_n3482_ | new_n3483_;
  assign new_n3485_ = ~new_n3065_ & \address[1] ;
  assign new_n3486_ = ~new_n3062_ & ~\address[1] ;
  assign \result[121]  = new_n3485_ | new_n3486_;
  assign new_n3488_ = ~new_n3054_ & \address[1] ;
  assign new_n3489_ = ~new_n3057_ & ~\address[1] ;
  assign \result[122]  = new_n3488_ | new_n3489_;
  assign new_n3491_ = ~new_n3050_ & \address[1] ;
  assign new_n3492_ = ~new_n3047_ & ~\address[1] ;
  assign \result[123]  = new_n3491_ | new_n3492_;
  assign new_n3494_ = ~new_n3092_ & \address[1] ;
  assign new_n3495_ = ~new_n3089_ & ~\address[1] ;
  assign \result[124]  = new_n3494_ | new_n3495_;
  assign new_n3497_ = ~new_n3107_ & \address[1] ;
  assign new_n3498_ = ~new_n3104_ & ~\address[1] ;
  assign \result[125]  = new_n3497_ | new_n3498_;
  assign new_n3500_ = ~new_n3100_ & \address[1] ;
  assign new_n3501_ = ~new_n3097_ & ~\address[1] ;
  assign \result[126]  = new_n3500_ | new_n3501_;
  assign new_n3503_ = ~new_n1213_ & new_n3120_;
  assign \result[127]  = new_n1784_ & ~new_n3503_;
  assign new_n3505_ = new_n1792_ & \address[1] ;
  assign new_n3506_ = new_n1787_ & ~\address[1] ;
  assign \address[0]  = new_n3505_ | new_n3506_;
endmodule


