module top ( 
    p0, q1, r2, s3, a, p1, q0, r3, s2, b, p2, q3, r0, s1, c, p3, q2, r1,
    s0, d, t0, u1, v2, w3, e, t1, u0, v3, w2, f, t2, u3, v0, w1, g, t3, u2,
    v1, w0, h, x0, y1, z2, i, x1, y0, z3, j, x2, y3, z0, k, x3, y2, z1, l,
    m, n, o, a1, b2, c3, d4, p, a0, b3, c2, e4, q, a3, b0, c1, r, a2, b1,
    c0, s, d0, e1, f2, g3, t, a4, d1, e0, f3, g2, u, b4, d2, e3, f0, g1, v,
    c4, d3, e2, f1, g0, w, h0, i1, j2, k3, x, h1, i0, j3, k2, y, h2, i3,
    j0, k1, z, h3, i2, j1, k0, l0, m1, n2, o3, l1, m0, n3, o2, l2, m3, n0,
    o1, l3, m2, n1, o0,
    t4, u5, v6, w7, t5, u4, v7, w6, t6, u7, v4, w5, t7, u6, v5, w4, p4, q5,
    r6, s7, p5, q4, r7, s6, p6, q7, r4, s5, p7, q6, r5, s4, x4, y5, z6, x5,
    y4, z7, x6, y7, z4, x7, y6, z5, e5, f6, g7, h8, d5, f7, g6, d6, e7, f4,
    g5, d7, e6, f5, g4, a5, b6, c7, b7, c6, a7, c5, a6, b5, l4, m5, n6, o7,
    a8, l5, m4, n7, o6, b8, l6, m7, n4, o5, c8, l7, m6, n5, o4, d8, h4, i5,
    j6, k7, e8, h5, i4, j7, k6, f8, h6, i7, j4, k5, g8, h7, i6, j5, k4  );
  input  p0, q1, r2, s3, a, p1, q0, r3, s2, b, p2, q3, r0, s1, c, p3, q2,
    r1, s0, d, t0, u1, v2, w3, e, t1, u0, v3, w2, f, t2, u3, v0, w1, g, t3,
    u2, v1, w0, h, x0, y1, z2, i, x1, y0, z3, j, x2, y3, z0, k, x3, y2, z1,
    l, m, n, o, a1, b2, c3, d4, p, a0, b3, c2, e4, q, a3, b0, c1, r, a2,
    b1, c0, s, d0, e1, f2, g3, t, a4, d1, e0, f3, g2, u, b4, d2, e3, f0,
    g1, v, c4, d3, e2, f1, g0, w, h0, i1, j2, k3, x, h1, i0, j3, k2, y, h2,
    i3, j0, k1, z, h3, i2, j1, k0, l0, m1, n2, o3, l1, m0, n3, o2, l2, m3,
    n0, o1, l3, m2, n1, o0;
  output t4, u5, v6, w7, t5, u4, v7, w6, t6, u7, v4, w5, t7, u6, v5, w4, p4,
    q5, r6, s7, p5, q4, r7, s6, p6, q7, r4, s5, p7, q6, r5, s4, x4, y5, z6,
    x5, y4, z7, x6, y7, z4, x7, y6, z5, e5, f6, g7, h8, d5, f7, g6, d6, e7,
    f4, g5, d7, e6, f5, g4, a5, b6, c7, b7, c6, a7, c5, a6, b5, l4, m5, n6,
    o7, a8, l5, m4, n7, o6, b8, l6, m7, n4, o5, c8, l7, m6, n5, o4, d8, h4,
    i5, j6, k7, e8, h5, i4, j7, k6, f8, h6, i7, j4, k5, g8, h7, i6, j5, k4;
  wire new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n342_, new_n343_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n529_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1055_,
    new_n1056_, new_n1057_, new_n1059_, new_n1061_, new_n1062_, new_n1063_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1076_, new_n1077_,
    new_n1079_, new_n1080_, new_n1081_, new_n1083_, new_n1085_, new_n1086_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1096_, new_n1097_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1122_, new_n1123_, new_n1125_, new_n1126_,
    new_n1127_, new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1199_,
    new_n1200_, new_n1202_, new_n1204_, new_n1205_, new_n1207_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1222_,
    new_n1223_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1237_,
    new_n1238_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1257_, new_n1260_,
    new_n1261_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1275_,
    new_n1276_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1284_, new_n1285_, new_n1287_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1302_, new_n1304_, new_n1305_, new_n1306_,
    new_n1308_, new_n1309_, new_n1311_, new_n1312_, new_n1313_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1327_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1346_;
  assign new_n243_ = d & f;
  assign new_n244_ = e & new_n243_;
  assign new_n245_ = a & new_n244_;
  assign new_n246_ = a & ~s1;
  assign new_n247_ = a & ~n;
  assign new_n248_ = a & r1;
  assign new_n249_ = ~new_n245_ & ~new_n246_;
  assign new_n250_ = ~new_n247_ & ~new_n248_;
  assign new_n251_ = new_n249_ & new_n250_;
  assign new_n252_ = o2 & ~new_n251_;
  assign new_n253_ = n2 & ~new_n251_;
  assign new_n254_ = ~new_n252_ & ~new_n253_;
  assign new_n255_ = z1 & o2;
  assign new_n256_ = r1 & new_n255_;
  assign new_n257_ = ~s1 & new_n256_;
  assign new_n258_ = ~p1 & new_n257_;
  assign new_n259_ = h2 & new_n258_;
  assign new_n260_ = ~g2 & ~h2;
  assign new_n261_ = f2 & new_n260_;
  assign new_n262_ = ~g2 & h2;
  assign new_n263_ = ~f2 & new_n262_;
  assign new_n264_ = ~new_n261_ & ~new_n263_;
  assign new_n265_ = o2 & l2;
  assign new_n266_ = ~r1 & new_n265_;
  assign new_n267_ = s1 & new_n266_;
  assign new_n268_ = ~p1 & new_n267_;
  assign new_n269_ = ~new_n264_ & new_n268_;
  assign new_n270_ = f2 & new_n269_;
  assign new_n271_ = f2 & new_n258_;
  assign new_n272_ = ~r1 & new_n255_;
  assign new_n273_ = s1 & new_n272_;
  assign new_n274_ = ~p1 & new_n273_;
  assign new_n275_ = h2 & new_n274_;
  assign new_n276_ = f2 & new_n274_;
  assign new_n277_ = r1 & new_n265_;
  assign new_n278_ = ~s1 & new_n277_;
  assign new_n279_ = ~p1 & new_n278_;
  assign new_n280_ = ~new_n264_ & new_n279_;
  assign new_n281_ = h2 & new_n280_;
  assign new_n282_ = f2 & new_n280_;
  assign new_n283_ = h2 & new_n269_;
  assign new_n284_ = ~new_n259_ & ~new_n270_;
  assign new_n285_ = ~new_n271_ & ~new_n275_;
  assign new_n286_ = new_n284_ & new_n285_;
  assign new_n287_ = ~new_n282_ & ~new_n283_;
  assign new_n288_ = ~new_n276_ & ~new_n281_;
  assign new_n289_ = new_n287_ & new_n288_;
  assign new_n290_ = new_n286_ & new_n289_;
  assign new_n291_ = s0 & u2;
  assign new_n292_ = u & new_n291_;
  assign new_n293_ = ~s0 & u2;
  assign new_n294_ = h0 & new_n293_;
  assign new_n295_ = y1 & x1;
  assign new_n296_ = m2 & new_n295_;
  assign new_n297_ = x2 & ~new_n296_;
  assign new_n298_ = u3 & ~i;
  assign new_n299_ = u3 & new_n291_;
  assign new_n300_ = ~u & new_n299_;
  assign new_n301_ = ~h & new_n300_;
  assign new_n302_ = ~j & d0;
  assign new_n303_ = ~l & ~d0;
  assign new_n304_ = x2 & ~h0;
  assign new_n305_ = ~d0 & new_n304_;
  assign new_n306_ = ~w2 & new_n305_;
  assign new_n307_ = ~m & new_n306_;
  assign new_n308_ = u2 & new_n307_;
  assign new_n309_ = ~s0 & new_n308_;
  assign new_n310_ = x2 & ~u;
  assign new_n311_ = ~d0 & new_n310_;
  assign new_n312_ = ~w2 & new_n311_;
  assign new_n313_ = ~m & new_n312_;
  assign new_n314_ = u2 & new_n313_;
  assign new_n315_ = s0 & new_n314_;
  assign new_n316_ = d0 & new_n304_;
  assign new_n317_ = ~w2 & new_n316_;
  assign new_n318_ = ~k & new_n317_;
  assign new_n319_ = u2 & new_n318_;
  assign new_n320_ = ~s0 & new_n319_;
  assign new_n321_ = u3 & new_n293_;
  assign new_n322_ = ~h0 & new_n321_;
  assign new_n323_ = ~h & new_n322_;
  assign new_n324_ = d0 & new_n310_;
  assign new_n325_ = ~w2 & new_n324_;
  assign new_n326_ = ~k & new_n325_;
  assign new_n327_ = u2 & new_n326_;
  assign new_n328_ = s0 & new_n327_;
  assign new_n329_ = g & ~new_n303_;
  assign new_n330_ = ~new_n298_ & ~new_n301_;
  assign new_n331_ = ~new_n302_ & new_n330_;
  assign new_n332_ = new_n329_ & new_n331_;
  assign new_n333_ = ~new_n323_ & ~new_n328_;
  assign new_n334_ = ~new_n309_ & ~new_n315_;
  assign new_n335_ = ~new_n320_ & new_n334_;
  assign new_n336_ = new_n333_ & new_n335_;
  assign new_n337_ = new_n332_ & new_n336_;
  assign new_n338_ = w2 & new_n337_;
  assign new_n339_ = w2 & ~x2;
  assign new_n340_ = ~new_n297_ & ~new_n338_;
  assign d8 = new_n339_ | ~new_n340_;
  assign new_n342_ = c2 & d8;
  assign new_n343_ = ~new_n292_ & ~new_n294_;
  assign j4 = new_n342_ | ~new_n343_;
  assign new_n345_ = ~new_n290_ & ~j4;
  assign new_n346_ = a & f0;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = r2 & new_n347_;
  assign new_n349_ = s0 & ~b2;
  assign new_n350_ = s0 & d8;
  assign new_n351_ = s1 & s0;
  assign new_n352_ = ~new_n349_ & ~new_n350_;
  assign new_n353_ = ~new_n351_ & new_n352_;
  assign new_n354_ = ~z3 & ~new_n353_;
  assign new_n355_ = ~d8 & new_n354_;
  assign new_n356_ = u2 & new_n355_;
  assign new_n357_ = n1 & d8;
  assign new_n358_ = ~s1 & n1;
  assign new_n359_ = ~b2 & n1;
  assign new_n360_ = r1 & n1;
  assign new_n361_ = ~new_n357_ & ~new_n358_;
  assign new_n362_ = ~new_n359_ & ~new_n360_;
  assign new_n363_ = new_n361_ & new_n362_;
  assign new_n364_ = ~z3 & ~new_n363_;
  assign new_n365_ = ~d8 & new_n364_;
  assign new_n366_ = v2 & new_n365_;
  assign new_n367_ = new_n296_ & new_n337_;
  assign new_n368_ = w2 & new_n367_;
  assign new_n369_ = ~z3 & ~y3;
  assign new_n370_ = ~d8 & new_n369_;
  assign new_n371_ = v2 & new_n370_;
  assign new_n372_ = ~s & ~l3;
  assign new_n373_ = ~d8 & new_n372_;
  assign new_n374_ = ~z3 & new_n373_;
  assign new_n375_ = u2 & new_n374_;
  assign new_n376_ = b2 & ~d8;
  assign new_n377_ = v1 & new_n376_;
  assign new_n378_ = i3 & ~new_n377_;
  assign new_n379_ = m3 & new_n378_;
  assign new_n380_ = ~h3 & new_n379_;
  assign new_n381_ = f3 & ~new_n377_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~i3 & ~new_n377_;
  assign new_n384_ = m3 & new_n383_;
  assign new_n385_ = h3 & new_n384_;
  assign new_n386_ = e3 & ~new_n377_;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_ = new_n382_ & new_n387_;
  assign new_n389_ = r1 & ~new_n290_;
  assign new_n390_ = ~new_n377_ & ~new_n388_;
  assign new_n391_ = ~new_n389_ & new_n390_;
  assign new_n392_ = g3 & new_n391_;
  assign new_n393_ = ~new_n388_ & new_n392_;
  assign new_n394_ = ~d8 & new_n393_;
  assign new_n395_ = ~new_n389_ & new_n394_;
  assign new_n396_ = y2 & new_n395_;
  assign new_n397_ = ~z3 & new_n396_;
  assign new_n398_ = ~new_n356_ & ~new_n366_;
  assign new_n399_ = ~new_n368_ & ~new_n371_;
  assign new_n400_ = new_n398_ & new_n399_;
  assign new_n401_ = ~new_n339_ & ~new_n375_;
  assign new_n402_ = ~new_n397_ & new_n401_;
  assign new_n403_ = new_n400_ & new_n402_;
  assign new_n404_ = ~new_n348_ & ~new_n403_;
  assign new_n405_ = ~n2 & ~new_n254_;
  assign new_n406_ = ~new_n404_ & new_n405_;
  assign new_n407_ = n2 & new_n254_;
  assign new_n408_ = ~new_n404_ & new_n407_;
  assign new_n409_ = s0 & u;
  assign new_n410_ = u2 & new_n409_;
  assign new_n411_ = ~t & new_n410_;
  assign new_n412_ = ~s0 & h0;
  assign new_n413_ = u2 & new_n412_;
  assign new_n414_ = ~g0 & new_n413_;
  assign new_n415_ = ~new_n411_ & ~new_n414_;
  assign i4 = d8 | ~new_n415_;
  assign h4 = v2 | d8;
  assign new_n418_ = i4 & ~h4;
  assign new_n419_ = new_n404_ & new_n418_;
  assign new_n420_ = y2 & ~new_n388_;
  assign new_n421_ = new_n404_ & new_n420_;
  assign new_n422_ = ~i4 & h4;
  assign new_n423_ = new_n404_ & new_n422_;
  assign new_n424_ = s0 & v;
  assign new_n425_ = ~i4 & new_n424_;
  assign new_n426_ = new_n404_ & new_n425_;
  assign new_n427_ = ~s0 & i0;
  assign new_n428_ = ~i4 & new_n427_;
  assign new_n429_ = new_n404_ & new_n428_;
  assign new_n430_ = ~new_n406_ & ~new_n408_;
  assign new_n431_ = ~new_n419_ & ~new_n421_;
  assign new_n432_ = new_n430_ & new_n431_;
  assign new_n433_ = ~new_n423_ & ~new_n426_;
  assign new_n434_ = ~new_n429_ & new_n433_;
  assign t4 = ~new_n432_ | ~new_n434_;
  assign new_n436_ = l2 & ~new_n264_;
  assign new_n437_ = u2 & ~new_n348_;
  assign new_n438_ = l0 & new_n437_;
  assign new_n439_ = ~s0 & l0;
  assign new_n440_ = ~t3 & ~o3;
  assign new_n441_ = ~n3 & new_n440_;
  assign new_n442_ = a2 & ~new_n441_;
  assign new_n443_ = l0 & ~new_n442_;
  assign new_n444_ = ~z1 & ~new_n443_;
  assign new_n445_ = ~new_n436_ & ~new_n438_;
  assign new_n446_ = ~new_n439_ & new_n445_;
  assign u5 = ~new_n444_ | ~new_n446_;
  assign v6 = ~y0 & ~z0;
  assign new_n449_ = ~z2 & ~a3;
  assign new_n450_ = k0 & ~new_n449_;
  assign new_n451_ = k0 & ~new_n442_;
  assign new_n452_ = h0 & k0;
  assign new_n453_ = ~new_n450_ & ~new_n451_;
  assign new_n454_ = ~l2 & ~new_n452_;
  assign t5 = ~new_n453_ | ~new_n454_;
  assign new_n456_ = o2 & new_n254_;
  assign new_n457_ = ~new_n404_ & new_n456_;
  assign new_n458_ = y2 & ~new_n382_;
  assign new_n459_ = ~new_n387_ & new_n458_;
  assign new_n460_ = new_n404_ & new_n459_;
  assign new_n461_ = n2 & o2;
  assign new_n462_ = ~new_n404_ & new_n461_;
  assign new_n463_ = ~o2 & new_n405_;
  assign new_n464_ = ~new_n404_ & new_n463_;
  assign new_n465_ = ~new_n457_ & ~new_n460_;
  assign new_n466_ = ~new_n419_ & new_n465_;
  assign new_n467_ = ~new_n423_ & ~new_n462_;
  assign new_n468_ = ~new_n464_ & new_n467_;
  assign u4 = ~new_n466_ | ~new_n468_;
  assign new_n470_ = ~p & ~q;
  assign new_n471_ = o & new_n470_;
  assign new_n472_ = l2 & new_n471_;
  assign new_n473_ = ~k2 & new_n472_;
  assign new_n474_ = ~x0 & ~z0;
  assign new_n475_ = y0 & new_n474_;
  assign new_n476_ = ~w0 & new_n475_;
  assign new_n477_ = x0 & ~z0;
  assign new_n478_ = ~y0 & new_n477_;
  assign new_n479_ = ~w0 & new_n478_;
  assign new_n480_ = w0 & z0;
  assign new_n481_ = ~new_n476_ & ~new_n479_;
  assign new_n482_ = ~new_n480_ & new_n481_;
  assign new_n483_ = u1 & ~z0;
  assign new_n484_ = ~x0 & new_n483_;
  assign new_n485_ = ~y0 & new_n484_;
  assign new_n486_ = ~w0 & new_n485_;
  assign new_n487_ = u1 & z0;
  assign new_n488_ = x0 & new_n487_;
  assign new_n489_ = ~y0 & new_n488_;
  assign new_n490_ = ~w0 & new_n489_;
  assign new_n491_ = y0 & new_n484_;
  assign new_n492_ = w0 & new_n491_;
  assign new_n493_ = y0 & new_n488_;
  assign new_n494_ = w0 & new_n493_;
  assign new_n495_ = ~new_n486_ & ~new_n490_;
  assign new_n496_ = ~new_n492_ & ~new_n494_;
  assign new_n497_ = new_n495_ & new_n496_;
  assign new_n498_ = new_n482_ & new_n497_;
  assign new_n499_ = j2 & new_n498_;
  assign t6 = new_n473_ | new_n499_;
  assign new_n501_ = n2 & new_n347_;
  assign new_n502_ = ~new_n403_ & new_n501_;
  assign new_n503_ = o2 & new_n347_;
  assign new_n504_ = r2 & new_n503_;
  assign new_n505_ = new_n347_ & ~new_n403_;
  assign new_n506_ = new_n251_ & new_n505_;
  assign new_n507_ = r2 & new_n501_;
  assign new_n508_ = new_n251_ & new_n347_;
  assign new_n509_ = r2 & new_n508_;
  assign new_n510_ = ~new_n403_ & new_n503_;
  assign new_n511_ = ~new_n502_ & ~new_n504_;
  assign new_n512_ = ~new_n506_ & new_n511_;
  assign new_n513_ = ~new_n507_ & ~new_n509_;
  assign new_n514_ = ~new_n510_ & new_n513_;
  assign v4 = ~new_n512_ | ~new_n514_;
  assign new_n516_ = j2 & ~new_n497_;
  assign new_n517_ = j2 & ~new_n482_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = l0 & new_n518_;
  assign new_n520_ = m0 & new_n519_;
  assign new_n521_ = k0 & new_n520_;
  assign new_n522_ = t0 & n3;
  assign new_n523_ = ~h0 & new_n522_;
  assign new_n524_ = new_n521_ & ~new_n523_;
  assign new_n525_ = new_n442_ & new_n524_;
  assign new_n526_ = j0 & new_n521_;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign w5 = n3 & ~new_n527_;
  assign new_n529_ = t0 & new_n497_;
  assign u6 = g0 & new_n529_;
  assign new_n531_ = h0 & ~l3;
  assign new_n532_ = t0 & new_n531_;
  assign new_n533_ = ~g0 & new_n532_;
  assign new_n534_ = ~q & l2;
  assign new_n535_ = ~o & new_n534_;
  assign new_n536_ = p & new_n535_;
  assign new_n537_ = ~new_n533_ & new_n536_;
  assign new_n538_ = h3 & new_n537_;
  assign new_n539_ = ~i3 & new_n537_;
  assign new_n540_ = ~y1 & m2;
  assign new_n541_ = ~w1 & new_n540_;
  assign new_n542_ = x1 & new_n541_;
  assign new_n543_ = ~new_n533_ & new_n542_;
  assign new_n544_ = p2 & l2;
  assign new_n545_ = p & new_n544_;
  assign new_n546_ = ~q & new_n545_;
  assign new_n547_ = ~new_n533_ & new_n546_;
  assign new_n548_ = m0 & ~new_n533_;
  assign new_n549_ = ~new_n547_ & ~new_n548_;
  assign new_n550_ = ~new_n538_ & ~new_n539_;
  assign new_n551_ = ~new_n543_ & new_n550_;
  assign v5 = ~new_n549_ | ~new_n551_;
  assign new_n553_ = ~b & ~new_n251_;
  assign new_n554_ = ~new_n404_ & new_n553_;
  assign new_n555_ = b & new_n251_;
  assign new_n556_ = ~new_n404_ & new_n555_;
  assign new_n557_ = d2 & new_n404_;
  assign new_n558_ = ~new_n554_ & ~new_n556_;
  assign w4 = new_n557_ | ~new_n558_;
  assign new_n560_ = z1 & ~f2;
  assign new_n561_ = ~t2 & new_n560_;
  assign new_n562_ = new_n348_ & new_n561_;
  assign new_n563_ = ~a & new_n562_;
  assign new_n564_ = z1 & ~g2;
  assign new_n565_ = t1 & new_n564_;
  assign new_n566_ = ~new_n403_ & new_n565_;
  assign new_n567_ = ~a & new_n566_;
  assign new_n568_ = ~new_n403_ & new_n561_;
  assign new_n569_ = ~a & new_n568_;
  assign new_n570_ = t1 & new_n560_;
  assign new_n571_ = new_n348_ & new_n570_;
  assign new_n572_ = ~a & new_n571_;
  assign new_n573_ = ~new_n403_ & new_n570_;
  assign new_n574_ = ~a & new_n573_;
  assign new_n575_ = ~t2 & new_n260_;
  assign new_n576_ = new_n348_ & new_n575_;
  assign new_n577_ = ~a & new_n576_;
  assign new_n578_ = l2 & new_n577_;
  assign new_n579_ = z1 & ~l2;
  assign new_n580_ = t1 & new_n579_;
  assign new_n581_ = ~new_n403_ & new_n580_;
  assign new_n582_ = ~a & new_n581_;
  assign new_n583_ = t1 & new_n260_;
  assign new_n584_ = new_n348_ & new_n583_;
  assign new_n585_ = ~a & new_n584_;
  assign new_n586_ = l2 & new_n585_;
  assign new_n587_ = ~t2 & new_n579_;
  assign new_n588_ = ~new_n403_ & new_n587_;
  assign new_n589_ = ~a & new_n588_;
  assign new_n590_ = new_n348_ & new_n580_;
  assign new_n591_ = ~a & new_n590_;
  assign new_n592_ = new_n348_ & new_n587_;
  assign new_n593_ = ~a & new_n592_;
  assign new_n594_ = ~f2 & ~g2;
  assign new_n595_ = ~t2 & new_n594_;
  assign new_n596_ = new_n348_ & new_n595_;
  assign new_n597_ = ~a & new_n596_;
  assign new_n598_ = l2 & new_n597_;
  assign new_n599_ = ~f2 & ~h2;
  assign new_n600_ = t1 & new_n599_;
  assign new_n601_ = ~new_n403_ & new_n600_;
  assign new_n602_ = ~a & new_n601_;
  assign new_n603_ = t1 & new_n594_;
  assign new_n604_ = new_n348_ & new_n603_;
  assign new_n605_ = ~a & new_n604_;
  assign new_n606_ = l2 & new_n605_;
  assign new_n607_ = ~t2 & new_n599_;
  assign new_n608_ = ~new_n403_ & new_n607_;
  assign new_n609_ = ~a & new_n608_;
  assign new_n610_ = ~new_n403_ & new_n575_;
  assign new_n611_ = ~a & new_n610_;
  assign new_n612_ = l2 & new_n611_;
  assign new_n613_ = new_n348_ & new_n600_;
  assign new_n614_ = ~a & new_n613_;
  assign new_n615_ = ~new_n403_ & new_n583_;
  assign new_n616_ = ~a & new_n615_;
  assign new_n617_ = l2 & new_n616_;
  assign new_n618_ = new_n348_ & new_n607_;
  assign new_n619_ = ~a & new_n618_;
  assign new_n620_ = ~new_n403_ & new_n595_;
  assign new_n621_ = ~a & new_n620_;
  assign new_n622_ = l2 & new_n621_;
  assign new_n623_ = z1 & ~h2;
  assign new_n624_ = t1 & new_n623_;
  assign new_n625_ = new_n348_ & new_n624_;
  assign new_n626_ = ~a & new_n625_;
  assign new_n627_ = ~new_n403_ & new_n603_;
  assign new_n628_ = ~a & new_n627_;
  assign new_n629_ = l2 & new_n628_;
  assign new_n630_ = ~t2 & new_n623_;
  assign new_n631_ = new_n348_ & new_n630_;
  assign new_n632_ = ~a & new_n631_;
  assign new_n633_ = ~new_n403_ & new_n630_;
  assign new_n634_ = ~a & new_n633_;
  assign new_n635_ = ~t2 & new_n564_;
  assign new_n636_ = new_n348_ & new_n635_;
  assign new_n637_ = ~a & new_n636_;
  assign new_n638_ = ~new_n403_ & new_n624_;
  assign new_n639_ = ~a & new_n638_;
  assign new_n640_ = ~new_n403_ & new_n635_;
  assign new_n641_ = ~a & new_n640_;
  assign new_n642_ = new_n348_ & new_n565_;
  assign new_n643_ = ~a & new_n642_;
  assign new_n644_ = ~new_n639_ & ~new_n641_;
  assign new_n645_ = ~new_n643_ & new_n644_;
  assign new_n646_ = ~new_n629_ & ~new_n632_;
  assign new_n647_ = ~new_n634_ & ~new_n637_;
  assign new_n648_ = new_n646_ & new_n647_;
  assign new_n649_ = new_n645_ & new_n648_;
  assign new_n650_ = ~new_n619_ & ~new_n622_;
  assign new_n651_ = ~new_n626_ & new_n650_;
  assign new_n652_ = ~new_n614_ & ~new_n617_;
  assign new_n653_ = ~new_n609_ & ~new_n612_;
  assign new_n654_ = new_n652_ & new_n653_;
  assign new_n655_ = new_n651_ & new_n654_;
  assign new_n656_ = new_n649_ & new_n655_;
  assign new_n657_ = ~new_n598_ & ~new_n602_;
  assign new_n658_ = ~new_n606_ & new_n657_;
  assign new_n659_ = ~new_n586_ & ~new_n589_;
  assign new_n660_ = ~new_n591_ & ~new_n593_;
  assign new_n661_ = new_n659_ & new_n660_;
  assign new_n662_ = new_n658_ & new_n661_;
  assign new_n663_ = ~new_n563_ & ~new_n567_;
  assign new_n664_ = ~new_n569_ & ~new_n572_;
  assign new_n665_ = new_n663_ & new_n664_;
  assign new_n666_ = ~new_n574_ & ~new_n578_;
  assign new_n667_ = ~new_n582_ & new_n666_;
  assign new_n668_ = new_n665_ & new_n667_;
  assign new_n669_ = new_n662_ & new_n668_;
  assign p4 = ~new_n656_ | ~new_n669_;
  assign new_n671_ = new_n442_ & ~new_n521_;
  assign new_n672_ = j0 & new_n523_;
  assign new_n673_ = ~i3 & h3;
  assign new_n674_ = i3 & ~h3;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = l2 & o0;
  assign new_n677_ = d3 & new_n676_;
  assign new_n678_ = new_n449_ & new_n677_;
  assign new_n679_ = z2 & new_n678_;
  assign new_n680_ = ~a3 & new_n678_;
  assign new_n681_ = ~d3 & new_n449_;
  assign new_n682_ = ~b3 & new_n681_;
  assign new_n683_ = ~c3 & new_n682_;
  assign new_n684_ = ~a3 & new_n683_;
  assign new_n685_ = ~new_n389_ & new_n449_;
  assign new_n686_ = ~c3 & new_n685_;
  assign new_n687_ = ~d3 & new_n686_;
  assign new_n688_ = ~b3 & new_n687_;
  assign new_n689_ = z2 & new_n683_;
  assign new_n690_ = o0 & new_n449_;
  assign new_n691_ = b3 & new_n690_;
  assign new_n692_ = ~c3 & new_n691_;
  assign new_n693_ = ~a3 & new_n692_;
  assign new_n694_ = l2 & new_n693_;
  assign new_n695_ = ~c3 & new_n690_;
  assign new_n696_ = ~new_n389_ & new_n695_;
  assign new_n697_ = b3 & new_n696_;
  assign new_n698_ = l2 & new_n697_;
  assign new_n699_ = ~new_n389_ & new_n676_;
  assign new_n700_ = new_n449_ & new_n699_;
  assign new_n701_ = d3 & new_n700_;
  assign new_n702_ = z2 & new_n692_;
  assign new_n703_ = l2 & new_n702_;
  assign new_n704_ = ~new_n688_ & ~new_n689_;
  assign new_n705_ = ~new_n679_ & ~new_n680_;
  assign new_n706_ = ~new_n684_ & new_n705_;
  assign new_n707_ = new_n704_ & new_n706_;
  assign new_n708_ = ~new_n701_ & ~new_n703_;
  assign new_n709_ = ~new_n694_ & ~new_n698_;
  assign new_n710_ = new_n708_ & new_n709_;
  assign new_n711_ = new_n707_ & new_n710_;
  assign new_n712_ = new_n685_ & new_n711_;
  assign new_n713_ = m3 & new_n712_;
  assign new_n714_ = i3 & new_n449_;
  assign new_n715_ = new_n711_ & new_n714_;
  assign new_n716_ = h3 & new_n715_;
  assign new_n717_ = ~new_n713_ & ~new_n716_;
  assign new_n718_ = ~new_n675_ & new_n717_;
  assign new_n719_ = t0 & ~new_n497_;
  assign new_n720_ = ~l2 & new_n719_;
  assign new_n721_ = g0 & new_n720_;
  assign new_n722_ = new_n442_ & new_n721_;
  assign new_n723_ = ~new_n471_ & ~new_n518_;
  assign new_n724_ = new_n482_ & ~new_n518_;
  assign new_n725_ = ~l2 & ~new_n518_;
  assign new_n726_ = new_n348_ & new_n442_;
  assign new_n727_ = t0 & new_n726_;
  assign new_n728_ = ~l3 & new_n727_;
  assign new_n729_ = t0 & new_n449_;
  assign new_n730_ = ~l3 & new_n729_;
  assign new_n731_ = new_n442_ & new_n730_;
  assign new_n732_ = ~h0 & new_n731_;
  assign new_n733_ = ~u2 & new_n442_;
  assign new_n734_ = t0 & new_n733_;
  assign new_n735_ = ~l3 & new_n734_;
  assign new_n736_ = ~s0 & d8;
  assign new_n737_ = ~h0 & new_n736_;
  assign new_n738_ = ~s0 & z3;
  assign new_n739_ = ~h0 & new_n738_;
  assign new_n740_ = ~u & new_n350_;
  assign new_n741_ = s0 & z3;
  assign new_n742_ = ~u & new_n741_;
  assign new_n743_ = ~new_n739_ & ~new_n740_;
  assign new_n744_ = ~new_n742_ & new_n743_;
  assign new_n745_ = ~new_n732_ & ~new_n735_;
  assign new_n746_ = ~new_n737_ & new_n745_;
  assign new_n747_ = new_n744_ & new_n746_;
  assign new_n748_ = ~new_n718_ & ~new_n722_;
  assign new_n749_ = ~new_n723_ & new_n748_;
  assign new_n750_ = ~new_n724_ & ~new_n725_;
  assign new_n751_ = ~new_n728_ & new_n750_;
  assign new_n752_ = new_n749_ & new_n751_;
  assign new_n753_ = new_n747_ & new_n752_;
  assign new_n754_ = new_n442_ & ~new_n753_;
  assign new_n755_ = j0 & ~new_n521_;
  assign new_n756_ = j0 & ~new_n753_;
  assign new_n757_ = new_n442_ & new_n523_;
  assign new_n758_ = ~new_n671_ & ~new_n672_;
  assign new_n759_ = ~new_n754_ & new_n758_;
  assign new_n760_ = ~new_n755_ & ~new_n756_;
  assign new_n761_ = ~new_n757_ & new_n760_;
  assign q5 = ~new_n759_ | ~new_n761_;
  assign new_n763_ = c3 & o0;
  assign new_n764_ = b3 & o0;
  assign new_n765_ = ~new_n763_ & ~new_n764_;
  assign new_n766_ = c3 & new_n711_;
  assign new_n767_ = new_n765_ & new_n766_;
  assign new_n768_ = b3 & new_n767_;
  assign new_n769_ = ~new_n389_ & new_n765_;
  assign new_n770_ = new_n711_ & new_n769_;
  assign new_n771_ = c3 & new_n770_;
  assign new_n772_ = a3 & ~new_n711_;
  assign new_n773_ = ~new_n768_ & ~new_n771_;
  assign r6 = new_n772_ | ~new_n773_;
  assign new_n775_ = g2 & ~h2;
  assign new_n776_ = g2 & l2;
  assign new_n777_ = f2 & ~h2;
  assign new_n778_ = f2 & l2;
  assign new_n779_ = ~h2 & ~l2;
  assign new_n780_ = ~new_n778_ & ~new_n779_;
  assign new_n781_ = ~new_n775_ & ~new_n776_;
  assign new_n782_ = ~new_n777_ & new_n781_;
  assign p5 = ~new_n780_ | ~new_n782_;
  assign new_n784_ = ~a & new_n599_;
  assign new_n785_ = ~t1 & new_n784_;
  assign new_n786_ = t2 & new_n785_;
  assign new_n787_ = t2 & a1;
  assign q4 = new_n786_ | new_n787_;
  assign new_n789_ = new_n296_ & ~new_n337_;
  assign new_n790_ = s1 & new_n789_;
  assign new_n791_ = ~r1 & new_n790_;
  assign new_n792_ = s1 & d4;
  assign new_n793_ = ~r1 & new_n792_;
  assign new_n794_ = s1 & d8;
  assign new_n795_ = ~r1 & new_n794_;
  assign new_n796_ = ~new_n791_ & ~new_n793_;
  assign r7 = new_n795_ | ~new_n796_;
  assign new_n798_ = ~o0 & new_n711_;
  assign new_n799_ = d3 & new_n798_;
  assign new_n800_ = c3 & ~new_n765_;
  assign s6 = new_n799_ | new_n800_;
  assign new_n802_ = i3 & ~new_n449_;
  assign new_n803_ = h3 & new_n802_;
  assign new_n804_ = ~new_n389_ & ~new_n711_;
  assign new_n805_ = ~new_n675_ & new_n804_;
  assign new_n806_ = m3 & new_n805_;
  assign new_n807_ = new_n711_ & new_n729_;
  assign new_n808_ = ~h0 & new_n807_;
  assign new_n809_ = ~new_n449_ & new_n808_;
  assign new_n810_ = i3 & ~new_n711_;
  assign new_n811_ = h3 & new_n810_;
  assign new_n812_ = ~new_n711_ & new_n808_;
  assign new_n813_ = ~new_n389_ & ~new_n449_;
  assign new_n814_ = ~new_n675_ & new_n813_;
  assign new_n815_ = m3 & new_n814_;
  assign new_n816_ = ~new_n803_ & ~new_n806_;
  assign new_n817_ = ~new_n809_ & new_n816_;
  assign new_n818_ = ~new_n811_ & ~new_n812_;
  assign new_n819_ = ~new_n815_ & new_n818_;
  assign new_n820_ = new_n817_ & new_n819_;
  assign new_n821_ = a3 & new_n711_;
  assign new_n822_ = new_n820_ & new_n821_;
  assign new_n823_ = z2 & new_n822_;
  assign new_n824_ = new_n711_ & new_n820_;
  assign new_n825_ = ~new_n389_ & new_n824_;
  assign new_n826_ = a3 & new_n825_;
  assign new_n827_ = new_n424_ & ~new_n820_;
  assign new_n828_ = ~u & new_n827_;
  assign new_n829_ = new_n427_ & ~new_n820_;
  assign new_n830_ = ~h0 & new_n829_;
  assign new_n831_ = ~new_n675_ & ~new_n820_;
  assign new_n832_ = ~s0 & new_n711_;
  assign new_n833_ = a3 & new_n832_;
  assign new_n834_ = ~new_n389_ & new_n833_;
  assign new_n835_ = h0 & new_n834_;
  assign new_n836_ = s0 & new_n711_;
  assign new_n837_ = a3 & new_n836_;
  assign new_n838_ = ~new_n389_ & new_n837_;
  assign new_n839_ = u & new_n838_;
  assign new_n840_ = z2 & new_n832_;
  assign new_n841_ = a3 & new_n840_;
  assign new_n842_ = h0 & new_n841_;
  assign new_n843_ = z2 & new_n836_;
  assign new_n844_ = a3 & new_n843_;
  assign new_n845_ = u & new_n844_;
  assign new_n846_ = ~s0 & ~new_n820_;
  assign new_n847_ = z2 & new_n846_;
  assign new_n848_ = a3 & new_n847_;
  assign new_n849_ = h0 & new_n848_;
  assign new_n850_ = ~s0 & ~new_n389_;
  assign new_n851_ = a3 & new_n850_;
  assign new_n852_ = ~new_n820_ & new_n851_;
  assign new_n853_ = h0 & new_n852_;
  assign new_n854_ = s0 & ~new_n820_;
  assign new_n855_ = z2 & new_n854_;
  assign new_n856_ = a3 & new_n855_;
  assign new_n857_ = u & new_n856_;
  assign new_n858_ = s0 & ~new_n389_;
  assign new_n859_ = a3 & new_n858_;
  assign new_n860_ = ~new_n820_ & new_n859_;
  assign new_n861_ = u & new_n860_;
  assign new_n862_ = ~new_n823_ & ~new_n826_;
  assign new_n863_ = ~new_n828_ & ~new_n830_;
  assign new_n864_ = new_n862_ & new_n863_;
  assign new_n865_ = ~new_n831_ & ~new_n835_;
  assign new_n866_ = ~new_n839_ & new_n865_;
  assign new_n867_ = new_n864_ & new_n866_;
  assign new_n868_ = ~new_n853_ & ~new_n857_;
  assign new_n869_ = ~new_n861_ & new_n868_;
  assign new_n870_ = ~new_n842_ & ~new_n845_;
  assign new_n871_ = ~new_n849_ & new_n870_;
  assign new_n872_ = new_n869_ & new_n871_;
  assign p6 = ~new_n867_ | ~new_n872_;
  assign new_n874_ = ~s1 & new_n789_;
  assign new_n875_ = ~s1 & d4;
  assign new_n876_ = ~s1 & d8;
  assign new_n877_ = ~new_n874_ & ~new_n875_;
  assign q7 = new_n876_ | ~new_n877_;
  assign new_n879_ = ~g1 & ~h1;
  assign new_n880_ = o0 & new_n879_;
  assign new_n881_ = ~f1 & new_n880_;
  assign new_n882_ = a & new_n881_;
  assign new_n883_ = g2 & new_n882_;
  assign new_n884_ = new_n264_ & new_n881_;
  assign new_n885_ = g2 & new_n884_;
  assign new_n886_ = h2 & new_n470_;
  assign new_n887_ = ~o & new_n886_;
  assign new_n888_ = ~l2 & new_n887_;
  assign new_n889_ = ~q1 & ~r1;
  assign new_n890_ = ~l2 & new_n889_;
  assign new_n891_ = ~h2 & new_n890_;
  assign new_n892_ = a & new_n891_;
  assign new_n893_ = ~s1 & new_n892_;
  assign new_n894_ = ~l2 & o0;
  assign new_n895_ = ~s1 & ~r1;
  assign new_n896_ = h2 & new_n895_;
  assign new_n897_ = ~q1 & new_n896_;
  assign new_n898_ = new_n264_ & new_n897_;
  assign new_n899_ = ~p & new_n898_;
  assign new_n900_ = ~q & new_n899_;
  assign new_n901_ = ~g2 & new_n900_;
  assign new_n902_ = ~o & new_n901_;
  assign new_n903_ = h2 & new_n879_;
  assign new_n904_ = ~f1 & new_n903_;
  assign new_n905_ = new_n264_ & new_n904_;
  assign new_n906_ = ~p & new_n905_;
  assign new_n907_ = ~q & new_n906_;
  assign new_n908_ = g2 & new_n907_;
  assign new_n909_ = ~o & new_n908_;
  assign new_n910_ = a & new_n897_;
  assign new_n911_ = ~p & new_n910_;
  assign new_n912_ = ~q & new_n911_;
  assign new_n913_ = ~g2 & new_n912_;
  assign new_n914_ = ~o & new_n913_;
  assign new_n915_ = a & new_n904_;
  assign new_n916_ = ~p & new_n915_;
  assign new_n917_ = ~q & new_n916_;
  assign new_n918_ = g2 & new_n917_;
  assign new_n919_ = ~o & new_n918_;
  assign new_n920_ = ~h2 & new_n895_;
  assign new_n921_ = ~q1 & new_n920_;
  assign new_n922_ = a & new_n921_;
  assign new_n923_ = ~g2 & new_n922_;
  assign new_n924_ = ~h2 & new_n879_;
  assign new_n925_ = ~f1 & new_n924_;
  assign new_n926_ = a & new_n925_;
  assign new_n927_ = ~s1 & new_n926_;
  assign new_n928_ = g2 & new_n927_;
  assign new_n929_ = ~q1 & new_n928_;
  assign new_n930_ = ~r1 & new_n929_;
  assign new_n931_ = o0 & new_n895_;
  assign new_n932_ = ~q1 & new_n931_;
  assign new_n933_ = a & new_n932_;
  assign new_n934_ = ~g2 & new_n933_;
  assign new_n935_ = new_n264_ & new_n932_;
  assign new_n936_ = ~g2 & new_n935_;
  assign new_n937_ = ~new_n883_ & ~new_n885_;
  assign new_n938_ = ~new_n888_ & ~new_n893_;
  assign new_n939_ = new_n937_ & new_n938_;
  assign new_n940_ = ~new_n894_ & ~new_n902_;
  assign new_n941_ = ~new_n909_ & new_n940_;
  assign new_n942_ = new_n939_ & new_n941_;
  assign new_n943_ = ~new_n930_ & ~new_n934_;
  assign new_n944_ = ~new_n936_ & new_n943_;
  assign new_n945_ = ~new_n914_ & ~new_n919_;
  assign new_n946_ = ~new_n923_ & new_n945_;
  assign new_n947_ = new_n944_ & new_n946_;
  assign r4 = ~new_n942_ | ~new_n947_;
  assign new_n949_ = ~o3 & new_n442_;
  assign s5 = new_n499_ | new_n949_;
  assign new_n951_ = a4 & ~d8;
  assign new_n952_ = ~new_n348_ & new_n951_;
  assign new_n953_ = ~new_n363_ & new_n952_;
  assign new_n954_ = a4 & new_n392_;
  assign new_n955_ = ~new_n348_ & new_n954_;
  assign new_n956_ = ~d8 & new_n955_;
  assign new_n957_ = ~new_n527_ & new_n952_;
  assign new_n958_ = e4 & i1;
  assign new_n959_ = new_n952_ & new_n958_;
  assign new_n960_ = ~v2 & new_n951_;
  assign new_n961_ = ~new_n363_ & new_n960_;
  assign new_n962_ = ~v2 & new_n353_;
  assign new_n963_ = ~d8 & new_n962_;
  assign new_n964_ = ~new_n392_ & new_n963_;
  assign new_n965_ = new_n958_ & new_n964_;
  assign new_n966_ = a4 & new_n965_;
  assign new_n967_ = s & new_n966_;
  assign new_n968_ = ~new_n527_ & new_n964_;
  assign new_n969_ = a4 & new_n968_;
  assign new_n970_ = l3 & new_n969_;
  assign new_n971_ = l3 & new_n966_;
  assign new_n972_ = y3 & ~new_n392_;
  assign new_n973_ = new_n363_ & new_n972_;
  assign new_n974_ = ~d8 & new_n973_;
  assign new_n975_ = ~new_n527_ & new_n974_;
  assign new_n976_ = s & new_n975_;
  assign new_n977_ = new_n353_ & new_n976_;
  assign new_n978_ = a4 & new_n977_;
  assign new_n979_ = y3 & new_n388_;
  assign new_n980_ = ~d8 & new_n979_;
  assign new_n981_ = new_n392_ & new_n980_;
  assign new_n982_ = new_n363_ & new_n981_;
  assign new_n983_ = a4 & new_n982_;
  assign new_n984_ = new_n958_ & new_n974_;
  assign new_n985_ = l3 & new_n984_;
  assign new_n986_ = new_n353_ & new_n985_;
  assign new_n987_ = a4 & new_n986_;
  assign new_n988_ = ~u2 & ~new_n392_;
  assign new_n989_ = new_n363_ & new_n988_;
  assign new_n990_ = ~d8 & new_n989_;
  assign new_n991_ = ~new_n527_ & new_n990_;
  assign new_n992_ = y3 & new_n991_;
  assign new_n993_ = a4 & new_n992_;
  assign new_n994_ = new_n958_ & new_n990_;
  assign new_n995_ = y3 & new_n994_;
  assign new_n996_ = a4 & new_n995_;
  assign new_n997_ = s & new_n969_;
  assign new_n998_ = l3 & new_n975_;
  assign new_n999_ = new_n353_ & new_n998_;
  assign new_n1000_ = a4 & new_n999_;
  assign new_n1001_ = y3 & ~y2;
  assign new_n1002_ = ~d8 & new_n1001_;
  assign new_n1003_ = new_n392_ & new_n1002_;
  assign new_n1004_ = new_n363_ & new_n1003_;
  assign new_n1005_ = a4 & new_n1004_;
  assign new_n1006_ = s & new_n984_;
  assign new_n1007_ = new_n353_ & new_n1006_;
  assign new_n1008_ = a4 & new_n1007_;
  assign new_n1009_ = y3 & new_n389_;
  assign new_n1010_ = ~d8 & new_n1009_;
  assign new_n1011_ = new_n392_ & new_n1010_;
  assign new_n1012_ = new_n363_ & new_n1011_;
  assign new_n1013_ = a4 & new_n1012_;
  assign new_n1014_ = ~v2 & ~u2;
  assign new_n1015_ = ~d8 & new_n1014_;
  assign new_n1016_ = ~new_n392_ & new_n1015_;
  assign new_n1017_ = new_n958_ & new_n1016_;
  assign new_n1018_ = a4 & new_n1017_;
  assign new_n1019_ = a4 & new_n388_;
  assign new_n1020_ = new_n392_ & new_n1019_;
  assign new_n1021_ = ~v2 & new_n1020_;
  assign new_n1022_ = ~d8 & new_n1021_;
  assign new_n1023_ = ~new_n527_ & new_n1016_;
  assign new_n1024_ = a4 & new_n1023_;
  assign new_n1025_ = ~y2 & a4;
  assign new_n1026_ = new_n392_ & new_n1025_;
  assign new_n1027_ = ~v2 & new_n1026_;
  assign new_n1028_ = ~d8 & new_n1027_;
  assign new_n1029_ = a4 & new_n389_;
  assign new_n1030_ = new_n392_ & new_n1029_;
  assign new_n1031_ = ~v2 & new_n1030_;
  assign new_n1032_ = ~d8 & new_n1031_;
  assign new_n1033_ = ~new_n1028_ & ~new_n1032_;
  assign new_n1034_ = ~new_n1018_ & ~new_n1022_;
  assign new_n1035_ = ~new_n1024_ & new_n1034_;
  assign new_n1036_ = new_n1033_ & new_n1035_;
  assign new_n1037_ = ~new_n1005_ & ~new_n1008_;
  assign new_n1038_ = ~new_n1013_ & new_n1037_;
  assign new_n1039_ = ~new_n996_ & ~new_n997_;
  assign new_n1040_ = ~new_n1000_ & new_n1039_;
  assign new_n1041_ = new_n1038_ & new_n1040_;
  assign new_n1042_ = new_n1036_ & new_n1041_;
  assign new_n1043_ = ~new_n983_ & ~new_n987_;
  assign new_n1044_ = ~new_n993_ & new_n1043_;
  assign new_n1045_ = ~new_n970_ & ~new_n971_;
  assign new_n1046_ = ~new_n978_ & new_n1045_;
  assign new_n1047_ = new_n1044_ & new_n1046_;
  assign new_n1048_ = ~new_n953_ & ~new_n956_;
  assign new_n1049_ = ~new_n957_ & new_n1048_;
  assign new_n1050_ = ~new_n959_ & ~new_n961_;
  assign new_n1051_ = ~new_n967_ & new_n1050_;
  assign new_n1052_ = new_n1049_ & new_n1051_;
  assign new_n1053_ = new_n1047_ & new_n1052_;
  assign p7 = ~new_n1042_ | ~new_n1053_;
  assign new_n1055_ = new_n711_ & new_n765_;
  assign new_n1056_ = b3 & new_n1055_;
  assign new_n1057_ = z2 & ~new_n711_;
  assign q6 = new_n1056_ | new_n1057_;
  assign new_n1059_ = ~new_n527_ & new_n753_;
  assign r5 = ~new_n533_ & new_n1059_;
  assign new_n1061_ = ~new_n290_ & j4;
  assign new_n1062_ = ~a & new_n1061_;
  assign new_n1063_ = ~a & f0;
  assign s4 = new_n1062_ | new_n1063_;
  assign new_n1065_ = b & ~new_n251_;
  assign new_n1066_ = ~c & new_n1065_;
  assign new_n1067_ = ~new_n404_ & new_n1066_;
  assign new_n1068_ = ~b & c;
  assign new_n1069_ = ~new_n404_ & new_n1068_;
  assign new_n1070_ = c & new_n251_;
  assign new_n1071_ = ~new_n404_ & new_n1070_;
  assign new_n1072_ = e2 & new_n404_;
  assign new_n1073_ = ~new_n1067_ & ~new_n1069_;
  assign new_n1074_ = ~new_n1071_ & ~new_n1072_;
  assign x4 = ~new_n1073_ | ~new_n1074_;
  assign new_n1076_ = t0 & l3;
  assign new_n1077_ = g0 & new_n1076_;
  assign y5 = ~new_n518_ | new_n1077_;
  assign new_n1079_ = k2 & ~l2;
  assign new_n1080_ = k2 & ~new_n471_;
  assign new_n1081_ = ~new_n1079_ & ~new_n1080_;
  assign x5 = new_n721_ | ~new_n1081_;
  assign new_n1083_ = v0 & ~x3;
  assign y4 = a | new_n1083_;
  assign new_n1085_ = k & ~d0;
  assign new_n1086_ = m & d0;
  assign z7 = new_n1085_ | new_n1086_;
  assign x6 = ~w0 & ~x0;
  assign y7 = p3 & j3;
  assign z4 = v0 & b4;
  assign new_n1091_ = r & k3;
  assign new_n1092_ = ~p3 & r;
  assign new_n1093_ = s2 & u0;
  assign new_n1094_ = ~new_n1091_ & ~new_n1092_;
  assign x7 = new_n1093_ | ~new_n1094_;
  assign new_n1096_ = ~k2 & ~new_n523_;
  assign new_n1097_ = ~i2 & ~d8;
  assign z5 = ~new_n1096_ | ~new_n1097_;
  assign new_n1099_ = ~e1 & l2;
  assign new_n1100_ = ~d1 & new_n1099_;
  assign new_n1101_ = ~p & q;
  assign new_n1102_ = n & new_n1101_;
  assign new_n1103_ = l2 & ~new_n1102_;
  assign e5 = new_n1100_ | new_n1103_;
  assign new_n1105_ = p2 & m2;
  assign new_n1106_ = q2 & m2;
  assign new_n1107_ = r0 & m2;
  assign new_n1108_ = ~new_n1105_ & ~new_n1106_;
  assign f6 = new_n1107_ | ~new_n1108_;
  assign new_n1110_ = y1 & m2;
  assign new_n1111_ = ~x1 & new_n1110_;
  assign new_n1112_ = ~q2 & new_n1111_;
  assign new_n1113_ = q2 & ~m2;
  assign new_n1114_ = p2 & new_n1113_;
  assign new_n1115_ = q & new_n1114_;
  assign new_n1116_ = ~p2 & new_n1111_;
  assign new_n1117_ = ~new_n1112_ & ~new_n1115_;
  assign new_n1118_ = ~new_n1116_ & new_n1117_;
  assign new_n1119_ = ~k1 & ~new_n1118_;
  assign new_n1120_ = q3 & new_n1118_;
  assign g7 = new_n1119_ | new_n1120_;
  assign new_n1122_ = ~w2 & d8;
  assign new_n1123_ = ~w2 & ~x2;
  assign h8 = new_n1122_ | new_n1123_;
  assign new_n1125_ = ~d1 & l2;
  assign new_n1126_ = ~e1 & new_n1125_;
  assign new_n1127_ = ~c1 & new_n1126_;
  assign d5 = new_n1103_ | new_n1127_;
  assign new_n1129_ = m1 & m2;
  assign f7 = ~new_n1108_ | new_n1129_;
  assign new_n1131_ = p & new_n1114_;
  assign new_n1132_ = ~q2 & m2;
  assign new_n1133_ = x1 & new_n1132_;
  assign new_n1134_ = ~y1 & new_n1133_;
  assign new_n1135_ = r0 & new_n1134_;
  assign new_n1136_ = ~p2 & m2;
  assign new_n1137_ = x1 & new_n1136_;
  assign new_n1138_ = ~y1 & new_n1137_;
  assign new_n1139_ = r0 & new_n1138_;
  assign new_n1140_ = ~new_n1135_ & ~new_n1139_;
  assign new_n1141_ = ~new_n1131_ & new_n1140_;
  assign new_n1142_ = ~p0 & ~new_n1141_;
  assign new_n1143_ = v3 & new_n1141_;
  assign g6 = new_n1142_ | new_n1143_;
  assign new_n1145_ = y3 & l3;
  assign new_n1146_ = z3 & new_n1145_;
  assign new_n1147_ = new_n958_ & new_n1146_;
  assign new_n1148_ = y3 & s;
  assign new_n1149_ = z3 & new_n1148_;
  assign new_n1150_ = new_n958_ & new_n1149_;
  assign e7 = new_n1147_ | new_n1150_;
  assign new_n1152_ = e0 & y;
  assign new_n1153_ = x & ~y;
  assign new_n1154_ = j1 & new_n1153_;
  assign new_n1155_ = e0 & ~x;
  assign new_n1156_ = ~new_n1152_ & ~new_n1154_;
  assign f4 = new_n1155_ | ~new_n1156_;
  assign g5 = new_n1099_ | new_n1103_;
  assign new_n1159_ = q2 & l2;
  assign new_n1160_ = p2 & new_n1159_;
  assign new_n1161_ = q & new_n1160_;
  assign new_n1162_ = q2 & ~new_n1161_;
  assign new_n1163_ = i1 & new_n1162_;
  assign new_n1164_ = ~s1 & m1;
  assign new_n1165_ = ~new_n1161_ & new_n1164_;
  assign new_n1166_ = i1 & new_n1165_;
  assign new_n1167_ = ~l2 & ~new_n1161_;
  assign new_n1168_ = i1 & new_n1167_;
  assign new_n1169_ = p2 & ~new_n1161_;
  assign new_n1170_ = i1 & new_n1169_;
  assign new_n1171_ = i1 & ~new_n1161_;
  assign new_n1172_ = ~q & new_n1171_;
  assign new_n1173_ = ~y3 & o1;
  assign new_n1174_ = ~new_n1161_ & new_n1173_;
  assign new_n1175_ = ~s1 & new_n1174_;
  assign new_n1176_ = m1 & new_n1175_;
  assign new_n1177_ = new_n290_ & new_n1174_;
  assign new_n1178_ = m1 & new_n1177_;
  assign new_n1179_ = ~y3 & ~new_n1161_;
  assign new_n1180_ = o1 & new_n1179_;
  assign new_n1181_ = q2 & new_n1180_;
  assign new_n1182_ = ~l2 & new_n1180_;
  assign new_n1183_ = p2 & new_n1180_;
  assign new_n1184_ = m1 & new_n290_;
  assign new_n1185_ = ~new_n1161_ & new_n1184_;
  assign new_n1186_ = i1 & new_n1185_;
  assign new_n1187_ = ~q & new_n1180_;
  assign new_n1188_ = ~new_n1183_ & ~new_n1186_;
  assign new_n1189_ = ~new_n1187_ & new_n1188_;
  assign new_n1190_ = ~new_n1178_ & ~new_n1181_;
  assign new_n1191_ = ~new_n1182_ & new_n1190_;
  assign new_n1192_ = new_n1189_ & new_n1191_;
  assign new_n1193_ = ~new_n1163_ & ~new_n1166_;
  assign new_n1194_ = ~new_n1168_ & new_n1193_;
  assign new_n1195_ = ~new_n1170_ & ~new_n1172_;
  assign new_n1196_ = ~new_n1176_ & new_n1195_;
  assign new_n1197_ = new_n1194_ & new_n1196_;
  assign d7 = ~new_n1192_ | ~new_n1197_;
  assign new_n1199_ = p2 & ~q2;
  assign new_n1200_ = ~p2 & q2;
  assign e6 = new_n1199_ | new_n1200_;
  assign new_n1202_ = ~c1 & new_n1099_;
  assign f5 = new_n1103_ | new_n1202_;
  assign new_n1204_ = p0 & ~y1;
  assign new_n1205_ = y1 & k1;
  assign g4 = new_n1204_ | new_n1205_;
  assign new_n1207_ = ~new_n1106_ & ~new_n1129_;
  assign b6 = new_n1107_ | ~new_n1207_;
  assign new_n1209_ = ~y3 & new_n290_;
  assign new_n1210_ = o1 & new_n1209_;
  assign new_n1211_ = ~new_n1161_ & new_n1210_;
  assign new_n1212_ = new_n290_ & ~new_n1161_;
  assign new_n1213_ = m1 & new_n1212_;
  assign new_n1214_ = ~s1 & ~y3;
  assign new_n1215_ = o1 & new_n1214_;
  assign new_n1216_ = ~new_n1161_ & new_n1215_;
  assign new_n1217_ = ~s1 & ~new_n1161_;
  assign new_n1218_ = m1 & new_n1217_;
  assign new_n1219_ = ~new_n1211_ & ~new_n1213_;
  assign new_n1220_ = ~new_n1216_ & ~new_n1218_;
  assign c7 = ~new_n1219_ | ~new_n1220_;
  assign new_n1222_ = x1 & m2;
  assign new_n1223_ = ~y1 & new_n1222_;
  assign c6 = w1 & new_n1223_;
  assign new_n1225_ = e1 & ~d1;
  assign new_n1226_ = ~e1 & d1;
  assign new_n1227_ = c1 & new_n1226_;
  assign new_n1228_ = ~c1 & e1;
  assign new_n1229_ = ~new_n1225_ & ~new_n1227_;
  assign c5 = new_n1228_ | ~new_n1229_;
  assign new_n1231_ = ~y & n0;
  assign new_n1232_ = ~x & y;
  assign new_n1233_ = e0 & new_n1232_;
  assign new_n1234_ = x & n0;
  assign new_n1235_ = ~new_n1231_ & ~new_n1233_;
  assign a6 = new_n1234_ | ~new_n1235_;
  assign new_n1237_ = c1 & ~d1;
  assign new_n1238_ = ~c1 & d1;
  assign b5 = new_n1237_ | new_n1238_;
  assign new_n1240_ = s1 & ~r1;
  assign new_n1241_ = ~d & new_n1240_;
  assign new_n1242_ = ~e & new_n1240_;
  assign new_n1243_ = ~e & b1;
  assign new_n1244_ = ~f & b1;
  assign new_n1245_ = ~d & b1;
  assign new_n1246_ = ~f & new_n1240_;
  assign new_n1247_ = ~new_n1241_ & ~new_n1242_;
  assign new_n1248_ = ~new_n1243_ & new_n1247_;
  assign new_n1249_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1250_ = ~new_n1246_ & new_n1249_;
  assign m5 = ~new_n1248_ | ~new_n1250_;
  assign new_n1252_ = i3 & ~new_n717_;
  assign new_n1253_ = ~i3 & new_n717_;
  assign new_n1254_ = h3 & new_n1253_;
  assign new_n1255_ = ~new_n1252_ & ~new_n1254_;
  assign n6 = new_n808_ | ~new_n1255_;
  assign new_n1257_ = ~new_n392_ & new_n441_;
  assign o7 = ~new_n363_ | new_n1257_;
  assign a8 = c4 | new_n789_;
  assign new_n1260_ = c1 & e1;
  assign new_n1261_ = d1 & new_n1260_;
  assign l5 = n & new_n1261_;
  assign n7 = new_n363_ & new_n392_;
  assign new_n1264_ = z2 & new_n824_;
  assign new_n1265_ = new_n675_ & new_n711_;
  assign new_n1266_ = z2 & new_n1265_;
  assign new_n1267_ = ~u & new_n854_;
  assign new_n1268_ = ~h0 & new_n846_;
  assign new_n1269_ = new_n675_ & ~new_n820_;
  assign new_n1270_ = z2 & new_n1269_;
  assign new_n1271_ = ~new_n1268_ & ~new_n1270_;
  assign new_n1272_ = ~new_n1264_ & ~new_n1266_;
  assign new_n1273_ = ~new_n1267_ & new_n1272_;
  assign o6 = ~new_n1271_ | ~new_n1273_;
  assign new_n1275_ = x2 & new_n337_;
  assign new_n1276_ = new_n296_ & new_n1275_;
  assign b8 = ~w2 & new_n1276_;
  assign new_n1278_ = ~i3 & m2;
  assign new_n1279_ = ~k2 & new_n1278_;
  assign new_n1280_ = p2 & ~k2;
  assign new_n1281_ = h3 & m2;
  assign new_n1282_ = ~k2 & new_n1281_;
  assign k6 = ~k2 & ~m0;
  assign new_n1284_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1285_ = ~new_n1282_ & ~k6;
  assign l6 = ~new_n1284_ | ~new_n1285_;
  assign new_n1287_ = new_n363_ & ~new_n392_;
  assign m7 = ~new_n441_ & new_n1287_;
  assign new_n1289_ = d1 & new_n1111_;
  assign new_n1290_ = e1 & new_n1289_;
  assign new_n1291_ = c1 & new_n1290_;
  assign new_n1292_ = ~n & new_n1111_;
  assign new_n1293_ = ~w1 & new_n296_;
  assign new_n1294_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1295_ = new_n1140_ & ~new_n1293_;
  assign n4 = ~new_n1294_ | ~new_n1295_;
  assign new_n1297_ = f2 & ~l2;
  assign new_n1298_ = h2 & new_n1297_;
  assign new_n1299_ = h2 & ~l2;
  assign new_n1300_ = ~g2 & new_n1299_;
  assign o5 = new_n1298_ | new_n1300_;
  assign new_n1302_ = w2 & ~new_n296_;
  assign c8 = ~a4 | new_n1302_;
  assign new_n1304_ = s & ~l3;
  assign new_n1305_ = u2 & new_n404_;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign l7 = new_n392_ | ~new_n1306_;
  assign new_n1308_ = h3 & ~new_n717_;
  assign new_n1309_ = ~new_n808_ & ~new_n1308_;
  assign m6 = new_n533_ | ~new_n1309_;
  assign new_n1311_ = g2 & ~l2;
  assign new_n1312_ = h2 & new_n1311_;
  assign new_n1313_ = ~f2 & new_n1312_;
  assign n5 = a | new_n1313_;
  assign o4 = w1 & new_n296_;
  assign i5 = new_n1103_ | new_n1125_;
  assign new_n1317_ = ~q2 & ~new_n389_;
  assign new_n1318_ = r0 & new_n1317_;
  assign new_n1319_ = ~l2 & ~new_n389_;
  assign new_n1320_ = r0 & new_n1319_;
  assign new_n1321_ = ~p2 & ~new_n389_;
  assign new_n1322_ = r0 & new_n1321_;
  assign new_n1323_ = ~new_n1318_ & ~new_n1320_;
  assign new_n1324_ = ~new_n533_ & ~new_n1322_;
  assign j6 = ~new_n1323_ | ~new_n1324_;
  assign k7 = i1 | new_n1111_;
  assign new_n1327_ = ~c1 & new_n1125_;
  assign h5 = new_n1103_ | new_n1327_;
  assign j7 = ~m1 & ~d8;
  assign new_n1330_ = ~p0 & q0;
  assign new_n1331_ = ~new_n1141_ & new_n1330_;
  assign new_n1332_ = p0 & ~q0;
  assign new_n1333_ = ~new_n1141_ & new_n1332_;
  assign new_n1334_ = w3 & new_n1141_;
  assign new_n1335_ = ~new_n1331_ & ~new_n1333_;
  assign h6 = new_n1334_ | ~new_n1335_;
  assign i7 = y3 & new_n958_;
  assign new_n1338_ = ~k1 & l1;
  assign new_n1339_ = ~new_n1118_ & new_n1338_;
  assign new_n1340_ = k1 & ~l1;
  assign new_n1341_ = ~new_n1118_ & new_n1340_;
  assign new_n1342_ = r3 & new_n1118_;
  assign new_n1343_ = ~new_n1339_ & ~new_n1341_;
  assign h7 = new_n1342_ | ~new_n1343_;
  assign i6 = l3 & ~new_n527_;
  assign new_n1346_ = ~c1 & l2;
  assign j5 = new_n1103_ | new_n1346_;
  assign d6 = ~p2;
  assign l4 = ~o3;
  assign w7 = c0;
  assign v7 = b0;
  assign w6 = y0;
  assign u7 = a0;
  assign t7 = z;
  assign s7 = w;
  assign z6 = v6;
  assign y6 = w0;
  assign a5 = m2;
  assign b7 = z0;
  assign a7 = y0;
  assign m4 = t3;
  assign e8 = x6;
  assign f8 = w0;
  assign k5 = l2;
  assign g8 = x0;
  assign k4 = s3;
endmodule

