module top ( 
    pp, pq, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pa1, pa0, pb0, pc1, pr, pb1, pc0, ps, pd0, pt, pd1, pe0, pu, pf0, pv,
    pg0, pw, ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pq0,
    pr0, ps0, pt0, pu0, pv0, pw0, px0, py0, pz0  );
  input  pp, pq, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po;
  output pa1, pa0, pb0, pc1, pr, pb1, pc0, ps, pd0, pt, pd1, pe0, pu, pf0, pv,
    pg0, pw, ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pq0,
    pr0, ps0, pt0, pu0, pv0, pw0, px0, py0, pz0;
  wire new_n57_, new_n58_, new_n59_, new_n60_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n83_, new_n84_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n350_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_;
  assign new_n57_ = pp & ~po;
  assign new_n58_ = ~pm & new_n57_;
  assign new_n59_ = ~pn & new_n58_;
  assign new_n60_ = pl & new_n59_;
  assign pa1 = pq & new_n60_;
  assign new_n62_ = pn & po;
  assign new_n63_ = ~pl & new_n62_;
  assign new_n64_ = ~pm & new_n63_;
  assign new_n65_ = pg & new_n64_;
  assign new_n66_ = pp & new_n65_;
  assign new_n67_ = pq & new_n66_;
  assign new_n68_ = ~pp & ~po;
  assign new_n69_ = ~pm & new_n68_;
  assign new_n70_ = pn & new_n69_;
  assign new_n71_ = ~pl & new_n70_;
  assign pc0 = pq & new_n71_;
  assign new_n73_ = ~pn & po;
  assign new_n74_ = ~pl & new_n73_;
  assign new_n75_ = pm & new_n74_;
  assign new_n76_ = pg & new_n75_;
  assign new_n77_ = ~pp & new_n76_;
  assign new_n78_ = ~pq & new_n77_;
  assign new_n79_ = ~pm & new_n74_;
  assign new_n80_ = ~pk & new_n79_;
  assign new_n81_ = pp & new_n80_;
  assign pb0 = pq & new_n81_;
  assign new_n83_ = ~new_n78_ & ~pb0;
  assign new_n84_ = ~new_n67_ & ~pc0;
  assign pa0 = ~new_n83_ | ~new_n84_;
  assign new_n86_ = ~pn & new_n69_;
  assign new_n87_ = pl & new_n86_;
  assign new_n88_ = ~pq & new_n87_;
  assign new_n89_ = pp & po;
  assign new_n90_ = pm & new_n89_;
  assign new_n91_ = pn & new_n90_;
  assign new_n92_ = ~pl & new_n91_;
  assign new_n93_ = pq & new_n92_;
  assign pc1 = new_n88_ | new_n93_;
  assign new_n95_ = ~pm & ~pn;
  assign new_n96_ = pe & new_n95_;
  assign new_n97_ = pl & new_n96_;
  assign new_n98_ = pa & new_n97_;
  assign new_n99_ = ~pq & new_n98_;
  assign new_n100_ = po & new_n99_;
  assign new_n101_ = ~pp & new_n100_;
  assign new_n102_ = ~pl & new_n96_;
  assign new_n103_ = pb & new_n102_;
  assign new_n104_ = pq & new_n103_;
  assign new_n105_ = ~po & new_n104_;
  assign new_n106_ = pp & new_n105_;
  assign new_n107_ = ~pi & pj;
  assign new_n108_ = pe & new_n107_;
  assign new_n109_ = ph & new_n108_;
  assign new_n110_ = ~pc & new_n109_;
  assign new_n111_ = ~pq & new_n110_;
  assign new_n112_ = pp & new_n111_;
  assign new_n113_ = pn & new_n112_;
  assign new_n114_ = po & new_n113_;
  assign new_n115_ = ~pl & new_n114_;
  assign new_n116_ = pm & new_n115_;
  assign new_n117_ = ~pf & new_n107_;
  assign new_n118_ = ph & new_n117_;
  assign new_n119_ = pe & new_n118_;
  assign new_n120_ = ~pq & new_n119_;
  assign new_n121_ = pp & new_n120_;
  assign new_n122_ = pn & new_n121_;
  assign new_n123_ = po & new_n122_;
  assign new_n124_ = ~pl & new_n123_;
  assign new_n125_ = pm & new_n124_;
  assign new_n126_ = pb & new_n109_;
  assign new_n127_ = ~pq & new_n126_;
  assign new_n128_ = pp & new_n127_;
  assign new_n129_ = pn & new_n128_;
  assign new_n130_ = po & new_n129_;
  assign new_n131_ = ~pl & new_n130_;
  assign new_n132_ = pm & new_n131_;
  assign new_n133_ = pm & new_n57_;
  assign new_n134_ = pn & new_n133_;
  assign new_n135_ = pl & new_n134_;
  assign new_n136_ = pq & new_n135_;
  assign new_n137_ = pn & ~po;
  assign new_n138_ = ~pl & new_n137_;
  assign new_n139_ = pm & new_n138_;
  assign new_n140_ = ~pg & new_n139_;
  assign new_n141_ = pp & new_n140_;
  assign new_n142_ = pq & new_n141_;
  assign new_n143_ = pl & new_n73_;
  assign new_n144_ = ~pm & new_n143_;
  assign new_n145_ = ~pg & new_n144_;
  assign new_n146_ = pp & new_n145_;
  assign new_n147_ = pq & new_n146_;
  assign new_n148_ = pm & new_n68_;
  assign new_n149_ = pn & new_n148_;
  assign new_n150_ = pl & new_n149_;
  assign new_n151_ = ~pq & new_n150_;
  assign new_n152_ = ~pm & new_n89_;
  assign new_n153_ = ~pn & new_n152_;
  assign new_n154_ = ~pl & new_n153_;
  assign new_n155_ = ~pq & new_n154_;
  assign new_n156_ = ~pp & po;
  assign new_n157_ = ~pm & new_n156_;
  assign new_n158_ = ~pn & new_n157_;
  assign new_n159_ = pl & new_n158_;
  assign new_n160_ = pq & new_n159_;
  assign new_n161_ = ~pl & new_n158_;
  assign new_n162_ = ~pq & new_n161_;
  assign new_n163_ = pl & new_n153_;
  assign new_n164_ = ~pq & new_n163_;
  assign new_n165_ = ~pq & new_n71_;
  assign new_n166_ = ~pn & new_n148_;
  assign new_n167_ = ~pl & new_n166_;
  assign new_n168_ = ~pq & new_n167_;
  assign new_n169_ = pm & new_n156_;
  assign new_n170_ = ~pn & new_n169_;
  assign new_n171_ = pl & new_n170_;
  assign new_n172_ = ~pq & new_n171_;
  assign new_n173_ = pn & new_n157_;
  assign new_n174_ = ~pl & new_n173_;
  assign new_n175_ = pq & new_n174_;
  assign new_n176_ = ~pq & new_n60_;
  assign new_n177_ = ~pn & new_n90_;
  assign new_n178_ = ~pl & new_n177_;
  assign new_n179_ = pq & new_n178_;
  assign new_n180_ = pf & new_n95_;
  assign new_n181_ = ~pl & new_n180_;
  assign new_n182_ = ~pb & new_n181_;
  assign new_n183_ = pq & new_n182_;
  assign new_n184_ = ~po & new_n183_;
  assign new_n185_ = pp & new_n184_;
  assign new_n186_ = ~pg & new_n75_;
  assign new_n187_ = pp & new_n186_;
  assign new_n188_ = ~pq & new_n187_;
  assign new_n189_ = ~pn & new_n133_;
  assign new_n190_ = pl & new_n189_;
  assign new_n191_ = pq & new_n190_;
  assign new_n192_ = ~pm & new_n138_;
  assign new_n193_ = pi & new_n192_;
  assign new_n194_ = pp & new_n193_;
  assign new_n195_ = pq & new_n194_;
  assign new_n196_ = pq & new_n161_;
  assign new_n197_ = ~pq & new_n174_;
  assign new_n198_ = ~pl & new_n59_;
  assign new_n199_ = ~pq & new_n198_;
  assign new_n200_ = ~pf & new_n192_;
  assign new_n201_ = pp & new_n200_;
  assign new_n202_ = ~pq & new_n201_;
  assign new_n203_ = pf & new_n192_;
  assign new_n204_ = pp & new_n203_;
  assign new_n205_ = ~pq & new_n204_;
  assign new_n206_ = pg & new_n144_;
  assign new_n207_ = pp & new_n206_;
  assign new_n208_ = pq & new_n207_;
  assign new_n209_ = ~pf & new_n95_;
  assign new_n210_ = ~pl & new_n209_;
  assign new_n211_ = pe & new_n210_;
  assign new_n212_ = pq & new_n211_;
  assign new_n213_ = ~po & new_n212_;
  assign new_n214_ = pp & new_n213_;
  assign new_n215_ = ~pn & ~po;
  assign new_n216_ = ~pl & new_n215_;
  assign new_n217_ = ~pm & new_n216_;
  assign new_n218_ = pc & new_n217_;
  assign new_n219_ = ~pp & new_n218_;
  assign new_n220_ = pq & new_n219_;
  assign new_n221_ = ~new_n78_ & ~new_n168_;
  assign new_n222_ = ~new_n164_ & ~new_n165_;
  assign new_n223_ = new_n221_ & new_n222_;
  assign new_n224_ = ~new_n160_ & ~new_n162_;
  assign new_n225_ = ~new_n151_ & ~new_n155_;
  assign new_n226_ = new_n224_ & new_n225_;
  assign new_n227_ = new_n223_ & new_n226_;
  assign new_n228_ = ~new_n142_ & ~new_n147_;
  assign new_n229_ = ~new_n67_ & ~new_n136_;
  assign new_n230_ = new_n228_ & new_n229_;
  assign new_n231_ = ~new_n125_ & ~new_n132_;
  assign new_n232_ = ~new_n101_ & ~new_n106_;
  assign new_n233_ = ~new_n116_ & new_n232_;
  assign new_n234_ = new_n231_ & new_n233_;
  assign new_n235_ = new_n230_ & new_n234_;
  assign new_n236_ = new_n227_ & new_n235_;
  assign new_n237_ = ~new_n214_ & ~new_n220_;
  assign new_n238_ = ~new_n205_ & ~new_n208_;
  assign new_n239_ = new_n237_ & new_n238_;
  assign new_n240_ = ~new_n196_ & ~new_n197_;
  assign new_n241_ = ~new_n199_ & ~new_n202_;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = new_n239_ & new_n242_;
  assign new_n244_ = ~new_n191_ & ~new_n195_;
  assign new_n245_ = ~new_n185_ & ~new_n188_;
  assign new_n246_ = new_n244_ & new_n245_;
  assign new_n247_ = ~new_n172_ & ~new_n175_;
  assign new_n248_ = ~new_n176_ & ~new_n179_;
  assign new_n249_ = new_n247_ & new_n248_;
  assign new_n250_ = new_n246_ & new_n249_;
  assign new_n251_ = new_n243_ & new_n250_;
  assign pr = ~new_n236_ | ~new_n251_;
  assign new_n253_ = pm & pn;
  assign new_n254_ = pj & new_n253_;
  assign new_n255_ = ~pl & new_n254_;
  assign new_n256_ = ph & new_n255_;
  assign new_n257_ = ~pq & new_n256_;
  assign new_n258_ = po & new_n257_;
  assign pb1 = ~pp & new_n258_;
  assign new_n260_ = ~pl & pm;
  assign new_n261_ = ~pf & new_n260_;
  assign new_n262_ = ~pi & new_n261_;
  assign new_n263_ = ~pe & new_n262_;
  assign new_n264_ = pp & new_n263_;
  assign new_n265_ = ~pq & new_n264_;
  assign new_n266_ = pn & new_n265_;
  assign new_n267_ = po & new_n266_;
  assign new_n268_ = ~pf & new_n215_;
  assign new_n269_ = ~pm & new_n268_;
  assign new_n270_ = ~pe & new_n269_;
  assign new_n271_ = pp & new_n270_;
  assign new_n272_ = pq & new_n271_;
  assign new_n273_ = ~pe & new_n260_;
  assign new_n274_ = ~pi & new_n273_;
  assign new_n275_ = pb & new_n274_;
  assign new_n276_ = pp & new_n275_;
  assign new_n277_ = ~pq & new_n276_;
  assign new_n278_ = pn & new_n277_;
  assign new_n279_ = po & new_n278_;
  assign new_n280_ = ~pc & new_n274_;
  assign new_n281_ = pp & new_n280_;
  assign new_n282_ = ~pq & new_n281_;
  assign new_n283_ = pn & new_n282_;
  assign new_n284_ = po & new_n283_;
  assign new_n285_ = pl & ~pm;
  assign new_n286_ = ~pe & new_n285_;
  assign new_n287_ = ~pf & new_n286_;
  assign new_n288_ = pa & new_n287_;
  assign new_n289_ = ~pp & new_n288_;
  assign new_n290_ = ~pq & new_n289_;
  assign new_n291_ = ~pn & new_n290_;
  assign new_n292_ = po & new_n291_;
  assign new_n293_ = ~pl & new_n86_;
  assign new_n294_ = ~pq & new_n293_;
  assign new_n295_ = pn & new_n152_;
  assign new_n296_ = pl & new_n295_;
  assign new_n297_ = ~pq & new_n296_;
  assign new_n298_ = ~pi & new_n253_;
  assign new_n299_ = ~pl & new_n298_;
  assign new_n300_ = ~ph & new_n299_;
  assign new_n301_ = po & new_n300_;
  assign new_n302_ = ~pq & new_n301_;
  assign new_n303_ = pm & new_n63_;
  assign new_n304_ = ~ph & new_n303_;
  assign new_n305_ = ~pp & new_n304_;
  assign new_n306_ = ~pq & new_n305_;
  assign new_n307_ = ~new_n284_ & ~new_n292_;
  assign new_n308_ = ~new_n267_ & ~new_n272_;
  assign new_n309_ = ~new_n279_ & new_n308_;
  assign new_n310_ = new_n307_ & new_n309_;
  assign new_n311_ = ~new_n302_ & ~new_n306_;
  assign new_n312_ = ~pa1 & ~new_n294_;
  assign new_n313_ = ~new_n297_ & new_n312_;
  assign new_n314_ = new_n311_ & new_n313_;
  assign ps = ~new_n310_ | ~new_n314_;
  assign new_n316_ = ph & ~pi;
  assign new_n317_ = pc & new_n316_;
  assign new_n318_ = pf & new_n317_;
  assign new_n319_ = ~pb & new_n318_;
  assign new_n320_ = ~pq & new_n319_;
  assign new_n321_ = pp & new_n320_;
  assign new_n322_ = pn & new_n321_;
  assign new_n323_ = po & new_n322_;
  assign new_n324_ = ~pl & new_n323_;
  assign new_n325_ = pm & new_n324_;
  assign new_n326_ = pl & new_n166_;
  assign new_n327_ = pq & new_n326_;
  assign new_n328_ = ~pq & po;
  assign new_n329_ = ~pm & new_n328_;
  assign new_n330_ = pn & new_n329_;
  assign new_n331_ = ~pl & new_n330_;
  assign new_n332_ = ~pq & ~po;
  assign new_n333_ = pm & new_n332_;
  assign new_n334_ = ~pn & new_n333_;
  assign new_n335_ = pl & new_n334_;
  assign new_n336_ = pn & new_n169_;
  assign new_n337_ = pl & new_n336_;
  assign new_n338_ = ~pq & new_n337_;
  assign new_n339_ = pp & ~pq;
  assign new_n340_ = pn & new_n339_;
  assign new_n341_ = ~po & new_n340_;
  assign new_n342_ = pm & new_n341_;
  assign new_n343_ = pq & new_n171_;
  assign new_n344_ = pm & new_n339_;
  assign new_n345_ = ~pn & new_n344_;
  assign new_n346_ = pl & new_n345_;
  assign new_n347_ = pl & new_n70_;
  assign new_n348_ = ~pq & new_n347_;
  assign pd1 = pq & new_n150_;
  assign new_n350_ = pq & new_n296_;
  assign pz0 = pq & new_n87_;
  assign new_n352_ = ~pl & new_n170_;
  assign new_n353_ = pq & new_n352_;
  assign new_n354_ = ~pl & new_n189_;
  assign new_n355_ = pq & new_n354_;
  assign new_n356_ = pl & new_n156_;
  assign new_n357_ = ~pn & new_n356_;
  assign new_n358_ = ~pa & new_n357_;
  assign new_n359_ = pk & new_n79_;
  assign new_n360_ = pp & new_n359_;
  assign new_n361_ = pq & new_n360_;
  assign new_n362_ = ~new_n279_ & ~new_n284_;
  assign new_n363_ = new_n308_ & new_n362_;
  assign new_n364_ = ~new_n358_ & ~new_n361_;
  assign new_n365_ = ~new_n302_ & ~new_n355_;
  assign new_n366_ = ~new_n297_ & new_n365_;
  assign new_n367_ = new_n364_ & new_n366_;
  assign new_n368_ = new_n363_ & new_n367_;
  assign new_n369_ = ~new_n88_ & ~new_n160_;
  assign new_n370_ = ~new_n353_ & new_n369_;
  assign new_n371_ = ~new_n147_ & ~new_n185_;
  assign new_n372_ = new_n370_ & new_n371_;
  assign new_n373_ = ~new_n350_ & ~pz0;
  assign new_n374_ = ~new_n306_ & ~pd1;
  assign new_n375_ = ~new_n164_ & new_n374_;
  assign new_n376_ = new_n373_ & new_n375_;
  assign new_n377_ = new_n372_ & new_n376_;
  assign new_n378_ = new_n368_ & new_n377_;
  assign new_n379_ = ~new_n191_ & ~new_n348_;
  assign new_n380_ = ~pa1 & ~new_n151_;
  assign new_n381_ = new_n379_ & new_n380_;
  assign new_n382_ = ~new_n343_ & ~new_n346_;
  assign new_n383_ = ~new_n176_ & ~new_n338_;
  assign new_n384_ = ~new_n342_ & new_n383_;
  assign new_n385_ = new_n382_ & new_n384_;
  assign new_n386_ = new_n381_ & new_n385_;
  assign new_n387_ = ~new_n132_ & ~new_n325_;
  assign new_n388_ = ~new_n116_ & ~new_n125_;
  assign new_n389_ = ~new_n292_ & new_n388_;
  assign new_n390_ = new_n387_ & new_n389_;
  assign new_n391_ = ~new_n172_ & ~new_n335_;
  assign new_n392_ = ~new_n208_ & ~new_n327_;
  assign new_n393_ = ~new_n331_ & new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = new_n390_ & new_n394_;
  assign new_n396_ = new_n386_ & new_n395_;
  assign pd0 = ~new_n378_ | ~new_n396_;
  assign new_n398_ = ~new_n199_ & ~new_n214_;
  assign new_n399_ = ~new_n220_ & new_n398_;
  assign new_n400_ = ~new_n147_ & ~new_n176_;
  assign new_n401_ = ~new_n196_ & new_n400_;
  assign new_n402_ = new_n399_ & new_n401_;
  assign new_n403_ = ~new_n136_ & ~new_n185_;
  assign new_n404_ = ~new_n142_ & new_n403_;
  assign new_n405_ = ~new_n191_ & ~new_n197_;
  assign new_n406_ = ~new_n188_ & ~new_n195_;
  assign new_n407_ = new_n405_ & new_n406_;
  assign new_n408_ = new_n404_ & new_n407_;
  assign new_n409_ = new_n402_ & new_n408_;
  assign new_n410_ = new_n232_ & new_n388_;
  assign new_n411_ = ~new_n132_ & ~new_n168_;
  assign new_n412_ = ~new_n172_ & new_n411_;
  assign new_n413_ = new_n410_ & new_n412_;
  assign new_n414_ = ~new_n155_ & ~new_n160_;
  assign new_n415_ = ~new_n162_ & new_n414_;
  assign new_n416_ = ~new_n164_ & ~new_n179_;
  assign new_n417_ = ~new_n151_ & ~new_n175_;
  assign new_n418_ = new_n416_ & new_n417_;
  assign new_n419_ = new_n415_ & new_n418_;
  assign new_n420_ = new_n413_ & new_n419_;
  assign pt = ~new_n409_ | ~new_n420_;
  assign new_n422_ = ~pj & ~pl;
  assign new_n423_ = pe & new_n422_;
  assign new_n424_ = ph & new_n423_;
  assign new_n425_ = ~pc & new_n424_;
  assign new_n426_ = po & new_n425_;
  assign new_n427_ = pp & new_n426_;
  assign new_n428_ = pm & new_n427_;
  assign new_n429_ = pn & new_n428_;
  assign new_n430_ = ~pf & new_n422_;
  assign new_n431_ = ph & new_n430_;
  assign new_n432_ = pe & new_n431_;
  assign new_n433_ = po & new_n432_;
  assign new_n434_ = pp & new_n433_;
  assign new_n435_ = pm & new_n434_;
  assign new_n436_ = pn & new_n435_;
  assign new_n437_ = ~pk & ~pl;
  assign new_n438_ = pg & new_n437_;
  assign new_n439_ = ~pi & new_n438_;
  assign new_n440_ = ~pc & new_n439_;
  assign new_n441_ = ~pq & new_n440_;
  assign new_n442_ = po & new_n441_;
  assign new_n443_ = pp & new_n442_;
  assign new_n444_ = pm & new_n443_;
  assign new_n445_ = ~pn & new_n444_;
  assign new_n446_ = pb & new_n424_;
  assign new_n447_ = po & new_n446_;
  assign new_n448_ = pp & new_n447_;
  assign new_n449_ = pm & new_n448_;
  assign new_n450_ = pn & new_n449_;
  assign new_n451_ = ~pm & pn;
  assign new_n452_ = ~pi & new_n451_;
  assign new_n453_ = ~pl & new_n452_;
  assign new_n454_ = ~pd & new_n453_;
  assign new_n455_ = pq & new_n454_;
  assign new_n456_ = ~po & new_n455_;
  assign new_n457_ = pp & new_n456_;
  assign new_n458_ = ~pq & new_n354_;
  assign new_n459_ = ~pp & ~pq;
  assign new_n460_ = pn & new_n459_;
  assign new_n461_ = po & new_n460_;
  assign new_n462_ = ~pm & new_n461_;
  assign new_n463_ = ~pp & pq;
  assign new_n464_ = pm & new_n463_;
  assign new_n465_ = ~po & new_n464_;
  assign new_n466_ = ~pl & new_n465_;
  assign new_n467_ = pn & new_n58_;
  assign new_n468_ = pl & new_n467_;
  assign new_n469_ = ~pq & new_n468_;
  assign new_n470_ = pi & new_n303_;
  assign new_n471_ = pp & new_n470_;
  assign new_n472_ = ~pq & new_n471_;
  assign new_n473_ = ~pl & new_n89_;
  assign new_n474_ = pn & new_n473_;
  assign new_n475_ = ~pg & new_n474_;
  assign new_n476_ = pq & new_n475_;
  assign new_n477_ = ~pl & new_n149_;
  assign new_n478_ = ~pq & new_n477_;
  assign new_n479_ = pp & pn;
  assign new_n480_ = ~pl & new_n479_;
  assign new_n481_ = pm & new_n480_;
  assign new_n482_ = pg & new_n481_;
  assign new_n483_ = pq & new_n482_;
  assign new_n484_ = ph & new_n303_;
  assign new_n485_ = ~pp & new_n484_;
  assign new_n486_ = ~pq & new_n485_;
  assign new_n487_ = ~pm & new_n463_;
  assign new_n488_ = pn & new_n487_;
  assign new_n489_ = pl & new_n488_;
  assign new_n490_ = ~pp & new_n186_;
  assign new_n491_ = ~pq & new_n490_;
  assign new_n492_ = ~new_n478_ & ~new_n483_;
  assign new_n493_ = ~pa1 & ~new_n476_;
  assign new_n494_ = new_n492_ & new_n493_;
  assign new_n495_ = ~new_n486_ & ~new_n489_;
  assign new_n496_ = ~new_n361_ & ~new_n491_;
  assign new_n497_ = new_n495_ & new_n496_;
  assign new_n498_ = new_n494_ & new_n497_;
  assign new_n499_ = ~new_n151_ & ~new_n350_;
  assign new_n500_ = ~new_n142_ & ~new_n472_;
  assign new_n501_ = new_n499_ & new_n500_;
  assign new_n502_ = ~new_n78_ & ~new_n191_;
  assign new_n503_ = ~new_n67_ & ~new_n188_;
  assign new_n504_ = ~new_n335_ & new_n503_;
  assign new_n505_ = new_n502_ & new_n504_;
  assign new_n506_ = new_n501_ & new_n505_;
  assign new_n507_ = new_n498_ & new_n506_;
  assign new_n508_ = ~new_n202_ & ~new_n469_;
  assign new_n509_ = ~new_n343_ & ~new_n466_;
  assign new_n510_ = new_n508_ & new_n509_;
  assign new_n511_ = ~new_n168_ & ~pd1;
  assign new_n512_ = ~new_n179_ & ~new_n462_;
  assign new_n513_ = new_n511_ & new_n512_;
  assign new_n514_ = new_n510_ & new_n513_;
  assign new_n515_ = ~new_n346_ & ~new_n458_;
  assign new_n516_ = ~new_n147_ & ~new_n457_;
  assign new_n517_ = new_n515_ & new_n516_;
  assign new_n518_ = ~new_n325_ & ~new_n450_;
  assign new_n519_ = ~new_n429_ & ~new_n436_;
  assign new_n520_ = ~new_n445_ & new_n519_;
  assign new_n521_ = new_n518_ & new_n520_;
  assign new_n522_ = new_n517_ & new_n521_;
  assign new_n523_ = new_n514_ & new_n522_;
  assign pe0 = ~new_n507_ | ~new_n523_;
  assign new_n525_ = pq & new_n477_;
  assign new_n526_ = pq & new_n347_;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = ~new_n458_ & new_n527_;
  assign new_n529_ = ~pc0 & ~new_n343_;
  assign new_n530_ = ~new_n350_ & new_n529_;
  assign pu = ~new_n528_ | ~new_n530_;
  assign new_n532_ = pf & new_n286_;
  assign new_n533_ = pa & new_n532_;
  assign new_n534_ = ~pq & new_n533_;
  assign new_n535_ = ~pn & new_n534_;
  assign new_n536_ = po & new_n535_;
  assign new_n537_ = ~pl & ~pm;
  assign new_n538_ = ~pe & new_n537_;
  assign new_n539_ = pf & new_n538_;
  assign new_n540_ = pb & new_n539_;
  assign new_n541_ = pp & new_n540_;
  assign new_n542_ = pq & new_n541_;
  assign new_n543_ = ~pn & new_n542_;
  assign new_n544_ = ~po & new_n543_;
  assign new_n545_ = pq & new_n468_;
  assign new_n546_ = pd & new_n453_;
  assign new_n547_ = pq & new_n546_;
  assign new_n548_ = ~po & new_n547_;
  assign new_n549_ = pp & new_n548_;
  assign new_n550_ = ~pl & new_n134_;
  assign new_n551_ = ~pq & new_n550_;
  assign new_n552_ = pm & ~pn;
  assign new_n553_ = pg & new_n552_;
  assign new_n554_ = ~pl & new_n553_;
  assign new_n555_ = pc & new_n554_;
  assign new_n556_ = ~pq & new_n555_;
  assign new_n557_ = po & new_n556_;
  assign new_n558_ = pp & new_n557_;
  assign new_n559_ = pi & new_n552_;
  assign new_n560_ = ~pl & new_n559_;
  assign new_n561_ = pg & new_n560_;
  assign new_n562_ = ~pq & new_n561_;
  assign new_n563_ = po & new_n562_;
  assign new_n564_ = pp & new_n563_;
  assign new_n565_ = pk & new_n552_;
  assign new_n566_ = ~pl & new_n565_;
  assign new_n567_ = pg & new_n566_;
  assign new_n568_ = ~pq & new_n567_;
  assign new_n569_ = po & new_n568_;
  assign new_n570_ = pp & new_n569_;
  assign new_n571_ = ~new_n348_ & ~new_n491_;
  assign new_n572_ = ~new_n486_ & new_n571_;
  assign new_n573_ = new_n519_ & new_n572_;
  assign new_n574_ = ~new_n476_ & ~new_n570_;
  assign new_n575_ = ~pc0 & ~new_n564_;
  assign new_n576_ = ~new_n483_ & new_n575_;
  assign new_n577_ = new_n574_ & new_n576_;
  assign new_n578_ = new_n573_ & new_n577_;
  assign new_n579_ = ~new_n172_ & ~new_n525_;
  assign new_n580_ = ~new_n165_ & ~pd1;
  assign new_n581_ = ~new_n472_ & new_n580_;
  assign new_n582_ = new_n579_ & new_n581_;
  assign new_n583_ = ~pa1 & ~new_n353_;
  assign new_n584_ = ~new_n478_ & ~new_n558_;
  assign new_n585_ = ~new_n202_ & new_n584_;
  assign new_n586_ = new_n583_ & new_n585_;
  assign new_n587_ = new_n582_ & new_n586_;
  assign new_n588_ = new_n578_ & new_n587_;
  assign new_n589_ = ~new_n195_ & ~new_n551_;
  assign new_n590_ = ~new_n147_ & ~new_n549_;
  assign new_n591_ = ~new_n462_ & new_n590_;
  assign new_n592_ = new_n589_ & new_n591_;
  assign new_n593_ = ~new_n179_ & ~new_n331_;
  assign new_n594_ = ~new_n164_ & ~new_n208_;
  assign new_n595_ = ~new_n355_ & new_n594_;
  assign new_n596_ = new_n593_ & new_n595_;
  assign new_n597_ = new_n592_ & new_n596_;
  assign new_n598_ = ~pb0 & ~new_n205_;
  assign new_n599_ = ~new_n88_ & ~new_n545_;
  assign new_n600_ = ~new_n136_ & new_n599_;
  assign new_n601_ = new_n598_ & new_n600_;
  assign new_n602_ = ~new_n325_ & ~new_n544_;
  assign new_n603_ = ~new_n175_ & new_n602_;
  assign new_n604_ = ~new_n450_ & ~new_n536_;
  assign new_n605_ = ~new_n445_ & new_n604_;
  assign new_n606_ = new_n603_ & new_n605_;
  assign new_n607_ = new_n601_ & new_n606_;
  assign new_n608_ = new_n597_ & new_n607_;
  assign pf0 = ~new_n588_ | ~new_n608_;
  assign new_n610_ = ~new_n526_ & ~new_n558_;
  assign new_n611_ = ~new_n208_ & ~new_n350_;
  assign new_n612_ = new_n610_ & new_n611_;
  assign new_n613_ = ~new_n343_ & ~new_n525_;
  assign new_n614_ = ~pc0 & ~new_n458_;
  assign new_n615_ = new_n613_ & new_n614_;
  assign new_n616_ = new_n612_ & new_n615_;
  assign new_n617_ = ~new_n67_ & ~new_n78_;
  assign new_n618_ = ~new_n165_ & ~new_n457_;
  assign new_n619_ = new_n617_ & new_n618_;
  assign new_n620_ = ~pb0 & ~new_n549_;
  assign new_n621_ = ~new_n564_ & ~new_n570_;
  assign new_n622_ = new_n620_ & new_n621_;
  assign new_n623_ = new_n619_ & new_n622_;
  assign pv = ~new_n616_ | ~new_n623_;
  assign new_n625_ = pl & new_n177_;
  assign new_n626_ = ~new_n272_ & ~new_n279_;
  assign new_n627_ = ~new_n284_ & new_n626_;
  assign new_n628_ = ~new_n302_ & ~new_n491_;
  assign new_n629_ = ~new_n267_ & new_n628_;
  assign new_n630_ = new_n627_ & new_n629_;
  assign new_n631_ = ~new_n338_ & ~new_n486_;
  assign new_n632_ = ~new_n327_ & new_n631_;
  assign new_n633_ = ~new_n185_ & ~new_n625_;
  assign new_n634_ = ~new_n549_ & new_n633_;
  assign new_n635_ = new_n632_ & new_n634_;
  assign new_n636_ = new_n630_ & new_n635_;
  assign new_n637_ = ~new_n472_ & ~new_n483_;
  assign new_n638_ = ~new_n155_ & new_n637_;
  assign new_n639_ = ~new_n162_ & ~new_n489_;
  assign new_n640_ = ~new_n564_ & new_n639_;
  assign new_n641_ = new_n638_ & new_n640_;
  assign new_n642_ = ~new_n195_ & ~new_n570_;
  assign new_n643_ = ~new_n545_ & new_n642_;
  assign new_n644_ = ~new_n172_ & ~new_n306_;
  assign new_n645_ = ~pa1 & ~new_n106_;
  assign new_n646_ = new_n644_ & new_n645_;
  assign new_n647_ = new_n643_ & new_n646_;
  assign new_n648_ = new_n641_ & new_n647_;
  assign new_n649_ = new_n636_ & new_n648_;
  assign new_n650_ = ~new_n214_ & ~new_n358_;
  assign new_n651_ = ~new_n164_ & new_n650_;
  assign new_n652_ = ~new_n142_ & ~new_n469_;
  assign new_n653_ = ~new_n558_ & new_n652_;
  assign new_n654_ = new_n651_ & new_n653_;
  assign new_n655_ = ~new_n136_ & ~new_n202_;
  assign new_n656_ = ~new_n297_ & new_n655_;
  assign new_n657_ = ~new_n101_ & ~new_n355_;
  assign new_n658_ = new_n369_ & new_n657_;
  assign new_n659_ = new_n656_ & new_n658_;
  assign new_n660_ = new_n654_ & new_n659_;
  assign new_n661_ = ~new_n343_ & ~new_n457_;
  assign new_n662_ = ~new_n551_ & new_n661_;
  assign new_n663_ = ~new_n346_ & ~new_n476_;
  assign new_n664_ = ~new_n188_ & new_n663_;
  assign new_n665_ = new_n662_ & new_n664_;
  assign new_n666_ = ~new_n292_ & ~new_n450_;
  assign new_n667_ = new_n519_ & new_n666_;
  assign new_n668_ = ~new_n191_ & ~new_n445_;
  assign new_n669_ = ~new_n196_ & new_n668_;
  assign new_n670_ = new_n667_ & new_n669_;
  assign new_n671_ = new_n665_ & new_n670_;
  assign new_n672_ = new_n660_ & new_n671_;
  assign pg0 = ~new_n649_ | ~new_n672_;
  assign new_n674_ = ~pl & pn;
  assign new_n675_ = ~pg & new_n674_;
  assign new_n676_ = ~pi & new_n675_;
  assign new_n677_ = ~pc & new_n676_;
  assign new_n678_ = pq & new_n677_;
  assign new_n679_ = po & new_n678_;
  assign new_n680_ = pp & new_n679_;
  assign new_n681_ = ~pb1 & ~new_n436_;
  assign new_n682_ = ~new_n361_ & ~new_n469_;
  assign new_n683_ = ~new_n466_ & new_n682_;
  assign new_n684_ = new_n681_ & new_n683_;
  assign new_n685_ = ~new_n353_ & ~new_n564_;
  assign new_n686_ = ~new_n343_ & ~new_n558_;
  assign new_n687_ = ~pz0 & new_n686_;
  assign new_n688_ = new_n685_ & new_n687_;
  assign new_n689_ = new_n684_ & new_n688_;
  assign new_n690_ = ~new_n188_ & ~new_n199_;
  assign new_n691_ = ~new_n205_ & ~new_n545_;
  assign new_n692_ = ~new_n172_ & new_n691_;
  assign new_n693_ = new_n690_ & new_n692_;
  assign new_n694_ = ~new_n93_ & ~new_n680_;
  assign new_n695_ = ~new_n458_ & new_n694_;
  assign new_n696_ = ~new_n176_ & ~new_n472_;
  assign new_n697_ = ~new_n88_ & new_n696_;
  assign new_n698_ = new_n695_ & new_n697_;
  assign new_n699_ = new_n693_ & new_n698_;
  assign new_n700_ = new_n689_ & new_n699_;
  assign new_n701_ = ~new_n220_ & ~new_n331_;
  assign new_n702_ = ~pc0 & ~new_n625_;
  assign new_n703_ = ~new_n151_ & new_n702_;
  assign new_n704_ = new_n701_ & new_n703_;
  assign new_n705_ = ~new_n445_ & ~new_n536_;
  assign new_n706_ = ~new_n160_ & new_n705_;
  assign new_n707_ = ~new_n429_ & ~new_n450_;
  assign new_n708_ = ~new_n544_ & new_n707_;
  assign new_n709_ = new_n706_ & new_n708_;
  assign new_n710_ = new_n704_ & new_n709_;
  assign new_n711_ = ~new_n164_ & ~new_n462_;
  assign new_n712_ = ~new_n155_ & ~pd1;
  assign new_n713_ = ~new_n327_ & new_n712_;
  assign new_n714_ = new_n711_ & new_n713_;
  assign new_n715_ = ~new_n175_ & ~new_n196_;
  assign new_n716_ = ~new_n549_ & new_n715_;
  assign new_n717_ = ~new_n142_ & ~new_n202_;
  assign new_n718_ = ~new_n570_ & new_n717_;
  assign new_n719_ = new_n716_ & new_n718_;
  assign new_n720_ = new_n714_ & new_n719_;
  assign new_n721_ = new_n710_ & new_n720_;
  assign ph0 = ~new_n700_ | ~new_n721_;
  assign new_n723_ = ~pc & new_n217_;
  assign new_n724_ = ~pp & new_n723_;
  assign new_n725_ = ~new_n125_ & ~new_n348_;
  assign new_n726_ = ~new_n294_ & ~new_n478_;
  assign new_n727_ = new_n725_ & new_n726_;
  assign new_n728_ = ~new_n327_ & ~new_n472_;
  assign new_n729_ = ~new_n165_ & ~new_n335_;
  assign new_n730_ = ~new_n199_ & new_n729_;
  assign new_n731_ = new_n728_ & new_n730_;
  assign new_n732_ = new_n727_ & new_n731_;
  assign new_n733_ = ~new_n188_ & ~new_n355_;
  assign new_n734_ = ~new_n151_ & ~new_n457_;
  assign new_n735_ = ~new_n155_ & new_n734_;
  assign new_n736_ = new_n733_ & new_n735_;
  assign new_n737_ = ~new_n458_ & ~new_n625_;
  assign new_n738_ = ~new_n136_ & ~new_n142_;
  assign new_n739_ = new_n737_ & new_n738_;
  assign new_n740_ = new_n736_ & new_n739_;
  assign new_n741_ = new_n732_ & new_n740_;
  assign new_n742_ = ~new_n162_ & ~new_n526_;
  assign new_n743_ = ~new_n168_ & ~new_n462_;
  assign new_n744_ = new_n742_ & new_n743_;
  assign new_n745_ = ~new_n325_ & ~new_n536_;
  assign new_n746_ = ~new_n116_ & ~new_n132_;
  assign new_n747_ = ~new_n544_ & new_n746_;
  assign new_n748_ = new_n745_ & new_n747_;
  assign new_n749_ = new_n744_ & new_n748_;
  assign new_n750_ = ~new_n185_ & ~new_n545_;
  assign new_n751_ = ~new_n176_ & ~new_n724_;
  assign new_n752_ = new_n750_ & new_n751_;
  assign new_n753_ = ~new_n172_ & ~new_n331_;
  assign new_n754_ = ~new_n175_ & ~new_n205_;
  assign new_n755_ = ~new_n164_ & new_n754_;
  assign new_n756_ = new_n753_ & new_n755_;
  assign new_n757_ = new_n752_ & new_n756_;
  assign new_n758_ = new_n749_ & new_n757_;
  assign pi0 = ~new_n741_ | ~new_n758_;
  assign new_n760_ = ~new_n67_ & ~new_n458_;
  assign new_n761_ = ~new_n78_ & ~new_n457_;
  assign new_n762_ = new_n760_ & new_n761_;
  assign new_n763_ = new_n622_ & new_n762_;
  assign new_n764_ = ~new_n350_ & ~new_n525_;
  assign new_n765_ = new_n529_ & new_n764_;
  assign new_n766_ = ~new_n208_ & ~new_n558_;
  assign new_n767_ = ~new_n526_ & new_n766_;
  assign new_n768_ = new_n765_ & new_n767_;
  assign py = ~new_n763_ | ~new_n768_;
  assign new_n770_ = ~new_n294_ & ~new_n306_;
  assign new_n771_ = ~new_n297_ & ~new_n338_;
  assign new_n772_ = new_n770_ & new_n771_;
  assign new_n773_ = ~new_n267_ & ~new_n302_;
  assign new_n774_ = ~new_n279_ & new_n773_;
  assign new_n775_ = new_n307_ & new_n774_;
  assign pj0 = ~new_n772_ | ~new_n775_;
  assign pz = new_n155_ | new_n162_;
  assign new_n778_ = ~new_n67_ & ~new_n151_;
  assign new_n779_ = ~new_n188_ & ~new_n292_;
  assign new_n780_ = new_n778_ & new_n779_;
  assign new_n781_ = ~pb1 & ~new_n267_;
  assign new_n782_ = new_n362_ & new_n781_;
  assign new_n783_ = new_n780_ & new_n782_;
  assign new_n784_ = ~new_n147_ & ~new_n172_;
  assign new_n785_ = new_n405_ & new_n784_;
  assign new_n786_ = ~new_n142_ & ~new_n195_;
  assign new_n787_ = ~new_n88_ & new_n786_;
  assign new_n788_ = new_n785_ & new_n787_;
  assign new_n789_ = new_n783_ & new_n788_;
  assign new_n790_ = ~new_n302_ & ~new_n338_;
  assign new_n791_ = ~new_n306_ & new_n790_;
  assign new_n792_ = ~new_n93_ & ~new_n294_;
  assign new_n793_ = new_n511_ & new_n792_;
  assign new_n794_ = new_n791_ & new_n793_;
  assign new_n795_ = ~new_n78_ & ~new_n160_;
  assign new_n796_ = ~new_n175_ & ~new_n208_;
  assign new_n797_ = new_n795_ & new_n796_;
  assign new_n798_ = ~new_n179_ & ~new_n297_;
  assign new_n799_ = new_n403_ & new_n798_;
  assign new_n800_ = new_n797_ & new_n799_;
  assign new_n801_ = new_n794_ & new_n800_;
  assign pk0 = ~new_n789_ | ~new_n801_;
  assign new_n803_ = ~pa1 & ~new_n202_;
  assign new_n804_ = ~new_n205_ & new_n803_;
  assign new_n805_ = ~new_n78_ & ~new_n199_;
  assign new_n806_ = ~pc0 & new_n805_;
  assign new_n807_ = new_n804_ & new_n806_;
  assign new_n808_ = ~new_n136_ & ~new_n165_;
  assign new_n809_ = ~new_n142_ & new_n808_;
  assign new_n810_ = ~new_n162_ & ~new_n191_;
  assign new_n811_ = ~new_n188_ & ~new_n197_;
  assign new_n812_ = new_n810_ & new_n811_;
  assign new_n813_ = new_n809_ & new_n812_;
  assign new_n814_ = new_n807_ & new_n813_;
  assign new_n815_ = ~pb0 & ~pz0;
  assign new_n816_ = ~new_n220_ & ~pd1;
  assign new_n817_ = new_n815_ & new_n816_;
  assign new_n818_ = ~new_n195_ & ~pb1;
  assign new_n819_ = ~new_n172_ & new_n818_;
  assign new_n820_ = new_n817_ & new_n819_;
  assign new_n821_ = ~new_n67_ & ~new_n160_;
  assign new_n822_ = ~new_n155_ & new_n821_;
  assign new_n823_ = ~new_n164_ & ~new_n168_;
  assign new_n824_ = ~new_n151_ & ~new_n179_;
  assign new_n825_ = new_n823_ & new_n824_;
  assign new_n826_ = new_n822_ & new_n825_;
  assign new_n827_ = new_n820_ & new_n826_;
  assign pl0 = ~new_n814_ | ~new_n827_;
  assign new_n829_ = ~new_n101_ & ~new_n214_;
  assign new_n830_ = ~new_n93_ & ~new_n220_;
  assign new_n831_ = ~new_n106_ & new_n830_;
  assign new_n832_ = new_n829_ & new_n831_;
  assign new_n833_ = ~new_n162_ & ~new_n172_;
  assign new_n834_ = ~new_n142_ & ~new_n160_;
  assign new_n835_ = ~new_n188_ & new_n834_;
  assign new_n836_ = new_n833_ & new_n835_;
  assign new_n837_ = new_n832_ & new_n836_;
  assign new_n838_ = ~new_n147_ & ~new_n155_;
  assign new_n839_ = ~new_n168_ & ~new_n197_;
  assign new_n840_ = ~new_n175_ & new_n839_;
  assign new_n841_ = new_n838_ & new_n840_;
  assign new_n842_ = ~new_n88_ & ~new_n208_;
  assign new_n843_ = ~new_n185_ & ~new_n196_;
  assign new_n844_ = ~new_n199_ & new_n843_;
  assign new_n845_ = new_n842_ & new_n844_;
  assign new_n846_ = new_n841_ & new_n845_;
  assign pm0 = ~new_n837_ | ~new_n846_;
  assign new_n848_ = ~new_n191_ & ~pb1;
  assign new_n849_ = new_n811_ & new_n848_;
  assign new_n850_ = ~new_n93_ & ~pz0;
  assign new_n851_ = ~pb0 & ~pd1;
  assign new_n852_ = new_n850_ & new_n851_;
  assign new_n853_ = new_n849_ & new_n852_;
  assign new_n854_ = ~new_n164_ & ~new_n172_;
  assign new_n855_ = ~new_n168_ & ~new_n195_;
  assign new_n856_ = new_n854_ & new_n855_;
  assign new_n857_ = ~new_n78_ & ~new_n136_;
  assign new_n858_ = ~new_n142_ & new_n857_;
  assign new_n859_ = new_n856_ & new_n858_;
  assign new_n860_ = new_n853_ & new_n859_;
  assign new_n861_ = ~pa1 & ~new_n208_;
  assign new_n862_ = ~new_n205_ & new_n861_;
  assign new_n863_ = ~pc0 & ~new_n88_;
  assign new_n864_ = ~new_n165_ & ~new_n179_;
  assign new_n865_ = new_n863_ & new_n864_;
  assign new_n866_ = new_n862_ & new_n865_;
  assign new_n867_ = ~new_n147_ & ~new_n175_;
  assign new_n868_ = ~new_n202_ & new_n867_;
  assign new_n869_ = ~new_n151_ & ~new_n185_;
  assign new_n870_ = new_n821_ & new_n869_;
  assign new_n871_ = new_n868_ & new_n870_;
  assign new_n872_ = new_n866_ & new_n871_;
  assign pn0 = ~new_n860_ | ~new_n872_;
  assign new_n874_ = ~new_n284_ & ~new_n302_;
  assign new_n875_ = ~new_n267_ & new_n874_;
  assign new_n876_ = ~new_n101_ & ~new_n306_;
  assign new_n877_ = ~pb1 & new_n876_;
  assign new_n878_ = new_n875_ & new_n877_;
  assign new_n879_ = ~new_n67_ & ~new_n294_;
  assign new_n880_ = ~new_n78_ & new_n879_;
  assign new_n881_ = ~new_n106_ & ~new_n179_;
  assign new_n882_ = ~new_n164_ & ~new_n214_;
  assign new_n883_ = new_n881_ & new_n882_;
  assign new_n884_ = new_n880_ & new_n883_;
  assign new_n885_ = new_n878_ & new_n884_;
  assign new_n886_ = ~new_n125_ & ~new_n279_;
  assign new_n887_ = new_n746_ & new_n886_;
  assign new_n888_ = ~new_n292_ & ~new_n297_;
  assign new_n889_ = ~new_n191_ & new_n888_;
  assign new_n890_ = new_n887_ & new_n889_;
  assign new_n891_ = ~new_n162_ & ~pz0;
  assign new_n892_ = ~new_n338_ & new_n891_;
  assign new_n893_ = ~pb0 & ~new_n220_;
  assign new_n894_ = ~new_n165_ & ~new_n195_;
  assign new_n895_ = new_n893_ & new_n894_;
  assign new_n896_ = new_n892_ & new_n895_;
  assign new_n897_ = new_n890_ & new_n896_;
  assign po0 = ~new_n885_ | ~new_n897_;
  assign new_n899_ = ~new_n350_ & new_n527_;
  assign new_n900_ = ~new_n208_ & new_n617_;
  assign new_n901_ = new_n899_ & new_n900_;
  assign new_n902_ = ~new_n160_ & ~new_n185_;
  assign new_n903_ = ~new_n136_ & new_n902_;
  assign new_n904_ = ~new_n172_ & ~new_n197_;
  assign new_n905_ = new_n244_ & new_n904_;
  assign new_n906_ = new_n903_ & new_n905_;
  assign new_n907_ = new_n901_ & new_n906_;
  assign new_n908_ = ~new_n151_ & ~new_n458_;
  assign new_n909_ = ~new_n147_ & new_n908_;
  assign new_n910_ = ~new_n142_ & ~new_n175_;
  assign new_n911_ = ~new_n188_ & new_n910_;
  assign new_n912_ = new_n909_ & new_n911_;
  assign new_n913_ = ~new_n549_ & ~new_n570_;
  assign new_n914_ = ~new_n558_ & ~new_n564_;
  assign new_n915_ = new_n913_ & new_n914_;
  assign new_n916_ = ~new_n168_ & ~new_n457_;
  assign new_n917_ = ~new_n179_ & new_n916_;
  assign new_n918_ = new_n915_ & new_n917_;
  assign new_n919_ = new_n912_ & new_n918_;
  assign pp0 = ~new_n907_ | ~new_n919_;
  assign new_n921_ = ~new_n205_ & ~new_n458_;
  assign new_n922_ = new_n527_ & new_n921_;
  assign new_n923_ = new_n915_ & new_n922_;
  assign new_n924_ = ~new_n155_ & ~new_n188_;
  assign new_n925_ = ~new_n151_ & ~new_n165_;
  assign new_n926_ = new_n924_ & new_n925_;
  assign new_n927_ = ~new_n172_ & ~new_n195_;
  assign new_n928_ = ~new_n168_ & ~new_n191_;
  assign new_n929_ = ~new_n343_ & new_n928_;
  assign new_n930_ = new_n927_ & new_n929_;
  assign new_n931_ = new_n926_ & new_n930_;
  assign new_n932_ = new_n923_ & new_n931_;
  assign new_n933_ = ~new_n162_ & ~new_n202_;
  assign new_n934_ = ~pc0 & ~new_n197_;
  assign new_n935_ = new_n933_ & new_n934_;
  assign new_n936_ = new_n229_ & new_n902_;
  assign new_n937_ = new_n935_ & new_n936_;
  assign new_n938_ = ~new_n78_ & ~new_n142_;
  assign new_n939_ = new_n248_ & new_n938_;
  assign new_n940_ = ~pb0 & ~new_n457_;
  assign new_n941_ = ~new_n116_ & new_n940_;
  assign new_n942_ = new_n231_ & new_n941_;
  assign new_n943_ = new_n939_ & new_n942_;
  assign new_n944_ = new_n937_ & new_n943_;
  assign pq0 = ~new_n932_ | ~new_n944_;
  assign new_n946_ = ~new_n208_ & ~new_n526_;
  assign new_n947_ = ~new_n205_ & new_n946_;
  assign new_n948_ = ~new_n202_ & ~new_n525_;
  assign new_n949_ = ~new_n350_ & new_n948_;
  assign new_n950_ = new_n947_ & new_n949_;
  assign new_n951_ = ~new_n165_ & ~new_n343_;
  assign new_n952_ = ~new_n147_ & new_n951_;
  assign new_n953_ = ~pc0 & ~new_n142_;
  assign new_n954_ = ~new_n175_ & new_n953_;
  assign new_n955_ = new_n952_ & new_n954_;
  assign new_n956_ = new_n950_ & new_n955_;
  assign new_n957_ = ~new_n155_ & new_n829_;
  assign new_n958_ = ~new_n106_ & new_n940_;
  assign new_n959_ = new_n957_ & new_n958_;
  assign new_n960_ = ~new_n162_ & ~new_n197_;
  assign new_n961_ = ~new_n179_ & new_n960_;
  assign new_n962_ = ~new_n172_ & ~new_n196_;
  assign new_n963_ = ~new_n188_ & new_n962_;
  assign new_n964_ = new_n961_ & new_n963_;
  assign new_n965_ = new_n959_ & new_n964_;
  assign pr0 = ~new_n956_ | ~new_n965_;
  assign new_n967_ = ~new_n132_ & ~new_n188_;
  assign new_n968_ = new_n908_ & new_n967_;
  assign new_n969_ = ~new_n457_ & ~new_n549_;
  assign new_n970_ = new_n388_ & new_n969_;
  assign new_n971_ = new_n968_ & new_n970_;
  assign new_n972_ = ~new_n78_ & new_n786_;
  assign new_n973_ = new_n785_ & new_n972_;
  assign new_n974_ = new_n971_ & new_n973_;
  assign new_n975_ = ~new_n526_ & ~new_n570_;
  assign new_n976_ = ~new_n564_ & new_n975_;
  assign new_n977_ = ~new_n168_ & ~new_n525_;
  assign new_n978_ = ~new_n350_ & ~new_n558_;
  assign new_n979_ = new_n977_ & new_n978_;
  assign new_n980_ = new_n976_ & new_n979_;
  assign new_n981_ = ~new_n175_ & ~new_n176_;
  assign new_n982_ = new_n902_ & new_n981_;
  assign new_n983_ = ~new_n179_ & ~new_n208_;
  assign new_n984_ = new_n229_ & new_n983_;
  assign new_n985_ = new_n982_ & new_n984_;
  assign new_n986_ = new_n980_ & new_n985_;
  assign ps0 = ~new_n974_ | ~new_n986_;
  assign new_n988_ = new_n231_ & ~new_n458_;
  assign new_n989_ = new_n233_ & new_n988_;
  assign new_n990_ = ~new_n162_ & ~new_n195_;
  assign new_n991_ = ~new_n168_ & new_n990_;
  assign new_n992_ = ~new_n191_ & ~new_n343_;
  assign new_n993_ = ~new_n165_ & new_n992_;
  assign new_n994_ = new_n991_ & new_n993_;
  assign new_n995_ = new_n989_ & new_n994_;
  assign new_n996_ = ~new_n160_ & new_n617_;
  assign new_n997_ = ~new_n164_ & ~new_n564_;
  assign new_n998_ = ~new_n558_ & new_n997_;
  assign new_n999_ = new_n996_ & new_n998_;
  assign new_n1000_ = ~pb0 & ~new_n214_;
  assign new_n1001_ = ~new_n220_ & ~new_n570_;
  assign new_n1002_ = ~new_n549_ & new_n1001_;
  assign new_n1003_ = new_n1000_ & new_n1002_;
  assign new_n1004_ = new_n999_ & new_n1003_;
  assign pt0 = ~new_n995_ | ~new_n1004_;
  assign new_n1006_ = ~new_n195_ & new_n811_;
  assign new_n1007_ = ~new_n191_ & new_n738_;
  assign new_n1008_ = new_n1006_ & new_n1007_;
  assign new_n1009_ = ~new_n220_ & ~new_n350_;
  assign new_n1010_ = new_n388_ & new_n1009_;
  assign new_n1011_ = ~new_n132_ & ~new_n179_;
  assign new_n1012_ = ~new_n175_ & new_n1011_;
  assign new_n1013_ = new_n1010_ & new_n1012_;
  assign new_n1014_ = new_n1008_ & new_n1013_;
  assign new_n1015_ = ~new_n78_ & new_n371_;
  assign new_n1016_ = ~new_n176_ & ~new_n208_;
  assign new_n1017_ = ~new_n199_ & new_n1016_;
  assign new_n1018_ = new_n1015_ & new_n1017_;
  assign new_n1019_ = ~new_n160_ & new_n778_;
  assign new_n1020_ = ~new_n168_ & ~new_n172_;
  assign new_n1021_ = ~new_n164_ & new_n1020_;
  assign new_n1022_ = new_n1019_ & new_n1021_;
  assign new_n1023_ = new_n1018_ & new_n1022_;
  assign pu0 = ~new_n1014_ | ~new_n1023_;
  assign new_n1025_ = ~new_n185_ & ~new_n343_;
  assign new_n1026_ = ~new_n78_ & new_n1025_;
  assign new_n1027_ = new_n527_ & new_n1026_;
  assign new_n1028_ = ~new_n188_ & ~new_n458_;
  assign new_n1029_ = ~new_n162_ & ~new_n175_;
  assign new_n1030_ = ~new_n67_ & new_n1029_;
  assign new_n1031_ = new_n1028_ & new_n1030_;
  assign new_n1032_ = new_n1027_ & new_n1031_;
  assign new_n1033_ = ~new_n136_ & ~new_n160_;
  assign new_n1034_ = ~new_n151_ & new_n1033_;
  assign new_n1035_ = new_n838_ & new_n1034_;
  assign new_n1036_ = ~new_n457_ & ~new_n570_;
  assign new_n1037_ = ~new_n142_ & new_n1036_;
  assign new_n1038_ = ~new_n549_ & new_n914_;
  assign new_n1039_ = new_n1037_ & new_n1038_;
  assign new_n1040_ = new_n1035_ & new_n1039_;
  assign pv0 = ~new_n1032_ | ~new_n1040_;
  assign new_n1042_ = ~new_n195_ & ~new_n197_;
  assign new_n1043_ = ~new_n172_ & ~new_n191_;
  assign new_n1044_ = new_n1042_ & new_n1043_;
  assign new_n1045_ = ~new_n196_ & ~new_n343_;
  assign new_n1046_ = ~new_n106_ & new_n1045_;
  assign new_n1047_ = new_n829_ & new_n1046_;
  assign pw0 = ~new_n1044_ | ~new_n1047_;
  assign new_n1049_ = new_n610_ & new_n621_;
  assign new_n1050_ = ~new_n196_ & ~new_n350_;
  assign new_n1051_ = ~new_n191_ & ~new_n525_;
  assign new_n1052_ = new_n1050_ & new_n1051_;
  assign new_n1053_ = new_n1049_ & new_n1052_;
  assign new_n1054_ = ~new_n172_ & ~new_n458_;
  assign new_n1055_ = new_n1042_ & new_n1054_;
  assign new_n1056_ = ~new_n106_ & new_n969_;
  assign new_n1057_ = new_n829_ & new_n1056_;
  assign new_n1058_ = new_n1055_ & new_n1057_;
  assign px0 = ~new_n1053_ | ~new_n1058_;
  assign new_n1060_ = ~pc0 & ~new_n205_;
  assign new_n1061_ = ~new_n558_ & new_n1060_;
  assign new_n1062_ = new_n976_ & new_n1061_;
  assign new_n1063_ = ~new_n185_ & ~new_n458_;
  assign new_n1064_ = ~new_n147_ & new_n1063_;
  assign new_n1065_ = ~new_n151_ & ~new_n525_;
  assign new_n1066_ = ~new_n136_ & new_n1065_;
  assign new_n1067_ = new_n1064_ & new_n1066_;
  assign new_n1068_ = new_n1062_ & new_n1067_;
  assign new_n1069_ = ~new_n162_ & new_n829_;
  assign new_n1070_ = new_n1056_ & new_n1069_;
  assign new_n1071_ = ~new_n175_ & new_n1042_;
  assign new_n1072_ = ~new_n172_ & ~new_n202_;
  assign new_n1073_ = ~new_n191_ & new_n1072_;
  assign new_n1074_ = new_n1071_ & new_n1073_;
  assign new_n1075_ = new_n1070_ & new_n1074_;
  assign py0 = ~new_n1068_ | ~new_n1075_;
  assign pw = pt;
  assign px = pt;
endmodule

