module top ( 
    p_127gat_18_, p_155gat_22_, p_120gat_17_, p_64gat_9_, p_106gat_15_,
    p_204gat_29_, p_1gat_0_, p_43gat_6_, p_85gat_12_, p_141gat_20_,
    p_183gat_26_, p_57gat_8_, p_148gat_21_, p_169gat_24_, p_225gat_32_,
    p_99gat_14_, p_230gat_37_, p_134gat_19_, p_162gat_23_, p_29gat_4_,
    p_78gat_11_, p_226gat_33_, p_22gat_3_, p_231gat_38_, p_36gat_5_,
    p_113gat_16_, p_8gat_1_, p_50gat_7_, p_227gat_34_, p_92gat_13_,
    p_197gat_28_, p_232gat_39_, p_233gat_40_, p_71gat_10_, p_190gat_27_,
    p_15gat_2_, p_228gat_35_, p_176gat_25_, p_218gat_31_, p_211gat_30_,
    p_229gat_36_,
    p_1332gat_585_, p_1331gat_572_, p_1334gat_577_, p_1354gat_562_,
    p_1352gat_570_, p_1336gat_586_, p_1330gat_576_, p_1335gat_573_,
    p_1353gat_566_, p_1329gat_580_, p_1328gat_584_, p_1342gat_559_,
    p_1351gat_557_, p_1333gat_581_, p_1349gat_565_, p_1350gat_561_,
    p_1348gat_569_, p_1347gat_556_, p_1341gat_563_, p_1325gat_579_,
    p_1326gat_575_, p_1344gat_568_, p_1324gat_583_, p_1343gat_555_,
    p_1345gat_564_, p_1337gat_582_, p_1327gat_571_, p_1340gat_567_,
    p_1346gat_560_, p_1339gat_574_, p_1355gat_558_, p_1338gat_578_  );
  input  p_127gat_18_, p_155gat_22_, p_120gat_17_, p_64gat_9_,
    p_106gat_15_, p_204gat_29_, p_1gat_0_, p_43gat_6_, p_85gat_12_,
    p_141gat_20_, p_183gat_26_, p_57gat_8_, p_148gat_21_, p_169gat_24_,
    p_225gat_32_, p_99gat_14_, p_230gat_37_, p_134gat_19_, p_162gat_23_,
    p_29gat_4_, p_78gat_11_, p_226gat_33_, p_22gat_3_, p_231gat_38_,
    p_36gat_5_, p_113gat_16_, p_8gat_1_, p_50gat_7_, p_227gat_34_,
    p_92gat_13_, p_197gat_28_, p_232gat_39_, p_233gat_40_, p_71gat_10_,
    p_190gat_27_, p_15gat_2_, p_228gat_35_, p_176gat_25_, p_218gat_31_,
    p_211gat_30_, p_229gat_36_;
  output p_1332gat_585_, p_1331gat_572_, p_1334gat_577_, p_1354gat_562_,
    p_1352gat_570_, p_1336gat_586_, p_1330gat_576_, p_1335gat_573_,
    p_1353gat_566_, p_1329gat_580_, p_1328gat_584_, p_1342gat_559_,
    p_1351gat_557_, p_1333gat_581_, p_1349gat_565_, p_1350gat_561_,
    p_1348gat_569_, p_1347gat_556_, p_1341gat_563_, p_1325gat_579_,
    p_1326gat_575_, p_1344gat_568_, p_1324gat_583_, p_1343gat_555_,
    p_1345gat_564_, p_1337gat_582_, p_1327gat_571_, p_1340gat_567_,
    p_1346gat_560_, p_1339gat_574_, p_1355gat_558_, p_1338gat_578_;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n453_, new_n454_, new_n455_, new_n456_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n581_, new_n582_,
    new_n583_, new_n584_;
  assign new_n74_ = p_106gat_15_ & p_99gat_14_;
  assign new_n75_ = p_106gat_15_ & ~new_n74_;
  assign new_n76_ = p_99gat_14_ & ~new_n74_;
  assign new_n77_ = ~new_n75_ & ~new_n76_;
  assign new_n78_ = p_85gat_12_ & p_92gat_13_;
  assign new_n79_ = p_92gat_13_ & ~new_n78_;
  assign new_n80_ = p_85gat_12_ & ~new_n78_;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = ~new_n77_ & ~new_n81_;
  assign new_n83_ = ~new_n77_ & ~new_n82_;
  assign new_n84_ = ~new_n81_ & ~new_n82_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = p_43gat_6_ & p_50gat_7_;
  assign new_n87_ = p_50gat_7_ & ~new_n86_;
  assign new_n88_ = p_43gat_6_ & ~new_n86_;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = p_29gat_4_ & p_36gat_5_;
  assign new_n91_ = p_36gat_5_ & ~new_n90_;
  assign new_n92_ = p_29gat_4_ & ~new_n90_;
  assign new_n93_ = ~new_n91_ & ~new_n92_;
  assign new_n94_ = ~new_n89_ & ~new_n93_;
  assign new_n95_ = ~new_n89_ & ~new_n94_;
  assign new_n96_ = ~new_n93_ & ~new_n94_;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~new_n85_ & ~new_n97_;
  assign new_n99_ = ~new_n85_ & ~new_n98_;
  assign new_n100_ = ~new_n97_ & ~new_n98_;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign new_n102_ = p_232gat_39_ & p_233gat_40_;
  assign new_n103_ = ~new_n101_ & new_n102_;
  assign new_n104_ = ~new_n101_ & ~new_n103_;
  assign new_n105_ = new_n102_ & ~new_n103_;
  assign new_n106_ = ~new_n104_ & ~new_n105_;
  assign new_n107_ = p_190gat_27_ & p_218gat_31_;
  assign new_n108_ = p_218gat_31_ & ~new_n107_;
  assign new_n109_ = p_190gat_27_ & ~new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = p_134gat_19_ & p_162gat_23_;
  assign new_n112_ = p_162gat_23_ & ~new_n111_;
  assign new_n113_ = p_134gat_19_ & ~new_n111_;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = ~new_n110_ & ~new_n114_;
  assign new_n116_ = ~new_n110_ & ~new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n115_;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = ~new_n106_ & ~new_n118_;
  assign new_n120_ = ~new_n106_ & ~new_n119_;
  assign new_n121_ = ~new_n118_ & ~new_n119_;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign new_n123_ = p_218gat_31_ & p_211gat_30_;
  assign new_n124_ = p_218gat_31_ & ~new_n123_;
  assign new_n125_ = p_211gat_30_ & ~new_n123_;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = p_204gat_29_ & p_197gat_28_;
  assign new_n128_ = p_204gat_29_ & ~new_n127_;
  assign new_n129_ = p_197gat_28_ & ~new_n127_;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = ~new_n126_ & ~new_n130_;
  assign new_n132_ = ~new_n126_ & ~new_n131_;
  assign new_n133_ = ~new_n130_ & ~new_n131_;
  assign new_n134_ = ~new_n132_ & ~new_n133_;
  assign new_n135_ = p_155gat_22_ & p_162gat_23_;
  assign new_n136_ = p_162gat_23_ & ~new_n135_;
  assign new_n137_ = p_155gat_22_ & ~new_n135_;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = p_141gat_20_ & p_148gat_21_;
  assign new_n140_ = p_148gat_21_ & ~new_n139_;
  assign new_n141_ = p_141gat_20_ & ~new_n139_;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign new_n143_ = ~new_n138_ & ~new_n142_;
  assign new_n144_ = ~new_n138_ & ~new_n143_;
  assign new_n145_ = ~new_n142_ & ~new_n143_;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~new_n134_ & ~new_n146_;
  assign new_n148_ = ~new_n134_ & ~new_n147_;
  assign new_n149_ = ~new_n146_ & ~new_n147_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = p_233gat_40_ & p_228gat_35_;
  assign new_n152_ = ~new_n150_ & new_n151_;
  assign new_n153_ = ~new_n150_ & ~new_n152_;
  assign new_n154_ = new_n151_ & ~new_n152_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = p_106gat_15_ & p_78gat_11_;
  assign new_n157_ = p_106gat_15_ & ~new_n156_;
  assign new_n158_ = p_78gat_11_ & ~new_n156_;
  assign new_n159_ = ~new_n157_ & ~new_n158_;
  assign new_n160_ = p_22gat_3_ & p_50gat_7_;
  assign new_n161_ = p_50gat_7_ & ~new_n160_;
  assign new_n162_ = p_22gat_3_ & ~new_n160_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = ~new_n159_ & ~new_n163_;
  assign new_n165_ = ~new_n159_ & ~new_n164_;
  assign new_n166_ = ~new_n163_ & ~new_n164_;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = ~new_n155_ & ~new_n167_;
  assign new_n169_ = ~new_n155_ & ~new_n168_;
  assign new_n170_ = ~new_n167_ & ~new_n168_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = p_183gat_26_ & p_190gat_27_;
  assign new_n173_ = p_190gat_27_ & ~new_n172_;
  assign new_n174_ = p_183gat_26_ & ~new_n172_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = p_169gat_24_ & p_176gat_25_;
  assign new_n177_ = p_176gat_25_ & ~new_n176_;
  assign new_n178_ = p_169gat_24_ & ~new_n176_;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = ~new_n175_ & ~new_n179_;
  assign new_n181_ = ~new_n175_ & ~new_n180_;
  assign new_n182_ = ~new_n179_ & ~new_n180_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = ~new_n134_ & ~new_n183_;
  assign new_n185_ = ~new_n134_ & ~new_n184_;
  assign new_n186_ = ~new_n183_ & ~new_n184_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = p_226gat_33_ & p_233gat_40_;
  assign new_n189_ = ~new_n187_ & new_n188_;
  assign new_n190_ = ~new_n187_ & ~new_n189_;
  assign new_n191_ = new_n188_ & ~new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = p_64gat_9_ & p_92gat_13_;
  assign new_n194_ = p_92gat_13_ & ~new_n193_;
  assign new_n195_ = p_64gat_9_ & ~new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = p_36gat_5_ & p_8gat_1_;
  assign new_n198_ = p_36gat_5_ & ~new_n197_;
  assign new_n199_ = p_8gat_1_ & ~new_n197_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = ~new_n196_ & ~new_n200_;
  assign new_n202_ = ~new_n196_ & ~new_n201_;
  assign new_n203_ = ~new_n200_ & ~new_n201_;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = ~new_n192_ & ~new_n204_;
  assign new_n206_ = ~new_n192_ & ~new_n205_;
  assign new_n207_ = ~new_n204_ & ~new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = p_127gat_18_ & p_134gat_19_;
  assign new_n210_ = p_134gat_19_ & ~new_n209_;
  assign new_n211_ = p_127gat_18_ & ~new_n209_;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign new_n213_ = p_120gat_17_ & p_113gat_16_;
  assign new_n214_ = p_120gat_17_ & ~new_n213_;
  assign new_n215_ = p_113gat_16_ & ~new_n213_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~new_n212_ & ~new_n216_;
  assign new_n218_ = ~new_n212_ & ~new_n217_;
  assign new_n219_ = ~new_n216_ & ~new_n217_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~new_n183_ & ~new_n220_;
  assign new_n222_ = ~new_n183_ & ~new_n221_;
  assign new_n223_ = ~new_n220_ & ~new_n221_;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = p_227gat_34_ & p_233gat_40_;
  assign new_n226_ = ~new_n224_ & new_n225_;
  assign new_n227_ = ~new_n224_ & ~new_n226_;
  assign new_n228_ = new_n225_ & ~new_n226_;
  assign new_n229_ = ~new_n227_ & ~new_n228_;
  assign new_n230_ = p_99gat_14_ & p_71gat_10_;
  assign new_n231_ = p_99gat_14_ & ~new_n230_;
  assign new_n232_ = p_71gat_10_ & ~new_n230_;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = p_43gat_6_ & p_15gat_2_;
  assign new_n235_ = p_43gat_6_ & ~new_n234_;
  assign new_n236_ = p_15gat_2_ & ~new_n234_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign new_n238_ = ~new_n233_ & ~new_n237_;
  assign new_n239_ = ~new_n233_ & ~new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n238_;
  assign new_n241_ = ~new_n239_ & ~new_n240_;
  assign new_n242_ = ~new_n229_ & ~new_n241_;
  assign new_n243_ = ~new_n229_ & ~new_n242_;
  assign new_n244_ = ~new_n241_ & ~new_n242_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = ~new_n146_ & ~new_n220_;
  assign new_n247_ = ~new_n146_ & ~new_n246_;
  assign new_n248_ = ~new_n220_ & ~new_n246_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = p_225gat_32_ & p_233gat_40_;
  assign new_n251_ = ~new_n249_ & new_n250_;
  assign new_n252_ = ~new_n249_ & ~new_n251_;
  assign new_n253_ = new_n250_ & ~new_n251_;
  assign new_n254_ = ~new_n252_ & ~new_n253_;
  assign new_n255_ = p_85gat_12_ & p_57gat_8_;
  assign new_n256_ = p_85gat_12_ & ~new_n255_;
  assign new_n257_ = p_57gat_8_ & ~new_n255_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = p_1gat_0_ & p_29gat_4_;
  assign new_n260_ = p_29gat_4_ & ~new_n259_;
  assign new_n261_ = p_1gat_0_ & ~new_n259_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = ~new_n258_ & ~new_n262_;
  assign new_n264_ = ~new_n258_ & ~new_n263_;
  assign new_n265_ = ~new_n262_ & ~new_n263_;
  assign new_n266_ = ~new_n264_ & ~new_n265_;
  assign new_n267_ = ~new_n254_ & ~new_n266_;
  assign new_n268_ = ~new_n254_ & ~new_n267_;
  assign new_n269_ = ~new_n266_ & ~new_n267_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = new_n171_ & new_n208_;
  assign new_n272_ = new_n245_ & new_n271_;
  assign new_n273_ = ~new_n270_ & new_n272_;
  assign new_n274_ = ~new_n245_ & new_n271_;
  assign new_n275_ = new_n270_ & new_n274_;
  assign new_n276_ = new_n171_ & ~new_n208_;
  assign new_n277_ = new_n245_ & new_n276_;
  assign new_n278_ = new_n270_ & new_n277_;
  assign new_n279_ = ~new_n171_ & new_n208_;
  assign new_n280_ = new_n245_ & new_n279_;
  assign new_n281_ = new_n270_ & new_n280_;
  assign new_n282_ = ~new_n273_ & ~new_n275_;
  assign new_n283_ = ~new_n278_ & new_n282_;
  assign new_n284_ = ~new_n281_ & new_n283_;
  assign new_n285_ = p_78gat_11_ & p_71gat_10_;
  assign new_n286_ = p_78gat_11_ & ~new_n285_;
  assign new_n287_ = p_71gat_10_ & ~new_n285_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = p_64gat_9_ & p_57gat_8_;
  assign new_n290_ = p_64gat_9_ & ~new_n289_;
  assign new_n291_ = p_57gat_8_ & ~new_n289_;
  assign new_n292_ = ~new_n290_ & ~new_n291_;
  assign new_n293_ = ~new_n288_ & ~new_n292_;
  assign new_n294_ = ~new_n288_ & ~new_n293_;
  assign new_n295_ = ~new_n292_ & ~new_n293_;
  assign new_n296_ = ~new_n294_ & ~new_n295_;
  assign new_n297_ = ~new_n85_ & ~new_n296_;
  assign new_n298_ = ~new_n85_ & ~new_n297_;
  assign new_n299_ = ~new_n296_ & ~new_n297_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = p_230gat_37_ & p_233gat_40_;
  assign new_n302_ = ~new_n300_ & new_n301_;
  assign new_n303_ = ~new_n300_ & ~new_n302_;
  assign new_n304_ = new_n301_ & ~new_n302_;
  assign new_n305_ = ~new_n303_ & ~new_n304_;
  assign new_n306_ = p_204gat_29_ & p_176gat_25_;
  assign new_n307_ = p_204gat_29_ & ~new_n306_;
  assign new_n308_ = p_176gat_25_ & ~new_n306_;
  assign new_n309_ = ~new_n307_ & ~new_n308_;
  assign new_n310_ = p_120gat_17_ & p_148gat_21_;
  assign new_n311_ = p_148gat_21_ & ~new_n310_;
  assign new_n312_ = p_120gat_17_ & ~new_n310_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign new_n314_ = ~new_n309_ & ~new_n313_;
  assign new_n315_ = ~new_n309_ & ~new_n314_;
  assign new_n316_ = ~new_n313_ & ~new_n314_;
  assign new_n317_ = ~new_n315_ & ~new_n316_;
  assign new_n318_ = ~new_n305_ & ~new_n317_;
  assign new_n319_ = ~new_n305_ & ~new_n318_;
  assign new_n320_ = ~new_n317_ & ~new_n318_;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = p_22gat_3_ & p_15gat_2_;
  assign new_n323_ = p_22gat_3_ & ~new_n322_;
  assign new_n324_ = p_15gat_2_ & ~new_n322_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = p_1gat_0_ & p_8gat_1_;
  assign new_n327_ = p_8gat_1_ & ~new_n326_;
  assign new_n328_ = p_1gat_0_ & ~new_n326_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~new_n325_ & ~new_n329_;
  assign new_n331_ = ~new_n325_ & ~new_n330_;
  assign new_n332_ = ~new_n329_ & ~new_n330_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_ = ~new_n296_ & ~new_n333_;
  assign new_n335_ = ~new_n296_ & ~new_n334_;
  assign new_n336_ = ~new_n333_ & ~new_n334_;
  assign new_n337_ = ~new_n335_ & ~new_n336_;
  assign new_n338_ = p_231gat_38_ & p_233gat_40_;
  assign new_n339_ = ~new_n337_ & new_n338_;
  assign new_n340_ = ~new_n337_ & ~new_n339_;
  assign new_n341_ = new_n338_ & ~new_n339_;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_ = p_183gat_26_ & p_211gat_30_;
  assign new_n344_ = p_211gat_30_ & ~new_n343_;
  assign new_n345_ = p_183gat_26_ & ~new_n343_;
  assign new_n346_ = ~new_n344_ & ~new_n345_;
  assign new_n347_ = p_127gat_18_ & p_155gat_22_;
  assign new_n348_ = p_155gat_22_ & ~new_n347_;
  assign new_n349_ = p_127gat_18_ & ~new_n347_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = ~new_n346_ & ~new_n350_;
  assign new_n352_ = ~new_n346_ & ~new_n351_;
  assign new_n353_ = ~new_n350_ & ~new_n351_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = ~new_n342_ & ~new_n354_;
  assign new_n356_ = ~new_n342_ & ~new_n355_;
  assign new_n357_ = ~new_n354_ & ~new_n355_;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = ~new_n97_ & ~new_n333_;
  assign new_n360_ = ~new_n97_ & ~new_n359_;
  assign new_n361_ = ~new_n333_ & ~new_n359_;
  assign new_n362_ = ~new_n360_ & ~new_n361_;
  assign new_n363_ = p_233gat_40_ & p_229gat_36_;
  assign new_n364_ = ~new_n362_ & new_n363_;
  assign new_n365_ = ~new_n362_ & ~new_n364_;
  assign new_n366_ = new_n363_ & ~new_n364_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = p_169gat_24_ & p_197gat_28_;
  assign new_n369_ = p_197gat_28_ & ~new_n368_;
  assign new_n370_ = p_169gat_24_ & ~new_n368_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = p_141gat_20_ & p_113gat_16_;
  assign new_n373_ = p_141gat_20_ & ~new_n372_;
  assign new_n374_ = p_113gat_16_ & ~new_n372_;
  assign new_n375_ = ~new_n373_ & ~new_n374_;
  assign new_n376_ = ~new_n371_ & ~new_n375_;
  assign new_n377_ = ~new_n371_ & ~new_n376_;
  assign new_n378_ = ~new_n375_ & ~new_n376_;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = ~new_n367_ & ~new_n379_;
  assign new_n381_ = ~new_n367_ & ~new_n380_;
  assign new_n382_ = ~new_n379_ & ~new_n380_;
  assign new_n383_ = ~new_n381_ & ~new_n382_;
  assign new_n384_ = new_n122_ & ~new_n284_;
  assign new_n385_ = ~new_n321_ & new_n384_;
  assign new_n386_ = ~new_n358_ & new_n385_;
  assign new_n387_ = new_n383_ & new_n386_;
  assign new_n388_ = ~new_n270_ & new_n387_;
  assign new_n389_ = p_57gat_8_ & new_n388_;
  assign new_n390_ = new_n388_ & ~new_n389_;
  assign new_n391_ = p_57gat_8_ & ~new_n389_;
  assign p_1332gat_585_ = new_n390_ | new_n391_;
  assign new_n393_ = ~new_n122_ & ~new_n284_;
  assign new_n394_ = new_n321_ & new_n393_;
  assign new_n395_ = new_n358_ & new_n394_;
  assign new_n396_ = ~new_n383_ & new_n395_;
  assign new_n397_ = ~new_n171_ & new_n396_;
  assign new_n398_ = p_50gat_7_ & new_n397_;
  assign new_n399_ = new_n397_ & ~new_n398_;
  assign new_n400_ = p_50gat_7_ & ~new_n398_;
  assign p_1331gat_572_ = new_n399_ | new_n400_;
  assign new_n402_ = ~new_n245_ & new_n387_;
  assign new_n403_ = p_71gat_10_ & new_n402_;
  assign new_n404_ = new_n402_ & ~new_n403_;
  assign new_n405_ = p_71gat_10_ & ~new_n403_;
  assign p_1334gat_577_ = new_n404_ | new_n405_;
  assign new_n407_ = new_n122_ & new_n321_;
  assign new_n408_ = new_n358_ & new_n407_;
  assign new_n409_ = ~new_n383_ & new_n408_;
  assign new_n410_ = ~new_n358_ & new_n407_;
  assign new_n411_ = new_n383_ & new_n410_;
  assign new_n412_ = new_n122_ & ~new_n321_;
  assign new_n413_ = new_n358_ & new_n412_;
  assign new_n414_ = new_n383_ & new_n413_;
  assign new_n415_ = ~new_n122_ & new_n321_;
  assign new_n416_ = new_n358_ & new_n415_;
  assign new_n417_ = new_n383_ & new_n416_;
  assign new_n418_ = ~new_n409_ & ~new_n411_;
  assign new_n419_ = ~new_n414_ & new_n418_;
  assign new_n420_ = ~new_n417_ & new_n419_;
  assign new_n421_ = ~new_n171_ & ~new_n420_;
  assign new_n422_ = ~new_n208_ & new_n421_;
  assign new_n423_ = new_n245_ & new_n422_;
  assign new_n424_ = new_n270_ & new_n423_;
  assign new_n425_ = ~new_n358_ & new_n424_;
  assign new_n426_ = p_211gat_30_ & new_n425_;
  assign new_n427_ = new_n425_ & ~new_n426_;
  assign new_n428_ = p_211gat_30_ & ~new_n426_;
  assign p_1354gat_562_ = new_n427_ | new_n428_;
  assign new_n430_ = ~new_n383_ & new_n424_;
  assign new_n431_ = p_197gat_28_ & new_n430_;
  assign new_n432_ = new_n430_ & ~new_n431_;
  assign new_n433_ = p_197gat_28_ & ~new_n431_;
  assign p_1352gat_570_ = new_n432_ | new_n433_;
  assign new_n435_ = ~new_n321_ & new_n393_;
  assign new_n436_ = new_n358_ & new_n435_;
  assign new_n437_ = new_n383_ & new_n436_;
  assign new_n438_ = ~new_n270_ & new_n437_;
  assign new_n439_ = p_85gat_12_ & new_n438_;
  assign new_n440_ = new_n438_ & ~new_n439_;
  assign new_n441_ = p_85gat_12_ & ~new_n439_;
  assign p_1336gat_586_ = new_n440_ | new_n441_;
  assign new_n443_ = ~new_n245_ & new_n396_;
  assign new_n444_ = p_43gat_6_ & new_n443_;
  assign new_n445_ = new_n443_ & ~new_n444_;
  assign new_n446_ = p_43gat_6_ & ~new_n444_;
  assign p_1330gat_576_ = new_n445_ | new_n446_;
  assign new_n448_ = ~new_n171_ & new_n387_;
  assign new_n449_ = p_78gat_11_ & new_n448_;
  assign new_n450_ = new_n448_ & ~new_n449_;
  assign new_n451_ = p_78gat_11_ & ~new_n449_;
  assign p_1335gat_573_ = new_n450_ | new_n451_;
  assign new_n453_ = ~new_n321_ & new_n424_;
  assign new_n454_ = p_204gat_29_ & new_n453_;
  assign new_n455_ = new_n453_ & ~new_n454_;
  assign new_n456_ = p_204gat_29_ & ~new_n454_;
  assign p_1353gat_566_ = new_n455_ | new_n456_;
  assign new_n458_ = ~new_n208_ & new_n396_;
  assign new_n459_ = p_36gat_5_ & new_n458_;
  assign new_n460_ = new_n458_ & ~new_n459_;
  assign new_n461_ = p_36gat_5_ & ~new_n459_;
  assign p_1329gat_580_ = new_n460_ | new_n461_;
  assign new_n463_ = ~new_n270_ & new_n396_;
  assign new_n464_ = p_29gat_4_ & new_n463_;
  assign new_n465_ = new_n463_ & ~new_n464_;
  assign new_n466_ = p_29gat_4_ & ~new_n464_;
  assign p_1328gat_584_ = new_n465_ | new_n466_;
  assign new_n468_ = new_n171_ & ~new_n420_;
  assign new_n469_ = new_n208_ & new_n468_;
  assign new_n470_ = ~new_n245_ & new_n469_;
  assign new_n471_ = ~new_n270_ & new_n470_;
  assign new_n472_ = ~new_n358_ & new_n471_;
  assign new_n473_ = p_127gat_18_ & new_n472_;
  assign new_n474_ = new_n472_ & ~new_n473_;
  assign new_n475_ = p_127gat_18_ & ~new_n473_;
  assign p_1342gat_559_ = new_n474_ | new_n475_;
  assign new_n477_ = ~new_n208_ & new_n468_;
  assign new_n478_ = ~new_n245_ & new_n477_;
  assign new_n479_ = new_n270_ & new_n478_;
  assign new_n480_ = ~new_n122_ & new_n479_;
  assign new_n481_ = p_190gat_27_ & new_n480_;
  assign new_n482_ = new_n480_ & ~new_n481_;
  assign new_n483_ = p_190gat_27_ & ~new_n481_;
  assign p_1351gat_557_ = new_n482_ | new_n483_;
  assign new_n485_ = ~new_n208_ & new_n387_;
  assign new_n486_ = p_64gat_9_ & new_n485_;
  assign new_n487_ = new_n485_ & ~new_n486_;
  assign new_n488_ = p_64gat_9_ & ~new_n486_;
  assign p_1333gat_581_ = new_n487_ | new_n488_;
  assign new_n490_ = ~new_n321_ & new_n479_;
  assign new_n491_ = p_176gat_25_ & new_n490_;
  assign new_n492_ = new_n490_ & ~new_n491_;
  assign new_n493_ = p_176gat_25_ & ~new_n491_;
  assign p_1349gat_565_ = new_n492_ | new_n493_;
  assign new_n495_ = ~new_n358_ & new_n479_;
  assign new_n496_ = p_183gat_26_ & new_n495_;
  assign new_n497_ = new_n495_ & ~new_n496_;
  assign new_n498_ = p_183gat_26_ & ~new_n496_;
  assign p_1350gat_561_ = new_n497_ | new_n498_;
  assign new_n500_ = ~new_n383_ & new_n479_;
  assign new_n501_ = p_169gat_24_ & new_n500_;
  assign new_n502_ = new_n500_ & ~new_n501_;
  assign new_n503_ = p_169gat_24_ & ~new_n501_;
  assign p_1348gat_569_ = new_n502_ | new_n503_;
  assign new_n505_ = new_n208_ & new_n421_;
  assign new_n506_ = new_n245_ & new_n505_;
  assign new_n507_ = ~new_n270_ & new_n506_;
  assign new_n508_ = ~new_n122_ & new_n507_;
  assign new_n509_ = p_162gat_23_ & new_n508_;
  assign new_n510_ = new_n508_ & ~new_n509_;
  assign new_n511_ = p_162gat_23_ & ~new_n509_;
  assign p_1347gat_556_ = new_n510_ | new_n511_;
  assign new_n513_ = ~new_n321_ & new_n471_;
  assign new_n514_ = p_120gat_17_ & new_n513_;
  assign new_n515_ = new_n513_ & ~new_n514_;
  assign new_n516_ = p_120gat_17_ & ~new_n514_;
  assign p_1341gat_563_ = new_n515_ | new_n516_;
  assign new_n518_ = new_n321_ & new_n384_;
  assign new_n519_ = ~new_n358_ & new_n518_;
  assign new_n520_ = ~new_n383_ & new_n519_;
  assign new_n521_ = ~new_n208_ & new_n520_;
  assign new_n522_ = p_8gat_1_ & new_n521_;
  assign new_n523_ = new_n521_ & ~new_n522_;
  assign new_n524_ = p_8gat_1_ & ~new_n522_;
  assign p_1325gat_579_ = new_n523_ | new_n524_;
  assign new_n526_ = ~new_n245_ & new_n520_;
  assign new_n527_ = p_15gat_2_ & new_n526_;
  assign new_n528_ = new_n526_ & ~new_n527_;
  assign new_n529_ = p_15gat_2_ & ~new_n527_;
  assign p_1326gat_575_ = new_n528_ | new_n529_;
  assign new_n531_ = ~new_n383_ & new_n507_;
  assign new_n532_ = p_141gat_20_ & new_n531_;
  assign new_n533_ = new_n531_ & ~new_n532_;
  assign new_n534_ = p_141gat_20_ & ~new_n532_;
  assign p_1344gat_568_ = new_n533_ | new_n534_;
  assign new_n536_ = ~new_n270_ & new_n520_;
  assign new_n537_ = p_1gat_0_ & new_n536_;
  assign new_n538_ = new_n536_ & ~new_n537_;
  assign new_n539_ = p_1gat_0_ & ~new_n537_;
  assign p_1324gat_583_ = new_n538_ | new_n539_;
  assign new_n541_ = ~new_n122_ & new_n471_;
  assign new_n542_ = p_134gat_19_ & new_n541_;
  assign new_n543_ = new_n541_ & ~new_n542_;
  assign new_n544_ = p_134gat_19_ & ~new_n542_;
  assign p_1343gat_555_ = new_n543_ | new_n544_;
  assign new_n546_ = ~new_n321_ & new_n507_;
  assign new_n547_ = p_148gat_21_ & new_n546_;
  assign new_n548_ = new_n546_ & ~new_n547_;
  assign new_n549_ = p_148gat_21_ & ~new_n547_;
  assign p_1345gat_564_ = new_n548_ | new_n549_;
  assign new_n551_ = ~new_n208_ & new_n437_;
  assign new_n552_ = p_92gat_13_ & new_n551_;
  assign new_n553_ = new_n551_ & ~new_n552_;
  assign new_n554_ = p_92gat_13_ & ~new_n552_;
  assign p_1337gat_582_ = new_n553_ | new_n554_;
  assign new_n556_ = ~new_n171_ & new_n520_;
  assign new_n557_ = p_22gat_3_ & new_n556_;
  assign new_n558_ = new_n556_ & ~new_n557_;
  assign new_n559_ = p_22gat_3_ & ~new_n557_;
  assign p_1327gat_571_ = new_n558_ | new_n559_;
  assign new_n561_ = ~new_n383_ & new_n471_;
  assign new_n562_ = p_113gat_16_ & new_n561_;
  assign new_n563_ = new_n561_ & ~new_n562_;
  assign new_n564_ = p_113gat_16_ & ~new_n562_;
  assign p_1340gat_567_ = new_n563_ | new_n564_;
  assign new_n566_ = ~new_n358_ & new_n507_;
  assign new_n567_ = p_155gat_22_ & new_n566_;
  assign new_n568_ = new_n566_ & ~new_n567_;
  assign new_n569_ = p_155gat_22_ & ~new_n567_;
  assign p_1346gat_560_ = new_n568_ | new_n569_;
  assign new_n571_ = ~new_n171_ & new_n437_;
  assign new_n572_ = p_106gat_15_ & new_n571_;
  assign new_n573_ = new_n571_ & ~new_n572_;
  assign new_n574_ = p_106gat_15_ & ~new_n572_;
  assign p_1339gat_574_ = new_n573_ | new_n574_;
  assign new_n576_ = ~new_n122_ & new_n424_;
  assign new_n577_ = p_218gat_31_ & new_n576_;
  assign new_n578_ = new_n576_ & ~new_n577_;
  assign new_n579_ = p_218gat_31_ & ~new_n577_;
  assign p_1355gat_558_ = new_n578_ | new_n579_;
  assign new_n581_ = ~new_n245_ & new_n437_;
  assign new_n582_ = p_99gat_14_ & new_n581_;
  assign new_n583_ = new_n581_ & ~new_n582_;
  assign new_n584_ = p_99gat_14_ & ~new_n582_;
  assign p_1338gat_578_ = new_n583_ | new_n584_;
endmodule

