module top ( 
    pdel1, pratr, pbull1, pbull0, pwatch, povacc, pverr_n, porwd_n,
    pvlenesr, pmmerr, paccrpy, pvacc, pcat4, pvst1, pcapsd, pcat3, pcat2,
    pcat1, plsd, pvst0, pcat0, pibt2, pkbg_n, pmarssr, pend, pvsumesr,
    pbull5, ppluto4, pstar2, pbull4, ppluto5, ppy, pstar3, pbull3,
    pcomppar, pibt1, pstar0, pbull2, pibt0, pstar1, ppluto0, pfbi, powl_n,
    ppluto1, piclr, ppluto2, pbull6, pcat5, ppluto3,
    pbull2_p, pend_p, pbull3_p, porwd_f, pbull4_p, ppluto3_p, pwatch_p,
    pbull5_p, pbull6_p, ppluto5_p, ppy_p, ppluto4_p, plsd_p, pvlenesr_p,
    pfbi_p, pstar1_p, pvsumesr_p, paccrpy_p, pkbg_f, pmarssr_p, pstar0_p,
    pstar3_p, pdel1_p, pstar2_p, pvst0_p, pcomppar_p, powl_f, psdo,
    pvst1_p, ppluto1_p, pratr_p, ppluto0_p, povacc_p, ppluto2_p, pbull0_p,
    pverr_f, pbull1_p  );
  input  pdel1, pratr, pbull1, pbull0, pwatch, povacc, pverr_n, porwd_n,
    pvlenesr, pmmerr, paccrpy, pvacc, pcat4, pvst1, pcapsd, pcat3, pcat2,
    pcat1, plsd, pvst0, pcat0, pibt2, pkbg_n, pmarssr, pend, pvsumesr,
    pbull5, ppluto4, pstar2, pbull4, ppluto5, ppy, pstar3, pbull3,
    pcomppar, pibt1, pstar0, pbull2, pibt0, pstar1, ppluto0, pfbi, powl_n,
    ppluto1, piclr, ppluto2, pbull6, pcat5, ppluto3;
  output pbull2_p, pend_p, pbull3_p, porwd_f, pbull4_p, ppluto3_p, pwatch_p,
    pbull5_p, pbull6_p, ppluto5_p, ppy_p, ppluto4_p, plsd_p, pvlenesr_p,
    pfbi_p, pstar1_p, pvsumesr_p, paccrpy_p, pkbg_f, pmarssr_p, pstar0_p,
    pstar3_p, pdel1_p, pstar2_p, pvst0_p, pcomppar_p, powl_f, psdo,
    pvst1_p, ppluto1_p, pratr_p, ppluto0_p, povacc_p, ppluto2_p, pbull0_p,
    pverr_f, pbull1_p;
  wire new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n166_,
    new_n167_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n196_, new_n197_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n220_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n256_, new_n258_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n274_, new_n276_,
    new_n277_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n298_,
    new_n299_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n308_, new_n309_, new_n310_, new_n311_, new_n313_,
    new_n314_, new_n316_, new_n317_, new_n318_, new_n320_, new_n321_,
    new_n323_, new_n324_, new_n327_, new_n328_, new_n330_, new_n331_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n342_, new_n343_, new_n344_;
  assign new_n87_ = pwatch & powl_n;
  assign new_n88_ = ~pbull2 & new_n87_;
  assign new_n89_ = pbull0 & new_n88_;
  assign new_n90_ = pbull1 & new_n89_;
  assign new_n91_ = ~pbull1 & powl_n;
  assign new_n92_ = ~pwatch & powl_n;
  assign new_n93_ = ~pbull0 & powl_n;
  assign new_n94_ = ~new_n91_ & ~new_n92_;
  assign new_n95_ = ~new_n93_ & new_n94_;
  assign new_n96_ = pbull2 & ~new_n95_;
  assign pbull2_p = new_n90_ | new_n96_;
  assign new_n98_ = pfbi & powl_n;
  assign new_n99_ = pstar0 & pstar1;
  assign new_n100_ = ~pstar2 & new_n99_;
  assign new_n101_ = new_n98_ & ~new_n100_;
  assign new_n102_ = pibt2 & ~pibt0;
  assign new_n103_ = pibt1 & new_n102_;
  assign new_n104_ = ~pcat4 & new_n103_;
  assign new_n105_ = pibt2 & pibt0;
  assign new_n106_ = ~pibt1 & new_n105_;
  assign new_n107_ = ~pcat3 & new_n106_;
  assign new_n108_ = ~pibt2 & pibt1;
  assign new_n109_ = ~pcat0 & new_n108_;
  assign new_n110_ = ~pibt0 & new_n109_;
  assign new_n111_ = pibt1 & new_n105_;
  assign new_n112_ = ~pcat5 & new_n111_;
  assign new_n113_ = pibt0 & new_n108_;
  assign new_n114_ = ~pcat1 & new_n113_;
  assign new_n115_ = ~pibt1 & new_n102_;
  assign new_n116_ = ~pcat2 & new_n115_;
  assign new_n117_ = ~new_n104_ & ~new_n107_;
  assign new_n118_ = ~new_n110_ & new_n117_;
  assign new_n119_ = ~new_n112_ & ~new_n114_;
  assign new_n120_ = ~new_n116_ & new_n119_;
  assign new_n121_ = new_n118_ & new_n120_;
  assign porwd_f = ~pwatch | new_n121_;
  assign new_n123_ = new_n98_ & ~porwd_f;
  assign new_n124_ = ~new_n101_ & ~new_n123_;
  assign new_n125_ = new_n98_ & new_n124_;
  assign new_n126_ = pend & powl_n;
  assign pend_p = new_n125_ | new_n126_;
  assign new_n128_ = pbull0 & pbull2;
  assign new_n129_ = pbull1 & pwatch;
  assign new_n130_ = new_n128_ & new_n129_;
  assign new_n131_ = ~pbull3 & new_n130_;
  assign new_n132_ = powl_n & new_n131_;
  assign new_n133_ = pbull3 & ~new_n130_;
  assign new_n134_ = powl_n & new_n133_;
  assign pbull3_p = new_n132_ | new_n134_;
  assign new_n136_ = ~pbull3 & powl_n;
  assign new_n137_ = pbull4 & new_n136_;
  assign new_n138_ = powl_n & ~new_n130_;
  assign new_n139_ = pbull4 & new_n138_;
  assign new_n140_ = pbull3 & new_n130_;
  assign new_n141_ = powl_n & new_n140_;
  assign new_n142_ = ~pbull4 & new_n141_;
  assign new_n143_ = ~new_n137_ & ~new_n139_;
  assign pbull4_p = new_n142_ | ~new_n143_;
  assign new_n145_ = pvst1 & new_n126_;
  assign new_n146_ = ~pkbg_n & powl_n;
  assign new_n147_ = ~pbull5 & pbull6;
  assign new_n148_ = ~pbull3 & new_n147_;
  assign new_n149_ = pbull4 & new_n148_;
  assign new_n150_ = ~pbull0 & new_n149_;
  assign new_n151_ = pbull1 & new_n150_;
  assign new_n152_ = ~pbull2 & new_n151_;
  assign new_n153_ = new_n87_ & new_n152_;
  assign new_n154_ = ~pcomppar & new_n126_;
  assign new_n155_ = ~pvst0 & new_n126_;
  assign new_n156_ = ~pmmerr & new_n155_;
  assign new_n157_ = ~new_n145_ & ~new_n146_;
  assign new_n158_ = ~new_n153_ & new_n157_;
  assign new_n159_ = ~new_n154_ & ~new_n156_;
  assign new_n160_ = new_n158_ & new_n159_;
  assign new_n161_ = pibt0 & ~new_n160_;
  assign new_n162_ = pibt2 & new_n161_;
  assign new_n163_ = ~pibt1 & new_n162_;
  assign new_n164_ = powl_n & ppluto3;
  assign ppluto3_p = new_n163_ | new_n164_;
  assign new_n166_ = povacc & powl_n;
  assign new_n167_ = ~pvacc & new_n166_;
  assign pwatch_p = new_n87_ | new_n167_;
  assign new_n169_ = pbull5 & new_n138_;
  assign new_n170_ = pbull4 & new_n141_;
  assign new_n171_ = ~pbull5 & new_n170_;
  assign new_n172_ = pbull5 & new_n136_;
  assign new_n173_ = pbull5 & pbull4_p;
  assign new_n174_ = ~new_n169_ & ~new_n171_;
  assign new_n175_ = ~new_n172_ & ~new_n173_;
  assign pbull5_p = ~new_n174_ | ~new_n175_;
  assign new_n177_ = powl_n & pbull6;
  assign new_n178_ = ~pbull4 & new_n177_;
  assign new_n179_ = ~pbull5 & new_n177_;
  assign new_n180_ = ~pbull2 & new_n177_;
  assign new_n181_ = ~pbull3 & new_n177_;
  assign new_n182_ = pbull6 & ~new_n95_;
  assign new_n183_ = pbull5 & new_n141_;
  assign new_n184_ = ~pbull6 & new_n183_;
  assign new_n185_ = pbull4 & new_n184_;
  assign new_n186_ = ~new_n95_ & new_n130_;
  assign new_n187_ = pbull4 & new_n186_;
  assign new_n188_ = pbull5 & new_n187_;
  assign new_n189_ = pbull3 & new_n188_;
  assign new_n190_ = ~new_n178_ & ~new_n179_;
  assign new_n191_ = ~new_n180_ & ~new_n181_;
  assign new_n192_ = new_n190_ & new_n191_;
  assign new_n193_ = ~new_n182_ & ~new_n185_;
  assign new_n194_ = ~new_n189_ & new_n193_;
  assign pbull6_p = ~new_n192_ | ~new_n194_;
  assign new_n196_ = pibt1 & new_n162_;
  assign new_n197_ = ppluto5 & powl_n;
  assign ppluto5_p = new_n196_ | new_n197_;
  assign new_n199_ = pfbi & ~piclr;
  assign new_n200_ = pdel1 & new_n199_;
  assign new_n201_ = ~pfbi & ~piclr;
  assign new_n202_ = ppy & new_n201_;
  assign ppy_p = new_n200_ | new_n202_;
  assign new_n204_ = ~pibt0 & ~new_n160_;
  assign new_n205_ = pibt2 & new_n204_;
  assign new_n206_ = pibt1 & new_n205_;
  assign new_n207_ = ppluto4 & powl_n;
  assign ppluto4_p = new_n206_ | new_n207_;
  assign new_n209_ = new_n87_ & ~new_n121_;
  assign new_n210_ = ~pstar3 & new_n209_;
  assign new_n211_ = new_n100_ & new_n210_;
  assign new_n212_ = pfbi & new_n211_;
  assign new_n213_ = plsd & powl_n;
  assign new_n214_ = ~pstar3 & new_n213_;
  assign new_n215_ = ~new_n100_ & new_n213_;
  assign new_n216_ = ~pfbi & new_n213_;
  assign new_n217_ = ~new_n212_ & ~new_n214_;
  assign new_n218_ = ~new_n215_ & ~new_n216_;
  assign plsd_p = ~new_n217_ | ~new_n218_;
  assign new_n220_ = pvlenesr & powl_n;
  assign pvlenesr_p = new_n146_ | new_n220_;
  assign new_n222_ = ~porwd_n & new_n101_;
  assign new_n223_ = pfbi & new_n101_;
  assign new_n224_ = ~porwd_n & new_n209_;
  assign new_n225_ = ~new_n98_ & ~new_n224_;
  assign new_n226_ = new_n209_ & ~new_n225_;
  assign new_n227_ = ~porwd_n & new_n226_;
  assign new_n228_ = ~new_n99_ & new_n226_;
  assign new_n229_ = pfbi & new_n209_;
  assign new_n230_ = powl_n & ~new_n99_;
  assign new_n231_ = ~new_n100_ & new_n230_;
  assign new_n232_ = pstar2 & new_n231_;
  assign new_n233_ = new_n224_ & new_n232_;
  assign new_n234_ = ~new_n99_ & new_n101_;
  assign new_n235_ = pfbi & new_n232_;
  assign new_n236_ = ~new_n222_ & ~new_n223_;
  assign new_n237_ = ~new_n227_ & ~new_n228_;
  assign new_n238_ = new_n236_ & new_n237_;
  assign new_n239_ = ~new_n234_ & ~new_n235_;
  assign new_n240_ = ~new_n229_ & ~new_n233_;
  assign new_n241_ = new_n239_ & new_n240_;
  assign pfbi_p = ~new_n238_ | ~new_n241_;
  assign new_n243_ = new_n98_ & ~new_n99_;
  assign new_n244_ = pstar0 & new_n243_;
  assign new_n245_ = ~pstar1 & new_n224_;
  assign new_n246_ = pstar0 & new_n245_;
  assign new_n247_ = pstar1 & new_n230_;
  assign new_n248_ = ~pstar0 & new_n247_;
  assign new_n249_ = ~porwd_n & ~porwd_f;
  assign new_n250_ = ~pfbi & ~new_n249_;
  assign new_n251_ = powl_n & new_n250_;
  assign new_n252_ = pstar1 & new_n251_;
  assign new_n253_ = ~new_n244_ & ~new_n246_;
  assign new_n254_ = ~new_n248_ & ~new_n252_;
  assign pstar1_p = ~new_n253_ | ~new_n254_;
  assign new_n256_ = pvsumesr & powl_n;
  assign pvsumesr_p = new_n145_ | new_n256_;
  assign new_n258_ = paccrpy & powl_n;
  assign paccrpy_p = new_n125_ | new_n258_;
  assign new_n260_ = ~pcat1 & new_n109_;
  assign new_n261_ = pwatch & new_n260_;
  assign new_n262_ = ~new_n100_ & new_n261_;
  assign new_n263_ = ~new_n100_ & ~porwd_f;
  assign new_n264_ = ~pstar3 & new_n261_;
  assign new_n265_ = ~pstar3 & ~porwd_f;
  assign new_n266_ = ~new_n262_ & ~new_n263_;
  assign new_n267_ = ~new_n264_ & ~new_n265_;
  assign new_n268_ = new_n266_ & new_n267_;
  assign new_n269_ = pkbg_n & ~new_n268_;
  assign new_n270_ = ~powl_n & ~new_n98_;
  assign new_n271_ = pkbg_n & new_n124_;
  assign new_n272_ = ~new_n269_ & ~new_n270_;
  assign pkbg_f = new_n271_ | ~new_n272_;
  assign new_n274_ = pmarssr & powl_n;
  assign pmarssr_p = new_n153_ | new_n274_;
  assign new_n276_ = pstar0 & new_n251_;
  assign new_n277_ = ~pstar0 & ~new_n225_;
  assign pstar0_p = new_n276_ | new_n277_;
  assign new_n279_ = ~pstar3 & new_n99_;
  assign new_n280_ = ~new_n225_ & new_n279_;
  assign new_n281_ = pstar2 & new_n280_;
  assign new_n282_ = pstar3 & new_n230_;
  assign new_n283_ = ~pstar2 & pstar3;
  assign new_n284_ = powl_n & new_n283_;
  assign new_n285_ = pstar3 & new_n251_;
  assign new_n286_ = ~new_n281_ & ~new_n282_;
  assign new_n287_ = ~new_n284_ & ~new_n285_;
  assign pstar3_p = ~new_n286_ | ~new_n287_;
  assign pdel1_p = pcapsd & ~piclr;
  assign new_n290_ = new_n98_ & new_n99_;
  assign new_n291_ = ~pstar2 & new_n290_;
  assign new_n292_ = new_n100_ & new_n224_;
  assign new_n293_ = pstar2 & new_n230_;
  assign new_n294_ = pstar2 & new_n251_;
  assign new_n295_ = ~new_n291_ & ~new_n292_;
  assign new_n296_ = ~new_n293_ & ~new_n294_;
  assign pstar2_p = ~new_n295_ | ~new_n296_;
  assign new_n298_ = pvst1 & new_n199_;
  assign new_n299_ = pvst0 & new_n201_;
  assign pvst0_p = new_n298_ | new_n299_;
  assign new_n301_ = pcomppar & powl_n;
  assign new_n302_ = ~pfbi & new_n301_;
  assign new_n303_ = ~pdel1 & new_n301_;
  assign new_n304_ = ~pcomppar & new_n98_;
  assign new_n305_ = pdel1 & new_n304_;
  assign new_n306_ = ~new_n302_ & ~new_n303_;
  assign pcomppar_p = new_n305_ | ~new_n306_;
  assign new_n308_ = pkbg_n & ~piclr;
  assign new_n309_ = ~pend & new_n308_;
  assign new_n310_ = ~new_n152_ & new_n309_;
  assign new_n311_ = ~pwatch & new_n309_;
  assign powl_f = new_n310_ | new_n311_;
  assign new_n313_ = ppy & new_n199_;
  assign new_n314_ = pvst1 & new_n201_;
  assign pvst1_p = new_n313_ | new_n314_;
  assign new_n316_ = new_n108_ & ~new_n160_;
  assign new_n317_ = pibt0 & new_n316_;
  assign new_n318_ = powl_n & ppluto1;
  assign ppluto1_p = new_n317_ | new_n318_;
  assign new_n320_ = pratr & powl_n;
  assign new_n321_ = ~new_n154_ & ~new_n320_;
  assign pratr_p = new_n156_ | ~new_n321_;
  assign new_n323_ = ~pibt0 & new_n316_;
  assign new_n324_ = ppluto0 & powl_n;
  assign ppluto0_p = new_n323_ | new_n324_;
  assign povacc_p = pvacc & ~piclr;
  assign new_n327_ = ~pibt1 & new_n205_;
  assign new_n328_ = powl_n & ppluto2;
  assign ppluto2_p = new_n327_ | new_n328_;
  assign new_n330_ = pbull0 & new_n92_;
  assign new_n331_ = ~pbull0 & new_n87_;
  assign pbull0_p = new_n330_ | new_n331_;
  assign new_n333_ = ~new_n152_ & ~new_n268_;
  assign new_n334_ = pverr_n & new_n333_;
  assign new_n335_ = ~pwatch & new_n124_;
  assign new_n336_ = pverr_n & new_n335_;
  assign new_n337_ = new_n124_ & ~new_n152_;
  assign new_n338_ = pverr_n & new_n337_;
  assign new_n339_ = ~new_n334_ & ~new_n336_;
  assign new_n340_ = ~new_n270_ & ~new_n338_;
  assign pverr_f = ~new_n339_ | ~new_n340_;
  assign new_n342_ = pbull0 & new_n87_;
  assign new_n343_ = ~pbull1 & new_n342_;
  assign new_n344_ = pbull1 & ~new_n95_;
  assign pbull1_p = new_n343_ | new_n344_;
  assign psdo = pvst0;
endmodule

