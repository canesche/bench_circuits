module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz, ph3,
    pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2, pm3,
    pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb, pp2,
    pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1,
    pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0,
    py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl,
    pm, pn, po,
    pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz,
    ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2,
    pm3, pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb,
    pp2, pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe,
    pt1, pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph,
    px0, py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1,
    pl, pm, pn, po;
  output pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5;
  wire new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n525_,
    new_n526_, new_n527_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1161_, new_n1162_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_;
  assign new_n235_ = ~pb0 & ~pv;
  assign new_n236_ = ps & new_n235_;
  assign new_n237_ = ~pv & ~pj1;
  assign new_n238_ = pb0 & ~pj1;
  assign new_n239_ = ~ps & ~pj1;
  assign new_n240_ = ~new_n236_ & ~new_n237_;
  assign new_n241_ = ~new_n238_ & ~new_n239_;
  assign new_n242_ = new_n240_ & new_n241_;
  assign pe5 = ~py1 & new_n242_;
  assign new_n244_ = pl2 & ~pm2;
  assign new_n245_ = pn2 & new_n244_;
  assign new_n246_ = ~pe0 & ~pf0;
  assign new_n247_ = pg0 & new_n246_;
  assign new_n248_ = ~po2 & new_n245_;
  assign new_n249_ = new_n247_ & new_n248_;
  assign new_n250_ = pp2 & new_n248_;
  assign new_n251_ = ~new_n249_ & ~new_n250_;
  assign new_n252_ = ~pk2 & new_n251_;
  assign new_n253_ = pk2 & ~new_n251_;
  assign new_n254_ = ~px1 & new_n253_;
  assign new_n255_ = ~new_n252_ & ~new_n254_;
  assign new_n256_ = ~py1 & new_n255_;
  assign new_n257_ = ~px1 & new_n256_;
  assign new_n258_ = pk2 & new_n256_;
  assign pf6 = new_n257_ | new_n258_;
  assign new_n260_ = ~pk1 & pe;
  assign new_n261_ = ~pe & ~pu0;
  assign new_n262_ = pd & new_n261_;
  assign new_n263_ = pc & ~pd;
  assign new_n264_ = ~pe & new_n263_;
  assign new_n265_ = ~pv2 & new_n264_;
  assign new_n266_ = ~new_n260_ & ~new_n262_;
  assign new_n267_ = ~new_n265_ & new_n266_;
  assign new_n268_ = ~pd & ~pe;
  assign new_n269_ = ~py1 & new_n267_;
  assign new_n270_ = ~new_n268_ & new_n269_;
  assign new_n271_ = ~pk2 & pl3;
  assign new_n272_ = ~pj2 & new_n271_;
  assign new_n273_ = pl3 & px1;
  assign new_n274_ = ~new_n272_ & ~new_n273_;
  assign new_n275_ = px1 & new_n274_;
  assign new_n276_ = ~pj2 & ~pk2;
  assign new_n277_ = new_n274_ & new_n276_;
  assign new_n278_ = ~pm3 & new_n274_;
  assign new_n279_ = ~new_n275_ & ~new_n277_;
  assign new_n280_ = ~new_n278_ & new_n279_;
  assign new_n281_ = new_n269_ & new_n280_;
  assign new_n282_ = pc & new_n269_;
  assign new_n283_ = ~new_n270_ & ~new_n281_;
  assign pg7 = new_n282_ | ~new_n283_;
  assign new_n285_ = ~pb0 & ~pu;
  assign new_n286_ = ps & new_n285_;
  assign new_n287_ = ~pu & ~pi1;
  assign new_n288_ = pb0 & ~pi1;
  assign new_n289_ = ~ps & ~pi1;
  assign new_n290_ = ~new_n286_ & ~new_n287_;
  assign new_n291_ = ~new_n288_ & ~new_n289_;
  assign new_n292_ = new_n290_ & new_n291_;
  assign pd5 = ~py1 & new_n292_;
  assign new_n294_ = ~pj1 & pe;
  assign new_n295_ = ~pt0 & ~pe;
  assign new_n296_ = pd & new_n295_;
  assign new_n297_ = ~pu2 & new_n264_;
  assign new_n298_ = ~new_n294_ & ~new_n296_;
  assign new_n299_ = ~new_n297_ & new_n298_;
  assign new_n300_ = ~py1 & new_n299_;
  assign new_n301_ = ~new_n268_ & new_n300_;
  assign new_n302_ = pk3 & ~pk2;
  assign new_n303_ = ~pj2 & new_n302_;
  assign new_n304_ = pk3 & px1;
  assign new_n305_ = ~new_n303_ & ~new_n304_;
  assign new_n306_ = px1 & new_n305_;
  assign new_n307_ = new_n276_ & new_n305_;
  assign new_n308_ = ~pl3 & new_n305_;
  assign new_n309_ = ~new_n306_ & ~new_n307_;
  assign new_n310_ = ~new_n308_ & new_n309_;
  assign new_n311_ = new_n300_ & new_n310_;
  assign new_n312_ = pc & new_n300_;
  assign new_n313_ = ~new_n301_ & ~new_n311_;
  assign pf7 = new_n312_ | ~new_n313_;
  assign new_n315_ = ~pc & ~pd;
  assign new_n316_ = ~pe & new_n315_;
  assign new_n317_ = px1 & new_n316_;
  assign new_n318_ = ~pl2 & new_n317_;
  assign new_n319_ = ~pe & px1;
  assign new_n320_ = ~pc & new_n319_;
  assign new_n321_ = ~pd & new_n320_;
  assign new_n322_ = ~py1 & ~new_n318_;
  assign new_n323_ = new_n321_ & new_n322_;
  assign new_n324_ = ~pl2 & new_n322_;
  assign pg6 = new_n323_ | new_n324_;
  assign new_n326_ = po2 & new_n244_;
  assign new_n327_ = pp2 & new_n244_;
  assign new_n328_ = ~pg0 & new_n244_;
  assign new_n329_ = ~new_n326_ & ~new_n327_;
  assign new_n330_ = ~new_n328_ & new_n329_;
  assign new_n331_ = pn2 & ~new_n330_;
  assign new_n332_ = pj2 & new_n331_;
  assign new_n333_ = ~pp2 & new_n332_;
  assign new_n334_ = ~po2 & new_n331_;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = ~py1 & ~new_n335_;
  assign new_n337_ = ~px1 & new_n336_;
  assign new_n338_ = pi2 & ~py1;
  assign pd6 = new_n337_ | new_n338_;
  assign new_n340_ = ~pi1 & pe;
  assign new_n341_ = ~ps0 & ~pe;
  assign new_n342_ = pd & new_n341_;
  assign new_n343_ = ~pt2 & new_n264_;
  assign new_n344_ = ~new_n340_ & ~new_n342_;
  assign new_n345_ = ~new_n343_ & new_n344_;
  assign new_n346_ = ~py1 & new_n345_;
  assign new_n347_ = ~new_n268_ & new_n346_;
  assign new_n348_ = pj3 & ~pk2;
  assign new_n349_ = ~pj2 & new_n348_;
  assign new_n350_ = pj3 & px1;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = px1 & new_n351_;
  assign new_n353_ = new_n276_ & new_n351_;
  assign new_n354_ = ~pk3 & new_n351_;
  assign new_n355_ = ~new_n352_ & ~new_n353_;
  assign new_n356_ = ~new_n354_ & new_n355_;
  assign new_n357_ = new_n346_ & new_n356_;
  assign new_n358_ = pc & new_n346_;
  assign new_n359_ = ~new_n347_ & ~new_n357_;
  assign pe7 = new_n358_ | ~new_n359_;
  assign new_n361_ = ~pb0 & ~px;
  assign new_n362_ = ps & new_n361_;
  assign new_n363_ = ~px & ~pl1;
  assign new_n364_ = pb0 & ~pl1;
  assign new_n365_ = ~ps & ~pl1;
  assign new_n366_ = ~new_n362_ & ~new_n363_;
  assign new_n367_ = ~new_n364_ & ~new_n365_;
  assign new_n368_ = new_n366_ & new_n367_;
  assign pg5 = ~py1 & new_n368_;
  assign new_n370_ = ~ph1 & pe;
  assign new_n371_ = ~pr0 & ~pe;
  assign new_n372_ = pd & new_n371_;
  assign new_n373_ = ~ps2 & new_n264_;
  assign new_n374_ = ~new_n370_ & ~new_n372_;
  assign new_n375_ = ~new_n373_ & new_n374_;
  assign new_n376_ = ~py1 & new_n375_;
  assign new_n377_ = ~new_n268_ & new_n376_;
  assign new_n378_ = ~pk2 & pi3;
  assign new_n379_ = ~pj2 & new_n378_;
  assign new_n380_ = pi3 & px1;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = px1 & new_n381_;
  assign new_n383_ = new_n276_ & new_n381_;
  assign new_n384_ = ~pj3 & new_n381_;
  assign new_n385_ = ~new_n382_ & ~new_n383_;
  assign new_n386_ = ~new_n384_ & new_n385_;
  assign new_n387_ = new_n376_ & new_n386_;
  assign new_n388_ = pc & new_n376_;
  assign new_n389_ = ~new_n377_ & ~new_n387_;
  assign pd7 = new_n388_ | ~new_n389_;
  assign new_n391_ = ~po2 & new_n244_;
  assign new_n392_ = pj2 & new_n244_;
  assign new_n393_ = ~new_n391_ & ~new_n392_;
  assign new_n394_ = ~po2 & new_n246_;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = pn2 & new_n395_;
  assign new_n397_ = ~pp2 & new_n396_;
  assign new_n398_ = pg0 & new_n397_;
  assign new_n399_ = po2 & new_n397_;
  assign new_n400_ = ~new_n398_ & ~new_n399_;
  assign new_n401_ = ~pj2 & new_n400_;
  assign new_n402_ = pj2 & ~new_n400_;
  assign new_n403_ = ~px1 & new_n402_;
  assign new_n404_ = ~new_n401_ & ~new_n403_;
  assign new_n405_ = ~py1 & new_n404_;
  assign new_n406_ = ~px1 & new_n405_;
  assign new_n407_ = pj2 & new_n405_;
  assign pe6 = new_n406_ | new_n407_;
  assign new_n409_ = ~pb0 & ~pw;
  assign new_n410_ = ps & new_n409_;
  assign new_n411_ = ~pw & ~pk1;
  assign new_n412_ = pb0 & ~pk1;
  assign new_n413_ = ~ps & ~pk1;
  assign new_n414_ = ~new_n410_ & ~new_n411_;
  assign new_n415_ = ~new_n412_ & ~new_n413_;
  assign new_n416_ = new_n414_ & new_n415_;
  assign pf5 = ~py1 & new_n416_;
  assign new_n418_ = ~pp & pr;
  assign new_n419_ = pi & new_n418_;
  assign new_n420_ = ~pp & ~pf1;
  assign new_n421_ = ~pr & ~pf1;
  assign new_n422_ = ~pf1 & ~pi;
  assign new_n423_ = ~new_n419_ & ~new_n420_;
  assign new_n424_ = ~new_n421_ & ~new_n422_;
  assign new_n425_ = new_n423_ & new_n424_;
  assign pa5 = ~py1 & new_n425_;
  assign pb6 = ph2 & ~pn0;
  assign new_n428_ = ~ph3 & ~pf;
  assign new_n429_ = ~pg & ph;
  assign new_n430_ = pf & new_n429_;
  assign new_n431_ = ~new_n428_ & ~new_n430_;
  assign new_n432_ = ~py1 & new_n431_;
  assign new_n433_ = ph & new_n432_;
  assign new_n434_ = ph3 & new_n432_;
  assign pc7 = new_n433_ | new_n434_;
  assign new_n436_ = ~pg3 & ~pf;
  assign new_n437_ = ~ph3 & ph;
  assign new_n438_ = pf & new_n437_;
  assign new_n439_ = ~new_n436_ & ~new_n438_;
  assign new_n440_ = ~py1 & new_n439_;
  assign new_n441_ = ph & new_n440_;
  assign new_n442_ = pg3 & new_n440_;
  assign pb7 = new_n441_ | new_n442_;
  assign pc6 = pl0 & ~pn0;
  assign new_n445_ = ~pf3 & ~pf;
  assign new_n446_ = ~pg3 & ph;
  assign new_n447_ = pf & new_n446_;
  assign new_n448_ = ~new_n445_ & ~new_n447_;
  assign new_n449_ = ~py1 & new_n448_;
  assign new_n450_ = ph & new_n449_;
  assign new_n451_ = pf3 & new_n449_;
  assign pa7 = new_n450_ | new_n451_;
  assign new_n453_ = ~pb0 & ~pt;
  assign new_n454_ = ps & new_n453_;
  assign new_n455_ = ~pt & ~ph1;
  assign new_n456_ = pb0 & ~ph1;
  assign new_n457_ = ~ps & ~ph1;
  assign new_n458_ = ~new_n454_ & ~new_n455_;
  assign new_n459_ = ~new_n456_ & ~new_n457_;
  assign new_n460_ = new_n458_ & new_n459_;
  assign pc5 = ~py1 & new_n460_;
  assign new_n462_ = ~pi0 & ~pj0;
  assign new_n463_ = ~pk0 & pl0;
  assign new_n464_ = pd2 & new_n463_;
  assign new_n465_ = new_n462_ & new_n464_;
  assign new_n466_ = ~ph0 & new_n465_;
  assign new_n467_ = ~pe4 & pi0;
  assign new_n468_ = pf4 & ~pj0;
  assign new_n469_ = pf4 & ~pg4;
  assign new_n470_ = ~pk0 & new_n469_;
  assign new_n471_ = pf4 & pg4;
  assign new_n472_ = pk0 & new_n471_;
  assign new_n473_ = ~pg4 & ~pk0;
  assign new_n474_ = ~pj0 & new_n473_;
  assign new_n475_ = pg4 & pk0;
  assign new_n476_ = ~pj0 & new_n475_;
  assign new_n477_ = ~new_n470_ & ~new_n472_;
  assign new_n478_ = ~new_n474_ & ~new_n476_;
  assign new_n479_ = new_n477_ & new_n478_;
  assign new_n480_ = ~new_n467_ & ~new_n468_;
  assign new_n481_ = ~new_n479_ & new_n480_;
  assign new_n482_ = pi0 & new_n481_;
  assign new_n483_ = ~ph0 & new_n482_;
  assign new_n484_ = ~pe4 & new_n481_;
  assign new_n485_ = ~ph0 & new_n484_;
  assign new_n486_ = ~pd4 & new_n482_;
  assign new_n487_ = ~pd4 & new_n484_;
  assign new_n488_ = ~new_n483_ & ~new_n485_;
  assign new_n489_ = ~new_n486_ & ~new_n487_;
  assign new_n490_ = new_n488_ & new_n489_;
  assign new_n491_ = ~pd4 & ~ph0;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = pc4 & new_n492_;
  assign new_n494_ = pb4 & new_n493_;
  assign new_n495_ = pa4 & new_n494_;
  assign new_n496_ = pz3 & new_n495_;
  assign new_n497_ = py3 & new_n496_;
  assign new_n498_ = ph4 & new_n497_;
  assign new_n499_ = ~new_n466_ & ~new_n498_;
  assign new_n500_ = ~pa2 & pf2;
  assign new_n501_ = new_n499_ & new_n500_;
  assign new_n502_ = ~pn0 & new_n501_;
  assign new_n503_ = ~pf2 & pe2;
  assign new_n504_ = ~pa2 & ~new_n498_;
  assign new_n505_ = ~new_n462_ & new_n504_;
  assign new_n506_ = ~new_n464_ & new_n504_;
  assign new_n507_ = ph0 & new_n504_;
  assign new_n508_ = ~new_n505_ & ~new_n506_;
  assign new_n509_ = ~new_n507_ & new_n508_;
  assign new_n510_ = new_n503_ & new_n509_;
  assign new_n511_ = ~pn0 & new_n510_;
  assign new_n512_ = ~pe2 & ~pn0;
  assign new_n513_ = pf2 & new_n512_;
  assign new_n514_ = ~new_n502_ & ~new_n511_;
  assign pa6 = new_n513_ | ~new_n514_;
  assign new_n516_ = ~pq & pr;
  assign new_n517_ = pi & new_n516_;
  assign new_n518_ = ~pq & ~pg1;
  assign new_n519_ = ~pr & ~pg1;
  assign new_n520_ = ~pg1 & ~pi;
  assign new_n521_ = ~new_n517_ & ~new_n518_;
  assign new_n522_ = ~new_n519_ & ~new_n520_;
  assign new_n523_ = new_n521_ & new_n522_;
  assign pb5 = ~py1 & new_n523_;
  assign new_n525_ = pg2 & ph2;
  assign new_n526_ = ~pn0 & new_n525_;
  assign new_n527_ = pc2 & ~pn0;
  assign pl4 = new_n526_ | new_n527_;
  assign new_n529_ = pb0 & ~pv;
  assign new_n530_ = ps & new_n529_;
  assign new_n531_ = ~pv & ~pr1;
  assign new_n532_ = ~pb0 & ~pr1;
  assign new_n533_ = ~ps & ~pr1;
  assign new_n534_ = ~new_n530_ & ~new_n531_;
  assign new_n535_ = ~new_n532_ & ~new_n533_;
  assign new_n536_ = new_n534_ & new_n535_;
  assign pm5 = ~py1 & new_n536_;
  assign new_n538_ = ~ps2 & ~pf;
  assign new_n539_ = ~pt2 & ~ph;
  assign new_n540_ = pf & new_n539_;
  assign new_n541_ = ~new_n538_ & ~new_n540_;
  assign new_n542_ = ~py1 & new_n541_;
  assign new_n543_ = ~ph & new_n542_;
  assign new_n544_ = ps2 & new_n542_;
  assign pn6 = new_n543_ | new_n544_;
  assign new_n546_ = ~ps1 & pe;
  assign new_n547_ = ~pc1 & ~pe;
  assign new_n548_ = pd & new_n547_;
  assign new_n549_ = ~pd3 & new_n264_;
  assign new_n550_ = ~new_n546_ & ~new_n548_;
  assign new_n551_ = ~new_n549_ & new_n550_;
  assign new_n552_ = ~py1 & new_n551_;
  assign new_n553_ = ~new_n268_ & new_n552_;
  assign new_n554_ = ~pk2 & pt3;
  assign new_n555_ = ~pj2 & new_n554_;
  assign new_n556_ = pt3 & px1;
  assign new_n557_ = ~new_n555_ & ~new_n556_;
  assign new_n558_ = px1 & new_n557_;
  assign new_n559_ = new_n276_ & new_n557_;
  assign new_n560_ = ~pu3 & new_n557_;
  assign new_n561_ = ~new_n558_ & ~new_n559_;
  assign new_n562_ = ~new_n560_ & new_n561_;
  assign new_n563_ = new_n552_ & new_n562_;
  assign new_n564_ = pc & new_n552_;
  assign new_n565_ = ~new_n553_ & ~new_n563_;
  assign po7 = new_n564_ | ~new_n565_;
  assign new_n567_ = pa4 & pz3;
  assign new_n568_ = pb4 & new_n567_;
  assign new_n569_ = ~pd4 & pc4;
  assign new_n570_ = pe4 & new_n569_;
  assign new_n571_ = new_n568_ & new_n570_;
  assign new_n572_ = py3 & new_n571_;
  assign new_n573_ = ~pl0 & ~pn0;
  assign new_n574_ = pz3 & py3;
  assign new_n575_ = new_n572_ & new_n573_;
  assign new_n576_ = ~new_n574_ & new_n575_;
  assign new_n577_ = pa4 & pb4;
  assign new_n578_ = pc4 & new_n577_;
  assign new_n579_ = new_n575_ & ~new_n578_;
  assign new_n580_ = pf4 & new_n573_;
  assign new_n581_ = ~new_n578_ & new_n580_;
  assign new_n582_ = ~pd4 & pe4;
  assign new_n583_ = pf4 & new_n582_;
  assign new_n584_ = new_n580_ & ~new_n583_;
  assign new_n585_ = ~new_n574_ & new_n580_;
  assign new_n586_ = new_n575_ & ~new_n583_;
  assign new_n587_ = ~new_n576_ & ~new_n579_;
  assign new_n588_ = ~new_n581_ & new_n587_;
  assign new_n589_ = ~new_n584_ & ~new_n585_;
  assign new_n590_ = ~new_n586_ & new_n589_;
  assign pa8 = ~new_n588_ | ~new_n590_;
  assign new_n592_ = pb0 & ~pu;
  assign new_n593_ = ps & new_n592_;
  assign new_n594_ = ~pu & ~pq1;
  assign new_n595_ = ~pb0 & ~pq1;
  assign new_n596_ = ~ps & ~pq1;
  assign new_n597_ = ~new_n593_ & ~new_n594_;
  assign new_n598_ = ~new_n595_ & ~new_n596_;
  assign new_n599_ = new_n597_ & new_n598_;
  assign pl5 = ~py1 & new_n599_;
  assign new_n601_ = ~pr & ~pj;
  assign new_n602_ = pi & new_n601_;
  assign new_n603_ = ~pr0 & ~pj;
  assign new_n604_ = pr & ~pr0;
  assign new_n605_ = ~pr0 & ~pi;
  assign new_n606_ = ~new_n602_ & ~new_n603_;
  assign new_n607_ = ~new_n604_ & ~new_n605_;
  assign new_n608_ = new_n606_ & new_n607_;
  assign pm4 = ~py1 & new_n608_;
  assign new_n610_ = ~pr1 & pe;
  assign new_n611_ = ~pb1 & ~pe;
  assign new_n612_ = pd & new_n611_;
  assign new_n613_ = ~pc3 & new_n264_;
  assign new_n614_ = ~new_n610_ & ~new_n612_;
  assign new_n615_ = ~new_n613_ & new_n614_;
  assign new_n616_ = ~py1 & new_n615_;
  assign new_n617_ = ~new_n268_ & new_n616_;
  assign new_n618_ = ~pk2 & ps3;
  assign new_n619_ = ~pj2 & new_n618_;
  assign new_n620_ = ps3 & px1;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = px1 & new_n621_;
  assign new_n623_ = new_n276_ & new_n621_;
  assign new_n624_ = ~pt3 & new_n621_;
  assign new_n625_ = ~new_n622_ & ~new_n623_;
  assign new_n626_ = ~new_n624_ & new_n625_;
  assign new_n627_ = new_n616_ & new_n626_;
  assign new_n628_ = pc & new_n616_;
  assign new_n629_ = ~new_n617_ & ~new_n627_;
  assign pn7 = new_n628_ | ~new_n629_;
  assign new_n631_ = ~pf & ~pt2;
  assign new_n632_ = ~pu2 & ~ph;
  assign new_n633_ = pf & new_n632_;
  assign new_n634_ = ~new_n631_ & ~new_n633_;
  assign new_n635_ = ~py1 & new_n634_;
  assign new_n636_ = ~ph & new_n635_;
  assign new_n637_ = pt2 & new_n635_;
  assign po6 = new_n636_ | new_n637_;
  assign new_n639_ = new_n578_ & new_n583_;
  assign new_n640_ = new_n574_ & new_n639_;
  assign new_n641_ = pa4 & new_n574_;
  assign new_n642_ = new_n573_ & new_n640_;
  assign new_n643_ = ~new_n641_ & new_n642_;
  assign new_n644_ = pb4 & pc4;
  assign new_n645_ = ~pd4 & new_n644_;
  assign new_n646_ = new_n642_ & ~new_n645_;
  assign new_n647_ = pg4 & new_n573_;
  assign new_n648_ = ~new_n645_ & new_n647_;
  assign new_n649_ = pe4 & pf4;
  assign new_n650_ = pg4 & new_n649_;
  assign new_n651_ = new_n647_ & ~new_n650_;
  assign new_n652_ = ~new_n641_ & new_n647_;
  assign new_n653_ = new_n642_ & ~new_n650_;
  assign new_n654_ = ~new_n643_ & ~new_n646_;
  assign new_n655_ = ~new_n648_ & new_n654_;
  assign new_n656_ = ~new_n651_ & ~new_n652_;
  assign new_n657_ = ~new_n653_ & new_n656_;
  assign pb8 = ~new_n655_ | ~new_n657_;
  assign new_n659_ = ~pq2 & px1;
  assign new_n660_ = ~pq2 & new_n335_;
  assign new_n661_ = ~pi2 & new_n660_;
  assign new_n662_ = ~new_n659_ & ~new_n661_;
  assign new_n663_ = ~py1 & new_n662_;
  assign new_n664_ = px1 & new_n663_;
  assign new_n665_ = ~pi2 & new_n335_;
  assign new_n666_ = new_n663_ & new_n665_;
  assign new_n667_ = ~pq2 & new_n663_;
  assign new_n668_ = ~new_n664_ & ~new_n666_;
  assign pl6 = new_n667_ | ~new_n668_;
  assign new_n670_ = ~pq1 & pe;
  assign new_n671_ = ~pa1 & ~pe;
  assign new_n672_ = pd & new_n671_;
  assign new_n673_ = ~pb3 & new_n264_;
  assign new_n674_ = ~new_n670_ & ~new_n672_;
  assign new_n675_ = ~new_n673_ & new_n674_;
  assign new_n676_ = ~py1 & new_n675_;
  assign new_n677_ = ~new_n268_ & new_n676_;
  assign new_n678_ = ~pk2 & pr3;
  assign new_n679_ = ~pj2 & new_n678_;
  assign new_n680_ = pr3 & px1;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = px1 & new_n681_;
  assign new_n683_ = new_n276_ & new_n681_;
  assign new_n684_ = ~ps3 & new_n681_;
  assign new_n685_ = ~new_n682_ & ~new_n683_;
  assign new_n686_ = ~new_n684_ & new_n685_;
  assign new_n687_ = new_n676_ & new_n686_;
  assign new_n688_ = pc & new_n676_;
  assign new_n689_ = ~new_n677_ & ~new_n687_;
  assign pm7 = new_n688_ | ~new_n689_;
  assign new_n691_ = ~pr & ~pk;
  assign new_n692_ = pi & new_n691_;
  assign new_n693_ = ~ps0 & ~pk;
  assign new_n694_ = pr & ~ps0;
  assign new_n695_ = ~ps0 & ~pi;
  assign new_n696_ = ~new_n692_ & ~new_n693_;
  assign new_n697_ = ~new_n694_ & ~new_n695_;
  assign new_n698_ = new_n696_ & new_n697_;
  assign pn4 = ~py1 & new_n698_;
  assign new_n700_ = pb0 & ~px;
  assign new_n701_ = ps & new_n700_;
  assign new_n702_ = ~px & ~pt1;
  assign new_n703_ = ~pb0 & ~pt1;
  assign new_n704_ = ~ps & ~pt1;
  assign new_n705_ = ~new_n701_ & ~new_n702_;
  assign new_n706_ = ~new_n703_ & ~new_n704_;
  assign new_n707_ = new_n705_ & new_n706_;
  assign po5 = ~py1 & new_n707_;
  assign new_n709_ = pb & ~new_n525_;
  assign new_n710_ = ~pn0 & new_n709_;
  assign new_n711_ = pl0 & new_n710_;
  assign new_n712_ = pd2 & new_n711_;
  assign new_n713_ = ph4 & new_n710_;
  assign pc8 = new_n712_ | new_n713_;
  assign new_n715_ = ~pp1 & pe;
  assign new_n716_ = ~pe & ~pz0;
  assign new_n717_ = pd & new_n716_;
  assign new_n718_ = ~pa3 & new_n264_;
  assign new_n719_ = ~new_n715_ & ~new_n717_;
  assign new_n720_ = ~new_n718_ & new_n719_;
  assign new_n721_ = ~py1 & new_n720_;
  assign new_n722_ = ~new_n268_ & new_n721_;
  assign new_n723_ = ~pk2 & pq3;
  assign new_n724_ = ~pj2 & new_n723_;
  assign new_n725_ = pq3 & px1;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = px1 & new_n726_;
  assign new_n728_ = new_n276_ & new_n726_;
  assign new_n729_ = ~pr3 & new_n726_;
  assign new_n730_ = ~new_n727_ & ~new_n728_;
  assign new_n731_ = ~new_n729_ & new_n730_;
  assign new_n732_ = new_n721_ & new_n731_;
  assign new_n733_ = pc & new_n721_;
  assign new_n734_ = ~new_n722_ & ~new_n732_;
  assign pl7 = new_n733_ | ~new_n734_;
  assign new_n736_ = pq2 & ~new_n665_;
  assign new_n737_ = ~px1 & new_n736_;
  assign new_n738_ = ~py1 & new_n737_;
  assign new_n739_ = px1 & new_n738_;
  assign new_n740_ = pr2 & pq2;
  assign new_n741_ = new_n738_ & ~new_n740_;
  assign new_n742_ = pr2 & ~py1;
  assign new_n743_ = ~new_n740_ & new_n742_;
  assign new_n744_ = new_n665_ & new_n742_;
  assign new_n745_ = px1 & new_n742_;
  assign new_n746_ = new_n665_ & new_n738_;
  assign new_n747_ = ~new_n739_ & ~new_n741_;
  assign new_n748_ = ~new_n743_ & new_n747_;
  assign new_n749_ = ~new_n744_ & ~new_n745_;
  assign new_n750_ = ~new_n746_ & new_n749_;
  assign pm6 = ~new_n748_ | ~new_n750_;
  assign new_n752_ = pb0 & ~pw;
  assign new_n753_ = ps & new_n752_;
  assign new_n754_ = ~pw & ~ps1;
  assign new_n755_ = ~pb0 & ~ps1;
  assign new_n756_ = ~ps & ~ps1;
  assign new_n757_ = ~new_n753_ & ~new_n754_;
  assign new_n758_ = ~new_n755_ & ~new_n756_;
  assign new_n759_ = new_n757_ & new_n758_;
  assign pn5 = ~py1 & new_n759_;
  assign new_n761_ = ~pr & ~pl;
  assign new_n762_ = pi & new_n761_;
  assign new_n763_ = ~pt0 & ~pl;
  assign new_n764_ = pr & ~pt0;
  assign new_n765_ = ~pt0 & ~pi;
  assign new_n766_ = ~new_n762_ & ~new_n763_;
  assign new_n767_ = ~new_n764_ & ~new_n765_;
  assign new_n768_ = new_n766_ & new_n767_;
  assign po4 = ~py1 & new_n768_;
  assign new_n770_ = ~pb0 & ~pz;
  assign new_n771_ = ps & new_n770_;
  assign new_n772_ = ~pz & ~pn1;
  assign new_n773_ = pb0 & ~pn1;
  assign new_n774_ = ~ps & ~pn1;
  assign new_n775_ = ~new_n771_ & ~new_n772_;
  assign new_n776_ = ~new_n773_ & ~new_n774_;
  assign new_n777_ = new_n775_ & new_n776_;
  assign pi5 = ~py1 & new_n777_;
  assign new_n779_ = pl2 & pm2;
  assign new_n780_ = pn2 & new_n779_;
  assign new_n781_ = ~new_n321_ & new_n780_;
  assign new_n782_ = ~py1 & new_n781_;
  assign new_n783_ = ~pl2 & new_n782_;
  assign new_n784_ = pn2 & pm2;
  assign new_n785_ = po2 & new_n784_;
  assign new_n786_ = new_n782_ & ~new_n785_;
  assign new_n787_ = po2 & ~py1;
  assign new_n788_ = ~new_n785_ & new_n787_;
  assign new_n789_ = new_n321_ & new_n787_;
  assign new_n790_ = ~pl2 & new_n787_;
  assign new_n791_ = new_n321_ & new_n782_;
  assign new_n792_ = ~new_n783_ & ~new_n786_;
  assign new_n793_ = ~new_n788_ & new_n792_;
  assign new_n794_ = ~new_n789_ & ~new_n790_;
  assign new_n795_ = ~new_n791_ & new_n794_;
  assign pj6 = ~new_n793_ | ~new_n795_;
  assign new_n797_ = ~po1 & pe;
  assign new_n798_ = ~pe & ~py0;
  assign new_n799_ = pd & new_n798_;
  assign new_n800_ = ~pz2 & new_n264_;
  assign new_n801_ = ~new_n797_ & ~new_n799_;
  assign new_n802_ = ~new_n800_ & new_n801_;
  assign new_n803_ = ~py1 & new_n802_;
  assign new_n804_ = ~new_n268_ & new_n803_;
  assign new_n805_ = ~pk2 & pp3;
  assign new_n806_ = ~pj2 & new_n805_;
  assign new_n807_ = pp3 & px1;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = px1 & new_n808_;
  assign new_n810_ = new_n276_ & new_n808_;
  assign new_n811_ = ~pq3 & new_n808_;
  assign new_n812_ = ~new_n809_ & ~new_n810_;
  assign new_n813_ = ~new_n811_ & new_n812_;
  assign new_n814_ = new_n803_ & new_n813_;
  assign new_n815_ = pc & new_n803_;
  assign new_n816_ = ~new_n804_ & ~new_n814_;
  assign pk7 = new_n815_ | ~new_n816_;
  assign new_n818_ = ~pb0 & ~py;
  assign new_n819_ = ps & new_n818_;
  assign new_n820_ = ~py & ~pm1;
  assign new_n821_ = pb0 & ~pm1;
  assign new_n822_ = ~ps & ~pm1;
  assign new_n823_ = ~new_n819_ & ~new_n820_;
  assign new_n824_ = ~new_n821_ & ~new_n822_;
  assign new_n825_ = new_n823_ & new_n824_;
  assign ph5 = ~py1 & new_n825_;
  assign pi4 = pa2 | ~px1;
  assign new_n828_ = ~pn1 & pe;
  assign new_n829_ = ~pe & ~px0;
  assign new_n830_ = pd & new_n829_;
  assign new_n831_ = ~py2 & new_n264_;
  assign new_n832_ = ~new_n828_ & ~new_n830_;
  assign new_n833_ = ~new_n831_ & new_n832_;
  assign new_n834_ = ~py1 & new_n833_;
  assign new_n835_ = ~new_n268_ & new_n834_;
  assign new_n836_ = ~pk2 & po3;
  assign new_n837_ = ~pj2 & new_n836_;
  assign new_n838_ = po3 & px1;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = px1 & new_n839_;
  assign new_n841_ = new_n276_ & new_n839_;
  assign new_n842_ = ~pp3 & new_n839_;
  assign new_n843_ = ~new_n840_ & ~new_n841_;
  assign new_n844_ = ~new_n842_ & new_n843_;
  assign new_n845_ = new_n834_ & new_n844_;
  assign new_n846_ = pc & new_n834_;
  assign new_n847_ = ~new_n835_ & ~new_n845_;
  assign pj7 = new_n846_ | ~new_n847_;
  assign new_n849_ = ~new_n321_ & new_n785_;
  assign new_n850_ = pl2 & new_n849_;
  assign new_n851_ = ~py1 & new_n850_;
  assign new_n852_ = ~new_n779_ & new_n851_;
  assign new_n853_ = pn2 & po2;
  assign new_n854_ = pp2 & new_n853_;
  assign new_n855_ = new_n851_ & ~new_n854_;
  assign new_n856_ = pp2 & ~py1;
  assign new_n857_ = ~new_n854_ & new_n856_;
  assign new_n858_ = new_n321_ & new_n856_;
  assign new_n859_ = ~new_n779_ & new_n856_;
  assign new_n860_ = new_n321_ & new_n851_;
  assign new_n861_ = ~new_n852_ & ~new_n855_;
  assign new_n862_ = ~new_n857_ & new_n861_;
  assign new_n863_ = ~new_n858_ & ~new_n859_;
  assign new_n864_ = ~new_n860_ & new_n863_;
  assign pk6 = ~new_n862_ | ~new_n864_;
  assign new_n866_ = ~pm2 & new_n319_;
  assign new_n867_ = ~pc & new_n866_;
  assign new_n868_ = ~pd & new_n867_;
  assign new_n869_ = ~py1 & ~new_n868_;
  assign new_n870_ = new_n321_ & new_n869_;
  assign new_n871_ = pm2 & new_n870_;
  assign new_n872_ = ~pm2 & new_n869_;
  assign new_n873_ = pl2 & new_n872_;
  assign new_n874_ = pl2 & new_n870_;
  assign new_n875_ = pm2 & new_n869_;
  assign new_n876_ = ~pl2 & new_n875_;
  assign new_n877_ = ~new_n871_ & ~new_n873_;
  assign new_n878_ = ~new_n874_ & ~new_n876_;
  assign ph6 = ~new_n877_ | ~new_n878_;
  assign new_n880_ = ~pm1 & pe;
  assign new_n881_ = ~pe & ~pw0;
  assign new_n882_ = pd & new_n881_;
  assign new_n883_ = ~px2 & new_n264_;
  assign new_n884_ = ~new_n880_ & ~new_n882_;
  assign new_n885_ = ~new_n883_ & new_n884_;
  assign new_n886_ = ~py1 & new_n885_;
  assign new_n887_ = ~new_n268_ & new_n886_;
  assign new_n888_ = ~pk2 & pn3;
  assign new_n889_ = ~pj2 & new_n888_;
  assign new_n890_ = pn3 & px1;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = px1 & new_n891_;
  assign new_n893_ = new_n276_ & new_n891_;
  assign new_n894_ = ~po3 & new_n891_;
  assign new_n895_ = ~new_n892_ & ~new_n893_;
  assign new_n896_ = ~new_n894_ & new_n895_;
  assign new_n897_ = new_n886_ & new_n896_;
  assign new_n898_ = pc & new_n886_;
  assign new_n899_ = ~new_n887_ & ~new_n897_;
  assign pi7 = new_n898_ | ~new_n899_;
  assign new_n901_ = ~po0 & px1;
  assign new_n902_ = ~po0 & ~new_n740_;
  assign new_n903_ = ~pi2 & ~po0;
  assign new_n904_ = ~new_n901_ & ~new_n902_;
  assign new_n905_ = ~new_n903_ & new_n904_;
  assign new_n906_ = new_n268_ & new_n905_;
  assign new_n907_ = ~pc & new_n906_;
  assign pj4 = py1 | new_n907_;
  assign new_n909_ = pb0 & ~pt;
  assign new_n910_ = ps & new_n909_;
  assign new_n911_ = ~pt & ~pp1;
  assign new_n912_ = ~pb0 & ~pp1;
  assign new_n913_ = ~ps & ~pp1;
  assign new_n914_ = ~new_n910_ & ~new_n911_;
  assign new_n915_ = ~new_n912_ & ~new_n913_;
  assign new_n916_ = new_n914_ & new_n915_;
  assign pk5 = ~py1 & new_n916_;
  assign new_n918_ = ~pl1 & pe;
  assign new_n919_ = ~pe & ~pv0;
  assign new_n920_ = pd & new_n919_;
  assign new_n921_ = ~pw2 & new_n264_;
  assign new_n922_ = ~new_n918_ & ~new_n920_;
  assign new_n923_ = ~new_n921_ & new_n922_;
  assign new_n924_ = ~py1 & new_n923_;
  assign new_n925_ = ~new_n268_ & new_n924_;
  assign new_n926_ = ~pk2 & pm3;
  assign new_n927_ = ~pj2 & new_n926_;
  assign new_n928_ = pm3 & px1;
  assign new_n929_ = ~new_n927_ & ~new_n928_;
  assign new_n930_ = px1 & new_n929_;
  assign new_n931_ = new_n276_ & new_n929_;
  assign new_n932_ = ~pn3 & new_n929_;
  assign new_n933_ = ~new_n930_ & ~new_n931_;
  assign new_n934_ = ~new_n932_ & new_n933_;
  assign new_n935_ = new_n924_ & new_n934_;
  assign new_n936_ = pc & new_n924_;
  assign new_n937_ = ~new_n925_ & ~new_n935_;
  assign ph7 = new_n936_ | ~new_n937_;
  assign new_n939_ = ~new_n321_ & new_n779_;
  assign new_n940_ = ~py1 & new_n939_;
  assign new_n941_ = ~pl2 & new_n940_;
  assign new_n942_ = ~new_n784_ & new_n940_;
  assign new_n943_ = pn2 & ~py1;
  assign new_n944_ = ~new_n784_ & new_n943_;
  assign new_n945_ = new_n321_ & new_n943_;
  assign new_n946_ = ~pl2 & new_n943_;
  assign new_n947_ = new_n321_ & new_n940_;
  assign new_n948_ = ~new_n941_ & ~new_n942_;
  assign new_n949_ = ~new_n944_ & new_n948_;
  assign new_n950_ = ~new_n945_ & ~new_n946_;
  assign new_n951_ = ~new_n947_ & new_n950_;
  assign pi6 = ~new_n949_ | ~new_n951_;
  assign new_n953_ = ~pa0 & ~pb0;
  assign new_n954_ = ps & new_n953_;
  assign new_n955_ = ~pa0 & ~po1;
  assign new_n956_ = pb0 & ~po1;
  assign new_n957_ = ~ps & ~po1;
  assign new_n958_ = ~new_n954_ & ~new_n955_;
  assign new_n959_ = ~new_n956_ & ~new_n957_;
  assign new_n960_ = new_n958_ & new_n959_;
  assign pj5 = ~py1 & new_n960_;
  assign new_n962_ = ~pa2 & ~pj2;
  assign new_n963_ = ~pk2 & new_n962_;
  assign new_n964_ = pi2 & pq2;
  assign new_n965_ = pi2 & pr2;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = ~pk0 & ~pl2;
  assign new_n968_ = ~pj0 & ~pk0;
  assign new_n969_ = ~pj0 & pl2;
  assign new_n970_ = ~new_n967_ & ~new_n968_;
  assign new_n971_ = ~pn2 & ~new_n969_;
  assign new_n972_ = new_n970_ & new_n971_;
  assign new_n973_ = ~po2 & ~pp2;
  assign new_n974_ = new_n972_ & new_n973_;
  assign new_n975_ = pm2 & new_n974_;
  assign new_n976_ = ~pi0 & ~pl2;
  assign new_n977_ = ~ph0 & ~pi0;
  assign new_n978_ = ~ph0 & pl2;
  assign new_n979_ = ~new_n976_ & ~new_n977_;
  assign new_n980_ = pn2 & ~new_n978_;
  assign new_n981_ = new_n979_ & new_n980_;
  assign new_n982_ = new_n974_ & new_n981_;
  assign new_n983_ = new_n973_ & new_n981_;
  assign new_n984_ = ~pm2 & new_n983_;
  assign new_n985_ = ~new_n975_ & ~new_n982_;
  assign new_n986_ = ~new_n984_ & new_n985_;
  assign new_n987_ = ~py1 & ~new_n986_;
  assign new_n988_ = new_n963_ & new_n966_;
  assign new_n989_ = new_n987_ & new_n988_;
  assign new_n990_ = ~pa2 & ~py1;
  assign new_n991_ = pd0 & new_n965_;
  assign new_n992_ = pi3 & pr2;
  assign new_n993_ = pd0 & new_n992_;
  assign new_n994_ = pi3 & ~pi2;
  assign new_n995_ = pi3 & pq2;
  assign new_n996_ = ~new_n991_ & ~new_n993_;
  assign new_n997_ = ~new_n994_ & new_n996_;
  assign new_n998_ = ~new_n964_ & ~new_n995_;
  assign new_n999_ = new_n997_ & new_n998_;
  assign new_n1000_ = pr2 & new_n999_;
  assign new_n1001_ = ~pi3 & new_n999_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~pi2 & new_n1002_;
  assign new_n1004_ = pk2 & new_n1003_;
  assign new_n1005_ = pj2 & new_n1003_;
  assign new_n1006_ = ~pq2 & new_n1002_;
  assign new_n1007_ = pj2 & new_n1006_;
  assign new_n1008_ = ~pr2 & ~pq2;
  assign new_n1009_ = pi2 & ~new_n1008_;
  assign new_n1010_ = new_n1006_ & new_n1009_;
  assign new_n1011_ = pk2 & new_n1006_;
  assign new_n1012_ = pr2 & pz1;
  assign new_n1013_ = pc0 & ~pr2;
  assign new_n1014_ = pc0 & pz1;
  assign new_n1015_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1016_ = ~new_n1014_ & new_n1015_;
  assign new_n1017_ = new_n1002_ & new_n1016_;
  assign new_n1018_ = pj2 & new_n1017_;
  assign new_n1019_ = new_n1009_ & new_n1017_;
  assign new_n1020_ = new_n1003_ & new_n1009_;
  assign new_n1021_ = pk2 & new_n1017_;
  assign new_n1022_ = ~new_n1004_ & ~new_n1005_;
  assign new_n1023_ = ~new_n1007_ & new_n1022_;
  assign new_n1024_ = ~new_n1010_ & ~new_n1011_;
  assign new_n1025_ = new_n1023_ & new_n1024_;
  assign new_n1026_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1027_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1028_ = new_n1026_ & new_n1027_;
  assign new_n1029_ = new_n1025_ & new_n1028_;
  assign new_n1030_ = new_n990_ & ~new_n1029_;
  assign new_n1031_ = ~px1 & new_n1030_;
  assign new_n1032_ = ~pm0 & new_n986_;
  assign new_n1033_ = pa2 & ~py1;
  assign new_n1034_ = new_n986_ & ~new_n1033_;
  assign new_n1035_ = ~px1 & ~new_n1033_;
  assign new_n1036_ = ~pd0 & new_n503_;
  assign new_n1037_ = pf2 & ~pe2;
  assign new_n1038_ = pd0 & new_n1037_;
  assign new_n1039_ = ~new_n1036_ & ~new_n1038_;
  assign new_n1040_ = ~px1 & new_n1039_;
  assign new_n1041_ = ~pm0 & ~px1;
  assign new_n1042_ = ~new_n990_ & ~new_n1033_;
  assign new_n1043_ = ~new_n990_ & new_n1039_;
  assign new_n1044_ = new_n986_ & new_n1039_;
  assign new_n1045_ = ~pm0 & ~new_n990_;
  assign new_n1046_ = ~new_n1032_ & ~new_n1034_;
  assign new_n1047_ = ~new_n1035_ & new_n1046_;
  assign new_n1048_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1049_ = new_n1047_ & new_n1048_;
  assign new_n1050_ = ~new_n1044_ & ~new_n1045_;
  assign new_n1051_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1052_ = new_n1050_ & new_n1051_;
  assign new_n1053_ = new_n1049_ & new_n1052_;
  assign new_n1054_ = ~new_n989_ & ~new_n1031_;
  assign pk4 = new_n1053_ | ~new_n1054_;
  assign new_n1056_ = ~pq & ~pr;
  assign new_n1057_ = pi & new_n1056_;
  assign new_n1058_ = ~pq & ~py0;
  assign new_n1059_ = pr & ~py0;
  assign new_n1060_ = ~pi & ~py0;
  assign new_n1061_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1062_ = ~new_n1059_ & ~new_n1060_;
  assign new_n1063_ = new_n1061_ & new_n1062_;
  assign pt4 = ~py1 & new_n1063_;
  assign new_n1065_ = ~py1 & ~pz1;
  assign new_n1066_ = pi3 & ~pr2;
  assign new_n1067_ = ~pi2 & ~new_n276_;
  assign new_n1068_ = pi3 & new_n1067_;
  assign new_n1069_ = pc0 & ~pd0;
  assign new_n1070_ = ~pd0 & ~pq2;
  assign new_n1071_ = ~new_n1013_ & ~new_n1069_;
  assign new_n1072_ = ~new_n1070_ & new_n1071_;
  assign new_n1073_ = new_n1009_ & new_n1072_;
  assign new_n1074_ = ~new_n1068_ & ~new_n1073_;
  assign new_n1075_ = ~new_n1066_ & new_n1074_;
  assign new_n1076_ = new_n986_ & new_n1075_;
  assign new_n1077_ = ~new_n276_ & new_n1075_;
  assign new_n1078_ = pq2 & new_n1074_;
  assign new_n1079_ = ~new_n276_ & new_n1078_;
  assign new_n1080_ = new_n1009_ & new_n1078_;
  assign new_n1081_ = new_n986_ & new_n1078_;
  assign new_n1082_ = new_n276_ & new_n1074_;
  assign new_n1083_ = ~new_n276_ & new_n1082_;
  assign new_n1084_ = new_n1009_ & new_n1082_;
  assign new_n1085_ = new_n1009_ & new_n1075_;
  assign new_n1086_ = new_n986_ & new_n1082_;
  assign new_n1087_ = ~new_n1076_ & ~new_n1077_;
  assign new_n1088_ = ~new_n1079_ & new_n1087_;
  assign new_n1089_ = ~new_n1080_ & ~new_n1081_;
  assign new_n1090_ = new_n1088_ & new_n1089_;
  assign new_n1091_ = ~new_n1085_ & ~new_n1086_;
  assign new_n1092_ = ~new_n1083_ & ~new_n1084_;
  assign new_n1093_ = new_n1091_ & new_n1092_;
  assign new_n1094_ = new_n1090_ & new_n1093_;
  assign new_n1095_ = new_n1065_ & new_n1094_;
  assign new_n1096_ = ~px1 & new_n1095_;
  assign new_n1097_ = ~pi3 & ~pr2;
  assign new_n1098_ = ~pi3 & new_n1067_;
  assign new_n1099_ = pd0 & ~px1;
  assign new_n1100_ = ~pc0 & new_n1099_;
  assign new_n1101_ = pd0 & ~pq2;
  assign new_n1102_ = ~px1 & new_n1101_;
  assign new_n1103_ = ~pr2 & ~px1;
  assign new_n1104_ = ~pc0 & new_n1103_;
  assign new_n1105_ = ~px1 & new_n1008_;
  assign new_n1106_ = ~pi2 & ~px1;
  assign new_n1107_ = ~new_n1100_ & ~new_n1102_;
  assign new_n1108_ = ~new_n1104_ & new_n1107_;
  assign new_n1109_ = ~new_n1105_ & ~new_n1106_;
  assign new_n1110_ = new_n1108_ & new_n1109_;
  assign new_n1111_ = ~new_n1098_ & ~new_n1110_;
  assign new_n1112_ = ~new_n1097_ & new_n1111_;
  assign new_n1113_ = ~new_n986_ & new_n1112_;
  assign new_n1114_ = ~new_n276_ & new_n1112_;
  assign new_n1115_ = pq2 & new_n1111_;
  assign new_n1116_ = ~new_n276_ & new_n1115_;
  assign new_n1117_ = new_n1009_ & new_n1115_;
  assign new_n1118_ = ~new_n986_ & new_n1115_;
  assign new_n1119_ = new_n276_ & new_n1111_;
  assign new_n1120_ = ~new_n276_ & new_n1119_;
  assign new_n1121_ = new_n1009_ & new_n1119_;
  assign new_n1122_ = new_n1009_ & new_n1112_;
  assign new_n1123_ = ~new_n986_ & new_n1119_;
  assign new_n1124_ = ~new_n1113_ & ~new_n1114_;
  assign new_n1125_ = ~new_n1116_ & new_n1124_;
  assign new_n1126_ = ~new_n1117_ & ~new_n1118_;
  assign new_n1127_ = new_n1125_ & new_n1126_;
  assign new_n1128_ = ~new_n1122_ & ~new_n1123_;
  assign new_n1129_ = ~new_n1120_ & ~new_n1121_;
  assign new_n1130_ = new_n1128_ & new_n1129_;
  assign new_n1131_ = new_n1127_ & new_n1130_;
  assign new_n1132_ = ~py1 & new_n1131_;
  assign new_n1133_ = pz1 & new_n1132_;
  assign new_n1134_ = ~py1 & ~px1;
  assign new_n1135_ = pi2 & new_n1134_;
  assign new_n1136_ = pq2 & new_n1135_;
  assign new_n1137_ = pr2 & new_n1136_;
  assign new_n1138_ = ~new_n1096_ & ~new_n1133_;
  assign pu5 = new_n1137_ | ~new_n1138_;
  assign new_n1140_ = ~pa3 & ~pf;
  assign new_n1141_ = ~pb3 & ph;
  assign new_n1142_ = pf & new_n1141_;
  assign new_n1143_ = ~new_n1140_ & ~new_n1142_;
  assign new_n1144_ = ~py1 & new_n1143_;
  assign new_n1145_ = ph & new_n1144_;
  assign new_n1146_ = pa3 & new_n1144_;
  assign pv6 = new_n1145_ | new_n1146_;
  assign new_n1148_ = new_n573_ & new_n641_;
  assign new_n1149_ = ~pz3 & new_n1148_;
  assign new_n1150_ = ~py3 & new_n1148_;
  assign new_n1151_ = pb4 & new_n573_;
  assign new_n1152_ = ~py3 & new_n1151_;
  assign new_n1153_ = ~new_n577_ & new_n1151_;
  assign new_n1154_ = ~pz3 & new_n1151_;
  assign new_n1155_ = ~new_n577_ & new_n1148_;
  assign new_n1156_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1157_ = ~new_n1152_ & new_n1156_;
  assign new_n1158_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1159_ = ~new_n1155_ & new_n1158_;
  assign pw7 = ~new_n1157_ | ~new_n1159_;
  assign new_n1161_ = ~px1 & new_n740_;
  assign new_n1162_ = pi2 & new_n1161_;
  assign pt5 = pn0 | new_n1162_;
  assign new_n1164_ = pr & ~pj;
  assign new_n1165_ = pi & new_n1164_;
  assign new_n1166_ = ~pj & ~pz0;
  assign new_n1167_ = ~pr & ~pz0;
  assign new_n1168_ = ~pi & ~pz0;
  assign new_n1169_ = ~new_n1165_ & ~new_n1166_;
  assign new_n1170_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1171_ = new_n1169_ & new_n1170_;
  assign pu4 = ~py1 & new_n1171_;
  assign new_n1173_ = py3 & new_n567_;
  assign new_n1174_ = ~pl0 & ~new_n1173_;
  assign new_n1175_ = ~pn0 & new_n1174_;
  assign new_n1176_ = py3 & new_n1175_;
  assign new_n1177_ = pz3 & new_n1176_;
  assign new_n1178_ = pa4 & new_n1175_;
  assign pv7 = new_n1177_ | new_n1178_;
  assign new_n1180_ = ~pb3 & ~pf;
  assign new_n1181_ = ~pc3 & ph;
  assign new_n1182_ = pf & new_n1181_;
  assign new_n1183_ = ~new_n1180_ & ~new_n1182_;
  assign new_n1184_ = ~py1 & new_n1183_;
  assign new_n1185_ = ph & new_n1184_;
  assign new_n1186_ = pb3 & new_n1184_;
  assign pw6 = new_n1185_ | new_n1186_;
  assign new_n1188_ = ~pf & ~py2;
  assign new_n1189_ = ~ph & ~pz2;
  assign new_n1190_ = pf & new_n1189_;
  assign new_n1191_ = ~new_n1188_ & ~new_n1190_;
  assign new_n1192_ = ~py1 & new_n1191_;
  assign new_n1193_ = ~ph & new_n1192_;
  assign new_n1194_ = py2 & new_n1192_;
  assign pt6 = new_n1193_ | new_n1194_;
  assign new_n1196_ = ~pl0 & ~new_n574_;
  assign new_n1197_ = ~pn0 & new_n1196_;
  assign new_n1198_ = py3 & new_n1197_;
  assign new_n1199_ = pz3 & new_n1197_;
  assign pu7 = new_n1198_ | new_n1199_;
  assign new_n1201_ = pr & ~pk;
  assign new_n1202_ = pi & new_n1201_;
  assign new_n1203_ = ~pa1 & ~pk;
  assign new_n1204_ = ~pa1 & ~pr;
  assign new_n1205_ = ~pa1 & ~pi;
  assign new_n1206_ = ~new_n1202_ & ~new_n1203_;
  assign new_n1207_ = ~new_n1204_ & ~new_n1205_;
  assign new_n1208_ = new_n1206_ & new_n1207_;
  assign pv4 = ~py1 & new_n1208_;
  assign new_n1210_ = pd4 & new_n644_;
  assign new_n1211_ = ~pe4 & ~pf4;
  assign new_n1212_ = ~pg4 & new_n1211_;
  assign new_n1213_ = new_n1210_ & new_n1212_;
  assign new_n1214_ = new_n641_ & new_n1213_;
  assign new_n1215_ = ~pf4 & ~pg4;
  assign new_n1216_ = pb2 & new_n1215_;
  assign new_n1217_ = py3 & new_n1216_;
  assign new_n1218_ = new_n573_ & new_n1214_;
  assign new_n1219_ = ~new_n1217_ & new_n1218_;
  assign new_n1220_ = ~new_n568_ & new_n1218_;
  assign new_n1221_ = pb2 & new_n573_;
  assign new_n1222_ = ~new_n568_ & new_n1221_;
  assign new_n1223_ = pd4 & pc4;
  assign new_n1224_ = ~pe4 & new_n1223_;
  assign new_n1225_ = new_n1221_ & ~new_n1224_;
  assign new_n1226_ = ~new_n1217_ & new_n1221_;
  assign new_n1227_ = new_n1218_ & ~new_n1224_;
  assign new_n1228_ = ~new_n1219_ & ~new_n1220_;
  assign new_n1229_ = ~new_n1222_ & new_n1228_;
  assign new_n1230_ = ~new_n1225_ & ~new_n1226_;
  assign new_n1231_ = ~new_n1227_ & new_n1230_;
  assign pw5 = ~new_n1229_ | ~new_n1231_;
  assign pt7 = ~py3 & new_n573_;
  assign new_n1234_ = ~pf & ~pz2;
  assign new_n1235_ = ~pg & ~ph;
  assign new_n1236_ = pf & new_n1235_;
  assign new_n1237_ = ~new_n1234_ & ~new_n1236_;
  assign new_n1238_ = ~py1 & new_n1237_;
  assign new_n1239_ = ~ph & new_n1238_;
  assign new_n1240_ = pz2 & new_n1238_;
  assign pu6 = new_n1239_ | new_n1240_;
  assign new_n1242_ = pa2 & ~pf2;
  assign new_n1243_ = pa2 & ~pe2;
  assign new_n1244_ = ~new_n498_ & ~new_n1242_;
  assign new_n1245_ = ~new_n1243_ & new_n1244_;
  assign new_n1246_ = ~new_n462_ & new_n1245_;
  assign new_n1247_ = ~new_n464_ & new_n1245_;
  assign new_n1248_ = ph0 & new_n1245_;
  assign new_n1249_ = ~new_n1246_ & ~new_n1247_;
  assign new_n1250_ = ~new_n1248_ & new_n1249_;
  assign pv5 = ~py1 & new_n1250_;
  assign new_n1252_ = pr & ~pl;
  assign new_n1253_ = pi & new_n1252_;
  assign new_n1254_ = ~pb1 & ~pl;
  assign new_n1255_ = ~pr & ~pb1;
  assign new_n1256_ = ~pb1 & ~pi;
  assign new_n1257_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1258_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1259_ = new_n1257_ & new_n1258_;
  assign pw4 = ~py1 & new_n1259_;
  assign new_n1261_ = ~pr & ~pm;
  assign new_n1262_ = pi & new_n1261_;
  assign new_n1263_ = ~pu0 & ~pm;
  assign new_n1264_ = pr & ~pu0;
  assign new_n1265_ = ~pu0 & ~pi;
  assign new_n1266_ = ~new_n1262_ & ~new_n1263_;
  assign new_n1267_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1268_ = new_n1266_ & new_n1267_;
  assign pp4 = ~py1 & new_n1268_;
  assign new_n1270_ = pb0 & ~pz;
  assign new_n1271_ = ps & new_n1270_;
  assign new_n1272_ = ~pz & ~pv1;
  assign new_n1273_ = ~pb0 & ~pv1;
  assign new_n1274_ = ~ps & ~pv1;
  assign new_n1275_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1276_ = ~new_n1273_ & ~new_n1274_;
  assign new_n1277_ = new_n1275_ & new_n1276_;
  assign pq5 = ~py1 & new_n1277_;
  assign new_n1279_ = ~pw2 & ~pf;
  assign new_n1280_ = ~ph & ~px2;
  assign new_n1281_ = pf & new_n1280_;
  assign new_n1282_ = ~new_n1279_ & ~new_n1281_;
  assign new_n1283_ = ~py1 & new_n1282_;
  assign new_n1284_ = ~ph & new_n1283_;
  assign new_n1285_ = pw2 & new_n1283_;
  assign pr6 = new_n1284_ | new_n1285_;
  assign new_n1287_ = pe & ~pw1;
  assign new_n1288_ = ~pg1 & ~pe;
  assign new_n1289_ = pd & new_n1288_;
  assign new_n1290_ = ~ph3 & new_n264_;
  assign new_n1291_ = ~new_n1287_ & ~new_n1289_;
  assign new_n1292_ = ~new_n1290_ & new_n1291_;
  assign new_n1293_ = ~py1 & new_n1292_;
  assign new_n1294_ = ~new_n268_ & new_n1293_;
  assign new_n1295_ = pk2 & ~px1;
  assign new_n1296_ = pj2 & ~px1;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = px3 & new_n1297_;
  assign new_n1299_ = new_n1293_ & new_n1298_;
  assign new_n1300_ = pc & new_n1293_;
  assign new_n1301_ = ~new_n1294_ & ~new_n1299_;
  assign ps7 = new_n1300_ | ~new_n1301_;
  assign new_n1303_ = pb0 & ~py;
  assign new_n1304_ = ps & new_n1303_;
  assign new_n1305_ = ~py & ~pu1;
  assign new_n1306_ = ~pb0 & ~pu1;
  assign new_n1307_ = ~ps & ~pu1;
  assign new_n1308_ = ~new_n1304_ & ~new_n1305_;
  assign new_n1309_ = ~new_n1306_ & ~new_n1307_;
  assign new_n1310_ = new_n1308_ & new_n1309_;
  assign pp5 = ~py1 & new_n1310_;
  assign new_n1312_ = ~pr & ~pn;
  assign new_n1313_ = pi & new_n1312_;
  assign new_n1314_ = ~pv0 & ~pn;
  assign new_n1315_ = pr & ~pv0;
  assign new_n1316_ = ~pv0 & ~pi;
  assign new_n1317_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1318_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1319_ = new_n1317_ & new_n1318_;
  assign pq4 = ~py1 & new_n1319_;
  assign new_n1321_ = pe & ~pv1;
  assign new_n1322_ = ~pf1 & ~pe;
  assign new_n1323_ = pd & new_n1322_;
  assign new_n1324_ = ~pg3 & new_n264_;
  assign new_n1325_ = ~new_n1321_ & ~new_n1323_;
  assign new_n1326_ = ~new_n1324_ & new_n1325_;
  assign new_n1327_ = ~py1 & new_n1326_;
  assign new_n1328_ = ~new_n268_ & new_n1327_;
  assign new_n1329_ = ~pk2 & pw3;
  assign new_n1330_ = ~pj2 & new_n1329_;
  assign new_n1331_ = pw3 & px1;
  assign new_n1332_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1333_ = px1 & new_n1332_;
  assign new_n1334_ = new_n276_ & new_n1332_;
  assign new_n1335_ = ~px3 & new_n1332_;
  assign new_n1336_ = ~new_n1333_ & ~new_n1334_;
  assign new_n1337_ = ~new_n1335_ & new_n1336_;
  assign new_n1338_ = new_n1327_ & new_n1337_;
  assign new_n1339_ = pc & new_n1327_;
  assign new_n1340_ = ~new_n1328_ & ~new_n1338_;
  assign pr7 = new_n1339_ | ~new_n1340_;
  assign new_n1342_ = ~pf & ~px2;
  assign new_n1343_ = ~ph & ~py2;
  assign new_n1344_ = pf & new_n1343_;
  assign new_n1345_ = ~new_n1342_ & ~new_n1344_;
  assign new_n1346_ = ~py1 & new_n1345_;
  assign new_n1347_ = ~ph & new_n1346_;
  assign new_n1348_ = px2 & new_n1346_;
  assign ps6 = new_n1347_ | new_n1348_;
  assign new_n1350_ = ~pf & ~pu2;
  assign new_n1351_ = ~pv2 & ~ph;
  assign new_n1352_ = pf & new_n1351_;
  assign new_n1353_ = ~new_n1350_ & ~new_n1352_;
  assign new_n1354_ = ~py1 & new_n1353_;
  assign new_n1355_ = ~ph & new_n1354_;
  assign new_n1356_ = pu2 & new_n1354_;
  assign pp6 = new_n1355_ | new_n1356_;
  assign new_n1358_ = ~pu1 & pe;
  assign new_n1359_ = ~pe1 & ~pe;
  assign new_n1360_ = pd & new_n1359_;
  assign new_n1361_ = ~pf3 & new_n264_;
  assign new_n1362_ = ~new_n1358_ & ~new_n1360_;
  assign new_n1363_ = ~new_n1361_ & new_n1362_;
  assign new_n1364_ = ~py1 & new_n1363_;
  assign new_n1365_ = ~new_n268_ & new_n1364_;
  assign new_n1366_ = ~pk2 & pv3;
  assign new_n1367_ = ~pj2 & new_n1366_;
  assign new_n1368_ = pv3 & px1;
  assign new_n1369_ = ~new_n1367_ & ~new_n1368_;
  assign new_n1370_ = px1 & new_n1369_;
  assign new_n1371_ = new_n276_ & new_n1369_;
  assign new_n1372_ = ~pw3 & new_n1369_;
  assign new_n1373_ = ~new_n1370_ & ~new_n1371_;
  assign new_n1374_ = ~new_n1372_ & new_n1373_;
  assign new_n1375_ = new_n1364_ & new_n1374_;
  assign new_n1376_ = pc & new_n1364_;
  assign new_n1377_ = ~new_n1365_ & ~new_n1375_;
  assign pq7 = new_n1376_ | ~new_n1377_;
  assign new_n1379_ = ~pr & ~po;
  assign new_n1380_ = pi & new_n1379_;
  assign new_n1381_ = ~pw0 & ~po;
  assign new_n1382_ = pr & ~pw0;
  assign new_n1383_ = ~pw0 & ~pi;
  assign new_n1384_ = ~new_n1380_ & ~new_n1381_;
  assign new_n1385_ = ~new_n1382_ & ~new_n1383_;
  assign new_n1386_ = new_n1384_ & new_n1385_;
  assign pr4 = ~py1 & new_n1386_;
  assign ps5 = py1 | new_n321_;
  assign new_n1389_ = pe & ~pt1;
  assign new_n1390_ = ~pd1 & ~pe;
  assign new_n1391_ = pd & new_n1390_;
  assign new_n1392_ = ~pe3 & new_n264_;
  assign new_n1393_ = ~new_n1389_ & ~new_n1391_;
  assign new_n1394_ = ~new_n1392_ & new_n1393_;
  assign new_n1395_ = ~py1 & new_n1394_;
  assign new_n1396_ = ~new_n268_ & new_n1395_;
  assign new_n1397_ = ~pk2 & pu3;
  assign new_n1398_ = ~pj2 & new_n1397_;
  assign new_n1399_ = pu3 & px1;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = px1 & new_n1400_;
  assign new_n1402_ = new_n276_ & new_n1400_;
  assign new_n1403_ = ~pv3 & new_n1400_;
  assign new_n1404_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1405_ = ~new_n1403_ & new_n1404_;
  assign new_n1406_ = new_n1395_ & new_n1405_;
  assign new_n1407_ = pc & new_n1395_;
  assign new_n1408_ = ~new_n1396_ & ~new_n1406_;
  assign pp7 = new_n1407_ | ~new_n1408_;
  assign new_n1410_ = ~pv2 & ~pf;
  assign new_n1411_ = ~pw2 & ~ph;
  assign new_n1412_ = pf & new_n1411_;
  assign new_n1413_ = ~new_n1410_ & ~new_n1412_;
  assign new_n1414_ = ~py1 & new_n1413_;
  assign new_n1415_ = ~ph & new_n1414_;
  assign new_n1416_ = pv2 & new_n1414_;
  assign pq6 = new_n1415_ | new_n1416_;
  assign new_n1418_ = ~pa0 & pb0;
  assign new_n1419_ = ps & new_n1418_;
  assign new_n1420_ = ~pa0 & ~pw1;
  assign new_n1421_ = ~pb0 & ~pw1;
  assign new_n1422_ = ~ps & ~pw1;
  assign new_n1423_ = ~new_n1419_ & ~new_n1420_;
  assign new_n1424_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1425_ = new_n1423_ & new_n1424_;
  assign pr5 = ~py1 & new_n1425_;
  assign new_n1427_ = ~pp & ~pr;
  assign new_n1428_ = pi & new_n1427_;
  assign new_n1429_ = ~pp & ~px0;
  assign new_n1430_ = pr & ~px0;
  assign new_n1431_ = ~px0 & ~pi;
  assign new_n1432_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1433_ = ~new_n1430_ & ~new_n1431_;
  assign new_n1434_ = new_n1432_ & new_n1433_;
  assign ps4 = ~py1 & new_n1434_;
  assign new_n1436_ = pr & ~pm;
  assign new_n1437_ = pi & new_n1436_;
  assign new_n1438_ = ~pc1 & ~pm;
  assign new_n1439_ = ~pc1 & ~pr;
  assign new_n1440_ = ~pc1 & ~pi;
  assign new_n1441_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1442_ = ~new_n1439_ & ~new_n1440_;
  assign new_n1443_ = new_n1441_ & new_n1442_;
  assign px4 = ~py1 & new_n1443_;
  assign new_n1445_ = ~pd2 & ~pl0;
  assign new_n1446_ = pb & ~new_n1445_;
  assign new_n1447_ = ~pn0 & new_n1446_;
  assign new_n1448_ = ~pg2 & new_n1447_;
  assign new_n1449_ = ~ph2 & new_n1447_;
  assign py5 = new_n1448_ | new_n1449_;
  assign new_n1451_ = ~pe3 & ~pf;
  assign new_n1452_ = ~pf3 & ph;
  assign new_n1453_ = pf & new_n1452_;
  assign new_n1454_ = ~new_n1451_ & ~new_n1453_;
  assign new_n1455_ = ~py1 & new_n1454_;
  assign new_n1456_ = ph & new_n1455_;
  assign new_n1457_ = pe3 & new_n1455_;
  assign pz6 = new_n1456_ | new_n1457_;
  assign new_n1459_ = new_n568_ & new_n1224_;
  assign new_n1460_ = new_n1217_ & new_n1459_;
  assign new_n1461_ = new_n527_ & ~new_n1460_;
  assign new_n1462_ = ~pl0 & new_n1461_;
  assign new_n1463_ = pb2 & ~pn0;
  assign new_n1464_ = ~pc2 & new_n1463_;
  assign new_n1465_ = ~pl0 & new_n1213_;
  assign new_n1466_ = new_n641_ & new_n1464_;
  assign new_n1467_ = new_n1465_ & new_n1466_;
  assign px5 = new_n1462_ | new_n1467_;
  assign new_n1469_ = pr & ~pn;
  assign new_n1470_ = pi & new_n1469_;
  assign new_n1471_ = ~pd1 & ~pn;
  assign new_n1472_ = ~pr & ~pd1;
  assign new_n1473_ = ~pd1 & ~pi;
  assign new_n1474_ = ~new_n1470_ & ~new_n1471_;
  assign new_n1475_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1476_ = new_n1474_ & new_n1475_;
  assign py4 = ~py1 & new_n1476_;
  assign new_n1478_ = new_n567_ & new_n645_;
  assign new_n1479_ = py3 & new_n1478_;
  assign new_n1480_ = new_n573_ & new_n1479_;
  assign new_n1481_ = ~py3 & new_n1480_;
  assign new_n1482_ = ~new_n568_ & new_n1480_;
  assign new_n1483_ = pe4 & new_n573_;
  assign new_n1484_ = ~new_n568_ & new_n1483_;
  assign new_n1485_ = ~new_n570_ & new_n1483_;
  assign new_n1486_ = ~py3 & new_n1483_;
  assign new_n1487_ = ~new_n570_ & new_n1480_;
  assign new_n1488_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1489_ = ~new_n1484_ & new_n1488_;
  assign new_n1490_ = ~new_n1485_ & ~new_n1486_;
  assign new_n1491_ = ~new_n1487_ & new_n1490_;
  assign pz7 = ~new_n1489_ | ~new_n1491_;
  assign new_n1493_ = ~pc3 & ~pf;
  assign new_n1494_ = ~pd3 & ph;
  assign new_n1495_ = pf & new_n1494_;
  assign new_n1496_ = ~new_n1493_ & ~new_n1495_;
  assign new_n1497_ = ~py1 & new_n1496_;
  assign new_n1498_ = ph & new_n1497_;
  assign new_n1499_ = pc3 & new_n1497_;
  assign px6 = new_n1498_ | new_n1499_;
  assign new_n1501_ = py3 & new_n578_;
  assign new_n1502_ = pz3 & new_n1501_;
  assign new_n1503_ = new_n573_ & new_n1502_;
  assign new_n1504_ = ~py3 & new_n1503_;
  assign new_n1505_ = ~new_n567_ & new_n1503_;
  assign new_n1506_ = pd4 & new_n573_;
  assign new_n1507_ = ~new_n567_ & new_n1506_;
  assign new_n1508_ = ~new_n1210_ & new_n1506_;
  assign new_n1509_ = ~py3 & new_n1506_;
  assign new_n1510_ = ~new_n1210_ & new_n1503_;
  assign new_n1511_ = ~new_n1504_ & ~new_n1505_;
  assign new_n1512_ = ~new_n1507_ & new_n1511_;
  assign new_n1513_ = ~new_n1508_ & ~new_n1509_;
  assign new_n1514_ = ~new_n1510_ & new_n1513_;
  assign py7 = ~new_n1512_ | ~new_n1514_;
  assign new_n1516_ = pr & ~po;
  assign new_n1517_ = pi & new_n1516_;
  assign new_n1518_ = ~pe1 & ~po;
  assign new_n1519_ = ~pr & ~pe1;
  assign new_n1520_ = ~pe1 & ~pi;
  assign new_n1521_ = ~new_n1517_ & ~new_n1518_;
  assign new_n1522_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1523_ = new_n1521_ & new_n1522_;
  assign pz4 = ~py1 & new_n1523_;
  assign new_n1525_ = py3 & new_n577_;
  assign new_n1526_ = pz3 & new_n1525_;
  assign new_n1527_ = new_n573_ & new_n1526_;
  assign new_n1528_ = ~pz3 & new_n1527_;
  assign new_n1529_ = ~py3 & new_n1527_;
  assign new_n1530_ = pc4 & new_n573_;
  assign new_n1531_ = ~py3 & new_n1530_;
  assign new_n1532_ = ~new_n578_ & new_n1530_;
  assign new_n1533_ = ~pz3 & new_n1530_;
  assign new_n1534_ = ~new_n578_ & new_n1527_;
  assign new_n1535_ = ~new_n1528_ & ~new_n1529_;
  assign new_n1536_ = ~new_n1531_ & new_n1535_;
  assign new_n1537_ = ~new_n1532_ & ~new_n1533_;
  assign new_n1538_ = ~new_n1534_ & new_n1537_;
  assign px7 = ~new_n1536_ | ~new_n1538_;
  assign new_n1540_ = ~pd3 & ~pf;
  assign new_n1541_ = ~pe3 & ph;
  assign new_n1542_ = pf & new_n1541_;
  assign new_n1543_ = ~new_n1540_ & ~new_n1542_;
  assign new_n1544_ = ~py1 & new_n1543_;
  assign new_n1545_ = ph & new_n1544_;
  assign new_n1546_ = pd3 & new_n1544_;
  assign py6 = new_n1545_ | new_n1546_;
  assign new_n1548_ = ~pe2 & new_n509_;
  assign new_n1549_ = ~pn0 & new_n1548_;
  assign new_n1550_ = ~pa2 & pe2;
  assign new_n1551_ = new_n499_ & new_n1550_;
  assign new_n1552_ = ~pn0 & new_n1551_;
  assign pz5 = new_n1549_ | new_n1552_;
endmodule

