module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pu, pv, pw, px, py, pz, pa, pb, pc, pd,
    pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pd0, pe0, pf0, pg0, ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0,
    pr0, ps0, pt0, pu0  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pu, pv, pw, px, py, pz, pa, pb,
    pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po;
  output pd0, pe0, pf0, pg0, ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0,
    pr0, ps0, pt0, pu0;
  wire new_n47_, new_n48_, new_n49_, new_n50_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n57_, new_n58_, new_n59_, new_n60_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n67_, new_n68_, new_n69_, new_n70_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_;
  assign new_n47_ = pc0 & ~pi;
  assign new_n48_ = ~pc0 & ~pu;
  assign new_n49_ = ~pu & ~pi;
  assign new_n50_ = ~new_n47_ & ~new_n48_;
  assign pd0 = new_n49_ | ~new_n50_;
  assign new_n52_ = pc0 & ~pj;
  assign new_n53_ = ~pc0 & ~pv;
  assign new_n54_ = ~pv & ~pj;
  assign new_n55_ = ~new_n52_ & ~new_n53_;
  assign pe0 = new_n54_ | ~new_n55_;
  assign new_n57_ = pc0 & ~pk;
  assign new_n58_ = ~pc0 & ~pw;
  assign new_n59_ = ~pw & ~pk;
  assign new_n60_ = ~new_n57_ & ~new_n58_;
  assign pf0 = new_n59_ | ~new_n60_;
  assign new_n62_ = pc0 & ~pl;
  assign new_n63_ = ~pc0 & ~px;
  assign new_n64_ = ~px & ~pl;
  assign new_n65_ = ~new_n62_ & ~new_n63_;
  assign pg0 = new_n64_ | ~new_n65_;
  assign new_n67_ = pc0 & ~pm;
  assign new_n68_ = ~pc0 & ~py;
  assign new_n69_ = ~py & ~pm;
  assign new_n70_ = ~new_n67_ & ~new_n68_;
  assign ph0 = new_n69_ | ~new_n70_;
  assign new_n72_ = pc0 & ~pn;
  assign new_n73_ = ~pc0 & ~pz;
  assign new_n74_ = ~pz & ~pn;
  assign new_n75_ = ~new_n72_ & ~new_n73_;
  assign pi0 = new_n74_ | ~new_n75_;
  assign new_n77_ = pc0 & ~po;
  assign new_n78_ = ~pa0 & ~pc0;
  assign new_n79_ = ~pa0 & ~po;
  assign new_n80_ = ~new_n77_ & ~new_n78_;
  assign pj0 = new_n79_ | ~new_n80_;
  assign new_n82_ = ~pp & pc0;
  assign new_n83_ = ~pb0 & ~pc0;
  assign new_n84_ = ~pp & ~pb0;
  assign new_n85_ = ~new_n82_ & ~new_n83_;
  assign pk0 = new_n84_ | ~new_n85_;
  assign new_n87_ = ~pq & pa;
  assign new_n88_ = pi & new_n87_;
  assign new_n89_ = ps & pa;
  assign new_n90_ = ~pq & new_n89_;
  assign new_n91_ = pr & pu;
  assign new_n92_ = pq & new_n91_;
  assign new_n93_ = ~pr & ~pu;
  assign new_n94_ = pq & new_n93_;
  assign new_n95_ = ~pq & ~ps;
  assign new_n96_ = pi & new_n95_;
  assign new_n97_ = ~pu & new_n89_;
  assign new_n98_ = ~pr & new_n97_;
  assign new_n99_ = ~pr & pa;
  assign new_n100_ = ~pu & new_n99_;
  assign new_n101_ = pi & new_n100_;
  assign new_n102_ = pr & pa;
  assign new_n103_ = pu & new_n102_;
  assign new_n104_ = pi & new_n103_;
  assign new_n105_ = pu & new_n89_;
  assign new_n106_ = pr & new_n105_;
  assign new_n107_ = ~ps & new_n91_;
  assign new_n108_ = pi & new_n107_;
  assign new_n109_ = ~ps & new_n93_;
  assign new_n110_ = pi & new_n109_;
  assign new_n111_ = ~new_n108_ & ~new_n110_;
  assign new_n112_ = ~new_n101_ & ~new_n104_;
  assign new_n113_ = ~new_n106_ & new_n112_;
  assign new_n114_ = new_n111_ & new_n113_;
  assign new_n115_ = ~new_n88_ & ~new_n90_;
  assign new_n116_ = ~new_n92_ & new_n115_;
  assign new_n117_ = ~new_n94_ & ~new_n96_;
  assign new_n118_ = ~new_n98_ & new_n117_;
  assign new_n119_ = new_n116_ & new_n118_;
  assign pm0 = ~new_n114_ | ~new_n119_;
  assign new_n121_ = ~pj & new_n95_;
  assign new_n122_ = ~pr & pv;
  assign new_n123_ = ~pu & new_n122_;
  assign new_n124_ = pq & new_n123_;
  assign new_n125_ = ~pq & ps;
  assign new_n126_ = ~pb & new_n125_;
  assign new_n127_ = ~new_n121_ & ~new_n124_;
  assign new_n128_ = ~new_n126_ & new_n127_;
  assign new_n129_ = ~pq & new_n128_;
  assign new_n130_ = new_n93_ & new_n128_;
  assign new_n131_ = pv & new_n128_;
  assign new_n132_ = ~new_n129_ & ~new_n130_;
  assign pn0 = new_n131_ | ~new_n132_;
  assign new_n134_ = ~pc & new_n125_;
  assign new_n135_ = ~pk & new_n95_;
  assign new_n136_ = ~pq & ~pk;
  assign new_n137_ = ~pc & new_n136_;
  assign new_n138_ = ~new_n134_ & ~new_n135_;
  assign new_n139_ = ~new_n137_ & new_n138_;
  assign new_n140_ = ~pv & pw;
  assign new_n141_ = pw & new_n139_;
  assign new_n142_ = ~new_n140_ & new_n141_;
  assign new_n143_ = ~pv & new_n93_;
  assign new_n144_ = new_n139_ & new_n143_;
  assign new_n145_ = pu & new_n144_;
  assign new_n146_ = pu & new_n141_;
  assign new_n147_ = pr & new_n141_;
  assign new_n148_ = ~pq & new_n139_;
  assign new_n149_ = pr & new_n144_;
  assign new_n150_ = ~new_n140_ & new_n144_;
  assign new_n151_ = ~new_n148_ & ~new_n149_;
  assign new_n152_ = ~new_n150_ & new_n151_;
  assign new_n153_ = ~new_n146_ & ~new_n147_;
  assign new_n154_ = ~new_n142_ & ~new_n145_;
  assign new_n155_ = new_n153_ & new_n154_;
  assign po0 = ~new_n152_ | ~new_n155_;
  assign new_n157_ = ~pd & new_n125_;
  assign new_n158_ = ~pl & new_n95_;
  assign new_n159_ = ~pq & ~pl;
  assign new_n160_ = ~pd & new_n159_;
  assign new_n161_ = ~new_n157_ & ~new_n158_;
  assign new_n162_ = ~new_n160_ & new_n161_;
  assign new_n163_ = ~pv & ~pw;
  assign new_n164_ = px & new_n163_;
  assign new_n165_ = px & new_n162_;
  assign new_n166_ = ~new_n164_ & new_n165_;
  assign new_n167_ = ~pu & ~pw;
  assign new_n168_ = ~pr & ~pv;
  assign new_n169_ = new_n167_ & new_n168_;
  assign new_n170_ = new_n162_ & new_n169_;
  assign new_n171_ = pu & new_n170_;
  assign new_n172_ = pu & new_n165_;
  assign new_n173_ = pr & new_n165_;
  assign new_n174_ = ~pq & new_n162_;
  assign new_n175_ = pr & new_n170_;
  assign new_n176_ = ~new_n164_ & new_n170_;
  assign new_n177_ = ~new_n174_ & ~new_n175_;
  assign new_n178_ = ~new_n176_ & new_n177_;
  assign new_n179_ = ~new_n172_ & ~new_n173_;
  assign new_n180_ = ~new_n166_ & ~new_n171_;
  assign new_n181_ = new_n179_ & new_n180_;
  assign pp0 = ~new_n178_ | ~new_n181_;
  assign new_n183_ = ~pe & new_n125_;
  assign new_n184_ = ~pm & new_n95_;
  assign new_n185_ = ~pq & ~pm;
  assign new_n186_ = ~pe & new_n185_;
  assign new_n187_ = ~new_n183_ & ~new_n184_;
  assign new_n188_ = ~new_n186_ & new_n187_;
  assign new_n189_ = ~pv & ~px;
  assign new_n190_ = ~pw & new_n189_;
  assign new_n191_ = py & new_n190_;
  assign new_n192_ = py & new_n188_;
  assign new_n193_ = ~new_n191_ & new_n192_;
  assign new_n194_ = ~pw & ~px;
  assign new_n195_ = ~pu & new_n194_;
  assign new_n196_ = new_n168_ & new_n195_;
  assign new_n197_ = new_n188_ & new_n196_;
  assign new_n198_ = pu & new_n197_;
  assign new_n199_ = pu & new_n192_;
  assign new_n200_ = pr & new_n192_;
  assign new_n201_ = ~pq & new_n188_;
  assign new_n202_ = pr & new_n197_;
  assign new_n203_ = ~new_n191_ & new_n197_;
  assign new_n204_ = ~new_n201_ & ~new_n202_;
  assign new_n205_ = ~new_n203_ & new_n204_;
  assign new_n206_ = ~new_n199_ & ~new_n200_;
  assign new_n207_ = ~new_n193_ & ~new_n198_;
  assign new_n208_ = new_n206_ & new_n207_;
  assign pq0 = ~new_n205_ | ~new_n208_;
  assign new_n210_ = ~pf & new_n125_;
  assign new_n211_ = ~pn & new_n95_;
  assign new_n212_ = ~pq & ~pn;
  assign new_n213_ = ~pf & new_n212_;
  assign new_n214_ = ~new_n210_ & ~new_n211_;
  assign new_n215_ = ~new_n213_ & new_n214_;
  assign new_n216_ = ~pw & ~py;
  assign new_n217_ = ~px & new_n216_;
  assign new_n218_ = pz & new_n217_;
  assign new_n219_ = pz & new_n215_;
  assign new_n220_ = ~new_n218_ & new_n219_;
  assign new_n221_ = ~py & new_n194_;
  assign new_n222_ = ~pu & new_n221_;
  assign new_n223_ = new_n168_ & new_n222_;
  assign new_n224_ = new_n215_ & new_n223_;
  assign new_n225_ = pr & new_n224_;
  assign new_n226_ = pr & new_n219_;
  assign new_n227_ = ~pu & ~pv;
  assign new_n228_ = new_n219_ & ~new_n227_;
  assign new_n229_ = ~pq & new_n215_;
  assign new_n230_ = new_n224_ & ~new_n227_;
  assign new_n231_ = ~new_n218_ & new_n224_;
  assign new_n232_ = ~new_n229_ & ~new_n230_;
  assign new_n233_ = ~new_n231_ & new_n232_;
  assign new_n234_ = ~new_n226_ & ~new_n228_;
  assign new_n235_ = ~new_n220_ & ~new_n225_;
  assign new_n236_ = new_n234_ & new_n235_;
  assign pr0 = ~new_n233_ | ~new_n236_;
  assign new_n238_ = ~pg & new_n125_;
  assign new_n239_ = ~po & new_n95_;
  assign new_n240_ = ~pq & ~po;
  assign new_n241_ = ~pg & new_n240_;
  assign new_n242_ = ~new_n238_ & ~new_n239_;
  assign new_n243_ = ~new_n241_ & new_n242_;
  assign new_n244_ = ~px & ~pz;
  assign new_n245_ = ~py & new_n244_;
  assign new_n246_ = pa0 & new_n245_;
  assign new_n247_ = pa0 & new_n243_;
  assign new_n248_ = ~new_n246_ & new_n247_;
  assign new_n249_ = ~pz & new_n217_;
  assign new_n250_ = ~pu & new_n249_;
  assign new_n251_ = new_n168_ & new_n250_;
  assign new_n252_ = new_n243_ & new_n251_;
  assign new_n253_ = pr & new_n252_;
  assign new_n254_ = pr & new_n247_;
  assign new_n255_ = ~pw & new_n227_;
  assign new_n256_ = new_n247_ & ~new_n255_;
  assign new_n257_ = ~pq & new_n243_;
  assign new_n258_ = new_n252_ & ~new_n255_;
  assign new_n259_ = ~new_n246_ & new_n252_;
  assign new_n260_ = ~new_n257_ & ~new_n258_;
  assign new_n261_ = ~new_n259_ & new_n260_;
  assign new_n262_ = ~new_n254_ & ~new_n256_;
  assign new_n263_ = ~new_n248_ & ~new_n253_;
  assign new_n264_ = new_n262_ & new_n263_;
  assign ps0 = ~new_n261_ | ~new_n264_;
  assign new_n266_ = ~ph & new_n125_;
  assign new_n267_ = ~pp & new_n95_;
  assign new_n268_ = ~pp & ~pq;
  assign new_n269_ = ~ph & new_n268_;
  assign new_n270_ = ~new_n266_ & ~new_n267_;
  assign new_n271_ = ~new_n269_ & new_n270_;
  assign new_n272_ = ~pa0 & ~py;
  assign new_n273_ = ~pz & new_n272_;
  assign new_n274_ = pb0 & new_n273_;
  assign new_n275_ = pb0 & new_n271_;
  assign new_n276_ = ~new_n274_ & new_n275_;
  assign new_n277_ = ~pa0 & new_n245_;
  assign new_n278_ = ~pu & new_n163_;
  assign new_n279_ = ~pr & new_n277_;
  assign new_n280_ = new_n278_ & new_n279_;
  assign new_n281_ = new_n271_ & new_n280_;
  assign new_n282_ = pr & new_n281_;
  assign new_n283_ = pr & new_n275_;
  assign new_n284_ = ~pv & new_n167_;
  assign new_n285_ = ~px & new_n284_;
  assign new_n286_ = new_n275_ & ~new_n285_;
  assign new_n287_ = ~pq & new_n271_;
  assign new_n288_ = new_n281_ & ~new_n285_;
  assign new_n289_ = ~new_n274_ & new_n281_;
  assign new_n290_ = ~new_n287_ & ~new_n288_;
  assign new_n291_ = ~new_n289_ & new_n290_;
  assign new_n292_ = ~new_n283_ & ~new_n286_;
  assign new_n293_ = ~new_n276_ & ~new_n282_;
  assign new_n294_ = new_n292_ & new_n293_;
  assign pt0 = ~new_n291_ | ~new_n294_;
  assign new_n296_ = ~pb0 & ~pz;
  assign new_n297_ = new_n272_ & new_n296_;
  assign new_n298_ = pu & ~pw;
  assign new_n299_ = new_n189_ & new_n298_;
  assign new_n300_ = ~pr & new_n297_;
  assign new_n301_ = new_n299_ & new_n300_;
  assign new_n302_ = pq & new_n301_;
  assign new_n303_ = pr & pc0;
  assign new_n304_ = pq & new_n303_;
  assign pu0 = new_n302_ | new_n304_;
  assign pl0 = pc0;
endmodule

