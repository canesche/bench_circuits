// Benchmark "testing" written by ABC on Thu Oct  8 22:16:45 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A107  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A107;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[168]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[177]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[187]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[196]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[207]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[216]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[226]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[236]_ , \new_[237]_ , \new_[241]_ ,
    \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ , \new_[246]_ ,
    \new_[249]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ , \new_[258]_ ,
    \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ , \new_[268]_ ,
    \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[277]_ , \new_[281]_ ,
    \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ , \new_[288]_ ,
    \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[297]_ , \new_[301]_ ,
    \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[307]_ , \new_[311]_ ,
    \new_[312]_ , \new_[313]_ , \new_[317]_ , \new_[318]_ , \new_[322]_ ,
    \new_[323]_ , \new_[324]_ , \new_[325]_ , \new_[326]_ , \new_[327]_ ,
    \new_[328]_ , \new_[331]_ , \new_[335]_ , \new_[336]_ , \new_[337]_ ,
    \new_[340]_ , \new_[344]_ , \new_[345]_ , \new_[346]_ , \new_[347]_ ,
    \new_[350]_ , \new_[354]_ , \new_[355]_ , \new_[356]_ , \new_[359]_ ,
    \new_[363]_ , \new_[364]_ , \new_[365]_ , \new_[366]_ , \new_[367]_ ,
    \new_[370]_ , \new_[374]_ , \new_[375]_ , \new_[376]_ , \new_[379]_ ,
    \new_[383]_ , \new_[384]_ , \new_[385]_ , \new_[386]_ , \new_[389]_ ,
    \new_[393]_ , \new_[394]_ , \new_[395]_ , \new_[399]_ , \new_[400]_ ,
    \new_[404]_ , \new_[405]_ , \new_[406]_ , \new_[407]_ , \new_[408]_ ,
    \new_[409]_ , \new_[412]_ , \new_[416]_ , \new_[417]_ , \new_[418]_ ,
    \new_[421]_ , \new_[425]_ , \new_[426]_ , \new_[427]_ , \new_[428]_ ,
    \new_[431]_ , \new_[435]_ , \new_[436]_ , \new_[437]_ , \new_[441]_ ,
    \new_[442]_ , \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ ,
    \new_[450]_ , \new_[453]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ ,
    \new_[462]_ , \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ ,
    \new_[472]_ , \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[482]_ ,
    \new_[483]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[498]_ , \new_[501]_ ,
    \new_[504]_ , \new_[507]_ , \new_[510]_ , \new_[513]_ , \new_[516]_ ,
    \new_[519]_ , \new_[522]_ , \new_[525]_ , \new_[529]_ , \new_[530]_ ,
    \new_[534]_ , \new_[535]_ , \new_[539]_ , \new_[540]_ , \new_[544]_ ,
    \new_[545]_ , \new_[549]_ , \new_[550]_ , \new_[554]_ , \new_[555]_ ,
    \new_[559]_ , \new_[560]_ , \new_[564]_ , \new_[565]_ , \new_[569]_ ,
    \new_[570]_ , \new_[574]_ , \new_[575]_ , \new_[579]_ , \new_[580]_ ,
    \new_[584]_ , \new_[585]_ , \new_[589]_ , \new_[590]_ , \new_[594]_ ,
    \new_[595]_ , \new_[599]_ , \new_[600]_ , \new_[604]_ , \new_[605]_ ,
    \new_[609]_ , \new_[610]_ , \new_[614]_ , \new_[615]_ , \new_[619]_ ,
    \new_[620]_ , \new_[624]_ , \new_[625]_ , \new_[629]_ , \new_[630]_ ,
    \new_[634]_ , \new_[635]_ , \new_[639]_ , \new_[640]_ , \new_[644]_ ,
    \new_[645]_ , \new_[649]_ , \new_[650]_ , \new_[654]_ , \new_[655]_ ,
    \new_[659]_ , \new_[660]_ , \new_[664]_ , \new_[665]_ , \new_[669]_ ,
    \new_[670]_ , \new_[674]_ , \new_[675]_ , \new_[679]_ , \new_[680]_ ,
    \new_[684]_ , \new_[685]_ , \new_[689]_ , \new_[690]_ , \new_[694]_ ,
    \new_[695]_ , \new_[699]_ , \new_[700]_ , \new_[704]_ , \new_[705]_ ,
    \new_[709]_ , \new_[710]_ , \new_[713]_ , \new_[716]_ , \new_[717]_ ,
    \new_[721]_ , \new_[722]_ , \new_[725]_ , \new_[728]_ , \new_[729]_ ,
    \new_[733]_ , \new_[734]_ , \new_[737]_ , \new_[740]_ , \new_[741]_ ,
    \new_[745]_ , \new_[746]_ , \new_[749]_ , \new_[752]_ , \new_[753]_ ,
    \new_[757]_ , \new_[758]_ , \new_[761]_ , \new_[764]_ , \new_[765]_ ,
    \new_[769]_ , \new_[770]_ , \new_[773]_ , \new_[776]_ , \new_[777]_ ,
    \new_[780]_ , \new_[783]_ , \new_[784]_ , \new_[787]_ , \new_[790]_ ,
    \new_[791]_ , \new_[794]_ , \new_[797]_ , \new_[798]_ , \new_[801]_ ,
    \new_[804]_ , \new_[805]_ , \new_[808]_ , \new_[811]_ , \new_[812]_ ,
    \new_[815]_ , \new_[818]_ , \new_[819]_ , \new_[822]_ , \new_[825]_ ,
    \new_[826]_ , \new_[829]_ , \new_[832]_ , \new_[833]_ , \new_[836]_ ,
    \new_[839]_ , \new_[840]_ , \new_[843]_ , \new_[846]_ , \new_[847]_ ,
    \new_[850]_ , \new_[853]_ , \new_[854]_ , \new_[857]_ , \new_[860]_ ,
    \new_[861]_ , \new_[864]_ , \new_[867]_ , \new_[868]_ , \new_[871]_ ,
    \new_[874]_ , \new_[875]_ , \new_[878]_ , \new_[881]_ , \new_[882]_ ,
    \new_[885]_ , \new_[888]_ , \new_[889]_ , \new_[892]_ , \new_[895]_ ,
    \new_[896]_ , \new_[899]_ , \new_[902]_ , \new_[903]_ , \new_[906]_ ,
    \new_[909]_ , \new_[910]_ , \new_[913]_ , \new_[916]_ , \new_[917]_ ,
    \new_[920]_ , \new_[923]_ , \new_[924]_ , \new_[927]_ , \new_[930]_ ,
    \new_[931]_ , \new_[934]_ , \new_[937]_ , \new_[938]_ , \new_[941]_ ,
    \new_[944]_ , \new_[945]_ , \new_[948]_ , \new_[951]_ , \new_[952]_ ,
    \new_[955]_ , \new_[958]_ , \new_[959]_ , \new_[962]_ , \new_[965]_ ,
    \new_[966]_ , \new_[969]_ , \new_[972]_ , \new_[973]_ , \new_[976]_ ,
    \new_[979]_ , \new_[980]_ , \new_[983]_ , \new_[986]_ , \new_[987]_ ,
    \new_[990]_ , \new_[993]_ , \new_[994]_ , \new_[997]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1004]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1011]_ , \new_[1014]_ , \new_[1015]_ , \new_[1018]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1025]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1032]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1039]_ , \new_[1042]_ , \new_[1043]_ , \new_[1046]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1053]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1060]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1067]_ , \new_[1070]_ , \new_[1071]_ , \new_[1074]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1081]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1088]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1095]_ , \new_[1098]_ , \new_[1099]_ , \new_[1102]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1109]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1116]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1123]_ , \new_[1126]_ , \new_[1127]_ , \new_[1130]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1137]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1144]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1151]_ , \new_[1154]_ , \new_[1155]_ , \new_[1158]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1165]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1172]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1179]_ , \new_[1182]_ , \new_[1183]_ , \new_[1186]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1193]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1200]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1207]_ , \new_[1210]_ , \new_[1211]_ , \new_[1214]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1221]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1228]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1235]_ , \new_[1238]_ , \new_[1239]_ , \new_[1242]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1249]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1256]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1263]_ , \new_[1266]_ , \new_[1267]_ , \new_[1270]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1277]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1284]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1291]_ , \new_[1294]_ , \new_[1295]_ , \new_[1298]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1305]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1312]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1319]_ , \new_[1322]_ , \new_[1323]_ , \new_[1326]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1333]_ , \new_[1337]_ ,
    \new_[1338]_ , \new_[1339]_ , \new_[1342]_ , \new_[1345]_ ,
    \new_[1346]_ , \new_[1349]_ , \new_[1353]_ , \new_[1354]_ ,
    \new_[1355]_ , \new_[1358]_ , \new_[1361]_ , \new_[1362]_ ,
    \new_[1365]_ , \new_[1369]_ , \new_[1370]_ , \new_[1371]_ ,
    \new_[1374]_ , \new_[1377]_ , \new_[1378]_ , \new_[1381]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1390]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1397]_ , \new_[1401]_ ,
    \new_[1402]_ , \new_[1403]_ , \new_[1406]_ , \new_[1409]_ ,
    \new_[1410]_ , \new_[1413]_ , \new_[1417]_ , \new_[1418]_ ,
    \new_[1419]_ , \new_[1422]_ , \new_[1425]_ , \new_[1426]_ ,
    \new_[1429]_ , \new_[1433]_ , \new_[1434]_ , \new_[1435]_ ,
    \new_[1438]_ , \new_[1441]_ , \new_[1442]_ , \new_[1445]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1454]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1461]_ , \new_[1465]_ ,
    \new_[1466]_ , \new_[1467]_ , \new_[1470]_ , \new_[1473]_ ,
    \new_[1474]_ , \new_[1477]_ , \new_[1481]_ , \new_[1482]_ ,
    \new_[1483]_ , \new_[1486]_ , \new_[1489]_ , \new_[1490]_ ,
    \new_[1493]_ , \new_[1497]_ , \new_[1498]_ , \new_[1499]_ ,
    \new_[1502]_ , \new_[1505]_ , \new_[1506]_ , \new_[1509]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1518]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1525]_ , \new_[1529]_ ,
    \new_[1530]_ , \new_[1531]_ , \new_[1534]_ , \new_[1537]_ ,
    \new_[1538]_ , \new_[1541]_ , \new_[1545]_ , \new_[1546]_ ,
    \new_[1547]_ , \new_[1550]_ , \new_[1553]_ , \new_[1554]_ ,
    \new_[1557]_ , \new_[1561]_ , \new_[1562]_ , \new_[1563]_ ,
    \new_[1566]_ , \new_[1569]_ , \new_[1570]_ , \new_[1573]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1582]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1589]_ , \new_[1593]_ ,
    \new_[1594]_ , \new_[1595]_ , \new_[1598]_ , \new_[1601]_ ,
    \new_[1602]_ , \new_[1605]_ , \new_[1609]_ , \new_[1610]_ ,
    \new_[1611]_ , \new_[1614]_ , \new_[1617]_ , \new_[1618]_ ,
    \new_[1621]_ , \new_[1625]_ , \new_[1626]_ , \new_[1627]_ ,
    \new_[1630]_ , \new_[1633]_ , \new_[1634]_ , \new_[1637]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1646]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1653]_ , \new_[1657]_ ,
    \new_[1658]_ , \new_[1659]_ , \new_[1662]_ , \new_[1665]_ ,
    \new_[1666]_ , \new_[1669]_ , \new_[1673]_ , \new_[1674]_ ,
    \new_[1675]_ , \new_[1678]_ , \new_[1681]_ , \new_[1682]_ ,
    \new_[1685]_ , \new_[1689]_ , \new_[1690]_ , \new_[1691]_ ,
    \new_[1694]_ , \new_[1697]_ , \new_[1698]_ , \new_[1701]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1710]_ ,
    \new_[1714]_ , \new_[1715]_ , \new_[1716]_ , \new_[1719]_ ,
    \new_[1723]_ , \new_[1724]_ , \new_[1725]_ , \new_[1728]_ ,
    \new_[1732]_ , \new_[1733]_ , \new_[1734]_ , \new_[1737]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1746]_ ,
    \new_[1750]_ , \new_[1751]_ , \new_[1752]_ , \new_[1755]_ ,
    \new_[1759]_ , \new_[1760]_ , \new_[1761]_ , \new_[1764]_ ,
    \new_[1768]_ , \new_[1769]_ , \new_[1770]_ , \new_[1773]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1782]_ ,
    \new_[1786]_ , \new_[1787]_ , \new_[1788]_ , \new_[1791]_ ,
    \new_[1795]_ , \new_[1796]_ , \new_[1797]_ , \new_[1800]_ ,
    \new_[1804]_ , \new_[1805]_ , \new_[1806]_ , \new_[1809]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1818]_ ,
    \new_[1822]_ , \new_[1823]_ , \new_[1824]_ , \new_[1827]_ ,
    \new_[1831]_ , \new_[1832]_ , \new_[1833]_ , \new_[1836]_ ,
    \new_[1840]_ , \new_[1841]_ , \new_[1842]_ , \new_[1845]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1854]_ ,
    \new_[1858]_ , \new_[1859]_ , \new_[1860]_ , \new_[1863]_ ,
    \new_[1867]_ , \new_[1868]_ , \new_[1869]_ , \new_[1872]_ ,
    \new_[1876]_ , \new_[1877]_ , \new_[1878]_ , \new_[1881]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1890]_ ,
    \new_[1894]_ , \new_[1895]_ , \new_[1896]_ , \new_[1899]_ ,
    \new_[1903]_ , \new_[1904]_ , \new_[1905]_ , \new_[1908]_ ,
    \new_[1912]_ , \new_[1913]_ , \new_[1914]_ , \new_[1917]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1926]_ ,
    \new_[1930]_ , \new_[1931]_ , \new_[1932]_ , \new_[1935]_ ,
    \new_[1939]_ , \new_[1940]_ , \new_[1941]_ , \new_[1944]_ ,
    \new_[1948]_ , \new_[1949]_ , \new_[1950]_ , \new_[1953]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1962]_ ,
    \new_[1966]_ , \new_[1967]_ , \new_[1968]_ , \new_[1971]_ ,
    \new_[1975]_ , \new_[1976]_ , \new_[1977]_ , \new_[1980]_ ,
    \new_[1984]_ , \new_[1985]_ , \new_[1986]_ , \new_[1989]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1998]_ ,
    \new_[2002]_ , \new_[2003]_ , \new_[2004]_ , \new_[2007]_ ,
    \new_[2011]_ , \new_[2012]_ , \new_[2013]_ , \new_[2016]_ ,
    \new_[2020]_ , \new_[2021]_ , \new_[2022]_ , \new_[2025]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2034]_ ,
    \new_[2038]_ , \new_[2039]_ , \new_[2040]_ , \new_[2043]_ ,
    \new_[2047]_ , \new_[2048]_ , \new_[2049]_ , \new_[2052]_ ,
    \new_[2056]_ , \new_[2057]_ , \new_[2058]_ , \new_[2061]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2070]_ ,
    \new_[2074]_ , \new_[2075]_ , \new_[2076]_ , \new_[2079]_ ,
    \new_[2083]_ , \new_[2084]_ , \new_[2085]_ , \new_[2088]_ ,
    \new_[2092]_ , \new_[2093]_ , \new_[2094]_ , \new_[2097]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2106]_ ,
    \new_[2110]_ , \new_[2111]_ , \new_[2112]_ , \new_[2115]_ ,
    \new_[2119]_ , \new_[2120]_ , \new_[2121]_ , \new_[2124]_ ,
    \new_[2128]_ , \new_[2129]_ , \new_[2130]_ , \new_[2133]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2142]_ ,
    \new_[2146]_ , \new_[2147]_ , \new_[2148]_ , \new_[2151]_ ,
    \new_[2155]_ , \new_[2156]_ , \new_[2157]_ , \new_[2160]_ ,
    \new_[2164]_ , \new_[2165]_ , \new_[2166]_ , \new_[2169]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2178]_ ,
    \new_[2182]_ , \new_[2183]_ , \new_[2184]_ , \new_[2187]_ ,
    \new_[2191]_ , \new_[2192]_ , \new_[2193]_ , \new_[2196]_ ,
    \new_[2200]_ , \new_[2201]_ , \new_[2202]_ , \new_[2205]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2214]_ ,
    \new_[2218]_ , \new_[2219]_ , \new_[2220]_ , \new_[2223]_ ,
    \new_[2227]_ , \new_[2228]_ , \new_[2229]_ , \new_[2232]_ ,
    \new_[2236]_ , \new_[2237]_ , \new_[2238]_ , \new_[2241]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2250]_ ,
    \new_[2254]_ , \new_[2255]_ , \new_[2256]_ , \new_[2259]_ ,
    \new_[2263]_ , \new_[2264]_ , \new_[2265]_ , \new_[2268]_ ,
    \new_[2272]_ , \new_[2273]_ , \new_[2274]_ , \new_[2277]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2286]_ ,
    \new_[2290]_ , \new_[2291]_ , \new_[2292]_ , \new_[2295]_ ,
    \new_[2299]_ , \new_[2300]_ , \new_[2301]_ , \new_[2304]_ ,
    \new_[2308]_ , \new_[2309]_ , \new_[2310]_ , \new_[2313]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2322]_ ,
    \new_[2326]_ , \new_[2327]_ , \new_[2328]_ , \new_[2331]_ ,
    \new_[2335]_ , \new_[2336]_ , \new_[2337]_ , \new_[2340]_ ,
    \new_[2344]_ , \new_[2345]_ , \new_[2346]_ , \new_[2349]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2358]_ ,
    \new_[2362]_ , \new_[2363]_ , \new_[2364]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2373]_ , \new_[2374]_ , \new_[2375]_ ,
    \new_[2378]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2388]_ , \new_[2389]_ , \new_[2393]_ , \new_[2394]_ ,
    \new_[2395]_ , \new_[2398]_ , \new_[2402]_ , \new_[2403]_ ,
    \new_[2404]_ , \new_[2408]_ , \new_[2409]_ , \new_[2413]_ ,
    \new_[2414]_ , \new_[2415]_ , \new_[2418]_ , \new_[2422]_ ,
    \new_[2423]_ , \new_[2424]_ , \new_[2428]_ , \new_[2429]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2438]_ ,
    \new_[2442]_ , \new_[2443]_ , \new_[2444]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2453]_ , \new_[2454]_ , \new_[2455]_ ,
    \new_[2458]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2468]_ , \new_[2469]_ , \new_[2473]_ , \new_[2474]_ ,
    \new_[2475]_ , \new_[2478]_ , \new_[2482]_ , \new_[2483]_ ,
    \new_[2484]_ , \new_[2488]_ , \new_[2489]_ , \new_[2493]_ ,
    \new_[2494]_ , \new_[2495]_ , \new_[2498]_ , \new_[2502]_ ,
    \new_[2503]_ , \new_[2504]_ , \new_[2508]_ , \new_[2509]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2518]_ ,
    \new_[2522]_ , \new_[2523]_ , \new_[2524]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2533]_ , \new_[2534]_ , \new_[2535]_ ,
    \new_[2538]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2548]_ , \new_[2549]_ , \new_[2553]_ , \new_[2554]_ ,
    \new_[2555]_ , \new_[2558]_ , \new_[2562]_ , \new_[2563]_ ,
    \new_[2564]_ , \new_[2568]_ , \new_[2569]_ , \new_[2573]_ ,
    \new_[2574]_ , \new_[2575]_ , \new_[2578]_ , \new_[2582]_ ,
    \new_[2583]_ , \new_[2584]_ , \new_[2588]_ , \new_[2589]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2598]_ ,
    \new_[2602]_ , \new_[2603]_ , \new_[2604]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2613]_ , \new_[2614]_ , \new_[2615]_ ,
    \new_[2618]_ , \new_[2622]_ , \new_[2623]_ , \new_[2624]_ ,
    \new_[2628]_ , \new_[2629]_ , \new_[2633]_ , \new_[2634]_ ,
    \new_[2635]_ , \new_[2638]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2648]_ , \new_[2649]_ , \new_[2653]_ ,
    \new_[2654]_ , \new_[2655]_ , \new_[2658]_ , \new_[2662]_ ,
    \new_[2663]_ , \new_[2664]_ , \new_[2668]_ , \new_[2669]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2678]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2693]_ , \new_[2694]_ , \new_[2695]_ ,
    \new_[2698]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2708]_ , \new_[2709]_ , \new_[2713]_ , \new_[2714]_ ,
    \new_[2715]_ , \new_[2718]_ , \new_[2722]_ , \new_[2723]_ ,
    \new_[2724]_ , \new_[2728]_ , \new_[2729]_ , \new_[2733]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2738]_ , \new_[2742]_ ,
    \new_[2743]_ , \new_[2744]_ , \new_[2748]_ , \new_[2749]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2758]_ ,
    \new_[2762]_ , \new_[2763]_ , \new_[2764]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2773]_ , \new_[2774]_ , \new_[2775]_ ,
    \new_[2778]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2788]_ , \new_[2789]_ , \new_[2793]_ , \new_[2794]_ ,
    \new_[2795]_ , \new_[2798]_ , \new_[2802]_ , \new_[2803]_ ,
    \new_[2804]_ , \new_[2808]_ , \new_[2809]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2815]_ , \new_[2818]_ , \new_[2822]_ ,
    \new_[2823]_ , \new_[2824]_ , \new_[2828]_ , \new_[2829]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2839]_ ,
    \new_[2840]_ , \new_[2844]_ , \new_[2845]_ , \new_[2846]_ ,
    \new_[2850]_ , \new_[2851]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2861]_ , \new_[2862]_ , \new_[2866]_ ,
    \new_[2867]_ , \new_[2868]_ , \new_[2872]_ , \new_[2873]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2883]_ ,
    \new_[2884]_ , \new_[2888]_ , \new_[2889]_ , \new_[2890]_ ,
    \new_[2894]_ , \new_[2895]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2905]_ , \new_[2906]_ , \new_[2910]_ ,
    \new_[2911]_ , \new_[2912]_ , \new_[2916]_ , \new_[2917]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2927]_ ,
    \new_[2928]_ , \new_[2932]_ , \new_[2933]_ , \new_[2934]_ ,
    \new_[2938]_ , \new_[2939]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2949]_ , \new_[2950]_ , \new_[2954]_ ,
    \new_[2955]_ , \new_[2956]_ , \new_[2960]_ , \new_[2961]_ ,
    \new_[2965]_ , \new_[2966]_ , \new_[2967]_ , \new_[2971]_ ,
    \new_[2972]_ , \new_[2976]_ , \new_[2977]_ , \new_[2978]_ ,
    \new_[2982]_ , \new_[2983]_ , \new_[2987]_ , \new_[2988]_ ,
    \new_[2989]_ , \new_[2993]_ , \new_[2994]_ , \new_[2998]_ ,
    \new_[2999]_ , \new_[3000]_ , \new_[3004]_ , \new_[3005]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3011]_ , \new_[3015]_ ,
    \new_[3016]_ , \new_[3020]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3026]_ , \new_[3027]_ , \new_[3031]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3037]_ , \new_[3038]_ , \new_[3042]_ ,
    \new_[3043]_ , \new_[3044]_ , \new_[3048]_ , \new_[3049]_ ,
    \new_[3053]_ , \new_[3054]_ , \new_[3055]_ , \new_[3059]_ ,
    \new_[3060]_ , \new_[3064]_ , \new_[3065]_ , \new_[3066]_ ,
    \new_[3070]_ , \new_[3071]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3081]_ , \new_[3082]_ , \new_[3086]_ ,
    \new_[3087]_ , \new_[3088]_ , \new_[3092]_ , \new_[3093]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ;
  assign A107 = \new_[493]_  | \new_[328]_ ;
  assign \new_[1]_  = \new_[3099]_  & \new_[3088]_ ;
  assign \new_[2]_  = \new_[3077]_  & \new_[3066]_ ;
  assign \new_[3]_  = \new_[3055]_  & \new_[3044]_ ;
  assign \new_[4]_  = \new_[3033]_  & \new_[3022]_ ;
  assign \new_[5]_  = \new_[3011]_  & \new_[3000]_ ;
  assign \new_[6]_  = \new_[2989]_  & \new_[2978]_ ;
  assign \new_[7]_  = \new_[2967]_  & \new_[2956]_ ;
  assign \new_[8]_  = \new_[2945]_  & \new_[2934]_ ;
  assign \new_[9]_  = \new_[2923]_  & \new_[2912]_ ;
  assign \new_[10]_  = \new_[2901]_  & \new_[2890]_ ;
  assign \new_[11]_  = \new_[2879]_  & \new_[2868]_ ;
  assign \new_[12]_  = \new_[2857]_  & \new_[2846]_ ;
  assign \new_[13]_  = \new_[2835]_  & \new_[2824]_ ;
  assign \new_[14]_  = \new_[2815]_  & \new_[2804]_ ;
  assign \new_[15]_  = \new_[2795]_  & \new_[2784]_ ;
  assign \new_[16]_  = \new_[2775]_  & \new_[2764]_ ;
  assign \new_[17]_  = \new_[2755]_  & \new_[2744]_ ;
  assign \new_[18]_  = \new_[2735]_  & \new_[2724]_ ;
  assign \new_[19]_  = \new_[2715]_  & \new_[2704]_ ;
  assign \new_[20]_  = \new_[2695]_  & \new_[2684]_ ;
  assign \new_[21]_  = \new_[2675]_  & \new_[2664]_ ;
  assign \new_[22]_  = \new_[2655]_  & \new_[2644]_ ;
  assign \new_[23]_  = \new_[2635]_  & \new_[2624]_ ;
  assign \new_[24]_  = \new_[2615]_  & \new_[2604]_ ;
  assign \new_[25]_  = \new_[2595]_  & \new_[2584]_ ;
  assign \new_[26]_  = \new_[2575]_  & \new_[2564]_ ;
  assign \new_[27]_  = \new_[2555]_  & \new_[2544]_ ;
  assign \new_[28]_  = \new_[2535]_  & \new_[2524]_ ;
  assign \new_[29]_  = \new_[2515]_  & \new_[2504]_ ;
  assign \new_[30]_  = \new_[2495]_  & \new_[2484]_ ;
  assign \new_[31]_  = \new_[2475]_  & \new_[2464]_ ;
  assign \new_[32]_  = \new_[2455]_  & \new_[2444]_ ;
  assign \new_[33]_  = \new_[2435]_  & \new_[2424]_ ;
  assign \new_[34]_  = \new_[2415]_  & \new_[2404]_ ;
  assign \new_[35]_  = \new_[2395]_  & \new_[2384]_ ;
  assign \new_[36]_  = \new_[2375]_  & \new_[2364]_ ;
  assign \new_[37]_  = \new_[2355]_  & \new_[2346]_ ;
  assign \new_[38]_  = \new_[2337]_  & \new_[2328]_ ;
  assign \new_[39]_  = \new_[2319]_  & \new_[2310]_ ;
  assign \new_[40]_  = \new_[2301]_  & \new_[2292]_ ;
  assign \new_[41]_  = \new_[2283]_  & \new_[2274]_ ;
  assign \new_[42]_  = \new_[2265]_  & \new_[2256]_ ;
  assign \new_[43]_  = \new_[2247]_  & \new_[2238]_ ;
  assign \new_[44]_  = \new_[2229]_  & \new_[2220]_ ;
  assign \new_[45]_  = \new_[2211]_  & \new_[2202]_ ;
  assign \new_[46]_  = \new_[2193]_  & \new_[2184]_ ;
  assign \new_[47]_  = \new_[2175]_  & \new_[2166]_ ;
  assign \new_[48]_  = \new_[2157]_  & \new_[2148]_ ;
  assign \new_[49]_  = \new_[2139]_  & \new_[2130]_ ;
  assign \new_[50]_  = \new_[2121]_  & \new_[2112]_ ;
  assign \new_[51]_  = \new_[2103]_  & \new_[2094]_ ;
  assign \new_[52]_  = \new_[2085]_  & \new_[2076]_ ;
  assign \new_[53]_  = \new_[2067]_  & \new_[2058]_ ;
  assign \new_[54]_  = \new_[2049]_  & \new_[2040]_ ;
  assign \new_[55]_  = \new_[2031]_  & \new_[2022]_ ;
  assign \new_[56]_  = \new_[2013]_  & \new_[2004]_ ;
  assign \new_[57]_  = \new_[1995]_  & \new_[1986]_ ;
  assign \new_[58]_  = \new_[1977]_  & \new_[1968]_ ;
  assign \new_[59]_  = \new_[1959]_  & \new_[1950]_ ;
  assign \new_[60]_  = \new_[1941]_  & \new_[1932]_ ;
  assign \new_[61]_  = \new_[1923]_  & \new_[1914]_ ;
  assign \new_[62]_  = \new_[1905]_  & \new_[1896]_ ;
  assign \new_[63]_  = \new_[1887]_  & \new_[1878]_ ;
  assign \new_[64]_  = \new_[1869]_  & \new_[1860]_ ;
  assign \new_[65]_  = \new_[1851]_  & \new_[1842]_ ;
  assign \new_[66]_  = \new_[1833]_  & \new_[1824]_ ;
  assign \new_[67]_  = \new_[1815]_  & \new_[1806]_ ;
  assign \new_[68]_  = \new_[1797]_  & \new_[1788]_ ;
  assign \new_[69]_  = \new_[1779]_  & \new_[1770]_ ;
  assign \new_[70]_  = \new_[1761]_  & \new_[1752]_ ;
  assign \new_[71]_  = \new_[1743]_  & \new_[1734]_ ;
  assign \new_[72]_  = \new_[1725]_  & \new_[1716]_ ;
  assign \new_[73]_  = \new_[1707]_  & \new_[1698]_ ;
  assign \new_[74]_  = \new_[1691]_  & \new_[1682]_ ;
  assign \new_[75]_  = \new_[1675]_  & \new_[1666]_ ;
  assign \new_[76]_  = \new_[1659]_  & \new_[1650]_ ;
  assign \new_[77]_  = \new_[1643]_  & \new_[1634]_ ;
  assign \new_[78]_  = \new_[1627]_  & \new_[1618]_ ;
  assign \new_[79]_  = \new_[1611]_  & \new_[1602]_ ;
  assign \new_[80]_  = \new_[1595]_  & \new_[1586]_ ;
  assign \new_[81]_  = \new_[1579]_  & \new_[1570]_ ;
  assign \new_[82]_  = \new_[1563]_  & \new_[1554]_ ;
  assign \new_[83]_  = \new_[1547]_  & \new_[1538]_ ;
  assign \new_[84]_  = \new_[1531]_  & \new_[1522]_ ;
  assign \new_[85]_  = \new_[1515]_  & \new_[1506]_ ;
  assign \new_[86]_  = \new_[1499]_  & \new_[1490]_ ;
  assign \new_[87]_  = \new_[1483]_  & \new_[1474]_ ;
  assign \new_[88]_  = \new_[1467]_  & \new_[1458]_ ;
  assign \new_[89]_  = \new_[1451]_  & \new_[1442]_ ;
  assign \new_[90]_  = \new_[1435]_  & \new_[1426]_ ;
  assign \new_[91]_  = \new_[1419]_  & \new_[1410]_ ;
  assign \new_[92]_  = \new_[1403]_  & \new_[1394]_ ;
  assign \new_[93]_  = \new_[1387]_  & \new_[1378]_ ;
  assign \new_[94]_  = \new_[1371]_  & \new_[1362]_ ;
  assign \new_[95]_  = \new_[1355]_  & \new_[1346]_ ;
  assign \new_[96]_  = \new_[1339]_  & \new_[1330]_ ;
  assign \new_[97]_  = \new_[1323]_  & \new_[1316]_ ;
  assign \new_[98]_  = \new_[1309]_  & \new_[1302]_ ;
  assign \new_[99]_  = \new_[1295]_  & \new_[1288]_ ;
  assign \new_[100]_  = \new_[1281]_  & \new_[1274]_ ;
  assign \new_[101]_  = \new_[1267]_  & \new_[1260]_ ;
  assign \new_[102]_  = \new_[1253]_  & \new_[1246]_ ;
  assign \new_[103]_  = \new_[1239]_  & \new_[1232]_ ;
  assign \new_[104]_  = \new_[1225]_  & \new_[1218]_ ;
  assign \new_[105]_  = \new_[1211]_  & \new_[1204]_ ;
  assign \new_[106]_  = \new_[1197]_  & \new_[1190]_ ;
  assign \new_[107]_  = \new_[1183]_  & \new_[1176]_ ;
  assign \new_[108]_  = \new_[1169]_  & \new_[1162]_ ;
  assign \new_[109]_  = \new_[1155]_  & \new_[1148]_ ;
  assign \new_[110]_  = \new_[1141]_  & \new_[1134]_ ;
  assign \new_[111]_  = \new_[1127]_  & \new_[1120]_ ;
  assign \new_[112]_  = \new_[1113]_  & \new_[1106]_ ;
  assign \new_[113]_  = \new_[1099]_  & \new_[1092]_ ;
  assign \new_[114]_  = \new_[1085]_  & \new_[1078]_ ;
  assign \new_[115]_  = \new_[1071]_  & \new_[1064]_ ;
  assign \new_[116]_  = \new_[1057]_  & \new_[1050]_ ;
  assign \new_[117]_  = \new_[1043]_  & \new_[1036]_ ;
  assign \new_[118]_  = \new_[1029]_  & \new_[1022]_ ;
  assign \new_[119]_  = \new_[1015]_  & \new_[1008]_ ;
  assign \new_[120]_  = \new_[1001]_  & \new_[994]_ ;
  assign \new_[121]_  = \new_[987]_  & \new_[980]_ ;
  assign \new_[122]_  = \new_[973]_  & \new_[966]_ ;
  assign \new_[123]_  = \new_[959]_  & \new_[952]_ ;
  assign \new_[124]_  = \new_[945]_  & \new_[938]_ ;
  assign \new_[125]_  = \new_[931]_  & \new_[924]_ ;
  assign \new_[126]_  = \new_[917]_  & \new_[910]_ ;
  assign \new_[127]_  = \new_[903]_  & \new_[896]_ ;
  assign \new_[128]_  = \new_[889]_  & \new_[882]_ ;
  assign \new_[129]_  = \new_[875]_  & \new_[868]_ ;
  assign \new_[130]_  = \new_[861]_  & \new_[854]_ ;
  assign \new_[131]_  = \new_[847]_  & \new_[840]_ ;
  assign \new_[132]_  = \new_[833]_  & \new_[826]_ ;
  assign \new_[133]_  = \new_[819]_  & \new_[812]_ ;
  assign \new_[134]_  = \new_[805]_  & \new_[798]_ ;
  assign \new_[135]_  = \new_[791]_  & \new_[784]_ ;
  assign \new_[136]_  = \new_[777]_  & \new_[770]_ ;
  assign \new_[137]_  = \new_[765]_  & \new_[758]_ ;
  assign \new_[138]_  = \new_[753]_  & \new_[746]_ ;
  assign \new_[139]_  = \new_[741]_  & \new_[734]_ ;
  assign \new_[140]_  = \new_[729]_  & \new_[722]_ ;
  assign \new_[141]_  = \new_[717]_  & \new_[710]_ ;
  assign \new_[142]_  = \new_[705]_  & \new_[700]_ ;
  assign \new_[143]_  = \new_[695]_  & \new_[690]_ ;
  assign \new_[144]_  = \new_[685]_  & \new_[680]_ ;
  assign \new_[145]_  = \new_[675]_  & \new_[670]_ ;
  assign \new_[146]_  = \new_[665]_  & \new_[660]_ ;
  assign \new_[147]_  = \new_[655]_  & \new_[650]_ ;
  assign \new_[148]_  = \new_[645]_  & \new_[640]_ ;
  assign \new_[149]_  = \new_[635]_  & \new_[630]_ ;
  assign \new_[150]_  = \new_[625]_  & \new_[620]_ ;
  assign \new_[151]_  = \new_[615]_  & \new_[610]_ ;
  assign \new_[152]_  = \new_[605]_  & \new_[600]_ ;
  assign \new_[153]_  = \new_[595]_  & \new_[590]_ ;
  assign \new_[154]_  = \new_[585]_  & \new_[580]_ ;
  assign \new_[155]_  = \new_[575]_  & \new_[570]_ ;
  assign \new_[156]_  = \new_[565]_  & \new_[560]_ ;
  assign \new_[157]_  = \new_[555]_  & \new_[550]_ ;
  assign \new_[158]_  = \new_[545]_  & \new_[540]_ ;
  assign \new_[159]_  = \new_[535]_  & \new_[530]_ ;
  assign \new_[160]_  = \new_[525]_  & \new_[522]_ ;
  assign \new_[161]_  = \new_[519]_  & \new_[516]_ ;
  assign \new_[162]_  = \new_[513]_  & \new_[510]_ ;
  assign \new_[163]_  = \new_[507]_  & \new_[504]_ ;
  assign \new_[164]_  = \new_[501]_  & \new_[498]_ ;
  assign \new_[165]_  = A266 & ~A265;
  assign \new_[168]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[172]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[173]_  = \new_[163]_  | \new_[172]_ ;
  assign \new_[174]_  = \new_[173]_  | \new_[168]_ ;
  assign \new_[177]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[181]_  = \new_[156]_  | \new_[157]_ ;
  assign \new_[182]_  = \new_[158]_  | \new_[181]_ ;
  assign \new_[183]_  = \new_[182]_  | \new_[177]_ ;
  assign \new_[184]_  = \new_[183]_  | \new_[174]_ ;
  assign \new_[187]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[191]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[192]_  = \new_[153]_  | \new_[191]_ ;
  assign \new_[193]_  = \new_[192]_  | \new_[187]_ ;
  assign \new_[196]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[200]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[201]_  = \new_[148]_  | \new_[200]_ ;
  assign \new_[202]_  = \new_[201]_  | \new_[196]_ ;
  assign \new_[203]_  = \new_[202]_  | \new_[193]_ ;
  assign \new_[204]_  = \new_[203]_  | \new_[184]_ ;
  assign \new_[207]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[211]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[212]_  = \new_[143]_  | \new_[211]_ ;
  assign \new_[213]_  = \new_[212]_  | \new_[207]_ ;
  assign \new_[216]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[220]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[221]_  = \new_[138]_  | \new_[220]_ ;
  assign \new_[222]_  = \new_[221]_  | \new_[216]_ ;
  assign \new_[223]_  = \new_[222]_  | \new_[213]_ ;
  assign \new_[226]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[230]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[231]_  = \new_[133]_  | \new_[230]_ ;
  assign \new_[232]_  = \new_[231]_  | \new_[226]_ ;
  assign \new_[236]_  = \new_[128]_  | \new_[129]_ ;
  assign \new_[237]_  = \new_[130]_  | \new_[236]_ ;
  assign \new_[241]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[242]_  = \new_[127]_  | \new_[241]_ ;
  assign \new_[243]_  = \new_[242]_  | \new_[237]_ ;
  assign \new_[244]_  = \new_[243]_  | \new_[232]_ ;
  assign \new_[245]_  = \new_[244]_  | \new_[223]_ ;
  assign \new_[246]_  = \new_[245]_  | \new_[204]_ ;
  assign \new_[249]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[253]_  = \new_[120]_  | \new_[121]_ ;
  assign \new_[254]_  = \new_[122]_  | \new_[253]_ ;
  assign \new_[255]_  = \new_[254]_  | \new_[249]_ ;
  assign \new_[258]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[262]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[263]_  = \new_[117]_  | \new_[262]_ ;
  assign \new_[264]_  = \new_[263]_  | \new_[258]_ ;
  assign \new_[265]_  = \new_[264]_  | \new_[255]_ ;
  assign \new_[268]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[272]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[273]_  = \new_[112]_  | \new_[272]_ ;
  assign \new_[274]_  = \new_[273]_  | \new_[268]_ ;
  assign \new_[277]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[281]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[282]_  = \new_[107]_  | \new_[281]_ ;
  assign \new_[283]_  = \new_[282]_  | \new_[277]_ ;
  assign \new_[284]_  = \new_[283]_  | \new_[274]_ ;
  assign \new_[285]_  = \new_[284]_  | \new_[265]_ ;
  assign \new_[288]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[292]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[293]_  = \new_[102]_  | \new_[292]_ ;
  assign \new_[294]_  = \new_[293]_  | \new_[288]_ ;
  assign \new_[297]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[301]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[302]_  = \new_[97]_  | \new_[301]_ ;
  assign \new_[303]_  = \new_[302]_  | \new_[297]_ ;
  assign \new_[304]_  = \new_[303]_  | \new_[294]_ ;
  assign \new_[307]_  = \new_[93]_  | \new_[94]_ ;
  assign \new_[311]_  = \new_[90]_  | \new_[91]_ ;
  assign \new_[312]_  = \new_[92]_  | \new_[311]_ ;
  assign \new_[313]_  = \new_[312]_  | \new_[307]_ ;
  assign \new_[317]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[318]_  = \new_[89]_  | \new_[317]_ ;
  assign \new_[322]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[323]_  = \new_[86]_  | \new_[322]_ ;
  assign \new_[324]_  = \new_[323]_  | \new_[318]_ ;
  assign \new_[325]_  = \new_[324]_  | \new_[313]_ ;
  assign \new_[326]_  = \new_[325]_  | \new_[304]_ ;
  assign \new_[327]_  = \new_[326]_  | \new_[285]_ ;
  assign \new_[328]_  = \new_[327]_  | \new_[246]_ ;
  assign \new_[331]_  = \new_[82]_  | \new_[83]_ ;
  assign \new_[335]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[336]_  = \new_[81]_  | \new_[335]_ ;
  assign \new_[337]_  = \new_[336]_  | \new_[331]_ ;
  assign \new_[340]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[344]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[345]_  = \new_[76]_  | \new_[344]_ ;
  assign \new_[346]_  = \new_[345]_  | \new_[340]_ ;
  assign \new_[347]_  = \new_[346]_  | \new_[337]_ ;
  assign \new_[350]_  = \new_[72]_  | \new_[73]_ ;
  assign \new_[354]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[355]_  = \new_[71]_  | \new_[354]_ ;
  assign \new_[356]_  = \new_[355]_  | \new_[350]_ ;
  assign \new_[359]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[363]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[364]_  = \new_[66]_  | \new_[363]_ ;
  assign \new_[365]_  = \new_[364]_  | \new_[359]_ ;
  assign \new_[366]_  = \new_[365]_  | \new_[356]_ ;
  assign \new_[367]_  = \new_[366]_  | \new_[347]_ ;
  assign \new_[370]_  = \new_[62]_  | \new_[63]_ ;
  assign \new_[374]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[375]_  = \new_[61]_  | \new_[374]_ ;
  assign \new_[376]_  = \new_[375]_  | \new_[370]_ ;
  assign \new_[379]_  = \new_[57]_  | \new_[58]_ ;
  assign \new_[383]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[384]_  = \new_[56]_  | \new_[383]_ ;
  assign \new_[385]_  = \new_[384]_  | \new_[379]_ ;
  assign \new_[386]_  = \new_[385]_  | \new_[376]_ ;
  assign \new_[389]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[393]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[394]_  = \new_[51]_  | \new_[393]_ ;
  assign \new_[395]_  = \new_[394]_  | \new_[389]_ ;
  assign \new_[399]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[400]_  = \new_[48]_  | \new_[399]_ ;
  assign \new_[404]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[405]_  = \new_[45]_  | \new_[404]_ ;
  assign \new_[406]_  = \new_[405]_  | \new_[400]_ ;
  assign \new_[407]_  = \new_[406]_  | \new_[395]_ ;
  assign \new_[408]_  = \new_[407]_  | \new_[386]_ ;
  assign \new_[409]_  = \new_[408]_  | \new_[367]_ ;
  assign \new_[412]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[416]_  = \new_[38]_  | \new_[39]_ ;
  assign \new_[417]_  = \new_[40]_  | \new_[416]_ ;
  assign \new_[418]_  = \new_[417]_  | \new_[412]_ ;
  assign \new_[421]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[425]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[426]_  = \new_[35]_  | \new_[425]_ ;
  assign \new_[427]_  = \new_[426]_  | \new_[421]_ ;
  assign \new_[428]_  = \new_[427]_  | \new_[418]_ ;
  assign \new_[431]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[435]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[436]_  = \new_[30]_  | \new_[435]_ ;
  assign \new_[437]_  = \new_[436]_  | \new_[431]_ ;
  assign \new_[441]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[442]_  = \new_[27]_  | \new_[441]_ ;
  assign \new_[446]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[447]_  = \new_[24]_  | \new_[446]_ ;
  assign \new_[448]_  = \new_[447]_  | \new_[442]_ ;
  assign \new_[449]_  = \new_[448]_  | \new_[437]_ ;
  assign \new_[450]_  = \new_[449]_  | \new_[428]_ ;
  assign \new_[453]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[457]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[458]_  = \new_[19]_  | \new_[457]_ ;
  assign \new_[459]_  = \new_[458]_  | \new_[453]_ ;
  assign \new_[462]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[466]_  = \new_[12]_  | \new_[13]_ ;
  assign \new_[467]_  = \new_[14]_  | \new_[466]_ ;
  assign \new_[468]_  = \new_[467]_  | \new_[462]_ ;
  assign \new_[469]_  = \new_[468]_  | \new_[459]_ ;
  assign \new_[472]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[476]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[477]_  = \new_[9]_  | \new_[476]_ ;
  assign \new_[478]_  = \new_[477]_  | \new_[472]_ ;
  assign \new_[482]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[483]_  = \new_[6]_  | \new_[482]_ ;
  assign \new_[487]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[488]_  = \new_[3]_  | \new_[487]_ ;
  assign \new_[489]_  = \new_[488]_  | \new_[483]_ ;
  assign \new_[490]_  = \new_[489]_  | \new_[478]_ ;
  assign \new_[491]_  = \new_[490]_  | \new_[469]_ ;
  assign \new_[492]_  = \new_[491]_  | \new_[450]_ ;
  assign \new_[493]_  = \new_[492]_  | \new_[409]_ ;
  assign \new_[498]_  = ~A266 & A265;
  assign \new_[501]_  = A268 & A267;
  assign \new_[504]_  = ~A266 & A265;
  assign \new_[507]_  = A269 & A267;
  assign \new_[510]_  = A200 & ~A199;
  assign \new_[513]_  = A233 & ~A232;
  assign \new_[516]_  = A166 & A168;
  assign \new_[519]_  = A233 & ~A232;
  assign \new_[522]_  = A167 & A168;
  assign \new_[525]_  = A233 & ~A232;
  assign \new_[529]_  = A232 & A200;
  assign \new_[530]_  = ~A199 & \new_[529]_ ;
  assign \new_[534]_  = A235 & A234;
  assign \new_[535]_  = ~A233 & \new_[534]_ ;
  assign \new_[539]_  = A232 & A200;
  assign \new_[540]_  = ~A199 & \new_[539]_ ;
  assign \new_[544]_  = A236 & A234;
  assign \new_[545]_  = ~A233 & \new_[544]_ ;
  assign \new_[549]_  = A201 & ~A200;
  assign \new_[550]_  = A199 & \new_[549]_ ;
  assign \new_[554]_  = A233 & ~A232;
  assign \new_[555]_  = A202 & \new_[554]_ ;
  assign \new_[559]_  = A201 & ~A200;
  assign \new_[560]_  = A199 & \new_[559]_ ;
  assign \new_[564]_  = A233 & ~A232;
  assign \new_[565]_  = A203 & \new_[564]_ ;
  assign \new_[569]_  = A232 & A166;
  assign \new_[570]_  = A168 & \new_[569]_ ;
  assign \new_[574]_  = A235 & A234;
  assign \new_[575]_  = ~A233 & \new_[574]_ ;
  assign \new_[579]_  = A232 & A166;
  assign \new_[580]_  = A168 & \new_[579]_ ;
  assign \new_[584]_  = A236 & A234;
  assign \new_[585]_  = ~A233 & \new_[584]_ ;
  assign \new_[589]_  = A199 & A166;
  assign \new_[590]_  = A168 & \new_[589]_ ;
  assign \new_[594]_  = A299 & ~A298;
  assign \new_[595]_  = A200 & \new_[594]_ ;
  assign \new_[599]_  = ~A200 & A166;
  assign \new_[600]_  = A168 & \new_[599]_ ;
  assign \new_[604]_  = A299 & ~A298;
  assign \new_[605]_  = ~A201 & \new_[604]_ ;
  assign \new_[609]_  = ~A199 & A166;
  assign \new_[610]_  = A168 & \new_[609]_ ;
  assign \new_[614]_  = A299 & ~A298;
  assign \new_[615]_  = ~A200 & \new_[614]_ ;
  assign \new_[619]_  = A232 & A167;
  assign \new_[620]_  = A168 & \new_[619]_ ;
  assign \new_[624]_  = A235 & A234;
  assign \new_[625]_  = ~A233 & \new_[624]_ ;
  assign \new_[629]_  = A232 & A167;
  assign \new_[630]_  = A168 & \new_[629]_ ;
  assign \new_[634]_  = A236 & A234;
  assign \new_[635]_  = ~A233 & \new_[634]_ ;
  assign \new_[639]_  = A199 & A167;
  assign \new_[640]_  = A168 & \new_[639]_ ;
  assign \new_[644]_  = A299 & ~A298;
  assign \new_[645]_  = A200 & \new_[644]_ ;
  assign \new_[649]_  = ~A200 & A167;
  assign \new_[650]_  = A168 & \new_[649]_ ;
  assign \new_[654]_  = A299 & ~A298;
  assign \new_[655]_  = ~A201 & \new_[654]_ ;
  assign \new_[659]_  = ~A199 & A167;
  assign \new_[660]_  = A168 & \new_[659]_ ;
  assign \new_[664]_  = A299 & ~A298;
  assign \new_[665]_  = ~A200 & \new_[664]_ ;
  assign \new_[669]_  = A167 & A169;
  assign \new_[670]_  = ~A170 & \new_[669]_ ;
  assign \new_[674]_  = A233 & ~A232;
  assign \new_[675]_  = A166 & \new_[674]_ ;
  assign \new_[679]_  = ~A167 & A169;
  assign \new_[680]_  = ~A170 & \new_[679]_ ;
  assign \new_[684]_  = A233 & ~A232;
  assign \new_[685]_  = ~A166 & \new_[684]_ ;
  assign \new_[689]_  = A167 & ~A169;
  assign \new_[690]_  = A170 & \new_[689]_ ;
  assign \new_[694]_  = A233 & ~A232;
  assign \new_[695]_  = ~A166 & \new_[694]_ ;
  assign \new_[699]_  = ~A167 & ~A169;
  assign \new_[700]_  = A170 & \new_[699]_ ;
  assign \new_[704]_  = A233 & ~A232;
  assign \new_[705]_  = A166 & \new_[704]_ ;
  assign \new_[709]_  = ~A200 & A166;
  assign \new_[710]_  = A168 & \new_[709]_ ;
  assign \new_[713]_  = ~A203 & ~A202;
  assign \new_[716]_  = A299 & ~A298;
  assign \new_[717]_  = \new_[716]_  & \new_[713]_ ;
  assign \new_[721]_  = ~A200 & A167;
  assign \new_[722]_  = A168 & \new_[721]_ ;
  assign \new_[725]_  = ~A203 & ~A202;
  assign \new_[728]_  = A299 & ~A298;
  assign \new_[729]_  = \new_[728]_  & \new_[725]_ ;
  assign \new_[733]_  = ~A166 & ~A167;
  assign \new_[734]_  = A170 & \new_[733]_ ;
  assign \new_[737]_  = A200 & ~A199;
  assign \new_[740]_  = A299 & ~A298;
  assign \new_[741]_  = \new_[740]_  & \new_[737]_ ;
  assign \new_[745]_  = ~A168 & A169;
  assign \new_[746]_  = A170 & \new_[745]_ ;
  assign \new_[749]_  = A200 & ~A199;
  assign \new_[752]_  = A299 & ~A298;
  assign \new_[753]_  = \new_[752]_  & \new_[749]_ ;
  assign \new_[757]_  = ~A166 & ~A167;
  assign \new_[758]_  = ~A169 & \new_[757]_ ;
  assign \new_[761]_  = A200 & ~A199;
  assign \new_[764]_  = A299 & ~A298;
  assign \new_[765]_  = \new_[764]_  & \new_[761]_ ;
  assign \new_[769]_  = ~A168 & ~A169;
  assign \new_[770]_  = ~A170 & \new_[769]_ ;
  assign \new_[773]_  = A200 & ~A199;
  assign \new_[776]_  = A299 & ~A298;
  assign \new_[777]_  = \new_[776]_  & \new_[773]_ ;
  assign \new_[780]_  = ~A200 & A199;
  assign \new_[783]_  = A202 & A201;
  assign \new_[784]_  = \new_[783]_  & \new_[780]_ ;
  assign \new_[787]_  = ~A233 & A232;
  assign \new_[790]_  = A235 & A234;
  assign \new_[791]_  = \new_[790]_  & \new_[787]_ ;
  assign \new_[794]_  = ~A200 & A199;
  assign \new_[797]_  = A202 & A201;
  assign \new_[798]_  = \new_[797]_  & \new_[794]_ ;
  assign \new_[801]_  = ~A233 & A232;
  assign \new_[804]_  = A236 & A234;
  assign \new_[805]_  = \new_[804]_  & \new_[801]_ ;
  assign \new_[808]_  = ~A200 & A199;
  assign \new_[811]_  = A203 & A201;
  assign \new_[812]_  = \new_[811]_  & \new_[808]_ ;
  assign \new_[815]_  = ~A233 & A232;
  assign \new_[818]_  = A235 & A234;
  assign \new_[819]_  = \new_[818]_  & \new_[815]_ ;
  assign \new_[822]_  = ~A200 & A199;
  assign \new_[825]_  = A203 & A201;
  assign \new_[826]_  = \new_[825]_  & \new_[822]_ ;
  assign \new_[829]_  = ~A233 & A232;
  assign \new_[832]_  = A236 & A234;
  assign \new_[833]_  = \new_[832]_  & \new_[829]_ ;
  assign \new_[836]_  = A166 & A168;
  assign \new_[839]_  = A200 & A199;
  assign \new_[840]_  = \new_[839]_  & \new_[836]_ ;
  assign \new_[843]_  = ~A299 & A298;
  assign \new_[846]_  = A301 & A300;
  assign \new_[847]_  = \new_[846]_  & \new_[843]_ ;
  assign \new_[850]_  = A166 & A168;
  assign \new_[853]_  = A200 & A199;
  assign \new_[854]_  = \new_[853]_  & \new_[850]_ ;
  assign \new_[857]_  = ~A299 & A298;
  assign \new_[860]_  = A302 & A300;
  assign \new_[861]_  = \new_[860]_  & \new_[857]_ ;
  assign \new_[864]_  = A166 & A168;
  assign \new_[867]_  = ~A201 & ~A200;
  assign \new_[868]_  = \new_[867]_  & \new_[864]_ ;
  assign \new_[871]_  = ~A299 & A298;
  assign \new_[874]_  = A301 & A300;
  assign \new_[875]_  = \new_[874]_  & \new_[871]_ ;
  assign \new_[878]_  = A166 & A168;
  assign \new_[881]_  = ~A201 & ~A200;
  assign \new_[882]_  = \new_[881]_  & \new_[878]_ ;
  assign \new_[885]_  = ~A299 & A298;
  assign \new_[888]_  = A302 & A300;
  assign \new_[889]_  = \new_[888]_  & \new_[885]_ ;
  assign \new_[892]_  = A166 & A168;
  assign \new_[895]_  = ~A200 & ~A199;
  assign \new_[896]_  = \new_[895]_  & \new_[892]_ ;
  assign \new_[899]_  = ~A299 & A298;
  assign \new_[902]_  = A301 & A300;
  assign \new_[903]_  = \new_[902]_  & \new_[899]_ ;
  assign \new_[906]_  = A166 & A168;
  assign \new_[909]_  = ~A200 & ~A199;
  assign \new_[910]_  = \new_[909]_  & \new_[906]_ ;
  assign \new_[913]_  = ~A299 & A298;
  assign \new_[916]_  = A302 & A300;
  assign \new_[917]_  = \new_[916]_  & \new_[913]_ ;
  assign \new_[920]_  = A167 & A168;
  assign \new_[923]_  = A200 & A199;
  assign \new_[924]_  = \new_[923]_  & \new_[920]_ ;
  assign \new_[927]_  = ~A299 & A298;
  assign \new_[930]_  = A301 & A300;
  assign \new_[931]_  = \new_[930]_  & \new_[927]_ ;
  assign \new_[934]_  = A167 & A168;
  assign \new_[937]_  = A200 & A199;
  assign \new_[938]_  = \new_[937]_  & \new_[934]_ ;
  assign \new_[941]_  = ~A299 & A298;
  assign \new_[944]_  = A302 & A300;
  assign \new_[945]_  = \new_[944]_  & \new_[941]_ ;
  assign \new_[948]_  = A167 & A168;
  assign \new_[951]_  = ~A201 & ~A200;
  assign \new_[952]_  = \new_[951]_  & \new_[948]_ ;
  assign \new_[955]_  = ~A299 & A298;
  assign \new_[958]_  = A301 & A300;
  assign \new_[959]_  = \new_[958]_  & \new_[955]_ ;
  assign \new_[962]_  = A167 & A168;
  assign \new_[965]_  = ~A201 & ~A200;
  assign \new_[966]_  = \new_[965]_  & \new_[962]_ ;
  assign \new_[969]_  = ~A299 & A298;
  assign \new_[972]_  = A302 & A300;
  assign \new_[973]_  = \new_[972]_  & \new_[969]_ ;
  assign \new_[976]_  = A167 & A168;
  assign \new_[979]_  = ~A200 & ~A199;
  assign \new_[980]_  = \new_[979]_  & \new_[976]_ ;
  assign \new_[983]_  = ~A299 & A298;
  assign \new_[986]_  = A301 & A300;
  assign \new_[987]_  = \new_[986]_  & \new_[983]_ ;
  assign \new_[990]_  = A167 & A168;
  assign \new_[993]_  = ~A200 & ~A199;
  assign \new_[994]_  = \new_[993]_  & \new_[990]_ ;
  assign \new_[997]_  = ~A299 & A298;
  assign \new_[1000]_  = A302 & A300;
  assign \new_[1001]_  = \new_[1000]_  & \new_[997]_ ;
  assign \new_[1004]_  = ~A168 & A169;
  assign \new_[1007]_  = ~A166 & A167;
  assign \new_[1008]_  = \new_[1007]_  & \new_[1004]_ ;
  assign \new_[1011]_  = A200 & ~A199;
  assign \new_[1014]_  = A299 & ~A298;
  assign \new_[1015]_  = \new_[1014]_  & \new_[1011]_ ;
  assign \new_[1018]_  = ~A168 & A169;
  assign \new_[1021]_  = A166 & ~A167;
  assign \new_[1022]_  = \new_[1021]_  & \new_[1018]_ ;
  assign \new_[1025]_  = A200 & ~A199;
  assign \new_[1028]_  = A299 & ~A298;
  assign \new_[1029]_  = \new_[1028]_  & \new_[1025]_ ;
  assign \new_[1032]_  = A169 & ~A170;
  assign \new_[1035]_  = A166 & A167;
  assign \new_[1036]_  = \new_[1035]_  & \new_[1032]_ ;
  assign \new_[1039]_  = ~A233 & A232;
  assign \new_[1042]_  = A235 & A234;
  assign \new_[1043]_  = \new_[1042]_  & \new_[1039]_ ;
  assign \new_[1046]_  = A169 & ~A170;
  assign \new_[1049]_  = A166 & A167;
  assign \new_[1050]_  = \new_[1049]_  & \new_[1046]_ ;
  assign \new_[1053]_  = ~A233 & A232;
  assign \new_[1056]_  = A236 & A234;
  assign \new_[1057]_  = \new_[1056]_  & \new_[1053]_ ;
  assign \new_[1060]_  = A169 & ~A170;
  assign \new_[1063]_  = A166 & A167;
  assign \new_[1064]_  = \new_[1063]_  & \new_[1060]_ ;
  assign \new_[1067]_  = A200 & A199;
  assign \new_[1070]_  = A299 & ~A298;
  assign \new_[1071]_  = \new_[1070]_  & \new_[1067]_ ;
  assign \new_[1074]_  = A169 & ~A170;
  assign \new_[1077]_  = A166 & A167;
  assign \new_[1078]_  = \new_[1077]_  & \new_[1074]_ ;
  assign \new_[1081]_  = ~A201 & ~A200;
  assign \new_[1084]_  = A299 & ~A298;
  assign \new_[1085]_  = \new_[1084]_  & \new_[1081]_ ;
  assign \new_[1088]_  = A169 & ~A170;
  assign \new_[1091]_  = A166 & A167;
  assign \new_[1092]_  = \new_[1091]_  & \new_[1088]_ ;
  assign \new_[1095]_  = ~A200 & ~A199;
  assign \new_[1098]_  = A299 & ~A298;
  assign \new_[1099]_  = \new_[1098]_  & \new_[1095]_ ;
  assign \new_[1102]_  = A169 & ~A170;
  assign \new_[1105]_  = ~A166 & ~A167;
  assign \new_[1106]_  = \new_[1105]_  & \new_[1102]_ ;
  assign \new_[1109]_  = ~A233 & A232;
  assign \new_[1112]_  = A235 & A234;
  assign \new_[1113]_  = \new_[1112]_  & \new_[1109]_ ;
  assign \new_[1116]_  = A169 & ~A170;
  assign \new_[1119]_  = ~A166 & ~A167;
  assign \new_[1120]_  = \new_[1119]_  & \new_[1116]_ ;
  assign \new_[1123]_  = ~A233 & A232;
  assign \new_[1126]_  = A236 & A234;
  assign \new_[1127]_  = \new_[1126]_  & \new_[1123]_ ;
  assign \new_[1130]_  = A169 & ~A170;
  assign \new_[1133]_  = ~A166 & ~A167;
  assign \new_[1134]_  = \new_[1133]_  & \new_[1130]_ ;
  assign \new_[1137]_  = A200 & A199;
  assign \new_[1140]_  = A299 & ~A298;
  assign \new_[1141]_  = \new_[1140]_  & \new_[1137]_ ;
  assign \new_[1144]_  = A169 & ~A170;
  assign \new_[1147]_  = ~A166 & ~A167;
  assign \new_[1148]_  = \new_[1147]_  & \new_[1144]_ ;
  assign \new_[1151]_  = ~A201 & ~A200;
  assign \new_[1154]_  = A299 & ~A298;
  assign \new_[1155]_  = \new_[1154]_  & \new_[1151]_ ;
  assign \new_[1158]_  = A169 & ~A170;
  assign \new_[1161]_  = ~A166 & ~A167;
  assign \new_[1162]_  = \new_[1161]_  & \new_[1158]_ ;
  assign \new_[1165]_  = ~A200 & ~A199;
  assign \new_[1168]_  = A299 & ~A298;
  assign \new_[1169]_  = \new_[1168]_  & \new_[1165]_ ;
  assign \new_[1172]_  = ~A168 & ~A169;
  assign \new_[1175]_  = A166 & A167;
  assign \new_[1176]_  = \new_[1175]_  & \new_[1172]_ ;
  assign \new_[1179]_  = A200 & ~A199;
  assign \new_[1182]_  = A299 & ~A298;
  assign \new_[1183]_  = \new_[1182]_  & \new_[1179]_ ;
  assign \new_[1186]_  = ~A169 & A170;
  assign \new_[1189]_  = ~A166 & A167;
  assign \new_[1190]_  = \new_[1189]_  & \new_[1186]_ ;
  assign \new_[1193]_  = ~A233 & A232;
  assign \new_[1196]_  = A235 & A234;
  assign \new_[1197]_  = \new_[1196]_  & \new_[1193]_ ;
  assign \new_[1200]_  = ~A169 & A170;
  assign \new_[1203]_  = ~A166 & A167;
  assign \new_[1204]_  = \new_[1203]_  & \new_[1200]_ ;
  assign \new_[1207]_  = ~A233 & A232;
  assign \new_[1210]_  = A236 & A234;
  assign \new_[1211]_  = \new_[1210]_  & \new_[1207]_ ;
  assign \new_[1214]_  = ~A169 & A170;
  assign \new_[1217]_  = ~A166 & A167;
  assign \new_[1218]_  = \new_[1217]_  & \new_[1214]_ ;
  assign \new_[1221]_  = A200 & A199;
  assign \new_[1224]_  = A299 & ~A298;
  assign \new_[1225]_  = \new_[1224]_  & \new_[1221]_ ;
  assign \new_[1228]_  = ~A169 & A170;
  assign \new_[1231]_  = ~A166 & A167;
  assign \new_[1232]_  = \new_[1231]_  & \new_[1228]_ ;
  assign \new_[1235]_  = ~A201 & ~A200;
  assign \new_[1238]_  = A299 & ~A298;
  assign \new_[1239]_  = \new_[1238]_  & \new_[1235]_ ;
  assign \new_[1242]_  = ~A169 & A170;
  assign \new_[1245]_  = ~A166 & A167;
  assign \new_[1246]_  = \new_[1245]_  & \new_[1242]_ ;
  assign \new_[1249]_  = ~A200 & ~A199;
  assign \new_[1252]_  = A299 & ~A298;
  assign \new_[1253]_  = \new_[1252]_  & \new_[1249]_ ;
  assign \new_[1256]_  = ~A169 & A170;
  assign \new_[1259]_  = A166 & ~A167;
  assign \new_[1260]_  = \new_[1259]_  & \new_[1256]_ ;
  assign \new_[1263]_  = ~A233 & A232;
  assign \new_[1266]_  = A235 & A234;
  assign \new_[1267]_  = \new_[1266]_  & \new_[1263]_ ;
  assign \new_[1270]_  = ~A169 & A170;
  assign \new_[1273]_  = A166 & ~A167;
  assign \new_[1274]_  = \new_[1273]_  & \new_[1270]_ ;
  assign \new_[1277]_  = ~A233 & A232;
  assign \new_[1280]_  = A236 & A234;
  assign \new_[1281]_  = \new_[1280]_  & \new_[1277]_ ;
  assign \new_[1284]_  = ~A169 & A170;
  assign \new_[1287]_  = A166 & ~A167;
  assign \new_[1288]_  = \new_[1287]_  & \new_[1284]_ ;
  assign \new_[1291]_  = A200 & A199;
  assign \new_[1294]_  = A299 & ~A298;
  assign \new_[1295]_  = \new_[1294]_  & \new_[1291]_ ;
  assign \new_[1298]_  = ~A169 & A170;
  assign \new_[1301]_  = A166 & ~A167;
  assign \new_[1302]_  = \new_[1301]_  & \new_[1298]_ ;
  assign \new_[1305]_  = ~A201 & ~A200;
  assign \new_[1308]_  = A299 & ~A298;
  assign \new_[1309]_  = \new_[1308]_  & \new_[1305]_ ;
  assign \new_[1312]_  = ~A169 & A170;
  assign \new_[1315]_  = A166 & ~A167;
  assign \new_[1316]_  = \new_[1315]_  & \new_[1312]_ ;
  assign \new_[1319]_  = ~A200 & ~A199;
  assign \new_[1322]_  = A299 & ~A298;
  assign \new_[1323]_  = \new_[1322]_  & \new_[1319]_ ;
  assign \new_[1326]_  = A166 & A168;
  assign \new_[1329]_  = ~A202 & ~A200;
  assign \new_[1330]_  = \new_[1329]_  & \new_[1326]_ ;
  assign \new_[1333]_  = A298 & ~A203;
  assign \new_[1337]_  = A301 & A300;
  assign \new_[1338]_  = ~A299 & \new_[1337]_ ;
  assign \new_[1339]_  = \new_[1338]_  & \new_[1333]_ ;
  assign \new_[1342]_  = A166 & A168;
  assign \new_[1345]_  = ~A202 & ~A200;
  assign \new_[1346]_  = \new_[1345]_  & \new_[1342]_ ;
  assign \new_[1349]_  = A298 & ~A203;
  assign \new_[1353]_  = A302 & A300;
  assign \new_[1354]_  = ~A299 & \new_[1353]_ ;
  assign \new_[1355]_  = \new_[1354]_  & \new_[1349]_ ;
  assign \new_[1358]_  = A167 & A168;
  assign \new_[1361]_  = ~A202 & ~A200;
  assign \new_[1362]_  = \new_[1361]_  & \new_[1358]_ ;
  assign \new_[1365]_  = A298 & ~A203;
  assign \new_[1369]_  = A301 & A300;
  assign \new_[1370]_  = ~A299 & \new_[1369]_ ;
  assign \new_[1371]_  = \new_[1370]_  & \new_[1365]_ ;
  assign \new_[1374]_  = A167 & A168;
  assign \new_[1377]_  = ~A202 & ~A200;
  assign \new_[1378]_  = \new_[1377]_  & \new_[1374]_ ;
  assign \new_[1381]_  = A298 & ~A203;
  assign \new_[1385]_  = A302 & A300;
  assign \new_[1386]_  = ~A299 & \new_[1385]_ ;
  assign \new_[1387]_  = \new_[1386]_  & \new_[1381]_ ;
  assign \new_[1390]_  = ~A167 & A170;
  assign \new_[1393]_  = ~A199 & ~A166;
  assign \new_[1394]_  = \new_[1393]_  & \new_[1390]_ ;
  assign \new_[1397]_  = A298 & A200;
  assign \new_[1401]_  = A301 & A300;
  assign \new_[1402]_  = ~A299 & \new_[1401]_ ;
  assign \new_[1403]_  = \new_[1402]_  & \new_[1397]_ ;
  assign \new_[1406]_  = ~A167 & A170;
  assign \new_[1409]_  = ~A199 & ~A166;
  assign \new_[1410]_  = \new_[1409]_  & \new_[1406]_ ;
  assign \new_[1413]_  = A298 & A200;
  assign \new_[1417]_  = A302 & A300;
  assign \new_[1418]_  = ~A299 & \new_[1417]_ ;
  assign \new_[1419]_  = \new_[1418]_  & \new_[1413]_ ;
  assign \new_[1422]_  = ~A167 & A170;
  assign \new_[1425]_  = A199 & ~A166;
  assign \new_[1426]_  = \new_[1425]_  & \new_[1422]_ ;
  assign \new_[1429]_  = A201 & ~A200;
  assign \new_[1433]_  = A299 & ~A298;
  assign \new_[1434]_  = A202 & \new_[1433]_ ;
  assign \new_[1435]_  = \new_[1434]_  & \new_[1429]_ ;
  assign \new_[1438]_  = ~A167 & A170;
  assign \new_[1441]_  = A199 & ~A166;
  assign \new_[1442]_  = \new_[1441]_  & \new_[1438]_ ;
  assign \new_[1445]_  = A201 & ~A200;
  assign \new_[1449]_  = A299 & ~A298;
  assign \new_[1450]_  = A203 & \new_[1449]_ ;
  assign \new_[1451]_  = \new_[1450]_  & \new_[1445]_ ;
  assign \new_[1454]_  = A169 & A170;
  assign \new_[1457]_  = ~A199 & ~A168;
  assign \new_[1458]_  = \new_[1457]_  & \new_[1454]_ ;
  assign \new_[1461]_  = A298 & A200;
  assign \new_[1465]_  = A301 & A300;
  assign \new_[1466]_  = ~A299 & \new_[1465]_ ;
  assign \new_[1467]_  = \new_[1466]_  & \new_[1461]_ ;
  assign \new_[1470]_  = A169 & A170;
  assign \new_[1473]_  = ~A199 & ~A168;
  assign \new_[1474]_  = \new_[1473]_  & \new_[1470]_ ;
  assign \new_[1477]_  = A298 & A200;
  assign \new_[1481]_  = A302 & A300;
  assign \new_[1482]_  = ~A299 & \new_[1481]_ ;
  assign \new_[1483]_  = \new_[1482]_  & \new_[1477]_ ;
  assign \new_[1486]_  = A169 & A170;
  assign \new_[1489]_  = A199 & ~A168;
  assign \new_[1490]_  = \new_[1489]_  & \new_[1486]_ ;
  assign \new_[1493]_  = A201 & ~A200;
  assign \new_[1497]_  = A299 & ~A298;
  assign \new_[1498]_  = A202 & \new_[1497]_ ;
  assign \new_[1499]_  = \new_[1498]_  & \new_[1493]_ ;
  assign \new_[1502]_  = A169 & A170;
  assign \new_[1505]_  = A199 & ~A168;
  assign \new_[1506]_  = \new_[1505]_  & \new_[1502]_ ;
  assign \new_[1509]_  = A201 & ~A200;
  assign \new_[1513]_  = A299 & ~A298;
  assign \new_[1514]_  = A203 & \new_[1513]_ ;
  assign \new_[1515]_  = \new_[1514]_  & \new_[1509]_ ;
  assign \new_[1518]_  = A169 & ~A170;
  assign \new_[1521]_  = A166 & A167;
  assign \new_[1522]_  = \new_[1521]_  & \new_[1518]_ ;
  assign \new_[1525]_  = ~A202 & ~A200;
  assign \new_[1529]_  = A299 & ~A298;
  assign \new_[1530]_  = ~A203 & \new_[1529]_ ;
  assign \new_[1531]_  = \new_[1530]_  & \new_[1525]_ ;
  assign \new_[1534]_  = A169 & ~A170;
  assign \new_[1537]_  = ~A166 & ~A167;
  assign \new_[1538]_  = \new_[1537]_  & \new_[1534]_ ;
  assign \new_[1541]_  = ~A202 & ~A200;
  assign \new_[1545]_  = A299 & ~A298;
  assign \new_[1546]_  = ~A203 & \new_[1545]_ ;
  assign \new_[1547]_  = \new_[1546]_  & \new_[1541]_ ;
  assign \new_[1550]_  = ~A167 & ~A169;
  assign \new_[1553]_  = ~A199 & ~A166;
  assign \new_[1554]_  = \new_[1553]_  & \new_[1550]_ ;
  assign \new_[1557]_  = A298 & A200;
  assign \new_[1561]_  = A301 & A300;
  assign \new_[1562]_  = ~A299 & \new_[1561]_ ;
  assign \new_[1563]_  = \new_[1562]_  & \new_[1557]_ ;
  assign \new_[1566]_  = ~A167 & ~A169;
  assign \new_[1569]_  = ~A199 & ~A166;
  assign \new_[1570]_  = \new_[1569]_  & \new_[1566]_ ;
  assign \new_[1573]_  = A298 & A200;
  assign \new_[1577]_  = A302 & A300;
  assign \new_[1578]_  = ~A299 & \new_[1577]_ ;
  assign \new_[1579]_  = \new_[1578]_  & \new_[1573]_ ;
  assign \new_[1582]_  = ~A167 & ~A169;
  assign \new_[1585]_  = A199 & ~A166;
  assign \new_[1586]_  = \new_[1585]_  & \new_[1582]_ ;
  assign \new_[1589]_  = A201 & ~A200;
  assign \new_[1593]_  = A299 & ~A298;
  assign \new_[1594]_  = A202 & \new_[1593]_ ;
  assign \new_[1595]_  = \new_[1594]_  & \new_[1589]_ ;
  assign \new_[1598]_  = ~A167 & ~A169;
  assign \new_[1601]_  = A199 & ~A166;
  assign \new_[1602]_  = \new_[1601]_  & \new_[1598]_ ;
  assign \new_[1605]_  = A201 & ~A200;
  assign \new_[1609]_  = A299 & ~A298;
  assign \new_[1610]_  = A203 & \new_[1609]_ ;
  assign \new_[1611]_  = \new_[1610]_  & \new_[1605]_ ;
  assign \new_[1614]_  = ~A169 & A170;
  assign \new_[1617]_  = ~A166 & A167;
  assign \new_[1618]_  = \new_[1617]_  & \new_[1614]_ ;
  assign \new_[1621]_  = ~A202 & ~A200;
  assign \new_[1625]_  = A299 & ~A298;
  assign \new_[1626]_  = ~A203 & \new_[1625]_ ;
  assign \new_[1627]_  = \new_[1626]_  & \new_[1621]_ ;
  assign \new_[1630]_  = ~A169 & A170;
  assign \new_[1633]_  = A166 & ~A167;
  assign \new_[1634]_  = \new_[1633]_  & \new_[1630]_ ;
  assign \new_[1637]_  = ~A202 & ~A200;
  assign \new_[1641]_  = A299 & ~A298;
  assign \new_[1642]_  = ~A203 & \new_[1641]_ ;
  assign \new_[1643]_  = \new_[1642]_  & \new_[1637]_ ;
  assign \new_[1646]_  = ~A169 & ~A170;
  assign \new_[1649]_  = ~A199 & ~A168;
  assign \new_[1650]_  = \new_[1649]_  & \new_[1646]_ ;
  assign \new_[1653]_  = A298 & A200;
  assign \new_[1657]_  = A301 & A300;
  assign \new_[1658]_  = ~A299 & \new_[1657]_ ;
  assign \new_[1659]_  = \new_[1658]_  & \new_[1653]_ ;
  assign \new_[1662]_  = ~A169 & ~A170;
  assign \new_[1665]_  = ~A199 & ~A168;
  assign \new_[1666]_  = \new_[1665]_  & \new_[1662]_ ;
  assign \new_[1669]_  = A298 & A200;
  assign \new_[1673]_  = A302 & A300;
  assign \new_[1674]_  = ~A299 & \new_[1673]_ ;
  assign \new_[1675]_  = \new_[1674]_  & \new_[1669]_ ;
  assign \new_[1678]_  = ~A169 & ~A170;
  assign \new_[1681]_  = A199 & ~A168;
  assign \new_[1682]_  = \new_[1681]_  & \new_[1678]_ ;
  assign \new_[1685]_  = A201 & ~A200;
  assign \new_[1689]_  = A299 & ~A298;
  assign \new_[1690]_  = A202 & \new_[1689]_ ;
  assign \new_[1691]_  = \new_[1690]_  & \new_[1685]_ ;
  assign \new_[1694]_  = ~A169 & ~A170;
  assign \new_[1697]_  = A199 & ~A168;
  assign \new_[1698]_  = \new_[1697]_  & \new_[1694]_ ;
  assign \new_[1701]_  = A201 & ~A200;
  assign \new_[1705]_  = A299 & ~A298;
  assign \new_[1706]_  = A203 & \new_[1705]_ ;
  assign \new_[1707]_  = \new_[1706]_  & \new_[1701]_ ;
  assign \new_[1710]_  = ~A168 & A169;
  assign \new_[1714]_  = ~A199 & ~A166;
  assign \new_[1715]_  = A167 & \new_[1714]_ ;
  assign \new_[1716]_  = \new_[1715]_  & \new_[1710]_ ;
  assign \new_[1719]_  = A298 & A200;
  assign \new_[1723]_  = A301 & A300;
  assign \new_[1724]_  = ~A299 & \new_[1723]_ ;
  assign \new_[1725]_  = \new_[1724]_  & \new_[1719]_ ;
  assign \new_[1728]_  = ~A168 & A169;
  assign \new_[1732]_  = ~A199 & ~A166;
  assign \new_[1733]_  = A167 & \new_[1732]_ ;
  assign \new_[1734]_  = \new_[1733]_  & \new_[1728]_ ;
  assign \new_[1737]_  = A298 & A200;
  assign \new_[1741]_  = A302 & A300;
  assign \new_[1742]_  = ~A299 & \new_[1741]_ ;
  assign \new_[1743]_  = \new_[1742]_  & \new_[1737]_ ;
  assign \new_[1746]_  = ~A168 & A169;
  assign \new_[1750]_  = A199 & ~A166;
  assign \new_[1751]_  = A167 & \new_[1750]_ ;
  assign \new_[1752]_  = \new_[1751]_  & \new_[1746]_ ;
  assign \new_[1755]_  = A201 & ~A200;
  assign \new_[1759]_  = A299 & ~A298;
  assign \new_[1760]_  = A202 & \new_[1759]_ ;
  assign \new_[1761]_  = \new_[1760]_  & \new_[1755]_ ;
  assign \new_[1764]_  = ~A168 & A169;
  assign \new_[1768]_  = A199 & ~A166;
  assign \new_[1769]_  = A167 & \new_[1768]_ ;
  assign \new_[1770]_  = \new_[1769]_  & \new_[1764]_ ;
  assign \new_[1773]_  = A201 & ~A200;
  assign \new_[1777]_  = A299 & ~A298;
  assign \new_[1778]_  = A203 & \new_[1777]_ ;
  assign \new_[1779]_  = \new_[1778]_  & \new_[1773]_ ;
  assign \new_[1782]_  = ~A168 & A169;
  assign \new_[1786]_  = ~A199 & A166;
  assign \new_[1787]_  = ~A167 & \new_[1786]_ ;
  assign \new_[1788]_  = \new_[1787]_  & \new_[1782]_ ;
  assign \new_[1791]_  = A298 & A200;
  assign \new_[1795]_  = A301 & A300;
  assign \new_[1796]_  = ~A299 & \new_[1795]_ ;
  assign \new_[1797]_  = \new_[1796]_  & \new_[1791]_ ;
  assign \new_[1800]_  = ~A168 & A169;
  assign \new_[1804]_  = ~A199 & A166;
  assign \new_[1805]_  = ~A167 & \new_[1804]_ ;
  assign \new_[1806]_  = \new_[1805]_  & \new_[1800]_ ;
  assign \new_[1809]_  = A298 & A200;
  assign \new_[1813]_  = A302 & A300;
  assign \new_[1814]_  = ~A299 & \new_[1813]_ ;
  assign \new_[1815]_  = \new_[1814]_  & \new_[1809]_ ;
  assign \new_[1818]_  = ~A168 & A169;
  assign \new_[1822]_  = A199 & A166;
  assign \new_[1823]_  = ~A167 & \new_[1822]_ ;
  assign \new_[1824]_  = \new_[1823]_  & \new_[1818]_ ;
  assign \new_[1827]_  = A201 & ~A200;
  assign \new_[1831]_  = A299 & ~A298;
  assign \new_[1832]_  = A202 & \new_[1831]_ ;
  assign \new_[1833]_  = \new_[1832]_  & \new_[1827]_ ;
  assign \new_[1836]_  = ~A168 & A169;
  assign \new_[1840]_  = A199 & A166;
  assign \new_[1841]_  = ~A167 & \new_[1840]_ ;
  assign \new_[1842]_  = \new_[1841]_  & \new_[1836]_ ;
  assign \new_[1845]_  = A201 & ~A200;
  assign \new_[1849]_  = A299 & ~A298;
  assign \new_[1850]_  = A203 & \new_[1849]_ ;
  assign \new_[1851]_  = \new_[1850]_  & \new_[1845]_ ;
  assign \new_[1854]_  = A169 & ~A170;
  assign \new_[1858]_  = A199 & A166;
  assign \new_[1859]_  = A167 & \new_[1858]_ ;
  assign \new_[1860]_  = \new_[1859]_  & \new_[1854]_ ;
  assign \new_[1863]_  = A298 & A200;
  assign \new_[1867]_  = A301 & A300;
  assign \new_[1868]_  = ~A299 & \new_[1867]_ ;
  assign \new_[1869]_  = \new_[1868]_  & \new_[1863]_ ;
  assign \new_[1872]_  = A169 & ~A170;
  assign \new_[1876]_  = A199 & A166;
  assign \new_[1877]_  = A167 & \new_[1876]_ ;
  assign \new_[1878]_  = \new_[1877]_  & \new_[1872]_ ;
  assign \new_[1881]_  = A298 & A200;
  assign \new_[1885]_  = A302 & A300;
  assign \new_[1886]_  = ~A299 & \new_[1885]_ ;
  assign \new_[1887]_  = \new_[1886]_  & \new_[1881]_ ;
  assign \new_[1890]_  = A169 & ~A170;
  assign \new_[1894]_  = ~A200 & A166;
  assign \new_[1895]_  = A167 & \new_[1894]_ ;
  assign \new_[1896]_  = \new_[1895]_  & \new_[1890]_ ;
  assign \new_[1899]_  = A298 & ~A201;
  assign \new_[1903]_  = A301 & A300;
  assign \new_[1904]_  = ~A299 & \new_[1903]_ ;
  assign \new_[1905]_  = \new_[1904]_  & \new_[1899]_ ;
  assign \new_[1908]_  = A169 & ~A170;
  assign \new_[1912]_  = ~A200 & A166;
  assign \new_[1913]_  = A167 & \new_[1912]_ ;
  assign \new_[1914]_  = \new_[1913]_  & \new_[1908]_ ;
  assign \new_[1917]_  = A298 & ~A201;
  assign \new_[1921]_  = A302 & A300;
  assign \new_[1922]_  = ~A299 & \new_[1921]_ ;
  assign \new_[1923]_  = \new_[1922]_  & \new_[1917]_ ;
  assign \new_[1926]_  = A169 & ~A170;
  assign \new_[1930]_  = ~A199 & A166;
  assign \new_[1931]_  = A167 & \new_[1930]_ ;
  assign \new_[1932]_  = \new_[1931]_  & \new_[1926]_ ;
  assign \new_[1935]_  = A298 & ~A200;
  assign \new_[1939]_  = A301 & A300;
  assign \new_[1940]_  = ~A299 & \new_[1939]_ ;
  assign \new_[1941]_  = \new_[1940]_  & \new_[1935]_ ;
  assign \new_[1944]_  = A169 & ~A170;
  assign \new_[1948]_  = ~A199 & A166;
  assign \new_[1949]_  = A167 & \new_[1948]_ ;
  assign \new_[1950]_  = \new_[1949]_  & \new_[1944]_ ;
  assign \new_[1953]_  = A298 & ~A200;
  assign \new_[1957]_  = A302 & A300;
  assign \new_[1958]_  = ~A299 & \new_[1957]_ ;
  assign \new_[1959]_  = \new_[1958]_  & \new_[1953]_ ;
  assign \new_[1962]_  = A169 & ~A170;
  assign \new_[1966]_  = A199 & ~A166;
  assign \new_[1967]_  = ~A167 & \new_[1966]_ ;
  assign \new_[1968]_  = \new_[1967]_  & \new_[1962]_ ;
  assign \new_[1971]_  = A298 & A200;
  assign \new_[1975]_  = A301 & A300;
  assign \new_[1976]_  = ~A299 & \new_[1975]_ ;
  assign \new_[1977]_  = \new_[1976]_  & \new_[1971]_ ;
  assign \new_[1980]_  = A169 & ~A170;
  assign \new_[1984]_  = A199 & ~A166;
  assign \new_[1985]_  = ~A167 & \new_[1984]_ ;
  assign \new_[1986]_  = \new_[1985]_  & \new_[1980]_ ;
  assign \new_[1989]_  = A298 & A200;
  assign \new_[1993]_  = A302 & A300;
  assign \new_[1994]_  = ~A299 & \new_[1993]_ ;
  assign \new_[1995]_  = \new_[1994]_  & \new_[1989]_ ;
  assign \new_[1998]_  = A169 & ~A170;
  assign \new_[2002]_  = ~A200 & ~A166;
  assign \new_[2003]_  = ~A167 & \new_[2002]_ ;
  assign \new_[2004]_  = \new_[2003]_  & \new_[1998]_ ;
  assign \new_[2007]_  = A298 & ~A201;
  assign \new_[2011]_  = A301 & A300;
  assign \new_[2012]_  = ~A299 & \new_[2011]_ ;
  assign \new_[2013]_  = \new_[2012]_  & \new_[2007]_ ;
  assign \new_[2016]_  = A169 & ~A170;
  assign \new_[2020]_  = ~A200 & ~A166;
  assign \new_[2021]_  = ~A167 & \new_[2020]_ ;
  assign \new_[2022]_  = \new_[2021]_  & \new_[2016]_ ;
  assign \new_[2025]_  = A298 & ~A201;
  assign \new_[2029]_  = A302 & A300;
  assign \new_[2030]_  = ~A299 & \new_[2029]_ ;
  assign \new_[2031]_  = \new_[2030]_  & \new_[2025]_ ;
  assign \new_[2034]_  = A169 & ~A170;
  assign \new_[2038]_  = ~A199 & ~A166;
  assign \new_[2039]_  = ~A167 & \new_[2038]_ ;
  assign \new_[2040]_  = \new_[2039]_  & \new_[2034]_ ;
  assign \new_[2043]_  = A298 & ~A200;
  assign \new_[2047]_  = A301 & A300;
  assign \new_[2048]_  = ~A299 & \new_[2047]_ ;
  assign \new_[2049]_  = \new_[2048]_  & \new_[2043]_ ;
  assign \new_[2052]_  = A169 & ~A170;
  assign \new_[2056]_  = ~A199 & ~A166;
  assign \new_[2057]_  = ~A167 & \new_[2056]_ ;
  assign \new_[2058]_  = \new_[2057]_  & \new_[2052]_ ;
  assign \new_[2061]_  = A298 & ~A200;
  assign \new_[2065]_  = A302 & A300;
  assign \new_[2066]_  = ~A299 & \new_[2065]_ ;
  assign \new_[2067]_  = \new_[2066]_  & \new_[2061]_ ;
  assign \new_[2070]_  = ~A168 & ~A169;
  assign \new_[2074]_  = ~A199 & A166;
  assign \new_[2075]_  = A167 & \new_[2074]_ ;
  assign \new_[2076]_  = \new_[2075]_  & \new_[2070]_ ;
  assign \new_[2079]_  = A298 & A200;
  assign \new_[2083]_  = A301 & A300;
  assign \new_[2084]_  = ~A299 & \new_[2083]_ ;
  assign \new_[2085]_  = \new_[2084]_  & \new_[2079]_ ;
  assign \new_[2088]_  = ~A168 & ~A169;
  assign \new_[2092]_  = ~A199 & A166;
  assign \new_[2093]_  = A167 & \new_[2092]_ ;
  assign \new_[2094]_  = \new_[2093]_  & \new_[2088]_ ;
  assign \new_[2097]_  = A298 & A200;
  assign \new_[2101]_  = A302 & A300;
  assign \new_[2102]_  = ~A299 & \new_[2101]_ ;
  assign \new_[2103]_  = \new_[2102]_  & \new_[2097]_ ;
  assign \new_[2106]_  = ~A168 & ~A169;
  assign \new_[2110]_  = A199 & A166;
  assign \new_[2111]_  = A167 & \new_[2110]_ ;
  assign \new_[2112]_  = \new_[2111]_  & \new_[2106]_ ;
  assign \new_[2115]_  = A201 & ~A200;
  assign \new_[2119]_  = A299 & ~A298;
  assign \new_[2120]_  = A202 & \new_[2119]_ ;
  assign \new_[2121]_  = \new_[2120]_  & \new_[2115]_ ;
  assign \new_[2124]_  = ~A168 & ~A169;
  assign \new_[2128]_  = A199 & A166;
  assign \new_[2129]_  = A167 & \new_[2128]_ ;
  assign \new_[2130]_  = \new_[2129]_  & \new_[2124]_ ;
  assign \new_[2133]_  = A201 & ~A200;
  assign \new_[2137]_  = A299 & ~A298;
  assign \new_[2138]_  = A203 & \new_[2137]_ ;
  assign \new_[2139]_  = \new_[2138]_  & \new_[2133]_ ;
  assign \new_[2142]_  = ~A169 & A170;
  assign \new_[2146]_  = A199 & ~A166;
  assign \new_[2147]_  = A167 & \new_[2146]_ ;
  assign \new_[2148]_  = \new_[2147]_  & \new_[2142]_ ;
  assign \new_[2151]_  = A298 & A200;
  assign \new_[2155]_  = A301 & A300;
  assign \new_[2156]_  = ~A299 & \new_[2155]_ ;
  assign \new_[2157]_  = \new_[2156]_  & \new_[2151]_ ;
  assign \new_[2160]_  = ~A169 & A170;
  assign \new_[2164]_  = A199 & ~A166;
  assign \new_[2165]_  = A167 & \new_[2164]_ ;
  assign \new_[2166]_  = \new_[2165]_  & \new_[2160]_ ;
  assign \new_[2169]_  = A298 & A200;
  assign \new_[2173]_  = A302 & A300;
  assign \new_[2174]_  = ~A299 & \new_[2173]_ ;
  assign \new_[2175]_  = \new_[2174]_  & \new_[2169]_ ;
  assign \new_[2178]_  = ~A169 & A170;
  assign \new_[2182]_  = ~A200 & ~A166;
  assign \new_[2183]_  = A167 & \new_[2182]_ ;
  assign \new_[2184]_  = \new_[2183]_  & \new_[2178]_ ;
  assign \new_[2187]_  = A298 & ~A201;
  assign \new_[2191]_  = A301 & A300;
  assign \new_[2192]_  = ~A299 & \new_[2191]_ ;
  assign \new_[2193]_  = \new_[2192]_  & \new_[2187]_ ;
  assign \new_[2196]_  = ~A169 & A170;
  assign \new_[2200]_  = ~A200 & ~A166;
  assign \new_[2201]_  = A167 & \new_[2200]_ ;
  assign \new_[2202]_  = \new_[2201]_  & \new_[2196]_ ;
  assign \new_[2205]_  = A298 & ~A201;
  assign \new_[2209]_  = A302 & A300;
  assign \new_[2210]_  = ~A299 & \new_[2209]_ ;
  assign \new_[2211]_  = \new_[2210]_  & \new_[2205]_ ;
  assign \new_[2214]_  = ~A169 & A170;
  assign \new_[2218]_  = ~A199 & ~A166;
  assign \new_[2219]_  = A167 & \new_[2218]_ ;
  assign \new_[2220]_  = \new_[2219]_  & \new_[2214]_ ;
  assign \new_[2223]_  = A298 & ~A200;
  assign \new_[2227]_  = A301 & A300;
  assign \new_[2228]_  = ~A299 & \new_[2227]_ ;
  assign \new_[2229]_  = \new_[2228]_  & \new_[2223]_ ;
  assign \new_[2232]_  = ~A169 & A170;
  assign \new_[2236]_  = ~A199 & ~A166;
  assign \new_[2237]_  = A167 & \new_[2236]_ ;
  assign \new_[2238]_  = \new_[2237]_  & \new_[2232]_ ;
  assign \new_[2241]_  = A298 & ~A200;
  assign \new_[2245]_  = A302 & A300;
  assign \new_[2246]_  = ~A299 & \new_[2245]_ ;
  assign \new_[2247]_  = \new_[2246]_  & \new_[2241]_ ;
  assign \new_[2250]_  = ~A169 & A170;
  assign \new_[2254]_  = A199 & A166;
  assign \new_[2255]_  = ~A167 & \new_[2254]_ ;
  assign \new_[2256]_  = \new_[2255]_  & \new_[2250]_ ;
  assign \new_[2259]_  = A298 & A200;
  assign \new_[2263]_  = A301 & A300;
  assign \new_[2264]_  = ~A299 & \new_[2263]_ ;
  assign \new_[2265]_  = \new_[2264]_  & \new_[2259]_ ;
  assign \new_[2268]_  = ~A169 & A170;
  assign \new_[2272]_  = A199 & A166;
  assign \new_[2273]_  = ~A167 & \new_[2272]_ ;
  assign \new_[2274]_  = \new_[2273]_  & \new_[2268]_ ;
  assign \new_[2277]_  = A298 & A200;
  assign \new_[2281]_  = A302 & A300;
  assign \new_[2282]_  = ~A299 & \new_[2281]_ ;
  assign \new_[2283]_  = \new_[2282]_  & \new_[2277]_ ;
  assign \new_[2286]_  = ~A169 & A170;
  assign \new_[2290]_  = ~A200 & A166;
  assign \new_[2291]_  = ~A167 & \new_[2290]_ ;
  assign \new_[2292]_  = \new_[2291]_  & \new_[2286]_ ;
  assign \new_[2295]_  = A298 & ~A201;
  assign \new_[2299]_  = A301 & A300;
  assign \new_[2300]_  = ~A299 & \new_[2299]_ ;
  assign \new_[2301]_  = \new_[2300]_  & \new_[2295]_ ;
  assign \new_[2304]_  = ~A169 & A170;
  assign \new_[2308]_  = ~A200 & A166;
  assign \new_[2309]_  = ~A167 & \new_[2308]_ ;
  assign \new_[2310]_  = \new_[2309]_  & \new_[2304]_ ;
  assign \new_[2313]_  = A298 & ~A201;
  assign \new_[2317]_  = A302 & A300;
  assign \new_[2318]_  = ~A299 & \new_[2317]_ ;
  assign \new_[2319]_  = \new_[2318]_  & \new_[2313]_ ;
  assign \new_[2322]_  = ~A169 & A170;
  assign \new_[2326]_  = ~A199 & A166;
  assign \new_[2327]_  = ~A167 & \new_[2326]_ ;
  assign \new_[2328]_  = \new_[2327]_  & \new_[2322]_ ;
  assign \new_[2331]_  = A298 & ~A200;
  assign \new_[2335]_  = A301 & A300;
  assign \new_[2336]_  = ~A299 & \new_[2335]_ ;
  assign \new_[2337]_  = \new_[2336]_  & \new_[2331]_ ;
  assign \new_[2340]_  = ~A169 & A170;
  assign \new_[2344]_  = ~A199 & A166;
  assign \new_[2345]_  = ~A167 & \new_[2344]_ ;
  assign \new_[2346]_  = \new_[2345]_  & \new_[2340]_ ;
  assign \new_[2349]_  = A298 & ~A200;
  assign \new_[2353]_  = A302 & A300;
  assign \new_[2354]_  = ~A299 & \new_[2353]_ ;
  assign \new_[2355]_  = \new_[2354]_  & \new_[2349]_ ;
  assign \new_[2358]_  = ~A167 & A170;
  assign \new_[2362]_  = ~A200 & A199;
  assign \new_[2363]_  = ~A166 & \new_[2362]_ ;
  assign \new_[2364]_  = \new_[2363]_  & \new_[2358]_ ;
  assign \new_[2368]_  = A298 & A202;
  assign \new_[2369]_  = A201 & \new_[2368]_ ;
  assign \new_[2373]_  = A301 & A300;
  assign \new_[2374]_  = ~A299 & \new_[2373]_ ;
  assign \new_[2375]_  = \new_[2374]_  & \new_[2369]_ ;
  assign \new_[2378]_  = ~A167 & A170;
  assign \new_[2382]_  = ~A200 & A199;
  assign \new_[2383]_  = ~A166 & \new_[2382]_ ;
  assign \new_[2384]_  = \new_[2383]_  & \new_[2378]_ ;
  assign \new_[2388]_  = A298 & A202;
  assign \new_[2389]_  = A201 & \new_[2388]_ ;
  assign \new_[2393]_  = A302 & A300;
  assign \new_[2394]_  = ~A299 & \new_[2393]_ ;
  assign \new_[2395]_  = \new_[2394]_  & \new_[2389]_ ;
  assign \new_[2398]_  = ~A167 & A170;
  assign \new_[2402]_  = ~A200 & A199;
  assign \new_[2403]_  = ~A166 & \new_[2402]_ ;
  assign \new_[2404]_  = \new_[2403]_  & \new_[2398]_ ;
  assign \new_[2408]_  = A298 & A203;
  assign \new_[2409]_  = A201 & \new_[2408]_ ;
  assign \new_[2413]_  = A301 & A300;
  assign \new_[2414]_  = ~A299 & \new_[2413]_ ;
  assign \new_[2415]_  = \new_[2414]_  & \new_[2409]_ ;
  assign \new_[2418]_  = ~A167 & A170;
  assign \new_[2422]_  = ~A200 & A199;
  assign \new_[2423]_  = ~A166 & \new_[2422]_ ;
  assign \new_[2424]_  = \new_[2423]_  & \new_[2418]_ ;
  assign \new_[2428]_  = A298 & A203;
  assign \new_[2429]_  = A201 & \new_[2428]_ ;
  assign \new_[2433]_  = A302 & A300;
  assign \new_[2434]_  = ~A299 & \new_[2433]_ ;
  assign \new_[2435]_  = \new_[2434]_  & \new_[2429]_ ;
  assign \new_[2438]_  = A169 & A170;
  assign \new_[2442]_  = ~A200 & A199;
  assign \new_[2443]_  = ~A168 & \new_[2442]_ ;
  assign \new_[2444]_  = \new_[2443]_  & \new_[2438]_ ;
  assign \new_[2448]_  = A298 & A202;
  assign \new_[2449]_  = A201 & \new_[2448]_ ;
  assign \new_[2453]_  = A301 & A300;
  assign \new_[2454]_  = ~A299 & \new_[2453]_ ;
  assign \new_[2455]_  = \new_[2454]_  & \new_[2449]_ ;
  assign \new_[2458]_  = A169 & A170;
  assign \new_[2462]_  = ~A200 & A199;
  assign \new_[2463]_  = ~A168 & \new_[2462]_ ;
  assign \new_[2464]_  = \new_[2463]_  & \new_[2458]_ ;
  assign \new_[2468]_  = A298 & A202;
  assign \new_[2469]_  = A201 & \new_[2468]_ ;
  assign \new_[2473]_  = A302 & A300;
  assign \new_[2474]_  = ~A299 & \new_[2473]_ ;
  assign \new_[2475]_  = \new_[2474]_  & \new_[2469]_ ;
  assign \new_[2478]_  = A169 & A170;
  assign \new_[2482]_  = ~A200 & A199;
  assign \new_[2483]_  = ~A168 & \new_[2482]_ ;
  assign \new_[2484]_  = \new_[2483]_  & \new_[2478]_ ;
  assign \new_[2488]_  = A298 & A203;
  assign \new_[2489]_  = A201 & \new_[2488]_ ;
  assign \new_[2493]_  = A301 & A300;
  assign \new_[2494]_  = ~A299 & \new_[2493]_ ;
  assign \new_[2495]_  = \new_[2494]_  & \new_[2489]_ ;
  assign \new_[2498]_  = A169 & A170;
  assign \new_[2502]_  = ~A200 & A199;
  assign \new_[2503]_  = ~A168 & \new_[2502]_ ;
  assign \new_[2504]_  = \new_[2503]_  & \new_[2498]_ ;
  assign \new_[2508]_  = A298 & A203;
  assign \new_[2509]_  = A201 & \new_[2508]_ ;
  assign \new_[2513]_  = A302 & A300;
  assign \new_[2514]_  = ~A299 & \new_[2513]_ ;
  assign \new_[2515]_  = \new_[2514]_  & \new_[2509]_ ;
  assign \new_[2518]_  = A169 & ~A170;
  assign \new_[2522]_  = ~A200 & A166;
  assign \new_[2523]_  = A167 & \new_[2522]_ ;
  assign \new_[2524]_  = \new_[2523]_  & \new_[2518]_ ;
  assign \new_[2528]_  = A298 & ~A203;
  assign \new_[2529]_  = ~A202 & \new_[2528]_ ;
  assign \new_[2533]_  = A301 & A300;
  assign \new_[2534]_  = ~A299 & \new_[2533]_ ;
  assign \new_[2535]_  = \new_[2534]_  & \new_[2529]_ ;
  assign \new_[2538]_  = A169 & ~A170;
  assign \new_[2542]_  = ~A200 & A166;
  assign \new_[2543]_  = A167 & \new_[2542]_ ;
  assign \new_[2544]_  = \new_[2543]_  & \new_[2538]_ ;
  assign \new_[2548]_  = A298 & ~A203;
  assign \new_[2549]_  = ~A202 & \new_[2548]_ ;
  assign \new_[2553]_  = A302 & A300;
  assign \new_[2554]_  = ~A299 & \new_[2553]_ ;
  assign \new_[2555]_  = \new_[2554]_  & \new_[2549]_ ;
  assign \new_[2558]_  = A169 & ~A170;
  assign \new_[2562]_  = ~A200 & ~A166;
  assign \new_[2563]_  = ~A167 & \new_[2562]_ ;
  assign \new_[2564]_  = \new_[2563]_  & \new_[2558]_ ;
  assign \new_[2568]_  = A298 & ~A203;
  assign \new_[2569]_  = ~A202 & \new_[2568]_ ;
  assign \new_[2573]_  = A301 & A300;
  assign \new_[2574]_  = ~A299 & \new_[2573]_ ;
  assign \new_[2575]_  = \new_[2574]_  & \new_[2569]_ ;
  assign \new_[2578]_  = A169 & ~A170;
  assign \new_[2582]_  = ~A200 & ~A166;
  assign \new_[2583]_  = ~A167 & \new_[2582]_ ;
  assign \new_[2584]_  = \new_[2583]_  & \new_[2578]_ ;
  assign \new_[2588]_  = A298 & ~A203;
  assign \new_[2589]_  = ~A202 & \new_[2588]_ ;
  assign \new_[2593]_  = A302 & A300;
  assign \new_[2594]_  = ~A299 & \new_[2593]_ ;
  assign \new_[2595]_  = \new_[2594]_  & \new_[2589]_ ;
  assign \new_[2598]_  = ~A167 & ~A169;
  assign \new_[2602]_  = ~A200 & A199;
  assign \new_[2603]_  = ~A166 & \new_[2602]_ ;
  assign \new_[2604]_  = \new_[2603]_  & \new_[2598]_ ;
  assign \new_[2608]_  = A298 & A202;
  assign \new_[2609]_  = A201 & \new_[2608]_ ;
  assign \new_[2613]_  = A301 & A300;
  assign \new_[2614]_  = ~A299 & \new_[2613]_ ;
  assign \new_[2615]_  = \new_[2614]_  & \new_[2609]_ ;
  assign \new_[2618]_  = ~A167 & ~A169;
  assign \new_[2622]_  = ~A200 & A199;
  assign \new_[2623]_  = ~A166 & \new_[2622]_ ;
  assign \new_[2624]_  = \new_[2623]_  & \new_[2618]_ ;
  assign \new_[2628]_  = A298 & A202;
  assign \new_[2629]_  = A201 & \new_[2628]_ ;
  assign \new_[2633]_  = A302 & A300;
  assign \new_[2634]_  = ~A299 & \new_[2633]_ ;
  assign \new_[2635]_  = \new_[2634]_  & \new_[2629]_ ;
  assign \new_[2638]_  = ~A167 & ~A169;
  assign \new_[2642]_  = ~A200 & A199;
  assign \new_[2643]_  = ~A166 & \new_[2642]_ ;
  assign \new_[2644]_  = \new_[2643]_  & \new_[2638]_ ;
  assign \new_[2648]_  = A298 & A203;
  assign \new_[2649]_  = A201 & \new_[2648]_ ;
  assign \new_[2653]_  = A301 & A300;
  assign \new_[2654]_  = ~A299 & \new_[2653]_ ;
  assign \new_[2655]_  = \new_[2654]_  & \new_[2649]_ ;
  assign \new_[2658]_  = ~A167 & ~A169;
  assign \new_[2662]_  = ~A200 & A199;
  assign \new_[2663]_  = ~A166 & \new_[2662]_ ;
  assign \new_[2664]_  = \new_[2663]_  & \new_[2658]_ ;
  assign \new_[2668]_  = A298 & A203;
  assign \new_[2669]_  = A201 & \new_[2668]_ ;
  assign \new_[2673]_  = A302 & A300;
  assign \new_[2674]_  = ~A299 & \new_[2673]_ ;
  assign \new_[2675]_  = \new_[2674]_  & \new_[2669]_ ;
  assign \new_[2678]_  = ~A169 & A170;
  assign \new_[2682]_  = ~A200 & ~A166;
  assign \new_[2683]_  = A167 & \new_[2682]_ ;
  assign \new_[2684]_  = \new_[2683]_  & \new_[2678]_ ;
  assign \new_[2688]_  = A298 & ~A203;
  assign \new_[2689]_  = ~A202 & \new_[2688]_ ;
  assign \new_[2693]_  = A301 & A300;
  assign \new_[2694]_  = ~A299 & \new_[2693]_ ;
  assign \new_[2695]_  = \new_[2694]_  & \new_[2689]_ ;
  assign \new_[2698]_  = ~A169 & A170;
  assign \new_[2702]_  = ~A200 & ~A166;
  assign \new_[2703]_  = A167 & \new_[2702]_ ;
  assign \new_[2704]_  = \new_[2703]_  & \new_[2698]_ ;
  assign \new_[2708]_  = A298 & ~A203;
  assign \new_[2709]_  = ~A202 & \new_[2708]_ ;
  assign \new_[2713]_  = A302 & A300;
  assign \new_[2714]_  = ~A299 & \new_[2713]_ ;
  assign \new_[2715]_  = \new_[2714]_  & \new_[2709]_ ;
  assign \new_[2718]_  = ~A169 & A170;
  assign \new_[2722]_  = ~A200 & A166;
  assign \new_[2723]_  = ~A167 & \new_[2722]_ ;
  assign \new_[2724]_  = \new_[2723]_  & \new_[2718]_ ;
  assign \new_[2728]_  = A298 & ~A203;
  assign \new_[2729]_  = ~A202 & \new_[2728]_ ;
  assign \new_[2733]_  = A301 & A300;
  assign \new_[2734]_  = ~A299 & \new_[2733]_ ;
  assign \new_[2735]_  = \new_[2734]_  & \new_[2729]_ ;
  assign \new_[2738]_  = ~A169 & A170;
  assign \new_[2742]_  = ~A200 & A166;
  assign \new_[2743]_  = ~A167 & \new_[2742]_ ;
  assign \new_[2744]_  = \new_[2743]_  & \new_[2738]_ ;
  assign \new_[2748]_  = A298 & ~A203;
  assign \new_[2749]_  = ~A202 & \new_[2748]_ ;
  assign \new_[2753]_  = A302 & A300;
  assign \new_[2754]_  = ~A299 & \new_[2753]_ ;
  assign \new_[2755]_  = \new_[2754]_  & \new_[2749]_ ;
  assign \new_[2758]_  = ~A169 & ~A170;
  assign \new_[2762]_  = ~A200 & A199;
  assign \new_[2763]_  = ~A168 & \new_[2762]_ ;
  assign \new_[2764]_  = \new_[2763]_  & \new_[2758]_ ;
  assign \new_[2768]_  = A298 & A202;
  assign \new_[2769]_  = A201 & \new_[2768]_ ;
  assign \new_[2773]_  = A301 & A300;
  assign \new_[2774]_  = ~A299 & \new_[2773]_ ;
  assign \new_[2775]_  = \new_[2774]_  & \new_[2769]_ ;
  assign \new_[2778]_  = ~A169 & ~A170;
  assign \new_[2782]_  = ~A200 & A199;
  assign \new_[2783]_  = ~A168 & \new_[2782]_ ;
  assign \new_[2784]_  = \new_[2783]_  & \new_[2778]_ ;
  assign \new_[2788]_  = A298 & A202;
  assign \new_[2789]_  = A201 & \new_[2788]_ ;
  assign \new_[2793]_  = A302 & A300;
  assign \new_[2794]_  = ~A299 & \new_[2793]_ ;
  assign \new_[2795]_  = \new_[2794]_  & \new_[2789]_ ;
  assign \new_[2798]_  = ~A169 & ~A170;
  assign \new_[2802]_  = ~A200 & A199;
  assign \new_[2803]_  = ~A168 & \new_[2802]_ ;
  assign \new_[2804]_  = \new_[2803]_  & \new_[2798]_ ;
  assign \new_[2808]_  = A298 & A203;
  assign \new_[2809]_  = A201 & \new_[2808]_ ;
  assign \new_[2813]_  = A301 & A300;
  assign \new_[2814]_  = ~A299 & \new_[2813]_ ;
  assign \new_[2815]_  = \new_[2814]_  & \new_[2809]_ ;
  assign \new_[2818]_  = ~A169 & ~A170;
  assign \new_[2822]_  = ~A200 & A199;
  assign \new_[2823]_  = ~A168 & \new_[2822]_ ;
  assign \new_[2824]_  = \new_[2823]_  & \new_[2818]_ ;
  assign \new_[2828]_  = A298 & A203;
  assign \new_[2829]_  = A201 & \new_[2828]_ ;
  assign \new_[2833]_  = A302 & A300;
  assign \new_[2834]_  = ~A299 & \new_[2833]_ ;
  assign \new_[2835]_  = \new_[2834]_  & \new_[2829]_ ;
  assign \new_[2839]_  = A167 & ~A168;
  assign \new_[2840]_  = A169 & \new_[2839]_ ;
  assign \new_[2844]_  = ~A200 & A199;
  assign \new_[2845]_  = ~A166 & \new_[2844]_ ;
  assign \new_[2846]_  = \new_[2845]_  & \new_[2840]_ ;
  assign \new_[2850]_  = A298 & A202;
  assign \new_[2851]_  = A201 & \new_[2850]_ ;
  assign \new_[2855]_  = A301 & A300;
  assign \new_[2856]_  = ~A299 & \new_[2855]_ ;
  assign \new_[2857]_  = \new_[2856]_  & \new_[2851]_ ;
  assign \new_[2861]_  = A167 & ~A168;
  assign \new_[2862]_  = A169 & \new_[2861]_ ;
  assign \new_[2866]_  = ~A200 & A199;
  assign \new_[2867]_  = ~A166 & \new_[2866]_ ;
  assign \new_[2868]_  = \new_[2867]_  & \new_[2862]_ ;
  assign \new_[2872]_  = A298 & A202;
  assign \new_[2873]_  = A201 & \new_[2872]_ ;
  assign \new_[2877]_  = A302 & A300;
  assign \new_[2878]_  = ~A299 & \new_[2877]_ ;
  assign \new_[2879]_  = \new_[2878]_  & \new_[2873]_ ;
  assign \new_[2883]_  = A167 & ~A168;
  assign \new_[2884]_  = A169 & \new_[2883]_ ;
  assign \new_[2888]_  = ~A200 & A199;
  assign \new_[2889]_  = ~A166 & \new_[2888]_ ;
  assign \new_[2890]_  = \new_[2889]_  & \new_[2884]_ ;
  assign \new_[2894]_  = A298 & A203;
  assign \new_[2895]_  = A201 & \new_[2894]_ ;
  assign \new_[2899]_  = A301 & A300;
  assign \new_[2900]_  = ~A299 & \new_[2899]_ ;
  assign \new_[2901]_  = \new_[2900]_  & \new_[2895]_ ;
  assign \new_[2905]_  = A167 & ~A168;
  assign \new_[2906]_  = A169 & \new_[2905]_ ;
  assign \new_[2910]_  = ~A200 & A199;
  assign \new_[2911]_  = ~A166 & \new_[2910]_ ;
  assign \new_[2912]_  = \new_[2911]_  & \new_[2906]_ ;
  assign \new_[2916]_  = A298 & A203;
  assign \new_[2917]_  = A201 & \new_[2916]_ ;
  assign \new_[2921]_  = A302 & A300;
  assign \new_[2922]_  = ~A299 & \new_[2921]_ ;
  assign \new_[2923]_  = \new_[2922]_  & \new_[2917]_ ;
  assign \new_[2927]_  = ~A167 & ~A168;
  assign \new_[2928]_  = A169 & \new_[2927]_ ;
  assign \new_[2932]_  = ~A200 & A199;
  assign \new_[2933]_  = A166 & \new_[2932]_ ;
  assign \new_[2934]_  = \new_[2933]_  & \new_[2928]_ ;
  assign \new_[2938]_  = A298 & A202;
  assign \new_[2939]_  = A201 & \new_[2938]_ ;
  assign \new_[2943]_  = A301 & A300;
  assign \new_[2944]_  = ~A299 & \new_[2943]_ ;
  assign \new_[2945]_  = \new_[2944]_  & \new_[2939]_ ;
  assign \new_[2949]_  = ~A167 & ~A168;
  assign \new_[2950]_  = A169 & \new_[2949]_ ;
  assign \new_[2954]_  = ~A200 & A199;
  assign \new_[2955]_  = A166 & \new_[2954]_ ;
  assign \new_[2956]_  = \new_[2955]_  & \new_[2950]_ ;
  assign \new_[2960]_  = A298 & A202;
  assign \new_[2961]_  = A201 & \new_[2960]_ ;
  assign \new_[2965]_  = A302 & A300;
  assign \new_[2966]_  = ~A299 & \new_[2965]_ ;
  assign \new_[2967]_  = \new_[2966]_  & \new_[2961]_ ;
  assign \new_[2971]_  = ~A167 & ~A168;
  assign \new_[2972]_  = A169 & \new_[2971]_ ;
  assign \new_[2976]_  = ~A200 & A199;
  assign \new_[2977]_  = A166 & \new_[2976]_ ;
  assign \new_[2978]_  = \new_[2977]_  & \new_[2972]_ ;
  assign \new_[2982]_  = A298 & A203;
  assign \new_[2983]_  = A201 & \new_[2982]_ ;
  assign \new_[2987]_  = A301 & A300;
  assign \new_[2988]_  = ~A299 & \new_[2987]_ ;
  assign \new_[2989]_  = \new_[2988]_  & \new_[2983]_ ;
  assign \new_[2993]_  = ~A167 & ~A168;
  assign \new_[2994]_  = A169 & \new_[2993]_ ;
  assign \new_[2998]_  = ~A200 & A199;
  assign \new_[2999]_  = A166 & \new_[2998]_ ;
  assign \new_[3000]_  = \new_[2999]_  & \new_[2994]_ ;
  assign \new_[3004]_  = A298 & A203;
  assign \new_[3005]_  = A201 & \new_[3004]_ ;
  assign \new_[3009]_  = A302 & A300;
  assign \new_[3010]_  = ~A299 & \new_[3009]_ ;
  assign \new_[3011]_  = \new_[3010]_  & \new_[3005]_ ;
  assign \new_[3015]_  = A167 & ~A168;
  assign \new_[3016]_  = ~A169 & \new_[3015]_ ;
  assign \new_[3020]_  = ~A200 & A199;
  assign \new_[3021]_  = A166 & \new_[3020]_ ;
  assign \new_[3022]_  = \new_[3021]_  & \new_[3016]_ ;
  assign \new_[3026]_  = A298 & A202;
  assign \new_[3027]_  = A201 & \new_[3026]_ ;
  assign \new_[3031]_  = A301 & A300;
  assign \new_[3032]_  = ~A299 & \new_[3031]_ ;
  assign \new_[3033]_  = \new_[3032]_  & \new_[3027]_ ;
  assign \new_[3037]_  = A167 & ~A168;
  assign \new_[3038]_  = ~A169 & \new_[3037]_ ;
  assign \new_[3042]_  = ~A200 & A199;
  assign \new_[3043]_  = A166 & \new_[3042]_ ;
  assign \new_[3044]_  = \new_[3043]_  & \new_[3038]_ ;
  assign \new_[3048]_  = A298 & A202;
  assign \new_[3049]_  = A201 & \new_[3048]_ ;
  assign \new_[3053]_  = A302 & A300;
  assign \new_[3054]_  = ~A299 & \new_[3053]_ ;
  assign \new_[3055]_  = \new_[3054]_  & \new_[3049]_ ;
  assign \new_[3059]_  = A167 & ~A168;
  assign \new_[3060]_  = ~A169 & \new_[3059]_ ;
  assign \new_[3064]_  = ~A200 & A199;
  assign \new_[3065]_  = A166 & \new_[3064]_ ;
  assign \new_[3066]_  = \new_[3065]_  & \new_[3060]_ ;
  assign \new_[3070]_  = A298 & A203;
  assign \new_[3071]_  = A201 & \new_[3070]_ ;
  assign \new_[3075]_  = A301 & A300;
  assign \new_[3076]_  = ~A299 & \new_[3075]_ ;
  assign \new_[3077]_  = \new_[3076]_  & \new_[3071]_ ;
  assign \new_[3081]_  = A167 & ~A168;
  assign \new_[3082]_  = ~A169 & \new_[3081]_ ;
  assign \new_[3086]_  = ~A200 & A199;
  assign \new_[3087]_  = A166 & \new_[3086]_ ;
  assign \new_[3088]_  = \new_[3087]_  & \new_[3082]_ ;
  assign \new_[3092]_  = A298 & A203;
  assign \new_[3093]_  = A201 & \new_[3092]_ ;
  assign \new_[3097]_  = A302 & A300;
  assign \new_[3098]_  = ~A299 & \new_[3097]_ ;
  assign \new_[3099]_  = \new_[3098]_  & \new_[3093]_ ;
endmodule


