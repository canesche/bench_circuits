module top ( 
    i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_  );
  input  i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_;
  wire new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_, new_n15_,
    new_n16_, new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_,
    new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_,
    new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_;
  assign new_n9_ = ~i_3_ & ~i_4_;
  assign new_n10_ = i_1_ & ~i_2_;
  assign new_n11_ = ~i_0_ & new_n10_;
  assign new_n12_ = new_n9_ & new_n11_;
  assign new_n13_ = i_3_ & ~i_4_;
  assign new_n14_ = ~i_1_ & ~i_2_;
  assign new_n15_ = ~i_0_ & new_n14_;
  assign new_n16_ = new_n13_ & new_n15_;
  assign new_n17_ = i_3_ & i_4_;
  assign new_n18_ = i_1_ & i_2_;
  assign new_n19_ = i_0_ & new_n18_;
  assign new_n20_ = new_n17_ & new_n19_;
  assign new_n21_ = ~new_n12_ & ~new_n16_;
  assign new_n22_ = ~new_n20_ & new_n21_;
  assign new_n23_ = ~i_0_ & new_n18_;
  assign new_n24_ = new_n13_ & new_n23_;
  assign new_n25_ = ~i_1_ & i_2_;
  assign new_n26_ = ~i_0_ & new_n25_;
  assign new_n27_ = new_n17_ & new_n26_;
  assign new_n28_ = new_n9_ & new_n26_;
  assign new_n29_ = new_n9_ & new_n19_;
  assign new_n30_ = ~new_n27_ & ~new_n28_;
  assign new_n31_ = ~new_n29_ & new_n30_;
  assign new_n32_ = new_n22_ & ~new_n24_;
  assign new_n33_ = new_n31_ & new_n32_;
  assign new_n34_ = i_0_ & new_n14_;
  assign new_n35_ = new_n9_ & new_n34_;
  assign new_n36_ = i_0_ & new_n25_;
  assign new_n37_ = new_n13_ & new_n36_;
  assign new_n38_ = ~i_3_ & i_4_;
  assign new_n39_ = i_0_ & new_n10_;
  assign new_n40_ = new_n38_ & new_n39_;
  assign new_n41_ = ~new_n35_ & ~new_n37_;
  assign new_n42_ = ~new_n40_ & new_n41_;
  assign new_n43_ = new_n23_ & new_n38_;
  assign new_n44_ = new_n13_ & new_n39_;
  assign new_n45_ = new_n11_ & new_n17_;
  assign new_n46_ = ~new_n43_ & ~new_n44_;
  assign new_n47_ = ~new_n45_ & new_n46_;
  assign new_n48_ = new_n36_ & new_n38_;
  assign new_n49_ = new_n15_ & new_n38_;
  assign new_n50_ = new_n17_ & new_n34_;
  assign new_n51_ = ~new_n48_ & ~new_n49_;
  assign new_n52_ = ~new_n50_ & new_n51_;
  assign new_n53_ = new_n42_ & new_n47_;
  assign new_n54_ = new_n52_ & new_n53_;
  assign o_1_ = ~new_n33_ | ~new_n54_;
  assign new_n56_ = ~i_3_ & i_1_;
  assign new_n57_ = ~i_0_ & new_n56_;
  assign new_n58_ = i_4_ & new_n57_;
  assign new_n59_ = i_3_ & i_2_;
  assign new_n60_ = ~i_1_ & new_n59_;
  assign new_n61_ = ~i_4_ & new_n60_;
  assign new_n62_ = ~new_n58_ & ~new_n61_;
  assign new_n63_ = ~i_4_ & new_n23_;
  assign new_n64_ = ~i_4_ & new_n39_;
  assign new_n65_ = i_3_ & new_n34_;
  assign new_n66_ = ~new_n63_ & ~new_n64_;
  assign new_n67_ = ~new_n65_ & new_n66_;
  assign new_n68_ = ~i_3_ & ~i_2_;
  assign new_n69_ = i_0_ & new_n68_;
  assign new_n70_ = i_4_ & new_n69_;
  assign new_n71_ = i_4_ & new_n26_;
  assign new_n72_ = ~i_3_ & i_2_;
  assign new_n73_ = i_0_ & new_n72_;
  assign new_n74_ = ~i_4_ & new_n73_;
  assign new_n75_ = ~new_n70_ & ~new_n71_;
  assign new_n76_ = ~new_n74_ & new_n75_;
  assign new_n77_ = i_3_ & ~i_2_;
  assign new_n78_ = i_1_ & new_n77_;
  assign new_n79_ = ~i_4_ & new_n78_;
  assign new_n80_ = ~i_0_ & new_n77_;
  assign new_n81_ = i_4_ & new_n80_;
  assign new_n82_ = ~i_1_ & new_n72_;
  assign new_n83_ = i_4_ & new_n82_;
  assign new_n84_ = ~new_n79_ & ~new_n81_;
  assign new_n85_ = ~new_n83_ & new_n84_;
  assign new_n86_ = new_n67_ & new_n76_;
  assign new_n87_ = new_n85_ & new_n86_;
  assign o_2_ = ~new_n62_ | ~new_n87_;
  assign new_n89_ = i_0_ & new_n59_;
  assign new_n90_ = i_4_ & new_n89_;
  assign new_n91_ = i_3_ & i_1_;
  assign new_n92_ = i_0_ & new_n91_;
  assign new_n93_ = i_4_ & new_n92_;
  assign new_n94_ = ~new_n90_ & ~new_n93_;
  assign new_n95_ = i_4_ & new_n19_;
  assign new_n96_ = i_3_ & new_n19_;
  assign new_n97_ = i_1_ & new_n59_;
  assign new_n98_ = i_4_ & new_n97_;
  assign new_n99_ = ~new_n95_ & ~new_n96_;
  assign new_n100_ = ~new_n98_ & new_n99_;
  assign o_0_ = ~new_n94_ | ~new_n100_;
endmodule

