module top ( 
    pp, pa0, pq, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0, px,
    pi0, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po,
    pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0  );
  input  pp, pa0, pq, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw,
    ph0, px, pi0, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl,
    pm, pn, po;
  output pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0;
  wire new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_;
  assign new_n45_ = pc & ~pd;
  assign new_n46_ = ~pi0 & pc;
  assign new_n47_ = ~pi0 & ~pd;
  assign new_n48_ = ~new_n45_ & ~new_n46_;
  assign new_n49_ = ~new_n47_ & new_n48_;
  assign new_n50_ = ~pd & new_n49_;
  assign new_n51_ = pc & new_n49_;
  assign new_n52_ = ph0 & new_n49_;
  assign new_n53_ = ~new_n50_ & ~new_n51_;
  assign new_n54_ = ~new_n52_ & new_n53_;
  assign new_n55_ = pd & new_n54_;
  assign new_n56_ = ~pc & new_n54_;
  assign new_n57_ = ~ph0 & new_n54_;
  assign new_n58_ = ~new_n55_ & ~new_n56_;
  assign pk0 = new_n57_ | ~new_n58_;
  assign new_n60_ = pi & ~pj;
  assign new_n61_ = pd & pe;
  assign new_n62_ = pe & ph;
  assign new_n63_ = pd & ph;
  assign new_n64_ = ~new_n61_ & ~new_n62_;
  assign new_n65_ = ~new_n63_ & new_n64_;
  assign new_n66_ = pe & new_n65_;
  assign new_n67_ = pd & new_n65_;
  assign new_n68_ = ph & new_n65_;
  assign new_n69_ = ~new_n66_ & ~new_n67_;
  assign new_n70_ = ~new_n68_ & new_n69_;
  assign new_n71_ = ~pe & new_n70_;
  assign new_n72_ = ~pd & new_n70_;
  assign new_n73_ = ~ph & new_n70_;
  assign new_n74_ = ~new_n71_ & ~new_n72_;
  assign new_n75_ = ~new_n73_ & new_n74_;
  assign new_n76_ = pc & new_n75_;
  assign new_n77_ = ~pd & pe;
  assign new_n78_ = ~pd & ph;
  assign new_n79_ = ~new_n62_ & ~new_n77_;
  assign new_n80_ = ~new_n78_ & new_n79_;
  assign new_n81_ = pe & new_n80_;
  assign new_n82_ = ~pd & new_n80_;
  assign new_n83_ = ph & new_n80_;
  assign new_n84_ = ~new_n81_ & ~new_n82_;
  assign new_n85_ = ~new_n83_ & new_n84_;
  assign new_n86_ = ~pe & new_n85_;
  assign new_n87_ = pd & new_n85_;
  assign new_n88_ = ~ph & new_n85_;
  assign new_n89_ = ~new_n86_ & ~new_n87_;
  assign new_n90_ = ~new_n88_ & new_n89_;
  assign new_n91_ = new_n75_ & new_n90_;
  assign new_n92_ = ~pc & new_n90_;
  assign new_n93_ = ~new_n76_ & ~new_n91_;
  assign new_n94_ = ~new_n92_ & new_n93_;
  assign new_n95_ = new_n60_ & ~new_n94_;
  assign new_n96_ = pb & new_n95_;
  assign new_n97_ = ~pe & ~ph;
  assign new_n98_ = ~pc & pg;
  assign new_n99_ = ~pd & pf;
  assign new_n100_ = ~new_n97_ & ~new_n98_;
  assign new_n101_ = ~new_n99_ & new_n100_;
  assign new_n102_ = ~pe & new_n101_;
  assign new_n103_ = ~ph & new_n101_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = pd & new_n104_;
  assign new_n106_ = ~pg & new_n105_;
  assign new_n107_ = pc & new_n105_;
  assign new_n108_ = ~pf & new_n104_;
  assign new_n109_ = pc & new_n108_;
  assign new_n110_ = pe & ~ph;
  assign new_n111_ = ~pf & new_n110_;
  assign new_n112_ = pd & new_n110_;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = pe & new_n113_;
  assign new_n115_ = ~pf & new_n114_;
  assign new_n116_ = pd & new_n114_;
  assign new_n117_ = ~ph & new_n113_;
  assign new_n118_ = pd & new_n117_;
  assign new_n119_ = ~new_n62_ & ~new_n97_;
  assign new_n120_ = new_n117_ & new_n119_;
  assign new_n121_ = ~pf & new_n117_;
  assign new_n122_ = new_n99_ & new_n113_;
  assign new_n123_ = pd & new_n122_;
  assign new_n124_ = new_n119_ & new_n122_;
  assign new_n125_ = new_n114_ & new_n119_;
  assign new_n126_ = ~pf & new_n122_;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_ = ~new_n123_ & ~new_n124_;
  assign new_n129_ = new_n127_ & new_n128_;
  assign new_n130_ = ~new_n115_ & ~new_n116_;
  assign new_n131_ = ~new_n118_ & new_n130_;
  assign new_n132_ = ~new_n120_ & ~new_n121_;
  assign new_n133_ = new_n131_ & new_n132_;
  assign new_n134_ = new_n129_ & new_n133_;
  assign new_n135_ = new_n108_ & new_n134_;
  assign new_n136_ = ~pg & new_n108_;
  assign new_n137_ = ~pg & ~ph;
  assign new_n138_ = ~pe & new_n137_;
  assign new_n139_ = ~pg & ph;
  assign new_n140_ = pe & new_n139_;
  assign new_n141_ = pc & new_n97_;
  assign new_n142_ = pc & new_n62_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = ~new_n138_ & ~new_n140_;
  assign new_n145_ = new_n143_ & new_n144_;
  assign new_n146_ = new_n104_ & new_n145_;
  assign new_n147_ = pc & new_n146_;
  assign new_n148_ = new_n134_ & new_n146_;
  assign new_n149_ = new_n105_ & new_n134_;
  assign new_n150_ = ~pg & new_n146_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = ~new_n147_ & ~new_n148_;
  assign new_n153_ = new_n151_ & new_n152_;
  assign new_n154_ = ~new_n106_ & ~new_n107_;
  assign new_n155_ = ~new_n109_ & new_n154_;
  assign new_n156_ = ~new_n135_ & ~new_n136_;
  assign new_n157_ = new_n155_ & new_n156_;
  assign new_n158_ = new_n153_ & new_n157_;
  assign new_n159_ = new_n60_ & new_n158_;
  assign new_n160_ = ~pb & new_n159_;
  assign pl0 = new_n96_ | new_n160_;
  assign new_n162_ = ~pa0 & pz;
  assign new_n163_ = ~pc0 & new_n162_;
  assign new_n164_ = pc & pd;
  assign new_n165_ = ~ps & ~px;
  assign new_n166_ = ~pt & ~py;
  assign new_n167_ = pr & pv;
  assign new_n168_ = pu & new_n167_;
  assign new_n169_ = pq & pw;
  assign new_n170_ = pp & new_n169_;
  assign new_n171_ = pq & pr;
  assign new_n172_ = pu & new_n171_;
  assign new_n173_ = pp & new_n167_;
  assign new_n174_ = pp & new_n171_;
  assign new_n175_ = pv & pw;
  assign new_n176_ = pu & new_n175_;
  assign new_n177_ = pu & new_n169_;
  assign new_n178_ = pp & new_n175_;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = ~new_n174_ & ~new_n176_;
  assign new_n181_ = new_n179_ & new_n180_;
  assign new_n182_ = ~new_n172_ & ~new_n173_;
  assign new_n183_ = ~new_n168_ & ~new_n170_;
  assign new_n184_ = new_n182_ & new_n183_;
  assign new_n185_ = new_n181_ & new_n184_;
  assign new_n186_ = ~new_n165_ & ~new_n166_;
  assign new_n187_ = ~new_n185_ & new_n186_;
  assign new_n188_ = ~new_n164_ & ~new_n187_;
  assign new_n189_ = new_n163_ & new_n188_;
  assign pm0 = pb & new_n189_;
  assign new_n191_ = ~pq & ~pv;
  assign new_n192_ = ~pr & ~pw;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = ~new_n165_ & new_n193_;
  assign new_n195_ = pp & new_n194_;
  assign new_n196_ = pt & new_n195_;
  assign new_n197_ = pu & new_n194_;
  assign new_n198_ = pt & new_n197_;
  assign new_n199_ = py & new_n195_;
  assign new_n200_ = py & new_n197_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~new_n196_ & ~new_n198_;
  assign new_n203_ = new_n201_ & new_n202_;
  assign new_n204_ = ~pd & new_n203_;
  assign new_n205_ = ~pp & ~pu;
  assign new_n206_ = ~new_n165_ & ~new_n192_;
  assign new_n207_ = ~new_n205_ & new_n206_;
  assign new_n208_ = pq & new_n207_;
  assign new_n209_ = pt & new_n208_;
  assign new_n210_ = pv & new_n207_;
  assign new_n211_ = pt & new_n210_;
  assign new_n212_ = py & new_n208_;
  assign new_n213_ = py & new_n210_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~new_n209_ & ~new_n211_;
  assign new_n216_ = new_n214_ & new_n215_;
  assign new_n217_ = ~pc & new_n216_;
  assign new_n218_ = ~new_n204_ & ~new_n217_;
  assign new_n219_ = pd0 & new_n218_;
  assign new_n220_ = new_n186_ & ~new_n205_;
  assign new_n221_ = pq & new_n220_;
  assign new_n222_ = pr & new_n221_;
  assign new_n223_ = pv & new_n220_;
  assign new_n224_ = pr & new_n223_;
  assign new_n225_ = pw & new_n221_;
  assign new_n226_ = pw & new_n223_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = ~new_n222_ & ~new_n224_;
  assign new_n229_ = new_n227_ & new_n228_;
  assign new_n230_ = ~pd & new_n229_;
  assign new_n231_ = ~pc & new_n229_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = pc0 & new_n232_;
  assign new_n234_ = ~pc0 & ~pd0;
  assign new_n235_ = ~pc0 & new_n218_;
  assign new_n236_ = pc0 & pd0;
  assign new_n237_ = ~pd0 & new_n232_;
  assign new_n238_ = new_n218_ & new_n232_;
  assign new_n239_ = ~new_n234_ & ~new_n235_;
  assign new_n240_ = ~new_n219_ & ~new_n233_;
  assign new_n241_ = new_n239_ & new_n240_;
  assign new_n242_ = ~new_n236_ & ~new_n237_;
  assign new_n243_ = ~new_n238_ & new_n242_;
  assign new_n244_ = new_n241_ & new_n243_;
  assign new_n245_ = new_n162_ & new_n244_;
  assign pn0 = pb & new_n245_;
  assign new_n247_ = px & new_n169_;
  assign new_n248_ = ps & new_n167_;
  assign new_n249_ = px & new_n171_;
  assign new_n250_ = ps & new_n169_;
  assign new_n251_ = ps & new_n171_;
  assign new_n252_ = px & new_n175_;
  assign new_n253_ = px & new_n167_;
  assign new_n254_ = ps & new_n175_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~new_n251_ & ~new_n252_;
  assign new_n257_ = new_n255_ & new_n256_;
  assign new_n258_ = ~new_n249_ & ~new_n250_;
  assign new_n259_ = ~new_n247_ & ~new_n248_;
  assign new_n260_ = new_n258_ & new_n259_;
  assign new_n261_ = new_n257_ & new_n260_;
  assign new_n262_ = ~new_n166_ & ~new_n205_;
  assign new_n263_ = ~new_n261_ & new_n262_;
  assign new_n264_ = ps & pv;
  assign new_n265_ = pu & new_n264_;
  assign new_n266_ = pq & px;
  assign new_n267_ = pp & new_n266_;
  assign new_n268_ = pq & ps;
  assign new_n269_ = pu & new_n268_;
  assign new_n270_ = pp & new_n264_;
  assign new_n271_ = pp & new_n268_;
  assign new_n272_ = pv & px;
  assign new_n273_ = pu & new_n272_;
  assign new_n274_ = pu & new_n266_;
  assign new_n275_ = pp & new_n272_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = ~new_n271_ & ~new_n273_;
  assign new_n278_ = new_n276_ & new_n277_;
  assign new_n279_ = ~new_n269_ & ~new_n270_;
  assign new_n280_ = ~new_n265_ & ~new_n267_;
  assign new_n281_ = new_n279_ & new_n280_;
  assign new_n282_ = new_n278_ & new_n281_;
  assign new_n283_ = ~new_n166_ & ~new_n192_;
  assign new_n284_ = ~new_n282_ & new_n283_;
  assign new_n285_ = new_n263_ & new_n284_;
  assign new_n286_ = pd0 & new_n284_;
  assign new_n287_ = pc0 & new_n263_;
  assign new_n288_ = ~new_n236_ & ~new_n287_;
  assign new_n289_ = ~new_n285_ & ~new_n286_;
  assign new_n290_ = new_n288_ & new_n289_;
  assign new_n291_ = ~pd & new_n290_;
  assign new_n292_ = pe0 & new_n291_;
  assign new_n293_ = pc & ~new_n292_;
  assign new_n294_ = ~pc0 & new_n293_;
  assign new_n295_ = pd0 & ~pe0;
  assign new_n296_ = new_n293_ & ~new_n295_;
  assign new_n297_ = ~pe0 & ~new_n292_;
  assign new_n298_ = ~new_n295_ & new_n297_;
  assign new_n299_ = new_n232_ & new_n297_;
  assign new_n300_ = ~pc0 & new_n297_;
  assign new_n301_ = ~pd0 & new_n216_;
  assign new_n302_ = ~new_n165_ & ~new_n191_;
  assign new_n303_ = ~new_n205_ & new_n302_;
  assign new_n304_ = pt & new_n303_;
  assign new_n305_ = pr & new_n304_;
  assign new_n306_ = py & new_n303_;
  assign new_n307_ = pr & new_n306_;
  assign new_n308_ = pw & new_n304_;
  assign new_n309_ = pw & new_n306_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~new_n305_ & ~new_n307_;
  assign new_n312_ = new_n310_ & new_n311_;
  assign new_n313_ = ~pc0 & new_n312_;
  assign new_n314_ = ~new_n301_ & ~new_n313_;
  assign new_n315_ = ~new_n292_ & new_n314_;
  assign new_n316_ = ~new_n295_ & new_n315_;
  assign new_n317_ = new_n232_ & new_n315_;
  assign new_n318_ = new_n232_ & new_n293_;
  assign new_n319_ = ~pc0 & new_n315_;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = ~new_n316_ & ~new_n317_;
  assign new_n322_ = new_n320_ & new_n321_;
  assign new_n323_ = ~new_n294_ & ~new_n296_;
  assign new_n324_ = ~new_n298_ & new_n323_;
  assign new_n325_ = ~new_n299_ & ~new_n300_;
  assign new_n326_ = new_n324_ & new_n325_;
  assign new_n327_ = new_n322_ & new_n326_;
  assign new_n328_ = new_n162_ & new_n327_;
  assign po0 = pb & new_n328_;
  assign new_n330_ = px & py;
  assign new_n331_ = ps & py;
  assign new_n332_ = pt & px;
  assign new_n333_ = ps & pt;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~new_n330_ & ~new_n331_;
  assign new_n336_ = new_n334_ & new_n335_;
  assign new_n337_ = pw & new_n330_;
  assign new_n338_ = pw & new_n332_;
  assign new_n339_ = pd0 & pe0;
  assign new_n340_ = pc0 & new_n339_;
  assign new_n341_ = ~new_n337_ & ~new_n338_;
  assign new_n342_ = ~new_n340_ & new_n341_;
  assign new_n343_ = new_n336_ & new_n342_;
  assign new_n344_ = ~pw & new_n343_;
  assign new_n345_ = ~ps & new_n343_;
  assign new_n346_ = ~pr & new_n342_;
  assign new_n347_ = ~ps & new_n346_;
  assign new_n348_ = new_n166_ & new_n346_;
  assign new_n349_ = ~pw & new_n346_;
  assign new_n350_ = new_n166_ & new_n343_;
  assign new_n351_ = ~new_n344_ & ~new_n345_;
  assign new_n352_ = ~new_n347_ & new_n351_;
  assign new_n353_ = ~new_n348_ & ~new_n349_;
  assign new_n354_ = ~new_n350_ & new_n353_;
  assign new_n355_ = new_n352_ & new_n354_;
  assign new_n356_ = pv & new_n355_;
  assign new_n357_ = pp & new_n356_;
  assign new_n358_ = pu & new_n356_;
  assign new_n359_ = pq & new_n355_;
  assign new_n360_ = pp & new_n359_;
  assign new_n361_ = pu & new_n359_;
  assign new_n362_ = pe0 & new_n236_;
  assign new_n363_ = new_n355_ & new_n362_;
  assign new_n364_ = ~new_n357_ & ~new_n358_;
  assign new_n365_ = ~new_n360_ & new_n364_;
  assign new_n366_ = ~new_n361_ & ~new_n363_;
  assign new_n367_ = new_n365_ & new_n366_;
  assign new_n368_ = ~pd & new_n367_;
  assign new_n369_ = pf0 & new_n368_;
  assign new_n370_ = pc & ~new_n369_;
  assign new_n371_ = ~pc0 & new_n370_;
  assign new_n372_ = ~pf0 & new_n339_;
  assign new_n373_ = new_n370_ & ~new_n372_;
  assign new_n374_ = ~pf0 & ~new_n369_;
  assign new_n375_ = ~new_n372_ & new_n374_;
  assign new_n376_ = new_n232_ & new_n374_;
  assign new_n377_ = ~pc0 & new_n374_;
  assign new_n378_ = ~pu & ~new_n362_;
  assign new_n379_ = ~pp & new_n378_;
  assign new_n380_ = ~pv & ~new_n362_;
  assign new_n381_ = ~pq & new_n380_;
  assign new_n382_ = pr & new_n186_;
  assign new_n383_ = ps & ~new_n166_;
  assign new_n384_ = pw & new_n383_;
  assign new_n385_ = ~pd0 & ~px;
  assign new_n386_ = ~pe0 & ~pw;
  assign new_n387_ = ~pc0 & ~px;
  assign new_n388_ = ~pd0 & ~pw;
  assign new_n389_ = ~pc0 & ~pw;
  assign new_n390_ = ~pd0 & ~py;
  assign new_n391_ = ~pt & new_n390_;
  assign new_n392_ = ~pe0 & ~py;
  assign new_n393_ = ~pt & new_n392_;
  assign new_n394_ = ~pe0 & ~px;
  assign new_n395_ = ~pc0 & ~py;
  assign new_n396_ = ~pt & new_n395_;
  assign new_n397_ = ~new_n394_ & ~new_n396_;
  assign new_n398_ = ~new_n391_ & ~new_n393_;
  assign new_n399_ = new_n397_ & new_n398_;
  assign new_n400_ = ~new_n385_ & ~new_n386_;
  assign new_n401_ = ~new_n387_ & new_n400_;
  assign new_n402_ = ~new_n388_ & ~new_n389_;
  assign new_n403_ = new_n401_ & new_n402_;
  assign new_n404_ = new_n399_ & new_n403_;
  assign new_n405_ = ~new_n382_ & ~new_n384_;
  assign new_n406_ = ~new_n404_ & new_n405_;
  assign new_n407_ = ~new_n379_ & ~new_n381_;
  assign new_n408_ = ~new_n406_ & new_n407_;
  assign new_n409_ = ~new_n369_ & new_n408_;
  assign new_n410_ = ~new_n372_ & new_n409_;
  assign new_n411_ = new_n232_ & new_n409_;
  assign new_n412_ = new_n232_ & new_n370_;
  assign new_n413_ = ~pc0 & new_n409_;
  assign new_n414_ = ~new_n412_ & ~new_n413_;
  assign new_n415_ = ~new_n410_ & ~new_n411_;
  assign new_n416_ = new_n414_ & new_n415_;
  assign new_n417_ = ~new_n371_ & ~new_n373_;
  assign new_n418_ = ~new_n375_ & new_n417_;
  assign new_n419_ = ~new_n376_ & ~new_n377_;
  assign new_n420_ = new_n418_ & new_n419_;
  assign new_n421_ = new_n416_ & new_n420_;
  assign new_n422_ = new_n162_ & new_n421_;
  assign pp0 = pb & new_n422_;
  assign new_n424_ = pr & px;
  assign new_n425_ = py & new_n424_;
  assign new_n426_ = ps & pw;
  assign new_n427_ = pt & new_n426_;
  assign new_n428_ = pr & ps;
  assign new_n429_ = py & new_n428_;
  assign new_n430_ = pt & new_n424_;
  assign new_n431_ = pt & new_n428_;
  assign new_n432_ = pw & px;
  assign new_n433_ = py & new_n432_;
  assign new_n434_ = py & new_n426_;
  assign new_n435_ = pt & new_n432_;
  assign new_n436_ = ~new_n434_ & ~new_n435_;
  assign new_n437_ = ~new_n431_ & ~new_n433_;
  assign new_n438_ = new_n436_ & new_n437_;
  assign new_n439_ = ~new_n429_ & ~new_n430_;
  assign new_n440_ = ~new_n425_ & ~new_n427_;
  assign new_n441_ = new_n439_ & new_n440_;
  assign new_n442_ = new_n438_ & new_n441_;
  assign new_n443_ = pv & ~new_n165_;
  assign new_n444_ = pw & new_n443_;
  assign new_n445_ = pt & new_n444_;
  assign new_n446_ = py & new_n444_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = new_n442_ & new_n447_;
  assign new_n449_ = ~pv & new_n448_;
  assign new_n450_ = ~pr & new_n448_;
  assign new_n451_ = ~pq & new_n447_;
  assign new_n452_ = ~pr & new_n451_;
  assign new_n453_ = new_n336_ & new_n451_;
  assign new_n454_ = ~pv & new_n451_;
  assign new_n455_ = new_n336_ & new_n448_;
  assign new_n456_ = ~new_n449_ & ~new_n450_;
  assign new_n457_ = ~new_n452_ & new_n456_;
  assign new_n458_ = ~new_n453_ & ~new_n454_;
  assign new_n459_ = ~new_n455_ & new_n458_;
  assign new_n460_ = new_n457_ & new_n459_;
  assign new_n461_ = pp & new_n460_;
  assign new_n462_ = ~new_n166_ & new_n206_;
  assign new_n463_ = pq & new_n462_;
  assign new_n464_ = pu & new_n463_;
  assign new_n465_ = pe0 & pf0;
  assign new_n466_ = pc0 & new_n465_;
  assign new_n467_ = pd0 & new_n466_;
  assign new_n468_ = pf0 & new_n362_;
  assign new_n469_ = ~pg0 & new_n468_;
  assign new_n470_ = ~pa0 & ~new_n469_;
  assign new_n471_ = ~pc & new_n470_;
  assign new_n472_ = ~pd & new_n470_;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign new_n474_ = pz & ~new_n473_;
  assign new_n475_ = pb & new_n474_;
  assign new_n476_ = new_n467_ & new_n475_;
  assign new_n477_ = ~pv & new_n476_;
  assign new_n478_ = ~pu & new_n476_;
  assign new_n479_ = ~pg0 & new_n475_;
  assign new_n480_ = ~pu & new_n479_;
  assign new_n481_ = new_n442_ & new_n479_;
  assign new_n482_ = ~pv & new_n479_;
  assign new_n483_ = new_n442_ & new_n476_;
  assign new_n484_ = ~new_n477_ & ~new_n478_;
  assign new_n485_ = ~new_n480_ & new_n484_;
  assign new_n486_ = ~new_n481_ & ~new_n482_;
  assign new_n487_ = ~new_n483_ & new_n486_;
  assign new_n488_ = new_n485_ & new_n487_;
  assign new_n489_ = ~new_n461_ & ~new_n464_;
  assign pq0 = new_n488_ | ~new_n489_;
  assign new_n491_ = ~pl & new_n333_;
  assign new_n492_ = pr & new_n491_;
  assign new_n493_ = ~pq & ~new_n492_;
  assign new_n494_ = ps & ~pm;
  assign new_n495_ = pt & new_n494_;
  assign new_n496_ = ~pr & ~new_n495_;
  assign new_n497_ = ps & ~po;
  assign new_n498_ = pt & ~pn;
  assign new_n499_ = ~new_n333_ & ~new_n497_;
  assign new_n500_ = ~new_n498_ & new_n499_;
  assign new_n501_ = ~new_n493_ & ~new_n496_;
  assign new_n502_ = ~new_n500_ & new_n501_;
  assign new_n503_ = pp & new_n502_;
  assign new_n504_ = pq & new_n333_;
  assign new_n505_ = pr & new_n504_;
  assign new_n506_ = ~pp & ~new_n505_;
  assign new_n507_ = ~pe0 & ~pf0;
  assign new_n508_ = ~pd0 & ~pf0;
  assign new_n509_ = ~pc0 & new_n508_;
  assign new_n510_ = pq & ~pk;
  assign new_n511_ = pr & new_n510_;
  assign new_n512_ = ps & new_n511_;
  assign new_n513_ = pt & new_n512_;
  assign new_n514_ = ~pr & ~pt;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign new_n516_ = pg0 & new_n515_;
  assign new_n517_ = pt & new_n516_;
  assign new_n518_ = pr & new_n517_;
  assign new_n519_ = ps & new_n516_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = ~new_n507_ & ~new_n509_;
  assign new_n522_ = ~new_n520_ & new_n521_;
  assign new_n523_ = new_n431_ & new_n522_;
  assign new_n524_ = ~pf0 & new_n523_;
  assign new_n525_ = ~pe0 & new_n523_;
  assign new_n526_ = pq & new_n522_;
  assign new_n527_ = ~pe0 & new_n526_;
  assign new_n528_ = new_n234_ & new_n526_;
  assign new_n529_ = ~pf0 & new_n526_;
  assign new_n530_ = new_n234_ & new_n523_;
  assign new_n531_ = ~new_n524_ & ~new_n525_;
  assign new_n532_ = ~new_n527_ & new_n531_;
  assign new_n533_ = ~new_n528_ & ~new_n529_;
  assign new_n534_ = ~new_n530_ & new_n533_;
  assign new_n535_ = new_n532_ & new_n534_;
  assign new_n536_ = ~new_n503_ & ~new_n506_;
  assign new_n537_ = ~new_n535_ & new_n536_;
  assign new_n538_ = ph0 & new_n537_;
  assign new_n539_ = ~pp & pk;
  assign new_n540_ = pq & new_n539_;
  assign new_n541_ = pe0 & ~new_n234_;
  assign new_n542_ = pf0 & new_n541_;
  assign new_n543_ = pc0 & pe0;
  assign new_n544_ = ~new_n339_ & ~new_n543_;
  assign new_n545_ = ~pf0 & new_n544_;
  assign new_n546_ = ~new_n542_ & ~new_n545_;
  assign new_n547_ = new_n540_ & new_n546_;
  assign new_n548_ = new_n431_ & new_n547_;
  assign new_n549_ = pp & pl;
  assign new_n550_ = ~pq & new_n549_;
  assign new_n551_ = new_n546_ & new_n550_;
  assign new_n552_ = new_n431_ & new_n551_;
  assign new_n553_ = pr & ~ps;
  assign new_n554_ = pt & new_n553_;
  assign new_n555_ = po & new_n251_;
  assign new_n556_ = pp & new_n555_;
  assign new_n557_ = ~pf0 & new_n234_;
  assign new_n558_ = new_n556_ & ~new_n557_;
  assign new_n559_ = ~pt & new_n558_;
  assign new_n560_ = new_n234_ & new_n559_;
  assign new_n561_ = pf0 & new_n560_;
  assign new_n562_ = ~pf0 & new_n559_;
  assign new_n563_ = pe0 & new_n562_;
  assign new_n564_ = pe0 & new_n560_;
  assign new_n565_ = pf0 & new_n559_;
  assign new_n566_ = ~pe0 & new_n565_;
  assign new_n567_ = ~new_n564_ & ~new_n566_;
  assign new_n568_ = ~new_n561_ & ~new_n563_;
  assign new_n569_ = new_n567_ & new_n568_;
  assign new_n570_ = pp & pm;
  assign new_n571_ = pq & new_n570_;
  assign new_n572_ = ~new_n554_ & new_n569_;
  assign new_n573_ = ~new_n571_ & new_n572_;
  assign new_n574_ = ~pr & ps;
  assign new_n575_ = pt & new_n574_;
  assign new_n576_ = new_n572_ & ~new_n575_;
  assign new_n577_ = pp & pn;
  assign new_n578_ = pq & new_n577_;
  assign new_n579_ = new_n569_ & ~new_n578_;
  assign new_n580_ = ~new_n571_ & new_n579_;
  assign new_n581_ = ~new_n575_ & new_n579_;
  assign new_n582_ = ~pe0 & new_n521_;
  assign new_n583_ = new_n234_ & new_n521_;
  assign new_n584_ = ~pf0 & new_n521_;
  assign new_n585_ = ~new_n582_ & ~new_n583_;
  assign new_n586_ = ~new_n584_ & new_n585_;
  assign new_n587_ = new_n569_ & new_n586_;
  assign new_n588_ = ~new_n573_ & ~new_n576_;
  assign new_n589_ = ~new_n580_ & new_n588_;
  assign new_n590_ = ~new_n581_ & ~new_n587_;
  assign new_n591_ = new_n589_ & new_n590_;
  assign new_n592_ = ~new_n548_ & ~new_n552_;
  assign new_n593_ = ~new_n591_ & new_n592_;
  assign new_n594_ = new_n537_ & new_n593_;
  assign new_n595_ = ~ph0 & new_n593_;
  assign new_n596_ = ~pg0 & new_n537_;
  assign new_n597_ = ~pg0 & ~ph0;
  assign new_n598_ = ~new_n538_ & ~new_n594_;
  assign new_n599_ = ~new_n595_ & new_n598_;
  assign new_n600_ = ~new_n596_ & ~new_n597_;
  assign new_n601_ = new_n599_ & new_n600_;
  assign new_n602_ = pa & new_n601_;
  assign pr0 = ~pa0 & new_n602_;
  assign new_n604_ = ~pq & ~new_n431_;
  assign new_n605_ = ~pg0 & new_n541_;
  assign new_n606_ = ~pr & ~ps;
  assign new_n607_ = ~pk & new_n431_;
  assign new_n608_ = pq & new_n607_;
  assign new_n609_ = pd0 & new_n465_;
  assign new_n610_ = ~pf0 & ~pg0;
  assign new_n611_ = ~new_n466_ & ~new_n609_;
  assign new_n612_ = ~new_n610_ & new_n611_;
  assign new_n613_ = ~new_n606_ & ~new_n608_;
  assign new_n614_ = ~new_n612_ & new_n613_;
  assign new_n615_ = ps & new_n614_;
  assign new_n616_ = pr & new_n615_;
  assign new_n617_ = pt & new_n614_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = ~new_n604_ & ~new_n605_;
  assign new_n620_ = ~new_n618_ & new_n619_;
  assign new_n621_ = new_n505_ & new_n620_;
  assign new_n622_ = ~pp & new_n621_;
  assign new_n623_ = ~pt & po;
  assign new_n624_ = ~ps & pn;
  assign new_n625_ = ~ps & ~pt;
  assign new_n626_ = ~new_n623_ & ~new_n624_;
  assign new_n627_ = ~new_n625_ & new_n626_;
  assign new_n628_ = new_n495_ & new_n627_;
  assign new_n629_ = new_n492_ & new_n628_;
  assign new_n630_ = pr & new_n627_;
  assign new_n631_ = new_n492_ & new_n630_;
  assign new_n632_ = pq & new_n628_;
  assign new_n633_ = pq & new_n630_;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = ~new_n629_ & ~new_n631_;
  assign new_n636_ = new_n634_ & new_n635_;
  assign new_n637_ = new_n621_ & new_n636_;
  assign new_n638_ = new_n620_ & new_n636_;
  assign new_n639_ = pp & new_n638_;
  assign new_n640_ = ~new_n622_ & ~new_n637_;
  assign new_n641_ = ~new_n639_ & new_n640_;
  assign new_n642_ = pi0 & new_n641_;
  assign new_n643_ = pt & ~pi0;
  assign new_n644_ = pk & new_n643_;
  assign new_n645_ = ~pp & new_n644_;
  assign new_n646_ = ~pp & ~new_n642_;
  assign new_n647_ = ~new_n645_ & new_n646_;
  assign new_n648_ = ~new_n251_ & new_n646_;
  assign new_n649_ = pi0 & ~new_n642_;
  assign new_n650_ = ~new_n251_ & new_n649_;
  assign new_n651_ = ~pg0 & new_n545_;
  assign new_n652_ = pf0 & pg0;
  assign new_n653_ = ~new_n234_ & new_n652_;
  assign new_n654_ = pe0 & new_n653_;
  assign new_n655_ = ~new_n651_ & ~new_n654_;
  assign new_n656_ = new_n649_ & new_n655_;
  assign new_n657_ = ~new_n645_ & new_n649_;
  assign new_n658_ = ~new_n496_ & ~new_n500_;
  assign new_n659_ = pq & new_n658_;
  assign new_n660_ = pr & ~pl;
  assign new_n661_ = ps & new_n660_;
  assign new_n662_ = pt & new_n661_;
  assign new_n663_ = ~new_n514_ & ~new_n606_;
  assign new_n664_ = ~new_n662_ & new_n663_;
  assign new_n665_ = ps & new_n664_;
  assign new_n666_ = pc0 & new_n665_;
  assign new_n667_ = pt & new_n664_;
  assign new_n668_ = pc0 & new_n667_;
  assign new_n669_ = pd0 & new_n665_;
  assign new_n670_ = pd0 & new_n667_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~new_n666_ & ~new_n668_;
  assign new_n673_ = new_n671_ & new_n672_;
  assign new_n674_ = ~new_n604_ & ~new_n659_;
  assign new_n675_ = ~new_n673_ & new_n674_;
  assign new_n676_ = new_n652_ & new_n675_;
  assign new_n677_ = pe0 & new_n676_;
  assign new_n678_ = ~pm & new_n333_;
  assign new_n679_ = ~pr & ~pm;
  assign new_n680_ = ~new_n514_ & ~new_n679_;
  assign new_n681_ = ~new_n606_ & ~new_n678_;
  assign new_n682_ = new_n680_ & new_n681_;
  assign new_n683_ = ps & new_n682_;
  assign new_n684_ = ~pc0 & new_n683_;
  assign new_n685_ = pt & new_n682_;
  assign new_n686_ = ~pc0 & new_n685_;
  assign new_n687_ = ~pe0 & new_n683_;
  assign new_n688_ = ~pe0 & new_n685_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = ~new_n684_ & ~new_n686_;
  assign new_n691_ = new_n689_ & new_n690_;
  assign new_n692_ = ~new_n339_ & ~new_n630_;
  assign new_n693_ = ~new_n691_ & new_n692_;
  assign new_n694_ = new_n610_ & new_n693_;
  assign new_n695_ = pq & new_n694_;
  assign new_n696_ = pl & new_n431_;
  assign new_n697_ = ~pq & new_n696_;
  assign new_n698_ = ~pd0 & new_n697_;
  assign new_n699_ = ~pc0 & new_n698_;
  assign new_n700_ = ~pe0 & new_n697_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = ~pf0 & ~new_n701_;
  assign new_n703_ = ~pg0 & new_n702_;
  assign new_n704_ = ~new_n677_ & ~new_n695_;
  assign new_n705_ = ~new_n703_ & new_n704_;
  assign new_n706_ = ~new_n642_ & new_n705_;
  assign new_n707_ = ~new_n251_ & new_n706_;
  assign new_n708_ = new_n655_ & new_n706_;
  assign new_n709_ = new_n646_ & new_n655_;
  assign new_n710_ = ~new_n645_ & new_n706_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = ~new_n707_ & ~new_n708_;
  assign new_n713_ = new_n711_ & new_n712_;
  assign new_n714_ = ~new_n647_ & ~new_n648_;
  assign new_n715_ = ~new_n650_ & new_n714_;
  assign new_n716_ = ~new_n656_ & ~new_n657_;
  assign new_n717_ = new_n715_ & new_n716_;
  assign new_n718_ = new_n713_ & new_n717_;
  assign new_n719_ = pa & new_n718_;
  assign ps0 = ~pa0 & new_n719_;
  assign pj0 = ~ph0;
endmodule

