// Benchmark "testing" written by ABC on Thu Oct  8 22:16:59 2020

module testing ( 
    A7979, A7978, A7977, A7976, A7975, A7974, A7912, A7911, A7910, A7909,
    A7908, A7907, A7845, A7844, A7843, A7842, A7841, A7840, A7778, A7777,
    A7776, A7775, A7774, A7773, A7711, A7710, A7709, A7708, A7707, A7706,
    A7644, A7643, A7642, A7641, A7640, A7639, A7577, A7576, A7575, A7574,
    A7573, A7572, A7510, A7509, A7508, A7507, A7506, A7505, A7443, A7442,
    A7441, A7440, A7439, A7438, A7376, A7375, A7374, A7373, A7372, A7371,
    A7309, A7308, A7307, A7306, A7305, A7304, A7242, A7241, A7240, A7239,
    A7238, A7237, A7175, A7174, A7173, A7172, A7171, A7170, A7108, A7107,
    A7106, A7105, A7104, A7103, A7041, A7040, A7039, A7038, A7037, A7036,
    A6974, A6973, A6972, A6971, A6970, A6969, A6907, A6906, A6905, A6904,
    A6903, A6902, A6840, A6839, A6838, A6837, A6836, A6835, A6773, A6772,
    A6771, A6770, A6769, A6768, A6706, A6705, A6704, A6703, A6702, A6701,
    A6639, A6638, A6637, A6636, A6635, A6634, A6572, A6571, A6570, A6569,
    A6568, A6567, A6505, A6504, A6503, A6502, A6501, A6500, A6438, A6437,
    A6436, A6435, A6434, A6433, A6371, A6370, A6369, A6368, A6367, A6366,
    A6304, A6303, A6302, A6301, A6300, A6299, A6237, A6236, A6235, A6234,
    A6233, A6232, A6170, A6169, A6168, A6167, A6166, A6165, A6103, A6102,
    A6101, A6100, A6099, A6098, A6036, A6035, A6034, A6033, A6032, A6031,
    A5969, A5968, A5967, A5966, A5965, A5964, A5902, A5901, A5900, A5899,
    A5898, A5897, A5835, A5834, A5833, A5832, A5831, A5830, A5768, A5767,
    A5766, A5765, A5764, A5763, A5701, A5700, A5699, A5698, A5697, A5696,
    A5629, A5630, A5631, A5632, A5633, A5634,
    A3161, A3160, A3159, A3158, A3157, A3156, A3094, A3093, A3092, A3091,
    A3090, A3089, A3027, A3026, A3025, A3024, A3023, A3022, A2960, A2959,
    A2958, A2957, A2956, A2955, A2893, A2892, A2891, A2890, A2889, A2888,
    A2826, A2825, A2824, A2823, A2822, A2821, A2759, A2758, A2757, A2756,
    A2755, A2754, A2692, A2691, A2690, A2689, A2688, A2687, A2625, A2624,
    A2623, A2622, A2621, A2620, A2558, A2557, A2556, A2555, A2554, A2553,
    A2491, A2490, A2489, A2488, A2487, A2486, A2424, A2423, A2422, A2421,
    A2420, A2419, A2357, A2356, A2355, A2354, A2353, A2352, A2290, A2289,
    A2288, A2287, A2286, A2285, A2223, A2222, A2221, A2220, A2219, A2218,
    A2156, A2155, A2154, A2153, A2152, A2151, A2089, A2088, A2087, A2086,
    A2085, A2084, A2022, A2021, A2020, A2019, A2018, A2017, A1955, A1954,
    A1953, A1952, A1951, A1950, A1888, A1887, A1886, A1885, A1884, A1883,
    A1821, A1820, A1819, A1818, A1817, A1816, A1754, A1753, A1752, A1751,
    A1750, A1749, A1687, A1686, A1685, A1684, A1683, A1682, A1620, A1619,
    A1618, A1617, A1616, A1615, A1553, A1552, A1551, A1550, A1549, A1548,
    A1486, A1485, A1484, A1483, A1482, A1481, A1419, A1418, A1417, A1416,
    A1415, A1414, A1352, A1351, A1350, A1349, A1348, A1347, A1285, A1284,
    A1283, A1282, A1281, A1280, A1218, A1217, A1216, A1215, A1214, A1213,
    A1151, A1150, A1149, A1148, A1147, A1146, A1084, A1083, A1082, A1081,
    A1080, A1079, A1017, A1016, A1015, A1014, A1013, A1012, A950, A949,
    A948, A947, A946, A945, A883, A882, A881, A880, A879, A878, A811, A812,
    A813, A814, A815, A816  );
  input  A7979, A7978, A7977, A7976, A7975, A7974, A7912, A7911, A7910,
    A7909, A7908, A7907, A7845, A7844, A7843, A7842, A7841, A7840, A7778,
    A7777, A7776, A7775, A7774, A7773, A7711, A7710, A7709, A7708, A7707,
    A7706, A7644, A7643, A7642, A7641, A7640, A7639, A7577, A7576, A7575,
    A7574, A7573, A7572, A7510, A7509, A7508, A7507, A7506, A7505, A7443,
    A7442, A7441, A7440, A7439, A7438, A7376, A7375, A7374, A7373, A7372,
    A7371, A7309, A7308, A7307, A7306, A7305, A7304, A7242, A7241, A7240,
    A7239, A7238, A7237, A7175, A7174, A7173, A7172, A7171, A7170, A7108,
    A7107, A7106, A7105, A7104, A7103, A7041, A7040, A7039, A7038, A7037,
    A7036, A6974, A6973, A6972, A6971, A6970, A6969, A6907, A6906, A6905,
    A6904, A6903, A6902, A6840, A6839, A6838, A6837, A6836, A6835, A6773,
    A6772, A6771, A6770, A6769, A6768, A6706, A6705, A6704, A6703, A6702,
    A6701, A6639, A6638, A6637, A6636, A6635, A6634, A6572, A6571, A6570,
    A6569, A6568, A6567, A6505, A6504, A6503, A6502, A6501, A6500, A6438,
    A6437, A6436, A6435, A6434, A6433, A6371, A6370, A6369, A6368, A6367,
    A6366, A6304, A6303, A6302, A6301, A6300, A6299, A6237, A6236, A6235,
    A6234, A6233, A6232, A6170, A6169, A6168, A6167, A6166, A6165, A6103,
    A6102, A6101, A6100, A6099, A6098, A6036, A6035, A6034, A6033, A6032,
    A6031, A5969, A5968, A5967, A5966, A5965, A5964, A5902, A5901, A5900,
    A5899, A5898, A5897, A5835, A5834, A5833, A5832, A5831, A5830, A5768,
    A5767, A5766, A5765, A5764, A5763, A5701, A5700, A5699, A5698, A5697,
    A5696, A5629, A5630, A5631, A5632, A5633, A5634;
  output A3161, A3160, A3159, A3158, A3157, A3156, A3094, A3093, A3092, A3091,
    A3090, A3089, A3027, A3026, A3025, A3024, A3023, A3022, A2960, A2959,
    A2958, A2957, A2956, A2955, A2893, A2892, A2891, A2890, A2889, A2888,
    A2826, A2825, A2824, A2823, A2822, A2821, A2759, A2758, A2757, A2756,
    A2755, A2754, A2692, A2691, A2690, A2689, A2688, A2687, A2625, A2624,
    A2623, A2622, A2621, A2620, A2558, A2557, A2556, A2555, A2554, A2553,
    A2491, A2490, A2489, A2488, A2487, A2486, A2424, A2423, A2422, A2421,
    A2420, A2419, A2357, A2356, A2355, A2354, A2353, A2352, A2290, A2289,
    A2288, A2287, A2286, A2285, A2223, A2222, A2221, A2220, A2219, A2218,
    A2156, A2155, A2154, A2153, A2152, A2151, A2089, A2088, A2087, A2086,
    A2085, A2084, A2022, A2021, A2020, A2019, A2018, A2017, A1955, A1954,
    A1953, A1952, A1951, A1950, A1888, A1887, A1886, A1885, A1884, A1883,
    A1821, A1820, A1819, A1818, A1817, A1816, A1754, A1753, A1752, A1751,
    A1750, A1749, A1687, A1686, A1685, A1684, A1683, A1682, A1620, A1619,
    A1618, A1617, A1616, A1615, A1553, A1552, A1551, A1550, A1549, A1548,
    A1486, A1485, A1484, A1483, A1482, A1481, A1419, A1418, A1417, A1416,
    A1415, A1414, A1352, A1351, A1350, A1349, A1348, A1347, A1285, A1284,
    A1283, A1282, A1281, A1280, A1218, A1217, A1216, A1215, A1214, A1213,
    A1151, A1150, A1149, A1148, A1147, A1146, A1084, A1083, A1082, A1081,
    A1080, A1079, A1017, A1016, A1015, A1014, A1013, A1012, A950, A949,
    A948, A947, A946, A945, A883, A882, A881, A880, A879, A878, A811, A812,
    A813, A814, A815, A816;
  wire new_A5695_, new_A5694_, new_A5693_, new_A5692_, new_A5691_,
    new_A5690_, new_A5689_, new_A5688_, new_A5687_, new_A5686_, new_A5685_,
    new_A5684_, new_A5683_, new_A5682_, new_A5681_, new_A5680_, new_A5679_,
    new_A5678_, new_A5677_, new_A5676_, new_A5675_, new_A5674_, new_A5673_,
    new_A5672_, new_A5671_, new_A5670_, new_A5669_, new_A5668_, new_A5667_,
    new_A5666_, new_A5665_, new_A5664_, new_A5663_, new_A5662_, new_A5661_,
    new_A5660_, new_A5659_, new_A5658_, new_A5657_, new_A5656_, new_A5655_,
    new_A5654_, new_A5653_, new_A5652_, new_A5651_, new_A5650_, new_A5649_,
    new_A5648_, new_A5647_, new_A5646_, new_A5645_, new_A5644_, new_A5643_,
    new_A5642_, new_A5641_, new_A5640_, new_A5639_, new_A5638_, new_A5637_,
    new_A5636_, new_A5635_, new_A5702_, new_A5703_, new_A5704_, new_A5705_,
    new_A5706_, new_A5707_, new_A5708_, new_A5709_, new_A5710_, new_A5711_,
    new_A5712_, new_A5713_, new_A5714_, new_A5715_, new_A5716_, new_A5717_,
    new_A5718_, new_A5719_, new_A5720_, new_A5721_, new_A5722_, new_A5723_,
    new_A5724_, new_A5725_, new_A5726_, new_A5727_, new_A5728_, new_A5729_,
    new_A5730_, new_A5731_, new_A5732_, new_A5733_, new_A5734_, new_A5735_,
    new_A5736_, new_A5737_, new_A5738_, new_A5739_, new_A5740_, new_A5741_,
    new_A5742_, new_A5743_, new_A5744_, new_A5745_, new_A5746_, new_A5747_,
    new_A5748_, new_A5749_, new_A5750_, new_A5751_, new_A5752_, new_A5753_,
    new_A5754_, new_A5755_, new_A5756_, new_A5757_, new_A5758_, new_A5759_,
    new_A5760_, new_A5761_, new_A5762_, new_A5769_, new_A5770_, new_A5771_,
    new_A5772_, new_A5773_, new_A5774_, new_A5775_, new_A5776_, new_A5777_,
    new_A5778_, new_A5779_, new_A5780_, new_A5781_, new_A5782_, new_A5783_,
    new_A5784_, new_A5785_, new_A5786_, new_A5787_, new_A5788_, new_A5789_,
    new_A5790_, new_A5791_, new_A5792_, new_A5793_, new_A5794_, new_A5795_,
    new_A5796_, new_A5797_, new_A5798_, new_A5799_, new_A5800_, new_A5801_,
    new_A5802_, new_A5803_, new_A5804_, new_A5805_, new_A5806_, new_A5807_,
    new_A5808_, new_A5809_, new_A5810_, new_A5811_, new_A5812_, new_A5813_,
    new_A5814_, new_A5815_, new_A5816_, new_A5817_, new_A5818_, new_A5819_,
    new_A5820_, new_A5821_, new_A5822_, new_A5823_, new_A5824_, new_A5825_,
    new_A5826_, new_A5827_, new_A5828_, new_A5829_, new_A5836_, new_A5837_,
    new_A5838_, new_A5839_, new_A5840_, new_A5841_, new_A5842_, new_A5843_,
    new_A5844_, new_A5845_, new_A5846_, new_A5847_, new_A5848_, new_A5849_,
    new_A5850_, new_A5851_, new_A5852_, new_A5853_, new_A5854_, new_A5855_,
    new_A5856_, new_A5857_, new_A5858_, new_A5859_, new_A5860_, new_A5861_,
    new_A5862_, new_A5863_, new_A5864_, new_A5865_, new_A5866_, new_A5867_,
    new_A5868_, new_A5869_, new_A5870_, new_A5871_, new_A5872_, new_A5873_,
    new_A5874_, new_A5875_, new_A5876_, new_A5877_, new_A5878_, new_A5879_,
    new_A5880_, new_A5881_, new_A5882_, new_A5883_, new_A5884_, new_A5885_,
    new_A5886_, new_A5887_, new_A5888_, new_A5889_, new_A5890_, new_A5891_,
    new_A5892_, new_A5893_, new_A5894_, new_A5895_, new_A5896_, new_A5903_,
    new_A5904_, new_A5905_, new_A5906_, new_A5907_, new_A5908_, new_A5909_,
    new_A5910_, new_A5911_, new_A5912_, new_A5913_, new_A5914_, new_A5915_,
    new_A5916_, new_A5917_, new_A5918_, new_A5919_, new_A5920_, new_A5921_,
    new_A5922_, new_A5923_, new_A5924_, new_A5925_, new_A5926_, new_A5927_,
    new_A5928_, new_A5929_, new_A5930_, new_A5931_, new_A5932_, new_A5933_,
    new_A5934_, new_A5935_, new_A5936_, new_A5937_, new_A5938_, new_A5939_,
    new_A5940_, new_A5941_, new_A5942_, new_A5943_, new_A5944_, new_A5945_,
    new_A5946_, new_A5947_, new_A5948_, new_A5949_, new_A5950_, new_A5951_,
    new_A5952_, new_A5953_, new_A5954_, new_A5955_, new_A5956_, new_A5957_,
    new_A5958_, new_A5959_, new_A5960_, new_A5961_, new_A5962_, new_A5963_,
    new_A5970_, new_A5971_, new_A5972_, new_A5973_, new_A5974_, new_A5975_,
    new_A5976_, new_A5977_, new_A5978_, new_A5979_, new_A5980_, new_A5981_,
    new_A5982_, new_A5983_, new_A5984_, new_A5985_, new_A5986_, new_A5987_,
    new_A5988_, new_A5989_, new_A5990_, new_A5991_, new_A5992_, new_A5993_,
    new_A5994_, new_A5995_, new_A5996_, new_A5997_, new_A5998_, new_A5999_,
    new_A6000_, new_A6001_, new_A6002_, new_A6003_, new_A6004_, new_A6005_,
    new_A6006_, new_A6007_, new_A6008_, new_A6009_, new_A6010_, new_A6011_,
    new_A6012_, new_A6013_, new_A6014_, new_A6015_, new_A6016_, new_A6017_,
    new_A6018_, new_A6019_, new_A6020_, new_A6021_, new_A6022_, new_A6023_,
    new_A6024_, new_A6025_, new_A6026_, new_A6027_, new_A6028_, new_A6029_,
    new_A6030_, new_A6037_, new_A6038_, new_A6039_, new_A6040_, new_A6041_,
    new_A6042_, new_A6043_, new_A6044_, new_A6045_, new_A6046_, new_A6047_,
    new_A6048_, new_A6049_, new_A6050_, new_A6051_, new_A6052_, new_A6053_,
    new_A6054_, new_A6055_, new_A6056_, new_A6057_, new_A6058_, new_A6059_,
    new_A6060_, new_A6061_, new_A6062_, new_A6063_, new_A6064_, new_A6065_,
    new_A6066_, new_A6067_, new_A6068_, new_A6069_, new_A6070_, new_A6071_,
    new_A6072_, new_A6073_, new_A6074_, new_A6075_, new_A6076_, new_A6077_,
    new_A6078_, new_A6079_, new_A6080_, new_A6081_, new_A6082_, new_A6083_,
    new_A6084_, new_A6085_, new_A6086_, new_A6087_, new_A6088_, new_A6089_,
    new_A6090_, new_A6091_, new_A6092_, new_A6093_, new_A6094_, new_A6095_,
    new_A6096_, new_A6097_, new_A6104_, new_A6105_, new_A6106_, new_A6107_,
    new_A6108_, new_A6109_, new_A6110_, new_A6111_, new_A6112_, new_A6113_,
    new_A6114_, new_A6115_, new_A6116_, new_A6117_, new_A6118_, new_A6119_,
    new_A6120_, new_A6121_, new_A6122_, new_A6123_, new_A6124_, new_A6125_,
    new_A6126_, new_A6127_, new_A6128_, new_A6129_, new_A6130_, new_A6131_,
    new_A6132_, new_A6133_, new_A6134_, new_A6135_, new_A6136_, new_A6137_,
    new_A6138_, new_A6139_, new_A6140_, new_A6141_, new_A6142_, new_A6143_,
    new_A6144_, new_A6145_, new_A6146_, new_A6147_, new_A6148_, new_A6149_,
    new_A6150_, new_A6151_, new_A6152_, new_A6153_, new_A6154_, new_A6155_,
    new_A6156_, new_A6157_, new_A6158_, new_A6159_, new_A6160_, new_A6161_,
    new_A6162_, new_A6163_, new_A6164_, new_A6171_, new_A6172_, new_A6173_,
    new_A6174_, new_A6175_, new_A6176_, new_A6177_, new_A6178_, new_A6179_,
    new_A6180_, new_A6181_, new_A6182_, new_A6183_, new_A6184_, new_A6185_,
    new_A6186_, new_A6187_, new_A6188_, new_A6189_, new_A6190_, new_A6191_,
    new_A6192_, new_A6193_, new_A6194_, new_A6195_, new_A6196_, new_A6197_,
    new_A6198_, new_A6199_, new_A6200_, new_A6201_, new_A6202_, new_A6203_,
    new_A6204_, new_A6205_, new_A6206_, new_A6207_, new_A6208_, new_A6209_,
    new_A6210_, new_A6211_, new_A6212_, new_A6213_, new_A6214_, new_A6215_,
    new_A6216_, new_A6217_, new_A6218_, new_A6219_, new_A6220_, new_A6221_,
    new_A6222_, new_A6223_, new_A6224_, new_A6225_, new_A6226_, new_A6227_,
    new_A6228_, new_A6229_, new_A6230_, new_A6231_, new_A6238_, new_A6239_,
    new_A6240_, new_A6241_, new_A6242_, new_A6243_, new_A6244_, new_A6245_,
    new_A6246_, new_A6247_, new_A6248_, new_A6249_, new_A6250_, new_A6251_,
    new_A6252_, new_A6253_, new_A6254_, new_A6255_, new_A6256_, new_A6257_,
    new_A6258_, new_A6259_, new_A6260_, new_A6261_, new_A6262_, new_A6263_,
    new_A6264_, new_A6265_, new_A6266_, new_A6267_, new_A6268_, new_A6269_,
    new_A6270_, new_A6271_, new_A6272_, new_A6273_, new_A6274_, new_A6275_,
    new_A6276_, new_A6277_, new_A6278_, new_A6279_, new_A6280_, new_A6281_,
    new_A6282_, new_A6283_, new_A6284_, new_A6285_, new_A6286_, new_A6287_,
    new_A6288_, new_A6289_, new_A6290_, new_A6291_, new_A6292_, new_A6293_,
    new_A6294_, new_A6295_, new_A6296_, new_A6297_, new_A6298_, new_A6305_,
    new_A6306_, new_A6307_, new_A6308_, new_A6309_, new_A6310_, new_A6311_,
    new_A6312_, new_A6313_, new_A6314_, new_A6315_, new_A6316_, new_A6317_,
    new_A6318_, new_A6319_, new_A6320_, new_A6321_, new_A6322_, new_A6323_,
    new_A6324_, new_A6325_, new_A6326_, new_A6327_, new_A6328_, new_A6329_,
    new_A6330_, new_A6331_, new_A6332_, new_A6333_, new_A6334_, new_A6335_,
    new_A6336_, new_A6337_, new_A6338_, new_A6339_, new_A6340_, new_A6341_,
    new_A6342_, new_A6343_, new_A6344_, new_A6345_, new_A6346_, new_A6347_,
    new_A6348_, new_A6349_, new_A6350_, new_A6351_, new_A6352_, new_A6353_,
    new_A6354_, new_A6355_, new_A6356_, new_A6357_, new_A6358_, new_A6359_,
    new_A6360_, new_A6361_, new_A6362_, new_A6363_, new_A6364_, new_A6365_,
    new_A6372_, new_A6373_, new_A6374_, new_A6375_, new_A6376_, new_A6377_,
    new_A6378_, new_A6379_, new_A6380_, new_A6381_, new_A6382_, new_A6383_,
    new_A6384_, new_A6385_, new_A6386_, new_A6387_, new_A6388_, new_A6389_,
    new_A6390_, new_A6391_, new_A6392_, new_A6393_, new_A6394_, new_A6395_,
    new_A6396_, new_A6397_, new_A6398_, new_A6399_, new_A6400_, new_A6401_,
    new_A6402_, new_A6403_, new_A6404_, new_A6405_, new_A6406_, new_A6407_,
    new_A6408_, new_A6409_, new_A6410_, new_A6411_, new_A6412_, new_A6413_,
    new_A6414_, new_A6415_, new_A6416_, new_A6417_, new_A6418_, new_A6419_,
    new_A6420_, new_A6421_, new_A6422_, new_A6423_, new_A6424_, new_A6425_,
    new_A6426_, new_A6427_, new_A6428_, new_A6429_, new_A6430_, new_A6431_,
    new_A6432_, new_A6439_, new_A6440_, new_A6441_, new_A6442_, new_A6443_,
    new_A6444_, new_A6445_, new_A6446_, new_A6447_, new_A6448_, new_A6449_,
    new_A6450_, new_A6451_, new_A6452_, new_A6453_, new_A6454_, new_A6455_,
    new_A6456_, new_A6457_, new_A6458_, new_A6459_, new_A6460_, new_A6461_,
    new_A6462_, new_A6463_, new_A6464_, new_A6465_, new_A6466_, new_A6467_,
    new_A6468_, new_A6469_, new_A6470_, new_A6471_, new_A6472_, new_A6473_,
    new_A6474_, new_A6475_, new_A6476_, new_A6477_, new_A6478_, new_A6479_,
    new_A6480_, new_A6481_, new_A6482_, new_A6483_, new_A6484_, new_A6485_,
    new_A6486_, new_A6487_, new_A6488_, new_A6489_, new_A6490_, new_A6491_,
    new_A6492_, new_A6493_, new_A6494_, new_A6495_, new_A6496_, new_A6497_,
    new_A6498_, new_A6499_, new_A6506_, new_A6507_, new_A6508_, new_A6509_,
    new_A6510_, new_A6511_, new_A6512_, new_A6513_, new_A6514_, new_A6515_,
    new_A6516_, new_A6517_, new_A6518_, new_A6519_, new_A6520_, new_A6521_,
    new_A6522_, new_A6523_, new_A6524_, new_A6525_, new_A6526_, new_A6527_,
    new_A6528_, new_A6529_, new_A6530_, new_A6531_, new_A6532_, new_A6533_,
    new_A6534_, new_A6535_, new_A6536_, new_A6537_, new_A6538_, new_A6539_,
    new_A6540_, new_A6541_, new_A6542_, new_A6543_, new_A6544_, new_A6545_,
    new_A6546_, new_A6547_, new_A6548_, new_A6549_, new_A6550_, new_A6551_,
    new_A6552_, new_A6553_, new_A6554_, new_A6555_, new_A6556_, new_A6557_,
    new_A6558_, new_A6559_, new_A6560_, new_A6561_, new_A6562_, new_A6563_,
    new_A6564_, new_A6565_, new_A6566_, new_A6573_, new_A6574_, new_A6575_,
    new_A6576_, new_A6577_, new_A6578_, new_A6579_, new_A6580_, new_A6581_,
    new_A6582_, new_A6583_, new_A6584_, new_A6585_, new_A6586_, new_A6587_,
    new_A6588_, new_A6589_, new_A6590_, new_A6591_, new_A6592_, new_A6593_,
    new_A6594_, new_A6595_, new_A6596_, new_A6597_, new_A6598_, new_A6599_,
    new_A6600_, new_A6601_, new_A6602_, new_A6603_, new_A6604_, new_A6605_,
    new_A6606_, new_A6607_, new_A6608_, new_A6609_, new_A6610_, new_A6611_,
    new_A6612_, new_A6613_, new_A6614_, new_A6615_, new_A6616_, new_A6617_,
    new_A6618_, new_A6619_, new_A6620_, new_A6621_, new_A6622_, new_A6623_,
    new_A6624_, new_A6625_, new_A6626_, new_A6627_, new_A6628_, new_A6629_,
    new_A6630_, new_A6631_, new_A6632_, new_A6633_, new_A6640_, new_A6641_,
    new_A6642_, new_A6643_, new_A6644_, new_A6645_, new_A6646_, new_A6647_,
    new_A6648_, new_A6649_, new_A6650_, new_A6651_, new_A6652_, new_A6653_,
    new_A6654_, new_A6655_, new_A6656_, new_A6657_, new_A6658_, new_A6659_,
    new_A6660_, new_A6661_, new_A6662_, new_A6663_, new_A6664_, new_A6665_,
    new_A6666_, new_A6667_, new_A6668_, new_A6669_, new_A6670_, new_A6671_,
    new_A6672_, new_A6673_, new_A6674_, new_A6675_, new_A6676_, new_A6677_,
    new_A6678_, new_A6679_, new_A6680_, new_A6681_, new_A6682_, new_A6683_,
    new_A6684_, new_A6685_, new_A6686_, new_A6687_, new_A6688_, new_A6689_,
    new_A6690_, new_A6691_, new_A6692_, new_A6693_, new_A6694_, new_A6695_,
    new_A6696_, new_A6697_, new_A6698_, new_A6699_, new_A6700_, new_A6707_,
    new_A6708_, new_A6709_, new_A6710_, new_A6711_, new_A6712_, new_A6713_,
    new_A6714_, new_A6715_, new_A6716_, new_A6717_, new_A6718_, new_A6719_,
    new_A6720_, new_A6721_, new_A6722_, new_A6723_, new_A6724_, new_A6725_,
    new_A6726_, new_A6727_, new_A6728_, new_A6729_, new_A6730_, new_A6731_,
    new_A6732_, new_A6733_, new_A6734_, new_A6735_, new_A6736_, new_A6737_,
    new_A6738_, new_A6739_, new_A6740_, new_A6741_, new_A6742_, new_A6743_,
    new_A6744_, new_A6745_, new_A6746_, new_A6747_, new_A6748_, new_A6749_,
    new_A6750_, new_A6751_, new_A6752_, new_A6753_, new_A6754_, new_A6755_,
    new_A6756_, new_A6757_, new_A6758_, new_A6759_, new_A6760_, new_A6761_,
    new_A6762_, new_A6763_, new_A6764_, new_A6765_, new_A6766_, new_A6767_,
    new_A6774_, new_A6775_, new_A6776_, new_A6777_, new_A6778_, new_A6779_,
    new_A6780_, new_A6781_, new_A6782_, new_A6783_, new_A6784_, new_A6785_,
    new_A6786_, new_A6787_, new_A6788_, new_A6789_, new_A6790_, new_A6791_,
    new_A6792_, new_A6793_, new_A6794_, new_A6795_, new_A6796_, new_A6797_,
    new_A6798_, new_A6799_, new_A6800_, new_A6801_, new_A6802_, new_A6803_,
    new_A6804_, new_A6805_, new_A6806_, new_A6807_, new_A6808_, new_A6809_,
    new_A6810_, new_A6811_, new_A6812_, new_A6813_, new_A6814_, new_A6815_,
    new_A6816_, new_A6817_, new_A6818_, new_A6819_, new_A6820_, new_A6821_,
    new_A6822_, new_A6823_, new_A6824_, new_A6825_, new_A6826_, new_A6827_,
    new_A6828_, new_A6829_, new_A6830_, new_A6831_, new_A6832_, new_A6833_,
    new_A6834_, new_A6841_, new_A6842_, new_A6843_, new_A6844_, new_A6845_,
    new_A6846_, new_A6847_, new_A6848_, new_A6849_, new_A6850_, new_A6851_,
    new_A6852_, new_A6853_, new_A6854_, new_A6855_, new_A6856_, new_A6857_,
    new_A6858_, new_A6859_, new_A6860_, new_A6861_, new_A6862_, new_A6863_,
    new_A6864_, new_A6865_, new_A6866_, new_A6867_, new_A6868_, new_A6869_,
    new_A6870_, new_A6871_, new_A6872_, new_A6873_, new_A6874_, new_A6875_,
    new_A6876_, new_A6877_, new_A6878_, new_A6879_, new_A6880_, new_A6881_,
    new_A6882_, new_A6883_, new_A6884_, new_A6885_, new_A6886_, new_A6887_,
    new_A6888_, new_A6889_, new_A6890_, new_A6891_, new_A6892_, new_A6893_,
    new_A6894_, new_A6895_, new_A6896_, new_A6897_, new_A6898_, new_A6899_,
    new_A6900_, new_A6901_, new_A6908_, new_A6909_, new_A6910_, new_A6911_,
    new_A6912_, new_A6913_, new_A6914_, new_A6915_, new_A6916_, new_A6917_,
    new_A6918_, new_A6919_, new_A6920_, new_A6921_, new_A6922_, new_A6923_,
    new_A6924_, new_A6925_, new_A6926_, new_A6927_, new_A6928_, new_A6929_,
    new_A6930_, new_A6931_, new_A6932_, new_A6933_, new_A6934_, new_A6935_,
    new_A6936_, new_A6937_, new_A6938_, new_A6939_, new_A6940_, new_A6941_,
    new_A6942_, new_A6943_, new_A6944_, new_A6945_, new_A6946_, new_A6947_,
    new_A6948_, new_A6949_, new_A6950_, new_A6951_, new_A6952_, new_A6953_,
    new_A6954_, new_A6955_, new_A6956_, new_A6957_, new_A6958_, new_A6959_,
    new_A6960_, new_A6961_, new_A6962_, new_A6963_, new_A6964_, new_A6965_,
    new_A6966_, new_A6967_, new_A6968_, new_A6975_, new_A6976_, new_A6977_,
    new_A6978_, new_A6979_, new_A6980_, new_A6981_, new_A6982_, new_A6983_,
    new_A6984_, new_A6985_, new_A6986_, new_A6987_, new_A6988_, new_A6989_,
    new_A6990_, new_A6991_, new_A6992_, new_A6993_, new_A6994_, new_A6995_,
    new_A6996_, new_A6997_, new_A6998_, new_A6999_, new_A7000_, new_A7001_,
    new_A7002_, new_A7003_, new_A7004_, new_A7005_, new_A7006_, new_A7007_,
    new_A7008_, new_A7009_, new_A7010_, new_A7011_, new_A7012_, new_A7013_,
    new_A7014_, new_A7015_, new_A7016_, new_A7017_, new_A7018_, new_A7019_,
    new_A7020_, new_A7021_, new_A7022_, new_A7023_, new_A7024_, new_A7025_,
    new_A7026_, new_A7027_, new_A7028_, new_A7029_, new_A7030_, new_A7031_,
    new_A7032_, new_A7033_, new_A7034_, new_A7035_, new_A7042_, new_A7043_,
    new_A7044_, new_A7045_, new_A7046_, new_A7047_, new_A7048_, new_A7049_,
    new_A7050_, new_A7051_, new_A7052_, new_A7053_, new_A7054_, new_A7055_,
    new_A7056_, new_A7057_, new_A7058_, new_A7059_, new_A7060_, new_A7061_,
    new_A7062_, new_A7063_, new_A7064_, new_A7065_, new_A7066_, new_A7067_,
    new_A7068_, new_A7069_, new_A7070_, new_A7071_, new_A7072_, new_A7073_,
    new_A7074_, new_A7075_, new_A7076_, new_A7077_, new_A7078_, new_A7079_,
    new_A7080_, new_A7081_, new_A7082_, new_A7083_, new_A7084_, new_A7085_,
    new_A7086_, new_A7087_, new_A7088_, new_A7089_, new_A7090_, new_A7091_,
    new_A7092_, new_A7093_, new_A7094_, new_A7095_, new_A7096_, new_A7097_,
    new_A7098_, new_A7099_, new_A7100_, new_A7101_, new_A7102_, new_A7109_,
    new_A7110_, new_A7111_, new_A7112_, new_A7113_, new_A7114_, new_A7115_,
    new_A7116_, new_A7117_, new_A7118_, new_A7119_, new_A7120_, new_A7121_,
    new_A7122_, new_A7123_, new_A7124_, new_A7125_, new_A7126_, new_A7127_,
    new_A7128_, new_A7129_, new_A7130_, new_A7131_, new_A7132_, new_A7133_,
    new_A7134_, new_A7135_, new_A7136_, new_A7137_, new_A7138_, new_A7139_,
    new_A7140_, new_A7141_, new_A7142_, new_A7143_, new_A7144_, new_A7145_,
    new_A7146_, new_A7147_, new_A7148_, new_A7149_, new_A7150_, new_A7151_,
    new_A7152_, new_A7153_, new_A7154_, new_A7155_, new_A7156_, new_A7157_,
    new_A7158_, new_A7159_, new_A7160_, new_A7161_, new_A7162_, new_A7163_,
    new_A7164_, new_A7165_, new_A7166_, new_A7167_, new_A7168_, new_A7169_,
    new_A7176_, new_A7177_, new_A7178_, new_A7179_, new_A7180_, new_A7181_,
    new_A7182_, new_A7183_, new_A7184_, new_A7185_, new_A7186_, new_A7187_,
    new_A7188_, new_A7189_, new_A7190_, new_A7191_, new_A7192_, new_A7193_,
    new_A7194_, new_A7195_, new_A7196_, new_A7197_, new_A7198_, new_A7199_,
    new_A7200_, new_A7201_, new_A7202_, new_A7203_, new_A7204_, new_A7205_,
    new_A7206_, new_A7207_, new_A7208_, new_A7209_, new_A7210_, new_A7211_,
    new_A7212_, new_A7213_, new_A7214_, new_A7215_, new_A7216_, new_A7217_,
    new_A7218_, new_A7219_, new_A7220_, new_A7221_, new_A7222_, new_A7223_,
    new_A7224_, new_A7225_, new_A7226_, new_A7227_, new_A7228_, new_A7229_,
    new_A7230_, new_A7231_, new_A7232_, new_A7233_, new_A7234_, new_A7235_,
    new_A7236_, new_A7243_, new_A7244_, new_A7245_, new_A7246_, new_A7247_,
    new_A7248_, new_A7249_, new_A7250_, new_A7251_, new_A7252_, new_A7253_,
    new_A7254_, new_A7255_, new_A7256_, new_A7257_, new_A7258_, new_A7259_,
    new_A7260_, new_A7261_, new_A7262_, new_A7263_, new_A7264_, new_A7265_,
    new_A7266_, new_A7267_, new_A7268_, new_A7269_, new_A7270_, new_A7271_,
    new_A7272_, new_A7273_, new_A7274_, new_A7275_, new_A7276_, new_A7277_,
    new_A7278_, new_A7279_, new_A7280_, new_A7281_, new_A7282_, new_A7283_,
    new_A7284_, new_A7285_, new_A7286_, new_A7287_, new_A7288_, new_A7289_,
    new_A7290_, new_A7291_, new_A7292_, new_A7293_, new_A7294_, new_A7295_,
    new_A7296_, new_A7297_, new_A7298_, new_A7299_, new_A7300_, new_A7301_,
    new_A7302_, new_A7303_, new_A7310_, new_A7311_, new_A7312_, new_A7313_,
    new_A7314_, new_A7315_, new_A7316_, new_A7317_, new_A7318_, new_A7319_,
    new_A7320_, new_A7321_, new_A7322_, new_A7323_, new_A7324_, new_A7325_,
    new_A7326_, new_A7327_, new_A7328_, new_A7329_, new_A7330_, new_A7331_,
    new_A7332_, new_A7333_, new_A7334_, new_A7335_, new_A7336_, new_A7337_,
    new_A7338_, new_A7339_, new_A7340_, new_A7341_, new_A7342_, new_A7343_,
    new_A7344_, new_A7345_, new_A7346_, new_A7347_, new_A7348_, new_A7349_,
    new_A7350_, new_A7351_, new_A7352_, new_A7353_, new_A7354_, new_A7355_,
    new_A7356_, new_A7357_, new_A7358_, new_A7359_, new_A7360_, new_A7361_,
    new_A7362_, new_A7363_, new_A7364_, new_A7365_, new_A7366_, new_A7367_,
    new_A7368_, new_A7369_, new_A7370_, new_A7377_, new_A7378_, new_A7379_,
    new_A7380_, new_A7381_, new_A7382_, new_A7383_, new_A7384_, new_A7385_,
    new_A7386_, new_A7387_, new_A7388_, new_A7389_, new_A7390_, new_A7391_,
    new_A7392_, new_A7393_, new_A7394_, new_A7395_, new_A7396_, new_A7397_,
    new_A7398_, new_A7399_, new_A7400_, new_A7401_, new_A7402_, new_A7403_,
    new_A7404_, new_A7405_, new_A7406_, new_A7407_, new_A7408_, new_A7409_,
    new_A7410_, new_A7411_, new_A7412_, new_A7413_, new_A7414_, new_A7415_,
    new_A7416_, new_A7417_, new_A7418_, new_A7419_, new_A7420_, new_A7421_,
    new_A7422_, new_A7423_, new_A7424_, new_A7425_, new_A7426_, new_A7427_,
    new_A7428_, new_A7429_, new_A7430_, new_A7431_, new_A7432_, new_A7433_,
    new_A7434_, new_A7435_, new_A7436_, new_A7437_, new_A7444_, new_A7445_,
    new_A7446_, new_A7447_, new_A7448_, new_A7449_, new_A7450_, new_A7451_,
    new_A7452_, new_A7453_, new_A7454_, new_A7455_, new_A7456_, new_A7457_,
    new_A7458_, new_A7459_, new_A7460_, new_A7461_, new_A7462_, new_A7463_,
    new_A7464_, new_A7465_, new_A7466_, new_A7467_, new_A7468_, new_A7469_,
    new_A7470_, new_A7471_, new_A7472_, new_A7473_, new_A7474_, new_A7475_,
    new_A7476_, new_A7477_, new_A7478_, new_A7479_, new_A7480_, new_A7481_,
    new_A7482_, new_A7483_, new_A7484_, new_A7485_, new_A7486_, new_A7487_,
    new_A7488_, new_A7489_, new_A7490_, new_A7491_, new_A7492_, new_A7493_,
    new_A7494_, new_A7495_, new_A7496_, new_A7497_, new_A7498_, new_A7499_,
    new_A7500_, new_A7501_, new_A7502_, new_A7503_, new_A7504_, new_A7511_,
    new_A7512_, new_A7513_, new_A7514_, new_A7515_, new_A7516_, new_A7517_,
    new_A7518_, new_A7519_, new_A7520_, new_A7521_, new_A7522_, new_A7523_,
    new_A7524_, new_A7525_, new_A7526_, new_A7527_, new_A7528_, new_A7529_,
    new_A7530_, new_A7531_, new_A7532_, new_A7533_, new_A7534_, new_A7535_,
    new_A7536_, new_A7537_, new_A7538_, new_A7539_, new_A7540_, new_A7541_,
    new_A7542_, new_A7543_, new_A7544_, new_A7545_, new_A7546_, new_A7547_,
    new_A7548_, new_A7549_, new_A7550_, new_A7551_, new_A7552_, new_A7553_,
    new_A7554_, new_A7555_, new_A7556_, new_A7557_, new_A7558_, new_A7559_,
    new_A7560_, new_A7561_, new_A7562_, new_A7563_, new_A7564_, new_A7565_,
    new_A7566_, new_A7567_, new_A7568_, new_A7569_, new_A7570_, new_A7571_,
    new_A7578_, new_A7579_, new_A7580_, new_A7581_, new_A7582_, new_A7583_,
    new_A7584_, new_A7585_, new_A7586_, new_A7587_, new_A7588_, new_A7589_,
    new_A7590_, new_A7591_, new_A7592_, new_A7593_, new_A7594_, new_A7595_,
    new_A7596_, new_A7597_, new_A7598_, new_A7599_, new_A7600_, new_A7601_,
    new_A7602_, new_A7603_, new_A7604_, new_A7605_, new_A7606_, new_A7607_,
    new_A7608_, new_A7609_, new_A7610_, new_A7611_, new_A7612_, new_A7613_,
    new_A7614_, new_A7615_, new_A7616_, new_A7617_, new_A7618_, new_A7619_,
    new_A7620_, new_A7621_, new_A7622_, new_A7623_, new_A7624_, new_A7625_,
    new_A7626_, new_A7627_, new_A7628_, new_A7629_, new_A7630_, new_A7631_,
    new_A7632_, new_A7633_, new_A7634_, new_A7635_, new_A7636_, new_A7637_,
    new_A7638_, new_A7645_, new_A7646_, new_A7647_, new_A7648_, new_A7649_,
    new_A7650_, new_A7651_, new_A7652_, new_A7653_, new_A7654_, new_A7655_,
    new_A7656_, new_A7657_, new_A7658_, new_A7659_, new_A7660_, new_A7661_,
    new_A7662_, new_A7663_, new_A7664_, new_A7665_, new_A7666_, new_A7667_,
    new_A7668_, new_A7669_, new_A7670_, new_A7671_, new_A7672_, new_A7673_,
    new_A7674_, new_A7675_, new_A7676_, new_A7677_, new_A7678_, new_A7679_,
    new_A7680_, new_A7681_, new_A7682_, new_A7683_, new_A7684_, new_A7685_,
    new_A7686_, new_A7687_, new_A7688_, new_A7689_, new_A7690_, new_A7691_,
    new_A7692_, new_A7693_, new_A7694_, new_A7695_, new_A7696_, new_A7697_,
    new_A7698_, new_A7699_, new_A7700_, new_A7701_, new_A7702_, new_A7703_,
    new_A7704_, new_A7705_, new_A7712_, new_A7713_, new_A7714_, new_A7715_,
    new_A7716_, new_A7717_, new_A7718_, new_A7719_, new_A7720_, new_A7721_,
    new_A7722_, new_A7723_, new_A7724_, new_A7725_, new_A7726_, new_A7727_,
    new_A7728_, new_A7729_, new_A7730_, new_A7731_, new_A7732_, new_A7733_,
    new_A7734_, new_A7735_, new_A7736_, new_A7737_, new_A7738_, new_A7739_,
    new_A7740_, new_A7741_, new_A7742_, new_A7743_, new_A7744_, new_A7745_,
    new_A7746_, new_A7747_, new_A7748_, new_A7749_, new_A7750_, new_A7751_,
    new_A7752_, new_A7753_, new_A7754_, new_A7755_, new_A7756_, new_A7757_,
    new_A7758_, new_A7759_, new_A7760_, new_A7761_, new_A7762_, new_A7763_,
    new_A7764_, new_A7765_, new_A7766_, new_A7767_, new_A7768_, new_A7769_,
    new_A7770_, new_A7771_, new_A7772_, new_A7779_, new_A7780_, new_A7781_,
    new_A7782_, new_A7783_, new_A7784_, new_A7785_, new_A7786_, new_A7787_,
    new_A7788_, new_A7789_, new_A7790_, new_A7791_, new_A7792_, new_A7793_,
    new_A7794_, new_A7795_, new_A7796_, new_A7797_, new_A7798_, new_A7799_,
    new_A7800_, new_A7801_, new_A7802_, new_A7803_, new_A7804_, new_A7805_,
    new_A7806_, new_A7807_, new_A7808_, new_A7809_, new_A7810_, new_A7811_,
    new_A7812_, new_A7813_, new_A7814_, new_A7815_, new_A7816_, new_A7817_,
    new_A7818_, new_A7819_, new_A7820_, new_A7821_, new_A7822_, new_A7823_,
    new_A7824_, new_A7825_, new_A7826_, new_A7827_, new_A7828_, new_A7829_,
    new_A7830_, new_A7831_, new_A7832_, new_A7833_, new_A7834_, new_A7835_,
    new_A7836_, new_A7837_, new_A7838_, new_A7839_, new_A7846_, new_A7847_,
    new_A7848_, new_A7849_, new_A7850_, new_A7851_, new_A7852_, new_A7853_,
    new_A7854_, new_A7855_, new_A7856_, new_A7857_, new_A7858_, new_A7859_,
    new_A7860_, new_A7861_, new_A7862_, new_A7863_, new_A7864_, new_A7865_,
    new_A7866_, new_A7867_, new_A7868_, new_A7869_, new_A7870_, new_A7871_,
    new_A7872_, new_A7873_, new_A7874_, new_A7875_, new_A7876_, new_A7877_,
    new_A7878_, new_A7879_, new_A7880_, new_A7881_, new_A7882_, new_A7883_,
    new_A7884_, new_A7885_, new_A7886_, new_A7887_, new_A7888_, new_A7889_,
    new_A7890_, new_A7891_, new_A7892_, new_A7893_, new_A7894_, new_A7895_,
    new_A7896_, new_A7897_, new_A7898_, new_A7899_, new_A7900_, new_A7901_,
    new_A7902_, new_A7903_, new_A7904_, new_A7905_, new_A7906_, new_A7913_,
    new_A7914_, new_A7915_, new_A7916_, new_A7917_, new_A7918_, new_A7919_,
    new_A7920_, new_A7921_, new_A7922_, new_A7923_, new_A7924_, new_A7925_,
    new_A7926_, new_A7927_, new_A7928_, new_A7929_, new_A7930_, new_A7931_,
    new_A7932_, new_A7933_, new_A7934_, new_A7935_, new_A7936_, new_A7937_,
    new_A7938_, new_A7939_, new_A7940_, new_A7941_, new_A7942_, new_A7943_,
    new_A7944_, new_A7945_, new_A7946_, new_A7947_, new_A7948_, new_A7949_,
    new_A7950_, new_A7951_, new_A7952_, new_A7953_, new_A7954_, new_A7955_,
    new_A7956_, new_A7957_, new_A7958_, new_A7959_, new_A7960_, new_A7961_,
    new_A7962_, new_A7963_, new_A7964_, new_A7965_, new_A7966_, new_A7967_,
    new_A7968_, new_A7969_, new_A7970_, new_A7971_, new_A7972_, new_A7973_,
    new_A7980_, new_A7981_, new_A7982_, new_A7983_, new_A7984_, new_A7985_,
    new_A7986_, new_A7987_, new_A7988_, new_A7989_, new_A7990_, new_A7991_,
    new_A7992_, new_A7993_, new_A7994_, new_A7995_, new_A7996_, new_A7997_,
    new_A7998_, new_A7999_, new_A8000_, new_A8001_, new_A8002_, new_A8003_,
    new_A8004_, new_A8005_, new_A8006_, new_A8007_, new_A8008_, new_A8009_,
    new_A8010_, new_A8011_, new_A8012_, new_A8013_, new_A8014_, new_A8015_,
    new_A8016_, new_A8017_, new_A8018_, new_A8019_, new_A8020_, new_A8021_,
    new_A8022_, new_A8023_, new_A8024_, new_A8025_, new_A8026_, new_A8027_,
    new_A8028_, new_A8029_, new_A8030_, new_A8031_, new_A8032_, new_A8033_,
    new_A8034_, new_A8035_, new_A8036_, new_A8037_, new_A8038_, new_A8039_,
    new_A8040_, new_A3283_, new_A3282_, new_A3281_, new_A3280_, new_A3279_,
    new_A3278_, new_A3277_, new_A3276_, new_A3275_, new_A3274_, new_A3273_,
    new_A3272_, new_A3271_, new_A3270_, new_A3269_, new_A3268_, new_A3267_,
    new_A3266_, new_A3265_, new_A3264_, new_A3263_, new_A3262_, new_A3261_,
    new_A3260_, new_A3259_, new_A3258_, new_A3257_, new_A3256_, new_A3255_,
    new_A3254_, new_A3253_, new_A3252_, new_A3251_, new_A3250_, new_A3249_,
    new_A3248_, new_A3247_, new_A3246_, new_A3245_, new_A3244_, new_A3243_,
    new_A3242_, new_A3241_, new_A3240_, new_A3239_, new_A3238_, new_A3237_,
    new_A3236_, new_A3235_, new_A3234_, new_A3233_, new_A3232_, new_A3231_,
    new_A3230_, new_A3229_, new_A3228_, new_A3227_, new_A3226_, new_A3225_,
    new_A3224_, new_A3223_, new_A3222_, new_A3221_, new_A3220_, new_A3219_,
    new_A3218_, new_A3217_, new_A3284_, new_A3285_, new_A3286_, new_A3287_,
    new_A3288_, new_A3289_, new_A3290_, new_A3291_, new_A3292_, new_A3293_,
    new_A3294_, new_A3295_, new_A3296_, new_A3297_, new_A3298_, new_A3299_,
    new_A3300_, new_A3301_, new_A3302_, new_A3303_, new_A3304_, new_A3305_,
    new_A3306_, new_A3307_, new_A3308_, new_A3309_, new_A3310_, new_A3311_,
    new_A3312_, new_A3313_, new_A3314_, new_A3315_, new_A3316_, new_A3317_,
    new_A3318_, new_A3319_, new_A3320_, new_A3321_, new_A3322_, new_A3323_,
    new_A3324_, new_A3325_, new_A3326_, new_A3327_, new_A3328_, new_A3329_,
    new_A3330_, new_A3331_, new_A3332_, new_A3333_, new_A3334_, new_A3335_,
    new_A3336_, new_A3337_, new_A3338_, new_A3339_, new_A3340_, new_A3341_,
    new_A3342_, new_A3343_, new_A3344_, new_A3345_, new_A3346_, new_A3347_,
    new_A3348_, new_A3349_, new_A3350_, new_A3351_, new_A3352_, new_A3353_,
    new_A3354_, new_A3355_, new_A3356_, new_A3357_, new_A3358_, new_A3359_,
    new_A3360_, new_A3361_, new_A3362_, new_A3363_, new_A3364_, new_A3365_,
    new_A3366_, new_A3367_, new_A3368_, new_A3369_, new_A3370_, new_A3371_,
    new_A3372_, new_A3373_, new_A3374_, new_A3375_, new_A3376_, new_A3377_,
    new_A3378_, new_A3379_, new_A3380_, new_A3381_, new_A3382_, new_A3383_,
    new_A3384_, new_A3385_, new_A3386_, new_A3387_, new_A3388_, new_A3389_,
    new_A3390_, new_A3391_, new_A3392_, new_A3393_, new_A3394_, new_A3395_,
    new_A3396_, new_A3397_, new_A3398_, new_A3399_, new_A3400_, new_A3401_,
    new_A3402_, new_A3403_, new_A3404_, new_A3405_, new_A3406_, new_A3407_,
    new_A3408_, new_A3409_, new_A3410_, new_A3411_, new_A3412_, new_A3413_,
    new_A3414_, new_A3415_, new_A3416_, new_A3417_, new_A3418_, new_A3419_,
    new_A3420_, new_A3421_, new_A3422_, new_A3423_, new_A3424_, new_A3425_,
    new_A3426_, new_A3427_, new_A3428_, new_A3429_, new_A3430_, new_A3431_,
    new_A3432_, new_A3433_, new_A3434_, new_A3435_, new_A3436_, new_A3437_,
    new_A3438_, new_A3439_, new_A3440_, new_A3441_, new_A3442_, new_A3443_,
    new_A3444_, new_A3445_, new_A3446_, new_A3447_, new_A3448_, new_A3449_,
    new_A3450_, new_A3451_, new_A3452_, new_A3453_, new_A3454_, new_A3455_,
    new_A3456_, new_A3457_, new_A3458_, new_A3459_, new_A3460_, new_A3461_,
    new_A3462_, new_A3463_, new_A3464_, new_A3465_, new_A3466_, new_A3467_,
    new_A3468_, new_A3469_, new_A3470_, new_A3471_, new_A3472_, new_A3473_,
    new_A3474_, new_A3475_, new_A3476_, new_A3477_, new_A3478_, new_A3479_,
    new_A3480_, new_A3481_, new_A3482_, new_A3483_, new_A3484_, new_A3485_,
    new_A3486_, new_A3487_, new_A3488_, new_A3489_, new_A3490_, new_A3491_,
    new_A3492_, new_A3493_, new_A3494_, new_A3495_, new_A3496_, new_A3497_,
    new_A3498_, new_A3499_, new_A3500_, new_A3501_, new_A3502_, new_A3503_,
    new_A3504_, new_A3505_, new_A3506_, new_A3507_, new_A3508_, new_A3509_,
    new_A3510_, new_A3511_, new_A3512_, new_A3513_, new_A3514_, new_A3515_,
    new_A3516_, new_A3517_, new_A3518_, new_A3519_, new_A3520_, new_A3521_,
    new_A3522_, new_A3523_, new_A3524_, new_A3525_, new_A3526_, new_A3527_,
    new_A3528_, new_A3529_, new_A3530_, new_A3531_, new_A3532_, new_A3533_,
    new_A3534_, new_A3535_, new_A3536_, new_A3537_, new_A3538_, new_A3539_,
    new_A3540_, new_A3541_, new_A3542_, new_A3543_, new_A3544_, new_A3545_,
    new_A3546_, new_A3547_, new_A3548_, new_A3549_, new_A3550_, new_A3551_,
    new_A3552_, new_A3553_, new_A3554_, new_A3555_, new_A3556_, new_A3557_,
    new_A3558_, new_A3559_, new_A3560_, new_A3561_, new_A3562_, new_A3563_,
    new_A3564_, new_A3565_, new_A3566_, new_A3567_, new_A3568_, new_A3569_,
    new_A3570_, new_A3571_, new_A3572_, new_A3573_, new_A3574_, new_A3575_,
    new_A3576_, new_A3577_, new_A3578_, new_A3579_, new_A3580_, new_A3581_,
    new_A3582_, new_A3583_, new_A3584_, new_A3585_, new_A3586_, new_A3587_,
    new_A3588_, new_A3589_, new_A3590_, new_A3591_, new_A3592_, new_A3593_,
    new_A3594_, new_A3595_, new_A3596_, new_A3597_, new_A3598_, new_A3599_,
    new_A3600_, new_A3601_, new_A3602_, new_A3603_, new_A3604_, new_A3605_,
    new_A3606_, new_A3607_, new_A3608_, new_A3609_, new_A3610_, new_A3611_,
    new_A3612_, new_A3613_, new_A3614_, new_A3615_, new_A3616_, new_A3617_,
    new_A3618_, new_A3619_, new_A3620_, new_A3621_, new_A3622_, new_A3623_,
    new_A3624_, new_A3625_, new_A3626_, new_A3627_, new_A3628_, new_A3629_,
    new_A3630_, new_A3631_, new_A3632_, new_A3633_, new_A3634_, new_A3635_,
    new_A3636_, new_A3637_, new_A3638_, new_A3639_, new_A3640_, new_A3641_,
    new_A3642_, new_A3643_, new_A3644_, new_A3645_, new_A3646_, new_A3647_,
    new_A3648_, new_A3649_, new_A3650_, new_A3651_, new_A3652_, new_A3653_,
    new_A3654_, new_A3655_, new_A3656_, new_A3657_, new_A3658_, new_A3659_,
    new_A3660_, new_A3661_, new_A3662_, new_A3663_, new_A3664_, new_A3665_,
    new_A3666_, new_A3667_, new_A3668_, new_A3669_, new_A3670_, new_A3671_,
    new_A3672_, new_A3673_, new_A3674_, new_A3675_, new_A3676_, new_A3677_,
    new_A3678_, new_A3679_, new_A3680_, new_A3681_, new_A3682_, new_A3683_,
    new_A3684_, new_A3685_, new_A3686_, new_A3687_, new_A3688_, new_A3689_,
    new_A3690_, new_A3691_, new_A3692_, new_A3693_, new_A3694_, new_A3695_,
    new_A3696_, new_A3697_, new_A3698_, new_A3699_, new_A3700_, new_A3701_,
    new_A3702_, new_A3703_, new_A3704_, new_A3705_, new_A3706_, new_A3707_,
    new_A3708_, new_A3709_, new_A3710_, new_A3711_, new_A3712_, new_A3713_,
    new_A3714_, new_A3715_, new_A3716_, new_A3717_, new_A3718_, new_A3719_,
    new_A3720_, new_A3721_, new_A3722_, new_A3723_, new_A3724_, new_A3725_,
    new_A3726_, new_A3727_, new_A3728_, new_A3729_, new_A3730_, new_A3731_,
    new_A3732_, new_A3733_, new_A3734_, new_A3735_, new_A3736_, new_A3737_,
    new_A3738_, new_A3739_, new_A3740_, new_A3741_, new_A3742_, new_A3743_,
    new_A3744_, new_A3745_, new_A3746_, new_A3747_, new_A3748_, new_A3749_,
    new_A3750_, new_A3751_, new_A3752_, new_A3753_, new_A3754_, new_A3755_,
    new_A3756_, new_A3757_, new_A3758_, new_A3759_, new_A3760_, new_A3761_,
    new_A3762_, new_A3763_, new_A3764_, new_A3765_, new_A3766_, new_A3767_,
    new_A3768_, new_A3769_, new_A3770_, new_A3771_, new_A3772_, new_A3773_,
    new_A3774_, new_A3775_, new_A3776_, new_A3777_, new_A3778_, new_A3779_,
    new_A3780_, new_A3781_, new_A3782_, new_A3783_, new_A3784_, new_A3785_,
    new_A3786_, new_A3787_, new_A3788_, new_A3789_, new_A3790_, new_A3791_,
    new_A3792_, new_A3793_, new_A3794_, new_A3795_, new_A3796_, new_A3797_,
    new_A3798_, new_A3799_, new_A3800_, new_A3801_, new_A3802_, new_A3803_,
    new_A3804_, new_A3805_, new_A3806_, new_A3807_, new_A3808_, new_A3809_,
    new_A3810_, new_A3811_, new_A3812_, new_A3813_, new_A3814_, new_A3815_,
    new_A3816_, new_A3817_, new_A3818_, new_A3819_, new_A3820_, new_A3821_,
    new_A3822_, new_A3823_, new_A3824_, new_A3825_, new_A3826_, new_A3827_,
    new_A3828_, new_A3829_, new_A3830_, new_A3831_, new_A3832_, new_A3833_,
    new_A3834_, new_A3835_, new_A3836_, new_A3837_, new_A3838_, new_A3839_,
    new_A3840_, new_A3841_, new_A3842_, new_A3843_, new_A3844_, new_A3845_,
    new_A3846_, new_A3847_, new_A3848_, new_A3849_, new_A3850_, new_A3851_,
    new_A3852_, new_A3853_, new_A3854_, new_A3855_, new_A3856_, new_A3857_,
    new_A3858_, new_A3859_, new_A3860_, new_A3861_, new_A3862_, new_A3863_,
    new_A3864_, new_A3865_, new_A3866_, new_A3867_, new_A3868_, new_A3869_,
    new_A3870_, new_A3871_, new_A3872_, new_A3873_, new_A3874_, new_A3875_,
    new_A3876_, new_A3877_, new_A3878_, new_A3879_, new_A3880_, new_A3881_,
    new_A3882_, new_A3883_, new_A3884_, new_A3885_, new_A3886_, new_A3887_,
    new_A3888_, new_A3889_, new_A3890_, new_A3891_, new_A3892_, new_A3893_,
    new_A3894_, new_A3895_, new_A3896_, new_A3897_, new_A3898_, new_A3899_,
    new_A3900_, new_A3901_, new_A3902_, new_A3903_, new_A3904_, new_A3905_,
    new_A3906_, new_A3907_, new_A3908_, new_A3909_, new_A3910_, new_A3911_,
    new_A3912_, new_A3913_, new_A3914_, new_A3915_, new_A3916_, new_A3917_,
    new_A3918_, new_A3919_, new_A3920_, new_A3921_, new_A3922_, new_A3923_,
    new_A3924_, new_A3925_, new_A3926_, new_A3927_, new_A3928_, new_A3929_,
    new_A3930_, new_A3931_, new_A3932_, new_A3933_, new_A3934_, new_A3935_,
    new_A3936_, new_A3937_, new_A3938_, new_A3939_, new_A3940_, new_A3941_,
    new_A3942_, new_A3943_, new_A3944_, new_A3945_, new_A3946_, new_A3947_,
    new_A3948_, new_A3949_, new_A3950_, new_A3951_, new_A3952_, new_A3953_,
    new_A3954_, new_A3955_, new_A3956_, new_A3957_, new_A3958_, new_A3959_,
    new_A3960_, new_A3961_, new_A3962_, new_A3963_, new_A3964_, new_A3965_,
    new_A3966_, new_A3967_, new_A3968_, new_A3969_, new_A3970_, new_A3971_,
    new_A3972_, new_A3973_, new_A3974_, new_A3975_, new_A3976_, new_A3977_,
    new_A3978_, new_A3979_, new_A3980_, new_A3981_, new_A3982_, new_A3983_,
    new_A3984_, new_A3985_, new_A3986_, new_A3987_, new_A3988_, new_A3989_,
    new_A3990_, new_A3991_, new_A3992_, new_A3993_, new_A3994_, new_A3995_,
    new_A3996_, new_A3997_, new_A3998_, new_A3999_, new_A4000_, new_A4001_,
    new_A4002_, new_A4003_, new_A4004_, new_A4005_, new_A4006_, new_A4007_,
    new_A4008_, new_A4009_, new_A4010_, new_A4011_, new_A4012_, new_A4013_,
    new_A4014_, new_A4015_, new_A4016_, new_A4017_, new_A4018_, new_A4019_,
    new_A4020_, new_A4021_, new_A4022_, new_A4023_, new_A4024_, new_A4025_,
    new_A4026_, new_A4027_, new_A4028_, new_A4029_, new_A4030_, new_A4031_,
    new_A4032_, new_A4033_, new_A4034_, new_A4035_, new_A4036_, new_A4037_,
    new_A4038_, new_A4039_, new_A4040_, new_A4041_, new_A4042_, new_A4043_,
    new_A4044_, new_A4045_, new_A4046_, new_A4047_, new_A4048_, new_A4049_,
    new_A4050_, new_A4051_, new_A4052_, new_A4053_, new_A4054_, new_A4055_,
    new_A4056_, new_A4057_, new_A4058_, new_A4059_, new_A4060_, new_A4061_,
    new_A4062_, new_A4063_, new_A4064_, new_A4065_, new_A4066_, new_A4067_,
    new_A4068_, new_A4069_, new_A4070_, new_A4071_, new_A4072_, new_A4073_,
    new_A4074_, new_A4075_, new_A4076_, new_A4077_, new_A4078_, new_A4079_,
    new_A4080_, new_A4081_, new_A4082_, new_A4083_, new_A4084_, new_A4085_,
    new_A4086_, new_A4087_, new_A4088_, new_A4089_, new_A4090_, new_A4091_,
    new_A4092_, new_A4093_, new_A4094_, new_A4095_, new_A4096_, new_A4097_,
    new_A4098_, new_A4099_, new_A4100_, new_A4101_, new_A4102_, new_A4103_,
    new_A4104_, new_A4105_, new_A4106_, new_A4107_, new_A4108_, new_A4109_,
    new_A4110_, new_A4111_, new_A4112_, new_A4113_, new_A4114_, new_A4115_,
    new_A4116_, new_A4117_, new_A4118_, new_A4119_, new_A4120_, new_A4121_,
    new_A4122_, new_A4123_, new_A4124_, new_A4125_, new_A4126_, new_A4127_,
    new_A4128_, new_A4129_, new_A4130_, new_A4131_, new_A4132_, new_A4133_,
    new_A4134_, new_A4135_, new_A4136_, new_A4137_, new_A4138_, new_A4139_,
    new_A4140_, new_A4141_, new_A4142_, new_A4143_, new_A4144_, new_A4145_,
    new_A4146_, new_A4147_, new_A4148_, new_A4149_, new_A4150_, new_A4151_,
    new_A4152_, new_A4153_, new_A4154_, new_A4155_, new_A4156_, new_A4157_,
    new_A4158_, new_A4159_, new_A4160_, new_A4161_, new_A4162_, new_A4163_,
    new_A4164_, new_A4165_, new_A4166_, new_A4167_, new_A4168_, new_A4169_,
    new_A4170_, new_A4171_, new_A4172_, new_A4173_, new_A4174_, new_A4175_,
    new_A4176_, new_A4177_, new_A4178_, new_A4179_, new_A4180_, new_A4181_,
    new_A4182_, new_A4183_, new_A4184_, new_A4185_, new_A4186_, new_A4187_,
    new_A4188_, new_A4189_, new_A4190_, new_A4191_, new_A4192_, new_A4193_,
    new_A4194_, new_A4195_, new_A4196_, new_A4197_, new_A4198_, new_A4199_,
    new_A4200_, new_A4201_, new_A4202_, new_A4203_, new_A4204_, new_A4205_,
    new_A4206_, new_A4207_, new_A4208_, new_A4209_, new_A4210_, new_A4211_,
    new_A4212_, new_A4213_, new_A4214_, new_A4215_, new_A4216_, new_A4217_,
    new_A4218_, new_A4219_, new_A4220_, new_A4221_, new_A4222_, new_A4223_,
    new_A4224_, new_A4225_, new_A4226_, new_A4227_, new_A4228_, new_A4229_,
    new_A4230_, new_A4231_, new_A4232_, new_A4233_, new_A4234_, new_A4235_,
    new_A4236_, new_A4237_, new_A4238_, new_A4239_, new_A4240_, new_A4241_,
    new_A4242_, new_A4243_, new_A4244_, new_A4245_, new_A4246_, new_A4247_,
    new_A4248_, new_A4249_, new_A4250_, new_A4251_, new_A4252_, new_A4253_,
    new_A4254_, new_A4255_, new_A4256_, new_A4257_, new_A4258_, new_A4259_,
    new_A4260_, new_A4261_, new_A4262_, new_A4263_, new_A4264_, new_A4265_,
    new_A4266_, new_A4267_, new_A4268_, new_A4269_, new_A4270_, new_A4271_,
    new_A4272_, new_A4273_, new_A4274_, new_A4275_, new_A4276_, new_A4277_,
    new_A4278_, new_A4279_, new_A4280_, new_A4281_, new_A4282_, new_A4283_,
    new_A4284_, new_A4285_, new_A4286_, new_A4287_, new_A4288_, new_A4289_,
    new_A4290_, new_A4291_, new_A4292_, new_A4293_, new_A4294_, new_A4295_,
    new_A4296_, new_A4297_, new_A4298_, new_A4299_, new_A4300_, new_A4301_,
    new_A4302_, new_A4303_, new_A4304_, new_A4305_, new_A4306_, new_A4307_,
    new_A4308_, new_A4309_, new_A4310_, new_A4311_, new_A4312_, new_A4313_,
    new_A4314_, new_A4315_, new_A4316_, new_A4317_, new_A4318_, new_A4319_,
    new_A4320_, new_A4321_, new_A4322_, new_A4323_, new_A4324_, new_A4325_,
    new_A4326_, new_A4327_, new_A4328_, new_A4329_, new_A4330_, new_A4331_,
    new_A4332_, new_A4333_, new_A4334_, new_A4335_, new_A4336_, new_A4337_,
    new_A4338_, new_A4339_, new_A4340_, new_A4341_, new_A4342_, new_A4343_,
    new_A4344_, new_A4345_, new_A4346_, new_A4347_, new_A4348_, new_A4349_,
    new_A4350_, new_A4351_, new_A4352_, new_A4353_, new_A4354_, new_A4355_,
    new_A4356_, new_A4357_, new_A4358_, new_A4359_, new_A4360_, new_A4361_,
    new_A4362_, new_A4363_, new_A4364_, new_A4365_, new_A4366_, new_A4367_,
    new_A4368_, new_A4369_, new_A4370_, new_A4371_, new_A4372_, new_A4373_,
    new_A4374_, new_A4375_, new_A4376_, new_A4377_, new_A4378_, new_A4379_,
    new_A4380_, new_A4381_, new_A4382_, new_A4383_, new_A4384_, new_A4385_,
    new_A4386_, new_A4387_, new_A4388_, new_A4389_, new_A4390_, new_A4391_,
    new_A4392_, new_A4393_, new_A4394_, new_A4395_, new_A4396_, new_A4397_,
    new_A4398_, new_A4399_, new_A4400_, new_A4401_, new_A4402_, new_A4403_,
    new_A4404_, new_A4405_, new_A4406_, new_A4407_, new_A4408_, new_A4409_,
    new_A4410_, new_A4411_, new_A4412_, new_A4413_, new_A4414_, new_A4415_,
    new_A4416_, new_A4417_, new_A4418_, new_A4419_, new_A4420_, new_A4421_,
    new_A4422_, new_A4423_, new_A4424_, new_A4425_, new_A4426_, new_A4427_,
    new_A4428_, new_A4429_, new_A4430_, new_A4431_, new_A4432_, new_A4433_,
    new_A4434_, new_A4435_, new_A4436_, new_A4437_, new_A4438_, new_A4439_,
    new_A4440_, new_A4441_, new_A4442_, new_A4443_, new_A4444_, new_A4445_,
    new_A4446_, new_A4447_, new_A4448_, new_A4449_, new_A4450_, new_A4451_,
    new_A4452_, new_A4453_, new_A4454_, new_A4455_, new_A4456_, new_A4457_,
    new_A4458_, new_A4459_, new_A4460_, new_A4461_, new_A4462_, new_A4463_,
    new_A4464_, new_A4465_, new_A4466_, new_A4467_, new_A4468_, new_A4469_,
    new_A4470_, new_A4471_, new_A4472_, new_A4473_, new_A4474_, new_A4475_,
    new_A4476_, new_A4477_, new_A4478_, new_A4479_, new_A4480_, new_A4481_,
    new_A4482_, new_A4483_, new_A4484_, new_A4485_, new_A4486_, new_A4487_,
    new_A4488_, new_A4489_, new_A4490_, new_A4491_, new_A4492_, new_A4493_,
    new_A4494_, new_A4495_, new_A4496_, new_A4497_, new_A4498_, new_A4499_,
    new_A4500_, new_A4501_, new_A4502_, new_A4503_, new_A4504_, new_A4505_,
    new_A4506_, new_A4507_, new_A4508_, new_A4509_, new_A4510_, new_A4511_,
    new_A4512_, new_A4513_, new_A4514_, new_A4515_, new_A4516_, new_A4517_,
    new_A4518_, new_A4519_, new_A4520_, new_A4521_, new_A4522_, new_A4523_,
    new_A4524_, new_A4525_, new_A4526_, new_A4527_, new_A4528_, new_A4529_,
    new_A4530_, new_A4531_, new_A4532_, new_A4533_, new_A4534_, new_A4535_,
    new_A4536_, new_A4537_, new_A4538_, new_A4539_, new_A4540_, new_A4541_,
    new_A4542_, new_A4543_, new_A4544_, new_A4545_, new_A4546_, new_A4547_,
    new_A4548_, new_A4549_, new_A4550_, new_A4551_, new_A4552_, new_A4553_,
    new_A4554_, new_A4555_, new_A4556_, new_A4557_, new_A4558_, new_A4559_,
    new_A4560_, new_A4561_, new_A4562_, new_A4563_, new_A4564_, new_A4565_,
    new_A4566_, new_A4567_, new_A4568_, new_A4569_, new_A4570_, new_A4571_,
    new_A4572_, new_A4573_, new_A4574_, new_A4575_, new_A4576_, new_A4577_,
    new_A4578_, new_A4579_, new_A4580_, new_A4581_, new_A4582_, new_A4583_,
    new_A4584_, new_A4585_, new_A4586_, new_A4587_, new_A4588_, new_A4589_,
    new_A4590_, new_A4591_, new_A4592_, new_A4593_, new_A4594_, new_A4595_,
    new_A4596_, new_A4597_, new_A4598_, new_A4599_, new_A4600_, new_A4601_,
    new_A4602_, new_A4603_, new_A4604_, new_A4605_, new_A4606_, new_A4607_,
    new_A4608_, new_A4609_, new_A4610_, new_A4611_, new_A4612_, new_A4613_,
    new_A4614_, new_A4615_, new_A4616_, new_A4617_, new_A4618_, new_A4619_,
    new_A4620_, new_A4621_, new_A4622_, new_A4623_, new_A4624_, new_A4625_,
    new_A4626_, new_A4627_, new_A4628_, new_A4629_, new_A4630_, new_A4631_,
    new_A4632_, new_A4633_, new_A4634_, new_A4635_, new_A4636_, new_A4637_,
    new_A4638_, new_A4639_, new_A4640_, new_A4641_, new_A4642_, new_A4643_,
    new_A4644_, new_A4645_, new_A4646_, new_A4647_, new_A4648_, new_A4649_,
    new_A4650_, new_A4651_, new_A4652_, new_A4653_, new_A4654_, new_A4655_,
    new_A4656_, new_A4657_, new_A4658_, new_A4659_, new_A4660_, new_A4661_,
    new_A4662_, new_A4663_, new_A4664_, new_A4665_, new_A4666_, new_A4667_,
    new_A4668_, new_A4669_, new_A4670_, new_A4671_, new_A4672_, new_A4673_,
    new_A4674_, new_A4675_, new_A4676_, new_A4677_, new_A4678_, new_A4679_,
    new_A4680_, new_A4681_, new_A4682_, new_A4683_, new_A4684_, new_A4685_,
    new_A4686_, new_A4687_, new_A4688_, new_A4689_, new_A4690_, new_A4691_,
    new_A4692_, new_A4693_, new_A4694_, new_A4695_, new_A4696_, new_A4697_,
    new_A4698_, new_A4699_, new_A4700_, new_A4701_, new_A4702_, new_A4703_,
    new_A4704_, new_A4705_, new_A4706_, new_A4707_, new_A4708_, new_A4709_,
    new_A4710_, new_A4711_, new_A4712_, new_A4713_, new_A4714_, new_A4715_,
    new_A4716_, new_A4717_, new_A4718_, new_A4719_, new_A4720_, new_A4721_,
    new_A4722_, new_A4723_, new_A4724_, new_A4725_, new_A4726_, new_A4727_,
    new_A4728_, new_A4729_, new_A4730_, new_A4731_, new_A4732_, new_A4733_,
    new_A4734_, new_A4735_, new_A4736_, new_A4737_, new_A4738_, new_A4739_,
    new_A4740_, new_A4741_, new_A4742_, new_A4743_, new_A4744_, new_A4745_,
    new_A4746_, new_A4747_, new_A4748_, new_A4749_, new_A4750_, new_A4751_,
    new_A4752_, new_A4753_, new_A4754_, new_A4755_, new_A4756_, new_A4757_,
    new_A4758_, new_A4759_, new_A4760_, new_A4761_, new_A4762_, new_A4763_,
    new_A4764_, new_A4765_, new_A4766_, new_A4767_, new_A4768_, new_A4769_,
    new_A4770_, new_A4771_, new_A4772_, new_A4773_, new_A4774_, new_A4775_,
    new_A4776_, new_A4777_, new_A4778_, new_A4779_, new_A4780_, new_A4781_,
    new_A4782_, new_A4783_, new_A4784_, new_A4785_, new_A4786_, new_A4787_,
    new_A4788_, new_A4789_, new_A4790_, new_A4791_, new_A4792_, new_A4793_,
    new_A4794_, new_A4795_, new_A4796_, new_A4797_, new_A4798_, new_A4799_,
    new_A4800_, new_A4801_, new_A4802_, new_A4803_, new_A4804_, new_A4805_,
    new_A4806_, new_A4807_, new_A4808_, new_A4809_, new_A4810_, new_A4811_,
    new_A4812_, new_A4813_, new_A4814_, new_A4815_, new_A4816_, new_A4817_,
    new_A4818_, new_A4819_, new_A4820_, new_A4821_, new_A4822_, new_A4823_,
    new_A4824_, new_A4825_, new_A4826_, new_A4827_, new_A4828_, new_A4829_,
    new_A4830_, new_A4831_, new_A4832_, new_A4833_, new_A4834_, new_A4835_,
    new_A4836_, new_A4837_, new_A4838_, new_A4839_, new_A4840_, new_A4841_,
    new_A4842_, new_A4843_, new_A4844_, new_A4845_, new_A4846_, new_A4847_,
    new_A4848_, new_A4849_, new_A4850_, new_A4851_, new_A4852_, new_A4853_,
    new_A4854_, new_A4855_, new_A4856_, new_A4857_, new_A4858_, new_A4859_,
    new_A4860_, new_A4861_, new_A4862_, new_A4863_, new_A4864_, new_A4865_,
    new_A4866_, new_A4867_, new_A4868_, new_A4869_, new_A4870_, new_A4871_,
    new_A4872_, new_A4873_, new_A4874_, new_A4875_, new_A4876_, new_A4877_,
    new_A4878_, new_A4879_, new_A4880_, new_A4881_, new_A4882_, new_A4883_,
    new_A4884_, new_A4885_, new_A4886_, new_A4887_, new_A4888_, new_A4889_,
    new_A4890_, new_A4891_, new_A4892_, new_A4893_, new_A4894_, new_A4895_,
    new_A4896_, new_A4897_, new_A4898_, new_A4899_, new_A4900_, new_A4901_,
    new_A4902_, new_A4903_, new_A4904_, new_A4905_, new_A4906_, new_A4907_,
    new_A4908_, new_A4909_, new_A4910_, new_A4911_, new_A4912_, new_A4913_,
    new_A4914_, new_A4915_, new_A4916_, new_A4917_, new_A4918_, new_A4919_,
    new_A4920_, new_A4921_, new_A4922_, new_A4923_, new_A4924_, new_A4925_,
    new_A4926_, new_A4927_, new_A4928_, new_A4929_, new_A4930_, new_A4931_,
    new_A4932_, new_A4933_, new_A4934_, new_A4935_, new_A4936_, new_A4937_,
    new_A4938_, new_A4939_, new_A4940_, new_A4941_, new_A4942_, new_A4943_,
    new_A4944_, new_A4945_, new_A4946_, new_A4947_, new_A4948_, new_A4949_,
    new_A4950_, new_A4951_, new_A4952_, new_A4953_, new_A4954_, new_A4955_,
    new_A4956_, new_A4957_, new_A4958_, new_A4959_, new_A4960_, new_A4961_,
    new_A4962_, new_A4963_, new_A4964_, new_A4965_, new_A4966_, new_A4967_,
    new_A4968_, new_A4969_, new_A4970_, new_A4971_, new_A4972_, new_A4973_,
    new_A4974_, new_A4975_, new_A4976_, new_A4977_, new_A4978_, new_A4979_,
    new_A4980_, new_A4981_, new_A4982_, new_A4983_, new_A4984_, new_A4985_,
    new_A4986_, new_A4987_, new_A4988_, new_A4989_, new_A4990_, new_A4991_,
    new_A4992_, new_A4993_, new_A4994_, new_A4995_, new_A4996_, new_A4997_,
    new_A4998_, new_A4999_, new_A5000_, new_A5001_, new_A5002_, new_A5003_,
    new_A5004_, new_A5005_, new_A5006_, new_A5007_, new_A5008_, new_A5009_,
    new_A5010_, new_A5011_, new_A5012_, new_A5013_, new_A5014_, new_A5015_,
    new_A5016_, new_A5017_, new_A5018_, new_A5019_, new_A5020_, new_A5021_,
    new_A5022_, new_A5023_, new_A5024_, new_A5025_, new_A5026_, new_A5027_,
    new_A5028_, new_A5029_, new_A5030_, new_A5031_, new_A5032_, new_A5033_,
    new_A5034_, new_A5035_, new_A5036_, new_A5037_, new_A5038_, new_A5039_,
    new_A5040_, new_A5041_, new_A5042_, new_A5043_, new_A5044_, new_A5045_,
    new_A5046_, new_A5047_, new_A5048_, new_A5049_, new_A5050_, new_A5051_,
    new_A5052_, new_A5053_, new_A5054_, new_A5055_, new_A5056_, new_A5057_,
    new_A5058_, new_A5059_, new_A5060_, new_A5061_, new_A5062_, new_A5063_,
    new_A5064_, new_A5065_, new_A5066_, new_A5067_, new_A5068_, new_A5069_,
    new_A5070_, new_A5071_, new_A5072_, new_A5073_, new_A5074_, new_A5075_,
    new_A5076_, new_A5077_, new_A5078_, new_A5079_, new_A5080_, new_A5081_,
    new_A5082_, new_A5083_, new_A5084_, new_A5085_, new_A5086_, new_A5087_,
    new_A5088_, new_A5089_, new_A5090_, new_A5091_, new_A5092_, new_A5093_,
    new_A5094_, new_A5095_, new_A5096_, new_A5097_, new_A5098_, new_A5099_,
    new_A5100_, new_A5101_, new_A5102_, new_A5103_, new_A5104_, new_A5105_,
    new_A5106_, new_A5107_, new_A5108_, new_A5109_, new_A5110_, new_A5111_,
    new_A5112_, new_A5113_, new_A5114_, new_A5115_, new_A5116_, new_A5117_,
    new_A5118_, new_A5119_, new_A5120_, new_A5121_, new_A5122_, new_A5123_,
    new_A5124_, new_A5125_, new_A5126_, new_A5127_, new_A5128_, new_A5129_,
    new_A5130_, new_A5131_, new_A5132_, new_A5133_, new_A5134_, new_A5135_,
    new_A5136_, new_A5137_, new_A5138_, new_A5139_, new_A5140_, new_A5141_,
    new_A5142_, new_A5143_, new_A5144_, new_A5145_, new_A5146_, new_A5147_,
    new_A5148_, new_A5149_, new_A5150_, new_A5151_, new_A5152_, new_A5153_,
    new_A5154_, new_A5155_, new_A5156_, new_A5157_, new_A5158_, new_A5159_,
    new_A5160_, new_A5161_, new_A5162_, new_A5163_, new_A5164_, new_A5165_,
    new_A5166_, new_A5167_, new_A5168_, new_A5169_, new_A5170_, new_A5171_,
    new_A5172_, new_A5173_, new_A5174_, new_A5175_, new_A5176_, new_A5177_,
    new_A5178_, new_A5179_, new_A5180_, new_A5181_, new_A5182_, new_A5183_,
    new_A5184_, new_A5185_, new_A5186_, new_A5187_, new_A5188_, new_A5189_,
    new_A5190_, new_A5191_, new_A5192_, new_A5193_, new_A5194_, new_A5195_,
    new_A5196_, new_A5197_, new_A5198_, new_A5199_, new_A5200_, new_A5201_,
    new_A5202_, new_A5203_, new_A5204_, new_A5205_, new_A5206_, new_A5207_,
    new_A5208_, new_A5209_, new_A5210_, new_A5211_, new_A5212_, new_A5213_,
    new_A5214_, new_A5215_, new_A5216_, new_A5217_, new_A5218_, new_A5219_,
    new_A5220_, new_A5221_, new_A5222_, new_A5223_, new_A5224_, new_A5225_,
    new_A5226_, new_A5227_, new_A5228_, new_A5229_, new_A5230_, new_A5231_,
    new_A5232_, new_A5233_, new_A5234_, new_A5235_, new_A5236_, new_A5237_,
    new_A5238_, new_A5239_, new_A5240_, new_A5241_, new_A5242_, new_A5243_,
    new_A5244_, new_A5245_, new_A5246_, new_A5247_, new_A5248_, new_A5249_,
    new_A5250_, new_A5251_, new_A5252_, new_A5253_, new_A5254_, new_A5255_,
    new_A5256_, new_A5257_, new_A5258_, new_A5259_, new_A5260_, new_A5261_,
    new_A5262_, new_A5263_, new_A5264_, new_A5265_, new_A5266_, new_A5267_,
    new_A5268_, new_A5269_, new_A5270_, new_A5271_, new_A5272_, new_A5273_,
    new_A5274_, new_A5275_, new_A5276_, new_A5277_, new_A5278_, new_A5279_,
    new_A5280_, new_A5281_, new_A5282_, new_A5283_, new_A5284_, new_A5285_,
    new_A5286_, new_A5287_, new_A5288_, new_A5289_, new_A5290_, new_A5291_,
    new_A5292_, new_A5293_, new_A5294_, new_A5295_, new_A5296_, new_A5297_,
    new_A5298_, new_A5299_, new_A5300_, new_A5301_, new_A5302_, new_A5303_,
    new_A5304_, new_A5305_, new_A5306_, new_A5307_, new_A5308_, new_A5309_,
    new_A5310_, new_A5311_, new_A5312_, new_A5313_, new_A5314_, new_A5315_,
    new_A5316_, new_A5317_, new_A5318_, new_A5319_, new_A5320_, new_A5321_,
    new_A5322_, new_A5323_, new_A5324_, new_A5325_, new_A5326_, new_A5327_,
    new_A5328_, new_A5329_, new_A5330_, new_A5331_, new_A5332_, new_A5333_,
    new_A5334_, new_A5335_, new_A5336_, new_A5337_, new_A5338_, new_A5339_,
    new_A5340_, new_A5341_, new_A5342_, new_A5343_, new_A5344_, new_A5345_,
    new_A5346_, new_A5347_, new_A5348_, new_A5349_, new_A5350_, new_A5351_,
    new_A5352_, new_A5353_, new_A5354_, new_A5355_, new_A5356_, new_A5357_,
    new_A5358_, new_A5359_, new_A5360_, new_A5361_, new_A5362_, new_A5363_,
    new_A5364_, new_A5365_, new_A5366_, new_A5367_, new_A5368_, new_A5369_,
    new_A5370_, new_A5371_, new_A5372_, new_A5373_, new_A5374_, new_A5375_,
    new_A5376_, new_A5377_, new_A5378_, new_A5379_, new_A5380_, new_A5381_,
    new_A5382_, new_A5383_, new_A5384_, new_A5385_, new_A5386_, new_A5387_,
    new_A5388_, new_A5389_, new_A5390_, new_A5391_, new_A5392_, new_A5393_,
    new_A5394_, new_A5395_, new_A5396_, new_A5397_, new_A5398_, new_A5399_,
    new_A5400_, new_A5401_, new_A5402_, new_A5403_, new_A5404_, new_A5405_,
    new_A5406_, new_A5407_, new_A5408_, new_A5409_, new_A5410_, new_A5411_,
    new_A5412_, new_A5413_, new_A5414_, new_A5415_, new_A5416_, new_A5417_,
    new_A5418_, new_A5419_, new_A5420_, new_A5421_, new_A5422_, new_A5423_,
    new_A5424_, new_A5425_, new_A5426_, new_A5427_, new_A5428_, new_A5429_,
    new_A5430_, new_A5431_, new_A5432_, new_A5433_, new_A5434_, new_A5435_,
    new_A5436_, new_A5437_, new_A5438_, new_A5439_, new_A5440_, new_A5441_,
    new_A5442_, new_A5443_, new_A5444_, new_A5445_, new_A5446_, new_A5447_,
    new_A5448_, new_A5449_, new_A5450_, new_A5451_, new_A5452_, new_A5453_,
    new_A5454_, new_A5455_, new_A5456_, new_A5457_, new_A5458_, new_A5459_,
    new_A5460_, new_A5461_, new_A5462_, new_A5463_, new_A5464_, new_A5465_,
    new_A5466_, new_A5467_, new_A5468_, new_A5469_, new_A5470_, new_A5471_,
    new_A5472_, new_A5473_, new_A5474_, new_A5475_, new_A5476_, new_A5477_,
    new_A5478_, new_A5479_, new_A5480_, new_A5481_, new_A5482_, new_A5483_,
    new_A5484_, new_A5485_, new_A5486_, new_A5487_, new_A5488_, new_A5489_,
    new_A5490_, new_A5491_, new_A5492_, new_A5493_, new_A5494_, new_A5495_,
    new_A5496_, new_A5497_, new_A5498_, new_A5499_, new_A5500_, new_A5501_,
    new_A5502_, new_A5503_, new_A5504_, new_A5505_, new_A5506_, new_A5507_,
    new_A5508_, new_A5509_, new_A5510_, new_A5511_, new_A5512_, new_A5513_,
    new_A5514_, new_A5515_, new_A5516_, new_A5517_, new_A5518_, new_A5519_,
    new_A5520_, new_A5521_, new_A5522_, new_A5523_, new_A5524_, new_A5525_,
    new_A5526_, new_A5527_, new_A5528_, new_A5529_, new_A5530_, new_A5531_,
    new_A5532_, new_A5533_, new_A5534_, new_A5535_, new_A5536_, new_A5537_,
    new_A5538_, new_A5539_, new_A5540_, new_A5541_, new_A5542_, new_A5543_,
    new_A5544_, new_A5545_, new_A5546_, new_A5547_, new_A5548_, new_A5549_,
    new_A5550_, new_A5551_, new_A5552_, new_A5553_, new_A5554_, new_A5555_,
    new_A5556_, new_A5557_, new_A5558_, new_A5559_, new_A5560_, new_A5561_,
    new_A5562_, new_A5563_, new_A5564_, new_A5565_, new_A5566_, new_A5567_,
    new_A5568_, new_A5569_, new_A5570_, new_A5571_, new_A5572_, new_A5573_,
    new_A5574_, new_A5575_, new_A5576_, new_A5577_, new_A5578_, new_A5579_,
    new_A5580_, new_A5581_, new_A5582_, new_A5583_, new_A5584_, new_A5585_,
    new_A5586_, new_A5587_, new_A5588_, new_A5589_, new_A5590_, new_A5591_,
    new_A5592_, new_A5593_, new_A5594_, new_A5595_, new_A5596_, new_A5597_,
    new_A5598_, new_A5599_, new_A5600_, new_A5601_, new_A5602_, new_A5603_,
    new_A5604_, new_A5605_, new_A5606_, new_A5607_, new_A5608_, new_A5609_,
    new_A5610_, new_A5611_, new_A5612_, new_A5613_, new_A5614_, new_A5615_,
    new_A5616_, new_A5617_, new_A5618_, new_A5619_, new_A5620_, new_A5621_,
    new_A5622_, new_A5623_, new_A5624_, new_A5625_, new_A5626_, new_A5627_,
    new_A5628_, new_A3216_, new_A3215_, new_A3214_, new_A3213_, new_A3212_,
    new_A3211_, new_A3210_, new_A3209_, new_A3208_, new_A3207_, new_A3206_,
    new_A3205_, new_A3204_, new_A3203_, new_A3202_, new_A3201_, new_A3200_,
    new_A3199_, new_A3198_, new_A3197_, new_A3196_, new_A3195_, new_A3194_,
    new_A3193_, new_A3192_, new_A3191_, new_A3190_, new_A3189_, new_A3188_,
    new_A3187_, new_A3186_, new_A3185_, new_A3184_, new_A3183_, new_A3182_,
    new_A3181_, new_A3180_, new_A3179_, new_A3178_, new_A3177_, new_A3176_,
    new_A3175_, new_A3174_, new_A3173_, new_A3172_, new_A3171_, new_A3170_,
    new_A3169_, new_A3168_, new_A3167_, new_A3166_, new_A3165_, new_A3164_,
    new_A3163_, new_A3162_, new_A3155_, new_A3154_, new_A3153_, new_A3152_,
    new_A3151_, new_A3150_, new_A3149_, new_A3148_, new_A3147_, new_A3146_,
    new_A3145_, new_A3144_, new_A3143_, new_A3142_, new_A3141_, new_A3140_,
    new_A3139_, new_A3138_, new_A3137_, new_A3136_, new_A3135_, new_A3134_,
    new_A3133_, new_A3132_, new_A3131_, new_A3130_, new_A3129_, new_A3128_,
    new_A3127_, new_A3126_, new_A3125_, new_A3124_, new_A3123_, new_A3122_,
    new_A3121_, new_A3120_, new_A3119_, new_A3118_, new_A3117_, new_A3116_,
    new_A3115_, new_A3114_, new_A3113_, new_A3112_, new_A3111_, new_A3110_,
    new_A3109_, new_A3108_, new_A3107_, new_A3106_, new_A3105_, new_A3104_,
    new_A3103_, new_A3102_, new_A3101_, new_A3100_, new_A3099_, new_A3098_,
    new_A3097_, new_A3096_, new_A3095_, new_A3088_, new_A3087_, new_A3086_,
    new_A3085_, new_A3084_, new_A3083_, new_A3082_, new_A3081_, new_A3080_,
    new_A3079_, new_A3078_, new_A3077_, new_A3076_, new_A3075_, new_A3074_,
    new_A3073_, new_A3072_, new_A3071_, new_A3070_, new_A3069_, new_A3068_,
    new_A3067_, new_A3066_, new_A3065_, new_A3064_, new_A3063_, new_A3062_,
    new_A3061_, new_A3060_, new_A3059_, new_A3058_, new_A3057_, new_A3056_,
    new_A3055_, new_A3054_, new_A3053_, new_A3052_, new_A3051_, new_A3050_,
    new_A3049_, new_A3048_, new_A3047_, new_A3046_, new_A3045_, new_A3044_,
    new_A3043_, new_A3042_, new_A3041_, new_A3040_, new_A3039_, new_A3038_,
    new_A3037_, new_A3036_, new_A3035_, new_A3034_, new_A3033_, new_A3032_,
    new_A3031_, new_A3030_, new_A3029_, new_A3028_, new_A3021_, new_A3020_,
    new_A3019_, new_A3018_, new_A3017_, new_A3016_, new_A3015_, new_A3014_,
    new_A3013_, new_A3012_, new_A3011_, new_A3010_, new_A3009_, new_A3008_,
    new_A3007_, new_A3006_, new_A3005_, new_A3004_, new_A3003_, new_A3002_,
    new_A3001_, new_A3000_, new_A2999_, new_A2998_, new_A2997_, new_A2996_,
    new_A2995_, new_A2994_, new_A2993_, new_A2992_, new_A2991_, new_A2990_,
    new_A2989_, new_A2988_, new_A2987_, new_A2986_, new_A2985_, new_A2984_,
    new_A2983_, new_A2982_, new_A2981_, new_A2980_, new_A2979_, new_A2978_,
    new_A2977_, new_A2976_, new_A2975_, new_A2974_, new_A2973_, new_A2972_,
    new_A2971_, new_A2970_, new_A2969_, new_A2968_, new_A2967_, new_A2966_,
    new_A2965_, new_A2964_, new_A2963_, new_A2962_, new_A2961_, new_A2954_,
    new_A2953_, new_A2952_, new_A2951_, new_A2950_, new_A2949_, new_A2948_,
    new_A2947_, new_A2946_, new_A2945_, new_A2944_, new_A2943_, new_A2942_,
    new_A2941_, new_A2940_, new_A2939_, new_A2938_, new_A2937_, new_A2936_,
    new_A2935_, new_A2934_, new_A2933_, new_A2932_, new_A2931_, new_A2930_,
    new_A2929_, new_A2928_, new_A2927_, new_A2926_, new_A2925_, new_A2924_,
    new_A2923_, new_A2922_, new_A2921_, new_A2920_, new_A2919_, new_A2918_,
    new_A2917_, new_A2916_, new_A2915_, new_A2914_, new_A2913_, new_A2912_,
    new_A2911_, new_A2910_, new_A2909_, new_A2908_, new_A2907_, new_A2906_,
    new_A2905_, new_A2904_, new_A2903_, new_A2902_, new_A2901_, new_A2900_,
    new_A2899_, new_A2898_, new_A2897_, new_A2896_, new_A2895_, new_A2894_,
    new_A2887_, new_A2886_, new_A2885_, new_A2884_, new_A2883_, new_A2882_,
    new_A2881_, new_A2880_, new_A2879_, new_A2878_, new_A2877_, new_A2876_,
    new_A2875_, new_A2874_, new_A2873_, new_A2872_, new_A2871_, new_A2870_,
    new_A2869_, new_A2868_, new_A2867_, new_A2866_, new_A2865_, new_A2864_,
    new_A2863_, new_A2862_, new_A2861_, new_A2860_, new_A2859_, new_A2858_,
    new_A2857_, new_A2856_, new_A2855_, new_A2854_, new_A2853_, new_A2852_,
    new_A2851_, new_A2850_, new_A2849_, new_A2848_, new_A2847_, new_A2846_,
    new_A2845_, new_A2844_, new_A2843_, new_A2842_, new_A2841_, new_A2840_,
    new_A2839_, new_A2838_, new_A2837_, new_A2836_, new_A2835_, new_A2834_,
    new_A2833_, new_A2832_, new_A2831_, new_A2830_, new_A2829_, new_A2828_,
    new_A2827_, new_A2820_, new_A2819_, new_A2818_, new_A2817_, new_A2816_,
    new_A2815_, new_A2814_, new_A2813_, new_A2812_, new_A2811_, new_A2810_,
    new_A2809_, new_A2808_, new_A2807_, new_A2806_, new_A2805_, new_A2804_,
    new_A2803_, new_A2802_, new_A2801_, new_A2800_, new_A2799_, new_A2798_,
    new_A2797_, new_A2796_, new_A2795_, new_A2794_, new_A2793_, new_A2792_,
    new_A2791_, new_A2790_, new_A2789_, new_A2788_, new_A2787_, new_A2786_,
    new_A2785_, new_A2784_, new_A2783_, new_A2782_, new_A2781_, new_A2780_,
    new_A2779_, new_A2778_, new_A2777_, new_A2776_, new_A2775_, new_A2774_,
    new_A2773_, new_A2772_, new_A2771_, new_A2770_, new_A2769_, new_A2768_,
    new_A2767_, new_A2766_, new_A2765_, new_A2764_, new_A2763_, new_A2762_,
    new_A2761_, new_A2760_, new_A2753_, new_A2752_, new_A2751_, new_A2750_,
    new_A2749_, new_A2748_, new_A2747_, new_A2746_, new_A2745_, new_A2744_,
    new_A2743_, new_A2742_, new_A2741_, new_A2740_, new_A2739_, new_A2738_,
    new_A2737_, new_A2736_, new_A2735_, new_A2734_, new_A2733_, new_A2732_,
    new_A2731_, new_A2730_, new_A2729_, new_A2728_, new_A2727_, new_A2726_,
    new_A2725_, new_A2724_, new_A2723_, new_A2722_, new_A2721_, new_A2720_,
    new_A2719_, new_A2718_, new_A2717_, new_A2716_, new_A2715_, new_A2714_,
    new_A2713_, new_A2712_, new_A2711_, new_A2710_, new_A2709_, new_A2708_,
    new_A2707_, new_A2706_, new_A2705_, new_A2704_, new_A2703_, new_A2702_,
    new_A2701_, new_A2700_, new_A2699_, new_A2698_, new_A2697_, new_A2696_,
    new_A2695_, new_A2694_, new_A2693_, new_A2686_, new_A2685_, new_A2684_,
    new_A2683_, new_A2682_, new_A2681_, new_A2680_, new_A2679_, new_A2678_,
    new_A2677_, new_A2676_, new_A2675_, new_A2674_, new_A2673_, new_A2672_,
    new_A2671_, new_A2670_, new_A2669_, new_A2668_, new_A2667_, new_A2666_,
    new_A2665_, new_A2664_, new_A2663_, new_A2662_, new_A2661_, new_A2660_,
    new_A2659_, new_A2658_, new_A2657_, new_A2656_, new_A2655_, new_A2654_,
    new_A2653_, new_A2652_, new_A2651_, new_A2650_, new_A2649_, new_A2648_,
    new_A2647_, new_A2646_, new_A2645_, new_A2644_, new_A2643_, new_A2642_,
    new_A2641_, new_A2640_, new_A2639_, new_A2638_, new_A2637_, new_A2636_,
    new_A2635_, new_A2634_, new_A2633_, new_A2632_, new_A2631_, new_A2630_,
    new_A2629_, new_A2628_, new_A2627_, new_A2626_, new_A2619_, new_A2618_,
    new_A2617_, new_A2616_, new_A2615_, new_A2614_, new_A2613_, new_A2612_,
    new_A2611_, new_A2610_, new_A2609_, new_A2608_, new_A2607_, new_A2606_,
    new_A2605_, new_A2604_, new_A2603_, new_A2602_, new_A2601_, new_A2600_,
    new_A2599_, new_A2598_, new_A2597_, new_A2596_, new_A2595_, new_A2594_,
    new_A2593_, new_A2592_, new_A2591_, new_A2590_, new_A2589_, new_A2588_,
    new_A2587_, new_A2586_, new_A2585_, new_A2584_, new_A2583_, new_A2582_,
    new_A2581_, new_A2580_, new_A2579_, new_A2578_, new_A2577_, new_A2576_,
    new_A2575_, new_A2574_, new_A2573_, new_A2572_, new_A2571_, new_A2570_,
    new_A2569_, new_A2568_, new_A2567_, new_A2566_, new_A2565_, new_A2564_,
    new_A2563_, new_A2562_, new_A2561_, new_A2560_, new_A2559_, new_A2552_,
    new_A2551_, new_A2550_, new_A2549_, new_A2548_, new_A2547_, new_A2546_,
    new_A2545_, new_A2544_, new_A2543_, new_A2542_, new_A2541_, new_A2540_,
    new_A2539_, new_A2538_, new_A2537_, new_A2536_, new_A2535_, new_A2534_,
    new_A2533_, new_A2532_, new_A2531_, new_A2530_, new_A2529_, new_A2528_,
    new_A2527_, new_A2526_, new_A2525_, new_A2524_, new_A2523_, new_A2522_,
    new_A2521_, new_A2520_, new_A2519_, new_A2518_, new_A2517_, new_A2516_,
    new_A2515_, new_A2514_, new_A2513_, new_A2512_, new_A2511_, new_A2510_,
    new_A2509_, new_A2508_, new_A2507_, new_A2506_, new_A2505_, new_A2504_,
    new_A2503_, new_A2502_, new_A2501_, new_A2500_, new_A2499_, new_A2498_,
    new_A2497_, new_A2496_, new_A2495_, new_A2494_, new_A2493_, new_A2492_,
    new_A2485_, new_A2484_, new_A2483_, new_A2482_, new_A2481_, new_A2480_,
    new_A2479_, new_A2478_, new_A2477_, new_A2476_, new_A2475_, new_A2474_,
    new_A2473_, new_A2472_, new_A2471_, new_A2470_, new_A2469_, new_A2468_,
    new_A2467_, new_A2466_, new_A2465_, new_A2464_, new_A2463_, new_A2462_,
    new_A2461_, new_A2460_, new_A2459_, new_A2458_, new_A2457_, new_A2456_,
    new_A2455_, new_A2454_, new_A2453_, new_A2452_, new_A2451_, new_A2450_,
    new_A2449_, new_A2448_, new_A2447_, new_A2446_, new_A2445_, new_A2444_,
    new_A2443_, new_A2442_, new_A2441_, new_A2440_, new_A2439_, new_A2438_,
    new_A2437_, new_A2436_, new_A2435_, new_A2434_, new_A2433_, new_A2432_,
    new_A2431_, new_A2430_, new_A2429_, new_A2428_, new_A2427_, new_A2426_,
    new_A2425_, new_A2418_, new_A2417_, new_A2416_, new_A2415_, new_A2414_,
    new_A2413_, new_A2412_, new_A2411_, new_A2410_, new_A2409_, new_A2408_,
    new_A2407_, new_A2406_, new_A2405_, new_A2404_, new_A2403_, new_A2402_,
    new_A2401_, new_A2400_, new_A2399_, new_A2398_, new_A2397_, new_A2396_,
    new_A2395_, new_A2394_, new_A2393_, new_A2392_, new_A2391_, new_A2390_,
    new_A2389_, new_A2388_, new_A2387_, new_A2386_, new_A2385_, new_A2384_,
    new_A2383_, new_A2382_, new_A2381_, new_A2380_, new_A2379_, new_A2378_,
    new_A2377_, new_A2376_, new_A2375_, new_A2374_, new_A2373_, new_A2372_,
    new_A2371_, new_A2370_, new_A2369_, new_A2368_, new_A2367_, new_A2366_,
    new_A2365_, new_A2364_, new_A2363_, new_A2362_, new_A2361_, new_A2360_,
    new_A2359_, new_A2358_, new_A2351_, new_A2350_, new_A2349_, new_A2348_,
    new_A2347_, new_A2346_, new_A2345_, new_A2344_, new_A2343_, new_A2342_,
    new_A2341_, new_A2340_, new_A2339_, new_A2338_, new_A2337_, new_A2336_,
    new_A2335_, new_A2334_, new_A2333_, new_A2332_, new_A2331_, new_A2330_,
    new_A2329_, new_A2328_, new_A2327_, new_A2326_, new_A2325_, new_A2324_,
    new_A2323_, new_A2322_, new_A2321_, new_A2320_, new_A2319_, new_A2318_,
    new_A2317_, new_A2316_, new_A2315_, new_A2314_, new_A2313_, new_A2312_,
    new_A2311_, new_A2310_, new_A2309_, new_A2308_, new_A2307_, new_A2306_,
    new_A2305_, new_A2304_, new_A2303_, new_A2302_, new_A2301_, new_A2300_,
    new_A2299_, new_A2298_, new_A2297_, new_A2296_, new_A2295_, new_A2294_,
    new_A2293_, new_A2292_, new_A2291_, new_A2284_, new_A2283_, new_A2282_,
    new_A2281_, new_A2280_, new_A2279_, new_A2278_, new_A2277_, new_A2276_,
    new_A2275_, new_A2274_, new_A2273_, new_A2272_, new_A2271_, new_A2270_,
    new_A2269_, new_A2268_, new_A2267_, new_A2266_, new_A2265_, new_A2264_,
    new_A2263_, new_A2262_, new_A2261_, new_A2260_, new_A2259_, new_A2258_,
    new_A2257_, new_A2256_, new_A2255_, new_A2254_, new_A2253_, new_A2252_,
    new_A2251_, new_A2250_, new_A2249_, new_A2248_, new_A2247_, new_A2246_,
    new_A2245_, new_A2244_, new_A2243_, new_A2242_, new_A2241_, new_A2240_,
    new_A2239_, new_A2238_, new_A2237_, new_A2236_, new_A2235_, new_A2234_,
    new_A2233_, new_A2232_, new_A2231_, new_A2230_, new_A2229_, new_A2228_,
    new_A2227_, new_A2226_, new_A2225_, new_A2224_, new_A2217_, new_A2216_,
    new_A2215_, new_A2214_, new_A2213_, new_A2212_, new_A2211_, new_A2210_,
    new_A2209_, new_A2208_, new_A2207_, new_A2206_, new_A2205_, new_A2204_,
    new_A2203_, new_A2202_, new_A2201_, new_A2200_, new_A2199_, new_A2198_,
    new_A2197_, new_A2196_, new_A2195_, new_A2194_, new_A2193_, new_A2192_,
    new_A2191_, new_A2190_, new_A2189_, new_A2188_, new_A2187_, new_A2186_,
    new_A2185_, new_A2184_, new_A2183_, new_A2182_, new_A2181_, new_A2180_,
    new_A2179_, new_A2178_, new_A2177_, new_A2176_, new_A2175_, new_A2174_,
    new_A2173_, new_A2172_, new_A2171_, new_A2170_, new_A2169_, new_A2168_,
    new_A2167_, new_A2166_, new_A2165_, new_A2164_, new_A2163_, new_A2162_,
    new_A2161_, new_A2160_, new_A2159_, new_A2158_, new_A2157_, new_A2150_,
    new_A2149_, new_A2148_, new_A2147_, new_A2146_, new_A2145_, new_A2144_,
    new_A2143_, new_A2142_, new_A2141_, new_A2140_, new_A2139_, new_A2138_,
    new_A2137_, new_A2136_, new_A2135_, new_A2134_, new_A2133_, new_A2132_,
    new_A2131_, new_A2130_, new_A2129_, new_A2128_, new_A2127_, new_A2126_,
    new_A2125_, new_A2124_, new_A2123_, new_A2122_, new_A2121_, new_A2120_,
    new_A2119_, new_A2118_, new_A2117_, new_A2116_, new_A2115_, new_A2114_,
    new_A2113_, new_A2112_, new_A2111_, new_A2110_, new_A2109_, new_A2108_,
    new_A2107_, new_A2106_, new_A2105_, new_A2104_, new_A2103_, new_A2102_,
    new_A2101_, new_A2100_, new_A2099_, new_A2098_, new_A2097_, new_A2096_,
    new_A2095_, new_A2094_, new_A2093_, new_A2092_, new_A2091_, new_A2090_,
    new_A2083_, new_A2082_, new_A2081_, new_A2080_, new_A2079_, new_A2078_,
    new_A2077_, new_A2076_, new_A2075_, new_A2074_, new_A2073_, new_A2072_,
    new_A2071_, new_A2070_, new_A2069_, new_A2068_, new_A2067_, new_A2066_,
    new_A2065_, new_A2064_, new_A2063_, new_A2062_, new_A2061_, new_A2060_,
    new_A2059_, new_A2058_, new_A2057_, new_A2056_, new_A2055_, new_A2054_,
    new_A2053_, new_A2052_, new_A2051_, new_A2050_, new_A2049_, new_A2048_,
    new_A2047_, new_A2046_, new_A2045_, new_A2044_, new_A2043_, new_A2042_,
    new_A2041_, new_A2040_, new_A2039_, new_A2038_, new_A2037_, new_A2036_,
    new_A2035_, new_A2034_, new_A2033_, new_A2032_, new_A2031_, new_A2030_,
    new_A2029_, new_A2028_, new_A2027_, new_A2026_, new_A2025_, new_A2024_,
    new_A2023_, new_A2016_, new_A2015_, new_A2014_, new_A2013_, new_A2012_,
    new_A2011_, new_A2010_, new_A2009_, new_A2008_, new_A2007_, new_A2006_,
    new_A2005_, new_A2004_, new_A2003_, new_A2002_, new_A2001_, new_A2000_,
    new_A1999_, new_A1998_, new_A1997_, new_A1996_, new_A1995_, new_A1994_,
    new_A1993_, new_A1992_, new_A1991_, new_A1990_, new_A1989_, new_A1988_,
    new_A1987_, new_A1986_, new_A1985_, new_A1984_, new_A1983_, new_A1982_,
    new_A1981_, new_A1980_, new_A1979_, new_A1978_, new_A1977_, new_A1976_,
    new_A1975_, new_A1974_, new_A1973_, new_A1972_, new_A1971_, new_A1970_,
    new_A1969_, new_A1968_, new_A1967_, new_A1966_, new_A1965_, new_A1964_,
    new_A1963_, new_A1962_, new_A1961_, new_A1960_, new_A1959_, new_A1958_,
    new_A1957_, new_A1956_, new_A1949_, new_A1948_, new_A1947_, new_A1946_,
    new_A1945_, new_A1944_, new_A1943_, new_A1942_, new_A1941_, new_A1940_,
    new_A1939_, new_A1938_, new_A1937_, new_A1936_, new_A1935_, new_A1934_,
    new_A1933_, new_A1932_, new_A1931_, new_A1930_, new_A1929_, new_A1928_,
    new_A1927_, new_A1926_, new_A1925_, new_A1924_, new_A1923_, new_A1922_,
    new_A1921_, new_A1920_, new_A1919_, new_A1918_, new_A1917_, new_A1916_,
    new_A1915_, new_A1914_, new_A1913_, new_A1912_, new_A1911_, new_A1910_,
    new_A1909_, new_A1908_, new_A1907_, new_A1906_, new_A1905_, new_A1904_,
    new_A1903_, new_A1902_, new_A1901_, new_A1900_, new_A1899_, new_A1898_,
    new_A1897_, new_A1896_, new_A1895_, new_A1894_, new_A1893_, new_A1892_,
    new_A1891_, new_A1890_, new_A1889_, new_A1882_, new_A1881_, new_A1880_,
    new_A1879_, new_A1878_, new_A1877_, new_A1876_, new_A1875_, new_A1874_,
    new_A1873_, new_A1872_, new_A1871_, new_A1870_, new_A1869_, new_A1868_,
    new_A1867_, new_A1866_, new_A1865_, new_A1864_, new_A1863_, new_A1862_,
    new_A1861_, new_A1860_, new_A1859_, new_A1858_, new_A1857_, new_A1856_,
    new_A1855_, new_A1854_, new_A1853_, new_A1852_, new_A1851_, new_A1850_,
    new_A1849_, new_A1848_, new_A1847_, new_A1846_, new_A1845_, new_A1844_,
    new_A1843_, new_A1842_, new_A1841_, new_A1840_, new_A1839_, new_A1838_,
    new_A1837_, new_A1836_, new_A1835_, new_A1834_, new_A1833_, new_A1832_,
    new_A1831_, new_A1830_, new_A1829_, new_A1828_, new_A1827_, new_A1826_,
    new_A1825_, new_A1824_, new_A1823_, new_A1822_, new_A1815_, new_A1814_,
    new_A1813_, new_A1812_, new_A1811_, new_A1810_, new_A1809_, new_A1808_,
    new_A1807_, new_A1806_, new_A1805_, new_A1804_, new_A1803_, new_A1802_,
    new_A1801_, new_A1800_, new_A1799_, new_A1798_, new_A1797_, new_A1796_,
    new_A1795_, new_A1794_, new_A1793_, new_A1792_, new_A1791_, new_A1790_,
    new_A1789_, new_A1788_, new_A1787_, new_A1786_, new_A1785_, new_A1784_,
    new_A1783_, new_A1782_, new_A1781_, new_A1780_, new_A1779_, new_A1778_,
    new_A1777_, new_A1776_, new_A1775_, new_A1774_, new_A1773_, new_A1772_,
    new_A1771_, new_A1770_, new_A1769_, new_A1768_, new_A1767_, new_A1766_,
    new_A1765_, new_A1764_, new_A1763_, new_A1762_, new_A1761_, new_A1760_,
    new_A1759_, new_A1758_, new_A1757_, new_A1756_, new_A1755_, new_A1748_,
    new_A1747_, new_A1746_, new_A1745_, new_A1744_, new_A1743_, new_A1742_,
    new_A1741_, new_A1740_, new_A1739_, new_A1738_, new_A1737_, new_A1736_,
    new_A1735_, new_A1734_, new_A1733_, new_A1732_, new_A1731_, new_A1730_,
    new_A1729_, new_A1728_, new_A1727_, new_A1726_, new_A1725_, new_A1724_,
    new_A1723_, new_A1722_, new_A1721_, new_A1720_, new_A1719_, new_A1718_,
    new_A1717_, new_A1716_, new_A1715_, new_A1714_, new_A1713_, new_A1712_,
    new_A1711_, new_A1710_, new_A1709_, new_A1708_, new_A1707_, new_A1706_,
    new_A1705_, new_A1704_, new_A1703_, new_A1702_, new_A1701_, new_A1700_,
    new_A1699_, new_A1698_, new_A1697_, new_A1696_, new_A1695_, new_A1694_,
    new_A1693_, new_A1692_, new_A1691_, new_A1690_, new_A1689_, new_A1688_,
    new_A1681_, new_A1680_, new_A1679_, new_A1678_, new_A1677_, new_A1676_,
    new_A1675_, new_A1674_, new_A1673_, new_A1672_, new_A1671_, new_A1670_,
    new_A1669_, new_A1668_, new_A1667_, new_A1666_, new_A1665_, new_A1664_,
    new_A1663_, new_A1662_, new_A1661_, new_A1660_, new_A1659_, new_A1658_,
    new_A1657_, new_A1656_, new_A1655_, new_A1654_, new_A1653_, new_A1652_,
    new_A1651_, new_A1650_, new_A1649_, new_A1648_, new_A1647_, new_A1646_,
    new_A1645_, new_A1644_, new_A1643_, new_A1642_, new_A1641_, new_A1640_,
    new_A1639_, new_A1638_, new_A1637_, new_A1636_, new_A1635_, new_A1634_,
    new_A1633_, new_A1632_, new_A1631_, new_A1630_, new_A1629_, new_A1628_,
    new_A1627_, new_A1626_, new_A1625_, new_A1624_, new_A1623_, new_A1622_,
    new_A1621_, new_A1614_, new_A1613_, new_A1612_, new_A1611_, new_A1610_,
    new_A1609_, new_A1608_, new_A1607_, new_A1606_, new_A1605_, new_A1604_,
    new_A1603_, new_A1602_, new_A1601_, new_A1600_, new_A1599_, new_A1598_,
    new_A1597_, new_A1596_, new_A1595_, new_A1594_, new_A1593_, new_A1592_,
    new_A1591_, new_A1590_, new_A1589_, new_A1588_, new_A1587_, new_A1586_,
    new_A1585_, new_A1584_, new_A1583_, new_A1582_, new_A1581_, new_A1580_,
    new_A1579_, new_A1578_, new_A1577_, new_A1576_, new_A1575_, new_A1574_,
    new_A1573_, new_A1572_, new_A1571_, new_A1570_, new_A1569_, new_A1568_,
    new_A1567_, new_A1566_, new_A1565_, new_A1564_, new_A1563_, new_A1562_,
    new_A1561_, new_A1560_, new_A1559_, new_A1558_, new_A1557_, new_A1556_,
    new_A1555_, new_A1554_, new_A1547_, new_A1546_, new_A1545_, new_A1544_,
    new_A1543_, new_A1542_, new_A1541_, new_A1540_, new_A1539_, new_A1538_,
    new_A1537_, new_A1536_, new_A1535_, new_A1534_, new_A1533_, new_A1532_,
    new_A1531_, new_A1530_, new_A1529_, new_A1528_, new_A1527_, new_A1526_,
    new_A1525_, new_A1524_, new_A1523_, new_A1522_, new_A1521_, new_A1520_,
    new_A1519_, new_A1518_, new_A1517_, new_A1516_, new_A1515_, new_A1514_,
    new_A1513_, new_A1512_, new_A1511_, new_A1510_, new_A1509_, new_A1508_,
    new_A1507_, new_A1506_, new_A1505_, new_A1504_, new_A1503_, new_A1502_,
    new_A1501_, new_A1500_, new_A1499_, new_A1498_, new_A1497_, new_A1496_,
    new_A1495_, new_A1494_, new_A1493_, new_A1492_, new_A1491_, new_A1490_,
    new_A1489_, new_A1488_, new_A1487_, new_A1480_, new_A1479_, new_A1478_,
    new_A1477_, new_A1476_, new_A1475_, new_A1474_, new_A1473_, new_A1472_,
    new_A1471_, new_A1470_, new_A1469_, new_A1468_, new_A1467_, new_A1466_,
    new_A1465_, new_A1464_, new_A1463_, new_A1462_, new_A1461_, new_A1460_,
    new_A1459_, new_A1458_, new_A1457_, new_A1456_, new_A1455_, new_A1454_,
    new_A1453_, new_A1452_, new_A1451_, new_A1450_, new_A1449_, new_A1448_,
    new_A1447_, new_A1446_, new_A1445_, new_A1444_, new_A1443_, new_A1442_,
    new_A1441_, new_A1440_, new_A1439_, new_A1438_, new_A1437_, new_A1436_,
    new_A1435_, new_A1434_, new_A1433_, new_A1432_, new_A1431_, new_A1430_,
    new_A1429_, new_A1428_, new_A1427_, new_A1426_, new_A1425_, new_A1424_,
    new_A1423_, new_A1422_, new_A1421_, new_A1420_, new_A1413_, new_A1412_,
    new_A1411_, new_A1410_, new_A1409_, new_A1408_, new_A1407_, new_A1406_,
    new_A1405_, new_A1404_, new_A1403_, new_A1402_, new_A1401_, new_A1400_,
    new_A1399_, new_A1398_, new_A1397_, new_A1396_, new_A1395_, new_A1394_,
    new_A1393_, new_A1392_, new_A1391_, new_A1390_, new_A1389_, new_A1388_,
    new_A1387_, new_A1386_, new_A1385_, new_A1384_, new_A1383_, new_A1382_,
    new_A1381_, new_A1380_, new_A1379_, new_A1378_, new_A1377_, new_A1376_,
    new_A1375_, new_A1374_, new_A1373_, new_A1372_, new_A1371_, new_A1370_,
    new_A1369_, new_A1368_, new_A1367_, new_A1366_, new_A1365_, new_A1364_,
    new_A1363_, new_A1362_, new_A1361_, new_A1360_, new_A1359_, new_A1358_,
    new_A1357_, new_A1356_, new_A1355_, new_A1354_, new_A1353_, new_A1346_,
    new_A1345_, new_A1344_, new_A1343_, new_A1342_, new_A1341_, new_A1340_,
    new_A1339_, new_A1338_, new_A1337_, new_A1336_, new_A1335_, new_A1334_,
    new_A1333_, new_A1332_, new_A1331_, new_A1330_, new_A1329_, new_A1328_,
    new_A1327_, new_A1326_, new_A1325_, new_A1324_, new_A1323_, new_A1322_,
    new_A1321_, new_A1320_, new_A1319_, new_A1318_, new_A1317_, new_A1316_,
    new_A1315_, new_A1314_, new_A1313_, new_A1312_, new_A1311_, new_A1310_,
    new_A1309_, new_A1308_, new_A1307_, new_A1306_, new_A1305_, new_A1304_,
    new_A1303_, new_A1302_, new_A1301_, new_A1300_, new_A1299_, new_A1298_,
    new_A1297_, new_A1296_, new_A1295_, new_A1294_, new_A1293_, new_A1292_,
    new_A1291_, new_A1290_, new_A1289_, new_A1288_, new_A1287_, new_A1286_,
    new_A1279_, new_A1278_, new_A1277_, new_A1276_, new_A1275_, new_A1274_,
    new_A1273_, new_A1272_, new_A1271_, new_A1270_, new_A1269_, new_A1268_,
    new_A1267_, new_A1266_, new_A1265_, new_A1264_, new_A1263_, new_A1262_,
    new_A1261_, new_A1260_, new_A1259_, new_A1258_, new_A1257_, new_A1256_,
    new_A1255_, new_A1254_, new_A1253_, new_A1252_, new_A1251_, new_A1250_,
    new_A1249_, new_A1248_, new_A1247_, new_A1246_, new_A1245_, new_A1244_,
    new_A1243_, new_A1242_, new_A1241_, new_A1240_, new_A1239_, new_A1238_,
    new_A1237_, new_A1236_, new_A1235_, new_A1234_, new_A1233_, new_A1232_,
    new_A1231_, new_A1230_, new_A1229_, new_A1228_, new_A1227_, new_A1226_,
    new_A1225_, new_A1224_, new_A1223_, new_A1222_, new_A1221_, new_A1220_,
    new_A1219_, new_A1212_, new_A1211_, new_A1210_, new_A1209_, new_A1208_,
    new_A1207_, new_A1206_, new_A1205_, new_A1204_, new_A1203_, new_A1202_,
    new_A1201_, new_A1200_, new_A1199_, new_A1198_, new_A1197_, new_A1196_,
    new_A1195_, new_A1194_, new_A1193_, new_A1192_, new_A1191_, new_A1190_,
    new_A1189_, new_A1188_, new_A1187_, new_A1186_, new_A1185_, new_A1184_,
    new_A1183_, new_A1182_, new_A1181_, new_A1180_, new_A1179_, new_A1178_,
    new_A1177_, new_A1176_, new_A1175_, new_A1174_, new_A1173_, new_A1172_,
    new_A1171_, new_A1170_, new_A1169_, new_A1168_, new_A1167_, new_A1166_,
    new_A1165_, new_A1164_, new_A1163_, new_A1162_, new_A1161_, new_A1160_,
    new_A1159_, new_A1158_, new_A1157_, new_A1156_, new_A1155_, new_A1154_,
    new_A1153_, new_A1152_, new_A1145_, new_A1144_, new_A1143_, new_A1142_,
    new_A1141_, new_A1140_, new_A1139_, new_A1138_, new_A1137_, new_A1136_,
    new_A1135_, new_A1134_, new_A1133_, new_A1132_, new_A1131_, new_A1130_,
    new_A1129_, new_A1128_, new_A1127_, new_A1126_, new_A1125_, new_A1124_,
    new_A1123_, new_A1122_, new_A1121_, new_A1120_, new_A1119_, new_A1118_,
    new_A1117_, new_A1116_, new_A1115_, new_A1114_, new_A1113_, new_A1112_,
    new_A1111_, new_A1110_, new_A1109_, new_A1108_, new_A1107_, new_A1106_,
    new_A1105_, new_A1104_, new_A1103_, new_A1102_, new_A1101_, new_A1100_,
    new_A1099_, new_A1098_, new_A1097_, new_A1096_, new_A1095_, new_A1094_,
    new_A1093_, new_A1092_, new_A1091_, new_A1090_, new_A1089_, new_A1088_,
    new_A1087_, new_A1086_, new_A1085_, new_A1078_, new_A1077_, new_A1076_,
    new_A1075_, new_A1074_, new_A1073_, new_A1072_, new_A1071_, new_A1070_,
    new_A1069_, new_A1068_, new_A1067_, new_A1066_, new_A1065_, new_A1064_,
    new_A1063_, new_A1062_, new_A1061_, new_A1060_, new_A1059_, new_A1058_,
    new_A1057_, new_A1056_, new_A1055_, new_A1054_, new_A1053_, new_A1052_,
    new_A1051_, new_A1050_, new_A1049_, new_A1048_, new_A1047_, new_A1046_,
    new_A1045_, new_A1044_, new_A1043_, new_A1042_, new_A1041_, new_A1040_,
    new_A1039_, new_A1038_, new_A1037_, new_A1036_, new_A1035_, new_A1034_,
    new_A1033_, new_A1032_, new_A1031_, new_A1030_, new_A1029_, new_A1028_,
    new_A1027_, new_A1026_, new_A1025_, new_A1024_, new_A1023_, new_A1022_,
    new_A1021_, new_A1020_, new_A1019_, new_A1018_, new_A1011_, new_A1010_,
    new_A1009_, new_A1008_, new_A1007_, new_A1006_, new_A1005_, new_A1004_,
    new_A1003_, new_A1002_, new_A1001_, new_A1000_, new_A999_, new_A998_,
    new_A997_, new_A996_, new_A995_, new_A994_, new_A993_, new_A992_,
    new_A991_, new_A990_, new_A989_, new_A988_, new_A987_, new_A986_,
    new_A985_, new_A984_, new_A983_, new_A982_, new_A981_, new_A980_,
    new_A979_, new_A978_, new_A977_, new_A976_, new_A975_, new_A974_,
    new_A973_, new_A972_, new_A971_, new_A970_, new_A969_, new_A968_,
    new_A967_, new_A966_, new_A965_, new_A964_, new_A963_, new_A962_,
    new_A961_, new_A960_, new_A959_, new_A958_, new_A957_, new_A956_,
    new_A955_, new_A954_, new_A953_, new_A952_, new_A951_, new_A944_,
    new_A943_, new_A942_, new_A941_, new_A940_, new_A939_, new_A938_,
    new_A937_, new_A936_, new_A935_, new_A934_, new_A933_, new_A932_,
    new_A931_, new_A930_, new_A929_, new_A928_, new_A927_, new_A926_,
    new_A925_, new_A924_, new_A923_, new_A922_, new_A921_, new_A920_,
    new_A919_, new_A918_, new_A917_, new_A916_, new_A915_, new_A914_,
    new_A913_, new_A912_, new_A911_, new_A910_, new_A909_, new_A908_,
    new_A907_, new_A906_, new_A905_, new_A904_, new_A903_, new_A902_,
    new_A901_, new_A900_, new_A899_, new_A898_, new_A897_, new_A896_,
    new_A895_, new_A894_, new_A893_, new_A892_, new_A891_, new_A890_,
    new_A889_, new_A888_, new_A887_, new_A886_, new_A885_, new_A884_,
    new_A877_, new_A876_, new_A875_, new_A874_, new_A873_, new_A872_,
    new_A805_, new_A806_, new_A807_, new_A808_, new_A809_, new_A810_,
    new_A817_, new_A818_, new_A819_, new_A820_, new_A821_, new_A822_,
    new_A823_, new_A824_, new_A825_, new_A826_, new_A827_, new_A828_,
    new_A829_, new_A830_, new_A831_, new_A832_, new_A833_, new_A834_,
    new_A835_, new_A836_, new_A837_, new_A838_, new_A839_, new_A840_,
    new_A841_, new_A842_, new_A843_, new_A844_, new_A845_, new_A846_,
    new_A847_, new_A848_, new_A849_, new_A850_, new_A851_, new_A852_,
    new_A853_, new_A854_, new_A855_, new_A856_, new_A857_, new_A858_,
    new_A859_, new_A860_, new_A861_, new_A862_, new_A863_, new_A864_,
    new_A865_, new_A866_, new_A867_, new_A868_, new_A869_, new_A870_,
    new_A871_;
  assign new_A5695_ = ~A5634 & new_A5648_;
  assign new_A5694_ = A5634 & ~new_A5648_;
  assign new_A5693_ = A5634 & ~new_A5648_;
  assign new_A5692_ = ~A5634 & ~new_A5648_;
  assign new_A5691_ = A5634 & new_A5648_;
  assign new_A5690_ = new_A5694_ | new_A5695_;
  assign new_A5689_ = ~A5634 & new_A5648_;
  assign new_A5688_ = new_A5692_ | new_A5693_;
  assign new_A5687_ = ~new_A5663_ & ~new_A5683_;
  assign new_A5686_ = new_A5663_ & new_A5683_;
  assign new_A5685_ = ~A5630 | ~new_A5655_;
  assign new_A5684_ = new_A5648_ & new_A5685_;
  assign new_A5683_ = A5631 | A5632;
  assign new_A5682_ = A5631 | new_A5648_;
  assign new_A5681_ = ~new_A5648_ & ~new_A5684_;
  assign new_A5680_ = new_A5648_ | new_A5685_;
  assign new_A5679_ = A5631 & ~A5632;
  assign new_A5678_ = ~A5631 & A5632;
  assign new_A5677_ = new_A5641_ | new_A5674_;
  assign new_A5676_ = ~new_A5641_ & ~new_A5675_;
  assign new_A5675_ = new_A5641_ & new_A5674_;
  assign new_A5674_ = ~A5630 | ~new_A5655_;
  assign new_A5673_ = ~A5631 & new_A5641_;
  assign new_A5672_ = A5631 & ~new_A5641_;
  assign new_A5671_ = A5633 & new_A5670_;
  assign new_A5670_ = new_A5689_ | new_A5688_;
  assign new_A5669_ = ~A5633 & new_A5668_;
  assign new_A5668_ = new_A5691_ | new_A5690_;
  assign new_A5667_ = A5633 | new_A5666_;
  assign new_A5666_ = new_A5687_ | new_A5686_;
  assign new_A5665_ = ~new_A5645_ & ~new_A5655_;
  assign new_A5664_ = new_A5645_ & new_A5655_;
  assign new_A5663_ = ~new_A5645_ | new_A5655_;
  assign new_A5662_ = A5629 & ~A5630;
  assign new_A5661_ = ~A5629 & A5630;
  assign new_A5660_ = new_A5682_ & ~new_A5683_;
  assign new_A5659_ = ~new_A5682_ & new_A5683_;
  assign new_A5658_ = ~new_A5681_ | ~new_A5680_;
  assign new_A5657_ = new_A5673_ | new_A5672_;
  assign new_A5656_ = new_A5679_ | new_A5678_;
  assign new_A5655_ = new_A5669_ | new_A5671_;
  assign new_A5654_ = ~new_A5676_ | ~new_A5677_;
  assign new_A5653_ = A5629 & ~A5630;
  assign new_A5652_ = new_A5643_ & ~new_A5655_;
  assign new_A5651_ = ~new_A5643_ & new_A5655_;
  assign new_A5650_ = ~new_A5641_ & new_A5667_;
  assign new_A5649_ = new_A5665_ | new_A5664_;
  assign new_A5648_ = new_A5662_ | new_A5661_;
  assign new_A5647_ = A5630 | new_A5663_;
  assign new_A5646_ = new_A5655_ & new_A5658_;
  assign new_A5645_ = new_A5660_ | new_A5659_;
  assign new_A5644_ = new_A5655_ & new_A5654_;
  assign new_A5643_ = new_A5657_ & new_A5656_;
  assign new_A5642_ = new_A5652_ | new_A5651_;
  assign new_A5641_ = A5630 | new_A5653_;
  assign new_A5640_ = new_A5641_ | new_A5650_;
  assign new_A5639_ = new_A5648_ & new_A5649_;
  assign new_A5638_ = new_A5648_ & new_A5647_;
  assign new_A5637_ = new_A5646_ | new_A5645_;
  assign new_A5636_ = new_A5644_ | new_A5643_;
  assign new_A5635_ = new_A5642_ & new_A5641_;
  assign new_A5702_ = new_A5709_ & new_A5708_;
  assign new_A5703_ = new_A5711_ | new_A5710_;
  assign new_A5704_ = new_A5713_ | new_A5712_;
  assign new_A5705_ = new_A5715_ & new_A5714_;
  assign new_A5706_ = new_A5715_ & new_A5716_;
  assign new_A5707_ = new_A5708_ | new_A5717_;
  assign new_A5708_ = A5697 | new_A5720_;
  assign new_A5709_ = new_A5719_ | new_A5718_;
  assign new_A5710_ = new_A5724_ & new_A5723_;
  assign new_A5711_ = new_A5722_ & new_A5721_;
  assign new_A5712_ = new_A5727_ | new_A5726_;
  assign new_A5713_ = new_A5722_ & new_A5725_;
  assign new_A5714_ = A5697 | new_A5730_;
  assign new_A5715_ = new_A5729_ | new_A5728_;
  assign new_A5716_ = new_A5732_ | new_A5731_;
  assign new_A5717_ = ~new_A5708_ & new_A5734_;
  assign new_A5718_ = ~new_A5710_ & new_A5722_;
  assign new_A5719_ = new_A5710_ & ~new_A5722_;
  assign new_A5720_ = A5696 & ~A5697;
  assign new_A5721_ = ~new_A5743_ | ~new_A5744_;
  assign new_A5722_ = new_A5736_ | new_A5738_;
  assign new_A5723_ = new_A5746_ | new_A5745_;
  assign new_A5724_ = new_A5740_ | new_A5739_;
  assign new_A5725_ = ~new_A5748_ | ~new_A5747_;
  assign new_A5726_ = ~new_A5749_ & new_A5750_;
  assign new_A5727_ = new_A5749_ & ~new_A5750_;
  assign new_A5728_ = ~A5696 & A5697;
  assign new_A5729_ = A5696 & ~A5697;
  assign new_A5730_ = ~new_A5712_ | new_A5722_;
  assign new_A5731_ = new_A5712_ & new_A5722_;
  assign new_A5732_ = ~new_A5712_ & ~new_A5722_;
  assign new_A5733_ = new_A5754_ | new_A5753_;
  assign new_A5734_ = A5700 | new_A5733_;
  assign new_A5735_ = new_A5758_ | new_A5757_;
  assign new_A5736_ = ~A5700 & new_A5735_;
  assign new_A5737_ = new_A5756_ | new_A5755_;
  assign new_A5738_ = A5700 & new_A5737_;
  assign new_A5739_ = A5698 & ~new_A5708_;
  assign new_A5740_ = ~A5698 & new_A5708_;
  assign new_A5741_ = ~A5697 | ~new_A5722_;
  assign new_A5742_ = new_A5708_ & new_A5741_;
  assign new_A5743_ = ~new_A5708_ & ~new_A5742_;
  assign new_A5744_ = new_A5708_ | new_A5741_;
  assign new_A5745_ = ~A5698 & A5699;
  assign new_A5746_ = A5698 & ~A5699;
  assign new_A5747_ = new_A5715_ | new_A5752_;
  assign new_A5748_ = ~new_A5715_ & ~new_A5751_;
  assign new_A5749_ = A5698 | new_A5715_;
  assign new_A5750_ = A5698 | A5699;
  assign new_A5751_ = new_A5715_ & new_A5752_;
  assign new_A5752_ = ~A5697 | ~new_A5722_;
  assign new_A5753_ = new_A5730_ & new_A5750_;
  assign new_A5754_ = ~new_A5730_ & ~new_A5750_;
  assign new_A5755_ = new_A5759_ | new_A5760_;
  assign new_A5756_ = ~A5701 & new_A5715_;
  assign new_A5757_ = new_A5761_ | new_A5762_;
  assign new_A5758_ = A5701 & new_A5715_;
  assign new_A5759_ = ~A5701 & ~new_A5715_;
  assign new_A5760_ = A5701 & ~new_A5715_;
  assign new_A5761_ = A5701 & ~new_A5715_;
  assign new_A5762_ = ~A5701 & new_A5715_;
  assign new_A5769_ = new_A5776_ & new_A5775_;
  assign new_A5770_ = new_A5778_ | new_A5777_;
  assign new_A5771_ = new_A5780_ | new_A5779_;
  assign new_A5772_ = new_A5782_ & new_A5781_;
  assign new_A5773_ = new_A5782_ & new_A5783_;
  assign new_A5774_ = new_A5775_ | new_A5784_;
  assign new_A5775_ = A5764 | new_A5787_;
  assign new_A5776_ = new_A5786_ | new_A5785_;
  assign new_A5777_ = new_A5791_ & new_A5790_;
  assign new_A5778_ = new_A5789_ & new_A5788_;
  assign new_A5779_ = new_A5794_ | new_A5793_;
  assign new_A5780_ = new_A5789_ & new_A5792_;
  assign new_A5781_ = A5764 | new_A5797_;
  assign new_A5782_ = new_A5796_ | new_A5795_;
  assign new_A5783_ = new_A5799_ | new_A5798_;
  assign new_A5784_ = ~new_A5775_ & new_A5801_;
  assign new_A5785_ = ~new_A5777_ & new_A5789_;
  assign new_A5786_ = new_A5777_ & ~new_A5789_;
  assign new_A5787_ = A5763 & ~A5764;
  assign new_A5788_ = ~new_A5810_ | ~new_A5811_;
  assign new_A5789_ = new_A5803_ | new_A5805_;
  assign new_A5790_ = new_A5813_ | new_A5812_;
  assign new_A5791_ = new_A5807_ | new_A5806_;
  assign new_A5792_ = ~new_A5815_ | ~new_A5814_;
  assign new_A5793_ = ~new_A5816_ & new_A5817_;
  assign new_A5794_ = new_A5816_ & ~new_A5817_;
  assign new_A5795_ = ~A5763 & A5764;
  assign new_A5796_ = A5763 & ~A5764;
  assign new_A5797_ = ~new_A5779_ | new_A5789_;
  assign new_A5798_ = new_A5779_ & new_A5789_;
  assign new_A5799_ = ~new_A5779_ & ~new_A5789_;
  assign new_A5800_ = new_A5821_ | new_A5820_;
  assign new_A5801_ = A5767 | new_A5800_;
  assign new_A5802_ = new_A5825_ | new_A5824_;
  assign new_A5803_ = ~A5767 & new_A5802_;
  assign new_A5804_ = new_A5823_ | new_A5822_;
  assign new_A5805_ = A5767 & new_A5804_;
  assign new_A5806_ = A5765 & ~new_A5775_;
  assign new_A5807_ = ~A5765 & new_A5775_;
  assign new_A5808_ = ~A5764 | ~new_A5789_;
  assign new_A5809_ = new_A5775_ & new_A5808_;
  assign new_A5810_ = ~new_A5775_ & ~new_A5809_;
  assign new_A5811_ = new_A5775_ | new_A5808_;
  assign new_A5812_ = ~A5765 & A5766;
  assign new_A5813_ = A5765 & ~A5766;
  assign new_A5814_ = new_A5782_ | new_A5819_;
  assign new_A5815_ = ~new_A5782_ & ~new_A5818_;
  assign new_A5816_ = A5765 | new_A5782_;
  assign new_A5817_ = A5765 | A5766;
  assign new_A5818_ = new_A5782_ & new_A5819_;
  assign new_A5819_ = ~A5764 | ~new_A5789_;
  assign new_A5820_ = new_A5797_ & new_A5817_;
  assign new_A5821_ = ~new_A5797_ & ~new_A5817_;
  assign new_A5822_ = new_A5826_ | new_A5827_;
  assign new_A5823_ = ~A5768 & new_A5782_;
  assign new_A5824_ = new_A5828_ | new_A5829_;
  assign new_A5825_ = A5768 & new_A5782_;
  assign new_A5826_ = ~A5768 & ~new_A5782_;
  assign new_A5827_ = A5768 & ~new_A5782_;
  assign new_A5828_ = A5768 & ~new_A5782_;
  assign new_A5829_ = ~A5768 & new_A5782_;
  assign new_A5836_ = new_A5843_ & new_A5842_;
  assign new_A5837_ = new_A5845_ | new_A5844_;
  assign new_A5838_ = new_A5847_ | new_A5846_;
  assign new_A5839_ = new_A5849_ & new_A5848_;
  assign new_A5840_ = new_A5849_ & new_A5850_;
  assign new_A5841_ = new_A5842_ | new_A5851_;
  assign new_A5842_ = A5831 | new_A5854_;
  assign new_A5843_ = new_A5853_ | new_A5852_;
  assign new_A5844_ = new_A5858_ & new_A5857_;
  assign new_A5845_ = new_A5856_ & new_A5855_;
  assign new_A5846_ = new_A5861_ | new_A5860_;
  assign new_A5847_ = new_A5856_ & new_A5859_;
  assign new_A5848_ = A5831 | new_A5864_;
  assign new_A5849_ = new_A5863_ | new_A5862_;
  assign new_A5850_ = new_A5866_ | new_A5865_;
  assign new_A5851_ = ~new_A5842_ & new_A5868_;
  assign new_A5852_ = ~new_A5844_ & new_A5856_;
  assign new_A5853_ = new_A5844_ & ~new_A5856_;
  assign new_A5854_ = A5830 & ~A5831;
  assign new_A5855_ = ~new_A5877_ | ~new_A5878_;
  assign new_A5856_ = new_A5870_ | new_A5872_;
  assign new_A5857_ = new_A5880_ | new_A5879_;
  assign new_A5858_ = new_A5874_ | new_A5873_;
  assign new_A5859_ = ~new_A5882_ | ~new_A5881_;
  assign new_A5860_ = ~new_A5883_ & new_A5884_;
  assign new_A5861_ = new_A5883_ & ~new_A5884_;
  assign new_A5862_ = ~A5830 & A5831;
  assign new_A5863_ = A5830 & ~A5831;
  assign new_A5864_ = ~new_A5846_ | new_A5856_;
  assign new_A5865_ = new_A5846_ & new_A5856_;
  assign new_A5866_ = ~new_A5846_ & ~new_A5856_;
  assign new_A5867_ = new_A5888_ | new_A5887_;
  assign new_A5868_ = A5834 | new_A5867_;
  assign new_A5869_ = new_A5892_ | new_A5891_;
  assign new_A5870_ = ~A5834 & new_A5869_;
  assign new_A5871_ = new_A5890_ | new_A5889_;
  assign new_A5872_ = A5834 & new_A5871_;
  assign new_A5873_ = A5832 & ~new_A5842_;
  assign new_A5874_ = ~A5832 & new_A5842_;
  assign new_A5875_ = ~A5831 | ~new_A5856_;
  assign new_A5876_ = new_A5842_ & new_A5875_;
  assign new_A5877_ = ~new_A5842_ & ~new_A5876_;
  assign new_A5878_ = new_A5842_ | new_A5875_;
  assign new_A5879_ = ~A5832 & A5833;
  assign new_A5880_ = A5832 & ~A5833;
  assign new_A5881_ = new_A5849_ | new_A5886_;
  assign new_A5882_ = ~new_A5849_ & ~new_A5885_;
  assign new_A5883_ = A5832 | new_A5849_;
  assign new_A5884_ = A5832 | A5833;
  assign new_A5885_ = new_A5849_ & new_A5886_;
  assign new_A5886_ = ~A5831 | ~new_A5856_;
  assign new_A5887_ = new_A5864_ & new_A5884_;
  assign new_A5888_ = ~new_A5864_ & ~new_A5884_;
  assign new_A5889_ = new_A5893_ | new_A5894_;
  assign new_A5890_ = ~A5835 & new_A5849_;
  assign new_A5891_ = new_A5895_ | new_A5896_;
  assign new_A5892_ = A5835 & new_A5849_;
  assign new_A5893_ = ~A5835 & ~new_A5849_;
  assign new_A5894_ = A5835 & ~new_A5849_;
  assign new_A5895_ = A5835 & ~new_A5849_;
  assign new_A5896_ = ~A5835 & new_A5849_;
  assign new_A5903_ = new_A5910_ & new_A5909_;
  assign new_A5904_ = new_A5912_ | new_A5911_;
  assign new_A5905_ = new_A5914_ | new_A5913_;
  assign new_A5906_ = new_A5916_ & new_A5915_;
  assign new_A5907_ = new_A5916_ & new_A5917_;
  assign new_A5908_ = new_A5909_ | new_A5918_;
  assign new_A5909_ = A5898 | new_A5921_;
  assign new_A5910_ = new_A5920_ | new_A5919_;
  assign new_A5911_ = new_A5925_ & new_A5924_;
  assign new_A5912_ = new_A5923_ & new_A5922_;
  assign new_A5913_ = new_A5928_ | new_A5927_;
  assign new_A5914_ = new_A5923_ & new_A5926_;
  assign new_A5915_ = A5898 | new_A5931_;
  assign new_A5916_ = new_A5930_ | new_A5929_;
  assign new_A5917_ = new_A5933_ | new_A5932_;
  assign new_A5918_ = ~new_A5909_ & new_A5935_;
  assign new_A5919_ = ~new_A5911_ & new_A5923_;
  assign new_A5920_ = new_A5911_ & ~new_A5923_;
  assign new_A5921_ = A5897 & ~A5898;
  assign new_A5922_ = ~new_A5944_ | ~new_A5945_;
  assign new_A5923_ = new_A5937_ | new_A5939_;
  assign new_A5924_ = new_A5947_ | new_A5946_;
  assign new_A5925_ = new_A5941_ | new_A5940_;
  assign new_A5926_ = ~new_A5949_ | ~new_A5948_;
  assign new_A5927_ = ~new_A5950_ & new_A5951_;
  assign new_A5928_ = new_A5950_ & ~new_A5951_;
  assign new_A5929_ = ~A5897 & A5898;
  assign new_A5930_ = A5897 & ~A5898;
  assign new_A5931_ = ~new_A5913_ | new_A5923_;
  assign new_A5932_ = new_A5913_ & new_A5923_;
  assign new_A5933_ = ~new_A5913_ & ~new_A5923_;
  assign new_A5934_ = new_A5955_ | new_A5954_;
  assign new_A5935_ = A5901 | new_A5934_;
  assign new_A5936_ = new_A5959_ | new_A5958_;
  assign new_A5937_ = ~A5901 & new_A5936_;
  assign new_A5938_ = new_A5957_ | new_A5956_;
  assign new_A5939_ = A5901 & new_A5938_;
  assign new_A5940_ = A5899 & ~new_A5909_;
  assign new_A5941_ = ~A5899 & new_A5909_;
  assign new_A5942_ = ~A5898 | ~new_A5923_;
  assign new_A5943_ = new_A5909_ & new_A5942_;
  assign new_A5944_ = ~new_A5909_ & ~new_A5943_;
  assign new_A5945_ = new_A5909_ | new_A5942_;
  assign new_A5946_ = ~A5899 & A5900;
  assign new_A5947_ = A5899 & ~A5900;
  assign new_A5948_ = new_A5916_ | new_A5953_;
  assign new_A5949_ = ~new_A5916_ & ~new_A5952_;
  assign new_A5950_ = A5899 | new_A5916_;
  assign new_A5951_ = A5899 | A5900;
  assign new_A5952_ = new_A5916_ & new_A5953_;
  assign new_A5953_ = ~A5898 | ~new_A5923_;
  assign new_A5954_ = new_A5931_ & new_A5951_;
  assign new_A5955_ = ~new_A5931_ & ~new_A5951_;
  assign new_A5956_ = new_A5960_ | new_A5961_;
  assign new_A5957_ = ~A5902 & new_A5916_;
  assign new_A5958_ = new_A5962_ | new_A5963_;
  assign new_A5959_ = A5902 & new_A5916_;
  assign new_A5960_ = ~A5902 & ~new_A5916_;
  assign new_A5961_ = A5902 & ~new_A5916_;
  assign new_A5962_ = A5902 & ~new_A5916_;
  assign new_A5963_ = ~A5902 & new_A5916_;
  assign new_A5970_ = new_A5977_ & new_A5976_;
  assign new_A5971_ = new_A5979_ | new_A5978_;
  assign new_A5972_ = new_A5981_ | new_A5980_;
  assign new_A5973_ = new_A5983_ & new_A5982_;
  assign new_A5974_ = new_A5983_ & new_A5984_;
  assign new_A5975_ = new_A5976_ | new_A5985_;
  assign new_A5976_ = A5965 | new_A5988_;
  assign new_A5977_ = new_A5987_ | new_A5986_;
  assign new_A5978_ = new_A5992_ & new_A5991_;
  assign new_A5979_ = new_A5990_ & new_A5989_;
  assign new_A5980_ = new_A5995_ | new_A5994_;
  assign new_A5981_ = new_A5990_ & new_A5993_;
  assign new_A5982_ = A5965 | new_A5998_;
  assign new_A5983_ = new_A5997_ | new_A5996_;
  assign new_A5984_ = new_A6000_ | new_A5999_;
  assign new_A5985_ = ~new_A5976_ & new_A6002_;
  assign new_A5986_ = ~new_A5978_ & new_A5990_;
  assign new_A5987_ = new_A5978_ & ~new_A5990_;
  assign new_A5988_ = A5964 & ~A5965;
  assign new_A5989_ = ~new_A6011_ | ~new_A6012_;
  assign new_A5990_ = new_A6004_ | new_A6006_;
  assign new_A5991_ = new_A6014_ | new_A6013_;
  assign new_A5992_ = new_A6008_ | new_A6007_;
  assign new_A5993_ = ~new_A6016_ | ~new_A6015_;
  assign new_A5994_ = ~new_A6017_ & new_A6018_;
  assign new_A5995_ = new_A6017_ & ~new_A6018_;
  assign new_A5996_ = ~A5964 & A5965;
  assign new_A5997_ = A5964 & ~A5965;
  assign new_A5998_ = ~new_A5980_ | new_A5990_;
  assign new_A5999_ = new_A5980_ & new_A5990_;
  assign new_A6000_ = ~new_A5980_ & ~new_A5990_;
  assign new_A6001_ = new_A6022_ | new_A6021_;
  assign new_A6002_ = A5968 | new_A6001_;
  assign new_A6003_ = new_A6026_ | new_A6025_;
  assign new_A6004_ = ~A5968 & new_A6003_;
  assign new_A6005_ = new_A6024_ | new_A6023_;
  assign new_A6006_ = A5968 & new_A6005_;
  assign new_A6007_ = A5966 & ~new_A5976_;
  assign new_A6008_ = ~A5966 & new_A5976_;
  assign new_A6009_ = ~A5965 | ~new_A5990_;
  assign new_A6010_ = new_A5976_ & new_A6009_;
  assign new_A6011_ = ~new_A5976_ & ~new_A6010_;
  assign new_A6012_ = new_A5976_ | new_A6009_;
  assign new_A6013_ = ~A5966 & A5967;
  assign new_A6014_ = A5966 & ~A5967;
  assign new_A6015_ = new_A5983_ | new_A6020_;
  assign new_A6016_ = ~new_A5983_ & ~new_A6019_;
  assign new_A6017_ = A5966 | new_A5983_;
  assign new_A6018_ = A5966 | A5967;
  assign new_A6019_ = new_A5983_ & new_A6020_;
  assign new_A6020_ = ~A5965 | ~new_A5990_;
  assign new_A6021_ = new_A5998_ & new_A6018_;
  assign new_A6022_ = ~new_A5998_ & ~new_A6018_;
  assign new_A6023_ = new_A6027_ | new_A6028_;
  assign new_A6024_ = ~A5969 & new_A5983_;
  assign new_A6025_ = new_A6029_ | new_A6030_;
  assign new_A6026_ = A5969 & new_A5983_;
  assign new_A6027_ = ~A5969 & ~new_A5983_;
  assign new_A6028_ = A5969 & ~new_A5983_;
  assign new_A6029_ = A5969 & ~new_A5983_;
  assign new_A6030_ = ~A5969 & new_A5983_;
  assign new_A6037_ = new_A6044_ & new_A6043_;
  assign new_A6038_ = new_A6046_ | new_A6045_;
  assign new_A6039_ = new_A6048_ | new_A6047_;
  assign new_A6040_ = new_A6050_ & new_A6049_;
  assign new_A6041_ = new_A6050_ & new_A6051_;
  assign new_A6042_ = new_A6043_ | new_A6052_;
  assign new_A6043_ = A6032 | new_A6055_;
  assign new_A6044_ = new_A6054_ | new_A6053_;
  assign new_A6045_ = new_A6059_ & new_A6058_;
  assign new_A6046_ = new_A6057_ & new_A6056_;
  assign new_A6047_ = new_A6062_ | new_A6061_;
  assign new_A6048_ = new_A6057_ & new_A6060_;
  assign new_A6049_ = A6032 | new_A6065_;
  assign new_A6050_ = new_A6064_ | new_A6063_;
  assign new_A6051_ = new_A6067_ | new_A6066_;
  assign new_A6052_ = ~new_A6043_ & new_A6069_;
  assign new_A6053_ = ~new_A6045_ & new_A6057_;
  assign new_A6054_ = new_A6045_ & ~new_A6057_;
  assign new_A6055_ = A6031 & ~A6032;
  assign new_A6056_ = ~new_A6078_ | ~new_A6079_;
  assign new_A6057_ = new_A6071_ | new_A6073_;
  assign new_A6058_ = new_A6081_ | new_A6080_;
  assign new_A6059_ = new_A6075_ | new_A6074_;
  assign new_A6060_ = ~new_A6083_ | ~new_A6082_;
  assign new_A6061_ = ~new_A6084_ & new_A6085_;
  assign new_A6062_ = new_A6084_ & ~new_A6085_;
  assign new_A6063_ = ~A6031 & A6032;
  assign new_A6064_ = A6031 & ~A6032;
  assign new_A6065_ = ~new_A6047_ | new_A6057_;
  assign new_A6066_ = new_A6047_ & new_A6057_;
  assign new_A6067_ = ~new_A6047_ & ~new_A6057_;
  assign new_A6068_ = new_A6089_ | new_A6088_;
  assign new_A6069_ = A6035 | new_A6068_;
  assign new_A6070_ = new_A6093_ | new_A6092_;
  assign new_A6071_ = ~A6035 & new_A6070_;
  assign new_A6072_ = new_A6091_ | new_A6090_;
  assign new_A6073_ = A6035 & new_A6072_;
  assign new_A6074_ = A6033 & ~new_A6043_;
  assign new_A6075_ = ~A6033 & new_A6043_;
  assign new_A6076_ = ~A6032 | ~new_A6057_;
  assign new_A6077_ = new_A6043_ & new_A6076_;
  assign new_A6078_ = ~new_A6043_ & ~new_A6077_;
  assign new_A6079_ = new_A6043_ | new_A6076_;
  assign new_A6080_ = ~A6033 & A6034;
  assign new_A6081_ = A6033 & ~A6034;
  assign new_A6082_ = new_A6050_ | new_A6087_;
  assign new_A6083_ = ~new_A6050_ & ~new_A6086_;
  assign new_A6084_ = A6033 | new_A6050_;
  assign new_A6085_ = A6033 | A6034;
  assign new_A6086_ = new_A6050_ & new_A6087_;
  assign new_A6087_ = ~A6032 | ~new_A6057_;
  assign new_A6088_ = new_A6065_ & new_A6085_;
  assign new_A6089_ = ~new_A6065_ & ~new_A6085_;
  assign new_A6090_ = new_A6094_ | new_A6095_;
  assign new_A6091_ = ~A6036 & new_A6050_;
  assign new_A6092_ = new_A6096_ | new_A6097_;
  assign new_A6093_ = A6036 & new_A6050_;
  assign new_A6094_ = ~A6036 & ~new_A6050_;
  assign new_A6095_ = A6036 & ~new_A6050_;
  assign new_A6096_ = A6036 & ~new_A6050_;
  assign new_A6097_ = ~A6036 & new_A6050_;
  assign new_A6104_ = new_A6111_ & new_A6110_;
  assign new_A6105_ = new_A6113_ | new_A6112_;
  assign new_A6106_ = new_A6115_ | new_A6114_;
  assign new_A6107_ = new_A6117_ & new_A6116_;
  assign new_A6108_ = new_A6117_ & new_A6118_;
  assign new_A6109_ = new_A6110_ | new_A6119_;
  assign new_A6110_ = A6099 | new_A6122_;
  assign new_A6111_ = new_A6121_ | new_A6120_;
  assign new_A6112_ = new_A6126_ & new_A6125_;
  assign new_A6113_ = new_A6124_ & new_A6123_;
  assign new_A6114_ = new_A6129_ | new_A6128_;
  assign new_A6115_ = new_A6124_ & new_A6127_;
  assign new_A6116_ = A6099 | new_A6132_;
  assign new_A6117_ = new_A6131_ | new_A6130_;
  assign new_A6118_ = new_A6134_ | new_A6133_;
  assign new_A6119_ = ~new_A6110_ & new_A6136_;
  assign new_A6120_ = ~new_A6112_ & new_A6124_;
  assign new_A6121_ = new_A6112_ & ~new_A6124_;
  assign new_A6122_ = A6098 & ~A6099;
  assign new_A6123_ = ~new_A6145_ | ~new_A6146_;
  assign new_A6124_ = new_A6138_ | new_A6140_;
  assign new_A6125_ = new_A6148_ | new_A6147_;
  assign new_A6126_ = new_A6142_ | new_A6141_;
  assign new_A6127_ = ~new_A6150_ | ~new_A6149_;
  assign new_A6128_ = ~new_A6151_ & new_A6152_;
  assign new_A6129_ = new_A6151_ & ~new_A6152_;
  assign new_A6130_ = ~A6098 & A6099;
  assign new_A6131_ = A6098 & ~A6099;
  assign new_A6132_ = ~new_A6114_ | new_A6124_;
  assign new_A6133_ = new_A6114_ & new_A6124_;
  assign new_A6134_ = ~new_A6114_ & ~new_A6124_;
  assign new_A6135_ = new_A6156_ | new_A6155_;
  assign new_A6136_ = A6102 | new_A6135_;
  assign new_A6137_ = new_A6160_ | new_A6159_;
  assign new_A6138_ = ~A6102 & new_A6137_;
  assign new_A6139_ = new_A6158_ | new_A6157_;
  assign new_A6140_ = A6102 & new_A6139_;
  assign new_A6141_ = A6100 & ~new_A6110_;
  assign new_A6142_ = ~A6100 & new_A6110_;
  assign new_A6143_ = ~A6099 | ~new_A6124_;
  assign new_A6144_ = new_A6110_ & new_A6143_;
  assign new_A6145_ = ~new_A6110_ & ~new_A6144_;
  assign new_A6146_ = new_A6110_ | new_A6143_;
  assign new_A6147_ = ~A6100 & A6101;
  assign new_A6148_ = A6100 & ~A6101;
  assign new_A6149_ = new_A6117_ | new_A6154_;
  assign new_A6150_ = ~new_A6117_ & ~new_A6153_;
  assign new_A6151_ = A6100 | new_A6117_;
  assign new_A6152_ = A6100 | A6101;
  assign new_A6153_ = new_A6117_ & new_A6154_;
  assign new_A6154_ = ~A6099 | ~new_A6124_;
  assign new_A6155_ = new_A6132_ & new_A6152_;
  assign new_A6156_ = ~new_A6132_ & ~new_A6152_;
  assign new_A6157_ = new_A6161_ | new_A6162_;
  assign new_A6158_ = ~A6103 & new_A6117_;
  assign new_A6159_ = new_A6163_ | new_A6164_;
  assign new_A6160_ = A6103 & new_A6117_;
  assign new_A6161_ = ~A6103 & ~new_A6117_;
  assign new_A6162_ = A6103 & ~new_A6117_;
  assign new_A6163_ = A6103 & ~new_A6117_;
  assign new_A6164_ = ~A6103 & new_A6117_;
  assign new_A6171_ = new_A6178_ & new_A6177_;
  assign new_A6172_ = new_A6180_ | new_A6179_;
  assign new_A6173_ = new_A6182_ | new_A6181_;
  assign new_A6174_ = new_A6184_ & new_A6183_;
  assign new_A6175_ = new_A6184_ & new_A6185_;
  assign new_A6176_ = new_A6177_ | new_A6186_;
  assign new_A6177_ = A6166 | new_A6189_;
  assign new_A6178_ = new_A6188_ | new_A6187_;
  assign new_A6179_ = new_A6193_ & new_A6192_;
  assign new_A6180_ = new_A6191_ & new_A6190_;
  assign new_A6181_ = new_A6196_ | new_A6195_;
  assign new_A6182_ = new_A6191_ & new_A6194_;
  assign new_A6183_ = A6166 | new_A6199_;
  assign new_A6184_ = new_A6198_ | new_A6197_;
  assign new_A6185_ = new_A6201_ | new_A6200_;
  assign new_A6186_ = ~new_A6177_ & new_A6203_;
  assign new_A6187_ = ~new_A6179_ & new_A6191_;
  assign new_A6188_ = new_A6179_ & ~new_A6191_;
  assign new_A6189_ = A6165 & ~A6166;
  assign new_A6190_ = ~new_A6212_ | ~new_A6213_;
  assign new_A6191_ = new_A6205_ | new_A6207_;
  assign new_A6192_ = new_A6215_ | new_A6214_;
  assign new_A6193_ = new_A6209_ | new_A6208_;
  assign new_A6194_ = ~new_A6217_ | ~new_A6216_;
  assign new_A6195_ = ~new_A6218_ & new_A6219_;
  assign new_A6196_ = new_A6218_ & ~new_A6219_;
  assign new_A6197_ = ~A6165 & A6166;
  assign new_A6198_ = A6165 & ~A6166;
  assign new_A6199_ = ~new_A6181_ | new_A6191_;
  assign new_A6200_ = new_A6181_ & new_A6191_;
  assign new_A6201_ = ~new_A6181_ & ~new_A6191_;
  assign new_A6202_ = new_A6223_ | new_A6222_;
  assign new_A6203_ = A6169 | new_A6202_;
  assign new_A6204_ = new_A6227_ | new_A6226_;
  assign new_A6205_ = ~A6169 & new_A6204_;
  assign new_A6206_ = new_A6225_ | new_A6224_;
  assign new_A6207_ = A6169 & new_A6206_;
  assign new_A6208_ = A6167 & ~new_A6177_;
  assign new_A6209_ = ~A6167 & new_A6177_;
  assign new_A6210_ = ~A6166 | ~new_A6191_;
  assign new_A6211_ = new_A6177_ & new_A6210_;
  assign new_A6212_ = ~new_A6177_ & ~new_A6211_;
  assign new_A6213_ = new_A6177_ | new_A6210_;
  assign new_A6214_ = ~A6167 & A6168;
  assign new_A6215_ = A6167 & ~A6168;
  assign new_A6216_ = new_A6184_ | new_A6221_;
  assign new_A6217_ = ~new_A6184_ & ~new_A6220_;
  assign new_A6218_ = A6167 | new_A6184_;
  assign new_A6219_ = A6167 | A6168;
  assign new_A6220_ = new_A6184_ & new_A6221_;
  assign new_A6221_ = ~A6166 | ~new_A6191_;
  assign new_A6222_ = new_A6199_ & new_A6219_;
  assign new_A6223_ = ~new_A6199_ & ~new_A6219_;
  assign new_A6224_ = new_A6228_ | new_A6229_;
  assign new_A6225_ = ~A6170 & new_A6184_;
  assign new_A6226_ = new_A6230_ | new_A6231_;
  assign new_A6227_ = A6170 & new_A6184_;
  assign new_A6228_ = ~A6170 & ~new_A6184_;
  assign new_A6229_ = A6170 & ~new_A6184_;
  assign new_A6230_ = A6170 & ~new_A6184_;
  assign new_A6231_ = ~A6170 & new_A6184_;
  assign new_A6238_ = new_A6245_ & new_A6244_;
  assign new_A6239_ = new_A6247_ | new_A6246_;
  assign new_A6240_ = new_A6249_ | new_A6248_;
  assign new_A6241_ = new_A6251_ & new_A6250_;
  assign new_A6242_ = new_A6251_ & new_A6252_;
  assign new_A6243_ = new_A6244_ | new_A6253_;
  assign new_A6244_ = A6233 | new_A6256_;
  assign new_A6245_ = new_A6255_ | new_A6254_;
  assign new_A6246_ = new_A6260_ & new_A6259_;
  assign new_A6247_ = new_A6258_ & new_A6257_;
  assign new_A6248_ = new_A6263_ | new_A6262_;
  assign new_A6249_ = new_A6258_ & new_A6261_;
  assign new_A6250_ = A6233 | new_A6266_;
  assign new_A6251_ = new_A6265_ | new_A6264_;
  assign new_A6252_ = new_A6268_ | new_A6267_;
  assign new_A6253_ = ~new_A6244_ & new_A6270_;
  assign new_A6254_ = ~new_A6246_ & new_A6258_;
  assign new_A6255_ = new_A6246_ & ~new_A6258_;
  assign new_A6256_ = A6232 & ~A6233;
  assign new_A6257_ = ~new_A6279_ | ~new_A6280_;
  assign new_A6258_ = new_A6272_ | new_A6274_;
  assign new_A6259_ = new_A6282_ | new_A6281_;
  assign new_A6260_ = new_A6276_ | new_A6275_;
  assign new_A6261_ = ~new_A6284_ | ~new_A6283_;
  assign new_A6262_ = ~new_A6285_ & new_A6286_;
  assign new_A6263_ = new_A6285_ & ~new_A6286_;
  assign new_A6264_ = ~A6232 & A6233;
  assign new_A6265_ = A6232 & ~A6233;
  assign new_A6266_ = ~new_A6248_ | new_A6258_;
  assign new_A6267_ = new_A6248_ & new_A6258_;
  assign new_A6268_ = ~new_A6248_ & ~new_A6258_;
  assign new_A6269_ = new_A6290_ | new_A6289_;
  assign new_A6270_ = A6236 | new_A6269_;
  assign new_A6271_ = new_A6294_ | new_A6293_;
  assign new_A6272_ = ~A6236 & new_A6271_;
  assign new_A6273_ = new_A6292_ | new_A6291_;
  assign new_A6274_ = A6236 & new_A6273_;
  assign new_A6275_ = A6234 & ~new_A6244_;
  assign new_A6276_ = ~A6234 & new_A6244_;
  assign new_A6277_ = ~A6233 | ~new_A6258_;
  assign new_A6278_ = new_A6244_ & new_A6277_;
  assign new_A6279_ = ~new_A6244_ & ~new_A6278_;
  assign new_A6280_ = new_A6244_ | new_A6277_;
  assign new_A6281_ = ~A6234 & A6235;
  assign new_A6282_ = A6234 & ~A6235;
  assign new_A6283_ = new_A6251_ | new_A6288_;
  assign new_A6284_ = ~new_A6251_ & ~new_A6287_;
  assign new_A6285_ = A6234 | new_A6251_;
  assign new_A6286_ = A6234 | A6235;
  assign new_A6287_ = new_A6251_ & new_A6288_;
  assign new_A6288_ = ~A6233 | ~new_A6258_;
  assign new_A6289_ = new_A6266_ & new_A6286_;
  assign new_A6290_ = ~new_A6266_ & ~new_A6286_;
  assign new_A6291_ = new_A6295_ | new_A6296_;
  assign new_A6292_ = ~A6237 & new_A6251_;
  assign new_A6293_ = new_A6297_ | new_A6298_;
  assign new_A6294_ = A6237 & new_A6251_;
  assign new_A6295_ = ~A6237 & ~new_A6251_;
  assign new_A6296_ = A6237 & ~new_A6251_;
  assign new_A6297_ = A6237 & ~new_A6251_;
  assign new_A6298_ = ~A6237 & new_A6251_;
  assign new_A6305_ = new_A6312_ & new_A6311_;
  assign new_A6306_ = new_A6314_ | new_A6313_;
  assign new_A6307_ = new_A6316_ | new_A6315_;
  assign new_A6308_ = new_A6318_ & new_A6317_;
  assign new_A6309_ = new_A6318_ & new_A6319_;
  assign new_A6310_ = new_A6311_ | new_A6320_;
  assign new_A6311_ = A6300 | new_A6323_;
  assign new_A6312_ = new_A6322_ | new_A6321_;
  assign new_A6313_ = new_A6327_ & new_A6326_;
  assign new_A6314_ = new_A6325_ & new_A6324_;
  assign new_A6315_ = new_A6330_ | new_A6329_;
  assign new_A6316_ = new_A6325_ & new_A6328_;
  assign new_A6317_ = A6300 | new_A6333_;
  assign new_A6318_ = new_A6332_ | new_A6331_;
  assign new_A6319_ = new_A6335_ | new_A6334_;
  assign new_A6320_ = ~new_A6311_ & new_A6337_;
  assign new_A6321_ = ~new_A6313_ & new_A6325_;
  assign new_A6322_ = new_A6313_ & ~new_A6325_;
  assign new_A6323_ = A6299 & ~A6300;
  assign new_A6324_ = ~new_A6346_ | ~new_A6347_;
  assign new_A6325_ = new_A6339_ | new_A6341_;
  assign new_A6326_ = new_A6349_ | new_A6348_;
  assign new_A6327_ = new_A6343_ | new_A6342_;
  assign new_A6328_ = ~new_A6351_ | ~new_A6350_;
  assign new_A6329_ = ~new_A6352_ & new_A6353_;
  assign new_A6330_ = new_A6352_ & ~new_A6353_;
  assign new_A6331_ = ~A6299 & A6300;
  assign new_A6332_ = A6299 & ~A6300;
  assign new_A6333_ = ~new_A6315_ | new_A6325_;
  assign new_A6334_ = new_A6315_ & new_A6325_;
  assign new_A6335_ = ~new_A6315_ & ~new_A6325_;
  assign new_A6336_ = new_A6357_ | new_A6356_;
  assign new_A6337_ = A6303 | new_A6336_;
  assign new_A6338_ = new_A6361_ | new_A6360_;
  assign new_A6339_ = ~A6303 & new_A6338_;
  assign new_A6340_ = new_A6359_ | new_A6358_;
  assign new_A6341_ = A6303 & new_A6340_;
  assign new_A6342_ = A6301 & ~new_A6311_;
  assign new_A6343_ = ~A6301 & new_A6311_;
  assign new_A6344_ = ~A6300 | ~new_A6325_;
  assign new_A6345_ = new_A6311_ & new_A6344_;
  assign new_A6346_ = ~new_A6311_ & ~new_A6345_;
  assign new_A6347_ = new_A6311_ | new_A6344_;
  assign new_A6348_ = ~A6301 & A6302;
  assign new_A6349_ = A6301 & ~A6302;
  assign new_A6350_ = new_A6318_ | new_A6355_;
  assign new_A6351_ = ~new_A6318_ & ~new_A6354_;
  assign new_A6352_ = A6301 | new_A6318_;
  assign new_A6353_ = A6301 | A6302;
  assign new_A6354_ = new_A6318_ & new_A6355_;
  assign new_A6355_ = ~A6300 | ~new_A6325_;
  assign new_A6356_ = new_A6333_ & new_A6353_;
  assign new_A6357_ = ~new_A6333_ & ~new_A6353_;
  assign new_A6358_ = new_A6362_ | new_A6363_;
  assign new_A6359_ = ~A6304 & new_A6318_;
  assign new_A6360_ = new_A6364_ | new_A6365_;
  assign new_A6361_ = A6304 & new_A6318_;
  assign new_A6362_ = ~A6304 & ~new_A6318_;
  assign new_A6363_ = A6304 & ~new_A6318_;
  assign new_A6364_ = A6304 & ~new_A6318_;
  assign new_A6365_ = ~A6304 & new_A6318_;
  assign new_A6372_ = new_A6379_ & new_A6378_;
  assign new_A6373_ = new_A6381_ | new_A6380_;
  assign new_A6374_ = new_A6383_ | new_A6382_;
  assign new_A6375_ = new_A6385_ & new_A6384_;
  assign new_A6376_ = new_A6385_ & new_A6386_;
  assign new_A6377_ = new_A6378_ | new_A6387_;
  assign new_A6378_ = A6367 | new_A6390_;
  assign new_A6379_ = new_A6389_ | new_A6388_;
  assign new_A6380_ = new_A6394_ & new_A6393_;
  assign new_A6381_ = new_A6392_ & new_A6391_;
  assign new_A6382_ = new_A6397_ | new_A6396_;
  assign new_A6383_ = new_A6392_ & new_A6395_;
  assign new_A6384_ = A6367 | new_A6400_;
  assign new_A6385_ = new_A6399_ | new_A6398_;
  assign new_A6386_ = new_A6402_ | new_A6401_;
  assign new_A6387_ = ~new_A6378_ & new_A6404_;
  assign new_A6388_ = ~new_A6380_ & new_A6392_;
  assign new_A6389_ = new_A6380_ & ~new_A6392_;
  assign new_A6390_ = A6366 & ~A6367;
  assign new_A6391_ = ~new_A6413_ | ~new_A6414_;
  assign new_A6392_ = new_A6406_ | new_A6408_;
  assign new_A6393_ = new_A6416_ | new_A6415_;
  assign new_A6394_ = new_A6410_ | new_A6409_;
  assign new_A6395_ = ~new_A6418_ | ~new_A6417_;
  assign new_A6396_ = ~new_A6419_ & new_A6420_;
  assign new_A6397_ = new_A6419_ & ~new_A6420_;
  assign new_A6398_ = ~A6366 & A6367;
  assign new_A6399_ = A6366 & ~A6367;
  assign new_A6400_ = ~new_A6382_ | new_A6392_;
  assign new_A6401_ = new_A6382_ & new_A6392_;
  assign new_A6402_ = ~new_A6382_ & ~new_A6392_;
  assign new_A6403_ = new_A6424_ | new_A6423_;
  assign new_A6404_ = A6370 | new_A6403_;
  assign new_A6405_ = new_A6428_ | new_A6427_;
  assign new_A6406_ = ~A6370 & new_A6405_;
  assign new_A6407_ = new_A6426_ | new_A6425_;
  assign new_A6408_ = A6370 & new_A6407_;
  assign new_A6409_ = A6368 & ~new_A6378_;
  assign new_A6410_ = ~A6368 & new_A6378_;
  assign new_A6411_ = ~A6367 | ~new_A6392_;
  assign new_A6412_ = new_A6378_ & new_A6411_;
  assign new_A6413_ = ~new_A6378_ & ~new_A6412_;
  assign new_A6414_ = new_A6378_ | new_A6411_;
  assign new_A6415_ = ~A6368 & A6369;
  assign new_A6416_ = A6368 & ~A6369;
  assign new_A6417_ = new_A6385_ | new_A6422_;
  assign new_A6418_ = ~new_A6385_ & ~new_A6421_;
  assign new_A6419_ = A6368 | new_A6385_;
  assign new_A6420_ = A6368 | A6369;
  assign new_A6421_ = new_A6385_ & new_A6422_;
  assign new_A6422_ = ~A6367 | ~new_A6392_;
  assign new_A6423_ = new_A6400_ & new_A6420_;
  assign new_A6424_ = ~new_A6400_ & ~new_A6420_;
  assign new_A6425_ = new_A6429_ | new_A6430_;
  assign new_A6426_ = ~A6371 & new_A6385_;
  assign new_A6427_ = new_A6431_ | new_A6432_;
  assign new_A6428_ = A6371 & new_A6385_;
  assign new_A6429_ = ~A6371 & ~new_A6385_;
  assign new_A6430_ = A6371 & ~new_A6385_;
  assign new_A6431_ = A6371 & ~new_A6385_;
  assign new_A6432_ = ~A6371 & new_A6385_;
  assign new_A6439_ = new_A6446_ & new_A6445_;
  assign new_A6440_ = new_A6448_ | new_A6447_;
  assign new_A6441_ = new_A6450_ | new_A6449_;
  assign new_A6442_ = new_A6452_ & new_A6451_;
  assign new_A6443_ = new_A6452_ & new_A6453_;
  assign new_A6444_ = new_A6445_ | new_A6454_;
  assign new_A6445_ = A6434 | new_A6457_;
  assign new_A6446_ = new_A6456_ | new_A6455_;
  assign new_A6447_ = new_A6461_ & new_A6460_;
  assign new_A6448_ = new_A6459_ & new_A6458_;
  assign new_A6449_ = new_A6464_ | new_A6463_;
  assign new_A6450_ = new_A6459_ & new_A6462_;
  assign new_A6451_ = A6434 | new_A6467_;
  assign new_A6452_ = new_A6466_ | new_A6465_;
  assign new_A6453_ = new_A6469_ | new_A6468_;
  assign new_A6454_ = ~new_A6445_ & new_A6471_;
  assign new_A6455_ = ~new_A6447_ & new_A6459_;
  assign new_A6456_ = new_A6447_ & ~new_A6459_;
  assign new_A6457_ = A6433 & ~A6434;
  assign new_A6458_ = ~new_A6480_ | ~new_A6481_;
  assign new_A6459_ = new_A6473_ | new_A6475_;
  assign new_A6460_ = new_A6483_ | new_A6482_;
  assign new_A6461_ = new_A6477_ | new_A6476_;
  assign new_A6462_ = ~new_A6485_ | ~new_A6484_;
  assign new_A6463_ = ~new_A6486_ & new_A6487_;
  assign new_A6464_ = new_A6486_ & ~new_A6487_;
  assign new_A6465_ = ~A6433 & A6434;
  assign new_A6466_ = A6433 & ~A6434;
  assign new_A6467_ = ~new_A6449_ | new_A6459_;
  assign new_A6468_ = new_A6449_ & new_A6459_;
  assign new_A6469_ = ~new_A6449_ & ~new_A6459_;
  assign new_A6470_ = new_A6491_ | new_A6490_;
  assign new_A6471_ = A6437 | new_A6470_;
  assign new_A6472_ = new_A6495_ | new_A6494_;
  assign new_A6473_ = ~A6437 & new_A6472_;
  assign new_A6474_ = new_A6493_ | new_A6492_;
  assign new_A6475_ = A6437 & new_A6474_;
  assign new_A6476_ = A6435 & ~new_A6445_;
  assign new_A6477_ = ~A6435 & new_A6445_;
  assign new_A6478_ = ~A6434 | ~new_A6459_;
  assign new_A6479_ = new_A6445_ & new_A6478_;
  assign new_A6480_ = ~new_A6445_ & ~new_A6479_;
  assign new_A6481_ = new_A6445_ | new_A6478_;
  assign new_A6482_ = ~A6435 & A6436;
  assign new_A6483_ = A6435 & ~A6436;
  assign new_A6484_ = new_A6452_ | new_A6489_;
  assign new_A6485_ = ~new_A6452_ & ~new_A6488_;
  assign new_A6486_ = A6435 | new_A6452_;
  assign new_A6487_ = A6435 | A6436;
  assign new_A6488_ = new_A6452_ & new_A6489_;
  assign new_A6489_ = ~A6434 | ~new_A6459_;
  assign new_A6490_ = new_A6467_ & new_A6487_;
  assign new_A6491_ = ~new_A6467_ & ~new_A6487_;
  assign new_A6492_ = new_A6496_ | new_A6497_;
  assign new_A6493_ = ~A6438 & new_A6452_;
  assign new_A6494_ = new_A6498_ | new_A6499_;
  assign new_A6495_ = A6438 & new_A6452_;
  assign new_A6496_ = ~A6438 & ~new_A6452_;
  assign new_A6497_ = A6438 & ~new_A6452_;
  assign new_A6498_ = A6438 & ~new_A6452_;
  assign new_A6499_ = ~A6438 & new_A6452_;
  assign new_A6506_ = new_A6513_ & new_A6512_;
  assign new_A6507_ = new_A6515_ | new_A6514_;
  assign new_A6508_ = new_A6517_ | new_A6516_;
  assign new_A6509_ = new_A6519_ & new_A6518_;
  assign new_A6510_ = new_A6519_ & new_A6520_;
  assign new_A6511_ = new_A6512_ | new_A6521_;
  assign new_A6512_ = A6501 | new_A6524_;
  assign new_A6513_ = new_A6523_ | new_A6522_;
  assign new_A6514_ = new_A6528_ & new_A6527_;
  assign new_A6515_ = new_A6526_ & new_A6525_;
  assign new_A6516_ = new_A6531_ | new_A6530_;
  assign new_A6517_ = new_A6526_ & new_A6529_;
  assign new_A6518_ = A6501 | new_A6534_;
  assign new_A6519_ = new_A6533_ | new_A6532_;
  assign new_A6520_ = new_A6536_ | new_A6535_;
  assign new_A6521_ = ~new_A6512_ & new_A6538_;
  assign new_A6522_ = ~new_A6514_ & new_A6526_;
  assign new_A6523_ = new_A6514_ & ~new_A6526_;
  assign new_A6524_ = A6500 & ~A6501;
  assign new_A6525_ = ~new_A6547_ | ~new_A6548_;
  assign new_A6526_ = new_A6540_ | new_A6542_;
  assign new_A6527_ = new_A6550_ | new_A6549_;
  assign new_A6528_ = new_A6544_ | new_A6543_;
  assign new_A6529_ = ~new_A6552_ | ~new_A6551_;
  assign new_A6530_ = ~new_A6553_ & new_A6554_;
  assign new_A6531_ = new_A6553_ & ~new_A6554_;
  assign new_A6532_ = ~A6500 & A6501;
  assign new_A6533_ = A6500 & ~A6501;
  assign new_A6534_ = ~new_A6516_ | new_A6526_;
  assign new_A6535_ = new_A6516_ & new_A6526_;
  assign new_A6536_ = ~new_A6516_ & ~new_A6526_;
  assign new_A6537_ = new_A6558_ | new_A6557_;
  assign new_A6538_ = A6504 | new_A6537_;
  assign new_A6539_ = new_A6562_ | new_A6561_;
  assign new_A6540_ = ~A6504 & new_A6539_;
  assign new_A6541_ = new_A6560_ | new_A6559_;
  assign new_A6542_ = A6504 & new_A6541_;
  assign new_A6543_ = A6502 & ~new_A6512_;
  assign new_A6544_ = ~A6502 & new_A6512_;
  assign new_A6545_ = ~A6501 | ~new_A6526_;
  assign new_A6546_ = new_A6512_ & new_A6545_;
  assign new_A6547_ = ~new_A6512_ & ~new_A6546_;
  assign new_A6548_ = new_A6512_ | new_A6545_;
  assign new_A6549_ = ~A6502 & A6503;
  assign new_A6550_ = A6502 & ~A6503;
  assign new_A6551_ = new_A6519_ | new_A6556_;
  assign new_A6552_ = ~new_A6519_ & ~new_A6555_;
  assign new_A6553_ = A6502 | new_A6519_;
  assign new_A6554_ = A6502 | A6503;
  assign new_A6555_ = new_A6519_ & new_A6556_;
  assign new_A6556_ = ~A6501 | ~new_A6526_;
  assign new_A6557_ = new_A6534_ & new_A6554_;
  assign new_A6558_ = ~new_A6534_ & ~new_A6554_;
  assign new_A6559_ = new_A6563_ | new_A6564_;
  assign new_A6560_ = ~A6505 & new_A6519_;
  assign new_A6561_ = new_A6565_ | new_A6566_;
  assign new_A6562_ = A6505 & new_A6519_;
  assign new_A6563_ = ~A6505 & ~new_A6519_;
  assign new_A6564_ = A6505 & ~new_A6519_;
  assign new_A6565_ = A6505 & ~new_A6519_;
  assign new_A6566_ = ~A6505 & new_A6519_;
  assign new_A6573_ = new_A6580_ & new_A6579_;
  assign new_A6574_ = new_A6582_ | new_A6581_;
  assign new_A6575_ = new_A6584_ | new_A6583_;
  assign new_A6576_ = new_A6586_ & new_A6585_;
  assign new_A6577_ = new_A6586_ & new_A6587_;
  assign new_A6578_ = new_A6579_ | new_A6588_;
  assign new_A6579_ = A6568 | new_A6591_;
  assign new_A6580_ = new_A6590_ | new_A6589_;
  assign new_A6581_ = new_A6595_ & new_A6594_;
  assign new_A6582_ = new_A6593_ & new_A6592_;
  assign new_A6583_ = new_A6598_ | new_A6597_;
  assign new_A6584_ = new_A6593_ & new_A6596_;
  assign new_A6585_ = A6568 | new_A6601_;
  assign new_A6586_ = new_A6600_ | new_A6599_;
  assign new_A6587_ = new_A6603_ | new_A6602_;
  assign new_A6588_ = ~new_A6579_ & new_A6605_;
  assign new_A6589_ = ~new_A6581_ & new_A6593_;
  assign new_A6590_ = new_A6581_ & ~new_A6593_;
  assign new_A6591_ = A6567 & ~A6568;
  assign new_A6592_ = ~new_A6614_ | ~new_A6615_;
  assign new_A6593_ = new_A6607_ | new_A6609_;
  assign new_A6594_ = new_A6617_ | new_A6616_;
  assign new_A6595_ = new_A6611_ | new_A6610_;
  assign new_A6596_ = ~new_A6619_ | ~new_A6618_;
  assign new_A6597_ = ~new_A6620_ & new_A6621_;
  assign new_A6598_ = new_A6620_ & ~new_A6621_;
  assign new_A6599_ = ~A6567 & A6568;
  assign new_A6600_ = A6567 & ~A6568;
  assign new_A6601_ = ~new_A6583_ | new_A6593_;
  assign new_A6602_ = new_A6583_ & new_A6593_;
  assign new_A6603_ = ~new_A6583_ & ~new_A6593_;
  assign new_A6604_ = new_A6625_ | new_A6624_;
  assign new_A6605_ = A6571 | new_A6604_;
  assign new_A6606_ = new_A6629_ | new_A6628_;
  assign new_A6607_ = ~A6571 & new_A6606_;
  assign new_A6608_ = new_A6627_ | new_A6626_;
  assign new_A6609_ = A6571 & new_A6608_;
  assign new_A6610_ = A6569 & ~new_A6579_;
  assign new_A6611_ = ~A6569 & new_A6579_;
  assign new_A6612_ = ~A6568 | ~new_A6593_;
  assign new_A6613_ = new_A6579_ & new_A6612_;
  assign new_A6614_ = ~new_A6579_ & ~new_A6613_;
  assign new_A6615_ = new_A6579_ | new_A6612_;
  assign new_A6616_ = ~A6569 & A6570;
  assign new_A6617_ = A6569 & ~A6570;
  assign new_A6618_ = new_A6586_ | new_A6623_;
  assign new_A6619_ = ~new_A6586_ & ~new_A6622_;
  assign new_A6620_ = A6569 | new_A6586_;
  assign new_A6621_ = A6569 | A6570;
  assign new_A6622_ = new_A6586_ & new_A6623_;
  assign new_A6623_ = ~A6568 | ~new_A6593_;
  assign new_A6624_ = new_A6601_ & new_A6621_;
  assign new_A6625_ = ~new_A6601_ & ~new_A6621_;
  assign new_A6626_ = new_A6630_ | new_A6631_;
  assign new_A6627_ = ~A6572 & new_A6586_;
  assign new_A6628_ = new_A6632_ | new_A6633_;
  assign new_A6629_ = A6572 & new_A6586_;
  assign new_A6630_ = ~A6572 & ~new_A6586_;
  assign new_A6631_ = A6572 & ~new_A6586_;
  assign new_A6632_ = A6572 & ~new_A6586_;
  assign new_A6633_ = ~A6572 & new_A6586_;
  assign new_A6640_ = new_A6647_ & new_A6646_;
  assign new_A6641_ = new_A6649_ | new_A6648_;
  assign new_A6642_ = new_A6651_ | new_A6650_;
  assign new_A6643_ = new_A6653_ & new_A6652_;
  assign new_A6644_ = new_A6653_ & new_A6654_;
  assign new_A6645_ = new_A6646_ | new_A6655_;
  assign new_A6646_ = A6635 | new_A6658_;
  assign new_A6647_ = new_A6657_ | new_A6656_;
  assign new_A6648_ = new_A6662_ & new_A6661_;
  assign new_A6649_ = new_A6660_ & new_A6659_;
  assign new_A6650_ = new_A6665_ | new_A6664_;
  assign new_A6651_ = new_A6660_ & new_A6663_;
  assign new_A6652_ = A6635 | new_A6668_;
  assign new_A6653_ = new_A6667_ | new_A6666_;
  assign new_A6654_ = new_A6670_ | new_A6669_;
  assign new_A6655_ = ~new_A6646_ & new_A6672_;
  assign new_A6656_ = ~new_A6648_ & new_A6660_;
  assign new_A6657_ = new_A6648_ & ~new_A6660_;
  assign new_A6658_ = A6634 & ~A6635;
  assign new_A6659_ = ~new_A6681_ | ~new_A6682_;
  assign new_A6660_ = new_A6674_ | new_A6676_;
  assign new_A6661_ = new_A6684_ | new_A6683_;
  assign new_A6662_ = new_A6678_ | new_A6677_;
  assign new_A6663_ = ~new_A6686_ | ~new_A6685_;
  assign new_A6664_ = ~new_A6687_ & new_A6688_;
  assign new_A6665_ = new_A6687_ & ~new_A6688_;
  assign new_A6666_ = ~A6634 & A6635;
  assign new_A6667_ = A6634 & ~A6635;
  assign new_A6668_ = ~new_A6650_ | new_A6660_;
  assign new_A6669_ = new_A6650_ & new_A6660_;
  assign new_A6670_ = ~new_A6650_ & ~new_A6660_;
  assign new_A6671_ = new_A6692_ | new_A6691_;
  assign new_A6672_ = A6638 | new_A6671_;
  assign new_A6673_ = new_A6696_ | new_A6695_;
  assign new_A6674_ = ~A6638 & new_A6673_;
  assign new_A6675_ = new_A6694_ | new_A6693_;
  assign new_A6676_ = A6638 & new_A6675_;
  assign new_A6677_ = A6636 & ~new_A6646_;
  assign new_A6678_ = ~A6636 & new_A6646_;
  assign new_A6679_ = ~A6635 | ~new_A6660_;
  assign new_A6680_ = new_A6646_ & new_A6679_;
  assign new_A6681_ = ~new_A6646_ & ~new_A6680_;
  assign new_A6682_ = new_A6646_ | new_A6679_;
  assign new_A6683_ = ~A6636 & A6637;
  assign new_A6684_ = A6636 & ~A6637;
  assign new_A6685_ = new_A6653_ | new_A6690_;
  assign new_A6686_ = ~new_A6653_ & ~new_A6689_;
  assign new_A6687_ = A6636 | new_A6653_;
  assign new_A6688_ = A6636 | A6637;
  assign new_A6689_ = new_A6653_ & new_A6690_;
  assign new_A6690_ = ~A6635 | ~new_A6660_;
  assign new_A6691_ = new_A6668_ & new_A6688_;
  assign new_A6692_ = ~new_A6668_ & ~new_A6688_;
  assign new_A6693_ = new_A6697_ | new_A6698_;
  assign new_A6694_ = ~A6639 & new_A6653_;
  assign new_A6695_ = new_A6699_ | new_A6700_;
  assign new_A6696_ = A6639 & new_A6653_;
  assign new_A6697_ = ~A6639 & ~new_A6653_;
  assign new_A6698_ = A6639 & ~new_A6653_;
  assign new_A6699_ = A6639 & ~new_A6653_;
  assign new_A6700_ = ~A6639 & new_A6653_;
  assign new_A6707_ = new_A6714_ & new_A6713_;
  assign new_A6708_ = new_A6716_ | new_A6715_;
  assign new_A6709_ = new_A6718_ | new_A6717_;
  assign new_A6710_ = new_A6720_ & new_A6719_;
  assign new_A6711_ = new_A6720_ & new_A6721_;
  assign new_A6712_ = new_A6713_ | new_A6722_;
  assign new_A6713_ = A6702 | new_A6725_;
  assign new_A6714_ = new_A6724_ | new_A6723_;
  assign new_A6715_ = new_A6729_ & new_A6728_;
  assign new_A6716_ = new_A6727_ & new_A6726_;
  assign new_A6717_ = new_A6732_ | new_A6731_;
  assign new_A6718_ = new_A6727_ & new_A6730_;
  assign new_A6719_ = A6702 | new_A6735_;
  assign new_A6720_ = new_A6734_ | new_A6733_;
  assign new_A6721_ = new_A6737_ | new_A6736_;
  assign new_A6722_ = ~new_A6713_ & new_A6739_;
  assign new_A6723_ = ~new_A6715_ & new_A6727_;
  assign new_A6724_ = new_A6715_ & ~new_A6727_;
  assign new_A6725_ = A6701 & ~A6702;
  assign new_A6726_ = ~new_A6748_ | ~new_A6749_;
  assign new_A6727_ = new_A6741_ | new_A6743_;
  assign new_A6728_ = new_A6751_ | new_A6750_;
  assign new_A6729_ = new_A6745_ | new_A6744_;
  assign new_A6730_ = ~new_A6753_ | ~new_A6752_;
  assign new_A6731_ = ~new_A6754_ & new_A6755_;
  assign new_A6732_ = new_A6754_ & ~new_A6755_;
  assign new_A6733_ = ~A6701 & A6702;
  assign new_A6734_ = A6701 & ~A6702;
  assign new_A6735_ = ~new_A6717_ | new_A6727_;
  assign new_A6736_ = new_A6717_ & new_A6727_;
  assign new_A6737_ = ~new_A6717_ & ~new_A6727_;
  assign new_A6738_ = new_A6759_ | new_A6758_;
  assign new_A6739_ = A6705 | new_A6738_;
  assign new_A6740_ = new_A6763_ | new_A6762_;
  assign new_A6741_ = ~A6705 & new_A6740_;
  assign new_A6742_ = new_A6761_ | new_A6760_;
  assign new_A6743_ = A6705 & new_A6742_;
  assign new_A6744_ = A6703 & ~new_A6713_;
  assign new_A6745_ = ~A6703 & new_A6713_;
  assign new_A6746_ = ~A6702 | ~new_A6727_;
  assign new_A6747_ = new_A6713_ & new_A6746_;
  assign new_A6748_ = ~new_A6713_ & ~new_A6747_;
  assign new_A6749_ = new_A6713_ | new_A6746_;
  assign new_A6750_ = ~A6703 & A6704;
  assign new_A6751_ = A6703 & ~A6704;
  assign new_A6752_ = new_A6720_ | new_A6757_;
  assign new_A6753_ = ~new_A6720_ & ~new_A6756_;
  assign new_A6754_ = A6703 | new_A6720_;
  assign new_A6755_ = A6703 | A6704;
  assign new_A6756_ = new_A6720_ & new_A6757_;
  assign new_A6757_ = ~A6702 | ~new_A6727_;
  assign new_A6758_ = new_A6735_ & new_A6755_;
  assign new_A6759_ = ~new_A6735_ & ~new_A6755_;
  assign new_A6760_ = new_A6764_ | new_A6765_;
  assign new_A6761_ = ~A6706 & new_A6720_;
  assign new_A6762_ = new_A6766_ | new_A6767_;
  assign new_A6763_ = A6706 & new_A6720_;
  assign new_A6764_ = ~A6706 & ~new_A6720_;
  assign new_A6765_ = A6706 & ~new_A6720_;
  assign new_A6766_ = A6706 & ~new_A6720_;
  assign new_A6767_ = ~A6706 & new_A6720_;
  assign new_A6774_ = new_A6781_ & new_A6780_;
  assign new_A6775_ = new_A6783_ | new_A6782_;
  assign new_A6776_ = new_A6785_ | new_A6784_;
  assign new_A6777_ = new_A6787_ & new_A6786_;
  assign new_A6778_ = new_A6787_ & new_A6788_;
  assign new_A6779_ = new_A6780_ | new_A6789_;
  assign new_A6780_ = A6769 | new_A6792_;
  assign new_A6781_ = new_A6791_ | new_A6790_;
  assign new_A6782_ = new_A6796_ & new_A6795_;
  assign new_A6783_ = new_A6794_ & new_A6793_;
  assign new_A6784_ = new_A6799_ | new_A6798_;
  assign new_A6785_ = new_A6794_ & new_A6797_;
  assign new_A6786_ = A6769 | new_A6802_;
  assign new_A6787_ = new_A6801_ | new_A6800_;
  assign new_A6788_ = new_A6804_ | new_A6803_;
  assign new_A6789_ = ~new_A6780_ & new_A6806_;
  assign new_A6790_ = ~new_A6782_ & new_A6794_;
  assign new_A6791_ = new_A6782_ & ~new_A6794_;
  assign new_A6792_ = A6768 & ~A6769;
  assign new_A6793_ = ~new_A6815_ | ~new_A6816_;
  assign new_A6794_ = new_A6808_ | new_A6810_;
  assign new_A6795_ = new_A6818_ | new_A6817_;
  assign new_A6796_ = new_A6812_ | new_A6811_;
  assign new_A6797_ = ~new_A6820_ | ~new_A6819_;
  assign new_A6798_ = ~new_A6821_ & new_A6822_;
  assign new_A6799_ = new_A6821_ & ~new_A6822_;
  assign new_A6800_ = ~A6768 & A6769;
  assign new_A6801_ = A6768 & ~A6769;
  assign new_A6802_ = ~new_A6784_ | new_A6794_;
  assign new_A6803_ = new_A6784_ & new_A6794_;
  assign new_A6804_ = ~new_A6784_ & ~new_A6794_;
  assign new_A6805_ = new_A6826_ | new_A6825_;
  assign new_A6806_ = A6772 | new_A6805_;
  assign new_A6807_ = new_A6830_ | new_A6829_;
  assign new_A6808_ = ~A6772 & new_A6807_;
  assign new_A6809_ = new_A6828_ | new_A6827_;
  assign new_A6810_ = A6772 & new_A6809_;
  assign new_A6811_ = A6770 & ~new_A6780_;
  assign new_A6812_ = ~A6770 & new_A6780_;
  assign new_A6813_ = ~A6769 | ~new_A6794_;
  assign new_A6814_ = new_A6780_ & new_A6813_;
  assign new_A6815_ = ~new_A6780_ & ~new_A6814_;
  assign new_A6816_ = new_A6780_ | new_A6813_;
  assign new_A6817_ = ~A6770 & A6771;
  assign new_A6818_ = A6770 & ~A6771;
  assign new_A6819_ = new_A6787_ | new_A6824_;
  assign new_A6820_ = ~new_A6787_ & ~new_A6823_;
  assign new_A6821_ = A6770 | new_A6787_;
  assign new_A6822_ = A6770 | A6771;
  assign new_A6823_ = new_A6787_ & new_A6824_;
  assign new_A6824_ = ~A6769 | ~new_A6794_;
  assign new_A6825_ = new_A6802_ & new_A6822_;
  assign new_A6826_ = ~new_A6802_ & ~new_A6822_;
  assign new_A6827_ = new_A6831_ | new_A6832_;
  assign new_A6828_ = ~A6773 & new_A6787_;
  assign new_A6829_ = new_A6833_ | new_A6834_;
  assign new_A6830_ = A6773 & new_A6787_;
  assign new_A6831_ = ~A6773 & ~new_A6787_;
  assign new_A6832_ = A6773 & ~new_A6787_;
  assign new_A6833_ = A6773 & ~new_A6787_;
  assign new_A6834_ = ~A6773 & new_A6787_;
  assign new_A6841_ = new_A6848_ & new_A6847_;
  assign new_A6842_ = new_A6850_ | new_A6849_;
  assign new_A6843_ = new_A6852_ | new_A6851_;
  assign new_A6844_ = new_A6854_ & new_A6853_;
  assign new_A6845_ = new_A6854_ & new_A6855_;
  assign new_A6846_ = new_A6847_ | new_A6856_;
  assign new_A6847_ = A6836 | new_A6859_;
  assign new_A6848_ = new_A6858_ | new_A6857_;
  assign new_A6849_ = new_A6863_ & new_A6862_;
  assign new_A6850_ = new_A6861_ & new_A6860_;
  assign new_A6851_ = new_A6866_ | new_A6865_;
  assign new_A6852_ = new_A6861_ & new_A6864_;
  assign new_A6853_ = A6836 | new_A6869_;
  assign new_A6854_ = new_A6868_ | new_A6867_;
  assign new_A6855_ = new_A6871_ | new_A6870_;
  assign new_A6856_ = ~new_A6847_ & new_A6873_;
  assign new_A6857_ = ~new_A6849_ & new_A6861_;
  assign new_A6858_ = new_A6849_ & ~new_A6861_;
  assign new_A6859_ = A6835 & ~A6836;
  assign new_A6860_ = ~new_A6882_ | ~new_A6883_;
  assign new_A6861_ = new_A6875_ | new_A6877_;
  assign new_A6862_ = new_A6885_ | new_A6884_;
  assign new_A6863_ = new_A6879_ | new_A6878_;
  assign new_A6864_ = ~new_A6887_ | ~new_A6886_;
  assign new_A6865_ = ~new_A6888_ & new_A6889_;
  assign new_A6866_ = new_A6888_ & ~new_A6889_;
  assign new_A6867_ = ~A6835 & A6836;
  assign new_A6868_ = A6835 & ~A6836;
  assign new_A6869_ = ~new_A6851_ | new_A6861_;
  assign new_A6870_ = new_A6851_ & new_A6861_;
  assign new_A6871_ = ~new_A6851_ & ~new_A6861_;
  assign new_A6872_ = new_A6893_ | new_A6892_;
  assign new_A6873_ = A6839 | new_A6872_;
  assign new_A6874_ = new_A6897_ | new_A6896_;
  assign new_A6875_ = ~A6839 & new_A6874_;
  assign new_A6876_ = new_A6895_ | new_A6894_;
  assign new_A6877_ = A6839 & new_A6876_;
  assign new_A6878_ = A6837 & ~new_A6847_;
  assign new_A6879_ = ~A6837 & new_A6847_;
  assign new_A6880_ = ~A6836 | ~new_A6861_;
  assign new_A6881_ = new_A6847_ & new_A6880_;
  assign new_A6882_ = ~new_A6847_ & ~new_A6881_;
  assign new_A6883_ = new_A6847_ | new_A6880_;
  assign new_A6884_ = ~A6837 & A6838;
  assign new_A6885_ = A6837 & ~A6838;
  assign new_A6886_ = new_A6854_ | new_A6891_;
  assign new_A6887_ = ~new_A6854_ & ~new_A6890_;
  assign new_A6888_ = A6837 | new_A6854_;
  assign new_A6889_ = A6837 | A6838;
  assign new_A6890_ = new_A6854_ & new_A6891_;
  assign new_A6891_ = ~A6836 | ~new_A6861_;
  assign new_A6892_ = new_A6869_ & new_A6889_;
  assign new_A6893_ = ~new_A6869_ & ~new_A6889_;
  assign new_A6894_ = new_A6898_ | new_A6899_;
  assign new_A6895_ = ~A6840 & new_A6854_;
  assign new_A6896_ = new_A6900_ | new_A6901_;
  assign new_A6897_ = A6840 & new_A6854_;
  assign new_A6898_ = ~A6840 & ~new_A6854_;
  assign new_A6899_ = A6840 & ~new_A6854_;
  assign new_A6900_ = A6840 & ~new_A6854_;
  assign new_A6901_ = ~A6840 & new_A6854_;
  assign new_A6908_ = new_A6915_ & new_A6914_;
  assign new_A6909_ = new_A6917_ | new_A6916_;
  assign new_A6910_ = new_A6919_ | new_A6918_;
  assign new_A6911_ = new_A6921_ & new_A6920_;
  assign new_A6912_ = new_A6921_ & new_A6922_;
  assign new_A6913_ = new_A6914_ | new_A6923_;
  assign new_A6914_ = A6903 | new_A6926_;
  assign new_A6915_ = new_A6925_ | new_A6924_;
  assign new_A6916_ = new_A6930_ & new_A6929_;
  assign new_A6917_ = new_A6928_ & new_A6927_;
  assign new_A6918_ = new_A6933_ | new_A6932_;
  assign new_A6919_ = new_A6928_ & new_A6931_;
  assign new_A6920_ = A6903 | new_A6936_;
  assign new_A6921_ = new_A6935_ | new_A6934_;
  assign new_A6922_ = new_A6938_ | new_A6937_;
  assign new_A6923_ = ~new_A6914_ & new_A6940_;
  assign new_A6924_ = ~new_A6916_ & new_A6928_;
  assign new_A6925_ = new_A6916_ & ~new_A6928_;
  assign new_A6926_ = A6902 & ~A6903;
  assign new_A6927_ = ~new_A6949_ | ~new_A6950_;
  assign new_A6928_ = new_A6942_ | new_A6944_;
  assign new_A6929_ = new_A6952_ | new_A6951_;
  assign new_A6930_ = new_A6946_ | new_A6945_;
  assign new_A6931_ = ~new_A6954_ | ~new_A6953_;
  assign new_A6932_ = ~new_A6955_ & new_A6956_;
  assign new_A6933_ = new_A6955_ & ~new_A6956_;
  assign new_A6934_ = ~A6902 & A6903;
  assign new_A6935_ = A6902 & ~A6903;
  assign new_A6936_ = ~new_A6918_ | new_A6928_;
  assign new_A6937_ = new_A6918_ & new_A6928_;
  assign new_A6938_ = ~new_A6918_ & ~new_A6928_;
  assign new_A6939_ = new_A6960_ | new_A6959_;
  assign new_A6940_ = A6906 | new_A6939_;
  assign new_A6941_ = new_A6964_ | new_A6963_;
  assign new_A6942_ = ~A6906 & new_A6941_;
  assign new_A6943_ = new_A6962_ | new_A6961_;
  assign new_A6944_ = A6906 & new_A6943_;
  assign new_A6945_ = A6904 & ~new_A6914_;
  assign new_A6946_ = ~A6904 & new_A6914_;
  assign new_A6947_ = ~A6903 | ~new_A6928_;
  assign new_A6948_ = new_A6914_ & new_A6947_;
  assign new_A6949_ = ~new_A6914_ & ~new_A6948_;
  assign new_A6950_ = new_A6914_ | new_A6947_;
  assign new_A6951_ = ~A6904 & A6905;
  assign new_A6952_ = A6904 & ~A6905;
  assign new_A6953_ = new_A6921_ | new_A6958_;
  assign new_A6954_ = ~new_A6921_ & ~new_A6957_;
  assign new_A6955_ = A6904 | new_A6921_;
  assign new_A6956_ = A6904 | A6905;
  assign new_A6957_ = new_A6921_ & new_A6958_;
  assign new_A6958_ = ~A6903 | ~new_A6928_;
  assign new_A6959_ = new_A6936_ & new_A6956_;
  assign new_A6960_ = ~new_A6936_ & ~new_A6956_;
  assign new_A6961_ = new_A6965_ | new_A6966_;
  assign new_A6962_ = ~A6907 & new_A6921_;
  assign new_A6963_ = new_A6967_ | new_A6968_;
  assign new_A6964_ = A6907 & new_A6921_;
  assign new_A6965_ = ~A6907 & ~new_A6921_;
  assign new_A6966_ = A6907 & ~new_A6921_;
  assign new_A6967_ = A6907 & ~new_A6921_;
  assign new_A6968_ = ~A6907 & new_A6921_;
  assign new_A6975_ = new_A6982_ & new_A6981_;
  assign new_A6976_ = new_A6984_ | new_A6983_;
  assign new_A6977_ = new_A6986_ | new_A6985_;
  assign new_A6978_ = new_A6988_ & new_A6987_;
  assign new_A6979_ = new_A6988_ & new_A6989_;
  assign new_A6980_ = new_A6981_ | new_A6990_;
  assign new_A6981_ = A6970 | new_A6993_;
  assign new_A6982_ = new_A6992_ | new_A6991_;
  assign new_A6983_ = new_A6997_ & new_A6996_;
  assign new_A6984_ = new_A6995_ & new_A6994_;
  assign new_A6985_ = new_A7000_ | new_A6999_;
  assign new_A6986_ = new_A6995_ & new_A6998_;
  assign new_A6987_ = A6970 | new_A7003_;
  assign new_A6988_ = new_A7002_ | new_A7001_;
  assign new_A6989_ = new_A7005_ | new_A7004_;
  assign new_A6990_ = ~new_A6981_ & new_A7007_;
  assign new_A6991_ = ~new_A6983_ & new_A6995_;
  assign new_A6992_ = new_A6983_ & ~new_A6995_;
  assign new_A6993_ = A6969 & ~A6970;
  assign new_A6994_ = ~new_A7016_ | ~new_A7017_;
  assign new_A6995_ = new_A7009_ | new_A7011_;
  assign new_A6996_ = new_A7019_ | new_A7018_;
  assign new_A6997_ = new_A7013_ | new_A7012_;
  assign new_A6998_ = ~new_A7021_ | ~new_A7020_;
  assign new_A6999_ = ~new_A7022_ & new_A7023_;
  assign new_A7000_ = new_A7022_ & ~new_A7023_;
  assign new_A7001_ = ~A6969 & A6970;
  assign new_A7002_ = A6969 & ~A6970;
  assign new_A7003_ = ~new_A6985_ | new_A6995_;
  assign new_A7004_ = new_A6985_ & new_A6995_;
  assign new_A7005_ = ~new_A6985_ & ~new_A6995_;
  assign new_A7006_ = new_A7027_ | new_A7026_;
  assign new_A7007_ = A6973 | new_A7006_;
  assign new_A7008_ = new_A7031_ | new_A7030_;
  assign new_A7009_ = ~A6973 & new_A7008_;
  assign new_A7010_ = new_A7029_ | new_A7028_;
  assign new_A7011_ = A6973 & new_A7010_;
  assign new_A7012_ = A6971 & ~new_A6981_;
  assign new_A7013_ = ~A6971 & new_A6981_;
  assign new_A7014_ = ~A6970 | ~new_A6995_;
  assign new_A7015_ = new_A6981_ & new_A7014_;
  assign new_A7016_ = ~new_A6981_ & ~new_A7015_;
  assign new_A7017_ = new_A6981_ | new_A7014_;
  assign new_A7018_ = ~A6971 & A6972;
  assign new_A7019_ = A6971 & ~A6972;
  assign new_A7020_ = new_A6988_ | new_A7025_;
  assign new_A7021_ = ~new_A6988_ & ~new_A7024_;
  assign new_A7022_ = A6971 | new_A6988_;
  assign new_A7023_ = A6971 | A6972;
  assign new_A7024_ = new_A6988_ & new_A7025_;
  assign new_A7025_ = ~A6970 | ~new_A6995_;
  assign new_A7026_ = new_A7003_ & new_A7023_;
  assign new_A7027_ = ~new_A7003_ & ~new_A7023_;
  assign new_A7028_ = new_A7032_ | new_A7033_;
  assign new_A7029_ = ~A6974 & new_A6988_;
  assign new_A7030_ = new_A7034_ | new_A7035_;
  assign new_A7031_ = A6974 & new_A6988_;
  assign new_A7032_ = ~A6974 & ~new_A6988_;
  assign new_A7033_ = A6974 & ~new_A6988_;
  assign new_A7034_ = A6974 & ~new_A6988_;
  assign new_A7035_ = ~A6974 & new_A6988_;
  assign new_A7042_ = new_A7049_ & new_A7048_;
  assign new_A7043_ = new_A7051_ | new_A7050_;
  assign new_A7044_ = new_A7053_ | new_A7052_;
  assign new_A7045_ = new_A7055_ & new_A7054_;
  assign new_A7046_ = new_A7055_ & new_A7056_;
  assign new_A7047_ = new_A7048_ | new_A7057_;
  assign new_A7048_ = A7037 | new_A7060_;
  assign new_A7049_ = new_A7059_ | new_A7058_;
  assign new_A7050_ = new_A7064_ & new_A7063_;
  assign new_A7051_ = new_A7062_ & new_A7061_;
  assign new_A7052_ = new_A7067_ | new_A7066_;
  assign new_A7053_ = new_A7062_ & new_A7065_;
  assign new_A7054_ = A7037 | new_A7070_;
  assign new_A7055_ = new_A7069_ | new_A7068_;
  assign new_A7056_ = new_A7072_ | new_A7071_;
  assign new_A7057_ = ~new_A7048_ & new_A7074_;
  assign new_A7058_ = ~new_A7050_ & new_A7062_;
  assign new_A7059_ = new_A7050_ & ~new_A7062_;
  assign new_A7060_ = A7036 & ~A7037;
  assign new_A7061_ = ~new_A7083_ | ~new_A7084_;
  assign new_A7062_ = new_A7076_ | new_A7078_;
  assign new_A7063_ = new_A7086_ | new_A7085_;
  assign new_A7064_ = new_A7080_ | new_A7079_;
  assign new_A7065_ = ~new_A7088_ | ~new_A7087_;
  assign new_A7066_ = ~new_A7089_ & new_A7090_;
  assign new_A7067_ = new_A7089_ & ~new_A7090_;
  assign new_A7068_ = ~A7036 & A7037;
  assign new_A7069_ = A7036 & ~A7037;
  assign new_A7070_ = ~new_A7052_ | new_A7062_;
  assign new_A7071_ = new_A7052_ & new_A7062_;
  assign new_A7072_ = ~new_A7052_ & ~new_A7062_;
  assign new_A7073_ = new_A7094_ | new_A7093_;
  assign new_A7074_ = A7040 | new_A7073_;
  assign new_A7075_ = new_A7098_ | new_A7097_;
  assign new_A7076_ = ~A7040 & new_A7075_;
  assign new_A7077_ = new_A7096_ | new_A7095_;
  assign new_A7078_ = A7040 & new_A7077_;
  assign new_A7079_ = A7038 & ~new_A7048_;
  assign new_A7080_ = ~A7038 & new_A7048_;
  assign new_A7081_ = ~A7037 | ~new_A7062_;
  assign new_A7082_ = new_A7048_ & new_A7081_;
  assign new_A7083_ = ~new_A7048_ & ~new_A7082_;
  assign new_A7084_ = new_A7048_ | new_A7081_;
  assign new_A7085_ = ~A7038 & A7039;
  assign new_A7086_ = A7038 & ~A7039;
  assign new_A7087_ = new_A7055_ | new_A7092_;
  assign new_A7088_ = ~new_A7055_ & ~new_A7091_;
  assign new_A7089_ = A7038 | new_A7055_;
  assign new_A7090_ = A7038 | A7039;
  assign new_A7091_ = new_A7055_ & new_A7092_;
  assign new_A7092_ = ~A7037 | ~new_A7062_;
  assign new_A7093_ = new_A7070_ & new_A7090_;
  assign new_A7094_ = ~new_A7070_ & ~new_A7090_;
  assign new_A7095_ = new_A7099_ | new_A7100_;
  assign new_A7096_ = ~A7041 & new_A7055_;
  assign new_A7097_ = new_A7101_ | new_A7102_;
  assign new_A7098_ = A7041 & new_A7055_;
  assign new_A7099_ = ~A7041 & ~new_A7055_;
  assign new_A7100_ = A7041 & ~new_A7055_;
  assign new_A7101_ = A7041 & ~new_A7055_;
  assign new_A7102_ = ~A7041 & new_A7055_;
  assign new_A7109_ = new_A7116_ & new_A7115_;
  assign new_A7110_ = new_A7118_ | new_A7117_;
  assign new_A7111_ = new_A7120_ | new_A7119_;
  assign new_A7112_ = new_A7122_ & new_A7121_;
  assign new_A7113_ = new_A7122_ & new_A7123_;
  assign new_A7114_ = new_A7115_ | new_A7124_;
  assign new_A7115_ = A7104 | new_A7127_;
  assign new_A7116_ = new_A7126_ | new_A7125_;
  assign new_A7117_ = new_A7131_ & new_A7130_;
  assign new_A7118_ = new_A7129_ & new_A7128_;
  assign new_A7119_ = new_A7134_ | new_A7133_;
  assign new_A7120_ = new_A7129_ & new_A7132_;
  assign new_A7121_ = A7104 | new_A7137_;
  assign new_A7122_ = new_A7136_ | new_A7135_;
  assign new_A7123_ = new_A7139_ | new_A7138_;
  assign new_A7124_ = ~new_A7115_ & new_A7141_;
  assign new_A7125_ = ~new_A7117_ & new_A7129_;
  assign new_A7126_ = new_A7117_ & ~new_A7129_;
  assign new_A7127_ = A7103 & ~A7104;
  assign new_A7128_ = ~new_A7150_ | ~new_A7151_;
  assign new_A7129_ = new_A7143_ | new_A7145_;
  assign new_A7130_ = new_A7153_ | new_A7152_;
  assign new_A7131_ = new_A7147_ | new_A7146_;
  assign new_A7132_ = ~new_A7155_ | ~new_A7154_;
  assign new_A7133_ = ~new_A7156_ & new_A7157_;
  assign new_A7134_ = new_A7156_ & ~new_A7157_;
  assign new_A7135_ = ~A7103 & A7104;
  assign new_A7136_ = A7103 & ~A7104;
  assign new_A7137_ = ~new_A7119_ | new_A7129_;
  assign new_A7138_ = new_A7119_ & new_A7129_;
  assign new_A7139_ = ~new_A7119_ & ~new_A7129_;
  assign new_A7140_ = new_A7161_ | new_A7160_;
  assign new_A7141_ = A7107 | new_A7140_;
  assign new_A7142_ = new_A7165_ | new_A7164_;
  assign new_A7143_ = ~A7107 & new_A7142_;
  assign new_A7144_ = new_A7163_ | new_A7162_;
  assign new_A7145_ = A7107 & new_A7144_;
  assign new_A7146_ = A7105 & ~new_A7115_;
  assign new_A7147_ = ~A7105 & new_A7115_;
  assign new_A7148_ = ~A7104 | ~new_A7129_;
  assign new_A7149_ = new_A7115_ & new_A7148_;
  assign new_A7150_ = ~new_A7115_ & ~new_A7149_;
  assign new_A7151_ = new_A7115_ | new_A7148_;
  assign new_A7152_ = ~A7105 & A7106;
  assign new_A7153_ = A7105 & ~A7106;
  assign new_A7154_ = new_A7122_ | new_A7159_;
  assign new_A7155_ = ~new_A7122_ & ~new_A7158_;
  assign new_A7156_ = A7105 | new_A7122_;
  assign new_A7157_ = A7105 | A7106;
  assign new_A7158_ = new_A7122_ & new_A7159_;
  assign new_A7159_ = ~A7104 | ~new_A7129_;
  assign new_A7160_ = new_A7137_ & new_A7157_;
  assign new_A7161_ = ~new_A7137_ & ~new_A7157_;
  assign new_A7162_ = new_A7166_ | new_A7167_;
  assign new_A7163_ = ~A7108 & new_A7122_;
  assign new_A7164_ = new_A7168_ | new_A7169_;
  assign new_A7165_ = A7108 & new_A7122_;
  assign new_A7166_ = ~A7108 & ~new_A7122_;
  assign new_A7167_ = A7108 & ~new_A7122_;
  assign new_A7168_ = A7108 & ~new_A7122_;
  assign new_A7169_ = ~A7108 & new_A7122_;
  assign new_A7176_ = new_A7183_ & new_A7182_;
  assign new_A7177_ = new_A7185_ | new_A7184_;
  assign new_A7178_ = new_A7187_ | new_A7186_;
  assign new_A7179_ = new_A7189_ & new_A7188_;
  assign new_A7180_ = new_A7189_ & new_A7190_;
  assign new_A7181_ = new_A7182_ | new_A7191_;
  assign new_A7182_ = A7171 | new_A7194_;
  assign new_A7183_ = new_A7193_ | new_A7192_;
  assign new_A7184_ = new_A7198_ & new_A7197_;
  assign new_A7185_ = new_A7196_ & new_A7195_;
  assign new_A7186_ = new_A7201_ | new_A7200_;
  assign new_A7187_ = new_A7196_ & new_A7199_;
  assign new_A7188_ = A7171 | new_A7204_;
  assign new_A7189_ = new_A7203_ | new_A7202_;
  assign new_A7190_ = new_A7206_ | new_A7205_;
  assign new_A7191_ = ~new_A7182_ & new_A7208_;
  assign new_A7192_ = ~new_A7184_ & new_A7196_;
  assign new_A7193_ = new_A7184_ & ~new_A7196_;
  assign new_A7194_ = A7170 & ~A7171;
  assign new_A7195_ = ~new_A7217_ | ~new_A7218_;
  assign new_A7196_ = new_A7210_ | new_A7212_;
  assign new_A7197_ = new_A7220_ | new_A7219_;
  assign new_A7198_ = new_A7214_ | new_A7213_;
  assign new_A7199_ = ~new_A7222_ | ~new_A7221_;
  assign new_A7200_ = ~new_A7223_ & new_A7224_;
  assign new_A7201_ = new_A7223_ & ~new_A7224_;
  assign new_A7202_ = ~A7170 & A7171;
  assign new_A7203_ = A7170 & ~A7171;
  assign new_A7204_ = ~new_A7186_ | new_A7196_;
  assign new_A7205_ = new_A7186_ & new_A7196_;
  assign new_A7206_ = ~new_A7186_ & ~new_A7196_;
  assign new_A7207_ = new_A7228_ | new_A7227_;
  assign new_A7208_ = A7174 | new_A7207_;
  assign new_A7209_ = new_A7232_ | new_A7231_;
  assign new_A7210_ = ~A7174 & new_A7209_;
  assign new_A7211_ = new_A7230_ | new_A7229_;
  assign new_A7212_ = A7174 & new_A7211_;
  assign new_A7213_ = A7172 & ~new_A7182_;
  assign new_A7214_ = ~A7172 & new_A7182_;
  assign new_A7215_ = ~A7171 | ~new_A7196_;
  assign new_A7216_ = new_A7182_ & new_A7215_;
  assign new_A7217_ = ~new_A7182_ & ~new_A7216_;
  assign new_A7218_ = new_A7182_ | new_A7215_;
  assign new_A7219_ = ~A7172 & A7173;
  assign new_A7220_ = A7172 & ~A7173;
  assign new_A7221_ = new_A7189_ | new_A7226_;
  assign new_A7222_ = ~new_A7189_ & ~new_A7225_;
  assign new_A7223_ = A7172 | new_A7189_;
  assign new_A7224_ = A7172 | A7173;
  assign new_A7225_ = new_A7189_ & new_A7226_;
  assign new_A7226_ = ~A7171 | ~new_A7196_;
  assign new_A7227_ = new_A7204_ & new_A7224_;
  assign new_A7228_ = ~new_A7204_ & ~new_A7224_;
  assign new_A7229_ = new_A7233_ | new_A7234_;
  assign new_A7230_ = ~A7175 & new_A7189_;
  assign new_A7231_ = new_A7235_ | new_A7236_;
  assign new_A7232_ = A7175 & new_A7189_;
  assign new_A7233_ = ~A7175 & ~new_A7189_;
  assign new_A7234_ = A7175 & ~new_A7189_;
  assign new_A7235_ = A7175 & ~new_A7189_;
  assign new_A7236_ = ~A7175 & new_A7189_;
  assign new_A7243_ = new_A7250_ & new_A7249_;
  assign new_A7244_ = new_A7252_ | new_A7251_;
  assign new_A7245_ = new_A7254_ | new_A7253_;
  assign new_A7246_ = new_A7256_ & new_A7255_;
  assign new_A7247_ = new_A7256_ & new_A7257_;
  assign new_A7248_ = new_A7249_ | new_A7258_;
  assign new_A7249_ = A7238 | new_A7261_;
  assign new_A7250_ = new_A7260_ | new_A7259_;
  assign new_A7251_ = new_A7265_ & new_A7264_;
  assign new_A7252_ = new_A7263_ & new_A7262_;
  assign new_A7253_ = new_A7268_ | new_A7267_;
  assign new_A7254_ = new_A7263_ & new_A7266_;
  assign new_A7255_ = A7238 | new_A7271_;
  assign new_A7256_ = new_A7270_ | new_A7269_;
  assign new_A7257_ = new_A7273_ | new_A7272_;
  assign new_A7258_ = ~new_A7249_ & new_A7275_;
  assign new_A7259_ = ~new_A7251_ & new_A7263_;
  assign new_A7260_ = new_A7251_ & ~new_A7263_;
  assign new_A7261_ = A7237 & ~A7238;
  assign new_A7262_ = ~new_A7284_ | ~new_A7285_;
  assign new_A7263_ = new_A7277_ | new_A7279_;
  assign new_A7264_ = new_A7287_ | new_A7286_;
  assign new_A7265_ = new_A7281_ | new_A7280_;
  assign new_A7266_ = ~new_A7289_ | ~new_A7288_;
  assign new_A7267_ = ~new_A7290_ & new_A7291_;
  assign new_A7268_ = new_A7290_ & ~new_A7291_;
  assign new_A7269_ = ~A7237 & A7238;
  assign new_A7270_ = A7237 & ~A7238;
  assign new_A7271_ = ~new_A7253_ | new_A7263_;
  assign new_A7272_ = new_A7253_ & new_A7263_;
  assign new_A7273_ = ~new_A7253_ & ~new_A7263_;
  assign new_A7274_ = new_A7295_ | new_A7294_;
  assign new_A7275_ = A7241 | new_A7274_;
  assign new_A7276_ = new_A7299_ | new_A7298_;
  assign new_A7277_ = ~A7241 & new_A7276_;
  assign new_A7278_ = new_A7297_ | new_A7296_;
  assign new_A7279_ = A7241 & new_A7278_;
  assign new_A7280_ = A7239 & ~new_A7249_;
  assign new_A7281_ = ~A7239 & new_A7249_;
  assign new_A7282_ = ~A7238 | ~new_A7263_;
  assign new_A7283_ = new_A7249_ & new_A7282_;
  assign new_A7284_ = ~new_A7249_ & ~new_A7283_;
  assign new_A7285_ = new_A7249_ | new_A7282_;
  assign new_A7286_ = ~A7239 & A7240;
  assign new_A7287_ = A7239 & ~A7240;
  assign new_A7288_ = new_A7256_ | new_A7293_;
  assign new_A7289_ = ~new_A7256_ & ~new_A7292_;
  assign new_A7290_ = A7239 | new_A7256_;
  assign new_A7291_ = A7239 | A7240;
  assign new_A7292_ = new_A7256_ & new_A7293_;
  assign new_A7293_ = ~A7238 | ~new_A7263_;
  assign new_A7294_ = new_A7271_ & new_A7291_;
  assign new_A7295_ = ~new_A7271_ & ~new_A7291_;
  assign new_A7296_ = new_A7300_ | new_A7301_;
  assign new_A7297_ = ~A7242 & new_A7256_;
  assign new_A7298_ = new_A7302_ | new_A7303_;
  assign new_A7299_ = A7242 & new_A7256_;
  assign new_A7300_ = ~A7242 & ~new_A7256_;
  assign new_A7301_ = A7242 & ~new_A7256_;
  assign new_A7302_ = A7242 & ~new_A7256_;
  assign new_A7303_ = ~A7242 & new_A7256_;
  assign new_A7310_ = new_A7317_ & new_A7316_;
  assign new_A7311_ = new_A7319_ | new_A7318_;
  assign new_A7312_ = new_A7321_ | new_A7320_;
  assign new_A7313_ = new_A7323_ & new_A7322_;
  assign new_A7314_ = new_A7323_ & new_A7324_;
  assign new_A7315_ = new_A7316_ | new_A7325_;
  assign new_A7316_ = A7305 | new_A7328_;
  assign new_A7317_ = new_A7327_ | new_A7326_;
  assign new_A7318_ = new_A7332_ & new_A7331_;
  assign new_A7319_ = new_A7330_ & new_A7329_;
  assign new_A7320_ = new_A7335_ | new_A7334_;
  assign new_A7321_ = new_A7330_ & new_A7333_;
  assign new_A7322_ = A7305 | new_A7338_;
  assign new_A7323_ = new_A7337_ | new_A7336_;
  assign new_A7324_ = new_A7340_ | new_A7339_;
  assign new_A7325_ = ~new_A7316_ & new_A7342_;
  assign new_A7326_ = ~new_A7318_ & new_A7330_;
  assign new_A7327_ = new_A7318_ & ~new_A7330_;
  assign new_A7328_ = A7304 & ~A7305;
  assign new_A7329_ = ~new_A7351_ | ~new_A7352_;
  assign new_A7330_ = new_A7344_ | new_A7346_;
  assign new_A7331_ = new_A7354_ | new_A7353_;
  assign new_A7332_ = new_A7348_ | new_A7347_;
  assign new_A7333_ = ~new_A7356_ | ~new_A7355_;
  assign new_A7334_ = ~new_A7357_ & new_A7358_;
  assign new_A7335_ = new_A7357_ & ~new_A7358_;
  assign new_A7336_ = ~A7304 & A7305;
  assign new_A7337_ = A7304 & ~A7305;
  assign new_A7338_ = ~new_A7320_ | new_A7330_;
  assign new_A7339_ = new_A7320_ & new_A7330_;
  assign new_A7340_ = ~new_A7320_ & ~new_A7330_;
  assign new_A7341_ = new_A7362_ | new_A7361_;
  assign new_A7342_ = A7308 | new_A7341_;
  assign new_A7343_ = new_A7366_ | new_A7365_;
  assign new_A7344_ = ~A7308 & new_A7343_;
  assign new_A7345_ = new_A7364_ | new_A7363_;
  assign new_A7346_ = A7308 & new_A7345_;
  assign new_A7347_ = A7306 & ~new_A7316_;
  assign new_A7348_ = ~A7306 & new_A7316_;
  assign new_A7349_ = ~A7305 | ~new_A7330_;
  assign new_A7350_ = new_A7316_ & new_A7349_;
  assign new_A7351_ = ~new_A7316_ & ~new_A7350_;
  assign new_A7352_ = new_A7316_ | new_A7349_;
  assign new_A7353_ = ~A7306 & A7307;
  assign new_A7354_ = A7306 & ~A7307;
  assign new_A7355_ = new_A7323_ | new_A7360_;
  assign new_A7356_ = ~new_A7323_ & ~new_A7359_;
  assign new_A7357_ = A7306 | new_A7323_;
  assign new_A7358_ = A7306 | A7307;
  assign new_A7359_ = new_A7323_ & new_A7360_;
  assign new_A7360_ = ~A7305 | ~new_A7330_;
  assign new_A7361_ = new_A7338_ & new_A7358_;
  assign new_A7362_ = ~new_A7338_ & ~new_A7358_;
  assign new_A7363_ = new_A7367_ | new_A7368_;
  assign new_A7364_ = ~A7309 & new_A7323_;
  assign new_A7365_ = new_A7369_ | new_A7370_;
  assign new_A7366_ = A7309 & new_A7323_;
  assign new_A7367_ = ~A7309 & ~new_A7323_;
  assign new_A7368_ = A7309 & ~new_A7323_;
  assign new_A7369_ = A7309 & ~new_A7323_;
  assign new_A7370_ = ~A7309 & new_A7323_;
  assign new_A7377_ = new_A7384_ & new_A7383_;
  assign new_A7378_ = new_A7386_ | new_A7385_;
  assign new_A7379_ = new_A7388_ | new_A7387_;
  assign new_A7380_ = new_A7390_ & new_A7389_;
  assign new_A7381_ = new_A7390_ & new_A7391_;
  assign new_A7382_ = new_A7383_ | new_A7392_;
  assign new_A7383_ = A7372 | new_A7395_;
  assign new_A7384_ = new_A7394_ | new_A7393_;
  assign new_A7385_ = new_A7399_ & new_A7398_;
  assign new_A7386_ = new_A7397_ & new_A7396_;
  assign new_A7387_ = new_A7402_ | new_A7401_;
  assign new_A7388_ = new_A7397_ & new_A7400_;
  assign new_A7389_ = A7372 | new_A7405_;
  assign new_A7390_ = new_A7404_ | new_A7403_;
  assign new_A7391_ = new_A7407_ | new_A7406_;
  assign new_A7392_ = ~new_A7383_ & new_A7409_;
  assign new_A7393_ = ~new_A7385_ & new_A7397_;
  assign new_A7394_ = new_A7385_ & ~new_A7397_;
  assign new_A7395_ = A7371 & ~A7372;
  assign new_A7396_ = ~new_A7418_ | ~new_A7419_;
  assign new_A7397_ = new_A7411_ | new_A7413_;
  assign new_A7398_ = new_A7421_ | new_A7420_;
  assign new_A7399_ = new_A7415_ | new_A7414_;
  assign new_A7400_ = ~new_A7423_ | ~new_A7422_;
  assign new_A7401_ = ~new_A7424_ & new_A7425_;
  assign new_A7402_ = new_A7424_ & ~new_A7425_;
  assign new_A7403_ = ~A7371 & A7372;
  assign new_A7404_ = A7371 & ~A7372;
  assign new_A7405_ = ~new_A7387_ | new_A7397_;
  assign new_A7406_ = new_A7387_ & new_A7397_;
  assign new_A7407_ = ~new_A7387_ & ~new_A7397_;
  assign new_A7408_ = new_A7429_ | new_A7428_;
  assign new_A7409_ = A7375 | new_A7408_;
  assign new_A7410_ = new_A7433_ | new_A7432_;
  assign new_A7411_ = ~A7375 & new_A7410_;
  assign new_A7412_ = new_A7431_ | new_A7430_;
  assign new_A7413_ = A7375 & new_A7412_;
  assign new_A7414_ = A7373 & ~new_A7383_;
  assign new_A7415_ = ~A7373 & new_A7383_;
  assign new_A7416_ = ~A7372 | ~new_A7397_;
  assign new_A7417_ = new_A7383_ & new_A7416_;
  assign new_A7418_ = ~new_A7383_ & ~new_A7417_;
  assign new_A7419_ = new_A7383_ | new_A7416_;
  assign new_A7420_ = ~A7373 & A7374;
  assign new_A7421_ = A7373 & ~A7374;
  assign new_A7422_ = new_A7390_ | new_A7427_;
  assign new_A7423_ = ~new_A7390_ & ~new_A7426_;
  assign new_A7424_ = A7373 | new_A7390_;
  assign new_A7425_ = A7373 | A7374;
  assign new_A7426_ = new_A7390_ & new_A7427_;
  assign new_A7427_ = ~A7372 | ~new_A7397_;
  assign new_A7428_ = new_A7405_ & new_A7425_;
  assign new_A7429_ = ~new_A7405_ & ~new_A7425_;
  assign new_A7430_ = new_A7434_ | new_A7435_;
  assign new_A7431_ = ~A7376 & new_A7390_;
  assign new_A7432_ = new_A7436_ | new_A7437_;
  assign new_A7433_ = A7376 & new_A7390_;
  assign new_A7434_ = ~A7376 & ~new_A7390_;
  assign new_A7435_ = A7376 & ~new_A7390_;
  assign new_A7436_ = A7376 & ~new_A7390_;
  assign new_A7437_ = ~A7376 & new_A7390_;
  assign new_A7444_ = new_A7451_ & new_A7450_;
  assign new_A7445_ = new_A7453_ | new_A7452_;
  assign new_A7446_ = new_A7455_ | new_A7454_;
  assign new_A7447_ = new_A7457_ & new_A7456_;
  assign new_A7448_ = new_A7457_ & new_A7458_;
  assign new_A7449_ = new_A7450_ | new_A7459_;
  assign new_A7450_ = A7439 | new_A7462_;
  assign new_A7451_ = new_A7461_ | new_A7460_;
  assign new_A7452_ = new_A7466_ & new_A7465_;
  assign new_A7453_ = new_A7464_ & new_A7463_;
  assign new_A7454_ = new_A7469_ | new_A7468_;
  assign new_A7455_ = new_A7464_ & new_A7467_;
  assign new_A7456_ = A7439 | new_A7472_;
  assign new_A7457_ = new_A7471_ | new_A7470_;
  assign new_A7458_ = new_A7474_ | new_A7473_;
  assign new_A7459_ = ~new_A7450_ & new_A7476_;
  assign new_A7460_ = ~new_A7452_ & new_A7464_;
  assign new_A7461_ = new_A7452_ & ~new_A7464_;
  assign new_A7462_ = A7438 & ~A7439;
  assign new_A7463_ = ~new_A7485_ | ~new_A7486_;
  assign new_A7464_ = new_A7478_ | new_A7480_;
  assign new_A7465_ = new_A7488_ | new_A7487_;
  assign new_A7466_ = new_A7482_ | new_A7481_;
  assign new_A7467_ = ~new_A7490_ | ~new_A7489_;
  assign new_A7468_ = ~new_A7491_ & new_A7492_;
  assign new_A7469_ = new_A7491_ & ~new_A7492_;
  assign new_A7470_ = ~A7438 & A7439;
  assign new_A7471_ = A7438 & ~A7439;
  assign new_A7472_ = ~new_A7454_ | new_A7464_;
  assign new_A7473_ = new_A7454_ & new_A7464_;
  assign new_A7474_ = ~new_A7454_ & ~new_A7464_;
  assign new_A7475_ = new_A7496_ | new_A7495_;
  assign new_A7476_ = A7442 | new_A7475_;
  assign new_A7477_ = new_A7500_ | new_A7499_;
  assign new_A7478_ = ~A7442 & new_A7477_;
  assign new_A7479_ = new_A7498_ | new_A7497_;
  assign new_A7480_ = A7442 & new_A7479_;
  assign new_A7481_ = A7440 & ~new_A7450_;
  assign new_A7482_ = ~A7440 & new_A7450_;
  assign new_A7483_ = ~A7439 | ~new_A7464_;
  assign new_A7484_ = new_A7450_ & new_A7483_;
  assign new_A7485_ = ~new_A7450_ & ~new_A7484_;
  assign new_A7486_ = new_A7450_ | new_A7483_;
  assign new_A7487_ = ~A7440 & A7441;
  assign new_A7488_ = A7440 & ~A7441;
  assign new_A7489_ = new_A7457_ | new_A7494_;
  assign new_A7490_ = ~new_A7457_ & ~new_A7493_;
  assign new_A7491_ = A7440 | new_A7457_;
  assign new_A7492_ = A7440 | A7441;
  assign new_A7493_ = new_A7457_ & new_A7494_;
  assign new_A7494_ = ~A7439 | ~new_A7464_;
  assign new_A7495_ = new_A7472_ & new_A7492_;
  assign new_A7496_ = ~new_A7472_ & ~new_A7492_;
  assign new_A7497_ = new_A7501_ | new_A7502_;
  assign new_A7498_ = ~A7443 & new_A7457_;
  assign new_A7499_ = new_A7503_ | new_A7504_;
  assign new_A7500_ = A7443 & new_A7457_;
  assign new_A7501_ = ~A7443 & ~new_A7457_;
  assign new_A7502_ = A7443 & ~new_A7457_;
  assign new_A7503_ = A7443 & ~new_A7457_;
  assign new_A7504_ = ~A7443 & new_A7457_;
  assign new_A7511_ = new_A7518_ & new_A7517_;
  assign new_A7512_ = new_A7520_ | new_A7519_;
  assign new_A7513_ = new_A7522_ | new_A7521_;
  assign new_A7514_ = new_A7524_ & new_A7523_;
  assign new_A7515_ = new_A7524_ & new_A7525_;
  assign new_A7516_ = new_A7517_ | new_A7526_;
  assign new_A7517_ = A7506 | new_A7529_;
  assign new_A7518_ = new_A7528_ | new_A7527_;
  assign new_A7519_ = new_A7533_ & new_A7532_;
  assign new_A7520_ = new_A7531_ & new_A7530_;
  assign new_A7521_ = new_A7536_ | new_A7535_;
  assign new_A7522_ = new_A7531_ & new_A7534_;
  assign new_A7523_ = A7506 | new_A7539_;
  assign new_A7524_ = new_A7538_ | new_A7537_;
  assign new_A7525_ = new_A7541_ | new_A7540_;
  assign new_A7526_ = ~new_A7517_ & new_A7543_;
  assign new_A7527_ = ~new_A7519_ & new_A7531_;
  assign new_A7528_ = new_A7519_ & ~new_A7531_;
  assign new_A7529_ = A7505 & ~A7506;
  assign new_A7530_ = ~new_A7552_ | ~new_A7553_;
  assign new_A7531_ = new_A7545_ | new_A7547_;
  assign new_A7532_ = new_A7555_ | new_A7554_;
  assign new_A7533_ = new_A7549_ | new_A7548_;
  assign new_A7534_ = ~new_A7557_ | ~new_A7556_;
  assign new_A7535_ = ~new_A7558_ & new_A7559_;
  assign new_A7536_ = new_A7558_ & ~new_A7559_;
  assign new_A7537_ = ~A7505 & A7506;
  assign new_A7538_ = A7505 & ~A7506;
  assign new_A7539_ = ~new_A7521_ | new_A7531_;
  assign new_A7540_ = new_A7521_ & new_A7531_;
  assign new_A7541_ = ~new_A7521_ & ~new_A7531_;
  assign new_A7542_ = new_A7563_ | new_A7562_;
  assign new_A7543_ = A7509 | new_A7542_;
  assign new_A7544_ = new_A7567_ | new_A7566_;
  assign new_A7545_ = ~A7509 & new_A7544_;
  assign new_A7546_ = new_A7565_ | new_A7564_;
  assign new_A7547_ = A7509 & new_A7546_;
  assign new_A7548_ = A7507 & ~new_A7517_;
  assign new_A7549_ = ~A7507 & new_A7517_;
  assign new_A7550_ = ~A7506 | ~new_A7531_;
  assign new_A7551_ = new_A7517_ & new_A7550_;
  assign new_A7552_ = ~new_A7517_ & ~new_A7551_;
  assign new_A7553_ = new_A7517_ | new_A7550_;
  assign new_A7554_ = ~A7507 & A7508;
  assign new_A7555_ = A7507 & ~A7508;
  assign new_A7556_ = new_A7524_ | new_A7561_;
  assign new_A7557_ = ~new_A7524_ & ~new_A7560_;
  assign new_A7558_ = A7507 | new_A7524_;
  assign new_A7559_ = A7507 | A7508;
  assign new_A7560_ = new_A7524_ & new_A7561_;
  assign new_A7561_ = ~A7506 | ~new_A7531_;
  assign new_A7562_ = new_A7539_ & new_A7559_;
  assign new_A7563_ = ~new_A7539_ & ~new_A7559_;
  assign new_A7564_ = new_A7568_ | new_A7569_;
  assign new_A7565_ = ~A7510 & new_A7524_;
  assign new_A7566_ = new_A7570_ | new_A7571_;
  assign new_A7567_ = A7510 & new_A7524_;
  assign new_A7568_ = ~A7510 & ~new_A7524_;
  assign new_A7569_ = A7510 & ~new_A7524_;
  assign new_A7570_ = A7510 & ~new_A7524_;
  assign new_A7571_ = ~A7510 & new_A7524_;
  assign new_A7578_ = new_A7585_ & new_A7584_;
  assign new_A7579_ = new_A7587_ | new_A7586_;
  assign new_A7580_ = new_A7589_ | new_A7588_;
  assign new_A7581_ = new_A7591_ & new_A7590_;
  assign new_A7582_ = new_A7591_ & new_A7592_;
  assign new_A7583_ = new_A7584_ | new_A7593_;
  assign new_A7584_ = A7573 | new_A7596_;
  assign new_A7585_ = new_A7595_ | new_A7594_;
  assign new_A7586_ = new_A7600_ & new_A7599_;
  assign new_A7587_ = new_A7598_ & new_A7597_;
  assign new_A7588_ = new_A7603_ | new_A7602_;
  assign new_A7589_ = new_A7598_ & new_A7601_;
  assign new_A7590_ = A7573 | new_A7606_;
  assign new_A7591_ = new_A7605_ | new_A7604_;
  assign new_A7592_ = new_A7608_ | new_A7607_;
  assign new_A7593_ = ~new_A7584_ & new_A7610_;
  assign new_A7594_ = ~new_A7586_ & new_A7598_;
  assign new_A7595_ = new_A7586_ & ~new_A7598_;
  assign new_A7596_ = A7572 & ~A7573;
  assign new_A7597_ = ~new_A7619_ | ~new_A7620_;
  assign new_A7598_ = new_A7612_ | new_A7614_;
  assign new_A7599_ = new_A7622_ | new_A7621_;
  assign new_A7600_ = new_A7616_ | new_A7615_;
  assign new_A7601_ = ~new_A7624_ | ~new_A7623_;
  assign new_A7602_ = ~new_A7625_ & new_A7626_;
  assign new_A7603_ = new_A7625_ & ~new_A7626_;
  assign new_A7604_ = ~A7572 & A7573;
  assign new_A7605_ = A7572 & ~A7573;
  assign new_A7606_ = ~new_A7588_ | new_A7598_;
  assign new_A7607_ = new_A7588_ & new_A7598_;
  assign new_A7608_ = ~new_A7588_ & ~new_A7598_;
  assign new_A7609_ = new_A7630_ | new_A7629_;
  assign new_A7610_ = A7576 | new_A7609_;
  assign new_A7611_ = new_A7634_ | new_A7633_;
  assign new_A7612_ = ~A7576 & new_A7611_;
  assign new_A7613_ = new_A7632_ | new_A7631_;
  assign new_A7614_ = A7576 & new_A7613_;
  assign new_A7615_ = A7574 & ~new_A7584_;
  assign new_A7616_ = ~A7574 & new_A7584_;
  assign new_A7617_ = ~A7573 | ~new_A7598_;
  assign new_A7618_ = new_A7584_ & new_A7617_;
  assign new_A7619_ = ~new_A7584_ & ~new_A7618_;
  assign new_A7620_ = new_A7584_ | new_A7617_;
  assign new_A7621_ = ~A7574 & A7575;
  assign new_A7622_ = A7574 & ~A7575;
  assign new_A7623_ = new_A7591_ | new_A7628_;
  assign new_A7624_ = ~new_A7591_ & ~new_A7627_;
  assign new_A7625_ = A7574 | new_A7591_;
  assign new_A7626_ = A7574 | A7575;
  assign new_A7627_ = new_A7591_ & new_A7628_;
  assign new_A7628_ = ~A7573 | ~new_A7598_;
  assign new_A7629_ = new_A7606_ & new_A7626_;
  assign new_A7630_ = ~new_A7606_ & ~new_A7626_;
  assign new_A7631_ = new_A7635_ | new_A7636_;
  assign new_A7632_ = ~A7577 & new_A7591_;
  assign new_A7633_ = new_A7637_ | new_A7638_;
  assign new_A7634_ = A7577 & new_A7591_;
  assign new_A7635_ = ~A7577 & ~new_A7591_;
  assign new_A7636_ = A7577 & ~new_A7591_;
  assign new_A7637_ = A7577 & ~new_A7591_;
  assign new_A7638_ = ~A7577 & new_A7591_;
  assign new_A7645_ = new_A7652_ & new_A7651_;
  assign new_A7646_ = new_A7654_ | new_A7653_;
  assign new_A7647_ = new_A7656_ | new_A7655_;
  assign new_A7648_ = new_A7658_ & new_A7657_;
  assign new_A7649_ = new_A7658_ & new_A7659_;
  assign new_A7650_ = new_A7651_ | new_A7660_;
  assign new_A7651_ = A7640 | new_A7663_;
  assign new_A7652_ = new_A7662_ | new_A7661_;
  assign new_A7653_ = new_A7667_ & new_A7666_;
  assign new_A7654_ = new_A7665_ & new_A7664_;
  assign new_A7655_ = new_A7670_ | new_A7669_;
  assign new_A7656_ = new_A7665_ & new_A7668_;
  assign new_A7657_ = A7640 | new_A7673_;
  assign new_A7658_ = new_A7672_ | new_A7671_;
  assign new_A7659_ = new_A7675_ | new_A7674_;
  assign new_A7660_ = ~new_A7651_ & new_A7677_;
  assign new_A7661_ = ~new_A7653_ & new_A7665_;
  assign new_A7662_ = new_A7653_ & ~new_A7665_;
  assign new_A7663_ = A7639 & ~A7640;
  assign new_A7664_ = ~new_A7686_ | ~new_A7687_;
  assign new_A7665_ = new_A7679_ | new_A7681_;
  assign new_A7666_ = new_A7689_ | new_A7688_;
  assign new_A7667_ = new_A7683_ | new_A7682_;
  assign new_A7668_ = ~new_A7691_ | ~new_A7690_;
  assign new_A7669_ = ~new_A7692_ & new_A7693_;
  assign new_A7670_ = new_A7692_ & ~new_A7693_;
  assign new_A7671_ = ~A7639 & A7640;
  assign new_A7672_ = A7639 & ~A7640;
  assign new_A7673_ = ~new_A7655_ | new_A7665_;
  assign new_A7674_ = new_A7655_ & new_A7665_;
  assign new_A7675_ = ~new_A7655_ & ~new_A7665_;
  assign new_A7676_ = new_A7697_ | new_A7696_;
  assign new_A7677_ = A7643 | new_A7676_;
  assign new_A7678_ = new_A7701_ | new_A7700_;
  assign new_A7679_ = ~A7643 & new_A7678_;
  assign new_A7680_ = new_A7699_ | new_A7698_;
  assign new_A7681_ = A7643 & new_A7680_;
  assign new_A7682_ = A7641 & ~new_A7651_;
  assign new_A7683_ = ~A7641 & new_A7651_;
  assign new_A7684_ = ~A7640 | ~new_A7665_;
  assign new_A7685_ = new_A7651_ & new_A7684_;
  assign new_A7686_ = ~new_A7651_ & ~new_A7685_;
  assign new_A7687_ = new_A7651_ | new_A7684_;
  assign new_A7688_ = ~A7641 & A7642;
  assign new_A7689_ = A7641 & ~A7642;
  assign new_A7690_ = new_A7658_ | new_A7695_;
  assign new_A7691_ = ~new_A7658_ & ~new_A7694_;
  assign new_A7692_ = A7641 | new_A7658_;
  assign new_A7693_ = A7641 | A7642;
  assign new_A7694_ = new_A7658_ & new_A7695_;
  assign new_A7695_ = ~A7640 | ~new_A7665_;
  assign new_A7696_ = new_A7673_ & new_A7693_;
  assign new_A7697_ = ~new_A7673_ & ~new_A7693_;
  assign new_A7698_ = new_A7702_ | new_A7703_;
  assign new_A7699_ = ~A7644 & new_A7658_;
  assign new_A7700_ = new_A7704_ | new_A7705_;
  assign new_A7701_ = A7644 & new_A7658_;
  assign new_A7702_ = ~A7644 & ~new_A7658_;
  assign new_A7703_ = A7644 & ~new_A7658_;
  assign new_A7704_ = A7644 & ~new_A7658_;
  assign new_A7705_ = ~A7644 & new_A7658_;
  assign new_A7712_ = new_A7719_ & new_A7718_;
  assign new_A7713_ = new_A7721_ | new_A7720_;
  assign new_A7714_ = new_A7723_ | new_A7722_;
  assign new_A7715_ = new_A7725_ & new_A7724_;
  assign new_A7716_ = new_A7725_ & new_A7726_;
  assign new_A7717_ = new_A7718_ | new_A7727_;
  assign new_A7718_ = A7707 | new_A7730_;
  assign new_A7719_ = new_A7729_ | new_A7728_;
  assign new_A7720_ = new_A7734_ & new_A7733_;
  assign new_A7721_ = new_A7732_ & new_A7731_;
  assign new_A7722_ = new_A7737_ | new_A7736_;
  assign new_A7723_ = new_A7732_ & new_A7735_;
  assign new_A7724_ = A7707 | new_A7740_;
  assign new_A7725_ = new_A7739_ | new_A7738_;
  assign new_A7726_ = new_A7742_ | new_A7741_;
  assign new_A7727_ = ~new_A7718_ & new_A7744_;
  assign new_A7728_ = ~new_A7720_ & new_A7732_;
  assign new_A7729_ = new_A7720_ & ~new_A7732_;
  assign new_A7730_ = A7706 & ~A7707;
  assign new_A7731_ = ~new_A7753_ | ~new_A7754_;
  assign new_A7732_ = new_A7746_ | new_A7748_;
  assign new_A7733_ = new_A7756_ | new_A7755_;
  assign new_A7734_ = new_A7750_ | new_A7749_;
  assign new_A7735_ = ~new_A7758_ | ~new_A7757_;
  assign new_A7736_ = ~new_A7759_ & new_A7760_;
  assign new_A7737_ = new_A7759_ & ~new_A7760_;
  assign new_A7738_ = ~A7706 & A7707;
  assign new_A7739_ = A7706 & ~A7707;
  assign new_A7740_ = ~new_A7722_ | new_A7732_;
  assign new_A7741_ = new_A7722_ & new_A7732_;
  assign new_A7742_ = ~new_A7722_ & ~new_A7732_;
  assign new_A7743_ = new_A7764_ | new_A7763_;
  assign new_A7744_ = A7710 | new_A7743_;
  assign new_A7745_ = new_A7768_ | new_A7767_;
  assign new_A7746_ = ~A7710 & new_A7745_;
  assign new_A7747_ = new_A7766_ | new_A7765_;
  assign new_A7748_ = A7710 & new_A7747_;
  assign new_A7749_ = A7708 & ~new_A7718_;
  assign new_A7750_ = ~A7708 & new_A7718_;
  assign new_A7751_ = ~A7707 | ~new_A7732_;
  assign new_A7752_ = new_A7718_ & new_A7751_;
  assign new_A7753_ = ~new_A7718_ & ~new_A7752_;
  assign new_A7754_ = new_A7718_ | new_A7751_;
  assign new_A7755_ = ~A7708 & A7709;
  assign new_A7756_ = A7708 & ~A7709;
  assign new_A7757_ = new_A7725_ | new_A7762_;
  assign new_A7758_ = ~new_A7725_ & ~new_A7761_;
  assign new_A7759_ = A7708 | new_A7725_;
  assign new_A7760_ = A7708 | A7709;
  assign new_A7761_ = new_A7725_ & new_A7762_;
  assign new_A7762_ = ~A7707 | ~new_A7732_;
  assign new_A7763_ = new_A7740_ & new_A7760_;
  assign new_A7764_ = ~new_A7740_ & ~new_A7760_;
  assign new_A7765_ = new_A7769_ | new_A7770_;
  assign new_A7766_ = ~A7711 & new_A7725_;
  assign new_A7767_ = new_A7771_ | new_A7772_;
  assign new_A7768_ = A7711 & new_A7725_;
  assign new_A7769_ = ~A7711 & ~new_A7725_;
  assign new_A7770_ = A7711 & ~new_A7725_;
  assign new_A7771_ = A7711 & ~new_A7725_;
  assign new_A7772_ = ~A7711 & new_A7725_;
  assign new_A7779_ = new_A7786_ & new_A7785_;
  assign new_A7780_ = new_A7788_ | new_A7787_;
  assign new_A7781_ = new_A7790_ | new_A7789_;
  assign new_A7782_ = new_A7792_ & new_A7791_;
  assign new_A7783_ = new_A7792_ & new_A7793_;
  assign new_A7784_ = new_A7785_ | new_A7794_;
  assign new_A7785_ = A7774 | new_A7797_;
  assign new_A7786_ = new_A7796_ | new_A7795_;
  assign new_A7787_ = new_A7801_ & new_A7800_;
  assign new_A7788_ = new_A7799_ & new_A7798_;
  assign new_A7789_ = new_A7804_ | new_A7803_;
  assign new_A7790_ = new_A7799_ & new_A7802_;
  assign new_A7791_ = A7774 | new_A7807_;
  assign new_A7792_ = new_A7806_ | new_A7805_;
  assign new_A7793_ = new_A7809_ | new_A7808_;
  assign new_A7794_ = ~new_A7785_ & new_A7811_;
  assign new_A7795_ = ~new_A7787_ & new_A7799_;
  assign new_A7796_ = new_A7787_ & ~new_A7799_;
  assign new_A7797_ = A7773 & ~A7774;
  assign new_A7798_ = ~new_A7820_ | ~new_A7821_;
  assign new_A7799_ = new_A7813_ | new_A7815_;
  assign new_A7800_ = new_A7823_ | new_A7822_;
  assign new_A7801_ = new_A7817_ | new_A7816_;
  assign new_A7802_ = ~new_A7825_ | ~new_A7824_;
  assign new_A7803_ = ~new_A7826_ & new_A7827_;
  assign new_A7804_ = new_A7826_ & ~new_A7827_;
  assign new_A7805_ = ~A7773 & A7774;
  assign new_A7806_ = A7773 & ~A7774;
  assign new_A7807_ = ~new_A7789_ | new_A7799_;
  assign new_A7808_ = new_A7789_ & new_A7799_;
  assign new_A7809_ = ~new_A7789_ & ~new_A7799_;
  assign new_A7810_ = new_A7831_ | new_A7830_;
  assign new_A7811_ = A7777 | new_A7810_;
  assign new_A7812_ = new_A7835_ | new_A7834_;
  assign new_A7813_ = ~A7777 & new_A7812_;
  assign new_A7814_ = new_A7833_ | new_A7832_;
  assign new_A7815_ = A7777 & new_A7814_;
  assign new_A7816_ = A7775 & ~new_A7785_;
  assign new_A7817_ = ~A7775 & new_A7785_;
  assign new_A7818_ = ~A7774 | ~new_A7799_;
  assign new_A7819_ = new_A7785_ & new_A7818_;
  assign new_A7820_ = ~new_A7785_ & ~new_A7819_;
  assign new_A7821_ = new_A7785_ | new_A7818_;
  assign new_A7822_ = ~A7775 & A7776;
  assign new_A7823_ = A7775 & ~A7776;
  assign new_A7824_ = new_A7792_ | new_A7829_;
  assign new_A7825_ = ~new_A7792_ & ~new_A7828_;
  assign new_A7826_ = A7775 | new_A7792_;
  assign new_A7827_ = A7775 | A7776;
  assign new_A7828_ = new_A7792_ & new_A7829_;
  assign new_A7829_ = ~A7774 | ~new_A7799_;
  assign new_A7830_ = new_A7807_ & new_A7827_;
  assign new_A7831_ = ~new_A7807_ & ~new_A7827_;
  assign new_A7832_ = new_A7836_ | new_A7837_;
  assign new_A7833_ = ~A7778 & new_A7792_;
  assign new_A7834_ = new_A7838_ | new_A7839_;
  assign new_A7835_ = A7778 & new_A7792_;
  assign new_A7836_ = ~A7778 & ~new_A7792_;
  assign new_A7837_ = A7778 & ~new_A7792_;
  assign new_A7838_ = A7778 & ~new_A7792_;
  assign new_A7839_ = ~A7778 & new_A7792_;
  assign new_A7846_ = new_A7853_ & new_A7852_;
  assign new_A7847_ = new_A7855_ | new_A7854_;
  assign new_A7848_ = new_A7857_ | new_A7856_;
  assign new_A7849_ = new_A7859_ & new_A7858_;
  assign new_A7850_ = new_A7859_ & new_A7860_;
  assign new_A7851_ = new_A7852_ | new_A7861_;
  assign new_A7852_ = A7841 | new_A7864_;
  assign new_A7853_ = new_A7863_ | new_A7862_;
  assign new_A7854_ = new_A7868_ & new_A7867_;
  assign new_A7855_ = new_A7866_ & new_A7865_;
  assign new_A7856_ = new_A7871_ | new_A7870_;
  assign new_A7857_ = new_A7866_ & new_A7869_;
  assign new_A7858_ = A7841 | new_A7874_;
  assign new_A7859_ = new_A7873_ | new_A7872_;
  assign new_A7860_ = new_A7876_ | new_A7875_;
  assign new_A7861_ = ~new_A7852_ & new_A7878_;
  assign new_A7862_ = ~new_A7854_ & new_A7866_;
  assign new_A7863_ = new_A7854_ & ~new_A7866_;
  assign new_A7864_ = A7840 & ~A7841;
  assign new_A7865_ = ~new_A7887_ | ~new_A7888_;
  assign new_A7866_ = new_A7880_ | new_A7882_;
  assign new_A7867_ = new_A7890_ | new_A7889_;
  assign new_A7868_ = new_A7884_ | new_A7883_;
  assign new_A7869_ = ~new_A7892_ | ~new_A7891_;
  assign new_A7870_ = ~new_A7893_ & new_A7894_;
  assign new_A7871_ = new_A7893_ & ~new_A7894_;
  assign new_A7872_ = ~A7840 & A7841;
  assign new_A7873_ = A7840 & ~A7841;
  assign new_A7874_ = ~new_A7856_ | new_A7866_;
  assign new_A7875_ = new_A7856_ & new_A7866_;
  assign new_A7876_ = ~new_A7856_ & ~new_A7866_;
  assign new_A7877_ = new_A7898_ | new_A7897_;
  assign new_A7878_ = A7844 | new_A7877_;
  assign new_A7879_ = new_A7902_ | new_A7901_;
  assign new_A7880_ = ~A7844 & new_A7879_;
  assign new_A7881_ = new_A7900_ | new_A7899_;
  assign new_A7882_ = A7844 & new_A7881_;
  assign new_A7883_ = A7842 & ~new_A7852_;
  assign new_A7884_ = ~A7842 & new_A7852_;
  assign new_A7885_ = ~A7841 | ~new_A7866_;
  assign new_A7886_ = new_A7852_ & new_A7885_;
  assign new_A7887_ = ~new_A7852_ & ~new_A7886_;
  assign new_A7888_ = new_A7852_ | new_A7885_;
  assign new_A7889_ = ~A7842 & A7843;
  assign new_A7890_ = A7842 & ~A7843;
  assign new_A7891_ = new_A7859_ | new_A7896_;
  assign new_A7892_ = ~new_A7859_ & ~new_A7895_;
  assign new_A7893_ = A7842 | new_A7859_;
  assign new_A7894_ = A7842 | A7843;
  assign new_A7895_ = new_A7859_ & new_A7896_;
  assign new_A7896_ = ~A7841 | ~new_A7866_;
  assign new_A7897_ = new_A7874_ & new_A7894_;
  assign new_A7898_ = ~new_A7874_ & ~new_A7894_;
  assign new_A7899_ = new_A7903_ | new_A7904_;
  assign new_A7900_ = ~A7845 & new_A7859_;
  assign new_A7901_ = new_A7905_ | new_A7906_;
  assign new_A7902_ = A7845 & new_A7859_;
  assign new_A7903_ = ~A7845 & ~new_A7859_;
  assign new_A7904_ = A7845 & ~new_A7859_;
  assign new_A7905_ = A7845 & ~new_A7859_;
  assign new_A7906_ = ~A7845 & new_A7859_;
  assign new_A7913_ = new_A7920_ & new_A7919_;
  assign new_A7914_ = new_A7922_ | new_A7921_;
  assign new_A7915_ = new_A7924_ | new_A7923_;
  assign new_A7916_ = new_A7926_ & new_A7925_;
  assign new_A7917_ = new_A7926_ & new_A7927_;
  assign new_A7918_ = new_A7919_ | new_A7928_;
  assign new_A7919_ = A7908 | new_A7931_;
  assign new_A7920_ = new_A7930_ | new_A7929_;
  assign new_A7921_ = new_A7935_ & new_A7934_;
  assign new_A7922_ = new_A7933_ & new_A7932_;
  assign new_A7923_ = new_A7938_ | new_A7937_;
  assign new_A7924_ = new_A7933_ & new_A7936_;
  assign new_A7925_ = A7908 | new_A7941_;
  assign new_A7926_ = new_A7940_ | new_A7939_;
  assign new_A7927_ = new_A7943_ | new_A7942_;
  assign new_A7928_ = ~new_A7919_ & new_A7945_;
  assign new_A7929_ = ~new_A7921_ & new_A7933_;
  assign new_A7930_ = new_A7921_ & ~new_A7933_;
  assign new_A7931_ = A7907 & ~A7908;
  assign new_A7932_ = ~new_A7954_ | ~new_A7955_;
  assign new_A7933_ = new_A7947_ | new_A7949_;
  assign new_A7934_ = new_A7957_ | new_A7956_;
  assign new_A7935_ = new_A7951_ | new_A7950_;
  assign new_A7936_ = ~new_A7959_ | ~new_A7958_;
  assign new_A7937_ = ~new_A7960_ & new_A7961_;
  assign new_A7938_ = new_A7960_ & ~new_A7961_;
  assign new_A7939_ = ~A7907 & A7908;
  assign new_A7940_ = A7907 & ~A7908;
  assign new_A7941_ = ~new_A7923_ | new_A7933_;
  assign new_A7942_ = new_A7923_ & new_A7933_;
  assign new_A7943_ = ~new_A7923_ & ~new_A7933_;
  assign new_A7944_ = new_A7965_ | new_A7964_;
  assign new_A7945_ = A7911 | new_A7944_;
  assign new_A7946_ = new_A7969_ | new_A7968_;
  assign new_A7947_ = ~A7911 & new_A7946_;
  assign new_A7948_ = new_A7967_ | new_A7966_;
  assign new_A7949_ = A7911 & new_A7948_;
  assign new_A7950_ = A7909 & ~new_A7919_;
  assign new_A7951_ = ~A7909 & new_A7919_;
  assign new_A7952_ = ~A7908 | ~new_A7933_;
  assign new_A7953_ = new_A7919_ & new_A7952_;
  assign new_A7954_ = ~new_A7919_ & ~new_A7953_;
  assign new_A7955_ = new_A7919_ | new_A7952_;
  assign new_A7956_ = ~A7909 & A7910;
  assign new_A7957_ = A7909 & ~A7910;
  assign new_A7958_ = new_A7926_ | new_A7963_;
  assign new_A7959_ = ~new_A7926_ & ~new_A7962_;
  assign new_A7960_ = A7909 | new_A7926_;
  assign new_A7961_ = A7909 | A7910;
  assign new_A7962_ = new_A7926_ & new_A7963_;
  assign new_A7963_ = ~A7908 | ~new_A7933_;
  assign new_A7964_ = new_A7941_ & new_A7961_;
  assign new_A7965_ = ~new_A7941_ & ~new_A7961_;
  assign new_A7966_ = new_A7970_ | new_A7971_;
  assign new_A7967_ = ~A7912 & new_A7926_;
  assign new_A7968_ = new_A7972_ | new_A7973_;
  assign new_A7969_ = A7912 & new_A7926_;
  assign new_A7970_ = ~A7912 & ~new_A7926_;
  assign new_A7971_ = A7912 & ~new_A7926_;
  assign new_A7972_ = A7912 & ~new_A7926_;
  assign new_A7973_ = ~A7912 & new_A7926_;
  assign new_A7980_ = new_A7987_ & new_A7986_;
  assign new_A7981_ = new_A7989_ | new_A7988_;
  assign new_A7982_ = new_A7991_ | new_A7990_;
  assign new_A7983_ = new_A7993_ & new_A7992_;
  assign new_A7984_ = new_A7993_ & new_A7994_;
  assign new_A7985_ = new_A7986_ | new_A7995_;
  assign new_A7986_ = A7975 | new_A7998_;
  assign new_A7987_ = new_A7997_ | new_A7996_;
  assign new_A7988_ = new_A8002_ & new_A8001_;
  assign new_A7989_ = new_A8000_ & new_A7999_;
  assign new_A7990_ = new_A8005_ | new_A8004_;
  assign new_A7991_ = new_A8000_ & new_A8003_;
  assign new_A7992_ = A7975 | new_A8008_;
  assign new_A7993_ = new_A8007_ | new_A8006_;
  assign new_A7994_ = new_A8010_ | new_A8009_;
  assign new_A7995_ = ~new_A7986_ & new_A8012_;
  assign new_A7996_ = ~new_A7988_ & new_A8000_;
  assign new_A7997_ = new_A7988_ & ~new_A8000_;
  assign new_A7998_ = A7974 & ~A7975;
  assign new_A7999_ = ~new_A8021_ | ~new_A8022_;
  assign new_A8000_ = new_A8014_ | new_A8016_;
  assign new_A8001_ = new_A8024_ | new_A8023_;
  assign new_A8002_ = new_A8018_ | new_A8017_;
  assign new_A8003_ = ~new_A8026_ | ~new_A8025_;
  assign new_A8004_ = ~new_A8027_ & new_A8028_;
  assign new_A8005_ = new_A8027_ & ~new_A8028_;
  assign new_A8006_ = ~A7974 & A7975;
  assign new_A8007_ = A7974 & ~A7975;
  assign new_A8008_ = ~new_A7990_ | new_A8000_;
  assign new_A8009_ = new_A7990_ & new_A8000_;
  assign new_A8010_ = ~new_A7990_ & ~new_A8000_;
  assign new_A8011_ = new_A8032_ | new_A8031_;
  assign new_A8012_ = A7978 | new_A8011_;
  assign new_A8013_ = new_A8036_ | new_A8035_;
  assign new_A8014_ = ~A7978 & new_A8013_;
  assign new_A8015_ = new_A8034_ | new_A8033_;
  assign new_A8016_ = A7978 & new_A8015_;
  assign new_A8017_ = A7976 & ~new_A7986_;
  assign new_A8018_ = ~A7976 & new_A7986_;
  assign new_A8019_ = ~A7975 | ~new_A8000_;
  assign new_A8020_ = new_A7986_ & new_A8019_;
  assign new_A8021_ = ~new_A7986_ & ~new_A8020_;
  assign new_A8022_ = new_A7986_ | new_A8019_;
  assign new_A8023_ = ~A7976 & A7977;
  assign new_A8024_ = A7976 & ~A7977;
  assign new_A8025_ = new_A7993_ | new_A8030_;
  assign new_A8026_ = ~new_A7993_ & ~new_A8029_;
  assign new_A8027_ = A7976 | new_A7993_;
  assign new_A8028_ = A7976 | A7977;
  assign new_A8029_ = new_A7993_ & new_A8030_;
  assign new_A8030_ = ~A7975 | ~new_A8000_;
  assign new_A8031_ = new_A8008_ & new_A8028_;
  assign new_A8032_ = ~new_A8008_ & ~new_A8028_;
  assign new_A8033_ = new_A8037_ | new_A8038_;
  assign new_A8034_ = ~A7979 & new_A7993_;
  assign new_A8035_ = new_A8039_ | new_A8040_;
  assign new_A8036_ = A7979 & new_A7993_;
  assign new_A8037_ = ~A7979 & ~new_A7993_;
  assign new_A8038_ = A7979 & ~new_A7993_;
  assign new_A8039_ = A7979 & ~new_A7993_;
  assign new_A8040_ = ~A7979 & new_A7993_;
  assign new_A3283_ = ~new_A3222_ & new_A3236_;
  assign new_A3282_ = new_A3222_ & ~new_A3236_;
  assign new_A3281_ = new_A3222_ & ~new_A3236_;
  assign new_A3280_ = ~new_A3222_ & ~new_A3236_;
  assign new_A3279_ = new_A3222_ & new_A3236_;
  assign new_A3278_ = new_A3282_ | new_A3283_;
  assign new_A3277_ = ~new_A3222_ & new_A3236_;
  assign new_A3276_ = new_A3280_ | new_A3281_;
  assign new_A3275_ = ~new_A3251_ & ~new_A3271_;
  assign new_A3274_ = new_A3251_ & new_A3271_;
  assign new_A3273_ = ~new_A3218_ | ~new_A3243_;
  assign new_A3272_ = new_A3236_ & new_A3273_;
  assign new_A3271_ = new_A3219_ | new_A3220_;
  assign new_A3270_ = new_A3219_ | new_A3236_;
  assign new_A3269_ = ~new_A3236_ & ~new_A3272_;
  assign new_A3268_ = new_A3236_ | new_A3273_;
  assign new_A3267_ = new_A3219_ & ~new_A3220_;
  assign new_A3266_ = ~new_A3219_ & new_A3220_;
  assign new_A3265_ = new_A3229_ | new_A3262_;
  assign new_A3264_ = ~new_A3229_ & ~new_A3263_;
  assign new_A3263_ = new_A3229_ & new_A3262_;
  assign new_A3262_ = ~new_A3218_ | ~new_A3243_;
  assign new_A3261_ = ~new_A3219_ & new_A3229_;
  assign new_A3260_ = new_A3219_ & ~new_A3229_;
  assign new_A3259_ = new_A3221_ & new_A3258_;
  assign new_A3258_ = new_A3277_ | new_A3276_;
  assign new_A3257_ = ~new_A3221_ & new_A3256_;
  assign new_A3256_ = new_A3279_ | new_A3278_;
  assign new_A3255_ = new_A3221_ | new_A3254_;
  assign new_A3254_ = new_A3275_ | new_A3274_;
  assign new_A3253_ = ~new_A3233_ & ~new_A3243_;
  assign new_A3252_ = new_A3233_ & new_A3243_;
  assign new_A3251_ = ~new_A3233_ | new_A3243_;
  assign new_A3250_ = new_A3217_ & ~new_A3218_;
  assign new_A3249_ = ~new_A3217_ & new_A3218_;
  assign new_A3248_ = new_A3270_ & ~new_A3271_;
  assign new_A3247_ = ~new_A3270_ & new_A3271_;
  assign new_A3246_ = ~new_A3269_ | ~new_A3268_;
  assign new_A3245_ = new_A3261_ | new_A3260_;
  assign new_A3244_ = new_A3267_ | new_A3266_;
  assign new_A3243_ = new_A3257_ | new_A3259_;
  assign new_A3242_ = ~new_A3264_ | ~new_A3265_;
  assign new_A3241_ = new_A3217_ & ~new_A3218_;
  assign new_A3240_ = new_A3231_ & ~new_A3243_;
  assign new_A3239_ = ~new_A3231_ & new_A3243_;
  assign new_A3238_ = ~new_A3229_ & new_A3255_;
  assign new_A3237_ = new_A3253_ | new_A3252_;
  assign new_A3236_ = new_A3250_ | new_A3249_;
  assign new_A3235_ = new_A3218_ | new_A3251_;
  assign new_A3234_ = new_A3243_ & new_A3246_;
  assign new_A3233_ = new_A3248_ | new_A3247_;
  assign new_A3232_ = new_A3243_ & new_A3242_;
  assign new_A3231_ = new_A3245_ & new_A3244_;
  assign new_A3230_ = new_A3240_ | new_A3239_;
  assign new_A3229_ = new_A3218_ | new_A3241_;
  assign new_A3228_ = new_A3229_ | new_A3238_;
  assign new_A3227_ = new_A3236_ & new_A3237_;
  assign new_A3226_ = new_A3236_ & new_A3235_;
  assign new_A3225_ = new_A3234_ | new_A3233_;
  assign new_A3224_ = new_A3232_ | new_A3231_;
  assign new_A3223_ = new_A3230_ & new_A3229_;
  assign new_A3222_ = new_A5640_;
  assign new_A3221_ = new_A5702_;
  assign new_A3220_ = new_A5769_;
  assign new_A3219_ = new_A5836_;
  assign new_A3218_ = new_A5903_;
  assign new_A3217_ = new_A5970_;
  assign new_A3284_ = new_A6037_;
  assign new_A3285_ = new_A6104_;
  assign new_A3286_ = new_A6171_;
  assign new_A3287_ = new_A6238_;
  assign new_A3288_ = new_A6305_;
  assign new_A3289_ = new_A6372_;
  assign new_A3290_ = new_A3297_ & new_A3296_;
  assign new_A3291_ = new_A3299_ | new_A3298_;
  assign new_A3292_ = new_A3301_ | new_A3300_;
  assign new_A3293_ = new_A3303_ & new_A3302_;
  assign new_A3294_ = new_A3303_ & new_A3304_;
  assign new_A3295_ = new_A3296_ | new_A3305_;
  assign new_A3296_ = new_A3285_ | new_A3308_;
  assign new_A3297_ = new_A3307_ | new_A3306_;
  assign new_A3298_ = new_A3312_ & new_A3311_;
  assign new_A3299_ = new_A3310_ & new_A3309_;
  assign new_A3300_ = new_A3315_ | new_A3314_;
  assign new_A3301_ = new_A3310_ & new_A3313_;
  assign new_A3302_ = new_A3285_ | new_A3318_;
  assign new_A3303_ = new_A3317_ | new_A3316_;
  assign new_A3304_ = new_A3320_ | new_A3319_;
  assign new_A3305_ = ~new_A3296_ & new_A3322_;
  assign new_A3306_ = ~new_A3298_ & new_A3310_;
  assign new_A3307_ = new_A3298_ & ~new_A3310_;
  assign new_A3308_ = new_A3284_ & ~new_A3285_;
  assign new_A3309_ = ~new_A3331_ | ~new_A3332_;
  assign new_A3310_ = new_A3324_ | new_A3326_;
  assign new_A3311_ = new_A3334_ | new_A3333_;
  assign new_A3312_ = new_A3328_ | new_A3327_;
  assign new_A3313_ = ~new_A3336_ | ~new_A3335_;
  assign new_A3314_ = ~new_A3337_ & new_A3338_;
  assign new_A3315_ = new_A3337_ & ~new_A3338_;
  assign new_A3316_ = ~new_A3284_ & new_A3285_;
  assign new_A3317_ = new_A3284_ & ~new_A3285_;
  assign new_A3318_ = ~new_A3300_ | new_A3310_;
  assign new_A3319_ = new_A3300_ & new_A3310_;
  assign new_A3320_ = ~new_A3300_ & ~new_A3310_;
  assign new_A3321_ = new_A3342_ | new_A3341_;
  assign new_A3322_ = new_A3288_ | new_A3321_;
  assign new_A3323_ = new_A3346_ | new_A3345_;
  assign new_A3324_ = ~new_A3288_ & new_A3323_;
  assign new_A3325_ = new_A3344_ | new_A3343_;
  assign new_A3326_ = new_A3288_ & new_A3325_;
  assign new_A3327_ = new_A3286_ & ~new_A3296_;
  assign new_A3328_ = ~new_A3286_ & new_A3296_;
  assign new_A3329_ = ~new_A3285_ | ~new_A3310_;
  assign new_A3330_ = new_A3296_ & new_A3329_;
  assign new_A3331_ = ~new_A3296_ & ~new_A3330_;
  assign new_A3332_ = new_A3296_ | new_A3329_;
  assign new_A3333_ = ~new_A3286_ & new_A3287_;
  assign new_A3334_ = new_A3286_ & ~new_A3287_;
  assign new_A3335_ = new_A3303_ | new_A3340_;
  assign new_A3336_ = ~new_A3303_ & ~new_A3339_;
  assign new_A3337_ = new_A3286_ | new_A3303_;
  assign new_A3338_ = new_A3286_ | new_A3287_;
  assign new_A3339_ = new_A3303_ & new_A3340_;
  assign new_A3340_ = ~new_A3285_ | ~new_A3310_;
  assign new_A3341_ = new_A3318_ & new_A3338_;
  assign new_A3342_ = ~new_A3318_ & ~new_A3338_;
  assign new_A3343_ = new_A3347_ | new_A3348_;
  assign new_A3344_ = ~new_A3289_ & new_A3303_;
  assign new_A3345_ = new_A3349_ | new_A3350_;
  assign new_A3346_ = new_A3289_ & new_A3303_;
  assign new_A3347_ = ~new_A3289_ & ~new_A3303_;
  assign new_A3348_ = new_A3289_ & ~new_A3303_;
  assign new_A3349_ = new_A3289_ & ~new_A3303_;
  assign new_A3350_ = ~new_A3289_ & new_A3303_;
  assign new_A3351_ = new_A6439_;
  assign new_A3352_ = new_A6506_;
  assign new_A3353_ = new_A6573_;
  assign new_A3354_ = new_A6640_;
  assign new_A3355_ = new_A6707_;
  assign new_A3356_ = new_A6774_;
  assign new_A3357_ = new_A3364_ & new_A3363_;
  assign new_A3358_ = new_A3366_ | new_A3365_;
  assign new_A3359_ = new_A3368_ | new_A3367_;
  assign new_A3360_ = new_A3370_ & new_A3369_;
  assign new_A3361_ = new_A3370_ & new_A3371_;
  assign new_A3362_ = new_A3363_ | new_A3372_;
  assign new_A3363_ = new_A3352_ | new_A3375_;
  assign new_A3364_ = new_A3374_ | new_A3373_;
  assign new_A3365_ = new_A3379_ & new_A3378_;
  assign new_A3366_ = new_A3377_ & new_A3376_;
  assign new_A3367_ = new_A3382_ | new_A3381_;
  assign new_A3368_ = new_A3377_ & new_A3380_;
  assign new_A3369_ = new_A3352_ | new_A3385_;
  assign new_A3370_ = new_A3384_ | new_A3383_;
  assign new_A3371_ = new_A3387_ | new_A3386_;
  assign new_A3372_ = ~new_A3363_ & new_A3389_;
  assign new_A3373_ = ~new_A3365_ & new_A3377_;
  assign new_A3374_ = new_A3365_ & ~new_A3377_;
  assign new_A3375_ = new_A3351_ & ~new_A3352_;
  assign new_A3376_ = ~new_A3398_ | ~new_A3399_;
  assign new_A3377_ = new_A3391_ | new_A3393_;
  assign new_A3378_ = new_A3401_ | new_A3400_;
  assign new_A3379_ = new_A3395_ | new_A3394_;
  assign new_A3380_ = ~new_A3403_ | ~new_A3402_;
  assign new_A3381_ = ~new_A3404_ & new_A3405_;
  assign new_A3382_ = new_A3404_ & ~new_A3405_;
  assign new_A3383_ = ~new_A3351_ & new_A3352_;
  assign new_A3384_ = new_A3351_ & ~new_A3352_;
  assign new_A3385_ = ~new_A3367_ | new_A3377_;
  assign new_A3386_ = new_A3367_ & new_A3377_;
  assign new_A3387_ = ~new_A3367_ & ~new_A3377_;
  assign new_A3388_ = new_A3409_ | new_A3408_;
  assign new_A3389_ = new_A3355_ | new_A3388_;
  assign new_A3390_ = new_A3413_ | new_A3412_;
  assign new_A3391_ = ~new_A3355_ & new_A3390_;
  assign new_A3392_ = new_A3411_ | new_A3410_;
  assign new_A3393_ = new_A3355_ & new_A3392_;
  assign new_A3394_ = new_A3353_ & ~new_A3363_;
  assign new_A3395_ = ~new_A3353_ & new_A3363_;
  assign new_A3396_ = ~new_A3352_ | ~new_A3377_;
  assign new_A3397_ = new_A3363_ & new_A3396_;
  assign new_A3398_ = ~new_A3363_ & ~new_A3397_;
  assign new_A3399_ = new_A3363_ | new_A3396_;
  assign new_A3400_ = ~new_A3353_ & new_A3354_;
  assign new_A3401_ = new_A3353_ & ~new_A3354_;
  assign new_A3402_ = new_A3370_ | new_A3407_;
  assign new_A3403_ = ~new_A3370_ & ~new_A3406_;
  assign new_A3404_ = new_A3353_ | new_A3370_;
  assign new_A3405_ = new_A3353_ | new_A3354_;
  assign new_A3406_ = new_A3370_ & new_A3407_;
  assign new_A3407_ = ~new_A3352_ | ~new_A3377_;
  assign new_A3408_ = new_A3385_ & new_A3405_;
  assign new_A3409_ = ~new_A3385_ & ~new_A3405_;
  assign new_A3410_ = new_A3414_ | new_A3415_;
  assign new_A3411_ = ~new_A3356_ & new_A3370_;
  assign new_A3412_ = new_A3416_ | new_A3417_;
  assign new_A3413_ = new_A3356_ & new_A3370_;
  assign new_A3414_ = ~new_A3356_ & ~new_A3370_;
  assign new_A3415_ = new_A3356_ & ~new_A3370_;
  assign new_A3416_ = new_A3356_ & ~new_A3370_;
  assign new_A3417_ = ~new_A3356_ & new_A3370_;
  assign new_A3418_ = new_A6841_;
  assign new_A3419_ = new_A6908_;
  assign new_A3420_ = new_A6975_;
  assign new_A3421_ = new_A7042_;
  assign new_A3422_ = new_A7109_;
  assign new_A3423_ = new_A7176_;
  assign new_A3424_ = new_A3431_ & new_A3430_;
  assign new_A3425_ = new_A3433_ | new_A3432_;
  assign new_A3426_ = new_A3435_ | new_A3434_;
  assign new_A3427_ = new_A3437_ & new_A3436_;
  assign new_A3428_ = new_A3437_ & new_A3438_;
  assign new_A3429_ = new_A3430_ | new_A3439_;
  assign new_A3430_ = new_A3419_ | new_A3442_;
  assign new_A3431_ = new_A3441_ | new_A3440_;
  assign new_A3432_ = new_A3446_ & new_A3445_;
  assign new_A3433_ = new_A3444_ & new_A3443_;
  assign new_A3434_ = new_A3449_ | new_A3448_;
  assign new_A3435_ = new_A3444_ & new_A3447_;
  assign new_A3436_ = new_A3419_ | new_A3452_;
  assign new_A3437_ = new_A3451_ | new_A3450_;
  assign new_A3438_ = new_A3454_ | new_A3453_;
  assign new_A3439_ = ~new_A3430_ & new_A3456_;
  assign new_A3440_ = ~new_A3432_ & new_A3444_;
  assign new_A3441_ = new_A3432_ & ~new_A3444_;
  assign new_A3442_ = new_A3418_ & ~new_A3419_;
  assign new_A3443_ = ~new_A3465_ | ~new_A3466_;
  assign new_A3444_ = new_A3458_ | new_A3460_;
  assign new_A3445_ = new_A3468_ | new_A3467_;
  assign new_A3446_ = new_A3462_ | new_A3461_;
  assign new_A3447_ = ~new_A3470_ | ~new_A3469_;
  assign new_A3448_ = ~new_A3471_ & new_A3472_;
  assign new_A3449_ = new_A3471_ & ~new_A3472_;
  assign new_A3450_ = ~new_A3418_ & new_A3419_;
  assign new_A3451_ = new_A3418_ & ~new_A3419_;
  assign new_A3452_ = ~new_A3434_ | new_A3444_;
  assign new_A3453_ = new_A3434_ & new_A3444_;
  assign new_A3454_ = ~new_A3434_ & ~new_A3444_;
  assign new_A3455_ = new_A3476_ | new_A3475_;
  assign new_A3456_ = new_A3422_ | new_A3455_;
  assign new_A3457_ = new_A3480_ | new_A3479_;
  assign new_A3458_ = ~new_A3422_ & new_A3457_;
  assign new_A3459_ = new_A3478_ | new_A3477_;
  assign new_A3460_ = new_A3422_ & new_A3459_;
  assign new_A3461_ = new_A3420_ & ~new_A3430_;
  assign new_A3462_ = ~new_A3420_ & new_A3430_;
  assign new_A3463_ = ~new_A3419_ | ~new_A3444_;
  assign new_A3464_ = new_A3430_ & new_A3463_;
  assign new_A3465_ = ~new_A3430_ & ~new_A3464_;
  assign new_A3466_ = new_A3430_ | new_A3463_;
  assign new_A3467_ = ~new_A3420_ & new_A3421_;
  assign new_A3468_ = new_A3420_ & ~new_A3421_;
  assign new_A3469_ = new_A3437_ | new_A3474_;
  assign new_A3470_ = ~new_A3437_ & ~new_A3473_;
  assign new_A3471_ = new_A3420_ | new_A3437_;
  assign new_A3472_ = new_A3420_ | new_A3421_;
  assign new_A3473_ = new_A3437_ & new_A3474_;
  assign new_A3474_ = ~new_A3419_ | ~new_A3444_;
  assign new_A3475_ = new_A3452_ & new_A3472_;
  assign new_A3476_ = ~new_A3452_ & ~new_A3472_;
  assign new_A3477_ = new_A3481_ | new_A3482_;
  assign new_A3478_ = ~new_A3423_ & new_A3437_;
  assign new_A3479_ = new_A3483_ | new_A3484_;
  assign new_A3480_ = new_A3423_ & new_A3437_;
  assign new_A3481_ = ~new_A3423_ & ~new_A3437_;
  assign new_A3482_ = new_A3423_ & ~new_A3437_;
  assign new_A3483_ = new_A3423_ & ~new_A3437_;
  assign new_A3484_ = ~new_A3423_ & new_A3437_;
  assign new_A3485_ = new_A7243_;
  assign new_A3486_ = new_A7310_;
  assign new_A3487_ = new_A7377_;
  assign new_A3488_ = new_A7444_;
  assign new_A3489_ = new_A7511_;
  assign new_A3490_ = new_A7578_;
  assign new_A3491_ = new_A3498_ & new_A3497_;
  assign new_A3492_ = new_A3500_ | new_A3499_;
  assign new_A3493_ = new_A3502_ | new_A3501_;
  assign new_A3494_ = new_A3504_ & new_A3503_;
  assign new_A3495_ = new_A3504_ & new_A3505_;
  assign new_A3496_ = new_A3497_ | new_A3506_;
  assign new_A3497_ = new_A3486_ | new_A3509_;
  assign new_A3498_ = new_A3508_ | new_A3507_;
  assign new_A3499_ = new_A3513_ & new_A3512_;
  assign new_A3500_ = new_A3511_ & new_A3510_;
  assign new_A3501_ = new_A3516_ | new_A3515_;
  assign new_A3502_ = new_A3511_ & new_A3514_;
  assign new_A3503_ = new_A3486_ | new_A3519_;
  assign new_A3504_ = new_A3518_ | new_A3517_;
  assign new_A3505_ = new_A3521_ | new_A3520_;
  assign new_A3506_ = ~new_A3497_ & new_A3523_;
  assign new_A3507_ = ~new_A3499_ & new_A3511_;
  assign new_A3508_ = new_A3499_ & ~new_A3511_;
  assign new_A3509_ = new_A3485_ & ~new_A3486_;
  assign new_A3510_ = ~new_A3532_ | ~new_A3533_;
  assign new_A3511_ = new_A3525_ | new_A3527_;
  assign new_A3512_ = new_A3535_ | new_A3534_;
  assign new_A3513_ = new_A3529_ | new_A3528_;
  assign new_A3514_ = ~new_A3537_ | ~new_A3536_;
  assign new_A3515_ = ~new_A3538_ & new_A3539_;
  assign new_A3516_ = new_A3538_ & ~new_A3539_;
  assign new_A3517_ = ~new_A3485_ & new_A3486_;
  assign new_A3518_ = new_A3485_ & ~new_A3486_;
  assign new_A3519_ = ~new_A3501_ | new_A3511_;
  assign new_A3520_ = new_A3501_ & new_A3511_;
  assign new_A3521_ = ~new_A3501_ & ~new_A3511_;
  assign new_A3522_ = new_A3543_ | new_A3542_;
  assign new_A3523_ = new_A3489_ | new_A3522_;
  assign new_A3524_ = new_A3547_ | new_A3546_;
  assign new_A3525_ = ~new_A3489_ & new_A3524_;
  assign new_A3526_ = new_A3545_ | new_A3544_;
  assign new_A3527_ = new_A3489_ & new_A3526_;
  assign new_A3528_ = new_A3487_ & ~new_A3497_;
  assign new_A3529_ = ~new_A3487_ & new_A3497_;
  assign new_A3530_ = ~new_A3486_ | ~new_A3511_;
  assign new_A3531_ = new_A3497_ & new_A3530_;
  assign new_A3532_ = ~new_A3497_ & ~new_A3531_;
  assign new_A3533_ = new_A3497_ | new_A3530_;
  assign new_A3534_ = ~new_A3487_ & new_A3488_;
  assign new_A3535_ = new_A3487_ & ~new_A3488_;
  assign new_A3536_ = new_A3504_ | new_A3541_;
  assign new_A3537_ = ~new_A3504_ & ~new_A3540_;
  assign new_A3538_ = new_A3487_ | new_A3504_;
  assign new_A3539_ = new_A3487_ | new_A3488_;
  assign new_A3540_ = new_A3504_ & new_A3541_;
  assign new_A3541_ = ~new_A3486_ | ~new_A3511_;
  assign new_A3542_ = new_A3519_ & new_A3539_;
  assign new_A3543_ = ~new_A3519_ & ~new_A3539_;
  assign new_A3544_ = new_A3548_ | new_A3549_;
  assign new_A3545_ = ~new_A3490_ & new_A3504_;
  assign new_A3546_ = new_A3550_ | new_A3551_;
  assign new_A3547_ = new_A3490_ & new_A3504_;
  assign new_A3548_ = ~new_A3490_ & ~new_A3504_;
  assign new_A3549_ = new_A3490_ & ~new_A3504_;
  assign new_A3550_ = new_A3490_ & ~new_A3504_;
  assign new_A3551_ = ~new_A3490_ & new_A3504_;
  assign new_A3552_ = new_A7645_;
  assign new_A3553_ = new_A7712_;
  assign new_A3554_ = new_A7779_;
  assign new_A3555_ = new_A7846_;
  assign new_A3556_ = new_A7913_;
  assign new_A3557_ = new_A7980_;
  assign new_A3558_ = new_A3565_ & new_A3564_;
  assign new_A3559_ = new_A3567_ | new_A3566_;
  assign new_A3560_ = new_A3569_ | new_A3568_;
  assign new_A3561_ = new_A3571_ & new_A3570_;
  assign new_A3562_ = new_A3571_ & new_A3572_;
  assign new_A3563_ = new_A3564_ | new_A3573_;
  assign new_A3564_ = new_A3553_ | new_A3576_;
  assign new_A3565_ = new_A3575_ | new_A3574_;
  assign new_A3566_ = new_A3580_ & new_A3579_;
  assign new_A3567_ = new_A3578_ & new_A3577_;
  assign new_A3568_ = new_A3583_ | new_A3582_;
  assign new_A3569_ = new_A3578_ & new_A3581_;
  assign new_A3570_ = new_A3553_ | new_A3586_;
  assign new_A3571_ = new_A3585_ | new_A3584_;
  assign new_A3572_ = new_A3588_ | new_A3587_;
  assign new_A3573_ = ~new_A3564_ & new_A3590_;
  assign new_A3574_ = ~new_A3566_ & new_A3578_;
  assign new_A3575_ = new_A3566_ & ~new_A3578_;
  assign new_A3576_ = new_A3552_ & ~new_A3553_;
  assign new_A3577_ = ~new_A3599_ | ~new_A3600_;
  assign new_A3578_ = new_A3592_ | new_A3594_;
  assign new_A3579_ = new_A3602_ | new_A3601_;
  assign new_A3580_ = new_A3596_ | new_A3595_;
  assign new_A3581_ = ~new_A3604_ | ~new_A3603_;
  assign new_A3582_ = ~new_A3605_ & new_A3606_;
  assign new_A3583_ = new_A3605_ & ~new_A3606_;
  assign new_A3584_ = ~new_A3552_ & new_A3553_;
  assign new_A3585_ = new_A3552_ & ~new_A3553_;
  assign new_A3586_ = ~new_A3568_ | new_A3578_;
  assign new_A3587_ = new_A3568_ & new_A3578_;
  assign new_A3588_ = ~new_A3568_ & ~new_A3578_;
  assign new_A3589_ = new_A3610_ | new_A3609_;
  assign new_A3590_ = new_A3556_ | new_A3589_;
  assign new_A3591_ = new_A3614_ | new_A3613_;
  assign new_A3592_ = ~new_A3556_ & new_A3591_;
  assign new_A3593_ = new_A3612_ | new_A3611_;
  assign new_A3594_ = new_A3556_ & new_A3593_;
  assign new_A3595_ = new_A3554_ & ~new_A3564_;
  assign new_A3596_ = ~new_A3554_ & new_A3564_;
  assign new_A3597_ = ~new_A3553_ | ~new_A3578_;
  assign new_A3598_ = new_A3564_ & new_A3597_;
  assign new_A3599_ = ~new_A3564_ & ~new_A3598_;
  assign new_A3600_ = new_A3564_ | new_A3597_;
  assign new_A3601_ = ~new_A3554_ & new_A3555_;
  assign new_A3602_ = new_A3554_ & ~new_A3555_;
  assign new_A3603_ = new_A3571_ | new_A3608_;
  assign new_A3604_ = ~new_A3571_ & ~new_A3607_;
  assign new_A3605_ = new_A3554_ | new_A3571_;
  assign new_A3606_ = new_A3554_ | new_A3555_;
  assign new_A3607_ = new_A3571_ & new_A3608_;
  assign new_A3608_ = ~new_A3553_ | ~new_A3578_;
  assign new_A3609_ = new_A3586_ & new_A3606_;
  assign new_A3610_ = ~new_A3586_ & ~new_A3606_;
  assign new_A3611_ = new_A3615_ | new_A3616_;
  assign new_A3612_ = ~new_A3557_ & new_A3571_;
  assign new_A3613_ = new_A3617_ | new_A3618_;
  assign new_A3614_ = new_A3557_ & new_A3571_;
  assign new_A3615_ = ~new_A3557_ & ~new_A3571_;
  assign new_A3616_ = new_A3557_ & ~new_A3571_;
  assign new_A3617_ = new_A3557_ & ~new_A3571_;
  assign new_A3618_ = ~new_A3557_ & new_A3571_;
  assign new_A3619_ = new_A5639_;
  assign new_A3620_ = new_A5703_;
  assign new_A3621_ = new_A5770_;
  assign new_A3622_ = new_A5837_;
  assign new_A3623_ = new_A5904_;
  assign new_A3624_ = new_A5971_;
  assign new_A3625_ = new_A3632_ & new_A3631_;
  assign new_A3626_ = new_A3634_ | new_A3633_;
  assign new_A3627_ = new_A3636_ | new_A3635_;
  assign new_A3628_ = new_A3638_ & new_A3637_;
  assign new_A3629_ = new_A3638_ & new_A3639_;
  assign new_A3630_ = new_A3631_ | new_A3640_;
  assign new_A3631_ = new_A3620_ | new_A3643_;
  assign new_A3632_ = new_A3642_ | new_A3641_;
  assign new_A3633_ = new_A3647_ & new_A3646_;
  assign new_A3634_ = new_A3645_ & new_A3644_;
  assign new_A3635_ = new_A3650_ | new_A3649_;
  assign new_A3636_ = new_A3645_ & new_A3648_;
  assign new_A3637_ = new_A3620_ | new_A3653_;
  assign new_A3638_ = new_A3652_ | new_A3651_;
  assign new_A3639_ = new_A3655_ | new_A3654_;
  assign new_A3640_ = ~new_A3631_ & new_A3657_;
  assign new_A3641_ = ~new_A3633_ & new_A3645_;
  assign new_A3642_ = new_A3633_ & ~new_A3645_;
  assign new_A3643_ = new_A3619_ & ~new_A3620_;
  assign new_A3644_ = ~new_A3666_ | ~new_A3667_;
  assign new_A3645_ = new_A3659_ | new_A3661_;
  assign new_A3646_ = new_A3669_ | new_A3668_;
  assign new_A3647_ = new_A3663_ | new_A3662_;
  assign new_A3648_ = ~new_A3671_ | ~new_A3670_;
  assign new_A3649_ = ~new_A3672_ & new_A3673_;
  assign new_A3650_ = new_A3672_ & ~new_A3673_;
  assign new_A3651_ = ~new_A3619_ & new_A3620_;
  assign new_A3652_ = new_A3619_ & ~new_A3620_;
  assign new_A3653_ = ~new_A3635_ | new_A3645_;
  assign new_A3654_ = new_A3635_ & new_A3645_;
  assign new_A3655_ = ~new_A3635_ & ~new_A3645_;
  assign new_A3656_ = new_A3677_ | new_A3676_;
  assign new_A3657_ = new_A3623_ | new_A3656_;
  assign new_A3658_ = new_A3681_ | new_A3680_;
  assign new_A3659_ = ~new_A3623_ & new_A3658_;
  assign new_A3660_ = new_A3679_ | new_A3678_;
  assign new_A3661_ = new_A3623_ & new_A3660_;
  assign new_A3662_ = new_A3621_ & ~new_A3631_;
  assign new_A3663_ = ~new_A3621_ & new_A3631_;
  assign new_A3664_ = ~new_A3620_ | ~new_A3645_;
  assign new_A3665_ = new_A3631_ & new_A3664_;
  assign new_A3666_ = ~new_A3631_ & ~new_A3665_;
  assign new_A3667_ = new_A3631_ | new_A3664_;
  assign new_A3668_ = ~new_A3621_ & new_A3622_;
  assign new_A3669_ = new_A3621_ & ~new_A3622_;
  assign new_A3670_ = new_A3638_ | new_A3675_;
  assign new_A3671_ = ~new_A3638_ & ~new_A3674_;
  assign new_A3672_ = new_A3621_ | new_A3638_;
  assign new_A3673_ = new_A3621_ | new_A3622_;
  assign new_A3674_ = new_A3638_ & new_A3675_;
  assign new_A3675_ = ~new_A3620_ | ~new_A3645_;
  assign new_A3676_ = new_A3653_ & new_A3673_;
  assign new_A3677_ = ~new_A3653_ & ~new_A3673_;
  assign new_A3678_ = new_A3682_ | new_A3683_;
  assign new_A3679_ = ~new_A3624_ & new_A3638_;
  assign new_A3680_ = new_A3684_ | new_A3685_;
  assign new_A3681_ = new_A3624_ & new_A3638_;
  assign new_A3682_ = ~new_A3624_ & ~new_A3638_;
  assign new_A3683_ = new_A3624_ & ~new_A3638_;
  assign new_A3684_ = new_A3624_ & ~new_A3638_;
  assign new_A3685_ = ~new_A3624_ & new_A3638_;
  assign new_A3686_ = new_A6038_;
  assign new_A3687_ = new_A6105_;
  assign new_A3688_ = new_A6172_;
  assign new_A3689_ = new_A6239_;
  assign new_A3690_ = new_A6306_;
  assign new_A3691_ = new_A6373_;
  assign new_A3692_ = new_A3699_ & new_A3698_;
  assign new_A3693_ = new_A3701_ | new_A3700_;
  assign new_A3694_ = new_A3703_ | new_A3702_;
  assign new_A3695_ = new_A3705_ & new_A3704_;
  assign new_A3696_ = new_A3705_ & new_A3706_;
  assign new_A3697_ = new_A3698_ | new_A3707_;
  assign new_A3698_ = new_A3687_ | new_A3710_;
  assign new_A3699_ = new_A3709_ | new_A3708_;
  assign new_A3700_ = new_A3714_ & new_A3713_;
  assign new_A3701_ = new_A3712_ & new_A3711_;
  assign new_A3702_ = new_A3717_ | new_A3716_;
  assign new_A3703_ = new_A3712_ & new_A3715_;
  assign new_A3704_ = new_A3687_ | new_A3720_;
  assign new_A3705_ = new_A3719_ | new_A3718_;
  assign new_A3706_ = new_A3722_ | new_A3721_;
  assign new_A3707_ = ~new_A3698_ & new_A3724_;
  assign new_A3708_ = ~new_A3700_ & new_A3712_;
  assign new_A3709_ = new_A3700_ & ~new_A3712_;
  assign new_A3710_ = new_A3686_ & ~new_A3687_;
  assign new_A3711_ = ~new_A3733_ | ~new_A3734_;
  assign new_A3712_ = new_A3726_ | new_A3728_;
  assign new_A3713_ = new_A3736_ | new_A3735_;
  assign new_A3714_ = new_A3730_ | new_A3729_;
  assign new_A3715_ = ~new_A3738_ | ~new_A3737_;
  assign new_A3716_ = ~new_A3739_ & new_A3740_;
  assign new_A3717_ = new_A3739_ & ~new_A3740_;
  assign new_A3718_ = ~new_A3686_ & new_A3687_;
  assign new_A3719_ = new_A3686_ & ~new_A3687_;
  assign new_A3720_ = ~new_A3702_ | new_A3712_;
  assign new_A3721_ = new_A3702_ & new_A3712_;
  assign new_A3722_ = ~new_A3702_ & ~new_A3712_;
  assign new_A3723_ = new_A3744_ | new_A3743_;
  assign new_A3724_ = new_A3690_ | new_A3723_;
  assign new_A3725_ = new_A3748_ | new_A3747_;
  assign new_A3726_ = ~new_A3690_ & new_A3725_;
  assign new_A3727_ = new_A3746_ | new_A3745_;
  assign new_A3728_ = new_A3690_ & new_A3727_;
  assign new_A3729_ = new_A3688_ & ~new_A3698_;
  assign new_A3730_ = ~new_A3688_ & new_A3698_;
  assign new_A3731_ = ~new_A3687_ | ~new_A3712_;
  assign new_A3732_ = new_A3698_ & new_A3731_;
  assign new_A3733_ = ~new_A3698_ & ~new_A3732_;
  assign new_A3734_ = new_A3698_ | new_A3731_;
  assign new_A3735_ = ~new_A3688_ & new_A3689_;
  assign new_A3736_ = new_A3688_ & ~new_A3689_;
  assign new_A3737_ = new_A3705_ | new_A3742_;
  assign new_A3738_ = ~new_A3705_ & ~new_A3741_;
  assign new_A3739_ = new_A3688_ | new_A3705_;
  assign new_A3740_ = new_A3688_ | new_A3689_;
  assign new_A3741_ = new_A3705_ & new_A3742_;
  assign new_A3742_ = ~new_A3687_ | ~new_A3712_;
  assign new_A3743_ = new_A3720_ & new_A3740_;
  assign new_A3744_ = ~new_A3720_ & ~new_A3740_;
  assign new_A3745_ = new_A3749_ | new_A3750_;
  assign new_A3746_ = ~new_A3691_ & new_A3705_;
  assign new_A3747_ = new_A3751_ | new_A3752_;
  assign new_A3748_ = new_A3691_ & new_A3705_;
  assign new_A3749_ = ~new_A3691_ & ~new_A3705_;
  assign new_A3750_ = new_A3691_ & ~new_A3705_;
  assign new_A3751_ = new_A3691_ & ~new_A3705_;
  assign new_A3752_ = ~new_A3691_ & new_A3705_;
  assign new_A3753_ = new_A6440_;
  assign new_A3754_ = new_A6507_;
  assign new_A3755_ = new_A6574_;
  assign new_A3756_ = new_A6641_;
  assign new_A3757_ = new_A6708_;
  assign new_A3758_ = new_A6775_;
  assign new_A3759_ = new_A3766_ & new_A3765_;
  assign new_A3760_ = new_A3768_ | new_A3767_;
  assign new_A3761_ = new_A3770_ | new_A3769_;
  assign new_A3762_ = new_A3772_ & new_A3771_;
  assign new_A3763_ = new_A3772_ & new_A3773_;
  assign new_A3764_ = new_A3765_ | new_A3774_;
  assign new_A3765_ = new_A3754_ | new_A3777_;
  assign new_A3766_ = new_A3776_ | new_A3775_;
  assign new_A3767_ = new_A3781_ & new_A3780_;
  assign new_A3768_ = new_A3779_ & new_A3778_;
  assign new_A3769_ = new_A3784_ | new_A3783_;
  assign new_A3770_ = new_A3779_ & new_A3782_;
  assign new_A3771_ = new_A3754_ | new_A3787_;
  assign new_A3772_ = new_A3786_ | new_A3785_;
  assign new_A3773_ = new_A3789_ | new_A3788_;
  assign new_A3774_ = ~new_A3765_ & new_A3791_;
  assign new_A3775_ = ~new_A3767_ & new_A3779_;
  assign new_A3776_ = new_A3767_ & ~new_A3779_;
  assign new_A3777_ = new_A3753_ & ~new_A3754_;
  assign new_A3778_ = ~new_A3800_ | ~new_A3801_;
  assign new_A3779_ = new_A3793_ | new_A3795_;
  assign new_A3780_ = new_A3803_ | new_A3802_;
  assign new_A3781_ = new_A3797_ | new_A3796_;
  assign new_A3782_ = ~new_A3805_ | ~new_A3804_;
  assign new_A3783_ = ~new_A3806_ & new_A3807_;
  assign new_A3784_ = new_A3806_ & ~new_A3807_;
  assign new_A3785_ = ~new_A3753_ & new_A3754_;
  assign new_A3786_ = new_A3753_ & ~new_A3754_;
  assign new_A3787_ = ~new_A3769_ | new_A3779_;
  assign new_A3788_ = new_A3769_ & new_A3779_;
  assign new_A3789_ = ~new_A3769_ & ~new_A3779_;
  assign new_A3790_ = new_A3811_ | new_A3810_;
  assign new_A3791_ = new_A3757_ | new_A3790_;
  assign new_A3792_ = new_A3815_ | new_A3814_;
  assign new_A3793_ = ~new_A3757_ & new_A3792_;
  assign new_A3794_ = new_A3813_ | new_A3812_;
  assign new_A3795_ = new_A3757_ & new_A3794_;
  assign new_A3796_ = new_A3755_ & ~new_A3765_;
  assign new_A3797_ = ~new_A3755_ & new_A3765_;
  assign new_A3798_ = ~new_A3754_ | ~new_A3779_;
  assign new_A3799_ = new_A3765_ & new_A3798_;
  assign new_A3800_ = ~new_A3765_ & ~new_A3799_;
  assign new_A3801_ = new_A3765_ | new_A3798_;
  assign new_A3802_ = ~new_A3755_ & new_A3756_;
  assign new_A3803_ = new_A3755_ & ~new_A3756_;
  assign new_A3804_ = new_A3772_ | new_A3809_;
  assign new_A3805_ = ~new_A3772_ & ~new_A3808_;
  assign new_A3806_ = new_A3755_ | new_A3772_;
  assign new_A3807_ = new_A3755_ | new_A3756_;
  assign new_A3808_ = new_A3772_ & new_A3809_;
  assign new_A3809_ = ~new_A3754_ | ~new_A3779_;
  assign new_A3810_ = new_A3787_ & new_A3807_;
  assign new_A3811_ = ~new_A3787_ & ~new_A3807_;
  assign new_A3812_ = new_A3816_ | new_A3817_;
  assign new_A3813_ = ~new_A3758_ & new_A3772_;
  assign new_A3814_ = new_A3818_ | new_A3819_;
  assign new_A3815_ = new_A3758_ & new_A3772_;
  assign new_A3816_ = ~new_A3758_ & ~new_A3772_;
  assign new_A3817_ = new_A3758_ & ~new_A3772_;
  assign new_A3818_ = new_A3758_ & ~new_A3772_;
  assign new_A3819_ = ~new_A3758_ & new_A3772_;
  assign new_A3820_ = new_A6842_;
  assign new_A3821_ = new_A6909_;
  assign new_A3822_ = new_A6976_;
  assign new_A3823_ = new_A7043_;
  assign new_A3824_ = new_A7110_;
  assign new_A3825_ = new_A7177_;
  assign new_A3826_ = new_A3833_ & new_A3832_;
  assign new_A3827_ = new_A3835_ | new_A3834_;
  assign new_A3828_ = new_A3837_ | new_A3836_;
  assign new_A3829_ = new_A3839_ & new_A3838_;
  assign new_A3830_ = new_A3839_ & new_A3840_;
  assign new_A3831_ = new_A3832_ | new_A3841_;
  assign new_A3832_ = new_A3821_ | new_A3844_;
  assign new_A3833_ = new_A3843_ | new_A3842_;
  assign new_A3834_ = new_A3848_ & new_A3847_;
  assign new_A3835_ = new_A3846_ & new_A3845_;
  assign new_A3836_ = new_A3851_ | new_A3850_;
  assign new_A3837_ = new_A3846_ & new_A3849_;
  assign new_A3838_ = new_A3821_ | new_A3854_;
  assign new_A3839_ = new_A3853_ | new_A3852_;
  assign new_A3840_ = new_A3856_ | new_A3855_;
  assign new_A3841_ = ~new_A3832_ & new_A3858_;
  assign new_A3842_ = ~new_A3834_ & new_A3846_;
  assign new_A3843_ = new_A3834_ & ~new_A3846_;
  assign new_A3844_ = new_A3820_ & ~new_A3821_;
  assign new_A3845_ = ~new_A3867_ | ~new_A3868_;
  assign new_A3846_ = new_A3860_ | new_A3862_;
  assign new_A3847_ = new_A3870_ | new_A3869_;
  assign new_A3848_ = new_A3864_ | new_A3863_;
  assign new_A3849_ = ~new_A3872_ | ~new_A3871_;
  assign new_A3850_ = ~new_A3873_ & new_A3874_;
  assign new_A3851_ = new_A3873_ & ~new_A3874_;
  assign new_A3852_ = ~new_A3820_ & new_A3821_;
  assign new_A3853_ = new_A3820_ & ~new_A3821_;
  assign new_A3854_ = ~new_A3836_ | new_A3846_;
  assign new_A3855_ = new_A3836_ & new_A3846_;
  assign new_A3856_ = ~new_A3836_ & ~new_A3846_;
  assign new_A3857_ = new_A3878_ | new_A3877_;
  assign new_A3858_ = new_A3824_ | new_A3857_;
  assign new_A3859_ = new_A3882_ | new_A3881_;
  assign new_A3860_ = ~new_A3824_ & new_A3859_;
  assign new_A3861_ = new_A3880_ | new_A3879_;
  assign new_A3862_ = new_A3824_ & new_A3861_;
  assign new_A3863_ = new_A3822_ & ~new_A3832_;
  assign new_A3864_ = ~new_A3822_ & new_A3832_;
  assign new_A3865_ = ~new_A3821_ | ~new_A3846_;
  assign new_A3866_ = new_A3832_ & new_A3865_;
  assign new_A3867_ = ~new_A3832_ & ~new_A3866_;
  assign new_A3868_ = new_A3832_ | new_A3865_;
  assign new_A3869_ = ~new_A3822_ & new_A3823_;
  assign new_A3870_ = new_A3822_ & ~new_A3823_;
  assign new_A3871_ = new_A3839_ | new_A3876_;
  assign new_A3872_ = ~new_A3839_ & ~new_A3875_;
  assign new_A3873_ = new_A3822_ | new_A3839_;
  assign new_A3874_ = new_A3822_ | new_A3823_;
  assign new_A3875_ = new_A3839_ & new_A3876_;
  assign new_A3876_ = ~new_A3821_ | ~new_A3846_;
  assign new_A3877_ = new_A3854_ & new_A3874_;
  assign new_A3878_ = ~new_A3854_ & ~new_A3874_;
  assign new_A3879_ = new_A3883_ | new_A3884_;
  assign new_A3880_ = ~new_A3825_ & new_A3839_;
  assign new_A3881_ = new_A3885_ | new_A3886_;
  assign new_A3882_ = new_A3825_ & new_A3839_;
  assign new_A3883_ = ~new_A3825_ & ~new_A3839_;
  assign new_A3884_ = new_A3825_ & ~new_A3839_;
  assign new_A3885_ = new_A3825_ & ~new_A3839_;
  assign new_A3886_ = ~new_A3825_ & new_A3839_;
  assign new_A3887_ = new_A7244_;
  assign new_A3888_ = new_A7311_;
  assign new_A3889_ = new_A7378_;
  assign new_A3890_ = new_A7445_;
  assign new_A3891_ = new_A7512_;
  assign new_A3892_ = new_A7579_;
  assign new_A3893_ = new_A3900_ & new_A3899_;
  assign new_A3894_ = new_A3902_ | new_A3901_;
  assign new_A3895_ = new_A3904_ | new_A3903_;
  assign new_A3896_ = new_A3906_ & new_A3905_;
  assign new_A3897_ = new_A3906_ & new_A3907_;
  assign new_A3898_ = new_A3899_ | new_A3908_;
  assign new_A3899_ = new_A3888_ | new_A3911_;
  assign new_A3900_ = new_A3910_ | new_A3909_;
  assign new_A3901_ = new_A3915_ & new_A3914_;
  assign new_A3902_ = new_A3913_ & new_A3912_;
  assign new_A3903_ = new_A3918_ | new_A3917_;
  assign new_A3904_ = new_A3913_ & new_A3916_;
  assign new_A3905_ = new_A3888_ | new_A3921_;
  assign new_A3906_ = new_A3920_ | new_A3919_;
  assign new_A3907_ = new_A3923_ | new_A3922_;
  assign new_A3908_ = ~new_A3899_ & new_A3925_;
  assign new_A3909_ = ~new_A3901_ & new_A3913_;
  assign new_A3910_ = new_A3901_ & ~new_A3913_;
  assign new_A3911_ = new_A3887_ & ~new_A3888_;
  assign new_A3912_ = ~new_A3934_ | ~new_A3935_;
  assign new_A3913_ = new_A3927_ | new_A3929_;
  assign new_A3914_ = new_A3937_ | new_A3936_;
  assign new_A3915_ = new_A3931_ | new_A3930_;
  assign new_A3916_ = ~new_A3939_ | ~new_A3938_;
  assign new_A3917_ = ~new_A3940_ & new_A3941_;
  assign new_A3918_ = new_A3940_ & ~new_A3941_;
  assign new_A3919_ = ~new_A3887_ & new_A3888_;
  assign new_A3920_ = new_A3887_ & ~new_A3888_;
  assign new_A3921_ = ~new_A3903_ | new_A3913_;
  assign new_A3922_ = new_A3903_ & new_A3913_;
  assign new_A3923_ = ~new_A3903_ & ~new_A3913_;
  assign new_A3924_ = new_A3945_ | new_A3944_;
  assign new_A3925_ = new_A3891_ | new_A3924_;
  assign new_A3926_ = new_A3949_ | new_A3948_;
  assign new_A3927_ = ~new_A3891_ & new_A3926_;
  assign new_A3928_ = new_A3947_ | new_A3946_;
  assign new_A3929_ = new_A3891_ & new_A3928_;
  assign new_A3930_ = new_A3889_ & ~new_A3899_;
  assign new_A3931_ = ~new_A3889_ & new_A3899_;
  assign new_A3932_ = ~new_A3888_ | ~new_A3913_;
  assign new_A3933_ = new_A3899_ & new_A3932_;
  assign new_A3934_ = ~new_A3899_ & ~new_A3933_;
  assign new_A3935_ = new_A3899_ | new_A3932_;
  assign new_A3936_ = ~new_A3889_ & new_A3890_;
  assign new_A3937_ = new_A3889_ & ~new_A3890_;
  assign new_A3938_ = new_A3906_ | new_A3943_;
  assign new_A3939_ = ~new_A3906_ & ~new_A3942_;
  assign new_A3940_ = new_A3889_ | new_A3906_;
  assign new_A3941_ = new_A3889_ | new_A3890_;
  assign new_A3942_ = new_A3906_ & new_A3943_;
  assign new_A3943_ = ~new_A3888_ | ~new_A3913_;
  assign new_A3944_ = new_A3921_ & new_A3941_;
  assign new_A3945_ = ~new_A3921_ & ~new_A3941_;
  assign new_A3946_ = new_A3950_ | new_A3951_;
  assign new_A3947_ = ~new_A3892_ & new_A3906_;
  assign new_A3948_ = new_A3952_ | new_A3953_;
  assign new_A3949_ = new_A3892_ & new_A3906_;
  assign new_A3950_ = ~new_A3892_ & ~new_A3906_;
  assign new_A3951_ = new_A3892_ & ~new_A3906_;
  assign new_A3952_ = new_A3892_ & ~new_A3906_;
  assign new_A3953_ = ~new_A3892_ & new_A3906_;
  assign new_A3954_ = new_A7646_;
  assign new_A3955_ = new_A7713_;
  assign new_A3956_ = new_A7780_;
  assign new_A3957_ = new_A7847_;
  assign new_A3958_ = new_A7914_;
  assign new_A3959_ = new_A7981_;
  assign new_A3960_ = new_A3967_ & new_A3966_;
  assign new_A3961_ = new_A3969_ | new_A3968_;
  assign new_A3962_ = new_A3971_ | new_A3970_;
  assign new_A3963_ = new_A3973_ & new_A3972_;
  assign new_A3964_ = new_A3973_ & new_A3974_;
  assign new_A3965_ = new_A3966_ | new_A3975_;
  assign new_A3966_ = new_A3955_ | new_A3978_;
  assign new_A3967_ = new_A3977_ | new_A3976_;
  assign new_A3968_ = new_A3982_ & new_A3981_;
  assign new_A3969_ = new_A3980_ & new_A3979_;
  assign new_A3970_ = new_A3985_ | new_A3984_;
  assign new_A3971_ = new_A3980_ & new_A3983_;
  assign new_A3972_ = new_A3955_ | new_A3988_;
  assign new_A3973_ = new_A3987_ | new_A3986_;
  assign new_A3974_ = new_A3990_ | new_A3989_;
  assign new_A3975_ = ~new_A3966_ & new_A3992_;
  assign new_A3976_ = ~new_A3968_ & new_A3980_;
  assign new_A3977_ = new_A3968_ & ~new_A3980_;
  assign new_A3978_ = new_A3954_ & ~new_A3955_;
  assign new_A3979_ = ~new_A4001_ | ~new_A4002_;
  assign new_A3980_ = new_A3994_ | new_A3996_;
  assign new_A3981_ = new_A4004_ | new_A4003_;
  assign new_A3982_ = new_A3998_ | new_A3997_;
  assign new_A3983_ = ~new_A4006_ | ~new_A4005_;
  assign new_A3984_ = ~new_A4007_ & new_A4008_;
  assign new_A3985_ = new_A4007_ & ~new_A4008_;
  assign new_A3986_ = ~new_A3954_ & new_A3955_;
  assign new_A3987_ = new_A3954_ & ~new_A3955_;
  assign new_A3988_ = ~new_A3970_ | new_A3980_;
  assign new_A3989_ = new_A3970_ & new_A3980_;
  assign new_A3990_ = ~new_A3970_ & ~new_A3980_;
  assign new_A3991_ = new_A4012_ | new_A4011_;
  assign new_A3992_ = new_A3958_ | new_A3991_;
  assign new_A3993_ = new_A4016_ | new_A4015_;
  assign new_A3994_ = ~new_A3958_ & new_A3993_;
  assign new_A3995_ = new_A4014_ | new_A4013_;
  assign new_A3996_ = new_A3958_ & new_A3995_;
  assign new_A3997_ = new_A3956_ & ~new_A3966_;
  assign new_A3998_ = ~new_A3956_ & new_A3966_;
  assign new_A3999_ = ~new_A3955_ | ~new_A3980_;
  assign new_A4000_ = new_A3966_ & new_A3999_;
  assign new_A4001_ = ~new_A3966_ & ~new_A4000_;
  assign new_A4002_ = new_A3966_ | new_A3999_;
  assign new_A4003_ = ~new_A3956_ & new_A3957_;
  assign new_A4004_ = new_A3956_ & ~new_A3957_;
  assign new_A4005_ = new_A3973_ | new_A4010_;
  assign new_A4006_ = ~new_A3973_ & ~new_A4009_;
  assign new_A4007_ = new_A3956_ | new_A3973_;
  assign new_A4008_ = new_A3956_ | new_A3957_;
  assign new_A4009_ = new_A3973_ & new_A4010_;
  assign new_A4010_ = ~new_A3955_ | ~new_A3980_;
  assign new_A4011_ = new_A3988_ & new_A4008_;
  assign new_A4012_ = ~new_A3988_ & ~new_A4008_;
  assign new_A4013_ = new_A4017_ | new_A4018_;
  assign new_A4014_ = ~new_A3959_ & new_A3973_;
  assign new_A4015_ = new_A4019_ | new_A4020_;
  assign new_A4016_ = new_A3959_ & new_A3973_;
  assign new_A4017_ = ~new_A3959_ & ~new_A3973_;
  assign new_A4018_ = new_A3959_ & ~new_A3973_;
  assign new_A4019_ = new_A3959_ & ~new_A3973_;
  assign new_A4020_ = ~new_A3959_ & new_A3973_;
  assign new_A4021_ = new_A5638_;
  assign new_A4022_ = new_A5704_;
  assign new_A4023_ = new_A5771_;
  assign new_A4024_ = new_A5838_;
  assign new_A4025_ = new_A5905_;
  assign new_A4026_ = new_A5972_;
  assign new_A4027_ = new_A4034_ & new_A4033_;
  assign new_A4028_ = new_A4036_ | new_A4035_;
  assign new_A4029_ = new_A4038_ | new_A4037_;
  assign new_A4030_ = new_A4040_ & new_A4039_;
  assign new_A4031_ = new_A4040_ & new_A4041_;
  assign new_A4032_ = new_A4033_ | new_A4042_;
  assign new_A4033_ = new_A4022_ | new_A4045_;
  assign new_A4034_ = new_A4044_ | new_A4043_;
  assign new_A4035_ = new_A4049_ & new_A4048_;
  assign new_A4036_ = new_A4047_ & new_A4046_;
  assign new_A4037_ = new_A4052_ | new_A4051_;
  assign new_A4038_ = new_A4047_ & new_A4050_;
  assign new_A4039_ = new_A4022_ | new_A4055_;
  assign new_A4040_ = new_A4054_ | new_A4053_;
  assign new_A4041_ = new_A4057_ | new_A4056_;
  assign new_A4042_ = ~new_A4033_ & new_A4059_;
  assign new_A4043_ = ~new_A4035_ & new_A4047_;
  assign new_A4044_ = new_A4035_ & ~new_A4047_;
  assign new_A4045_ = new_A4021_ & ~new_A4022_;
  assign new_A4046_ = ~new_A4068_ | ~new_A4069_;
  assign new_A4047_ = new_A4061_ | new_A4063_;
  assign new_A4048_ = new_A4071_ | new_A4070_;
  assign new_A4049_ = new_A4065_ | new_A4064_;
  assign new_A4050_ = ~new_A4073_ | ~new_A4072_;
  assign new_A4051_ = ~new_A4074_ & new_A4075_;
  assign new_A4052_ = new_A4074_ & ~new_A4075_;
  assign new_A4053_ = ~new_A4021_ & new_A4022_;
  assign new_A4054_ = new_A4021_ & ~new_A4022_;
  assign new_A4055_ = ~new_A4037_ | new_A4047_;
  assign new_A4056_ = new_A4037_ & new_A4047_;
  assign new_A4057_ = ~new_A4037_ & ~new_A4047_;
  assign new_A4058_ = new_A4079_ | new_A4078_;
  assign new_A4059_ = new_A4025_ | new_A4058_;
  assign new_A4060_ = new_A4083_ | new_A4082_;
  assign new_A4061_ = ~new_A4025_ & new_A4060_;
  assign new_A4062_ = new_A4081_ | new_A4080_;
  assign new_A4063_ = new_A4025_ & new_A4062_;
  assign new_A4064_ = new_A4023_ & ~new_A4033_;
  assign new_A4065_ = ~new_A4023_ & new_A4033_;
  assign new_A4066_ = ~new_A4022_ | ~new_A4047_;
  assign new_A4067_ = new_A4033_ & new_A4066_;
  assign new_A4068_ = ~new_A4033_ & ~new_A4067_;
  assign new_A4069_ = new_A4033_ | new_A4066_;
  assign new_A4070_ = ~new_A4023_ & new_A4024_;
  assign new_A4071_ = new_A4023_ & ~new_A4024_;
  assign new_A4072_ = new_A4040_ | new_A4077_;
  assign new_A4073_ = ~new_A4040_ & ~new_A4076_;
  assign new_A4074_ = new_A4023_ | new_A4040_;
  assign new_A4075_ = new_A4023_ | new_A4024_;
  assign new_A4076_ = new_A4040_ & new_A4077_;
  assign new_A4077_ = ~new_A4022_ | ~new_A4047_;
  assign new_A4078_ = new_A4055_ & new_A4075_;
  assign new_A4079_ = ~new_A4055_ & ~new_A4075_;
  assign new_A4080_ = new_A4084_ | new_A4085_;
  assign new_A4081_ = ~new_A4026_ & new_A4040_;
  assign new_A4082_ = new_A4086_ | new_A4087_;
  assign new_A4083_ = new_A4026_ & new_A4040_;
  assign new_A4084_ = ~new_A4026_ & ~new_A4040_;
  assign new_A4085_ = new_A4026_ & ~new_A4040_;
  assign new_A4086_ = new_A4026_ & ~new_A4040_;
  assign new_A4087_ = ~new_A4026_ & new_A4040_;
  assign new_A4088_ = new_A6039_;
  assign new_A4089_ = new_A6106_;
  assign new_A4090_ = new_A6173_;
  assign new_A4091_ = new_A6240_;
  assign new_A4092_ = new_A6307_;
  assign new_A4093_ = new_A6374_;
  assign new_A4094_ = new_A4101_ & new_A4100_;
  assign new_A4095_ = new_A4103_ | new_A4102_;
  assign new_A4096_ = new_A4105_ | new_A4104_;
  assign new_A4097_ = new_A4107_ & new_A4106_;
  assign new_A4098_ = new_A4107_ & new_A4108_;
  assign new_A4099_ = new_A4100_ | new_A4109_;
  assign new_A4100_ = new_A4089_ | new_A4112_;
  assign new_A4101_ = new_A4111_ | new_A4110_;
  assign new_A4102_ = new_A4116_ & new_A4115_;
  assign new_A4103_ = new_A4114_ & new_A4113_;
  assign new_A4104_ = new_A4119_ | new_A4118_;
  assign new_A4105_ = new_A4114_ & new_A4117_;
  assign new_A4106_ = new_A4089_ | new_A4122_;
  assign new_A4107_ = new_A4121_ | new_A4120_;
  assign new_A4108_ = new_A4124_ | new_A4123_;
  assign new_A4109_ = ~new_A4100_ & new_A4126_;
  assign new_A4110_ = ~new_A4102_ & new_A4114_;
  assign new_A4111_ = new_A4102_ & ~new_A4114_;
  assign new_A4112_ = new_A4088_ & ~new_A4089_;
  assign new_A4113_ = ~new_A4135_ | ~new_A4136_;
  assign new_A4114_ = new_A4128_ | new_A4130_;
  assign new_A4115_ = new_A4138_ | new_A4137_;
  assign new_A4116_ = new_A4132_ | new_A4131_;
  assign new_A4117_ = ~new_A4140_ | ~new_A4139_;
  assign new_A4118_ = ~new_A4141_ & new_A4142_;
  assign new_A4119_ = new_A4141_ & ~new_A4142_;
  assign new_A4120_ = ~new_A4088_ & new_A4089_;
  assign new_A4121_ = new_A4088_ & ~new_A4089_;
  assign new_A4122_ = ~new_A4104_ | new_A4114_;
  assign new_A4123_ = new_A4104_ & new_A4114_;
  assign new_A4124_ = ~new_A4104_ & ~new_A4114_;
  assign new_A4125_ = new_A4146_ | new_A4145_;
  assign new_A4126_ = new_A4092_ | new_A4125_;
  assign new_A4127_ = new_A4150_ | new_A4149_;
  assign new_A4128_ = ~new_A4092_ & new_A4127_;
  assign new_A4129_ = new_A4148_ | new_A4147_;
  assign new_A4130_ = new_A4092_ & new_A4129_;
  assign new_A4131_ = new_A4090_ & ~new_A4100_;
  assign new_A4132_ = ~new_A4090_ & new_A4100_;
  assign new_A4133_ = ~new_A4089_ | ~new_A4114_;
  assign new_A4134_ = new_A4100_ & new_A4133_;
  assign new_A4135_ = ~new_A4100_ & ~new_A4134_;
  assign new_A4136_ = new_A4100_ | new_A4133_;
  assign new_A4137_ = ~new_A4090_ & new_A4091_;
  assign new_A4138_ = new_A4090_ & ~new_A4091_;
  assign new_A4139_ = new_A4107_ | new_A4144_;
  assign new_A4140_ = ~new_A4107_ & ~new_A4143_;
  assign new_A4141_ = new_A4090_ | new_A4107_;
  assign new_A4142_ = new_A4090_ | new_A4091_;
  assign new_A4143_ = new_A4107_ & new_A4144_;
  assign new_A4144_ = ~new_A4089_ | ~new_A4114_;
  assign new_A4145_ = new_A4122_ & new_A4142_;
  assign new_A4146_ = ~new_A4122_ & ~new_A4142_;
  assign new_A4147_ = new_A4151_ | new_A4152_;
  assign new_A4148_ = ~new_A4093_ & new_A4107_;
  assign new_A4149_ = new_A4153_ | new_A4154_;
  assign new_A4150_ = new_A4093_ & new_A4107_;
  assign new_A4151_ = ~new_A4093_ & ~new_A4107_;
  assign new_A4152_ = new_A4093_ & ~new_A4107_;
  assign new_A4153_ = new_A4093_ & ~new_A4107_;
  assign new_A4154_ = ~new_A4093_ & new_A4107_;
  assign new_A4155_ = new_A6441_;
  assign new_A4156_ = new_A6508_;
  assign new_A4157_ = new_A6575_;
  assign new_A4158_ = new_A6642_;
  assign new_A4159_ = new_A6709_;
  assign new_A4160_ = new_A6776_;
  assign new_A4161_ = new_A4168_ & new_A4167_;
  assign new_A4162_ = new_A4170_ | new_A4169_;
  assign new_A4163_ = new_A4172_ | new_A4171_;
  assign new_A4164_ = new_A4174_ & new_A4173_;
  assign new_A4165_ = new_A4174_ & new_A4175_;
  assign new_A4166_ = new_A4167_ | new_A4176_;
  assign new_A4167_ = new_A4156_ | new_A4179_;
  assign new_A4168_ = new_A4178_ | new_A4177_;
  assign new_A4169_ = new_A4183_ & new_A4182_;
  assign new_A4170_ = new_A4181_ & new_A4180_;
  assign new_A4171_ = new_A4186_ | new_A4185_;
  assign new_A4172_ = new_A4181_ & new_A4184_;
  assign new_A4173_ = new_A4156_ | new_A4189_;
  assign new_A4174_ = new_A4188_ | new_A4187_;
  assign new_A4175_ = new_A4191_ | new_A4190_;
  assign new_A4176_ = ~new_A4167_ & new_A4193_;
  assign new_A4177_ = ~new_A4169_ & new_A4181_;
  assign new_A4178_ = new_A4169_ & ~new_A4181_;
  assign new_A4179_ = new_A4155_ & ~new_A4156_;
  assign new_A4180_ = ~new_A4202_ | ~new_A4203_;
  assign new_A4181_ = new_A4195_ | new_A4197_;
  assign new_A4182_ = new_A4205_ | new_A4204_;
  assign new_A4183_ = new_A4199_ | new_A4198_;
  assign new_A4184_ = ~new_A4207_ | ~new_A4206_;
  assign new_A4185_ = ~new_A4208_ & new_A4209_;
  assign new_A4186_ = new_A4208_ & ~new_A4209_;
  assign new_A4187_ = ~new_A4155_ & new_A4156_;
  assign new_A4188_ = new_A4155_ & ~new_A4156_;
  assign new_A4189_ = ~new_A4171_ | new_A4181_;
  assign new_A4190_ = new_A4171_ & new_A4181_;
  assign new_A4191_ = ~new_A4171_ & ~new_A4181_;
  assign new_A4192_ = new_A4213_ | new_A4212_;
  assign new_A4193_ = new_A4159_ | new_A4192_;
  assign new_A4194_ = new_A4217_ | new_A4216_;
  assign new_A4195_ = ~new_A4159_ & new_A4194_;
  assign new_A4196_ = new_A4215_ | new_A4214_;
  assign new_A4197_ = new_A4159_ & new_A4196_;
  assign new_A4198_ = new_A4157_ & ~new_A4167_;
  assign new_A4199_ = ~new_A4157_ & new_A4167_;
  assign new_A4200_ = ~new_A4156_ | ~new_A4181_;
  assign new_A4201_ = new_A4167_ & new_A4200_;
  assign new_A4202_ = ~new_A4167_ & ~new_A4201_;
  assign new_A4203_ = new_A4167_ | new_A4200_;
  assign new_A4204_ = ~new_A4157_ & new_A4158_;
  assign new_A4205_ = new_A4157_ & ~new_A4158_;
  assign new_A4206_ = new_A4174_ | new_A4211_;
  assign new_A4207_ = ~new_A4174_ & ~new_A4210_;
  assign new_A4208_ = new_A4157_ | new_A4174_;
  assign new_A4209_ = new_A4157_ | new_A4158_;
  assign new_A4210_ = new_A4174_ & new_A4211_;
  assign new_A4211_ = ~new_A4156_ | ~new_A4181_;
  assign new_A4212_ = new_A4189_ & new_A4209_;
  assign new_A4213_ = ~new_A4189_ & ~new_A4209_;
  assign new_A4214_ = new_A4218_ | new_A4219_;
  assign new_A4215_ = ~new_A4160_ & new_A4174_;
  assign new_A4216_ = new_A4220_ | new_A4221_;
  assign new_A4217_ = new_A4160_ & new_A4174_;
  assign new_A4218_ = ~new_A4160_ & ~new_A4174_;
  assign new_A4219_ = new_A4160_ & ~new_A4174_;
  assign new_A4220_ = new_A4160_ & ~new_A4174_;
  assign new_A4221_ = ~new_A4160_ & new_A4174_;
  assign new_A4222_ = new_A6843_;
  assign new_A4223_ = new_A6910_;
  assign new_A4224_ = new_A6977_;
  assign new_A4225_ = new_A7044_;
  assign new_A4226_ = new_A7111_;
  assign new_A4227_ = new_A7178_;
  assign new_A4228_ = new_A4235_ & new_A4234_;
  assign new_A4229_ = new_A4237_ | new_A4236_;
  assign new_A4230_ = new_A4239_ | new_A4238_;
  assign new_A4231_ = new_A4241_ & new_A4240_;
  assign new_A4232_ = new_A4241_ & new_A4242_;
  assign new_A4233_ = new_A4234_ | new_A4243_;
  assign new_A4234_ = new_A4223_ | new_A4246_;
  assign new_A4235_ = new_A4245_ | new_A4244_;
  assign new_A4236_ = new_A4250_ & new_A4249_;
  assign new_A4237_ = new_A4248_ & new_A4247_;
  assign new_A4238_ = new_A4253_ | new_A4252_;
  assign new_A4239_ = new_A4248_ & new_A4251_;
  assign new_A4240_ = new_A4223_ | new_A4256_;
  assign new_A4241_ = new_A4255_ | new_A4254_;
  assign new_A4242_ = new_A4258_ | new_A4257_;
  assign new_A4243_ = ~new_A4234_ & new_A4260_;
  assign new_A4244_ = ~new_A4236_ & new_A4248_;
  assign new_A4245_ = new_A4236_ & ~new_A4248_;
  assign new_A4246_ = new_A4222_ & ~new_A4223_;
  assign new_A4247_ = ~new_A4269_ | ~new_A4270_;
  assign new_A4248_ = new_A4262_ | new_A4264_;
  assign new_A4249_ = new_A4272_ | new_A4271_;
  assign new_A4250_ = new_A4266_ | new_A4265_;
  assign new_A4251_ = ~new_A4274_ | ~new_A4273_;
  assign new_A4252_ = ~new_A4275_ & new_A4276_;
  assign new_A4253_ = new_A4275_ & ~new_A4276_;
  assign new_A4254_ = ~new_A4222_ & new_A4223_;
  assign new_A4255_ = new_A4222_ & ~new_A4223_;
  assign new_A4256_ = ~new_A4238_ | new_A4248_;
  assign new_A4257_ = new_A4238_ & new_A4248_;
  assign new_A4258_ = ~new_A4238_ & ~new_A4248_;
  assign new_A4259_ = new_A4280_ | new_A4279_;
  assign new_A4260_ = new_A4226_ | new_A4259_;
  assign new_A4261_ = new_A4284_ | new_A4283_;
  assign new_A4262_ = ~new_A4226_ & new_A4261_;
  assign new_A4263_ = new_A4282_ | new_A4281_;
  assign new_A4264_ = new_A4226_ & new_A4263_;
  assign new_A4265_ = new_A4224_ & ~new_A4234_;
  assign new_A4266_ = ~new_A4224_ & new_A4234_;
  assign new_A4267_ = ~new_A4223_ | ~new_A4248_;
  assign new_A4268_ = new_A4234_ & new_A4267_;
  assign new_A4269_ = ~new_A4234_ & ~new_A4268_;
  assign new_A4270_ = new_A4234_ | new_A4267_;
  assign new_A4271_ = ~new_A4224_ & new_A4225_;
  assign new_A4272_ = new_A4224_ & ~new_A4225_;
  assign new_A4273_ = new_A4241_ | new_A4278_;
  assign new_A4274_ = ~new_A4241_ & ~new_A4277_;
  assign new_A4275_ = new_A4224_ | new_A4241_;
  assign new_A4276_ = new_A4224_ | new_A4225_;
  assign new_A4277_ = new_A4241_ & new_A4278_;
  assign new_A4278_ = ~new_A4223_ | ~new_A4248_;
  assign new_A4279_ = new_A4256_ & new_A4276_;
  assign new_A4280_ = ~new_A4256_ & ~new_A4276_;
  assign new_A4281_ = new_A4285_ | new_A4286_;
  assign new_A4282_ = ~new_A4227_ & new_A4241_;
  assign new_A4283_ = new_A4287_ | new_A4288_;
  assign new_A4284_ = new_A4227_ & new_A4241_;
  assign new_A4285_ = ~new_A4227_ & ~new_A4241_;
  assign new_A4286_ = new_A4227_ & ~new_A4241_;
  assign new_A4287_ = new_A4227_ & ~new_A4241_;
  assign new_A4288_ = ~new_A4227_ & new_A4241_;
  assign new_A4289_ = new_A7245_;
  assign new_A4290_ = new_A7312_;
  assign new_A4291_ = new_A7379_;
  assign new_A4292_ = new_A7446_;
  assign new_A4293_ = new_A7513_;
  assign new_A4294_ = new_A7580_;
  assign new_A4295_ = new_A4302_ & new_A4301_;
  assign new_A4296_ = new_A4304_ | new_A4303_;
  assign new_A4297_ = new_A4306_ | new_A4305_;
  assign new_A4298_ = new_A4308_ & new_A4307_;
  assign new_A4299_ = new_A4308_ & new_A4309_;
  assign new_A4300_ = new_A4301_ | new_A4310_;
  assign new_A4301_ = new_A4290_ | new_A4313_;
  assign new_A4302_ = new_A4312_ | new_A4311_;
  assign new_A4303_ = new_A4317_ & new_A4316_;
  assign new_A4304_ = new_A4315_ & new_A4314_;
  assign new_A4305_ = new_A4320_ | new_A4319_;
  assign new_A4306_ = new_A4315_ & new_A4318_;
  assign new_A4307_ = new_A4290_ | new_A4323_;
  assign new_A4308_ = new_A4322_ | new_A4321_;
  assign new_A4309_ = new_A4325_ | new_A4324_;
  assign new_A4310_ = ~new_A4301_ & new_A4327_;
  assign new_A4311_ = ~new_A4303_ & new_A4315_;
  assign new_A4312_ = new_A4303_ & ~new_A4315_;
  assign new_A4313_ = new_A4289_ & ~new_A4290_;
  assign new_A4314_ = ~new_A4336_ | ~new_A4337_;
  assign new_A4315_ = new_A4329_ | new_A4331_;
  assign new_A4316_ = new_A4339_ | new_A4338_;
  assign new_A4317_ = new_A4333_ | new_A4332_;
  assign new_A4318_ = ~new_A4341_ | ~new_A4340_;
  assign new_A4319_ = ~new_A4342_ & new_A4343_;
  assign new_A4320_ = new_A4342_ & ~new_A4343_;
  assign new_A4321_ = ~new_A4289_ & new_A4290_;
  assign new_A4322_ = new_A4289_ & ~new_A4290_;
  assign new_A4323_ = ~new_A4305_ | new_A4315_;
  assign new_A4324_ = new_A4305_ & new_A4315_;
  assign new_A4325_ = ~new_A4305_ & ~new_A4315_;
  assign new_A4326_ = new_A4347_ | new_A4346_;
  assign new_A4327_ = new_A4293_ | new_A4326_;
  assign new_A4328_ = new_A4351_ | new_A4350_;
  assign new_A4329_ = ~new_A4293_ & new_A4328_;
  assign new_A4330_ = new_A4349_ | new_A4348_;
  assign new_A4331_ = new_A4293_ & new_A4330_;
  assign new_A4332_ = new_A4291_ & ~new_A4301_;
  assign new_A4333_ = ~new_A4291_ & new_A4301_;
  assign new_A4334_ = ~new_A4290_ | ~new_A4315_;
  assign new_A4335_ = new_A4301_ & new_A4334_;
  assign new_A4336_ = ~new_A4301_ & ~new_A4335_;
  assign new_A4337_ = new_A4301_ | new_A4334_;
  assign new_A4338_ = ~new_A4291_ & new_A4292_;
  assign new_A4339_ = new_A4291_ & ~new_A4292_;
  assign new_A4340_ = new_A4308_ | new_A4345_;
  assign new_A4341_ = ~new_A4308_ & ~new_A4344_;
  assign new_A4342_ = new_A4291_ | new_A4308_;
  assign new_A4343_ = new_A4291_ | new_A4292_;
  assign new_A4344_ = new_A4308_ & new_A4345_;
  assign new_A4345_ = ~new_A4290_ | ~new_A4315_;
  assign new_A4346_ = new_A4323_ & new_A4343_;
  assign new_A4347_ = ~new_A4323_ & ~new_A4343_;
  assign new_A4348_ = new_A4352_ | new_A4353_;
  assign new_A4349_ = ~new_A4294_ & new_A4308_;
  assign new_A4350_ = new_A4354_ | new_A4355_;
  assign new_A4351_ = new_A4294_ & new_A4308_;
  assign new_A4352_ = ~new_A4294_ & ~new_A4308_;
  assign new_A4353_ = new_A4294_ & ~new_A4308_;
  assign new_A4354_ = new_A4294_ & ~new_A4308_;
  assign new_A4355_ = ~new_A4294_ & new_A4308_;
  assign new_A4356_ = new_A7647_;
  assign new_A4357_ = new_A7714_;
  assign new_A4358_ = new_A7781_;
  assign new_A4359_ = new_A7848_;
  assign new_A4360_ = new_A7915_;
  assign new_A4361_ = new_A7982_;
  assign new_A4362_ = new_A4369_ & new_A4368_;
  assign new_A4363_ = new_A4371_ | new_A4370_;
  assign new_A4364_ = new_A4373_ | new_A4372_;
  assign new_A4365_ = new_A4375_ & new_A4374_;
  assign new_A4366_ = new_A4375_ & new_A4376_;
  assign new_A4367_ = new_A4368_ | new_A4377_;
  assign new_A4368_ = new_A4357_ | new_A4380_;
  assign new_A4369_ = new_A4379_ | new_A4378_;
  assign new_A4370_ = new_A4384_ & new_A4383_;
  assign new_A4371_ = new_A4382_ & new_A4381_;
  assign new_A4372_ = new_A4387_ | new_A4386_;
  assign new_A4373_ = new_A4382_ & new_A4385_;
  assign new_A4374_ = new_A4357_ | new_A4390_;
  assign new_A4375_ = new_A4389_ | new_A4388_;
  assign new_A4376_ = new_A4392_ | new_A4391_;
  assign new_A4377_ = ~new_A4368_ & new_A4394_;
  assign new_A4378_ = ~new_A4370_ & new_A4382_;
  assign new_A4379_ = new_A4370_ & ~new_A4382_;
  assign new_A4380_ = new_A4356_ & ~new_A4357_;
  assign new_A4381_ = ~new_A4403_ | ~new_A4404_;
  assign new_A4382_ = new_A4396_ | new_A4398_;
  assign new_A4383_ = new_A4406_ | new_A4405_;
  assign new_A4384_ = new_A4400_ | new_A4399_;
  assign new_A4385_ = ~new_A4408_ | ~new_A4407_;
  assign new_A4386_ = ~new_A4409_ & new_A4410_;
  assign new_A4387_ = new_A4409_ & ~new_A4410_;
  assign new_A4388_ = ~new_A4356_ & new_A4357_;
  assign new_A4389_ = new_A4356_ & ~new_A4357_;
  assign new_A4390_ = ~new_A4372_ | new_A4382_;
  assign new_A4391_ = new_A4372_ & new_A4382_;
  assign new_A4392_ = ~new_A4372_ & ~new_A4382_;
  assign new_A4393_ = new_A4414_ | new_A4413_;
  assign new_A4394_ = new_A4360_ | new_A4393_;
  assign new_A4395_ = new_A4418_ | new_A4417_;
  assign new_A4396_ = ~new_A4360_ & new_A4395_;
  assign new_A4397_ = new_A4416_ | new_A4415_;
  assign new_A4398_ = new_A4360_ & new_A4397_;
  assign new_A4399_ = new_A4358_ & ~new_A4368_;
  assign new_A4400_ = ~new_A4358_ & new_A4368_;
  assign new_A4401_ = ~new_A4357_ | ~new_A4382_;
  assign new_A4402_ = new_A4368_ & new_A4401_;
  assign new_A4403_ = ~new_A4368_ & ~new_A4402_;
  assign new_A4404_ = new_A4368_ | new_A4401_;
  assign new_A4405_ = ~new_A4358_ & new_A4359_;
  assign new_A4406_ = new_A4358_ & ~new_A4359_;
  assign new_A4407_ = new_A4375_ | new_A4412_;
  assign new_A4408_ = ~new_A4375_ & ~new_A4411_;
  assign new_A4409_ = new_A4358_ | new_A4375_;
  assign new_A4410_ = new_A4358_ | new_A4359_;
  assign new_A4411_ = new_A4375_ & new_A4412_;
  assign new_A4412_ = ~new_A4357_ | ~new_A4382_;
  assign new_A4413_ = new_A4390_ & new_A4410_;
  assign new_A4414_ = ~new_A4390_ & ~new_A4410_;
  assign new_A4415_ = new_A4419_ | new_A4420_;
  assign new_A4416_ = ~new_A4361_ & new_A4375_;
  assign new_A4417_ = new_A4421_ | new_A4422_;
  assign new_A4418_ = new_A4361_ & new_A4375_;
  assign new_A4419_ = ~new_A4361_ & ~new_A4375_;
  assign new_A4420_ = new_A4361_ & ~new_A4375_;
  assign new_A4421_ = new_A4361_ & ~new_A4375_;
  assign new_A4422_ = ~new_A4361_ & new_A4375_;
  assign new_A4423_ = new_A5637_;
  assign new_A4424_ = new_A5705_;
  assign new_A4425_ = new_A5772_;
  assign new_A4426_ = new_A5839_;
  assign new_A4427_ = new_A5906_;
  assign new_A4428_ = new_A5973_;
  assign new_A4429_ = new_A4436_ & new_A4435_;
  assign new_A4430_ = new_A4438_ | new_A4437_;
  assign new_A4431_ = new_A4440_ | new_A4439_;
  assign new_A4432_ = new_A4442_ & new_A4441_;
  assign new_A4433_ = new_A4442_ & new_A4443_;
  assign new_A4434_ = new_A4435_ | new_A4444_;
  assign new_A4435_ = new_A4424_ | new_A4447_;
  assign new_A4436_ = new_A4446_ | new_A4445_;
  assign new_A4437_ = new_A4451_ & new_A4450_;
  assign new_A4438_ = new_A4449_ & new_A4448_;
  assign new_A4439_ = new_A4454_ | new_A4453_;
  assign new_A4440_ = new_A4449_ & new_A4452_;
  assign new_A4441_ = new_A4424_ | new_A4457_;
  assign new_A4442_ = new_A4456_ | new_A4455_;
  assign new_A4443_ = new_A4459_ | new_A4458_;
  assign new_A4444_ = ~new_A4435_ & new_A4461_;
  assign new_A4445_ = ~new_A4437_ & new_A4449_;
  assign new_A4446_ = new_A4437_ & ~new_A4449_;
  assign new_A4447_ = new_A4423_ & ~new_A4424_;
  assign new_A4448_ = ~new_A4470_ | ~new_A4471_;
  assign new_A4449_ = new_A4463_ | new_A4465_;
  assign new_A4450_ = new_A4473_ | new_A4472_;
  assign new_A4451_ = new_A4467_ | new_A4466_;
  assign new_A4452_ = ~new_A4475_ | ~new_A4474_;
  assign new_A4453_ = ~new_A4476_ & new_A4477_;
  assign new_A4454_ = new_A4476_ & ~new_A4477_;
  assign new_A4455_ = ~new_A4423_ & new_A4424_;
  assign new_A4456_ = new_A4423_ & ~new_A4424_;
  assign new_A4457_ = ~new_A4439_ | new_A4449_;
  assign new_A4458_ = new_A4439_ & new_A4449_;
  assign new_A4459_ = ~new_A4439_ & ~new_A4449_;
  assign new_A4460_ = new_A4481_ | new_A4480_;
  assign new_A4461_ = new_A4427_ | new_A4460_;
  assign new_A4462_ = new_A4485_ | new_A4484_;
  assign new_A4463_ = ~new_A4427_ & new_A4462_;
  assign new_A4464_ = new_A4483_ | new_A4482_;
  assign new_A4465_ = new_A4427_ & new_A4464_;
  assign new_A4466_ = new_A4425_ & ~new_A4435_;
  assign new_A4467_ = ~new_A4425_ & new_A4435_;
  assign new_A4468_ = ~new_A4424_ | ~new_A4449_;
  assign new_A4469_ = new_A4435_ & new_A4468_;
  assign new_A4470_ = ~new_A4435_ & ~new_A4469_;
  assign new_A4471_ = new_A4435_ | new_A4468_;
  assign new_A4472_ = ~new_A4425_ & new_A4426_;
  assign new_A4473_ = new_A4425_ & ~new_A4426_;
  assign new_A4474_ = new_A4442_ | new_A4479_;
  assign new_A4475_ = ~new_A4442_ & ~new_A4478_;
  assign new_A4476_ = new_A4425_ | new_A4442_;
  assign new_A4477_ = new_A4425_ | new_A4426_;
  assign new_A4478_ = new_A4442_ & new_A4479_;
  assign new_A4479_ = ~new_A4424_ | ~new_A4449_;
  assign new_A4480_ = new_A4457_ & new_A4477_;
  assign new_A4481_ = ~new_A4457_ & ~new_A4477_;
  assign new_A4482_ = new_A4486_ | new_A4487_;
  assign new_A4483_ = ~new_A4428_ & new_A4442_;
  assign new_A4484_ = new_A4488_ | new_A4489_;
  assign new_A4485_ = new_A4428_ & new_A4442_;
  assign new_A4486_ = ~new_A4428_ & ~new_A4442_;
  assign new_A4487_ = new_A4428_ & ~new_A4442_;
  assign new_A4488_ = new_A4428_ & ~new_A4442_;
  assign new_A4489_ = ~new_A4428_ & new_A4442_;
  assign new_A4490_ = new_A6040_;
  assign new_A4491_ = new_A6107_;
  assign new_A4492_ = new_A6174_;
  assign new_A4493_ = new_A6241_;
  assign new_A4494_ = new_A6308_;
  assign new_A4495_ = new_A6375_;
  assign new_A4496_ = new_A4503_ & new_A4502_;
  assign new_A4497_ = new_A4505_ | new_A4504_;
  assign new_A4498_ = new_A4507_ | new_A4506_;
  assign new_A4499_ = new_A4509_ & new_A4508_;
  assign new_A4500_ = new_A4509_ & new_A4510_;
  assign new_A4501_ = new_A4502_ | new_A4511_;
  assign new_A4502_ = new_A4491_ | new_A4514_;
  assign new_A4503_ = new_A4513_ | new_A4512_;
  assign new_A4504_ = new_A4518_ & new_A4517_;
  assign new_A4505_ = new_A4516_ & new_A4515_;
  assign new_A4506_ = new_A4521_ | new_A4520_;
  assign new_A4507_ = new_A4516_ & new_A4519_;
  assign new_A4508_ = new_A4491_ | new_A4524_;
  assign new_A4509_ = new_A4523_ | new_A4522_;
  assign new_A4510_ = new_A4526_ | new_A4525_;
  assign new_A4511_ = ~new_A4502_ & new_A4528_;
  assign new_A4512_ = ~new_A4504_ & new_A4516_;
  assign new_A4513_ = new_A4504_ & ~new_A4516_;
  assign new_A4514_ = new_A4490_ & ~new_A4491_;
  assign new_A4515_ = ~new_A4537_ | ~new_A4538_;
  assign new_A4516_ = new_A4530_ | new_A4532_;
  assign new_A4517_ = new_A4540_ | new_A4539_;
  assign new_A4518_ = new_A4534_ | new_A4533_;
  assign new_A4519_ = ~new_A4542_ | ~new_A4541_;
  assign new_A4520_ = ~new_A4543_ & new_A4544_;
  assign new_A4521_ = new_A4543_ & ~new_A4544_;
  assign new_A4522_ = ~new_A4490_ & new_A4491_;
  assign new_A4523_ = new_A4490_ & ~new_A4491_;
  assign new_A4524_ = ~new_A4506_ | new_A4516_;
  assign new_A4525_ = new_A4506_ & new_A4516_;
  assign new_A4526_ = ~new_A4506_ & ~new_A4516_;
  assign new_A4527_ = new_A4548_ | new_A4547_;
  assign new_A4528_ = new_A4494_ | new_A4527_;
  assign new_A4529_ = new_A4552_ | new_A4551_;
  assign new_A4530_ = ~new_A4494_ & new_A4529_;
  assign new_A4531_ = new_A4550_ | new_A4549_;
  assign new_A4532_ = new_A4494_ & new_A4531_;
  assign new_A4533_ = new_A4492_ & ~new_A4502_;
  assign new_A4534_ = ~new_A4492_ & new_A4502_;
  assign new_A4535_ = ~new_A4491_ | ~new_A4516_;
  assign new_A4536_ = new_A4502_ & new_A4535_;
  assign new_A4537_ = ~new_A4502_ & ~new_A4536_;
  assign new_A4538_ = new_A4502_ | new_A4535_;
  assign new_A4539_ = ~new_A4492_ & new_A4493_;
  assign new_A4540_ = new_A4492_ & ~new_A4493_;
  assign new_A4541_ = new_A4509_ | new_A4546_;
  assign new_A4542_ = ~new_A4509_ & ~new_A4545_;
  assign new_A4543_ = new_A4492_ | new_A4509_;
  assign new_A4544_ = new_A4492_ | new_A4493_;
  assign new_A4545_ = new_A4509_ & new_A4546_;
  assign new_A4546_ = ~new_A4491_ | ~new_A4516_;
  assign new_A4547_ = new_A4524_ & new_A4544_;
  assign new_A4548_ = ~new_A4524_ & ~new_A4544_;
  assign new_A4549_ = new_A4553_ | new_A4554_;
  assign new_A4550_ = ~new_A4495_ & new_A4509_;
  assign new_A4551_ = new_A4555_ | new_A4556_;
  assign new_A4552_ = new_A4495_ & new_A4509_;
  assign new_A4553_ = ~new_A4495_ & ~new_A4509_;
  assign new_A4554_ = new_A4495_ & ~new_A4509_;
  assign new_A4555_ = new_A4495_ & ~new_A4509_;
  assign new_A4556_ = ~new_A4495_ & new_A4509_;
  assign new_A4557_ = new_A6442_;
  assign new_A4558_ = new_A6509_;
  assign new_A4559_ = new_A6576_;
  assign new_A4560_ = new_A6643_;
  assign new_A4561_ = new_A6710_;
  assign new_A4562_ = new_A6777_;
  assign new_A4563_ = new_A4570_ & new_A4569_;
  assign new_A4564_ = new_A4572_ | new_A4571_;
  assign new_A4565_ = new_A4574_ | new_A4573_;
  assign new_A4566_ = new_A4576_ & new_A4575_;
  assign new_A4567_ = new_A4576_ & new_A4577_;
  assign new_A4568_ = new_A4569_ | new_A4578_;
  assign new_A4569_ = new_A4558_ | new_A4581_;
  assign new_A4570_ = new_A4580_ | new_A4579_;
  assign new_A4571_ = new_A4585_ & new_A4584_;
  assign new_A4572_ = new_A4583_ & new_A4582_;
  assign new_A4573_ = new_A4588_ | new_A4587_;
  assign new_A4574_ = new_A4583_ & new_A4586_;
  assign new_A4575_ = new_A4558_ | new_A4591_;
  assign new_A4576_ = new_A4590_ | new_A4589_;
  assign new_A4577_ = new_A4593_ | new_A4592_;
  assign new_A4578_ = ~new_A4569_ & new_A4595_;
  assign new_A4579_ = ~new_A4571_ & new_A4583_;
  assign new_A4580_ = new_A4571_ & ~new_A4583_;
  assign new_A4581_ = new_A4557_ & ~new_A4558_;
  assign new_A4582_ = ~new_A4604_ | ~new_A4605_;
  assign new_A4583_ = new_A4597_ | new_A4599_;
  assign new_A4584_ = new_A4607_ | new_A4606_;
  assign new_A4585_ = new_A4601_ | new_A4600_;
  assign new_A4586_ = ~new_A4609_ | ~new_A4608_;
  assign new_A4587_ = ~new_A4610_ & new_A4611_;
  assign new_A4588_ = new_A4610_ & ~new_A4611_;
  assign new_A4589_ = ~new_A4557_ & new_A4558_;
  assign new_A4590_ = new_A4557_ & ~new_A4558_;
  assign new_A4591_ = ~new_A4573_ | new_A4583_;
  assign new_A4592_ = new_A4573_ & new_A4583_;
  assign new_A4593_ = ~new_A4573_ & ~new_A4583_;
  assign new_A4594_ = new_A4615_ | new_A4614_;
  assign new_A4595_ = new_A4561_ | new_A4594_;
  assign new_A4596_ = new_A4619_ | new_A4618_;
  assign new_A4597_ = ~new_A4561_ & new_A4596_;
  assign new_A4598_ = new_A4617_ | new_A4616_;
  assign new_A4599_ = new_A4561_ & new_A4598_;
  assign new_A4600_ = new_A4559_ & ~new_A4569_;
  assign new_A4601_ = ~new_A4559_ & new_A4569_;
  assign new_A4602_ = ~new_A4558_ | ~new_A4583_;
  assign new_A4603_ = new_A4569_ & new_A4602_;
  assign new_A4604_ = ~new_A4569_ & ~new_A4603_;
  assign new_A4605_ = new_A4569_ | new_A4602_;
  assign new_A4606_ = ~new_A4559_ & new_A4560_;
  assign new_A4607_ = new_A4559_ & ~new_A4560_;
  assign new_A4608_ = new_A4576_ | new_A4613_;
  assign new_A4609_ = ~new_A4576_ & ~new_A4612_;
  assign new_A4610_ = new_A4559_ | new_A4576_;
  assign new_A4611_ = new_A4559_ | new_A4560_;
  assign new_A4612_ = new_A4576_ & new_A4613_;
  assign new_A4613_ = ~new_A4558_ | ~new_A4583_;
  assign new_A4614_ = new_A4591_ & new_A4611_;
  assign new_A4615_ = ~new_A4591_ & ~new_A4611_;
  assign new_A4616_ = new_A4620_ | new_A4621_;
  assign new_A4617_ = ~new_A4562_ & new_A4576_;
  assign new_A4618_ = new_A4622_ | new_A4623_;
  assign new_A4619_ = new_A4562_ & new_A4576_;
  assign new_A4620_ = ~new_A4562_ & ~new_A4576_;
  assign new_A4621_ = new_A4562_ & ~new_A4576_;
  assign new_A4622_ = new_A4562_ & ~new_A4576_;
  assign new_A4623_ = ~new_A4562_ & new_A4576_;
  assign new_A4624_ = new_A6844_;
  assign new_A4625_ = new_A6911_;
  assign new_A4626_ = new_A6978_;
  assign new_A4627_ = new_A7045_;
  assign new_A4628_ = new_A7112_;
  assign new_A4629_ = new_A7179_;
  assign new_A4630_ = new_A4637_ & new_A4636_;
  assign new_A4631_ = new_A4639_ | new_A4638_;
  assign new_A4632_ = new_A4641_ | new_A4640_;
  assign new_A4633_ = new_A4643_ & new_A4642_;
  assign new_A4634_ = new_A4643_ & new_A4644_;
  assign new_A4635_ = new_A4636_ | new_A4645_;
  assign new_A4636_ = new_A4625_ | new_A4648_;
  assign new_A4637_ = new_A4647_ | new_A4646_;
  assign new_A4638_ = new_A4652_ & new_A4651_;
  assign new_A4639_ = new_A4650_ & new_A4649_;
  assign new_A4640_ = new_A4655_ | new_A4654_;
  assign new_A4641_ = new_A4650_ & new_A4653_;
  assign new_A4642_ = new_A4625_ | new_A4658_;
  assign new_A4643_ = new_A4657_ | new_A4656_;
  assign new_A4644_ = new_A4660_ | new_A4659_;
  assign new_A4645_ = ~new_A4636_ & new_A4662_;
  assign new_A4646_ = ~new_A4638_ & new_A4650_;
  assign new_A4647_ = new_A4638_ & ~new_A4650_;
  assign new_A4648_ = new_A4624_ & ~new_A4625_;
  assign new_A4649_ = ~new_A4671_ | ~new_A4672_;
  assign new_A4650_ = new_A4664_ | new_A4666_;
  assign new_A4651_ = new_A4674_ | new_A4673_;
  assign new_A4652_ = new_A4668_ | new_A4667_;
  assign new_A4653_ = ~new_A4676_ | ~new_A4675_;
  assign new_A4654_ = ~new_A4677_ & new_A4678_;
  assign new_A4655_ = new_A4677_ & ~new_A4678_;
  assign new_A4656_ = ~new_A4624_ & new_A4625_;
  assign new_A4657_ = new_A4624_ & ~new_A4625_;
  assign new_A4658_ = ~new_A4640_ | new_A4650_;
  assign new_A4659_ = new_A4640_ & new_A4650_;
  assign new_A4660_ = ~new_A4640_ & ~new_A4650_;
  assign new_A4661_ = new_A4682_ | new_A4681_;
  assign new_A4662_ = new_A4628_ | new_A4661_;
  assign new_A4663_ = new_A4686_ | new_A4685_;
  assign new_A4664_ = ~new_A4628_ & new_A4663_;
  assign new_A4665_ = new_A4684_ | new_A4683_;
  assign new_A4666_ = new_A4628_ & new_A4665_;
  assign new_A4667_ = new_A4626_ & ~new_A4636_;
  assign new_A4668_ = ~new_A4626_ & new_A4636_;
  assign new_A4669_ = ~new_A4625_ | ~new_A4650_;
  assign new_A4670_ = new_A4636_ & new_A4669_;
  assign new_A4671_ = ~new_A4636_ & ~new_A4670_;
  assign new_A4672_ = new_A4636_ | new_A4669_;
  assign new_A4673_ = ~new_A4626_ & new_A4627_;
  assign new_A4674_ = new_A4626_ & ~new_A4627_;
  assign new_A4675_ = new_A4643_ | new_A4680_;
  assign new_A4676_ = ~new_A4643_ & ~new_A4679_;
  assign new_A4677_ = new_A4626_ | new_A4643_;
  assign new_A4678_ = new_A4626_ | new_A4627_;
  assign new_A4679_ = new_A4643_ & new_A4680_;
  assign new_A4680_ = ~new_A4625_ | ~new_A4650_;
  assign new_A4681_ = new_A4658_ & new_A4678_;
  assign new_A4682_ = ~new_A4658_ & ~new_A4678_;
  assign new_A4683_ = new_A4687_ | new_A4688_;
  assign new_A4684_ = ~new_A4629_ & new_A4643_;
  assign new_A4685_ = new_A4689_ | new_A4690_;
  assign new_A4686_ = new_A4629_ & new_A4643_;
  assign new_A4687_ = ~new_A4629_ & ~new_A4643_;
  assign new_A4688_ = new_A4629_ & ~new_A4643_;
  assign new_A4689_ = new_A4629_ & ~new_A4643_;
  assign new_A4690_ = ~new_A4629_ & new_A4643_;
  assign new_A4691_ = new_A7246_;
  assign new_A4692_ = new_A7313_;
  assign new_A4693_ = new_A7380_;
  assign new_A4694_ = new_A7447_;
  assign new_A4695_ = new_A7514_;
  assign new_A4696_ = new_A7581_;
  assign new_A4697_ = new_A4704_ & new_A4703_;
  assign new_A4698_ = new_A4706_ | new_A4705_;
  assign new_A4699_ = new_A4708_ | new_A4707_;
  assign new_A4700_ = new_A4710_ & new_A4709_;
  assign new_A4701_ = new_A4710_ & new_A4711_;
  assign new_A4702_ = new_A4703_ | new_A4712_;
  assign new_A4703_ = new_A4692_ | new_A4715_;
  assign new_A4704_ = new_A4714_ | new_A4713_;
  assign new_A4705_ = new_A4719_ & new_A4718_;
  assign new_A4706_ = new_A4717_ & new_A4716_;
  assign new_A4707_ = new_A4722_ | new_A4721_;
  assign new_A4708_ = new_A4717_ & new_A4720_;
  assign new_A4709_ = new_A4692_ | new_A4725_;
  assign new_A4710_ = new_A4724_ | new_A4723_;
  assign new_A4711_ = new_A4727_ | new_A4726_;
  assign new_A4712_ = ~new_A4703_ & new_A4729_;
  assign new_A4713_ = ~new_A4705_ & new_A4717_;
  assign new_A4714_ = new_A4705_ & ~new_A4717_;
  assign new_A4715_ = new_A4691_ & ~new_A4692_;
  assign new_A4716_ = ~new_A4738_ | ~new_A4739_;
  assign new_A4717_ = new_A4731_ | new_A4733_;
  assign new_A4718_ = new_A4741_ | new_A4740_;
  assign new_A4719_ = new_A4735_ | new_A4734_;
  assign new_A4720_ = ~new_A4743_ | ~new_A4742_;
  assign new_A4721_ = ~new_A4744_ & new_A4745_;
  assign new_A4722_ = new_A4744_ & ~new_A4745_;
  assign new_A4723_ = ~new_A4691_ & new_A4692_;
  assign new_A4724_ = new_A4691_ & ~new_A4692_;
  assign new_A4725_ = ~new_A4707_ | new_A4717_;
  assign new_A4726_ = new_A4707_ & new_A4717_;
  assign new_A4727_ = ~new_A4707_ & ~new_A4717_;
  assign new_A4728_ = new_A4749_ | new_A4748_;
  assign new_A4729_ = new_A4695_ | new_A4728_;
  assign new_A4730_ = new_A4753_ | new_A4752_;
  assign new_A4731_ = ~new_A4695_ & new_A4730_;
  assign new_A4732_ = new_A4751_ | new_A4750_;
  assign new_A4733_ = new_A4695_ & new_A4732_;
  assign new_A4734_ = new_A4693_ & ~new_A4703_;
  assign new_A4735_ = ~new_A4693_ & new_A4703_;
  assign new_A4736_ = ~new_A4692_ | ~new_A4717_;
  assign new_A4737_ = new_A4703_ & new_A4736_;
  assign new_A4738_ = ~new_A4703_ & ~new_A4737_;
  assign new_A4739_ = new_A4703_ | new_A4736_;
  assign new_A4740_ = ~new_A4693_ & new_A4694_;
  assign new_A4741_ = new_A4693_ & ~new_A4694_;
  assign new_A4742_ = new_A4710_ | new_A4747_;
  assign new_A4743_ = ~new_A4710_ & ~new_A4746_;
  assign new_A4744_ = new_A4693_ | new_A4710_;
  assign new_A4745_ = new_A4693_ | new_A4694_;
  assign new_A4746_ = new_A4710_ & new_A4747_;
  assign new_A4747_ = ~new_A4692_ | ~new_A4717_;
  assign new_A4748_ = new_A4725_ & new_A4745_;
  assign new_A4749_ = ~new_A4725_ & ~new_A4745_;
  assign new_A4750_ = new_A4754_ | new_A4755_;
  assign new_A4751_ = ~new_A4696_ & new_A4710_;
  assign new_A4752_ = new_A4756_ | new_A4757_;
  assign new_A4753_ = new_A4696_ & new_A4710_;
  assign new_A4754_ = ~new_A4696_ & ~new_A4710_;
  assign new_A4755_ = new_A4696_ & ~new_A4710_;
  assign new_A4756_ = new_A4696_ & ~new_A4710_;
  assign new_A4757_ = ~new_A4696_ & new_A4710_;
  assign new_A4758_ = new_A7648_;
  assign new_A4759_ = new_A7715_;
  assign new_A4760_ = new_A7782_;
  assign new_A4761_ = new_A7849_;
  assign new_A4762_ = new_A7916_;
  assign new_A4763_ = new_A7983_;
  assign new_A4764_ = new_A4771_ & new_A4770_;
  assign new_A4765_ = new_A4773_ | new_A4772_;
  assign new_A4766_ = new_A4775_ | new_A4774_;
  assign new_A4767_ = new_A4777_ & new_A4776_;
  assign new_A4768_ = new_A4777_ & new_A4778_;
  assign new_A4769_ = new_A4770_ | new_A4779_;
  assign new_A4770_ = new_A4759_ | new_A4782_;
  assign new_A4771_ = new_A4781_ | new_A4780_;
  assign new_A4772_ = new_A4786_ & new_A4785_;
  assign new_A4773_ = new_A4784_ & new_A4783_;
  assign new_A4774_ = new_A4789_ | new_A4788_;
  assign new_A4775_ = new_A4784_ & new_A4787_;
  assign new_A4776_ = new_A4759_ | new_A4792_;
  assign new_A4777_ = new_A4791_ | new_A4790_;
  assign new_A4778_ = new_A4794_ | new_A4793_;
  assign new_A4779_ = ~new_A4770_ & new_A4796_;
  assign new_A4780_ = ~new_A4772_ & new_A4784_;
  assign new_A4781_ = new_A4772_ & ~new_A4784_;
  assign new_A4782_ = new_A4758_ & ~new_A4759_;
  assign new_A4783_ = ~new_A4805_ | ~new_A4806_;
  assign new_A4784_ = new_A4798_ | new_A4800_;
  assign new_A4785_ = new_A4808_ | new_A4807_;
  assign new_A4786_ = new_A4802_ | new_A4801_;
  assign new_A4787_ = ~new_A4810_ | ~new_A4809_;
  assign new_A4788_ = ~new_A4811_ & new_A4812_;
  assign new_A4789_ = new_A4811_ & ~new_A4812_;
  assign new_A4790_ = ~new_A4758_ & new_A4759_;
  assign new_A4791_ = new_A4758_ & ~new_A4759_;
  assign new_A4792_ = ~new_A4774_ | new_A4784_;
  assign new_A4793_ = new_A4774_ & new_A4784_;
  assign new_A4794_ = ~new_A4774_ & ~new_A4784_;
  assign new_A4795_ = new_A4816_ | new_A4815_;
  assign new_A4796_ = new_A4762_ | new_A4795_;
  assign new_A4797_ = new_A4820_ | new_A4819_;
  assign new_A4798_ = ~new_A4762_ & new_A4797_;
  assign new_A4799_ = new_A4818_ | new_A4817_;
  assign new_A4800_ = new_A4762_ & new_A4799_;
  assign new_A4801_ = new_A4760_ & ~new_A4770_;
  assign new_A4802_ = ~new_A4760_ & new_A4770_;
  assign new_A4803_ = ~new_A4759_ | ~new_A4784_;
  assign new_A4804_ = new_A4770_ & new_A4803_;
  assign new_A4805_ = ~new_A4770_ & ~new_A4804_;
  assign new_A4806_ = new_A4770_ | new_A4803_;
  assign new_A4807_ = ~new_A4760_ & new_A4761_;
  assign new_A4808_ = new_A4760_ & ~new_A4761_;
  assign new_A4809_ = new_A4777_ | new_A4814_;
  assign new_A4810_ = ~new_A4777_ & ~new_A4813_;
  assign new_A4811_ = new_A4760_ | new_A4777_;
  assign new_A4812_ = new_A4760_ | new_A4761_;
  assign new_A4813_ = new_A4777_ & new_A4814_;
  assign new_A4814_ = ~new_A4759_ | ~new_A4784_;
  assign new_A4815_ = new_A4792_ & new_A4812_;
  assign new_A4816_ = ~new_A4792_ & ~new_A4812_;
  assign new_A4817_ = new_A4821_ | new_A4822_;
  assign new_A4818_ = ~new_A4763_ & new_A4777_;
  assign new_A4819_ = new_A4823_ | new_A4824_;
  assign new_A4820_ = new_A4763_ & new_A4777_;
  assign new_A4821_ = ~new_A4763_ & ~new_A4777_;
  assign new_A4822_ = new_A4763_ & ~new_A4777_;
  assign new_A4823_ = new_A4763_ & ~new_A4777_;
  assign new_A4824_ = ~new_A4763_ & new_A4777_;
  assign new_A4825_ = new_A5636_;
  assign new_A4826_ = new_A5706_;
  assign new_A4827_ = new_A5773_;
  assign new_A4828_ = new_A5840_;
  assign new_A4829_ = new_A5907_;
  assign new_A4830_ = new_A5974_;
  assign new_A4831_ = new_A4838_ & new_A4837_;
  assign new_A4832_ = new_A4840_ | new_A4839_;
  assign new_A4833_ = new_A4842_ | new_A4841_;
  assign new_A4834_ = new_A4844_ & new_A4843_;
  assign new_A4835_ = new_A4844_ & new_A4845_;
  assign new_A4836_ = new_A4837_ | new_A4846_;
  assign new_A4837_ = new_A4826_ | new_A4849_;
  assign new_A4838_ = new_A4848_ | new_A4847_;
  assign new_A4839_ = new_A4853_ & new_A4852_;
  assign new_A4840_ = new_A4851_ & new_A4850_;
  assign new_A4841_ = new_A4856_ | new_A4855_;
  assign new_A4842_ = new_A4851_ & new_A4854_;
  assign new_A4843_ = new_A4826_ | new_A4859_;
  assign new_A4844_ = new_A4858_ | new_A4857_;
  assign new_A4845_ = new_A4861_ | new_A4860_;
  assign new_A4846_ = ~new_A4837_ & new_A4863_;
  assign new_A4847_ = ~new_A4839_ & new_A4851_;
  assign new_A4848_ = new_A4839_ & ~new_A4851_;
  assign new_A4849_ = new_A4825_ & ~new_A4826_;
  assign new_A4850_ = ~new_A4872_ | ~new_A4873_;
  assign new_A4851_ = new_A4865_ | new_A4867_;
  assign new_A4852_ = new_A4875_ | new_A4874_;
  assign new_A4853_ = new_A4869_ | new_A4868_;
  assign new_A4854_ = ~new_A4877_ | ~new_A4876_;
  assign new_A4855_ = ~new_A4878_ & new_A4879_;
  assign new_A4856_ = new_A4878_ & ~new_A4879_;
  assign new_A4857_ = ~new_A4825_ & new_A4826_;
  assign new_A4858_ = new_A4825_ & ~new_A4826_;
  assign new_A4859_ = ~new_A4841_ | new_A4851_;
  assign new_A4860_ = new_A4841_ & new_A4851_;
  assign new_A4861_ = ~new_A4841_ & ~new_A4851_;
  assign new_A4862_ = new_A4883_ | new_A4882_;
  assign new_A4863_ = new_A4829_ | new_A4862_;
  assign new_A4864_ = new_A4887_ | new_A4886_;
  assign new_A4865_ = ~new_A4829_ & new_A4864_;
  assign new_A4866_ = new_A4885_ | new_A4884_;
  assign new_A4867_ = new_A4829_ & new_A4866_;
  assign new_A4868_ = new_A4827_ & ~new_A4837_;
  assign new_A4869_ = ~new_A4827_ & new_A4837_;
  assign new_A4870_ = ~new_A4826_ | ~new_A4851_;
  assign new_A4871_ = new_A4837_ & new_A4870_;
  assign new_A4872_ = ~new_A4837_ & ~new_A4871_;
  assign new_A4873_ = new_A4837_ | new_A4870_;
  assign new_A4874_ = ~new_A4827_ & new_A4828_;
  assign new_A4875_ = new_A4827_ & ~new_A4828_;
  assign new_A4876_ = new_A4844_ | new_A4881_;
  assign new_A4877_ = ~new_A4844_ & ~new_A4880_;
  assign new_A4878_ = new_A4827_ | new_A4844_;
  assign new_A4879_ = new_A4827_ | new_A4828_;
  assign new_A4880_ = new_A4844_ & new_A4881_;
  assign new_A4881_ = ~new_A4826_ | ~new_A4851_;
  assign new_A4882_ = new_A4859_ & new_A4879_;
  assign new_A4883_ = ~new_A4859_ & ~new_A4879_;
  assign new_A4884_ = new_A4888_ | new_A4889_;
  assign new_A4885_ = ~new_A4830_ & new_A4844_;
  assign new_A4886_ = new_A4890_ | new_A4891_;
  assign new_A4887_ = new_A4830_ & new_A4844_;
  assign new_A4888_ = ~new_A4830_ & ~new_A4844_;
  assign new_A4889_ = new_A4830_ & ~new_A4844_;
  assign new_A4890_ = new_A4830_ & ~new_A4844_;
  assign new_A4891_ = ~new_A4830_ & new_A4844_;
  assign new_A4892_ = new_A6041_;
  assign new_A4893_ = new_A6108_;
  assign new_A4894_ = new_A6175_;
  assign new_A4895_ = new_A6242_;
  assign new_A4896_ = new_A6309_;
  assign new_A4897_ = new_A6376_;
  assign new_A4898_ = new_A4905_ & new_A4904_;
  assign new_A4899_ = new_A4907_ | new_A4906_;
  assign new_A4900_ = new_A4909_ | new_A4908_;
  assign new_A4901_ = new_A4911_ & new_A4910_;
  assign new_A4902_ = new_A4911_ & new_A4912_;
  assign new_A4903_ = new_A4904_ | new_A4913_;
  assign new_A4904_ = new_A4893_ | new_A4916_;
  assign new_A4905_ = new_A4915_ | new_A4914_;
  assign new_A4906_ = new_A4920_ & new_A4919_;
  assign new_A4907_ = new_A4918_ & new_A4917_;
  assign new_A4908_ = new_A4923_ | new_A4922_;
  assign new_A4909_ = new_A4918_ & new_A4921_;
  assign new_A4910_ = new_A4893_ | new_A4926_;
  assign new_A4911_ = new_A4925_ | new_A4924_;
  assign new_A4912_ = new_A4928_ | new_A4927_;
  assign new_A4913_ = ~new_A4904_ & new_A4930_;
  assign new_A4914_ = ~new_A4906_ & new_A4918_;
  assign new_A4915_ = new_A4906_ & ~new_A4918_;
  assign new_A4916_ = new_A4892_ & ~new_A4893_;
  assign new_A4917_ = ~new_A4939_ | ~new_A4940_;
  assign new_A4918_ = new_A4932_ | new_A4934_;
  assign new_A4919_ = new_A4942_ | new_A4941_;
  assign new_A4920_ = new_A4936_ | new_A4935_;
  assign new_A4921_ = ~new_A4944_ | ~new_A4943_;
  assign new_A4922_ = ~new_A4945_ & new_A4946_;
  assign new_A4923_ = new_A4945_ & ~new_A4946_;
  assign new_A4924_ = ~new_A4892_ & new_A4893_;
  assign new_A4925_ = new_A4892_ & ~new_A4893_;
  assign new_A4926_ = ~new_A4908_ | new_A4918_;
  assign new_A4927_ = new_A4908_ & new_A4918_;
  assign new_A4928_ = ~new_A4908_ & ~new_A4918_;
  assign new_A4929_ = new_A4950_ | new_A4949_;
  assign new_A4930_ = new_A4896_ | new_A4929_;
  assign new_A4931_ = new_A4954_ | new_A4953_;
  assign new_A4932_ = ~new_A4896_ & new_A4931_;
  assign new_A4933_ = new_A4952_ | new_A4951_;
  assign new_A4934_ = new_A4896_ & new_A4933_;
  assign new_A4935_ = new_A4894_ & ~new_A4904_;
  assign new_A4936_ = ~new_A4894_ & new_A4904_;
  assign new_A4937_ = ~new_A4893_ | ~new_A4918_;
  assign new_A4938_ = new_A4904_ & new_A4937_;
  assign new_A4939_ = ~new_A4904_ & ~new_A4938_;
  assign new_A4940_ = new_A4904_ | new_A4937_;
  assign new_A4941_ = ~new_A4894_ & new_A4895_;
  assign new_A4942_ = new_A4894_ & ~new_A4895_;
  assign new_A4943_ = new_A4911_ | new_A4948_;
  assign new_A4944_ = ~new_A4911_ & ~new_A4947_;
  assign new_A4945_ = new_A4894_ | new_A4911_;
  assign new_A4946_ = new_A4894_ | new_A4895_;
  assign new_A4947_ = new_A4911_ & new_A4948_;
  assign new_A4948_ = ~new_A4893_ | ~new_A4918_;
  assign new_A4949_ = new_A4926_ & new_A4946_;
  assign new_A4950_ = ~new_A4926_ & ~new_A4946_;
  assign new_A4951_ = new_A4955_ | new_A4956_;
  assign new_A4952_ = ~new_A4897_ & new_A4911_;
  assign new_A4953_ = new_A4957_ | new_A4958_;
  assign new_A4954_ = new_A4897_ & new_A4911_;
  assign new_A4955_ = ~new_A4897_ & ~new_A4911_;
  assign new_A4956_ = new_A4897_ & ~new_A4911_;
  assign new_A4957_ = new_A4897_ & ~new_A4911_;
  assign new_A4958_ = ~new_A4897_ & new_A4911_;
  assign new_A4959_ = new_A6443_;
  assign new_A4960_ = new_A6510_;
  assign new_A4961_ = new_A6577_;
  assign new_A4962_ = new_A6644_;
  assign new_A4963_ = new_A6711_;
  assign new_A4964_ = new_A6778_;
  assign new_A4965_ = new_A4972_ & new_A4971_;
  assign new_A4966_ = new_A4974_ | new_A4973_;
  assign new_A4967_ = new_A4976_ | new_A4975_;
  assign new_A4968_ = new_A4978_ & new_A4977_;
  assign new_A4969_ = new_A4978_ & new_A4979_;
  assign new_A4970_ = new_A4971_ | new_A4980_;
  assign new_A4971_ = new_A4960_ | new_A4983_;
  assign new_A4972_ = new_A4982_ | new_A4981_;
  assign new_A4973_ = new_A4987_ & new_A4986_;
  assign new_A4974_ = new_A4985_ & new_A4984_;
  assign new_A4975_ = new_A4990_ | new_A4989_;
  assign new_A4976_ = new_A4985_ & new_A4988_;
  assign new_A4977_ = new_A4960_ | new_A4993_;
  assign new_A4978_ = new_A4992_ | new_A4991_;
  assign new_A4979_ = new_A4995_ | new_A4994_;
  assign new_A4980_ = ~new_A4971_ & new_A4997_;
  assign new_A4981_ = ~new_A4973_ & new_A4985_;
  assign new_A4982_ = new_A4973_ & ~new_A4985_;
  assign new_A4983_ = new_A4959_ & ~new_A4960_;
  assign new_A4984_ = ~new_A5006_ | ~new_A5007_;
  assign new_A4985_ = new_A4999_ | new_A5001_;
  assign new_A4986_ = new_A5009_ | new_A5008_;
  assign new_A4987_ = new_A5003_ | new_A5002_;
  assign new_A4988_ = ~new_A5011_ | ~new_A5010_;
  assign new_A4989_ = ~new_A5012_ & new_A5013_;
  assign new_A4990_ = new_A5012_ & ~new_A5013_;
  assign new_A4991_ = ~new_A4959_ & new_A4960_;
  assign new_A4992_ = new_A4959_ & ~new_A4960_;
  assign new_A4993_ = ~new_A4975_ | new_A4985_;
  assign new_A4994_ = new_A4975_ & new_A4985_;
  assign new_A4995_ = ~new_A4975_ & ~new_A4985_;
  assign new_A4996_ = new_A5017_ | new_A5016_;
  assign new_A4997_ = new_A4963_ | new_A4996_;
  assign new_A4998_ = new_A5021_ | new_A5020_;
  assign new_A4999_ = ~new_A4963_ & new_A4998_;
  assign new_A5000_ = new_A5019_ | new_A5018_;
  assign new_A5001_ = new_A4963_ & new_A5000_;
  assign new_A5002_ = new_A4961_ & ~new_A4971_;
  assign new_A5003_ = ~new_A4961_ & new_A4971_;
  assign new_A5004_ = ~new_A4960_ | ~new_A4985_;
  assign new_A5005_ = new_A4971_ & new_A5004_;
  assign new_A5006_ = ~new_A4971_ & ~new_A5005_;
  assign new_A5007_ = new_A4971_ | new_A5004_;
  assign new_A5008_ = ~new_A4961_ & new_A4962_;
  assign new_A5009_ = new_A4961_ & ~new_A4962_;
  assign new_A5010_ = new_A4978_ | new_A5015_;
  assign new_A5011_ = ~new_A4978_ & ~new_A5014_;
  assign new_A5012_ = new_A4961_ | new_A4978_;
  assign new_A5013_ = new_A4961_ | new_A4962_;
  assign new_A5014_ = new_A4978_ & new_A5015_;
  assign new_A5015_ = ~new_A4960_ | ~new_A4985_;
  assign new_A5016_ = new_A4993_ & new_A5013_;
  assign new_A5017_ = ~new_A4993_ & ~new_A5013_;
  assign new_A5018_ = new_A5022_ | new_A5023_;
  assign new_A5019_ = ~new_A4964_ & new_A4978_;
  assign new_A5020_ = new_A5024_ | new_A5025_;
  assign new_A5021_ = new_A4964_ & new_A4978_;
  assign new_A5022_ = ~new_A4964_ & ~new_A4978_;
  assign new_A5023_ = new_A4964_ & ~new_A4978_;
  assign new_A5024_ = new_A4964_ & ~new_A4978_;
  assign new_A5025_ = ~new_A4964_ & new_A4978_;
  assign new_A5026_ = new_A6845_;
  assign new_A5027_ = new_A6912_;
  assign new_A5028_ = new_A6979_;
  assign new_A5029_ = new_A7046_;
  assign new_A5030_ = new_A7113_;
  assign new_A5031_ = new_A7180_;
  assign new_A5032_ = new_A5039_ & new_A5038_;
  assign new_A5033_ = new_A5041_ | new_A5040_;
  assign new_A5034_ = new_A5043_ | new_A5042_;
  assign new_A5035_ = new_A5045_ & new_A5044_;
  assign new_A5036_ = new_A5045_ & new_A5046_;
  assign new_A5037_ = new_A5038_ | new_A5047_;
  assign new_A5038_ = new_A5027_ | new_A5050_;
  assign new_A5039_ = new_A5049_ | new_A5048_;
  assign new_A5040_ = new_A5054_ & new_A5053_;
  assign new_A5041_ = new_A5052_ & new_A5051_;
  assign new_A5042_ = new_A5057_ | new_A5056_;
  assign new_A5043_ = new_A5052_ & new_A5055_;
  assign new_A5044_ = new_A5027_ | new_A5060_;
  assign new_A5045_ = new_A5059_ | new_A5058_;
  assign new_A5046_ = new_A5062_ | new_A5061_;
  assign new_A5047_ = ~new_A5038_ & new_A5064_;
  assign new_A5048_ = ~new_A5040_ & new_A5052_;
  assign new_A5049_ = new_A5040_ & ~new_A5052_;
  assign new_A5050_ = new_A5026_ & ~new_A5027_;
  assign new_A5051_ = ~new_A5073_ | ~new_A5074_;
  assign new_A5052_ = new_A5066_ | new_A5068_;
  assign new_A5053_ = new_A5076_ | new_A5075_;
  assign new_A5054_ = new_A5070_ | new_A5069_;
  assign new_A5055_ = ~new_A5078_ | ~new_A5077_;
  assign new_A5056_ = ~new_A5079_ & new_A5080_;
  assign new_A5057_ = new_A5079_ & ~new_A5080_;
  assign new_A5058_ = ~new_A5026_ & new_A5027_;
  assign new_A5059_ = new_A5026_ & ~new_A5027_;
  assign new_A5060_ = ~new_A5042_ | new_A5052_;
  assign new_A5061_ = new_A5042_ & new_A5052_;
  assign new_A5062_ = ~new_A5042_ & ~new_A5052_;
  assign new_A5063_ = new_A5084_ | new_A5083_;
  assign new_A5064_ = new_A5030_ | new_A5063_;
  assign new_A5065_ = new_A5088_ | new_A5087_;
  assign new_A5066_ = ~new_A5030_ & new_A5065_;
  assign new_A5067_ = new_A5086_ | new_A5085_;
  assign new_A5068_ = new_A5030_ & new_A5067_;
  assign new_A5069_ = new_A5028_ & ~new_A5038_;
  assign new_A5070_ = ~new_A5028_ & new_A5038_;
  assign new_A5071_ = ~new_A5027_ | ~new_A5052_;
  assign new_A5072_ = new_A5038_ & new_A5071_;
  assign new_A5073_ = ~new_A5038_ & ~new_A5072_;
  assign new_A5074_ = new_A5038_ | new_A5071_;
  assign new_A5075_ = ~new_A5028_ & new_A5029_;
  assign new_A5076_ = new_A5028_ & ~new_A5029_;
  assign new_A5077_ = new_A5045_ | new_A5082_;
  assign new_A5078_ = ~new_A5045_ & ~new_A5081_;
  assign new_A5079_ = new_A5028_ | new_A5045_;
  assign new_A5080_ = new_A5028_ | new_A5029_;
  assign new_A5081_ = new_A5045_ & new_A5082_;
  assign new_A5082_ = ~new_A5027_ | ~new_A5052_;
  assign new_A5083_ = new_A5060_ & new_A5080_;
  assign new_A5084_ = ~new_A5060_ & ~new_A5080_;
  assign new_A5085_ = new_A5089_ | new_A5090_;
  assign new_A5086_ = ~new_A5031_ & new_A5045_;
  assign new_A5087_ = new_A5091_ | new_A5092_;
  assign new_A5088_ = new_A5031_ & new_A5045_;
  assign new_A5089_ = ~new_A5031_ & ~new_A5045_;
  assign new_A5090_ = new_A5031_ & ~new_A5045_;
  assign new_A5091_ = new_A5031_ & ~new_A5045_;
  assign new_A5092_ = ~new_A5031_ & new_A5045_;
  assign new_A5093_ = new_A7247_;
  assign new_A5094_ = new_A7314_;
  assign new_A5095_ = new_A7381_;
  assign new_A5096_ = new_A7448_;
  assign new_A5097_ = new_A7515_;
  assign new_A5098_ = new_A7582_;
  assign new_A5099_ = new_A5106_ & new_A5105_;
  assign new_A5100_ = new_A5108_ | new_A5107_;
  assign new_A5101_ = new_A5110_ | new_A5109_;
  assign new_A5102_ = new_A5112_ & new_A5111_;
  assign new_A5103_ = new_A5112_ & new_A5113_;
  assign new_A5104_ = new_A5105_ | new_A5114_;
  assign new_A5105_ = new_A5094_ | new_A5117_;
  assign new_A5106_ = new_A5116_ | new_A5115_;
  assign new_A5107_ = new_A5121_ & new_A5120_;
  assign new_A5108_ = new_A5119_ & new_A5118_;
  assign new_A5109_ = new_A5124_ | new_A5123_;
  assign new_A5110_ = new_A5119_ & new_A5122_;
  assign new_A5111_ = new_A5094_ | new_A5127_;
  assign new_A5112_ = new_A5126_ | new_A5125_;
  assign new_A5113_ = new_A5129_ | new_A5128_;
  assign new_A5114_ = ~new_A5105_ & new_A5131_;
  assign new_A5115_ = ~new_A5107_ & new_A5119_;
  assign new_A5116_ = new_A5107_ & ~new_A5119_;
  assign new_A5117_ = new_A5093_ & ~new_A5094_;
  assign new_A5118_ = ~new_A5140_ | ~new_A5141_;
  assign new_A5119_ = new_A5133_ | new_A5135_;
  assign new_A5120_ = new_A5143_ | new_A5142_;
  assign new_A5121_ = new_A5137_ | new_A5136_;
  assign new_A5122_ = ~new_A5145_ | ~new_A5144_;
  assign new_A5123_ = ~new_A5146_ & new_A5147_;
  assign new_A5124_ = new_A5146_ & ~new_A5147_;
  assign new_A5125_ = ~new_A5093_ & new_A5094_;
  assign new_A5126_ = new_A5093_ & ~new_A5094_;
  assign new_A5127_ = ~new_A5109_ | new_A5119_;
  assign new_A5128_ = new_A5109_ & new_A5119_;
  assign new_A5129_ = ~new_A5109_ & ~new_A5119_;
  assign new_A5130_ = new_A5151_ | new_A5150_;
  assign new_A5131_ = new_A5097_ | new_A5130_;
  assign new_A5132_ = new_A5155_ | new_A5154_;
  assign new_A5133_ = ~new_A5097_ & new_A5132_;
  assign new_A5134_ = new_A5153_ | new_A5152_;
  assign new_A5135_ = new_A5097_ & new_A5134_;
  assign new_A5136_ = new_A5095_ & ~new_A5105_;
  assign new_A5137_ = ~new_A5095_ & new_A5105_;
  assign new_A5138_ = ~new_A5094_ | ~new_A5119_;
  assign new_A5139_ = new_A5105_ & new_A5138_;
  assign new_A5140_ = ~new_A5105_ & ~new_A5139_;
  assign new_A5141_ = new_A5105_ | new_A5138_;
  assign new_A5142_ = ~new_A5095_ & new_A5096_;
  assign new_A5143_ = new_A5095_ & ~new_A5096_;
  assign new_A5144_ = new_A5112_ | new_A5149_;
  assign new_A5145_ = ~new_A5112_ & ~new_A5148_;
  assign new_A5146_ = new_A5095_ | new_A5112_;
  assign new_A5147_ = new_A5095_ | new_A5096_;
  assign new_A5148_ = new_A5112_ & new_A5149_;
  assign new_A5149_ = ~new_A5094_ | ~new_A5119_;
  assign new_A5150_ = new_A5127_ & new_A5147_;
  assign new_A5151_ = ~new_A5127_ & ~new_A5147_;
  assign new_A5152_ = new_A5156_ | new_A5157_;
  assign new_A5153_ = ~new_A5098_ & new_A5112_;
  assign new_A5154_ = new_A5158_ | new_A5159_;
  assign new_A5155_ = new_A5098_ & new_A5112_;
  assign new_A5156_ = ~new_A5098_ & ~new_A5112_;
  assign new_A5157_ = new_A5098_ & ~new_A5112_;
  assign new_A5158_ = new_A5098_ & ~new_A5112_;
  assign new_A5159_ = ~new_A5098_ & new_A5112_;
  assign new_A5160_ = new_A7649_;
  assign new_A5161_ = new_A7716_;
  assign new_A5162_ = new_A7783_;
  assign new_A5163_ = new_A7850_;
  assign new_A5164_ = new_A7917_;
  assign new_A5165_ = new_A7984_;
  assign new_A5166_ = new_A5173_ & new_A5172_;
  assign new_A5167_ = new_A5175_ | new_A5174_;
  assign new_A5168_ = new_A5177_ | new_A5176_;
  assign new_A5169_ = new_A5179_ & new_A5178_;
  assign new_A5170_ = new_A5179_ & new_A5180_;
  assign new_A5171_ = new_A5172_ | new_A5181_;
  assign new_A5172_ = new_A5161_ | new_A5184_;
  assign new_A5173_ = new_A5183_ | new_A5182_;
  assign new_A5174_ = new_A5188_ & new_A5187_;
  assign new_A5175_ = new_A5186_ & new_A5185_;
  assign new_A5176_ = new_A5191_ | new_A5190_;
  assign new_A5177_ = new_A5186_ & new_A5189_;
  assign new_A5178_ = new_A5161_ | new_A5194_;
  assign new_A5179_ = new_A5193_ | new_A5192_;
  assign new_A5180_ = new_A5196_ | new_A5195_;
  assign new_A5181_ = ~new_A5172_ & new_A5198_;
  assign new_A5182_ = ~new_A5174_ & new_A5186_;
  assign new_A5183_ = new_A5174_ & ~new_A5186_;
  assign new_A5184_ = new_A5160_ & ~new_A5161_;
  assign new_A5185_ = ~new_A5207_ | ~new_A5208_;
  assign new_A5186_ = new_A5200_ | new_A5202_;
  assign new_A5187_ = new_A5210_ | new_A5209_;
  assign new_A5188_ = new_A5204_ | new_A5203_;
  assign new_A5189_ = ~new_A5212_ | ~new_A5211_;
  assign new_A5190_ = ~new_A5213_ & new_A5214_;
  assign new_A5191_ = new_A5213_ & ~new_A5214_;
  assign new_A5192_ = ~new_A5160_ & new_A5161_;
  assign new_A5193_ = new_A5160_ & ~new_A5161_;
  assign new_A5194_ = ~new_A5176_ | new_A5186_;
  assign new_A5195_ = new_A5176_ & new_A5186_;
  assign new_A5196_ = ~new_A5176_ & ~new_A5186_;
  assign new_A5197_ = new_A5218_ | new_A5217_;
  assign new_A5198_ = new_A5164_ | new_A5197_;
  assign new_A5199_ = new_A5222_ | new_A5221_;
  assign new_A5200_ = ~new_A5164_ & new_A5199_;
  assign new_A5201_ = new_A5220_ | new_A5219_;
  assign new_A5202_ = new_A5164_ & new_A5201_;
  assign new_A5203_ = new_A5162_ & ~new_A5172_;
  assign new_A5204_ = ~new_A5162_ & new_A5172_;
  assign new_A5205_ = ~new_A5161_ | ~new_A5186_;
  assign new_A5206_ = new_A5172_ & new_A5205_;
  assign new_A5207_ = ~new_A5172_ & ~new_A5206_;
  assign new_A5208_ = new_A5172_ | new_A5205_;
  assign new_A5209_ = ~new_A5162_ & new_A5163_;
  assign new_A5210_ = new_A5162_ & ~new_A5163_;
  assign new_A5211_ = new_A5179_ | new_A5216_;
  assign new_A5212_ = ~new_A5179_ & ~new_A5215_;
  assign new_A5213_ = new_A5162_ | new_A5179_;
  assign new_A5214_ = new_A5162_ | new_A5163_;
  assign new_A5215_ = new_A5179_ & new_A5216_;
  assign new_A5216_ = ~new_A5161_ | ~new_A5186_;
  assign new_A5217_ = new_A5194_ & new_A5214_;
  assign new_A5218_ = ~new_A5194_ & ~new_A5214_;
  assign new_A5219_ = new_A5223_ | new_A5224_;
  assign new_A5220_ = ~new_A5165_ & new_A5179_;
  assign new_A5221_ = new_A5225_ | new_A5226_;
  assign new_A5222_ = new_A5165_ & new_A5179_;
  assign new_A5223_ = ~new_A5165_ & ~new_A5179_;
  assign new_A5224_ = new_A5165_ & ~new_A5179_;
  assign new_A5225_ = new_A5165_ & ~new_A5179_;
  assign new_A5226_ = ~new_A5165_ & new_A5179_;
  assign new_A5227_ = new_A5635_;
  assign new_A5228_ = new_A5707_;
  assign new_A5229_ = new_A5774_;
  assign new_A5230_ = new_A5841_;
  assign new_A5231_ = new_A5908_;
  assign new_A5232_ = new_A5975_;
  assign new_A5233_ = new_A5240_ & new_A5239_;
  assign new_A5234_ = new_A5242_ | new_A5241_;
  assign new_A5235_ = new_A5244_ | new_A5243_;
  assign new_A5236_ = new_A5246_ & new_A5245_;
  assign new_A5237_ = new_A5246_ & new_A5247_;
  assign new_A5238_ = new_A5239_ | new_A5248_;
  assign new_A5239_ = new_A5228_ | new_A5251_;
  assign new_A5240_ = new_A5250_ | new_A5249_;
  assign new_A5241_ = new_A5255_ & new_A5254_;
  assign new_A5242_ = new_A5253_ & new_A5252_;
  assign new_A5243_ = new_A5258_ | new_A5257_;
  assign new_A5244_ = new_A5253_ & new_A5256_;
  assign new_A5245_ = new_A5228_ | new_A5261_;
  assign new_A5246_ = new_A5260_ | new_A5259_;
  assign new_A5247_ = new_A5263_ | new_A5262_;
  assign new_A5248_ = ~new_A5239_ & new_A5265_;
  assign new_A5249_ = ~new_A5241_ & new_A5253_;
  assign new_A5250_ = new_A5241_ & ~new_A5253_;
  assign new_A5251_ = new_A5227_ & ~new_A5228_;
  assign new_A5252_ = ~new_A5274_ | ~new_A5275_;
  assign new_A5253_ = new_A5267_ | new_A5269_;
  assign new_A5254_ = new_A5277_ | new_A5276_;
  assign new_A5255_ = new_A5271_ | new_A5270_;
  assign new_A5256_ = ~new_A5279_ | ~new_A5278_;
  assign new_A5257_ = ~new_A5280_ & new_A5281_;
  assign new_A5258_ = new_A5280_ & ~new_A5281_;
  assign new_A5259_ = ~new_A5227_ & new_A5228_;
  assign new_A5260_ = new_A5227_ & ~new_A5228_;
  assign new_A5261_ = ~new_A5243_ | new_A5253_;
  assign new_A5262_ = new_A5243_ & new_A5253_;
  assign new_A5263_ = ~new_A5243_ & ~new_A5253_;
  assign new_A5264_ = new_A5285_ | new_A5284_;
  assign new_A5265_ = new_A5231_ | new_A5264_;
  assign new_A5266_ = new_A5289_ | new_A5288_;
  assign new_A5267_ = ~new_A5231_ & new_A5266_;
  assign new_A5268_ = new_A5287_ | new_A5286_;
  assign new_A5269_ = new_A5231_ & new_A5268_;
  assign new_A5270_ = new_A5229_ & ~new_A5239_;
  assign new_A5271_ = ~new_A5229_ & new_A5239_;
  assign new_A5272_ = ~new_A5228_ | ~new_A5253_;
  assign new_A5273_ = new_A5239_ & new_A5272_;
  assign new_A5274_ = ~new_A5239_ & ~new_A5273_;
  assign new_A5275_ = new_A5239_ | new_A5272_;
  assign new_A5276_ = ~new_A5229_ & new_A5230_;
  assign new_A5277_ = new_A5229_ & ~new_A5230_;
  assign new_A5278_ = new_A5246_ | new_A5283_;
  assign new_A5279_ = ~new_A5246_ & ~new_A5282_;
  assign new_A5280_ = new_A5229_ | new_A5246_;
  assign new_A5281_ = new_A5229_ | new_A5230_;
  assign new_A5282_ = new_A5246_ & new_A5283_;
  assign new_A5283_ = ~new_A5228_ | ~new_A5253_;
  assign new_A5284_ = new_A5261_ & new_A5281_;
  assign new_A5285_ = ~new_A5261_ & ~new_A5281_;
  assign new_A5286_ = new_A5290_ | new_A5291_;
  assign new_A5287_ = ~new_A5232_ & new_A5246_;
  assign new_A5288_ = new_A5292_ | new_A5293_;
  assign new_A5289_ = new_A5232_ & new_A5246_;
  assign new_A5290_ = ~new_A5232_ & ~new_A5246_;
  assign new_A5291_ = new_A5232_ & ~new_A5246_;
  assign new_A5292_ = new_A5232_ & ~new_A5246_;
  assign new_A5293_ = ~new_A5232_ & new_A5246_;
  assign new_A5294_ = new_A6042_;
  assign new_A5295_ = new_A6109_;
  assign new_A5296_ = new_A6176_;
  assign new_A5297_ = new_A6243_;
  assign new_A5298_ = new_A6310_;
  assign new_A5299_ = new_A6377_;
  assign new_A5300_ = new_A5307_ & new_A5306_;
  assign new_A5301_ = new_A5309_ | new_A5308_;
  assign new_A5302_ = new_A5311_ | new_A5310_;
  assign new_A5303_ = new_A5313_ & new_A5312_;
  assign new_A5304_ = new_A5313_ & new_A5314_;
  assign new_A5305_ = new_A5306_ | new_A5315_;
  assign new_A5306_ = new_A5295_ | new_A5318_;
  assign new_A5307_ = new_A5317_ | new_A5316_;
  assign new_A5308_ = new_A5322_ & new_A5321_;
  assign new_A5309_ = new_A5320_ & new_A5319_;
  assign new_A5310_ = new_A5325_ | new_A5324_;
  assign new_A5311_ = new_A5320_ & new_A5323_;
  assign new_A5312_ = new_A5295_ | new_A5328_;
  assign new_A5313_ = new_A5327_ | new_A5326_;
  assign new_A5314_ = new_A5330_ | new_A5329_;
  assign new_A5315_ = ~new_A5306_ & new_A5332_;
  assign new_A5316_ = ~new_A5308_ & new_A5320_;
  assign new_A5317_ = new_A5308_ & ~new_A5320_;
  assign new_A5318_ = new_A5294_ & ~new_A5295_;
  assign new_A5319_ = ~new_A5341_ | ~new_A5342_;
  assign new_A5320_ = new_A5334_ | new_A5336_;
  assign new_A5321_ = new_A5344_ | new_A5343_;
  assign new_A5322_ = new_A5338_ | new_A5337_;
  assign new_A5323_ = ~new_A5346_ | ~new_A5345_;
  assign new_A5324_ = ~new_A5347_ & new_A5348_;
  assign new_A5325_ = new_A5347_ & ~new_A5348_;
  assign new_A5326_ = ~new_A5294_ & new_A5295_;
  assign new_A5327_ = new_A5294_ & ~new_A5295_;
  assign new_A5328_ = ~new_A5310_ | new_A5320_;
  assign new_A5329_ = new_A5310_ & new_A5320_;
  assign new_A5330_ = ~new_A5310_ & ~new_A5320_;
  assign new_A5331_ = new_A5352_ | new_A5351_;
  assign new_A5332_ = new_A5298_ | new_A5331_;
  assign new_A5333_ = new_A5356_ | new_A5355_;
  assign new_A5334_ = ~new_A5298_ & new_A5333_;
  assign new_A5335_ = new_A5354_ | new_A5353_;
  assign new_A5336_ = new_A5298_ & new_A5335_;
  assign new_A5337_ = new_A5296_ & ~new_A5306_;
  assign new_A5338_ = ~new_A5296_ & new_A5306_;
  assign new_A5339_ = ~new_A5295_ | ~new_A5320_;
  assign new_A5340_ = new_A5306_ & new_A5339_;
  assign new_A5341_ = ~new_A5306_ & ~new_A5340_;
  assign new_A5342_ = new_A5306_ | new_A5339_;
  assign new_A5343_ = ~new_A5296_ & new_A5297_;
  assign new_A5344_ = new_A5296_ & ~new_A5297_;
  assign new_A5345_ = new_A5313_ | new_A5350_;
  assign new_A5346_ = ~new_A5313_ & ~new_A5349_;
  assign new_A5347_ = new_A5296_ | new_A5313_;
  assign new_A5348_ = new_A5296_ | new_A5297_;
  assign new_A5349_ = new_A5313_ & new_A5350_;
  assign new_A5350_ = ~new_A5295_ | ~new_A5320_;
  assign new_A5351_ = new_A5328_ & new_A5348_;
  assign new_A5352_ = ~new_A5328_ & ~new_A5348_;
  assign new_A5353_ = new_A5357_ | new_A5358_;
  assign new_A5354_ = ~new_A5299_ & new_A5313_;
  assign new_A5355_ = new_A5359_ | new_A5360_;
  assign new_A5356_ = new_A5299_ & new_A5313_;
  assign new_A5357_ = ~new_A5299_ & ~new_A5313_;
  assign new_A5358_ = new_A5299_ & ~new_A5313_;
  assign new_A5359_ = new_A5299_ & ~new_A5313_;
  assign new_A5360_ = ~new_A5299_ & new_A5313_;
  assign new_A5361_ = new_A6444_;
  assign new_A5362_ = new_A6511_;
  assign new_A5363_ = new_A6578_;
  assign new_A5364_ = new_A6645_;
  assign new_A5365_ = new_A6712_;
  assign new_A5366_ = new_A6779_;
  assign new_A5367_ = new_A5374_ & new_A5373_;
  assign new_A5368_ = new_A5376_ | new_A5375_;
  assign new_A5369_ = new_A5378_ | new_A5377_;
  assign new_A5370_ = new_A5380_ & new_A5379_;
  assign new_A5371_ = new_A5380_ & new_A5381_;
  assign new_A5372_ = new_A5373_ | new_A5382_;
  assign new_A5373_ = new_A5362_ | new_A5385_;
  assign new_A5374_ = new_A5384_ | new_A5383_;
  assign new_A5375_ = new_A5389_ & new_A5388_;
  assign new_A5376_ = new_A5387_ & new_A5386_;
  assign new_A5377_ = new_A5392_ | new_A5391_;
  assign new_A5378_ = new_A5387_ & new_A5390_;
  assign new_A5379_ = new_A5362_ | new_A5395_;
  assign new_A5380_ = new_A5394_ | new_A5393_;
  assign new_A5381_ = new_A5397_ | new_A5396_;
  assign new_A5382_ = ~new_A5373_ & new_A5399_;
  assign new_A5383_ = ~new_A5375_ & new_A5387_;
  assign new_A5384_ = new_A5375_ & ~new_A5387_;
  assign new_A5385_ = new_A5361_ & ~new_A5362_;
  assign new_A5386_ = ~new_A5408_ | ~new_A5409_;
  assign new_A5387_ = new_A5401_ | new_A5403_;
  assign new_A5388_ = new_A5411_ | new_A5410_;
  assign new_A5389_ = new_A5405_ | new_A5404_;
  assign new_A5390_ = ~new_A5413_ | ~new_A5412_;
  assign new_A5391_ = ~new_A5414_ & new_A5415_;
  assign new_A5392_ = new_A5414_ & ~new_A5415_;
  assign new_A5393_ = ~new_A5361_ & new_A5362_;
  assign new_A5394_ = new_A5361_ & ~new_A5362_;
  assign new_A5395_ = ~new_A5377_ | new_A5387_;
  assign new_A5396_ = new_A5377_ & new_A5387_;
  assign new_A5397_ = ~new_A5377_ & ~new_A5387_;
  assign new_A5398_ = new_A5419_ | new_A5418_;
  assign new_A5399_ = new_A5365_ | new_A5398_;
  assign new_A5400_ = new_A5423_ | new_A5422_;
  assign new_A5401_ = ~new_A5365_ & new_A5400_;
  assign new_A5402_ = new_A5421_ | new_A5420_;
  assign new_A5403_ = new_A5365_ & new_A5402_;
  assign new_A5404_ = new_A5363_ & ~new_A5373_;
  assign new_A5405_ = ~new_A5363_ & new_A5373_;
  assign new_A5406_ = ~new_A5362_ | ~new_A5387_;
  assign new_A5407_ = new_A5373_ & new_A5406_;
  assign new_A5408_ = ~new_A5373_ & ~new_A5407_;
  assign new_A5409_ = new_A5373_ | new_A5406_;
  assign new_A5410_ = ~new_A5363_ & new_A5364_;
  assign new_A5411_ = new_A5363_ & ~new_A5364_;
  assign new_A5412_ = new_A5380_ | new_A5417_;
  assign new_A5413_ = ~new_A5380_ & ~new_A5416_;
  assign new_A5414_ = new_A5363_ | new_A5380_;
  assign new_A5415_ = new_A5363_ | new_A5364_;
  assign new_A5416_ = new_A5380_ & new_A5417_;
  assign new_A5417_ = ~new_A5362_ | ~new_A5387_;
  assign new_A5418_ = new_A5395_ & new_A5415_;
  assign new_A5419_ = ~new_A5395_ & ~new_A5415_;
  assign new_A5420_ = new_A5424_ | new_A5425_;
  assign new_A5421_ = ~new_A5366_ & new_A5380_;
  assign new_A5422_ = new_A5426_ | new_A5427_;
  assign new_A5423_ = new_A5366_ & new_A5380_;
  assign new_A5424_ = ~new_A5366_ & ~new_A5380_;
  assign new_A5425_ = new_A5366_ & ~new_A5380_;
  assign new_A5426_ = new_A5366_ & ~new_A5380_;
  assign new_A5427_ = ~new_A5366_ & new_A5380_;
  assign new_A5428_ = new_A6846_;
  assign new_A5429_ = new_A6913_;
  assign new_A5430_ = new_A6980_;
  assign new_A5431_ = new_A7047_;
  assign new_A5432_ = new_A7114_;
  assign new_A5433_ = new_A7181_;
  assign new_A5434_ = new_A5441_ & new_A5440_;
  assign new_A5435_ = new_A5443_ | new_A5442_;
  assign new_A5436_ = new_A5445_ | new_A5444_;
  assign new_A5437_ = new_A5447_ & new_A5446_;
  assign new_A5438_ = new_A5447_ & new_A5448_;
  assign new_A5439_ = new_A5440_ | new_A5449_;
  assign new_A5440_ = new_A5429_ | new_A5452_;
  assign new_A5441_ = new_A5451_ | new_A5450_;
  assign new_A5442_ = new_A5456_ & new_A5455_;
  assign new_A5443_ = new_A5454_ & new_A5453_;
  assign new_A5444_ = new_A5459_ | new_A5458_;
  assign new_A5445_ = new_A5454_ & new_A5457_;
  assign new_A5446_ = new_A5429_ | new_A5462_;
  assign new_A5447_ = new_A5461_ | new_A5460_;
  assign new_A5448_ = new_A5464_ | new_A5463_;
  assign new_A5449_ = ~new_A5440_ & new_A5466_;
  assign new_A5450_ = ~new_A5442_ & new_A5454_;
  assign new_A5451_ = new_A5442_ & ~new_A5454_;
  assign new_A5452_ = new_A5428_ & ~new_A5429_;
  assign new_A5453_ = ~new_A5475_ | ~new_A5476_;
  assign new_A5454_ = new_A5468_ | new_A5470_;
  assign new_A5455_ = new_A5478_ | new_A5477_;
  assign new_A5456_ = new_A5472_ | new_A5471_;
  assign new_A5457_ = ~new_A5480_ | ~new_A5479_;
  assign new_A5458_ = ~new_A5481_ & new_A5482_;
  assign new_A5459_ = new_A5481_ & ~new_A5482_;
  assign new_A5460_ = ~new_A5428_ & new_A5429_;
  assign new_A5461_ = new_A5428_ & ~new_A5429_;
  assign new_A5462_ = ~new_A5444_ | new_A5454_;
  assign new_A5463_ = new_A5444_ & new_A5454_;
  assign new_A5464_ = ~new_A5444_ & ~new_A5454_;
  assign new_A5465_ = new_A5486_ | new_A5485_;
  assign new_A5466_ = new_A5432_ | new_A5465_;
  assign new_A5467_ = new_A5490_ | new_A5489_;
  assign new_A5468_ = ~new_A5432_ & new_A5467_;
  assign new_A5469_ = new_A5488_ | new_A5487_;
  assign new_A5470_ = new_A5432_ & new_A5469_;
  assign new_A5471_ = new_A5430_ & ~new_A5440_;
  assign new_A5472_ = ~new_A5430_ & new_A5440_;
  assign new_A5473_ = ~new_A5429_ | ~new_A5454_;
  assign new_A5474_ = new_A5440_ & new_A5473_;
  assign new_A5475_ = ~new_A5440_ & ~new_A5474_;
  assign new_A5476_ = new_A5440_ | new_A5473_;
  assign new_A5477_ = ~new_A5430_ & new_A5431_;
  assign new_A5478_ = new_A5430_ & ~new_A5431_;
  assign new_A5479_ = new_A5447_ | new_A5484_;
  assign new_A5480_ = ~new_A5447_ & ~new_A5483_;
  assign new_A5481_ = new_A5430_ | new_A5447_;
  assign new_A5482_ = new_A5430_ | new_A5431_;
  assign new_A5483_ = new_A5447_ & new_A5484_;
  assign new_A5484_ = ~new_A5429_ | ~new_A5454_;
  assign new_A5485_ = new_A5462_ & new_A5482_;
  assign new_A5486_ = ~new_A5462_ & ~new_A5482_;
  assign new_A5487_ = new_A5491_ | new_A5492_;
  assign new_A5488_ = ~new_A5433_ & new_A5447_;
  assign new_A5489_ = new_A5493_ | new_A5494_;
  assign new_A5490_ = new_A5433_ & new_A5447_;
  assign new_A5491_ = ~new_A5433_ & ~new_A5447_;
  assign new_A5492_ = new_A5433_ & ~new_A5447_;
  assign new_A5493_ = new_A5433_ & ~new_A5447_;
  assign new_A5494_ = ~new_A5433_ & new_A5447_;
  assign new_A5495_ = new_A7248_;
  assign new_A5496_ = new_A7315_;
  assign new_A5497_ = new_A7382_;
  assign new_A5498_ = new_A7449_;
  assign new_A5499_ = new_A7516_;
  assign new_A5500_ = new_A7583_;
  assign new_A5501_ = new_A5508_ & new_A5507_;
  assign new_A5502_ = new_A5510_ | new_A5509_;
  assign new_A5503_ = new_A5512_ | new_A5511_;
  assign new_A5504_ = new_A5514_ & new_A5513_;
  assign new_A5505_ = new_A5514_ & new_A5515_;
  assign new_A5506_ = new_A5507_ | new_A5516_;
  assign new_A5507_ = new_A5496_ | new_A5519_;
  assign new_A5508_ = new_A5518_ | new_A5517_;
  assign new_A5509_ = new_A5523_ & new_A5522_;
  assign new_A5510_ = new_A5521_ & new_A5520_;
  assign new_A5511_ = new_A5526_ | new_A5525_;
  assign new_A5512_ = new_A5521_ & new_A5524_;
  assign new_A5513_ = new_A5496_ | new_A5529_;
  assign new_A5514_ = new_A5528_ | new_A5527_;
  assign new_A5515_ = new_A5531_ | new_A5530_;
  assign new_A5516_ = ~new_A5507_ & new_A5533_;
  assign new_A5517_ = ~new_A5509_ & new_A5521_;
  assign new_A5518_ = new_A5509_ & ~new_A5521_;
  assign new_A5519_ = new_A5495_ & ~new_A5496_;
  assign new_A5520_ = ~new_A5542_ | ~new_A5543_;
  assign new_A5521_ = new_A5535_ | new_A5537_;
  assign new_A5522_ = new_A5545_ | new_A5544_;
  assign new_A5523_ = new_A5539_ | new_A5538_;
  assign new_A5524_ = ~new_A5547_ | ~new_A5546_;
  assign new_A5525_ = ~new_A5548_ & new_A5549_;
  assign new_A5526_ = new_A5548_ & ~new_A5549_;
  assign new_A5527_ = ~new_A5495_ & new_A5496_;
  assign new_A5528_ = new_A5495_ & ~new_A5496_;
  assign new_A5529_ = ~new_A5511_ | new_A5521_;
  assign new_A5530_ = new_A5511_ & new_A5521_;
  assign new_A5531_ = ~new_A5511_ & ~new_A5521_;
  assign new_A5532_ = new_A5553_ | new_A5552_;
  assign new_A5533_ = new_A5499_ | new_A5532_;
  assign new_A5534_ = new_A5557_ | new_A5556_;
  assign new_A5535_ = ~new_A5499_ & new_A5534_;
  assign new_A5536_ = new_A5555_ | new_A5554_;
  assign new_A5537_ = new_A5499_ & new_A5536_;
  assign new_A5538_ = new_A5497_ & ~new_A5507_;
  assign new_A5539_ = ~new_A5497_ & new_A5507_;
  assign new_A5540_ = ~new_A5496_ | ~new_A5521_;
  assign new_A5541_ = new_A5507_ & new_A5540_;
  assign new_A5542_ = ~new_A5507_ & ~new_A5541_;
  assign new_A5543_ = new_A5507_ | new_A5540_;
  assign new_A5544_ = ~new_A5497_ & new_A5498_;
  assign new_A5545_ = new_A5497_ & ~new_A5498_;
  assign new_A5546_ = new_A5514_ | new_A5551_;
  assign new_A5547_ = ~new_A5514_ & ~new_A5550_;
  assign new_A5548_ = new_A5497_ | new_A5514_;
  assign new_A5549_ = new_A5497_ | new_A5498_;
  assign new_A5550_ = new_A5514_ & new_A5551_;
  assign new_A5551_ = ~new_A5496_ | ~new_A5521_;
  assign new_A5552_ = new_A5529_ & new_A5549_;
  assign new_A5553_ = ~new_A5529_ & ~new_A5549_;
  assign new_A5554_ = new_A5558_ | new_A5559_;
  assign new_A5555_ = ~new_A5500_ & new_A5514_;
  assign new_A5556_ = new_A5560_ | new_A5561_;
  assign new_A5557_ = new_A5500_ & new_A5514_;
  assign new_A5558_ = ~new_A5500_ & ~new_A5514_;
  assign new_A5559_ = new_A5500_ & ~new_A5514_;
  assign new_A5560_ = new_A5500_ & ~new_A5514_;
  assign new_A5561_ = ~new_A5500_ & new_A5514_;
  assign new_A5562_ = new_A7650_;
  assign new_A5563_ = new_A7717_;
  assign new_A5564_ = new_A7784_;
  assign new_A5565_ = new_A7851_;
  assign new_A5566_ = new_A7918_;
  assign new_A5567_ = new_A7985_;
  assign new_A5568_ = new_A5575_ & new_A5574_;
  assign new_A5569_ = new_A5577_ | new_A5576_;
  assign new_A5570_ = new_A5579_ | new_A5578_;
  assign new_A5571_ = new_A5581_ & new_A5580_;
  assign new_A5572_ = new_A5581_ & new_A5582_;
  assign new_A5573_ = new_A5574_ | new_A5583_;
  assign new_A5574_ = new_A5563_ | new_A5586_;
  assign new_A5575_ = new_A5585_ | new_A5584_;
  assign new_A5576_ = new_A5590_ & new_A5589_;
  assign new_A5577_ = new_A5588_ & new_A5587_;
  assign new_A5578_ = new_A5593_ | new_A5592_;
  assign new_A5579_ = new_A5588_ & new_A5591_;
  assign new_A5580_ = new_A5563_ | new_A5596_;
  assign new_A5581_ = new_A5595_ | new_A5594_;
  assign new_A5582_ = new_A5598_ | new_A5597_;
  assign new_A5583_ = ~new_A5574_ & new_A5600_;
  assign new_A5584_ = ~new_A5576_ & new_A5588_;
  assign new_A5585_ = new_A5576_ & ~new_A5588_;
  assign new_A5586_ = new_A5562_ & ~new_A5563_;
  assign new_A5587_ = ~new_A5609_ | ~new_A5610_;
  assign new_A5588_ = new_A5602_ | new_A5604_;
  assign new_A5589_ = new_A5612_ | new_A5611_;
  assign new_A5590_ = new_A5606_ | new_A5605_;
  assign new_A5591_ = ~new_A5614_ | ~new_A5613_;
  assign new_A5592_ = ~new_A5615_ & new_A5616_;
  assign new_A5593_ = new_A5615_ & ~new_A5616_;
  assign new_A5594_ = ~new_A5562_ & new_A5563_;
  assign new_A5595_ = new_A5562_ & ~new_A5563_;
  assign new_A5596_ = ~new_A5578_ | new_A5588_;
  assign new_A5597_ = new_A5578_ & new_A5588_;
  assign new_A5598_ = ~new_A5578_ & ~new_A5588_;
  assign new_A5599_ = new_A5620_ | new_A5619_;
  assign new_A5600_ = new_A5566_ | new_A5599_;
  assign new_A5601_ = new_A5624_ | new_A5623_;
  assign new_A5602_ = ~new_A5566_ & new_A5601_;
  assign new_A5603_ = new_A5622_ | new_A5621_;
  assign new_A5604_ = new_A5566_ & new_A5603_;
  assign new_A5605_ = new_A5564_ & ~new_A5574_;
  assign new_A5606_ = ~new_A5564_ & new_A5574_;
  assign new_A5607_ = ~new_A5563_ | ~new_A5588_;
  assign new_A5608_ = new_A5574_ & new_A5607_;
  assign new_A5609_ = ~new_A5574_ & ~new_A5608_;
  assign new_A5610_ = new_A5574_ | new_A5607_;
  assign new_A5611_ = ~new_A5564_ & new_A5565_;
  assign new_A5612_ = new_A5564_ & ~new_A5565_;
  assign new_A5613_ = new_A5581_ | new_A5618_;
  assign new_A5614_ = ~new_A5581_ & ~new_A5617_;
  assign new_A5615_ = new_A5564_ | new_A5581_;
  assign new_A5616_ = new_A5564_ | new_A5565_;
  assign new_A5617_ = new_A5581_ & new_A5618_;
  assign new_A5618_ = ~new_A5563_ | ~new_A5588_;
  assign new_A5619_ = new_A5596_ & new_A5616_;
  assign new_A5620_ = ~new_A5596_ & ~new_A5616_;
  assign new_A5621_ = new_A5625_ | new_A5626_;
  assign new_A5622_ = ~new_A5567_ & new_A5581_;
  assign new_A5623_ = new_A5627_ | new_A5628_;
  assign new_A5624_ = new_A5567_ & new_A5581_;
  assign new_A5625_ = ~new_A5567_ & ~new_A5581_;
  assign new_A5626_ = new_A5567_ & ~new_A5581_;
  assign new_A5627_ = new_A5567_ & ~new_A5581_;
  assign new_A5628_ = ~new_A5567_ & new_A5581_;
  assign new_A3216_ = ~new_A3155_ & new_A3169_;
  assign new_A3215_ = new_A3155_ & ~new_A3169_;
  assign new_A3214_ = new_A3155_ & ~new_A3169_;
  assign new_A3213_ = ~new_A3155_ & ~new_A3169_;
  assign new_A3212_ = new_A3155_ & new_A3169_;
  assign new_A3211_ = new_A3215_ | new_A3216_;
  assign new_A3210_ = ~new_A3155_ & new_A3169_;
  assign new_A3209_ = new_A3213_ | new_A3214_;
  assign new_A3208_ = ~new_A3184_ & ~new_A3204_;
  assign new_A3207_ = new_A3184_ & new_A3204_;
  assign new_A3206_ = ~new_A3151_ | ~new_A3176_;
  assign new_A3205_ = new_A3169_ & new_A3206_;
  assign new_A3204_ = new_A3152_ | new_A3153_;
  assign new_A3203_ = new_A3152_ | new_A3169_;
  assign new_A3202_ = ~new_A3169_ & ~new_A3205_;
  assign new_A3201_ = new_A3169_ | new_A3206_;
  assign new_A3200_ = new_A3152_ & ~new_A3153_;
  assign new_A3199_ = ~new_A3152_ & new_A3153_;
  assign new_A3198_ = new_A3162_ | new_A3195_;
  assign new_A3197_ = ~new_A3162_ & ~new_A3196_;
  assign new_A3196_ = new_A3162_ & new_A3195_;
  assign new_A3195_ = ~new_A3151_ | ~new_A3176_;
  assign new_A3194_ = ~new_A3152_ & new_A3162_;
  assign new_A3193_ = new_A3152_ & ~new_A3162_;
  assign new_A3192_ = new_A3154_ & new_A3191_;
  assign new_A3191_ = new_A3210_ | new_A3209_;
  assign new_A3190_ = ~new_A3154_ & new_A3189_;
  assign new_A3189_ = new_A3212_ | new_A3211_;
  assign new_A3188_ = new_A3154_ | new_A3187_;
  assign new_A3187_ = new_A3208_ | new_A3207_;
  assign new_A3186_ = ~new_A3166_ & ~new_A3176_;
  assign new_A3185_ = new_A3166_ & new_A3176_;
  assign new_A3184_ = ~new_A3166_ | new_A3176_;
  assign new_A3183_ = new_A3150_ & ~new_A3151_;
  assign new_A3182_ = ~new_A3150_ & new_A3151_;
  assign new_A3181_ = new_A3203_ & ~new_A3204_;
  assign new_A3180_ = ~new_A3203_ & new_A3204_;
  assign new_A3179_ = ~new_A3202_ | ~new_A3201_;
  assign new_A3178_ = new_A3194_ | new_A3193_;
  assign new_A3177_ = new_A3200_ | new_A3199_;
  assign new_A3176_ = new_A3190_ | new_A3192_;
  assign new_A3175_ = ~new_A3197_ | ~new_A3198_;
  assign new_A3174_ = new_A3150_ & ~new_A3151_;
  assign new_A3173_ = new_A3164_ & ~new_A3176_;
  assign new_A3172_ = ~new_A3164_ & new_A3176_;
  assign new_A3171_ = ~new_A3162_ & new_A3188_;
  assign new_A3170_ = new_A3186_ | new_A3185_;
  assign new_A3169_ = new_A3183_ | new_A3182_;
  assign new_A3168_ = new_A3151_ | new_A3184_;
  assign new_A3167_ = new_A3176_ & new_A3179_;
  assign new_A3166_ = new_A3181_ | new_A3180_;
  assign new_A3165_ = new_A3176_ & new_A3175_;
  assign new_A3164_ = new_A3178_ & new_A3177_;
  assign new_A3163_ = new_A3173_ | new_A3172_;
  assign new_A3162_ = new_A3151_ | new_A3174_;
  assign A3161 = new_A3162_ | new_A3171_;
  assign A3160 = new_A3169_ & new_A3170_;
  assign A3159 = new_A3169_ & new_A3168_;
  assign A3158 = new_A3167_ | new_A3166_;
  assign A3157 = new_A3165_ | new_A3164_;
  assign A3156 = new_A3163_ & new_A3162_;
  assign new_A3155_ = new_A5573_;
  assign new_A3154_ = new_A5506_;
  assign new_A3153_ = new_A5439_;
  assign new_A3152_ = new_A5372_;
  assign new_A3151_ = new_A5305_;
  assign new_A3150_ = new_A5238_;
  assign new_A3149_ = ~new_A3088_ & new_A3102_;
  assign new_A3148_ = new_A3088_ & ~new_A3102_;
  assign new_A3147_ = new_A3088_ & ~new_A3102_;
  assign new_A3146_ = ~new_A3088_ & ~new_A3102_;
  assign new_A3145_ = new_A3088_ & new_A3102_;
  assign new_A3144_ = new_A3148_ | new_A3149_;
  assign new_A3143_ = ~new_A3088_ & new_A3102_;
  assign new_A3142_ = new_A3146_ | new_A3147_;
  assign new_A3141_ = ~new_A3117_ & ~new_A3137_;
  assign new_A3140_ = new_A3117_ & new_A3137_;
  assign new_A3139_ = ~new_A3084_ | ~new_A3109_;
  assign new_A3138_ = new_A3102_ & new_A3139_;
  assign new_A3137_ = new_A3085_ | new_A3086_;
  assign new_A3136_ = new_A3085_ | new_A3102_;
  assign new_A3135_ = ~new_A3102_ & ~new_A3138_;
  assign new_A3134_ = new_A3102_ | new_A3139_;
  assign new_A3133_ = new_A3085_ & ~new_A3086_;
  assign new_A3132_ = ~new_A3085_ & new_A3086_;
  assign new_A3131_ = new_A3095_ | new_A3128_;
  assign new_A3130_ = ~new_A3095_ & ~new_A3129_;
  assign new_A3129_ = new_A3095_ & new_A3128_;
  assign new_A3128_ = ~new_A3084_ | ~new_A3109_;
  assign new_A3127_ = ~new_A3085_ & new_A3095_;
  assign new_A3126_ = new_A3085_ & ~new_A3095_;
  assign new_A3125_ = new_A3087_ & new_A3124_;
  assign new_A3124_ = new_A3143_ | new_A3142_;
  assign new_A3123_ = ~new_A3087_ & new_A3122_;
  assign new_A3122_ = new_A3145_ | new_A3144_;
  assign new_A3121_ = new_A3087_ | new_A3120_;
  assign new_A3120_ = new_A3141_ | new_A3140_;
  assign new_A3119_ = ~new_A3099_ & ~new_A3109_;
  assign new_A3118_ = new_A3099_ & new_A3109_;
  assign new_A3117_ = ~new_A3099_ | new_A3109_;
  assign new_A3116_ = new_A3083_ & ~new_A3084_;
  assign new_A3115_ = ~new_A3083_ & new_A3084_;
  assign new_A3114_ = new_A3136_ & ~new_A3137_;
  assign new_A3113_ = ~new_A3136_ & new_A3137_;
  assign new_A3112_ = ~new_A3135_ | ~new_A3134_;
  assign new_A3111_ = new_A3127_ | new_A3126_;
  assign new_A3110_ = new_A3133_ | new_A3132_;
  assign new_A3109_ = new_A3123_ | new_A3125_;
  assign new_A3108_ = ~new_A3130_ | ~new_A3131_;
  assign new_A3107_ = new_A3083_ & ~new_A3084_;
  assign new_A3106_ = new_A3097_ & ~new_A3109_;
  assign new_A3105_ = ~new_A3097_ & new_A3109_;
  assign new_A3104_ = ~new_A3095_ & new_A3121_;
  assign new_A3103_ = new_A3119_ | new_A3118_;
  assign new_A3102_ = new_A3116_ | new_A3115_;
  assign new_A3101_ = new_A3084_ | new_A3117_;
  assign new_A3100_ = new_A3109_ & new_A3112_;
  assign new_A3099_ = new_A3114_ | new_A3113_;
  assign new_A3098_ = new_A3109_ & new_A3108_;
  assign new_A3097_ = new_A3111_ & new_A3110_;
  assign new_A3096_ = new_A3106_ | new_A3105_;
  assign new_A3095_ = new_A3084_ | new_A3107_;
  assign A3094 = new_A3095_ | new_A3104_;
  assign A3093 = new_A3102_ & new_A3103_;
  assign A3092 = new_A3102_ & new_A3101_;
  assign A3091 = new_A3100_ | new_A3099_;
  assign A3090 = new_A3098_ | new_A3097_;
  assign A3089 = new_A3096_ & new_A3095_;
  assign new_A3088_ = new_A5171_;
  assign new_A3087_ = new_A5104_;
  assign new_A3086_ = new_A5037_;
  assign new_A3085_ = new_A4970_;
  assign new_A3084_ = new_A4903_;
  assign new_A3083_ = new_A4836_;
  assign new_A3082_ = ~new_A3021_ & new_A3035_;
  assign new_A3081_ = new_A3021_ & ~new_A3035_;
  assign new_A3080_ = new_A3021_ & ~new_A3035_;
  assign new_A3079_ = ~new_A3021_ & ~new_A3035_;
  assign new_A3078_ = new_A3021_ & new_A3035_;
  assign new_A3077_ = new_A3081_ | new_A3082_;
  assign new_A3076_ = ~new_A3021_ & new_A3035_;
  assign new_A3075_ = new_A3079_ | new_A3080_;
  assign new_A3074_ = ~new_A3050_ & ~new_A3070_;
  assign new_A3073_ = new_A3050_ & new_A3070_;
  assign new_A3072_ = ~new_A3017_ | ~new_A3042_;
  assign new_A3071_ = new_A3035_ & new_A3072_;
  assign new_A3070_ = new_A3018_ | new_A3019_;
  assign new_A3069_ = new_A3018_ | new_A3035_;
  assign new_A3068_ = ~new_A3035_ & ~new_A3071_;
  assign new_A3067_ = new_A3035_ | new_A3072_;
  assign new_A3066_ = new_A3018_ & ~new_A3019_;
  assign new_A3065_ = ~new_A3018_ & new_A3019_;
  assign new_A3064_ = new_A3028_ | new_A3061_;
  assign new_A3063_ = ~new_A3028_ & ~new_A3062_;
  assign new_A3062_ = new_A3028_ & new_A3061_;
  assign new_A3061_ = ~new_A3017_ | ~new_A3042_;
  assign new_A3060_ = ~new_A3018_ & new_A3028_;
  assign new_A3059_ = new_A3018_ & ~new_A3028_;
  assign new_A3058_ = new_A3020_ & new_A3057_;
  assign new_A3057_ = new_A3076_ | new_A3075_;
  assign new_A3056_ = ~new_A3020_ & new_A3055_;
  assign new_A3055_ = new_A3078_ | new_A3077_;
  assign new_A3054_ = new_A3020_ | new_A3053_;
  assign new_A3053_ = new_A3074_ | new_A3073_;
  assign new_A3052_ = ~new_A3032_ & ~new_A3042_;
  assign new_A3051_ = new_A3032_ & new_A3042_;
  assign new_A3050_ = ~new_A3032_ | new_A3042_;
  assign new_A3049_ = new_A3016_ & ~new_A3017_;
  assign new_A3048_ = ~new_A3016_ & new_A3017_;
  assign new_A3047_ = new_A3069_ & ~new_A3070_;
  assign new_A3046_ = ~new_A3069_ & new_A3070_;
  assign new_A3045_ = ~new_A3068_ | ~new_A3067_;
  assign new_A3044_ = new_A3060_ | new_A3059_;
  assign new_A3043_ = new_A3066_ | new_A3065_;
  assign new_A3042_ = new_A3056_ | new_A3058_;
  assign new_A3041_ = ~new_A3063_ | ~new_A3064_;
  assign new_A3040_ = new_A3016_ & ~new_A3017_;
  assign new_A3039_ = new_A3030_ & ~new_A3042_;
  assign new_A3038_ = ~new_A3030_ & new_A3042_;
  assign new_A3037_ = ~new_A3028_ & new_A3054_;
  assign new_A3036_ = new_A3052_ | new_A3051_;
  assign new_A3035_ = new_A3049_ | new_A3048_;
  assign new_A3034_ = new_A3017_ | new_A3050_;
  assign new_A3033_ = new_A3042_ & new_A3045_;
  assign new_A3032_ = new_A3047_ | new_A3046_;
  assign new_A3031_ = new_A3042_ & new_A3041_;
  assign new_A3030_ = new_A3044_ & new_A3043_;
  assign new_A3029_ = new_A3039_ | new_A3038_;
  assign new_A3028_ = new_A3017_ | new_A3040_;
  assign A3027 = new_A3028_ | new_A3037_;
  assign A3026 = new_A3035_ & new_A3036_;
  assign A3025 = new_A3035_ & new_A3034_;
  assign A3024 = new_A3033_ | new_A3032_;
  assign A3023 = new_A3031_ | new_A3030_;
  assign A3022 = new_A3029_ & new_A3028_;
  assign new_A3021_ = new_A4769_;
  assign new_A3020_ = new_A4702_;
  assign new_A3019_ = new_A4635_;
  assign new_A3018_ = new_A4568_;
  assign new_A3017_ = new_A4501_;
  assign new_A3016_ = new_A4434_;
  assign new_A3015_ = ~new_A2954_ & new_A2968_;
  assign new_A3014_ = new_A2954_ & ~new_A2968_;
  assign new_A3013_ = new_A2954_ & ~new_A2968_;
  assign new_A3012_ = ~new_A2954_ & ~new_A2968_;
  assign new_A3011_ = new_A2954_ & new_A2968_;
  assign new_A3010_ = new_A3014_ | new_A3015_;
  assign new_A3009_ = ~new_A2954_ & new_A2968_;
  assign new_A3008_ = new_A3012_ | new_A3013_;
  assign new_A3007_ = ~new_A2983_ & ~new_A3003_;
  assign new_A3006_ = new_A2983_ & new_A3003_;
  assign new_A3005_ = ~new_A2950_ | ~new_A2975_;
  assign new_A3004_ = new_A2968_ & new_A3005_;
  assign new_A3003_ = new_A2951_ | new_A2952_;
  assign new_A3002_ = new_A2951_ | new_A2968_;
  assign new_A3001_ = ~new_A2968_ & ~new_A3004_;
  assign new_A3000_ = new_A2968_ | new_A3005_;
  assign new_A2999_ = new_A2951_ & ~new_A2952_;
  assign new_A2998_ = ~new_A2951_ & new_A2952_;
  assign new_A2997_ = new_A2961_ | new_A2994_;
  assign new_A2996_ = ~new_A2961_ & ~new_A2995_;
  assign new_A2995_ = new_A2961_ & new_A2994_;
  assign new_A2994_ = ~new_A2950_ | ~new_A2975_;
  assign new_A2993_ = ~new_A2951_ & new_A2961_;
  assign new_A2992_ = new_A2951_ & ~new_A2961_;
  assign new_A2991_ = new_A2953_ & new_A2990_;
  assign new_A2990_ = new_A3009_ | new_A3008_;
  assign new_A2989_ = ~new_A2953_ & new_A2988_;
  assign new_A2988_ = new_A3011_ | new_A3010_;
  assign new_A2987_ = new_A2953_ | new_A2986_;
  assign new_A2986_ = new_A3007_ | new_A3006_;
  assign new_A2985_ = ~new_A2965_ & ~new_A2975_;
  assign new_A2984_ = new_A2965_ & new_A2975_;
  assign new_A2983_ = ~new_A2965_ | new_A2975_;
  assign new_A2982_ = new_A2949_ & ~new_A2950_;
  assign new_A2981_ = ~new_A2949_ & new_A2950_;
  assign new_A2980_ = new_A3002_ & ~new_A3003_;
  assign new_A2979_ = ~new_A3002_ & new_A3003_;
  assign new_A2978_ = ~new_A3001_ | ~new_A3000_;
  assign new_A2977_ = new_A2993_ | new_A2992_;
  assign new_A2976_ = new_A2999_ | new_A2998_;
  assign new_A2975_ = new_A2989_ | new_A2991_;
  assign new_A2974_ = ~new_A2996_ | ~new_A2997_;
  assign new_A2973_ = new_A2949_ & ~new_A2950_;
  assign new_A2972_ = new_A2963_ & ~new_A2975_;
  assign new_A2971_ = ~new_A2963_ & new_A2975_;
  assign new_A2970_ = ~new_A2961_ & new_A2987_;
  assign new_A2969_ = new_A2985_ | new_A2984_;
  assign new_A2968_ = new_A2982_ | new_A2981_;
  assign new_A2967_ = new_A2950_ | new_A2983_;
  assign new_A2966_ = new_A2975_ & new_A2978_;
  assign new_A2965_ = new_A2980_ | new_A2979_;
  assign new_A2964_ = new_A2975_ & new_A2974_;
  assign new_A2963_ = new_A2977_ & new_A2976_;
  assign new_A2962_ = new_A2972_ | new_A2971_;
  assign new_A2961_ = new_A2950_ | new_A2973_;
  assign A2960 = new_A2961_ | new_A2970_;
  assign A2959 = new_A2968_ & new_A2969_;
  assign A2958 = new_A2968_ & new_A2967_;
  assign A2957 = new_A2966_ | new_A2965_;
  assign A2956 = new_A2964_ | new_A2963_;
  assign A2955 = new_A2962_ & new_A2961_;
  assign new_A2954_ = new_A4367_;
  assign new_A2953_ = new_A4300_;
  assign new_A2952_ = new_A4233_;
  assign new_A2951_ = new_A4166_;
  assign new_A2950_ = new_A4099_;
  assign new_A2949_ = new_A4032_;
  assign new_A2948_ = ~new_A2887_ & new_A2901_;
  assign new_A2947_ = new_A2887_ & ~new_A2901_;
  assign new_A2946_ = new_A2887_ & ~new_A2901_;
  assign new_A2945_ = ~new_A2887_ & ~new_A2901_;
  assign new_A2944_ = new_A2887_ & new_A2901_;
  assign new_A2943_ = new_A2947_ | new_A2948_;
  assign new_A2942_ = ~new_A2887_ & new_A2901_;
  assign new_A2941_ = new_A2945_ | new_A2946_;
  assign new_A2940_ = ~new_A2916_ & ~new_A2936_;
  assign new_A2939_ = new_A2916_ & new_A2936_;
  assign new_A2938_ = ~new_A2883_ | ~new_A2908_;
  assign new_A2937_ = new_A2901_ & new_A2938_;
  assign new_A2936_ = new_A2884_ | new_A2885_;
  assign new_A2935_ = new_A2884_ | new_A2901_;
  assign new_A2934_ = ~new_A2901_ & ~new_A2937_;
  assign new_A2933_ = new_A2901_ | new_A2938_;
  assign new_A2932_ = new_A2884_ & ~new_A2885_;
  assign new_A2931_ = ~new_A2884_ & new_A2885_;
  assign new_A2930_ = new_A2894_ | new_A2927_;
  assign new_A2929_ = ~new_A2894_ & ~new_A2928_;
  assign new_A2928_ = new_A2894_ & new_A2927_;
  assign new_A2927_ = ~new_A2883_ | ~new_A2908_;
  assign new_A2926_ = ~new_A2884_ & new_A2894_;
  assign new_A2925_ = new_A2884_ & ~new_A2894_;
  assign new_A2924_ = new_A2886_ & new_A2923_;
  assign new_A2923_ = new_A2942_ | new_A2941_;
  assign new_A2922_ = ~new_A2886_ & new_A2921_;
  assign new_A2921_ = new_A2944_ | new_A2943_;
  assign new_A2920_ = new_A2886_ | new_A2919_;
  assign new_A2919_ = new_A2940_ | new_A2939_;
  assign new_A2918_ = ~new_A2898_ & ~new_A2908_;
  assign new_A2917_ = new_A2898_ & new_A2908_;
  assign new_A2916_ = ~new_A2898_ | new_A2908_;
  assign new_A2915_ = new_A2882_ & ~new_A2883_;
  assign new_A2914_ = ~new_A2882_ & new_A2883_;
  assign new_A2913_ = new_A2935_ & ~new_A2936_;
  assign new_A2912_ = ~new_A2935_ & new_A2936_;
  assign new_A2911_ = ~new_A2934_ | ~new_A2933_;
  assign new_A2910_ = new_A2926_ | new_A2925_;
  assign new_A2909_ = new_A2932_ | new_A2931_;
  assign new_A2908_ = new_A2922_ | new_A2924_;
  assign new_A2907_ = ~new_A2929_ | ~new_A2930_;
  assign new_A2906_ = new_A2882_ & ~new_A2883_;
  assign new_A2905_ = new_A2896_ & ~new_A2908_;
  assign new_A2904_ = ~new_A2896_ & new_A2908_;
  assign new_A2903_ = ~new_A2894_ & new_A2920_;
  assign new_A2902_ = new_A2918_ | new_A2917_;
  assign new_A2901_ = new_A2915_ | new_A2914_;
  assign new_A2900_ = new_A2883_ | new_A2916_;
  assign new_A2899_ = new_A2908_ & new_A2911_;
  assign new_A2898_ = new_A2913_ | new_A2912_;
  assign new_A2897_ = new_A2908_ & new_A2907_;
  assign new_A2896_ = new_A2910_ & new_A2909_;
  assign new_A2895_ = new_A2905_ | new_A2904_;
  assign new_A2894_ = new_A2883_ | new_A2906_;
  assign A2893 = new_A2894_ | new_A2903_;
  assign A2892 = new_A2901_ & new_A2902_;
  assign A2891 = new_A2901_ & new_A2900_;
  assign A2890 = new_A2899_ | new_A2898_;
  assign A2889 = new_A2897_ | new_A2896_;
  assign A2888 = new_A2895_ & new_A2894_;
  assign new_A2887_ = new_A3965_;
  assign new_A2886_ = new_A3898_;
  assign new_A2885_ = new_A3831_;
  assign new_A2884_ = new_A3764_;
  assign new_A2883_ = new_A3697_;
  assign new_A2882_ = new_A3630_;
  assign new_A2881_ = ~new_A2820_ & new_A2834_;
  assign new_A2880_ = new_A2820_ & ~new_A2834_;
  assign new_A2879_ = new_A2820_ & ~new_A2834_;
  assign new_A2878_ = ~new_A2820_ & ~new_A2834_;
  assign new_A2877_ = new_A2820_ & new_A2834_;
  assign new_A2876_ = new_A2880_ | new_A2881_;
  assign new_A2875_ = ~new_A2820_ & new_A2834_;
  assign new_A2874_ = new_A2878_ | new_A2879_;
  assign new_A2873_ = ~new_A2849_ & ~new_A2869_;
  assign new_A2872_ = new_A2849_ & new_A2869_;
  assign new_A2871_ = ~new_A2816_ | ~new_A2841_;
  assign new_A2870_ = new_A2834_ & new_A2871_;
  assign new_A2869_ = new_A2817_ | new_A2818_;
  assign new_A2868_ = new_A2817_ | new_A2834_;
  assign new_A2867_ = ~new_A2834_ & ~new_A2870_;
  assign new_A2866_ = new_A2834_ | new_A2871_;
  assign new_A2865_ = new_A2817_ & ~new_A2818_;
  assign new_A2864_ = ~new_A2817_ & new_A2818_;
  assign new_A2863_ = new_A2827_ | new_A2860_;
  assign new_A2862_ = ~new_A2827_ & ~new_A2861_;
  assign new_A2861_ = new_A2827_ & new_A2860_;
  assign new_A2860_ = ~new_A2816_ | ~new_A2841_;
  assign new_A2859_ = ~new_A2817_ & new_A2827_;
  assign new_A2858_ = new_A2817_ & ~new_A2827_;
  assign new_A2857_ = new_A2819_ & new_A2856_;
  assign new_A2856_ = new_A2875_ | new_A2874_;
  assign new_A2855_ = ~new_A2819_ & new_A2854_;
  assign new_A2854_ = new_A2877_ | new_A2876_;
  assign new_A2853_ = new_A2819_ | new_A2852_;
  assign new_A2852_ = new_A2873_ | new_A2872_;
  assign new_A2851_ = ~new_A2831_ & ~new_A2841_;
  assign new_A2850_ = new_A2831_ & new_A2841_;
  assign new_A2849_ = ~new_A2831_ | new_A2841_;
  assign new_A2848_ = new_A2815_ & ~new_A2816_;
  assign new_A2847_ = ~new_A2815_ & new_A2816_;
  assign new_A2846_ = new_A2868_ & ~new_A2869_;
  assign new_A2845_ = ~new_A2868_ & new_A2869_;
  assign new_A2844_ = ~new_A2867_ | ~new_A2866_;
  assign new_A2843_ = new_A2859_ | new_A2858_;
  assign new_A2842_ = new_A2865_ | new_A2864_;
  assign new_A2841_ = new_A2855_ | new_A2857_;
  assign new_A2840_ = ~new_A2862_ | ~new_A2863_;
  assign new_A2839_ = new_A2815_ & ~new_A2816_;
  assign new_A2838_ = new_A2829_ & ~new_A2841_;
  assign new_A2837_ = ~new_A2829_ & new_A2841_;
  assign new_A2836_ = ~new_A2827_ & new_A2853_;
  assign new_A2835_ = new_A2851_ | new_A2850_;
  assign new_A2834_ = new_A2848_ | new_A2847_;
  assign new_A2833_ = new_A2816_ | new_A2849_;
  assign new_A2832_ = new_A2841_ & new_A2844_;
  assign new_A2831_ = new_A2846_ | new_A2845_;
  assign new_A2830_ = new_A2841_ & new_A2840_;
  assign new_A2829_ = new_A2843_ & new_A2842_;
  assign new_A2828_ = new_A2838_ | new_A2837_;
  assign new_A2827_ = new_A2816_ | new_A2839_;
  assign A2826 = new_A2827_ | new_A2836_;
  assign A2825 = new_A2834_ & new_A2835_;
  assign A2824 = new_A2834_ & new_A2833_;
  assign A2823 = new_A2832_ | new_A2831_;
  assign A2822 = new_A2830_ | new_A2829_;
  assign A2821 = new_A2828_ & new_A2827_;
  assign new_A2820_ = new_A3563_;
  assign new_A2819_ = new_A3496_;
  assign new_A2818_ = new_A3429_;
  assign new_A2817_ = new_A3362_;
  assign new_A2816_ = new_A3295_;
  assign new_A2815_ = new_A3223_;
  assign new_A2814_ = ~new_A2753_ & new_A2767_;
  assign new_A2813_ = new_A2753_ & ~new_A2767_;
  assign new_A2812_ = new_A2753_ & ~new_A2767_;
  assign new_A2811_ = ~new_A2753_ & ~new_A2767_;
  assign new_A2810_ = new_A2753_ & new_A2767_;
  assign new_A2809_ = new_A2813_ | new_A2814_;
  assign new_A2808_ = ~new_A2753_ & new_A2767_;
  assign new_A2807_ = new_A2811_ | new_A2812_;
  assign new_A2806_ = ~new_A2782_ & ~new_A2802_;
  assign new_A2805_ = new_A2782_ & new_A2802_;
  assign new_A2804_ = ~new_A2749_ | ~new_A2774_;
  assign new_A2803_ = new_A2767_ & new_A2804_;
  assign new_A2802_ = new_A2750_ | new_A2751_;
  assign new_A2801_ = new_A2750_ | new_A2767_;
  assign new_A2800_ = ~new_A2767_ & ~new_A2803_;
  assign new_A2799_ = new_A2767_ | new_A2804_;
  assign new_A2798_ = new_A2750_ & ~new_A2751_;
  assign new_A2797_ = ~new_A2750_ & new_A2751_;
  assign new_A2796_ = new_A2760_ | new_A2793_;
  assign new_A2795_ = ~new_A2760_ & ~new_A2794_;
  assign new_A2794_ = new_A2760_ & new_A2793_;
  assign new_A2793_ = ~new_A2749_ | ~new_A2774_;
  assign new_A2792_ = ~new_A2750_ & new_A2760_;
  assign new_A2791_ = new_A2750_ & ~new_A2760_;
  assign new_A2790_ = new_A2752_ & new_A2789_;
  assign new_A2789_ = new_A2808_ | new_A2807_;
  assign new_A2788_ = ~new_A2752_ & new_A2787_;
  assign new_A2787_ = new_A2810_ | new_A2809_;
  assign new_A2786_ = new_A2752_ | new_A2785_;
  assign new_A2785_ = new_A2806_ | new_A2805_;
  assign new_A2784_ = ~new_A2764_ & ~new_A2774_;
  assign new_A2783_ = new_A2764_ & new_A2774_;
  assign new_A2782_ = ~new_A2764_ | new_A2774_;
  assign new_A2781_ = new_A2748_ & ~new_A2749_;
  assign new_A2780_ = ~new_A2748_ & new_A2749_;
  assign new_A2779_ = new_A2801_ & ~new_A2802_;
  assign new_A2778_ = ~new_A2801_ & new_A2802_;
  assign new_A2777_ = ~new_A2800_ | ~new_A2799_;
  assign new_A2776_ = new_A2792_ | new_A2791_;
  assign new_A2775_ = new_A2798_ | new_A2797_;
  assign new_A2774_ = new_A2788_ | new_A2790_;
  assign new_A2773_ = ~new_A2795_ | ~new_A2796_;
  assign new_A2772_ = new_A2748_ & ~new_A2749_;
  assign new_A2771_ = new_A2762_ & ~new_A2774_;
  assign new_A2770_ = ~new_A2762_ & new_A2774_;
  assign new_A2769_ = ~new_A2760_ & new_A2786_;
  assign new_A2768_ = new_A2784_ | new_A2783_;
  assign new_A2767_ = new_A2781_ | new_A2780_;
  assign new_A2766_ = new_A2749_ | new_A2782_;
  assign new_A2765_ = new_A2774_ & new_A2777_;
  assign new_A2764_ = new_A2779_ | new_A2778_;
  assign new_A2763_ = new_A2774_ & new_A2773_;
  assign new_A2762_ = new_A2776_ & new_A2775_;
  assign new_A2761_ = new_A2771_ | new_A2770_;
  assign new_A2760_ = new_A2749_ | new_A2772_;
  assign A2759 = new_A2760_ | new_A2769_;
  assign A2758 = new_A2767_ & new_A2768_;
  assign A2757 = new_A2767_ & new_A2766_;
  assign A2756 = new_A2765_ | new_A2764_;
  assign A2755 = new_A2763_ | new_A2762_;
  assign A2754 = new_A2761_ & new_A2760_;
  assign new_A2753_ = new_A5572_;
  assign new_A2752_ = new_A5505_;
  assign new_A2751_ = new_A5438_;
  assign new_A2750_ = new_A5371_;
  assign new_A2749_ = new_A5304_;
  assign new_A2748_ = new_A5237_;
  assign new_A2747_ = ~new_A2686_ & new_A2700_;
  assign new_A2746_ = new_A2686_ & ~new_A2700_;
  assign new_A2745_ = new_A2686_ & ~new_A2700_;
  assign new_A2744_ = ~new_A2686_ & ~new_A2700_;
  assign new_A2743_ = new_A2686_ & new_A2700_;
  assign new_A2742_ = new_A2746_ | new_A2747_;
  assign new_A2741_ = ~new_A2686_ & new_A2700_;
  assign new_A2740_ = new_A2744_ | new_A2745_;
  assign new_A2739_ = ~new_A2715_ & ~new_A2735_;
  assign new_A2738_ = new_A2715_ & new_A2735_;
  assign new_A2737_ = ~new_A2682_ | ~new_A2707_;
  assign new_A2736_ = new_A2700_ & new_A2737_;
  assign new_A2735_ = new_A2683_ | new_A2684_;
  assign new_A2734_ = new_A2683_ | new_A2700_;
  assign new_A2733_ = ~new_A2700_ & ~new_A2736_;
  assign new_A2732_ = new_A2700_ | new_A2737_;
  assign new_A2731_ = new_A2683_ & ~new_A2684_;
  assign new_A2730_ = ~new_A2683_ & new_A2684_;
  assign new_A2729_ = new_A2693_ | new_A2726_;
  assign new_A2728_ = ~new_A2693_ & ~new_A2727_;
  assign new_A2727_ = new_A2693_ & new_A2726_;
  assign new_A2726_ = ~new_A2682_ | ~new_A2707_;
  assign new_A2725_ = ~new_A2683_ & new_A2693_;
  assign new_A2724_ = new_A2683_ & ~new_A2693_;
  assign new_A2723_ = new_A2685_ & new_A2722_;
  assign new_A2722_ = new_A2741_ | new_A2740_;
  assign new_A2721_ = ~new_A2685_ & new_A2720_;
  assign new_A2720_ = new_A2743_ | new_A2742_;
  assign new_A2719_ = new_A2685_ | new_A2718_;
  assign new_A2718_ = new_A2739_ | new_A2738_;
  assign new_A2717_ = ~new_A2697_ & ~new_A2707_;
  assign new_A2716_ = new_A2697_ & new_A2707_;
  assign new_A2715_ = ~new_A2697_ | new_A2707_;
  assign new_A2714_ = new_A2681_ & ~new_A2682_;
  assign new_A2713_ = ~new_A2681_ & new_A2682_;
  assign new_A2712_ = new_A2734_ & ~new_A2735_;
  assign new_A2711_ = ~new_A2734_ & new_A2735_;
  assign new_A2710_ = ~new_A2733_ | ~new_A2732_;
  assign new_A2709_ = new_A2725_ | new_A2724_;
  assign new_A2708_ = new_A2731_ | new_A2730_;
  assign new_A2707_ = new_A2721_ | new_A2723_;
  assign new_A2706_ = ~new_A2728_ | ~new_A2729_;
  assign new_A2705_ = new_A2681_ & ~new_A2682_;
  assign new_A2704_ = new_A2695_ & ~new_A2707_;
  assign new_A2703_ = ~new_A2695_ & new_A2707_;
  assign new_A2702_ = ~new_A2693_ & new_A2719_;
  assign new_A2701_ = new_A2717_ | new_A2716_;
  assign new_A2700_ = new_A2714_ | new_A2713_;
  assign new_A2699_ = new_A2682_ | new_A2715_;
  assign new_A2698_ = new_A2707_ & new_A2710_;
  assign new_A2697_ = new_A2712_ | new_A2711_;
  assign new_A2696_ = new_A2707_ & new_A2706_;
  assign new_A2695_ = new_A2709_ & new_A2708_;
  assign new_A2694_ = new_A2704_ | new_A2703_;
  assign new_A2693_ = new_A2682_ | new_A2705_;
  assign A2692 = new_A2693_ | new_A2702_;
  assign A2691 = new_A2700_ & new_A2701_;
  assign A2690 = new_A2700_ & new_A2699_;
  assign A2689 = new_A2698_ | new_A2697_;
  assign A2688 = new_A2696_ | new_A2695_;
  assign A2687 = new_A2694_ & new_A2693_;
  assign new_A2686_ = new_A5170_;
  assign new_A2685_ = new_A5103_;
  assign new_A2684_ = new_A5036_;
  assign new_A2683_ = new_A4969_;
  assign new_A2682_ = new_A4902_;
  assign new_A2681_ = new_A4835_;
  assign new_A2680_ = ~new_A2619_ & new_A2633_;
  assign new_A2679_ = new_A2619_ & ~new_A2633_;
  assign new_A2678_ = new_A2619_ & ~new_A2633_;
  assign new_A2677_ = ~new_A2619_ & ~new_A2633_;
  assign new_A2676_ = new_A2619_ & new_A2633_;
  assign new_A2675_ = new_A2679_ | new_A2680_;
  assign new_A2674_ = ~new_A2619_ & new_A2633_;
  assign new_A2673_ = new_A2677_ | new_A2678_;
  assign new_A2672_ = ~new_A2648_ & ~new_A2668_;
  assign new_A2671_ = new_A2648_ & new_A2668_;
  assign new_A2670_ = ~new_A2615_ | ~new_A2640_;
  assign new_A2669_ = new_A2633_ & new_A2670_;
  assign new_A2668_ = new_A2616_ | new_A2617_;
  assign new_A2667_ = new_A2616_ | new_A2633_;
  assign new_A2666_ = ~new_A2633_ & ~new_A2669_;
  assign new_A2665_ = new_A2633_ | new_A2670_;
  assign new_A2664_ = new_A2616_ & ~new_A2617_;
  assign new_A2663_ = ~new_A2616_ & new_A2617_;
  assign new_A2662_ = new_A2626_ | new_A2659_;
  assign new_A2661_ = ~new_A2626_ & ~new_A2660_;
  assign new_A2660_ = new_A2626_ & new_A2659_;
  assign new_A2659_ = ~new_A2615_ | ~new_A2640_;
  assign new_A2658_ = ~new_A2616_ & new_A2626_;
  assign new_A2657_ = new_A2616_ & ~new_A2626_;
  assign new_A2656_ = new_A2618_ & new_A2655_;
  assign new_A2655_ = new_A2674_ | new_A2673_;
  assign new_A2654_ = ~new_A2618_ & new_A2653_;
  assign new_A2653_ = new_A2676_ | new_A2675_;
  assign new_A2652_ = new_A2618_ | new_A2651_;
  assign new_A2651_ = new_A2672_ | new_A2671_;
  assign new_A2650_ = ~new_A2630_ & ~new_A2640_;
  assign new_A2649_ = new_A2630_ & new_A2640_;
  assign new_A2648_ = ~new_A2630_ | new_A2640_;
  assign new_A2647_ = new_A2614_ & ~new_A2615_;
  assign new_A2646_ = ~new_A2614_ & new_A2615_;
  assign new_A2645_ = new_A2667_ & ~new_A2668_;
  assign new_A2644_ = ~new_A2667_ & new_A2668_;
  assign new_A2643_ = ~new_A2666_ | ~new_A2665_;
  assign new_A2642_ = new_A2658_ | new_A2657_;
  assign new_A2641_ = new_A2664_ | new_A2663_;
  assign new_A2640_ = new_A2654_ | new_A2656_;
  assign new_A2639_ = ~new_A2661_ | ~new_A2662_;
  assign new_A2638_ = new_A2614_ & ~new_A2615_;
  assign new_A2637_ = new_A2628_ & ~new_A2640_;
  assign new_A2636_ = ~new_A2628_ & new_A2640_;
  assign new_A2635_ = ~new_A2626_ & new_A2652_;
  assign new_A2634_ = new_A2650_ | new_A2649_;
  assign new_A2633_ = new_A2647_ | new_A2646_;
  assign new_A2632_ = new_A2615_ | new_A2648_;
  assign new_A2631_ = new_A2640_ & new_A2643_;
  assign new_A2630_ = new_A2645_ | new_A2644_;
  assign new_A2629_ = new_A2640_ & new_A2639_;
  assign new_A2628_ = new_A2642_ & new_A2641_;
  assign new_A2627_ = new_A2637_ | new_A2636_;
  assign new_A2626_ = new_A2615_ | new_A2638_;
  assign A2625 = new_A2626_ | new_A2635_;
  assign A2624 = new_A2633_ & new_A2634_;
  assign A2623 = new_A2633_ & new_A2632_;
  assign A2622 = new_A2631_ | new_A2630_;
  assign A2621 = new_A2629_ | new_A2628_;
  assign A2620 = new_A2627_ & new_A2626_;
  assign new_A2619_ = new_A4768_;
  assign new_A2618_ = new_A4701_;
  assign new_A2617_ = new_A4634_;
  assign new_A2616_ = new_A4567_;
  assign new_A2615_ = new_A4500_;
  assign new_A2614_ = new_A4433_;
  assign new_A2613_ = ~new_A2552_ & new_A2566_;
  assign new_A2612_ = new_A2552_ & ~new_A2566_;
  assign new_A2611_ = new_A2552_ & ~new_A2566_;
  assign new_A2610_ = ~new_A2552_ & ~new_A2566_;
  assign new_A2609_ = new_A2552_ & new_A2566_;
  assign new_A2608_ = new_A2612_ | new_A2613_;
  assign new_A2607_ = ~new_A2552_ & new_A2566_;
  assign new_A2606_ = new_A2610_ | new_A2611_;
  assign new_A2605_ = ~new_A2581_ & ~new_A2601_;
  assign new_A2604_ = new_A2581_ & new_A2601_;
  assign new_A2603_ = ~new_A2548_ | ~new_A2573_;
  assign new_A2602_ = new_A2566_ & new_A2603_;
  assign new_A2601_ = new_A2549_ | new_A2550_;
  assign new_A2600_ = new_A2549_ | new_A2566_;
  assign new_A2599_ = ~new_A2566_ & ~new_A2602_;
  assign new_A2598_ = new_A2566_ | new_A2603_;
  assign new_A2597_ = new_A2549_ & ~new_A2550_;
  assign new_A2596_ = ~new_A2549_ & new_A2550_;
  assign new_A2595_ = new_A2559_ | new_A2592_;
  assign new_A2594_ = ~new_A2559_ & ~new_A2593_;
  assign new_A2593_ = new_A2559_ & new_A2592_;
  assign new_A2592_ = ~new_A2548_ | ~new_A2573_;
  assign new_A2591_ = ~new_A2549_ & new_A2559_;
  assign new_A2590_ = new_A2549_ & ~new_A2559_;
  assign new_A2589_ = new_A2551_ & new_A2588_;
  assign new_A2588_ = new_A2607_ | new_A2606_;
  assign new_A2587_ = ~new_A2551_ & new_A2586_;
  assign new_A2586_ = new_A2609_ | new_A2608_;
  assign new_A2585_ = new_A2551_ | new_A2584_;
  assign new_A2584_ = new_A2605_ | new_A2604_;
  assign new_A2583_ = ~new_A2563_ & ~new_A2573_;
  assign new_A2582_ = new_A2563_ & new_A2573_;
  assign new_A2581_ = ~new_A2563_ | new_A2573_;
  assign new_A2580_ = new_A2547_ & ~new_A2548_;
  assign new_A2579_ = ~new_A2547_ & new_A2548_;
  assign new_A2578_ = new_A2600_ & ~new_A2601_;
  assign new_A2577_ = ~new_A2600_ & new_A2601_;
  assign new_A2576_ = ~new_A2599_ | ~new_A2598_;
  assign new_A2575_ = new_A2591_ | new_A2590_;
  assign new_A2574_ = new_A2597_ | new_A2596_;
  assign new_A2573_ = new_A2587_ | new_A2589_;
  assign new_A2572_ = ~new_A2594_ | ~new_A2595_;
  assign new_A2571_ = new_A2547_ & ~new_A2548_;
  assign new_A2570_ = new_A2561_ & ~new_A2573_;
  assign new_A2569_ = ~new_A2561_ & new_A2573_;
  assign new_A2568_ = ~new_A2559_ & new_A2585_;
  assign new_A2567_ = new_A2583_ | new_A2582_;
  assign new_A2566_ = new_A2580_ | new_A2579_;
  assign new_A2565_ = new_A2548_ | new_A2581_;
  assign new_A2564_ = new_A2573_ & new_A2576_;
  assign new_A2563_ = new_A2578_ | new_A2577_;
  assign new_A2562_ = new_A2573_ & new_A2572_;
  assign new_A2561_ = new_A2575_ & new_A2574_;
  assign new_A2560_ = new_A2570_ | new_A2569_;
  assign new_A2559_ = new_A2548_ | new_A2571_;
  assign A2558 = new_A2559_ | new_A2568_;
  assign A2557 = new_A2566_ & new_A2567_;
  assign A2556 = new_A2566_ & new_A2565_;
  assign A2555 = new_A2564_ | new_A2563_;
  assign A2554 = new_A2562_ | new_A2561_;
  assign A2553 = new_A2560_ & new_A2559_;
  assign new_A2552_ = new_A4366_;
  assign new_A2551_ = new_A4299_;
  assign new_A2550_ = new_A4232_;
  assign new_A2549_ = new_A4165_;
  assign new_A2548_ = new_A4098_;
  assign new_A2547_ = new_A4031_;
  assign new_A2546_ = ~new_A2485_ & new_A2499_;
  assign new_A2545_ = new_A2485_ & ~new_A2499_;
  assign new_A2544_ = new_A2485_ & ~new_A2499_;
  assign new_A2543_ = ~new_A2485_ & ~new_A2499_;
  assign new_A2542_ = new_A2485_ & new_A2499_;
  assign new_A2541_ = new_A2545_ | new_A2546_;
  assign new_A2540_ = ~new_A2485_ & new_A2499_;
  assign new_A2539_ = new_A2543_ | new_A2544_;
  assign new_A2538_ = ~new_A2514_ & ~new_A2534_;
  assign new_A2537_ = new_A2514_ & new_A2534_;
  assign new_A2536_ = ~new_A2481_ | ~new_A2506_;
  assign new_A2535_ = new_A2499_ & new_A2536_;
  assign new_A2534_ = new_A2482_ | new_A2483_;
  assign new_A2533_ = new_A2482_ | new_A2499_;
  assign new_A2532_ = ~new_A2499_ & ~new_A2535_;
  assign new_A2531_ = new_A2499_ | new_A2536_;
  assign new_A2530_ = new_A2482_ & ~new_A2483_;
  assign new_A2529_ = ~new_A2482_ & new_A2483_;
  assign new_A2528_ = new_A2492_ | new_A2525_;
  assign new_A2527_ = ~new_A2492_ & ~new_A2526_;
  assign new_A2526_ = new_A2492_ & new_A2525_;
  assign new_A2525_ = ~new_A2481_ | ~new_A2506_;
  assign new_A2524_ = ~new_A2482_ & new_A2492_;
  assign new_A2523_ = new_A2482_ & ~new_A2492_;
  assign new_A2522_ = new_A2484_ & new_A2521_;
  assign new_A2521_ = new_A2540_ | new_A2539_;
  assign new_A2520_ = ~new_A2484_ & new_A2519_;
  assign new_A2519_ = new_A2542_ | new_A2541_;
  assign new_A2518_ = new_A2484_ | new_A2517_;
  assign new_A2517_ = new_A2538_ | new_A2537_;
  assign new_A2516_ = ~new_A2496_ & ~new_A2506_;
  assign new_A2515_ = new_A2496_ & new_A2506_;
  assign new_A2514_ = ~new_A2496_ | new_A2506_;
  assign new_A2513_ = new_A2480_ & ~new_A2481_;
  assign new_A2512_ = ~new_A2480_ & new_A2481_;
  assign new_A2511_ = new_A2533_ & ~new_A2534_;
  assign new_A2510_ = ~new_A2533_ & new_A2534_;
  assign new_A2509_ = ~new_A2532_ | ~new_A2531_;
  assign new_A2508_ = new_A2524_ | new_A2523_;
  assign new_A2507_ = new_A2530_ | new_A2529_;
  assign new_A2506_ = new_A2520_ | new_A2522_;
  assign new_A2505_ = ~new_A2527_ | ~new_A2528_;
  assign new_A2504_ = new_A2480_ & ~new_A2481_;
  assign new_A2503_ = new_A2494_ & ~new_A2506_;
  assign new_A2502_ = ~new_A2494_ & new_A2506_;
  assign new_A2501_ = ~new_A2492_ & new_A2518_;
  assign new_A2500_ = new_A2516_ | new_A2515_;
  assign new_A2499_ = new_A2513_ | new_A2512_;
  assign new_A2498_ = new_A2481_ | new_A2514_;
  assign new_A2497_ = new_A2506_ & new_A2509_;
  assign new_A2496_ = new_A2511_ | new_A2510_;
  assign new_A2495_ = new_A2506_ & new_A2505_;
  assign new_A2494_ = new_A2508_ & new_A2507_;
  assign new_A2493_ = new_A2503_ | new_A2502_;
  assign new_A2492_ = new_A2481_ | new_A2504_;
  assign A2491 = new_A2492_ | new_A2501_;
  assign A2490 = new_A2499_ & new_A2500_;
  assign A2489 = new_A2499_ & new_A2498_;
  assign A2488 = new_A2497_ | new_A2496_;
  assign A2487 = new_A2495_ | new_A2494_;
  assign A2486 = new_A2493_ & new_A2492_;
  assign new_A2485_ = new_A3964_;
  assign new_A2484_ = new_A3897_;
  assign new_A2483_ = new_A3830_;
  assign new_A2482_ = new_A3763_;
  assign new_A2481_ = new_A3696_;
  assign new_A2480_ = new_A3629_;
  assign new_A2479_ = ~new_A2418_ & new_A2432_;
  assign new_A2478_ = new_A2418_ & ~new_A2432_;
  assign new_A2477_ = new_A2418_ & ~new_A2432_;
  assign new_A2476_ = ~new_A2418_ & ~new_A2432_;
  assign new_A2475_ = new_A2418_ & new_A2432_;
  assign new_A2474_ = new_A2478_ | new_A2479_;
  assign new_A2473_ = ~new_A2418_ & new_A2432_;
  assign new_A2472_ = new_A2476_ | new_A2477_;
  assign new_A2471_ = ~new_A2447_ & ~new_A2467_;
  assign new_A2470_ = new_A2447_ & new_A2467_;
  assign new_A2469_ = ~new_A2414_ | ~new_A2439_;
  assign new_A2468_ = new_A2432_ & new_A2469_;
  assign new_A2467_ = new_A2415_ | new_A2416_;
  assign new_A2466_ = new_A2415_ | new_A2432_;
  assign new_A2465_ = ~new_A2432_ & ~new_A2468_;
  assign new_A2464_ = new_A2432_ | new_A2469_;
  assign new_A2463_ = new_A2415_ & ~new_A2416_;
  assign new_A2462_ = ~new_A2415_ & new_A2416_;
  assign new_A2461_ = new_A2425_ | new_A2458_;
  assign new_A2460_ = ~new_A2425_ & ~new_A2459_;
  assign new_A2459_ = new_A2425_ & new_A2458_;
  assign new_A2458_ = ~new_A2414_ | ~new_A2439_;
  assign new_A2457_ = ~new_A2415_ & new_A2425_;
  assign new_A2456_ = new_A2415_ & ~new_A2425_;
  assign new_A2455_ = new_A2417_ & new_A2454_;
  assign new_A2454_ = new_A2473_ | new_A2472_;
  assign new_A2453_ = ~new_A2417_ & new_A2452_;
  assign new_A2452_ = new_A2475_ | new_A2474_;
  assign new_A2451_ = new_A2417_ | new_A2450_;
  assign new_A2450_ = new_A2471_ | new_A2470_;
  assign new_A2449_ = ~new_A2429_ & ~new_A2439_;
  assign new_A2448_ = new_A2429_ & new_A2439_;
  assign new_A2447_ = ~new_A2429_ | new_A2439_;
  assign new_A2446_ = new_A2413_ & ~new_A2414_;
  assign new_A2445_ = ~new_A2413_ & new_A2414_;
  assign new_A2444_ = new_A2466_ & ~new_A2467_;
  assign new_A2443_ = ~new_A2466_ & new_A2467_;
  assign new_A2442_ = ~new_A2465_ | ~new_A2464_;
  assign new_A2441_ = new_A2457_ | new_A2456_;
  assign new_A2440_ = new_A2463_ | new_A2462_;
  assign new_A2439_ = new_A2453_ | new_A2455_;
  assign new_A2438_ = ~new_A2460_ | ~new_A2461_;
  assign new_A2437_ = new_A2413_ & ~new_A2414_;
  assign new_A2436_ = new_A2427_ & ~new_A2439_;
  assign new_A2435_ = ~new_A2427_ & new_A2439_;
  assign new_A2434_ = ~new_A2425_ & new_A2451_;
  assign new_A2433_ = new_A2449_ | new_A2448_;
  assign new_A2432_ = new_A2446_ | new_A2445_;
  assign new_A2431_ = new_A2414_ | new_A2447_;
  assign new_A2430_ = new_A2439_ & new_A2442_;
  assign new_A2429_ = new_A2444_ | new_A2443_;
  assign new_A2428_ = new_A2439_ & new_A2438_;
  assign new_A2427_ = new_A2441_ & new_A2440_;
  assign new_A2426_ = new_A2436_ | new_A2435_;
  assign new_A2425_ = new_A2414_ | new_A2437_;
  assign A2424 = new_A2425_ | new_A2434_;
  assign A2423 = new_A2432_ & new_A2433_;
  assign A2422 = new_A2432_ & new_A2431_;
  assign A2421 = new_A2430_ | new_A2429_;
  assign A2420 = new_A2428_ | new_A2427_;
  assign A2419 = new_A2426_ & new_A2425_;
  assign new_A2418_ = new_A3562_;
  assign new_A2417_ = new_A3495_;
  assign new_A2416_ = new_A3428_;
  assign new_A2415_ = new_A3361_;
  assign new_A2414_ = new_A3294_;
  assign new_A2413_ = new_A3224_;
  assign new_A2412_ = ~new_A2351_ & new_A2365_;
  assign new_A2411_ = new_A2351_ & ~new_A2365_;
  assign new_A2410_ = new_A2351_ & ~new_A2365_;
  assign new_A2409_ = ~new_A2351_ & ~new_A2365_;
  assign new_A2408_ = new_A2351_ & new_A2365_;
  assign new_A2407_ = new_A2411_ | new_A2412_;
  assign new_A2406_ = ~new_A2351_ & new_A2365_;
  assign new_A2405_ = new_A2409_ | new_A2410_;
  assign new_A2404_ = ~new_A2380_ & ~new_A2400_;
  assign new_A2403_ = new_A2380_ & new_A2400_;
  assign new_A2402_ = ~new_A2347_ | ~new_A2372_;
  assign new_A2401_ = new_A2365_ & new_A2402_;
  assign new_A2400_ = new_A2348_ | new_A2349_;
  assign new_A2399_ = new_A2348_ | new_A2365_;
  assign new_A2398_ = ~new_A2365_ & ~new_A2401_;
  assign new_A2397_ = new_A2365_ | new_A2402_;
  assign new_A2396_ = new_A2348_ & ~new_A2349_;
  assign new_A2395_ = ~new_A2348_ & new_A2349_;
  assign new_A2394_ = new_A2358_ | new_A2391_;
  assign new_A2393_ = ~new_A2358_ & ~new_A2392_;
  assign new_A2392_ = new_A2358_ & new_A2391_;
  assign new_A2391_ = ~new_A2347_ | ~new_A2372_;
  assign new_A2390_ = ~new_A2348_ & new_A2358_;
  assign new_A2389_ = new_A2348_ & ~new_A2358_;
  assign new_A2388_ = new_A2350_ & new_A2387_;
  assign new_A2387_ = new_A2406_ | new_A2405_;
  assign new_A2386_ = ~new_A2350_ & new_A2385_;
  assign new_A2385_ = new_A2408_ | new_A2407_;
  assign new_A2384_ = new_A2350_ | new_A2383_;
  assign new_A2383_ = new_A2404_ | new_A2403_;
  assign new_A2382_ = ~new_A2362_ & ~new_A2372_;
  assign new_A2381_ = new_A2362_ & new_A2372_;
  assign new_A2380_ = ~new_A2362_ | new_A2372_;
  assign new_A2379_ = new_A2346_ & ~new_A2347_;
  assign new_A2378_ = ~new_A2346_ & new_A2347_;
  assign new_A2377_ = new_A2399_ & ~new_A2400_;
  assign new_A2376_ = ~new_A2399_ & new_A2400_;
  assign new_A2375_ = ~new_A2398_ | ~new_A2397_;
  assign new_A2374_ = new_A2390_ | new_A2389_;
  assign new_A2373_ = new_A2396_ | new_A2395_;
  assign new_A2372_ = new_A2386_ | new_A2388_;
  assign new_A2371_ = ~new_A2393_ | ~new_A2394_;
  assign new_A2370_ = new_A2346_ & ~new_A2347_;
  assign new_A2369_ = new_A2360_ & ~new_A2372_;
  assign new_A2368_ = ~new_A2360_ & new_A2372_;
  assign new_A2367_ = ~new_A2358_ & new_A2384_;
  assign new_A2366_ = new_A2382_ | new_A2381_;
  assign new_A2365_ = new_A2379_ | new_A2378_;
  assign new_A2364_ = new_A2347_ | new_A2380_;
  assign new_A2363_ = new_A2372_ & new_A2375_;
  assign new_A2362_ = new_A2377_ | new_A2376_;
  assign new_A2361_ = new_A2372_ & new_A2371_;
  assign new_A2360_ = new_A2374_ & new_A2373_;
  assign new_A2359_ = new_A2369_ | new_A2368_;
  assign new_A2358_ = new_A2347_ | new_A2370_;
  assign A2357 = new_A2358_ | new_A2367_;
  assign A2356 = new_A2365_ & new_A2366_;
  assign A2355 = new_A2365_ & new_A2364_;
  assign A2354 = new_A2363_ | new_A2362_;
  assign A2353 = new_A2361_ | new_A2360_;
  assign A2352 = new_A2359_ & new_A2358_;
  assign new_A2351_ = new_A5571_;
  assign new_A2350_ = new_A5504_;
  assign new_A2349_ = new_A5437_;
  assign new_A2348_ = new_A5370_;
  assign new_A2347_ = new_A5303_;
  assign new_A2346_ = new_A5236_;
  assign new_A2345_ = ~new_A2284_ & new_A2298_;
  assign new_A2344_ = new_A2284_ & ~new_A2298_;
  assign new_A2343_ = new_A2284_ & ~new_A2298_;
  assign new_A2342_ = ~new_A2284_ & ~new_A2298_;
  assign new_A2341_ = new_A2284_ & new_A2298_;
  assign new_A2340_ = new_A2344_ | new_A2345_;
  assign new_A2339_ = ~new_A2284_ & new_A2298_;
  assign new_A2338_ = new_A2342_ | new_A2343_;
  assign new_A2337_ = ~new_A2313_ & ~new_A2333_;
  assign new_A2336_ = new_A2313_ & new_A2333_;
  assign new_A2335_ = ~new_A2280_ | ~new_A2305_;
  assign new_A2334_ = new_A2298_ & new_A2335_;
  assign new_A2333_ = new_A2281_ | new_A2282_;
  assign new_A2332_ = new_A2281_ | new_A2298_;
  assign new_A2331_ = ~new_A2298_ & ~new_A2334_;
  assign new_A2330_ = new_A2298_ | new_A2335_;
  assign new_A2329_ = new_A2281_ & ~new_A2282_;
  assign new_A2328_ = ~new_A2281_ & new_A2282_;
  assign new_A2327_ = new_A2291_ | new_A2324_;
  assign new_A2326_ = ~new_A2291_ & ~new_A2325_;
  assign new_A2325_ = new_A2291_ & new_A2324_;
  assign new_A2324_ = ~new_A2280_ | ~new_A2305_;
  assign new_A2323_ = ~new_A2281_ & new_A2291_;
  assign new_A2322_ = new_A2281_ & ~new_A2291_;
  assign new_A2321_ = new_A2283_ & new_A2320_;
  assign new_A2320_ = new_A2339_ | new_A2338_;
  assign new_A2319_ = ~new_A2283_ & new_A2318_;
  assign new_A2318_ = new_A2341_ | new_A2340_;
  assign new_A2317_ = new_A2283_ | new_A2316_;
  assign new_A2316_ = new_A2337_ | new_A2336_;
  assign new_A2315_ = ~new_A2295_ & ~new_A2305_;
  assign new_A2314_ = new_A2295_ & new_A2305_;
  assign new_A2313_ = ~new_A2295_ | new_A2305_;
  assign new_A2312_ = new_A2279_ & ~new_A2280_;
  assign new_A2311_ = ~new_A2279_ & new_A2280_;
  assign new_A2310_ = new_A2332_ & ~new_A2333_;
  assign new_A2309_ = ~new_A2332_ & new_A2333_;
  assign new_A2308_ = ~new_A2331_ | ~new_A2330_;
  assign new_A2307_ = new_A2323_ | new_A2322_;
  assign new_A2306_ = new_A2329_ | new_A2328_;
  assign new_A2305_ = new_A2319_ | new_A2321_;
  assign new_A2304_ = ~new_A2326_ | ~new_A2327_;
  assign new_A2303_ = new_A2279_ & ~new_A2280_;
  assign new_A2302_ = new_A2293_ & ~new_A2305_;
  assign new_A2301_ = ~new_A2293_ & new_A2305_;
  assign new_A2300_ = ~new_A2291_ & new_A2317_;
  assign new_A2299_ = new_A2315_ | new_A2314_;
  assign new_A2298_ = new_A2312_ | new_A2311_;
  assign new_A2297_ = new_A2280_ | new_A2313_;
  assign new_A2296_ = new_A2305_ & new_A2308_;
  assign new_A2295_ = new_A2310_ | new_A2309_;
  assign new_A2294_ = new_A2305_ & new_A2304_;
  assign new_A2293_ = new_A2307_ & new_A2306_;
  assign new_A2292_ = new_A2302_ | new_A2301_;
  assign new_A2291_ = new_A2280_ | new_A2303_;
  assign A2290 = new_A2291_ | new_A2300_;
  assign A2289 = new_A2298_ & new_A2299_;
  assign A2288 = new_A2298_ & new_A2297_;
  assign A2287 = new_A2296_ | new_A2295_;
  assign A2286 = new_A2294_ | new_A2293_;
  assign A2285 = new_A2292_ & new_A2291_;
  assign new_A2284_ = new_A5169_;
  assign new_A2283_ = new_A5102_;
  assign new_A2282_ = new_A5035_;
  assign new_A2281_ = new_A4968_;
  assign new_A2280_ = new_A4901_;
  assign new_A2279_ = new_A4834_;
  assign new_A2278_ = ~new_A2217_ & new_A2231_;
  assign new_A2277_ = new_A2217_ & ~new_A2231_;
  assign new_A2276_ = new_A2217_ & ~new_A2231_;
  assign new_A2275_ = ~new_A2217_ & ~new_A2231_;
  assign new_A2274_ = new_A2217_ & new_A2231_;
  assign new_A2273_ = new_A2277_ | new_A2278_;
  assign new_A2272_ = ~new_A2217_ & new_A2231_;
  assign new_A2271_ = new_A2275_ | new_A2276_;
  assign new_A2270_ = ~new_A2246_ & ~new_A2266_;
  assign new_A2269_ = new_A2246_ & new_A2266_;
  assign new_A2268_ = ~new_A2213_ | ~new_A2238_;
  assign new_A2267_ = new_A2231_ & new_A2268_;
  assign new_A2266_ = new_A2214_ | new_A2215_;
  assign new_A2265_ = new_A2214_ | new_A2231_;
  assign new_A2264_ = ~new_A2231_ & ~new_A2267_;
  assign new_A2263_ = new_A2231_ | new_A2268_;
  assign new_A2262_ = new_A2214_ & ~new_A2215_;
  assign new_A2261_ = ~new_A2214_ & new_A2215_;
  assign new_A2260_ = new_A2224_ | new_A2257_;
  assign new_A2259_ = ~new_A2224_ & ~new_A2258_;
  assign new_A2258_ = new_A2224_ & new_A2257_;
  assign new_A2257_ = ~new_A2213_ | ~new_A2238_;
  assign new_A2256_ = ~new_A2214_ & new_A2224_;
  assign new_A2255_ = new_A2214_ & ~new_A2224_;
  assign new_A2254_ = new_A2216_ & new_A2253_;
  assign new_A2253_ = new_A2272_ | new_A2271_;
  assign new_A2252_ = ~new_A2216_ & new_A2251_;
  assign new_A2251_ = new_A2274_ | new_A2273_;
  assign new_A2250_ = new_A2216_ | new_A2249_;
  assign new_A2249_ = new_A2270_ | new_A2269_;
  assign new_A2248_ = ~new_A2228_ & ~new_A2238_;
  assign new_A2247_ = new_A2228_ & new_A2238_;
  assign new_A2246_ = ~new_A2228_ | new_A2238_;
  assign new_A2245_ = new_A2212_ & ~new_A2213_;
  assign new_A2244_ = ~new_A2212_ & new_A2213_;
  assign new_A2243_ = new_A2265_ & ~new_A2266_;
  assign new_A2242_ = ~new_A2265_ & new_A2266_;
  assign new_A2241_ = ~new_A2264_ | ~new_A2263_;
  assign new_A2240_ = new_A2256_ | new_A2255_;
  assign new_A2239_ = new_A2262_ | new_A2261_;
  assign new_A2238_ = new_A2252_ | new_A2254_;
  assign new_A2237_ = ~new_A2259_ | ~new_A2260_;
  assign new_A2236_ = new_A2212_ & ~new_A2213_;
  assign new_A2235_ = new_A2226_ & ~new_A2238_;
  assign new_A2234_ = ~new_A2226_ & new_A2238_;
  assign new_A2233_ = ~new_A2224_ & new_A2250_;
  assign new_A2232_ = new_A2248_ | new_A2247_;
  assign new_A2231_ = new_A2245_ | new_A2244_;
  assign new_A2230_ = new_A2213_ | new_A2246_;
  assign new_A2229_ = new_A2238_ & new_A2241_;
  assign new_A2228_ = new_A2243_ | new_A2242_;
  assign new_A2227_ = new_A2238_ & new_A2237_;
  assign new_A2226_ = new_A2240_ & new_A2239_;
  assign new_A2225_ = new_A2235_ | new_A2234_;
  assign new_A2224_ = new_A2213_ | new_A2236_;
  assign A2223 = new_A2224_ | new_A2233_;
  assign A2222 = new_A2231_ & new_A2232_;
  assign A2221 = new_A2231_ & new_A2230_;
  assign A2220 = new_A2229_ | new_A2228_;
  assign A2219 = new_A2227_ | new_A2226_;
  assign A2218 = new_A2225_ & new_A2224_;
  assign new_A2217_ = new_A4767_;
  assign new_A2216_ = new_A4700_;
  assign new_A2215_ = new_A4633_;
  assign new_A2214_ = new_A4566_;
  assign new_A2213_ = new_A4499_;
  assign new_A2212_ = new_A4432_;
  assign new_A2211_ = ~new_A2150_ & new_A2164_;
  assign new_A2210_ = new_A2150_ & ~new_A2164_;
  assign new_A2209_ = new_A2150_ & ~new_A2164_;
  assign new_A2208_ = ~new_A2150_ & ~new_A2164_;
  assign new_A2207_ = new_A2150_ & new_A2164_;
  assign new_A2206_ = new_A2210_ | new_A2211_;
  assign new_A2205_ = ~new_A2150_ & new_A2164_;
  assign new_A2204_ = new_A2208_ | new_A2209_;
  assign new_A2203_ = ~new_A2179_ & ~new_A2199_;
  assign new_A2202_ = new_A2179_ & new_A2199_;
  assign new_A2201_ = ~new_A2146_ | ~new_A2171_;
  assign new_A2200_ = new_A2164_ & new_A2201_;
  assign new_A2199_ = new_A2147_ | new_A2148_;
  assign new_A2198_ = new_A2147_ | new_A2164_;
  assign new_A2197_ = ~new_A2164_ & ~new_A2200_;
  assign new_A2196_ = new_A2164_ | new_A2201_;
  assign new_A2195_ = new_A2147_ & ~new_A2148_;
  assign new_A2194_ = ~new_A2147_ & new_A2148_;
  assign new_A2193_ = new_A2157_ | new_A2190_;
  assign new_A2192_ = ~new_A2157_ & ~new_A2191_;
  assign new_A2191_ = new_A2157_ & new_A2190_;
  assign new_A2190_ = ~new_A2146_ | ~new_A2171_;
  assign new_A2189_ = ~new_A2147_ & new_A2157_;
  assign new_A2188_ = new_A2147_ & ~new_A2157_;
  assign new_A2187_ = new_A2149_ & new_A2186_;
  assign new_A2186_ = new_A2205_ | new_A2204_;
  assign new_A2185_ = ~new_A2149_ & new_A2184_;
  assign new_A2184_ = new_A2207_ | new_A2206_;
  assign new_A2183_ = new_A2149_ | new_A2182_;
  assign new_A2182_ = new_A2203_ | new_A2202_;
  assign new_A2181_ = ~new_A2161_ & ~new_A2171_;
  assign new_A2180_ = new_A2161_ & new_A2171_;
  assign new_A2179_ = ~new_A2161_ | new_A2171_;
  assign new_A2178_ = new_A2145_ & ~new_A2146_;
  assign new_A2177_ = ~new_A2145_ & new_A2146_;
  assign new_A2176_ = new_A2198_ & ~new_A2199_;
  assign new_A2175_ = ~new_A2198_ & new_A2199_;
  assign new_A2174_ = ~new_A2197_ | ~new_A2196_;
  assign new_A2173_ = new_A2189_ | new_A2188_;
  assign new_A2172_ = new_A2195_ | new_A2194_;
  assign new_A2171_ = new_A2185_ | new_A2187_;
  assign new_A2170_ = ~new_A2192_ | ~new_A2193_;
  assign new_A2169_ = new_A2145_ & ~new_A2146_;
  assign new_A2168_ = new_A2159_ & ~new_A2171_;
  assign new_A2167_ = ~new_A2159_ & new_A2171_;
  assign new_A2166_ = ~new_A2157_ & new_A2183_;
  assign new_A2165_ = new_A2181_ | new_A2180_;
  assign new_A2164_ = new_A2178_ | new_A2177_;
  assign new_A2163_ = new_A2146_ | new_A2179_;
  assign new_A2162_ = new_A2171_ & new_A2174_;
  assign new_A2161_ = new_A2176_ | new_A2175_;
  assign new_A2160_ = new_A2171_ & new_A2170_;
  assign new_A2159_ = new_A2173_ & new_A2172_;
  assign new_A2158_ = new_A2168_ | new_A2167_;
  assign new_A2157_ = new_A2146_ | new_A2169_;
  assign A2156 = new_A2157_ | new_A2166_;
  assign A2155 = new_A2164_ & new_A2165_;
  assign A2154 = new_A2164_ & new_A2163_;
  assign A2153 = new_A2162_ | new_A2161_;
  assign A2152 = new_A2160_ | new_A2159_;
  assign A2151 = new_A2158_ & new_A2157_;
  assign new_A2150_ = new_A4365_;
  assign new_A2149_ = new_A4298_;
  assign new_A2148_ = new_A4231_;
  assign new_A2147_ = new_A4164_;
  assign new_A2146_ = new_A4097_;
  assign new_A2145_ = new_A4030_;
  assign new_A2144_ = ~new_A2083_ & new_A2097_;
  assign new_A2143_ = new_A2083_ & ~new_A2097_;
  assign new_A2142_ = new_A2083_ & ~new_A2097_;
  assign new_A2141_ = ~new_A2083_ & ~new_A2097_;
  assign new_A2140_ = new_A2083_ & new_A2097_;
  assign new_A2139_ = new_A2143_ | new_A2144_;
  assign new_A2138_ = ~new_A2083_ & new_A2097_;
  assign new_A2137_ = new_A2141_ | new_A2142_;
  assign new_A2136_ = ~new_A2112_ & ~new_A2132_;
  assign new_A2135_ = new_A2112_ & new_A2132_;
  assign new_A2134_ = ~new_A2079_ | ~new_A2104_;
  assign new_A2133_ = new_A2097_ & new_A2134_;
  assign new_A2132_ = new_A2080_ | new_A2081_;
  assign new_A2131_ = new_A2080_ | new_A2097_;
  assign new_A2130_ = ~new_A2097_ & ~new_A2133_;
  assign new_A2129_ = new_A2097_ | new_A2134_;
  assign new_A2128_ = new_A2080_ & ~new_A2081_;
  assign new_A2127_ = ~new_A2080_ & new_A2081_;
  assign new_A2126_ = new_A2090_ | new_A2123_;
  assign new_A2125_ = ~new_A2090_ & ~new_A2124_;
  assign new_A2124_ = new_A2090_ & new_A2123_;
  assign new_A2123_ = ~new_A2079_ | ~new_A2104_;
  assign new_A2122_ = ~new_A2080_ & new_A2090_;
  assign new_A2121_ = new_A2080_ & ~new_A2090_;
  assign new_A2120_ = new_A2082_ & new_A2119_;
  assign new_A2119_ = new_A2138_ | new_A2137_;
  assign new_A2118_ = ~new_A2082_ & new_A2117_;
  assign new_A2117_ = new_A2140_ | new_A2139_;
  assign new_A2116_ = new_A2082_ | new_A2115_;
  assign new_A2115_ = new_A2136_ | new_A2135_;
  assign new_A2114_ = ~new_A2094_ & ~new_A2104_;
  assign new_A2113_ = new_A2094_ & new_A2104_;
  assign new_A2112_ = ~new_A2094_ | new_A2104_;
  assign new_A2111_ = new_A2078_ & ~new_A2079_;
  assign new_A2110_ = ~new_A2078_ & new_A2079_;
  assign new_A2109_ = new_A2131_ & ~new_A2132_;
  assign new_A2108_ = ~new_A2131_ & new_A2132_;
  assign new_A2107_ = ~new_A2130_ | ~new_A2129_;
  assign new_A2106_ = new_A2122_ | new_A2121_;
  assign new_A2105_ = new_A2128_ | new_A2127_;
  assign new_A2104_ = new_A2118_ | new_A2120_;
  assign new_A2103_ = ~new_A2125_ | ~new_A2126_;
  assign new_A2102_ = new_A2078_ & ~new_A2079_;
  assign new_A2101_ = new_A2092_ & ~new_A2104_;
  assign new_A2100_ = ~new_A2092_ & new_A2104_;
  assign new_A2099_ = ~new_A2090_ & new_A2116_;
  assign new_A2098_ = new_A2114_ | new_A2113_;
  assign new_A2097_ = new_A2111_ | new_A2110_;
  assign new_A2096_ = new_A2079_ | new_A2112_;
  assign new_A2095_ = new_A2104_ & new_A2107_;
  assign new_A2094_ = new_A2109_ | new_A2108_;
  assign new_A2093_ = new_A2104_ & new_A2103_;
  assign new_A2092_ = new_A2106_ & new_A2105_;
  assign new_A2091_ = new_A2101_ | new_A2100_;
  assign new_A2090_ = new_A2079_ | new_A2102_;
  assign A2089 = new_A2090_ | new_A2099_;
  assign A2088 = new_A2097_ & new_A2098_;
  assign A2087 = new_A2097_ & new_A2096_;
  assign A2086 = new_A2095_ | new_A2094_;
  assign A2085 = new_A2093_ | new_A2092_;
  assign A2084 = new_A2091_ & new_A2090_;
  assign new_A2083_ = new_A3963_;
  assign new_A2082_ = new_A3896_;
  assign new_A2081_ = new_A3829_;
  assign new_A2080_ = new_A3762_;
  assign new_A2079_ = new_A3695_;
  assign new_A2078_ = new_A3628_;
  assign new_A2077_ = ~new_A2016_ & new_A2030_;
  assign new_A2076_ = new_A2016_ & ~new_A2030_;
  assign new_A2075_ = new_A2016_ & ~new_A2030_;
  assign new_A2074_ = ~new_A2016_ & ~new_A2030_;
  assign new_A2073_ = new_A2016_ & new_A2030_;
  assign new_A2072_ = new_A2076_ | new_A2077_;
  assign new_A2071_ = ~new_A2016_ & new_A2030_;
  assign new_A2070_ = new_A2074_ | new_A2075_;
  assign new_A2069_ = ~new_A2045_ & ~new_A2065_;
  assign new_A2068_ = new_A2045_ & new_A2065_;
  assign new_A2067_ = ~new_A2012_ | ~new_A2037_;
  assign new_A2066_ = new_A2030_ & new_A2067_;
  assign new_A2065_ = new_A2013_ | new_A2014_;
  assign new_A2064_ = new_A2013_ | new_A2030_;
  assign new_A2063_ = ~new_A2030_ & ~new_A2066_;
  assign new_A2062_ = new_A2030_ | new_A2067_;
  assign new_A2061_ = new_A2013_ & ~new_A2014_;
  assign new_A2060_ = ~new_A2013_ & new_A2014_;
  assign new_A2059_ = new_A2023_ | new_A2056_;
  assign new_A2058_ = ~new_A2023_ & ~new_A2057_;
  assign new_A2057_ = new_A2023_ & new_A2056_;
  assign new_A2056_ = ~new_A2012_ | ~new_A2037_;
  assign new_A2055_ = ~new_A2013_ & new_A2023_;
  assign new_A2054_ = new_A2013_ & ~new_A2023_;
  assign new_A2053_ = new_A2015_ & new_A2052_;
  assign new_A2052_ = new_A2071_ | new_A2070_;
  assign new_A2051_ = ~new_A2015_ & new_A2050_;
  assign new_A2050_ = new_A2073_ | new_A2072_;
  assign new_A2049_ = new_A2015_ | new_A2048_;
  assign new_A2048_ = new_A2069_ | new_A2068_;
  assign new_A2047_ = ~new_A2027_ & ~new_A2037_;
  assign new_A2046_ = new_A2027_ & new_A2037_;
  assign new_A2045_ = ~new_A2027_ | new_A2037_;
  assign new_A2044_ = new_A2011_ & ~new_A2012_;
  assign new_A2043_ = ~new_A2011_ & new_A2012_;
  assign new_A2042_ = new_A2064_ & ~new_A2065_;
  assign new_A2041_ = ~new_A2064_ & new_A2065_;
  assign new_A2040_ = ~new_A2063_ | ~new_A2062_;
  assign new_A2039_ = new_A2055_ | new_A2054_;
  assign new_A2038_ = new_A2061_ | new_A2060_;
  assign new_A2037_ = new_A2051_ | new_A2053_;
  assign new_A2036_ = ~new_A2058_ | ~new_A2059_;
  assign new_A2035_ = new_A2011_ & ~new_A2012_;
  assign new_A2034_ = new_A2025_ & ~new_A2037_;
  assign new_A2033_ = ~new_A2025_ & new_A2037_;
  assign new_A2032_ = ~new_A2023_ & new_A2049_;
  assign new_A2031_ = new_A2047_ | new_A2046_;
  assign new_A2030_ = new_A2044_ | new_A2043_;
  assign new_A2029_ = new_A2012_ | new_A2045_;
  assign new_A2028_ = new_A2037_ & new_A2040_;
  assign new_A2027_ = new_A2042_ | new_A2041_;
  assign new_A2026_ = new_A2037_ & new_A2036_;
  assign new_A2025_ = new_A2039_ & new_A2038_;
  assign new_A2024_ = new_A2034_ | new_A2033_;
  assign new_A2023_ = new_A2012_ | new_A2035_;
  assign A2022 = new_A2023_ | new_A2032_;
  assign A2021 = new_A2030_ & new_A2031_;
  assign A2020 = new_A2030_ & new_A2029_;
  assign A2019 = new_A2028_ | new_A2027_;
  assign A2018 = new_A2026_ | new_A2025_;
  assign A2017 = new_A2024_ & new_A2023_;
  assign new_A2016_ = new_A3561_;
  assign new_A2015_ = new_A3494_;
  assign new_A2014_ = new_A3427_;
  assign new_A2013_ = new_A3360_;
  assign new_A2012_ = new_A3293_;
  assign new_A2011_ = new_A3225_;
  assign new_A2010_ = ~new_A1949_ & new_A1963_;
  assign new_A2009_ = new_A1949_ & ~new_A1963_;
  assign new_A2008_ = new_A1949_ & ~new_A1963_;
  assign new_A2007_ = ~new_A1949_ & ~new_A1963_;
  assign new_A2006_ = new_A1949_ & new_A1963_;
  assign new_A2005_ = new_A2009_ | new_A2010_;
  assign new_A2004_ = ~new_A1949_ & new_A1963_;
  assign new_A2003_ = new_A2007_ | new_A2008_;
  assign new_A2002_ = ~new_A1978_ & ~new_A1998_;
  assign new_A2001_ = new_A1978_ & new_A1998_;
  assign new_A2000_ = ~new_A1945_ | ~new_A1970_;
  assign new_A1999_ = new_A1963_ & new_A2000_;
  assign new_A1998_ = new_A1946_ | new_A1947_;
  assign new_A1997_ = new_A1946_ | new_A1963_;
  assign new_A1996_ = ~new_A1963_ & ~new_A1999_;
  assign new_A1995_ = new_A1963_ | new_A2000_;
  assign new_A1994_ = new_A1946_ & ~new_A1947_;
  assign new_A1993_ = ~new_A1946_ & new_A1947_;
  assign new_A1992_ = new_A1956_ | new_A1989_;
  assign new_A1991_ = ~new_A1956_ & ~new_A1990_;
  assign new_A1990_ = new_A1956_ & new_A1989_;
  assign new_A1989_ = ~new_A1945_ | ~new_A1970_;
  assign new_A1988_ = ~new_A1946_ & new_A1956_;
  assign new_A1987_ = new_A1946_ & ~new_A1956_;
  assign new_A1986_ = new_A1948_ & new_A1985_;
  assign new_A1985_ = new_A2004_ | new_A2003_;
  assign new_A1984_ = ~new_A1948_ & new_A1983_;
  assign new_A1983_ = new_A2006_ | new_A2005_;
  assign new_A1982_ = new_A1948_ | new_A1981_;
  assign new_A1981_ = new_A2002_ | new_A2001_;
  assign new_A1980_ = ~new_A1960_ & ~new_A1970_;
  assign new_A1979_ = new_A1960_ & new_A1970_;
  assign new_A1978_ = ~new_A1960_ | new_A1970_;
  assign new_A1977_ = new_A1944_ & ~new_A1945_;
  assign new_A1976_ = ~new_A1944_ & new_A1945_;
  assign new_A1975_ = new_A1997_ & ~new_A1998_;
  assign new_A1974_ = ~new_A1997_ & new_A1998_;
  assign new_A1973_ = ~new_A1996_ | ~new_A1995_;
  assign new_A1972_ = new_A1988_ | new_A1987_;
  assign new_A1971_ = new_A1994_ | new_A1993_;
  assign new_A1970_ = new_A1984_ | new_A1986_;
  assign new_A1969_ = ~new_A1991_ | ~new_A1992_;
  assign new_A1968_ = new_A1944_ & ~new_A1945_;
  assign new_A1967_ = new_A1958_ & ~new_A1970_;
  assign new_A1966_ = ~new_A1958_ & new_A1970_;
  assign new_A1965_ = ~new_A1956_ & new_A1982_;
  assign new_A1964_ = new_A1980_ | new_A1979_;
  assign new_A1963_ = new_A1977_ | new_A1976_;
  assign new_A1962_ = new_A1945_ | new_A1978_;
  assign new_A1961_ = new_A1970_ & new_A1973_;
  assign new_A1960_ = new_A1975_ | new_A1974_;
  assign new_A1959_ = new_A1970_ & new_A1969_;
  assign new_A1958_ = new_A1972_ & new_A1971_;
  assign new_A1957_ = new_A1967_ | new_A1966_;
  assign new_A1956_ = new_A1945_ | new_A1968_;
  assign A1955 = new_A1956_ | new_A1965_;
  assign A1954 = new_A1963_ & new_A1964_;
  assign A1953 = new_A1963_ & new_A1962_;
  assign A1952 = new_A1961_ | new_A1960_;
  assign A1951 = new_A1959_ | new_A1958_;
  assign A1950 = new_A1957_ & new_A1956_;
  assign new_A1949_ = new_A5570_;
  assign new_A1948_ = new_A5503_;
  assign new_A1947_ = new_A5436_;
  assign new_A1946_ = new_A5369_;
  assign new_A1945_ = new_A5302_;
  assign new_A1944_ = new_A5235_;
  assign new_A1943_ = ~new_A1882_ & new_A1896_;
  assign new_A1942_ = new_A1882_ & ~new_A1896_;
  assign new_A1941_ = new_A1882_ & ~new_A1896_;
  assign new_A1940_ = ~new_A1882_ & ~new_A1896_;
  assign new_A1939_ = new_A1882_ & new_A1896_;
  assign new_A1938_ = new_A1942_ | new_A1943_;
  assign new_A1937_ = ~new_A1882_ & new_A1896_;
  assign new_A1936_ = new_A1940_ | new_A1941_;
  assign new_A1935_ = ~new_A1911_ & ~new_A1931_;
  assign new_A1934_ = new_A1911_ & new_A1931_;
  assign new_A1933_ = ~new_A1878_ | ~new_A1903_;
  assign new_A1932_ = new_A1896_ & new_A1933_;
  assign new_A1931_ = new_A1879_ | new_A1880_;
  assign new_A1930_ = new_A1879_ | new_A1896_;
  assign new_A1929_ = ~new_A1896_ & ~new_A1932_;
  assign new_A1928_ = new_A1896_ | new_A1933_;
  assign new_A1927_ = new_A1879_ & ~new_A1880_;
  assign new_A1926_ = ~new_A1879_ & new_A1880_;
  assign new_A1925_ = new_A1889_ | new_A1922_;
  assign new_A1924_ = ~new_A1889_ & ~new_A1923_;
  assign new_A1923_ = new_A1889_ & new_A1922_;
  assign new_A1922_ = ~new_A1878_ | ~new_A1903_;
  assign new_A1921_ = ~new_A1879_ & new_A1889_;
  assign new_A1920_ = new_A1879_ & ~new_A1889_;
  assign new_A1919_ = new_A1881_ & new_A1918_;
  assign new_A1918_ = new_A1937_ | new_A1936_;
  assign new_A1917_ = ~new_A1881_ & new_A1916_;
  assign new_A1916_ = new_A1939_ | new_A1938_;
  assign new_A1915_ = new_A1881_ | new_A1914_;
  assign new_A1914_ = new_A1935_ | new_A1934_;
  assign new_A1913_ = ~new_A1893_ & ~new_A1903_;
  assign new_A1912_ = new_A1893_ & new_A1903_;
  assign new_A1911_ = ~new_A1893_ | new_A1903_;
  assign new_A1910_ = new_A1877_ & ~new_A1878_;
  assign new_A1909_ = ~new_A1877_ & new_A1878_;
  assign new_A1908_ = new_A1930_ & ~new_A1931_;
  assign new_A1907_ = ~new_A1930_ & new_A1931_;
  assign new_A1906_ = ~new_A1929_ | ~new_A1928_;
  assign new_A1905_ = new_A1921_ | new_A1920_;
  assign new_A1904_ = new_A1927_ | new_A1926_;
  assign new_A1903_ = new_A1917_ | new_A1919_;
  assign new_A1902_ = ~new_A1924_ | ~new_A1925_;
  assign new_A1901_ = new_A1877_ & ~new_A1878_;
  assign new_A1900_ = new_A1891_ & ~new_A1903_;
  assign new_A1899_ = ~new_A1891_ & new_A1903_;
  assign new_A1898_ = ~new_A1889_ & new_A1915_;
  assign new_A1897_ = new_A1913_ | new_A1912_;
  assign new_A1896_ = new_A1910_ | new_A1909_;
  assign new_A1895_ = new_A1878_ | new_A1911_;
  assign new_A1894_ = new_A1903_ & new_A1906_;
  assign new_A1893_ = new_A1908_ | new_A1907_;
  assign new_A1892_ = new_A1903_ & new_A1902_;
  assign new_A1891_ = new_A1905_ & new_A1904_;
  assign new_A1890_ = new_A1900_ | new_A1899_;
  assign new_A1889_ = new_A1878_ | new_A1901_;
  assign A1888 = new_A1889_ | new_A1898_;
  assign A1887 = new_A1896_ & new_A1897_;
  assign A1886 = new_A1896_ & new_A1895_;
  assign A1885 = new_A1894_ | new_A1893_;
  assign A1884 = new_A1892_ | new_A1891_;
  assign A1883 = new_A1890_ & new_A1889_;
  assign new_A1882_ = new_A5168_;
  assign new_A1881_ = new_A5101_;
  assign new_A1880_ = new_A5034_;
  assign new_A1879_ = new_A4967_;
  assign new_A1878_ = new_A4900_;
  assign new_A1877_ = new_A4833_;
  assign new_A1876_ = ~new_A1815_ & new_A1829_;
  assign new_A1875_ = new_A1815_ & ~new_A1829_;
  assign new_A1874_ = new_A1815_ & ~new_A1829_;
  assign new_A1873_ = ~new_A1815_ & ~new_A1829_;
  assign new_A1872_ = new_A1815_ & new_A1829_;
  assign new_A1871_ = new_A1875_ | new_A1876_;
  assign new_A1870_ = ~new_A1815_ & new_A1829_;
  assign new_A1869_ = new_A1873_ | new_A1874_;
  assign new_A1868_ = ~new_A1844_ & ~new_A1864_;
  assign new_A1867_ = new_A1844_ & new_A1864_;
  assign new_A1866_ = ~new_A1811_ | ~new_A1836_;
  assign new_A1865_ = new_A1829_ & new_A1866_;
  assign new_A1864_ = new_A1812_ | new_A1813_;
  assign new_A1863_ = new_A1812_ | new_A1829_;
  assign new_A1862_ = ~new_A1829_ & ~new_A1865_;
  assign new_A1861_ = new_A1829_ | new_A1866_;
  assign new_A1860_ = new_A1812_ & ~new_A1813_;
  assign new_A1859_ = ~new_A1812_ & new_A1813_;
  assign new_A1858_ = new_A1822_ | new_A1855_;
  assign new_A1857_ = ~new_A1822_ & ~new_A1856_;
  assign new_A1856_ = new_A1822_ & new_A1855_;
  assign new_A1855_ = ~new_A1811_ | ~new_A1836_;
  assign new_A1854_ = ~new_A1812_ & new_A1822_;
  assign new_A1853_ = new_A1812_ & ~new_A1822_;
  assign new_A1852_ = new_A1814_ & new_A1851_;
  assign new_A1851_ = new_A1870_ | new_A1869_;
  assign new_A1850_ = ~new_A1814_ & new_A1849_;
  assign new_A1849_ = new_A1872_ | new_A1871_;
  assign new_A1848_ = new_A1814_ | new_A1847_;
  assign new_A1847_ = new_A1868_ | new_A1867_;
  assign new_A1846_ = ~new_A1826_ & ~new_A1836_;
  assign new_A1845_ = new_A1826_ & new_A1836_;
  assign new_A1844_ = ~new_A1826_ | new_A1836_;
  assign new_A1843_ = new_A1810_ & ~new_A1811_;
  assign new_A1842_ = ~new_A1810_ & new_A1811_;
  assign new_A1841_ = new_A1863_ & ~new_A1864_;
  assign new_A1840_ = ~new_A1863_ & new_A1864_;
  assign new_A1839_ = ~new_A1862_ | ~new_A1861_;
  assign new_A1838_ = new_A1854_ | new_A1853_;
  assign new_A1837_ = new_A1860_ | new_A1859_;
  assign new_A1836_ = new_A1850_ | new_A1852_;
  assign new_A1835_ = ~new_A1857_ | ~new_A1858_;
  assign new_A1834_ = new_A1810_ & ~new_A1811_;
  assign new_A1833_ = new_A1824_ & ~new_A1836_;
  assign new_A1832_ = ~new_A1824_ & new_A1836_;
  assign new_A1831_ = ~new_A1822_ & new_A1848_;
  assign new_A1830_ = new_A1846_ | new_A1845_;
  assign new_A1829_ = new_A1843_ | new_A1842_;
  assign new_A1828_ = new_A1811_ | new_A1844_;
  assign new_A1827_ = new_A1836_ & new_A1839_;
  assign new_A1826_ = new_A1841_ | new_A1840_;
  assign new_A1825_ = new_A1836_ & new_A1835_;
  assign new_A1824_ = new_A1838_ & new_A1837_;
  assign new_A1823_ = new_A1833_ | new_A1832_;
  assign new_A1822_ = new_A1811_ | new_A1834_;
  assign A1821 = new_A1822_ | new_A1831_;
  assign A1820 = new_A1829_ & new_A1830_;
  assign A1819 = new_A1829_ & new_A1828_;
  assign A1818 = new_A1827_ | new_A1826_;
  assign A1817 = new_A1825_ | new_A1824_;
  assign A1816 = new_A1823_ & new_A1822_;
  assign new_A1815_ = new_A4766_;
  assign new_A1814_ = new_A4699_;
  assign new_A1813_ = new_A4632_;
  assign new_A1812_ = new_A4565_;
  assign new_A1811_ = new_A4498_;
  assign new_A1810_ = new_A4431_;
  assign new_A1809_ = ~new_A1748_ & new_A1762_;
  assign new_A1808_ = new_A1748_ & ~new_A1762_;
  assign new_A1807_ = new_A1748_ & ~new_A1762_;
  assign new_A1806_ = ~new_A1748_ & ~new_A1762_;
  assign new_A1805_ = new_A1748_ & new_A1762_;
  assign new_A1804_ = new_A1808_ | new_A1809_;
  assign new_A1803_ = ~new_A1748_ & new_A1762_;
  assign new_A1802_ = new_A1806_ | new_A1807_;
  assign new_A1801_ = ~new_A1777_ & ~new_A1797_;
  assign new_A1800_ = new_A1777_ & new_A1797_;
  assign new_A1799_ = ~new_A1744_ | ~new_A1769_;
  assign new_A1798_ = new_A1762_ & new_A1799_;
  assign new_A1797_ = new_A1745_ | new_A1746_;
  assign new_A1796_ = new_A1745_ | new_A1762_;
  assign new_A1795_ = ~new_A1762_ & ~new_A1798_;
  assign new_A1794_ = new_A1762_ | new_A1799_;
  assign new_A1793_ = new_A1745_ & ~new_A1746_;
  assign new_A1792_ = ~new_A1745_ & new_A1746_;
  assign new_A1791_ = new_A1755_ | new_A1788_;
  assign new_A1790_ = ~new_A1755_ & ~new_A1789_;
  assign new_A1789_ = new_A1755_ & new_A1788_;
  assign new_A1788_ = ~new_A1744_ | ~new_A1769_;
  assign new_A1787_ = ~new_A1745_ & new_A1755_;
  assign new_A1786_ = new_A1745_ & ~new_A1755_;
  assign new_A1785_ = new_A1747_ & new_A1784_;
  assign new_A1784_ = new_A1803_ | new_A1802_;
  assign new_A1783_ = ~new_A1747_ & new_A1782_;
  assign new_A1782_ = new_A1805_ | new_A1804_;
  assign new_A1781_ = new_A1747_ | new_A1780_;
  assign new_A1780_ = new_A1801_ | new_A1800_;
  assign new_A1779_ = ~new_A1759_ & ~new_A1769_;
  assign new_A1778_ = new_A1759_ & new_A1769_;
  assign new_A1777_ = ~new_A1759_ | new_A1769_;
  assign new_A1776_ = new_A1743_ & ~new_A1744_;
  assign new_A1775_ = ~new_A1743_ & new_A1744_;
  assign new_A1774_ = new_A1796_ & ~new_A1797_;
  assign new_A1773_ = ~new_A1796_ & new_A1797_;
  assign new_A1772_ = ~new_A1795_ | ~new_A1794_;
  assign new_A1771_ = new_A1787_ | new_A1786_;
  assign new_A1770_ = new_A1793_ | new_A1792_;
  assign new_A1769_ = new_A1783_ | new_A1785_;
  assign new_A1768_ = ~new_A1790_ | ~new_A1791_;
  assign new_A1767_ = new_A1743_ & ~new_A1744_;
  assign new_A1766_ = new_A1757_ & ~new_A1769_;
  assign new_A1765_ = ~new_A1757_ & new_A1769_;
  assign new_A1764_ = ~new_A1755_ & new_A1781_;
  assign new_A1763_ = new_A1779_ | new_A1778_;
  assign new_A1762_ = new_A1776_ | new_A1775_;
  assign new_A1761_ = new_A1744_ | new_A1777_;
  assign new_A1760_ = new_A1769_ & new_A1772_;
  assign new_A1759_ = new_A1774_ | new_A1773_;
  assign new_A1758_ = new_A1769_ & new_A1768_;
  assign new_A1757_ = new_A1771_ & new_A1770_;
  assign new_A1756_ = new_A1766_ | new_A1765_;
  assign new_A1755_ = new_A1744_ | new_A1767_;
  assign A1754 = new_A1755_ | new_A1764_;
  assign A1753 = new_A1762_ & new_A1763_;
  assign A1752 = new_A1762_ & new_A1761_;
  assign A1751 = new_A1760_ | new_A1759_;
  assign A1750 = new_A1758_ | new_A1757_;
  assign A1749 = new_A1756_ & new_A1755_;
  assign new_A1748_ = new_A4364_;
  assign new_A1747_ = new_A4297_;
  assign new_A1746_ = new_A4230_;
  assign new_A1745_ = new_A4163_;
  assign new_A1744_ = new_A4096_;
  assign new_A1743_ = new_A4029_;
  assign new_A1742_ = ~new_A1681_ & new_A1695_;
  assign new_A1741_ = new_A1681_ & ~new_A1695_;
  assign new_A1740_ = new_A1681_ & ~new_A1695_;
  assign new_A1739_ = ~new_A1681_ & ~new_A1695_;
  assign new_A1738_ = new_A1681_ & new_A1695_;
  assign new_A1737_ = new_A1741_ | new_A1742_;
  assign new_A1736_ = ~new_A1681_ & new_A1695_;
  assign new_A1735_ = new_A1739_ | new_A1740_;
  assign new_A1734_ = ~new_A1710_ & ~new_A1730_;
  assign new_A1733_ = new_A1710_ & new_A1730_;
  assign new_A1732_ = ~new_A1677_ | ~new_A1702_;
  assign new_A1731_ = new_A1695_ & new_A1732_;
  assign new_A1730_ = new_A1678_ | new_A1679_;
  assign new_A1729_ = new_A1678_ | new_A1695_;
  assign new_A1728_ = ~new_A1695_ & ~new_A1731_;
  assign new_A1727_ = new_A1695_ | new_A1732_;
  assign new_A1726_ = new_A1678_ & ~new_A1679_;
  assign new_A1725_ = ~new_A1678_ & new_A1679_;
  assign new_A1724_ = new_A1688_ | new_A1721_;
  assign new_A1723_ = ~new_A1688_ & ~new_A1722_;
  assign new_A1722_ = new_A1688_ & new_A1721_;
  assign new_A1721_ = ~new_A1677_ | ~new_A1702_;
  assign new_A1720_ = ~new_A1678_ & new_A1688_;
  assign new_A1719_ = new_A1678_ & ~new_A1688_;
  assign new_A1718_ = new_A1680_ & new_A1717_;
  assign new_A1717_ = new_A1736_ | new_A1735_;
  assign new_A1716_ = ~new_A1680_ & new_A1715_;
  assign new_A1715_ = new_A1738_ | new_A1737_;
  assign new_A1714_ = new_A1680_ | new_A1713_;
  assign new_A1713_ = new_A1734_ | new_A1733_;
  assign new_A1712_ = ~new_A1692_ & ~new_A1702_;
  assign new_A1711_ = new_A1692_ & new_A1702_;
  assign new_A1710_ = ~new_A1692_ | new_A1702_;
  assign new_A1709_ = new_A1676_ & ~new_A1677_;
  assign new_A1708_ = ~new_A1676_ & new_A1677_;
  assign new_A1707_ = new_A1729_ & ~new_A1730_;
  assign new_A1706_ = ~new_A1729_ & new_A1730_;
  assign new_A1705_ = ~new_A1728_ | ~new_A1727_;
  assign new_A1704_ = new_A1720_ | new_A1719_;
  assign new_A1703_ = new_A1726_ | new_A1725_;
  assign new_A1702_ = new_A1716_ | new_A1718_;
  assign new_A1701_ = ~new_A1723_ | ~new_A1724_;
  assign new_A1700_ = new_A1676_ & ~new_A1677_;
  assign new_A1699_ = new_A1690_ & ~new_A1702_;
  assign new_A1698_ = ~new_A1690_ & new_A1702_;
  assign new_A1697_ = ~new_A1688_ & new_A1714_;
  assign new_A1696_ = new_A1712_ | new_A1711_;
  assign new_A1695_ = new_A1709_ | new_A1708_;
  assign new_A1694_ = new_A1677_ | new_A1710_;
  assign new_A1693_ = new_A1702_ & new_A1705_;
  assign new_A1692_ = new_A1707_ | new_A1706_;
  assign new_A1691_ = new_A1702_ & new_A1701_;
  assign new_A1690_ = new_A1704_ & new_A1703_;
  assign new_A1689_ = new_A1699_ | new_A1698_;
  assign new_A1688_ = new_A1677_ | new_A1700_;
  assign A1687 = new_A1688_ | new_A1697_;
  assign A1686 = new_A1695_ & new_A1696_;
  assign A1685 = new_A1695_ & new_A1694_;
  assign A1684 = new_A1693_ | new_A1692_;
  assign A1683 = new_A1691_ | new_A1690_;
  assign A1682 = new_A1689_ & new_A1688_;
  assign new_A1681_ = new_A3962_;
  assign new_A1680_ = new_A3895_;
  assign new_A1679_ = new_A3828_;
  assign new_A1678_ = new_A3761_;
  assign new_A1677_ = new_A3694_;
  assign new_A1676_ = new_A3627_;
  assign new_A1675_ = ~new_A1614_ & new_A1628_;
  assign new_A1674_ = new_A1614_ & ~new_A1628_;
  assign new_A1673_ = new_A1614_ & ~new_A1628_;
  assign new_A1672_ = ~new_A1614_ & ~new_A1628_;
  assign new_A1671_ = new_A1614_ & new_A1628_;
  assign new_A1670_ = new_A1674_ | new_A1675_;
  assign new_A1669_ = ~new_A1614_ & new_A1628_;
  assign new_A1668_ = new_A1672_ | new_A1673_;
  assign new_A1667_ = ~new_A1643_ & ~new_A1663_;
  assign new_A1666_ = new_A1643_ & new_A1663_;
  assign new_A1665_ = ~new_A1610_ | ~new_A1635_;
  assign new_A1664_ = new_A1628_ & new_A1665_;
  assign new_A1663_ = new_A1611_ | new_A1612_;
  assign new_A1662_ = new_A1611_ | new_A1628_;
  assign new_A1661_ = ~new_A1628_ & ~new_A1664_;
  assign new_A1660_ = new_A1628_ | new_A1665_;
  assign new_A1659_ = new_A1611_ & ~new_A1612_;
  assign new_A1658_ = ~new_A1611_ & new_A1612_;
  assign new_A1657_ = new_A1621_ | new_A1654_;
  assign new_A1656_ = ~new_A1621_ & ~new_A1655_;
  assign new_A1655_ = new_A1621_ & new_A1654_;
  assign new_A1654_ = ~new_A1610_ | ~new_A1635_;
  assign new_A1653_ = ~new_A1611_ & new_A1621_;
  assign new_A1652_ = new_A1611_ & ~new_A1621_;
  assign new_A1651_ = new_A1613_ & new_A1650_;
  assign new_A1650_ = new_A1669_ | new_A1668_;
  assign new_A1649_ = ~new_A1613_ & new_A1648_;
  assign new_A1648_ = new_A1671_ | new_A1670_;
  assign new_A1647_ = new_A1613_ | new_A1646_;
  assign new_A1646_ = new_A1667_ | new_A1666_;
  assign new_A1645_ = ~new_A1625_ & ~new_A1635_;
  assign new_A1644_ = new_A1625_ & new_A1635_;
  assign new_A1643_ = ~new_A1625_ | new_A1635_;
  assign new_A1642_ = new_A1609_ & ~new_A1610_;
  assign new_A1641_ = ~new_A1609_ & new_A1610_;
  assign new_A1640_ = new_A1662_ & ~new_A1663_;
  assign new_A1639_ = ~new_A1662_ & new_A1663_;
  assign new_A1638_ = ~new_A1661_ | ~new_A1660_;
  assign new_A1637_ = new_A1653_ | new_A1652_;
  assign new_A1636_ = new_A1659_ | new_A1658_;
  assign new_A1635_ = new_A1649_ | new_A1651_;
  assign new_A1634_ = ~new_A1656_ | ~new_A1657_;
  assign new_A1633_ = new_A1609_ & ~new_A1610_;
  assign new_A1632_ = new_A1623_ & ~new_A1635_;
  assign new_A1631_ = ~new_A1623_ & new_A1635_;
  assign new_A1630_ = ~new_A1621_ & new_A1647_;
  assign new_A1629_ = new_A1645_ | new_A1644_;
  assign new_A1628_ = new_A1642_ | new_A1641_;
  assign new_A1627_ = new_A1610_ | new_A1643_;
  assign new_A1626_ = new_A1635_ & new_A1638_;
  assign new_A1625_ = new_A1640_ | new_A1639_;
  assign new_A1624_ = new_A1635_ & new_A1634_;
  assign new_A1623_ = new_A1637_ & new_A1636_;
  assign new_A1622_ = new_A1632_ | new_A1631_;
  assign new_A1621_ = new_A1610_ | new_A1633_;
  assign A1620 = new_A1621_ | new_A1630_;
  assign A1619 = new_A1628_ & new_A1629_;
  assign A1618 = new_A1628_ & new_A1627_;
  assign A1617 = new_A1626_ | new_A1625_;
  assign A1616 = new_A1624_ | new_A1623_;
  assign A1615 = new_A1622_ & new_A1621_;
  assign new_A1614_ = new_A3560_;
  assign new_A1613_ = new_A3493_;
  assign new_A1612_ = new_A3426_;
  assign new_A1611_ = new_A3359_;
  assign new_A1610_ = new_A3292_;
  assign new_A1609_ = new_A3226_;
  assign new_A1608_ = ~new_A1547_ & new_A1561_;
  assign new_A1607_ = new_A1547_ & ~new_A1561_;
  assign new_A1606_ = new_A1547_ & ~new_A1561_;
  assign new_A1605_ = ~new_A1547_ & ~new_A1561_;
  assign new_A1604_ = new_A1547_ & new_A1561_;
  assign new_A1603_ = new_A1607_ | new_A1608_;
  assign new_A1602_ = ~new_A1547_ & new_A1561_;
  assign new_A1601_ = new_A1605_ | new_A1606_;
  assign new_A1600_ = ~new_A1576_ & ~new_A1596_;
  assign new_A1599_ = new_A1576_ & new_A1596_;
  assign new_A1598_ = ~new_A1543_ | ~new_A1568_;
  assign new_A1597_ = new_A1561_ & new_A1598_;
  assign new_A1596_ = new_A1544_ | new_A1545_;
  assign new_A1595_ = new_A1544_ | new_A1561_;
  assign new_A1594_ = ~new_A1561_ & ~new_A1597_;
  assign new_A1593_ = new_A1561_ | new_A1598_;
  assign new_A1592_ = new_A1544_ & ~new_A1545_;
  assign new_A1591_ = ~new_A1544_ & new_A1545_;
  assign new_A1590_ = new_A1554_ | new_A1587_;
  assign new_A1589_ = ~new_A1554_ & ~new_A1588_;
  assign new_A1588_ = new_A1554_ & new_A1587_;
  assign new_A1587_ = ~new_A1543_ | ~new_A1568_;
  assign new_A1586_ = ~new_A1544_ & new_A1554_;
  assign new_A1585_ = new_A1544_ & ~new_A1554_;
  assign new_A1584_ = new_A1546_ & new_A1583_;
  assign new_A1583_ = new_A1602_ | new_A1601_;
  assign new_A1582_ = ~new_A1546_ & new_A1581_;
  assign new_A1581_ = new_A1604_ | new_A1603_;
  assign new_A1580_ = new_A1546_ | new_A1579_;
  assign new_A1579_ = new_A1600_ | new_A1599_;
  assign new_A1578_ = ~new_A1558_ & ~new_A1568_;
  assign new_A1577_ = new_A1558_ & new_A1568_;
  assign new_A1576_ = ~new_A1558_ | new_A1568_;
  assign new_A1575_ = new_A1542_ & ~new_A1543_;
  assign new_A1574_ = ~new_A1542_ & new_A1543_;
  assign new_A1573_ = new_A1595_ & ~new_A1596_;
  assign new_A1572_ = ~new_A1595_ & new_A1596_;
  assign new_A1571_ = ~new_A1594_ | ~new_A1593_;
  assign new_A1570_ = new_A1586_ | new_A1585_;
  assign new_A1569_ = new_A1592_ | new_A1591_;
  assign new_A1568_ = new_A1582_ | new_A1584_;
  assign new_A1567_ = ~new_A1589_ | ~new_A1590_;
  assign new_A1566_ = new_A1542_ & ~new_A1543_;
  assign new_A1565_ = new_A1556_ & ~new_A1568_;
  assign new_A1564_ = ~new_A1556_ & new_A1568_;
  assign new_A1563_ = ~new_A1554_ & new_A1580_;
  assign new_A1562_ = new_A1578_ | new_A1577_;
  assign new_A1561_ = new_A1575_ | new_A1574_;
  assign new_A1560_ = new_A1543_ | new_A1576_;
  assign new_A1559_ = new_A1568_ & new_A1571_;
  assign new_A1558_ = new_A1573_ | new_A1572_;
  assign new_A1557_ = new_A1568_ & new_A1567_;
  assign new_A1556_ = new_A1570_ & new_A1569_;
  assign new_A1555_ = new_A1565_ | new_A1564_;
  assign new_A1554_ = new_A1543_ | new_A1566_;
  assign A1553 = new_A1554_ | new_A1563_;
  assign A1552 = new_A1561_ & new_A1562_;
  assign A1551 = new_A1561_ & new_A1560_;
  assign A1550 = new_A1559_ | new_A1558_;
  assign A1549 = new_A1557_ | new_A1556_;
  assign A1548 = new_A1555_ & new_A1554_;
  assign new_A1547_ = new_A5569_;
  assign new_A1546_ = new_A5502_;
  assign new_A1545_ = new_A5435_;
  assign new_A1544_ = new_A5368_;
  assign new_A1543_ = new_A5301_;
  assign new_A1542_ = new_A5234_;
  assign new_A1541_ = ~new_A1480_ & new_A1494_;
  assign new_A1540_ = new_A1480_ & ~new_A1494_;
  assign new_A1539_ = new_A1480_ & ~new_A1494_;
  assign new_A1538_ = ~new_A1480_ & ~new_A1494_;
  assign new_A1537_ = new_A1480_ & new_A1494_;
  assign new_A1536_ = new_A1540_ | new_A1541_;
  assign new_A1535_ = ~new_A1480_ & new_A1494_;
  assign new_A1534_ = new_A1538_ | new_A1539_;
  assign new_A1533_ = ~new_A1509_ & ~new_A1529_;
  assign new_A1532_ = new_A1509_ & new_A1529_;
  assign new_A1531_ = ~new_A1476_ | ~new_A1501_;
  assign new_A1530_ = new_A1494_ & new_A1531_;
  assign new_A1529_ = new_A1477_ | new_A1478_;
  assign new_A1528_ = new_A1477_ | new_A1494_;
  assign new_A1527_ = ~new_A1494_ & ~new_A1530_;
  assign new_A1526_ = new_A1494_ | new_A1531_;
  assign new_A1525_ = new_A1477_ & ~new_A1478_;
  assign new_A1524_ = ~new_A1477_ & new_A1478_;
  assign new_A1523_ = new_A1487_ | new_A1520_;
  assign new_A1522_ = ~new_A1487_ & ~new_A1521_;
  assign new_A1521_ = new_A1487_ & new_A1520_;
  assign new_A1520_ = ~new_A1476_ | ~new_A1501_;
  assign new_A1519_ = ~new_A1477_ & new_A1487_;
  assign new_A1518_ = new_A1477_ & ~new_A1487_;
  assign new_A1517_ = new_A1479_ & new_A1516_;
  assign new_A1516_ = new_A1535_ | new_A1534_;
  assign new_A1515_ = ~new_A1479_ & new_A1514_;
  assign new_A1514_ = new_A1537_ | new_A1536_;
  assign new_A1513_ = new_A1479_ | new_A1512_;
  assign new_A1512_ = new_A1533_ | new_A1532_;
  assign new_A1511_ = ~new_A1491_ & ~new_A1501_;
  assign new_A1510_ = new_A1491_ & new_A1501_;
  assign new_A1509_ = ~new_A1491_ | new_A1501_;
  assign new_A1508_ = new_A1475_ & ~new_A1476_;
  assign new_A1507_ = ~new_A1475_ & new_A1476_;
  assign new_A1506_ = new_A1528_ & ~new_A1529_;
  assign new_A1505_ = ~new_A1528_ & new_A1529_;
  assign new_A1504_ = ~new_A1527_ | ~new_A1526_;
  assign new_A1503_ = new_A1519_ | new_A1518_;
  assign new_A1502_ = new_A1525_ | new_A1524_;
  assign new_A1501_ = new_A1515_ | new_A1517_;
  assign new_A1500_ = ~new_A1522_ | ~new_A1523_;
  assign new_A1499_ = new_A1475_ & ~new_A1476_;
  assign new_A1498_ = new_A1489_ & ~new_A1501_;
  assign new_A1497_ = ~new_A1489_ & new_A1501_;
  assign new_A1496_ = ~new_A1487_ & new_A1513_;
  assign new_A1495_ = new_A1511_ | new_A1510_;
  assign new_A1494_ = new_A1508_ | new_A1507_;
  assign new_A1493_ = new_A1476_ | new_A1509_;
  assign new_A1492_ = new_A1501_ & new_A1504_;
  assign new_A1491_ = new_A1506_ | new_A1505_;
  assign new_A1490_ = new_A1501_ & new_A1500_;
  assign new_A1489_ = new_A1503_ & new_A1502_;
  assign new_A1488_ = new_A1498_ | new_A1497_;
  assign new_A1487_ = new_A1476_ | new_A1499_;
  assign A1486 = new_A1487_ | new_A1496_;
  assign A1485 = new_A1494_ & new_A1495_;
  assign A1484 = new_A1494_ & new_A1493_;
  assign A1483 = new_A1492_ | new_A1491_;
  assign A1482 = new_A1490_ | new_A1489_;
  assign A1481 = new_A1488_ & new_A1487_;
  assign new_A1480_ = new_A5167_;
  assign new_A1479_ = new_A5100_;
  assign new_A1478_ = new_A5033_;
  assign new_A1477_ = new_A4966_;
  assign new_A1476_ = new_A4899_;
  assign new_A1475_ = new_A4832_;
  assign new_A1474_ = ~new_A1413_ & new_A1427_;
  assign new_A1473_ = new_A1413_ & ~new_A1427_;
  assign new_A1472_ = new_A1413_ & ~new_A1427_;
  assign new_A1471_ = ~new_A1413_ & ~new_A1427_;
  assign new_A1470_ = new_A1413_ & new_A1427_;
  assign new_A1469_ = new_A1473_ | new_A1474_;
  assign new_A1468_ = ~new_A1413_ & new_A1427_;
  assign new_A1467_ = new_A1471_ | new_A1472_;
  assign new_A1466_ = ~new_A1442_ & ~new_A1462_;
  assign new_A1465_ = new_A1442_ & new_A1462_;
  assign new_A1464_ = ~new_A1409_ | ~new_A1434_;
  assign new_A1463_ = new_A1427_ & new_A1464_;
  assign new_A1462_ = new_A1410_ | new_A1411_;
  assign new_A1461_ = new_A1410_ | new_A1427_;
  assign new_A1460_ = ~new_A1427_ & ~new_A1463_;
  assign new_A1459_ = new_A1427_ | new_A1464_;
  assign new_A1458_ = new_A1410_ & ~new_A1411_;
  assign new_A1457_ = ~new_A1410_ & new_A1411_;
  assign new_A1456_ = new_A1420_ | new_A1453_;
  assign new_A1455_ = ~new_A1420_ & ~new_A1454_;
  assign new_A1454_ = new_A1420_ & new_A1453_;
  assign new_A1453_ = ~new_A1409_ | ~new_A1434_;
  assign new_A1452_ = ~new_A1410_ & new_A1420_;
  assign new_A1451_ = new_A1410_ & ~new_A1420_;
  assign new_A1450_ = new_A1412_ & new_A1449_;
  assign new_A1449_ = new_A1468_ | new_A1467_;
  assign new_A1448_ = ~new_A1412_ & new_A1447_;
  assign new_A1447_ = new_A1470_ | new_A1469_;
  assign new_A1446_ = new_A1412_ | new_A1445_;
  assign new_A1445_ = new_A1466_ | new_A1465_;
  assign new_A1444_ = ~new_A1424_ & ~new_A1434_;
  assign new_A1443_ = new_A1424_ & new_A1434_;
  assign new_A1442_ = ~new_A1424_ | new_A1434_;
  assign new_A1441_ = new_A1408_ & ~new_A1409_;
  assign new_A1440_ = ~new_A1408_ & new_A1409_;
  assign new_A1439_ = new_A1461_ & ~new_A1462_;
  assign new_A1438_ = ~new_A1461_ & new_A1462_;
  assign new_A1437_ = ~new_A1460_ | ~new_A1459_;
  assign new_A1436_ = new_A1452_ | new_A1451_;
  assign new_A1435_ = new_A1458_ | new_A1457_;
  assign new_A1434_ = new_A1448_ | new_A1450_;
  assign new_A1433_ = ~new_A1455_ | ~new_A1456_;
  assign new_A1432_ = new_A1408_ & ~new_A1409_;
  assign new_A1431_ = new_A1422_ & ~new_A1434_;
  assign new_A1430_ = ~new_A1422_ & new_A1434_;
  assign new_A1429_ = ~new_A1420_ & new_A1446_;
  assign new_A1428_ = new_A1444_ | new_A1443_;
  assign new_A1427_ = new_A1441_ | new_A1440_;
  assign new_A1426_ = new_A1409_ | new_A1442_;
  assign new_A1425_ = new_A1434_ & new_A1437_;
  assign new_A1424_ = new_A1439_ | new_A1438_;
  assign new_A1423_ = new_A1434_ & new_A1433_;
  assign new_A1422_ = new_A1436_ & new_A1435_;
  assign new_A1421_ = new_A1431_ | new_A1430_;
  assign new_A1420_ = new_A1409_ | new_A1432_;
  assign A1419 = new_A1420_ | new_A1429_;
  assign A1418 = new_A1427_ & new_A1428_;
  assign A1417 = new_A1427_ & new_A1426_;
  assign A1416 = new_A1425_ | new_A1424_;
  assign A1415 = new_A1423_ | new_A1422_;
  assign A1414 = new_A1421_ & new_A1420_;
  assign new_A1413_ = new_A4765_;
  assign new_A1412_ = new_A4698_;
  assign new_A1411_ = new_A4631_;
  assign new_A1410_ = new_A4564_;
  assign new_A1409_ = new_A4497_;
  assign new_A1408_ = new_A4430_;
  assign new_A1407_ = ~new_A1346_ & new_A1360_;
  assign new_A1406_ = new_A1346_ & ~new_A1360_;
  assign new_A1405_ = new_A1346_ & ~new_A1360_;
  assign new_A1404_ = ~new_A1346_ & ~new_A1360_;
  assign new_A1403_ = new_A1346_ & new_A1360_;
  assign new_A1402_ = new_A1406_ | new_A1407_;
  assign new_A1401_ = ~new_A1346_ & new_A1360_;
  assign new_A1400_ = new_A1404_ | new_A1405_;
  assign new_A1399_ = ~new_A1375_ & ~new_A1395_;
  assign new_A1398_ = new_A1375_ & new_A1395_;
  assign new_A1397_ = ~new_A1342_ | ~new_A1367_;
  assign new_A1396_ = new_A1360_ & new_A1397_;
  assign new_A1395_ = new_A1343_ | new_A1344_;
  assign new_A1394_ = new_A1343_ | new_A1360_;
  assign new_A1393_ = ~new_A1360_ & ~new_A1396_;
  assign new_A1392_ = new_A1360_ | new_A1397_;
  assign new_A1391_ = new_A1343_ & ~new_A1344_;
  assign new_A1390_ = ~new_A1343_ & new_A1344_;
  assign new_A1389_ = new_A1353_ | new_A1386_;
  assign new_A1388_ = ~new_A1353_ & ~new_A1387_;
  assign new_A1387_ = new_A1353_ & new_A1386_;
  assign new_A1386_ = ~new_A1342_ | ~new_A1367_;
  assign new_A1385_ = ~new_A1343_ & new_A1353_;
  assign new_A1384_ = new_A1343_ & ~new_A1353_;
  assign new_A1383_ = new_A1345_ & new_A1382_;
  assign new_A1382_ = new_A1401_ | new_A1400_;
  assign new_A1381_ = ~new_A1345_ & new_A1380_;
  assign new_A1380_ = new_A1403_ | new_A1402_;
  assign new_A1379_ = new_A1345_ | new_A1378_;
  assign new_A1378_ = new_A1399_ | new_A1398_;
  assign new_A1377_ = ~new_A1357_ & ~new_A1367_;
  assign new_A1376_ = new_A1357_ & new_A1367_;
  assign new_A1375_ = ~new_A1357_ | new_A1367_;
  assign new_A1374_ = new_A1341_ & ~new_A1342_;
  assign new_A1373_ = ~new_A1341_ & new_A1342_;
  assign new_A1372_ = new_A1394_ & ~new_A1395_;
  assign new_A1371_ = ~new_A1394_ & new_A1395_;
  assign new_A1370_ = ~new_A1393_ | ~new_A1392_;
  assign new_A1369_ = new_A1385_ | new_A1384_;
  assign new_A1368_ = new_A1391_ | new_A1390_;
  assign new_A1367_ = new_A1381_ | new_A1383_;
  assign new_A1366_ = ~new_A1388_ | ~new_A1389_;
  assign new_A1365_ = new_A1341_ & ~new_A1342_;
  assign new_A1364_ = new_A1355_ & ~new_A1367_;
  assign new_A1363_ = ~new_A1355_ & new_A1367_;
  assign new_A1362_ = ~new_A1353_ & new_A1379_;
  assign new_A1361_ = new_A1377_ | new_A1376_;
  assign new_A1360_ = new_A1374_ | new_A1373_;
  assign new_A1359_ = new_A1342_ | new_A1375_;
  assign new_A1358_ = new_A1367_ & new_A1370_;
  assign new_A1357_ = new_A1372_ | new_A1371_;
  assign new_A1356_ = new_A1367_ & new_A1366_;
  assign new_A1355_ = new_A1369_ & new_A1368_;
  assign new_A1354_ = new_A1364_ | new_A1363_;
  assign new_A1353_ = new_A1342_ | new_A1365_;
  assign A1352 = new_A1353_ | new_A1362_;
  assign A1351 = new_A1360_ & new_A1361_;
  assign A1350 = new_A1360_ & new_A1359_;
  assign A1349 = new_A1358_ | new_A1357_;
  assign A1348 = new_A1356_ | new_A1355_;
  assign A1347 = new_A1354_ & new_A1353_;
  assign new_A1346_ = new_A4363_;
  assign new_A1345_ = new_A4296_;
  assign new_A1344_ = new_A4229_;
  assign new_A1343_ = new_A4162_;
  assign new_A1342_ = new_A4095_;
  assign new_A1341_ = new_A4028_;
  assign new_A1340_ = ~new_A1279_ & new_A1293_;
  assign new_A1339_ = new_A1279_ & ~new_A1293_;
  assign new_A1338_ = new_A1279_ & ~new_A1293_;
  assign new_A1337_ = ~new_A1279_ & ~new_A1293_;
  assign new_A1336_ = new_A1279_ & new_A1293_;
  assign new_A1335_ = new_A1339_ | new_A1340_;
  assign new_A1334_ = ~new_A1279_ & new_A1293_;
  assign new_A1333_ = new_A1337_ | new_A1338_;
  assign new_A1332_ = ~new_A1308_ & ~new_A1328_;
  assign new_A1331_ = new_A1308_ & new_A1328_;
  assign new_A1330_ = ~new_A1275_ | ~new_A1300_;
  assign new_A1329_ = new_A1293_ & new_A1330_;
  assign new_A1328_ = new_A1276_ | new_A1277_;
  assign new_A1327_ = new_A1276_ | new_A1293_;
  assign new_A1326_ = ~new_A1293_ & ~new_A1329_;
  assign new_A1325_ = new_A1293_ | new_A1330_;
  assign new_A1324_ = new_A1276_ & ~new_A1277_;
  assign new_A1323_ = ~new_A1276_ & new_A1277_;
  assign new_A1322_ = new_A1286_ | new_A1319_;
  assign new_A1321_ = ~new_A1286_ & ~new_A1320_;
  assign new_A1320_ = new_A1286_ & new_A1319_;
  assign new_A1319_ = ~new_A1275_ | ~new_A1300_;
  assign new_A1318_ = ~new_A1276_ & new_A1286_;
  assign new_A1317_ = new_A1276_ & ~new_A1286_;
  assign new_A1316_ = new_A1278_ & new_A1315_;
  assign new_A1315_ = new_A1334_ | new_A1333_;
  assign new_A1314_ = ~new_A1278_ & new_A1313_;
  assign new_A1313_ = new_A1336_ | new_A1335_;
  assign new_A1312_ = new_A1278_ | new_A1311_;
  assign new_A1311_ = new_A1332_ | new_A1331_;
  assign new_A1310_ = ~new_A1290_ & ~new_A1300_;
  assign new_A1309_ = new_A1290_ & new_A1300_;
  assign new_A1308_ = ~new_A1290_ | new_A1300_;
  assign new_A1307_ = new_A1274_ & ~new_A1275_;
  assign new_A1306_ = ~new_A1274_ & new_A1275_;
  assign new_A1305_ = new_A1327_ & ~new_A1328_;
  assign new_A1304_ = ~new_A1327_ & new_A1328_;
  assign new_A1303_ = ~new_A1326_ | ~new_A1325_;
  assign new_A1302_ = new_A1318_ | new_A1317_;
  assign new_A1301_ = new_A1324_ | new_A1323_;
  assign new_A1300_ = new_A1314_ | new_A1316_;
  assign new_A1299_ = ~new_A1321_ | ~new_A1322_;
  assign new_A1298_ = new_A1274_ & ~new_A1275_;
  assign new_A1297_ = new_A1288_ & ~new_A1300_;
  assign new_A1296_ = ~new_A1288_ & new_A1300_;
  assign new_A1295_ = ~new_A1286_ & new_A1312_;
  assign new_A1294_ = new_A1310_ | new_A1309_;
  assign new_A1293_ = new_A1307_ | new_A1306_;
  assign new_A1292_ = new_A1275_ | new_A1308_;
  assign new_A1291_ = new_A1300_ & new_A1303_;
  assign new_A1290_ = new_A1305_ | new_A1304_;
  assign new_A1289_ = new_A1300_ & new_A1299_;
  assign new_A1288_ = new_A1302_ & new_A1301_;
  assign new_A1287_ = new_A1297_ | new_A1296_;
  assign new_A1286_ = new_A1275_ | new_A1298_;
  assign A1285 = new_A1286_ | new_A1295_;
  assign A1284 = new_A1293_ & new_A1294_;
  assign A1283 = new_A1293_ & new_A1292_;
  assign A1282 = new_A1291_ | new_A1290_;
  assign A1281 = new_A1289_ | new_A1288_;
  assign A1280 = new_A1287_ & new_A1286_;
  assign new_A1279_ = new_A3961_;
  assign new_A1278_ = new_A3894_;
  assign new_A1277_ = new_A3827_;
  assign new_A1276_ = new_A3760_;
  assign new_A1275_ = new_A3693_;
  assign new_A1274_ = new_A3626_;
  assign new_A1273_ = ~new_A1212_ & new_A1226_;
  assign new_A1272_ = new_A1212_ & ~new_A1226_;
  assign new_A1271_ = new_A1212_ & ~new_A1226_;
  assign new_A1270_ = ~new_A1212_ & ~new_A1226_;
  assign new_A1269_ = new_A1212_ & new_A1226_;
  assign new_A1268_ = new_A1272_ | new_A1273_;
  assign new_A1267_ = ~new_A1212_ & new_A1226_;
  assign new_A1266_ = new_A1270_ | new_A1271_;
  assign new_A1265_ = ~new_A1241_ & ~new_A1261_;
  assign new_A1264_ = new_A1241_ & new_A1261_;
  assign new_A1263_ = ~new_A1208_ | ~new_A1233_;
  assign new_A1262_ = new_A1226_ & new_A1263_;
  assign new_A1261_ = new_A1209_ | new_A1210_;
  assign new_A1260_ = new_A1209_ | new_A1226_;
  assign new_A1259_ = ~new_A1226_ & ~new_A1262_;
  assign new_A1258_ = new_A1226_ | new_A1263_;
  assign new_A1257_ = new_A1209_ & ~new_A1210_;
  assign new_A1256_ = ~new_A1209_ & new_A1210_;
  assign new_A1255_ = new_A1219_ | new_A1252_;
  assign new_A1254_ = ~new_A1219_ & ~new_A1253_;
  assign new_A1253_ = new_A1219_ & new_A1252_;
  assign new_A1252_ = ~new_A1208_ | ~new_A1233_;
  assign new_A1251_ = ~new_A1209_ & new_A1219_;
  assign new_A1250_ = new_A1209_ & ~new_A1219_;
  assign new_A1249_ = new_A1211_ & new_A1248_;
  assign new_A1248_ = new_A1267_ | new_A1266_;
  assign new_A1247_ = ~new_A1211_ & new_A1246_;
  assign new_A1246_ = new_A1269_ | new_A1268_;
  assign new_A1245_ = new_A1211_ | new_A1244_;
  assign new_A1244_ = new_A1265_ | new_A1264_;
  assign new_A1243_ = ~new_A1223_ & ~new_A1233_;
  assign new_A1242_ = new_A1223_ & new_A1233_;
  assign new_A1241_ = ~new_A1223_ | new_A1233_;
  assign new_A1240_ = new_A1207_ & ~new_A1208_;
  assign new_A1239_ = ~new_A1207_ & new_A1208_;
  assign new_A1238_ = new_A1260_ & ~new_A1261_;
  assign new_A1237_ = ~new_A1260_ & new_A1261_;
  assign new_A1236_ = ~new_A1259_ | ~new_A1258_;
  assign new_A1235_ = new_A1251_ | new_A1250_;
  assign new_A1234_ = new_A1257_ | new_A1256_;
  assign new_A1233_ = new_A1247_ | new_A1249_;
  assign new_A1232_ = ~new_A1254_ | ~new_A1255_;
  assign new_A1231_ = new_A1207_ & ~new_A1208_;
  assign new_A1230_ = new_A1221_ & ~new_A1233_;
  assign new_A1229_ = ~new_A1221_ & new_A1233_;
  assign new_A1228_ = ~new_A1219_ & new_A1245_;
  assign new_A1227_ = new_A1243_ | new_A1242_;
  assign new_A1226_ = new_A1240_ | new_A1239_;
  assign new_A1225_ = new_A1208_ | new_A1241_;
  assign new_A1224_ = new_A1233_ & new_A1236_;
  assign new_A1223_ = new_A1238_ | new_A1237_;
  assign new_A1222_ = new_A1233_ & new_A1232_;
  assign new_A1221_ = new_A1235_ & new_A1234_;
  assign new_A1220_ = new_A1230_ | new_A1229_;
  assign new_A1219_ = new_A1208_ | new_A1231_;
  assign A1218 = new_A1219_ | new_A1228_;
  assign A1217 = new_A1226_ & new_A1227_;
  assign A1216 = new_A1226_ & new_A1225_;
  assign A1215 = new_A1224_ | new_A1223_;
  assign A1214 = new_A1222_ | new_A1221_;
  assign A1213 = new_A1220_ & new_A1219_;
  assign new_A1212_ = new_A3559_;
  assign new_A1211_ = new_A3492_;
  assign new_A1210_ = new_A3425_;
  assign new_A1209_ = new_A3358_;
  assign new_A1208_ = new_A3291_;
  assign new_A1207_ = new_A3227_;
  assign new_A1206_ = ~new_A1145_ & new_A1159_;
  assign new_A1205_ = new_A1145_ & ~new_A1159_;
  assign new_A1204_ = new_A1145_ & ~new_A1159_;
  assign new_A1203_ = ~new_A1145_ & ~new_A1159_;
  assign new_A1202_ = new_A1145_ & new_A1159_;
  assign new_A1201_ = new_A1205_ | new_A1206_;
  assign new_A1200_ = ~new_A1145_ & new_A1159_;
  assign new_A1199_ = new_A1203_ | new_A1204_;
  assign new_A1198_ = ~new_A1174_ & ~new_A1194_;
  assign new_A1197_ = new_A1174_ & new_A1194_;
  assign new_A1196_ = ~new_A1141_ | ~new_A1166_;
  assign new_A1195_ = new_A1159_ & new_A1196_;
  assign new_A1194_ = new_A1142_ | new_A1143_;
  assign new_A1193_ = new_A1142_ | new_A1159_;
  assign new_A1192_ = ~new_A1159_ & ~new_A1195_;
  assign new_A1191_ = new_A1159_ | new_A1196_;
  assign new_A1190_ = new_A1142_ & ~new_A1143_;
  assign new_A1189_ = ~new_A1142_ & new_A1143_;
  assign new_A1188_ = new_A1152_ | new_A1185_;
  assign new_A1187_ = ~new_A1152_ & ~new_A1186_;
  assign new_A1186_ = new_A1152_ & new_A1185_;
  assign new_A1185_ = ~new_A1141_ | ~new_A1166_;
  assign new_A1184_ = ~new_A1142_ & new_A1152_;
  assign new_A1183_ = new_A1142_ & ~new_A1152_;
  assign new_A1182_ = new_A1144_ & new_A1181_;
  assign new_A1181_ = new_A1200_ | new_A1199_;
  assign new_A1180_ = ~new_A1144_ & new_A1179_;
  assign new_A1179_ = new_A1202_ | new_A1201_;
  assign new_A1178_ = new_A1144_ | new_A1177_;
  assign new_A1177_ = new_A1198_ | new_A1197_;
  assign new_A1176_ = ~new_A1156_ & ~new_A1166_;
  assign new_A1175_ = new_A1156_ & new_A1166_;
  assign new_A1174_ = ~new_A1156_ | new_A1166_;
  assign new_A1173_ = new_A1140_ & ~new_A1141_;
  assign new_A1172_ = ~new_A1140_ & new_A1141_;
  assign new_A1171_ = new_A1193_ & ~new_A1194_;
  assign new_A1170_ = ~new_A1193_ & new_A1194_;
  assign new_A1169_ = ~new_A1192_ | ~new_A1191_;
  assign new_A1168_ = new_A1184_ | new_A1183_;
  assign new_A1167_ = new_A1190_ | new_A1189_;
  assign new_A1166_ = new_A1180_ | new_A1182_;
  assign new_A1165_ = ~new_A1187_ | ~new_A1188_;
  assign new_A1164_ = new_A1140_ & ~new_A1141_;
  assign new_A1163_ = new_A1154_ & ~new_A1166_;
  assign new_A1162_ = ~new_A1154_ & new_A1166_;
  assign new_A1161_ = ~new_A1152_ & new_A1178_;
  assign new_A1160_ = new_A1176_ | new_A1175_;
  assign new_A1159_ = new_A1173_ | new_A1172_;
  assign new_A1158_ = new_A1141_ | new_A1174_;
  assign new_A1157_ = new_A1166_ & new_A1169_;
  assign new_A1156_ = new_A1171_ | new_A1170_;
  assign new_A1155_ = new_A1166_ & new_A1165_;
  assign new_A1154_ = new_A1168_ & new_A1167_;
  assign new_A1153_ = new_A1163_ | new_A1162_;
  assign new_A1152_ = new_A1141_ | new_A1164_;
  assign A1151 = new_A1152_ | new_A1161_;
  assign A1150 = new_A1159_ & new_A1160_;
  assign A1149 = new_A1159_ & new_A1158_;
  assign A1148 = new_A1157_ | new_A1156_;
  assign A1147 = new_A1155_ | new_A1154_;
  assign A1146 = new_A1153_ & new_A1152_;
  assign new_A1145_ = new_A5568_;
  assign new_A1144_ = new_A5501_;
  assign new_A1143_ = new_A5434_;
  assign new_A1142_ = new_A5367_;
  assign new_A1141_ = new_A5300_;
  assign new_A1140_ = new_A5233_;
  assign new_A1139_ = ~new_A1078_ & new_A1092_;
  assign new_A1138_ = new_A1078_ & ~new_A1092_;
  assign new_A1137_ = new_A1078_ & ~new_A1092_;
  assign new_A1136_ = ~new_A1078_ & ~new_A1092_;
  assign new_A1135_ = new_A1078_ & new_A1092_;
  assign new_A1134_ = new_A1138_ | new_A1139_;
  assign new_A1133_ = ~new_A1078_ & new_A1092_;
  assign new_A1132_ = new_A1136_ | new_A1137_;
  assign new_A1131_ = ~new_A1107_ & ~new_A1127_;
  assign new_A1130_ = new_A1107_ & new_A1127_;
  assign new_A1129_ = ~new_A1074_ | ~new_A1099_;
  assign new_A1128_ = new_A1092_ & new_A1129_;
  assign new_A1127_ = new_A1075_ | new_A1076_;
  assign new_A1126_ = new_A1075_ | new_A1092_;
  assign new_A1125_ = ~new_A1092_ & ~new_A1128_;
  assign new_A1124_ = new_A1092_ | new_A1129_;
  assign new_A1123_ = new_A1075_ & ~new_A1076_;
  assign new_A1122_ = ~new_A1075_ & new_A1076_;
  assign new_A1121_ = new_A1085_ | new_A1118_;
  assign new_A1120_ = ~new_A1085_ & ~new_A1119_;
  assign new_A1119_ = new_A1085_ & new_A1118_;
  assign new_A1118_ = ~new_A1074_ | ~new_A1099_;
  assign new_A1117_ = ~new_A1075_ & new_A1085_;
  assign new_A1116_ = new_A1075_ & ~new_A1085_;
  assign new_A1115_ = new_A1077_ & new_A1114_;
  assign new_A1114_ = new_A1133_ | new_A1132_;
  assign new_A1113_ = ~new_A1077_ & new_A1112_;
  assign new_A1112_ = new_A1135_ | new_A1134_;
  assign new_A1111_ = new_A1077_ | new_A1110_;
  assign new_A1110_ = new_A1131_ | new_A1130_;
  assign new_A1109_ = ~new_A1089_ & ~new_A1099_;
  assign new_A1108_ = new_A1089_ & new_A1099_;
  assign new_A1107_ = ~new_A1089_ | new_A1099_;
  assign new_A1106_ = new_A1073_ & ~new_A1074_;
  assign new_A1105_ = ~new_A1073_ & new_A1074_;
  assign new_A1104_ = new_A1126_ & ~new_A1127_;
  assign new_A1103_ = ~new_A1126_ & new_A1127_;
  assign new_A1102_ = ~new_A1125_ | ~new_A1124_;
  assign new_A1101_ = new_A1117_ | new_A1116_;
  assign new_A1100_ = new_A1123_ | new_A1122_;
  assign new_A1099_ = new_A1113_ | new_A1115_;
  assign new_A1098_ = ~new_A1120_ | ~new_A1121_;
  assign new_A1097_ = new_A1073_ & ~new_A1074_;
  assign new_A1096_ = new_A1087_ & ~new_A1099_;
  assign new_A1095_ = ~new_A1087_ & new_A1099_;
  assign new_A1094_ = ~new_A1085_ & new_A1111_;
  assign new_A1093_ = new_A1109_ | new_A1108_;
  assign new_A1092_ = new_A1106_ | new_A1105_;
  assign new_A1091_ = new_A1074_ | new_A1107_;
  assign new_A1090_ = new_A1099_ & new_A1102_;
  assign new_A1089_ = new_A1104_ | new_A1103_;
  assign new_A1088_ = new_A1099_ & new_A1098_;
  assign new_A1087_ = new_A1101_ & new_A1100_;
  assign new_A1086_ = new_A1096_ | new_A1095_;
  assign new_A1085_ = new_A1074_ | new_A1097_;
  assign A1084 = new_A1085_ | new_A1094_;
  assign A1083 = new_A1092_ & new_A1093_;
  assign A1082 = new_A1092_ & new_A1091_;
  assign A1081 = new_A1090_ | new_A1089_;
  assign A1080 = new_A1088_ | new_A1087_;
  assign A1079 = new_A1086_ & new_A1085_;
  assign new_A1078_ = new_A5166_;
  assign new_A1077_ = new_A5099_;
  assign new_A1076_ = new_A5032_;
  assign new_A1075_ = new_A4965_;
  assign new_A1074_ = new_A4898_;
  assign new_A1073_ = new_A4831_;
  assign new_A1072_ = ~new_A1011_ & new_A1025_;
  assign new_A1071_ = new_A1011_ & ~new_A1025_;
  assign new_A1070_ = new_A1011_ & ~new_A1025_;
  assign new_A1069_ = ~new_A1011_ & ~new_A1025_;
  assign new_A1068_ = new_A1011_ & new_A1025_;
  assign new_A1067_ = new_A1071_ | new_A1072_;
  assign new_A1066_ = ~new_A1011_ & new_A1025_;
  assign new_A1065_ = new_A1069_ | new_A1070_;
  assign new_A1064_ = ~new_A1040_ & ~new_A1060_;
  assign new_A1063_ = new_A1040_ & new_A1060_;
  assign new_A1062_ = ~new_A1007_ | ~new_A1032_;
  assign new_A1061_ = new_A1025_ & new_A1062_;
  assign new_A1060_ = new_A1008_ | new_A1009_;
  assign new_A1059_ = new_A1008_ | new_A1025_;
  assign new_A1058_ = ~new_A1025_ & ~new_A1061_;
  assign new_A1057_ = new_A1025_ | new_A1062_;
  assign new_A1056_ = new_A1008_ & ~new_A1009_;
  assign new_A1055_ = ~new_A1008_ & new_A1009_;
  assign new_A1054_ = new_A1018_ | new_A1051_;
  assign new_A1053_ = ~new_A1018_ & ~new_A1052_;
  assign new_A1052_ = new_A1018_ & new_A1051_;
  assign new_A1051_ = ~new_A1007_ | ~new_A1032_;
  assign new_A1050_ = ~new_A1008_ & new_A1018_;
  assign new_A1049_ = new_A1008_ & ~new_A1018_;
  assign new_A1048_ = new_A1010_ & new_A1047_;
  assign new_A1047_ = new_A1066_ | new_A1065_;
  assign new_A1046_ = ~new_A1010_ & new_A1045_;
  assign new_A1045_ = new_A1068_ | new_A1067_;
  assign new_A1044_ = new_A1010_ | new_A1043_;
  assign new_A1043_ = new_A1064_ | new_A1063_;
  assign new_A1042_ = ~new_A1022_ & ~new_A1032_;
  assign new_A1041_ = new_A1022_ & new_A1032_;
  assign new_A1040_ = ~new_A1022_ | new_A1032_;
  assign new_A1039_ = new_A1006_ & ~new_A1007_;
  assign new_A1038_ = ~new_A1006_ & new_A1007_;
  assign new_A1037_ = new_A1059_ & ~new_A1060_;
  assign new_A1036_ = ~new_A1059_ & new_A1060_;
  assign new_A1035_ = ~new_A1058_ | ~new_A1057_;
  assign new_A1034_ = new_A1050_ | new_A1049_;
  assign new_A1033_ = new_A1056_ | new_A1055_;
  assign new_A1032_ = new_A1046_ | new_A1048_;
  assign new_A1031_ = ~new_A1053_ | ~new_A1054_;
  assign new_A1030_ = new_A1006_ & ~new_A1007_;
  assign new_A1029_ = new_A1020_ & ~new_A1032_;
  assign new_A1028_ = ~new_A1020_ & new_A1032_;
  assign new_A1027_ = ~new_A1018_ & new_A1044_;
  assign new_A1026_ = new_A1042_ | new_A1041_;
  assign new_A1025_ = new_A1039_ | new_A1038_;
  assign new_A1024_ = new_A1007_ | new_A1040_;
  assign new_A1023_ = new_A1032_ & new_A1035_;
  assign new_A1022_ = new_A1037_ | new_A1036_;
  assign new_A1021_ = new_A1032_ & new_A1031_;
  assign new_A1020_ = new_A1034_ & new_A1033_;
  assign new_A1019_ = new_A1029_ | new_A1028_;
  assign new_A1018_ = new_A1007_ | new_A1030_;
  assign A1017 = new_A1018_ | new_A1027_;
  assign A1016 = new_A1025_ & new_A1026_;
  assign A1015 = new_A1025_ & new_A1024_;
  assign A1014 = new_A1023_ | new_A1022_;
  assign A1013 = new_A1021_ | new_A1020_;
  assign A1012 = new_A1019_ & new_A1018_;
  assign new_A1011_ = new_A4764_;
  assign new_A1010_ = new_A4697_;
  assign new_A1009_ = new_A4630_;
  assign new_A1008_ = new_A4563_;
  assign new_A1007_ = new_A4496_;
  assign new_A1006_ = new_A4429_;
  assign new_A1005_ = ~new_A944_ & new_A958_;
  assign new_A1004_ = new_A944_ & ~new_A958_;
  assign new_A1003_ = new_A944_ & ~new_A958_;
  assign new_A1002_ = ~new_A944_ & ~new_A958_;
  assign new_A1001_ = new_A944_ & new_A958_;
  assign new_A1000_ = new_A1004_ | new_A1005_;
  assign new_A999_ = ~new_A944_ & new_A958_;
  assign new_A998_ = new_A1002_ | new_A1003_;
  assign new_A997_ = ~new_A973_ & ~new_A993_;
  assign new_A996_ = new_A973_ & new_A993_;
  assign new_A995_ = ~new_A940_ | ~new_A965_;
  assign new_A994_ = new_A958_ & new_A995_;
  assign new_A993_ = new_A941_ | new_A942_;
  assign new_A992_ = new_A941_ | new_A958_;
  assign new_A991_ = ~new_A958_ & ~new_A994_;
  assign new_A990_ = new_A958_ | new_A995_;
  assign new_A989_ = new_A941_ & ~new_A942_;
  assign new_A988_ = ~new_A941_ & new_A942_;
  assign new_A987_ = new_A951_ | new_A984_;
  assign new_A986_ = ~new_A951_ & ~new_A985_;
  assign new_A985_ = new_A951_ & new_A984_;
  assign new_A984_ = ~new_A940_ | ~new_A965_;
  assign new_A983_ = ~new_A941_ & new_A951_;
  assign new_A982_ = new_A941_ & ~new_A951_;
  assign new_A981_ = new_A943_ & new_A980_;
  assign new_A980_ = new_A999_ | new_A998_;
  assign new_A979_ = ~new_A943_ & new_A978_;
  assign new_A978_ = new_A1001_ | new_A1000_;
  assign new_A977_ = new_A943_ | new_A976_;
  assign new_A976_ = new_A997_ | new_A996_;
  assign new_A975_ = ~new_A955_ & ~new_A965_;
  assign new_A974_ = new_A955_ & new_A965_;
  assign new_A973_ = ~new_A955_ | new_A965_;
  assign new_A972_ = new_A939_ & ~new_A940_;
  assign new_A971_ = ~new_A939_ & new_A940_;
  assign new_A970_ = new_A992_ & ~new_A993_;
  assign new_A969_ = ~new_A992_ & new_A993_;
  assign new_A968_ = ~new_A991_ | ~new_A990_;
  assign new_A967_ = new_A983_ | new_A982_;
  assign new_A966_ = new_A989_ | new_A988_;
  assign new_A965_ = new_A979_ | new_A981_;
  assign new_A964_ = ~new_A986_ | ~new_A987_;
  assign new_A963_ = new_A939_ & ~new_A940_;
  assign new_A962_ = new_A953_ & ~new_A965_;
  assign new_A961_ = ~new_A953_ & new_A965_;
  assign new_A960_ = ~new_A951_ & new_A977_;
  assign new_A959_ = new_A975_ | new_A974_;
  assign new_A958_ = new_A972_ | new_A971_;
  assign new_A957_ = new_A940_ | new_A973_;
  assign new_A956_ = new_A965_ & new_A968_;
  assign new_A955_ = new_A970_ | new_A969_;
  assign new_A954_ = new_A965_ & new_A964_;
  assign new_A953_ = new_A967_ & new_A966_;
  assign new_A952_ = new_A962_ | new_A961_;
  assign new_A951_ = new_A940_ | new_A963_;
  assign A950 = new_A951_ | new_A960_;
  assign A949 = new_A958_ & new_A959_;
  assign A948 = new_A958_ & new_A957_;
  assign A947 = new_A956_ | new_A955_;
  assign A946 = new_A954_ | new_A953_;
  assign A945 = new_A952_ & new_A951_;
  assign new_A944_ = new_A4362_;
  assign new_A943_ = new_A4295_;
  assign new_A942_ = new_A4228_;
  assign new_A941_ = new_A4161_;
  assign new_A940_ = new_A4094_;
  assign new_A939_ = new_A4027_;
  assign new_A938_ = ~new_A877_ & new_A891_;
  assign new_A937_ = new_A877_ & ~new_A891_;
  assign new_A936_ = new_A877_ & ~new_A891_;
  assign new_A935_ = ~new_A877_ & ~new_A891_;
  assign new_A934_ = new_A877_ & new_A891_;
  assign new_A933_ = new_A937_ | new_A938_;
  assign new_A932_ = ~new_A877_ & new_A891_;
  assign new_A931_ = new_A935_ | new_A936_;
  assign new_A930_ = ~new_A906_ & ~new_A926_;
  assign new_A929_ = new_A906_ & new_A926_;
  assign new_A928_ = ~new_A873_ | ~new_A898_;
  assign new_A927_ = new_A891_ & new_A928_;
  assign new_A926_ = new_A874_ | new_A875_;
  assign new_A925_ = new_A874_ | new_A891_;
  assign new_A924_ = ~new_A891_ & ~new_A927_;
  assign new_A923_ = new_A891_ | new_A928_;
  assign new_A922_ = new_A874_ & ~new_A875_;
  assign new_A921_ = ~new_A874_ & new_A875_;
  assign new_A920_ = new_A884_ | new_A917_;
  assign new_A919_ = ~new_A884_ & ~new_A918_;
  assign new_A918_ = new_A884_ & new_A917_;
  assign new_A917_ = ~new_A873_ | ~new_A898_;
  assign new_A916_ = ~new_A874_ & new_A884_;
  assign new_A915_ = new_A874_ & ~new_A884_;
  assign new_A914_ = new_A876_ & new_A913_;
  assign new_A913_ = new_A932_ | new_A931_;
  assign new_A912_ = ~new_A876_ & new_A911_;
  assign new_A911_ = new_A934_ | new_A933_;
  assign new_A910_ = new_A876_ | new_A909_;
  assign new_A909_ = new_A930_ | new_A929_;
  assign new_A908_ = ~new_A888_ & ~new_A898_;
  assign new_A907_ = new_A888_ & new_A898_;
  assign new_A906_ = ~new_A888_ | new_A898_;
  assign new_A905_ = new_A872_ & ~new_A873_;
  assign new_A904_ = ~new_A872_ & new_A873_;
  assign new_A903_ = new_A925_ & ~new_A926_;
  assign new_A902_ = ~new_A925_ & new_A926_;
  assign new_A901_ = ~new_A924_ | ~new_A923_;
  assign new_A900_ = new_A916_ | new_A915_;
  assign new_A899_ = new_A922_ | new_A921_;
  assign new_A898_ = new_A912_ | new_A914_;
  assign new_A897_ = ~new_A919_ | ~new_A920_;
  assign new_A896_ = new_A872_ & ~new_A873_;
  assign new_A895_ = new_A886_ & ~new_A898_;
  assign new_A894_ = ~new_A886_ & new_A898_;
  assign new_A893_ = ~new_A884_ & new_A910_;
  assign new_A892_ = new_A908_ | new_A907_;
  assign new_A891_ = new_A905_ | new_A904_;
  assign new_A890_ = new_A873_ | new_A906_;
  assign new_A889_ = new_A898_ & new_A901_;
  assign new_A888_ = new_A903_ | new_A902_;
  assign new_A887_ = new_A898_ & new_A897_;
  assign new_A886_ = new_A900_ & new_A899_;
  assign new_A885_ = new_A895_ | new_A894_;
  assign new_A884_ = new_A873_ | new_A896_;
  assign A883 = new_A884_ | new_A893_;
  assign A882 = new_A891_ & new_A892_;
  assign A881 = new_A891_ & new_A890_;
  assign A880 = new_A889_ | new_A888_;
  assign A879 = new_A887_ | new_A886_;
  assign A878 = new_A885_ & new_A884_;
  assign new_A877_ = new_A3960_;
  assign new_A876_ = new_A3893_;
  assign new_A875_ = new_A3826_;
  assign new_A874_ = new_A3759_;
  assign new_A873_ = new_A3692_;
  assign new_A872_ = new_A3625_;
  assign new_A805_ = new_A3558_;
  assign new_A806_ = new_A3491_;
  assign new_A807_ = new_A3424_;
  assign new_A808_ = new_A3357_;
  assign new_A809_ = new_A3290_;
  assign new_A810_ = new_A3228_;
  assign A811 = new_A818_ & new_A817_;
  assign A812 = new_A820_ | new_A819_;
  assign A813 = new_A822_ | new_A821_;
  assign A814 = new_A824_ & new_A823_;
  assign A815 = new_A824_ & new_A825_;
  assign A816 = new_A817_ | new_A826_;
  assign new_A817_ = new_A806_ | new_A829_;
  assign new_A818_ = new_A828_ | new_A827_;
  assign new_A819_ = new_A833_ & new_A832_;
  assign new_A820_ = new_A831_ & new_A830_;
  assign new_A821_ = new_A836_ | new_A835_;
  assign new_A822_ = new_A831_ & new_A834_;
  assign new_A823_ = new_A806_ | new_A839_;
  assign new_A824_ = new_A838_ | new_A837_;
  assign new_A825_ = new_A841_ | new_A840_;
  assign new_A826_ = ~new_A817_ & new_A843_;
  assign new_A827_ = ~new_A819_ & new_A831_;
  assign new_A828_ = new_A819_ & ~new_A831_;
  assign new_A829_ = new_A805_ & ~new_A806_;
  assign new_A830_ = ~new_A852_ | ~new_A853_;
  assign new_A831_ = new_A845_ | new_A847_;
  assign new_A832_ = new_A855_ | new_A854_;
  assign new_A833_ = new_A849_ | new_A848_;
  assign new_A834_ = ~new_A857_ | ~new_A856_;
  assign new_A835_ = ~new_A858_ & new_A859_;
  assign new_A836_ = new_A858_ & ~new_A859_;
  assign new_A837_ = ~new_A805_ & new_A806_;
  assign new_A838_ = new_A805_ & ~new_A806_;
  assign new_A839_ = ~new_A821_ | new_A831_;
  assign new_A840_ = new_A821_ & new_A831_;
  assign new_A841_ = ~new_A821_ & ~new_A831_;
  assign new_A842_ = new_A863_ | new_A862_;
  assign new_A843_ = new_A809_ | new_A842_;
  assign new_A844_ = new_A867_ | new_A866_;
  assign new_A845_ = ~new_A809_ & new_A844_;
  assign new_A846_ = new_A865_ | new_A864_;
  assign new_A847_ = new_A809_ & new_A846_;
  assign new_A848_ = new_A807_ & ~new_A817_;
  assign new_A849_ = ~new_A807_ & new_A817_;
  assign new_A850_ = ~new_A806_ | ~new_A831_;
  assign new_A851_ = new_A817_ & new_A850_;
  assign new_A852_ = ~new_A817_ & ~new_A851_;
  assign new_A853_ = new_A817_ | new_A850_;
  assign new_A854_ = ~new_A807_ & new_A808_;
  assign new_A855_ = new_A807_ & ~new_A808_;
  assign new_A856_ = new_A824_ | new_A861_;
  assign new_A857_ = ~new_A824_ & ~new_A860_;
  assign new_A858_ = new_A807_ | new_A824_;
  assign new_A859_ = new_A807_ | new_A808_;
  assign new_A860_ = new_A824_ & new_A861_;
  assign new_A861_ = ~new_A806_ | ~new_A831_;
  assign new_A862_ = new_A839_ & new_A859_;
  assign new_A863_ = ~new_A839_ & ~new_A859_;
  assign new_A864_ = new_A868_ | new_A869_;
  assign new_A865_ = ~new_A810_ & new_A824_;
  assign new_A866_ = new_A870_ | new_A871_;
  assign new_A867_ = new_A810_ & new_A824_;
  assign new_A868_ = ~new_A810_ & ~new_A824_;
  assign new_A869_ = new_A810_ & ~new_A824_;
  assign new_A870_ = new_A810_ & ~new_A824_;
  assign new_A871_ = ~new_A810_ & new_A824_;
endmodule


