// Benchmark "systemcaes" written by ABC on Thu Oct  8 22:04:26 2020

module systemcaes ( clock, 
    clk, reset, load_i, decrypt_i, \data_i[0] , \data_i[1] , \data_i[2] ,
    \data_i[3] , \data_i[4] , \data_i[5] , \data_i[6] , \data_i[7] ,
    \data_i[8] , \data_i[9] , \data_i[10] , \data_i[11] , \data_i[12] ,
    \data_i[13] , \data_i[14] , \data_i[15] , \data_i[16] , \data_i[17] ,
    \data_i[18] , \data_i[19] , \data_i[20] , \data_i[21] , \data_i[22] ,
    \data_i[23] , \data_i[24] , \data_i[25] , \data_i[26] , \data_i[27] ,
    \data_i[28] , \data_i[29] , \data_i[30] , \data_i[31] , \data_i[32] ,
    \data_i[33] , \data_i[34] , \data_i[35] , \data_i[36] , \data_i[37] ,
    \data_i[38] , \data_i[39] , \data_i[40] , \data_i[41] , \data_i[42] ,
    \data_i[43] , \data_i[44] , \data_i[45] , \data_i[46] , \data_i[47] ,
    \data_i[48] , \data_i[49] , \data_i[50] , \data_i[51] , \data_i[52] ,
    \data_i[53] , \data_i[54] , \data_i[55] , \data_i[56] , \data_i[57] ,
    \data_i[58] , \data_i[59] , \data_i[60] , \data_i[61] , \data_i[62] ,
    \data_i[63] , \data_i[64] , \data_i[65] , \data_i[66] , \data_i[67] ,
    \data_i[68] , \data_i[69] , \data_i[70] , \data_i[71] , \data_i[72] ,
    \data_i[73] , \data_i[74] , \data_i[75] , \data_i[76] , \data_i[77] ,
    \data_i[78] , \data_i[79] , \data_i[80] , \data_i[81] , \data_i[82] ,
    \data_i[83] , \data_i[84] , \data_i[85] , \data_i[86] , \data_i[87] ,
    \data_i[88] , \data_i[89] , \data_i[90] , \data_i[91] , \data_i[92] ,
    \data_i[93] , \data_i[94] , \data_i[95] , \data_i[96] , \data_i[97] ,
    \data_i[98] , \data_i[99] , \data_i[100] , \data_i[101] ,
    \data_i[102] , \data_i[103] , \data_i[104] , \data_i[105] ,
    \data_i[106] , \data_i[107] , \data_i[108] , \data_i[109] ,
    \data_i[110] , \data_i[111] , \data_i[112] , \data_i[113] ,
    \data_i[114] , \data_i[115] , \data_i[116] , \data_i[117] ,
    \data_i[118] , \data_i[119] , \data_i[120] , \data_i[121] ,
    \data_i[122] , \data_i[123] , \data_i[124] , \data_i[125] ,
    \data_i[126] , \data_i[127] , \key_i[0] , \key_i[1] , \key_i[2] ,
    \key_i[3] , \key_i[4] , \key_i[5] , \key_i[6] , \key_i[7] , \key_i[8] ,
    \key_i[9] , \key_i[10] , \key_i[11] , \key_i[12] , \key_i[13] ,
    \key_i[14] , \key_i[15] , \key_i[16] , \key_i[17] , \key_i[18] ,
    \key_i[19] , \key_i[20] , \key_i[21] , \key_i[22] , \key_i[23] ,
    \key_i[24] , \key_i[25] , \key_i[26] , \key_i[27] , \key_i[28] ,
    \key_i[29] , \key_i[30] , \key_i[31] , \key_i[32] , \key_i[33] ,
    \key_i[34] , \key_i[35] , \key_i[36] , \key_i[37] , \key_i[38] ,
    \key_i[39] , \key_i[40] , \key_i[41] , \key_i[42] , \key_i[43] ,
    \key_i[44] , \key_i[45] , \key_i[46] , \key_i[47] , \key_i[48] ,
    \key_i[49] , \key_i[50] , \key_i[51] , \key_i[52] , \key_i[53] ,
    \key_i[54] , \key_i[55] , \key_i[56] , \key_i[57] , \key_i[58] ,
    \key_i[59] , \key_i[60] , \key_i[61] , \key_i[62] , \key_i[63] ,
    \key_i[64] , \key_i[65] , \key_i[66] , \key_i[67] , \key_i[68] ,
    \key_i[69] , \key_i[70] , \key_i[71] , \key_i[72] , \key_i[73] ,
    \key_i[74] , \key_i[75] , \key_i[76] , \key_i[77] , \key_i[78] ,
    \key_i[79] , \key_i[80] , \key_i[81] , \key_i[82] , \key_i[83] ,
    \key_i[84] , \key_i[85] , \key_i[86] , \key_i[87] , \key_i[88] ,
    \key_i[89] , \key_i[90] , \key_i[91] , \key_i[92] , \key_i[93] ,
    \key_i[94] , \key_i[95] , \key_i[96] , \key_i[97] , \key_i[98] ,
    \key_i[99] , \key_i[100] , \key_i[101] , \key_i[102] , \key_i[103] ,
    \key_i[104] , \key_i[105] , \key_i[106] , \key_i[107] , \key_i[108] ,
    \key_i[109] , \key_i[110] , \key_i[111] , \key_i[112] , \key_i[113] ,
    \key_i[114] , \key_i[115] , \key_i[116] , \key_i[117] , \key_i[118] ,
    \key_i[119] , \key_i[120] , \key_i[121] , \key_i[122] , \key_i[123] ,
    \key_i[124] , \key_i[125] , \key_i[126] , \key_i[127] ,
    ready_o, \data_o[0] , \data_o[1] , \data_o[2] , \data_o[3] ,
    \data_o[4] , \data_o[5] , \data_o[6] , \data_o[7] , \data_o[8] ,
    \data_o[9] , \data_o[10] , \data_o[11] , \data_o[12] , \data_o[13] ,
    \data_o[14] , \data_o[15] , \data_o[16] , \data_o[17] , \data_o[18] ,
    \data_o[19] , \data_o[20] , \data_o[21] , \data_o[22] , \data_o[23] ,
    \data_o[24] , \data_o[25] , \data_o[26] , \data_o[27] , \data_o[28] ,
    \data_o[29] , \data_o[30] , \data_o[31] , \data_o[32] , \data_o[33] ,
    \data_o[34] , \data_o[35] , \data_o[36] , \data_o[37] , \data_o[38] ,
    \data_o[39] , \data_o[40] , \data_o[41] , \data_o[42] , \data_o[43] ,
    \data_o[44] , \data_o[45] , \data_o[46] , \data_o[47] , \data_o[48] ,
    \data_o[49] , \data_o[50] , \data_o[51] , \data_o[52] , \data_o[53] ,
    \data_o[54] , \data_o[55] , \data_o[56] , \data_o[57] , \data_o[58] ,
    \data_o[59] , \data_o[60] , \data_o[61] , \data_o[62] , \data_o[63] ,
    \data_o[64] , \data_o[65] , \data_o[66] , \data_o[67] , \data_o[68] ,
    \data_o[69] , \data_o[70] , \data_o[71] , \data_o[72] , \data_o[73] ,
    \data_o[74] , \data_o[75] , \data_o[76] , \data_o[77] , \data_o[78] ,
    \data_o[79] , \data_o[80] , \data_o[81] , \data_o[82] , \data_o[83] ,
    \data_o[84] , \data_o[85] , \data_o[86] , \data_o[87] , \data_o[88] ,
    \data_o[89] , \data_o[90] , \data_o[91] , \data_o[92] , \data_o[93] ,
    \data_o[94] , \data_o[95] , \data_o[96] , \data_o[97] , \data_o[98] ,
    \data_o[99] , \data_o[100] , \data_o[101] , \data_o[102] ,
    \data_o[103] , \data_o[104] , \data_o[105] , \data_o[106] ,
    \data_o[107] , \data_o[108] , \data_o[109] , \data_o[110] ,
    \data_o[111] , \data_o[112] , \data_o[113] , \data_o[114] ,
    \data_o[115] , \data_o[116] , \data_o[117] , \data_o[118] ,
    \data_o[119] , \data_o[120] , \data_o[121] , \data_o[122] ,
    \data_o[123] , \data_o[124] , \data_o[125] , \data_o[126] ,
    \data_o[127]   );
  input  clock;
  input  clk, reset, load_i, decrypt_i, \data_i[0] , \data_i[1] ,
    \data_i[2] , \data_i[3] , \data_i[4] , \data_i[5] , \data_i[6] ,
    \data_i[7] , \data_i[8] , \data_i[9] , \data_i[10] , \data_i[11] ,
    \data_i[12] , \data_i[13] , \data_i[14] , \data_i[15] , \data_i[16] ,
    \data_i[17] , \data_i[18] , \data_i[19] , \data_i[20] , \data_i[21] ,
    \data_i[22] , \data_i[23] , \data_i[24] , \data_i[25] , \data_i[26] ,
    \data_i[27] , \data_i[28] , \data_i[29] , \data_i[30] , \data_i[31] ,
    \data_i[32] , \data_i[33] , \data_i[34] , \data_i[35] , \data_i[36] ,
    \data_i[37] , \data_i[38] , \data_i[39] , \data_i[40] , \data_i[41] ,
    \data_i[42] , \data_i[43] , \data_i[44] , \data_i[45] , \data_i[46] ,
    \data_i[47] , \data_i[48] , \data_i[49] , \data_i[50] , \data_i[51] ,
    \data_i[52] , \data_i[53] , \data_i[54] , \data_i[55] , \data_i[56] ,
    \data_i[57] , \data_i[58] , \data_i[59] , \data_i[60] , \data_i[61] ,
    \data_i[62] , \data_i[63] , \data_i[64] , \data_i[65] , \data_i[66] ,
    \data_i[67] , \data_i[68] , \data_i[69] , \data_i[70] , \data_i[71] ,
    \data_i[72] , \data_i[73] , \data_i[74] , \data_i[75] , \data_i[76] ,
    \data_i[77] , \data_i[78] , \data_i[79] , \data_i[80] , \data_i[81] ,
    \data_i[82] , \data_i[83] , \data_i[84] , \data_i[85] , \data_i[86] ,
    \data_i[87] , \data_i[88] , \data_i[89] , \data_i[90] , \data_i[91] ,
    \data_i[92] , \data_i[93] , \data_i[94] , \data_i[95] , \data_i[96] ,
    \data_i[97] , \data_i[98] , \data_i[99] , \data_i[100] , \data_i[101] ,
    \data_i[102] , \data_i[103] , \data_i[104] , \data_i[105] ,
    \data_i[106] , \data_i[107] , \data_i[108] , \data_i[109] ,
    \data_i[110] , \data_i[111] , \data_i[112] , \data_i[113] ,
    \data_i[114] , \data_i[115] , \data_i[116] , \data_i[117] ,
    \data_i[118] , \data_i[119] , \data_i[120] , \data_i[121] ,
    \data_i[122] , \data_i[123] , \data_i[124] , \data_i[125] ,
    \data_i[126] , \data_i[127] , \key_i[0] , \key_i[1] , \key_i[2] ,
    \key_i[3] , \key_i[4] , \key_i[5] , \key_i[6] , \key_i[7] , \key_i[8] ,
    \key_i[9] , \key_i[10] , \key_i[11] , \key_i[12] , \key_i[13] ,
    \key_i[14] , \key_i[15] , \key_i[16] , \key_i[17] , \key_i[18] ,
    \key_i[19] , \key_i[20] , \key_i[21] , \key_i[22] , \key_i[23] ,
    \key_i[24] , \key_i[25] , \key_i[26] , \key_i[27] , \key_i[28] ,
    \key_i[29] , \key_i[30] , \key_i[31] , \key_i[32] , \key_i[33] ,
    \key_i[34] , \key_i[35] , \key_i[36] , \key_i[37] , \key_i[38] ,
    \key_i[39] , \key_i[40] , \key_i[41] , \key_i[42] , \key_i[43] ,
    \key_i[44] , \key_i[45] , \key_i[46] , \key_i[47] , \key_i[48] ,
    \key_i[49] , \key_i[50] , \key_i[51] , \key_i[52] , \key_i[53] ,
    \key_i[54] , \key_i[55] , \key_i[56] , \key_i[57] , \key_i[58] ,
    \key_i[59] , \key_i[60] , \key_i[61] , \key_i[62] , \key_i[63] ,
    \key_i[64] , \key_i[65] , \key_i[66] , \key_i[67] , \key_i[68] ,
    \key_i[69] , \key_i[70] , \key_i[71] , \key_i[72] , \key_i[73] ,
    \key_i[74] , \key_i[75] , \key_i[76] , \key_i[77] , \key_i[78] ,
    \key_i[79] , \key_i[80] , \key_i[81] , \key_i[82] , \key_i[83] ,
    \key_i[84] , \key_i[85] , \key_i[86] , \key_i[87] , \key_i[88] ,
    \key_i[89] , \key_i[90] , \key_i[91] , \key_i[92] , \key_i[93] ,
    \key_i[94] , \key_i[95] , \key_i[96] , \key_i[97] , \key_i[98] ,
    \key_i[99] , \key_i[100] , \key_i[101] , \key_i[102] , \key_i[103] ,
    \key_i[104] , \key_i[105] , \key_i[106] , \key_i[107] , \key_i[108] ,
    \key_i[109] , \key_i[110] , \key_i[111] , \key_i[112] , \key_i[113] ,
    \key_i[114] , \key_i[115] , \key_i[116] , \key_i[117] , \key_i[118] ,
    \key_i[119] , \key_i[120] , \key_i[121] , \key_i[122] , \key_i[123] ,
    \key_i[124] , \key_i[125] , \key_i[126] , \key_i[127] ;
  output ready_o, \data_o[0] , \data_o[1] , \data_o[2] , \data_o[3] ,
    \data_o[4] , \data_o[5] , \data_o[6] , \data_o[7] , \data_o[8] ,
    \data_o[9] , \data_o[10] , \data_o[11] , \data_o[12] , \data_o[13] ,
    \data_o[14] , \data_o[15] , \data_o[16] , \data_o[17] , \data_o[18] ,
    \data_o[19] , \data_o[20] , \data_o[21] , \data_o[22] , \data_o[23] ,
    \data_o[24] , \data_o[25] , \data_o[26] , \data_o[27] , \data_o[28] ,
    \data_o[29] , \data_o[30] , \data_o[31] , \data_o[32] , \data_o[33] ,
    \data_o[34] , \data_o[35] , \data_o[36] , \data_o[37] , \data_o[38] ,
    \data_o[39] , \data_o[40] , \data_o[41] , \data_o[42] , \data_o[43] ,
    \data_o[44] , \data_o[45] , \data_o[46] , \data_o[47] , \data_o[48] ,
    \data_o[49] , \data_o[50] , \data_o[51] , \data_o[52] , \data_o[53] ,
    \data_o[54] , \data_o[55] , \data_o[56] , \data_o[57] , \data_o[58] ,
    \data_o[59] , \data_o[60] , \data_o[61] , \data_o[62] , \data_o[63] ,
    \data_o[64] , \data_o[65] , \data_o[66] , \data_o[67] , \data_o[68] ,
    \data_o[69] , \data_o[70] , \data_o[71] , \data_o[72] , \data_o[73] ,
    \data_o[74] , \data_o[75] , \data_o[76] , \data_o[77] , \data_o[78] ,
    \data_o[79] , \data_o[80] , \data_o[81] , \data_o[82] , \data_o[83] ,
    \data_o[84] , \data_o[85] , \data_o[86] , \data_o[87] , \data_o[88] ,
    \data_o[89] , \data_o[90] , \data_o[91] , \data_o[92] , \data_o[93] ,
    \data_o[94] , \data_o[95] , \data_o[96] , \data_o[97] , \data_o[98] ,
    \data_o[99] , \data_o[100] , \data_o[101] , \data_o[102] ,
    \data_o[103] , \data_o[104] , \data_o[105] , \data_o[106] ,
    \data_o[107] , \data_o[108] , \data_o[109] , \data_o[110] ,
    \data_o[111] , \data_o[112] , \data_o[113] , \data_o[114] ,
    \data_o[115] , \data_o[116] , \data_o[117] , \data_o[118] ,
    \data_o[119] , \data_o[120] , \data_o[121] , \data_o[122] ,
    \data_o[123] , \data_o[124] , \data_o[125] , \data_o[126] ,
    \data_o[127] ;
  reg \\ks1_key_reg_reg[11] , \\ks1_key_reg_reg[12] ,
    \\ks1_key_reg_reg[13] , \\ks1_key_reg_reg[14] , \\ks1_key_reg_reg[15] ,
    \\sbox1_to_invert_reg[1] , \\sbox1_to_invert_reg[3] ,
    \\sbox1_to_invert_reg[2] , \\sbox1_to_invert_reg[0] ,
    \\ks1_key_reg_reg[8] , \\ks1_key_reg_reg[10] , \\ks1_key_reg_reg[9] ,
    \\ks1_key_reg_reg[43] , \\ks1_key_reg_reg[44] , \\ks1_key_reg_reg[45] ,
    \\ks1_key_reg_reg[46] , \\ks1_key_reg_reg[47] , \\ks1_key_reg_reg[40] ,
    \\sub1_data_reg_reg[109] , \\sub1_data_reg_reg[110] ,
    \\sub1_data_reg_reg[13] , \\sub1_data_reg_reg[14] ,
    \\sub1_data_reg_reg[45] , \\sub1_data_reg_reg[46] ,
    \\sub1_data_reg_reg[77] , \\sub1_data_reg_reg[78] ,
    \\sub1_data_reg_reg[102] , \\sub1_data_reg_reg[101] ,
    \\sub1_data_reg_reg[118] , \\sub1_data_reg_reg[117] ,
    \\sub1_data_reg_reg[21] , \\sub1_data_reg_reg[22] ,
    \\sub1_data_reg_reg[37] , \\sub1_data_reg_reg[38] ,
    \\sub1_data_reg_reg[53] , \\sub1_data_reg_reg[54] ,
    \\sub1_data_reg_reg[5] , \\sub1_data_reg_reg[6] ,
    \\sub1_data_reg_reg[70] , \\sub1_data_reg_reg[69] ,
    \\sub1_data_reg_reg[85] , \\sub1_data_reg_reg[86] ,
    \\ks1_key_reg_reg[42] , \\ks1_key_reg_reg[41] , \\ks1_key_reg_reg[76] ,
    \\ks1_key_reg_reg[75] , \\ks1_key_reg_reg[74] , \\ks1_key_reg_reg[73] ,
    \\ks1_key_reg_reg[77] , \\ks1_key_reg_reg[78] ,
    \\sub1_data_reg_reg[125] , \\sub1_data_reg_reg[126] ,
    \\sub1_data_reg_reg[29] , \\sub1_data_reg_reg[94] ,
    \\sub1_data_reg_reg[30] , \\sub1_data_reg_reg[93] ,
    \\ks1_key_reg_reg[72] , \\ks1_key_reg_reg[79] ,
    \\sub1_data_reg_reg[104] , \\sub1_data_reg_reg[40] ,
    \\sub1_data_reg_reg[72] , \\sub1_data_reg_reg[8] ,
    \\sub1_data_reg_reg[0] , \\sub1_data_reg_reg[112] ,
    \\sub1_data_reg_reg[16] , \\sub1_data_reg_reg[64] ,
    \\sub1_data_reg_reg[80] , \\sub1_data_reg_reg[96] ,
    \\sub1_data_reg_reg[48] , \\sub1_data_reg_reg[61] ,
    \\sub1_data_reg_reg[62] , \\ks1_col_reg[21] , \\ks1_col_reg[22] ,
    \\sub1_data_reg_reg[107] , \\sub1_data_reg_reg[108] ,
    \\sub1_data_reg_reg[111] , \\sub1_data_reg_reg[11] ,
    \\sub1_data_reg_reg[12] , \\sub1_data_reg_reg[15] ,
    \\sub1_data_reg_reg[44] , \\sub1_data_reg_reg[43] ,
    \\sub1_data_reg_reg[47] , \\sub1_data_reg_reg[75] ,
    \\sub1_data_reg_reg[76] , \\sub1_data_reg_reg[79] ,
    \\sub1_data_reg_reg[103] , \\sub1_data_reg_reg[115] ,
    \\sub1_data_reg_reg[116] , \\sub1_data_reg_reg[119] ,
    \\sub1_data_reg_reg[20] , \\sub1_data_reg_reg[19] ,
    \\sub1_data_reg_reg[23] , \\sub1_data_reg_reg[32] ,
    \\sub1_data_reg_reg[4] , \\sub1_data_reg_reg[51] ,
    \\sub1_data_reg_reg[52] , \\sub1_data_reg_reg[55] ,
    \\sub1_data_reg_reg[36] , \\sub1_data_reg_reg[68] ,
    \\sub1_data_reg_reg[67] , \\sub1_data_reg_reg[3] ,
    \\sub1_data_reg_reg[7] , \\sub1_data_reg_reg[71] ,
    \\sub1_data_reg_reg[84] , \\sub1_data_reg_reg[83] ,
    \\sub1_data_reg_reg[87] , \\sub1_data_reg_reg[120] ,
    \\sub1_data_reg_reg[24] , \\sub1_data_reg_reg[56] ,
    \\sub1_data_reg_reg[88] , \\sbox1_alph_reg[2] , \\ks1_col_reg[30] ,
    \\sub1_data_reg_reg[100] , \\ks1_col_reg[6] , \\ks1_col_reg[5] ,
    \\sub1_data_reg_reg[35] , \\sub1_data_reg_reg[39] , \\ks1_col_reg[29] ,
    \\sub1_data_reg_reg[99] , \\sub1_data_reg_reg[123] ,
    \\sub1_data_reg_reg[124] , \\sub1_data_reg_reg[127] ,
    \\sub1_data_reg_reg[27] , \\sub1_data_reg_reg[28] ,
    \\sub1_data_reg_reg[31] , \\sub1_data_reg_reg[59] ,
    \\sub1_data_reg_reg[60] , \\sub1_data_reg_reg[63] ,
    \\sub1_data_reg_reg[95] , \\sub1_data_reg_reg[91] ,
    \\sub1_data_reg_reg[92] , \\ks1_col_reg[16] , \\sbox1_alph_reg[0] ,
    \\ks1_key_reg_reg[107] , \\ks1_key_reg_reg[108] , \\ks1_col_reg[20] ,
    \\ks1_key_reg_reg[104] , \\ks1_col_reg[23] , \\ks1_col_reg[19] ,
    \\sub1_data_reg_reg[106] , \\sub1_data_reg_reg[10] ,
    \\sub1_data_reg_reg[74] , \\sub1_data_reg_reg[42] ,
    \\sub1_data_reg_reg[114] , \\ks1_col_reg[24] , \\ks1_col_reg[3] ,
    \\ks1_col_reg[4] , \\sub1_data_reg_reg[18] , \\sub1_data_reg_reg[2] ,
    \\sub1_data_reg_reg[50] , \\sub1_data_reg_reg[66] ,
    \\sub1_data_reg_reg[82] , \\sub1_data_reg_reg[98] , \\ks1_col_reg[0] ,
    \\ks1_col_reg[28] , \\ks1_key_reg_reg[111] , \\ks1_col_reg[27] ,
    \\ks1_col_reg[31] , \\sub1_data_reg_reg[34] , \\ks1_col_reg[7] ,
    \\sub1_data_reg_reg[122] , \\sub1_data_reg_reg[26] ,
    \\sub1_data_reg_reg[58] , \\sub1_data_reg_reg[90] ,
    \\sbox1_ah_reg_reg[2] , \\sbox1_alph_reg[1] , \\ks1_key_reg_reg[110] ,
    \\ks1_key_reg_reg[109] , \\sub1_data_reg_reg[105] ,
    \\sub1_data_reg_reg[41] , \\sub1_data_reg_reg[73] ,
    \\sub1_data_reg_reg[9] , \\sub1_data_reg_reg[17] ,
    \\sub1_data_reg_reg[1] , \\sub1_data_reg_reg[65] ,
    \\sub1_data_reg_reg[97] , \\ks1_key_reg_reg[105] , \\ks1_col_reg[18] ,
    \\sbox1_ah_reg_reg[0] , \\sub1_data_reg_reg[81] ,
    \\sub1_data_reg_reg[49] , \\sub1_data_reg_reg[113] ,
    \\sub1_data_reg_reg[33] , \\sub1_data_reg_reg[57] ,
    \\sub1_data_reg_reg[89] , \\sub1_data_reg_reg[25] , \\ks1_col_reg[26] ,
    \\sub1_data_reg_reg[121] , \\ks1_key_reg_reg[106] , \\ks1_col_reg[2] ,
    \\sbox1_ah_reg_reg[1] , \\ks1_col_reg[17] , \\sbox1_alph_reg[3] ,
    \\ks1_col_reg[25] , \\ks1_col_reg[1] , \\sbox1_ah_reg_reg[3] ,
    \\ks1_key_reg_reg[28] , \\ks1_key_reg_reg[27] , \\ks1_key_reg_reg[29] ,
    \\ks1_key_reg_reg[30] , \\ks1_key_reg_reg[24] , \\ks1_key_reg_reg[31] ,
    \\ks1_key_reg_reg[25] , \\ks1_key_reg_reg[26] , \\ks1_key_reg_reg[60] ,
    \\ks1_key_reg_reg[2] , \\ks1_key_reg_reg[3] , \\ks1_key_reg_reg[4] ,
    \\ks1_key_reg_reg[5] , \\ks1_key_reg_reg[6] , \\ks1_key_reg_reg[0] ,
    \\ks1_key_reg_reg[1] , \\ks1_key_reg_reg[23] , \\ks1_key_reg_reg[7] ,
    \\ks1_key_reg_reg[61] , \\ks1_key_reg_reg[59] , \\ks1_key_reg_reg[17] ,
    \\ks1_key_reg_reg[16] , \\ks1_key_reg_reg[19] , \\ks1_key_reg_reg[18] ,
    \\ks1_key_reg_reg[21] , \\ks1_key_reg_reg[22] , \\ks1_key_reg_reg[20] ,
    \\ks1_key_reg_reg[57] , \\ks1_key_reg_reg[58] , \\ks1_key_reg_reg[63] ,
    \\ks1_key_reg_reg[62] , \\ks1_key_reg_reg[56] , \\ks1_key_reg_reg[92] ,
    \\ks1_key_reg_reg[32] , \\ks1_key_reg_reg[33] , \\ks1_key_reg_reg[34] ,
    \\ks1_key_reg_reg[35] , \\ks1_key_reg_reg[36] , \\ks1_key_reg_reg[38] ,
    \\ks1_key_reg_reg[39] , \\ks1_key_reg_reg[55] , \\ks1_key_reg_reg[37] ,
    \\ks1_key_reg_reg[91] , \\ks1_key_reg_reg[93] , \\ks1_key_reg_reg[49] ,
    \\ks1_key_reg_reg[50] , \\ks1_key_reg_reg[51] , \\ks1_key_reg_reg[52] ,
    \\ks1_key_reg_reg[54] , \\ks1_key_reg_reg[48] , \\ks1_key_reg_reg[53] ,
    \\ks1_key_reg_reg[90] , \\ks1_key_reg_reg[88] , \\ks1_key_reg_reg[94] ,
    \\ks1_key_reg_reg[95] , \\ks1_key_reg_reg[89] , \\ks1_key_reg_reg[69] ,
    \\addroundkey_data_reg_reg[60] , \\addroundkey_data_reg_reg[111] ,
    \\addroundkey_data_reg_reg[63] , \\addroundkey_data_reg_reg[6] ,
    \\addroundkey_data_reg_reg[76] , \\addroundkey_data_reg_reg[25] ,
    \\addroundkey_data_reg_reg[77] , \\addroundkey_data_reg_reg[78] ,
    \\addroundkey_data_reg_reg[79] , \\addroundkey_data_reg_reg[26] ,
    \\addroundkey_data_reg_reg[29] , \\addroundkey_data_reg_reg[8] ,
    \\addroundkey_data_reg_reg[105] , \\addroundkey_data_reg_reg[0] ,
    \\addroundkey_data_reg_reg[106] , \\addroundkey_data_reg_reg[107] ,
    \\addroundkey_data_reg_reg[122] , \\addroundkey_data_reg_reg[3] ,
    \\addroundkey_data_reg_reg[41] , \\addroundkey_data_reg_reg[123] ,
    \\addroundkey_data_reg_reg[42] , \\addroundkey_data_reg_reg[43] ,
    \\addroundkey_data_reg_reg[44] , \\addroundkey_data_reg_reg[108] ,
    \\addroundkey_data_reg_reg[125] , \\addroundkey_data_reg_reg[46] ,
    \\addroundkey_data_reg_reg[47] , \\addroundkey_data_reg_reg[126] ,
    \\addroundkey_data_reg_reg[127] , \\addroundkey_data_reg_reg[10] ,
    \\addroundkey_data_reg_reg[13] , \\addroundkey_data_reg_reg[110] ,
    \\addroundkey_data_reg_reg[58] , \\addroundkey_data_reg_reg[57] ,
    \\addroundkey_data_reg_reg[59] , \\ks1_key_reg_reg[124] ,
    \\ks1_key_reg_reg[64] , \\ks1_key_reg_reg[65] , \\ks1_key_reg_reg[67] ,
    \\ks1_key_reg_reg[66] , \\ks1_key_reg_reg[68] , \\ks1_key_reg_reg[70] ,
    \\ks1_key_reg_reg[71] , \\ks1_key_reg_reg[87] ,
    \\addroundkey_data_reg_reg[5] , \\ks1_key_reg_reg[81] ,
    \\addroundkey_data_reg_reg[40] , \\addroundkey_data_reg_reg[124] ,
    \\addroundkey_data_reg_reg[61] , \\addroundkey_data_reg_reg[62] ,
    \\addroundkey_data_reg_reg[1] , \\addroundkey_data_reg_reg[73] ,
    \\addroundkey_data_reg_reg[74] , \\addroundkey_data_reg_reg[24] ,
    \\addroundkey_data_reg_reg[72] , \\addroundkey_data_reg_reg[7] ,
    \\addroundkey_data_reg_reg[28] , \\addroundkey_data_reg_reg[104] ,
    \\addroundkey_data_reg_reg[30] , \\addroundkey_data_reg_reg[2] ,
    \\addroundkey_data_reg_reg[31] , \\addroundkey_data_reg_reg[90] ,
    \\addroundkey_data_reg_reg[91] , \\addroundkey_data_reg_reg[92] ,
    \\addroundkey_data_reg_reg[34] , \\addroundkey_data_reg_reg[93] ,
    \\addroundkey_data_reg_reg[11] , \\addroundkey_data_reg_reg[94] ,
    \\addroundkey_data_reg_reg[95] , \\addroundkey_data_reg_reg[120] ,
    \\addroundkey_data_reg_reg[9] , \\addroundkey_data_reg_reg[121] ,
    \\addroundkey_data_reg_reg[45] , \\addroundkey_data_reg_reg[4] ,
    \\addroundkey_data_reg_reg[12] , \\addroundkey_data_reg_reg[109] ,
    \\addroundkey_data_reg_reg[14] , \\addroundkey_data_reg_reg[56] ,
    \\addroundkey_data_reg_reg[15] , \\ks1_key_reg_reg[125] ,
    \\ks1_key_reg_reg[123] , \\ks1_key_reg_reg[80] ,
    \\ks1_key_reg_reg[83] , \\ks1_key_reg_reg[84] , \\ks1_key_reg_reg[85] ,
    \\ks1_key_reg_reg[82] , \\ks1_key_reg_reg[86] ,
    \\addroundkey_data_reg_reg[27] , \\addroundkey_data_reg_reg[75] ,
    \\addroundkey_data_reg_reg[100] , \\addroundkey_data_reg_reg[33] ,
    \\addroundkey_data_reg_reg[103] , \\addroundkey_data_reg_reg[98] ,
    \\addroundkey_data_reg_reg[35] , \\mix1_data_reg_reg[100] ,
    \\mix1_data_reg_reg[108] , \\mix1_data_reg_reg[116] ,
    \\mix1_data_reg_reg[124] , \\addroundkey_data_reg_reg[101] ,
    \\addroundkey_data_reg_reg[112] , \\addroundkey_data_reg_reg[64] ,
    \\addroundkey_data_reg_reg[65] , \\addroundkey_data_reg_reg[20] ,
    \\addroundkey_data_reg_reg[66] , \\addroundkey_data_reg_reg[67] ,
    \\addroundkey_data_reg_reg[21] , \\addroundkey_data_reg_reg[69] ,
    \\addroundkey_data_reg_reg[22] , \\addroundkey_data_reg_reg[70] ,
    \\addroundkey_data_reg_reg[102] , \\addroundkey_data_reg_reg[23] ,
    \\addroundkey_data_reg_reg[115] , \\addroundkey_data_reg_reg[116] ,
    \\addroundkey_data_reg_reg[80] , \\addroundkey_data_reg_reg[81] ,
    \\addroundkey_data_reg_reg[83] , \\addroundkey_data_reg_reg[85] ,
    \\addroundkey_data_reg_reg[86] , \\addroundkey_data_reg_reg[84] ,
    \\addroundkey_data_reg_reg[87] , \\addroundkey_data_reg_reg[88] ,
    \\addroundkey_data_reg_reg[32] , \\addroundkey_data_reg_reg[119] ,
    \\addroundkey_data_reg_reg[96] , \\addroundkey_data_reg_reg[97] ,
    \\addroundkey_data_reg_reg[36] , \\addroundkey_data_reg_reg[99] ,
    \\addroundkey_data_reg_reg[37] , \\addroundkey_data_reg_reg[38] ,
    \\addroundkey_data_reg_reg[39] , \\addroundkey_data_reg_reg[49] ,
    \\addroundkey_data_reg_reg[52] , \\addroundkey_data_reg_reg[55] ,
    \\addroundkey_data_reg_reg[17] , \\ks1_key_reg_reg[120] ,
    \\ks1_key_reg_reg[121] , \\ks1_key_reg_reg[127] ,
    \\addroundkey_round_reg[0] , \\addroundkey_data_reg_reg[118] ,
    \\addroundkey_data_reg_reg[89] , \\addroundkey_data_reg_reg[117] ,
    \\ks1_key_reg_reg[126] , \\addroundkey_data_reg_reg[82] ,
    \\ks1_key_reg_reg[122] , \\addroundkey_data_reg_reg[114] ,
    \\addroundkey_data_reg_reg[54] , \\addroundkey_data_reg_reg[71] ,
    \\addroundkey_data_reg_reg[16] , \\addroundkey_data_reg_reg[68] ,
    \\addroundkey_data_reg_reg[53] , \\addroundkey_data_reg_reg[113] ,
    \\addroundkey_data_reg_reg[19] , \\addroundkey_data_reg_reg[51] ,
    \\addroundkey_data_reg_reg[50] , \\addroundkey_data_reg_reg[18] ,
    \\addroundkey_data_reg_reg[48] , \\ks1_key_reg_reg[97] ,
    \\mix1_data_reg_reg[107] , \\mix1_data_reg_reg[115] ,
    \\mix1_data_reg_reg[99] , \\ks1_key_reg_reg[96] ,
    \\ks1_key_reg_reg[98] , \\ks1_key_reg_reg[100] ,
    \\ks1_key_reg_reg[101] , \\ks1_key_reg_reg[102] ,
    \\ks1_key_reg_reg[103] , \\ks1_key_reg_reg[119] ,
    \\mix1_data_reg_reg[123] , \\ks1_key_reg_reg[113] ,
    \\mix1_data_reg_reg[36] , \\mix1_data_reg_reg[44] ,
    \\mix1_data_reg_reg[60] , \\mix1_data_reg_reg[68] ,
    \\mix1_data_reg_reg[52] , \\mix1_data_reg_reg[84] ,
    \\mix1_data_reg_reg[76] , \\mix1_data_reg_reg[92] ,
    \\ks1_key_reg_reg[112] , \\ks1_key_reg_reg[115] ,
    \\ks1_key_reg_reg[116] , \\ks1_key_reg_reg[114] ,
    \\ks1_key_reg_reg[118] , addroundkey_ready_o_reg,
    \\ks1_key_reg_reg[117] , \\ks1_key_reg_reg[99] ,
    \\mix1_data_reg_reg[105] , \\mix1_data_reg_reg[106] ,
    \\mix1_data_reg_reg[113] , \\mix1_data_reg_reg[114] ,
    \\mix1_data_reg_reg[121] , \\mix1_data_reg_reg[122] ,
    \\mix1_data_reg_reg[35] , \\mix1_data_reg_reg[43] ,
    \\mix1_data_reg_reg[51] , \\mix1_data_reg_reg[59] ,
    \\mix1_data_reg_reg[67] , \\mix1_data_reg_reg[75] ,
    \\mix1_data_reg_reg[97] , \\mix1_data_reg_reg[98] ,
    \\mix1_data_reg_reg[91] , \\mix1_data_reg_reg[83] ,
    \\mix1_data_reg_reg[120] , \\mix1_data_reg_reg[117] ,
    \\mix1_data_reg_reg[125] , \\mix1_data_reg_reg[118] ,
    \\mix1_data_reg_reg[104] , \\mix1_data_reg_reg[112] ,
    \\mix1_data_reg_reg[96] , \\mix1_data_reg_reg[126] ,
    \\mix1_data_reg_reg[110] , \\mix1_data_reg_reg[102] ,
    \\mix1_data_reg_reg[109] , \\mix1_data_reg_reg[101] ,
    \\mix1_data_o_reg_reg[12] , \\mix1_data_o_reg_reg[20] ,
    \\mix1_data_o_reg_reg[28] , \\mix1_data_o_reg_reg[4] ,
    \\mix1_data_reg_reg[33] , \\mix1_data_reg_reg[34] ,
    \\mix1_data_reg_reg[42] , \\mix1_data_reg_reg[41] ,
    \\mix1_data_reg_reg[49] , \\mix1_data_reg_reg[50] ,
    \\mix1_data_reg_reg[57] , \\mix1_data_reg_reg[58] ,
    \\mix1_data_reg_reg[65] , \\mix1_data_reg_reg[66] ,
    \\mix1_data_reg_reg[74] , \\mix1_data_reg_reg[73] ,
    \\mix1_data_reg_reg[81] , \\mix1_data_reg_reg[82] ,
    \\mix1_data_reg_reg[89] , \\mix1_data_reg_reg[90] ,
    \\mix1_data_reg_reg[61] , \\mix1_data_reg_reg[62] ,
    \\mix1_data_reg_reg[69] , \\mix1_data_reg_reg[45] ,
    \\mix1_data_reg_reg[37] , \\mix1_data_reg_reg[53] ,
    \\mix1_data_reg_reg[77] , \\mix1_data_o_reg_reg[3] ,
    \\mix1_data_reg_reg[38] , \\mix1_data_reg_reg[46] ,
    \\mix1_data_reg_reg[54] , \\mix1_data_reg_reg[70] ,
    \\mix1_data_reg_reg[78] , \\mix1_data_reg_reg[86] ,
    \\mix1_data_reg_reg[94] , \\mix1_data_reg_reg[32] ,
    \\mix1_data_reg_reg[48] , \\mix1_data_reg_reg[56] ,
    \\mix1_data_reg_reg[64] , \\mix1_data_reg_reg[88] ,
    \\mix1_data_reg_reg[80] , \\mix1_data_reg_reg[72] ,
    \\mix1_data_reg_reg[40] , \\mix1_data_o_reg_reg[27] ,
    \\mix1_data_o_reg_reg[11] , \\mix1_data_o_reg_reg[19] ,
    \\mix1_data_reg_reg[85] , \\mix1_data_reg_reg[93] ,
    \\mix1_data_reg_reg[103] , \\mix1_data_reg_reg[111] ,
    \\mix1_data_reg_reg[127] , \\mix1_data_reg_reg[119] ,
    \\mix1_data_o_reg_reg[17] , \\mix1_data_o_reg_reg[18] ,
    \\mix1_data_o_reg_reg[1] , \\mix1_data_o_reg_reg[25] ,
    \\mix1_data_o_reg_reg[26] , \\mix1_data_o_reg_reg[9] ,
    \\mix1_data_o_reg_reg[2] , \\mix1_data_o_reg_reg[10] ,
    \\mix1_data_reg_reg[79] , \\mix1_data_o_reg_reg[8] ,
    \\mix1_data_reg_reg[55] , \\mix1_data_reg_reg[71] ,
    \\mix1_data_o_reg_reg[13] , \\mix1_data_o_reg_reg[21] ,
    \\mix1_data_reg_reg[63] , \\mix1_data_o_reg_reg[22] ,
    \\mix1_data_o_reg_reg[30] , \\mix1_data_o_reg_reg[16] ,
    \\mix1_data_reg_reg[47] , \\mix1_data_reg_reg[39] ,
    \\mix1_data_o_reg_reg[6] , \\mix1_data_o_reg_reg[14] ,
    \\mix1_data_o_reg_reg[0] , \\mix1_data_o_reg_reg[24] ,
    \\mix1_data_reg_reg[95] , \\mix1_data_o_reg_reg[29] ,
    \\mix1_data_o_reg_reg[5] , \\mix1_data_reg_reg[87] ,
    \\mix1_data_o_reg_reg[7] , \\mix1_data_o_reg_reg[23] ,
    \\mix1_data_o_reg_reg[31] , \\mix1_data_o_reg_reg[15] ,
    \\addroundkey_round_reg[1] , \\addroundkey_round_reg[3] ,
    \\addroundkey_round_reg[2] , \\ks1_state_reg[0] , \\ks1_state_reg[2] ,
    \\round_reg[1] , \\round_reg[2] , \\round_reg[0] , \\round_reg[3] ,
    addroundkey_start_i_reg, \\mix1_state_reg[0] , \\mix1_state_reg[1] ,
    state_reg, \\sub1_state_reg[0] , ready_o_reg, \\sub1_state_reg[3] ,
    \\sub1_state_reg[2] , \\sub1_state_reg[1] , \\sub1_state_reg[4] ,
    \\mix1_data_o_reg_reg[104] , \\mix1_data_o_reg_reg[102] ,
    \\mix1_data_o_reg_reg[105] , \\mix1_data_o_reg_reg[108] ,
    \\mix1_data_o_reg_reg[110] , \\mix1_data_o_reg_reg[112] ,
    \\mix1_data_o_reg_reg[45] , \\mix1_data_o_reg_reg[67] ,
    \\mix1_data_o_reg_reg[70] , \\mix1_data_o_reg_reg[85] ,
    \\mix1_data_o_reg_reg[98] , \\mix1_data_o_reg_reg[82] ,
    \\mix1_data_o_reg_reg[99] , \\mix1_data_o_reg_reg[72] ,
    \\mix1_data_o_reg_reg[48] , \\mix1_data_o_reg_reg[91] ,
    \\mix1_data_o_reg_reg[69] , \\mix1_data_o_reg_reg[57] ,
    \\mix1_data_o_reg_reg[33] , \\mix1_data_o_reg_reg[65] ,
    \\mix1_data_o_reg_reg[71] , \\mix1_data_o_reg_reg[93] ,
    \\mix1_data_o_reg_reg[106] , \\mix1_data_o_reg_reg[77] ,
    \\mix1_data_o_reg_reg[78] , \\mix1_data_o_reg_reg[122] ,
    \\mix1_data_o_reg_reg[64] , \\mix1_data_o_reg_reg[49] ,
    \\mix1_data_o_reg_reg[116] , \\mix1_data_o_reg_reg[86] ,
    \\mix1_data_o_reg_reg[88] , \\mix1_data_o_reg_reg[89] ,
    \\mix1_data_o_reg_reg[126] , \\mix1_data_o_reg_reg[90] ,
    \\mix1_data_o_reg_reg[74] , \\mix1_data_o_reg_reg[56] ,
    \\mix1_data_o_reg_reg[47] , \\mix1_data_o_reg_reg[97] ,
    \\mix1_data_o_reg_reg[43] , \\mix1_data_o_reg_reg[76] ,
    \\mix1_data_o_reg_reg[37] , \\mix1_data_o_reg_reg[84] ,
    \\mix1_data_o_reg_reg[103] , \\mix1_data_o_reg_reg[109] ,
    \\mix1_data_o_reg_reg[53] , \\mix1_data_o_reg_reg[119] ,
    \\mix1_data_o_reg_reg[125] , \\mix1_data_o_reg_reg[36] ,
    \\mix1_data_o_reg_reg[39] , \\mix1_data_o_reg_reg[55] ,
    \\mix1_data_o_reg_reg[62] , \\mix1_data_o_reg_reg[96] ,
    \\mix1_data_o_reg_reg[115] , \\mix1_data_o_reg_reg[46] ,
    \\mix1_data_o_reg_reg[80] , \\mix1_data_o_reg_reg[123] ,
    \\mix1_data_o_reg_reg[83] , \\mix1_data_o_reg_reg[58] ,
    \\mix1_data_o_reg_reg[68] , \\mix1_data_o_reg_reg[101] ,
    \\mix1_data_o_reg_reg[118] , \\mix1_data_o_reg_reg[52] ,
    \\mix1_data_o_reg_reg[59] , \\mix1_data_o_reg_reg[87] ,
    \\mix1_data_o_reg_reg[51] , \\mix1_data_o_reg_reg[66] ,
    \\mix1_data_o_reg_reg[81] , \\mix1_data_o_reg_reg[107] ,
    \\mix1_data_o_reg_reg[44] , \\mix1_data_o_reg_reg[42] ,
    \\mix1_data_o_reg_reg[94] , \\mix1_data_o_reg_reg[54] ,
    \\mix1_data_o_reg_reg[50] , \\mix1_data_o_reg_reg[124] ,
    \\mix1_data_o_reg_reg[32] , \\mix1_data_o_reg_reg[75] ,
    \\mix1_data_o_reg_reg[61] , \\mix1_data_o_reg_reg[63] ,
    \\mix1_data_o_reg_reg[120] , \\mix1_data_o_reg_reg[40] ,
    \\mix1_data_o_reg_reg[111] , \\mix1_data_o_reg_reg[34] ,
    \\mix1_data_o_reg_reg[113] , \\mix1_data_o_reg_reg[41] ,
    \\mix1_data_o_reg_reg[121] , \\mix1_data_o_reg_reg[92] ,
    \\mix1_data_o_reg_reg[117] , \\mix1_data_o_reg_reg[60] ,
    \\mix1_data_o_reg_reg[114] , \\mix1_data_o_reg_reg[38] ,
    \\mix1_data_o_reg_reg[73] , \\mix1_data_o_reg_reg[127] ,
    \\mix1_data_o_reg_reg[95] , \\mix1_data_o_reg_reg[79] ,
    \\mix1_data_o_reg_reg[35] , \\mix1_data_o_reg_reg[100] ,
    ks1_ready_o_reg, mix1_ready_o_reg, first_round_reg_reg,
    \\ks1_state_reg[1] , sub1_ready_o_reg;
  wire \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1072]_ , \new_[1076]_ ,
    \new_[1078]_ , \new_[1079]_ , \new_[1080]_ , \new_[1082]_ ,
    \new_[1083]_ , \new_[1084]_ , \new_[1085]_ , \new_[1086]_ ,
    \new_[1087]_ , \new_[1088]_ , \new_[1089]_ , \new_[1090]_ ,
    \new_[1091]_ , \new_[1092]_ , \new_[1093]_ , \new_[1094]_ ,
    \new_[1095]_ , \new_[1096]_ , \new_[1097]_ , \new_[1098]_ ,
    \new_[1099]_ , \new_[1100]_ , \new_[1101]_ , \new_[1102]_ ,
    \new_[1103]_ , \new_[1104]_ , \new_[1105]_ , \new_[1106]_ ,
    \new_[1107]_ , \new_[1108]_ , \new_[1109]_ , \new_[1110]_ ,
    \new_[1111]_ , \new_[1112]_ , \new_[1113]_ , \new_[1114]_ ,
    \new_[1115]_ , \new_[1116]_ , \new_[1117]_ , \new_[1118]_ ,
    \new_[1119]_ , \new_[1120]_ , \new_[1121]_ , \new_[1122]_ ,
    \new_[1123]_ , \new_[1124]_ , \new_[1125]_ , \new_[1126]_ ,
    \new_[1127]_ , \new_[1128]_ , \new_[1129]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1176]_ , \new_[1177]_ , \new_[1178]_ , \new_[1179]_ ,
    \new_[1180]_ , \new_[1181]_ , \new_[1182]_ , \new_[1183]_ ,
    \new_[1184]_ , \new_[1185]_ , \new_[1186]_ , \new_[1187]_ ,
    \new_[1188]_ , \new_[1189]_ , \new_[1190]_ , \new_[1191]_ ,
    \new_[1192]_ , \new_[1193]_ , \new_[1194]_ , \new_[1195]_ ,
    \new_[1196]_ , \new_[1197]_ , \new_[1198]_ , \new_[1199]_ ,
    \new_[1200]_ , \new_[1201]_ , \new_[1202]_ , \new_[1203]_ ,
    \new_[1204]_ , \new_[1205]_ , \new_[1206]_ , \new_[1207]_ ,
    \new_[1208]_ , \new_[1209]_ , \new_[1210]_ , \new_[1211]_ ,
    \new_[1212]_ , \new_[1213]_ , \new_[1214]_ , \new_[1215]_ ,
    \new_[1216]_ , \new_[1217]_ , \new_[1218]_ , \new_[1219]_ ,
    \new_[1220]_ , \new_[1221]_ , \new_[1222]_ , \new_[1223]_ ,
    \new_[1224]_ , \new_[1225]_ , \new_[1226]_ , \new_[1227]_ ,
    \new_[1228]_ , \new_[1231]_ , \new_[1232]_ , \new_[1233]_ ,
    \new_[1234]_ , \new_[1235]_ , \new_[1236]_ , \new_[1237]_ ,
    \new_[1238]_ , \new_[1239]_ , \new_[1240]_ , \new_[1241]_ ,
    \new_[1242]_ , \new_[1243]_ , \new_[1244]_ , \new_[1245]_ ,
    \new_[1246]_ , \new_[1247]_ , \new_[1248]_ , \new_[1249]_ ,
    \new_[1250]_ , \new_[1251]_ , \new_[1252]_ , \new_[1253]_ ,
    \new_[1254]_ , \new_[1255]_ , \new_[1256]_ , \new_[1257]_ ,
    \new_[1258]_ , \new_[1259]_ , \new_[1260]_ , \new_[1261]_ ,
    \new_[1262]_ , \new_[1263]_ , \new_[1264]_ , \new_[1265]_ ,
    \new_[1266]_ , \new_[1267]_ , \new_[1268]_ , \new_[1269]_ ,
    \new_[1270]_ , \new_[1272]_ , \new_[1274]_ , \new_[1279]_ ,
    \new_[1280]_ , \new_[1281]_ , \new_[1282]_ , \new_[1283]_ ,
    \new_[1284]_ , \new_[1285]_ , \new_[1286]_ , \new_[1287]_ ,
    \new_[1289]_ , \new_[1297]_ , \new_[1298]_ , \new_[1299]_ ,
    \new_[1300]_ , \new_[1305]_ , \new_[1306]_ , \new_[1307]_ ,
    \new_[1308]_ , \new_[1309]_ , \new_[1310]_ , \new_[1311]_ ,
    \new_[1312]_ , \new_[1313]_ , \new_[1314]_ , \new_[1315]_ ,
    \new_[1316]_ , \new_[1317]_ , \new_[1318]_ , \new_[1319]_ ,
    \new_[1320]_ , \new_[1321]_ , \new_[1322]_ , \new_[1323]_ ,
    \new_[1324]_ , \new_[1331]_ , \new_[1332]_ , \new_[1333]_ ,
    \new_[1343]_ , \new_[1355]_ , \new_[1356]_ , \new_[1357]_ ,
    \new_[1358]_ , \new_[1375]_ , \new_[1377]_ , \new_[1378]_ ,
    \new_[1379]_ , \new_[1380]_ , \new_[1381]_ , \new_[1382]_ ,
    \new_[1383]_ , \new_[1384]_ , \new_[1385]_ , \new_[1386]_ ,
    \new_[1387]_ , \new_[1388]_ , \new_[1389]_ , \new_[1390]_ ,
    \new_[1391]_ , \new_[1392]_ , \new_[1393]_ , \new_[1394]_ ,
    \new_[1395]_ , \new_[1408]_ , \new_[1409]_ , \new_[1410]_ ,
    \new_[1411]_ , \new_[1414]_ , \new_[1416]_ , \new_[1417]_ ,
    \new_[1418]_ , \new_[1419]_ , \new_[1420]_ , \new_[1421]_ ,
    \new_[1422]_ , \new_[1423]_ , \new_[1424]_ , \new_[1425]_ ,
    \new_[1426]_ , \new_[1427]_ , \new_[1428]_ , \new_[1429]_ ,
    \new_[1430]_ , \new_[1431]_ , \new_[1432]_ , \new_[1433]_ ,
    \new_[1434]_ , \new_[1435]_ , \new_[1436]_ , \new_[1437]_ ,
    \new_[1438]_ , \new_[1439]_ , \new_[1440]_ , \new_[1441]_ ,
    \new_[1442]_ , \new_[1443]_ , \new_[1444]_ , \new_[1453]_ ,
    \new_[1454]_ , \new_[1455]_ , \new_[1456]_ , \new_[1457]_ ,
    \new_[1458]_ , \new_[1459]_ , \new_[1460]_ , \new_[1461]_ ,
    \new_[1462]_ , \new_[1463]_ , \new_[1464]_ , \new_[1465]_ ,
    \new_[1466]_ , \new_[1467]_ , \new_[1468]_ , \new_[1469]_ ,
    \new_[1470]_ , \new_[1471]_ , \new_[1472]_ , \new_[1473]_ ,
    \new_[1474]_ , \new_[1475]_ , \new_[1476]_ , \new_[1477]_ ,
    \new_[1478]_ , \new_[1479]_ , \new_[1480]_ , \new_[1481]_ ,
    \new_[1482]_ , \new_[1483]_ , \new_[1484]_ , \new_[1485]_ ,
    \new_[1486]_ , \new_[1487]_ , \new_[1488]_ , \new_[1489]_ ,
    \new_[1490]_ , \new_[1491]_ , \new_[1492]_ , \new_[1493]_ ,
    \new_[1494]_ , \new_[1495]_ , \new_[1496]_ , \new_[1497]_ ,
    \new_[1498]_ , \new_[1499]_ , \new_[1500]_ , \new_[1501]_ ,
    \new_[1502]_ , \new_[1503]_ , \new_[1504]_ , \new_[1505]_ ,
    \new_[1506]_ , \new_[1507]_ , \new_[1508]_ , \new_[1512]_ ,
    \new_[1520]_ , \new_[1521]_ , \new_[1522]_ , \new_[1530]_ ,
    \new_[1535]_ , \new_[1536]_ , \new_[1537]_ , \new_[1538]_ ,
    \new_[1539]_ , \new_[1540]_ , \new_[1541]_ , \new_[1542]_ ,
    \new_[1543]_ , \new_[1544]_ , \new_[1545]_ , \new_[1546]_ ,
    \new_[1548]_ , \new_[1549]_ , \new_[1550]_ , \new_[1551]_ ,
    \new_[1552]_ , \new_[1553]_ , \new_[1554]_ , \new_[1555]_ ,
    \new_[1556]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1577]_ ,
    \new_[1582]_ , \new_[1583]_ , \new_[1584]_ , \new_[1585]_ ,
    \new_[1586]_ , \new_[1587]_ , \new_[1588]_ , \new_[1590]_ ,
    \new_[1591]_ , \new_[1592]_ , \new_[1593]_ , \new_[1594]_ ,
    \new_[1595]_ , \new_[1596]_ , \new_[1604]_ , \new_[1605]_ ,
    \new_[1606]_ , \new_[1607]_ , \new_[1608]_ , \new_[1609]_ ,
    \new_[1610]_ , \new_[1611]_ , \new_[1612]_ , \new_[1613]_ ,
    \new_[1614]_ , \new_[1615]_ , \new_[1616]_ , \new_[1617]_ ,
    \new_[1618]_ , \new_[1619]_ , \new_[1620]_ , \new_[1621]_ ,
    \new_[1622]_ , \new_[1623]_ , \new_[1624]_ , \new_[1625]_ ,
    \new_[1626]_ , \new_[1627]_ , \new_[1628]_ , \new_[1629]_ ,
    \new_[1630]_ , \new_[1631]_ , \new_[1632]_ , \new_[1633]_ ,
    \new_[1634]_ , \new_[1635]_ , \new_[1636]_ , \new_[1637]_ ,
    \new_[1638]_ , \new_[1639]_ , \new_[1640]_ , \new_[1641]_ ,
    \new_[1642]_ , \new_[1643]_ , \new_[1644]_ , \new_[1645]_ ,
    \new_[1646]_ , \new_[1647]_ , \new_[1648]_ , \new_[1649]_ ,
    \new_[1650]_ , \new_[1651]_ , \new_[1652]_ , \new_[1653]_ ,
    \new_[1654]_ , \new_[1655]_ , \new_[1656]_ , \new_[1657]_ ,
    \new_[1658]_ , \new_[1659]_ , \new_[1661]_ , \new_[1662]_ ,
    \new_[1663]_ , \new_[1664]_ , \new_[1666]_ , \new_[1667]_ ,
    \new_[1668]_ , \new_[1669]_ , \new_[1672]_ , \new_[1673]_ ,
    \new_[1674]_ , \new_[1675]_ , \new_[1676]_ , \new_[1677]_ ,
    \new_[1678]_ , \new_[1679]_ , \new_[1680]_ , \new_[1681]_ ,
    \new_[1682]_ , \new_[1683]_ , \new_[1684]_ , \new_[1685]_ ,
    \new_[1686]_ , \new_[1687]_ , \new_[1688]_ , \new_[1689]_ ,
    \new_[1690]_ , \new_[1691]_ , \new_[1692]_ , \new_[1693]_ ,
    \new_[1694]_ , \new_[1695]_ , \new_[1696]_ , \new_[1697]_ ,
    \new_[1698]_ , \new_[1699]_ , \new_[1700]_ , \new_[1701]_ ,
    \new_[1702]_ , \new_[1703]_ , \new_[1704]_ , \new_[1706]_ ,
    \new_[1707]_ , \new_[1709]_ , \new_[1710]_ , \new_[1711]_ ,
    \new_[1712]_ , \new_[1713]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1720]_ , \new_[1721]_ ,
    \new_[1722]_ , \new_[1723]_ , \new_[1724]_ , \new_[1729]_ ,
    \new_[1730]_ , \new_[1731]_ , \new_[1732]_ , \new_[1733]_ ,
    \new_[1734]_ , \new_[1735]_ , \new_[1736]_ , \new_[1737]_ ,
    \new_[1738]_ , \new_[1739]_ , \new_[1740]_ , \new_[1741]_ ,
    \new_[1742]_ , \new_[1743]_ , \new_[1744]_ , \new_[1745]_ ,
    \new_[1746]_ , \new_[1747]_ , \new_[1748]_ , \new_[1749]_ ,
    \new_[1750]_ , \new_[1751]_ , \new_[1752]_ , \new_[1753]_ ,
    \new_[1754]_ , \new_[1756]_ , \new_[1758]_ , \new_[1759]_ ,
    \new_[1760]_ , \new_[1761]_ , \new_[1762]_ , \new_[1763]_ ,
    \new_[1764]_ , \new_[1765]_ , \new_[1766]_ , \new_[1767]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1805]_ ,
    \new_[1806]_ , \new_[1807]_ , \new_[1808]_ , \new_[1809]_ ,
    \new_[1810]_ , \new_[1811]_ , \new_[1812]_ , \new_[1813]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1816]_ , \new_[1817]_ ,
    \new_[1818]_ , \new_[1819]_ , \new_[1820]_ , \new_[1821]_ ,
    \new_[1822]_ , \new_[1823]_ , \new_[1824]_ , \new_[1825]_ ,
    \new_[1826]_ , \new_[1827]_ , \new_[1828]_ , \new_[1829]_ ,
    \new_[1830]_ , \new_[1831]_ , \new_[1832]_ , \new_[1833]_ ,
    \new_[1834]_ , \new_[1835]_ , \new_[1836]_ , \new_[1837]_ ,
    \new_[1838]_ , \new_[1839]_ , \new_[1840]_ , \new_[1841]_ ,
    \new_[1843]_ , \new_[1844]_ , \new_[1845]_ , \new_[1846]_ ,
    \new_[1848]_ , \new_[1849]_ , \new_[1850]_ , \new_[1851]_ ,
    \new_[1852]_ , \new_[1853]_ , \new_[1854]_ , \new_[1855]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1932]_ , \new_[1933]_ ,
    \new_[1934]_ , \new_[1935]_ , \new_[1936]_ , \new_[1937]_ ,
    \new_[1938]_ , \new_[1939]_ , \new_[1940]_ , \new_[1941]_ ,
    \new_[1942]_ , \new_[1943]_ , \new_[1944]_ , \new_[1945]_ ,
    \new_[1946]_ , \new_[1947]_ , \new_[1948]_ , \new_[1949]_ ,
    \new_[1950]_ , \new_[1951]_ , \new_[1952]_ , \new_[1953]_ ,
    \new_[1954]_ , \new_[1955]_ , \new_[1957]_ , \new_[1958]_ ,
    \new_[1959]_ , \new_[1960]_ , \new_[1961]_ , \new_[1962]_ ,
    \new_[1963]_ , \new_[1964]_ , \new_[1965]_ , \new_[1966]_ ,
    \new_[1967]_ , \new_[1968]_ , \new_[1969]_ , \new_[1970]_ ,
    \new_[1971]_ , \new_[1972]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1993]_ ,
    \new_[1994]_ , \new_[2004]_ , \new_[2005]_ , \new_[2006]_ ,
    \new_[2007]_ , \new_[2008]_ , \new_[2009]_ , \new_[2010]_ ,
    \new_[2011]_ , \new_[2012]_ , \new_[2013]_ , \new_[2014]_ ,
    \new_[2015]_ , \new_[2017]_ , \new_[2025]_ , \new_[2026]_ ,
    \new_[2027]_ , \new_[2028]_ , \new_[2029]_ , \new_[2030]_ ,
    \new_[2031]_ , \new_[2032]_ , \new_[2033]_ , \new_[2034]_ ,
    \new_[2035]_ , \new_[2036]_ , \new_[2037]_ , \new_[2038]_ ,
    \new_[2039]_ , \new_[2040]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2060]_ , \new_[2061]_ ,
    \new_[2062]_ , \new_[2063]_ , \new_[2064]_ , \new_[2066]_ ,
    \new_[2067]_ , \new_[2068]_ , \new_[2069]_ , \new_[2070]_ ,
    \new_[2080]_ , \new_[2081]_ , \new_[2082]_ , \new_[2083]_ ,
    \new_[2084]_ , \new_[2085]_ , \new_[2086]_ , \new_[2087]_ ,
    \new_[2088]_ , \new_[2089]_ , \new_[2090]_ , \new_[2091]_ ,
    \new_[2092]_ , \new_[2093]_ , \new_[2094]_ , \new_[2095]_ ,
    \new_[2131]_ , \new_[2132]_ , \new_[2133]_ , \new_[2134]_ ,
    \new_[2135]_ , \new_[2136]_ , \new_[2137]_ , \new_[2138]_ ,
    \new_[2139]_ , \new_[2142]_ , \new_[2143]_ , \new_[2151]_ ,
    \new_[2152]_ , \new_[2153]_ , \new_[2154]_ , \new_[2155]_ ,
    \new_[2156]_ , \new_[2157]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2196]_ , \new_[2197]_ ,
    \new_[2198]_ , \new_[2199]_ , \new_[2200]_ , \new_[2201]_ ,
    \new_[2202]_ , \new_[2203]_ , \new_[2209]_ , \new_[2210]_ ,
    \new_[2211]_ , \new_[2212]_ , \new_[2213]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2224]_ , \new_[2225]_ ,
    \new_[2226]_ , \new_[2227]_ , \new_[2264]_ , \new_[2265]_ ,
    \new_[2266]_ , \new_[2267]_ , \new_[2271]_ , \new_[2273]_ ,
    \new_[2275]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2289]_ ,
    \new_[2290]_ , \new_[2291]_ , \new_[2301]_ , \new_[2302]_ ,
    \new_[2344]_ , \new_[2345]_ , \new_[2346]_ , \new_[2347]_ ,
    \new_[2348]_ , \new_[2349]_ , \new_[2350]_ , \new_[2351]_ ,
    \new_[2352]_ , \new_[2353]_ , \new_[2354]_ , \new_[2355]_ ,
    \new_[2356]_ , \new_[2357]_ , \new_[2358]_ , \new_[2359]_ ,
    \new_[2362]_ , \new_[2363]_ , \new_[2364]_ , \new_[2365]_ ,
    \new_[2366]_ , \new_[2367]_ , \new_[2368]_ , \new_[2411]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2439]_ , \new_[2440]_ , \new_[2441]_ ,
    \new_[2442]_ , \new_[2461]_ , \new_[2501]_ , \new_[2502]_ ,
    \new_[2503]_ , \new_[2504]_ , \new_[2505]_ , \new_[2506]_ ,
    \new_[2507]_ , \new_[2508]_ , \new_[2509]_ , \new_[2510]_ ,
    \new_[2511]_ , \new_[2512]_ , \new_[2513]_ , \new_[2514]_ ,
    \new_[2515]_ , \new_[2516]_ , \new_[2517]_ , \new_[2518]_ ,
    \new_[2519]_ , \new_[2520]_ , \new_[2521]_ , \new_[2522]_ ,
    \new_[2523]_ , \new_[2524]_ , \new_[2525]_ , \new_[2526]_ ,
    \new_[2527]_ , \new_[2528]_ , \new_[2529]_ , \new_[2530]_ ,
    \new_[2531]_ , \new_[2532]_ , \new_[2533]_ , \new_[2534]_ ,
    \new_[2535]_ , \new_[2536]_ , \new_[2537]_ , \new_[2538]_ ,
    \new_[2539]_ , \new_[2540]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2543]_ , \new_[2544]_ , \new_[2545]_ , \new_[2546]_ ,
    \new_[2547]_ , \new_[2548]_ , \new_[2549]_ , \new_[2550]_ ,
    \new_[2551]_ , \new_[2552]_ , \new_[2557]_ , \new_[2558]_ ,
    \new_[2559]_ , \new_[2568]_ , \new_[2569]_ , \new_[2570]_ ,
    \new_[2571]_ , \new_[2572]_ , \new_[2573]_ , \new_[2574]_ ,
    \new_[2575]_ , \new_[2576]_ , \new_[2577]_ , \new_[2578]_ ,
    \new_[2579]_ , \new_[2580]_ , \new_[2581]_ , \new_[2582]_ ,
    \new_[2583]_ , \new_[2584]_ , \new_[2585]_ , \new_[2586]_ ,
    \new_[2587]_ , \new_[2588]_ , \new_[2589]_ , \new_[2590]_ ,
    \new_[2591]_ , \new_[2592]_ , \new_[2593]_ , \new_[2594]_ ,
    \new_[2595]_ , \new_[2596]_ , \new_[2597]_ , \new_[2598]_ ,
    \new_[2599]_ , \new_[2600]_ , \new_[2601]_ , \new_[2602]_ ,
    \new_[2603]_ , \new_[2604]_ , \new_[2605]_ , \new_[2606]_ ,
    \new_[2607]_ , \new_[2608]_ , \new_[2609]_ , \new_[2610]_ ,
    \new_[2611]_ , \new_[2612]_ , \new_[2613]_ , \new_[2614]_ ,
    \new_[2615]_ , \new_[2616]_ , \new_[2617]_ , \new_[2618]_ ,
    \new_[2619]_ , \new_[2620]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2626]_ , \new_[2627]_ ,
    \new_[2628]_ , \new_[2629]_ , \new_[2630]_ , \new_[2631]_ ,
    \new_[2632]_ , \new_[2633]_ , \new_[2634]_ , \new_[2635]_ ,
    \new_[2636]_ , \new_[2637]_ , \new_[2638]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2641]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2650]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2653]_ , \new_[2654]_ , \new_[2655]_ ,
    \new_[2656]_ , \new_[2657]_ , \new_[2658]_ , \new_[2659]_ ,
    \new_[2660]_ , \new_[2661]_ , \new_[2662]_ , \new_[2663]_ ,
    \new_[2664]_ , \new_[2665]_ , \new_[2666]_ , \new_[2675]_ ,
    \new_[2676]_ , \new_[2684]_ , \new_[2685]_ , \new_[2686]_ ,
    \new_[2687]_ , \new_[2688]_ , \new_[2689]_ , \new_[2690]_ ,
    \new_[2691]_ , \new_[2692]_ , \new_[2693]_ , \new_[2694]_ ,
    \new_[2695]_ , \new_[2696]_ , \new_[2697]_ , \new_[2698]_ ,
    \new_[2699]_ , \new_[2700]_ , \new_[2701]_ , \new_[2702]_ ,
    \new_[2703]_ , \new_[2704]_ , \new_[2705]_ , \new_[2706]_ ,
    \new_[2707]_ , \new_[2708]_ , \new_[2709]_ , \new_[2710]_ ,
    \new_[2711]_ , \new_[2712]_ , \new_[2713]_ , \new_[2714]_ ,
    \new_[2715]_ , \new_[2716]_ , \new_[2717]_ , \new_[2718]_ ,
    \new_[2719]_ , \new_[2720]_ , \new_[2721]_ , \new_[2722]_ ,
    \new_[2723]_ , \new_[2724]_ , \new_[2725]_ , \new_[2726]_ ,
    \new_[2727]_ , \new_[2728]_ , \new_[2729]_ , \new_[2730]_ ,
    \new_[2731]_ , \new_[2732]_ , \new_[2733]_ , \new_[2734]_ ,
    \new_[2735]_ , \new_[2736]_ , \new_[2737]_ , \new_[2738]_ ,
    \new_[2739]_ , \new_[2740]_ , \new_[2741]_ , \new_[2742]_ ,
    \new_[2743]_ , \new_[2744]_ , \new_[2745]_ , \new_[2746]_ ,
    \new_[2747]_ , \new_[2748]_ , \new_[2749]_ , \new_[2750]_ ,
    \new_[2751]_ , \new_[2752]_ , \new_[2753]_ , \new_[2754]_ ,
    \new_[2755]_ , \new_[2756]_ , \new_[2757]_ , \new_[2758]_ ,
    \new_[2759]_ , \new_[2760]_ , \new_[2761]_ , \new_[2762]_ ,
    \new_[2763]_ , \new_[2764]_ , \new_[2765]_ , \new_[2766]_ ,
    \new_[2767]_ , \new_[2768]_ , \new_[2769]_ , \new_[2770]_ ,
    \new_[2771]_ , \new_[2772]_ , \new_[2773]_ , \new_[2774]_ ,
    \new_[2775]_ , \new_[2776]_ , \new_[2777]_ , \new_[2778]_ ,
    \new_[2779]_ , \new_[2780]_ , \new_[2781]_ , \new_[2782]_ ,
    \new_[2783]_ , \new_[2784]_ , \new_[2785]_ , \new_[2786]_ ,
    \new_[2787]_ , \new_[2788]_ , \new_[2789]_ , \new_[2790]_ ,
    \new_[2791]_ , \new_[2792]_ , \new_[2793]_ , \new_[2794]_ ,
    \new_[2795]_ , \new_[2796]_ , \new_[2797]_ , \new_[2798]_ ,
    \new_[2799]_ , \new_[2800]_ , \new_[2801]_ , \new_[2802]_ ,
    \new_[2803]_ , \new_[2804]_ , \new_[2805]_ , \new_[2806]_ ,
    \new_[2807]_ , \new_[2808]_ , \new_[2809]_ , \new_[2810]_ ,
    \new_[2827]_ , \new_[2828]_ , \new_[2829]_ , \new_[2830]_ ,
    \new_[2831]_ , \new_[2833]_ , \new_[2834]_ , \new_[2835]_ ,
    \new_[2839]_ , \new_[2840]_ , \new_[2841]_ , \new_[2842]_ ,
    \new_[2843]_ , \new_[2844]_ , \new_[2845]_ , \new_[2846]_ ,
    \new_[2847]_ , \new_[2848]_ , \new_[2849]_ , \new_[2850]_ ,
    \new_[2851]_ , \new_[2852]_ , \new_[2853]_ , \new_[2854]_ ,
    \new_[2855]_ , \new_[2856]_ , \new_[2857]_ , \new_[2858]_ ,
    \new_[2859]_ , \new_[2860]_ , \new_[2861]_ , \new_[2862]_ ,
    \new_[2863]_ , \new_[2864]_ , \new_[2865]_ , \new_[2866]_ ,
    \new_[2867]_ , \new_[2868]_ , \new_[2869]_ , \new_[2870]_ ,
    \new_[2871]_ , \new_[2872]_ , \new_[2873]_ , \new_[2874]_ ,
    \new_[2875]_ , \new_[2876]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2880]_ , \new_[2881]_ , \new_[2882]_ ,
    \new_[2883]_ , \new_[2884]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2888]_ , \new_[2889]_ , \new_[2890]_ ,
    \new_[2891]_ , \new_[2892]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2896]_ , \new_[2897]_ , \new_[2898]_ ,
    \new_[2899]_ , \new_[2900]_ , \new_[2901]_ , \new_[2902]_ ,
    \new_[2903]_ , \new_[2904]_ , \new_[2905]_ , \new_[2906]_ ,
    \new_[2907]_ , \new_[2908]_ , \new_[2909]_ , \new_[2910]_ ,
    \new_[2911]_ , \new_[2912]_ , \new_[2913]_ , \new_[2914]_ ,
    \new_[2915]_ , \new_[2916]_ , \new_[2917]_ , \new_[2918]_ ,
    \new_[2923]_ , \new_[2924]_ , \new_[2925]_ , \new_[2926]_ ,
    \new_[2931]_ , \new_[2932]_ , \new_[2933]_ , \new_[2934]_ ,
    \new_[2935]_ , \new_[2936]_ , \new_[2937]_ , \new_[2938]_ ,
    \new_[2939]_ , \new_[2940]_ , \new_[2941]_ , \new_[2942]_ ,
    \new_[2943]_ , \new_[2944]_ , \new_[2945]_ , \new_[2946]_ ,
    \new_[2947]_ , \new_[2948]_ , \new_[2949]_ , \new_[2950]_ ,
    \new_[2951]_ , \new_[2952]_ , \new_[2953]_ , \new_[2954]_ ,
    \new_[2955]_ , \new_[2956]_ , \new_[2957]_ , \new_[2958]_ ,
    \new_[2959]_ , \new_[2960]_ , \new_[2961]_ , \new_[2962]_ ,
    \new_[2963]_ , \new_[2964]_ , \new_[2965]_ , \new_[2966]_ ,
    \new_[2967]_ , \new_[2968]_ , \new_[2969]_ , \new_[2970]_ ,
    \new_[2971]_ , \new_[2972]_ , \new_[2973]_ , \new_[2974]_ ,
    \new_[2975]_ , \new_[2993]_ , \new_[2994]_ , \new_[2995]_ ,
    \new_[2996]_ , \new_[2997]_ , \new_[2998]_ , \new_[2999]_ ,
    \new_[3000]_ , \new_[3001]_ , \new_[3002]_ , \new_[3003]_ ,
    \new_[3004]_ , \new_[3005]_ , \new_[3006]_ , \new_[3007]_ ,
    \new_[3008]_ , \new_[3009]_ , \new_[3010]_ , \new_[3011]_ ,
    \new_[3012]_ , \new_[3013]_ , \new_[3014]_ , \new_[3015]_ ,
    \new_[3016]_ , \new_[3017]_ , \new_[3018]_ , \new_[3019]_ ,
    \new_[3020]_ , \new_[3021]_ , \new_[3022]_ , \new_[3023]_ ,
    \new_[3024]_ , \new_[3025]_ , \new_[3026]_ , \new_[3027]_ ,
    \new_[3028]_ , \new_[3029]_ , \new_[3030]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3033]_ , \new_[3034]_ , \new_[3035]_ ,
    \new_[3036]_ , \new_[3037]_ , \new_[3038]_ , \new_[3039]_ ,
    \new_[3040]_ , \new_[3041]_ , \new_[3042]_ , \new_[3043]_ ,
    \new_[3044]_ , \new_[3045]_ , \new_[3050]_ , \new_[3051]_ ,
    \new_[3052]_ , \new_[3053]_ , \new_[3054]_ , \new_[3055]_ ,
    \new_[3056]_ , \new_[3057]_ , \new_[3058]_ , \new_[3059]_ ,
    \new_[3060]_ , \new_[3061]_ , \new_[3062]_ , \new_[3063]_ ,
    \new_[3064]_ , \new_[3065]_ , \new_[3066]_ , \new_[3067]_ ,
    \new_[3068]_ , \new_[3069]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3073]_ , \new_[3074]_ , \new_[3075]_ ,
    \new_[3076]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3090]_ , \new_[3091]_ ,
    \new_[3092]_ , \new_[3093]_ , \new_[3094]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ,
    \new_[3100]_ , \new_[3101]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3105]_ , \new_[3106]_ , \new_[3107]_ ,
    \new_[3108]_ , \new_[3109]_ , \new_[3110]_ , \new_[3111]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3114]_ , \new_[3115]_ ,
    \new_[3116]_ , \new_[3117]_ , \new_[3118]_ , \new_[3119]_ ,
    \new_[3120]_ , \new_[3121]_ , \new_[3122]_ , \new_[3123]_ ,
    \new_[3124]_ , \new_[3125]_ , \new_[3126]_ , \new_[3127]_ ,
    \new_[3128]_ , \new_[3129]_ , \new_[3130]_ , \new_[3131]_ ,
    \new_[3132]_ , \new_[3133]_ , \new_[3134]_ , \new_[3135]_ ,
    \new_[3136]_ , \new_[3137]_ , \new_[3138]_ , \new_[3139]_ ,
    \new_[3140]_ , \new_[3141]_ , \new_[3142]_ , \new_[3143]_ ,
    \new_[3144]_ , \new_[3145]_ , \new_[3146]_ , \new_[3147]_ ,
    \new_[3148]_ , \new_[3149]_ , \new_[3150]_ , \new_[3151]_ ,
    \new_[3152]_ , \new_[3153]_ , \new_[3154]_ , \new_[3155]_ ,
    \new_[3156]_ , \new_[3157]_ , \new_[3158]_ , \new_[3159]_ ,
    \new_[3160]_ , \new_[3161]_ , \new_[3162]_ , \new_[3163]_ ,
    \new_[3164]_ , \new_[3165]_ , \new_[3166]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3169]_ , \new_[3170]_ , \new_[3171]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3177]_ , \new_[3178]_ , \new_[3179]_ ,
    \new_[3180]_ , \new_[3181]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3184]_ , \new_[3185]_ , \new_[3186]_ , \new_[3187]_ ,
    \new_[3188]_ , \new_[3189]_ , \new_[3190]_ , \new_[3191]_ ,
    \new_[3192]_ , \new_[3194]_ , \new_[3196]_ , \new_[3197]_ ,
    \new_[3199]_ , \new_[3201]_ , \new_[3202]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3208]_ , \new_[3209]_ ,
    \new_[3211]_ , \new_[3212]_ , \new_[3213]_ , \new_[3214]_ ,
    \new_[3216]_ , \new_[3217]_ , \new_[3218]_ , \new_[3219]_ ,
    \new_[3220]_ , \new_[3221]_ , \new_[3222]_ , \new_[3223]_ ,
    \new_[3224]_ , \new_[3225]_ , \new_[3226]_ , \new_[3227]_ ,
    \new_[3228]_ , \new_[3229]_ , \new_[3230]_ , \new_[3231]_ ,
    \new_[3232]_ , \new_[3233]_ , \new_[3234]_ , \new_[3235]_ ,
    \new_[3236]_ , \new_[3237]_ , \new_[3238]_ , \new_[3239]_ ,
    \new_[3240]_ , \new_[3241]_ , \new_[3242]_ , \new_[3243]_ ,
    \new_[3244]_ , \new_[3245]_ , \new_[3246]_ , \new_[3247]_ ,
    \new_[3248]_ , \new_[3249]_ , \new_[3250]_ , \new_[3251]_ ,
    \new_[3252]_ , \new_[3253]_ , \new_[3254]_ , \new_[3255]_ ,
    \new_[3256]_ , \new_[3257]_ , \new_[3258]_ , \new_[3259]_ ,
    \new_[3260]_ , \new_[3261]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3265]_ , \new_[3266]_ , \new_[3267]_ ,
    \new_[3268]_ , \new_[3269]_ , \new_[3270]_ , \new_[3271]_ ,
    \new_[3272]_ , \new_[3273]_ , \new_[3274]_ , \new_[3275]_ ,
    \new_[3276]_ , \new_[3277]_ , \new_[3278]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3282]_ , \new_[3283]_ ,
    \new_[3284]_ , \new_[3285]_ , \new_[3286]_ , \new_[3287]_ ,
    \new_[3288]_ , \new_[3289]_ , \new_[3290]_ , \new_[3291]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3302]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3306]_ , \new_[3307]_ ,
    \new_[3308]_ , \new_[3309]_ , \new_[3310]_ , \new_[3315]_ ,
    \new_[3316]_ , \new_[3317]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3321]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3324]_ , \new_[3325]_ , \new_[3326]_ , \new_[3327]_ ,
    \new_[3328]_ , \new_[3329]_ , \new_[3330]_ , \new_[3331]_ ,
    \new_[3332]_ , \new_[3333]_ , \new_[3334]_ , \new_[3335]_ ,
    \new_[3336]_ , \new_[3337]_ , \new_[3338]_ , \new_[3339]_ ,
    \new_[3340]_ , \new_[3341]_ , \new_[3342]_ , \new_[3343]_ ,
    \new_[3344]_ , \new_[3345]_ , \new_[3346]_ , \new_[3347]_ ,
    \new_[3348]_ , \new_[3349]_ , \new_[3350]_ , \new_[3351]_ ,
    \new_[3352]_ , \new_[3353]_ , \new_[3354]_ , \new_[3355]_ ,
    \new_[3356]_ , \new_[3357]_ , \new_[3358]_ , \new_[3359]_ ,
    \new_[3360]_ , \new_[3361]_ , \new_[3362]_ , \new_[3363]_ ,
    \new_[3364]_ , \new_[3365]_ , \new_[3366]_ , \new_[3367]_ ,
    \new_[3368]_ , \new_[3369]_ , \new_[3370]_ , \new_[3371]_ ,
    \new_[3372]_ , \new_[3373]_ , \new_[3374]_ , \new_[3375]_ ,
    \new_[3376]_ , \new_[3377]_ , \new_[3378]_ , \new_[3379]_ ,
    \new_[3380]_ , \new_[3381]_ , \new_[3382]_ , \new_[3383]_ ,
    \new_[3384]_ , \new_[3385]_ , \new_[3386]_ , \new_[3387]_ ,
    \new_[3388]_ , \new_[3389]_ , \new_[3390]_ , \new_[3391]_ ,
    \new_[3392]_ , \new_[3393]_ , \new_[3394]_ , \new_[3395]_ ,
    \new_[3396]_ , \new_[3397]_ , \new_[3398]_ , \new_[3399]_ ,
    \new_[3400]_ , \new_[3401]_ , \new_[3402]_ , \new_[3403]_ ,
    \new_[3404]_ , \new_[3405]_ , \new_[3406]_ , \new_[3407]_ ,
    \new_[3408]_ , \new_[3409]_ , \new_[3410]_ , \new_[3411]_ ,
    \new_[3412]_ , \new_[3413]_ , \new_[3414]_ , \new_[3415]_ ,
    \new_[3416]_ , \new_[3417]_ , \new_[3418]_ , \new_[3419]_ ,
    \new_[3420]_ , \new_[3421]_ , \new_[3422]_ , \new_[3423]_ ,
    \new_[3424]_ , \new_[3425]_ , \new_[3426]_ , \new_[3427]_ ,
    \new_[3428]_ , \new_[3429]_ , \new_[3430]_ , \new_[3431]_ ,
    \new_[3432]_ , \new_[3433]_ , \new_[3434]_ , \new_[3435]_ ,
    \new_[3436]_ , \new_[3437]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3441]_ , \new_[3442]_ , \new_[3443]_ ,
    \new_[3444]_ , \new_[3445]_ , \new_[3446]_ , \new_[3447]_ ,
    \new_[3448]_ , \new_[3449]_ , \new_[3450]_ , \new_[3451]_ ,
    \new_[3452]_ , \new_[3453]_ , \new_[3454]_ , \new_[3455]_ ,
    \new_[3456]_ , \new_[3457]_ , \new_[3458]_ , \new_[3459]_ ,
    \new_[3460]_ , \new_[3461]_ , \new_[3462]_ , \new_[3463]_ ,
    \new_[3464]_ , \new_[3465]_ , \new_[3466]_ , \new_[3467]_ ,
    \new_[3468]_ , \new_[3469]_ , \new_[3470]_ , \new_[3471]_ ,
    \new_[3472]_ , \new_[3473]_ , \new_[3474]_ , \new_[3475]_ ,
    \new_[3476]_ , \new_[3477]_ , \new_[3478]_ , \new_[3479]_ ,
    \new_[3480]_ , \new_[3481]_ , \new_[3482]_ , \new_[3483]_ ,
    \new_[3484]_ , \new_[3485]_ , \new_[3486]_ , \new_[3487]_ ,
    \new_[3488]_ , \new_[3489]_ , \new_[3490]_ , \new_[3491]_ ,
    \new_[3492]_ , \new_[3493]_ , \new_[3494]_ , \new_[3495]_ ,
    \new_[3496]_ , \new_[3497]_ , \new_[3498]_ , \new_[3499]_ ,
    \new_[3500]_ , \new_[3501]_ , \new_[3502]_ , \new_[3503]_ ,
    \new_[3504]_ , \new_[3505]_ , \new_[3506]_ , \new_[3507]_ ,
    \new_[3508]_ , \new_[3513]_ , \new_[3514]_ , \new_[3515]_ ,
    \new_[3516]_ , \new_[3517]_ , \new_[3518]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3521]_ , \new_[3522]_ , \new_[3523]_ ,
    \new_[3524]_ , \new_[3525]_ , \new_[3526]_ , \new_[3527]_ ,
    \new_[3528]_ , \new_[3529]_ , \new_[3530]_ , \new_[3531]_ ,
    \new_[3532]_ , \new_[3533]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3536]_ , \new_[3537]_ , \new_[3538]_ , \new_[3539]_ ,
    \new_[3540]_ , \new_[3549]_ , \new_[3550]_ , \new_[3551]_ ,
    \new_[3552]_ , \new_[3553]_ , \new_[3554]_ , \new_[3555]_ ,
    \new_[3556]_ , \new_[3557]_ , \new_[3558]_ , \new_[3559]_ ,
    \new_[3560]_ , \new_[3561]_ , \new_[3562]_ , \new_[3563]_ ,
    \new_[3564]_ , \new_[3565]_ , \new_[3566]_ , \new_[3567]_ ,
    \new_[3568]_ , \new_[3569]_ , \new_[3570]_ , \new_[3571]_ ,
    \new_[3572]_ , \new_[3573]_ , \new_[3574]_ , \new_[3575]_ ,
    \new_[3576]_ , \new_[3577]_ , \new_[3578]_ , \new_[3579]_ ,
    \new_[3580]_ , \new_[3581]_ , \new_[3582]_ , \new_[3583]_ ,
    \new_[3584]_ , \new_[3585]_ , \new_[3586]_ , \new_[3587]_ ,
    \new_[3588]_ , \new_[3589]_ , \new_[3590]_ , \new_[3591]_ ,
    \new_[3592]_ , \new_[3593]_ , \new_[3594]_ , \new_[3595]_ ,
    \new_[3596]_ , \new_[3597]_ , \new_[3598]_ , \new_[3599]_ ,
    \new_[3600]_ , \new_[3601]_ , \new_[3602]_ , \new_[3603]_ ,
    \new_[3604]_ , \new_[3605]_ , \new_[3606]_ , \new_[3607]_ ,
    \new_[3608]_ , \new_[3609]_ , \new_[3610]_ , \new_[3611]_ ,
    \new_[3612]_ , \new_[3613]_ , \new_[3614]_ , \new_[3615]_ ,
    \new_[3616]_ , \new_[3617]_ , \new_[3618]_ , \new_[3619]_ ,
    \new_[3620]_ , \new_[3621]_ , \new_[3622]_ , \new_[3623]_ ,
    \new_[3624]_ , \new_[3625]_ , \new_[3626]_ , \new_[3627]_ ,
    \new_[3628]_ , \new_[3629]_ , \new_[3630]_ , \new_[3631]_ ,
    \new_[3632]_ , \new_[3633]_ , \new_[3642]_ , \new_[3647]_ ,
    \new_[3648]_ , \new_[3649]_ , \new_[3650]_ , \new_[3651]_ ,
    \new_[3652]_ , \new_[3653]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3656]_ , \new_[3657]_ , \new_[3658]_ , \new_[3659]_ ,
    \new_[3660]_ , \new_[3661]_ , \new_[3662]_ , \new_[3663]_ ,
    \new_[3664]_ , \new_[3665]_ , \new_[3666]_ , \new_[3667]_ ,
    \new_[3668]_ , \new_[3669]_ , \new_[3670]_ , \new_[3671]_ ,
    \new_[3672]_ , \new_[3673]_ , \new_[3674]_ , \new_[3675]_ ,
    \new_[3680]_ , \new_[3681]_ , \new_[3682]_ , \new_[3683]_ ,
    \new_[3684]_ , \new_[3685]_ , \new_[3686]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3690]_ , \new_[3691]_ ,
    \new_[3692]_ , \new_[3693]_ , \new_[3694]_ , \new_[3695]_ ,
    \new_[3696]_ , \new_[3697]_ , \new_[3698]_ , \new_[3699]_ ,
    \new_[3700]_ , \new_[3701]_ , \new_[3702]_ , \new_[3703]_ ,
    \new_[3704]_ , \new_[3705]_ , \new_[3706]_ , \new_[3707]_ ,
    \new_[3708]_ , \new_[3709]_ , \new_[3710]_ , \new_[3711]_ ,
    \new_[3712]_ , \new_[3713]_ , \new_[3714]_ , \new_[3715]_ ,
    \new_[3716]_ , \new_[3717]_ , \new_[3718]_ , \new_[3719]_ ,
    \new_[3720]_ , \new_[3721]_ , \new_[3722]_ , \new_[3723]_ ,
    \new_[3724]_ , \new_[3725]_ , \new_[3726]_ , \new_[3727]_ ,
    \new_[3728]_ , \new_[3729]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3732]_ , \new_[3733]_ , \new_[3734]_ , \new_[3735]_ ,
    \new_[3736]_ , \new_[3737]_ , \new_[3738]_ , \new_[3739]_ ,
    \new_[3740]_ , \new_[3741]_ , \new_[3742]_ , \new_[3743]_ ,
    \new_[3744]_ , \new_[3745]_ , \new_[3746]_ , \new_[3747]_ ,
    \new_[3748]_ , \new_[3749]_ , \new_[3750]_ , \new_[3751]_ ,
    \new_[3752]_ , \new_[3753]_ , \new_[3754]_ , \new_[3755]_ ,
    \new_[3756]_ , \new_[3757]_ , \new_[3758]_ , \new_[3759]_ ,
    \new_[3760]_ , \new_[3761]_ , \new_[3762]_ , \new_[3763]_ ,
    \new_[3764]_ , \new_[3765]_ , \new_[3766]_ , \new_[3767]_ ,
    \new_[3768]_ , \new_[3769]_ , \new_[3770]_ , \new_[3771]_ ,
    \new_[3772]_ , \new_[3773]_ , \new_[3774]_ , \new_[3775]_ ,
    \new_[3776]_ , \new_[3777]_ , \new_[3778]_ , \new_[3779]_ ,
    \new_[3780]_ , \new_[3781]_ , \new_[3782]_ , \new_[3783]_ ,
    \new_[3784]_ , \new_[3785]_ , \new_[3786]_ , \new_[3787]_ ,
    \new_[3788]_ , \new_[3789]_ , \new_[3790]_ , \new_[3791]_ ,
    \new_[3792]_ , \new_[3793]_ , \new_[3794]_ , \new_[3795]_ ,
    \new_[3796]_ , \new_[3797]_ , \new_[3798]_ , \new_[3799]_ ,
    \new_[3800]_ , \new_[3801]_ , \new_[3802]_ , \new_[3803]_ ,
    \new_[3804]_ , \new_[3805]_ , \new_[3806]_ , \new_[3807]_ ,
    \new_[3808]_ , \new_[3809]_ , \new_[3810]_ , \new_[3811]_ ,
    \new_[3812]_ , \new_[3813]_ , \new_[3814]_ , \new_[3815]_ ,
    \new_[3816]_ , \new_[3821]_ , \new_[3822]_ , \new_[3823]_ ,
    \new_[3824]_ , \new_[3825]_ , \new_[3826]_ , \new_[3827]_ ,
    \new_[3828]_ , \new_[3829]_ , \new_[3830]_ , \new_[3831]_ ,
    \new_[3832]_ , \new_[3833]_ , \new_[3834]_ , \new_[3835]_ ,
    \new_[3836]_ , \new_[3837]_ , \new_[3838]_ , \new_[3839]_ ,
    \new_[3840]_ , \new_[3841]_ , \new_[3842]_ , \new_[3843]_ ,
    \new_[3844]_ , \new_[3845]_ , \new_[3846]_ , \new_[3847]_ ,
    \new_[3848]_ , \new_[3849]_ , \new_[3850]_ , \new_[3851]_ ,
    \new_[3852]_ , \new_[3853]_ , \new_[3854]_ , \new_[3855]_ ,
    \new_[3856]_ , \new_[3857]_ , \new_[3858]_ , \new_[3859]_ ,
    \new_[3860]_ , \new_[3861]_ , \new_[3862]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3865]_ , \new_[3866]_ , \new_[3867]_ ,
    \new_[3868]_ , \new_[3869]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3872]_ , \new_[3873]_ , \new_[3874]_ , \new_[3875]_ ,
    \new_[3876]_ , \new_[3877]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3880]_ , \new_[3881]_ , \new_[3882]_ , \new_[3883]_ ,
    \new_[3884]_ , \new_[3885]_ , \new_[3886]_ , \new_[3887]_ ,
    \new_[3888]_ , \new_[3889]_ , \new_[3890]_ , \new_[3891]_ ,
    \new_[3892]_ , \new_[3893]_ , \new_[3894]_ , \new_[3895]_ ,
    \new_[3896]_ , \new_[3897]_ , \new_[3898]_ , \new_[3899]_ ,
    \new_[3900]_ , \new_[3901]_ , \new_[3902]_ , \new_[3903]_ ,
    \new_[3904]_ , \new_[3905]_ , \new_[3906]_ , \new_[3907]_ ,
    \new_[3908]_ , \new_[3909]_ , \new_[3910]_ , \new_[3911]_ ,
    \new_[3912]_ , \new_[3913]_ , \new_[3914]_ , \new_[3915]_ ,
    \new_[3916]_ , \new_[3917]_ , \new_[3918]_ , \new_[3919]_ ,
    \new_[3920]_ , \new_[3921]_ , \new_[3922]_ , \new_[3923]_ ,
    \new_[3924]_ , \new_[3925]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3928]_ , \new_[3929]_ , \new_[3930]_ , \new_[3931]_ ,
    \new_[3932]_ , \new_[3933]_ , \new_[3934]_ , \new_[3935]_ ,
    \new_[3936]_ , \new_[3937]_ , \new_[3938]_ , \new_[3939]_ ,
    \new_[3940]_ , \new_[3941]_ , \new_[3942]_ , \new_[3943]_ ,
    \new_[3944]_ , \new_[3945]_ , \new_[3946]_ , \new_[3947]_ ,
    \new_[3948]_ , \new_[3949]_ , \new_[3950]_ , \new_[3951]_ ,
    \new_[3952]_ , \new_[3953]_ , \new_[3954]_ , \new_[3955]_ ,
    \new_[3956]_ , \new_[3957]_ , \new_[3958]_ , \new_[3959]_ ,
    \new_[3960]_ , \new_[3961]_ , \new_[3962]_ , \new_[3963]_ ,
    \new_[3964]_ , \new_[3965]_ , \new_[3966]_ , \new_[3967]_ ,
    \new_[3968]_ , \new_[3969]_ , \new_[3970]_ , \new_[3971]_ ,
    \new_[3972]_ , \new_[3973]_ , \new_[3974]_ , \new_[3975]_ ,
    \new_[3976]_ , \new_[3977]_ , \new_[3978]_ , \new_[3979]_ ,
    \new_[3980]_ , \new_[3981]_ , \new_[3982]_ , \new_[3983]_ ,
    \new_[3984]_ , \new_[3985]_ , \new_[3986]_ , \new_[3987]_ ,
    \new_[3988]_ , \new_[3989]_ , \new_[3990]_ , \new_[3991]_ ,
    \new_[3992]_ , \new_[3993]_ , \new_[3994]_ , \new_[3995]_ ,
    \new_[3996]_ , \new_[3997]_ , \new_[3998]_ , \new_[3999]_ ,
    \new_[4000]_ , \new_[4001]_ , \new_[4002]_ , \new_[4003]_ ,
    \new_[4004]_ , \new_[4005]_ , \new_[4006]_ , \new_[4007]_ ,
    \new_[4008]_ , \new_[4009]_ , \new_[4010]_ , \new_[4011]_ ,
    \new_[4012]_ , \new_[4013]_ , \new_[4014]_ , \new_[4015]_ ,
    \new_[4016]_ , \new_[4017]_ , \new_[4018]_ , \new_[4019]_ ,
    \new_[4020]_ , \new_[4021]_ , \new_[4022]_ , \new_[4023]_ ,
    \new_[4024]_ , \new_[4025]_ , \new_[4026]_ , \new_[4027]_ ,
    \new_[4028]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4033]_ , \new_[4034]_ , \new_[4035]_ ,
    \new_[4036]_ , \new_[4037]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4041]_ , \new_[4042]_ , \new_[4043]_ ,
    \new_[4044]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4048]_ , \new_[4049]_ , \new_[4050]_ , \new_[4051]_ ,
    \new_[4052]_ , \new_[4053]_ , \new_[4054]_ , \new_[4055]_ ,
    \new_[4056]_ , \new_[4057]_ , \new_[4058]_ , \new_[4059]_ ,
    \new_[4060]_ , \new_[4061]_ , \new_[4062]_ , \new_[4063]_ ,
    \new_[4064]_ , \new_[4065]_ , \new_[4066]_ , \new_[4067]_ ,
    \new_[4068]_ , \new_[4069]_ , \new_[4070]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4074]_ , \new_[4075]_ ,
    \new_[4076]_ , \new_[4077]_ , \new_[4078]_ , \new_[4079]_ ,
    \new_[4080]_ , \new_[4081]_ , \new_[4082]_ , \new_[4083]_ ,
    \new_[4084]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4088]_ , \new_[4089]_ , \new_[4090]_ , \new_[4091]_ ,
    \new_[4092]_ , \new_[4093]_ , \new_[4094]_ , \new_[4095]_ ,
    \new_[4096]_ , \new_[4097]_ , \new_[4098]_ , \new_[4099]_ ,
    \new_[4100]_ , \new_[4101]_ , \new_[4102]_ , \new_[4103]_ ,
    \new_[4104]_ , \new_[4105]_ , \new_[4106]_ , \new_[4107]_ ,
    \new_[4108]_ , \new_[4109]_ , \new_[4110]_ , \new_[4111]_ ,
    \new_[4112]_ , \new_[4113]_ , \new_[4114]_ , \new_[4115]_ ,
    \new_[4116]_ , \new_[4117]_ , \new_[4118]_ , \new_[4119]_ ,
    \new_[4120]_ , \new_[4121]_ , \new_[4122]_ , \new_[4123]_ ,
    \new_[4124]_ , \new_[4125]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4128]_ , \new_[4129]_ , \new_[4130]_ , \new_[4131]_ ,
    \new_[4132]_ , \new_[4133]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4136]_ , \new_[4137]_ , \new_[4138]_ , \new_[4139]_ ,
    \new_[4140]_ , \new_[4141]_ , \new_[4142]_ , \new_[4143]_ ,
    \new_[4144]_ , \new_[4149]_ , \new_[4150]_ , \new_[4151]_ ,
    \new_[4152]_ , \new_[4153]_ , \new_[4154]_ , \new_[4155]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4160]_ , \new_[4161]_ , \new_[4162]_ , \new_[4163]_ ,
    \new_[4164]_ , \new_[4165]_ , \new_[4166]_ , \new_[4167]_ ,
    \new_[4168]_ , \new_[4169]_ , \new_[4170]_ , \new_[4171]_ ,
    \new_[4172]_ , \new_[4173]_ , \new_[4174]_ , \new_[4175]_ ,
    \new_[4176]_ , \new_[4177]_ , \new_[4178]_ , \new_[4179]_ ,
    \new_[4180]_ , \new_[4181]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4184]_ , \new_[4185]_ , \new_[4186]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4192]_ , \new_[4193]_ , \new_[4194]_ , \new_[4195]_ ,
    \new_[4196]_ , \new_[4197]_ , \new_[4198]_ , \new_[4199]_ ,
    \new_[4200]_ , \new_[4201]_ , \new_[4202]_ , \new_[4203]_ ,
    \new_[4204]_ , \new_[4205]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4208]_ , \new_[4209]_ , \new_[4210]_ , \new_[4211]_ ,
    \new_[4212]_ , \new_[4213]_ , \new_[4214]_ , \new_[4215]_ ,
    \new_[4216]_ , \new_[4217]_ , \new_[4218]_ , \new_[4219]_ ,
    \new_[4220]_ , \new_[4221]_ , \new_[4222]_ , \new_[4223]_ ,
    \new_[4224]_ , \new_[4225]_ , \new_[4226]_ , \new_[4227]_ ,
    \new_[4228]_ , \new_[4229]_ , \new_[4230]_ , \new_[4232]_ ,
    \new_[4234]_ , \new_[4235]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4238]_ , \new_[4239]_ , \new_[4240]_ , \new_[4241]_ ,
    \new_[4242]_ , \new_[4243]_ , \new_[4244]_ , \new_[4245]_ ,
    \new_[4246]_ , \new_[4247]_ , \new_[4248]_ , \new_[4249]_ ,
    \new_[4250]_ , \new_[4251]_ , \new_[4252]_ , \new_[4253]_ ,
    \new_[4254]_ , \new_[4255]_ , \new_[4256]_ , \new_[4257]_ ,
    \new_[4258]_ , \new_[4259]_ , \new_[4260]_ , \new_[4261]_ ,
    \new_[4262]_ , \new_[4263]_ , \new_[4264]_ , \new_[4265]_ ,
    \new_[4266]_ , \new_[4267]_ , \new_[4268]_ , \new_[4269]_ ,
    \new_[4270]_ , \new_[4271]_ , \new_[4272]_ , \new_[4273]_ ,
    \new_[4274]_ , \new_[4275]_ , \new_[4276]_ , \new_[4277]_ ,
    \new_[4278]_ , \new_[4279]_ , \new_[4281]_ , \new_[4282]_ ,
    \new_[4283]_ , \new_[4284]_ , \new_[4285]_ , \new_[4286]_ ,
    \new_[4287]_ , \new_[4288]_ , \new_[4289]_ , \new_[4290]_ ,
    \new_[4291]_ , \new_[4292]_ , \new_[4293]_ , \new_[4294]_ ,
    \new_[4295]_ , \new_[4296]_ , \new_[4297]_ , \new_[4298]_ ,
    \new_[4299]_ , \new_[4300]_ , \new_[4301]_ , \new_[4302]_ ,
    \new_[4303]_ , \new_[4304]_ , \new_[4305]_ , \new_[4306]_ ,
    \new_[4307]_ , \new_[4308]_ , \new_[4309]_ , \new_[4310]_ ,
    \new_[4311]_ , \new_[4312]_ , \new_[4313]_ , \new_[4314]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4320]_ , \new_[4321]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4325]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4328]_ , \new_[4329]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4332]_ , \new_[4333]_ , \new_[4334]_ ,
    \new_[4335]_ , \new_[4336]_ , \new_[4337]_ , \new_[4338]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4341]_ , \new_[4342]_ ,
    \new_[4343]_ , \new_[4344]_ , \new_[4345]_ , \new_[4346]_ ,
    \new_[4347]_ , \new_[4348]_ , \new_[4349]_ , \new_[4350]_ ,
    \new_[4351]_ , \new_[4352]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4356]_ , \new_[4357]_ , \new_[4358]_ ,
    \new_[4359]_ , \new_[4360]_ , \new_[4361]_ , \new_[4362]_ ,
    \new_[4363]_ , \new_[4364]_ , \new_[4365]_ , \new_[4366]_ ,
    \new_[4367]_ , \new_[4368]_ , \new_[4369]_ , \new_[4370]_ ,
    \new_[4371]_ , \new_[4372]_ , \new_[4373]_ , \new_[4374]_ ,
    \new_[4375]_ , \new_[4376]_ , \new_[4377]_ , \new_[4378]_ ,
    \new_[4379]_ , \new_[4380]_ , \new_[4381]_ , \new_[4382]_ ,
    \new_[4383]_ , \new_[4384]_ , \new_[4385]_ , \new_[4386]_ ,
    \new_[4387]_ , \new_[4388]_ , \new_[4389]_ , \new_[4390]_ ,
    \new_[4391]_ , \new_[4392]_ , \new_[4393]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4396]_ , \new_[4397]_ , \new_[4398]_ ,
    \new_[4399]_ , \new_[4400]_ , \new_[4401]_ , \new_[4402]_ ,
    \new_[4403]_ , \new_[4404]_ , \new_[4405]_ , \new_[4406]_ ,
    \new_[4407]_ , \new_[4408]_ , \new_[4409]_ , \new_[4410]_ ,
    \new_[4411]_ , \new_[4412]_ , \new_[4413]_ , \new_[4414]_ ,
    \new_[4415]_ , \new_[4416]_ , \new_[4417]_ , \new_[4418]_ ,
    \new_[4419]_ , \new_[4420]_ , \new_[4421]_ , \new_[4422]_ ,
    \new_[4423]_ , \new_[4424]_ , \new_[4425]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4430]_ ,
    \new_[4431]_ , \new_[4432]_ , \new_[4433]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4437]_ , \new_[4438]_ ,
    \new_[4439]_ , \new_[4440]_ , \new_[4441]_ , \new_[4442]_ ,
    \new_[4443]_ , \new_[4444]_ , \new_[4445]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4448]_ , \new_[4449]_ , \new_[4450]_ ,
    \new_[4451]_ , \new_[4452]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4455]_ , \new_[4456]_ , \new_[4457]_ , \new_[4458]_ ,
    \new_[4459]_ , \new_[4460]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4464]_ , \new_[4465]_ , \new_[4466]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4471]_ , \new_[4472]_ , \new_[4473]_ , \new_[4474]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4477]_ , \new_[4478]_ ,
    \new_[4479]_ , \new_[4480]_ , \new_[4481]_ , \new_[4482]_ ,
    \new_[4483]_ , \new_[4484]_ , \new_[4485]_ , \new_[4486]_ ,
    \new_[4487]_ , \new_[4488]_ , \new_[4489]_ , \new_[4490]_ ,
    \new_[4491]_ , \new_[4492]_ , \new_[4493]_ , \new_[4494]_ ,
    \new_[4495]_ , \new_[4496]_ , \new_[4497]_ , \new_[4498]_ ,
    \new_[4499]_ , \new_[4500]_ , \new_[4501]_ , \new_[4502]_ ,
    \new_[4503]_ , \new_[4506]_ , \new_[4507]_ , \new_[4508]_ ,
    \new_[4509]_ , \new_[4510]_ , \new_[4511]_ , \new_[4512]_ ,
    \new_[4513]_ , \new_[4514]_ , \new_[4515]_ , \new_[4516]_ ,
    \new_[4517]_ , \new_[4518]_ , \new_[4519]_ , \new_[4520]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4523]_ , \new_[4524]_ ,
    \new_[4525]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4529]_ , \new_[4530]_ , \new_[4531]_ , \new_[4532]_ ,
    \new_[4533]_ , \new_[4534]_ , \new_[4535]_ , \new_[4536]_ ,
    \new_[4537]_ , \new_[4538]_ , \new_[4539]_ , \new_[4540]_ ,
    \new_[4541]_ , \new_[4542]_ , \new_[4543]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4547]_ , \new_[4548]_ ,
    \new_[4549]_ , \new_[4550]_ , \new_[4551]_ , \new_[4552]_ ,
    \new_[4553]_ , \new_[4554]_ , \new_[4555]_ , \new_[4556]_ ,
    \new_[4557]_ , \new_[4558]_ , \new_[4559]_ , \new_[4560]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4565]_ , \new_[4566]_ , \new_[4567]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4570]_ , \new_[4571]_ , \new_[4572]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4578]_ , \new_[4579]_ , \new_[4580]_ ,
    \new_[4581]_ , \new_[4582]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4586]_ , \new_[4587]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4590]_ , \new_[4591]_ , \new_[4592]_ ,
    \new_[4593]_ , \new_[4594]_ , \new_[4595]_ , \new_[4596]_ ,
    \new_[4597]_ , \new_[4598]_ , \new_[4599]_ , \new_[4600]_ ,
    \new_[4601]_ , \new_[4602]_ , \new_[4603]_ , \new_[4604]_ ,
    \new_[4605]_ , \new_[4606]_ , \new_[4607]_ , \new_[4608]_ ,
    \new_[4609]_ , \new_[4610]_ , \new_[4611]_ , \new_[4612]_ ,
    \new_[4613]_ , \new_[4614]_ , \new_[4615]_ , \new_[4616]_ ,
    \new_[4617]_ , \new_[4618]_ , \new_[4619]_ , \new_[4620]_ ,
    \new_[4621]_ , \new_[4622]_ , \new_[4623]_ , \new_[4624]_ ,
    \new_[4625]_ , \new_[4626]_ , \new_[4627]_ , \new_[4628]_ ,
    \new_[4629]_ , \new_[4630]_ , \new_[4631]_ , \new_[4632]_ ,
    \new_[4633]_ , \new_[4634]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4637]_ , \new_[4638]_ , \new_[4639]_ , \new_[4640]_ ,
    \new_[4641]_ , \new_[4642]_ , \new_[4643]_ , \new_[4644]_ ,
    \new_[4645]_ , \new_[4646]_ , \new_[4647]_ , \new_[4648]_ ,
    \new_[4649]_ , \new_[4650]_ , \new_[4651]_ , \new_[4652]_ ,
    \new_[4653]_ , \new_[4654]_ , \new_[4655]_ , \new_[4656]_ ,
    \new_[4657]_ , \new_[4658]_ , \new_[4659]_ , \new_[4660]_ ,
    \new_[4661]_ , \new_[4662]_ , \new_[4663]_ , \new_[4664]_ ,
    \new_[4665]_ , \new_[4666]_ , \new_[4667]_ , \new_[4668]_ ,
    \new_[4669]_ , \new_[4670]_ , \new_[4671]_ , \new_[4672]_ ,
    \new_[4673]_ , \new_[4674]_ , \new_[4675]_ , \new_[4676]_ ,
    \new_[4677]_ , \new_[4678]_ , \new_[4679]_ , \new_[4680]_ ,
    \new_[4681]_ , \new_[4682]_ , \new_[4683]_ , \new_[4684]_ ,
    \new_[4685]_ , \new_[4686]_ , \new_[4687]_ , \new_[4688]_ ,
    \new_[4689]_ , \new_[4690]_ , \new_[4691]_ , \new_[4692]_ ,
    \new_[4693]_ , \new_[4694]_ , \new_[4695]_ , \new_[4696]_ ,
    \new_[4697]_ , \new_[4698]_ , \new_[4699]_ , \new_[4700]_ ,
    \new_[4701]_ , \new_[4702]_ , \new_[4703]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4706]_ , \new_[4707]_ , \new_[4708]_ ,
    \new_[4709]_ , \new_[4710]_ , \new_[4711]_ , \new_[4712]_ ,
    \new_[4713]_ , \new_[4714]_ , \new_[4715]_ , \new_[4716]_ ,
    \new_[4717]_ , \new_[4718]_ , \new_[4719]_ , \new_[4720]_ ,
    \new_[4721]_ , \new_[4722]_ , \new_[4723]_ , \new_[4724]_ ,
    \new_[4725]_ , \new_[4726]_ , \new_[4727]_ , \new_[4728]_ ,
    \new_[4729]_ , \new_[4730]_ , \new_[4731]_ , \new_[4732]_ ,
    \new_[4733]_ , \new_[4734]_ , \new_[4735]_ , \new_[4736]_ ,
    \new_[4737]_ , \new_[4738]_ , \new_[4739]_ , \new_[4740]_ ,
    \new_[4741]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4746]_ , \new_[4747]_ , \new_[4748]_ ,
    \new_[4749]_ , \new_[4750]_ , \new_[4751]_ , \new_[4752]_ ,
    \new_[4753]_ , \new_[4754]_ , \new_[4755]_ , \new_[4756]_ ,
    \new_[4757]_ , \new_[4758]_ , \new_[4759]_ , \new_[4760]_ ,
    \new_[4761]_ , \new_[4762]_ , \new_[4763]_ , \new_[4764]_ ,
    \new_[4765]_ , \new_[4766]_ , \new_[4767]_ , \new_[4768]_ ,
    \new_[4769]_ , \new_[4770]_ , \new_[4771]_ , \new_[4772]_ ,
    \new_[4773]_ , \new_[4774]_ , \new_[4775]_ , \new_[4776]_ ,
    \new_[4777]_ , \new_[4778]_ , \new_[4779]_ , \new_[4780]_ ,
    \new_[4781]_ , \new_[4782]_ , \new_[4783]_ , \new_[4784]_ ,
    \new_[4785]_ , \new_[4786]_ , \new_[4787]_ , \new_[4788]_ ,
    \new_[4789]_ , \new_[4790]_ , \new_[4791]_ , \new_[4792]_ ,
    \new_[4793]_ , \new_[4794]_ , \new_[4795]_ , \new_[4796]_ ,
    \new_[4797]_ , \new_[4798]_ , \new_[4799]_ , \new_[4800]_ ,
    \new_[4801]_ , \new_[4802]_ , \new_[4803]_ , \new_[4804]_ ,
    \new_[4805]_ , \new_[4806]_ , \new_[4807]_ , \new_[4808]_ ,
    \new_[4809]_ , \new_[4810]_ , \new_[4811]_ , \new_[4812]_ ,
    \new_[4813]_ , \new_[4814]_ , \new_[4815]_ , \new_[4816]_ ,
    \new_[4817]_ , \new_[4818]_ , \new_[4819]_ , \new_[4820]_ ,
    \new_[4821]_ , \new_[4822]_ , \new_[4823]_ , \new_[4824]_ ,
    \new_[4825]_ , \new_[4826]_ , \new_[4827]_ , \new_[4828]_ ,
    \new_[4829]_ , \new_[4830]_ , \new_[4831]_ , \new_[4832]_ ,
    \new_[4833]_ , \new_[4834]_ , \new_[4835]_ , \new_[4836]_ ,
    \new_[4837]_ , \new_[4838]_ , \new_[4839]_ , \new_[4840]_ ,
    \new_[4841]_ , \new_[4842]_ , \new_[4843]_ , \new_[4844]_ ,
    \new_[4845]_ , \new_[4846]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4850]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4853]_ , \new_[4854]_ , \new_[4855]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4858]_ , \new_[4859]_ , \new_[4860]_ ,
    \new_[4861]_ , \new_[4862]_ , \new_[4863]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4869]_ , \new_[4870]_ , \new_[4871]_ , \new_[4872]_ ,
    \new_[4873]_ , \new_[4874]_ , \new_[4875]_ , \new_[4876]_ ,
    \new_[4877]_ , \new_[4878]_ , \new_[4879]_ , \new_[4880]_ ,
    \new_[4881]_ , \new_[4882]_ , \new_[4883]_ , \new_[4884]_ ,
    \new_[4885]_ , \new_[4886]_ , \new_[4887]_ , \new_[4888]_ ,
    \new_[4889]_ , \new_[4890]_ , \new_[4891]_ , \new_[4892]_ ,
    \new_[4893]_ , \new_[4894]_ , \new_[4895]_ , \new_[4896]_ ,
    \new_[4897]_ , \new_[4898]_ , \new_[4899]_ , \new_[4900]_ ,
    \new_[4901]_ , \new_[4902]_ , \new_[4903]_ , \new_[4904]_ ,
    \new_[4905]_ , \new_[4906]_ , \new_[4907]_ , \new_[4908]_ ,
    \new_[4909]_ , \new_[4910]_ , \new_[4911]_ , \new_[4912]_ ,
    \new_[4913]_ , \new_[4914]_ , \new_[4915]_ , \new_[4916]_ ,
    \new_[4917]_ , \new_[4918]_ , \new_[4919]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4923]_ , \new_[4924]_ ,
    \new_[4925]_ , \new_[4926]_ , \new_[4927]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4933]_ , \new_[4934]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4940]_ ,
    \new_[4941]_ , \new_[4942]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4947]_ , \new_[4948]_ ,
    \new_[4949]_ , \new_[4950]_ , \new_[4951]_ , \new_[4952]_ ,
    \new_[4953]_ , \new_[4954]_ , \new_[4955]_ , \new_[4956]_ ,
    \new_[4957]_ , \new_[4958]_ , \new_[4959]_ , \new_[4960]_ ,
    \new_[4961]_ , \new_[4962]_ , \new_[4963]_ , \new_[4964]_ ,
    \new_[4965]_ , \new_[4966]_ , \new_[4967]_ , \new_[4968]_ ,
    \new_[4969]_ , \new_[4970]_ , \new_[4971]_ , \new_[4972]_ ,
    \new_[4973]_ , \new_[4974]_ , \new_[4975]_ , \new_[4976]_ ,
    \new_[4977]_ , \new_[4978]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4981]_ , \new_[4982]_ , \new_[4983]_ , \new_[4984]_ ,
    \new_[4985]_ , \new_[4986]_ , \new_[4987]_ , \new_[4988]_ ,
    \new_[4989]_ , \new_[4990]_ , \new_[4991]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4994]_ , \new_[4995]_ , \new_[4996]_ ,
    \new_[4997]_ , \new_[4998]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5003]_ , \new_[5004]_ ,
    \new_[5005]_ , \new_[5006]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5010]_ , \new_[5011]_ , \new_[5012]_ ,
    \new_[5013]_ , \new_[5014]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5017]_ , \new_[5018]_ , \new_[5019]_ , \new_[5020]_ ,
    \new_[5021]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5027]_ , \new_[5028]_ ,
    \new_[5029]_ , \new_[5030]_ , \new_[5031]_ , \new_[5032]_ ,
    \new_[5033]_ , \new_[5034]_ , \new_[5035]_ , \new_[5036]_ ,
    \new_[5037]_ , \new_[5038]_ , \new_[5039]_ , \new_[5040]_ ,
    \new_[5041]_ , \new_[5042]_ , \new_[5043]_ , \new_[5044]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5048]_ ,
    \new_[5049]_ , \new_[5050]_ , \new_[5051]_ , \new_[5052]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5055]_ , \new_[5056]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5067]_ , \new_[5068]_ ,
    \new_[5069]_ , \new_[5070]_ , \new_[5071]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5075]_ , \new_[5076]_ ,
    \new_[5077]_ , \new_[5078]_ , \new_[5079]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5082]_ , \new_[5083]_ , \new_[5084]_ ,
    \new_[5085]_ , \new_[5086]_ , \new_[5087]_ , \new_[5088]_ ,
    \new_[5089]_ , \new_[5090]_ , \new_[5091]_ , \new_[5092]_ ,
    \new_[5093]_ , \new_[5094]_ , \new_[5095]_ , \new_[5096]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5099]_ , \new_[5100]_ ,
    \new_[5101]_ , \new_[5102]_ , \new_[5103]_ , \new_[5104]_ ,
    \new_[5105]_ , \new_[5106]_ , \new_[5107]_ , \new_[5108]_ ,
    \new_[5109]_ , \new_[5110]_ , \new_[5111]_ , \new_[5112]_ ,
    \new_[5113]_ , \new_[5114]_ , \new_[5115]_ , \new_[5116]_ ,
    \new_[5117]_ , \new_[5118]_ , \new_[5119]_ , \new_[5120]_ ,
    \new_[5121]_ , \new_[5122]_ , \new_[5123]_ , \new_[5124]_ ,
    \new_[5125]_ , \new_[5126]_ , \new_[5127]_ , \new_[5128]_ ,
    \new_[5129]_ , \new_[5130]_ , \new_[5131]_ , \new_[5132]_ ,
    \new_[5133]_ , \new_[5134]_ , \new_[5135]_ , \new_[5136]_ ,
    \new_[5137]_ , \new_[5138]_ , \new_[5139]_ , \new_[5140]_ ,
    \new_[5141]_ , \new_[5142]_ , \new_[5143]_ , \new_[5144]_ ,
    \new_[5145]_ , \new_[5146]_ , \new_[5147]_ , \new_[5148]_ ,
    \new_[5149]_ , \new_[5150]_ , \new_[5151]_ , \new_[5152]_ ,
    \new_[5153]_ , \new_[5154]_ , \new_[5155]_ , \new_[5156]_ ,
    \new_[5157]_ , \new_[5158]_ , \new_[5159]_ , \new_[5160]_ ,
    \new_[5161]_ , \new_[5162]_ , \new_[5163]_ , \new_[5164]_ ,
    \new_[5165]_ , \new_[5166]_ , \new_[5167]_ , \new_[5168]_ ,
    \new_[5169]_ , \new_[5170]_ , \new_[5171]_ , \new_[5172]_ ,
    \new_[5173]_ , \new_[5174]_ , \new_[5175]_ , \new_[5176]_ ,
    \new_[5177]_ , \new_[5178]_ , \new_[5179]_ , \new_[5180]_ ,
    \new_[5181]_ , \new_[5182]_ , \new_[5183]_ , \new_[5184]_ ,
    \new_[5185]_ , \new_[5186]_ , \new_[5187]_ , \new_[5188]_ ,
    \new_[5189]_ , \new_[5190]_ , \new_[5191]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5194]_ , \new_[5195]_ , \new_[5196]_ ,
    \new_[5197]_ , \new_[5198]_ , \new_[5199]_ , \new_[5200]_ ,
    \new_[5201]_ , \new_[5202]_ , \new_[5203]_ , \new_[5204]_ ,
    \new_[5205]_ , \new_[5206]_ , \new_[5207]_ , \new_[5208]_ ,
    \new_[5209]_ , \new_[5210]_ , \new_[5211]_ , \new_[5212]_ ,
    \new_[5213]_ , \new_[5214]_ , \new_[5215]_ , \new_[5216]_ ,
    \new_[5217]_ , \new_[5218]_ , \new_[5219]_ , \new_[5220]_ ,
    \new_[5221]_ , \new_[5222]_ , \new_[5223]_ , \new_[5224]_ ,
    \new_[5225]_ , \new_[5226]_ , \new_[5227]_ , \new_[5228]_ ,
    \new_[5229]_ , \new_[5230]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5233]_ , \new_[5234]_ , \new_[5235]_ , \new_[5236]_ ,
    \new_[5237]_ , \new_[5238]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5242]_ , \new_[5243]_ , \new_[5244]_ ,
    \new_[5245]_ , \new_[5246]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5249]_ , \new_[5250]_ , \new_[5251]_ , \new_[5252]_ ,
    \new_[5253]_ , \new_[5254]_ , \new_[5255]_ , \new_[5256]_ ,
    \new_[5257]_ , \new_[5258]_ , \new_[5259]_ , \new_[5260]_ ,
    \new_[5261]_ , \new_[5262]_ , \new_[5263]_ , \new_[5264]_ ,
    \new_[5265]_ , \new_[5266]_ , \new_[5267]_ , \new_[5268]_ ,
    \new_[5269]_ , \new_[5270]_ , \new_[5271]_ , \new_[5272]_ ,
    \new_[5273]_ , \new_[5274]_ , \new_[5275]_ , \new_[5276]_ ,
    \new_[5277]_ , \new_[5278]_ , \new_[5279]_ , \new_[5280]_ ,
    \new_[5281]_ , \new_[5282]_ , \new_[5283]_ , \new_[5284]_ ,
    \new_[5285]_ , \new_[5286]_ , \new_[5287]_ , \new_[5288]_ ,
    \new_[5289]_ , \new_[5290]_ , \new_[5291]_ , \new_[5292]_ ,
    \new_[5293]_ , \new_[5294]_ , \new_[5295]_ , \new_[5296]_ ,
    \new_[5297]_ , \new_[5298]_ , \new_[5299]_ , \new_[5300]_ ,
    \new_[5301]_ , \new_[5302]_ , \new_[5303]_ , \new_[5304]_ ,
    \new_[5305]_ , \new_[5306]_ , \new_[5307]_ , \new_[5308]_ ,
    \new_[5309]_ , \new_[5310]_ , \new_[5311]_ , \new_[5312]_ ,
    \new_[5313]_ , \new_[5314]_ , \new_[5315]_ , \new_[5316]_ ,
    \new_[5317]_ , \new_[5318]_ , \new_[5319]_ , \new_[5320]_ ,
    \new_[5321]_ , \new_[5322]_ , \new_[5323]_ , \new_[5324]_ ,
    \new_[5325]_ , \new_[5326]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5329]_ , \new_[5330]_ , \new_[5331]_ , \new_[5332]_ ,
    \new_[5333]_ , \new_[5334]_ , \new_[5335]_ , \new_[5336]_ ,
    \new_[5337]_ , \new_[5338]_ , \new_[5339]_ , \new_[5340]_ ,
    \new_[5341]_ , \new_[5342]_ , \new_[5343]_ , \new_[5344]_ ,
    \new_[5345]_ , \new_[5346]_ , \new_[5347]_ , \new_[5348]_ ,
    \new_[5349]_ , \new_[5350]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5355]_ , \new_[5356]_ ,
    \new_[5357]_ , \new_[5358]_ , \new_[5359]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5362]_ , \new_[5363]_ , \new_[5364]_ ,
    \new_[5365]_ , \new_[5366]_ , \new_[5367]_ , \new_[5368]_ ,
    \new_[5369]_ , \new_[5370]_ , \new_[5371]_ , \new_[5372]_ ,
    \new_[5373]_ , \new_[5374]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5377]_ , \new_[5378]_ , \new_[5379]_ , \new_[5380]_ ,
    \new_[5381]_ , \new_[5382]_ , \new_[5383]_ , \new_[5384]_ ,
    \new_[5385]_ , \new_[5386]_ , \new_[5387]_ , \new_[5388]_ ,
    \new_[5389]_ , \new_[5390]_ , \new_[5391]_ , \new_[5392]_ ,
    \new_[5393]_ , \new_[5394]_ , \new_[5395]_ , \new_[5396]_ ,
    \new_[5397]_ , \new_[5398]_ , \new_[5399]_ , \new_[5400]_ ,
    \new_[5401]_ , \new_[5402]_ , \new_[5403]_ , \new_[5404]_ ,
    \new_[5405]_ , \new_[5406]_ , \new_[5407]_ , \new_[5408]_ ,
    \new_[5409]_ , \new_[5410]_ , \new_[5411]_ , \new_[5412]_ ,
    \new_[5413]_ , \new_[5414]_ , \new_[5415]_ , \new_[5416]_ ,
    \new_[5417]_ , \new_[5418]_ , \new_[5419]_ , \new_[5420]_ ,
    \new_[5421]_ , \new_[5422]_ , \new_[5423]_ , \new_[5424]_ ,
    \new_[5425]_ , \new_[5426]_ , \new_[5427]_ , \new_[5428]_ ,
    \new_[5429]_ , \new_[5430]_ , \new_[5433]_ , \new_[5434]_ ,
    \new_[5435]_ , \new_[5436]_ , \new_[5437]_ , \new_[5438]_ ,
    \new_[5439]_ , \new_[5440]_ , \new_[5441]_ , \new_[5442]_ ,
    \new_[5443]_ , \new_[5444]_ , \new_[5445]_ , \new_[5446]_ ,
    \new_[5447]_ , \new_[5448]_ , \new_[5449]_ , \new_[5450]_ ,
    \new_[5451]_ , \new_[5452]_ , \new_[5453]_ , \new_[5454]_ ,
    \new_[5455]_ , \new_[5456]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5459]_ , \new_[5460]_ , \new_[5461]_ , \new_[5462]_ ,
    \new_[5463]_ , \new_[5464]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5468]_ , \new_[5469]_ , \new_[5470]_ ,
    \new_[5471]_ , \new_[5472]_ , \new_[5473]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5476]_ , \new_[5477]_ , \new_[5478]_ ,
    \new_[5479]_ , \new_[5481]_ , \new_[5482]_ , \new_[5483]_ ,
    \new_[5484]_ , \new_[5485]_ , \new_[5486]_ , \new_[5487]_ ,
    \new_[5488]_ , \new_[5489]_ , \new_[5490]_ , \new_[5491]_ ,
    \new_[5492]_ , \new_[5493]_ , \new_[5494]_ , \new_[5495]_ ,
    \new_[5496]_ , \new_[5497]_ , \new_[5498]_ , \new_[5499]_ ,
    \new_[5500]_ , \new_[5501]_ , \new_[5502]_ , \new_[5503]_ ,
    \new_[5504]_ , \new_[5505]_ , \new_[5506]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5513]_ , \new_[5514]_ , \new_[5515]_ ,
    \new_[5516]_ , \new_[5517]_ , \new_[5518]_ , \new_[5519]_ ,
    \new_[5520]_ , \new_[5521]_ , \new_[5522]_ , \new_[5523]_ ,
    \new_[5524]_ , \new_[5525]_ , \new_[5526]_ , \new_[5527]_ ,
    \new_[5528]_ , \new_[5529]_ , \new_[5530]_ , \new_[5531]_ ,
    \new_[5532]_ , \new_[5533]_ , \new_[5534]_ , \new_[5535]_ ,
    \new_[5536]_ , \new_[5537]_ , \new_[5538]_ , \new_[5539]_ ,
    \new_[5540]_ , \new_[5541]_ , \new_[5542]_ , \new_[5543]_ ,
    \new_[5544]_ , \new_[5545]_ , \new_[5546]_ , \new_[5547]_ ,
    \new_[5549]_ , \new_[5550]_ , \new_[5551]_ , \new_[5552]_ ,
    \new_[5553]_ , \new_[5554]_ , \new_[5555]_ , \new_[5556]_ ,
    \new_[5557]_ , \new_[5558]_ , \new_[5559]_ , \new_[5560]_ ,
    \new_[5561]_ , \new_[5562]_ , \new_[5563]_ , \new_[5564]_ ,
    \new_[5565]_ , \new_[5566]_ , \new_[5567]_ , \new_[5568]_ ,
    \new_[5569]_ , \new_[5570]_ , \new_[5571]_ , \new_[5572]_ ,
    \new_[5573]_ , \new_[5574]_ , \new_[5575]_ , \new_[5576]_ ,
    \new_[5577]_ , \new_[5578]_ , \new_[5579]_ , \new_[5580]_ ,
    \new_[5581]_ , \new_[5582]_ , \new_[5583]_ , \new_[5584]_ ,
    \new_[5585]_ , \new_[5586]_ , \new_[5587]_ , \new_[5588]_ ,
    \new_[5589]_ , \new_[5590]_ , \new_[5591]_ , \new_[5592]_ ,
    \new_[5593]_ , \new_[5594]_ , \new_[5595]_ , \new_[5596]_ ,
    \new_[5597]_ , \new_[5598]_ , \new_[5599]_ , \new_[5600]_ ,
    \new_[5601]_ , \new_[5602]_ , \new_[5603]_ , \new_[5604]_ ,
    \new_[5605]_ , \new_[5606]_ , \new_[5607]_ , \new_[5608]_ ,
    \new_[5609]_ , \new_[5610]_ , \new_[5611]_ , \new_[5612]_ ,
    \new_[5613]_ , \new_[5614]_ , \new_[5615]_ , \new_[5617]_ ,
    \new_[5618]_ , \new_[5619]_ , \new_[5620]_ , \new_[5621]_ ,
    \new_[5622]_ , \new_[5623]_ , \new_[5624]_ , \new_[5625]_ ,
    \new_[5626]_ , \new_[5627]_ , \new_[5628]_ , \new_[5629]_ ,
    \new_[5630]_ , \new_[5631]_ , \new_[5632]_ , \new_[5633]_ ,
    \new_[5634]_ , \new_[5635]_ , \new_[5636]_ , \new_[5637]_ ,
    \new_[5638]_ , \new_[5639]_ , \new_[5640]_ , \new_[5641]_ ,
    \new_[5642]_ , \new_[5643]_ , \new_[5644]_ , \new_[5645]_ ,
    \new_[5646]_ , \new_[5647]_ , \new_[5648]_ , \new_[5649]_ ,
    \new_[5650]_ , \new_[5651]_ , \new_[5652]_ , \new_[5653]_ ,
    \new_[5654]_ , \new_[5655]_ , \new_[5656]_ , \new_[5657]_ ,
    \new_[5658]_ , \new_[5659]_ , \new_[5660]_ , \new_[5661]_ ,
    \new_[5662]_ , \new_[5663]_ , \new_[5664]_ , \new_[5665]_ ,
    \new_[5666]_ , \new_[5667]_ , \new_[5668]_ , \new_[5669]_ ,
    \new_[5670]_ , \new_[5671]_ , \new_[5672]_ , \new_[5673]_ ,
    \new_[5674]_ , \new_[5675]_ , \new_[5676]_ , \new_[5677]_ ,
    \new_[5678]_ , \new_[5679]_ , \new_[5680]_ , \new_[5681]_ ,
    \new_[5682]_ , \new_[5683]_ , \new_[5684]_ , \new_[5685]_ ,
    \new_[5686]_ , \new_[5687]_ , \new_[5688]_ , \new_[5689]_ ,
    \new_[5690]_ , \new_[5691]_ , \new_[5692]_ , \new_[5693]_ ,
    \new_[5694]_ , \new_[5695]_ , \new_[5696]_ , \new_[5697]_ ,
    \new_[5698]_ , \new_[5699]_ , \new_[5700]_ , \new_[5701]_ ,
    \new_[5702]_ , \new_[5703]_ , \new_[5704]_ , \new_[5705]_ ,
    \new_[5706]_ , \new_[5707]_ , \new_[5708]_ , \new_[5709]_ ,
    \new_[5710]_ , \new_[5711]_ , \new_[5712]_ , \new_[5713]_ ,
    \new_[5714]_ , \new_[5715]_ , \new_[5716]_ , \new_[5717]_ ,
    \new_[5718]_ , \new_[5719]_ , \new_[5720]_ , \new_[5721]_ ,
    \new_[5722]_ , \new_[5723]_ , \new_[5724]_ , \new_[5725]_ ,
    \new_[5726]_ , \new_[5727]_ , \new_[5728]_ , \new_[5729]_ ,
    \new_[5730]_ , \new_[5731]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5734]_ , \new_[5735]_ , \new_[5736]_ , \new_[5737]_ ,
    \new_[5738]_ , \new_[5739]_ , \new_[5740]_ , \new_[5741]_ ,
    \new_[5742]_ , \new_[5743]_ , \new_[5744]_ , \new_[5745]_ ,
    \new_[5746]_ , \new_[5747]_ , \new_[5748]_ , \new_[5749]_ ,
    \new_[5750]_ , \new_[5751]_ , \new_[5752]_ , \new_[5753]_ ,
    \new_[5754]_ , \new_[5755]_ , \new_[5756]_ , \new_[5757]_ ,
    \new_[5759]_ , \new_[5760]_ , \new_[5761]_ , \new_[5762]_ ,
    \new_[5763]_ , \new_[5764]_ , \new_[5765]_ , \new_[5766]_ ,
    \new_[5767]_ , \new_[5768]_ , \new_[5769]_ , \new_[5770]_ ,
    \new_[5771]_ , \new_[5772]_ , \new_[5773]_ , \new_[5774]_ ,
    \new_[5775]_ , \new_[5776]_ , \new_[5777]_ , \new_[5778]_ ,
    \new_[5779]_ , \new_[5780]_ , \new_[5781]_ , \new_[5782]_ ,
    \new_[5783]_ , \new_[5784]_ , \new_[5785]_ , \new_[5787]_ ,
    \new_[5788]_ , \new_[5789]_ , \new_[5790]_ , \new_[5791]_ ,
    \new_[5792]_ , \new_[5793]_ , \new_[5794]_ , \new_[5795]_ ,
    \new_[5796]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5800]_ , \new_[5801]_ , \new_[5802]_ , \new_[5803]_ ,
    \new_[5804]_ , \new_[5805]_ , \new_[5806]_ , \new_[5807]_ ,
    \new_[5808]_ , \new_[5809]_ , \new_[5810]_ , \new_[5811]_ ,
    \new_[5812]_ , \new_[5813]_ , \new_[5814]_ , \new_[5815]_ ,
    \new_[5816]_ , \new_[5817]_ , \new_[5818]_ , \new_[5819]_ ,
    \new_[5820]_ , \new_[5821]_ , \new_[5822]_ , \new_[5823]_ ,
    \new_[5824]_ , \new_[5825]_ , \new_[5826]_ , \new_[5827]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5830]_ , \new_[5831]_ ,
    \new_[5832]_ , \new_[5833]_ , \new_[5834]_ , \new_[5835]_ ,
    \new_[5836]_ , \new_[5837]_ , \new_[5838]_ , \new_[5839]_ ,
    \new_[5840]_ , \new_[5841]_ , \new_[5842]_ , \new_[5843]_ ,
    \new_[5844]_ , \new_[5845]_ , \new_[5846]_ , \new_[5847]_ ,
    \new_[5848]_ , \new_[5849]_ , \new_[5850]_ , \new_[5851]_ ,
    \new_[5852]_ , \new_[5853]_ , \new_[5854]_ , \new_[5855]_ ,
    \new_[5856]_ , \new_[5857]_ , \new_[5858]_ , \new_[5859]_ ,
    \new_[5860]_ , \new_[5861]_ , \new_[5862]_ , \new_[5863]_ ,
    \new_[5864]_ , \new_[5865]_ , \new_[5866]_ , \new_[5867]_ ,
    \new_[5868]_ , \new_[5869]_ , \new_[5870]_ , \new_[5871]_ ,
    \new_[5872]_ , \new_[5873]_ , \new_[5874]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5877]_ , \new_[5878]_ , \new_[5879]_ ,
    \new_[5880]_ , \new_[5881]_ , \new_[5882]_ , \new_[5883]_ ,
    \new_[5884]_ , \new_[5885]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5888]_ , \new_[5889]_ , \new_[5890]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5896]_ , \new_[5897]_ , \new_[5898]_ , \new_[5899]_ ,
    \new_[5900]_ , \new_[5901]_ , \new_[5902]_ , \new_[5903]_ ,
    \new_[5904]_ , \new_[5905]_ , \new_[5906]_ , \new_[5907]_ ,
    \new_[5908]_ , \new_[5910]_ , \new_[5911]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5914]_ , \new_[5915]_ , \new_[5916]_ ,
    \new_[5917]_ , \new_[5918]_ , \new_[5919]_ , \new_[5920]_ ,
    \new_[5921]_ , \new_[5922]_ , \new_[5923]_ , \new_[5924]_ ,
    \new_[5926]_ , \new_[5927]_ , \new_[5928]_ , \new_[5929]_ ,
    \new_[5930]_ , \new_[5931]_ , \new_[5932]_ , \new_[5933]_ ,
    \new_[5934]_ , \new_[5935]_ , \new_[5936]_ , \new_[5937]_ ,
    \new_[5938]_ , \new_[5939]_ , \new_[5940]_ , \new_[5941]_ ,
    \new_[5942]_ , \new_[5943]_ , \new_[5944]_ , \new_[5945]_ ,
    \new_[5946]_ , \new_[5947]_ , \new_[5948]_ , \new_[5949]_ ,
    \new_[5950]_ , \new_[5951]_ , \new_[5952]_ , \new_[5953]_ ,
    \new_[5954]_ , \new_[5955]_ , \new_[5956]_ , \new_[5957]_ ,
    \new_[5958]_ , \new_[5959]_ , \new_[5960]_ , \new_[5961]_ ,
    \new_[5962]_ , \new_[5963]_ , \new_[5964]_ , \new_[5965]_ ,
    \new_[5966]_ , \new_[5967]_ , \new_[5968]_ , \new_[5969]_ ,
    \new_[5970]_ , \new_[5971]_ , \new_[5972]_ , \new_[5973]_ ,
    \new_[5974]_ , \new_[5975]_ , \new_[5976]_ , \new_[5977]_ ,
    \new_[5978]_ , \new_[5979]_ , \new_[5980]_ , \new_[5981]_ ,
    \new_[5982]_ , \new_[5983]_ , \new_[5984]_ , \new_[5985]_ ,
    \new_[5986]_ , \new_[5987]_ , \new_[5988]_ , \new_[5989]_ ,
    \new_[5990]_ , \new_[5991]_ , \new_[5992]_ , \new_[5994]_ ,
    \new_[5995]_ , \new_[5996]_ , \new_[5997]_ , \new_[5998]_ ,
    \new_[5999]_ , \new_[6001]_ , \new_[6002]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6005]_ , \new_[6006]_ , \new_[6007]_ ,
    \new_[6008]_ , \new_[6009]_ , \new_[6010]_ , \new_[6011]_ ,
    \new_[6012]_ , \new_[6013]_ , \new_[6014]_ , \new_[6015]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6022]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6028]_ , \new_[6029]_ , \new_[6030]_ , \new_[6031]_ ,
    \new_[6032]_ , \new_[6033]_ , \new_[6034]_ , \new_[6035]_ ,
    \new_[6036]_ , \new_[6037]_ , \new_[6038]_ , \new_[6039]_ ,
    \new_[6040]_ , \new_[6041]_ , \new_[6042]_ , \new_[6043]_ ,
    \new_[6044]_ , \new_[6045]_ , \new_[6046]_ , \new_[6047]_ ,
    \new_[6048]_ , \new_[6049]_ , \new_[6050]_ , \new_[6051]_ ,
    \new_[6052]_ , \new_[6053]_ , \new_[6054]_ , \new_[6055]_ ,
    \new_[6056]_ , \new_[6057]_ , \new_[6058]_ , \new_[6059]_ ,
    \new_[6060]_ , \new_[6061]_ , \new_[6062]_ , \new_[6063]_ ,
    \new_[6064]_ , \new_[6065]_ , \new_[6066]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6069]_ , \new_[6070]_ , \new_[6071]_ ,
    \new_[6072]_ , \new_[6073]_ , \new_[6074]_ , \new_[6076]_ ,
    \new_[6077]_ , \new_[6078]_ , \new_[6079]_ , \new_[6080]_ ,
    \new_[6081]_ , \new_[6082]_ , \new_[6083]_ , \new_[6084]_ ,
    \new_[6085]_ , \new_[6086]_ , \new_[6087]_ , \new_[6088]_ ,
    \new_[6089]_ , \new_[6090]_ , \new_[6091]_ , \new_[6092]_ ,
    \new_[6093]_ , \new_[6094]_ , \new_[6095]_ , \new_[6096]_ ,
    \new_[6097]_ , \new_[6098]_ , \new_[6099]_ , \new_[6100]_ ,
    \new_[6101]_ , \new_[6102]_ , \new_[6103]_ , \new_[6104]_ ,
    \new_[6105]_ , \new_[6106]_ , \new_[6107]_ , \new_[6108]_ ,
    \new_[6109]_ , \new_[6110]_ , \new_[6111]_ , \new_[6112]_ ,
    \new_[6113]_ , \new_[6114]_ , \new_[6115]_ , \new_[6116]_ ,
    \new_[6117]_ , \new_[6118]_ , \new_[6119]_ , \new_[6120]_ ,
    \new_[6121]_ , \new_[6122]_ , \new_[6123]_ , \new_[6124]_ ,
    \new_[6125]_ , \new_[6126]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6130]_ , \new_[6131]_ , \new_[6132]_ ,
    \new_[6133]_ , \new_[6134]_ , \new_[6135]_ , \new_[6136]_ ,
    \new_[6137]_ , \new_[6138]_ , \new_[6139]_ , \new_[6140]_ ,
    \new_[6141]_ , \new_[6142]_ , \new_[6143]_ , \new_[6144]_ ,
    \new_[6145]_ , \new_[6146]_ , \new_[6147]_ , \new_[6148]_ ,
    \new_[6149]_ , \new_[6150]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6155]_ , \new_[6158]_ , \new_[6159]_ ,
    \new_[6160]_ , \new_[6161]_ , \new_[6162]_ , \new_[6163]_ ,
    \new_[6164]_ , \new_[6165]_ , \new_[6166]_ , \new_[6167]_ ,
    \new_[6168]_ , \new_[6169]_ , \new_[6170]_ , \new_[6171]_ ,
    \new_[6172]_ , \new_[6173]_ , \new_[6174]_ , \new_[6175]_ ,
    \new_[6176]_ , \new_[6177]_ , \new_[6178]_ , \new_[6179]_ ,
    \new_[6180]_ , \new_[6181]_ , \new_[6182]_ , \new_[6183]_ ,
    \new_[6184]_ , \new_[6185]_ , \new_[6186]_ , \new_[6187]_ ,
    \new_[6188]_ , \new_[6189]_ , \new_[6190]_ , \new_[6191]_ ,
    \new_[6192]_ , \new_[6193]_ , \new_[6194]_ , \new_[6195]_ ,
    \new_[6196]_ , \new_[6197]_ , \new_[6198]_ , \new_[6199]_ ,
    \new_[6200]_ , \new_[6201]_ , \new_[6202]_ , \new_[6203]_ ,
    \new_[6204]_ , \new_[6205]_ , \new_[6206]_ , \new_[6207]_ ,
    \new_[6208]_ , \new_[6209]_ , \new_[6210]_ , \new_[6211]_ ,
    \new_[6212]_ , \new_[6213]_ , \new_[6214]_ , \new_[6215]_ ,
    \new_[6216]_ , \new_[6217]_ , \new_[6218]_ , \new_[6219]_ ,
    \new_[6220]_ , \new_[6221]_ , \new_[6222]_ , \new_[6223]_ ,
    \new_[6224]_ , \new_[6225]_ , \new_[6226]_ , \new_[6227]_ ,
    \new_[6228]_ , \new_[6229]_ , \new_[6230]_ , \new_[6231]_ ,
    \new_[6232]_ , \new_[6233]_ , \new_[6234]_ , \new_[6235]_ ,
    \new_[6236]_ , \new_[6237]_ , \new_[6238]_ , \new_[6239]_ ,
    \new_[6240]_ , \new_[6241]_ , \new_[6242]_ , \new_[6243]_ ,
    \new_[6244]_ , \new_[6245]_ , \new_[6246]_ , \new_[6247]_ ,
    \new_[6248]_ , \new_[6249]_ , \new_[6250]_ , \new_[6251]_ ,
    \new_[6252]_ , \new_[6253]_ , \new_[6254]_ , \new_[6255]_ ,
    \new_[6256]_ , \new_[6257]_ , \new_[6258]_ , \new_[6259]_ ,
    \new_[6260]_ , \new_[6261]_ , \new_[6262]_ , \new_[6263]_ ,
    \new_[6264]_ , \new_[6265]_ , \new_[6266]_ , \new_[6267]_ ,
    \new_[6268]_ , \new_[6269]_ , \new_[6270]_ , \new_[6271]_ ,
    \new_[6272]_ , \new_[6273]_ , \new_[6274]_ , \new_[6275]_ ,
    \new_[6276]_ , \new_[6277]_ , \new_[6278]_ , \new_[6279]_ ,
    \new_[6280]_ , \new_[6281]_ , \new_[6282]_ , \new_[6283]_ ,
    \new_[6284]_ , \new_[6285]_ , \new_[6286]_ , \new_[6287]_ ,
    \new_[6288]_ , \new_[6289]_ , \new_[6290]_ , \new_[6291]_ ,
    \new_[6292]_ , \new_[6293]_ , \new_[6294]_ , \new_[6295]_ ,
    \new_[6296]_ , \new_[6297]_ , \new_[6298]_ , \new_[6299]_ ,
    \new_[6300]_ , \new_[6301]_ , \new_[6302]_ , \new_[6303]_ ,
    \new_[6304]_ , \new_[6305]_ , \new_[6306]_ , \new_[6307]_ ,
    \new_[6308]_ , \new_[6309]_ , \new_[6310]_ , \new_[6311]_ ,
    \new_[6312]_ , \new_[6313]_ , \new_[6314]_ , \new_[6315]_ ,
    \new_[6316]_ , \new_[6317]_ , \new_[6318]_ , \new_[6319]_ ,
    \new_[6320]_ , \new_[6321]_ , \new_[6322]_ , \new_[6323]_ ,
    \new_[6324]_ , \new_[6325]_ , \new_[6326]_ , \new_[6327]_ ,
    \new_[6328]_ , \new_[6329]_ , \new_[6330]_ , \new_[6331]_ ,
    \new_[6332]_ , \new_[6333]_ , \new_[6334]_ , \new_[6335]_ ,
    \new_[6336]_ , \new_[6337]_ , \new_[6338]_ , \new_[6339]_ ,
    \new_[6340]_ , \new_[6341]_ , \new_[6342]_ , \new_[6343]_ ,
    \new_[6344]_ , \new_[6345]_ , \new_[6346]_ , \new_[6347]_ ,
    \new_[6348]_ , \new_[6349]_ , \new_[6350]_ , \new_[6351]_ ,
    \new_[6352]_ , \new_[6353]_ , \new_[6354]_ , \new_[6355]_ ,
    \new_[6356]_ , \new_[6357]_ , \new_[6358]_ , \new_[6359]_ ,
    \new_[6360]_ , \new_[6361]_ , \new_[6362]_ , \new_[6363]_ ,
    \new_[6364]_ , \new_[6365]_ , \new_[6366]_ , \new_[6367]_ ,
    \new_[6368]_ , \new_[6369]_ , \new_[6370]_ , \new_[6371]_ ,
    \new_[6372]_ , \new_[6373]_ , \new_[6374]_ , \new_[6375]_ ,
    \new_[6376]_ , \new_[6377]_ , \new_[6378]_ , \new_[6379]_ ,
    \new_[6380]_ , \new_[6381]_ , \new_[6382]_ , \new_[6383]_ ,
    \new_[6384]_ , \new_[6385]_ , \new_[6386]_ , \new_[6387]_ ,
    \new_[6388]_ , \new_[6389]_ , \new_[6390]_ , \new_[6391]_ ,
    \new_[6392]_ , \new_[6393]_ , \new_[6394]_ , \new_[6395]_ ,
    \new_[6396]_ , \new_[6397]_ , \new_[6398]_ , \new_[6399]_ ,
    \new_[6400]_ , \new_[6401]_ , \new_[6402]_ , \new_[6403]_ ,
    \new_[6404]_ , \new_[6405]_ , \new_[6406]_ , \new_[6407]_ ,
    \new_[6408]_ , \new_[6409]_ , \new_[6410]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6413]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6416]_ , \new_[6417]_ , \new_[6418]_ , \new_[6419]_ ,
    \new_[6420]_ , \new_[6421]_ , \new_[6422]_ , \new_[6423]_ ,
    \new_[6424]_ , \new_[6425]_ , \new_[6426]_ , \new_[6427]_ ,
    \new_[6428]_ , \new_[6429]_ , \new_[6430]_ , \new_[6431]_ ,
    \new_[6432]_ , \new_[6433]_ , \new_[6434]_ , \new_[6435]_ ,
    \new_[6436]_ , \new_[6437]_ , \new_[6438]_ , \new_[6439]_ ,
    \new_[6440]_ , \new_[6441]_ , \new_[6442]_ , \new_[6443]_ ,
    \new_[6444]_ , \new_[6445]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6449]_ , \new_[6450]_ , \new_[6451]_ ,
    \new_[6452]_ , \new_[6453]_ , \new_[6454]_ , \new_[6455]_ ,
    \new_[6456]_ , \new_[6457]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6460]_ , \new_[6461]_ , \new_[6462]_ , \new_[6463]_ ,
    \new_[6464]_ , \new_[6465]_ , \new_[6466]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6470]_ , \new_[6471]_ ,
    \new_[6472]_ , \new_[6473]_ , \new_[6474]_ , \new_[6475]_ ,
    \new_[6476]_ , \new_[6477]_ , \new_[6478]_ , \new_[6479]_ ,
    \new_[6480]_ , \new_[6481]_ , \new_[6482]_ , \new_[6483]_ ,
    \new_[6484]_ , \new_[6485]_ , \new_[6486]_ , \new_[6487]_ ,
    \new_[6488]_ , \new_[6489]_ , \new_[6490]_ , \new_[6491]_ ,
    \new_[6492]_ , \new_[6493]_ , \new_[6494]_ , \new_[6495]_ ,
    \new_[6496]_ , \new_[6497]_ , \new_[6498]_ , \new_[6499]_ ,
    \new_[6500]_ , \new_[6501]_ , \new_[6502]_ , \new_[6503]_ ,
    \new_[6504]_ , \new_[6505]_ , \new_[6506]_ , \new_[6507]_ ,
    \new_[6508]_ , \new_[6509]_ , \new_[6510]_ , \new_[6511]_ ,
    \new_[6512]_ , \new_[6513]_ , \new_[6514]_ , \new_[6515]_ ,
    \new_[6516]_ , \new_[6517]_ , \new_[6518]_ , \new_[6519]_ ,
    \new_[6520]_ , \new_[6521]_ , \new_[6522]_ , \new_[6523]_ ,
    \new_[6524]_ , \new_[6525]_ , \new_[6526]_ , \new_[6527]_ ,
    \new_[6528]_ , \new_[6529]_ , \new_[6530]_ , \new_[6531]_ ,
    \new_[6532]_ , \new_[6533]_ , \new_[6534]_ , \new_[6535]_ ,
    \new_[6536]_ , \new_[6537]_ , \new_[6538]_ , \new_[6539]_ ,
    \new_[6540]_ , \new_[6541]_ , \new_[6542]_ , \new_[6543]_ ,
    \new_[6544]_ , \new_[6545]_ , \new_[6546]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6549]_ , \new_[6550]_ , \new_[6551]_ ,
    \new_[6552]_ , \new_[6553]_ , \new_[6554]_ , \new_[6555]_ ,
    \new_[6556]_ , \new_[6557]_ , \new_[6558]_ , \new_[6559]_ ,
    \new_[6560]_ , \new_[6561]_ , \new_[6562]_ , \new_[6563]_ ,
    \new_[6564]_ , \new_[6565]_ , \new_[6566]_ , \new_[6567]_ ,
    \new_[6568]_ , \new_[6569]_ , \new_[6570]_ , \new_[6571]_ ,
    \new_[6572]_ , \new_[6573]_ , \new_[6574]_ , \new_[6575]_ ,
    \new_[6576]_ , \new_[6577]_ , \new_[6578]_ , \new_[6579]_ ,
    \new_[6580]_ , \new_[6581]_ , \new_[6582]_ , \new_[6583]_ ,
    \new_[6584]_ , \new_[6585]_ , \new_[6586]_ , \new_[6587]_ ,
    \new_[6588]_ , \new_[6589]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6592]_ , \new_[6593]_ , \new_[6594]_ , \new_[6595]_ ,
    \new_[6596]_ , \new_[6597]_ , \new_[6598]_ , \new_[6599]_ ,
    \new_[6600]_ , \new_[6601]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6608]_ , \new_[6609]_ , \new_[6610]_ , \new_[6611]_ ,
    \new_[6612]_ , \new_[6613]_ , \new_[6614]_ , \new_[6615]_ ,
    \new_[6616]_ , \new_[6617]_ , \new_[6618]_ , \new_[6619]_ ,
    \new_[6620]_ , \new_[6621]_ , \new_[6622]_ , \new_[6623]_ ,
    \new_[6624]_ , \new_[6625]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6628]_ , \new_[6629]_ , \new_[6630]_ , \new_[6631]_ ,
    \new_[6632]_ , \new_[6633]_ , \new_[6634]_ , \new_[6635]_ ,
    \new_[6636]_ , \new_[6637]_ , \new_[6638]_ , \new_[6639]_ ,
    \new_[6640]_ , \new_[6641]_ , \new_[6642]_ , \new_[6643]_ ,
    \new_[6644]_ , \new_[6645]_ , \new_[6646]_ , \new_[6647]_ ,
    \new_[6648]_ , \new_[6649]_ , \new_[6650]_ , \new_[6651]_ ,
    \new_[6652]_ , \new_[6653]_ , \new_[6654]_ , \new_[6655]_ ,
    \new_[6656]_ , \new_[6657]_ , \new_[6658]_ , \new_[6659]_ ,
    \new_[6660]_ , \new_[6661]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6664]_ , \new_[6665]_ , \new_[6666]_ , \new_[6667]_ ,
    \new_[6668]_ , \new_[6669]_ , \new_[6670]_ , \new_[6671]_ ,
    \new_[6672]_ , \new_[6673]_ , \new_[6674]_ , \new_[6675]_ ,
    \new_[6676]_ , \new_[6677]_ , \new_[6678]_ , \new_[6679]_ ,
    \new_[6680]_ , \new_[6681]_ , \new_[6682]_ , \new_[6683]_ ,
    \new_[6684]_ , \new_[6685]_ , \new_[6686]_ , \new_[6687]_ ,
    \new_[6688]_ , \new_[6689]_ , \new_[6690]_ , \new_[6691]_ ,
    \new_[6692]_ , \new_[6693]_ , \new_[6694]_ , \new_[6695]_ ,
    \new_[6696]_ , \new_[6697]_ , \new_[6698]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6701]_ , \new_[6702]_ , \new_[6703]_ ,
    \new_[6704]_ , \new_[6705]_ , \new_[6706]_ , \new_[6707]_ ,
    \new_[6708]_ , \new_[6709]_ , \new_[6710]_ , \new_[6711]_ ,
    \new_[6712]_ , \new_[6713]_ , \new_[6714]_ , \new_[6715]_ ,
    \new_[6716]_ , \new_[6717]_ , \new_[6718]_ , \new_[6719]_ ,
    \new_[6720]_ , \new_[6721]_ , \new_[6722]_ , \new_[6723]_ ,
    \new_[6724]_ , \new_[6725]_ , \new_[6726]_ , \new_[6727]_ ,
    \new_[6728]_ , \new_[6729]_ , \new_[6730]_ , \new_[6731]_ ,
    \new_[6732]_ , \new_[6733]_ , \new_[6734]_ , \new_[6735]_ ,
    \new_[6736]_ , \new_[6737]_ , \new_[6738]_ , \new_[6739]_ ,
    \new_[6740]_ , \new_[6741]_ , \new_[6742]_ , \new_[6743]_ ,
    \new_[6744]_ , \new_[6745]_ , \new_[6746]_ , \new_[6747]_ ,
    \new_[6748]_ , \new_[6749]_ , \new_[6750]_ , \new_[6751]_ ,
    \new_[6752]_ , \new_[6753]_ , \new_[6754]_ , \new_[6755]_ ,
    \new_[6756]_ , \new_[6757]_ , \new_[6758]_ , \new_[6760]_ ,
    \new_[6761]_ , \new_[6762]_ , \new_[6763]_ , \new_[6764]_ ,
    \new_[6766]_ , \new_[6767]_ , \new_[6768]_ , \new_[6769]_ ,
    \new_[6770]_ , \new_[6771]_ , \new_[6772]_ , \new_[6773]_ ,
    \new_[6774]_ , \new_[6775]_ , \new_[6776]_ , \new_[6777]_ ,
    \new_[6778]_ , \new_[6779]_ , \new_[6780]_ , \new_[6784]_ ,
    \new_[6785]_ , \new_[6786]_ , \new_[6787]_ , \new_[6788]_ ,
    \new_[6789]_ , \new_[6790]_ , \new_[6791]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6795]_ , \new_[6796]_ ,
    \new_[6797]_ , \new_[6798]_ , \new_[6799]_ , \new_[6800]_ ,
    \new_[6801]_ , \new_[6802]_ , \new_[6803]_ , \new_[6804]_ ,
    \new_[6805]_ , \new_[6806]_ , \new_[6807]_ , \new_[6808]_ ,
    \new_[6809]_ , \new_[6810]_ , \new_[6811]_ , \new_[6812]_ ,
    \new_[6813]_ , \new_[6814]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6817]_ , \new_[6818]_ , \new_[6819]_ , \new_[6820]_ ,
    \new_[6821]_ , \new_[6822]_ , \new_[6823]_ , \new_[6824]_ ,
    \new_[6825]_ , \new_[6826]_ , \new_[6827]_ , \new_[6828]_ ,
    \new_[6829]_ , \new_[6830]_ , \new_[6831]_ , \new_[6832]_ ,
    \new_[6860]_ , \new_[6861]_ , \new_[6862]_ , \new_[6863]_ ,
    \new_[6864]_ , \new_[6865]_ , \new_[6866]_ , \new_[6867]_ ,
    \new_[6868]_ , \new_[6869]_ , \new_[6870]_ , \new_[6871]_ ,
    \new_[6872]_ , \new_[6873]_ , \new_[6874]_ , \new_[6875]_ ,
    \new_[6876]_ , \new_[6877]_ , \new_[6878]_ , \new_[6879]_ ,
    \new_[6880]_ , \new_[6881]_ , \new_[6882]_ , \new_[6883]_ ,
    \new_[6884]_ , \new_[6885]_ , \new_[6886]_ , \new_[6887]_ ,
    \new_[6888]_ , \new_[6889]_ , \new_[6890]_ , \new_[6891]_ ,
    \new_[6892]_ , \new_[6893]_ , \new_[6894]_ , \new_[6895]_ ,
    \new_[6896]_ , \new_[6897]_ , \new_[6898]_ , \new_[6899]_ ,
    \new_[6900]_ , \new_[6901]_ , \new_[6902]_ , \new_[6903]_ ,
    \new_[6904]_ , \new_[6905]_ , \new_[6906]_ , \new_[6907]_ ,
    \new_[6908]_ , \new_[6909]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6913]_ , \new_[6914]_ , \new_[6915]_ , \new_[6918]_ ,
    \new_[6919]_ , \new_[6920]_ , \new_[6921]_ , \new_[6923]_ ,
    \new_[6924]_ , \new_[6925]_ , \new_[6926]_ , \new_[6928]_ ,
    \new_[6929]_ , \new_[6931]_ , \new_[6932]_ , \new_[6933]_ ,
    \new_[6934]_ , \new_[6935]_ , \new_[6936]_ , \new_[6937]_ ,
    \new_[6938]_ , \new_[6939]_ , \new_[6943]_ , \new_[6947]_ ,
    \new_[6949]_ , \new_[6950]_ , \new_[6951]_ , \new_[6952]_ ,
    \new_[6953]_ , \new_[6954]_ , \new_[6955]_ , \new_[6956]_ ,
    \new_[6957]_ , \new_[6958]_ , \new_[7006]_ , \new_[7007]_ ,
    \new_[7008]_ , \new_[7009]_ , \new_[7010]_ , \new_[7011]_ ,
    \new_[7012]_ , \new_[7013]_ , \new_[7014]_ , \new_[7015]_ ,
    \new_[7016]_ , \new_[7017]_ , \new_[7018]_ , \new_[7019]_ ,
    \new_[7020]_ , \new_[7021]_ , \new_[7022]_ , \new_[7023]_ ,
    \new_[7024]_ , \new_[7025]_ , \new_[7026]_ , \new_[7027]_ ,
    \new_[7028]_ , \new_[7029]_ , \new_[7030]_ , \new_[7031]_ ,
    \new_[7032]_ , \new_[7033]_ , \new_[7035]_ , \new_[7036]_ ,
    \new_[7037]_ , \new_[7038]_ , \new_[7039]_ , \new_[7040]_ ,
    \new_[7041]_ , \new_[7042]_ , \new_[7044]_ , \new_[7045]_ ,
    \new_[7046]_ , \new_[7047]_ , \new_[7048]_ , \new_[7049]_ ,
    \new_[7050]_ , \new_[7051]_ , \new_[7052]_ , \new_[7053]_ ,
    \new_[7054]_ , \new_[7055]_ , \new_[7056]_ , \new_[7058]_ ,
    \new_[7059]_ , \new_[7060]_ , \new_[7061]_ , \new_[7062]_ ,
    \new_[7063]_ , \new_[7064]_ , \new_[7065]_ , \new_[7067]_ ,
    \new_[7068]_ , \new_[7069]_ , \new_[7070]_ , \new_[7071]_ ,
    \new_[7072]_ , \new_[7073]_ , \new_[7074]_ , \new_[7075]_ ,
    \new_[7076]_ , \new_[7077]_ , \new_[7078]_ , \new_[7079]_ ,
    \new_[7080]_ , \new_[7081]_ , \new_[7082]_ , \new_[7083]_ ,
    \new_[7084]_ , \new_[7085]_ , \new_[7086]_ , \new_[7087]_ ,
    \new_[7088]_ , \new_[7089]_ , \new_[7090]_ , \new_[7091]_ ,
    \new_[7092]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7096]_ , \new_[7097]_ , \new_[7098]_ , \new_[7099]_ ,
    \new_[7100]_ , \new_[7101]_ , \new_[7102]_ , \new_[7103]_ ,
    \new_[7104]_ , \new_[7105]_ , \new_[7106]_ , \new_[7107]_ ,
    \new_[7108]_ , \new_[7109]_ , \new_[7110]_ , \new_[7111]_ ,
    \new_[7112]_ , \new_[7113]_ , \new_[7114]_ , \new_[7115]_ ,
    \new_[7116]_ , \new_[7117]_ , \new_[7118]_ , \new_[7119]_ ,
    \new_[7120]_ , \new_[7121]_ , \new_[7122]_ , \new_[7123]_ ,
    \new_[7124]_ , \new_[7125]_ , \new_[7126]_ , \new_[7127]_ ,
    \new_[7128]_ , \new_[7129]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7135]_ ,
    \new_[7136]_ , \new_[7137]_ , \new_[7138]_ , \new_[7139]_ ,
    \new_[7140]_ , \new_[7141]_ , \new_[7142]_ , \new_[7143]_ ,
    \new_[7144]_ , \new_[7145]_ , \new_[7146]_ , \new_[7147]_ ,
    \new_[7148]_ , \new_[7149]_ , \new_[7150]_ , \new_[7151]_ ,
    \new_[7152]_ , \new_[7153]_ , \new_[7154]_ , \new_[7155]_ ,
    \new_[7156]_ , \new_[7157]_ , \new_[7158]_ , \new_[7159]_ ,
    \new_[7160]_ , \new_[7161]_ , \new_[7162]_ , \new_[7163]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7169]_ , \new_[7170]_ , \new_[7171]_ ,
    \new_[7172]_ , \new_[7173]_ , \new_[7174]_ , \new_[7175]_ ,
    \new_[7176]_ , \new_[7177]_ , \new_[7178]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7182]_ , \new_[7183]_ ,
    \new_[7184]_ , \new_[7185]_ , \new_[7186]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7192]_ , \new_[7193]_ , \new_[7194]_ , \new_[7195]_ ,
    \new_[7196]_ , \new_[7197]_ , \new_[7198]_ , \new_[7199]_ ,
    \new_[7200]_ , \new_[7201]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7205]_ , \new_[7206]_ , \new_[7207]_ ,
    \new_[7208]_ , \new_[7209]_ , \new_[7210]_ , \new_[7211]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7215]_ ,
    \new_[7216]_ , \new_[7217]_ , \new_[7218]_ , \new_[7219]_ ,
    \new_[7220]_ , \new_[7221]_ , \new_[7222]_ , \new_[7223]_ ,
    \new_[7224]_ , \new_[7225]_ , \new_[7226]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7230]_ , \new_[7231]_ ,
    \new_[7232]_ , \new_[7233]_ , \new_[7234]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7244]_ , \new_[7245]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7248]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7255]_ ,
    \new_[7256]_ , \new_[7257]_ , \new_[7258]_ , \new_[7259]_ ,
    \new_[7260]_ , \new_[7261]_ , \new_[7262]_ , \new_[7263]_ ,
    \new_[7264]_ , \new_[7265]_ , \new_[7266]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7270]_ , \new_[7271]_ ,
    \new_[7272]_ , \new_[7273]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7276]_ , \new_[7277]_ , \new_[7278]_ , \new_[7279]_ ,
    \new_[7280]_ , \new_[7281]_ , \new_[7282]_ , \new_[7283]_ ,
    \new_[7284]_ , \new_[7285]_ , \new_[7286]_ , \new_[7287]_ ,
    \new_[7288]_ , \new_[7289]_ , \new_[7290]_ , \new_[7291]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7294]_ , \new_[7295]_ ,
    \new_[7296]_ , \new_[7297]_ , \new_[7298]_ , \new_[7299]_ ,
    \new_[7300]_ , \new_[7301]_ , \new_[7302]_ , \new_[7303]_ ,
    \new_[7304]_ , \new_[7305]_ , \new_[7306]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7312]_ , \new_[7313]_ , \new_[7314]_ , \new_[7315]_ ,
    \new_[7316]_ , \new_[7317]_ , \new_[7318]_ , \new_[7319]_ ,
    \new_[7320]_ , \new_[7321]_ , \new_[7322]_ , \new_[7323]_ ,
    \new_[7324]_ , \new_[7325]_ , \new_[7326]_ , \new_[7327]_ ,
    \new_[7328]_ , \new_[7329]_ , \new_[7330]_ , \new_[7331]_ ,
    \new_[7332]_ , \new_[7333]_ , \new_[7334]_ , \new_[7335]_ ,
    \new_[7336]_ , \new_[7337]_ , \new_[7338]_ , \new_[7339]_ ,
    \new_[7340]_ , \new_[7341]_ , \new_[7342]_ , \new_[7343]_ ,
    \new_[7344]_ , \new_[7345]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7348]_ , \new_[7349]_ , \new_[7350]_ , \new_[7351]_ ,
    \new_[7352]_ , \new_[7353]_ , \new_[7354]_ , \new_[7355]_ ,
    \new_[7356]_ , \new_[7357]_ , \new_[7358]_ , \new_[7359]_ ,
    \new_[7360]_ , \new_[7361]_ , \new_[7362]_ , \new_[7363]_ ,
    \new_[7364]_ , \new_[7365]_ , \new_[7366]_ , \new_[7367]_ ,
    \new_[7368]_ , \new_[7369]_ , \new_[7370]_ , \new_[7371]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7374]_ , \new_[7375]_ ,
    \new_[7376]_ , \new_[7377]_ , \new_[7378]_ , \new_[7379]_ ,
    \new_[7380]_ , \new_[7381]_ , \new_[7382]_ , \new_[7383]_ ,
    \new_[7384]_ , \new_[7385]_ , \new_[7386]_ , \new_[7387]_ ,
    \new_[7388]_ , \new_[7389]_ , \new_[7390]_ , \new_[7391]_ ,
    \new_[7392]_ , \new_[7393]_ , \new_[7394]_ , \new_[7395]_ ,
    \new_[7396]_ , \new_[7397]_ , \new_[7398]_ , \new_[7399]_ ,
    \new_[7400]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7404]_ , \new_[7405]_ , \new_[7406]_ , \new_[7407]_ ,
    \new_[7408]_ , \new_[7409]_ , \new_[7410]_ , \new_[7411]_ ,
    \new_[7412]_ , \new_[7413]_ , \new_[7414]_ , \new_[7415]_ ,
    \new_[7416]_ , \new_[7417]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7422]_ , \new_[7423]_ ,
    \new_[7424]_ , \new_[7425]_ , \new_[7426]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7429]_ , \new_[7430]_ , \new_[7431]_ ,
    \new_[7432]_ , \new_[7433]_ , \new_[7434]_ , \new_[7435]_ ,
    \new_[7436]_ , \new_[7437]_ , \new_[7438]_ , \new_[7439]_ ,
    \new_[7440]_ , \new_[7441]_ , \new_[7442]_ , \new_[7444]_ ,
    \new_[7445]_ , \new_[7446]_ , \new_[7447]_ , \new_[7448]_ ,
    \new_[7449]_ , \new_[7450]_ , \new_[7451]_ , \new_[7452]_ ,
    \new_[7453]_ , \new_[7454]_ , \new_[7455]_ , \new_[7456]_ ,
    \new_[7457]_ , \new_[7458]_ , \new_[7459]_ , \new_[7460]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7465]_ , \new_[7466]_ , \new_[7467]_ , \new_[7468]_ ,
    \new_[7469]_ , \new_[7470]_ , \new_[7471]_ , \new_[7472]_ ,
    \new_[7473]_ , \new_[7474]_ , \new_[7475]_ , \new_[7476]_ ,
    \new_[7477]_ , \new_[7478]_ , \new_[7479]_ , \new_[7480]_ ,
    \new_[7481]_ , \new_[7482]_ , \new_[7483]_ , \new_[7484]_ ,
    \new_[7485]_ , \new_[7486]_ , \new_[7487]_ , \new_[7488]_ ,
    \new_[7489]_ , \new_[7490]_ , \new_[7491]_ , \new_[7492]_ ,
    \new_[7493]_ , \new_[7494]_ , \new_[7495]_ , \new_[7496]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7499]_ , \new_[7500]_ ,
    \new_[7501]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7506]_ , \new_[7507]_ , \new_[7508]_ ,
    \new_[7509]_ , \new_[7510]_ , \new_[7511]_ , \new_[7512]_ ,
    \new_[7513]_ , \new_[7514]_ , \new_[7515]_ , \new_[7516]_ ,
    \new_[7517]_ , \new_[7518]_ , \new_[7519]_ , \new_[7520]_ ,
    \new_[7521]_ , \new_[7522]_ , \new_[7523]_ , \new_[7524]_ ,
    \new_[7525]_ , \new_[7526]_ , \new_[7527]_ , \new_[7528]_ ,
    \new_[7529]_ , \new_[7530]_ , \new_[7531]_ , \new_[7532]_ ,
    \new_[7533]_ , \new_[7534]_ , \new_[7535]_ , \new_[7536]_ ,
    \new_[7537]_ , \new_[7538]_ , \new_[7539]_ , \new_[7540]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7543]_ , \new_[7544]_ ,
    \new_[7545]_ , \new_[7546]_ , \new_[7547]_ , \new_[7548]_ ,
    \new_[7549]_ , \new_[7550]_ , \new_[7551]_ , \new_[7552]_ ,
    \new_[7553]_ , \new_[7554]_ , \new_[7555]_ , \new_[7556]_ ,
    \new_[7557]_ , \new_[7558]_ , \new_[7559]_ , \new_[7560]_ ,
    \new_[7561]_ , \new_[7562]_ , \new_[7563]_ , \new_[7564]_ ,
    \new_[7565]_ , \new_[7566]_ , \new_[7568]_ , \new_[7569]_ ,
    \new_[7570]_ , \new_[7571]_ , \new_[7572]_ , \new_[7573]_ ,
    \new_[7574]_ , \new_[7575]_ , \new_[7576]_ , \new_[7577]_ ,
    \new_[7578]_ , \new_[7579]_ , \new_[7580]_ , \new_[7581]_ ,
    \new_[7582]_ , \new_[7583]_ , \new_[7584]_ , \new_[7585]_ ,
    \new_[7586]_ , \new_[7587]_ , \new_[7588]_ , \new_[7589]_ ,
    \new_[7590]_ , \new_[7591]_ , \new_[7592]_ , \new_[7593]_ ,
    \new_[7594]_ , \new_[7595]_ , \new_[7596]_ , \new_[7597]_ ,
    \new_[7598]_ , \new_[7599]_ , \new_[7600]_ , \new_[7602]_ ,
    \new_[7603]_ , \new_[7604]_ , \new_[7605]_ , \new_[7606]_ ,
    \new_[7607]_ , \new_[7609]_ , \new_[7610]_ , \new_[7611]_ ,
    \new_[7612]_ , \new_[7613]_ , \new_[7614]_ , \new_[7615]_ ,
    \new_[7616]_ , \new_[7617]_ , \new_[7618]_ , \new_[7619]_ ,
    \new_[7620]_ , \new_[7621]_ , \new_[7622]_ , \new_[7623]_ ,
    \new_[7624]_ , \new_[7625]_ , \new_[7626]_ , \new_[7627]_ ,
    \new_[7628]_ , \new_[7629]_ , \new_[7631]_ , \new_[7632]_ ,
    \new_[7633]_ , \new_[7634]_ , \new_[7635]_ , \new_[7636]_ ,
    \new_[7637]_ , \new_[7638]_ , \new_[7639]_ , \new_[7640]_ ,
    \new_[7641]_ , \new_[7642]_ , \new_[7643]_ , \new_[7644]_ ,
    \new_[7645]_ , \new_[7646]_ , \new_[7647]_ , \new_[7648]_ ,
    \new_[7649]_ , \new_[7650]_ , \new_[7651]_ , \new_[7652]_ ,
    \new_[7653]_ , \new_[7654]_ , \new_[7655]_ , \new_[7656]_ ,
    \new_[7657]_ , \new_[7658]_ , \new_[7659]_ , \new_[7660]_ ,
    \new_[7661]_ , \new_[7662]_ , \new_[7663]_ , \new_[7664]_ ,
    \new_[7665]_ , \new_[7666]_ , \new_[7667]_ , \new_[7668]_ ,
    \new_[7669]_ , \new_[7670]_ , \new_[7671]_ , \new_[7672]_ ,
    \new_[7673]_ , \new_[7674]_ , \new_[7675]_ , \new_[7676]_ ,
    \new_[7677]_ , \new_[7678]_ , \new_[7679]_ , \new_[7680]_ ,
    \new_[7681]_ , \new_[7682]_ , \new_[7683]_ , \new_[7684]_ ,
    \new_[7685]_ , \new_[7686]_ , \new_[7687]_ , \new_[7688]_ ,
    \new_[7689]_ , \new_[7690]_ , \new_[7691]_ , \new_[7692]_ ,
    \new_[7693]_ , \new_[7694]_ , \new_[7695]_ , \new_[7696]_ ,
    \new_[7697]_ , \new_[7698]_ , \new_[7699]_ , \new_[7700]_ ,
    \new_[7701]_ , \new_[7702]_ , \new_[7703]_ , \new_[7704]_ ,
    \new_[7705]_ , \new_[7706]_ , \new_[7707]_ , \new_[7708]_ ,
    \new_[7709]_ , \new_[7710]_ , \new_[7711]_ , \new_[7712]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7715]_ , \new_[7716]_ ,
    \new_[7717]_ , \new_[7718]_ , \new_[7719]_ , \new_[7720]_ ,
    \new_[7721]_ , \new_[7722]_ , \new_[7723]_ , \new_[7724]_ ,
    \new_[7725]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7733]_ , \new_[7734]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7737]_ , \new_[7738]_ , \new_[7739]_ , \new_[7740]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7748]_ ,
    \new_[7749]_ , \new_[7750]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7754]_ , \new_[7755]_ , \new_[7756]_ ,
    \new_[7757]_ , \new_[7758]_ , \new_[7759]_ , \new_[7760]_ ,
    \new_[7761]_ , \new_[7762]_ , \new_[7763]_ , \new_[7764]_ ,
    \new_[7765]_ , \new_[7766]_ , \new_[7767]_ , \new_[7768]_ ,
    \new_[7769]_ , \new_[7770]_ , \new_[7771]_ , \new_[7772]_ ,
    \new_[7773]_ , \new_[7774]_ , \new_[7775]_ , \new_[7776]_ ,
    \new_[7777]_ , \new_[7778]_ , \new_[7779]_ , \new_[7780]_ ,
    \new_[7781]_ , \new_[7782]_ , \new_[7783]_ , \new_[7784]_ ,
    \new_[7785]_ , \new_[7786]_ , \new_[7787]_ , \new_[7788]_ ,
    \new_[7789]_ , \new_[7790]_ , \new_[7791]_ , \new_[7792]_ ,
    \new_[7793]_ , \new_[7794]_ , \new_[7795]_ , \new_[7796]_ ,
    \new_[7797]_ , \new_[7798]_ , \new_[7799]_ , \new_[7800]_ ,
    \new_[7801]_ , \new_[7802]_ , \new_[7803]_ , \new_[7804]_ ,
    \new_[7805]_ , \new_[7806]_ , \new_[7807]_ , \new_[7808]_ ,
    \new_[7809]_ , \new_[7810]_ , \new_[7811]_ , \new_[7812]_ ,
    \new_[7813]_ , \new_[7814]_ , \new_[7815]_ , \new_[7816]_ ,
    \new_[7817]_ , \new_[7818]_ , \new_[7819]_ , \new_[7820]_ ,
    \new_[7821]_ , \new_[7822]_ , \new_[7823]_ , \new_[7824]_ ,
    \new_[7825]_ , \new_[7826]_ , \new_[7827]_ , \new_[7828]_ ,
    \new_[7829]_ , \new_[7830]_ , \new_[7831]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7834]_ , \new_[7835]_ , \new_[7836]_ ,
    \new_[7837]_ , \new_[7838]_ , \new_[7839]_ , \new_[7840]_ ,
    \new_[7841]_ , \new_[7842]_ , \new_[7843]_ , \new_[7844]_ ,
    \new_[7845]_ , \new_[7846]_ , \new_[7847]_ , \new_[7848]_ ,
    \new_[7849]_ , \new_[7850]_ , \new_[7851]_ , \new_[7852]_ ,
    \new_[7853]_ , \new_[7854]_ , \new_[7855]_ , \new_[7856]_ ,
    \new_[7857]_ , \new_[7858]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7863]_ , \new_[7864]_ ,
    \new_[7865]_ , \new_[7866]_ , \new_[7867]_ , \new_[7868]_ ,
    \new_[7869]_ , \new_[7870]_ , \new_[7871]_ , \new_[7872]_ ,
    \new_[7873]_ , \new_[7874]_ , \new_[7875]_ , \new_[7876]_ ,
    \new_[7877]_ , \new_[7878]_ , \new_[7879]_ , \new_[7880]_ ,
    \new_[7881]_ , \new_[7882]_ , \new_[7883]_ , \new_[7884]_ ,
    \new_[7885]_ , \new_[7886]_ , \new_[7887]_ , \new_[7888]_ ,
    \new_[7889]_ , \new_[7890]_ , \new_[7891]_ , \new_[7892]_ ,
    \new_[7893]_ , \new_[7894]_ , \new_[7895]_ , \new_[7896]_ ,
    \new_[7897]_ , \new_[7898]_ , \new_[7899]_ , \new_[7900]_ ,
    \new_[7901]_ , \new_[7902]_ , \new_[7903]_ , \new_[7904]_ ,
    \new_[7905]_ , \new_[7906]_ , \new_[7907]_ , \new_[7908]_ ,
    \new_[7909]_ , \new_[7910]_ , \new_[7911]_ , \new_[7912]_ ,
    \new_[7913]_ , \new_[7914]_ , \new_[7915]_ , \new_[7916]_ ,
    \new_[7917]_ , \new_[7918]_ , \new_[7919]_ , \new_[7920]_ ,
    \new_[7921]_ , \new_[7922]_ , \new_[7923]_ , \new_[7924]_ ,
    \new_[7925]_ , \new_[7926]_ , \new_[7927]_ , \new_[7928]_ ,
    \new_[7929]_ , \new_[7930]_ , \new_[7931]_ , \new_[7932]_ ,
    \new_[7933]_ , \new_[7934]_ , \new_[7935]_ , \new_[7936]_ ,
    \new_[7937]_ , \new_[7938]_ , \new_[7939]_ , \new_[7940]_ ,
    \new_[7941]_ , \new_[7942]_ , \new_[7943]_ , \new_[7944]_ ,
    \new_[7945]_ , \new_[7946]_ , \new_[7947]_ , \new_[7948]_ ,
    \new_[7949]_ , \new_[7950]_ , \new_[7951]_ , \new_[7952]_ ,
    \new_[7953]_ , \new_[7954]_ , \new_[7955]_ , \new_[7956]_ ,
    \new_[7957]_ , \new_[7958]_ , \new_[7959]_ , \new_[7960]_ ,
    \new_[7961]_ , \new_[7962]_ , \new_[7963]_ , \new_[7964]_ ,
    \new_[7965]_ , \new_[7966]_ , \new_[7967]_ , \new_[7968]_ ,
    \new_[7969]_ , \new_[7970]_ , \new_[7971]_ , \new_[7972]_ ,
    \new_[7973]_ , \new_[7974]_ , \new_[7975]_ , \new_[7976]_ ,
    \new_[7977]_ , \new_[7978]_ , \new_[7979]_ , \new_[7980]_ ,
    \new_[7981]_ , \new_[7982]_ , \new_[7983]_ , \new_[7984]_ ,
    \new_[7985]_ , \new_[7986]_ , \new_[7987]_ , \new_[7988]_ ,
    \new_[7989]_ , \new_[7990]_ , \new_[7991]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7994]_ , \new_[7995]_ , \new_[7996]_ ,
    \new_[7997]_ , \new_[7998]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8005]_ , \new_[8006]_ , \new_[8007]_ , \new_[8008]_ ,
    \new_[8009]_ , \new_[8010]_ , \new_[8011]_ , \new_[8012]_ ,
    \new_[8013]_ , \new_[8014]_ , \new_[8015]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8018]_ , \new_[8019]_ , \new_[8020]_ ,
    \new_[8021]_ , \new_[8022]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8025]_ , \new_[8026]_ , \new_[8027]_ , \new_[8028]_ ,
    \new_[8029]_ , \new_[8030]_ , \new_[8031]_ , \new_[8032]_ ,
    \new_[8033]_ , \new_[8034]_ , \new_[8035]_ , \new_[8036]_ ,
    \new_[8037]_ , \new_[8038]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8041]_ , \new_[8042]_ , \new_[8043]_ , \new_[8044]_ ,
    \new_[8045]_ , \new_[8046]_ , \new_[8047]_ , \new_[8048]_ ,
    \new_[8049]_ , \new_[8050]_ , \new_[8051]_ , \new_[8052]_ ,
    \new_[8053]_ , \new_[8054]_ , \new_[8055]_ , \new_[8056]_ ,
    \new_[8057]_ , \new_[8058]_ , \new_[8059]_ , \new_[8060]_ ,
    \new_[8061]_ , \new_[8062]_ , \new_[8063]_ , \new_[8064]_ ,
    \new_[8065]_ , \new_[8066]_ , \new_[8067]_ , \new_[8068]_ ,
    \new_[8069]_ , \new_[8070]_ , \new_[8071]_ , \new_[8072]_ ,
    \new_[8073]_ , \new_[8074]_ , \new_[8075]_ , \new_[8076]_ ,
    \new_[8077]_ , \new_[8078]_ , \new_[8079]_ , \new_[8080]_ ,
    \new_[8081]_ , \new_[8082]_ , \new_[8083]_ , \new_[8084]_ ,
    \new_[8085]_ , \new_[8086]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8089]_ , \new_[8090]_ , \new_[8091]_ , \new_[8092]_ ,
    \new_[8093]_ , \new_[8094]_ , \new_[8095]_ , \new_[8096]_ ,
    \new_[8097]_ , \new_[8098]_ , \new_[8099]_ , \new_[8100]_ ,
    \new_[8101]_ , \new_[8102]_ , \new_[8103]_ , \new_[8104]_ ,
    \new_[8105]_ , \new_[8106]_ , \new_[8107]_ , \new_[8108]_ ,
    \new_[8109]_ , \new_[8110]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8113]_ , \new_[8114]_ , \new_[8115]_ , \new_[8116]_ ,
    \new_[8117]_ , \new_[8118]_ , \new_[8119]_ , \new_[8120]_ ,
    \new_[8121]_ , \new_[8122]_ , \new_[8123]_ , \new_[8124]_ ,
    \new_[8125]_ , \new_[8126]_ , \new_[8127]_ , \new_[8128]_ ,
    \new_[8129]_ , \new_[8130]_ , \new_[8131]_ , \new_[8132]_ ,
    \new_[8133]_ , \new_[8134]_ , \new_[8135]_ , \new_[8136]_ ,
    \new_[8137]_ , \new_[8138]_ , \new_[8139]_ , \new_[8140]_ ,
    \new_[8141]_ , \new_[8142]_ , \new_[8143]_ , \new_[8144]_ ,
    \new_[8145]_ , \new_[8146]_ , \new_[8147]_ , \new_[8148]_ ,
    \new_[8149]_ , \new_[8150]_ , \new_[8151]_ , \new_[8152]_ ,
    \new_[8153]_ , \new_[8154]_ , \new_[8155]_ , \new_[8156]_ ,
    \new_[8157]_ , \new_[8158]_ , \new_[8159]_ , \new_[8160]_ ,
    \new_[8161]_ , \new_[8162]_ , \new_[8163]_ , \new_[8164]_ ,
    \new_[8165]_ , \new_[8166]_ , \new_[8167]_ , \new_[8168]_ ,
    \new_[8169]_ , \new_[8170]_ , \new_[8171]_ , \new_[8172]_ ,
    \new_[8173]_ , \new_[8174]_ , \new_[8175]_ , \new_[8176]_ ,
    \new_[8177]_ , \new_[8178]_ , \new_[8179]_ , \new_[8180]_ ,
    \new_[8181]_ , \new_[8182]_ , \new_[8183]_ , \new_[8184]_ ,
    \new_[8185]_ , \new_[8186]_ , \new_[8187]_ , \new_[8188]_ ,
    \new_[8189]_ , \new_[8190]_ , \new_[8191]_ , \new_[8192]_ ,
    \new_[8193]_ , \new_[8194]_ , \new_[8195]_ , \new_[8196]_ ,
    \new_[8197]_ , \new_[8198]_ , \new_[8199]_ , \new_[8201]_ ,
    \new_[8202]_ , \new_[8203]_ , \new_[8204]_ , \new_[8205]_ ,
    \new_[8206]_ , \new_[8207]_ , \new_[8208]_ , \new_[8209]_ ,
    \new_[8210]_ , \new_[8211]_ , \new_[8212]_ , \new_[8213]_ ,
    \new_[8214]_ , \new_[8215]_ , \new_[8216]_ , \new_[8217]_ ,
    \new_[8218]_ , \new_[8219]_ , \new_[8220]_ , \new_[8221]_ ,
    \new_[8222]_ , \new_[8223]_ , \new_[8224]_ , \new_[8225]_ ,
    \new_[8226]_ , \new_[8227]_ , \new_[8228]_ , \new_[8229]_ ,
    \new_[8230]_ , \new_[8231]_ , \new_[8232]_ , \new_[8233]_ ,
    \new_[8234]_ , \new_[8235]_ , \new_[8236]_ , \new_[8237]_ ,
    \new_[8238]_ , \new_[8239]_ , \new_[8240]_ , \new_[8241]_ ,
    \new_[8242]_ , \new_[8243]_ , \new_[8244]_ , \new_[8245]_ ,
    \new_[8246]_ , \new_[8247]_ , \new_[8248]_ , \new_[8249]_ ,
    \new_[8250]_ , \new_[8251]_ , \new_[8252]_ , \new_[8253]_ ,
    \new_[8254]_ , \new_[8255]_ , \new_[8256]_ , \new_[8257]_ ,
    \new_[8258]_ , \new_[8259]_ , \new_[8260]_ , \new_[8261]_ ,
    \new_[8262]_ , \new_[8263]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8266]_ , \new_[8267]_ , \new_[8268]_ , \new_[8269]_ ,
    \new_[8270]_ , \new_[8271]_ , \new_[8272]_ , \new_[8273]_ ,
    \new_[8274]_ , \new_[8275]_ , \new_[8276]_ , \new_[8277]_ ,
    \new_[8278]_ , \new_[8279]_ , \new_[8280]_ , \new_[8281]_ ,
    \new_[8282]_ , \new_[8283]_ , \new_[8284]_ , \new_[8285]_ ,
    \new_[8286]_ , \new_[8287]_ , \new_[8288]_ , \new_[8289]_ ,
    \new_[8290]_ , \new_[8291]_ , \new_[8292]_ , \new_[8293]_ ,
    \new_[8294]_ , \new_[8295]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8302]_ , \new_[8303]_ , \new_[8304]_ , \new_[8305]_ ,
    \new_[8306]_ , \new_[8307]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8310]_ , \new_[8311]_ , \new_[8312]_ , \new_[8313]_ ,
    \new_[8314]_ , \new_[8315]_ , \new_[8316]_ , \new_[8317]_ ,
    \new_[8319]_ , \new_[8320]_ , \new_[8321]_ , \new_[8322]_ ,
    \new_[8323]_ , \new_[8324]_ , \new_[8325]_ , \new_[8326]_ ,
    \new_[8327]_ , \new_[8328]_ , \new_[8329]_ , \new_[8330]_ ,
    \new_[8331]_ , \new_[8332]_ , \new_[8333]_ , \new_[8334]_ ,
    \new_[8335]_ , \new_[8336]_ , \new_[8337]_ , \new_[8338]_ ,
    \new_[8339]_ , \new_[8341]_ , \new_[8342]_ , \new_[8343]_ ,
    \new_[8344]_ , \new_[8345]_ , \new_[8346]_ , \new_[8347]_ ,
    \new_[8348]_ , \new_[8349]_ , \new_[8350]_ , \new_[8351]_ ,
    \new_[8352]_ , \new_[8353]_ , \new_[8354]_ , \new_[8355]_ ,
    \new_[8356]_ , \new_[8357]_ , \new_[8358]_ , \new_[8359]_ ,
    \new_[8360]_ , \new_[8361]_ , \new_[8362]_ , \new_[8363]_ ,
    \new_[8364]_ , \new_[8365]_ , \new_[8366]_ , \new_[8367]_ ,
    \new_[8368]_ , \new_[8369]_ , \new_[8370]_ , \new_[8371]_ ,
    \new_[8372]_ , \new_[8373]_ , \new_[8374]_ , \new_[8375]_ ,
    \new_[8376]_ , \new_[8377]_ , \new_[8378]_ , \new_[8379]_ ,
    \new_[8380]_ , \new_[8381]_ , \new_[8382]_ , \new_[8383]_ ,
    \new_[8384]_ , \new_[8385]_ , \new_[8386]_ , \new_[8387]_ ,
    \new_[8388]_ , \new_[8389]_ , \new_[8390]_ , \new_[8391]_ ,
    \new_[8392]_ , \new_[8393]_ , \new_[8394]_ , \new_[8395]_ ,
    \new_[8396]_ , \new_[8397]_ , \new_[8398]_ , \new_[8399]_ ,
    \new_[8400]_ , \new_[8401]_ , \new_[8402]_ , \new_[8403]_ ,
    \new_[8404]_ , \new_[8405]_ , \new_[8406]_ , \new_[8408]_ ,
    \new_[8409]_ , \new_[8410]_ , \new_[8411]_ , \new_[8412]_ ,
    \new_[8413]_ , \new_[8414]_ , \new_[8415]_ , \new_[8416]_ ,
    \new_[8417]_ , \new_[8418]_ , \new_[8419]_ , \new_[8420]_ ,
    \new_[8421]_ , \new_[8422]_ , \new_[8423]_ , \new_[8424]_ ,
    \new_[8425]_ , \new_[8426]_ , \new_[8427]_ , \new_[8428]_ ,
    \new_[8429]_ , \new_[8430]_ , \new_[8431]_ , \new_[8432]_ ,
    \new_[8433]_ , \new_[8434]_ , \new_[8435]_ , \new_[8436]_ ,
    \new_[8437]_ , \new_[8438]_ , \new_[8439]_ , \new_[8440]_ ,
    \new_[8441]_ , \new_[8442]_ , \new_[8443]_ , \new_[8444]_ ,
    \new_[8445]_ , \new_[8446]_ , \new_[8447]_ , \new_[8448]_ ,
    \new_[8449]_ , \new_[8450]_ , \new_[8451]_ , \new_[8452]_ ,
    \new_[8453]_ , \new_[8454]_ , \new_[8455]_ , \new_[8456]_ ,
    \new_[8457]_ , \new_[8458]_ , \new_[8459]_ , \new_[8460]_ ,
    \new_[8461]_ , \new_[8462]_ , \new_[8463]_ , \new_[8464]_ ,
    \new_[8465]_ , \new_[8466]_ , \new_[8467]_ , \new_[8468]_ ,
    \new_[8469]_ , \new_[8470]_ , \new_[8471]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8474]_ , \new_[8475]_ , \new_[8476]_ ,
    \new_[8477]_ , \new_[8478]_ , \new_[8479]_ , \new_[8480]_ ,
    \new_[8481]_ , \new_[8482]_ , \new_[8483]_ , \new_[8484]_ ,
    \new_[8485]_ , \new_[8486]_ , \new_[8487]_ , \new_[8488]_ ,
    \new_[8489]_ , \new_[8490]_ , \new_[8491]_ , \new_[8492]_ ,
    \new_[8493]_ , \new_[8494]_ , \new_[8495]_ , \new_[8496]_ ,
    \new_[8497]_ , \new_[8498]_ , \new_[8499]_ , \new_[8500]_ ,
    \new_[8501]_ , \new_[8502]_ , \new_[8503]_ , \new_[8504]_ ,
    \new_[8505]_ , \new_[8506]_ , \new_[8507]_ , \new_[8508]_ ,
    \new_[8509]_ , \new_[8510]_ , \new_[8511]_ , \new_[8512]_ ,
    \new_[8513]_ , \new_[8514]_ , \new_[8515]_ , \new_[8516]_ ,
    \new_[8517]_ , \new_[8518]_ , \new_[8519]_ , \new_[8520]_ ,
    \new_[8521]_ , \new_[8522]_ , \new_[8523]_ , \new_[8524]_ ,
    \new_[8525]_ , \new_[8526]_ , \new_[8527]_ , \new_[8528]_ ,
    \new_[8529]_ , \new_[8530]_ , \new_[8531]_ , \new_[8532]_ ,
    \new_[8533]_ , \new_[8534]_ , \new_[8535]_ , \new_[8536]_ ,
    \new_[8537]_ , \new_[8538]_ , \new_[8539]_ , \new_[8540]_ ,
    \new_[8541]_ , \new_[8543]_ , \new_[8544]_ , \new_[8546]_ ,
    \new_[8547]_ , \new_[8548]_ , \new_[8550]_ , \new_[8551]_ ,
    \new_[8553]_ , \new_[8554]_ , \new_[8555]_ , \new_[8556]_ ,
    \new_[8557]_ , \new_[8558]_ , \new_[8559]_ , \new_[8560]_ ,
    \new_[8561]_ , \new_[8562]_ , \new_[8563]_ , \new_[8564]_ ,
    \new_[8565]_ , \new_[8566]_ , \new_[8567]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8570]_ , \new_[8571]_ , \new_[8572]_ ,
    \new_[8573]_ , \new_[8575]_ , \new_[8576]_ , \new_[8578]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8581]_ , \new_[8582]_ ,
    \new_[8583]_ , \new_[8584]_ , \new_[8585]_ , \new_[8586]_ ,
    \new_[8587]_ , \new_[8588]_ , \new_[8589]_ , \new_[8590]_ ,
    \new_[8591]_ , \new_[8592]_ , \new_[8593]_ , \new_[8594]_ ,
    \new_[8595]_ , \new_[8597]_ , \new_[8598]_ , \new_[8599]_ ,
    \new_[8600]_ , \new_[8601]_ , \new_[8602]_ , \new_[8603]_ ,
    \new_[8604]_ , \new_[8605]_ , \new_[8607]_ , \new_[8608]_ ,
    \new_[8609]_ , \new_[8610]_ , \new_[8611]_ , \new_[8612]_ ,
    \new_[8613]_ , \new_[8614]_ , \new_[8615]_ , \new_[8617]_ ,
    \new_[8618]_ , \new_[8619]_ , \new_[8620]_ , \new_[8621]_ ,
    \new_[8622]_ , \new_[8623]_ , \new_[8624]_ , \new_[8625]_ ,
    \new_[8626]_ , \new_[8627]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8631]_ , \new_[8632]_ , \new_[8633]_ , \new_[8634]_ ,
    \new_[8635]_ , \new_[8636]_ , \new_[8637]_ , \new_[8638]_ ,
    \new_[8639]_ , \new_[8640]_ , \new_[8641]_ , \new_[8642]_ ,
    \new_[8643]_ , \new_[8644]_ , \new_[8645]_ , \new_[8646]_ ,
    \new_[8647]_ , \new_[8648]_ , \new_[8650]_ , \new_[8651]_ ,
    \new_[8652]_ , \new_[8653]_ , \new_[8654]_ , \new_[8655]_ ,
    \new_[8656]_ , \new_[8657]_ , \new_[8658]_ , \new_[8659]_ ,
    \new_[8660]_ , \new_[8661]_ , \new_[8662]_ , \new_[8663]_ ,
    \new_[8664]_ , \new_[8665]_ , \new_[8666]_ , \new_[8667]_ ,
    \new_[8668]_ , \new_[8669]_ , \new_[8670]_ , \new_[8671]_ ,
    \new_[8672]_ , \new_[8673]_ , \new_[8674]_ , \new_[8675]_ ,
    \new_[8676]_ , \new_[8677]_ , \new_[8678]_ , \new_[8679]_ ,
    \new_[8680]_ , \new_[8681]_ , \new_[8682]_ , \new_[8683]_ ,
    \new_[8684]_ , \new_[8685]_ , \new_[8686]_ , \new_[8687]_ ,
    \new_[8688]_ , \new_[8689]_ , \new_[8690]_ , \new_[8691]_ ,
    \new_[8692]_ , \new_[8693]_ , \new_[8694]_ , \new_[8695]_ ,
    \new_[8696]_ , \new_[8697]_ , \new_[8698]_ , \new_[8699]_ ,
    \new_[8700]_ , \new_[8701]_ , \new_[8702]_ , \new_[8703]_ ,
    \new_[8704]_ , \new_[8705]_ , \new_[8706]_ , \new_[8707]_ ,
    \new_[8708]_ , \new_[8709]_ , \new_[8710]_ , \new_[8711]_ ,
    \new_[8712]_ , \new_[8713]_ , \new_[8714]_ , \new_[8715]_ ,
    \new_[8716]_ , \new_[8717]_ , \new_[8718]_ , \new_[8719]_ ,
    \new_[8720]_ , \new_[8721]_ , \new_[8722]_ , \new_[8723]_ ,
    \new_[8724]_ , \new_[8725]_ , \new_[8726]_ , \new_[8727]_ ,
    \new_[8728]_ , \new_[8729]_ , \new_[8730]_ , \new_[8731]_ ,
    \new_[8732]_ , \new_[8733]_ , \new_[8734]_ , \new_[8735]_ ,
    \new_[8736]_ , \new_[8737]_ , \new_[8738]_ , \new_[8739]_ ,
    \new_[8740]_ , \new_[8741]_ , \new_[8742]_ , \new_[8743]_ ,
    \new_[8744]_ , \new_[8745]_ , \new_[8746]_ , \new_[8747]_ ,
    \new_[8748]_ , \new_[8749]_ , \new_[8750]_ , \new_[8751]_ ,
    \new_[8752]_ , \new_[8753]_ , \new_[8754]_ , \new_[8755]_ ,
    \new_[8756]_ , \new_[8757]_ , \new_[8758]_ , \new_[8759]_ ,
    \new_[8760]_ , \new_[8761]_ , \new_[8762]_ , \new_[8763]_ ,
    \new_[8764]_ , \new_[8765]_ , \new_[8766]_ , \new_[8767]_ ,
    \new_[8768]_ , \new_[8769]_ , \new_[8770]_ , \new_[8771]_ ,
    \new_[8772]_ , \new_[8773]_ , \new_[8774]_ , \new_[8775]_ ,
    \new_[8776]_ , \new_[8777]_ , \new_[8778]_ , \new_[8779]_ ,
    \new_[8780]_ , \new_[8781]_ , \new_[8782]_ , \new_[8783]_ ,
    \new_[8784]_ , \new_[8785]_ , \new_[8786]_ , \new_[8787]_ ,
    \new_[8788]_ , \new_[8789]_ , \new_[8790]_ , \new_[8791]_ ,
    \new_[8792]_ , \new_[8793]_ , \new_[8794]_ , \new_[8795]_ ,
    \new_[8796]_ , \new_[8797]_ , \new_[8798]_ , \new_[8799]_ ,
    \new_[8800]_ , \new_[8801]_ , \new_[8802]_ , \new_[8803]_ ,
    \new_[8804]_ , \new_[8805]_ , \new_[8806]_ , \new_[8807]_ ,
    \new_[8808]_ , \new_[8809]_ , \new_[8810]_ , \new_[8811]_ ,
    \new_[8812]_ , \new_[8813]_ , \new_[8814]_ , \new_[8815]_ ,
    \new_[8816]_ , \new_[8817]_ , \new_[8818]_ , \new_[8819]_ ,
    \new_[8820]_ , \new_[8821]_ , \new_[8822]_ , \new_[8823]_ ,
    \new_[8824]_ , \new_[8825]_ , \new_[8826]_ , \new_[8827]_ ,
    \new_[8828]_ , \new_[8829]_ , \new_[8830]_ , \new_[8831]_ ,
    \new_[8832]_ , \new_[8833]_ , \new_[8834]_ , \new_[8835]_ ,
    \new_[8836]_ , \new_[8837]_ , \new_[8839]_ , \new_[8840]_ ,
    \new_[8841]_ , \new_[8842]_ , \new_[8843]_ , \new_[8844]_ ,
    \new_[8845]_ , \new_[8847]_ , \new_[8848]_ , \new_[8849]_ ,
    \new_[8850]_ , \new_[8851]_ , \new_[8852]_ , \new_[8853]_ ,
    \new_[8854]_ , \new_[8855]_ , \new_[8856]_ , \new_[8857]_ ,
    \new_[8858]_ , \new_[8859]_ , \new_[8860]_ , \new_[8861]_ ,
    \new_[8862]_ , \new_[8863]_ , \new_[8864]_ , \new_[8865]_ ,
    \new_[8866]_ , \new_[8867]_ , \new_[8868]_ , \new_[8869]_ ,
    \new_[8870]_ , \new_[8871]_ , \new_[8872]_ , \new_[8873]_ ,
    \new_[8874]_ , \new_[8875]_ , \new_[8876]_ , \new_[8877]_ ,
    \new_[8878]_ , \new_[8879]_ , \new_[8880]_ , \new_[8881]_ ,
    \new_[8882]_ , \new_[8883]_ , \new_[8884]_ , \new_[8885]_ ,
    \new_[8886]_ , \new_[8887]_ , \new_[8888]_ , \new_[8889]_ ,
    \new_[8890]_ , \new_[8891]_ , \new_[8892]_ , \new_[8893]_ ,
    \new_[8894]_ , \new_[8895]_ , \new_[8896]_ , \new_[8897]_ ,
    \new_[8898]_ , \new_[8899]_ , \new_[8900]_ , \new_[8901]_ ,
    \new_[8902]_ , \new_[8903]_ , \new_[8904]_ , \new_[8905]_ ,
    \new_[8906]_ , \new_[8907]_ , \new_[8908]_ , \new_[8909]_ ,
    \new_[8910]_ , \new_[8911]_ , \new_[8912]_ , \new_[8913]_ ,
    \new_[8914]_ , \new_[8915]_ , \new_[8916]_ , \new_[8917]_ ,
    \new_[8918]_ , \new_[8919]_ , \new_[8920]_ , \new_[8921]_ ,
    \new_[8922]_ , \new_[8923]_ , \new_[8924]_ , \new_[8925]_ ,
    \new_[8926]_ , \new_[8927]_ , \new_[8928]_ , \new_[8929]_ ,
    \new_[8930]_ , \new_[8931]_ , \new_[8932]_ , \new_[8933]_ ,
    \new_[8934]_ , \new_[8935]_ , \new_[8936]_ , \new_[8937]_ ,
    \new_[8938]_ , \new_[8939]_ , \new_[8940]_ , \new_[8941]_ ,
    \new_[8942]_ , \new_[8943]_ , \new_[8944]_ , \new_[8945]_ ,
    \new_[8946]_ , \new_[8947]_ , \new_[8948]_ , \new_[8949]_ ,
    \new_[8950]_ , \new_[8951]_ , \new_[8952]_ , \new_[8953]_ ,
    \new_[8954]_ , \new_[8955]_ , \new_[8956]_ , \new_[8957]_ ,
    \new_[8958]_ , \new_[8959]_ , \new_[8960]_ , \new_[8961]_ ,
    \new_[8962]_ , \new_[8963]_ , \new_[8964]_ , \new_[8965]_ ,
    \new_[8966]_ , \new_[8967]_ , \new_[8968]_ , \new_[8969]_ ,
    \new_[8970]_ , \new_[8971]_ , \new_[8972]_ , \new_[8973]_ ,
    \new_[8974]_ , \new_[8975]_ , \new_[8976]_ , \new_[8977]_ ,
    \new_[8978]_ , \new_[8979]_ , \new_[8981]_ , \new_[8982]_ ,
    \new_[8983]_ , \new_[8984]_ , \new_[8985]_ , \new_[8986]_ ,
    \new_[8987]_ , \new_[8988]_ , \new_[8989]_ , \new_[8990]_ ,
    \new_[8991]_ , \new_[8992]_ , \new_[8993]_ , \new_[8994]_ ,
    \new_[8995]_ , \new_[8996]_ , \new_[8997]_ , \new_[8998]_ ,
    \new_[8999]_ , \new_[9000]_ , \new_[9001]_ , \new_[9002]_ ,
    \new_[9003]_ , \new_[9004]_ , \new_[9005]_ , \new_[9006]_ ,
    \new_[9007]_ , \new_[9008]_ , \new_[9009]_ , \new_[9010]_ ,
    \new_[9011]_ , \new_[9013]_ , \new_[9014]_ , \new_[9015]_ ,
    \new_[9016]_ , \new_[9017]_ , \new_[9018]_ , \new_[9019]_ , n780, n785,
    n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840, n845,
    n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900, n905,
    n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960, n965,
    n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015, n1020,
    n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070,
    n1075, n1080, n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1120,
    n1125, n1130, n1135, n1140, n1145, n1150, n1155, n1160, n1165, n1170,
    n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220,
    n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270,
    n1275, n1280, n1285, n1290, n1295, n1300, n1305, n1310, n1315, n1320,
    n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365, n1370,
    n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415, n1420,
    n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465, n1470,
    n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515, n1520,
    n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570,
    n1575, n1580, n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620,
    n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670,
    n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720,
    n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770,
    n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820,
    n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870,
    n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920,
    n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970,
    n1975, n1980, n1985, n1990, n1995, n2000, n2005, n2010, n2015, n2020,
    n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070,
    n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120,
    n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165, n2170,
    n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210, n2215, n2220,
    n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260, n2265, n2270,
    n2275, n2280, n2285, n2290, n2295, n2300, n2305, n2310, n2315, n2320,
    n2325, n2330, n2335, n2340, n2345, n2350, n2355, n2360, n2365, n2370,
    n2375, n2380, n2385, n2390, n2395, n2400, n2405, n2410, n2415, n2420,
    n2425, n2430, n2435, n2440, n2445, n2450, n2455, n2460, n2465, n2470,
    n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520,
    n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570,
    n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620,
    n2625, n2630, n2635, n2640, n2645, n2650, n2655, n2660, n2665, n2670,
    n2675, n2680, n2685, n2690, n2695, n2700, n2705, n2710, n2715, n2720,
    n2725, n2730, n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770,
    n2775, n2780, n2785, n2790, n2795, n2800, n2805, n2810, n2815, n2820,
    n2825, n2830, n2835, n2840, n2845, n2850, n2855, n2860, n2865, n2870,
    n2875, n2880, n2885, n2890, n2895, n2900, n2905, n2910, n2915, n2920,
    n2925, n2930, n2935, n2940, n2945, n2950, n2955, n2960, n2965, n2970,
    n2975, n2980, n2985, n2990, n2995, n3000, n3005, n3010, n3015, n3020,
    n3025, n3030, n3035, n3040, n3045, n3050, n3055, n3060, n3065, n3070,
    n3075, n3080, n3085, n3090, n3095, n3100, n3105, n3110, n3115, n3120,
    n3125, n3130, n3135, n3140, n3145, n3150, n3155, n3160, n3165, n3170,
    n3175, n3180, n3185, n3190, n3195, n3200, n3205, n3210, n3215, n3220,
    n3225, n3230, n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270,
    n3275, n3280, n3285, n3290, n3295, n3300, n3305, n3310, n3315, n3320,
    n3325, n3330, n3335, n3340, n3345, n3350, n3355, n3360, n3365, n3370,
    n3375, n3380, n3385, n3390, n3395, n3400, n3405, n3410, n3415, n3420,
    n3425, n3430, n3435, n3440, n3445, n3450, n3455, n3460, n3465, n3470,
    n3475, n3480, n3485, n3490, n3495, n3500, n3505, n3510, n3515, n3520,
    n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570,
    n3575, n3580, n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620,
    n3625, n3630, n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670,
    n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720,
    n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770,
    n3775, n3780, n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820,
    n3825, n3830, n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3870,
    n3875, n3880, n3885, n3890, n3895, n3900, n3905, n3910, n3915, n3920,
    n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3960, n3965, n3970,
    n3975, n3980, n3985, n3990, n3995, n4000, n4005, n4010, n4015, n4020,
    n4025, n4030, n4035, n4040, n4045, n4050, n4055, n4060, n4065, n4070,
    n4075, n4080, n4085, n4090, n4095, n4100, n4105, n4110, n4115, n4120,
    n4125;
  assign \new_[1061]_  = \\ks1_key_reg_reg[11] ;
  assign \new_[1062]_  = \\ks1_key_reg_reg[12] ;
  assign \new_[1063]_  = \\ks1_key_reg_reg[13] ;
  assign \new_[1064]_  = \\ks1_key_reg_reg[14] ;
  assign \new_[1065]_  = \\ks1_key_reg_reg[15] ;
  assign \new_[1066]_  = \\sbox1_to_invert_reg[1] ;
  assign \new_[1067]_  = \\sbox1_to_invert_reg[3] ;
  assign \new_[1068]_  = \\sbox1_to_invert_reg[2] ;
  assign \new_[1069]_  = \\sbox1_to_invert_reg[0] ;
  assign \new_[1070]_  = \\ks1_key_reg_reg[8] ;
  assign n795 = ~\new_[1078]_  | ~\new_[7121]_ ;
  assign \new_[1072]_  = \\ks1_key_reg_reg[10] ;
  assign n805 = \new_[1297]_  ? \new_[1087]_  : \new_[1231]_ ;
  assign n810 = \new_[8642]_  ? \new_[1088]_  : \new_[1124]_ ;
  assign n815 = \new_[1093]_  ? \new_[1086]_  : \new_[1091]_ ;
  assign \new_[1076]_  = \\ks1_key_reg_reg[9] ;
  assign n825 = ~\new_[8844]_  | ~\new_[7113]_ ;
  assign \new_[1078]_  = ~\new_[8852]_  | ~\new_[1085]_ ;
  assign \new_[1079]_  = \\ks1_key_reg_reg[43] ;
  assign \new_[1080]_  = \\ks1_key_reg_reg[44] ;
  assign n830 = ~\new_[1090]_  | ~\new_[6936]_ ;
  assign \new_[1082]_  = \\ks1_key_reg_reg[45] ;
  assign \new_[1083]_  = \\ks1_key_reg_reg[46] ;
  assign \new_[1084]_  = \\ks1_key_reg_reg[47] ;
  assign \new_[1085]_  = ~\new_[1092]_  | (~n855 & ~\new_[8382]_ );
  assign \new_[1086]_  = \new_[1904]_  ? \new_[1121]_  : \new_[1882]_ ;
  assign \new_[1087]_  = \new_[1176]_  ? \new_[1120]_  : \new_[1129]_ ;
  assign \new_[1088]_  = \new_[1298]_  ? \new_[1122]_  : \new_[1357]_ ;
  assign \new_[1089]_  = \\ks1_key_reg_reg[40] ;
  assign \new_[1090]_  = ~\new_[1123]_  | ~n4105;
  assign \new_[1091]_  = ~\new_[1093]_ ;
  assign \new_[1092]_  = ~n855 | ~\new_[8382]_ ;
  assign \new_[1093]_  = \new_[8702]_  ? \new_[1177]_  : \new_[1454]_ ;
  assign \new_[1094]_  = \\sub1_data_reg_reg[109] ;
  assign \new_[1095]_  = \\sub1_data_reg_reg[110] ;
  assign \new_[1096]_  = \\sub1_data_reg_reg[13] ;
  assign \new_[1097]_  = \\sub1_data_reg_reg[14] ;
  assign \new_[1098]_  = \\sub1_data_reg_reg[45] ;
  assign \new_[1099]_  = \\sub1_data_reg_reg[46] ;
  assign \new_[1100]_  = \\sub1_data_reg_reg[77] ;
  assign \new_[1101]_  = \\sub1_data_reg_reg[78] ;
  assign \new_[1102]_  = \\sub1_data_reg_reg[102] ;
  assign \new_[1103]_  = \\sub1_data_reg_reg[101] ;
  assign \new_[1104]_  = \\sub1_data_reg_reg[118] ;
  assign \new_[1105]_  = \\sub1_data_reg_reg[117] ;
  assign \new_[1106]_  = \\sub1_data_reg_reg[21] ;
  assign \new_[1107]_  = \\sub1_data_reg_reg[22] ;
  assign \new_[1108]_  = \\sub1_data_reg_reg[37] ;
  assign \new_[1109]_  = \\sub1_data_reg_reg[38] ;
  assign \new_[1110]_  = \\sub1_data_reg_reg[53] ;
  assign \new_[1111]_  = \\sub1_data_reg_reg[54] ;
  assign \new_[1112]_  = \\sub1_data_reg_reg[5] ;
  assign \new_[1113]_  = \\sub1_data_reg_reg[6] ;
  assign \new_[1114]_  = \\sub1_data_reg_reg[70] ;
  assign \new_[1115]_  = \\sub1_data_reg_reg[69] ;
  assign \new_[1116]_  = \\sub1_data_reg_reg[85] ;
  assign \new_[1117]_  = \\sub1_data_reg_reg[86] ;
  assign \new_[1118]_  = \\ks1_key_reg_reg[42] ;
  assign \new_[1119]_  = \\ks1_key_reg_reg[41] ;
  assign \new_[1120]_  = ~\new_[1178]_  | ~\new_[1179]_ ;
  assign \new_[1121]_  = ~\new_[1180]_  | ~\new_[1182]_ ;
  assign \new_[1122]_  = ~\new_[1183]_  | ~\new_[1184]_ ;
  assign \new_[1123]_  = ~\new_[1185]_  | (~n990 & ~\new_[4619]_ );
  assign \new_[1124]_  = ~\new_[8642]_ ;
  assign \new_[1125]_  = \\ks1_key_reg_reg[76] ;
  assign \new_[1126]_  = \\ks1_key_reg_reg[75] ;
  assign \new_[1127]_  = ~\\ks1_key_reg_reg[74] ;
  assign \new_[1128]_  = ~\\ks1_key_reg_reg[73] ;
  assign \new_[1129]_  = ~\new_[1176]_ ;
  assign n855 = ~\new_[1228]_  | ~\new_[1280]_ ;
  assign n910 = ~\new_[1421]_  | ~\new_[1256]_ ;
  assign \new_[1132]_  = \\ks1_key_reg_reg[77] ;
  assign \new_[1133]_  = \\ks1_key_reg_reg[78] ;
  assign \new_[1134]_  = \\sub1_data_reg_reg[125] ;
  assign \new_[1135]_  = \\sub1_data_reg_reg[126] ;
  assign \new_[1136]_  = \\sub1_data_reg_reg[29] ;
  assign \new_[1137]_  = \\sub1_data_reg_reg[94] ;
  assign \new_[1138]_  = \\sub1_data_reg_reg[30] ;
  assign \new_[1139]_  = \\sub1_data_reg_reg[93] ;
  assign \new_[1140]_  = \\ks1_key_reg_reg[72] ;
  assign \new_[1141]_  = \\ks1_key_reg_reg[79] ;
  assign \new_[1142]_  = \\sub1_data_reg_reg[104] ;
  assign \new_[1143]_  = \\sub1_data_reg_reg[40] ;
  assign \new_[1144]_  = \\sub1_data_reg_reg[72] ;
  assign \new_[1145]_  = \\sub1_data_reg_reg[8] ;
  assign \new_[1146]_  = ~\\sub1_data_reg_reg[0] ;
  assign \new_[1147]_  = \\sub1_data_reg_reg[112] ;
  assign \new_[1148]_  = \\sub1_data_reg_reg[16] ;
  assign \new_[1149]_  = \\sub1_data_reg_reg[64] ;
  assign \new_[1150]_  = \\sub1_data_reg_reg[80] ;
  assign \new_[1151]_  = \\sub1_data_reg_reg[96] ;
  assign \new_[1152]_  = \\sub1_data_reg_reg[48] ;
  assign n915 = ~\new_[1419]_  | ~\new_[1255]_ ;
  assign n925 = ~\new_[6697]_  | ~\new_[1257]_ ;
  assign n920 = ~\new_[6695]_  | ~\new_[1258]_ ;
  assign n930 = ~\new_[6693]_  | ~\new_[1259]_ ;
  assign n935 = ~\new_[6696]_  | ~\new_[1260]_ ;
  assign n940 = ~\new_[1417]_  | ~\new_[1261]_ ;
  assign n945 = ~\new_[1416]_  | ~\new_[1262]_ ;
  assign n950 = ~\new_[6526]_  | ~\new_[1263]_ ;
  assign n955 = ~\new_[6524]_  | ~\new_[1264]_ ;
  assign n960 = ~\new_[6692]_  | ~\new_[1265]_ ;
  assign n965 = ~\new_[6691]_  | ~\new_[1267]_ ;
  assign n975 = ~\new_[6525]_  | ~\new_[1266]_ ;
  assign n970 = ~\new_[6527]_  | ~\new_[1268]_ ;
  assign n980 = ~\new_[6522]_  | ~\new_[1269]_ ;
  assign n985 = ~\new_[6523]_  | ~\new_[1270]_ ;
  assign n870 = ~\new_[1279]_  | ~\new_[6192]_ ;
  assign n875 = ~\new_[1281]_  | ~\new_[6191]_ ;
  assign n880 = ~\new_[1282]_  | ~\new_[6189]_ ;
  assign n885 = ~\new_[1283]_  | ~\new_[6188]_ ;
  assign n890 = ~\new_[1284]_  | ~\new_[6193]_ ;
  assign n895 = ~\new_[1285]_  | ~\new_[6190]_ ;
  assign n900 = ~\new_[1286]_  | ~\new_[6151]_ ;
  assign n905 = ~\new_[1287]_  | ~\new_[6194]_ ;
  assign \new_[1176]_  = \new_[1711]_  ? \new_[1355]_  : \new_[1594]_ ;
  assign \new_[1177]_  = \new_[1880]_  ? \new_[1356]_  : \new_[1846]_ ;
  assign \new_[1178]_  = ~\new_[1274]_  | ~\new_[1944]_ ;
  assign \new_[1179]_  = ~\new_[1272]_  | ~\new_[1932]_ ;
  assign \new_[1180]_  = ~\new_[1274]_  | ~\new_[1545]_ ;
  assign \new_[1181]_  = \new_[8981]_  ? \new_[8425]_  : \new_[8982]_ ;
  assign \new_[1182]_  = ~\new_[1272]_  | ~\new_[8428]_ ;
  assign \new_[1183]_  = ~\new_[1274]_  | ~\new_[1232]_ ;
  assign \new_[1184]_  = ~\new_[1272]_  | ~\new_[8425]_ ;
  assign \new_[1185]_  = ~n990 | ~\new_[4619]_ ;
  assign \new_[1186]_  = \\sub1_data_reg_reg[61] ;
  assign \new_[1187]_  = \\sub1_data_reg_reg[62] ;
  assign \new_[1188]_  = ~\\ks1_col_reg[21] ;
  assign \new_[1189]_  = ~\\ks1_col_reg[22] ;
  assign \new_[1190]_  = \\sub1_data_reg_reg[107] ;
  assign \new_[1191]_  = \\sub1_data_reg_reg[108] ;
  assign \new_[1192]_  = \\sub1_data_reg_reg[111] ;
  assign \new_[1193]_  = \\sub1_data_reg_reg[11] ;
  assign \new_[1194]_  = \\sub1_data_reg_reg[12] ;
  assign \new_[1195]_  = \\sub1_data_reg_reg[15] ;
  assign \new_[1196]_  = \\sub1_data_reg_reg[44] ;
  assign \new_[1197]_  = \\sub1_data_reg_reg[43] ;
  assign \new_[1198]_  = \\sub1_data_reg_reg[47] ;
  assign \new_[1199]_  = \\sub1_data_reg_reg[75] ;
  assign \new_[1200]_  = \\sub1_data_reg_reg[76] ;
  assign \new_[1201]_  = \\sub1_data_reg_reg[79] ;
  assign \new_[1202]_  = \\sub1_data_reg_reg[103] ;
  assign \new_[1203]_  = \\sub1_data_reg_reg[115] ;
  assign \new_[1204]_  = \\sub1_data_reg_reg[116] ;
  assign \new_[1205]_  = \\sub1_data_reg_reg[119] ;
  assign \new_[1206]_  = \\sub1_data_reg_reg[20] ;
  assign \new_[1207]_  = \\sub1_data_reg_reg[19] ;
  assign \new_[1208]_  = \\sub1_data_reg_reg[23] ;
  assign \new_[1209]_  = \\sub1_data_reg_reg[32] ;
  assign \new_[1210]_  = \\sub1_data_reg_reg[4] ;
  assign \new_[1211]_  = \\sub1_data_reg_reg[51] ;
  assign \new_[1212]_  = \\sub1_data_reg_reg[52] ;
  assign \new_[1213]_  = \\sub1_data_reg_reg[55] ;
  assign \new_[1214]_  = \\sub1_data_reg_reg[36] ;
  assign \new_[1215]_  = \\sub1_data_reg_reg[68] ;
  assign \new_[1216]_  = \\sub1_data_reg_reg[67] ;
  assign \new_[1217]_  = \\sub1_data_reg_reg[3] ;
  assign \new_[1218]_  = \\sub1_data_reg_reg[7] ;
  assign \new_[1219]_  = \\sub1_data_reg_reg[71] ;
  assign \new_[1220]_  = \\sub1_data_reg_reg[84] ;
  assign \new_[1221]_  = \\sub1_data_reg_reg[83] ;
  assign \new_[1222]_  = \\sub1_data_reg_reg[87] ;
  assign \new_[1223]_  = \\sub1_data_reg_reg[120] ;
  assign \new_[1224]_  = \\sub1_data_reg_reg[24] ;
  assign \new_[1225]_  = \\sub1_data_reg_reg[56] ;
  assign \new_[1226]_  = \\sub1_data_reg_reg[88] ;
  assign \new_[1227]_  = \\sbox1_alph_reg[2] ;
  assign \new_[1228]_  = ~\new_[1331]_  | ~\new_[2957]_ ;
  assign n1015 = ~\new_[6925]_  | ~\new_[1332]_ ;
  assign n1010 = ~\new_[7062]_  | ~\new_[1333]_ ;
  assign \new_[1231]_  = ~\new_[1297]_ ;
  assign \new_[1232]_  = ~\new_[8425]_ ;
  assign \new_[1233]_  = ~\\ks1_col_reg[30] ;
  assign \new_[1234]_  = \\sub1_data_reg_reg[100] ;
  assign \new_[1235]_  = ~\\ks1_col_reg[6] ;
  assign \new_[1236]_  = ~\\ks1_col_reg[5] ;
  assign \new_[1237]_  = \\sub1_data_reg_reg[35] ;
  assign \new_[1238]_  = \\sub1_data_reg_reg[39] ;
  assign \new_[1239]_  = ~\\ks1_col_reg[29] ;
  assign \new_[1240]_  = \\sub1_data_reg_reg[99] ;
  assign \new_[1241]_  = \\sub1_data_reg_reg[123] ;
  assign \new_[1242]_  = \\sub1_data_reg_reg[124] ;
  assign \new_[1243]_  = \\sub1_data_reg_reg[127] ;
  assign \new_[1244]_  = \\sub1_data_reg_reg[27] ;
  assign \new_[1245]_  = \\sub1_data_reg_reg[28] ;
  assign \new_[1246]_  = \\sub1_data_reg_reg[31] ;
  assign \new_[1247]_  = \\sub1_data_reg_reg[59] ;
  assign \new_[1248]_  = \\sub1_data_reg_reg[60] ;
  assign \new_[1249]_  = \\sub1_data_reg_reg[63] ;
  assign \new_[1250]_  = \\sub1_data_reg_reg[95] ;
  assign \new_[1251]_  = \\sub1_data_reg_reg[91] ;
  assign \new_[1252]_  = \\sub1_data_reg_reg[92] ;
  assign \new_[1253]_  = ~\\ks1_col_reg[16] ;
  assign \new_[1254]_  = \\sbox1_alph_reg[0] ;
  assign \new_[1255]_  = ~\new_[6670]_  & ~\new_[1418]_ ;
  assign \new_[1256]_  = ~\new_[6513]_  & ~\new_[1422]_ ;
  assign \new_[1257]_  = ~\new_[6516]_  & ~\new_[1425]_ ;
  assign \new_[1258]_  = ~\new_[6622]_  & ~\new_[1426]_ ;
  assign \new_[1259]_  = ~\new_[6680]_  & ~\new_[1429]_ ;
  assign \new_[1260]_  = ~\new_[6679]_  & ~\new_[1430]_ ;
  assign \new_[1261]_  = ~\new_[6689]_  & ~\new_[1431]_ ;
  assign \new_[1262]_  = ~\new_[6685]_  & ~\new_[1432]_ ;
  assign \new_[1263]_  = ~\new_[6686]_  & ~\new_[1435]_ ;
  assign \new_[1264]_  = ~\new_[6447]_  & ~\new_[1436]_ ;
  assign \new_[1265]_  = ~\new_[6577]_  & ~\new_[1437]_ ;
  assign \new_[1266]_  = ~\new_[6582]_  & ~\new_[1438]_ ;
  assign \new_[1267]_  = ~\new_[6684]_  & ~\new_[1439]_ ;
  assign \new_[1268]_  = ~\new_[6688]_  & ~\new_[1440]_ ;
  assign \new_[1269]_  = ~\new_[6517]_  & ~\new_[1443]_ ;
  assign \new_[1270]_  = ~\new_[6690]_  & ~\new_[1444]_ ;
  assign n1035 = ~\new_[6472]_  | (~\new_[1496]_  & ~\new_[6825]_ );
  assign \new_[1272]_  = \new_[8983]_  ? \new_[8453]_  : \new_[8979]_ ;
  assign n1030 = ~\new_[6463]_  | (~\new_[1495]_  & ~\new_[6803]_ );
  assign \new_[1274]_  = \new_[8979]_  ? \new_[8453]_  : \new_[8983]_ ;
  assign n1040 = ~\new_[6474]_  | (~\new_[1499]_  & ~\new_[6825]_ );
  assign n1050 = ~\new_[6477]_  | (~\new_[1500]_  & ~\new_[6803]_ );
  assign n1055 = ~\new_[6462]_  | (~\new_[1507]_  & ~\new_[6809]_ );
  assign n1045 = ~\new_[6460]_  | (~\new_[1508]_  & ~\new_[6825]_ );
  assign \new_[1279]_  = ~\new_[1423]_  & (~\new_[7564]_  | ~\new_[1098]_ );
  assign \new_[1280]_  = ~n1025 | ~\new_[3077]_ ;
  assign \new_[1281]_  = ~\new_[1424]_  & (~\new_[7564]_  | ~\new_[1099]_ );
  assign \new_[1282]_  = ~\new_[1427]_  & (~\new_[7564]_  | ~\new_[1100]_ );
  assign \new_[1283]_  = ~\new_[1428]_  & (~\new_[7564]_  | ~\new_[1101]_ );
  assign \new_[1284]_  = ~\new_[1433]_  & (~\new_[7564]_  | ~\new_[1094]_ );
  assign \new_[1285]_  = ~\new_[1434]_  & (~\new_[7564]_  | ~\new_[1095]_ );
  assign \new_[1286]_  = ~\new_[1441]_  & (~\new_[7564]_  | ~\new_[1096]_ );
  assign \new_[1287]_  = ~\new_[1442]_  & (~\new_[7564]_  | ~\new_[1097]_ );
  assign n990 = ~\new_[8815]_  | ~\new_[1522]_ ;
  assign \new_[1289]_  = ~\new_[1414]_  & (~\new_[1537]_  | ~\new_[1712]_ );
  assign n1090 = ~\new_[1389]_  | (~\new_[7077]_  & ~\new_[7646]_ );
  assign n1095 = ~\new_[1390]_  | (~\new_[6911]_  & ~\new_[7646]_ );
  assign n1100 = ~\new_[1391]_  | (~\new_[6903]_  & ~\new_[7559]_ );
  assign n1120 = ~\new_[1392]_  | (~\new_[7069]_  & ~\new_[7497]_ );
  assign n1105 = ~\new_[1393]_  | (~\new_[7071]_  & ~\new_[7498]_ );
  assign n1110 = ~\new_[1394]_  | (~\new_[7076]_  & ~\new_[7559]_ );
  assign n1115 = ~\new_[1395]_  | (~\new_[1586]_  & ~\new_[7497]_ );
  assign \new_[1297]_  = \new_[1766]_  ^ \new_[1536]_ ;
  assign \new_[1298]_  = ~\new_[1357]_ ;
  assign \new_[1299]_  = ~\new_[8600]_  | ~n1065;
  assign \new_[1300]_  = ~n1060 | ~\new_[2995]_ ;
  assign n1070 = ~\new_[1408]_  | ~\new_[6510]_ ;
  assign n1075 = ~\new_[1409]_  | ~\new_[6683]_ ;
  assign n1080 = ~\new_[1410]_  | ~\new_[6512]_ ;
  assign n1085 = ~\new_[1411]_  | ~\new_[6520]_ ;
  assign \new_[1305]_  = ~\\ks1_key_reg_reg[107] ;
  assign \new_[1306]_  = ~\\ks1_key_reg_reg[108] ;
  assign \new_[1307]_  = ~\\ks1_col_reg[20] ;
  assign \new_[1308]_  = ~\\ks1_key_reg_reg[104] ;
  assign \new_[1309]_  = ~\\ks1_col_reg[23] ;
  assign \new_[1310]_  = ~\\ks1_col_reg[19] ;
  assign \new_[1311]_  = \\sub1_data_reg_reg[106] ;
  assign \new_[1312]_  = \\sub1_data_reg_reg[10] ;
  assign \new_[1313]_  = \\sub1_data_reg_reg[74] ;
  assign \new_[1314]_  = \\sub1_data_reg_reg[42] ;
  assign \new_[1315]_  = \\sub1_data_reg_reg[114] ;
  assign \new_[1316]_  = ~\\ks1_col_reg[24] ;
  assign \new_[1317]_  = ~\\ks1_col_reg[3] ;
  assign \new_[1318]_  = ~\\ks1_col_reg[4] ;
  assign \new_[1319]_  = \\sub1_data_reg_reg[18] ;
  assign \new_[1320]_  = \\sub1_data_reg_reg[2] ;
  assign \new_[1321]_  = \\sub1_data_reg_reg[50] ;
  assign \new_[1322]_  = \\sub1_data_reg_reg[66] ;
  assign \new_[1323]_  = \\sub1_data_reg_reg[82] ;
  assign \new_[1324]_  = \\sub1_data_reg_reg[98] ;
  assign n1310 = ~\new_[6471]_  | (~\new_[1582]_  & ~\new_[7427]_ );
  assign n1315 = ~\new_[6468]_  | (~\new_[1583]_  & ~\new_[7427]_ );
  assign n1320 = ~\new_[6567]_  | (~\new_[1584]_  & ~\new_[6803]_ );
  assign n1325 = ~\new_[6486]_  | (~\new_[1585]_  & ~\new_[6803]_ );
  assign n1125 = ~\new_[6469]_  | (~\new_[1555]_  & ~\new_[6803]_ );
  assign n1130 = ~\new_[6475]_  | (~\new_[1556]_  & ~\new_[6824]_ );
  assign \new_[1331]_  = ~n1025;
  assign \new_[1332]_  = ~\new_[8608]_  | ~n4105;
  assign \new_[1333]_  = ~\new_[1535]_  | ~n4105;
  assign n1205 = ~\new_[1479]_  | (~\new_[1740]_  & ~\new_[7479]_ );
  assign n1210 = ~\new_[1481]_  | (~\new_[6787]_  & ~\new_[7479]_ );
  assign n1215 = ~\new_[1482]_  | (~\new_[7081]_  & ~\new_[7479]_ );
  assign n1220 = ~\new_[1483]_  | (~\new_[6909]_  & ~\new_[7559]_ );
  assign n1230 = ~\new_[1468]_  | (~\new_[6913]_  & ~\new_[7479]_ );
  assign n1225 = ~\new_[1469]_  | (~\new_[6928]_  & ~\new_[7559]_ );
  assign n1235 = ~\new_[1470]_  | (~\new_[6937]_  & ~\new_[7559]_ );
  assign n1265 = ~\new_[1471]_  | (~\new_[1745]_  & ~\new_[7498]_ );
  assign n1280 = ~\new_[1472]_  | (~\new_[7078]_  & ~\new_[7498]_ );
  assign \new_[1343]_  = ~\\ks1_col_reg[0] ;
  assign n1245 = ~\new_[1473]_  | (~\new_[6753]_  & ~\new_[7497]_ );
  assign n1250 = ~\new_[1474]_  | (~\new_[7011]_  & ~\new_[7494]_ );
  assign n1255 = ~\new_[1475]_  | (~\new_[7080]_  & ~\new_[7494]_ );
  assign n1260 = ~\new_[1476]_  | (~\new_[6923]_  & ~\new_[7646]_ );
  assign n1275 = ~\new_[1485]_  | (~\new_[6760]_  & ~\new_[7497]_ );
  assign n1270 = ~\new_[1486]_  | (~\new_[7063]_  & ~\new_[7494]_ );
  assign n1290 = ~\new_[1487]_  | (~\new_[6905]_  & ~\new_[7494]_ );
  assign n1285 = ~\new_[1477]_  | (~\new_[7033]_  & ~\new_[7559]_ );
  assign n1300 = ~\new_[1488]_  | (~\new_[7072]_  & ~\new_[7497]_ );
  assign n1295 = ~\new_[1489]_  | (~\new_[7064]_  & ~\new_[7497]_ );
  assign n1305 = ~\new_[1490]_  | (~\new_[7073]_  & ~\new_[7494]_ );
  assign \new_[1355]_  = ~\new_[8512]_  | ~\new_[8705]_ ;
  assign \new_[1356]_  = ~\new_[8512]_  | ~\new_[8979]_ ;
  assign \new_[1357]_  = ~\new_[8512]_  | ~n1755;
  assign \new_[1358]_  = ~\new_[1512]_  | ~\new_[2842]_ ;
  assign n1145 = ~\new_[1491]_  | ~\new_[6674]_ ;
  assign n1150 = ~\new_[1492]_  | ~\new_[6612]_ ;
  assign n1155 = ~\new_[1493]_  | ~\new_[6673]_ ;
  assign n1160 = ~\new_[1494]_  | ~\new_[6604]_ ;
  assign n1135 = ~\new_[1478]_  | (~\new_[7635]_  & ~\new_[1188]_ );
  assign n1165 = ~\new_[1497]_  | ~\new_[6687]_ ;
  assign n1140 = ~\new_[1480]_  | (~\new_[7635]_  & ~\new_[1189]_ );
  assign n1170 = ~\new_[1498]_  | ~\new_[6677]_ ;
  assign n1180 = ~\new_[1501]_  | ~\new_[6682]_ ;
  assign n1175 = ~\new_[1502]_  | ~\new_[6678]_ ;
  assign n1185 = ~\new_[1503]_  | ~\new_[6669]_ ;
  assign n1190 = ~\new_[1504]_  | ~\new_[6521]_ ;
  assign n1195 = ~\new_[1505]_  | ~\new_[6519]_ ;
  assign n1200 = ~\new_[1506]_  | ~\new_[6675]_ ;
  assign n1240 = ~\new_[1484]_  | (~\new_[1688]_  & ~\new_[6825]_ );
  assign n1330 = \new_[1941]_  ^ n1600;
  assign \new_[1375]_  = ~\\ks1_col_reg[28] ;
  assign n1440 = \new_[1593]_  ^ n1670;
  assign \new_[1377]_  = \new_[1932]_  ^ \new_[1593]_ ;
  assign \new_[1378]_  = ~\\ks1_key_reg_reg[111] ;
  assign \new_[1379]_  = ~\\ks1_col_reg[27] ;
  assign \new_[1380]_  = ~\\ks1_col_reg[31] ;
  assign \new_[1381]_  = \\sub1_data_reg_reg[34] ;
  assign \new_[1382]_  = ~\\ks1_col_reg[7] ;
  assign \new_[1383]_  = \\sub1_data_reg_reg[122] ;
  assign \new_[1384]_  = \\sub1_data_reg_reg[26] ;
  assign \new_[1385]_  = \\sub1_data_reg_reg[58] ;
  assign \new_[1386]_  = \\sub1_data_reg_reg[90] ;
  assign \new_[1387]_  = \\sbox1_ah_reg_reg[2] ;
  assign \new_[1388]_  = \\sbox1_alph_reg[1] ;
  assign \new_[1389]_  = ~\new_[1561]_  & (~\new_[7116]_  | ~\new_[8026]_ );
  assign \new_[1390]_  = ~\new_[1563]_  & (~\new_[6832]_  | ~\new_[1147]_ );
  assign \new_[1391]_  = ~\new_[1564]_  & (~\new_[6832]_  | ~\new_[1148]_ );
  assign \new_[1392]_  = ~\new_[1566]_  & (~\new_[7114]_  | ~\new_[1152]_ );
  assign \new_[1393]_  = ~\new_[1567]_  & (~\new_[6832]_  | ~\new_[1149]_ );
  assign \new_[1394]_  = ~\new_[1569]_  & (~\new_[6832]_  | ~\new_[1150]_ );
  assign \new_[1395]_  = ~\new_[1571]_  & (~\new_[7114]_  | ~\new_[1151]_ );
  assign n1375 = ~\new_[6464]_  | (~\new_[1693]_  & ~\new_[6825]_ );
  assign n1380 = ~\new_[6563]_  | (~\new_[1694]_  & ~\new_[6825]_ );
  assign n1385 = ~\new_[6564]_  | (~\new_[1695]_  & ~\new_[7427]_ );
  assign n1390 = ~\new_[6482]_  | (~\new_[1696]_  & ~\new_[7427]_ );
  assign n1395 = ~\new_[6478]_  | (~\new_[1697]_  & ~\new_[6825]_ );
  assign n1400 = ~\new_[6476]_  | (~\new_[1698]_  & ~\new_[6803]_ );
  assign n1405 = ~\new_[6481]_  | (~\new_[1699]_  & ~\new_[6824]_ );
  assign n1410 = ~\new_[6484]_  | (~\new_[1700]_  & ~\new_[6824]_ );
  assign n1415 = ~\new_[6479]_  | (~\new_[1701]_  & ~\new_[6809]_ );
  assign n1425 = ~\new_[6467]_  | (~\new_[1702]_  & ~\new_[6809]_ );
  assign n1430 = ~\new_[6483]_  | (~\new_[1703]_  & ~\new_[6825]_ );
  assign n1420 = ~\new_[6461]_  | (~\new_[1704]_  & ~\new_[6825]_ );
  assign \new_[1408]_  = ~\new_[1562]_  & (~\new_[7564]_  | ~\new_[1143]_ );
  assign \new_[1409]_  = ~\new_[1565]_  & (~\new_[7270]_  | ~\new_[1142]_ );
  assign \new_[1410]_  = ~\new_[1568]_  & (~\new_[7270]_  | ~\new_[1145]_ );
  assign \new_[1411]_  = ~\new_[1570]_  & (~\new_[7270]_  | ~\new_[1144]_ );
  assign n1025 = ~\new_[8609]_  | ~\new_[1692]_ ;
  assign n1060 = ~\new_[1512]_ ;
  assign \new_[1414]_  = ~\new_[1537]_  & ~\new_[1712]_ ;
  assign n1435 = ~\new_[1577]_  | (~\new_[7635]_  & ~\new_[1253]_ );
  assign \new_[1416]_  = ~\new_[1560]_  | ~\new_[7564]_ ;
  assign \new_[1417]_  = ~\new_[1559]_  | ~\new_[7564]_ ;
  assign \new_[1418]_  = ~\new_[6824]_  & (~\new_[6166]_  | ~\new_[1605]_ );
  assign \new_[1419]_  = ~\new_[1553]_  | ~\new_[7564]_ ;
  assign \new_[1420]_  = ~\new_[1588]_  | ~\new_[1713]_ ;
  assign \new_[1421]_  = ~\new_[1554]_  | ~\new_[7564]_ ;
  assign \new_[1422]_  = ~\new_[6824]_  & (~\new_[6167]_  | ~\new_[1606]_ );
  assign \new_[1423]_  = ~\new_[6954]_  & (~\new_[6002]_  | ~\new_[1610]_ );
  assign \new_[1424]_  = ~\new_[6954]_  & (~\new_[6004]_  | ~\new_[1611]_ );
  assign \new_[1425]_  = ~\new_[6954]_  & (~\new_[6006]_  | ~\new_[1616]_ );
  assign \new_[1426]_  = ~\new_[6954]_  & (~\new_[6007]_  | ~\new_[1617]_ );
  assign \new_[1427]_  = ~\new_[6954]_  & (~\new_[5957]_  | ~\new_[1623]_ );
  assign \new_[1428]_  = ~\new_[6954]_  & (~\new_[5958]_  | ~\new_[1624]_ );
  assign \new_[1429]_  = ~\new_[6954]_  & (~\new_[6090]_  | ~\new_[1661]_ );
  assign \new_[1430]_  = ~\new_[6954]_  & (~\new_[6091]_  | ~\new_[1662]_ );
  assign \new_[1431]_  = ~\new_[6954]_  & (~\new_[6003]_  | ~\new_[1663]_ );
  assign \new_[1432]_  = ~\new_[6954]_  & (~\new_[6029]_  | ~\new_[1664]_ );
  assign \new_[1433]_  = ~\new_[6954]_  & (~\new_[6010]_  | ~\new_[1635]_ );
  assign \new_[1434]_  = ~\new_[6954]_  & (~\new_[6008]_  | ~\new_[1636]_ );
  assign \new_[1435]_  = ~\new_[6824]_  & (~\new_[6022]_  | ~\new_[1666]_ );
  assign \new_[1436]_  = ~\new_[6824]_  & (~\new_[6016]_  | ~\new_[1667]_ );
  assign \new_[1437]_  = ~\new_[6824]_  & (~\new_[6023]_  | ~\new_[1668]_ );
  assign \new_[1438]_  = ~\new_[6824]_  & (~\new_[6001]_  | ~\new_[1644]_ );
  assign \new_[1439]_  = ~\new_[6824]_  & (~\new_[6025]_  | ~\new_[1669]_ );
  assign \new_[1440]_  = ~\new_[6824]_  & (~\new_[6026]_  | ~\new_[1645]_ );
  assign \new_[1441]_  = ~\new_[6954]_  & (~\new_[6005]_  | ~\new_[1649]_ );
  assign \new_[1442]_  = ~\new_[6954]_  & (~\new_[6028]_  | ~\new_[1650]_ );
  assign \new_[1443]_  = ~\new_[6954]_  & (~\new_[6024]_  | ~\new_[1655]_ );
  assign \new_[1444]_  = ~\new_[6954]_  & (~\new_[6020]_  | ~\new_[1657]_ );
  assign n1335 = ~\new_[1546]_  | (~\new_[7614]_  & ~\new_[1233]_ );
  assign n1345 = ~\new_[1549]_  | (~\new_[7635]_  & ~\new_[1235]_ );
  assign n1365 = ~\new_[1544]_  | (~\new_[7614]_  & ~\new_[1239]_ );
  assign n1350 = ~\new_[1548]_  | (~\new_[7635]_  & ~\new_[1236]_ );
  assign n1355 = ~\new_[1550]_  | (~\new_[1731]_  & ~\new_[6809]_ );
  assign n1360 = ~\new_[1551]_  | (~\new_[1732]_  & ~\new_[6809]_ );
  assign n1340 = ~\new_[1543]_  | (~\new_[1739]_  & ~\new_[6809]_ );
  assign n1370 = ~\new_[1552]_  | (~\new_[1741]_  & ~\new_[6809]_ );
  assign \new_[1453]_  = \new_[1903]_  ^ \new_[1706]_ ;
  assign \new_[1454]_  = ~\new_[8702]_ ;
  assign \new_[1455]_  = \\ks1_key_reg_reg[110] ;
  assign \new_[1456]_  = \\ks1_key_reg_reg[109] ;
  assign \new_[1457]_  = \\sub1_data_reg_reg[105] ;
  assign \new_[1458]_  = \\sub1_data_reg_reg[41] ;
  assign \new_[1459]_  = \\sub1_data_reg_reg[73] ;
  assign \new_[1460]_  = \\sub1_data_reg_reg[9] ;
  assign \new_[1461]_  = \\sub1_data_reg_reg[17] ;
  assign \new_[1462]_  = ~\\sub1_data_reg_reg[1] ;
  assign \new_[1463]_  = \\sub1_data_reg_reg[65] ;
  assign \new_[1464]_  = \\sub1_data_reg_reg[97] ;
  assign \new_[1465]_  = ~\\ks1_key_reg_reg[105] ;
  assign \new_[1466]_  = ~\\ks1_col_reg[18] ;
  assign \new_[1467]_  = \\sbox1_ah_reg_reg[0] ;
  assign \new_[1468]_  = ~\new_[1626]_  & (~\new_[6832]_  | ~\new_[1207]_ );
  assign \new_[1469]_  = ~\new_[1627]_  & (~\new_[7114]_  | ~\new_[1206]_ );
  assign \new_[1470]_  = ~\new_[1628]_  & (~\new_[7116]_  | ~\new_[1208]_ );
  assign \new_[1471]_  = ~\new_[1631]_  & (~\new_[7114]_  | ~\new_[1214]_ );
  assign \new_[1472]_  = ~\new_[1632]_  & (~\new_[7116]_  | ~\new_[1217]_ );
  assign \new_[1473]_  = ~\new_[1638]_  & (~\new_[7116]_  | ~\new_[1210]_ );
  assign \new_[1474]_  = ~\new_[1639]_  & (~\new_[6832]_  | ~\new_[1211]_ );
  assign \new_[1475]_  = ~\new_[1640]_  & (~\new_[6832]_  | ~\new_[1212]_ );
  assign \new_[1476]_  = ~\new_[1641]_  & (~\new_[6832]_  | ~\new_[1213]_ );
  assign \new_[1477]_  = ~\new_[1652]_  & (~\new_[7116]_  | ~\new_[1218]_ );
  assign \new_[1478]_  = ~\new_[1604]_  & (~\new_[6957]_  | ~\new_[7955]_ );
  assign \new_[1479]_  = ~\new_[1607]_  & (~\new_[6832]_  | ~\new_[1202]_ );
  assign \new_[1480]_  = ~\new_[1613]_  & (~\new_[6957]_  | ~\new_[7947]_ );
  assign \new_[1481]_  = ~\new_[1614]_  & (~\new_[6832]_  | ~\new_[1203]_ );
  assign \new_[1482]_  = ~\new_[1615]_  & (~\new_[6832]_  | ~\new_[1204]_ );
  assign \new_[1483]_  = ~\new_[1618]_  & (~\new_[6832]_  | ~\new_[1205]_ );
  assign \new_[1484]_  = (~\new_[1744]_  | ~\new_[7606]_ ) & (~\new_[7114]_  | ~\new_[1209]_ );
  assign \new_[1485]_  = ~\new_[1642]_  & (~\new_[6832]_  | ~\new_[1216]_ );
  assign \new_[1486]_  = ~\new_[1643]_  & (~\new_[7114]_  | ~\new_[1215]_ );
  assign \new_[1487]_  = ~\new_[1646]_  & (~\new_[6832]_  | ~\new_[1219]_ );
  assign \new_[1488]_  = ~\new_[1653]_  & (~\new_[6832]_  | ~\new_[1221]_ );
  assign \new_[1489]_  = ~\new_[1654]_  & (~\new_[6832]_  | ~\new_[1220]_ );
  assign \new_[1490]_  = ~\new_[1656]_  & (~\new_[6832]_  | ~\new_[1222]_ );
  assign \new_[1491]_  = ~\new_[1608]_  & (~\new_[7270]_  | ~\new_[1197]_ );
  assign \new_[1492]_  = ~\new_[1609]_  & (~\new_[7270]_  | ~\new_[1196]_ );
  assign \new_[1493]_  = ~\new_[1612]_  & (~\new_[7270]_  | ~\new_[1198]_ );
  assign \new_[1494]_  = ~\new_[1619]_  & (~\new_[7564]_  | ~\new_[1199]_ );
  assign \new_[1495]_  = ~\new_[1620]_  & (~\new_[1134]_  | ~\new_[6363]_ );
  assign \new_[1496]_  = ~\new_[1621]_  & (~\new_[1135]_  | ~\new_[6363]_ );
  assign \new_[1497]_  = ~\new_[1622]_  & (~\new_[7270]_  | ~\new_[1200]_ );
  assign \new_[1498]_  = ~\new_[1625]_  & (~\new_[7270]_  | ~\new_[1201]_ );
  assign \new_[1499]_  = ~\new_[1629]_  & (~\new_[1136]_  | ~\new_[6357]_ );
  assign \new_[1500]_  = ~\new_[1630]_  & (~\new_[1138]_  | ~\new_[6357]_ );
  assign \new_[1501]_  = ~\new_[1633]_  & (~\new_[7564]_  | ~\new_[1190]_ );
  assign \new_[1502]_  = ~\new_[1634]_  & (~\new_[7270]_  | ~\new_[1191]_ );
  assign \new_[1503]_  = ~\new_[1637]_  & (~\new_[7270]_  | ~\new_[1192]_ );
  assign \new_[1504]_  = ~\new_[1647]_  & (~\new_[7270]_  | ~\new_[1193]_ );
  assign \new_[1505]_  = ~\new_[1648]_  & (~\new_[7564]_  | ~\new_[1194]_ );
  assign \new_[1506]_  = ~\new_[1651]_  & (~\new_[7564]_  | ~\new_[1195]_ );
  assign \new_[1507]_  = ~\new_[1658]_  & (~\new_[1139]_  | ~\new_[6358]_ );
  assign \new_[1508]_  = ~\new_[1659]_  & (~\new_[1137]_  | ~\new_[6358]_ );
  assign n1450 = \new_[8004]_  ? \new_[7470]_  : \new_[8271]_ ;
  assign n1445 = \new_[7971]_  ? \new_[7597]_  : \new_[8287]_ ;
  assign n1460 = \new_[7949]_  ? \new_[7597]_  : \new_[1743]_ ;
  assign \new_[1512]_  = \new_[3075]_  ? \new_[1743]_  : \new_[2954]_ ;
  assign n1495 = ~\new_[1678]_  | (~\new_[6766]_  & ~\new_[7494]_ );
  assign n1515 = ~\new_[1672]_  | (~\new_[6807]_  & ~\new_[7494]_ );
  assign n1520 = ~\new_[1673]_  | (~\new_[7070]_  & ~\new_[7479]_ );
  assign n1525 = ~\new_[1674]_  | (~\new_[6918]_  & ~\new_[7497]_ );
  assign n1530 = ~\new_[1681]_  | (~\new_[6904]_  & ~\new_[7559]_ );
  assign n1535 = ~\new_[1682]_  | (~\new_[6926]_  & ~\new_[7498]_ );
  assign n1540 = ~\new_[1683]_  | (~\new_[1845]_  & ~\new_[7498]_ );
  assign \new_[1520]_  = \\sub1_data_reg_reg[81] ;
  assign \new_[1521]_  = \\sub1_data_reg_reg[49] ;
  assign \new_[1522]_  = ~\new_[8819]_  | ~\new_[8748]_ ;
  assign n1475 = ~\new_[1686]_  | ~\new_[6617]_ ;
  assign n1545 = ~\new_[1675]_  | (~\new_[7635]_  & ~\new_[1343]_ );
  assign n1470 = ~\new_[1676]_  | (~\new_[7635]_  & ~\new_[1310]_ );
  assign n1455 = ~\new_[1677]_  | (~\new_[7635]_  & ~\new_[1307]_ );
  assign n1480 = ~\new_[1687]_  | ~\new_[6672]_ ;
  assign n1465 = ~\new_[1679]_  | (~\new_[7635]_  & ~\new_[1309]_ );
  assign n1500 = ~\new_[1680]_  | (~\new_[7614]_  & ~\new_[1316]_ );
  assign \new_[1530]_  = \\sub1_data_reg_reg[113] ;
  assign n1505 = ~\new_[1684]_  | (~\new_[7635]_  & ~\new_[1317]_ );
  assign n1510 = ~\new_[1685]_  | (~\new_[7635]_  & ~\new_[1318]_ );
  assign n1490 = ~\new_[1689]_  | ~\new_[6681]_ ;
  assign n1485 = ~\new_[1690]_  | ~\new_[6518]_ ;
  assign \new_[1535]_  = ~\new_[8823]_ ;
  assign \new_[1536]_  = ~\new_[8981]_  | ~\new_[1923]_ ;
  assign \new_[1537]_  = ~\new_[1710]_  & ~\new_[1767]_ ;
  assign \new_[1538]_  = \\sub1_data_reg_reg[33] ;
  assign \new_[1539]_  = ~\\sub1_data_reg_reg[57] ;
  assign \new_[1540]_  = ~\\sub1_data_reg_reg[89] ;
  assign \new_[1541]_  = ~\\sub1_data_reg_reg[25] ;
  assign \new_[1542]_  = ~\\ks1_col_reg[26] ;
  assign \new_[1543]_  = (~\new_[1780]_  | ~\new_[7606]_ ) & (~\new_[7116]_  | ~\new_[1234]_ );
  assign \new_[1544]_  = (~\new_[6957]_  | ~\new_[8120]_ ) & (~\new_[8162]_  | ~\new_[7821]_ );
  assign \new_[1545]_  = ~\new_[8428]_ ;
  assign \new_[1546]_  = (~\new_[6957]_  | ~\new_[8027]_ ) & (~\new_[8172]_  | ~\new_[7821]_ );
  assign n1605 = \new_[8707]_  ^ n1730;
  assign \new_[1548]_  = (~\new_[6955]_  | ~\new_[8095]_ ) & (~\new_[8162]_  | ~\new_[7631]_ );
  assign \new_[1549]_  = (~\new_[6955]_  | ~\new_[8134]_ ) & (~\new_[8172]_  | ~\new_[7631]_ );
  assign \new_[1550]_  = (~\new_[1806]_  | ~\new_[7606]_ ) & (~\new_[7116]_  | ~\new_[1237]_ );
  assign \new_[1551]_  = (~\new_[1807]_  | ~\new_[7606]_ ) & (~\new_[7114]_  | ~\new_[1238]_ );
  assign \new_[1552]_  = (~\new_[1803]_  | ~\new_[7606]_ ) & (~\new_[7114]_  | ~\new_[1240]_ );
  assign \new_[1553]_  = \new_[8162]_  ? \new_[7569]_  : \new_[1115]_ ;
  assign \new_[1554]_  = \new_[8172]_  ? \new_[7569]_  : \new_[1114]_ ;
  assign \new_[1555]_  = ~\new_[1717]_  & (~\new_[1186]_  | ~\new_[6361]_ );
  assign \new_[1556]_  = ~\new_[1718]_  & (~\new_[1187]_  | ~\new_[6361]_ );
  assign n1555 = \new_[7984]_  ? \new_[7470]_  : \new_[1805]_ ;
  assign \new_[1558]_  = ~\\sub1_data_reg_reg[121] ;
  assign \new_[1559]_  = \new_[1115]_  ? \new_[7569]_  : \new_[8162]_ ;
  assign \new_[1560]_  = \new_[1114]_  ? \new_[7569]_  : \new_[8172]_ ;
  assign \new_[1561]_  = ~\new_[6954]_  & (~\new_[6084]_  | ~\new_[1756]_ );
  assign \new_[1562]_  = ~\new_[1729]_  & ~\new_[6803]_ ;
  assign \new_[1563]_  = ~\new_[1730]_  & ~\new_[6824]_ ;
  assign \new_[1564]_  = ~\new_[6954]_  & (~\new_[6089]_  | ~\new_[1758]_ );
  assign \new_[1565]_  = ~\new_[1733]_  & ~\new_[7427]_ ;
  assign \new_[1566]_  = ~\new_[6803]_  & (~\new_[6019]_  | ~\new_[1759]_ );
  assign \new_[1567]_  = ~\new_[1734]_  & ~\new_[6703]_ ;
  assign \new_[1568]_  = ~\new_[1735]_  & ~\new_[6803]_ ;
  assign \new_[1569]_  = ~\new_[1736]_  & ~\new_[6703]_ ;
  assign \new_[1570]_  = ~\new_[1737]_  & ~\new_[6808]_ ;
  assign \new_[1571]_  = ~\new_[1738]_  & ~\new_[6703]_ ;
  assign n1560 = ~\new_[1721]_  | (~\new_[7614]_  & ~\new_[1379]_ );
  assign n1550 = ~\new_[1722]_  | (~\new_[7614]_  & ~\new_[1375]_ );
  assign n1565 = ~\new_[1723]_  | (~\new_[7614]_  & ~\new_[1380]_ );
  assign n1575 = ~\new_[1724]_  | (~\new_[7635]_  & ~\new_[1382]_ );
  assign n1570 = ~\new_[1720]_  | (~\new_[1844]_  & ~\new_[6825]_ );
  assign \new_[1577]_  = ~\new_[1746]_  & (~\new_[6957]_  | ~\new_[8056]_ );
  assign n1580 = ~\new_[6473]_  | (~\new_[1762]_  & ~\new_[6824]_ );
  assign n1585 = ~\new_[6553]_  | (~\new_[1763]_  & ~\new_[6825]_ );
  assign n1590 = ~\new_[6465]_  | (~\new_[1764]_  & ~\new_[6825]_ );
  assign n1595 = ~\new_[6466]_  | (~\new_[1765]_  & ~\new_[6809]_ );
  assign \new_[1582]_  = ~\new_[1748]_  & (~\new_[1223]_  | ~\new_[6363]_ );
  assign \new_[1583]_  = ~\new_[1749]_  & (~\new_[1224]_  | ~\new_[6357]_ );
  assign \new_[1584]_  = ~\new_[1750]_  & (~\new_[1225]_  | ~\new_[6361]_ );
  assign \new_[1585]_  = ~\new_[1707]_  & (~\new_[1226]_  | ~\new_[6358]_ );
  assign \new_[1586]_  = ~\new_[1747]_  & (~\new_[1149]_  | ~\new_[7569]_ );
  assign \new_[1587]_  = ~\new_[1716]_  | ~\new_[2996]_ ;
  assign \new_[1588]_  = ~\new_[8516]_ ;
  assign n1665 = ~\new_[1760]_  | (~\new_[7635]_  & ~\new_[1466]_ );
  assign \new_[1590]_  = ~\\ks1_key_reg_reg[106] ;
  assign \new_[1591]_  = ~\\ks1_col_reg[2] ;
  assign \new_[1592]_  = \\sbox1_ah_reg_reg[1] ;
  assign \new_[1593]_  = ~\new_[1710]_ ;
  assign \new_[1594]_  = ~\new_[1711]_ ;
  assign \new_[1595]_  = ~\new_[1713]_ ;
  assign \new_[1596]_  = ~\\ks1_col_reg[17] ;
  assign n1685 = ~\new_[1769]_  | (~\new_[6907]_  & ~\new_[7497]_ );
  assign n1640 = ~\new_[1770]_  | (~\new_[6805]_  & ~\new_[7494]_ );
  assign n1645 = ~\new_[1771]_  | (~\new_[6939]_  & ~\new_[7479]_ );
  assign n1680 = ~\new_[1772]_  | (~\new_[7068]_  & ~\new_[7479]_ );
  assign n1650 = ~\new_[1773]_  | (~\new_[6906]_  & ~\new_[7479]_ );
  assign n1675 = ~\new_[1774]_  | (~\new_[7082]_  & ~\new_[7559]_ );
  assign n1655 = ~\new_[1775]_  | (~\new_[1895]_  & ~\new_[7646]_ );
  assign \new_[1604]_  = ~\new_[8161]_  & ~\new_[7826]_ ;
  assign \new_[1605]_  = ~\new_[8162]_  | ~\new_[6394]_ ;
  assign \new_[1606]_  = ~\new_[8172]_  | ~\new_[6394]_ ;
  assign \new_[1607]_  = ~\new_[1781]_  & ~\new_[6703]_ ;
  assign \new_[1608]_  = ~\new_[1782]_  & ~\new_[6808]_ ;
  assign \new_[1609]_  = ~\new_[1783]_  & ~\new_[6808]_ ;
  assign \new_[1610]_  = ~\new_[8162]_  | ~\new_[6360]_ ;
  assign \new_[1611]_  = ~\new_[8172]_  | ~\new_[6360]_ ;
  assign \new_[1612]_  = ~\new_[1784]_  & ~\new_[6803]_ ;
  assign \new_[1613]_  = ~\new_[8171]_  & ~\new_[7826]_ ;
  assign \new_[1614]_  = ~\new_[1785]_  & ~\new_[6703]_ ;
  assign \new_[1615]_  = ~\new_[1786]_  & ~\new_[6808]_ ;
  assign \new_[1616]_  = ~\new_[8162]_  | ~\new_[6368]_ ;
  assign \new_[1617]_  = ~\new_[8172]_  | ~\new_[6368]_ ;
  assign \new_[1618]_  = ~\new_[1787]_  & ~\new_[6703]_ ;
  assign \new_[1619]_  = ~\new_[1788]_  & ~\new_[6703]_ ;
  assign \new_[1620]_  = ~\new_[8161]_  & ~\new_[6363]_ ;
  assign \new_[1621]_  = ~\new_[8171]_  & ~\new_[6363]_ ;
  assign \new_[1622]_  = ~\new_[1789]_  & ~\new_[6808]_ ;
  assign \new_[1623]_  = ~\new_[8162]_  | ~\new_[6356]_ ;
  assign \new_[1624]_  = ~\new_[8172]_  | ~\new_[6356]_ ;
  assign \new_[1625]_  = ~\new_[1790]_  & ~\new_[6808]_ ;
  assign \new_[1626]_  = ~\new_[6954]_  & (~\new_[6085]_  | ~\new_[1832]_ );
  assign \new_[1627]_  = ~\new_[6954]_  & (~\new_[6088]_  | ~\new_[1833]_ );
  assign \new_[1628]_  = ~\new_[6954]_  & (~\new_[6074]_  | ~\new_[1834]_ );
  assign \new_[1629]_  = ~\new_[8161]_  & ~\new_[6357]_ ;
  assign \new_[1630]_  = ~\new_[8171]_  & ~\new_[6357]_ ;
  assign \new_[1631]_  = ~\new_[6954]_  & (~\new_[6017]_  | ~\new_[1835]_ );
  assign \new_[1632]_  = ~\new_[6803]_  & (~\new_[6027]_  | ~\new_[1840]_ );
  assign \new_[1633]_  = ~\new_[1791]_  & ~\new_[6703]_ ;
  assign \new_[1634]_  = ~\new_[1792]_  & ~\new_[7427]_ ;
  assign \new_[1635]_  = ~\new_[8162]_  | ~\new_[6365]_ ;
  assign \new_[1636]_  = ~\new_[8172]_  | ~\new_[6365]_ ;
  assign \new_[1637]_  = ~\new_[1793]_  & ~\new_[6703]_ ;
  assign \new_[1638]_  = ~\new_[6954]_  & (~\new_[6018]_  | ~\new_[1841]_ );
  assign \new_[1639]_  = ~\new_[6954]_  & (~\new_[5999]_  | ~\new_[1836]_ );
  assign \new_[1640]_  = ~\new_[6954]_  & (~\new_[6021]_  | ~\new_[1837]_ );
  assign \new_[1641]_  = ~\new_[6803]_  & (~\new_[6009]_  | ~\new_[1838]_ );
  assign \new_[1642]_  = ~\new_[1794]_  & ~\new_[6703]_ ;
  assign \new_[1643]_  = ~\new_[1795]_  & ~\new_[6703]_ ;
  assign \new_[1644]_  = ~\new_[8162]_  | ~\new_[6362]_ ;
  assign \new_[1645]_  = ~\new_[8172]_  | ~\new_[6362]_ ;
  assign \new_[1646]_  = ~\new_[1796]_  & ~\new_[6703]_ ;
  assign \new_[1647]_  = ~\new_[1797]_  & ~\new_[6808]_ ;
  assign \new_[1648]_  = ~\new_[1798]_  & ~\new_[7427]_ ;
  assign \new_[1649]_  = ~\new_[8162]_  | ~\new_[6359]_ ;
  assign \new_[1650]_  = ~\new_[8172]_  | ~\new_[6359]_ ;
  assign \new_[1651]_  = ~\new_[1799]_  & ~\new_[6703]_ ;
  assign \new_[1652]_  = ~\new_[6803]_  & (~\new_[6015]_  | ~\new_[1839]_ );
  assign \new_[1653]_  = ~\new_[1800]_  & ~\new_[6703]_ ;
  assign \new_[1654]_  = ~\new_[1801]_  & ~\new_[6824]_ ;
  assign \new_[1655]_  = ~\new_[8162]_  | ~\new_[6366]_ ;
  assign \new_[1656]_  = ~\new_[1802]_  & ~\new_[6824]_ ;
  assign \new_[1657]_  = ~\new_[8172]_  | ~\new_[6366]_ ;
  assign \new_[1658]_  = ~\new_[8161]_  & ~\new_[6358]_ ;
  assign \new_[1659]_  = ~\new_[8171]_  & ~\new_[6358]_ ;
  assign n1620 = ~\new_[1776]_  | ~\new_[6671]_ ;
  assign \new_[1661]_  = ~\new_[8162]_  | ~\new_[6172]_ ;
  assign \new_[1662]_  = ~\new_[8172]_  | ~\new_[6172]_ ;
  assign \new_[1663]_  = ~\new_[8162]_  | ~\new_[6367]_ ;
  assign \new_[1664]_  = ~\new_[8172]_  | ~\new_[6367]_ ;
  assign n1625 = ~\new_[1777]_  | ~\new_[6676]_ ;
  assign \new_[1666]_  = ~\new_[8162]_  | ~\new_[6354]_ ;
  assign \new_[1667]_  = ~\new_[8172]_  | ~\new_[6354]_ ;
  assign \new_[1668]_  = ~\new_[8162]_  | ~\new_[6355]_ ;
  assign \new_[1669]_  = ~\new_[8172]_  | ~\new_[6355]_ ;
  assign n1630 = ~\new_[1778]_  | ~\new_[6514]_ ;
  assign n1635 = ~\new_[1779]_  | ~\new_[6515]_ ;
  assign \new_[1672]_  = ~\new_[1818]_  & (~\new_[7114]_  | ~\new_[1319]_ );
  assign \new_[1673]_  = ~\new_[1821]_  & (~\new_[7116]_  | ~\new_[1320]_ );
  assign \new_[1674]_  = ~\new_[1824]_  & (~\new_[7114]_  | ~\new_[1321]_ );
  assign \new_[1675]_  = (~\new_[6955]_  | ~\new_[7954]_ ) & (~\new_[8170]_  | ~\new_[7631]_ );
  assign \new_[1676]_  = ~\new_[1808]_  & (~\new_[6957]_  | ~\new_[8140]_ );
  assign \new_[1677]_  = ~\new_[1809]_  & (~\new_[6957]_  | ~\new_[8038]_ );
  assign \new_[1678]_  = ~\new_[1814]_  & (~\new_[6832]_  | ~\new_[1315]_ );
  assign \new_[1679]_  = ~\new_[1810]_  & (~\new_[6957]_  | ~\new_[7997]_ );
  assign \new_[1680]_  = (~\new_[6957]_  | ~\new_[8041]_ ) & (~\new_[8170]_  | ~\new_[7821]_ );
  assign \new_[1681]_  = ~\new_[1828]_  & (~\new_[6832]_  | ~\new_[1322]_ );
  assign \new_[1682]_  = ~\new_[1830]_  & (~\new_[6832]_  | ~\new_[1323]_ );
  assign \new_[1683]_  = ~\new_[1754]_  & (~\new_[7116]_  | ~\new_[1324]_ );
  assign \new_[1684]_  = (~\new_[6955]_  | ~\new_[8012]_ ) & (~\new_[8984]_  | ~\new_[7631]_ );
  assign \new_[1685]_  = (~\new_[6955]_  | ~\new_[8079]_ ) & (~\new_[1896]_  | ~\new_[7631]_ );
  assign \new_[1686]_  = ~\new_[1812]_  & (~\new_[7564]_  | ~\new_[1314]_ );
  assign \new_[1687]_  = ~\new_[1813]_  & (~\new_[7270]_  | ~\new_[1313]_ );
  assign \new_[1688]_  = ~\new_[6014]_  & (~\new_[8170]_  | ~\new_[6367]_ );
  assign \new_[1689]_  = ~\new_[1823]_  & (~\new_[7564]_  | ~\new_[1311]_ );
  assign \new_[1690]_  = ~\new_[1829]_  & (~\new_[7270]_  | ~\new_[1312]_ );
  assign \new_[1691]_  = ~n1615 | ~\new_[3099]_ ;
  assign \new_[1692]_  = ~n1610 | ~\new_[8615]_ ;
  assign \new_[1693]_  = ~\new_[1815]_  & (~\new_[1241]_  | ~\new_[6363]_ );
  assign \new_[1694]_  = ~\new_[1816]_  & (~\new_[1242]_  | ~\new_[6363]_ );
  assign \new_[1695]_  = ~\new_[1817]_  & (~\new_[6363]_  | ~\new_[1243]_ );
  assign \new_[1696]_  = ~\new_[1819]_  & (~\new_[1244]_  | ~\new_[6357]_ );
  assign \new_[1697]_  = ~\new_[1820]_  & (~\new_[1245]_  | ~\new_[6357]_ );
  assign \new_[1698]_  = ~\new_[1822]_  & (~\new_[6357]_  | ~\new_[1246]_ );
  assign \new_[1699]_  = ~\new_[1825]_  & (~\new_[1247]_  | ~\new_[6361]_ );
  assign \new_[1700]_  = ~\new_[1826]_  & (~\new_[1248]_  | ~\new_[6361]_ );
  assign \new_[1701]_  = ~\new_[1827]_  & (~\new_[6361]_  | ~\new_[1249]_ );
  assign \new_[1702]_  = ~\new_[1751]_  & (~\new_[1251]_  | ~\new_[6358]_ );
  assign \new_[1703]_  = ~\new_[1752]_  & (~\new_[1252]_  | ~\new_[6358]_ );
  assign \new_[1704]_  = ~\new_[1753]_  & (~\new_[6358]_  | ~\new_[1250]_ );
  assign n1660 = \new_[7986]_  ? \new_[7470]_  : \new_[1899]_ ;
  assign \new_[1706]_  = ~\new_[8979]_  | ~\new_[1932]_ ;
  assign \new_[1707]_  = ~\new_[8169]_  & ~\new_[6358]_ ;
  assign n1710 = ~\new_[1843]_  | (~\new_[7614]_  & ~\new_[1542]_ );
  assign \new_[1709]_  = \\sbox1_alph_reg[3] ;
  assign \new_[1710]_  = ~\new_[8515]_ ;
  assign \new_[1711]_  = ~\new_[1848]_  | ~\new_[8707]_ ;
  assign \new_[1712]_  = ~\new_[8705]_  | ~\new_[1945]_ ;
  assign \new_[1713]_  = ~\new_[8705]_  | ~\new_[1941]_ ;
  assign n1670 = ~\new_[1767]_ ;
  assign \new_[1715]_  = ~\\ks1_col_reg[25] ;
  assign \new_[1716]_  = ~\new_[9013]_ ;
  assign \new_[1717]_  = ~\new_[8161]_  & ~\new_[6361]_ ;
  assign \new_[1718]_  = ~\new_[8171]_  & ~\new_[6361]_ ;
  assign n1690 = ~\new_[1849]_  | (~\new_[1894]_  & ~\new_[6825]_ );
  assign \new_[1720]_  = (~\new_[1874]_  | ~\new_[7606]_ ) & (~\new_[7116]_  | ~\new_[1381]_ );
  assign \new_[1721]_  = (~\new_[6957]_  | ~\new_[7959]_ ) & (~\new_[8984]_  | ~\new_[7821]_ );
  assign \new_[1722]_  = (~\new_[6957]_  | ~\new_[8096]_ ) & (~\new_[1896]_  | ~\new_[7821]_ );
  assign \new_[1723]_  = (~\new_[6957]_  | ~\new_[8050]_ ) & (~\new_[1898]_  | ~\new_[7821]_ );
  assign \new_[1724]_  = (~\new_[6955]_  | ~\new_[8045]_ ) & (~\new_[1898]_  | ~\new_[7631]_ );
  assign n1715 = ~\new_[6431]_  | (~\new_[1859]_  & ~\new_[6825]_ );
  assign n1705 = ~\new_[6470]_  | (~\new_[1860]_  & ~\new_[6825]_ );
  assign n1695 = ~\new_[6480]_  | (~\new_[1861]_  & ~\new_[6825]_ );
  assign n1700 = ~\new_[6485]_  | (~\new_[1862]_  & ~\new_[6803]_ );
  assign \new_[1729]_  = (~\new_[8170]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1142]_ );
  assign \new_[1730]_  = (~\new_[8170]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1147]_ );
  assign \new_[1731]_  = (~\new_[8984]_  | ~\new_[6367]_ ) & (~\new_[6173]_  | ~\new_[1237]_ );
  assign \new_[1732]_  = (~\new_[1898]_  | ~\new_[6367]_ ) & (~\new_[6173]_  | ~\new_[1238]_ );
  assign \new_[1733]_  = (~\new_[8170]_  | ~\new_[6365]_ ) & (~\new_[1143]_  | ~\new_[6436]_ );
  assign \new_[1734]_  = (~\new_[8170]_  | ~\new_[6362]_ ) & (~\new_[6417]_  | ~\new_[1149]_ );
  assign \new_[1735]_  = (~\new_[8170]_  | ~\new_[6359]_ ) & (~\new_[6170]_  | ~\new_[1144]_ );
  assign \new_[1736]_  = (~\new_[8170]_  | ~\new_[6366]_ ) & (~\new_[1150]_  | ~\new_[6435]_ );
  assign \new_[1737]_  = (~\new_[8170]_  | ~\new_[6356]_ ) & (~\new_[1145]_  | ~\new_[6092]_ );
  assign \new_[1738]_  = (~\new_[8170]_  | ~\new_[6394]_ ) & (~\new_[1151]_  | ~\new_[6453]_ );
  assign \new_[1739]_  = (~\new_[1896]_  | ~\new_[6394]_ ) & (~\new_[1234]_  | ~\new_[6453]_ );
  assign \new_[1740]_  = ~\new_[1850]_  & (~\new_[1219]_  | ~\new_[7632]_ );
  assign \new_[1741]_  = (~\new_[8984]_  | ~\new_[6394]_ ) & (~\new_[6453]_  | ~\new_[1240]_ );
  assign \new_[1742]_  = ~\new_[1805]_ ;
  assign \new_[1743]_  = ~\new_[1831]_  | ~\new_[1854]_ ;
  assign \new_[1744]_  = \new_[1149]_  ? \new_[7569]_  : \new_[8170]_ ;
  assign \new_[1745]_  = (~\new_[1896]_  | ~\new_[7632]_ ) & (~\new_[1215]_  | ~\new_[7738]_ );
  assign \new_[1746]_  = ~\new_[8169]_  & ~\new_[7826]_ ;
  assign \new_[1747]_  = ~\new_[8169]_  & ~\new_[7569]_ ;
  assign \new_[1748]_  = ~\new_[8169]_  & ~\new_[6363]_ ;
  assign \new_[1749]_  = ~\new_[8169]_  & ~\new_[6357]_ ;
  assign \new_[1750]_  = ~\new_[8169]_  & ~\new_[6361]_ ;
  assign \new_[1751]_  = ~\new_[8985]_  & ~\new_[6358]_ ;
  assign \new_[1752]_  = ~\new_[1872]_  & ~\new_[6358]_ ;
  assign \new_[1753]_  = ~\new_[1914]_  & ~\new_[6358]_ ;
  assign \new_[1754]_  = ~\new_[1863]_  & ~\new_[6954]_ ;
  assign n1735 = ~\new_[1857]_  | (~\new_[7635]_  & ~\new_[1596]_ );
  assign \new_[1756]_  = ~\new_[8170]_  | ~\new_[6355]_ ;
  assign n1725 = ~\new_[1858]_  | (~\new_[7635]_  & ~\new_[1591]_ );
  assign \new_[1758]_  = ~\new_[8170]_  | ~\new_[6172]_ ;
  assign \new_[1759]_  = ~\new_[8170]_  | ~\new_[6354]_ ;
  assign \new_[1760]_  = ~\new_[1875]_  & (~\new_[6957]_  | ~\new_[8083]_ );
  assign \new_[1761]_  = ~\\ks1_col_reg[1] ;
  assign \new_[1762]_  = ~\new_[1877]_  & (~\new_[1383]_  | ~\new_[6363]_ );
  assign \new_[1763]_  = ~\new_[1878]_  & (~\new_[1384]_  | ~\new_[6357]_ );
  assign \new_[1764]_  = ~\new_[1879]_  & (~\new_[1385]_  | ~\new_[6361]_ );
  assign \new_[1765]_  = ~\new_[1876]_  & (~\new_[1386]_  | ~\new_[6358]_ );
  assign \new_[1766]_  = ~\new_[1881]_  | ~n1755;
  assign \new_[1767]_  = ~\new_[1848]_ ;
  assign n1730 = \new_[8705]_ ;
  assign \new_[1769]_  = ~\new_[1884]_  & (~\new_[6832]_  | ~\new_[1530]_ );
  assign \new_[1770]_  = ~\new_[1885]_  & (~\new_[6832]_  | ~\new_[1461]_ );
  assign \new_[1771]_  = ~\new_[1886]_  & (~\new_[7116]_  | ~\new_[8068]_ );
  assign \new_[1772]_  = ~\new_[1888]_  & (~\new_[7114]_  | ~\new_[1521]_ );
  assign \new_[1773]_  = ~\new_[1889]_  & (~\new_[6832]_  | ~\new_[1463]_ );
  assign \new_[1774]_  = ~\new_[1891]_  & (~\new_[6832]_  | ~\new_[1520]_ );
  assign \new_[1775]_  = ~\new_[1852]_  & (~\new_[7116]_  | ~\new_[1464]_ );
  assign \new_[1776]_  = ~\new_[1883]_  & (~\new_[7270]_  | ~\new_[1458]_ );
  assign \new_[1777]_  = ~\new_[1887]_  & (~\new_[7270]_  | ~\new_[1457]_ );
  assign \new_[1778]_  = ~\new_[1890]_  & (~\new_[7270]_  | ~\new_[1460]_ );
  assign \new_[1779]_  = ~\new_[1853]_  & (~\new_[7564]_  | ~\new_[1459]_ );
  assign \new_[1780]_  = \new_[1896]_  ? \new_[7632]_  : \new_[1215]_ ;
  assign \new_[1781]_  = (~\new_[1898]_  | ~\new_[6394]_ ) & (~\new_[1202]_  | ~\new_[6453]_ );
  assign \new_[1782]_  = (~\new_[8984]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1190]_ );
  assign \new_[1783]_  = (~\new_[1896]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1191]_ );
  assign \new_[1784]_  = (~\new_[1898]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1192]_ );
  assign \new_[1785]_  = (~\new_[8984]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1203]_ );
  assign \new_[1786]_  = (~\new_[1896]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1204]_ );
  assign \new_[1787]_  = (~\new_[1898]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1205]_ );
  assign \new_[1788]_  = (~\new_[8984]_  | ~\new_[6356]_ ) & (~\new_[1193]_  | ~\new_[6092]_ );
  assign \new_[1789]_  = (~\new_[1896]_  | ~\new_[6356]_ ) & (~\new_[1194]_  | ~\new_[6092]_ );
  assign \new_[1790]_  = (~\new_[1898]_  | ~\new_[6356]_ ) & (~\new_[1195]_  | ~\new_[6092]_ );
  assign \new_[1791]_  = (~\new_[8984]_  | ~\new_[6365]_ ) & (~\new_[1197]_  | ~\new_[6436]_ );
  assign \new_[1792]_  = (~\new_[1896]_  | ~\new_[6365]_ ) & (~\new_[1196]_  | ~\new_[6436]_ );
  assign \new_[1793]_  = (~\new_[1898]_  | ~\new_[6365]_ ) & (~\new_[6436]_  | ~\new_[1198]_ );
  assign \new_[1794]_  = (~\new_[8984]_  | ~\new_[6362]_ ) & (~\new_[6417]_  | ~\new_[1216]_ );
  assign \new_[1795]_  = (~\new_[1896]_  | ~\new_[6362]_ ) & (~\new_[1215]_  | ~\new_[6417]_ );
  assign \new_[1796]_  = (~\new_[1898]_  | ~\new_[6362]_ ) & (~\new_[6417]_  | ~\new_[1219]_ );
  assign \new_[1797]_  = (~\new_[8984]_  | ~\new_[6359]_ ) & (~\new_[1199]_  | ~\new_[6170]_ );
  assign \new_[1798]_  = (~\new_[1896]_  | ~\new_[6359]_ ) & (~\new_[1200]_  | ~\new_[6170]_ );
  assign \new_[1799]_  = (~\new_[1898]_  | ~\new_[6359]_ ) & (~\new_[6170]_  | ~\new_[1201]_ );
  assign \new_[1800]_  = (~\new_[8984]_  | ~\new_[6366]_ ) & (~\new_[1221]_  | ~\new_[6435]_ );
  assign \new_[1801]_  = (~\new_[1896]_  | ~\new_[6366]_ ) & (~\new_[1220]_  | ~\new_[6435]_ );
  assign \new_[1802]_  = (~\new_[1898]_  | ~\new_[6366]_ ) & (~\new_[6435]_  | ~\new_[1222]_ );
  assign \new_[1803]_  = \new_[8984]_  ? \new_[7569]_  : \new_[1216]_ ;
  assign n1720 = \new_[8075]_  ? \new_[7597]_  : \new_[9004]_ ;
  assign \new_[1805]_  = ~\new_[1855]_  | ~\new_[1892]_ ;
  assign \new_[1806]_  = \new_[1216]_  ? \new_[7632]_  : \new_[8984]_ ;
  assign \new_[1807]_  = \new_[1219]_  ? \new_[7569]_  : \new_[1898]_ ;
  assign \new_[1808]_  = ~\new_[8985]_  & ~\new_[7826]_ ;
  assign \new_[1809]_  = ~\new_[1872]_  & ~\new_[7826]_ ;
  assign \new_[1810]_  = ~\new_[1914]_  & ~\new_[7826]_ ;
  assign \new_[1811]_  = ~\new_[1873]_  | ~\new_[2955]_ ;
  assign \new_[1812]_  = ~\new_[1864]_  & ~\new_[6808]_ ;
  assign \new_[1813]_  = ~\new_[1865]_  & ~\new_[6803]_ ;
  assign \new_[1814]_  = ~\new_[1867]_  & ~\new_[6808]_ ;
  assign \new_[1815]_  = ~\new_[8985]_  & ~\new_[6363]_ ;
  assign \new_[1816]_  = ~\new_[1872]_  & ~\new_[6363]_ ;
  assign \new_[1817]_  = ~\new_[1914]_  & ~\new_[6363]_ ;
  assign \new_[1818]_  = ~\new_[6954]_  & (~\new_[6083]_  | ~\new_[1900]_ );
  assign \new_[1819]_  = ~\new_[8985]_  & ~\new_[6357]_ ;
  assign \new_[1820]_  = ~\new_[1872]_  & ~\new_[6357]_ ;
  assign \new_[1821]_  = ~\new_[6954]_  & (~\new_[6013]_  | ~\new_[1901]_ );
  assign \new_[1822]_  = ~\new_[1914]_  & ~\new_[6357]_ ;
  assign \new_[1823]_  = ~\new_[1868]_  & ~\new_[7427]_ ;
  assign \new_[1824]_  = ~\new_[6803]_  & (~\new_[6012]_  | ~\new_[1902]_ );
  assign \new_[1825]_  = ~\new_[8985]_  & ~\new_[6361]_ ;
  assign \new_[1826]_  = ~\new_[1872]_  & ~\new_[6361]_ ;
  assign \new_[1827]_  = ~\new_[1914]_  & ~\new_[6361]_ ;
  assign \new_[1828]_  = ~\new_[1869]_  & ~\new_[6824]_ ;
  assign \new_[1829]_  = ~\new_[1871]_  & ~\new_[6803]_ ;
  assign \new_[1830]_  = ~\new_[1870]_  & ~\new_[6808]_ ;
  assign \new_[1831]_  = ~\new_[8209]_  | ~\new_[3355]_ ;
  assign \new_[1832]_  = ~\new_[8984]_  | ~\new_[6172]_ ;
  assign \new_[1833]_  = ~\new_[1896]_  | ~\new_[6172]_ ;
  assign \new_[1834]_  = ~\new_[1898]_  | ~\new_[6172]_ ;
  assign \new_[1835]_  = ~\new_[1896]_  | ~\new_[6367]_ ;
  assign \new_[1836]_  = ~\new_[8984]_  | ~\new_[6354]_ ;
  assign \new_[1837]_  = ~\new_[1896]_  | ~\new_[6354]_ ;
  assign \new_[1838]_  = ~\new_[1898]_  | ~\new_[6354]_ ;
  assign \new_[1839]_  = ~\new_[1898]_  | ~\new_[6355]_ ;
  assign \new_[1840]_  = ~\new_[8984]_  | ~\new_[6355]_ ;
  assign \new_[1841]_  = ~\new_[1896]_  | ~\new_[6355]_ ;
  assign n1745 = ~\new_[1893]_  | (~\new_[7614]_  & ~\new_[1715]_ );
  assign \new_[1843]_  = (~\new_[6957]_  | ~\new_[8023]_ ) & (~\new_[1929]_  | ~\new_[7821]_ );
  assign \new_[1844]_  = (~\new_[1929]_  | ~\new_[6367]_ ) & (~\new_[6173]_  | ~\new_[1381]_ );
  assign \new_[1845]_  = (~\new_[1929]_  | ~\new_[7738]_ ) & (~\new_[1322]_  | ~\new_[7569]_ );
  assign \new_[1846]_  = ~\new_[1880]_ ;
  assign n1740 = \new_[1945]_  ^ n1755;
  assign \new_[1848]_  = ~\new_[8455]_ ;
  assign \new_[1849]_  = (~\new_[1916]_  | ~\new_[7606]_ ) & (~\new_[7114]_  | ~\new_[1538]_ );
  assign \new_[1850]_  = \new_[1898]_  & \new_[7738]_ ;
  assign \new_[1851]_  = ~\new_[3076]_  | ~\new_[1899]_ ;
  assign \new_[1852]_  = ~\new_[1912]_  & ~\new_[6954]_ ;
  assign \new_[1853]_  = ~\new_[1913]_  & ~\new_[6808]_ ;
  assign \new_[1854]_  = ~\new_[8168]_  | ~\new_[3098]_ ;
  assign \new_[1855]_  = ~\new_[1915]_  | ~\new_[3536]_ ;
  assign n1750 = ~\new_[1905]_  | (~\new_[7635]_  & ~\new_[1761]_ );
  assign \new_[1857]_  = ~\new_[1918]_  & (~\new_[6957]_  | ~\new_[8029]_ );
  assign \new_[1858]_  = (~\new_[6955]_  | ~\new_[8142]_ ) & (~\new_[1929]_  | ~\new_[7631]_ );
  assign \new_[1859]_  = ~\new_[1919]_  & (~\new_[8101]_  | ~\new_[6363]_ );
  assign \new_[1860]_  = ~\new_[1920]_  & (~\new_[8053]_  | ~\new_[6357]_ );
  assign \new_[1861]_  = ~\new_[1921]_  & (~\new_[8020]_  | ~\new_[6361]_ );
  assign \new_[1862]_  = ~\new_[1917]_  & (~\new_[7939]_  | ~\new_[6358]_ );
  assign \new_[1863]_  = (~\new_[1929]_  | ~\new_[6394]_ ) & (~\new_[1324]_  | ~\new_[6453]_ );
  assign \new_[1864]_  = (~\new_[1929]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1311]_ );
  assign \new_[1865]_  = (~\new_[1929]_  | ~\new_[6356]_ ) & (~\new_[1312]_  | ~\new_[6092]_ );
  assign \new_[1866]_  = \\sbox1_ah_reg_reg[3] ;
  assign \new_[1867]_  = (~\new_[1929]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1315]_ );
  assign \new_[1868]_  = (~\new_[1929]_  | ~\new_[6365]_ ) & (~\new_[1314]_  | ~\new_[6436]_ );
  assign \new_[1869]_  = (~\new_[1929]_  | ~\new_[6362]_ ) & (~\new_[6417]_  | ~\new_[1322]_ );
  assign \new_[1870]_  = (~\new_[1929]_  | ~\new_[6366]_ ) & (~\new_[1323]_  | ~\new_[6435]_ );
  assign \new_[1871]_  = (~\new_[1929]_  | ~\new_[6359]_ ) & (~\new_[1313]_  | ~\new_[6170]_ );
  assign \new_[1872]_  = ~\new_[1896]_ ;
  assign \new_[1873]_  = ~\new_[1899]_ ;
  assign \new_[1874]_  = \new_[1322]_  ? \new_[7632]_  : \new_[1929]_ ;
  assign \new_[1875]_  = ~\new_[1922]_  & ~\new_[7826]_ ;
  assign \new_[1876]_  = ~\new_[1922]_  & ~\new_[6358]_ ;
  assign \new_[1877]_  = ~\new_[1934]_  & ~\new_[6363]_ ;
  assign \new_[1878]_  = ~\new_[1922]_  & ~\new_[6357]_ ;
  assign \new_[1879]_  = ~\new_[1934]_  & ~\new_[6361]_ ;
  assign \new_[1880]_  = ~\new_[1923]_  | ~\new_[8518]_ ;
  assign \new_[1881]_  = \new_[1932]_  ^ \new_[8707]_ ;
  assign \new_[1882]_  = ~\new_[1904]_ ;
  assign \new_[1883]_  = ~\new_[1906]_  & ~\new_[6808]_ ;
  assign \new_[1884]_  = ~\new_[1907]_  & ~\new_[6808]_ ;
  assign \new_[1885]_  = ~\new_[6803]_  & (~\new_[6086]_  | ~\new_[1926]_ );
  assign \new_[1886]_  = ~\new_[6954]_  & (~\new_[6087]_  | ~\new_[1927]_ );
  assign \new_[1887]_  = ~\new_[1908]_  & ~\new_[6808]_ ;
  assign \new_[1888]_  = ~\new_[6954]_  & (~\new_[6011]_  | ~\new_[1928]_ );
  assign \new_[1889]_  = ~\new_[1909]_  & ~\new_[6703]_ ;
  assign \new_[1890]_  = ~\new_[1910]_  & ~\new_[6808]_ ;
  assign \new_[1891]_  = ~\new_[1911]_  & ~\new_[6703]_ ;
  assign \new_[1892]_  = ~\new_[1924]_  | ~\new_[3359]_ ;
  assign \new_[1893]_  = (~\new_[6957]_  | ~\new_[8024]_ ) & (~\new_[1938]_  | ~\new_[7821]_ );
  assign \new_[1894]_  = (~\new_[1938]_  | ~\new_[6367]_ ) & (~\new_[6173]_  | ~\new_[1538]_ );
  assign \new_[1895]_  = (~\new_[1938]_  | ~\new_[7738]_ ) & (~\new_[1463]_  | ~\new_[7569]_ );
  assign \new_[1896]_  = \new_[8190]_ ;
  assign \new_[1897]_  = ~\new_[8190]_ ;
  assign \new_[1898]_  = ~\new_[1914]_ ;
  assign \new_[1899]_  = ~\new_[1925]_  | ~\new_[1933]_ ;
  assign \new_[1900]_  = ~\new_[1929]_  | ~\new_[6172]_ ;
  assign \new_[1901]_  = ~\new_[1929]_  | ~\new_[6355]_ ;
  assign \new_[1902]_  = ~\new_[1929]_  | ~\new_[6354]_ ;
  assign \new_[1903]_  = ~n1755 | ~\new_[8707]_ ;
  assign \new_[1904]_  = \new_[8707]_  ^ \new_[1945]_ ;
  assign \new_[1905]_  = (~\new_[6955]_  | ~\new_[8111]_ ) & (~\new_[1939]_  | ~\new_[7631]_ );
  assign \new_[1906]_  = (~\new_[1939]_  | ~\new_[6360]_ ) & (~\new_[6454]_  | ~\new_[1457]_ );
  assign \new_[1907]_  = (~\new_[1938]_  | ~\new_[6368]_ ) & (~\new_[6434]_  | ~\new_[1530]_ );
  assign \new_[1908]_  = (~\new_[1939]_  | ~\new_[6365]_ ) & (~\new_[1458]_  | ~\new_[6436]_ );
  assign \new_[1909]_  = (~\new_[1938]_  | ~\new_[6362]_ ) & (~\new_[6417]_  | ~\new_[1463]_ );
  assign \new_[1910]_  = (~\new_[1939]_  | ~\new_[6359]_ ) & (~\new_[6170]_  | ~\new_[1459]_ );
  assign \new_[1911]_  = (~\new_[1938]_  | ~\new_[6366]_ ) & (~\new_[1520]_  | ~\new_[6435]_ );
  assign \new_[1912]_  = (~\new_[1939]_  | ~\new_[6394]_ ) & (~\new_[1464]_  | ~\new_[6453]_ );
  assign \new_[1913]_  = (~\new_[1939]_  | ~\new_[6356]_ ) & (~\new_[6092]_  | ~\new_[1460]_ );
  assign \new_[1914]_  = \new_[1924]_ ;
  assign \new_[1915]_  = ~\new_[1924]_ ;
  assign \new_[1916]_  = \new_[1463]_  ? \new_[7569]_  : \new_[1939]_ ;
  assign \new_[1917]_  = ~\new_[1936]_  & ~\new_[6358]_ ;
  assign \new_[1918]_  = ~\new_[1936]_  & ~\new_[7826]_ ;
  assign \new_[1919]_  = ~\new_[1935]_  & ~\new_[6363]_ ;
  assign \new_[1920]_  = ~\new_[1936]_  & ~\new_[6357]_ ;
  assign \new_[1921]_  = ~\new_[1935]_  & ~\new_[6361]_ ;
  assign \new_[1922]_  = ~\new_[1929]_ ;
  assign \new_[1923]_  = \new_[1941]_  ^ \new_[8513]_ ;
  assign \new_[1924]_  = ~\new_[8214]_ ;
  assign \new_[1925]_  = ~\new_[1940]_  | ~\new_[3356]_ ;
  assign \new_[1926]_  = ~\new_[1939]_  | ~\new_[6172]_ ;
  assign \new_[1927]_  = ~\new_[1939]_  | ~\new_[6355]_ ;
  assign \new_[1928]_  = ~\new_[1939]_  | ~\new_[6354]_ ;
  assign \new_[1929]_  = ~\new_[1934]_ ;
  assign \new_[1930]_  = \new_[1986]_  ? \new_[8431]_  : \new_[2010]_ ;
  assign n1755 = ~\new_[8446]_ ;
  assign \new_[1932]_  = ~\new_[1944]_ ;
  assign \new_[1933]_  = ~\new_[8260]_  | ~\new_[3535]_ ;
  assign \new_[1934]_  = \new_[8766]_ ;
  assign \new_[1935]_  = ~\new_[1938]_ ;
  assign \new_[1936]_  = ~\new_[1939]_ ;
  assign \new_[1937]_  = ~\new_[8432]_ ;
  assign \new_[1938]_  = \new_[8259]_ ;
  assign \new_[1939]_  = \new_[8259]_ ;
  assign \new_[1940]_  = ~\new_[8260]_ ;
  assign \new_[1941]_  = ~\new_[1944]_ ;
  assign \new_[1942]_  = \\ks1_key_reg_reg[28] ;
  assign \new_[1943]_  = ~\new_[1968]_  | ~\new_[1954]_ ;
  assign \new_[1944]_  = ~\new_[1948]_ ;
  assign \new_[1945]_  = ~\new_[8514]_ ;
  assign \new_[1946]_  = \\ks1_key_reg_reg[27] ;
  assign \new_[1947]_  = \\ks1_key_reg_reg[29] ;
  assign \new_[1948]_  = ~\new_[1972]_  | ~\new_[1985]_ ;
  assign \new_[1949]_  = \\ks1_key_reg_reg[30] ;
  assign \new_[1950]_  = \\ks1_key_reg_reg[24] ;
  assign \new_[1951]_  = \\ks1_key_reg_reg[31] ;
  assign \new_[1952]_  = \\ks1_key_reg_reg[25] ;
  assign \new_[1953]_  = ~\new_[8165]_  | ~\new_[8215]_ ;
  assign \new_[1954]_  = ~\new_[8164]_  | ~\new_[8876]_ ;
  assign \new_[1955]_  = \\ks1_key_reg_reg[26] ;
  assign n1760 = \new_[1942]_  ? \new_[7597]_  : \new_[2017]_ ;
  assign \new_[1957]_  = ~\new_[2036]_  | ~\new_[1994]_ ;
  assign \new_[1958]_  = ~\\ks1_key_reg_reg[60] ;
  assign \new_[1959]_  = \\ks1_key_reg_reg[2] ;
  assign \new_[1960]_  = \\ks1_key_reg_reg[3] ;
  assign \new_[1961]_  = \\ks1_key_reg_reg[4] ;
  assign \new_[1962]_  = \\ks1_key_reg_reg[5] ;
  assign \new_[1963]_  = \\ks1_key_reg_reg[6] ;
  assign \new_[1964]_  = \\ks1_key_reg_reg[0] ;
  assign \new_[1965]_  = \\ks1_key_reg_reg[1] ;
  assign \new_[1966]_  = \\ks1_key_reg_reg[23] ;
  assign \new_[1967]_  = ~\new_[2012]_  | ~\new_[8166]_ ;
  assign \new_[1968]_  = ~\new_[8166]_  | ~\new_[2013]_ ;
  assign \new_[1969]_  = \\ks1_key_reg_reg[7] ;
  assign \new_[1970]_  = ~\new_[2011]_  | ~\new_[2050]_ ;
  assign \new_[1971]_  = ~\new_[2014]_  | ~\new_[8347]_ ;
  assign \new_[1972]_  = ~\new_[2050]_  | ~\new_[2015]_ ;
  assign n1765 = \new_[1946]_  ? \new_[7597]_  : \new_[2039]_ ;
  assign n1770 = \new_[1947]_  ? \new_[7470]_  : \new_[2040]_ ;
  assign \new_[1975]_  = ~\\ks1_key_reg_reg[61] ;
  assign \new_[1976]_  = ~\\ks1_key_reg_reg[59] ;
  assign \new_[1977]_  = \\ks1_key_reg_reg[17] ;
  assign \new_[1978]_  = \\ks1_key_reg_reg[16] ;
  assign \new_[1979]_  = \\ks1_key_reg_reg[19] ;
  assign \new_[1980]_  = \\ks1_key_reg_reg[18] ;
  assign \new_[1981]_  = \\ks1_key_reg_reg[21] ;
  assign \new_[1982]_  = \\ks1_key_reg_reg[22] ;
  assign \new_[1983]_  = ~\new_[8580]_  | ~\new_[8585]_ ;
  assign \new_[1984]_  = ~\new_[8430]_  | ~\new_[2038]_ ;
  assign \new_[1985]_  = ~\new_[2038]_  | ~\new_[2037]_ ;
  assign \new_[1986]_  = ~\new_[2010]_ ;
  assign \new_[1987]_  = ~\new_[8429]_ ;
  assign n1785 = \new_[1951]_  ? \new_[7597]_  : \new_[2061]_ ;
  assign n1775 = \new_[1949]_  ? \new_[7597]_  : \new_[2060]_ ;
  assign n1780 = \new_[1950]_  ? \new_[7597]_  : \new_[2062]_ ;
  assign n1790 = \new_[1952]_  ? \new_[7597]_  : \new_[2053]_ ;
  assign n1795 = \new_[1955]_  ? \new_[7470]_  : \new_[2054]_ ;
  assign \new_[1993]_  = \\ks1_key_reg_reg[20] ;
  assign \new_[1994]_  = ~\new_[8347]_ ;
  assign n1810 = \new_[1960]_  ? \new_[7597]_  : \new_[2080]_ ;
  assign n1815 = \new_[1961]_  ? \new_[7597]_  : \new_[2081]_ ;
  assign n1820 = \new_[1962]_  ? \new_[7470]_  : \new_[2082]_ ;
  assign n1825 = \new_[1963]_  ? \new_[7597]_  : \new_[2083]_ ;
  assign n1845 = \new_[1969]_  ? \new_[7597]_  : \new_[2084]_ ;
  assign n1830 = \new_[1964]_  ? \new_[8843]_  : \new_[2085]_ ;
  assign n1835 = \new_[1965]_  ? \new_[7597]_  : \new_[2086]_ ;
  assign n1840 = \new_[1966]_  ? \new_[7597]_  : \new_[2087]_ ;
  assign n1805 = \new_[1959]_  ? \new_[7597]_  : \new_[2088]_ ;
  assign \new_[2004]_  = ~\\ks1_key_reg_reg[57] ;
  assign \new_[2005]_  = ~\\ks1_key_reg_reg[58] ;
  assign \new_[2006]_  = ~\\ks1_key_reg_reg[63] ;
  assign \new_[2007]_  = ~\\ks1_key_reg_reg[62] ;
  assign \new_[2008]_  = ~\new_[8655]_  | ~\new_[4464]_ ;
  assign \new_[2009]_  = ~\\ks1_key_reg_reg[56] ;
  assign \new_[2010]_  = \new_[2094]_  ? \new_[8373]_  : \new_[8387]_ ;
  assign \new_[2011]_  = ~\new_[8430]_ ;
  assign \new_[2012]_  = ~\new_[8215]_ ;
  assign \new_[2013]_  = ~\new_[8876]_ ;
  assign \new_[2014]_  = ~\new_[2036]_ ;
  assign \new_[2015]_  = ~\new_[2037]_ ;
  assign n1800 = (~\new_[2064]_  & ~\new_[8343]_ ) | (~\new_[7410]_  & ~\new_[1958]_ );
  assign \new_[2017]_  = \new_[9017]_  ^ \new_[2064]_ ;
  assign n1865 = \new_[1978]_  ? \new_[7597]_  : \new_[2151]_ ;
  assign n1860 = \new_[1977]_  ? \new_[7470]_  : \new_[2152]_ ;
  assign n1875 = \new_[1980]_  ? \new_[7597]_  : \new_[2153]_ ;
  assign n1870 = \new_[1979]_  ? \new_[7470]_  : \new_[2154]_ ;
  assign n1890 = \new_[1993]_  ? \new_[7597]_  : \new_[2155]_ ;
  assign n1880 = \new_[1981]_  ? \new_[7597]_  : \new_[2156]_ ;
  assign n1885 = \new_[1982]_  ? \new_[7597]_  : \new_[2157]_ ;
  assign \new_[2025]_  = ~\\ks1_key_reg_reg[92] ;
  assign \new_[2026]_  = ~\\ks1_key_reg_reg[32] ;
  assign \new_[2027]_  = ~\\ks1_key_reg_reg[33] ;
  assign \new_[2028]_  = ~\\ks1_key_reg_reg[34] ;
  assign \new_[2029]_  = ~\\ks1_key_reg_reg[35] ;
  assign \new_[2030]_  = ~\\ks1_key_reg_reg[36] ;
  assign \new_[2031]_  = ~\\ks1_key_reg_reg[38] ;
  assign \new_[2032]_  = ~\\ks1_key_reg_reg[39] ;
  assign \new_[2033]_  = ~\\ks1_key_reg_reg[55] ;
  assign \new_[2034]_  = ~\\ks1_key_reg_reg[37] ;
  assign \new_[2035]_  = ~\new_[8368]_  | ~\new_[4542]_ ;
  assign \new_[2036]_  = ~\new_[2092]_  | ~\new_[2663]_ ;
  assign \new_[2037]_  = ~\new_[2093]_  | ~\new_[2664]_ ;
  assign \new_[2038]_  = ~\new_[2050]_ ;
  assign \new_[2039]_  = \new_[8396]_  ^ \new_[2142]_ ;
  assign \new_[2040]_  = \new_[4524]_  ^ \new_[2143]_ ;
  assign n1855 = \new_[7957]_  ? \new_[7470]_  : \new_[2142]_ ;
  assign n1850 = \new_[8001]_  ? \new_[7597]_  : \new_[2143]_ ;
  assign \new_[2043]_  = \\ks1_key_reg_reg[91] ;
  assign \new_[2044]_  = ~\\ks1_key_reg_reg[93] ;
  assign \new_[2045]_  = ~\\ks1_key_reg_reg[49] ;
  assign \new_[2046]_  = ~\\ks1_key_reg_reg[50] ;
  assign \new_[2047]_  = ~\\ks1_key_reg_reg[51] ;
  assign \new_[2048]_  = ~\\ks1_key_reg_reg[52] ;
  assign \new_[2049]_  = ~\\ks1_key_reg_reg[54] ;
  assign \new_[2050]_  = ~\new_[8718]_  | ~\new_[2557]_ ;
  assign \new_[2051]_  = ~\\ks1_key_reg_reg[48] ;
  assign \new_[2052]_  = ~\\ks1_key_reg_reg[53] ;
  assign \new_[2053]_  = \new_[8277]_  ^ \new_[2212]_ ;
  assign \new_[2054]_  = \new_[4515]_  ^ \new_[2213]_ ;
  assign n1895 = \new_[8124]_  ? \new_[7470]_  : \new_[2212]_ ;
  assign n1900 = \new_[8055]_  ? \new_[7470]_  : \new_[2213]_ ;
  assign n1915 = \new_[8000]_  ? \new_[7597]_  : \new_[2211]_ ;
  assign n1910 = \new_[8005]_  ? \new_[7597]_  : \new_[2209]_ ;
  assign n1905 = \new_[7941]_  ? \new_[7597]_  : \new_[2210]_ ;
  assign \new_[2060]_  = \new_[8358]_  ^ \new_[2209]_ ;
  assign \new_[2061]_  = \new_[4507]_  ^ \new_[2210]_ ;
  assign \new_[2062]_  = \new_[4514]_  ^ \new_[2211]_ ;
  assign \new_[2063]_  = \new_[2810]_  ^ \new_[8383]_ ;
  assign \new_[2064]_  = \new_[2970]_  ^ \new_[2275]_ ;
  assign n1920 = \new_[8151]_  ? \new_[7597]_  : \new_[2275]_ ;
  assign \new_[2066]_  = ~\\ks1_key_reg_reg[90] ;
  assign \new_[2067]_  = \\ks1_key_reg_reg[88] ;
  assign \new_[2068]_  = \\ks1_key_reg_reg[94] ;
  assign \new_[2069]_  = \\ks1_key_reg_reg[95] ;
  assign \new_[2070]_  = \\ks1_key_reg_reg[89] ;
  assign n1925 = (~\new_[2287]_  & ~\new_[7573]_ ) | (~\new_[7469]_  & ~\new_[2026]_ );
  assign n1930 = (~\new_[2289]_  & ~\new_[7573]_ ) | (~\new_[7410]_  & ~\new_[2027]_ );
  assign n1935 = (~\new_[2291]_  & ~\new_[7573]_ ) | (~\new_[7469]_  & ~\new_[2028]_ );
  assign n1940 = (~\new_[2282]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2029]_ );
  assign n1945 = (~\new_[2283]_  & ~\new_[8343]_ ) | (~\new_[7597]_  & ~\new_[2030]_ );
  assign n1965 = (~\new_[2284]_  & ~\new_[7573]_ ) | (~\new_[7597]_  & ~\new_[2034]_ );
  assign n1950 = (~\new_[2285]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2031]_ );
  assign n1955 = (~\new_[2286]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2032]_ );
  assign n1960 = (~\new_[2290]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2033]_ );
  assign \new_[2080]_  = \new_[4508]_  ^ \new_[2282]_ ;
  assign \new_[2081]_  = \new_[4432]_  ^ \new_[2283]_ ;
  assign \new_[2082]_  = \new_[8878]_  ^ \new_[2284]_ ;
  assign \new_[2083]_  = \new_[8250]_  ^ \new_[2285]_ ;
  assign \new_[2084]_  = \new_[4435]_  ^ \new_[2286]_ ;
  assign \new_[2085]_  = \new_[4618]_  ^ \new_[2287]_ ;
  assign \new_[2086]_  = \new_[8968]_  ^ \new_[2289]_ ;
  assign \new_[2087]_  = \new_[4513]_  ^ \new_[2290]_ ;
  assign \new_[2088]_  = \new_[4617]_  ^ \new_[2291]_ ;
  assign \new_[2089]_  = ~\new_[8854]_ ;
  assign \new_[2090]_  = ~\new_[8339]_ ;
  assign \new_[2091]_  = ~\new_[2217]_  | ~\new_[8725]_ ;
  assign \new_[2092]_  = ~\new_[2160]_  | ~\new_[8725]_ ;
  assign \new_[2093]_  = ~\new_[2161]_  | ~\new_[8725]_ ;
  assign \new_[2094]_  = ~\new_[2159]_  & (~\new_[2442]_  | ~\new_[2355]_ );
  assign \new_[2095]_  = \\ks1_key_reg_reg[69] ;
  assign \data_o[60]  = \\addroundkey_data_reg_reg[60] ;
  assign \data_o[111]  = \\addroundkey_data_reg_reg[111] ;
  assign \data_o[63]  = \\addroundkey_data_reg_reg[63] ;
  assign \data_o[6]  = \\addroundkey_data_reg_reg[6] ;
  assign \data_o[76]  = \\addroundkey_data_reg_reg[76] ;
  assign \data_o[25]  = \\addroundkey_data_reg_reg[25] ;
  assign \data_o[77]  = \\addroundkey_data_reg_reg[77] ;
  assign \data_o[78]  = \\addroundkey_data_reg_reg[78] ;
  assign \data_o[79]  = \\addroundkey_data_reg_reg[79] ;
  assign \data_o[26]  = \\addroundkey_data_reg_reg[26] ;
  assign \data_o[29]  = \\addroundkey_data_reg_reg[29] ;
  assign \data_o[8]  = \\addroundkey_data_reg_reg[8] ;
  assign \data_o[105]  = \\addroundkey_data_reg_reg[105] ;
  assign \data_o[0]  = \\addroundkey_data_reg_reg[0] ;
  assign \data_o[106]  = \\addroundkey_data_reg_reg[106] ;
  assign \data_o[107]  = \\addroundkey_data_reg_reg[107] ;
  assign \data_o[122]  = \\addroundkey_data_reg_reg[122] ;
  assign \data_o[3]  = \\addroundkey_data_reg_reg[3] ;
  assign \data_o[41]  = \\addroundkey_data_reg_reg[41] ;
  assign \data_o[123]  = \\addroundkey_data_reg_reg[123] ;
  assign \data_o[42]  = \\addroundkey_data_reg_reg[42] ;
  assign \data_o[43]  = \\addroundkey_data_reg_reg[43] ;
  assign \data_o[44]  = \\addroundkey_data_reg_reg[44] ;
  assign \data_o[108]  = \\addroundkey_data_reg_reg[108] ;
  assign \data_o[125]  = \\addroundkey_data_reg_reg[125] ;
  assign \data_o[46]  = \\addroundkey_data_reg_reg[46] ;
  assign \data_o[47]  = \\addroundkey_data_reg_reg[47] ;
  assign \data_o[126]  = \\addroundkey_data_reg_reg[126] ;
  assign \data_o[127]  = \\addroundkey_data_reg_reg[127] ;
  assign \data_o[10]  = \\addroundkey_data_reg_reg[10] ;
  assign \data_o[13]  = \\addroundkey_data_reg_reg[13] ;
  assign \data_o[110]  = \\addroundkey_data_reg_reg[110] ;
  assign \data_o[58]  = \\addroundkey_data_reg_reg[58] ;
  assign \data_o[57]  = \\addroundkey_data_reg_reg[57] ;
  assign \data_o[59]  = \\addroundkey_data_reg_reg[59] ;
  assign \new_[2131]_  = \\ks1_key_reg_reg[124] ;
  assign \new_[2132]_  = \\ks1_key_reg_reg[64] ;
  assign \new_[2133]_  = \\ks1_key_reg_reg[65] ;
  assign \new_[2134]_  = \\ks1_key_reg_reg[67] ;
  assign \new_[2135]_  = \\ks1_key_reg_reg[66] ;
  assign \new_[2136]_  = \\ks1_key_reg_reg[68] ;
  assign \new_[2137]_  = \\ks1_key_reg_reg[70] ;
  assign \new_[2138]_  = \\ks1_key_reg_reg[71] ;
  assign \new_[2139]_  = \\ks1_key_reg_reg[87] ;
  assign n1970 = \new_[2043]_  ? \new_[7597]_  : \new_[2358]_ ;
  assign n1975 = (~\new_[2359]_  & ~\new_[8343]_ ) | (~\new_[7410]_  & ~\new_[2044]_ );
  assign \new_[2142]_  = \new_[2969]_  ^ \new_[2358]_ ;
  assign \new_[2143]_  = \new_[3079]_  ^ \new_[2359]_ ;
  assign n2005 = (~\new_[2362]_  & ~\new_[8343]_ ) | (~\new_[7410]_  & ~\new_[2051]_ );
  assign n1980 = (~\new_[2363]_  & ~\new_[7573]_ ) | (~\new_[7410]_  & ~\new_[2045]_ );
  assign n1985 = (~\new_[2364]_  & ~\new_[7573]_ ) | (~\new_[7410]_  & ~\new_[2046]_ );
  assign n1990 = (~\new_[2365]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2047]_ );
  assign n1995 = (~\new_[2366]_  & ~\new_[7573]_ ) | (~\new_[7410]_  & ~\new_[2048]_ );
  assign n2010 = (~\new_[2367]_  & ~\new_[8343]_ ) | (~\new_[7597]_  & ~\new_[2052]_ );
  assign n2000 = (~\new_[2368]_  & ~\new_[7573]_ ) | (~\new_[7597]_  & ~\new_[2049]_ );
  assign \new_[2151]_  = \new_[8785]_  ^ \new_[2362]_ ;
  assign \new_[2152]_  = \new_[8330]_  ^ \new_[2363]_ ;
  assign \new_[2153]_  = \new_[4620]_  ^ \new_[2364]_ ;
  assign \new_[2154]_  = \new_[8278]_  ^ \new_[2365]_ ;
  assign \new_[2155]_  = \new_[8312]_  ^ \new_[2366]_ ;
  assign \new_[2156]_  = \new_[4438]_  ^ \new_[2367]_ ;
  assign \new_[2157]_  = \new_[8297]_  ^ \new_[2368]_ ;
  assign \data_o[5]  = \\addroundkey_data_reg_reg[5] ;
  assign \new_[2159]_  = ~\new_[2442]_  & ~\new_[2355]_ ;
  assign \new_[2160]_  = \new_[3292]_  ? \new_[8447]_  : \new_[3041]_ ;
  assign \new_[2161]_  = \new_[8385]_  ? \new_[8447]_  : \new_[8387]_ ;
  assign \new_[2162]_  = \\ks1_key_reg_reg[81] ;
  assign \data_o[40]  = \\addroundkey_data_reg_reg[40] ;
  assign \data_o[124]  = \\addroundkey_data_reg_reg[124] ;
  assign \data_o[61]  = \\addroundkey_data_reg_reg[61] ;
  assign \data_o[62]  = \\addroundkey_data_reg_reg[62] ;
  assign \data_o[1]  = \\addroundkey_data_reg_reg[1] ;
  assign \data_o[73]  = \\addroundkey_data_reg_reg[73] ;
  assign \data_o[74]  = \\addroundkey_data_reg_reg[74] ;
  assign \data_o[24]  = \\addroundkey_data_reg_reg[24] ;
  assign \data_o[72]  = \\addroundkey_data_reg_reg[72] ;
  assign \data_o[7]  = \\addroundkey_data_reg_reg[7] ;
  assign \data_o[28]  = \\addroundkey_data_reg_reg[28] ;
  assign \data_o[104]  = \\addroundkey_data_reg_reg[104] ;
  assign \data_o[30]  = \\addroundkey_data_reg_reg[30] ;
  assign \data_o[2]  = \\addroundkey_data_reg_reg[2] ;
  assign \data_o[31]  = \\addroundkey_data_reg_reg[31] ;
  assign \data_o[90]  = \\addroundkey_data_reg_reg[90] ;
  assign \data_o[91]  = \\addroundkey_data_reg_reg[91] ;
  assign \data_o[92]  = \\addroundkey_data_reg_reg[92] ;
  assign \data_o[34]  = \\addroundkey_data_reg_reg[34] ;
  assign \data_o[93]  = \\addroundkey_data_reg_reg[93] ;
  assign \data_o[11]  = \\addroundkey_data_reg_reg[11] ;
  assign \data_o[94]  = \\addroundkey_data_reg_reg[94] ;
  assign \data_o[95]  = \\addroundkey_data_reg_reg[95] ;
  assign \data_o[120]  = \\addroundkey_data_reg_reg[120] ;
  assign \data_o[9]  = \\addroundkey_data_reg_reg[9] ;
  assign \data_o[121]  = \\addroundkey_data_reg_reg[121] ;
  assign \data_o[45]  = \\addroundkey_data_reg_reg[45] ;
  assign \data_o[4]  = \\addroundkey_data_reg_reg[4] ;
  assign \data_o[12]  = \\addroundkey_data_reg_reg[12] ;
  assign \data_o[109]  = \\addroundkey_data_reg_reg[109] ;
  assign \data_o[14]  = \\addroundkey_data_reg_reg[14] ;
  assign \data_o[56]  = \\addroundkey_data_reg_reg[56] ;
  assign \data_o[15]  = \\addroundkey_data_reg_reg[15] ;
  assign \new_[2196]_  = \\ks1_key_reg_reg[125] ;
  assign \new_[2197]_  = \\ks1_key_reg_reg[123] ;
  assign \new_[2198]_  = \\ks1_key_reg_reg[80] ;
  assign \new_[2199]_  = \\ks1_key_reg_reg[83] ;
  assign \new_[2200]_  = \\ks1_key_reg_reg[84] ;
  assign \new_[2201]_  = \\ks1_key_reg_reg[85] ;
  assign \new_[2202]_  = \\ks1_key_reg_reg[82] ;
  assign \new_[2203]_  = \\ks1_key_reg_reg[86] ;
  assign n2020 = \new_[2067]_  ? \new_[7597]_  : \new_[2441]_ ;
  assign n2035 = \new_[2070]_  ? \new_[7597]_  : \new_[2432]_ ;
  assign n2015 = (~\new_[2433]_  & ~\new_[8343]_ ) | (~\new_[7469]_  & ~\new_[2066]_ );
  assign n2025 = \new_[2068]_  ? \new_[8843]_  : \new_[2439]_ ;
  assign n2030 = \new_[2069]_  ? \new_[7597]_  : \new_[2440]_ ;
  assign \new_[2209]_  = \new_[2834]_  ^ \new_[2439]_ ;
  assign \new_[2210]_  = \new_[2835]_  ^ \new_[2440]_ ;
  assign \new_[2211]_  = \new_[2967]_  ^ \new_[2441]_ ;
  assign \new_[2212]_  = \new_[2968]_  ^ \new_[2432]_ ;
  assign \new_[2213]_  = \new_[3078]_  ^ \new_[2433]_ ;
  assign \data_o[27]  = \\addroundkey_data_reg_reg[27] ;
  assign \data_o[75]  = \\addroundkey_data_reg_reg[75] ;
  assign \new_[2216]_  = ~\new_[8629]_ ;
  assign \new_[2217]_  = \new_[3293]_  ? \new_[2427]_  : \new_[3042]_ ;
  assign \new_[2218]_  = \new_[3003]_  ^ \new_[8721]_ ;
  assign \data_o[100]  = \\addroundkey_data_reg_reg[100] ;
  assign \data_o[33]  = \\addroundkey_data_reg_reg[33] ;
  assign \data_o[103]  = \\addroundkey_data_reg_reg[103] ;
  assign \data_o[98]  = \\addroundkey_data_reg_reg[98] ;
  assign \data_o[35]  = \\addroundkey_data_reg_reg[35] ;
  assign \new_[2224]_  = ~\\mix1_data_reg_reg[100] ;
  assign \new_[2225]_  = ~\\mix1_data_reg_reg[108] ;
  assign \new_[2226]_  = ~\\mix1_data_reg_reg[116] ;
  assign \new_[2227]_  = ~\\mix1_data_reg_reg[124] ;
  assign \data_o[101]  = \\addroundkey_data_reg_reg[101] ;
  assign \data_o[112]  = \\addroundkey_data_reg_reg[112] ;
  assign \data_o[64]  = \\addroundkey_data_reg_reg[64] ;
  assign \data_o[65]  = \\addroundkey_data_reg_reg[65] ;
  assign \data_o[20]  = \\addroundkey_data_reg_reg[20] ;
  assign \data_o[66]  = \\addroundkey_data_reg_reg[66] ;
  assign \data_o[67]  = \\addroundkey_data_reg_reg[67] ;
  assign \data_o[21]  = \\addroundkey_data_reg_reg[21] ;
  assign \data_o[69]  = \\addroundkey_data_reg_reg[69] ;
  assign \data_o[22]  = \\addroundkey_data_reg_reg[22] ;
  assign \data_o[70]  = \\addroundkey_data_reg_reg[70] ;
  assign \data_o[102]  = \\addroundkey_data_reg_reg[102] ;
  assign \data_o[23]  = \\addroundkey_data_reg_reg[23] ;
  assign \data_o[115]  = \\addroundkey_data_reg_reg[115] ;
  assign \data_o[116]  = \\addroundkey_data_reg_reg[116] ;
  assign \data_o[80]  = \\addroundkey_data_reg_reg[80] ;
  assign \data_o[81]  = \\addroundkey_data_reg_reg[81] ;
  assign \data_o[83]  = \\addroundkey_data_reg_reg[83] ;
  assign \data_o[85]  = \\addroundkey_data_reg_reg[85] ;
  assign \data_o[86]  = \\addroundkey_data_reg_reg[86] ;
  assign \data_o[84]  = \\addroundkey_data_reg_reg[84] ;
  assign \data_o[87]  = \\addroundkey_data_reg_reg[87] ;
  assign \data_o[88]  = \\addroundkey_data_reg_reg[88] ;
  assign \data_o[32]  = \\addroundkey_data_reg_reg[32] ;
  assign \data_o[119]  = \\addroundkey_data_reg_reg[119] ;
  assign \data_o[96]  = \\addroundkey_data_reg_reg[96] ;
  assign \data_o[97]  = \\addroundkey_data_reg_reg[97] ;
  assign \data_o[36]  = \\addroundkey_data_reg_reg[36] ;
  assign \data_o[99]  = \\addroundkey_data_reg_reg[99] ;
  assign \data_o[37]  = \\addroundkey_data_reg_reg[37] ;
  assign \data_o[38]  = \\addroundkey_data_reg_reg[38] ;
  assign \data_o[39]  = \\addroundkey_data_reg_reg[39] ;
  assign \data_o[49]  = \\addroundkey_data_reg_reg[49] ;
  assign \data_o[52]  = \\addroundkey_data_reg_reg[52] ;
  assign \data_o[55]  = \\addroundkey_data_reg_reg[55] ;
  assign \data_o[17]  = \\addroundkey_data_reg_reg[17] ;
  assign \new_[2264]_  = \\ks1_key_reg_reg[120] ;
  assign \new_[2265]_  = \\ks1_key_reg_reg[121] ;
  assign \new_[2266]_  = \\ks1_key_reg_reg[127] ;
  assign \new_[2267]_  = \\addroundkey_round_reg[0] ;
  assign \data_o[118]  = \\addroundkey_data_reg_reg[118] ;
  assign \data_o[89]  = \\addroundkey_data_reg_reg[89] ;
  assign \data_o[117]  = \\addroundkey_data_reg_reg[117] ;
  assign \new_[2271]_  = \\ks1_key_reg_reg[126] ;
  assign \data_o[82]  = \\addroundkey_data_reg_reg[82] ;
  assign \new_[2273]_  = \\ks1_key_reg_reg[122] ;
  assign n2220 = \new_[2131]_  ? \new_[7597]_  : \new_[2559]_ ;
  assign \new_[2275]_  = \new_[3375]_  ^ \new_[2559]_ ;
  assign \data_o[114]  = \\addroundkey_data_reg_reg[114] ;
  assign \data_o[54]  = \\addroundkey_data_reg_reg[54] ;
  assign \data_o[71]  = \\addroundkey_data_reg_reg[71] ;
  assign \data_o[16]  = \\addroundkey_data_reg_reg[16] ;
  assign \data_o[68]  = \\addroundkey_data_reg_reg[68] ;
  assign \data_o[53]  = \\addroundkey_data_reg_reg[53] ;
  assign \new_[2282]_  = \new_[2839]_  ^ \new_[2568]_ ;
  assign \new_[2283]_  = \new_[2840]_  ^ \new_[2569]_ ;
  assign \new_[2284]_  = \new_[2841]_  ^ \new_[2570]_ ;
  assign \new_[2285]_  = \new_[2993]_  ^ \new_[2571]_ ;
  assign \new_[2286]_  = \new_[2994]_  ^ \new_[2572]_ ;
  assign \new_[2287]_  = \new_[2573]_  ^ \new_[2956]_ ;
  assign \data_o[113]  = \\addroundkey_data_reg_reg[113] ;
  assign \new_[2289]_  = \new_[2574]_  ^ \new_[2962]_ ;
  assign \new_[2290]_  = \new_[2575]_  ^ \new_[2966]_ ;
  assign \new_[2291]_  = \new_[2576]_  ^ \new_[2971]_ ;
  assign n2225 = \new_[2132]_  ? \new_[7470]_  : \new_[2573]_ ;
  assign n2230 = \new_[2133]_  ? \new_[7470]_  : \new_[2574]_ ;
  assign n2240 = \new_[2135]_  ? \new_[7470]_  : \new_[2576]_ ;
  assign n2235 = \new_[2134]_  ? \new_[7470]_  : \new_[2568]_ ;
  assign n2245 = \new_[2136]_  ? \new_[7470]_  : \new_[2569]_ ;
  assign n2040 = \new_[2095]_  ? \new_[7470]_  : \new_[2570]_ ;
  assign n2250 = \new_[2137]_  ? \new_[7597]_  : \new_[2571]_ ;
  assign n2255 = \new_[2138]_  ? \new_[7470]_  : \new_[2572]_ ;
  assign n2260 = \new_[2139]_  ? \new_[7597]_  : \new_[2575]_ ;
  assign \new_[2301]_  = ~\new_[8877]_  | ~\new_[8582]_ ;
  assign \new_[2302]_  = ~\new_[8216]_  | ~\new_[8583]_ ;
  assign n2055 = ~\new_[2502]_  | (~\new_[3741]_  & ~\new_[8961]_ );
  assign \data_o[19]  = \\addroundkey_data_reg_reg[19] ;
  assign \data_o[51]  = \\addroundkey_data_reg_reg[51] ;
  assign n2060 = ~\new_[2503]_  | (~\new_[3742]_  & ~\new_[8955]_ );
  assign \data_o[50]  = \\addroundkey_data_reg_reg[50] ;
  assign \data_o[18]  = \\addroundkey_data_reg_reg[18] ;
  assign n2070 = ~\new_[2505]_  | (~\new_[3743]_  & ~\new_[8957]_ );
  assign n2065 = ~\new_[2504]_  | (~\new_[3744]_  & ~\new_[8961]_ );
  assign n2075 = ~\new_[2506]_  | (~\new_[3745]_  & ~\new_[8957]_ );
  assign n2090 = ~\new_[2508]_  | (~\new_[3746]_  & ~\new_[8957]_ );
  assign n2080 = ~\new_[2507]_  | (~\new_[3747]_  & ~\new_[8961]_ );
  assign n2085 = ~\new_[2509]_  | (~\new_[3748]_  & ~\new_[8957]_ );
  assign n2095 = ~\new_[2510]_  | (~\new_[3749]_  & ~\new_[8961]_ );
  assign n2100 = ~\new_[2511]_  | (~\new_[3750]_  & ~\new_[8958]_ );
  assign n2105 = ~\new_[2512]_  | (~\new_[3751]_  & ~\new_[8957]_ );
  assign n2115 = ~\new_[2514]_  | (~\new_[3752]_  & ~\new_[8958]_ );
  assign n2125 = ~\new_[2515]_  | (~\new_[3753]_  & ~\new_[8961]_ );
  assign n2130 = ~\new_[2513]_  | (~\new_[3754]_  & ~\new_[8958]_ );
  assign n2110 = ~\new_[2533]_  | (~\new_[3755]_  & ~\new_[8957]_ );
  assign n2140 = ~\new_[2516]_  | (~\new_[3756]_  & ~\new_[8957]_ );
  assign n2135 = ~\new_[2517]_  | (~\new_[3758]_  & ~\new_[8961]_ );
  assign n2175 = ~\new_[2525]_  | (~\new_[3766]_  & ~\new_[8961]_ );
  assign n2145 = ~\new_[2518]_  | (~\new_[3760]_  & ~\new_[8961]_ );
  assign n2150 = ~\new_[2519]_  | (~\new_[3762]_  & ~\new_[8958]_ );
  assign n2120 = ~\new_[2520]_  | (~\new_[3757]_  & ~\new_[8961]_ );
  assign n2165 = ~\new_[2522]_  | (~\new_[3764]_  & ~\new_[8961]_ );
  assign n2155 = ~\new_[2521]_  | (~\new_[3763]_  & ~\new_[8956]_ );
  assign n2160 = ~\new_[2526]_  | (~\new_[3767]_  & ~\new_[8958]_ );
  assign n2170 = ~\new_[2523]_  | (~\new_[3765]_  & ~\new_[8958]_ );
  assign n2180 = ~\new_[2524]_  | (~\new_[3761]_  & ~\new_[8960]_ );
  assign n2185 = ~\new_[2527]_  | (~\new_[3768]_  & ~\new_[8960]_ );
  assign \data_o[48]  = \\addroundkey_data_reg_reg[48] ;
  assign n2190 = ~\new_[2529]_  | (~\new_[3770]_  & ~\new_[8961]_ );
  assign n2195 = ~\new_[2528]_  | (~\new_[3769]_  & ~\new_[8956]_ );
  assign n2200 = ~\new_[2530]_  | (~\new_[3771]_  & ~\new_[8960]_ );
  assign n2210 = ~\new_[2531]_  | (~\new_[3772]_  & ~\new_[8958]_ );
  assign n2205 = ~\new_[2532]_  | (~\new_[3773]_  & ~\new_[8957]_ );
  assign n2215 = ~\new_[2534]_  | (~\new_[3774]_  & ~\new_[8961]_ );
  assign n2050 = ~\new_[2501]_  | (~\new_[3776]_  & ~\new_[8961]_ );
  assign n2265 = ~\new_[2535]_  | (~\new_[3775]_  & ~\new_[8958]_ );
  assign n2045 = ~\new_[2536]_  | (~\new_[3777]_  & ~\new_[8958]_ );
  assign \new_[2344]_  = \\ks1_key_reg_reg[97] ;
  assign \new_[2345]_  = ~\\mix1_data_reg_reg[107] ;
  assign \new_[2346]_  = ~\\mix1_data_reg_reg[115] ;
  assign \new_[2347]_  = ~\\mix1_data_reg_reg[99] ;
  assign \new_[2348]_  = \\ks1_key_reg_reg[96] ;
  assign \new_[2349]_  = \\ks1_key_reg_reg[98] ;
  assign \new_[2350]_  = \\ks1_key_reg_reg[100] ;
  assign \new_[2351]_  = \\ks1_key_reg_reg[101] ;
  assign \new_[2352]_  = \\ks1_key_reg_reg[102] ;
  assign \new_[2353]_  = \\ks1_key_reg_reg[103] ;
  assign \new_[2354]_  = \\ks1_key_reg_reg[119] ;
  assign \new_[2355]_  = ~\new_[2427]_ ;
  assign \new_[2356]_  = ~\\mix1_data_reg_reg[123] ;
  assign \new_[2357]_  = ~\new_[2558]_  | ~\new_[8724]_ ;
  assign \new_[2358]_  = \new_[3374]_  ^ \new_[2676]_ ;
  assign \new_[2359]_  = \new_[3102]_  ^ \new_[2675]_ ;
  assign n2445 = \new_[2197]_  ? \new_[7597]_  : \new_[2676]_ ;
  assign n2440 = \new_[2196]_  ? \new_[7597]_  : \new_[2675]_ ;
  assign \new_[2362]_  = \new_[2684]_  ^ \new_[2958]_ ;
  assign \new_[2363]_  = \new_[2685]_  ^ \new_[2959]_ ;
  assign \new_[2364]_  = \new_[2686]_  ^ \new_[2960]_ ;
  assign \new_[2365]_  = \new_[2687]_  ^ \new_[2961]_ ;
  assign \new_[2366]_  = \new_[2688]_  ^ \new_[2963]_ ;
  assign \new_[2367]_  = \new_[2689]_  ^ \new_[2964]_ ;
  assign \new_[2368]_  = \new_[2690]_  ^ \new_[2965]_ ;
  assign n2450 = \new_[2198]_  ? \new_[7470]_  : \new_[2684]_ ;
  assign n2270 = \new_[2162]_  ? \new_[7597]_  : \new_[2685]_ ;
  assign n2470 = \new_[2202]_  ? \new_[7470]_  : \new_[2686]_ ;
  assign n2455 = \new_[2199]_  ? \new_[7597]_  : \new_[2687]_ ;
  assign n2460 = \new_[2200]_  ? \new_[7470]_  : \new_[2688]_ ;
  assign n2465 = \new_[2201]_  ? \new_[7597]_  : \new_[2689]_ ;
  assign n2475 = \new_[2203]_  ? \new_[7470]_  : \new_[2690]_ ;
  assign n2285 = ~\new_[2578]_  | (~\new_[3897]_  & ~\new_[8960]_ );
  assign n2290 = ~\new_[2579]_  | (~\new_[3898]_  & ~\new_[8957]_ );
  assign n2295 = ~\new_[2580]_  | (~\new_[3899]_  & ~\new_[8958]_ );
  assign n2315 = ~\new_[2581]_  | (~\new_[3900]_  & ~\new_[8955]_ );
  assign n2310 = ~\new_[2583]_  | (~\new_[3902]_  & ~\new_[8956]_ );
  assign n2300 = ~\new_[2582]_  | (~\new_[3901]_  & ~\new_[8956]_ );
  assign n2305 = ~\new_[2584]_  | (~\new_[3903]_  & ~\new_[8957]_ );
  assign n2485 = ~\new_[2585]_  | (~\new_[3904]_  & ~\new_[8961]_ );
  assign n2480 = ~\new_[2586]_  | (~\new_[3905]_  & ~\new_[8961]_ );
  assign n2320 = ~\new_[2587]_  | (~\new_[3906]_  & ~\new_[8958]_ );
  assign n2325 = ~\new_[2588]_  | (~\new_[3907]_  & ~\new_[8961]_ );
  assign n2340 = ~\new_[2589]_  | (~\new_[3908]_  & ~\new_[8958]_ );
  assign n2335 = ~\new_[2590]_  | (~\new_[3909]_  & ~\new_[8958]_ );
  assign n2345 = ~\new_[2591]_  | (~\new_[3911]_  & ~\new_[8956]_ );
  assign n2330 = ~\new_[2595]_  | (~\new_[3910]_  & ~\new_[8958]_ );
  assign n2350 = ~\new_[2592]_  | (~\new_[3912]_  & ~\new_[8958]_ );
  assign n2355 = ~\new_[2593]_  | (~\new_[3913]_  & ~\new_[8961]_ );
  assign n2375 = ~\new_[2599]_  | (~\new_[3915]_  & ~\new_[8958]_ );
  assign n2360 = ~\new_[2594]_  | (~\new_[3914]_  & ~\new_[8961]_ );
  assign n2370 = ~\new_[2597]_  | (~\new_[3916]_  & ~\new_[8961]_ );
  assign n2365 = ~\new_[2596]_  | (~\new_[3917]_  & ~\new_[8961]_ );
  assign n2380 = ~\new_[2598]_  | (~\new_[3918]_  & ~\new_[8961]_ );
  assign n2385 = ~\new_[2600]_  | (~\new_[3919]_  & ~\new_[8961]_ );
  assign n2390 = ~\new_[2601]_  | (~\new_[3920]_  & ~\new_[8958]_ );
  assign n2400 = ~\new_[2603]_  | (~\new_[3921]_  & ~\new_[8961]_ );
  assign n2395 = ~\new_[2602]_  | (~\new_[3922]_  & ~\new_[8958]_ );
  assign n2275 = ~\new_[2604]_  | (~\new_[3923]_  & ~\new_[8958]_ );
  assign n2280 = ~\new_[2605]_  | (~\new_[3924]_  & ~\new_[8961]_ );
  assign n2405 = ~\new_[2606]_  | (~\new_[3925]_  & ~\new_[8961]_ );
  assign n2420 = ~\new_[2609]_  | (~\new_[3926]_  & ~\new_[8955]_ );
  assign n2410 = ~\new_[2607]_  | (~\new_[3927]_  & ~\new_[8958]_ );
  assign n2415 = ~\new_[2608]_  | (~\new_[3928]_  & ~\new_[8958]_ );
  assign n2425 = ~\new_[2610]_  | (~\new_[3929]_  & ~\new_[8961]_ );
  assign n2435 = ~\new_[2612]_  | (~\new_[3930]_  & ~\new_[8958]_ );
  assign n2430 = ~\new_[2611]_  | (~\new_[3931]_  & ~\new_[8958]_ );
  assign \new_[2411]_  = \\ks1_key_reg_reg[113] ;
  assign n2730 = ~\new_[4446]_  | ~\new_[5143]_  | ~\new_[2803]_ ;
  assign \new_[2413]_  = ~\\mix1_data_reg_reg[36] ;
  assign \new_[2414]_  = ~\\mix1_data_reg_reg[44] ;
  assign \new_[2415]_  = ~\\mix1_data_reg_reg[60] ;
  assign \new_[2416]_  = ~\\mix1_data_reg_reg[68] ;
  assign \new_[2417]_  = ~\\mix1_data_reg_reg[52] ;
  assign \new_[2418]_  = ~\\mix1_data_reg_reg[84] ;
  assign \new_[2419]_  = ~\\mix1_data_reg_reg[76] ;
  assign \new_[2420]_  = ~\\mix1_data_reg_reg[92] ;
  assign \new_[2421]_  = \\ks1_key_reg_reg[112] ;
  assign \new_[2422]_  = \\ks1_key_reg_reg[115] ;
  assign \new_[2423]_  = \\ks1_key_reg_reg[116] ;
  assign \new_[2424]_  = \\ks1_key_reg_reg[114] ;
  assign \new_[2425]_  = \\ks1_key_reg_reg[118] ;
  assign \new_[2426]_  = addroundkey_ready_o_reg;
  assign \new_[2427]_  = ~\new_[2804]_  | ~\new_[2661]_ ;
  assign n2515 = ~\new_[2662]_  | ~\new_[7240]_ ;
  assign n2520 = ~\new_[8464]_  | ~\new_[7171]_ ;
  assign n2525 = ~\new_[8474]_  | ~\new_[7184]_ ;
  assign n2530 = ~\new_[8459]_  | ~\new_[7226]_ ;
  assign \new_[2432]_  = \new_[3373]_  ^ \new_[2830]_ ;
  assign \new_[2433]_  = \new_[3101]_  ^ \new_[2831]_ ;
  assign n2715 = \new_[2264]_  ? \new_[7597]_  : \new_[2827]_ ;
  assign n2720 = \new_[2265]_  ? \new_[7597]_  : \new_[2830]_ ;
  assign n2760 = \new_[2273]_  ? \new_[7470]_  : \new_[2831]_ ;
  assign n2750 = \new_[2271]_  ? \new_[7597]_  : \new_[2828]_ ;
  assign n2725 = \new_[2266]_  ? \new_[7470]_  : \new_[2829]_ ;
  assign \new_[2439]_  = \new_[3348]_  ^ \new_[2828]_ ;
  assign \new_[2440]_  = \new_[3349]_  ^ \new_[2829]_ ;
  assign \new_[2441]_  = \new_[3372]_  ^ \new_[2827]_ ;
  assign \new_[2442]_  = ~\new_[2558]_ ;
  assign n2540 = ~\new_[2697]_  | (~\new_[4010]_  & ~\new_[8957]_ );
  assign n2800 = ~\new_[2693]_  | (~\new_[4009]_  & ~\new_[8960]_ );
  assign n2545 = ~\new_[2694]_  | (~\new_[4011]_  & ~\new_[8958]_ );
  assign n2535 = ~\new_[2708]_  | (~\new_[4012]_  & ~\new_[8956]_ );
  assign n2550 = ~\new_[2696]_  | (~\new_[4013]_  & ~\new_[8958]_ );
  assign n2560 = ~\new_[2698]_  | (~\new_[4014]_  & ~\new_[8956]_ );
  assign n2555 = ~\new_[2700]_  | (~\new_[4015]_  & ~\new_[8957]_ );
  assign n2565 = ~\new_[2699]_  | (~\new_[4017]_  & ~\new_[8957]_ );
  assign n2795 = ~\new_[2701]_  | (~\new_[4016]_  & ~\new_[8958]_ );
  assign n2570 = ~\new_[2703]_  | (~\new_[4019]_  & ~\new_[8960]_ );
  assign n2785 = ~\new_[2702]_  | (~\new_[4018]_  & ~\new_[8961]_ );
  assign n2575 = ~\new_[2704]_  | (~\new_[4020]_  & ~\new_[8961]_ );
  assign n2590 = ~\new_[2713]_  | (~\new_[4026]_  & ~\new_[8960]_ );
  assign n2765 = ~\new_[2711]_  | (~\new_[4023]_  & ~\new_[8958]_ );
  assign n2580 = ~\new_[2707]_  | (~\new_[4021]_  & ~\new_[8958]_ );
  assign n2585 = ~\new_[2706]_  | (~\new_[4022]_  & ~\new_[8961]_ );
  assign n2775 = ~\new_[2709]_  | (~\new_[4024]_  & ~\new_[8955]_ );
  assign n2595 = ~\new_[2710]_  | (~\new_[4025]_  & ~\new_[8958]_ );
  assign \new_[2461]_  = \\ks1_key_reg_reg[117] ;
  assign n2600 = ~\new_[2712]_  | (~\new_[4027]_  & ~\new_[8956]_ );
  assign n2500 = ~\new_[2720]_  | (~\new_[4029]_  & ~\new_[8956]_ );
  assign n2605 = ~\new_[2715]_  | (~\new_[4028]_  & ~\new_[8961]_ );
  assign n2745 = ~\new_[2719]_  | (~\new_[4032]_  & ~\new_[8961]_ );
  assign n2610 = ~\new_[2714]_  | (~\new_[4030]_  & ~\new_[8961]_ );
  assign n2615 = ~\new_[2716]_  | (~\new_[4031]_  & ~\new_[8958]_ );
  assign n2755 = ~\new_[2717]_  | (~\new_[4033]_  & ~\new_[8958]_ );
  assign n2620 = ~\new_[2718]_  | (~\new_[4034]_  & ~\new_[8961]_ );
  assign n2635 = ~\new_[2721]_  | (~\new_[4035]_  & ~\new_[8957]_ );
  assign n2735 = ~\new_[2723]_  | (~\new_[4036]_  & ~\new_[8957]_ );
  assign n2625 = ~\new_[2722]_  | (~\new_[4037]_  & ~\new_[8961]_ );
  assign n2630 = ~\new_[2724]_  | (~\new_[4038]_  & ~\new_[8961]_ );
  assign n2640 = ~\new_[2725]_  | (~\new_[4039]_  & ~\new_[8961]_ );
  assign n2645 = ~\new_[2726]_  | (~\new_[4040]_  & ~\new_[8961]_ );
  assign n2655 = ~\new_[2729]_  | (~\new_[4042]_  & ~\new_[8960]_ );
  assign n2740 = ~\new_[2727]_  | (~\new_[4041]_  & ~\new_[8961]_ );
  assign n2650 = ~\new_[2728]_  | (~\new_[4043]_  & ~\new_[8961]_ );
  assign n2495 = ~\new_[2730]_  | (~\new_[4044]_  & ~\new_[8958]_ );
  assign n2510 = ~\new_[2732]_  | (~\new_[4045]_  & ~\new_[8958]_ );
  assign n2660 = ~\new_[2731]_  | (~\new_[4046]_  & ~\new_[8961]_ );
  assign n2670 = ~\new_[2735]_  | (~\new_[4048]_  & ~\new_[8960]_ );
  assign n2665 = ~\new_[2733]_  | (~\new_[4047]_  & ~\new_[8961]_ );
  assign n2505 = ~\new_[2734]_  | (~\new_[4049]_  & ~\new_[8960]_ );
  assign n2680 = ~\new_[2737]_  | (~\new_[4051]_  & ~\new_[8958]_ );
  assign n2675 = ~\new_[2736]_  | (~\new_[4050]_  & ~\new_[8958]_ );
  assign n2685 = ~\new_[2738]_  | (~\new_[4052]_  & ~\new_[8958]_ );
  assign n2690 = ~\new_[2739]_  | (~\new_[4053]_  & ~\new_[8956]_ );
  assign n2820 = ~\new_[2695]_  | (~\new_[4054]_  & ~\new_[8961]_ );
  assign n2695 = ~\new_[2740]_  | (~\new_[4055]_  & ~\new_[8958]_ );
  assign n2810 = ~\new_[2741]_  | (~\new_[4056]_  & ~\new_[8958]_ );
  assign n2805 = ~\new_[2742]_  | (~\new_[4057]_  & ~\new_[8958]_ );
  assign n2700 = ~\new_[2743]_  | (~\new_[4058]_  & ~\new_[8956]_ );
  assign n2790 = ~\new_[2744]_  | (~\new_[4059]_  & ~\new_[8956]_ );
  assign n2490 = ~\new_[2705]_  | (~\new_[4063]_  & ~\new_[8961]_ );
  assign n2770 = ~\new_[2745]_  | (~\new_[4060]_  & ~\new_[8958]_ );
  assign n2705 = ~\new_[2746]_  | (~\new_[4061]_  & ~\new_[8957]_ );
  assign n2780 = ~\new_[2747]_  | (~\new_[4062]_  & ~\new_[8961]_ );
  assign n2710 = ~\new_[2748]_  | (~\new_[4064]_  & ~\new_[8960]_ );
  assign n2815 = ~\new_[2692]_  | (~\new_[4065]_  & ~\new_[8960]_ );
  assign \new_[2501]_  = ~\new_[2614]_  | ~\new_[8955]_ ;
  assign \new_[2502]_  = ~\new_[2615]_  | ~\new_[8955]_ ;
  assign \new_[2503]_  = ~\new_[2616]_  | ~\new_[8955]_ ;
  assign \new_[2504]_  = ~\new_[2623]_  | ~\new_[8955]_ ;
  assign \new_[2505]_  = ~\new_[2622]_  | ~\new_[8955]_ ;
  assign \new_[2506]_  = ~\new_[2613]_  | ~\new_[8958]_ ;
  assign \new_[2507]_  = ~\new_[2625]_  | ~\new_[8956]_ ;
  assign \new_[2508]_  = ~\new_[2624]_  | ~\new_[8960]_ ;
  assign \new_[2509]_  = ~\new_[2691]_  | ~\new_[8956]_ ;
  assign \new_[2510]_  = ~\new_[2629]_  | ~\new_[8956]_ ;
  assign \new_[2511]_  = ~\new_[2631]_  | ~\new_[8956]_ ;
  assign \new_[2512]_  = ~\new_[2632]_  | ~\new_[8958]_ ;
  assign \new_[2513]_  = ~\new_[2634]_  | ~\new_[8958]_ ;
  assign \new_[2514]_  = ~\new_[2635]_  | ~\new_[8956]_ ;
  assign \new_[2515]_  = ~\new_[2633]_  | ~\new_[8957]_ ;
  assign \new_[2516]_  = ~\new_[2637]_  | ~\new_[8955]_ ;
  assign \new_[2517]_  = ~\new_[2636]_  | ~\new_[8956]_ ;
  assign \new_[2518]_  = ~\new_[2638]_  | ~\new_[8955]_ ;
  assign \new_[2519]_  = ~\new_[2640]_  | ~\new_[8955]_ ;
  assign \new_[2520]_  = ~\new_[2641]_  | ~\new_[8955]_ ;
  assign \new_[2521]_  = ~\new_[2642]_  | ~\new_[8955]_ ;
  assign \new_[2522]_  = ~\new_[2643]_  | ~\new_[8955]_ ;
  assign \new_[2523]_  = ~\new_[2645]_  | ~\new_[8955]_ ;
  assign \new_[2524]_  = ~\new_[2646]_  | ~\new_[8960]_ ;
  assign \new_[2525]_  = ~\new_[2639]_  | ~\new_[8960]_ ;
  assign \new_[2526]_  = ~\new_[2644]_  | ~\new_[8956]_ ;
  assign \new_[2527]_  = ~\new_[2647]_  | ~\new_[8956]_ ;
  assign \new_[2528]_  = ~\new_[2648]_  | ~\new_[8958]_ ;
  assign \new_[2529]_  = ~\new_[2649]_  | ~\new_[8955]_ ;
  assign \new_[2530]_  = ~\new_[2652]_  | ~\new_[8955]_ ;
  assign \new_[2531]_  = ~\new_[2650]_  | ~\new_[8958]_ ;
  assign \new_[2532]_  = ~\new_[2654]_  | ~\new_[8955]_ ;
  assign \new_[2533]_  = ~\new_[2651]_  | ~\new_[8955]_ ;
  assign \new_[2534]_  = ~\new_[2655]_  | ~\new_[8955]_ ;
  assign \new_[2535]_  = ~\new_[2656]_  | ~\new_[8955]_ ;
  assign \new_[2536]_  = ~\new_[2657]_  | ~\new_[8958]_ ;
  assign \new_[2537]_  = \\ks1_key_reg_reg[99] ;
  assign \new_[2538]_  = ~\\mix1_data_reg_reg[105] ;
  assign \new_[2539]_  = ~\\mix1_data_reg_reg[106] ;
  assign \new_[2540]_  = ~\\mix1_data_reg_reg[113] ;
  assign \new_[2541]_  = ~\\mix1_data_reg_reg[114] ;
  assign \new_[2542]_  = ~\\mix1_data_reg_reg[121] ;
  assign \new_[2543]_  = ~\\mix1_data_reg_reg[122] ;
  assign \new_[2544]_  = ~\\mix1_data_reg_reg[35] ;
  assign \new_[2545]_  = ~\\mix1_data_reg_reg[43] ;
  assign \new_[2546]_  = ~\\mix1_data_reg_reg[51] ;
  assign \new_[2547]_  = ~\\mix1_data_reg_reg[59] ;
  assign \new_[2548]_  = ~\\mix1_data_reg_reg[67] ;
  assign \new_[2549]_  = ~\\mix1_data_reg_reg[75] ;
  assign \new_[2550]_  = ~\\mix1_data_reg_reg[97] ;
  assign \new_[2551]_  = ~\\mix1_data_reg_reg[98] ;
  assign \new_[2552]_  = ~\\mix1_data_reg_reg[91] ;
  assign n2830 = ~\new_[8435]_  | ~\new_[7238]_ ;
  assign n2835 = ~\new_[2806]_  | ~\new_[7342]_ ;
  assign n2880 = ~\new_[8708]_  | ~\new_[7399]_ ;
  assign n2840 = ~\new_[2809]_  | ~\new_[7195]_ ;
  assign \new_[2557]_  = ~\new_[3003]_  | ~\new_[8724]_ ;
  assign \new_[2558]_  = ~\new_[2666]_ ;
  assign \new_[2559]_  = \new_[2933]_  ^ \new_[3517]_ ;
  assign n2845 = \new_[2348]_  ? \new_[7470]_  : \new_[2942]_ ;
  assign n2825 = \new_[2344]_  ? \new_[7597]_  : \new_[2950]_ ;
  assign n2850 = \new_[2349]_  ? \new_[7470]_  : \new_[2951]_ ;
  assign n2855 = \new_[2350]_  ? \new_[7470]_  : \new_[2944]_ ;
  assign n2860 = \new_[2351]_  ? \new_[7470]_  : \new_[2945]_ ;
  assign n2865 = \new_[2352]_  ? \new_[7597]_  : \new_[2946]_ ;
  assign n2870 = \new_[2353]_  ? \new_[7470]_  : \new_[2947]_ ;
  assign n2875 = \new_[2354]_  ? \new_[7470]_  : \new_[2949]_ ;
  assign \new_[2568]_  = ~\new_[2833]_  | (~\new_[3060]_  & ~\new_[3319]_ );
  assign \new_[2569]_  = \new_[2944]_  ^ \new_[3074]_ ;
  assign \new_[2570]_  = \new_[2945]_  ^ \new_[3322]_ ;
  assign \new_[2571]_  = \new_[2946]_  ^ \new_[3323]_ ;
  assign \new_[2572]_  = \new_[2947]_  ^ \new_[3324]_ ;
  assign \new_[2573]_  = \new_[3360]_  ^ \new_[2942]_ ;
  assign \new_[2574]_  = \new_[3367]_  ^ \new_[2950]_ ;
  assign \new_[2575]_  = \new_[3371]_  ^ \new_[2949]_ ;
  assign \new_[2576]_  = \new_[3380]_  ^ \new_[2951]_ ;
  assign \new_[2577]_  = ~\\mix1_data_reg_reg[83] ;
  assign \new_[2578]_  = ~\new_[2749]_  | ~\new_[8955]_ ;
  assign \new_[2579]_  = ~\new_[2750]_  | ~\new_[8955]_ ;
  assign \new_[2580]_  = ~\new_[2751]_  | ~\new_[8960]_ ;
  assign \new_[2581]_  = ~\new_[2752]_  | ~\new_[8955]_ ;
  assign \new_[2582]_  = ~\new_[2754]_  | ~\new_[8960]_ ;
  assign \new_[2583]_  = ~\new_[2805]_  | ~\new_[8955]_ ;
  assign \new_[2584]_  = ~\new_[2802]_  | ~\new_[8960]_ ;
  assign \new_[2585]_  = ~\new_[2753]_  | ~\new_[8960]_ ;
  assign \new_[2586]_  = ~\new_[2760]_  | ~\new_[8955]_ ;
  assign \new_[2587]_  = ~\new_[2759]_  | ~\new_[8956]_ ;
  assign \new_[2588]_  = ~\new_[2777]_  | ~\new_[8955]_ ;
  assign \new_[2589]_  = ~\new_[2778]_  | ~\new_[8956]_ ;
  assign \new_[2590]_  = ~\new_[2779]_  | ~\new_[8958]_ ;
  assign \new_[2591]_  = ~\new_[2780]_  | ~\new_[8955]_ ;
  assign \new_[2592]_  = ~\new_[2781]_  | ~\new_[8956]_ ;
  assign \new_[2593]_  = ~\new_[2782]_  | ~\new_[8955]_ ;
  assign \new_[2594]_  = ~\new_[2783]_  | ~\new_[8955]_ ;
  assign \new_[2595]_  = ~\new_[2784]_  | ~\new_[8956]_ ;
  assign \new_[2596]_  = ~\new_[2788]_  | ~\new_[8955]_ ;
  assign \new_[2597]_  = ~\new_[2785]_  | ~\new_[8955]_ ;
  assign \new_[2598]_  = ~\new_[2787]_  | ~\new_[8958]_ ;
  assign \new_[2599]_  = ~\new_[2786]_  | ~\new_[8956]_ ;
  assign \new_[2600]_  = ~\new_[2789]_  | ~\new_[8956]_ ;
  assign \new_[2601]_  = ~\new_[2790]_  | ~\new_[8956]_ ;
  assign \new_[2602]_  = ~\new_[2791]_  | ~\new_[8955]_ ;
  assign \new_[2603]_  = ~\new_[2792]_  | ~\new_[8955]_ ;
  assign \new_[2604]_  = ~\new_[2793]_  | ~\new_[8956]_ ;
  assign \new_[2605]_  = ~\new_[2794]_  | ~\new_[8955]_ ;
  assign \new_[2606]_  = ~\new_[2795]_  | ~\new_[8955]_ ;
  assign \new_[2607]_  = ~\new_[2796]_  | ~\new_[8955]_ ;
  assign \new_[2608]_  = ~\new_[2797]_  | ~\new_[8955]_ ;
  assign \new_[2609]_  = ~\new_[2798]_  | ~\new_[8958]_ ;
  assign \new_[2610]_  = ~\new_[2799]_  | ~\new_[8956]_ ;
  assign \new_[2611]_  = ~\new_[2800]_  | ~\new_[8955]_ ;
  assign \new_[2612]_  = ~\new_[2801]_  | ~\new_[8958]_ ;
  assign \new_[2613]_  = ~\new_[3150]_  | (~\new_[3009]_  & ~\new_[4798]_ );
  assign \new_[2614]_  = ~\new_[3118]_  | (~\new_[3004]_  & ~\new_[4798]_ );
  assign \new_[2615]_  = ~\new_[3120]_  | (~\new_[3005]_  & ~\new_[4798]_ );
  assign \new_[2616]_  = ~\new_[3135]_  | (~\new_[3006]_  & ~\new_[4798]_ );
  assign \new_[2617]_  = ~\\mix1_data_reg_reg[120] ;
  assign \new_[2618]_  = ~\\mix1_data_reg_reg[117] ;
  assign \new_[2619]_  = ~\\mix1_data_reg_reg[125] ;
  assign \new_[2620]_  = ~\\mix1_data_reg_reg[118] ;
  assign n2955 = ~\new_[8955]_  | (~\new_[7269]_  & ~\new_[4797]_ );
  assign \new_[2622]_  = ~\new_[3147]_  | (~\new_[3008]_  & ~\new_[4798]_ );
  assign \new_[2623]_  = ~\new_[3146]_  | (~\new_[3007]_  & ~\new_[4798]_ );
  assign \new_[2624]_  = ~\new_[3152]_  | (~\new_[3011]_  & ~\new_[4798]_ );
  assign \new_[2625]_  = ~\new_[3151]_  | (~\new_[3010]_  & ~\new_[4798]_ );
  assign \new_[2626]_  = ~\\mix1_data_reg_reg[104] ;
  assign \new_[2627]_  = ~\\mix1_data_reg_reg[112] ;
  assign \new_[2628]_  = ~\\mix1_data_reg_reg[96] ;
  assign \new_[2629]_  = ~\new_[3160]_  | (~\new_[3013]_  & ~\new_[4798]_ );
  assign \new_[2630]_  = ~\\mix1_data_reg_reg[126] ;
  assign \new_[2631]_  = ~\new_[3170]_  | (~\new_[3014]_  & ~\new_[4798]_ );
  assign \new_[2632]_  = ~\new_[3115]_  | (~\new_[3016]_  & ~\new_[4798]_ );
  assign \new_[2633]_  = ~\new_[3204]_  | (~\new_[3015]_  & ~\new_[4798]_ );
  assign \new_[2634]_  = ~\new_[3202]_  | (~\new_[3018]_  & ~\new_[4798]_ );
  assign \new_[2635]_  = ~\new_[3205]_  | (~\new_[3017]_  & ~\new_[4798]_ );
  assign \new_[2636]_  = ~\new_[3208]_  | (~\new_[3019]_  & ~\new_[4798]_ );
  assign \new_[2637]_  = ~\new_[3209]_  | (~\new_[3020]_  & ~\new_[3675]_ );
  assign \new_[2638]_  = ~\new_[3211]_  | (~\new_[3021]_  & ~\new_[3675]_ );
  assign \new_[2639]_  = ~\new_[3221]_  | (~\new_[3022]_  & ~\new_[4798]_ );
  assign \new_[2640]_  = ~\new_[3214]_  | (~\new_[3023]_  & ~\new_[4798]_ );
  assign \new_[2641]_  = ~\new_[3216]_  | (~\new_[3024]_  & ~\new_[4798]_ );
  assign \new_[2642]_  = ~\new_[3217]_  | (~\new_[3025]_  & ~\new_[4798]_ );
  assign \new_[2643]_  = ~\new_[3219]_  | (~\new_[3026]_  & ~\new_[4798]_ );
  assign \new_[2644]_  = ~\new_[3212]_  | (~\new_[3029]_  & ~\new_[4798]_ );
  assign \new_[2645]_  = ~\new_[3213]_  | (~\new_[3027]_  & ~\new_[4798]_ );
  assign \new_[2646]_  = ~\new_[3220]_  | (~\new_[3028]_  & ~\new_[4798]_ );
  assign \new_[2647]_  = ~\new_[3226]_  | (~\new_[3030]_  & ~\new_[4798]_ );
  assign \new_[2648]_  = ~\new_[3234]_  | (~\new_[3032]_  & ~\new_[3675]_ );
  assign \new_[2649]_  = ~\new_[3239]_  | (~\new_[3033]_  & ~\new_[4798]_ );
  assign \new_[2650]_  = ~\new_[3243]_  | (~\new_[3034]_  & ~\new_[4798]_ );
  assign \new_[2651]_  = ~\new_[3229]_  | (~\new_[3031]_  & ~\new_[4798]_ );
  assign \new_[2652]_  = ~\new_[3246]_  | (~\new_[3036]_  & ~\new_[4798]_ );
  assign \new_[2653]_  = ~\\mix1_data_reg_reg[110] ;
  assign \new_[2654]_  = ~\new_[3244]_  | (~\new_[3035]_  & ~\new_[4798]_ );
  assign \new_[2655]_  = ~\new_[3247]_  | (~\new_[3037]_  & ~\new_[4798]_ );
  assign \new_[2656]_  = ~\new_[3248]_  | (~\new_[3038]_  & ~\new_[4798]_ );
  assign \new_[2657]_  = ~\new_[3250]_  | (~\new_[3039]_  & ~\new_[4798]_ );
  assign \new_[2658]_  = ~\\mix1_data_reg_reg[102] ;
  assign \new_[2659]_  = ~\\mix1_data_reg_reg[109] ;
  assign \new_[2660]_  = ~\\mix1_data_reg_reg[101] ;
  assign \new_[2661]_  = ~\new_[2923]_  | ~\new_[3291]_ ;
  assign \new_[2662]_  = (~\new_[3073]_  | ~\new_[8713]_ ) & (~\new_[7960]_  | ~\new_[8716]_ );
  assign \new_[2663]_  = ~\new_[3293]_  | ~\new_[8724]_ ;
  assign \new_[2664]_  = ~\new_[3292]_  | ~\new_[8373]_ ;
  assign \new_[2665]_  = ~\new_[3291]_  | ~\new_[8373]_ ;
  assign \new_[2666]_  = ~\new_[8388]_ ;
  assign n2890 = ~\new_[2937]_  | ~\new_[7255]_ ;
  assign n2895 = ~\new_[2938]_  | ~\new_[7285]_ ;
  assign n2910 = ~\new_[2939]_  | ~\new_[7288]_ ;
  assign n2900 = ~\new_[2940]_  | ~\new_[7345]_ ;
  assign n2905 = ~\new_[2941]_  | ~\new_[7340]_ ;
  assign n2920 = ~\new_[2943]_  | ~\new_[7360]_ ;
  assign n2915 = ~\new_[2948]_  | ~\new_[7337]_ ;
  assign n2925 = ~\new_[2952]_  | ~\new_[7328]_ ;
  assign \new_[2675]_  = \new_[3044]_  ^ \new_[3518]_ ;
  assign \new_[2676]_  = \new_[3045]_  ^ \new_[3308]_ ;
  assign n2885 = \new_[2411]_  ? \new_[7597]_  : \new_[3061]_ ;
  assign n2930 = \new_[2421]_  ? \new_[7470]_  : \new_[3064]_ ;
  assign n2945 = \new_[2424]_  ? \new_[7470]_  : \new_[3065]_ ;
  assign n2940 = \new_[2423]_  ? \new_[8843]_  : \new_[3067]_ ;
  assign n2960 = \new_[2461]_  ? \new_[7597]_  : \new_[3063]_ ;
  assign n2950 = \new_[2425]_  ? \new_[7597]_  : \new_[3068]_ ;
  assign n2935 = \new_[2422]_  ? \new_[8843]_  : \new_[3069]_ ;
  assign \new_[2684]_  = \new_[3362]_  ^ \new_[3064]_ ;
  assign \new_[2685]_  = \new_[3363]_  ^ \new_[3061]_ ;
  assign \new_[2686]_  = \new_[3364]_  ^ \new_[3065]_ ;
  assign \new_[2687]_  = \new_[3365]_  ^ \new_[3069]_ ;
  assign \new_[2688]_  = \new_[3368]_  ^ \new_[3067]_ ;
  assign \new_[2689]_  = \new_[3369]_  ^ \new_[3063]_ ;
  assign \new_[2690]_  = \new_[3370]_  ^ \new_[3068]_ ;
  assign \new_[2691]_  = ~\new_[3153]_  | (~\new_[3012]_  & ~\new_[4798]_ );
  assign \new_[2692]_  = ~\new_[2843]_  | ~\new_[8957]_ ;
  assign \new_[2693]_  = ~\new_[2845]_  | ~\new_[8955]_ ;
  assign \new_[2694]_  = ~\new_[2846]_  | ~\new_[8956]_ ;
  assign \new_[2695]_  = ~\new_[2909]_  | ~\new_[8960]_ ;
  assign \new_[2696]_  = ~\new_[2847]_  | ~\new_[8956]_ ;
  assign \new_[2697]_  = ~\new_[2848]_  | ~\new_[8955]_ ;
  assign \new_[2698]_  = ~\new_[2849]_  | ~\new_[8955]_ ;
  assign \new_[2699]_  = ~\new_[2850]_  | ~\new_[8958]_ ;
  assign \new_[2700]_  = ~\new_[2851]_  | ~\new_[8958]_ ;
  assign \new_[2701]_  = ~\new_[2856]_  | ~\new_[8960]_ ;
  assign \new_[2702]_  = ~\new_[2853]_  | ~\new_[8957]_ ;
  assign \new_[2703]_  = ~\new_[2854]_  | ~\new_[8957]_ ;
  assign \new_[2704]_  = ~\new_[2855]_  | ~\new_[8960]_ ;
  assign \new_[2705]_  = ~\new_[2844]_  | ~\new_[8955]_ ;
  assign \new_[2706]_  = ~\new_[2857]_  | ~\new_[8955]_ ;
  assign \new_[2707]_  = ~\new_[2858]_  | ~\new_[8958]_ ;
  assign \new_[2708]_  = ~\new_[2859]_  | ~\new_[8955]_ ;
  assign \new_[2709]_  = ~\new_[2860]_  | ~\new_[8955]_ ;
  assign \new_[2710]_  = ~\new_[2863]_  | ~\new_[8958]_ ;
  assign \new_[2711]_  = ~\new_[2865]_  | ~\new_[8958]_ ;
  assign \new_[2712]_  = ~\new_[2871]_  | ~\new_[8958]_ ;
  assign \new_[2713]_  = ~\new_[2925]_  | ~\new_[8960]_ ;
  assign \new_[2714]_  = ~\new_[2875]_  | ~\new_[8956]_ ;
  assign \new_[2715]_  = ~\new_[2924]_  | ~\new_[8956]_ ;
  assign \new_[2716]_  = ~\new_[2852]_  | ~\new_[8955]_ ;
  assign \new_[2717]_  = ~\new_[2886]_  | ~\new_[8956]_ ;
  assign \new_[2718]_  = ~\new_[2888]_  | ~\new_[8955]_ ;
  assign \new_[2719]_  = ~\new_[2887]_  | ~\new_[8955]_ ;
  assign \new_[2720]_  = ~\new_[2892]_  | ~\new_[8955]_ ;
  assign \new_[2721]_  = ~\new_[2889]_  | ~\new_[8955]_ ;
  assign \new_[2722]_  = ~\new_[2890]_  | ~\new_[8955]_ ;
  assign \new_[2723]_  = ~\new_[2893]_  | ~\new_[8955]_ ;
  assign \new_[2724]_  = ~\new_[2891]_  | ~\new_[8958]_ ;
  assign \new_[2725]_  = ~\new_[2894]_  | ~\new_[8958]_ ;
  assign \new_[2726]_  = ~\new_[2895]_  | ~\new_[8960]_ ;
  assign \new_[2727]_  = ~\new_[2896]_  | ~\new_[8960]_ ;
  assign \new_[2728]_  = ~\new_[2897]_  | ~\new_[8956]_ ;
  assign \new_[2729]_  = ~\new_[2898]_  | ~\new_[8958]_ ;
  assign \new_[2730]_  = ~\new_[2899]_  | ~\new_[8958]_ ;
  assign \new_[2731]_  = ~\new_[2900]_  | ~\new_[8958]_ ;
  assign \new_[2732]_  = ~\new_[2901]_  | ~\new_[8956]_ ;
  assign \new_[2733]_  = ~\new_[2902]_  | ~\new_[8956]_ ;
  assign \new_[2734]_  = ~\new_[2904]_  | ~\new_[8955]_ ;
  assign \new_[2735]_  = ~\new_[2903]_  | ~\new_[8960]_ ;
  assign \new_[2736]_  = ~\new_[2905]_  | ~\new_[8956]_ ;
  assign \new_[2737]_  = ~\new_[2906]_  | ~\new_[8960]_ ;
  assign \new_[2738]_  = ~\new_[2907]_  | ~\new_[8956]_ ;
  assign \new_[2739]_  = ~\new_[2908]_  | ~\new_[8955]_ ;
  assign \new_[2740]_  = ~\new_[2910]_  | ~\new_[8955]_ ;
  assign \new_[2741]_  = ~\new_[2911]_  | ~\new_[8955]_ ;
  assign \new_[2742]_  = ~\new_[2912]_  | ~\new_[8955]_ ;
  assign \new_[2743]_  = ~\new_[2913]_  | ~\new_[8960]_ ;
  assign \new_[2744]_  = ~\new_[2914]_  | ~\new_[8958]_ ;
  assign \new_[2745]_  = ~\new_[2915]_  | ~\new_[8958]_ ;
  assign \new_[2746]_  = ~\new_[2916]_  | ~\new_[8955]_ ;
  assign \new_[2747]_  = ~\new_[2917]_  | ~\new_[8955]_ ;
  assign \new_[2748]_  = ~\new_[2918]_  | ~\new_[8958]_ ;
  assign \new_[2749]_  = ~\new_[3116]_  | (~\new_[3255]_  & ~\new_[4798]_ );
  assign \new_[2750]_  = ~\new_[3119]_  | (~\new_[3256]_  & ~\new_[4798]_ );
  assign \new_[2751]_  = ~\new_[3124]_  | (~\new_[3258]_  & ~\new_[4798]_ );
  assign \new_[2752]_  = ~\new_[3139]_  | (~\new_[3259]_  & ~\new_[4798]_ );
  assign \new_[2753]_  = ~\new_[3145]_  | (~\new_[3263]_  & ~\new_[4798]_ );
  assign \new_[2754]_  = ~\new_[3142]_  | (~\new_[3260]_  & ~\new_[3675]_ );
  assign \new_[2755]_  = \\mix1_data_o_reg_reg[12] ;
  assign \new_[2756]_  = \\mix1_data_o_reg_reg[20] ;
  assign \new_[2757]_  = \\mix1_data_o_reg_reg[28] ;
  assign \new_[2758]_  = \\mix1_data_o_reg_reg[4] ;
  assign \new_[2759]_  = ~\new_[3222]_  | (~\new_[3264]_  & ~\new_[4798]_ );
  assign \new_[2760]_  = ~\new_[3154]_  | (~\new_[3265]_  & ~\new_[3675]_ );
  assign \new_[2761]_  = ~\\mix1_data_reg_reg[33] ;
  assign \new_[2762]_  = ~\\mix1_data_reg_reg[34] ;
  assign \new_[2763]_  = ~\\mix1_data_reg_reg[42] ;
  assign \new_[2764]_  = ~\\mix1_data_reg_reg[41] ;
  assign \new_[2765]_  = ~\\mix1_data_reg_reg[49] ;
  assign \new_[2766]_  = ~\\mix1_data_reg_reg[50] ;
  assign \new_[2767]_  = ~\\mix1_data_reg_reg[57] ;
  assign \new_[2768]_  = ~\\mix1_data_reg_reg[58] ;
  assign \new_[2769]_  = ~\\mix1_data_reg_reg[65] ;
  assign \new_[2770]_  = ~\\mix1_data_reg_reg[66] ;
  assign \new_[2771]_  = ~\\mix1_data_reg_reg[74] ;
  assign \new_[2772]_  = ~\\mix1_data_reg_reg[73] ;
  assign \new_[2773]_  = ~\\mix1_data_reg_reg[81] ;
  assign \new_[2774]_  = ~\\mix1_data_reg_reg[82] ;
  assign \new_[2775]_  = ~\\mix1_data_reg_reg[89] ;
  assign \new_[2776]_  = ~\\mix1_data_reg_reg[90] ;
  assign \new_[2777]_  = ~\new_[3158]_  | (~\new_[3266]_  & ~\new_[4798]_ );
  assign \new_[2778]_  = ~\new_[3191]_  | (~\new_[3267]_  & ~\new_[4798]_ );
  assign \new_[2779]_  = ~\new_[3165]_  | (~\new_[3268]_  & ~\new_[4798]_ );
  assign \new_[2780]_  = ~\new_[3169]_  | (~\new_[3269]_  & ~\new_[4798]_ );
  assign \new_[2781]_  = ~\new_[3171]_  | (~\new_[3270]_  & ~\new_[4798]_ );
  assign \new_[2782]_  = ~\new_[3175]_  | (~\new_[3271]_  & ~\new_[4798]_ );
  assign \new_[2783]_  = ~\new_[3176]_  | (~\new_[3273]_  & ~\new_[4798]_ );
  assign \new_[2784]_  = ~\new_[3174]_  | (~\new_[3272]_  & ~\new_[4798]_ );
  assign \new_[2785]_  = ~\new_[3178]_  | (~\new_[3274]_  & ~\new_[4798]_ );
  assign \new_[2786]_  = ~\new_[3181]_  | (~\new_[3277]_  & ~\new_[4798]_ );
  assign \new_[2787]_  = ~\new_[3179]_  | (~\new_[3275]_  & ~\new_[4798]_ );
  assign \new_[2788]_  = ~\new_[3180]_  | (~\new_[3276]_  & ~\new_[4798]_ );
  assign \new_[2789]_  = ~\new_[3182]_  | (~\new_[3278]_  & ~\new_[4798]_ );
  assign \new_[2790]_  = ~\new_[3189]_  | (~\new_[3279]_  & ~\new_[3675]_ );
  assign \new_[2791]_  = ~\new_[3192]_  | (~\new_[3280]_  & ~\new_[4798]_ );
  assign \new_[2792]_  = ~\new_[3197]_  | (~\new_[3281]_  & ~\new_[4798]_ );
  assign \new_[2793]_  = ~\new_[3206]_  | (~\new_[3282]_  & ~\new_[4798]_ );
  assign \new_[2794]_  = ~\new_[3218]_  | (~\new_[3283]_  & ~\new_[4798]_ );
  assign \new_[2795]_  = ~\new_[3223]_  | (~\new_[3284]_  & ~\new_[4798]_ );
  assign \new_[2796]_  = ~\new_[3227]_  | (~\new_[3285]_  & ~\new_[4798]_ );
  assign \new_[2797]_  = ~\new_[3230]_  | (~\new_[3286]_  & ~\new_[4798]_ );
  assign \new_[2798]_  = ~\new_[3231]_  | (~\new_[3287]_  & ~\new_[4798]_ );
  assign \new_[2799]_  = ~\new_[3238]_  | (~\new_[3288]_  & ~\new_[4798]_ );
  assign \new_[2800]_  = ~\new_[3241]_  | (~\new_[3289]_  & ~\new_[4798]_ );
  assign \new_[2801]_  = ~\new_[3242]_  | (~\new_[3290]_  & ~\new_[4798]_ );
  assign \new_[2802]_  = ~\new_[3143]_  | (~\new_[3261]_  & ~\new_[4798]_ );
  assign \new_[2803]_  = \new_[5764]_  | \new_[8954]_ ;
  assign \new_[2804]_  = ~\new_[3003]_  | ~\new_[3040]_ ;
  assign \new_[2805]_  = ~\new_[3144]_  | (~\new_[3262]_  & ~\new_[4798]_ );
  assign \new_[2806]_  = (~\new_[3320]_  | ~\new_[8713]_ ) & (~\new_[8003]_  | ~\new_[8716]_ );
  assign \new_[2807]_  = ~\new_[3041]_  | ~\new_[3293]_ ;
  assign \new_[2808]_  = ~\new_[3292]_  | ~\new_[3042]_ ;
  assign \new_[2809]_  = (~\new_[3321]_  | ~\new_[8713]_ ) & (~\new_[8716]_  | ~\new_[8070]_ );
  assign \new_[2810]_  = ~\new_[3291]_ ;
  assign n2970 = ~\new_[3050]_  | ~\new_[7091]_ ;
  assign n2975 = ~\new_[3051]_  | ~\new_[7152]_ ;
  assign n2980 = ~\new_[3052]_  | ~\new_[7367]_ ;
  assign n2985 = ~\new_[3053]_  | ~\new_[7326]_ ;
  assign n2990 = ~\new_[3054]_  | ~\new_[7402]_ ;
  assign n2995 = ~\new_[8586]_  | ~\new_[7180]_ ;
  assign n3000 = ~\new_[3055]_  | ~\new_[7316]_ ;
  assign n3005 = ~\new_[3056]_  | ~\new_[7369]_ ;
  assign n3010 = ~\new_[3057]_  | ~\new_[7401]_ ;
  assign n3015 = ~\new_[3058]_  | ~\new_[7394]_ ;
  assign n3020 = ~\new_[3059]_  | ~\new_[7155]_ ;
  assign n3025 = ~\new_[3062]_  | ~\new_[7317]_ ;
  assign n3045 = ~\new_[3066]_  | ~\new_[7249]_ ;
  assign n3040 = ~\new_[3070]_  | ~\new_[7150]_ ;
  assign n3035 = ~\new_[3072]_  | ~\new_[7185]_ ;
  assign n3030 = ~\new_[3071]_  | ~\new_[7343]_ ;
  assign \new_[2827]_  = \new_[3630]_  ^ \new_[3305]_ ;
  assign \new_[2828]_  = \new_[3622]_  ^ \new_[3309]_ ;
  assign \new_[2829]_  = \new_[3623]_  ^ \new_[3310]_ ;
  assign \new_[2830]_  = \new_[3303]_  ^ \new_[3306]_ ;
  assign \new_[2831]_  = \new_[3302]_  ^ \new_[3307]_ ;
  assign n2965 = \new_[2537]_  ? \new_[7597]_  : \new_[3319]_ ;
  assign \new_[2833]_  = ~\new_[3060]_  | ~\new_[3319]_ ;
  assign \new_[2834]_  = ~\new_[3080]_  | (~\new_[4143]_  & ~\new_[6053]_ );
  assign \new_[2835]_  = ~\new_[3081]_  | (~\new_[4143]_  & ~\new_[6054]_ );
  assign n3075 = ~\new_[3111]_  | ~\new_[7197]_ ;
  assign n3050 = ~\new_[3112]_  | ~\new_[7257]_ ;
  assign n3080 = ~\new_[3113]_  | ~\new_[7243]_ ;
  assign \new_[2839]_  = (~\new_[4235]_  | ~\new_[8958]_ ) & (~\new_[6739]_  | ~\new_[8964]_ );
  assign \new_[2840]_  = (~\new_[3858]_  | ~\new_[8958]_ ) & (~\new_[6583]_  | ~\new_[8964]_ );
  assign \new_[2841]_  = (~\new_[4236]_  | ~\new_[8961]_ ) & (~\new_[6603]_  | ~\new_[8964]_ );
  assign \new_[2842]_  = ~\new_[2995]_ ;
  assign \new_[2843]_  = ~\new_[3117]_  | (~\new_[3411]_  & ~\new_[4798]_ );
  assign \new_[2844]_  = ~\new_[3114]_  | (~\new_[3413]_  & ~\new_[4798]_ );
  assign \new_[2845]_  = ~\new_[3121]_  | (~\new_[3412]_  & ~\new_[4798]_ );
  assign \new_[2846]_  = ~\new_[3122]_  | (~\new_[3414]_  & ~\new_[4798]_ );
  assign \new_[2847]_  = ~\new_[3123]_  | (~\new_[3415]_  & ~\new_[4798]_ );
  assign \new_[2848]_  = ~\new_[3125]_  | (~\new_[3416]_  & ~\new_[4798]_ );
  assign \new_[2849]_  = ~\new_[3126]_  | (~\new_[3417]_  & ~\new_[4798]_ );
  assign \new_[2850]_  = ~\new_[3128]_  | (~\new_[3418]_  & ~\new_[4798]_ );
  assign \new_[2851]_  = ~\new_[3129]_  | (~\new_[3419]_  & ~\new_[4798]_ );
  assign \new_[2852]_  = ~\new_[3157]_  | (~\new_[3434]_  & ~\new_[4798]_ );
  assign \new_[2853]_  = ~\new_[3130]_  | (~\new_[3420]_  & ~\new_[4798]_ );
  assign \new_[2854]_  = ~\new_[3132]_  | (~\new_[3422]_  & ~\new_[4798]_ );
  assign \new_[2855]_  = ~\new_[3131]_  | (~\new_[3421]_  & ~\new_[4798]_ );
  assign \new_[2856]_  = ~\new_[3133]_  | (~\new_[3423]_  & ~\new_[4798]_ );
  assign \new_[2857]_  = ~\new_[3136]_  | (~\new_[3425]_  & ~\new_[4798]_ );
  assign \new_[2858]_  = ~\new_[3137]_  | (~\new_[3426]_  & ~\new_[4798]_ );
  assign \new_[2859]_  = ~\new_[3134]_  | (~\new_[3424]_  & ~\new_[4798]_ );
  assign \new_[2860]_  = ~\new_[3138]_  | (~\new_[3427]_  & ~\new_[4798]_ );
  assign \new_[2861]_  = ~\\mix1_data_reg_reg[61] ;
  assign \new_[2862]_  = ~\\mix1_data_reg_reg[62] ;
  assign \new_[2863]_  = ~\new_[3140]_  | (~\new_[3428]_  & ~\new_[4798]_ );
  assign \new_[2864]_  = ~\\mix1_data_reg_reg[69] ;
  assign \new_[2865]_  = ~\new_[3141]_  | (~\new_[3429]_  & ~\new_[4798]_ );
  assign \new_[2866]_  = ~\\mix1_data_reg_reg[45] ;
  assign \new_[2867]_  = ~\\mix1_data_reg_reg[37] ;
  assign \new_[2868]_  = ~\\mix1_data_reg_reg[53] ;
  assign \new_[2869]_  = ~\\mix1_data_reg_reg[77] ;
  assign \new_[2870]_  = \\mix1_data_o_reg_reg[3] ;
  assign \new_[2871]_  = ~\new_[3148]_  | (~\new_[3431]_  & ~\new_[4798]_ );
  assign \new_[2872]_  = ~\\mix1_data_reg_reg[38] ;
  assign \new_[2873]_  = ~\\mix1_data_reg_reg[46] ;
  assign \new_[2874]_  = ~\\mix1_data_reg_reg[54] ;
  assign \new_[2875]_  = ~\new_[3156]_  | (~\new_[3433]_  & ~\new_[4798]_ );
  assign \new_[2876]_  = ~\\mix1_data_reg_reg[70] ;
  assign \new_[2877]_  = ~\\mix1_data_reg_reg[78] ;
  assign \new_[2878]_  = ~\\mix1_data_reg_reg[86] ;
  assign \new_[2879]_  = ~\\mix1_data_reg_reg[94] ;
  assign \new_[2880]_  = ~\\mix1_data_reg_reg[32] ;
  assign \new_[2881]_  = ~\\mix1_data_reg_reg[48] ;
  assign \new_[2882]_  = ~\\mix1_data_reg_reg[56] ;
  assign \new_[2883]_  = ~\\mix1_data_reg_reg[64] ;
  assign \new_[2884]_  = ~\\mix1_data_reg_reg[88] ;
  assign \new_[2885]_  = ~\\mix1_data_reg_reg[80] ;
  assign \new_[2886]_  = ~\new_[3159]_  | (~\new_[3435]_  & ~\new_[4798]_ );
  assign \new_[2887]_  = ~\new_[3155]_  | (~\new_[3438]_  & ~\new_[4798]_ );
  assign \new_[2888]_  = ~\new_[3161]_  | (~\new_[3436]_  & ~\new_[4798]_ );
  assign \new_[2889]_  = ~\new_[3183]_  | (~\new_[3439]_  & ~\new_[4798]_ );
  assign \new_[2890]_  = ~\new_[3163]_  | (~\new_[3440]_  & ~\new_[4798]_ );
  assign \new_[2891]_  = ~\new_[3127]_  | (~\new_[3441]_  & ~\new_[4798]_ );
  assign \new_[2892]_  = ~\new_[3162]_  | (~\new_[3437]_  & ~\new_[4798]_ );
  assign \new_[2893]_  = ~\new_[3166]_  | (~\new_[3444]_  & ~\new_[4798]_ );
  assign \new_[2894]_  = ~\new_[3164]_  | (~\new_[3442]_  & ~\new_[3675]_ );
  assign \new_[2895]_  = ~\new_[3167]_  | (~\new_[3445]_  & ~\new_[4798]_ );
  assign \new_[2896]_  = ~\new_[3168]_  | (~\new_[3446]_  & ~\new_[4798]_ );
  assign \new_[2897]_  = ~\new_[3172]_  | (~\new_[3447]_  & ~\new_[4798]_ );
  assign \new_[2898]_  = ~\new_[3173]_  | (~\new_[3448]_  & ~\new_[4798]_ );
  assign \new_[2899]_  = ~\new_[3177]_  | (~\new_[3449]_  & ~\new_[4798]_ );
  assign \new_[2900]_  = ~\new_[3184]_  | (~\new_[3450]_  & ~\new_[4798]_ );
  assign \new_[2901]_  = ~\new_[3185]_  | (~\new_[3451]_  & ~\new_[4798]_ );
  assign \new_[2902]_  = ~\new_[3186]_  | (~\new_[3452]_  & ~\new_[3675]_ );
  assign \new_[2903]_  = ~\new_[3188]_  | (~\new_[3454]_  & ~\new_[4798]_ );
  assign \new_[2904]_  = ~\new_[3187]_  | (~\new_[3453]_  & ~\new_[4798]_ );
  assign \new_[2905]_  = ~\new_[3190]_  | (~\new_[3455]_  & ~\new_[3675]_ );
  assign \new_[2906]_  = ~\new_[3194]_  | (~\new_[3456]_  & ~\new_[4798]_ );
  assign \new_[2907]_  = ~\new_[3196]_  | (~\new_[3457]_  & ~\new_[4798]_ );
  assign \new_[2908]_  = ~\new_[3199]_  | (~\new_[3458]_  & ~\new_[4798]_ );
  assign \new_[2909]_  = ~\new_[3224]_  | (~\new_[3459]_  & ~\new_[3675]_ );
  assign \new_[2910]_  = ~\new_[3225]_  | (~\new_[3460]_  & ~\new_[3675]_ );
  assign \new_[2911]_  = ~\new_[3228]_  | (~\new_[3461]_  & ~\new_[4798]_ );
  assign \new_[2912]_  = ~\new_[3232]_  | (~\new_[3463]_  & ~\new_[3675]_ );
  assign \new_[2913]_  = ~\new_[3233]_  | (~\new_[3462]_  & ~\new_[4798]_ );
  assign \new_[2914]_  = ~\new_[3236]_  | (~\new_[3464]_  & ~\new_[4798]_ );
  assign \new_[2915]_  = ~\new_[3237]_  | (~\new_[3465]_  & ~\new_[4798]_ );
  assign \new_[2916]_  = ~\new_[3240]_  | (~\new_[3466]_  & ~\new_[4798]_ );
  assign \new_[2917]_  = ~\new_[3245]_  | (~\new_[3467]_  & ~\new_[4798]_ );
  assign \new_[2918]_  = ~\new_[3249]_  | (~\new_[3468]_  & ~\new_[4798]_ );
  assign n3105 = ~\new_[3251]_  | ~\new_[7221]_ ;
  assign n3100 = ~\new_[3252]_  | ~\new_[7381]_ ;
  assign n3055 = ~\new_[3253]_  | ~\new_[7215]_ ;
  assign n3060 = ~\new_[3254]_  | ~\new_[7380]_ ;
  assign \new_[2923]_  = ~\new_[3003]_ ;
  assign \new_[2924]_  = ~\new_[3201]_  | (~\new_[3432]_  & ~\new_[4798]_ );
  assign \new_[2925]_  = ~\new_[3149]_  | (~\new_[3430]_  & ~\new_[4798]_ );
  assign \new_[2926]_  = ~\\mix1_data_reg_reg[72] ;
  assign n3095 = ~\new_[3315]_  | ~\new_[7158]_ ;
  assign n3090 = ~\new_[3316]_  | ~\new_[7165]_ ;
  assign n3065 = ~\new_[3317]_  | ~\new_[7307]_ ;
  assign n3085 = ~\new_[3318]_  | ~\new_[7325]_ ;
  assign \new_[2931]_  = ~\\mix1_data_reg_reg[40] ;
  assign \new_[2932]_  = \\mix1_data_o_reg_reg[27] ;
  assign \new_[2933]_  = \new_[3304]_  & \new_[3520]_ ;
  assign \new_[2934]_  = \\mix1_data_o_reg_reg[11] ;
  assign \new_[2935]_  = \\mix1_data_o_reg_reg[19] ;
  assign \new_[2936]_  = ~\\mix1_data_reg_reg[85] ;
  assign \new_[2937]_  = ~\new_[3090]_  & (~\new_[8114]_  | ~\new_[7645]_ );
  assign \new_[2938]_  = ~\new_[3091]_  & (~\new_[8093]_  | ~\new_[7645]_ );
  assign \new_[2939]_  = ~\new_[3092]_  & (~\new_[7945]_  | ~\new_[7645]_ );
  assign \new_[2940]_  = ~\new_[3093]_  & (~\new_[7981]_  | ~\new_[7645]_ );
  assign \new_[2941]_  = ~\new_[3094]_  & (~\new_[8032]_  | ~\new_[7499]_ );
  assign \new_[2942]_  = \new_[1343]_  ^ \new_[3350]_ ;
  assign \new_[2943]_  = ~\new_[3095]_  & (~\new_[8065]_  | ~\new_[7499]_ );
  assign \new_[2944]_  = \new_[1318]_  ^ \new_[3351]_ ;
  assign \new_[2945]_  = \new_[1236]_  ^ \new_[3352]_ ;
  assign \new_[2946]_  = \new_[1235]_  ^ \new_[3353]_ ;
  assign \new_[2947]_  = \new_[1382]_  ^ \new_[3354]_ ;
  assign \new_[2948]_  = ~\new_[3096]_  & (~\new_[8076]_  | ~\new_[7499]_ );
  assign \new_[2949]_  = \new_[1309]_  ^ \new_[3361]_ ;
  assign \new_[2950]_  = \new_[1761]_  ^ \new_[3366]_ ;
  assign \new_[2951]_  = \new_[1591]_  ^ \new_[3379]_ ;
  assign \new_[2952]_  = ~\new_[3097]_  & (~\new_[7977]_  | ~\new_[7499]_ );
  assign \new_[2953]_  = ~\\mix1_data_reg_reg[93] ;
  assign \new_[2954]_  = ~\new_[3075]_ ;
  assign \new_[2955]_  = ~\new_[3076]_ ;
  assign \new_[2956]_  = ~\new_[3325]_  & (~\new_[4332]_  | ~\new_[6062]_ );
  assign \new_[2957]_  = ~\new_[3077]_ ;
  assign \new_[2958]_  = ~\new_[3326]_  & (~\new_[4332]_  | ~\new_[6055]_ );
  assign \new_[2959]_  = ~\new_[3327]_  & (~\new_[4332]_  | ~\new_[6065]_ );
  assign \new_[2960]_  = ~\new_[3328]_  & (~\new_[4332]_  | ~\new_[6137]_ );
  assign \new_[2961]_  = ~\new_[3329]_  & (~\new_[4332]_  | ~\new_[6064]_ );
  assign \new_[2962]_  = ~\new_[3330]_  & (~\new_[4332]_  | ~\new_[6138]_ );
  assign \new_[2963]_  = ~\new_[3331]_  & (~\new_[4332]_  | ~\new_[6061]_ );
  assign \new_[2964]_  = ~\new_[3332]_  & (~\new_[4332]_  | ~\new_[6057]_ );
  assign \new_[2965]_  = ~\new_[3333]_  & (~\new_[4332]_  | ~\new_[6069]_ );
  assign \new_[2966]_  = ~\new_[3334]_  & (~\new_[4332]_  | ~\new_[6067]_ );
  assign \new_[2967]_  = ~\new_[3335]_  | (~\new_[4143]_  & ~\new_[6059]_ );
  assign \new_[2968]_  = ~\new_[3336]_  | (~\new_[4143]_  & ~\new_[6068]_ );
  assign \new_[2969]_  = ~\new_[3337]_  | (~\new_[4143]_  & ~\new_[6056]_ );
  assign \new_[2970]_  = ~\new_[3338]_  & (~\new_[4332]_  | ~\new_[6066]_ );
  assign \new_[2971]_  = ~\new_[3339]_  & (~\new_[4332]_  | ~\new_[6135]_ );
  assign \new_[2972]_  = ~\new_[4165]_  & ~\new_[8962]_ ;
  assign \new_[2973]_  = ~\new_[4149]_  & ~\new_[8954]_ ;
  assign \new_[2974]_  = ~\new_[4158]_  & ~\new_[8964]_ ;
  assign \new_[2975]_  = ~\new_[3966]_  & ~\new_[8954]_ ;
  assign n3070 = ~\new_[3110]_  | ~\new_[7163]_ ;
  assign n3130 = ~\new_[3390]_  | ~\new_[7186]_ ;
  assign n3135 = ~\new_[3391]_  | ~\new_[7283]_ ;
  assign n3145 = ~\new_[3392]_  | ~\new_[7376]_ ;
  assign n3140 = ~\new_[3393]_  | ~\new_[7309]_ ;
  assign n3150 = ~\new_[3394]_  | ~\new_[7157]_ ;
  assign n3155 = ~\new_[3395]_  | ~\new_[7388]_ ;
  assign n3160 = ~\new_[3396]_  | ~\new_[7164]_ ;
  assign n3165 = ~\new_[3397]_  | ~\new_[7358]_ ;
  assign n3170 = ~\new_[3398]_  | ~\new_[7191]_ ;
  assign n3175 = ~\new_[3399]_  | ~\new_[7242]_ ;
  assign n3185 = ~\new_[3400]_  | ~\new_[7211]_ ;
  assign n3180 = ~\new_[3401]_  | ~\new_[7324]_ ;
  assign n3190 = ~\new_[3402]_  | ~\new_[7225]_ ;
  assign n3195 = ~\new_[3403]_  | ~\new_[7108]_ ;
  assign n3200 = ~\new_[3404]_  | ~\new_[7154]_ ;
  assign n3205 = ~\new_[3405]_  | ~\new_[7212]_ ;
  assign \new_[2993]_  = (~\new_[3859]_  | ~\new_[8961]_ ) & (~\new_[6734]_  | ~\new_[8964]_ );
  assign \new_[2994]_  = (~\new_[3860]_  | ~\new_[8961]_ ) & (~\new_[6737]_  | ~\new_[8964]_ );
  assign \new_[2995]_  = (~\new_[3861]_  | ~\new_[8958]_ ) & (~\new_[6736]_  | ~\new_[8962]_ );
  assign \new_[2996]_  = ~\new_[3099]_ ;
  assign \new_[2997]_  = ~\new_[3100]_ ;
  assign \new_[2998]_  = ~\\mix1_data_reg_reg[103] ;
  assign \new_[2999]_  = ~\\mix1_data_reg_reg[111] ;
  assign \new_[3000]_  = ~\\mix1_data_reg_reg[127] ;
  assign \new_[3001]_  = ~\\mix1_data_reg_reg[119] ;
  assign \new_[3002]_  = ~\new_[3469]_  | ~\new_[8661]_ ;
  assign \new_[3003]_  = ~\new_[3506]_  | ~\new_[4320]_ ;
  assign \new_[3004]_  = ~\new_[3470]_  & (~\new_[5597]_  | ~\data_o[111] );
  assign \new_[3005]_  = ~\new_[3471]_  & (~\new_[5597]_  | ~\data_o[63] );
  assign \new_[3006]_  = ~\new_[3472]_  & (~\new_[5549]_  | ~\data_o[6] );
  assign \new_[3007]_  = ~\new_[3473]_  & (~\new_[5550]_  | ~\data_o[76] );
  assign \new_[3008]_  = ~\new_[3474]_  & (~\new_[5549]_  | ~\data_o[25] );
  assign \new_[3009]_  = ~\new_[3475]_  & (~\new_[5597]_  | ~\data_o[77] );
  assign \new_[3010]_  = ~\new_[3476]_  & (~\new_[5549]_  | ~\data_o[78] );
  assign \new_[3011]_  = ~\new_[3477]_  & (~\new_[5597]_  | ~\data_o[26] );
  assign \new_[3012]_  = ~\new_[3478]_  & (~\new_[5549]_  | ~\data_o[79] );
  assign \new_[3013]_  = ~\new_[3479]_  & (~\new_[5549]_  | ~\data_o[29] );
  assign \new_[3014]_  = ~\new_[3480]_  & (~\new_[5550]_  | ~\data_o[8] );
  assign \new_[3015]_  = ~\new_[3484]_  & (~\new_[5549]_  | ~\data_o[122] );
  assign \new_[3016]_  = ~\new_[3481]_  & (~\new_[5606]_  | ~\data_o[105] );
  assign \new_[3017]_  = ~\new_[3483]_  & (~\new_[5550]_  | ~\data_o[106] );
  assign \new_[3018]_  = ~\new_[3482]_  & (~\new_[5549]_  | ~\data_o[3] );
  assign \new_[3019]_  = ~\new_[3485]_  & (~\new_[5597]_  | ~\data_o[41] );
  assign \new_[3020]_  = ~\new_[3486]_  & (~\new_[5597]_  | ~\data_o[123] );
  assign \new_[3021]_  = ~\new_[3487]_  & (~\new_[5550]_  | ~\data_o[42] );
  assign \new_[3022]_  = ~\new_[3493]_  & (~\new_[5550]_  | ~\data_o[47] );
  assign \new_[3023]_  = ~\new_[3488]_  & (~\new_[5550]_  | ~\data_o[43] );
  assign \new_[3024]_  = ~\new_[3490]_  & (~\new_[5549]_  | ~\data_o[107] );
  assign \new_[3025]_  = ~\new_[3489]_  & (~\new_[5597]_  | ~\data_o[44] );
  assign \new_[3026]_  = ~\new_[3491]_  & (~\new_[5550]_  | ~\data_o[125] );
  assign \new_[3027]_  = ~\new_[3492]_  & (~\new_[5606]_  | ~\data_o[46] );
  assign \new_[3028]_  = ~\new_[3494]_  & (~\new_[5606]_  | ~\data_o[126] );
  assign \new_[3029]_  = ~\new_[3495]_  & (~\new_[5606]_  | ~\data_o[108] );
  assign \new_[3030]_  = ~\new_[3496]_  & (~\new_[5549]_  | ~\data_o[127] );
  assign \new_[3031]_  = ~\new_[3498]_  & (~\new_[5597]_  | ~\data_o[0] );
  assign \new_[3032]_  = ~\new_[3497]_  & (~\new_[5606]_  | ~\data_o[13] );
  assign \new_[3033]_  = ~\new_[3499]_  & (~\new_[5597]_  | ~\data_o[10] );
  assign \new_[3034]_  = ~\new_[3500]_  & (~\new_[5549]_  | ~\data_o[57] );
  assign \new_[3035]_  = ~\new_[3501]_  & (~\new_[5597]_  | ~\data_o[58] );
  assign \new_[3036]_  = ~\new_[3502]_  & (~\new_[5549]_  | ~\data_o[110] );
  assign \new_[3037]_  = ~\new_[3503]_  & (~\new_[5549]_  | ~\data_o[59] );
  assign \new_[3038]_  = ~\new_[3504]_  & (~\new_[5597]_  | ~\data_o[5] );
  assign \new_[3039]_  = ~\new_[3505]_  & (~\new_[5549]_  | ~\data_o[60] );
  assign \new_[3040]_  = ~\new_[3291]_ ;
  assign \new_[3041]_  = ~\new_[3292]_ ;
  assign \new_[3042]_  = ~\new_[3293]_ ;
  assign \new_[3043]_  = ~\new_[3516]_  | ~\new_[8489]_ ;
  assign \new_[3044]_  = ~\new_[3521]_  & ~\new_[3620]_ ;
  assign \new_[3045]_  = ~\new_[3624]_  & (~\new_[4227]_  | ~\new_[3629]_ );
  assign n3110 = ~\new_[7415]_  | (~\new_[3557]_  & ~\new_[7560]_ );
  assign n3115 = ~\new_[7526]_  | (~\new_[3558]_  & ~\new_[7560]_ );
  assign n3120 = ~\new_[7478]_  | (~\new_[3559]_  & ~\new_[7560]_ );
  assign n3125 = ~\new_[7490]_  | (~\new_[3560]_  & ~\new_[7560]_ );
  assign \new_[3050]_  = (~\new_[3562]_  | ~\new_[8713]_ ) & (~\new_[8063]_  | ~\new_[8716]_ );
  assign \new_[3051]_  = (~\new_[3563]_  | ~\new_[8713]_ ) & (~\new_[8019]_  | ~\new_[8716]_ );
  assign \new_[3052]_  = (~\new_[3564]_  | ~\new_[7825]_ ) & (~\new_[7976]_  | ~\new_[8716]_ );
  assign \new_[3053]_  = (~\new_[3565]_  | ~\new_[8713]_ ) & (~\new_[8074]_  | ~\new_[8716]_ );
  assign \new_[3054]_  = (~\new_[3566]_  | ~\new_[7825]_ ) & (~\new_[7990]_  | ~\new_[8716]_ );
  assign \new_[3055]_  = ~\new_[3340]_  & (~\new_[8143]_  | ~\new_[7645]_ );
  assign \new_[3056]_  = ~\new_[3341]_  & (~\new_[8033]_  | ~\new_[7645]_ );
  assign \new_[3057]_  = ~\new_[3342]_  & (~\new_[8039]_  | ~\new_[7645]_ );
  assign \new_[3058]_  = ~\new_[3343]_  & (~\new_[8154]_  | ~\new_[7645]_ );
  assign \new_[3059]_  = ~\new_[3344]_  & (~\new_[8010]_  | ~\new_[7499]_ );
  assign \new_[3060]_  = ~\new_[3407]_  & (~\new_[4134]_  | ~\new_[8960]_ );
  assign \new_[3061]_  = \new_[1596]_  ^ \new_[3539]_ ;
  assign \new_[3062]_  = ~\new_[3345]_  & (~\new_[7972]_  | ~\new_[7499]_ );
  assign \new_[3063]_  = \new_[1188]_  ^ \new_[3533]_ ;
  assign \new_[3064]_  = \new_[1253]_  ^ \new_[3537]_ ;
  assign \new_[3065]_  = \new_[1466]_  ^ \new_[3538]_ ;
  assign \new_[3066]_  = ~\new_[3346]_  & (~\new_[7978]_  | ~\new_[7499]_ );
  assign \new_[3067]_  = \new_[1307]_  ^ \new_[3534]_ ;
  assign \new_[3068]_  = \new_[1189]_  ^ \new_[3540]_ ;
  assign \new_[3069]_  = \new_[1310]_  ^ \new_[3532]_ ;
  assign \new_[3070]_  = ~\new_[3347]_  & (~\new_[8100]_  | ~\new_[7499]_ );
  assign \new_[3071]_  = (~\new_[3567]_  | ~\new_[8713]_ ) & (~\new_[8021]_  | ~\new_[8716]_ );
  assign \new_[3072]_  = (~\new_[3568]_  | ~\new_[7825]_ ) & (~\new_[8102]_  | ~\new_[8716]_ );
  assign \new_[3073]_  = ~\new_[3529]_  | (~\new_[8710]_  & ~\new_[2224]_ );
  assign \new_[3074]_  = ~\new_[3522]_  | (~\new_[4143]_  & ~\new_[6133]_ );
  assign \new_[3075]_  = ~\new_[3523]_  & ~\new_[3971]_ ;
  assign \new_[3076]_  = ~\new_[3524]_  & (~\new_[4332]_  | ~\new_[6215]_ );
  assign \new_[3077]_  = ~\new_[3526]_  & ~\new_[3569]_ ;
  assign \new_[3078]_  = ~\new_[3527]_  & (~\new_[4332]_  | ~\new_[6058]_ );
  assign \new_[3079]_  = ~\new_[3528]_  & (~\new_[3983]_  | ~\new_[6060]_ );
  assign \new_[3080]_  = ~\new_[3759]_  | ~\new_[8961]_ ;
  assign \new_[3081]_  = ~\new_[3787]_  | ~\new_[8961]_ ;
  assign n3250 = ~\new_[3549]_  | ~\new_[7335]_ ;
  assign n3255 = ~\new_[3550]_  | ~\new_[7363]_ ;
  assign n3260 = ~\new_[3551]_  | ~\new_[7371]_ ;
  assign n3215 = ~\new_[3552]_  | ~\new_[7355]_ ;
  assign n3265 = ~\new_[3553]_  | ~\new_[7198]_ ;
  assign n3270 = ~\new_[3554]_  | ~\new_[7177]_ ;
  assign n3275 = ~\new_[3555]_  | ~\new_[7183]_ ;
  assign n3280 = ~\new_[3556]_  | ~\new_[7318]_ ;
  assign \new_[3090]_  = ~\new_[3560]_  & ~\new_[7829]_ ;
  assign \new_[3091]_  = ~\new_[3557]_  & ~\new_[7829]_ ;
  assign \new_[3092]_  = ~\new_[3558]_  & ~\new_[7829]_ ;
  assign \new_[3093]_  = ~\new_[3559]_  & ~\new_[7829]_ ;
  assign \new_[3094]_  = ~\new_[3560]_  & ~\new_[8562]_ ;
  assign \new_[3095]_  = ~\new_[3557]_  & ~\new_[8562]_ ;
  assign \new_[3096]_  = ~\new_[3558]_  & ~\new_[8562]_ ;
  assign \new_[3097]_  = ~\new_[3559]_  & ~\new_[8562]_ ;
  assign \new_[3098]_  = ~\new_[3355]_ ;
  assign \new_[3099]_  = (~\new_[4155]_  | ~\new_[8958]_ ) & (~\new_[6762]_  | ~\new_[8959]_ );
  assign \new_[3100]_  = (~\new_[4249]_  | ~\new_[8961]_ ) & (~\new_[7041]_  | ~\new_[8964]_ );
  assign \new_[3101]_  = (~\new_[4353]_  | ~\new_[8961]_ ) & (~\new_[6899]_  | ~\new_[8964]_ );
  assign \new_[3102]_  = (~\new_[4354]_  | ~\new_[8961]_ ) & (~\new_[6898]_  | ~\new_[8962]_ );
  assign \new_[3103]_  = \\mix1_data_o_reg_reg[17] ;
  assign \new_[3104]_  = \\mix1_data_o_reg_reg[18] ;
  assign \new_[3105]_  = \\mix1_data_o_reg_reg[1] ;
  assign \new_[3106]_  = \\mix1_data_o_reg_reg[25] ;
  assign \new_[3107]_  = \\mix1_data_o_reg_reg[26] ;
  assign \new_[3108]_  = \\mix1_data_o_reg_reg[9] ;
  assign \new_[3109]_  = \\mix1_data_o_reg_reg[2] ;
  assign \new_[3110]_  = (~\new_[3680]_  | ~\new_[7825]_ ) & (~\new_[8040]_  | ~\new_[8716]_ );
  assign \new_[3111]_  = (~\new_[3681]_  | ~\new_[8713]_ ) & (~\new_[8036]_  | ~\new_[8716]_ );
  assign \new_[3112]_  = (~\new_[3682]_  | ~\new_[8713]_ ) & (~\new_[8112]_  | ~\new_[8716]_ );
  assign \new_[3113]_  = (~\new_[3683]_  | ~\new_[8713]_ ) & (~\new_[8015]_  | ~\new_[8716]_ );
  assign \new_[3114]_  = ~\new_[3888]_  | ~\data_o[100] ;
  assign \new_[3115]_  = ~\new_[3888]_  | ~\data_o[105] ;
  assign \new_[3116]_  = ~\new_[3888]_  | ~\data_o[61] ;
  assign \new_[3117]_  = ~\new_[3886]_  | ~\data_o[18] ;
  assign \new_[3118]_  = ~\new_[3886]_  | ~\data_o[111] ;
  assign \new_[3119]_  = ~\new_[3888]_  | ~\data_o[62] ;
  assign \new_[3120]_  = ~\new_[3888]_  | ~\data_o[63] ;
  assign \new_[3121]_  = ~\new_[3887]_  | ~\data_o[19] ;
  assign \new_[3122]_  = ~\new_[3887]_  | ~\data_o[64] ;
  assign \new_[3123]_  = ~\new_[3887]_  | ~\data_o[65] ;
  assign \new_[3124]_  = ~\new_[3887]_  | ~\data_o[1] ;
  assign \new_[3125]_  = ~\new_[3886]_  | ~\data_o[112] ;
  assign \new_[3126]_  = ~\new_[3886]_  | ~\data_o[66] ;
  assign \new_[3127]_  = ~\new_[3888]_  | ~\data_o[86] ;
  assign \new_[3128]_  = ~\new_[3888]_  | ~\data_o[67] ;
  assign \new_[3129]_  = ~\new_[3887]_  | ~\data_o[20] ;
  assign \new_[3130]_  = ~\new_[3887]_  | ~\data_o[68] ;
  assign \new_[3131]_  = ~\new_[3886]_  | ~\data_o[69] ;
  assign \new_[3132]_  = ~\new_[3886]_  | ~\data_o[21] ;
  assign \new_[3133]_  = ~\new_[3887]_  | ~\data_o[113] ;
  assign \new_[3134]_  = ~\new_[3887]_  | ~\data_o[101] ;
  assign \new_[3135]_  = ~\new_[3888]_  | ~\data_o[6] ;
  assign \new_[3136]_  = ~\new_[3888]_  | ~\data_o[70] ;
  assign \new_[3137]_  = ~\new_[3887]_  | ~\data_o[22] ;
  assign \new_[3138]_  = ~\new_[3887]_  | ~\data_o[71] ;
  assign \new_[3139]_  = ~\new_[3887]_  | ~\data_o[72] ;
  assign \new_[3140]_  = ~\new_[3887]_  | ~\data_o[23] ;
  assign \new_[3141]_  = ~\new_[3888]_  | ~\data_o[114] ;
  assign \new_[3142]_  = ~\new_[3888]_  | ~\data_o[73] ;
  assign \new_[3143]_  = ~\new_[3886]_  | ~\data_o[74] ;
  assign \new_[3144]_  = ~\new_[3886]_  | ~\data_o[24] ;
  assign \new_[3145]_  = ~\new_[3886]_  | ~\data_o[75] ;
  assign \new_[3146]_  = ~\new_[3886]_  | ~\data_o[76] ;
  assign \new_[3147]_  = ~\new_[3888]_  | ~\data_o[25] ;
  assign \new_[3148]_  = ~\new_[3888]_  | ~\data_o[115] ;
  assign \new_[3149]_  = ~\new_[3886]_  | ~\data_o[102] ;
  assign \new_[3150]_  = ~\new_[3886]_  | ~\data_o[77] ;
  assign \new_[3151]_  = ~\new_[3886]_  | ~\data_o[78] ;
  assign \new_[3152]_  = ~\new_[3886]_  | ~\data_o[26] ;
  assign \new_[3153]_  = ~\new_[3887]_  | ~\data_o[79] ;
  assign \new_[3154]_  = ~\new_[3887]_  | ~\data_o[27] ;
  assign \new_[3155]_  = ~\new_[3888]_  | ~\data_o[117] ;
  assign \new_[3156]_  = ~\new_[3888]_  | ~\data_o[80] ;
  assign \new_[3157]_  = ~\new_[3888]_  | ~\data_o[81] ;
  assign \new_[3158]_  = ~\new_[3888]_  | ~\data_o[28] ;
  assign \new_[3159]_  = ~\new_[3888]_  | ~\data_o[82] ;
  assign \new_[3160]_  = ~\new_[3886]_  | ~\data_o[29] ;
  assign \new_[3161]_  = ~\new_[3886]_  | ~\data_o[83] ;
  assign \new_[3162]_  = ~\new_[3888]_  | ~\data_o[103] ;
  assign \new_[3163]_  = ~\new_[3888]_  | ~\data_o[85] ;
  assign \new_[3164]_  = ~\new_[3888]_  | ~\data_o[87] ;
  assign \new_[3165]_  = ~\new_[3888]_  | ~\data_o[30] ;
  assign \new_[3166]_  = ~\new_[3888]_  | ~\data_o[118] ;
  assign \new_[3167]_  = ~\new_[3888]_  | ~\data_o[88] ;
  assign \new_[3168]_  = ~\new_[3886]_  | ~\data_o[89] ;
  assign \new_[3169]_  = ~\new_[3886]_  | ~\data_o[31] ;
  assign \new_[3170]_  = ~\new_[3887]_  | ~\data_o[8] ;
  assign \new_[3171]_  = ~\new_[3887]_  | ~\data_o[90] ;
  assign \new_[3172]_  = ~\new_[3888]_  | ~\data_o[32] ;
  assign \new_[3173]_  = ~\new_[3888]_  | ~\data_o[119] ;
  assign \new_[3174]_  = ~\new_[3887]_  | ~\data_o[104] ;
  assign \new_[3175]_  = ~\new_[3887]_  | ~\data_o[91] ;
  assign \new_[3176]_  = ~\new_[3888]_  | ~\data_o[92] ;
  assign \new_[3177]_  = ~\new_[3888]_  | ~\data_o[33] ;
  assign \new_[3178]_  = ~\new_[3888]_  | ~\data_o[93] ;
  assign \new_[3179]_  = ~\new_[3888]_  | ~\data_o[94] ;
  assign \new_[3180]_  = ~\new_[3886]_  | ~\data_o[34] ;
  assign \new_[3181]_  = ~\new_[3886]_  | ~\data_o[11] ;
  assign \new_[3182]_  = ~\new_[3888]_  | ~\data_o[95] ;
  assign \new_[3183]_  = ~\new_[3888]_  | ~\data_o[84] ;
  assign \new_[3184]_  = ~\new_[3887]_  | ~\data_o[96] ;
  assign \new_[3185]_  = ~\new_[3887]_  | ~\data_o[35] ;
  assign \new_[3186]_  = ~\new_[3887]_  | ~\data_o[97] ;
  assign \new_[3187]_  = ~\new_[3887]_  | ~\data_o[98] ;
  assign \new_[3188]_  = ~\new_[3886]_  | ~\data_o[36] ;
  assign \new_[3189]_  = ~\new_[3886]_  | ~\data_o[120] ;
  assign \new_[3190]_  = ~\new_[3886]_  | ~\data_o[99] ;
  assign \new_[3191]_  = ~\new_[3886]_  | ~\data_o[2] ;
  assign \new_[3192]_  = ~\new_[3888]_  | ~\data_o[9] ;
  assign n3285 = ~\new_[3577]_  | ~\new_[7220]_ ;
  assign \new_[3194]_  = ~\new_[3888]_  | ~\data_o[37] ;
  assign n3320 = ~\new_[3571]_  | ~\new_[7331]_ ;
  assign \new_[3196]_  = ~\new_[3887]_  | ~\data_o[38] ;
  assign \new_[3197]_  = ~\new_[3887]_  | ~\data_o[121] ;
  assign n3290 = ~\new_[3572]_  | ~\new_[7109]_ ;
  assign \new_[3199]_  = ~\new_[3888]_  | ~\data_o[39] ;
  assign n3295 = ~\new_[3573]_  | ~\new_[7258]_ ;
  assign \new_[3201]_  = ~\new_[3888]_  | ~\data_o[116] ;
  assign \new_[3202]_  = ~\new_[3886]_  | ~\data_o[3] ;
  assign n3300 = ~\new_[3574]_  | ~\new_[7189]_ ;
  assign \new_[3204]_  = ~\new_[3886]_  | ~\data_o[122] ;
  assign \new_[3205]_  = ~\new_[3888]_  | ~\data_o[106] ;
  assign \new_[3206]_  = ~\new_[3888]_  | ~\data_o[40] ;
  assign n3315 = ~\new_[3575]_  | ~\new_[7194]_ ;
  assign \new_[3208]_  = ~\new_[3886]_  | ~\data_o[41] ;
  assign \new_[3209]_  = ~\new_[3886]_  | ~\data_o[123] ;
  assign n3310 = ~\new_[3576]_  | ~\new_[7247]_ ;
  assign \new_[3211]_  = ~\new_[3888]_  | ~\data_o[42] ;
  assign \new_[3212]_  = ~\new_[3888]_  | ~\data_o[108] ;
  assign \new_[3213]_  = ~\new_[3887]_  | ~\data_o[46] ;
  assign \new_[3214]_  = ~\new_[3887]_  | ~\data_o[43] ;
  assign n3305 = ~\new_[3578]_  | ~\new_[7166]_ ;
  assign \new_[3216]_  = ~\new_[3888]_  | ~\data_o[107] ;
  assign \new_[3217]_  = ~\new_[3888]_  | ~\data_o[44] ;
  assign \new_[3218]_  = ~\new_[3888]_  | ~\data_o[124] ;
  assign \new_[3219]_  = ~\new_[3888]_  | ~\data_o[125] ;
  assign \new_[3220]_  = ~\new_[3888]_  | ~\data_o[126] ;
  assign \new_[3221]_  = ~\new_[3888]_  | ~\data_o[47] ;
  assign \new_[3222]_  = ~\new_[3887]_  | ~\data_o[7] ;
  assign \new_[3223]_  = ~\new_[3887]_  | ~\data_o[45] ;
  assign \new_[3224]_  = ~\new_[3888]_  | ~\data_o[48] ;
  assign \new_[3225]_  = ~\new_[3888]_  | ~\data_o[49] ;
  assign \new_[3226]_  = ~\new_[3888]_  | ~\data_o[127] ;
  assign \new_[3227]_  = ~\new_[3888]_  | ~\data_o[4] ;
  assign \new_[3228]_  = ~\new_[3888]_  | ~\data_o[50] ;
  assign \new_[3229]_  = ~\new_[3888]_  | ~\data_o[0] ;
  assign \new_[3230]_  = ~\new_[3887]_  | ~\data_o[12] ;
  assign \new_[3231]_  = ~\new_[3887]_  | ~\data_o[109] ;
  assign \new_[3232]_  = ~\new_[3888]_  | ~\data_o[51] ;
  assign \new_[3233]_  = ~\new_[3888]_  | ~\data_o[52] ;
  assign \new_[3234]_  = ~\new_[3888]_  | ~\data_o[13] ;
  assign \new_[3235]_  = ~\new_[8888]_  | ~\new_[8660]_ ;
  assign \new_[3236]_  = ~\new_[3888]_  | ~\data_o[53] ;
  assign \new_[3237]_  = ~\new_[3888]_  | ~\data_o[54] ;
  assign \new_[3238]_  = ~\new_[3888]_  | ~\data_o[14] ;
  assign \new_[3239]_  = ~\new_[3887]_  | ~\data_o[10] ;
  assign \new_[3240]_  = ~\new_[3887]_  | ~\data_o[55] ;
  assign \new_[3241]_  = ~\new_[3888]_  | ~\data_o[56] ;
  assign \new_[3242]_  = ~\new_[3888]_  | ~\data_o[15] ;
  assign \new_[3243]_  = ~\new_[3888]_  | ~\data_o[57] ;
  assign \new_[3244]_  = ~\new_[3888]_  | ~\data_o[58] ;
  assign \new_[3245]_  = ~\new_[3888]_  | ~\data_o[16] ;
  assign \new_[3246]_  = ~\new_[3888]_  | ~\data_o[110] ;
  assign \new_[3247]_  = ~\new_[3886]_  | ~\data_o[59] ;
  assign \new_[3248]_  = ~\new_[3886]_  | ~\data_o[5] ;
  assign \new_[3249]_  = ~\new_[3886]_  | ~\data_o[17] ;
  assign \new_[3250]_  = ~\new_[3886]_  | ~\data_o[60] ;
  assign \new_[3251]_  = (~\new_[3827]_  | ~\new_[8713]_ ) & (~\new_[8066]_  | ~\new_[8716]_ );
  assign \new_[3252]_  = (~\new_[3828]_  | ~\new_[7825]_ ) & (~\new_[7988]_  | ~\new_[8716]_ );
  assign \new_[3253]_  = (~\new_[3829]_  | ~\new_[8713]_ ) & (~\new_[8002]_  | ~\new_[8716]_ );
  assign \new_[3254]_  = (~\new_[3830]_  | ~\new_[7825]_ ) & (~\new_[8117]_  | ~\new_[8716]_ );
  assign \new_[3255]_  = ~\new_[3579]_  & (~\new_[5606]_  | ~\data_o[61] );
  assign \new_[3256]_  = ~\new_[3580]_  & (~\new_[5597]_  | ~\data_o[62] );
  assign \new_[3257]_  = \\mix1_data_o_reg_reg[10] ;
  assign \new_[3258]_  = ~\new_[3581]_  & (~\new_[5549]_  | ~\data_o[1] );
  assign \new_[3259]_  = ~\new_[3582]_  & (~\new_[5549]_  | ~\data_o[72] );
  assign \new_[3260]_  = ~\new_[3583]_  & (~\new_[5549]_  | ~\data_o[73] );
  assign \new_[3261]_  = ~\new_[3585]_  & (~\new_[5550]_  | ~\data_o[74] );
  assign \new_[3262]_  = ~\new_[3584]_  & (~\new_[5606]_  | ~\data_o[24] );
  assign \new_[3263]_  = ~\new_[3586]_  & (~\new_[5550]_  | ~\data_o[75] );
  assign \new_[3264]_  = ~\new_[3587]_  & (~\new_[5597]_  | ~\data_o[7] );
  assign \new_[3265]_  = ~\new_[3588]_  & (~\new_[5550]_  | ~\data_o[27] );
  assign \new_[3266]_  = ~\new_[3589]_  & (~\new_[5606]_  | ~\data_o[28] );
  assign \new_[3267]_  = ~\new_[3590]_  & (~\new_[5597]_  | ~\data_o[2] );
  assign \new_[3268]_  = ~\new_[3591]_  & (~\new_[5549]_  | ~\data_o[30] );
  assign \new_[3269]_  = ~\new_[3592]_  & (~\new_[5606]_  | ~\data_o[31] );
  assign \new_[3270]_  = ~\new_[3593]_  & (~\new_[5597]_  | ~\data_o[90] );
  assign \new_[3271]_  = ~\new_[3594]_  & (~\new_[5597]_  | ~\data_o[91] );
  assign \new_[3272]_  = ~\new_[3595]_  & (~\new_[5549]_  | ~\data_o[104] );
  assign \new_[3273]_  = ~\new_[3596]_  & (~\new_[5597]_  | ~\data_o[92] );
  assign \new_[3274]_  = ~\new_[3597]_  & (~\new_[5597]_  | ~\data_o[93] );
  assign \new_[3275]_  = ~\new_[3598]_  & (~\new_[5606]_  | ~\data_o[94] );
  assign \new_[3276]_  = ~\new_[3599]_  & (~\new_[5549]_  | ~\data_o[34] );
  assign \new_[3277]_  = ~\new_[3600]_  & (~\new_[5549]_  | ~\data_o[11] );
  assign \new_[3278]_  = ~\new_[3601]_  & (~\new_[5550]_  | ~\data_o[95] );
  assign \new_[3279]_  = ~\new_[3602]_  & (~\new_[5597]_  | ~\data_o[120] );
  assign \new_[3280]_  = ~\new_[3603]_  & (~\new_[5549]_  | ~\data_o[9] );
  assign \new_[3281]_  = ~\new_[3604]_  & (~\new_[5549]_  | ~\data_o[121] );
  assign \new_[3282]_  = ~\new_[3605]_  & (~\new_[5597]_  | ~\data_o[40] );
  assign \new_[3283]_  = ~\new_[3606]_  & (~\new_[5550]_  | ~\data_o[124] );
  assign \new_[3284]_  = ~\new_[3607]_  & (~\new_[5549]_  | ~\data_o[45] );
  assign \new_[3285]_  = ~\new_[3608]_  & (~\new_[5550]_  | ~\data_o[4] );
  assign \new_[3286]_  = ~\new_[3609]_  & (~\new_[5597]_  | ~\data_o[12] );
  assign \new_[3287]_  = ~\new_[3610]_  & (~\new_[5606]_  | ~\data_o[109] );
  assign \new_[3288]_  = ~\new_[3611]_  & (~\new_[5597]_  | ~\data_o[14] );
  assign \new_[3289]_  = ~\new_[3612]_  & (~\new_[5597]_  | ~\data_o[56] );
  assign \new_[3290]_  = ~\new_[3613]_  & (~\new_[5549]_  | ~\data_o[15] );
  assign \new_[3291]_  = ~\new_[4322]_  | ~\new_[3614]_ ;
  assign \new_[3292]_  = ~\new_[4421]_  | ~\new_[3615]_ ;
  assign \new_[3293]_  = ~\new_[4324]_  | ~\new_[3616]_ ;
  assign n3230 = ~\new_[3617]_  | ~\new_[7346]_ ;
  assign n3225 = ~\new_[3618]_  | ~\new_[7199]_ ;
  assign n3235 = ~\new_[3619]_  | ~\new_[7354]_ ;
  assign n3210 = ~\new_[3621]_  | ~\new_[7289]_ ;
  assign n3220 = ~\new_[3625]_  | ~\new_[7162]_ ;
  assign n3240 = ~\new_[3626]_  | ~\new_[7173]_ ;
  assign n3340 = ~\new_[3627]_  | ~\new_[7179]_ ;
  assign n3345 = ~\new_[3628]_  | ~\new_[7090]_ ;
  assign \new_[3302]_  = ~\new_[3620]_  & (~\new_[3825]_  | ~\new_[3839]_ );
  assign \new_[3303]_  = ~\new_[3624]_  & (~\new_[3839]_  | ~\new_[4135]_ );
  assign \new_[3304]_  = ~\new_[3624]_  & (~\new_[4227]_  | ~\new_[3976]_ );
  assign \new_[3305]_  = \new_[8041]_  ^ \new_[3831]_ ;
  assign \new_[3306]_  = \new_[8024]_  ^ \new_[3832]_ ;
  assign \new_[3307]_  = \new_[8023]_  ^ \new_[3833]_ ;
  assign \new_[3308]_  = \new_[7959]_  ^ \new_[3834]_ ;
  assign \new_[3309]_  = \new_[8027]_  ^ \new_[3835]_ ;
  assign \new_[3310]_  = \new_[8050]_  ^ \new_[3836]_ ;
  assign n3330 = ~\new_[7449]_  | (~\new_[3647]_  & ~\new_[7560]_ );
  assign n3335 = ~\new_[7542]_  | (~\new_[3649]_  & ~\new_[7560]_ );
  assign n3325 = ~\new_[7473]_  | (~\new_[3651]_  & ~\new_[7560]_ );
  assign n3245 = ~\new_[7434]_  | (~\new_[3653]_  & ~\new_[7560]_ );
  assign \new_[3315]_  = (~\new_[3655]_  | ~\new_[8713]_ ) & (~\new_[8085]_  | ~\new_[8716]_ );
  assign \new_[3316]_  = (~\new_[3656]_  | ~\new_[8713]_ ) & (~\new_[7948]_  | ~\new_[8716]_ );
  assign \new_[3317]_  = (~\new_[3657]_  | ~\new_[7825]_ ) & (~\new_[8118]_  | ~\new_[8716]_ );
  assign \new_[3318]_  = (~\new_[3658]_  | ~\new_[8713]_ ) & (~\new_[7966]_  | ~\new_[8716]_ );
  assign \new_[3319]_  = \new_[1317]_  ^ \new_[3642]_ ;
  assign \new_[3320]_  = ~\new_[3530]_  | (~\new_[8710]_  & ~\new_[2346]_ );
  assign \new_[3321]_  = ~\new_[3531]_  | (~\new_[8710]_  & ~\new_[2347]_ );
  assign \new_[3322]_  = ~\new_[3631]_  | (~\new_[4143]_  & ~\new_[6140]_ );
  assign \new_[3323]_  = ~\new_[3632]_  | (~\new_[4143]_  & ~\new_[6070]_ );
  assign \new_[3324]_  = ~\new_[3633]_  | (~\new_[4143]_  & ~\new_[6134]_ );
  assign \new_[3325]_  = ~\new_[4186]_  & ~\new_[8954]_ ;
  assign \new_[3326]_  = ~\new_[4137]_  & ~\new_[8954]_ ;
  assign \new_[3327]_  = ~\new_[3847]_  & ~\new_[8954]_ ;
  assign \new_[3328]_  = ~\new_[4138]_  & ~\new_[8954]_ ;
  assign \new_[3329]_  = ~\new_[4139]_  & ~\new_[8954]_ ;
  assign \new_[3330]_  = ~\new_[4140]_  & ~\new_[8954]_ ;
  assign \new_[3331]_  = ~\new_[4141]_  & ~\new_[8954]_ ;
  assign \new_[3332]_  = ~\new_[3848]_  & ~\new_[8954]_ ;
  assign \new_[3333]_  = ~\new_[3849]_  & ~\new_[8954]_ ;
  assign \new_[3334]_  = ~\new_[4142]_  & ~\new_[8954]_ ;
  assign \new_[3335]_  = \new_[3850]_  | \new_[8963]_ ;
  assign \new_[3336]_  = \new_[3851]_  | \new_[8963]_ ;
  assign \new_[3337]_  = \new_[3853]_  | \new_[8963]_ ;
  assign \new_[3338]_  = ~\new_[3854]_  & ~\new_[8964]_ ;
  assign \new_[3339]_  = ~\new_[3856]_  & ~\new_[8964]_ ;
  assign \new_[3340]_  = ~\new_[3653]_  & ~\new_[7829]_ ;
  assign \new_[3341]_  = ~\new_[3647]_  & ~\new_[7829]_ ;
  assign \new_[3342]_  = ~\new_[3649]_  & ~\new_[7829]_ ;
  assign \new_[3343]_  = ~\new_[3651]_  & ~\new_[7829]_ ;
  assign \new_[3344]_  = ~\new_[3653]_  & ~\new_[8562]_ ;
  assign \new_[3345]_  = ~\new_[3647]_  & ~\new_[8562]_ ;
  assign \new_[3346]_  = ~\new_[3649]_  & ~\new_[8562]_ ;
  assign \new_[3347]_  = ~\new_[3651]_  & ~\new_[8562]_ ;
  assign \new_[3348]_  = (~\new_[4333]_  & ~\new_[8962]_ ) | (~\new_[6741]_  & ~\new_[8960]_ );
  assign \new_[3349]_  = (~\new_[4334]_  & ~\new_[8962]_ ) | (~\new_[6608]_  & ~\new_[8960]_ );
  assign \new_[3350]_  = (~\new_[4339]_  | ~\new_[8961]_ ) & (~\new_[7045]_  | ~\new_[8964]_ );
  assign \new_[3351]_  = (~\new_[4337]_  | ~\new_[8961]_ ) & (~\new_[7140]_  | ~\new_[8963]_ );
  assign \new_[3352]_  = (~\new_[4341]_  | ~\new_[8961]_ ) & (~\new_[7119]_  | ~\new_[8964]_ );
  assign \new_[3353]_  = (~\new_[4342]_  | ~\new_[8961]_ ) & (~\new_[7149]_  | ~\new_[8964]_ );
  assign \new_[3354]_  = (~\new_[4343]_  | ~\new_[8961]_ ) & (~\new_[7142]_  | ~\new_[8964]_ );
  assign \new_[3355]_  = (~\new_[4344]_  | ~\new_[8961]_ ) & (~\new_[7143]_  | ~\new_[8963]_ );
  assign \new_[3356]_  = ~\new_[3535]_ ;
  assign \new_[3357]_  = ~\new_[8267]_ ;
  assign \new_[3358]_  = ~\new_[8231]_ ;
  assign \new_[3359]_  = ~\new_[3536]_ ;
  assign \new_[3360]_  = (~\new_[4239]_  & ~\new_[8962]_ ) | (~\new_[7051]_  & ~\new_[8961]_ );
  assign \new_[3361]_  = (~\new_[4245]_  | ~\new_[8961]_ ) & (~\new_[7144]_  | ~\new_[8964]_ );
  assign \new_[3362]_  = (~\new_[4250]_  & ~\new_[8962]_ ) | (~\new_[6924]_  & ~\new_[8961]_ );
  assign \new_[3363]_  = (~\new_[4251]_  & ~\new_[8962]_ ) | (~\new_[6735]_  & ~\new_[8961]_ );
  assign \new_[3364]_  = (~\new_[4252]_  & ~\new_[8962]_ ) | (~\new_[6738]_  & ~\new_[8961]_ );
  assign \new_[3365]_  = (~\new_[4253]_  & ~\new_[8962]_ ) | (~\new_[7055]_  & ~\new_[8961]_ );
  assign \new_[3366]_  = (~\new_[4351]_  | ~\new_[8961]_ ) & (~\new_[7058]_  | ~\new_[8964]_ );
  assign \new_[3367]_  = (~\new_[4254]_  & ~\new_[8962]_ ) | (~\new_[7059]_  & ~\new_[8961]_ );
  assign \new_[3368]_  = (~\new_[4255]_  & ~\new_[8962]_ ) | (~\new_[7048]_  & ~\new_[8961]_ );
  assign \new_[3369]_  = (~\new_[4256]_  & ~\new_[8962]_ ) | (~\new_[7039]_  & ~\new_[8961]_ );
  assign \new_[3370]_  = (~\new_[4257]_  & ~\new_[8964]_ ) | (~\new_[7053]_  & ~\new_[8961]_ );
  assign \new_[3371]_  = (~\new_[4258]_  & ~\new_[8963]_ ) | (~\new_[7060]_  & ~\new_[8961]_ );
  assign \new_[3372]_  = (~\new_[4352]_  & ~\new_[8962]_ ) | (~\new_[6742]_  & ~\new_[8960]_ );
  assign \new_[3373]_  = (~\new_[4259]_  & ~\new_[8962]_ ) | (~\new_[6743]_  & ~\new_[8960]_ );
  assign \new_[3374]_  = (~\new_[4260]_  & ~\new_[8962]_ ) | (~\new_[6744]_  & ~\new_[8961]_ );
  assign \new_[3375]_  = (~\new_[4261]_  & ~\new_[8962]_ ) | (~\new_[7040]_  & ~\new_[8961]_ );
  assign \new_[3376]_  = ~\\mix1_data_reg_reg[79] ;
  assign \new_[3377]_  = \\mix1_data_o_reg_reg[8] ;
  assign \new_[3378]_  = ~\\mix1_data_reg_reg[55] ;
  assign \new_[3379]_  = (~\new_[4355]_  | ~\new_[8961]_ ) & (~\new_[7037]_  | ~\new_[8964]_ );
  assign \new_[3380]_  = (~\new_[4262]_  & ~\new_[8963]_ ) | (~\new_[6740]_  & ~\new_[8961]_ );
  assign \new_[3381]_  = ~\\mix1_data_reg_reg[71] ;
  assign \new_[3382]_  = \\mix1_data_o_reg_reg[13] ;
  assign \new_[3383]_  = \\mix1_data_o_reg_reg[21] ;
  assign \new_[3384]_  = ~\\mix1_data_reg_reg[63] ;
  assign \new_[3385]_  = \\mix1_data_o_reg_reg[22] ;
  assign \new_[3386]_  = \\mix1_data_o_reg_reg[30] ;
  assign \new_[3387]_  = \\mix1_data_o_reg_reg[16] ;
  assign \new_[3388]_  = ~\\mix1_data_reg_reg[47] ;
  assign \new_[3389]_  = ~\\mix1_data_reg_reg[39] ;
  assign \new_[3390]_  = ~\new_[3659]_  & (~\new_[8016]_  | ~\new_[7645]_ );
  assign \new_[3391]_  = ~\new_[3660]_  & (~\new_[8099]_  | ~\new_[7645]_ );
  assign \new_[3392]_  = ~\new_[3661]_  & (~\new_[8044]_  | ~\new_[7645]_ );
  assign \new_[3393]_  = ~\new_[3662]_  & (~\new_[8007]_  | ~\new_[7645]_ );
  assign \new_[3394]_  = ~\new_[3663]_  & (~\new_[8090]_  | ~\new_[7645]_ );
  assign \new_[3395]_  = ~\new_[3664]_  & (~\new_[8128]_  | ~\new_[7645]_ );
  assign \new_[3396]_  = ~\new_[3665]_  & (~\new_[8062]_  | ~\new_[7645]_ );
  assign \new_[3397]_  = ~\new_[3666]_  & (~\new_[8048]_  | ~\new_[7645]_ );
  assign \new_[3398]_  = ~\new_[3667]_  & (~\new_[8067]_  | ~\new_[7499]_ );
  assign \new_[3399]_  = ~\new_[3668]_  & (~\new_[8129]_  | ~\new_[7499]_ );
  assign \new_[3400]_  = ~\new_[3669]_  & (~\new_[7940]_  | ~\new_[7499]_ );
  assign \new_[3401]_  = ~\new_[3670]_  & (~\new_[7938]_  | ~\new_[7499]_ );
  assign \new_[3402]_  = ~\new_[3671]_  & (~\new_[8126]_  | ~\new_[7499]_ );
  assign \new_[3403]_  = ~\new_[3672]_  & (~\new_[7998]_  | ~\new_[7499]_ );
  assign \new_[3404]_  = ~\new_[3673]_  & (~\new_[8081]_  | ~\new_[7499]_ );
  assign \new_[3405]_  = ~\new_[3674]_  & (~\new_[8091]_  | ~\new_[7499]_ );
  assign \new_[3406]_  = \\mix1_data_o_reg_reg[6] ;
  assign \new_[3407]_  = ~\new_[6602]_  & ~\new_[8965]_ ;
  assign \new_[3408]_  = ~\new_[8891]_  | ~\new_[4361]_ ;
  assign \new_[3409]_  = \\mix1_data_o_reg_reg[14] ;
  assign \new_[3410]_  = \\mix1_data_o_reg_reg[0] ;
  assign \new_[3411]_  = ~\new_[3684]_  & (~\new_[5606]_  | ~\data_o[18] );
  assign \new_[3412]_  = ~\new_[3686]_  & (~\new_[5597]_  | ~\data_o[19] );
  assign \new_[3413]_  = ~\new_[3685]_  & (~\new_[5549]_  | ~\data_o[100] );
  assign \new_[3414]_  = ~\new_[3687]_  & (~\new_[5597]_  | ~\data_o[64] );
  assign \new_[3415]_  = ~\new_[3688]_  & (~\new_[5549]_  | ~\data_o[65] );
  assign \new_[3416]_  = ~\new_[3689]_  & (~\new_[5597]_  | ~\data_o[112] );
  assign \new_[3417]_  = ~\new_[3690]_  & (~\new_[5597]_  | ~\data_o[66] );
  assign \new_[3418]_  = ~\new_[3691]_  & (~\new_[5549]_  | ~\data_o[67] );
  assign \new_[3419]_  = ~\new_[3692]_  & (~\new_[5549]_  | ~\data_o[20] );
  assign \new_[3420]_  = ~\new_[3693]_  & (~\new_[5549]_  | ~\data_o[68] );
  assign \new_[3421]_  = ~\new_[3694]_  & (~\new_[5597]_  | ~\data_o[69] );
  assign \new_[3422]_  = ~\new_[3696]_  & (~\new_[5606]_  | ~\data_o[21] );
  assign \new_[3423]_  = ~\new_[3695]_  & (~\new_[5549]_  | ~\data_o[113] );
  assign \new_[3424]_  = ~\new_[3697]_  & (~\new_[5550]_  | ~\data_o[101] );
  assign \new_[3425]_  = ~\new_[3698]_  & (~\new_[5606]_  | ~\data_o[70] );
  assign \new_[3426]_  = ~\new_[3699]_  & (~\new_[5606]_  | ~\data_o[22] );
  assign \new_[3427]_  = ~\new_[3700]_  & (~\new_[5597]_  | ~\data_o[71] );
  assign \new_[3428]_  = ~\new_[3702]_  & (~\new_[5550]_  | ~\data_o[23] );
  assign \new_[3429]_  = ~\new_[3701]_  & (~\new_[5549]_  | ~\data_o[114] );
  assign \new_[3430]_  = ~\new_[3704]_  & (~\new_[5606]_  | ~\data_o[102] );
  assign \new_[3431]_  = ~\new_[3703]_  & (~\new_[5606]_  | ~\data_o[115] );
  assign \new_[3432]_  = ~\new_[3705]_  & (~\new_[5549]_  | ~\data_o[116] );
  assign \new_[3433]_  = ~\new_[3706]_  & (~\new_[5549]_  | ~\data_o[80] );
  assign \new_[3434]_  = ~\new_[3707]_  & (~\new_[5597]_  | ~\data_o[81] );
  assign \new_[3435]_  = ~\new_[3708]_  & (~\new_[5597]_  | ~\data_o[82] );
  assign \new_[3436]_  = ~\new_[3709]_  & (~\new_[5549]_  | ~\data_o[83] );
  assign \new_[3437]_  = ~\new_[3710]_  & (~\new_[5549]_  | ~\data_o[103] );
  assign \new_[3438]_  = ~\new_[3711]_  & (~\new_[5597]_  | ~\data_o[117] );
  assign \new_[3439]_  = ~\new_[3712]_  & (~\new_[5550]_  | ~\data_o[84] );
  assign \new_[3440]_  = ~\new_[3713]_  & (~\new_[5549]_  | ~\data_o[85] );
  assign \new_[3441]_  = ~\new_[3714]_  & (~\new_[5549]_  | ~\data_o[86] );
  assign \new_[3442]_  = ~\new_[3715]_  & (~\new_[5549]_  | ~\data_o[87] );
  assign \new_[3443]_  = \\mix1_data_o_reg_reg[24] ;
  assign \new_[3444]_  = ~\new_[3716]_  & (~\new_[5550]_  | ~\data_o[118] );
  assign \new_[3445]_  = ~\new_[3717]_  & (~\new_[5550]_  | ~\data_o[88] );
  assign \new_[3446]_  = ~\new_[3718]_  & (~\new_[5549]_  | ~\data_o[89] );
  assign \new_[3447]_  = ~\new_[3719]_  & (~\new_[5549]_  | ~\data_o[32] );
  assign \new_[3448]_  = ~\new_[3720]_  & (~\new_[5606]_  | ~\data_o[119] );
  assign \new_[3449]_  = ~\new_[3721]_  & (~\new_[5597]_  | ~\data_o[33] );
  assign \new_[3450]_  = ~\new_[3723]_  & (~\new_[5597]_  | ~\data_o[96] );
  assign \new_[3451]_  = ~\new_[3724]_  & (~\new_[5550]_  | ~\data_o[35] );
  assign \new_[3452]_  = ~\new_[3725]_  & (~\new_[5550]_  | ~\data_o[97] );
  assign \new_[3453]_  = ~\new_[3727]_  & (~\new_[5597]_  | ~\data_o[98] );
  assign \new_[3454]_  = ~\new_[3726]_  & (~\new_[5549]_  | ~\data_o[36] );
  assign \new_[3455]_  = ~\new_[3728]_  & (~\new_[5549]_  | ~\data_o[99] );
  assign \new_[3456]_  = ~\new_[3729]_  & (~\new_[5549]_  | ~\data_o[37] );
  assign \new_[3457]_  = ~\new_[3730]_  & (~\new_[5549]_  | ~\data_o[38] );
  assign \new_[3458]_  = ~\new_[3722]_  & (~\new_[5550]_  | ~\data_o[39] );
  assign \new_[3459]_  = ~\new_[3734]_  & (~\new_[5597]_  | ~\data_o[48] );
  assign \new_[3460]_  = ~\new_[3731]_  & (~\new_[5549]_  | ~\data_o[49] );
  assign \new_[3461]_  = ~\new_[3732]_  & (~\new_[5550]_  | ~\data_o[50] );
  assign \new_[3462]_  = ~\new_[3735]_  & (~\new_[5549]_  | ~\data_o[52] );
  assign \new_[3463]_  = ~\new_[3733]_  & (~\new_[5550]_  | ~\data_o[51] );
  assign \new_[3464]_  = ~\new_[3736]_  & (~\new_[5549]_  | ~\data_o[53] );
  assign \new_[3465]_  = ~\new_[3737]_  & (~\new_[5550]_  | ~\data_o[54] );
  assign \new_[3466]_  = ~\new_[3738]_  & (~\new_[5549]_  | ~\data_o[55] );
  assign \new_[3467]_  = ~\new_[3739]_  & (~\new_[5606]_  | ~\data_o[16] );
  assign \new_[3468]_  = ~\new_[3740]_  & (~\new_[5606]_  | ~\data_o[17] );
  assign \new_[3469]_  = ~\new_[8888]_ ;
  assign \new_[3470]_  = ~\new_[3778]_  & ~\new_[5551]_ ;
  assign \new_[3471]_  = ~\new_[3779]_  & ~\new_[5553]_ ;
  assign \new_[3472]_  = ~\new_[3780]_  & ~\new_[5552]_ ;
  assign \new_[3473]_  = ~\new_[3781]_  & ~\new_[5552]_ ;
  assign \new_[3474]_  = ~\new_[3782]_  & ~\new_[5552]_ ;
  assign \new_[3475]_  = ~\new_[3783]_  & ~\new_[5553]_ ;
  assign \new_[3476]_  = ~\new_[3784]_  & ~\new_[5606]_ ;
  assign \new_[3477]_  = ~\new_[3785]_  & ~\new_[5606]_ ;
  assign \new_[3478]_  = ~\new_[3786]_  & ~\new_[5606]_ ;
  assign \new_[3479]_  = ~\new_[3788]_  & ~\new_[5552]_ ;
  assign \new_[3480]_  = ~\new_[3789]_  & ~\new_[5552]_ ;
  assign \new_[3481]_  = ~\new_[3790]_  & ~\new_[5551]_ ;
  assign \new_[3482]_  = ~\new_[3791]_  & ~\new_[5606]_ ;
  assign \new_[3483]_  = ~\new_[3793]_  & ~\new_[5552]_ ;
  assign \new_[3484]_  = ~\new_[3792]_  & ~\new_[5553]_ ;
  assign \new_[3485]_  = ~\new_[3794]_  & ~\new_[5551]_ ;
  assign \new_[3486]_  = ~\new_[3795]_  & ~\new_[5551]_ ;
  assign \new_[3487]_  = ~\new_[3796]_  & ~\new_[5551]_ ;
  assign \new_[3488]_  = ~\new_[3797]_  & ~\new_[5606]_ ;
  assign \new_[3489]_  = ~\new_[3799]_  & ~\new_[5552]_ ;
  assign \new_[3490]_  = ~\new_[3798]_  & ~\new_[5551]_ ;
  assign \new_[3491]_  = ~\new_[3800]_  & ~\new_[5553]_ ;
  assign \new_[3492]_  = ~\new_[3801]_  & ~\new_[5553]_ ;
  assign \new_[3493]_  = ~\new_[3803]_  & ~\new_[5552]_ ;
  assign \new_[3494]_  = ~\new_[3804]_  & ~\new_[5553]_ ;
  assign \new_[3495]_  = ~\new_[3802]_  & ~\new_[5553]_ ;
  assign \new_[3496]_  = ~\new_[3805]_  & ~\new_[5553]_ ;
  assign \new_[3497]_  = ~\new_[3806]_  & ~\new_[5606]_ ;
  assign \new_[3498]_  = ~\new_[3808]_  & ~\new_[5553]_ ;
  assign \new_[3499]_  = ~\new_[3807]_  & ~\new_[5552]_ ;
  assign \new_[3500]_  = ~\new_[3809]_  & ~\new_[5551]_ ;
  assign \new_[3501]_  = ~\new_[3810]_  & ~\new_[5552]_ ;
  assign \new_[3502]_  = ~\new_[3811]_  & ~\new_[5552]_ ;
  assign \new_[3503]_  = ~\new_[3812]_  & ~\new_[5606]_ ;
  assign \new_[3504]_  = ~\new_[3813]_  & ~\new_[5552]_ ;
  assign \new_[3505]_  = ~\new_[3814]_  & ~\new_[5606]_ ;
  assign \new_[3506]_  = (~\new_[3969]_  | ~\new_[8489]_ ) & (~\new_[4465]_  | ~\new_[5794]_ );
  assign \new_[3507]_  = ~\new_[8374]_  | ~\new_[8489]_ ;
  assign \new_[3508]_  = ~\new_[3815]_  | ~\new_[8489]_ ;
  assign n3350 = ~\new_[3821]_  | ~\new_[7382]_ ;
  assign n3355 = ~\new_[3822]_  | ~\new_[7368]_ ;
  assign n3365 = ~\new_[3823]_  | ~\new_[7375]_ ;
  assign n3360 = ~\new_[3824]_  | ~\new_[7336]_ ;
  assign \new_[3513]_  = ~\\mix1_data_reg_reg[95] ;
  assign \new_[3514]_  = \\mix1_data_o_reg_reg[29] ;
  assign \new_[3515]_  = \\mix1_data_o_reg_reg[5] ;
  assign \new_[3516]_  = ~\new_[3816]_  | ~\new_[4326]_ ;
  assign \new_[3517]_  = \new_[8096]_  ^ \new_[3973]_ ;
  assign \new_[3518]_  = \new_[8120]_  ^ \new_[3977]_ ;
  assign \new_[3519]_  = ~\\mix1_data_reg_reg[87] ;
  assign \new_[3520]_  = ~\new_[3620]_ ;
  assign \new_[3521]_  = ~\new_[4227]_  & ~\new_[3826]_ ;
  assign \new_[3522]_  = ~\new_[4164]_  | ~\new_[8960]_ ;
  assign \new_[3523]_  = ~\new_[4229]_  & ~\new_[8964]_ ;
  assign \new_[3524]_  = ~\new_[4234]_  & ~\new_[8954]_ ;
  assign \new_[3525]_  = ~\new_[3868]_  & ~\new_[8963]_ ;
  assign \new_[3526]_  = ~\new_[3884]_  & ~\new_[8954]_ ;
  assign \new_[3527]_  = ~\new_[3852]_  & ~\new_[8964]_ ;
  assign \new_[3528]_  = ~\new_[3855]_  & ~\new_[8954]_ ;
  assign \new_[3529]_  = ~\new_[6160]_  | ~\new_[3654]_ ;
  assign \new_[3530]_  = ~\new_[6160]_  | ~\new_[3865]_ ;
  assign \new_[3531]_  = ~\new_[8710]_  | ~\new_[3867]_ ;
  assign \new_[3532]_  = (~\new_[4336]_  | ~\new_[8961]_ ) & (~\new_[7112]_  | ~\new_[8964]_ );
  assign \new_[3533]_  = (~\new_[4350]_  | ~\new_[8961]_ ) & (~\new_[7050]_  | ~\new_[8964]_ );
  assign \new_[3534]_  = (~\new_[4238]_  | ~\new_[8961]_ ) & (~\new_[7100]_  | ~\new_[8964]_ );
  assign \new_[3535]_  = (~\new_[4345]_  | ~\new_[8961]_ ) & (~\new_[7148]_  | ~\new_[8962]_ );
  assign \new_[3536]_  = (~\new_[4348]_  | ~\new_[8965]_ ) & (~\new_[7141]_  | ~\new_[8963]_ );
  assign \new_[3537]_  = (~\new_[4338]_  | ~\new_[8961]_ ) & (~\new_[7044]_  | ~\new_[8964]_ );
  assign \new_[3538]_  = (~\new_[4237]_  | ~\new_[8961]_ ) & (~\new_[7052]_  | ~\new_[8964]_ );
  assign \new_[3539]_  = (~\new_[4242]_  | ~\new_[8961]_ ) & (~\new_[7046]_  | ~\new_[8964]_ );
  assign \new_[3540]_  = (~\new_[4349]_  | ~\new_[8961]_ ) & (~\new_[7095]_  | ~\new_[8964]_ );
  assign n3405 = ~\new_[7459]_  | (~\new_[3997]_  & ~\new_[7560]_ );
  assign n3370 = ~\new_[7557]_  | (~\new_[3998]_  & ~\new_[7560]_ );
  assign n3375 = ~\new_[7411]_  | (~\new_[3999]_  & ~\new_[7560]_ );
  assign n3380 = ~\new_[7474]_  | (~\new_[4000]_  & ~\new_[7560]_ );
  assign n3385 = ~\new_[7501]_  | (~\new_[4001]_  & ~\new_[7560]_ );
  assign n3390 = ~\new_[7409]_  | (~\new_[4002]_  & ~\new_[7560]_ );
  assign n3400 = ~\new_[7511]_  | (~\new_[4003]_  & ~\new_[7560]_ );
  assign n3395 = ~\new_[7419]_  | (~\new_[4004]_  & ~\new_[7560]_ );
  assign \new_[3549]_  = ~\new_[3876]_  & (~\new_[7974]_  | ~\new_[7645]_ );
  assign \new_[3550]_  = ~\new_[3877]_  & (~\new_[7969]_  | ~\new_[7645]_ );
  assign \new_[3551]_  = ~\new_[3878]_  & (~\new_[8061]_  | ~\new_[7645]_ );
  assign \new_[3552]_  = ~\new_[3879]_  & (~\new_[8089]_  | ~\new_[7645]_ );
  assign \new_[3553]_  = ~\new_[3880]_  & (~\new_[8042]_  | ~\new_[7499]_ );
  assign \new_[3554]_  = ~\new_[3881]_  & (~\new_[8088]_  | ~\new_[7499]_ );
  assign \new_[3555]_  = ~\new_[3882]_  & (~\new_[8136]_  | ~\new_[7499]_ );
  assign \new_[3556]_  = ~\new_[3883]_  & (~\new_[8082]_  | ~\new_[7499]_ );
  assign \new_[3557]_  = ~\new_[3648]_ ;
  assign \new_[3558]_  = ~\new_[3650]_ ;
  assign \new_[3559]_  = ~\new_[3652]_ ;
  assign \new_[3560]_  = ~\new_[3654]_ ;
  assign \new_[3561]_  = ~\new_[4143]_  & (~\new_[6141]_  | ~\new_[6145]_ );
  assign \new_[3562]_  = ~\new_[3869]_  | (~\new_[6159]_  & ~\new_[2538]_ );
  assign \new_[3563]_  = ~\new_[3870]_  | (~\new_[6147]_  & ~\new_[2539]_ );
  assign \new_[3564]_  = ~\new_[3871]_  | (~\new_[6147]_  & ~\new_[2540]_ );
  assign \new_[3565]_  = ~\new_[3872]_  | (~\new_[6159]_  & ~\new_[2541]_ );
  assign \new_[3566]_  = ~\new_[3873]_  | (~\new_[6159]_  & ~\new_[2542]_ );
  assign \new_[3567]_  = ~\new_[3874]_  | (~\new_[6147]_  & ~\new_[2550]_ );
  assign \new_[3568]_  = ~\new_[3875]_  | (~\new_[6159]_  & ~\new_[2551]_ );
  assign \new_[3569]_  = ~\new_[4143]_  & (~\new_[6142]_  | ~\new_[6146]_ );
  assign \new_[3570]_  = ~\new_[4143]_  & (~\new_[6143]_  | ~\new_[6144]_ );
  assign \new_[3571]_  = ~\new_[3890]_  & (~\new_[8145]_  | ~\new_[7645]_ );
  assign \new_[3572]_  = ~\new_[3891]_  & (~\new_[8030]_  | ~\new_[7645]_ );
  assign \new_[3573]_  = ~\new_[3892]_  & (~\new_[8054]_  | ~\new_[7645]_ );
  assign \new_[3574]_  = ~\new_[3893]_  & (~\new_[8043]_  | ~\new_[7499]_ );
  assign \new_[3575]_  = ~\new_[3894]_  & (~\new_[7992]_  | ~\new_[7499]_ );
  assign \new_[3576]_  = ~\new_[3895]_  & (~\new_[8144]_  | ~\new_[7499]_ );
  assign \new_[3577]_  = ~\new_[3889]_  & (~\new_[8155]_  | ~\new_[7645]_ );
  assign \new_[3578]_  = ~\new_[3896]_  & (~\new_[8110]_  | ~\new_[7499]_ );
  assign \new_[3579]_  = ~\new_[3932]_  & ~\new_[5552]_ ;
  assign \new_[3580]_  = ~\new_[3933]_  & ~\new_[5552]_ ;
  assign \new_[3581]_  = ~\new_[3934]_  & ~\new_[5551]_ ;
  assign \new_[3582]_  = ~\new_[3936]_  & ~\new_[5606]_ ;
  assign \new_[3583]_  = ~\new_[3937]_  & ~\new_[5553]_ ;
  assign \new_[3584]_  = ~\new_[3939]_  & ~\new_[5606]_ ;
  assign \new_[3585]_  = ~\new_[3938]_  & ~\new_[5551]_ ;
  assign \new_[3586]_  = ~\new_[3940]_  & ~\new_[5552]_ ;
  assign \new_[3587]_  = ~\new_[3942]_  & ~\new_[5551]_ ;
  assign \new_[3588]_  = ~\new_[3943]_  & ~\new_[5551]_ ;
  assign \new_[3589]_  = ~\new_[3944]_  & ~\new_[5606]_ ;
  assign \new_[3590]_  = ~\new_[3945]_  & ~\new_[5606]_ ;
  assign \new_[3591]_  = ~\new_[3946]_  & ~\new_[5606]_ ;
  assign \new_[3592]_  = ~\new_[3947]_  & ~\new_[5552]_ ;
  assign \new_[3593]_  = ~\new_[3948]_  & ~\new_[5552]_ ;
  assign \new_[3594]_  = ~\new_[3935]_  & ~\new_[5552]_ ;
  assign \new_[3595]_  = ~\new_[3950]_  & ~\new_[5606]_ ;
  assign \new_[3596]_  = ~\new_[3949]_  & ~\new_[5606]_ ;
  assign \new_[3597]_  = ~\new_[3951]_  & ~\new_[5552]_ ;
  assign \new_[3598]_  = ~\new_[3952]_  & ~\new_[5551]_ ;
  assign \new_[3599]_  = ~\new_[3953]_  & ~\new_[5606]_ ;
  assign \new_[3600]_  = ~\new_[3954]_  & ~\new_[5553]_ ;
  assign \new_[3601]_  = ~\new_[3955]_  & ~\new_[5551]_ ;
  assign \new_[3602]_  = ~\new_[3956]_  & ~\new_[5552]_ ;
  assign \new_[3603]_  = ~\new_[3957]_  & ~\new_[5551]_ ;
  assign \new_[3604]_  = ~\new_[3958]_  & ~\new_[5606]_ ;
  assign \new_[3605]_  = ~\new_[3959]_  & ~\new_[5551]_ ;
  assign \new_[3606]_  = ~\new_[3960]_  & ~\new_[5551]_ ;
  assign \new_[3607]_  = ~\new_[3961]_  & ~\new_[5552]_ ;
  assign \new_[3608]_  = ~\new_[3962]_  & ~\new_[5606]_ ;
  assign \new_[3609]_  = ~\new_[3963]_  & ~\new_[5606]_ ;
  assign \new_[3610]_  = ~\new_[3964]_  & ~\new_[5553]_ ;
  assign \new_[3611]_  = ~\new_[3965]_  & ~\new_[5552]_ ;
  assign \new_[3612]_  = ~\new_[3967]_  & ~\new_[5552]_ ;
  assign \new_[3613]_  = ~\new_[3968]_  & ~\new_[5553]_ ;
  assign \new_[3614]_  = ~\new_[3970]_  | ~\new_[8489]_ ;
  assign \new_[3615]_  = ~\new_[8389]_  | ~\new_[8489]_ ;
  assign \new_[3616]_  = ~\new_[8415]_  | ~\new_[8489]_ ;
  assign \new_[3617]_  = ~\new_[3837]_  & (~\new_[7942]_  | ~\new_[7645]_ );
  assign \new_[3618]_  = ~\new_[3838]_  & (~\new_[8035]_  | ~\new_[7645]_ );
  assign \new_[3619]_  = ~\new_[3840]_  & (~\new_[7985]_  | ~\new_[7645]_ );
  assign \new_[3620]_  = ~\new_[4227]_  & ~\new_[3975]_ ;
  assign \new_[3621]_  = ~\new_[3841]_  & (~\new_[8116]_  | ~\new_[7645]_ );
  assign \new_[3622]_  = ~\new_[4330]_  | ~\new_[3976]_ ;
  assign \new_[3623]_  = \new_[4330]_  | \new_[3975]_ ;
  assign \new_[3624]_  = ~\new_[3974]_  & ~\new_[4135]_ ;
  assign \new_[3625]_  = ~\new_[3842]_  & (~\new_[8092]_  | ~\new_[7499]_ );
  assign \new_[3626]_  = ~\new_[3843]_  & (~\new_[8025]_  | ~\new_[7499]_ );
  assign \new_[3627]_  = ~\new_[3844]_  & (~\new_[8147]_  | ~\new_[7499]_ );
  assign \new_[3628]_  = ~\new_[3845]_  & (~\new_[8133]_  | ~\new_[7499]_ );
  assign \new_[3629]_  = ~\new_[3826]_ ;
  assign \new_[3630]_  = ~\new_[4227]_  | ~\new_[4225]_  | ~\new_[4413]_ ;
  assign \new_[3631]_  = ~\new_[4157]_  | ~\new_[8960]_ ;
  assign \new_[3632]_  = ~\new_[4144]_  | ~\new_[8960]_ ;
  assign \new_[3633]_  = ~\new_[4136]_  | ~\new_[8960]_ ;
  assign n3465 = ~\new_[3984]_  | ~\new_[7344]_ ;
  assign n3460 = ~\new_[3985]_  | ~\new_[7233]_ ;
  assign n3420 = ~\new_[3986]_  | ~\new_[7293]_ ;
  assign n3440 = ~\new_[3987]_  | ~\new_[7362]_ ;
  assign n3425 = ~\new_[3988]_  | ~\new_[7188]_ ;
  assign n3410 = ~\new_[3989]_  | ~\new_[7334]_ ;
  assign n3505 = ~\new_[3990]_  | ~\new_[7253]_ ;
  assign n3490 = ~\new_[3991]_  | ~\new_[7352]_ ;
  assign \new_[3642]_  = (~\new_[4444]_  | ~\new_[8961]_ ) & (~\new_[7111]_  | ~\new_[8963]_ );
  assign n3475 = ~\new_[7440]_  | (~\new_[4167]_  & ~\new_[7560]_ );
  assign n3445 = ~\new_[7457]_  | (~\new_[4170]_  & ~\new_[7560]_ );
  assign n3450 = ~\new_[7556]_  | (~\new_[4175]_  & ~\new_[7560]_ );
  assign n3470 = ~\new_[7532]_  | (~\new_[4176]_  & ~\new_[7560]_ );
  assign \new_[3647]_  = ~\new_[3864]_ ;
  assign \new_[3648]_  = \new_[4997]_  ? \new_[7583]_  : \new_[4178]_ ;
  assign \new_[3649]_  = ~\new_[3865]_ ;
  assign \new_[3650]_  = \new_[4999]_  ? \new_[7583]_  : \new_[4179]_ ;
  assign \new_[3651]_  = ~\new_[3866]_ ;
  assign \new_[3652]_  = \new_[5001]_  ? \new_[7583]_  : \new_[4180]_ ;
  assign \new_[3653]_  = ~\new_[3867]_ ;
  assign \new_[3654]_  = \new_[5003]_  ? \new_[7632]_  : \new_[4181]_ ;
  assign \new_[3655]_  = ~\new_[3992]_  | (~\new_[8710]_  & ~\new_[2658]_ );
  assign \new_[3656]_  = ~\new_[3993]_  | (~\new_[6162]_  & ~\new_[2653]_ );
  assign \new_[3657]_  = ~\new_[3994]_  | (~\new_[8710]_  & ~\new_[2620]_ );
  assign \new_[3658]_  = ~\new_[3995]_  | (~\new_[8710]_  & ~\new_[2630]_ );
  assign \new_[3659]_  = ~\new_[4000]_  & ~\new_[7829]_ ;
  assign \new_[3660]_  = ~\new_[4003]_  & ~\new_[7829]_ ;
  assign \new_[3661]_  = ~\new_[4004]_  & ~\new_[7829]_ ;
  assign \new_[3662]_  = ~\new_[3997]_  & ~\new_[7829]_ ;
  assign \new_[3663]_  = ~\new_[3998]_  & ~\new_[7829]_ ;
  assign \new_[3664]_  = ~\new_[3999]_  & ~\new_[7829]_ ;
  assign \new_[3665]_  = ~\new_[4001]_  & ~\new_[7829]_ ;
  assign \new_[3666]_  = ~\new_[4002]_  & ~\new_[7829]_ ;
  assign \new_[3667]_  = ~\new_[4000]_  & ~\new_[8562]_ ;
  assign \new_[3668]_  = ~\new_[4003]_  & ~\new_[8562]_ ;
  assign \new_[3669]_  = ~\new_[4004]_  & ~\new_[8562]_ ;
  assign \new_[3670]_  = ~\new_[3997]_  & ~\new_[8562]_ ;
  assign \new_[3671]_  = ~\new_[3998]_  & ~\new_[8562]_ ;
  assign \new_[3672]_  = ~\new_[3999]_  & ~\new_[8562]_ ;
  assign \new_[3673]_  = ~\new_[4001]_  & ~\new_[8562]_ ;
  assign \new_[3674]_  = ~\new_[4002]_  & ~\new_[8562]_ ;
  assign \new_[3675]_  = ~\new_[5114]_ ;
  assign n3480 = ~\new_[7543]_  | (~\new_[4182]_  & ~\new_[7560]_ );
  assign n3455 = ~\new_[7432]_  | (~\new_[4183]_  & ~\new_[7560]_ );
  assign n3485 = ~\new_[7485]_  | (~\new_[4184]_  & ~\new_[7560]_ );
  assign n3415 = ~\new_[7429]_  | (~\new_[4185]_  & ~\new_[7560]_ );
  assign \new_[3680]_  = ~\new_[4005]_  | (~\new_[8710]_  & ~\new_[2626]_ );
  assign \new_[3681]_  = ~\new_[4006]_  | (~\new_[8710]_  & ~\new_[2627]_ );
  assign \new_[3682]_  = ~\new_[4007]_  | (~\new_[6162]_  & ~\new_[2617]_ );
  assign \new_[3683]_  = ~\new_[4008]_  | (~\new_[8710]_  & ~\new_[2628]_ );
  assign \new_[3684]_  = ~\new_[4066]_  & ~\new_[5606]_ ;
  assign \new_[3685]_  = ~\new_[4067]_  & ~\new_[5551]_ ;
  assign \new_[3686]_  = ~\new_[4068]_  & ~\new_[5551]_ ;
  assign \new_[3687]_  = ~\new_[4069]_  & ~\new_[5553]_ ;
  assign \new_[3688]_  = ~\new_[4070]_  & ~\new_[5551]_ ;
  assign \new_[3689]_  = ~\new_[4071]_  & ~\new_[5553]_ ;
  assign \new_[3690]_  = ~\new_[4072]_  & ~\new_[5553]_ ;
  assign \new_[3691]_  = ~\new_[4073]_  & ~\new_[5552]_ ;
  assign \new_[3692]_  = ~\new_[4074]_  & ~\new_[5606]_ ;
  assign \new_[3693]_  = ~\new_[4075]_  & ~\new_[5553]_ ;
  assign \new_[3694]_  = ~\new_[4076]_  & ~\new_[5606]_ ;
  assign \new_[3695]_  = ~\new_[4078]_  & ~\new_[5553]_ ;
  assign \new_[3696]_  = ~\new_[4077]_  & ~\new_[5552]_ ;
  assign \new_[3697]_  = ~\new_[4079]_  & ~\new_[5551]_ ;
  assign \new_[3698]_  = ~\new_[4080]_  & ~\new_[5606]_ ;
  assign \new_[3699]_  = ~\new_[4081]_  & ~\new_[5606]_ ;
  assign \new_[3700]_  = ~\new_[4082]_  & ~\new_[5553]_ ;
  assign \new_[3701]_  = ~\new_[4084]_  & ~\new_[5606]_ ;
  assign \new_[3702]_  = ~\new_[4083]_  & ~\new_[5553]_ ;
  assign \new_[3703]_  = ~\new_[4085]_  & ~\new_[5552]_ ;
  assign \new_[3704]_  = ~\new_[4086]_  & ~\new_[5553]_ ;
  assign \new_[3705]_  = ~\new_[4087]_  & ~\new_[5553]_ ;
  assign \new_[3706]_  = ~\new_[4088]_  & ~\new_[5606]_ ;
  assign \new_[3707]_  = ~\new_[4089]_  & ~\new_[5551]_ ;
  assign \new_[3708]_  = ~\new_[4090]_  & ~\new_[5551]_ ;
  assign \new_[3709]_  = ~\new_[4091]_  & ~\new_[5553]_ ;
  assign \new_[3710]_  = ~\new_[4094]_  & ~\new_[5553]_ ;
  assign \new_[3711]_  = ~\new_[4092]_  & ~\new_[5552]_ ;
  assign \new_[3712]_  = ~\new_[4093]_  & ~\new_[5552]_ ;
  assign \new_[3713]_  = ~\new_[4095]_  & ~\new_[5551]_ ;
  assign \new_[3714]_  = ~\new_[4096]_  & ~\new_[5606]_ ;
  assign \new_[3715]_  = ~\new_[4097]_  & ~\new_[5552]_ ;
  assign \new_[3716]_  = ~\new_[4098]_  & ~\new_[5606]_ ;
  assign \new_[3717]_  = ~\new_[4099]_  & ~\new_[5551]_ ;
  assign \new_[3718]_  = ~\new_[4100]_  & ~\new_[5551]_ ;
  assign \new_[3719]_  = ~\new_[4101]_  & ~\new_[5551]_ ;
  assign \new_[3720]_  = ~\new_[4102]_  & ~\new_[5606]_ ;
  assign \new_[3721]_  = ~\new_[4103]_  & ~\new_[5551]_ ;
  assign \new_[3722]_  = ~\new_[4112]_  & ~\new_[5551]_ ;
  assign \new_[3723]_  = ~\new_[4104]_  & ~\new_[5553]_ ;
  assign \new_[3724]_  = ~\new_[4105]_  & ~\new_[5552]_ ;
  assign \new_[3725]_  = ~\new_[4106]_  & ~\new_[5553]_ ;
  assign \new_[3726]_  = ~\new_[4108]_  & ~\new_[5551]_ ;
  assign \new_[3727]_  = ~\new_[4107]_  & ~\new_[5552]_ ;
  assign \new_[3728]_  = ~\new_[4109]_  & ~\new_[5551]_ ;
  assign \new_[3729]_  = ~\new_[4110]_  & ~\new_[5553]_ ;
  assign \new_[3730]_  = ~\new_[4111]_  & ~\new_[5606]_ ;
  assign \new_[3731]_  = ~\new_[4114]_  & ~\new_[5551]_ ;
  assign \new_[3732]_  = ~\new_[4115]_  & ~\new_[5553]_ ;
  assign \new_[3733]_  = ~\new_[4116]_  & ~\new_[5552]_ ;
  assign \new_[3734]_  = ~\new_[4113]_  & ~\new_[5551]_ ;
  assign \new_[3735]_  = ~\new_[4117]_  & ~\new_[5606]_ ;
  assign \new_[3736]_  = ~\new_[4118]_  & ~\new_[5553]_ ;
  assign \new_[3737]_  = ~\new_[4119]_  & ~\new_[5606]_ ;
  assign \new_[3738]_  = ~\new_[4120]_  & ~\new_[5553]_ ;
  assign \new_[3739]_  = ~\new_[4121]_  & ~\new_[5553]_ ;
  assign \new_[3740]_  = ~\new_[4122]_  & ~\new_[5553]_ ;
  assign \new_[3741]_  = \key_i[63]  ^ \new_[4187]_ ;
  assign \new_[3742]_  = \key_i[6]  ^ \new_[4188]_ ;
  assign \new_[3743]_  = \key_i[25]  ^ \new_[4189]_ ;
  assign \new_[3744]_  = \key_i[76]  ^ \new_[4190]_ ;
  assign \new_[3745]_  = \key_i[77]  ^ \new_[4191]_ ;
  assign \new_[3746]_  = \key_i[26]  ^ \new_[4192]_ ;
  assign \new_[3747]_  = \key_i[78]  ^ \new_[4193]_ ;
  assign \new_[3748]_  = \key_i[79]  ^ \new_[4194]_ ;
  assign \new_[3749]_  = \key_i[29]  ^ \new_[4195]_ ;
  assign \new_[3750]_  = \key_i[8]  ^ \new_[4196]_ ;
  assign \new_[3751]_  = \key_i[105]  ^ \new_[4197]_ ;
  assign \new_[3752]_  = \key_i[106]  ^ \new_[4198]_ ;
  assign \new_[3753]_  = \key_i[122]  ^ \new_[4199]_ ;
  assign \new_[3754]_  = \key_i[3]  ^ \new_[4200]_ ;
  assign \new_[3755]_  = \key_i[0]  ^ \new_[4201]_ ;
  assign \new_[3756]_  = \key_i[123]  ^ \new_[4202]_ ;
  assign \new_[3757]_  = \key_i[107]  ^ \new_[4204]_ ;
  assign \new_[3758]_  = \key_i[41]  ^ \new_[4203]_ ;
  assign \new_[3759]_  = ~\new_[3972]_ ;
  assign \new_[3760]_  = \key_i[42]  ^ \new_[4205]_ ;
  assign \new_[3761]_  = \key_i[126]  ^ \new_[4211]_ ;
  assign \new_[3762]_  = \key_i[43]  ^ \new_[4206]_ ;
  assign \new_[3763]_  = \key_i[44]  ^ \new_[4207]_ ;
  assign \new_[3764]_  = \key_i[125]  ^ \new_[4208]_ ;
  assign \new_[3765]_  = \key_i[46]  ^ \new_[4210]_ ;
  assign \new_[3766]_  = \key_i[47]  ^ \new_[4212]_ ;
  assign \new_[3767]_  = \key_i[108]  ^ \new_[4209]_ ;
  assign \new_[3768]_  = \key_i[127]  ^ \new_[4213]_ ;
  assign \new_[3769]_  = \key_i[13]  ^ \new_[4214]_ ;
  assign \new_[3770]_  = \key_i[10]  ^ \new_[4215]_ ;
  assign \new_[3771]_  = \key_i[110]  ^ \new_[4216]_ ;
  assign \new_[3772]_  = \key_i[57]  ^ \new_[4217]_ ;
  assign \new_[3773]_  = \key_i[58]  ^ \new_[4218]_ ;
  assign \new_[3774]_  = \key_i[59]  ^ \new_[4219]_ ;
  assign \new_[3775]_  = \key_i[5]  ^ \new_[4220]_ ;
  assign \new_[3776]_  = \key_i[111]  ^ \new_[4221]_ ;
  assign \new_[3777]_  = \key_i[60]  ^ \new_[4222]_ ;
  assign \new_[3778]_  = \new_[7984]_  ^ \new_[4221]_ ;
  assign \new_[3779]_  = \new_[7941]_  ^ \new_[4187]_ ;
  assign \new_[3780]_  = \new_[1963]_  ^ \new_[4188]_ ;
  assign \new_[3781]_  = \new_[1125]_  ^ \new_[4190]_ ;
  assign \new_[3782]_  = \new_[1952]_  ^ \new_[4189]_ ;
  assign \new_[3783]_  = \new_[1132]_  ^ \new_[4191]_ ;
  assign \new_[3784]_  = \new_[1133]_  ^ \new_[4193]_ ;
  assign \new_[3785]_  = \new_[1955]_  ^ \new_[4192]_ ;
  assign \new_[3786]_  = \new_[1141]_  ^ \new_[4194]_ ;
  assign \new_[3787]_  = ~\new_[3941]_ ;
  assign \new_[3788]_  = \new_[1947]_  ^ \new_[4195]_ ;
  assign \new_[3789]_  = \new_[1070]_  ^ \new_[4196]_ ;
  assign \new_[3790]_  = \new_[7986]_  ^ \new_[4197]_ ;
  assign \new_[3791]_  = \new_[1960]_  ^ \new_[4200]_ ;
  assign \new_[3792]_  = \new_[2273]_  ^ \new_[4199]_ ;
  assign \new_[3793]_  = \new_[8075]_  ^ \new_[4198]_ ;
  assign \new_[3794]_  = \new_[1119]_  ^ \new_[4203]_ ;
  assign \new_[3795]_  = \new_[2197]_  ^ \new_[4202]_ ;
  assign \new_[3796]_  = \new_[1118]_  ^ \new_[4205]_ ;
  assign \new_[3797]_  = \new_[1079]_  ^ \new_[4206]_ ;
  assign \new_[3798]_  = \new_[7971]_  ^ \new_[4204]_ ;
  assign \new_[3799]_  = \new_[1080]_  ^ \new_[4207]_ ;
  assign \new_[3800]_  = \new_[2196]_  ^ \new_[4208]_ ;
  assign \new_[3801]_  = \new_[1083]_  ^ \new_[4210]_ ;
  assign \new_[3802]_  = \new_[8004]_  ^ \new_[4209]_ ;
  assign \new_[3803]_  = \new_[1084]_  ^ \new_[4212]_ ;
  assign \new_[3804]_  = \new_[2271]_  ^ \new_[4211]_ ;
  assign \new_[3805]_  = \new_[2266]_  ^ \new_[4213]_ ;
  assign \new_[3806]_  = \new_[1063]_  ^ \new_[4214]_ ;
  assign \new_[3807]_  = \new_[1072]_  ^ \new_[4215]_ ;
  assign \new_[3808]_  = \new_[1964]_  ^ \new_[4201]_ ;
  assign \new_[3809]_  = \new_[8124]_  ^ \new_[4217]_ ;
  assign \new_[3810]_  = \new_[8055]_  ^ \new_[4218]_ ;
  assign \new_[3811]_  = \new_[1455]_  ^ \new_[4216]_ ;
  assign \new_[3812]_  = \new_[7957]_  ^ \new_[4219]_ ;
  assign \new_[3813]_  = \new_[1962]_  ^ \new_[4220]_ ;
  assign \new_[3814]_  = \new_[8028]_  ^ \new_[4222]_ ;
  assign \new_[3815]_  = ~\new_[4223]_  | ~\new_[4422]_  | ~\new_[4466]_ ;
  assign \new_[3816]_  = ~\new_[4123]_  & (~\new_[4512]_  | ~\new_[7631]_ );
  assign n3430 = ~\new_[7463]_  | (~\new_[4150]_  & ~\new_[7560]_ );
  assign n3435 = ~\new_[7453]_  | (~\new_[4151]_  & ~\new_[7560]_ );
  assign n3495 = ~\new_[7452]_  | (~\new_[4152]_  & ~\new_[7560]_ );
  assign n3500 = ~\new_[7509]_  | (~\new_[4156]_  & ~\new_[7560]_ );
  assign \new_[3821]_  = (~\new_[4159]_  | ~\new_[8713]_ ) & (~\new_[7983]_  | ~\new_[8716]_ );
  assign \new_[3822]_  = (~\new_[4160]_  | ~\new_[8713]_ ) & (~\new_[8073]_  | ~\new_[8716]_ );
  assign \new_[3823]_  = (~\new_[4161]_  | ~\new_[8713]_ ) & (~\new_[8149]_  | ~\new_[8716]_ );
  assign \new_[3824]_  = (~\new_[4162]_  | ~\new_[7825]_ ) & (~\new_[8069]_  | ~\new_[8716]_ );
  assign \new_[3825]_  = ~\new_[4331]_  & ~\new_[4135]_ ;
  assign \new_[3826]_  = ~\new_[4135]_  | ~\new_[3980]_ ;
  assign \new_[3827]_  = ~\new_[4130]_  | (~\new_[6162]_  & ~\new_[2660]_ );
  assign \new_[3828]_  = ~\new_[4131]_  | (~\new_[6162]_  & ~\new_[2659]_ );
  assign \new_[3829]_  = ~\new_[3978]_  | (~\new_[6162]_  & ~\new_[2618]_ );
  assign \new_[3830]_  = ~\new_[3979]_  | (~\new_[6147]_  & ~\new_[2619]_ );
  assign \new_[3831]_  = ~\new_[4124]_  & (~\new_[4332]_  | ~\new_[6895]_ );
  assign \new_[3832]_  = ~\new_[4125]_  & (~\new_[4332]_  | ~\new_[6896]_ );
  assign \new_[3833]_  = ~\new_[4126]_  & (~\new_[4332]_  | ~\new_[6897]_ );
  assign \new_[3834]_  = ~\new_[4127]_  & (~\new_[4332]_  | ~\new_[7145]_ );
  assign \new_[3835]_  = ~\new_[4128]_  & (~\new_[4332]_  | ~\new_[7089]_ );
  assign \new_[3836]_  = ~\new_[4129]_  & (~\new_[4332]_  | ~\new_[6894]_ );
  assign \new_[3837]_  = ~\new_[4156]_  & ~\new_[7829]_ ;
  assign \new_[3838]_  = ~\new_[4150]_  & ~\new_[7829]_ ;
  assign \new_[3839]_  = \new_[4413]_  & \new_[4330]_ ;
  assign \new_[3840]_  = ~\new_[4151]_  & ~\new_[7829]_ ;
  assign \new_[3841]_  = ~\new_[4152]_  & ~\new_[7829]_ ;
  assign \new_[3842]_  = ~\new_[4156]_  & ~\new_[8562]_ ;
  assign \new_[3843]_  = ~\new_[4150]_  & ~\new_[8562]_ ;
  assign \new_[3844]_  = ~\new_[4151]_  & ~\new_[8562]_ ;
  assign \new_[3845]_  = ~\new_[4152]_  & ~\new_[8562]_ ;
  assign \new_[3846]_  = \\mix1_data_o_reg_reg[7] ;
  assign \new_[3847]_  = (~\key_i[49]  | ~\new_[4798]_ ) & (~\new_[8141]_  | ~\new_[8726]_ );
  assign \new_[3848]_  = (~\key_i[53]  | ~\new_[4798]_ ) & (~\new_[7993]_  | ~\new_[8726]_ );
  assign \new_[3849]_  = (~\key_i[54]  | ~\new_[4798]_ ) & (~\new_[8122]_  | ~\new_[8726]_ );
  assign \new_[3850]_  = (~\key_i[56]  | ~\new_[4798]_ ) & (~\new_[8000]_  | ~\new_[8726]_ );
  assign \new_[3851]_  = (~\key_i[57]  | ~\new_[4798]_ ) & (~\new_[8124]_  | ~\new_[8726]_ );
  assign \new_[3852]_  = (~\key_i[58]  | ~\new_[4798]_ ) & (~\new_[8055]_  | ~\new_[8726]_ );
  assign \new_[3853]_  = (~\key_i[59]  | ~\new_[4798]_ ) & (~\new_[7957]_  | ~\new_[8726]_ );
  assign \new_[3854]_  = (~\key_i[60]  | ~\new_[4798]_ ) & (~\new_[8028]_  | ~\new_[8726]_ );
  assign \new_[3855]_  = (~\key_i[61]  | ~\new_[4798]_ ) & (~\new_[8001]_  | ~\new_[8726]_ );
  assign \new_[3856]_  = (~\key_i[34]  | ~\new_[4798]_ ) & (~\new_[7980]_  | ~\new_[8726]_ );
  assign \new_[3857]_  = \\mix1_data_o_reg_reg[23] ;
  assign \new_[3858]_  = \key_i[36]  ? \new_[5114]_  : \new_[5603]_ ;
  assign \new_[3859]_  = \key_i[38]  ? \new_[5114]_  : \new_[5601]_ ;
  assign \new_[3860]_  = \key_i[39]  ? \new_[5114]_  : \new_[5605]_ ;
  assign \new_[3861]_  = \key_i[40]  ? \new_[5114]_  : \new_[5602]_ ;
  assign \new_[3862]_  = \key_i[41]  ? \new_[5114]_  : \new_[5604]_ ;
  assign \new_[3863]_  = \\mix1_data_o_reg_reg[31] ;
  assign \new_[3864]_  = \new_[5129]_  ? \new_[7583]_  : \new_[4276]_ ;
  assign \new_[3865]_  = \new_[5132]_  ? \new_[7632]_  : \new_[4277]_ ;
  assign \new_[3866]_  = \new_[5135]_  ? \new_[7583]_  : \new_[4278]_ ;
  assign \new_[3867]_  = \new_[5138]_  ? \new_[7632]_  : \new_[4279]_ ;
  assign \new_[3868]_  = (~\key_i[45]  | ~\new_[4798]_ ) & (~\new_[1082]_  | ~\new_[8726]_ );
  assign \new_[3869]_  = ~\new_[6161]_  | ~\new_[4177]_ ;
  assign \new_[3870]_  = ~\new_[6161]_  | ~\new_[4166]_ ;
  assign \new_[3871]_  = ~\new_[6162]_  | ~\new_[4169]_ ;
  assign \new_[3872]_  = ~\new_[6162]_  | ~\new_[4168]_ ;
  assign \new_[3873]_  = ~\new_[6162]_  | ~\new_[4171]_ ;
  assign \new_[3874]_  = ~\new_[6162]_  | ~\new_[4172]_ ;
  assign \new_[3875]_  = ~\new_[6162]_  | ~\new_[4174]_ ;
  assign \new_[3876]_  = ~\new_[4176]_  & ~\new_[7829]_ ;
  assign \new_[3877]_  = ~\new_[4167]_  & ~\new_[7829]_ ;
  assign \new_[3878]_  = ~\new_[4170]_  & ~\new_[7829]_ ;
  assign \new_[3879]_  = ~\new_[4175]_  & ~\new_[7829]_ ;
  assign \new_[3880]_  = ~\new_[4176]_  & ~\new_[8562]_ ;
  assign \new_[3881]_  = ~\new_[4167]_  & ~\new_[8562]_ ;
  assign \new_[3882]_  = ~\new_[4170]_  & ~\new_[8562]_ ;
  assign \new_[3883]_  = ~\new_[4175]_  & ~\new_[8562]_ ;
  assign \new_[3884]_  = (~\key_i[46]  | ~\new_[4798]_ ) & (~\new_[1083]_  | ~\new_[8726]_ );
  assign \new_[3885]_  = \\mix1_data_o_reg_reg[15] ;
  assign \new_[3886]_  = ~\new_[5114]_ ;
  assign \new_[3887]_  = ~\new_[5114]_ ;
  assign \new_[3888]_  = ~\new_[5114]_ ;
  assign \new_[3889]_  = ~\new_[4182]_  & ~\new_[7829]_ ;
  assign \new_[3890]_  = ~\new_[4185]_  & ~\new_[7829]_ ;
  assign \new_[3891]_  = ~\new_[4183]_  & ~\new_[7829]_ ;
  assign \new_[3892]_  = ~\new_[4184]_  & ~\new_[7829]_ ;
  assign \new_[3893]_  = ~\new_[4182]_  & ~\new_[8562]_ ;
  assign \new_[3894]_  = ~\new_[4185]_  & ~\new_[8562]_ ;
  assign \new_[3895]_  = ~\new_[4183]_  & ~\new_[8562]_ ;
  assign \new_[3896]_  = ~\new_[4184]_  & ~\new_[8562]_ ;
  assign \new_[3897]_  = \key_i[61]  ^ \new_[4285]_ ;
  assign \new_[3898]_  = \key_i[62]  ^ \new_[4286]_ ;
  assign \new_[3899]_  = \key_i[1]  ^ \new_[4287]_ ;
  assign \new_[3900]_  = \key_i[72]  ^ \new_[4288]_ ;
  assign \new_[3901]_  = \key_i[73]  ^ \new_[4289]_ ;
  assign \new_[3902]_  = \key_i[24]  ^ \new_[4290]_ ;
  assign \new_[3903]_  = \key_i[74]  ^ \new_[4291]_ ;
  assign \new_[3904]_  = \key_i[75]  ^ \new_[4292]_ ;
  assign \new_[3905]_  = \key_i[27]  ^ \new_[4293]_ ;
  assign \new_[3906]_  = \key_i[7]  ^ \new_[4294]_ ;
  assign \new_[3907]_  = \key_i[28]  ^ \new_[4295]_ ;
  assign \new_[3908]_  = \key_i[2]  ^ \new_[4296]_ ;
  assign \new_[3909]_  = \key_i[30]  ^ \new_[4297]_ ;
  assign \new_[3910]_  = \key_i[104]  ^ \new_[4298]_ ;
  assign \new_[3911]_  = \key_i[31]  ^ \new_[4299]_ ;
  assign \new_[3912]_  = \key_i[90]  ^ \new_[4300]_ ;
  assign \new_[3913]_  = \key_i[91]  ^ \new_[4302]_ ;
  assign \new_[3914]_  = \key_i[92]  ^ \new_[4303]_ ;
  assign \new_[3915]_  = \key_i[11]  ^ \new_[4304]_ ;
  assign \new_[3916]_  = \key_i[93]  ^ \new_[4305]_ ;
  assign \new_[3917]_  = \key_i[34]  ^ \new_[4306]_ ;
  assign \new_[3918]_  = \key_i[94]  ^ \new_[4307]_ ;
  assign \new_[3919]_  = \key_i[95]  ^ \new_[4308]_ ;
  assign \new_[3920]_  = \key_i[120]  ^ \new_[4309]_ ;
  assign \new_[3921]_  = \key_i[121]  ^ \new_[4311]_ ;
  assign \new_[3922]_  = \key_i[9]  ^ \new_[4310]_ ;
  assign \new_[3923]_  = \key_i[40]  ^ \new_[4301]_ ;
  assign \new_[3924]_  = \key_i[124]  ^ \new_[4312]_ ;
  assign \new_[3925]_  = \key_i[45]  ^ \new_[4313]_ ;
  assign \new_[3926]_  = \key_i[109]  ^ \new_[4314]_ ;
  assign \new_[3927]_  = \key_i[4]  ^ \new_[4315]_ ;
  assign \new_[3928]_  = \key_i[12]  ^ \new_[4316]_ ;
  assign \new_[3929]_  = \key_i[14]  ^ \new_[4317]_ ;
  assign \new_[3930]_  = \key_i[15]  ^ \new_[4318]_ ;
  assign \new_[3931]_  = \key_i[56]  ^ \new_[4319]_ ;
  assign \new_[3932]_  = \new_[8001]_  ^ \new_[4285]_ ;
  assign \new_[3933]_  = \new_[8005]_  ^ \new_[4286]_ ;
  assign \new_[3934]_  = \new_[1965]_  ^ \new_[4287]_ ;
  assign \new_[3935]_  = \new_[2043]_  ^ \new_[4302]_ ;
  assign \new_[3936]_  = \new_[1140]_  ^ \new_[4288]_ ;
  assign \new_[3937]_  = \new_[8119]_  ^ \new_[4289]_ ;
  assign \new_[3938]_  = \new_[8130]_  ^ \new_[4291]_ ;
  assign \new_[3939]_  = \new_[1950]_  ^ \new_[4290]_ ;
  assign \new_[3940]_  = \new_[1126]_  ^ \new_[4292]_ ;
  assign \new_[3941]_  = (~\key_i[63]  | ~\new_[4798]_ ) & (~\new_[7941]_  | ~\new_[8726]_ );
  assign \new_[3942]_  = \new_[1969]_  ^ \new_[4294]_ ;
  assign \new_[3943]_  = \new_[1946]_  ^ \new_[4293]_ ;
  assign \new_[3944]_  = \new_[1942]_  ^ \new_[4295]_ ;
  assign \new_[3945]_  = \new_[1959]_  ^ \new_[4296]_ ;
  assign \new_[3946]_  = \new_[1949]_  ^ \new_[4297]_ ;
  assign \new_[3947]_  = \new_[1951]_  ^ \new_[4299]_ ;
  assign \new_[3948]_  = \new_[8037]_  ^ \new_[4300]_ ;
  assign \new_[3949]_  = \new_[8151]_  ^ \new_[4303]_ ;
  assign \new_[3950]_  = \new_[7949]_  ^ \new_[4298]_ ;
  assign \new_[3951]_  = \new_[8094]_  ^ \new_[4305]_ ;
  assign \new_[3952]_  = \new_[2068]_  ^ \new_[4307]_ ;
  assign \new_[3953]_  = \new_[7980]_  ^ \new_[4306]_ ;
  assign \new_[3954]_  = \new_[1061]_  ^ \new_[4304]_ ;
  assign \new_[3955]_  = \new_[2069]_  ^ \new_[4308]_ ;
  assign \new_[3956]_  = \new_[2264]_  ^ \new_[4309]_ ;
  assign \new_[3957]_  = \new_[1076]_  ^ \new_[4310]_ ;
  assign \new_[3958]_  = \new_[2265]_  ^ \new_[4311]_ ;
  assign \new_[3959]_  = \new_[1089]_  ^ \new_[4301]_ ;
  assign \new_[3960]_  = \new_[2131]_  ^ \new_[4312]_ ;
  assign \new_[3961]_  = \new_[1082]_  ^ \new_[4313]_ ;
  assign \new_[3962]_  = \new_[1961]_  ^ \new_[4315]_ ;
  assign \new_[3963]_  = \new_[1062]_  ^ \new_[4316]_ ;
  assign \new_[3964]_  = \new_[1456]_  ^ \new_[4314]_ ;
  assign \new_[3965]_  = \new_[1064]_  ^ \new_[4317]_ ;
  assign \new_[3966]_  = (~\key_i[47]  | ~\new_[4798]_ ) & (~\new_[1084]_  | ~\new_[8726]_ );
  assign \new_[3967]_  = \new_[8000]_  ^ \new_[4319]_ ;
  assign \new_[3968]_  = \new_[1065]_  ^ \new_[4318]_ ;
  assign \new_[3969]_  = ~\new_[4427]_  | ~\new_[4429]_  | ~\new_[4328]_  | ~\new_[4426]_ ;
  assign \new_[3970]_  = ~\new_[4428]_  | ~\new_[4424]_  | ~\new_[4425]_  | ~\new_[4423]_ ;
  assign \new_[3971]_  = ~\new_[4143]_  & (~\new_[6565]_  | ~\new_[6216]_ );
  assign \new_[3972]_  = (~\key_i[62]  | ~\new_[4798]_ ) & (~\new_[8005]_  | ~\new_[8726]_ );
  assign \new_[3973]_  = ~\new_[4163]_  & (~\new_[4226]_  | ~\new_[8961]_ );
  assign \new_[3974]_  = ~\new_[4227]_  | ~\new_[4132]_ ;
  assign \new_[3975]_  = ~\new_[4135]_  | ~\new_[4132]_ ;
  assign \new_[3976]_  = ~\new_[4135]_  & ~\new_[4133]_ ;
  assign \new_[3977]_  = ~\new_[4224]_  & (~\new_[4332]_  | ~\new_[7147]_ );
  assign \new_[3978]_  = ~\new_[6160]_  | ~\new_[4241]_ ;
  assign \new_[3979]_  = ~\new_[6161]_  | ~\new_[4244]_ ;
  assign \new_[3980]_  = ~\new_[4133]_ ;
  assign \new_[3981]_  = \\addroundkey_round_reg[1] ;
  assign \new_[3982]_  = \\addroundkey_round_reg[3] ;
  assign \new_[3983]_  = ~\new_[4143]_ ;
  assign \new_[3984]_  = ~\new_[4263]_  & (~\new_[8059]_  | ~\new_[7645]_ );
  assign \new_[3985]_  = ~\new_[4264]_  & (~\new_[8087]_  | ~\new_[7645]_ );
  assign \new_[3986]_  = ~\new_[4265]_  & (~\new_[8132]_  | ~\new_[7645]_ );
  assign \new_[3987]_  = ~\new_[4266]_  & (~\new_[7645]_  | ~\new_[8080]_ );
  assign \new_[3988]_  = ~\new_[4267]_  & (~\new_[8127]_  | ~\new_[7499]_ );
  assign \new_[3989]_  = ~\new_[4268]_  & (~\new_[7956]_  | ~\new_[7499]_ );
  assign \new_[3990]_  = ~\new_[4269]_  & (~\new_[8152]_  | ~\new_[7499]_ );
  assign \new_[3991]_  = ~\new_[4270]_  & (~\new_[7499]_  | ~\new_[8104]_ );
  assign \new_[3992]_  = ~\new_[6161]_  | ~\new_[4275]_ ;
  assign \new_[3993]_  = ~\new_[6161]_  | ~\new_[4272]_ ;
  assign \new_[3994]_  = ~\new_[6162]_  | ~\new_[4273]_ ;
  assign \new_[3995]_  = ~\new_[6160]_  | ~\new_[4274]_ ;
  assign \new_[3996]_  = \\addroundkey_round_reg[2] ;
  assign \new_[3997]_  = ~\new_[4166]_ ;
  assign \new_[3998]_  = ~\new_[4169]_ ;
  assign \new_[3999]_  = ~\new_[4168]_ ;
  assign \new_[4000]_  = ~\new_[4172]_ ;
  assign \new_[4001]_  = ~\new_[4171]_ ;
  assign \new_[4002]_  = ~\new_[4173]_ ;
  assign \new_[4003]_  = ~\new_[4174]_ ;
  assign \new_[4004]_  = ~\new_[4177]_ ;
  assign \new_[4005]_  = ~\new_[6162]_  | ~\new_[4284]_ ;
  assign \new_[4006]_  = ~\new_[8710]_  | ~\new_[4282]_ ;
  assign \new_[4007]_  = ~\new_[6160]_  | ~\new_[4283]_ ;
  assign \new_[4008]_  = ~\new_[8710]_  | ~\new_[4281]_ ;
  assign \new_[4009]_  = \key_i[19]  ^ \new_[4363]_ ;
  assign \new_[4010]_  = \key_i[112]  ^ \new_[4364]_ ;
  assign \new_[4011]_  = \key_i[64]  ^ \new_[4365]_ ;
  assign \new_[4012]_  = \key_i[101]  ^ \new_[4366]_ ;
  assign \new_[4013]_  = \key_i[65]  ^ \new_[4367]_ ;
  assign \new_[4014]_  = \key_i[66]  ^ \new_[4368]_ ;
  assign \new_[4015]_  = \key_i[20]  ^ \new_[4369]_ ;
  assign \new_[4016]_  = \key_i[113]  ^ \new_[4371]_ ;
  assign \new_[4017]_  = \key_i[67]  ^ \new_[4370]_ ;
  assign \new_[4018]_  = \key_i[68]  ^ \new_[4372]_ ;
  assign \new_[4019]_  = \key_i[21]  ^ \new_[4373]_ ;
  assign \new_[4020]_  = \key_i[69]  ^ \new_[4374]_ ;
  assign \new_[4021]_  = \key_i[22]  ^ \new_[4375]_ ;
  assign \new_[4022]_  = \key_i[70]  ^ \new_[4376]_ ;
  assign \new_[4023]_  = \key_i[114]  ^ \new_[4377]_ ;
  assign \new_[4024]_  = \key_i[71]  ^ \new_[4378]_ ;
  assign \new_[4025]_  = \key_i[23]  ^ \new_[4379]_ ;
  assign \new_[4026]_  = \key_i[102]  ^ \new_[4381]_ ;
  assign \new_[4027]_  = \key_i[115]  ^ \new_[4380]_ ;
  assign \new_[4028]_  = \key_i[116]  ^ \new_[4382]_ ;
  assign \new_[4029]_  = \key_i[103]  ^ \new_[4383]_ ;
  assign \new_[4030]_  = \key_i[80]  ^ \new_[4384]_ ;
  assign \new_[4031]_  = \key_i[81]  ^ \new_[4385]_ ;
  assign \new_[4032]_  = \key_i[117]  ^ \new_[4386]_ ;
  assign \new_[4033]_  = \key_i[82]  ^ \new_[4387]_ ;
  assign \new_[4034]_  = \key_i[83]  ^ \new_[4388]_ ;
  assign \new_[4035]_  = \key_i[84]  ^ \new_[4389]_ ;
  assign \new_[4036]_  = \key_i[118]  ^ \new_[4391]_ ;
  assign \new_[4037]_  = \key_i[85]  ^ \new_[4390]_ ;
  assign \new_[4038]_  = \key_i[86]  ^ \new_[4392]_ ;
  assign \new_[4039]_  = \key_i[87]  ^ \new_[4393]_ ;
  assign \new_[4040]_  = \key_i[88]  ^ \new_[4394]_ ;
  assign \new_[4041]_  = \key_i[89]  ^ \new_[4395]_ ;
  assign \new_[4042]_  = \key_i[119]  ^ \new_[4396]_ ;
  assign \new_[4043]_  = \key_i[32]  ^ \new_[4397]_ ;
  assign \new_[4044]_  = \key_i[33]  ^ \new_[4398]_ ;
  assign \new_[4045]_  = \key_i[35]  ^ \new_[4399]_ ;
  assign \new_[4046]_  = \key_i[96]  ^ \new_[4400]_ ;
  assign \new_[4047]_  = \key_i[97]  ^ \new_[4401]_ ;
  assign \new_[4048]_  = \key_i[36]  ^ \new_[4402]_ ;
  assign \new_[4049]_  = \key_i[98]  ^ \new_[4403]_ ;
  assign \new_[4050]_  = \key_i[99]  ^ \new_[4404]_ ;
  assign \new_[4051]_  = \key_i[37]  ^ \new_[4405]_ ;
  assign \new_[4052]_  = \key_i[38]  ^ \new_[4406]_ ;
  assign \new_[4053]_  = \key_i[39]  ^ \new_[4407]_ ;
  assign \new_[4054]_  = \key_i[48]  ^ \new_[4408]_ ;
  assign \new_[4055]_  = \key_i[49]  ^ \new_[4409]_ ;
  assign \new_[4056]_  = \key_i[50]  ^ \new_[4410]_ ;
  assign \new_[4057]_  = \key_i[51]  ^ \new_[4411]_ ;
  assign \new_[4058]_  = \key_i[52]  ^ \new_[4412]_ ;
  assign \new_[4059]_  = \key_i[53]  ^ \new_[4414]_ ;
  assign \new_[4060]_  = \key_i[54]  ^ \new_[4415]_ ;
  assign \new_[4061]_  = \key_i[55]  ^ \new_[4416]_ ;
  assign \new_[4062]_  = \key_i[16]  ^ \new_[4417]_ ;
  assign \new_[4063]_  = \key_i[100]  ^ \new_[4418]_ ;
  assign \new_[4064]_  = \key_i[17]  ^ \new_[4419]_ ;
  assign \new_[4065]_  = \key_i[18]  ^ \new_[4420]_ ;
  assign \new_[4066]_  = \new_[1980]_  ^ \new_[4420]_ ;
  assign \new_[4067]_  = \new_[2350]_  ^ \new_[4418]_ ;
  assign \new_[4068]_  = \new_[1979]_  ^ \new_[4363]_ ;
  assign \new_[4069]_  = \new_[2132]_  ^ \new_[4365]_ ;
  assign \new_[4070]_  = \new_[2133]_  ^ \new_[4367]_ ;
  assign \new_[4071]_  = \new_[2421]_  ^ \new_[4364]_ ;
  assign \new_[4072]_  = \new_[2135]_  ^ \new_[4368]_ ;
  assign \new_[4073]_  = \new_[2134]_  ^ \new_[4370]_ ;
  assign \new_[4074]_  = \new_[1993]_  ^ \new_[4369]_ ;
  assign \new_[4075]_  = \new_[2136]_  ^ \new_[4372]_ ;
  assign \new_[4076]_  = \new_[2095]_  ^ \new_[4374]_ ;
  assign \new_[4077]_  = \new_[1981]_  ^ \new_[4373]_ ;
  assign \new_[4078]_  = \new_[2411]_  ^ \new_[4371]_ ;
  assign \new_[4079]_  = \new_[2351]_  ^ \new_[4366]_ ;
  assign \new_[4080]_  = \new_[2137]_  ^ \new_[4376]_ ;
  assign \new_[4081]_  = \new_[1982]_  ^ \new_[4375]_ ;
  assign \new_[4082]_  = \new_[2138]_  ^ \new_[4378]_ ;
  assign \new_[4083]_  = \new_[1966]_  ^ \new_[4379]_ ;
  assign \new_[4084]_  = \new_[2424]_  ^ \new_[4377]_ ;
  assign \new_[4085]_  = \new_[2422]_  ^ \new_[4380]_ ;
  assign \new_[4086]_  = \new_[2352]_  ^ \new_[4381]_ ;
  assign \new_[4087]_  = \new_[2423]_  ^ \new_[4382]_ ;
  assign \new_[4088]_  = \new_[2198]_  ^ \new_[4384]_ ;
  assign \new_[4089]_  = \new_[2162]_  ^ \new_[4385]_ ;
  assign \new_[4090]_  = \new_[2202]_  ^ \new_[4387]_ ;
  assign \new_[4091]_  = \new_[2199]_  ^ \new_[4388]_ ;
  assign \new_[4092]_  = \new_[2461]_  ^ \new_[4386]_ ;
  assign \new_[4093]_  = \new_[2200]_  ^ \new_[4389]_ ;
  assign \new_[4094]_  = \new_[2353]_  ^ \new_[4383]_ ;
  assign \new_[4095]_  = \new_[2201]_  ^ \new_[4390]_ ;
  assign \new_[4096]_  = \new_[2203]_  ^ \new_[4392]_ ;
  assign \new_[4097]_  = \new_[2139]_  ^ \new_[4393]_ ;
  assign \new_[4098]_  = \new_[2425]_  ^ \new_[4391]_ ;
  assign \new_[4099]_  = \new_[2067]_  ^ \new_[4394]_ ;
  assign \new_[4100]_  = \new_[2070]_  ^ \new_[4395]_ ;
  assign \new_[4101]_  = \new_[7973]_  ^ \new_[4397]_ ;
  assign \new_[4102]_  = \new_[2354]_  ^ \new_[4396]_ ;
  assign \new_[4103]_  = \new_[7968]_  ^ \new_[4398]_ ;
  assign \new_[4104]_  = \new_[2348]_  ^ \new_[4400]_ ;
  assign \new_[4105]_  = \new_[7991]_  ^ \new_[4399]_ ;
  assign \new_[4106]_  = \new_[2344]_  ^ \new_[4401]_ ;
  assign \new_[4107]_  = \new_[2349]_  ^ \new_[4403]_ ;
  assign \new_[4108]_  = \new_[8064]_  ^ \new_[4402]_ ;
  assign \new_[4109]_  = \new_[2537]_  ^ \new_[4404]_ ;
  assign \new_[4110]_  = \new_[8109]_  ^ \new_[4405]_ ;
  assign \new_[4111]_  = \new_[8156]_  ^ \new_[4406]_ ;
  assign \new_[4112]_  = \new_[8150]_  ^ \new_[4407]_ ;
  assign \new_[4113]_  = \new_[8008]_  ^ \new_[4408]_ ;
  assign \new_[4114]_  = \new_[8141]_  ^ \new_[4409]_ ;
  assign \new_[4115]_  = \new_[8011]_  ^ \new_[4410]_ ;
  assign \new_[4116]_  = \new_[8057]_  ^ \new_[4411]_ ;
  assign \new_[4117]_  = \new_[8138]_  ^ \new_[4412]_ ;
  assign \new_[4118]_  = \new_[7993]_  ^ \new_[4414]_ ;
  assign \new_[4119]_  = \new_[8122]_  ^ \new_[4415]_ ;
  assign \new_[4120]_  = \new_[8009]_  ^ \new_[4416]_ ;
  assign \new_[4121]_  = \new_[1978]_  ^ \new_[4417]_ ;
  assign \new_[4122]_  = \new_[1977]_  ^ \new_[4419]_ ;
  assign \new_[4123]_  = ~\new_[4430]_  | ~\new_[4327]_ ;
  assign \new_[4124]_  = ~\new_[4518]_  & ~\new_[8964]_ ;
  assign \new_[4125]_  = ~\new_[4517]_  & ~\new_[8964]_ ;
  assign \new_[4126]_  = ~\new_[4519]_  & ~\new_[8964]_ ;
  assign \new_[4127]_  = ~\new_[4525]_  & ~\new_[8964]_ ;
  assign \new_[4128]_  = ~\new_[4570]_  & ~\new_[8964]_ ;
  assign \new_[4129]_  = ~\new_[4516]_  & ~\new_[8964]_ ;
  assign \new_[4130]_  = ~\new_[6162]_  | ~\new_[4247]_ ;
  assign \new_[4131]_  = ~\new_[8710]_  | ~\new_[4240]_ ;
  assign \new_[4132]_  = \new_[4331]_  & \new_[4413]_ ;
  assign \new_[4133]_  = \new_[4331]_  | \new_[4413]_ ;
  assign \new_[4134]_  = ~\new_[4715]_  | ~\new_[4360]_ ;
  assign \new_[4135]_  = ~\new_[4225]_ ;
  assign \new_[4136]_  = ~\new_[4228]_ ;
  assign \new_[4137]_  = (~\key_i[48]  | ~\new_[4798]_ ) & (~\new_[8008]_  | ~\new_[8726]_ );
  assign \new_[4138]_  = (~\key_i[50]  | ~\new_[4798]_ ) & (~\new_[8011]_  | ~\new_[8726]_ );
  assign \new_[4139]_  = (~\key_i[51]  | ~\new_[4798]_ ) & (~\new_[8057]_  | ~\new_[8726]_ );
  assign \new_[4140]_  = (~\key_i[33]  | ~\new_[4798]_ ) & (~\new_[7968]_  | ~\new_[8726]_ );
  assign \new_[4141]_  = (~\key_i[52]  | ~\new_[4798]_ ) & (~\new_[8138]_  | ~\new_[8726]_ );
  assign \new_[4142]_  = (~\key_i[55]  | ~\new_[4798]_ ) & (~\new_[8009]_  | ~\new_[8726]_ );
  assign \new_[4143]_  = ~\new_[4332]_ ;
  assign \new_[4144]_  = ~\new_[4246]_ ;
  assign n3525 = ~\new_[7460]_  | (~\new_[4448]_  & ~\new_[7560]_ );
  assign n3515 = ~\new_[7458]_  | (~\new_[4449]_  & ~\new_[7560]_ );
  assign n3520 = ~\new_[7437]_  | (~\new_[4450]_  & ~\new_[7560]_ );
  assign n3510 = ~\new_[7420]_  | (~\new_[4451]_  & ~\new_[7560]_ );
  assign \new_[4149]_  = (~\key_i[43]  | ~\new_[4798]_ ) & (~\new_[1079]_  | ~\new_[8726]_ );
  assign \new_[4150]_  = ~\new_[4240]_ ;
  assign \new_[4151]_  = ~\new_[4241]_ ;
  assign \new_[4152]_  = ~\new_[4244]_ ;
  assign \new_[4153]_  = \new_[5737]_  ? \new_[4798]_  : \key_i[75] ;
  assign \new_[4154]_  = \new_[5735]_  ? \new_[4798]_  : \key_i[76] ;
  assign \new_[4155]_  = \new_[5738]_  ? \new_[4798]_  : \key_i[77] ;
  assign \new_[4156]_  = ~\new_[4247]_ ;
  assign \new_[4157]_  = ~\new_[4232]_ ;
  assign \new_[4158]_  = (~\key_i[44]  | ~\new_[4798]_ ) & (~\new_[1080]_  | ~\new_[8726]_ );
  assign \new_[4159]_  = ~\new_[4356]_  | (~\new_[8710]_  & ~\new_[2998]_ );
  assign \new_[4160]_  = ~\new_[4357]_  | (~\new_[8710]_  & ~\new_[2999]_ );
  assign \new_[4161]_  = ~\new_[4358]_  | (~\new_[8710]_  & ~\new_[3001]_ );
  assign \new_[4162]_  = ~\new_[4359]_  | (~\new_[8710]_  & ~\new_[3000]_ );
  assign \new_[4163]_  = ~\new_[7146]_  & ~\new_[8965]_ ;
  assign \new_[4164]_  = ~\new_[4271]_ ;
  assign \new_[4165]_  = (~\key_i[42]  | ~\new_[4798]_ ) & (~\new_[1118]_  | ~\new_[8726]_ );
  assign \new_[4166]_  = \new_[4996]_  ? \new_[7632]_  : \new_[4452]_ ;
  assign \new_[4167]_  = ~\new_[4272]_ ;
  assign \new_[4168]_  = \new_[4998]_  ? \new_[7632]_  : \new_[4455]_ ;
  assign \new_[4169]_  = \new_[4731]_  ? \new_[7632]_  : \new_[4454]_ ;
  assign \new_[4170]_  = ~\new_[4273]_ ;
  assign \new_[4171]_  = \new_[4733]_  ? \new_[7632]_  : \new_[4458]_ ;
  assign \new_[4172]_  = \new_[4732]_  ? \new_[7632]_  : \new_[4456]_ ;
  assign \new_[4173]_  = \new_[5000]_  ? \new_[7632]_  : \new_[4459]_ ;
  assign \new_[4174]_  = \new_[5002]_  ? \new_[7632]_  : \new_[4461]_ ;
  assign \new_[4175]_  = ~\new_[4274]_ ;
  assign \new_[4176]_  = ~\new_[4275]_ ;
  assign \new_[4177]_  = \new_[4734]_  ? \new_[7632]_  : \new_[4463]_ ;
  assign \new_[4178]_  = \new_[4453]_  ^ \new_[4719]_ ;
  assign \new_[4179]_  = \new_[4457]_  ^ \new_[4720]_ ;
  assign \new_[4180]_  = \new_[4460]_  ^ \new_[4719]_ ;
  assign \new_[4181]_  = \new_[4462]_  ^ \new_[4720]_ ;
  assign \new_[4182]_  = ~\new_[4281]_ ;
  assign \new_[4183]_  = ~\new_[4282]_ ;
  assign \new_[4184]_  = ~\new_[4283]_ ;
  assign \new_[4185]_  = ~\new_[4284]_ ;
  assign \new_[4186]_  = (~\key_i[32]  | ~\new_[4798]_ ) & (~\new_[7973]_  | ~\new_[8726]_ );
  assign \new_[4187]_  = \new_[5561]_  ? \new_[7888]_  : \new_[4468]_ ;
  assign \new_[4188]_  = \new_[5569]_  ? \new_[7878]_  : \new_[4470]_ ;
  assign \new_[4189]_  = \new_[5562]_  ? \new_[7882]_  : \new_[4471]_ ;
  assign \new_[4190]_  = \new_[5563]_  ? \new_[7882]_  : \new_[4472]_ ;
  assign \new_[4191]_  = \new_[5565]_  ? \new_[7885]_  : \new_[4473]_ ;
  assign \new_[4192]_  = \new_[5566]_  ? \new_[7885]_  : \new_[4474]_ ;
  assign \new_[4193]_  = \new_[5567]_  ? \new_[7884]_  : \new_[4475]_ ;
  assign \new_[4194]_  = \new_[5568]_  ? \new_[7878]_  : \new_[4476]_ ;
  assign \new_[4195]_  = \new_[5571]_  ? \new_[7885]_  : \new_[4477]_ ;
  assign \new_[4196]_  = \new_[5564]_  ? \new_[7882]_  : \new_[4479]_ ;
  assign \new_[4197]_  = \new_[5586]_  ? \new_[7884]_  : \new_[4480]_ ;
  assign \new_[4198]_  = \new_[5572]_  ? \new_[7884]_  : \new_[4469]_ ;
  assign \new_[4199]_  = \new_[5573]_  ? \new_[7884]_  : \new_[4478]_ ;
  assign \new_[4200]_  = \new_[5574]_  ? \new_[7888]_  : \new_[4481]_ ;
  assign \new_[4201]_  = \new_[5570]_  ? \new_[7888]_  : \new_[4489]_ ;
  assign \new_[4202]_  = \new_[5575]_  ? \new_[7888]_  : \new_[4482]_ ;
  assign \new_[4203]_  = \new_[5577]_  ? \new_[7885]_  : \new_[4483]_ ;
  assign \new_[4204]_  = \new_[5578]_  ? \new_[7885]_  : \new_[4484]_ ;
  assign \new_[4205]_  = \new_[5581]_  ? \new_[7885]_  : \new_[4485]_ ;
  assign \new_[4206]_  = \new_[5583]_  ? \new_[7884]_  : \new_[4487]_ ;
  assign \new_[4207]_  = \new_[5584]_  ? \new_[7882]_  : \new_[4493]_ ;
  assign \new_[4208]_  = \new_[5579]_  ? \new_[7885]_  : \new_[4491]_ ;
  assign \new_[4209]_  = \new_[5576]_  ? \new_[7885]_  : \new_[4486]_ ;
  assign \new_[4210]_  = \new_[5580]_  ? \new_[7882]_  : \new_[4490]_ ;
  assign \new_[4211]_  = \new_[5582]_  ? \new_[7884]_  : \new_[4492]_ ;
  assign \new_[4212]_  = \new_[5585]_  ? \new_[7888]_  : \new_[4488]_ ;
  assign \new_[4213]_  = \new_[5588]_  ? \new_[7882]_  : \new_[4494]_ ;
  assign \new_[4214]_  = \new_[5587]_  ? \new_[7878]_  : \new_[4495]_ ;
  assign \new_[4215]_  = \new_[5589]_  ? \new_[7882]_  : \new_[4496]_ ;
  assign \new_[4216]_  = \new_[5590]_  ? \new_[7882]_  : \new_[4497]_ ;
  assign \new_[4217]_  = \new_[5591]_  ? \new_[7888]_  : \new_[4498]_ ;
  assign \new_[4218]_  = \new_[5592]_  ? \new_[7884]_  : \new_[4499]_ ;
  assign \new_[4219]_  = \new_[5593]_  ? \new_[7884]_  : \new_[4500]_ ;
  assign \new_[4220]_  = \new_[5594]_  ? \new_[7884]_  : \new_[4501]_ ;
  assign \new_[4221]_  = \new_[5595]_  ? \new_[7884]_  : \new_[4502]_ ;
  assign \new_[4222]_  = \new_[5596]_  ? \new_[7884]_  : \new_[4503]_ ;
  assign \new_[4223]_  = ~\new_[4467]_  & (~\new_[4436]_  | ~\new_[8329]_ );
  assign \new_[4224]_  = ~\new_[4522]_  & ~\new_[8964]_ ;
  assign \new_[4225]_  = ~\new_[4523]_  | ~\new_[4446]_ ;
  assign \new_[4226]_  = ~\new_[4716]_  | ~\new_[4447]_ ;
  assign \new_[4227]_  = ~\new_[4330]_ ;
  assign \new_[4228]_  = (~\key_i[71]  | ~\new_[4798]_ ) & (~\new_[2138]_  | ~\new_[8726]_ );
  assign \new_[4229]_  = (~\key_i[72]  | ~\new_[4798]_ ) & (~\new_[1140]_  | ~\new_[8726]_ );
  assign \new_[4230]_  = \\ks1_state_reg[0] ;
  assign n3530 = \new_[4441]_  | \new_[4624]_ ;
  assign \new_[4232]_  = (~\key_i[69]  | ~\new_[4798]_ ) & (~\new_[2095]_  | ~\new_[8726]_ );
  assign n3535 = \new_[4442]_  | \new_[4626]_ ;
  assign \new_[4234]_  = (~\new_[8726]_  | ~\new_[8119]_ ) & (~\key_i[73]  | ~\new_[4798]_ );
  assign \new_[4235]_  = \key_i[35]  ? \new_[5114]_  : \new_[5599]_ ;
  assign \new_[4236]_  = \key_i[37]  ? \new_[5114]_  : \new_[5600]_ ;
  assign \new_[4237]_  = \key_i[114]  ? \new_[5114]_  : \new_[5865]_ ;
  assign \new_[4238]_  = \key_i[116]  ? \new_[5114]_  : \new_[5812]_ ;
  assign \new_[4239]_  = (~\new_[5768]_  | ~\new_[5114]_ ) & (~\key_i[64]  | ~\new_[4798]_ );
  assign \new_[4240]_  = \new_[5289]_  ? \new_[7632]_  : \new_[4530]_ ;
  assign \new_[4241]_  = \new_[5290]_  ? \new_[7632]_  : \new_[4531]_ ;
  assign \new_[4242]_  = \key_i[113]  ? \new_[5114]_  : \new_[5813]_ ;
  assign \new_[4243]_  = \new_[5736]_  ? \new_[4798]_  : \key_i[74] ;
  assign \new_[4244]_  = \new_[5291]_  ? \new_[7583]_  : \new_[4532]_ ;
  assign \new_[4245]_  = \key_i[119]  ? \new_[5114]_  : \new_[5868]_ ;
  assign \new_[4246]_  = (~\key_i[70]  | ~\new_[4798]_ ) & (~\new_[2137]_  | ~\new_[8726]_ );
  assign \new_[4247]_  = \new_[5292]_  ? \new_[7632]_  : \new_[4533]_ ;
  assign \new_[4248]_  = \new_[5734]_  ? \new_[4798]_  : \key_i[78] ;
  assign \new_[4249]_  = \new_[5739]_  ? \new_[4798]_  : \key_i[79] ;
  assign \new_[4250]_  = (~\new_[5740]_  | ~\new_[5114]_ ) & (~\key_i[80]  | ~\new_[3675]_ );
  assign \new_[4251]_  = (~\new_[5731]_  | ~\new_[5114]_ ) & (~\key_i[81]  | ~\new_[3675]_ );
  assign \new_[4252]_  = (~\new_[5741]_  | ~\new_[5114]_ ) & (~\key_i[82]  | ~\new_[4798]_ );
  assign \new_[4253]_  = (~\new_[5742]_  | ~\new_[5114]_ ) & (~\key_i[83]  | ~\new_[4798]_ );
  assign \new_[4254]_  = (~\new_[5769]_  | ~\new_[5114]_ ) & (~\key_i[65]  | ~\new_[4798]_ );
  assign \new_[4255]_  = (~\new_[5743]_  | ~\new_[5114]_ ) & (~\key_i[84]  | ~\new_[4798]_ );
  assign \new_[4256]_  = (~\new_[5744]_  | ~\new_[5114]_ ) & (~\key_i[85]  | ~\new_[4798]_ );
  assign \new_[4257]_  = (~\new_[5745]_  | ~\new_[5114]_ ) & (~\key_i[86]  | ~\new_[4798]_ );
  assign \new_[4258]_  = (~\new_[5770]_  | ~\new_[5114]_ ) & (~\key_i[87]  | ~\new_[4798]_ );
  assign \new_[4259]_  = (~\new_[5746]_  | ~\new_[5114]_ ) & (~\key_i[89]  | ~\new_[3675]_ );
  assign \new_[4260]_  = (~\new_[5748]_  | ~\new_[5114]_ ) & (~\key_i[91]  | ~\new_[3675]_ );
  assign \new_[4261]_  = (~\new_[5771]_  | ~\new_[5114]_ ) & (~\key_i[92]  | ~\new_[3675]_ );
  assign \new_[4262]_  = (~\new_[5767]_  | ~\new_[5114]_ ) & (~\key_i[66]  | ~\new_[3675]_ );
  assign \new_[4263]_  = ~\new_[4451]_  & ~\new_[7829]_ ;
  assign \new_[4264]_  = ~\new_[4448]_  & ~\new_[7829]_ ;
  assign \new_[4265]_  = ~\new_[4449]_  & ~\new_[7829]_ ;
  assign \new_[4266]_  = ~\new_[4450]_  & ~\new_[7829]_ ;
  assign \new_[4267]_  = ~\new_[4451]_  & ~\new_[8562]_ ;
  assign \new_[4268]_  = ~\new_[4448]_  & ~\new_[8562]_ ;
  assign \new_[4269]_  = ~\new_[4449]_  & ~\new_[8562]_ ;
  assign \new_[4270]_  = ~\new_[4450]_  & ~\new_[8562]_ ;
  assign \new_[4271]_  = (~\key_i[68]  | ~\new_[4798]_ ) & (~\new_[2136]_  | ~\new_[8726]_ );
  assign \new_[4272]_  = \new_[5369]_  ? \new_[7632]_  : \new_[4535]_ ;
  assign \new_[4273]_  = \new_[5371]_  ? \new_[7632]_  : \new_[4537]_ ;
  assign \new_[4274]_  = \new_[5373]_  ? \new_[7583]_  : \new_[4539]_ ;
  assign \new_[4275]_  = \new_[5375]_  ? \new_[7632]_  : \new_[4541]_ ;
  assign \new_[4276]_  = \new_[4992]_  ^ \new_[4534]_ ;
  assign \new_[4277]_  = \new_[4993]_  ^ \new_[4536]_ ;
  assign \new_[4278]_  = \new_[4992]_  ^ \new_[4538]_ ;
  assign \new_[4279]_  = \new_[4993]_  ^ \new_[4540]_ ;
  assign n3540 = \new_[4443]_  | \new_[4625]_ ;
  assign \new_[4281]_  = \new_[4820]_  ? \new_[7632]_  : \new_[4543]_ ;
  assign \new_[4282]_  = \new_[4828]_  ? \new_[7632]_  : \new_[4544]_ ;
  assign \new_[4283]_  = \new_[4824]_  ? \new_[7632]_  : \new_[4545]_ ;
  assign \new_[4284]_  = \new_[4821]_  ? \new_[7632]_  : \new_[4546]_ ;
  assign \new_[4285]_  = \new_[5622]_  ? \new_[7885]_  : \new_[4547]_ ;
  assign \new_[4286]_  = \new_[5624]_  ? \new_[7882]_  : \new_[4548]_ ;
  assign \new_[4287]_  = \new_[5623]_  ? \new_[7888]_  : \new_[4549]_ ;
  assign \new_[4288]_  = \new_[5629]_  ? \new_[7885]_  : \new_[4550]_ ;
  assign \new_[4289]_  = \new_[5630]_  ? \new_[7884]_  : \new_[4551]_ ;
  assign \new_[4290]_  = \new_[5631]_  ? \new_[7884]_  : \new_[4552]_ ;
  assign \new_[4291]_  = \new_[5632]_  ? \new_[7882]_  : \new_[4553]_ ;
  assign \new_[4292]_  = \new_[5634]_  ? \new_[7884]_  : \new_[4554]_ ;
  assign \new_[4293]_  = \new_[5628]_  ? \new_[7878]_  : \new_[4555]_ ;
  assign \new_[4294]_  = \new_[5626]_  ? \new_[7884]_  : \new_[4579]_ ;
  assign \new_[4295]_  = \new_[5637]_  ? \new_[7878]_  : \new_[4556]_ ;
  assign \new_[4296]_  = \new_[5633]_  ? \new_[7878]_  : \new_[4558]_ ;
  assign \new_[4297]_  = \new_[5625]_  ? \new_[7884]_  : \new_[4559]_ ;
  assign \new_[4298]_  = \new_[5651]_  ? \new_[7885]_  : \new_[4560]_ ;
  assign \new_[4299]_  = \new_[5642]_  ? \new_[7882]_  : \new_[4561]_ ;
  assign \new_[4300]_  = \new_[5635]_  ? \new_[7888]_  : \new_[4562]_ ;
  assign \new_[4301]_  = \new_[5627]_  ? \new_[7884]_  : \new_[4573]_ ;
  assign \new_[4302]_  = \new_[5640]_  ? \new_[7882]_  : \new_[4563]_ ;
  assign \new_[4303]_  = \new_[5653]_  ? \new_[7882]_  : \new_[4564]_ ;
  assign \new_[4304]_  = \new_[5636]_  ? \new_[7882]_  : \new_[4565]_ ;
  assign \new_[4305]_  = \new_[8235]_  ? \new_[7888]_  : \new_[4566]_ ;
  assign \new_[4306]_  = \new_[5638]_  ? \new_[7885]_  : \new_[4567]_ ;
  assign \new_[4307]_  = \new_[5639]_  ? \new_[7878]_  : \new_[4568]_ ;
  assign \new_[4308]_  = \new_[5641]_  ? \new_[7882]_  : \new_[4557]_ ;
  assign \new_[4309]_  = \new_[5643]_  ? \new_[7888]_  : \new_[4569]_ ;
  assign \new_[4310]_  = \new_[5644]_  ? \new_[7884]_  : \new_[4571]_ ;
  assign \new_[4311]_  = \new_[5645]_  ? \new_[7884]_  : \new_[4572]_ ;
  assign \new_[4312]_  = \new_[5646]_  ? \new_[7884]_  : \new_[4575]_ ;
  assign \new_[4313]_  = \new_[5647]_  ? \new_[7878]_  : \new_[4574]_ ;
  assign \new_[4314]_  = \new_[5648]_  ? \new_[7878]_  : \new_[4577]_ ;
  assign \new_[4315]_  = \new_[5649]_  ? \new_[7884]_  : \new_[4576]_ ;
  assign \new_[4316]_  = \new_[5650]_  ? \new_[7885]_  : \new_[4578]_ ;
  assign \new_[4317]_  = \new_[5652]_  ? \new_[7884]_  : \new_[4580]_ ;
  assign \new_[4318]_  = \new_[5654]_  ? \new_[7884]_  : \new_[4581]_ ;
  assign \new_[4319]_  = \new_[5655]_  ? \new_[7882]_  : \new_[4582]_ ;
  assign \new_[4320]_  = ~\new_[7025]_  | ~\new_[7604]_  | ~\new_[4329]_  | ~\new_[6636]_ ;
  assign \new_[4321]_  = \new_[5614]_  | \new_[8489]_ ;
  assign \new_[4322]_  = \new_[5668]_  | \new_[8489]_ ;
  assign \new_[4323]_  = \new_[5667]_  | \new_[8489]_ ;
  assign \new_[4324]_  = \new_[5756]_  | \new_[8489]_ ;
  assign \new_[4325]_  = \new_[5615]_  | \new_[8489]_ ;
  assign \new_[4326]_  = ~\new_[8176]_  | ~\new_[8378]_ ;
  assign \new_[4327]_  = ~\new_[4433]_  | ~\new_[8422]_ ;
  assign \new_[4328]_  = ~\new_[4440]_  | ~\new_[8329]_ ;
  assign \new_[4329]_  = ~\new_[8489]_ ;
  assign \new_[4330]_  = \new_[4520]_  | \new_[4624]_ ;
  assign \new_[4331]_  = \new_[4521]_  | \new_[4626]_ ;
  assign \new_[4332]_  = ~\new_[4797]_  | ~\new_[8965]_ ;
  assign \new_[4333]_  = (~\new_[5729]_  | ~\new_[5114]_ ) & (~\key_i[94]  | ~\new_[4798]_ );
  assign \new_[4334]_  = (~\new_[5730]_  | ~\new_[5114]_ ) & (~\key_i[95]  | ~\new_[4798]_ );
  assign \new_[4335]_  = \key_i[107]  ? \new_[5114]_  : \new_[5861]_ ;
  assign \new_[4336]_  = \key_i[115]  ? \new_[5114]_  : \new_[5809]_ ;
  assign \new_[4337]_  = \key_i[100]  ? \new_[5114]_  : \new_[5805]_ ;
  assign \new_[4338]_  = \key_i[112]  ? \new_[5114]_  : \new_[5867]_ ;
  assign \new_[4339]_  = \key_i[96]  ? \new_[5114]_  : \new_[5864]_ ;
  assign \new_[4340]_  = \key_i[108]  ? \new_[5114]_  : \new_[5863]_ ;
  assign \new_[4341]_  = \key_i[101]  ? \new_[5114]_  : \new_[5810]_ ;
  assign \new_[4342]_  = \key_i[102]  ? \new_[5114]_  : \new_[5807]_ ;
  assign \new_[4343]_  = \key_i[103]  ? \new_[5114]_  : \new_[5804]_ ;
  assign \new_[4344]_  = \key_i[104]  ? \new_[5114]_  : \new_[5808]_ ;
  assign \new_[4345]_  = \key_i[105]  ? \new_[5114]_  : \new_[5862]_ ;
  assign \new_[4346]_  = (~\new_[5811]_  | ~\new_[5114]_ ) & (~\key_i[109]  | ~\new_[3675]_ );
  assign \new_[4347]_  = (~\new_[5806]_  | ~\new_[5114]_ ) & (~\key_i[110]  | ~\new_[3675]_ );
  assign \new_[4348]_  = \key_i[111]  ? \new_[5114]_  : \new_[5866]_ ;
  assign \new_[4349]_  = \key_i[118]  ? \new_[5114]_  : \new_[5860]_ ;
  assign \new_[4350]_  = \key_i[117]  ? \new_[5114]_  : \new_[5814]_ ;
  assign \new_[4351]_  = \key_i[97]  ? \new_[5114]_  : \new_[5869]_ ;
  assign \new_[4352]_  = (~\new_[5732]_  | ~\new_[5114]_ ) & (~\key_i[88]  | ~\new_[4798]_ );
  assign \new_[4353]_  = \key_i[90]  ? \new_[5114]_  : \new_[5747]_ ;
  assign \new_[4354]_  = \key_i[93]  ? \new_[5114]_  : \new_[5733]_ ;
  assign \new_[4355]_  = \key_i[98]  ? \new_[5114]_  : \new_[5870]_ ;
  assign \new_[4356]_  = ~\new_[6161]_  | ~\new_[4529]_ ;
  assign \new_[4357]_  = ~\new_[6162]_  | ~\new_[4526]_ ;
  assign \new_[4358]_  = ~\new_[6162]_  | ~\new_[4527]_ ;
  assign \new_[4359]_  = ~\new_[6162]_  | ~\new_[4528]_ ;
  assign \new_[4360]_  = ~\new_[4622]_  & (~\key_i[67]  | ~\new_[4798]_ );
  assign \new_[4361]_  = ~\new_[8828]_ ;
  assign \new_[4362]_  = \\ks1_state_reg[2] ;
  assign \new_[4363]_  = \new_[5673]_  ? \new_[7878]_  : \new_[4629]_ ;
  assign \new_[4364]_  = \new_[5674]_  ? \new_[7888]_  : \new_[4630]_ ;
  assign \new_[4365]_  = \new_[5710]_  ? \new_[7882]_  : \new_[4631]_ ;
  assign \new_[4366]_  = \new_[5694]_  ? \new_[7884]_  : \new_[4635]_ ;
  assign \new_[4367]_  = \new_[5675]_  ? \new_[7882]_  : \new_[4632]_ ;
  assign \new_[4368]_  = \new_[5676]_  ? \new_[7885]_  : \new_[4633]_ ;
  assign \new_[4369]_  = \new_[5678]_  ? \new_[7884]_  : \new_[4634]_ ;
  assign \new_[4370]_  = \new_[5679]_  ? \new_[7885]_  : \new_[4636]_ ;
  assign \new_[4371]_  = \new_[5680]_  ? \new_[7884]_  : \new_[4637]_ ;
  assign \new_[4372]_  = \new_[5681]_  ? \new_[7878]_  : \new_[4638]_ ;
  assign \new_[4373]_  = \new_[5682]_  ? \new_[7884]_  : \new_[4639]_ ;
  assign \new_[4374]_  = \new_[5683]_  ? \new_[7884]_  : \new_[4640]_ ;
  assign \new_[4375]_  = \new_[5684]_  ? \new_[7888]_  : \new_[4641]_ ;
  assign \new_[4376]_  = \new_[5685]_  ? \new_[7884]_  : \new_[4642]_ ;
  assign \new_[4377]_  = \new_[5686]_  ? \new_[7882]_  : \new_[4643]_ ;
  assign \new_[4378]_  = \new_[5687]_  ? \new_[7884]_  : \new_[4644]_ ;
  assign \new_[4379]_  = \new_[5688]_  ? \new_[7884]_  : \new_[4645]_ ;
  assign \new_[4380]_  = \new_[5689]_  ? \new_[7878]_  : \new_[4647]_ ;
  assign \new_[4381]_  = \new_[5726]_  ? \new_[7888]_  : \new_[4646]_ ;
  assign \new_[4382]_  = \new_[5696]_  ? \new_[7878]_  : \new_[4648]_ ;
  assign \new_[4383]_  = \new_[5690]_  ? \new_[7884]_  : \new_[4649]_ ;
  assign \new_[4384]_  = \new_[5691]_  ? \new_[7884]_  : \new_[4650]_ ;
  assign \new_[4385]_  = \new_[5714]_  ? \new_[7882]_  : \new_[4651]_ ;
  assign \new_[4386]_  = \new_[5692]_  ? \new_[7882]_  : \new_[4652]_ ;
  assign \new_[4387]_  = \new_[5693]_  ? \new_[7885]_  : \new_[4653]_ ;
  assign \new_[4388]_  = \new_[5695]_  ? \new_[7884]_  : \new_[4654]_ ;
  assign \new_[4389]_  = \new_[5728]_  ? \new_[7882]_  : \new_[4675]_ ;
  assign \new_[4390]_  = \new_[5703]_  ? \new_[7878]_  : \new_[4656]_ ;
  assign \new_[4391]_  = \new_[5697]_  ? \new_[7884]_  : \new_[4657]_ ;
  assign \new_[4392]_  = \new_[5698]_  ? \new_[7888]_  : \new_[4658]_ ;
  assign \new_[4393]_  = \new_[5699]_  ? \new_[7882]_  : \new_[4659]_ ;
  assign \new_[4394]_  = \new_[5700]_  ? \new_[7882]_  : \new_[4660]_ ;
  assign \new_[4395]_  = \new_[5701]_  ? \new_[7884]_  : \new_[4655]_ ;
  assign \new_[4396]_  = \new_[5702]_  ? \new_[7882]_  : \new_[4661]_ ;
  assign \new_[4397]_  = \new_[5704]_  ? \new_[7884]_  : \new_[4662]_ ;
  assign \new_[4398]_  = \new_[5705]_  ? \new_[7878]_  : \new_[4663]_ ;
  assign \new_[4399]_  = \new_[5706]_  ? \new_[7884]_  : \new_[4664]_ ;
  assign \new_[4400]_  = \new_[5672]_  ? \new_[7888]_  : \new_[4665]_ ;
  assign \new_[4401]_  = \new_[5707]_  ? \new_[7884]_  : \new_[4666]_ ;
  assign \new_[4402]_  = \new_[5725]_  ? \new_[7884]_  : \new_[4667]_ ;
  assign \new_[4403]_  = \new_[5708]_  ? \new_[7884]_  : \new_[4668]_ ;
  assign \new_[4404]_  = \new_[5709]_  ? \new_[7878]_  : \new_[4669]_ ;
  assign \new_[4405]_  = \new_[5677]_  ? \new_[7884]_  : \new_[4670]_ ;
  assign \new_[4406]_  = \new_[5711]_  ? \new_[7884]_  : \new_[4671]_ ;
  assign \new_[4407]_  = \new_[5712]_  ? \new_[7884]_  : \new_[4672]_ ;
  assign \new_[4408]_  = \new_[5713]_  ? \new_[7882]_  : \new_[4673]_ ;
  assign \new_[4409]_  = \new_[5715]_  ? \new_[7882]_  : \new_[4674]_ ;
  assign \new_[4410]_  = \new_[5716]_  ? \new_[7882]_  : \new_[4676]_ ;
  assign \new_[4411]_  = \new_[5717]_  ? \new_[7882]_  : \new_[4677]_ ;
  assign \new_[4412]_  = \new_[5718]_  ? \new_[7882]_  : \new_[4678]_ ;
  assign \new_[4413]_  = ~\new_[4625]_  & (~\new_[5961]_  | ~\new_[4627]_ );
  assign \new_[4414]_  = \new_[5719]_  ? \new_[7884]_  : \new_[4679]_ ;
  assign \new_[4415]_  = \new_[5720]_  ? \new_[7884]_  : \new_[4680]_ ;
  assign \new_[4416]_  = \new_[5721]_  ? \new_[7884]_  : \new_[4681]_ ;
  assign \new_[4417]_  = \new_[5722]_  ? \new_[7888]_  : \new_[4682]_ ;
  assign \new_[4418]_  = \new_[5723]_  ? \new_[7882]_  : \new_[4683]_ ;
  assign \new_[4419]_  = \new_[5724]_  ? \new_[7884]_  : \new_[4684]_ ;
  assign \new_[4420]_  = \new_[5727]_  ? \new_[7882]_  : \new_[4628]_ ;
  assign \new_[4421]_  = \new_[5757]_  | \new_[8489]_ ;
  assign \new_[4422]_  = ~\new_[8847]_  | ~\new_[8378]_ ;
  assign \new_[4423]_  = ~\new_[4510]_  | ~\new_[8378]_ ;
  assign \new_[4424]_  = ~\new_[4511]_  | ~\new_[8329]_ ;
  assign \new_[4425]_  = ~\new_[4506]_  | ~\new_[8422]_ ;
  assign \new_[4426]_  = ~\new_[4509]_  | ~\new_[8422]_ ;
  assign \new_[4427]_  = ~\new_[8840]_  | ~\new_[8378]_ ;
  assign \new_[4428]_  = ~\new_[4515]_  | ~\new_[8424]_ ;
  assign \new_[4429]_  = ~\new_[4507]_  | ~\new_[8424]_ ;
  assign \new_[4430]_  = ~\new_[4524]_  | ~\new_[8424]_ ;
  assign \new_[4431]_  = ~\new_[4508]_ ;
  assign \new_[4432]_  = ~\new_[8423]_ ;
  assign \new_[4433]_  = ~\new_[8878]_ ;
  assign \new_[4434]_  = ~\new_[8250]_ ;
  assign \new_[4435]_  = ~\new_[4509]_ ;
  assign \new_[4436]_  = ~\new_[8785]_ ;
  assign \new_[4437]_  = ~\new_[8312]_ ;
  assign \new_[4438]_  = ~\new_[4512]_ ;
  assign \new_[4439]_  = ~\new_[8297]_ ;
  assign \new_[4440]_  = ~\new_[4513]_ ;
  assign \new_[4441]_  = \new_[5765]_  & \new_[4627]_ ;
  assign \new_[4442]_  = \new_[5849]_  & \new_[4627]_ ;
  assign \new_[4443]_  = \new_[5857]_  & \new_[4627]_ ;
  assign \new_[4444]_  = \key_i[99]  ? \new_[5114]_  : \new_[5859]_ ;
  assign \new_[4445]_  = \key_i[106]  ? \new_[5114]_  : \new_[5832]_ ;
  assign \new_[4446]_  = ~\new_[8964]_  | ~\new_[7923]_ ;
  assign \new_[4447]_  = ~\new_[4623]_  & (~\key_i[124]  | ~\new_[3675]_ );
  assign \new_[4448]_  = ~\new_[4526]_ ;
  assign \new_[4449]_  = ~\new_[4527]_ ;
  assign \new_[4450]_  = ~\new_[4528]_ ;
  assign \new_[4451]_  = ~\new_[4529]_ ;
  assign \new_[4452]_  = \new_[5128]_  ^ \new_[4722]_ ;
  assign \new_[4453]_  = \new_[8636]_  ^ \new_[4723]_ ;
  assign \new_[4454]_  = \new_[8523]_  ^ \new_[4731]_ ;
  assign \new_[4455]_  = \new_[5131]_  ^ \new_[4724]_ ;
  assign \new_[4456]_  = \new_[8523]_  ^ \new_[4732]_ ;
  assign \new_[4457]_  = \new_[8601]_  ^ \new_[4725]_ ;
  assign \new_[4458]_  = \new_[8494]_  ^ \new_[4733]_ ;
  assign \new_[4459]_  = \new_[5128]_  ^ \new_[4726]_ ;
  assign \new_[4460]_  = \new_[5251]_  ^ \new_[4730]_ ;
  assign \new_[4461]_  = \new_[5131]_  ^ \new_[4727]_ ;
  assign \new_[4462]_  = \new_[8751]_  ^ \new_[4728]_ ;
  assign \new_[4463]_  = \new_[8494]_  ^ \new_[4734]_ ;
  assign \new_[4464]_  = ~\new_[4542]_ ;
  assign \new_[4465]_  = \new_[8490]_  & \new_[7259]_ ;
  assign \new_[4466]_  = \new_[4618]_  | \new_[7826]_ ;
  assign \new_[4467]_  = ~\new_[4621]_  & ~\new_[8418]_ ;
  assign \new_[4468]_  = ~\new_[4685]_  & (~\new_[7097]_  | ~\new_[1249]_ );
  assign \new_[4469]_  = ~\new_[4592]_  & (~\new_[6785]_  | ~\new_[1311]_ );
  assign \new_[4470]_  = ~\new_[4686]_  & (~\new_[6770]_  | ~\new_[1113]_ );
  assign \new_[4471]_  = ~\new_[4583]_  & (~\new_[6770]_  | ~\new_[8053]_ );
  assign \new_[4472]_  = ~\new_[4584]_  & (~\new_[6770]_  | ~\new_[1200]_ );
  assign \new_[4473]_  = ~\new_[4585]_  & (~\new_[6770]_  | ~\new_[1100]_ );
  assign \new_[4474]_  = ~\new_[4586]_  & (~\new_[6770]_  | ~\new_[1384]_ );
  assign \new_[4475]_  = ~\new_[4587]_  & (~\new_[6770]_  | ~\new_[1101]_ );
  assign \new_[4476]_  = ~\new_[4588]_  & (~\new_[6770]_  | ~\new_[1201]_ );
  assign \new_[4477]_  = ~\new_[4589]_  & (~\new_[6785]_  | ~\new_[1136]_ );
  assign \new_[4478]_  = ~\new_[4593]_  & (~\new_[6785]_  | ~\new_[1383]_ );
  assign \new_[4479]_  = ~\new_[4590]_  & (~\new_[6770]_  | ~\new_[1145]_ );
  assign \new_[4480]_  = ~\new_[4591]_  & (~\new_[6770]_  | ~\new_[1457]_ );
  assign \new_[4481]_  = ~\new_[4594]_  & (~\new_[6770]_  | ~\new_[1217]_ );
  assign \new_[4482]_  = ~\new_[4595]_  & (~\new_[6785]_  | ~\new_[1241]_ );
  assign \new_[4483]_  = ~\new_[4596]_  & (~\new_[6785]_  | ~\new_[1458]_ );
  assign \new_[4484]_  = ~\new_[4597]_  & (~\new_[6785]_  | ~\new_[1190]_ );
  assign \new_[4485]_  = ~\new_[4598]_  & (~\new_[6785]_  | ~\new_[1314]_ );
  assign \new_[4486]_  = ~\new_[4601]_  & (~\new_[6785]_  | ~\new_[1191]_ );
  assign \new_[4487]_  = ~\new_[4599]_  & (~\new_[6785]_  | ~\new_[1197]_ );
  assign \new_[4488]_  = ~\new_[4605]_  & (~\new_[7097]_  | ~\new_[1198]_ );
  assign \new_[4489]_  = ~\new_[4603]_  & (~\new_[7097]_  | ~\new_[8026]_ );
  assign \new_[4490]_  = ~\new_[4604]_  & (~\new_[6770]_  | ~\new_[1099]_ );
  assign \new_[4491]_  = ~\new_[4602]_  & (~\new_[6785]_  | ~\new_[1134]_ );
  assign \new_[4492]_  = ~\new_[4606]_  & (~\new_[6785]_  | ~\new_[1135]_ );
  assign \new_[4493]_  = ~\new_[4600]_  & (~\new_[6785]_  | ~\new_[1196]_ );
  assign \new_[4494]_  = ~\new_[4607]_  & (~\new_[6770]_  | ~\new_[1243]_ );
  assign \new_[4495]_  = ~\new_[4608]_  & (~\new_[6785]_  | ~\new_[1096]_ );
  assign \new_[4496]_  = ~\new_[4609]_  & (~\new_[6770]_  | ~\new_[1312]_ );
  assign \new_[4497]_  = ~\new_[4611]_  & (~\new_[6770]_  | ~\new_[1095]_ );
  assign \new_[4498]_  = ~\new_[4610]_  & (~\new_[6770]_  | ~\new_[8020]_ );
  assign \new_[4499]_  = ~\new_[4612]_  & (~\new_[6770]_  | ~\new_[1385]_ );
  assign \new_[4500]_  = ~\new_[4613]_  & (~\new_[6786]_  | ~\new_[1247]_ );
  assign \new_[4501]_  = ~\new_[4614]_  & (~\new_[6786]_  | ~\new_[1112]_ );
  assign \new_[4502]_  = ~\new_[4615]_  & (~\new_[6770]_  | ~\new_[1192]_ );
  assign \new_[4503]_  = ~\new_[4616]_  & (~\new_[6763]_  | ~\new_[1248]_ );
  assign n3545 = ~\new_[7598]_  | ~\new_[8418]_ ;
  assign n3550 = ~\new_[4721]_  | (~\new_[7826]_  & ~\new_[7843]_ );
  assign \new_[4506]_  = ~\new_[4617]_ ;
  assign \new_[4507]_  = ~\new_[5071]_  | (~\new_[4782]_  & ~\new_[9001]_ );
  assign \new_[4508]_  = (~\new_[4783]_  | ~\new_[8965]_ ) & (~\new_[7475]_  | ~\new_[8967]_ );
  assign \new_[4509]_  = ~\new_[4943]_  | (~\new_[4785]_  & ~\new_[9001]_ );
  assign \new_[4510]_  = ~\new_[4619]_ ;
  assign \new_[4511]_  = ~\new_[4620]_ ;
  assign \new_[4512]_  = ~\new_[4892]_  | (~\new_[4792]_  & ~\new_[8967]_ );
  assign \new_[4513]_  = (~\new_[4793]_  | ~\new_[9000]_ ) & (~\new_[7570]_  | ~\new_[9001]_ );
  assign \new_[4514]_  = ~\new_[4621]_ ;
  assign \new_[4515]_  = ~\new_[4953]_  | (~\new_[4795]_  & ~\new_[9001]_ );
  assign \new_[4516]_  = (~\key_i[127]  | ~\new_[4798]_ ) & (~\new_[2266]_  | ~\new_[8726]_ );
  assign \new_[4517]_  = (~\key_i[121]  | ~\new_[4798]_ ) & (~\new_[2265]_  | ~\new_[8726]_ );
  assign \new_[4518]_  = (~\key_i[120]  | ~\new_[4798]_ ) & (~\new_[2264]_  | ~\new_[8726]_ );
  assign \new_[4519]_  = (~\key_i[122]  | ~\new_[4798]_ ) & (~\new_[2273]_  | ~\new_[8726]_ );
  assign \new_[4520]_  = ~\new_[4718]_  & (~\new_[6101]_  | ~\new_[6036]_ );
  assign \new_[4521]_  = ~\new_[4718]_  & (~\new_[6171]_  | ~\new_[6197]_ );
  assign \new_[4522]_  = (~\key_i[125]  | ~\new_[4798]_ ) & (~\new_[2196]_  | ~\new_[8726]_ );
  assign \new_[4523]_  = ~\new_[4717]_  | ~\new_[8965]_ ;
  assign \new_[4524]_  = ~\new_[4894]_  | (~\new_[4796]_  & ~\new_[8967]_ );
  assign \new_[4525]_  = (~\key_i[123]  | ~\new_[4798]_ ) & (~\new_[2197]_  | ~\new_[8726]_ );
  assign \new_[4526]_  = \new_[5370]_  ? \new_[7632]_  : \new_[4800]_ ;
  assign \new_[4527]_  = \new_[5372]_  ? \new_[7632]_  : \new_[4802]_ ;
  assign \new_[4528]_  = \new_[5374]_  ? \new_[7583]_  : \new_[4804]_ ;
  assign \new_[4529]_  = \new_[5376]_  ? \new_[7632]_  : \new_[4806]_ ;
  assign \new_[4530]_  = \new_[4809]_  ^ \new_[4799]_ ;
  assign \new_[4531]_  = \new_[4812]_  ^ \new_[4801]_ ;
  assign \new_[4532]_  = \new_[4815]_  ^ \new_[4803]_ ;
  assign \new_[4533]_  = \new_[4818]_  ^ \new_[4805]_ ;
  assign \new_[4534]_  = \new_[4822]_  ^ \new_[4808]_ ;
  assign \new_[4535]_  = \new_[5117]_  ^ \new_[4810]_ ;
  assign \new_[4536]_  = \new_[4823]_  ^ \new_[4811]_ ;
  assign \new_[4537]_  = \new_[5120]_  ^ \new_[4813]_ ;
  assign \new_[4538]_  = \new_[4825]_  ^ \new_[4814]_ ;
  assign \new_[4539]_  = \new_[5123]_  ^ \new_[4816]_ ;
  assign \new_[4540]_  = \new_[4826]_  ^ \new_[4817]_ ;
  assign \new_[4541]_  = \new_[5126]_  ^ \new_[4819]_ ;
  assign \new_[4542]_  = \new_[5619]_  ? \new_[4807]_  : \new_[5670]_ ;
  assign \new_[4543]_  = \new_[8526]_  ^ \new_[4820]_ ;
  assign \new_[4544]_  = \new_[8526]_  ^ \new_[4828]_ ;
  assign \new_[4545]_  = \new_[8498]_  ^ \new_[4824]_ ;
  assign \new_[4546]_  = \new_[8498]_  ^ \new_[4821]_ ;
  assign \new_[4547]_  = ~\new_[4736]_  & (~\new_[6770]_  | ~\new_[1186]_ );
  assign \new_[4548]_  = ~\new_[4737]_  & (~\new_[6770]_  | ~\new_[1187]_ );
  assign \new_[4549]_  = ~\new_[4738]_  & (~\new_[6770]_  | ~\new_[8068]_ );
  assign \new_[4550]_  = ~\new_[4739]_  & (~\new_[6770]_  | ~\new_[1144]_ );
  assign \new_[4551]_  = ~\new_[4740]_  & (~\new_[6785]_  | ~\new_[1459]_ );
  assign \new_[4552]_  = ~\new_[4741]_  & (~\new_[6770]_  | ~\new_[1224]_ );
  assign \new_[4553]_  = ~\new_[4742]_  & (~\new_[6785]_  | ~\new_[1313]_ );
  assign \new_[4554]_  = ~\new_[4687]_  & (~\new_[6770]_  | ~\new_[1199]_ );
  assign \new_[4555]_  = ~\new_[4688]_  & (~\new_[6770]_  | ~\new_[1244]_ );
  assign \new_[4556]_  = ~\new_[4690]_  & (~\new_[6770]_  | ~\new_[1245]_ );
  assign \new_[4557]_  = ~\new_[4691]_  & (~\new_[6770]_  | ~\new_[1250]_ );
  assign \new_[4558]_  = ~\new_[4692]_  & (~\new_[6785]_  | ~\new_[1320]_ );
  assign \new_[4559]_  = ~\new_[4693]_  & (~\new_[6785]_  | ~\new_[1138]_ );
  assign \new_[4560]_  = ~\new_[4694]_  & (~\new_[6785]_  | ~\new_[1142]_ );
  assign \new_[4561]_  = ~\new_[4695]_  & (~\new_[6785]_  | ~\new_[1246]_ );
  assign \new_[4562]_  = ~\new_[4696]_  & (~\new_[6770]_  | ~\new_[1386]_ );
  assign \new_[4563]_  = ~\new_[4697]_  & (~\new_[6770]_  | ~\new_[1251]_ );
  assign \new_[4564]_  = ~\new_[4698]_  & (~\new_[6770]_  | ~\new_[1252]_ );
  assign \new_[4565]_  = ~\new_[4700]_  & (~\new_[6770]_  | ~\new_[1193]_ );
  assign \new_[4566]_  = ~\new_[4699]_  & (~\new_[6770]_  | ~\new_[1139]_ );
  assign \new_[4567]_  = ~\new_[4701]_  & (~\new_[6763]_  | ~\new_[1381]_ );
  assign \new_[4568]_  = ~\new_[4702]_  & (~\new_[6770]_  | ~\new_[1137]_ );
  assign \new_[4569]_  = ~\new_[4703]_  & (~\new_[6770]_  | ~\new_[1223]_ );
  assign \new_[4570]_  = (~\key_i[126]  | ~\new_[4798]_ ) & (~\new_[2271]_  | ~\new_[8726]_ );
  assign \new_[4571]_  = ~\new_[4704]_  & (~\new_[6763]_  | ~\new_[1460]_ );
  assign \new_[4572]_  = ~\new_[4705]_  & (~\new_[6770]_  | ~\new_[8101]_ );
  assign \new_[4573]_  = ~\new_[4706]_  & (~\new_[6785]_  | ~\new_[1143]_ );
  assign \new_[4574]_  = ~\new_[4708]_  & (~\new_[7097]_  | ~\new_[1098]_ );
  assign \new_[4575]_  = ~\new_[4707]_  & (~\new_[6770]_  | ~\new_[1242]_ );
  assign \new_[4576]_  = ~\new_[4710]_  & (~\new_[6785]_  | ~\new_[1210]_ );
  assign \new_[4577]_  = ~\new_[4709]_  & (~\new_[6785]_  | ~\new_[1094]_ );
  assign \new_[4578]_  = ~\new_[4711]_  & (~\new_[6785]_  | ~\new_[1194]_ );
  assign \new_[4579]_  = ~\new_[4689]_  & (~\new_[6785]_  | ~\new_[1218]_ );
  assign \new_[4580]_  = ~\new_[4712]_  & (~\new_[6770]_  | ~\new_[1097]_ );
  assign \new_[4581]_  = ~\new_[4713]_  & (~\new_[6785]_  | ~\new_[1195]_ );
  assign \new_[4582]_  = ~\new_[4714]_  & (~\new_[6785]_  | ~\new_[1225]_ );
  assign \new_[4583]_  = ~\new_[6774]_  & (~\new_[4959]_  | ~\new_[4851]_ );
  assign \new_[4584]_  = ~\new_[6774]_  & (~\new_[4984]_  | ~\new_[4852]_ );
  assign \new_[4585]_  = ~\new_[6774]_  & (~\new_[4960]_  | ~\new_[4853]_ );
  assign \new_[4586]_  = ~\new_[6774]_  & (~\new_[4962]_  | ~\new_[4854]_ );
  assign \new_[4587]_  = ~\new_[6784]_  & (~\new_[4963]_  | ~\new_[4855]_ );
  assign \new_[4588]_  = ~\new_[6774]_  & (~\new_[4964]_  | ~\new_[4856]_ );
  assign \new_[4589]_  = ~\new_[6784]_  & (~\new_[4961]_  | ~\new_[4857]_ );
  assign \new_[4590]_  = ~\new_[6784]_  & (~\new_[4965]_  | ~\new_[4858]_ );
  assign \new_[4591]_  = ~\new_[6774]_  & (~\new_[4968]_  | ~\new_[4859]_ );
  assign \new_[4592]_  = ~\new_[6774]_  & (~\new_[4969]_  | ~\new_[4862]_ );
  assign \new_[4593]_  = ~\new_[6774]_  & (~\new_[4970]_  | ~\new_[4860]_ );
  assign \new_[4594]_  = ~\new_[6784]_  & (~\new_[4967]_  | ~\new_[4861]_ );
  assign \new_[4595]_  = ~\new_[6784]_  & (~\new_[4971]_  | ~\new_[4863]_ );
  assign \new_[4596]_  = ~\new_[6784]_  & (~\new_[4972]_  | ~\new_[4864]_ );
  assign \new_[4597]_  = ~\new_[6784]_  & (~\new_[4975]_  | ~\new_[4866]_ );
  assign \new_[4598]_  = ~\new_[6774]_  & (~\new_[4973]_  | ~\new_[4865]_ );
  assign \new_[4599]_  = ~\new_[6784]_  & (~\new_[4977]_  | ~\new_[4867]_ );
  assign \new_[4600]_  = ~\new_[6764]_  & (~\new_[4976]_  | ~\new_[4868]_ );
  assign \new_[4601]_  = ~\new_[6784]_  & (~\new_[4979]_  | ~\new_[4872]_ );
  assign \new_[4602]_  = ~\new_[7097]_  & (~\new_[4978]_  | ~\new_[4869]_ );
  assign \new_[4603]_  = ~\new_[6774]_  & (~\new_[4966]_  | ~\new_[4875]_ );
  assign \new_[4604]_  = ~\new_[6774]_  & (~\new_[4974]_  | ~\new_[4873]_ );
  assign \new_[4605]_  = ~\new_[6764]_  & (~\new_[4957]_  | ~\new_[4871]_ );
  assign \new_[4606]_  = ~\new_[6774]_  & (~\new_[4980]_  | ~\new_[4870]_ );
  assign \new_[4607]_  = ~\new_[6784]_  & (~\new_[4981]_  | ~\new_[4874]_ );
  assign \new_[4608]_  = ~\new_[6784]_  & (~\new_[4982]_  | ~\new_[4876]_ );
  assign \new_[4609]_  = ~\new_[6784]_  & (~\new_[4983]_  | ~\new_[4877]_ );
  assign \new_[4610]_  = ~\new_[6784]_  & (~\new_[4985]_  | ~\new_[4878]_ );
  assign \new_[4611]_  = ~\new_[6784]_  & (~\new_[4986]_  | ~\new_[4880]_ );
  assign \new_[4612]_  = ~\new_[6774]_  & (~\new_[4987]_  | ~\new_[4879]_ );
  assign \new_[4613]_  = ~\new_[6774]_  & (~\new_[4988]_  | ~\new_[4881]_ );
  assign \new_[4614]_  = ~\new_[6774]_  & (~\new_[4989]_  | ~\new_[4882]_ );
  assign \new_[4615]_  = ~\new_[6784]_  & (~\new_[4991]_  | ~\new_[4848]_ );
  assign \new_[4616]_  = ~\new_[6774]_  & (~\new_[4990]_  | ~\new_[4883]_ );
  assign \new_[4617]_  = (~\new_[4885]_  | ~\new_[8966]_ ) & (~\new_[7568]_  | ~\new_[8967]_ );
  assign \new_[4618]_  = (~\new_[4887]_  | ~\new_[8966]_ ) & (~\new_[7649]_  | ~\new_[9001]_ );
  assign \new_[4619]_  = (~\new_[4886]_  | ~\new_[9000]_ ) & (~\new_[7575]_  | ~\new_[9001]_ );
  assign \new_[4620]_  = (~\new_[4888]_  | ~\new_[9000]_ ) & (~\new_[7578]_  | ~\new_[9001]_ );
  assign \new_[4621]_  = (~\new_[4890]_  | ~\new_[8966]_ ) & (~\new_[7651]_  | ~\new_[8967]_ );
  assign \new_[4622]_  = ~\new_[6602]_  & ~\new_[4797]_ ;
  assign \new_[4623]_  = ~\new_[7146]_  & ~\new_[4797]_ ;
  assign \new_[4624]_  = \new_[8964]_  & \new_[7928]_ ;
  assign \new_[4625]_  = \new_[8967]_  & \new_[7916]_ ;
  assign \new_[4626]_  = \new_[8967]_  & \new_[7918]_ ;
  assign \new_[4627]_  = ~\new_[4718]_ ;
  assign \new_[4628]_  = ~\new_[4829]_  & (~\new_[6786]_  | ~\new_[1319]_ );
  assign \new_[4629]_  = ~\new_[4830]_  & (~\new_[6786]_  | ~\new_[1207]_ );
  assign \new_[4630]_  = ~\new_[4832]_  & (~\new_[6786]_  | ~\new_[1147]_ );
  assign \new_[4631]_  = ~\new_[4831]_  & (~\new_[6786]_  | ~\new_[1149]_ );
  assign \new_[4632]_  = ~\new_[4833]_  & (~\new_[6786]_  | ~\new_[1463]_ );
  assign \new_[4633]_  = ~\new_[4834]_  & (~\new_[6786]_  | ~\new_[1322]_ );
  assign \new_[4634]_  = ~\new_[4835]_  & (~\new_[6786]_  | ~\new_[1206]_ );
  assign \new_[4635]_  = ~\new_[4841]_  & (~\new_[6786]_  | ~\new_[1103]_ );
  assign \new_[4636]_  = ~\new_[4836]_  & (~\new_[6786]_  | ~\new_[1216]_ );
  assign \new_[4637]_  = ~\new_[4838]_  & (~\new_[6763]_  | ~\new_[1530]_ );
  assign \new_[4638]_  = ~\new_[4837]_  & (~\new_[6785]_  | ~\new_[1215]_ );
  assign \new_[4639]_  = ~\new_[4839]_  & (~\new_[6786]_  | ~\new_[1106]_ );
  assign \new_[4640]_  = ~\new_[4840]_  & (~\new_[6786]_  | ~\new_[1115]_ );
  assign \new_[4641]_  = ~\new_[4842]_  & (~\new_[6786]_  | ~\new_[1107]_ );
  assign \new_[4642]_  = ~\new_[4843]_  & (~\new_[6786]_  | ~\new_[1114]_ );
  assign \new_[4643]_  = ~\new_[4845]_  & (~\new_[6786]_  | ~\new_[1315]_ );
  assign \new_[4644]_  = ~\new_[4844]_  & (~\new_[6786]_  | ~\new_[1219]_ );
  assign \new_[4645]_  = ~\new_[4846]_  & (~\new_[6786]_  | ~\new_[1208]_ );
  assign \new_[4646]_  = ~\new_[4847]_  & (~\new_[6786]_  | ~\new_[1102]_ );
  assign \new_[4647]_  = ~\new_[4743]_  & (~\new_[6785]_  | ~\new_[1203]_ );
  assign \new_[4648]_  = ~\new_[4744]_  & (~\new_[6786]_  | ~\new_[1204]_ );
  assign \new_[4649]_  = ~\new_[4747]_  & (~\new_[6786]_  | ~\new_[1202]_ );
  assign \new_[4650]_  = ~\new_[4745]_  & (~\new_[6785]_  | ~\new_[1150]_ );
  assign \new_[4651]_  = ~\new_[4746]_  & (~\new_[6786]_  | ~\new_[1520]_ );
  assign \new_[4652]_  = ~\new_[4749]_  & (~\new_[6786]_  | ~\new_[1105]_ );
  assign \new_[4653]_  = ~\new_[4748]_  & (~\new_[6786]_  | ~\new_[1323]_ );
  assign \new_[4654]_  = ~\new_[4750]_  & (~\new_[6786]_  | ~\new_[1221]_ );
  assign \new_[4655]_  = ~\new_[4756]_  & (~\new_[6785]_  | ~\new_[7939]_ );
  assign \new_[4656]_  = ~\new_[4751]_  & (~\new_[6786]_  | ~\new_[1116]_ );
  assign \new_[4657]_  = ~\new_[4753]_  & (~\new_[6786]_  | ~\new_[1104]_ );
  assign \new_[4658]_  = ~\new_[4752]_  & (~\new_[6786]_  | ~\new_[1117]_ );
  assign \new_[4659]_  = ~\new_[4754]_  & (~\new_[6786]_  | ~\new_[1222]_ );
  assign \new_[4660]_  = ~\new_[4755]_  & (~\new_[6785]_  | ~\new_[1226]_ );
  assign \new_[4661]_  = ~\new_[4757]_  & (~\new_[6786]_  | ~\new_[1205]_ );
  assign \new_[4662]_  = ~\new_[4758]_  & (~\new_[6786]_  | ~\new_[1209]_ );
  assign \new_[4663]_  = ~\new_[4759]_  & (~\new_[6786]_  | ~\new_[1538]_ );
  assign \new_[4664]_  = ~\new_[4760]_  & (~\new_[6786]_  | ~\new_[1237]_ );
  assign \new_[4665]_  = ~\new_[4761]_  & (~\new_[6785]_  | ~\new_[1151]_ );
  assign \new_[4666]_  = ~\new_[4762]_  & (~\new_[6786]_  | ~\new_[1464]_ );
  assign \new_[4667]_  = ~\new_[4763]_  & (~\new_[6786]_  | ~\new_[1214]_ );
  assign \new_[4668]_  = ~\new_[4764]_  & (~\new_[6786]_  | ~\new_[1324]_ );
  assign \new_[4669]_  = ~\new_[4765]_  & (~\new_[6786]_  | ~\new_[1240]_ );
  assign \new_[4670]_  = ~\new_[4766]_  & (~\new_[6786]_  | ~\new_[1108]_ );
  assign \new_[4671]_  = ~\new_[4767]_  & (~\new_[6785]_  | ~\new_[1109]_ );
  assign \new_[4672]_  = ~\new_[4768]_  & (~\new_[6786]_  | ~\new_[1238]_ );
  assign \new_[4673]_  = ~\new_[4769]_  & (~\new_[6786]_  | ~\new_[1152]_ );
  assign \new_[4674]_  = ~\new_[4770]_  & (~\new_[6786]_  | ~\new_[1521]_ );
  assign \new_[4675]_  = ~\new_[4771]_  & (~\new_[6786]_  | ~\new_[1220]_ );
  assign \new_[4676]_  = ~\new_[4772]_  & (~\new_[6786]_  | ~\new_[1321]_ );
  assign \new_[4677]_  = ~\new_[4773]_  & (~\new_[6786]_  | ~\new_[1211]_ );
  assign \new_[4678]_  = ~\new_[4774]_  & (~\new_[6786]_  | ~\new_[1212]_ );
  assign \new_[4679]_  = ~\new_[4775]_  & (~\new_[6786]_  | ~\new_[1110]_ );
  assign \new_[4680]_  = ~\new_[4776]_  & (~\new_[6763]_  | ~\new_[1111]_ );
  assign \new_[4681]_  = ~\new_[4777]_  & (~\new_[6786]_  | ~\new_[1213]_ );
  assign \new_[4682]_  = ~\new_[4778]_  & (~\new_[6785]_  | ~\new_[1148]_ );
  assign \new_[4683]_  = ~\new_[4779]_  & (~\new_[6786]_  | ~\new_[1234]_ );
  assign \new_[4684]_  = ~\new_[4780]_  & (~\new_[6763]_  | ~\new_[1461]_ );
  assign \new_[4685]_  = ~\new_[6774]_  & (~\new_[4956]_  | ~\new_[4849]_ );
  assign \new_[4686]_  = ~\new_[6774]_  & (~\new_[4958]_  | ~\new_[4850]_ );
  assign \new_[4687]_  = ~\new_[6763]_  & (~\new_[5086]_  | ~\new_[4906]_ );
  assign \new_[4688]_  = ~\new_[6774]_  & (~\new_[5087]_  | ~\new_[4907]_ );
  assign \new_[4689]_  = ~\new_[6784]_  & (~\new_[5088]_  | ~\new_[4908]_ );
  assign \new_[4690]_  = ~\new_[6784]_  & (~\new_[5089]_  | ~\new_[4909]_ );
  assign \new_[4691]_  = ~\new_[6764]_  & (~\new_[5101]_  | ~\new_[4921]_ );
  assign \new_[4692]_  = ~\new_[6784]_  & (~\new_[5090]_  | ~\new_[4910]_ );
  assign \new_[4693]_  = ~\new_[6784]_  & (~\new_[5091]_  | ~\new_[4911]_ );
  assign \new_[4694]_  = ~\new_[6784]_  & (~\new_[5093]_  | ~\new_[4913]_ );
  assign \new_[4695]_  = ~\new_[6784]_  & (~\new_[5092]_  | ~\new_[4912]_ );
  assign \new_[4696]_  = ~\new_[6784]_  & (~\new_[5094]_  | ~\new_[4914]_ );
  assign \new_[4697]_  = ~\new_[6784]_  & (~\new_[5095]_  | ~\new_[4915]_ );
  assign \new_[4698]_  = ~\new_[6774]_  & (~\new_[5096]_  | ~\new_[4916]_ );
  assign \new_[4699]_  = ~\new_[6784]_  & (~\new_[5098]_  | ~\new_[4917]_ );
  assign \new_[4700]_  = ~\new_[6774]_  & (~\new_[5099]_  | ~\new_[4920]_ );
  assign \new_[4701]_  = ~\new_[6764]_  & (~\new_[5100]_  | ~\new_[4919]_ );
  assign \new_[4702]_  = ~\new_[6774]_  & (~\new_[5097]_  | ~\new_[4918]_ );
  assign \new_[4703]_  = ~\new_[6774]_  & (~\new_[5102]_  | ~\new_[4922]_ );
  assign \new_[4704]_  = ~\new_[6785]_  & (~\new_[5103]_  | ~\new_[4923]_ );
  assign \new_[4705]_  = ~\new_[6784]_  & (~\new_[5104]_  | ~\new_[4924]_ );
  assign \new_[4706]_  = ~\new_[6774]_  & (~\new_[5105]_  | ~\new_[4925]_ );
  assign \new_[4707]_  = ~\new_[6764]_  & (~\new_[5106]_  | ~\new_[4927]_ );
  assign \new_[4708]_  = ~\new_[6784]_  & (~\new_[5107]_  | ~\new_[4926]_ );
  assign \new_[4709]_  = ~\new_[6784]_  & (~\new_[5109]_  | ~\new_[4930]_ );
  assign \new_[4710]_  = ~\new_[6774]_  & (~\new_[5108]_  | ~\new_[4928]_ );
  assign \new_[4711]_  = ~\new_[6774]_  & (~\new_[5110]_  | ~\new_[4929]_ );
  assign \new_[4712]_  = ~\new_[6784]_  & (~\new_[5111]_  | ~\new_[4931]_ );
  assign \new_[4713]_  = ~\new_[6784]_  & (~\new_[5112]_  | ~\new_[4933]_ );
  assign \new_[4714]_  = ~\new_[6784]_  & (~\new_[5113]_  | ~\new_[4932]_ );
  assign \new_[4715]_  = ~\new_[2134]_  | ~\new_[8726]_ ;
  assign \new_[4716]_  = ~\new_[2131]_  | ~\new_[8726]_ ;
  assign \new_[4717]_  = ~\new_[5114]_  | ~\new_[6198]_  | ~\new_[6035]_ ;
  assign \new_[4718]_  = ~\new_[5114]_  | ~\new_[8965]_ ;
  assign \new_[4719]_  = \new_[5486]_  ^ \new_[8495]_ ;
  assign \new_[4720]_  = \new_[5487]_  ^ \new_[8523]_ ;
  assign \new_[4721]_  = ~\new_[4362]_  | ~\new_[4884]_  | ~\new_[7843]_ ;
  assign \new_[4722]_  = \new_[8496]_  ^ \new_[4996]_ ;
  assign \new_[4723]_  = \new_[5251]_  ^ \new_[4997]_ ;
  assign \new_[4724]_  = \new_[8527]_  ^ \new_[4998]_ ;
  assign \new_[4725]_  = \new_[8751]_  ^ \new_[4999]_ ;
  assign \new_[4726]_  = \new_[5000]_  ^ \new_[8496]_ ;
  assign \new_[4727]_  = \new_[8527]_  ^ \new_[5002]_ ;
  assign \new_[4728]_  = \new_[8601]_  ^ \new_[5003]_ ;
  assign \new_[4729]_  = ~\new_[8411]_ ;
  assign \new_[4730]_  = \new_[8636]_  ^ \new_[5001]_ ;
  assign \new_[4731]_  = \new_[5007]_  ^ \new_[4895]_ ;
  assign \new_[4732]_  = \new_[5006]_  ^ \new_[4896]_ ;
  assign \new_[4733]_  = \new_[5009]_  ^ \new_[4898]_ ;
  assign \new_[4734]_  = \new_[5011]_  ^ \new_[4897]_ ;
  assign \new_[4735]_  = ~\new_[8660]_ ;
  assign \new_[4736]_  = ~\new_[6774]_  & (~\new_[5079]_  | ~\new_[4899]_ );
  assign \new_[4737]_  = ~\new_[6774]_  & (~\new_[5080]_  | ~\new_[4900]_ );
  assign \new_[4738]_  = ~\new_[6774]_  & (~\new_[5081]_  | ~\new_[4901]_ );
  assign \new_[4739]_  = ~\new_[6774]_  & (~\new_[5082]_  | ~\new_[4902]_ );
  assign \new_[4740]_  = ~\new_[6774]_  & (~\new_[5083]_  | ~\new_[4903]_ );
  assign \new_[4741]_  = ~\new_[6774]_  & (~\new_[5084]_  | ~\new_[4905]_ );
  assign \new_[4742]_  = ~\new_[7097]_  & (~\new_[5085]_  | ~\new_[4904]_ );
  assign \new_[4743]_  = ~\new_[6764]_  & (~\new_[5164]_  | ~\new_[5032]_ );
  assign \new_[4744]_  = ~\new_[6763]_  & (~\new_[5165]_  | ~\new_[5034]_ );
  assign \new_[4745]_  = ~\new_[6763]_  & (~\new_[5166]_  | ~\new_[5035]_ );
  assign \new_[4746]_  = ~\new_[6764]_  & (~\new_[5167]_  | ~\new_[5036]_ );
  assign \new_[4747]_  = ~\new_[6763]_  & (~\new_[5168]_  | ~\new_[5040]_ );
  assign \new_[4748]_  = ~\new_[7097]_  & (~\new_[5169]_  | ~\new_[5037]_ );
  assign \new_[4749]_  = ~\new_[6764]_  & (~\new_[5170]_  | ~\new_[5039]_ );
  assign \new_[4750]_  = ~\new_[6764]_  & (~\new_[5155]_  | ~\new_[5038]_ );
  assign \new_[4751]_  = ~\new_[6764]_  & (~\new_[5171]_  | ~\new_[5041]_ );
  assign \new_[4752]_  = ~\new_[7097]_  & (~\new_[5172]_  | ~\new_[5019]_ );
  assign \new_[4753]_  = ~\new_[7097]_  & (~\new_[5173]_  | ~\new_[5043]_ );
  assign \new_[4754]_  = ~\new_[6763]_  & (~\new_[5174]_  | ~\new_[5042]_ );
  assign \new_[4755]_  = ~\new_[6784]_  & (~\new_[5185]_  | ~\new_[5044]_ );
  assign \new_[4756]_  = ~\new_[6784]_  & (~\new_[5175]_  | ~\new_[5045]_ );
  assign \new_[4757]_  = ~\new_[6763]_  & (~\new_[5176]_  | ~\new_[5047]_ );
  assign \new_[4758]_  = ~\new_[6764]_  & (~\new_[5177]_  | ~\new_[5048]_ );
  assign \new_[4759]_  = ~\new_[6763]_  & (~\new_[5178]_  | ~\new_[5049]_ );
  assign \new_[4760]_  = ~\new_[6763]_  & (~\new_[5179]_  | ~\new_[5050]_ );
  assign \new_[4761]_  = ~\new_[6764]_  & (~\new_[5180]_  | ~\new_[5051]_ );
  assign \new_[4762]_  = ~\new_[6764]_  & (~\new_[5181]_  | ~\new_[5052]_ );
  assign \new_[4763]_  = ~\new_[6763]_  & (~\new_[5182]_  | ~\new_[5053]_ );
  assign \new_[4764]_  = ~\new_[6763]_  & (~\new_[5183]_  | ~\new_[5054]_ );
  assign \new_[4765]_  = ~\new_[6763]_  & (~\new_[5188]_  | ~\new_[5055]_ );
  assign \new_[4766]_  = ~\new_[6764]_  & (~\new_[5184]_  | ~\new_[5056]_ );
  assign \new_[4767]_  = ~\new_[6763]_  & (~\new_[5186]_  | ~\new_[5057]_ );
  assign \new_[4768]_  = ~\new_[6763]_  & (~\new_[5187]_  | ~\new_[5058]_ );
  assign \new_[4769]_  = ~\new_[7097]_  & (~\new_[5190]_  | ~\new_[5059]_ );
  assign \new_[4770]_  = ~\new_[6764]_  & (~\new_[5191]_  | ~\new_[5060]_ );
  assign \new_[4771]_  = ~\new_[6764]_  & (~\new_[5189]_  | ~\new_[5046]_ );
  assign \new_[4772]_  = ~\new_[6763]_  & (~\new_[5192]_  | ~\new_[5061]_ );
  assign \new_[4773]_  = ~\new_[6764]_  & (~\new_[5193]_  | ~\new_[5062]_ );
  assign \new_[4774]_  = ~\new_[6763]_  & (~\new_[5194]_  | ~\new_[5063]_ );
  assign \new_[4775]_  = ~\new_[6764]_  & (~\new_[5195]_  | ~\new_[5064]_ );
  assign \new_[4776]_  = ~\new_[6763]_  & (~\new_[5196]_  | ~\new_[5065]_ );
  assign \new_[4777]_  = ~\new_[6763]_  & (~\new_[5197]_  | ~\new_[5066]_ );
  assign \new_[4778]_  = ~\new_[6763]_  & (~\new_[5198]_  | ~\new_[5067]_ );
  assign \new_[4779]_  = ~\new_[6764]_  & (~\new_[5200]_  | ~\new_[5013]_ );
  assign \new_[4780]_  = ~\new_[6763]_  & (~\new_[5199]_  | ~\new_[5068]_ );
  assign \new_[4781]_  = ~\new_[4935]_  & (~\new_[6499]_  | ~\new_[5115]_ );
  assign \new_[4782]_  = ~\new_[4936]_  & (~\new_[6500]_  | ~\new_[5202]_ );
  assign \new_[4783]_  = \new_[4937]_  | \new_[4938]_ ;
  assign \new_[4784]_  = ~\new_[4940]_  & (~\new_[6502]_  | ~\new_[8310]_ );
  assign \new_[4785]_  = ~\new_[4944]_  & (~\new_[6507]_  | ~\new_[8310]_ );
  assign \new_[4786]_  = (~\new_[6385]_  | ~\new_[8727]_ ) & (~\key_i[8]  | ~\new_[5253]_ );
  assign \new_[4787]_  = \new_[5073]_  | \new_[4946]_ ;
  assign \new_[4788]_  = \new_[5074]_  | \new_[4947]_ ;
  assign \new_[4789]_  = \key_i[13]  ? \new_[8727]_  : \new_[6505]_ ;
  assign \new_[4790]_  = ~\new_[4948]_  & (~\new_[6506]_  | ~\new_[8310]_ );
  assign \new_[4791]_  = \new_[4949]_  | \new_[4950]_ ;
  assign \new_[4792]_  = (~\new_[6186]_  | ~\new_[5114]_ ) & (~\key_i[21]  | ~\new_[5253]_ );
  assign \new_[4793]_  = ~\new_[4951]_  | (~\new_[6384]_  & ~\new_[8307]_ );
  assign \new_[4794]_  = ~\new_[4952]_  & (~\new_[6503]_  | ~\new_[5115]_ );
  assign \new_[4795]_  = ~\new_[4954]_  & (~\new_[6508]_  | ~\new_[5202]_ );
  assign \new_[4796]_  = ~\new_[4955]_  & (~\new_[6509]_  | ~\new_[5115]_ );
  assign \new_[4797]_  = ~\new_[5114]_  | ~\new_[8993]_ ;
  assign \new_[4798]_  = ~\new_[5114]_ ;
  assign \new_[4799]_  = \new_[5289]_  ^ \new_[5116]_ ;
  assign \new_[4800]_  = \new_[5243]_  ^ \new_[5118]_ ;
  assign \new_[4801]_  = \new_[5290]_  ^ \new_[5119]_ ;
  assign \new_[4802]_  = \new_[5245]_  ^ \new_[5121]_ ;
  assign \new_[4803]_  = \new_[5291]_  ^ \new_[5122]_ ;
  assign \new_[4804]_  = \new_[5243]_  ^ \new_[5124]_ ;
  assign \new_[4805]_  = \new_[5292]_  ^ \new_[5125]_ ;
  assign \new_[4806]_  = \new_[5245]_  ^ \new_[5127]_ ;
  assign \new_[4807]_  = \new_[5306]_  ^ \new_[8163]_ ;
  assign \new_[4808]_  = \new_[8739]_  ^ \new_[5129]_ ;
  assign \new_[4809]_  = \new_[5130]_  ^ \new_[8758]_ ;
  assign \new_[4810]_  = \new_[5429]_  ^ \new_[5141]_ ;
  assign \new_[4811]_  = \new_[5310]_  ^ \new_[5132]_ ;
  assign \new_[4812]_  = \new_[8790]_  ^ \new_[5133]_ ;
  assign \new_[4813]_  = \new_[5430]_  ^ \new_[5134]_ ;
  assign \new_[4814]_  = \new_[8691]_  ^ \new_[5135]_ ;
  assign \new_[4815]_  = \new_[5136]_  ^ \new_[8736]_ ;
  assign \new_[4816]_  = \new_[5429]_  ^ \new_[5137]_ ;
  assign \new_[4817]_  = \new_[5308]_  ^ \new_[5138]_ ;
  assign \new_[4818]_  = \new_[8441]_  ^ \new_[5139]_ ;
  assign \new_[4819]_  = \new_[5430]_  ^ \new_[5140]_ ;
  assign \new_[4820]_  = \new_[8797]_  ^ \new_[5004]_ ;
  assign \new_[4821]_  = \new_[8857]_  ^ \new_[5005]_ ;
  assign \new_[4822]_  = \new_[8762]_  ^ \new_[5011]_ ;
  assign \new_[4823]_  = \new_[8797]_  ^ \new_[5007]_ ;
  assign \new_[4824]_  = \new_[8762]_  ^ \new_[5008]_ ;
  assign \new_[4825]_  = \new_[8857]_  ^ \new_[5009]_ ;
  assign \new_[4826]_  = \new_[8444]_  ^ \new_[5006]_ ;
  assign \new_[4827]_  = ~\new_[8661]_ ;
  assign \new_[4828]_  = \new_[8444]_  ^ \new_[5010]_ ;
  assign \new_[4829]_  = ~\new_[6764]_  & (~\new_[5144]_  | ~\new_[5012]_ );
  assign \new_[4830]_  = ~\new_[6763]_  & (~\new_[5145]_  | ~\new_[5014]_ );
  assign \new_[4831]_  = ~\new_[6763]_  & (~\new_[5146]_  | ~\new_[5015]_ );
  assign \new_[4832]_  = ~\new_[6764]_  & (~\new_[5147]_  | ~\new_[5016]_ );
  assign \new_[4833]_  = ~\new_[6763]_  & (~\new_[5148]_  | ~\new_[5017]_ );
  assign \new_[4834]_  = ~\new_[6763]_  & (~\new_[5149]_  | ~\new_[5018]_ );
  assign \new_[4835]_  = ~\new_[6764]_  & (~\new_[5150]_  | ~\new_[5020]_ );
  assign \new_[4836]_  = ~\new_[6764]_  & (~\new_[5151]_  | ~\new_[5021]_ );
  assign \new_[4837]_  = ~\new_[6764]_  & (~\new_[5153]_  | ~\new_[5022]_ );
  assign \new_[4838]_  = ~\new_[6764]_  & (~\new_[5154]_  | ~\new_[5023]_ );
  assign \new_[4839]_  = ~\new_[6763]_  & (~\new_[5156]_  | ~\new_[5024]_ );
  assign \new_[4840]_  = ~\new_[6764]_  & (~\new_[5157]_  | ~\new_[5025]_ );
  assign \new_[4841]_  = ~\new_[6764]_  & (~\new_[5152]_  | ~\new_[5026]_ );
  assign \new_[4842]_  = ~\new_[6763]_  & (~\new_[5158]_  | ~\new_[5028]_ );
  assign \new_[4843]_  = ~\new_[6764]_  & (~\new_[5159]_  | ~\new_[5027]_ );
  assign \new_[4844]_  = ~\new_[6764]_  & (~\new_[5160]_  | ~\new_[5029]_ );
  assign \new_[4845]_  = ~\new_[6764]_  & (~\new_[5161]_  | ~\new_[5031]_ );
  assign \new_[4846]_  = ~\new_[6764]_  & (~\new_[5162]_  | ~\new_[5030]_ );
  assign \new_[4847]_  = ~\new_[6764]_  & (~\new_[5163]_  | ~\new_[5033]_ );
  assign \new_[4848]_  = (~\new_[7673]_  | ~\new_[6788]_ ) & (~\new_[5239]_  | ~\new_[6914]_ );
  assign \new_[4849]_  = (~\new_[7666]_  | ~\new_[7115]_ ) & (~\new_[5204]_  | ~\new_[6638]_ );
  assign \new_[4850]_  = (~\new_[7772]_  | ~\new_[6788]_ ) & (~\new_[5223]_  | ~\new_[6638]_ );
  assign \new_[4851]_  = (~\new_[7665]_  | ~\new_[6788]_ ) & (~\new_[5205]_  | ~\new_[6638]_ );
  assign \new_[4852]_  = (~\new_[7677]_  | ~\new_[6788]_ ) & (~\new_[5206]_  | ~\new_[6638]_ );
  assign \new_[4853]_  = (~\new_[7758]_  | ~\new_[6788]_ ) & (~\new_[5207]_  | ~\new_[6638]_ );
  assign \new_[4854]_  = (~\new_[7783]_  | ~\new_[6788]_ ) & (~\new_[5211]_  | ~\new_[6638]_ );
  assign \new_[4855]_  = (~\new_[7704]_  | ~\new_[6788]_ ) & (~\new_[5208]_  | ~\new_[6914]_ );
  assign \new_[4856]_  = (~\new_[7712]_  | ~\new_[6788]_ ) & (~\new_[5209]_  | ~\new_[6914]_ );
  assign \new_[4857]_  = (~\new_[7714]_  | ~\new_[6788]_ ) & (~\new_[5210]_  | ~\new_[6638]_ );
  assign \new_[4858]_  = (~\new_[7778]_  | ~\new_[6788]_ ) & (~\new_[5212]_  | ~\new_[6638]_ );
  assign \new_[4859]_  = (~\new_[7775]_  | ~\new_[6788]_ ) & (~\new_[5213]_  | ~\new_[6638]_ );
  assign \new_[4860]_  = (~\new_[7803]_  | ~\new_[6788]_ ) & (~\new_[5215]_  | ~\new_[6638]_ );
  assign \new_[4861]_  = (~\new_[7812]_  | ~\new_[6788]_ ) & (~\new_[5216]_  | ~\new_[6638]_ );
  assign \new_[4862]_  = (~\new_[7808]_  | ~\new_[6788]_ ) & (~\new_[5214]_  | ~\new_[6638]_ );
  assign \new_[4863]_  = (~\new_[7749]_  | ~\new_[6788]_ ) & (~\new_[5218]_  | ~\new_[6638]_ );
  assign \new_[4864]_  = (~\new_[7806]_  | ~\new_[6788]_ ) & (~\new_[5219]_  | ~\new_[6638]_ );
  assign \new_[4865]_  = (~\new_[7723]_  | ~\new_[6788]_ ) & (~\new_[5220]_  | ~\new_[6638]_ );
  assign \new_[4866]_  = (~\new_[7667]_  | ~\new_[6788]_ ) & (~\new_[5221]_  | ~\new_[6638]_ );
  assign \new_[4867]_  = (~\new_[7782]_  | ~\new_[7115]_ ) & (~\new_[5222]_  | ~\new_[6638]_ );
  assign \new_[4868]_  = (~\new_[7777]_  | ~\new_[6788]_ ) & (~\new_[5235]_  | ~\new_[6638]_ );
  assign \new_[4869]_  = (~\new_[7695]_  | ~\new_[7115]_ ) & (~\new_[5226]_  | ~\new_[6638]_ );
  assign \new_[4870]_  = (~\new_[7737]_  | ~\new_[6788]_ ) & (~\new_[5228]_  | ~\new_[6638]_ );
  assign \new_[4871]_  = (~\new_[7801]_  | ~\new_[6788]_ ) & (~\new_[5224]_  | ~\new_[6638]_ );
  assign \new_[4872]_  = (~\new_[7670]_  | ~\new_[7115]_ ) & (~\new_[5227]_  | ~\new_[6638]_ );
  assign \new_[4873]_  = (~\new_[7684]_  | ~\new_[6788]_ ) & (~\new_[5217]_  | ~\new_[6638]_ );
  assign \new_[4874]_  = (~\new_[7750]_  | ~\new_[6788]_ ) & (~\new_[5229]_  | ~\new_[6638]_ );
  assign \new_[4875]_  = (~\new_[7633]_  | ~\new_[6788]_ ) & (~\new_[5225]_  | ~\new_[6638]_ );
  assign \new_[4876]_  = (~\new_[7787]_  | ~\new_[6788]_ ) & (~\new_[5230]_  | ~\new_[6638]_ );
  assign \new_[4877]_  = (~\new_[7746]_  | ~\new_[6788]_ ) & (~\new_[5231]_  | ~\new_[6638]_ );
  assign \new_[4878]_  = (~\new_[7647]_  | ~\new_[6788]_ ) & (~\new_[5232]_  | ~\new_[6638]_ );
  assign \new_[4879]_  = (~\new_[7717]_  | ~\new_[6788]_ ) & (~\new_[5234]_  | ~\new_[6638]_ );
  assign \new_[4880]_  = (~\new_[7692]_  | ~\new_[6788]_ ) & (~\new_[5233]_  | ~\new_[6638]_ );
  assign \new_[4881]_  = (~\new_[7685]_  | ~\new_[6788]_ ) & (~\new_[5236]_  | ~\new_[6638]_ );
  assign \new_[4882]_  = (~\new_[7811]_  | ~\new_[6788]_ ) & (~\new_[5237]_  | ~\new_[6914]_ );
  assign \new_[4883]_  = (~\new_[7689]_  | ~\new_[6788]_ ) & (~\new_[5238]_  | ~\new_[6638]_ );
  assign \new_[4884]_  = ~\new_[4934]_ ;
  assign \new_[4885]_  = \new_[5069]_  | \new_[5070]_ ;
  assign \new_[4886]_  = ~\new_[5072]_  | (~\new_[6386]_  & ~\new_[8307]_ );
  assign \new_[4887]_  = (~\new_[6387]_  & ~\new_[5203]_ ) | (~\new_[8135]_  & ~\new_[5202]_ );
  assign \new_[4888]_  = ~\new_[5076]_  | (~\new_[6388]_  & ~\new_[5201]_ );
  assign \new_[4889]_  = \new_[5077]_  | \new_[5078]_ ;
  assign \new_[4890]_  = (~\new_[6383]_  & ~\new_[5253]_ ) | (~\new_[8131]_  & ~\new_[8308]_ );
  assign \new_[4891]_  = \new_[7596]_  | \new_[9000]_ ;
  assign \new_[4892]_  = ~\new_[7562]_  | ~\new_[9001]_ ;
  assign \new_[4893]_  = \new_[7612]_  | \new_[9002]_ ;
  assign \new_[4894]_  = \new_[7611]_  | \new_[9002]_ ;
  assign \new_[4895]_  = \new_[8637]_  ^ \new_[8751]_ ;
  assign \new_[4896]_  = \new_[8754]_  ^ \new_[8601]_ ;
  assign \new_[4897]_  = \new_[8753]_  ^ \new_[5251]_ ;
  assign \new_[4898]_  = \new_[8602]_  ^ \new_[8636]_ ;
  assign \new_[4899]_  = (~\new_[7793]_  | ~\new_[6788]_ ) & (~\new_[5254]_  | ~\new_[6637]_ );
  assign \new_[4900]_  = (~\new_[7736]_  | ~\new_[6788]_ ) & (~\new_[5255]_  | ~\new_[6637]_ );
  assign \new_[4901]_  = (~\new_[7663]_  | ~\new_[6788]_ ) & (~\new_[5256]_  | ~\new_[6638]_ );
  assign \new_[4902]_  = (~\new_[7766]_  | ~\new_[6788]_ ) & (~\new_[5257]_  | ~\new_[6914]_ );
  assign \new_[4903]_  = (~\new_[7686]_  | ~\new_[6788]_ ) & (~\new_[5258]_  | ~\new_[6638]_ );
  assign \new_[4904]_  = (~\new_[7726]_  | ~\new_[6788]_ ) & (~\new_[5260]_  | ~\new_[6638]_ );
  assign \new_[4905]_  = (~\new_[7671]_  | ~\new_[6788]_ ) & (~\new_[5259]_  | ~\new_[6638]_ );
  assign \new_[4906]_  = (~\new_[7715]_  | ~\new_[6788]_ ) & (~\new_[5261]_  | ~\new_[6638]_ );
  assign \new_[4907]_  = (~\new_[7724]_  | ~\new_[6788]_ ) & (~\new_[5288]_  | ~\new_[6638]_ );
  assign \new_[4908]_  = (~\new_[7813]_  | ~\new_[6788]_ ) & (~\new_[5284]_  | ~\new_[6638]_ );
  assign \new_[4909]_  = (~\new_[7794]_  | ~\new_[6788]_ ) & (~\new_[5262]_  | ~\new_[6638]_ );
  assign \new_[4910]_  = (~\new_[7789]_  | ~\new_[6788]_ ) & (~\new_[5263]_  | ~\new_[6914]_ );
  assign \new_[4911]_  = (~\new_[7733]_  | ~\new_[6788]_ ) & (~\new_[5264]_  | ~\new_[6638]_ );
  assign \new_[4912]_  = (~\new_[7707]_  | ~\new_[6788]_ ) & (~\new_[5265]_  | ~\new_[6638]_ );
  assign \new_[4913]_  = (~\new_[7810]_  | ~\new_[6788]_ ) & (~\new_[5266]_  | ~\new_[6638]_ );
  assign \new_[4914]_  = (~\new_[7759]_  | ~\new_[6788]_ ) & (~\new_[5267]_  | ~\new_[6638]_ );
  assign \new_[4915]_  = (~\new_[7776]_  | ~\new_[6788]_ ) & (~\new_[5268]_  | ~\new_[6638]_ );
  assign \new_[4916]_  = (~\new_[7795]_  | ~\new_[6788]_ ) & (~\new_[5269]_  | ~\new_[6637]_ );
  assign \new_[4917]_  = (~\new_[7753]_  | ~\new_[6788]_ ) & (~\new_[5270]_  | ~\new_[6637]_ );
  assign \new_[4918]_  = (~\new_[7700]_  | ~\new_[6788]_ ) & (~\new_[5273]_  | ~\new_[6638]_ );
  assign \new_[4919]_  = (~\new_[7719]_  | ~\new_[6788]_ ) & (~\new_[5272]_  | ~\new_[6780]_ );
  assign \new_[4920]_  = (~\new_[7732]_  | ~\new_[6788]_ ) & (~\new_[5271]_  | ~\new_[6638]_ );
  assign \new_[4921]_  = (~\new_[7734]_  | ~\new_[6788]_ ) & (~\new_[5274]_  | ~\new_[6638]_ );
  assign \new_[4922]_  = (~\new_[7796]_  | ~\new_[6788]_ ) & (~\new_[5275]_  | ~\new_[6638]_ );
  assign \new_[4923]_  = (~\new_[7809]_  | ~\new_[6788]_ ) & (~\new_[5276]_  | ~\new_[6637]_ );
  assign \new_[4924]_  = (~\new_[7644]_  | ~\new_[6788]_ ) & (~\new_[5277]_  | ~\new_[6638]_ );
  assign \new_[4925]_  = (~\new_[7773]_  | ~\new_[6788]_ ) & (~\new_[5278]_  | ~\new_[6638]_ );
  assign \new_[4926]_  = (~\new_[7745]_  | ~\new_[6788]_ ) & (~\new_[5279]_  | ~\new_[6638]_ );
  assign \new_[4927]_  = (~\new_[7739]_  | ~\new_[6788]_ ) & (~\new_[5280]_  | ~\new_[6638]_ );
  assign \new_[4928]_  = (~\new_[7669]_  | ~\new_[6788]_ ) & (~\new_[5281]_  | ~\new_[6914]_ );
  assign \new_[4929]_  = (~\new_[7774]_  | ~\new_[6788]_ ) & (~\new_[5283]_  | ~\new_[6638]_ );
  assign \new_[4930]_  = (~\new_[7756]_  | ~\new_[6788]_ ) & (~\new_[5282]_  | ~\new_[6638]_ );
  assign \new_[4931]_  = (~\new_[7731]_  | ~\new_[6788]_ ) & (~\new_[5285]_  | ~\new_[6638]_ );
  assign \new_[4932]_  = (~\new_[7786]_  | ~\new_[6788]_ ) & (~\new_[5287]_  | ~\new_[6638]_ );
  assign \new_[4933]_  = (~\new_[7699]_  | ~\new_[6788]_ ) & (~\new_[5286]_  | ~\new_[6638]_ );
  assign \new_[4934]_  = ~\new_[5249]_  | ~\new_[5143]_ ;
  assign \new_[4935]_  = \key_i[30]  & \new_[5203]_ ;
  assign \new_[4936]_  = \key_i[31]  & \new_[5201]_ ;
  assign \new_[4937]_  = \key_i[3]  & \new_[5201]_ ;
  assign \new_[4938]_  = ~\new_[8307]_  & (~\new_[6811]_  | ~\new_[6531]_ );
  assign \new_[4939]_  = \new_[7661]_  | \new_[9002]_ ;
  assign \new_[4940]_  = \key_i[4]  & \new_[5203]_ ;
  assign \new_[4941]_  = ~\key_i[5]  | ~\new_[5203]_ ;
  assign \new_[4942]_  = ~\new_[6504]_  | ~\new_[8308]_ ;
  assign \new_[4943]_  = \new_[7641]_  | \new_[9000]_ ;
  assign \new_[4944]_  = \key_i[7]  & \new_[5203]_ ;
  assign \new_[4945]_  = \key_i[9]  & \new_[5203]_ ;
  assign \new_[4946]_  = ~\new_[5203]_  & (~\new_[6756]_  | ~\new_[6537]_ );
  assign \new_[4947]_  = ~\new_[8401]_  & (~\new_[6769]_  | ~\new_[6710]_ );
  assign \new_[4948]_  = \key_i[15]  & \new_[8307]_ ;
  assign \new_[4949]_  = \key_i[17]  & \new_[5201]_ ;
  assign \new_[4950]_  = ~\new_[5201]_  & (~\new_[6810]_  | ~\new_[6528]_ );
  assign \new_[4951]_  = \new_[7964]_  | \new_[8308]_ ;
  assign \new_[4952]_  = \key_i[25]  & \new_[5203]_ ;
  assign \new_[4953]_  = \new_[7652]_  | \new_[9000]_ ;
  assign \new_[4954]_  = \key_i[26]  & \new_[5203]_ ;
  assign \new_[4955]_  = \key_i[29]  & \new_[5203]_ ;
  assign \new_[4956]_  = ~\new_[6919]_  | ~\new_[5204]_ ;
  assign \new_[4957]_  = ~\new_[6919]_  | ~\new_[5224]_ ;
  assign \new_[4958]_  = ~\new_[6745]_  | ~\new_[5223]_ ;
  assign \new_[4959]_  = ~\new_[6745]_  | ~\new_[5205]_ ;
  assign \new_[4960]_  = ~\new_[6745]_  | ~\new_[5207]_ ;
  assign \new_[4961]_  = ~\new_[6919]_  | ~\new_[5210]_ ;
  assign \new_[4962]_  = ~\new_[6745]_  | ~\new_[5211]_ ;
  assign \new_[4963]_  = ~\new_[6745]_  | ~\new_[5208]_ ;
  assign \new_[4964]_  = ~\new_[6745]_  | ~\new_[5209]_ ;
  assign \new_[4965]_  = ~\new_[6919]_  | ~\new_[5212]_ ;
  assign \new_[4966]_  = ~\new_[6642]_  | ~\new_[5225]_ ;
  assign \new_[4967]_  = ~\new_[6919]_  | ~\new_[5216]_ ;
  assign \new_[4968]_  = ~\new_[6919]_  | ~\new_[5213]_ ;
  assign \new_[4969]_  = ~\new_[6919]_  | ~\new_[5214]_ ;
  assign \new_[4970]_  = ~\new_[6919]_  | ~\new_[5215]_ ;
  assign \new_[4971]_  = ~\new_[6745]_  | ~\new_[5218]_ ;
  assign \new_[4972]_  = ~\new_[6745]_  | ~\new_[5219]_ ;
  assign \new_[4973]_  = ~\new_[6919]_  | ~\new_[5220]_ ;
  assign \new_[4974]_  = ~\new_[6919]_  | ~\new_[5217]_ ;
  assign \new_[4975]_  = ~\new_[6745]_  | ~\new_[5221]_ ;
  assign \new_[4976]_  = ~\new_[6745]_  | ~\new_[5235]_ ;
  assign \new_[4977]_  = ~\new_[6919]_  | ~\new_[5222]_ ;
  assign \new_[4978]_  = ~\new_[6919]_  | ~\new_[5226]_ ;
  assign \new_[4979]_  = ~\new_[6745]_  | ~\new_[5227]_ ;
  assign \new_[4980]_  = ~\new_[6642]_  | ~\new_[5228]_ ;
  assign \new_[4981]_  = ~\new_[6642]_  | ~\new_[5229]_ ;
  assign \new_[4982]_  = ~\new_[6919]_  | ~\new_[5230]_ ;
  assign \new_[4983]_  = ~\new_[6745]_  | ~\new_[5231]_ ;
  assign \new_[4984]_  = ~\new_[6919]_  | ~\new_[5206]_ ;
  assign \new_[4985]_  = ~\new_[6919]_  | ~\new_[5232]_ ;
  assign \new_[4986]_  = ~\new_[6745]_  | ~\new_[5233]_ ;
  assign \new_[4987]_  = ~\new_[6642]_  | ~\new_[5234]_ ;
  assign \new_[4988]_  = ~\new_[6642]_  | ~\new_[5236]_ ;
  assign \new_[4989]_  = ~\new_[6919]_  | ~\new_[5237]_ ;
  assign \new_[4990]_  = ~\new_[6919]_  | ~\new_[5238]_ ;
  assign \new_[4991]_  = ~\new_[6745]_  | ~\new_[5239]_ ;
  assign \new_[4992]_  = \new_[5250]_  ^ \new_[8498]_ ;
  assign \new_[4993]_  = \new_[5252]_  ^ \new_[8526]_ ;
  assign \new_[4994]_  = ~\new_[5240]_  | ~\new_[5379]_ ;
  assign \new_[4995]_  = \new_[5240]_  | \new_[5379]_ ;
  assign \new_[4996]_  = \new_[5294]_  ^ \new_[8636]_ ;
  assign \new_[4997]_  = \new_[5242]_  ^ \new_[5296]_ ;
  assign \new_[4998]_  = \new_[5297]_  ^ \new_[8601]_ ;
  assign \new_[4999]_  = \new_[5244]_  ^ \new_[5299]_ ;
  assign \new_[5000]_  = \new_[5300]_  ^ \new_[5251]_ ;
  assign \new_[5001]_  = \new_[5246]_  ^ \new_[5302]_ ;
  assign \new_[5002]_  = \new_[5303]_  ^ \new_[8751]_ ;
  assign \new_[5003]_  = \new_[5247]_  ^ \new_[5305]_ ;
  assign \new_[5004]_  = \new_[8741]_  ^ \new_[5308]_ ;
  assign \new_[5005]_  = \new_[8693]_  ^ \new_[8739]_ ;
  assign \new_[5006]_  = \new_[8797]_  ^ \new_[5310]_ ;
  assign \new_[5007]_  = \new_[8444]_  ^ \new_[5308]_ ;
  assign \new_[5008]_  = \new_[8740]_  ^ \new_[8691]_ ;
  assign \new_[5009]_  = \new_[8762]_  ^ \new_[8739]_ ;
  assign \new_[5010]_  = \new_[8692]_  ^ \new_[5310]_ ;
  assign \new_[5011]_  = \new_[8857]_  ^ \new_[8691]_ ;
  assign \new_[5012]_  = (~\new_[7697]_  | ~\new_[6788]_ ) & (~\new_[5312]_  | ~\new_[6780]_ );
  assign \new_[5013]_  = (~\new_[7790]_  | ~\new_[6788]_ ) & (~\new_[5368]_  | ~\new_[6780]_ );
  assign \new_[5014]_  = (~\new_[7703]_  | ~\new_[6788]_ ) & (~\new_[5313]_  | ~\new_[6780]_ );
  assign \new_[5015]_  = (~\new_[7798]_  | ~\new_[6788]_ ) & (~\new_[5314]_  | ~\new_[6780]_ );
  assign \new_[5016]_  = (~\new_[7721]_  | ~\new_[6788]_ ) & (~\new_[5315]_  | ~\new_[6914]_ );
  assign \new_[5017]_  = (~\new_[7781]_  | ~\new_[6788]_ ) & (~\new_[5316]_  | ~\new_[6780]_ );
  assign \new_[5018]_  = (~\new_[7748]_  | ~\new_[6788]_ ) & (~\new_[5318]_  | ~\new_[6780]_ );
  assign \new_[5019]_  = (~\new_[7744]_  | ~\new_[6788]_ ) & (~\new_[5340]_  | ~\new_[6637]_ );
  assign \new_[5020]_  = (~\new_[7706]_  | ~\new_[6788]_ ) & (~\new_[5322]_  | ~\new_[6780]_ );
  assign \new_[5021]_  = (~\new_[7696]_  | ~\new_[6788]_ ) & (~\new_[5323]_  | ~\new_[6780]_ );
  assign \new_[5022]_  = (~\new_[7784]_  | ~\new_[6788]_ ) & (~\new_[5325]_  | ~\new_[6780]_ );
  assign \new_[5023]_  = (~\new_[7702]_  | ~\new_[6788]_ ) & (~\new_[5326]_  | ~\new_[6914]_ );
  assign \new_[5024]_  = (~\new_[7705]_  | ~\new_[6788]_ ) & (~\new_[5319]_  | ~\new_[6914]_ );
  assign \new_[5025]_  = (~\new_[7804]_  | ~\new_[6788]_ ) & (~\new_[5327]_  | ~\new_[6914]_ );
  assign \new_[5026]_  = (~\new_[7771]_  | ~\new_[6788]_ ) & (~\new_[5324]_  | ~\new_[6637]_ );
  assign \new_[5027]_  = (~\new_[7701]_  | ~\new_[6788]_ ) & (~\new_[5337]_  | ~\new_[6780]_ );
  assign \new_[5028]_  = (~\new_[7807]_  | ~\new_[6788]_ ) & (~\new_[5329]_  | ~\new_[6637]_ );
  assign \new_[5029]_  = (~\new_[7672]_  | ~\new_[6788]_ ) & (~\new_[5330]_  | ~\new_[6780]_ );
  assign \new_[5030]_  = (~\new_[7741]_  | ~\new_[6788]_ ) & (~\new_[5332]_  | ~\new_[6780]_ );
  assign \new_[5031]_  = (~\new_[7805]_  | ~\new_[6788]_ ) & (~\new_[5331]_  | ~\new_[6780]_ );
  assign \new_[5032]_  = (~\new_[7718]_  | ~\new_[6788]_ ) & (~\new_[5334]_  | ~\new_[6914]_ );
  assign \new_[5033]_  = (~\new_[7797]_  | ~\new_[6788]_ ) & (~\new_[5333]_  | ~\new_[6914]_ );
  assign \new_[5034]_  = (~\new_[7708]_  | ~\new_[6788]_ ) & (~\new_[5335]_  | ~\new_[6637]_ );
  assign \new_[5035]_  = (~\new_[7763]_  | ~\new_[6788]_ ) & (~\new_[5347]_  | ~\new_[6780]_ );
  assign \new_[5036]_  = (~\new_[7716]_  | ~\new_[6788]_ ) & (~\new_[5336]_  | ~\new_[6780]_ );
  assign \new_[5037]_  = (~\new_[7713]_  | ~\new_[6788]_ ) & (~\new_[5357]_  | ~\new_[6780]_ );
  assign \new_[5038]_  = (~\new_[7693]_  | ~\new_[6788]_ ) & (~\new_[5317]_  | ~\new_[6780]_ );
  assign \new_[5039]_  = (~\new_[7687]_  | ~\new_[6788]_ ) & (~\new_[5328]_  | ~\new_[6637]_ );
  assign \new_[5040]_  = (~\new_[7785]_  | ~\new_[6788]_ ) & (~\new_[5320]_  | ~\new_[6780]_ );
  assign \new_[5041]_  = (~\new_[7791]_  | ~\new_[6788]_ ) & (~\new_[5339]_  | ~\new_[6637]_ );
  assign \new_[5042]_  = (~\new_[7740]_  | ~\new_[6788]_ ) & (~\new_[5341]_  | ~\new_[6914]_ );
  assign \new_[5043]_  = (~\new_[7792]_  | ~\new_[6788]_ ) & (~\new_[5321]_  | ~\new_[6780]_ );
  assign \new_[5044]_  = (~\new_[7725]_  | ~\new_[6788]_ ) & (~\new_[5342]_  | ~\new_[6638]_ );
  assign \new_[5045]_  = (~\new_[7638]_  | ~\new_[6788]_ ) & (~\new_[5343]_  | ~\new_[6638]_ );
  assign \new_[5046]_  = (~\new_[7711]_  | ~\new_[6788]_ ) & (~\new_[5338]_  | ~\new_[6780]_ );
  assign \new_[5047]_  = (~\new_[7735]_  | ~\new_[6788]_ ) & (~\new_[5344]_  | ~\new_[6780]_ );
  assign \new_[5048]_  = (~\new_[7799]_  | ~\new_[6788]_ ) & (~\new_[5345]_  | ~\new_[6780]_ );
  assign \new_[5049]_  = (~\new_[7802]_  | ~\new_[6788]_ ) & (~\new_[5346]_  | ~\new_[6780]_ );
  assign \new_[5050]_  = (~\new_[7788]_  | ~\new_[6788]_ ) & (~\new_[5348]_  | ~\new_[6780]_ );
  assign \new_[5051]_  = (~\new_[7720]_  | ~\new_[6788]_ ) & (~\new_[5349]_  | ~\new_[6780]_ );
  assign \new_[5052]_  = (~\new_[7800]_  | ~\new_[6788]_ ) & (~\new_[5350]_  | ~\new_[6914]_ );
  assign \new_[5053]_  = (~\new_[7709]_  | ~\new_[6788]_ ) & (~\new_[5351]_  | ~\new_[6637]_ );
  assign \new_[5054]_  = (~\new_[7698]_  | ~\new_[6788]_ ) & (~\new_[5352]_  | ~\new_[6780]_ );
  assign \new_[5055]_  = (~\new_[7678]_  | ~\new_[6788]_ ) & (~\new_[5356]_  | ~\new_[6637]_ );
  assign \new_[5056]_  = (~\new_[7742]_  | ~\new_[6788]_ ) & (~\new_[5353]_  | ~\new_[6780]_ );
  assign \new_[5057]_  = (~\new_[7674]_  | ~\new_[6788]_ ) & (~\new_[5354]_  | ~\new_[6637]_ );
  assign \new_[5058]_  = (~\new_[7754]_  | ~\new_[6788]_ ) & (~\new_[5355]_  | ~\new_[6780]_ );
  assign \new_[5059]_  = (~\new_[7755]_  | ~\new_[6788]_ ) & (~\new_[5358]_  | ~\new_[6780]_ );
  assign \new_[5060]_  = (~\new_[7743]_  | ~\new_[6788]_ ) & (~\new_[5359]_  | ~\new_[6780]_ );
  assign \new_[5061]_  = (~\new_[7722]_  | ~\new_[6788]_ ) & (~\new_[5360]_  | ~\new_[6780]_ );
  assign \new_[5062]_  = (~\new_[7728]_  | ~\new_[6788]_ ) & (~\new_[5361]_  | ~\new_[6780]_ );
  assign \new_[5063]_  = (~\new_[7757]_  | ~\new_[6788]_ ) & (~\new_[5362]_  | ~\new_[6780]_ );
  assign \new_[5064]_  = (~\new_[7710]_  | ~\new_[6788]_ ) & (~\new_[5363]_  | ~\new_[6637]_ );
  assign \new_[5065]_  = (~\new_[7780]_  | ~\new_[6788]_ ) & (~\new_[5364]_  | ~\new_[6780]_ );
  assign \new_[5066]_  = (~\new_[7779]_  | ~\new_[6788]_ ) & (~\new_[5365]_  | ~\new_[6637]_ );
  assign \new_[5067]_  = (~\new_[7680]_  | ~\new_[6788]_ ) & (~\new_[5366]_  | ~\new_[6914]_ );
  assign \new_[5068]_  = (~\new_[7691]_  | ~\new_[6788]_ ) & (~\new_[5367]_  | ~\new_[6780]_ );
  assign \new_[5069]_  = \key_i[2]  & \new_[5253]_ ;
  assign \new_[5070]_  = ~\new_[5253]_  & (~\new_[6818]_  | ~\new_[6698]_ );
  assign \new_[5071]_  = \new_[7642]_  | \new_[8965]_ ;
  assign \new_[5072]_  = \new_[8146]_  | \new_[8727]_ ;
  assign \new_[5073]_  = \key_i[11]  & \new_[5253]_ ;
  assign \new_[5074]_  = \key_i[12]  & \new_[8307]_ ;
  assign \new_[5075]_  = \new_[7594]_  | \new_[8880]_ ;
  assign \new_[5076]_  = \new_[8159]_  | \new_[8727]_ ;
  assign \new_[5077]_  = \key_i[1]  & \new_[8307]_ ;
  assign \new_[5078]_  = ~\new_[5253]_  & (~\new_[6816]_  | ~\new_[6707]_ );
  assign \new_[5079]_  = ~\new_[6745]_  | ~\new_[5254]_ ;
  assign \new_[5080]_  = ~\new_[6919]_  | ~\new_[5255]_ ;
  assign \new_[5081]_  = ~\new_[6919]_  | ~\new_[5256]_ ;
  assign \new_[5082]_  = ~\new_[6745]_  | ~\new_[5257]_ ;
  assign \new_[5083]_  = ~\new_[6745]_  | ~\new_[5258]_ ;
  assign \new_[5084]_  = ~\new_[6919]_  | ~\new_[5259]_ ;
  assign \new_[5085]_  = ~\new_[6919]_  | ~\new_[5260]_ ;
  assign \new_[5086]_  = ~\new_[6919]_  | ~\new_[5261]_ ;
  assign \new_[5087]_  = ~\new_[6919]_  | ~\new_[5288]_ ;
  assign \new_[5088]_  = ~\new_[6919]_  | ~\new_[5284]_ ;
  assign \new_[5089]_  = ~\new_[6919]_  | ~\new_[5262]_ ;
  assign \new_[5090]_  = ~\new_[6919]_  | ~\new_[5263]_ ;
  assign \new_[5091]_  = ~\new_[6745]_  | ~\new_[5264]_ ;
  assign \new_[5092]_  = ~\new_[6919]_  | ~\new_[5265]_ ;
  assign \new_[5093]_  = ~\new_[6919]_  | ~\new_[5266]_ ;
  assign \new_[5094]_  = ~\new_[6745]_  | ~\new_[5267]_ ;
  assign \new_[5095]_  = ~\new_[6642]_  | ~\new_[5268]_ ;
  assign \new_[5096]_  = ~\new_[6745]_  | ~\new_[5269]_ ;
  assign \new_[5097]_  = ~\new_[6745]_  | ~\new_[5273]_ ;
  assign \new_[5098]_  = ~\new_[6919]_  | ~\new_[5270]_ ;
  assign \new_[5099]_  = ~\new_[6745]_  | ~\new_[5271]_ ;
  assign \new_[5100]_  = ~\new_[6642]_  | ~\new_[5272]_ ;
  assign \new_[5101]_  = ~\new_[6745]_  | ~\new_[5274]_ ;
  assign \new_[5102]_  = ~\new_[6919]_  | ~\new_[5275]_ ;
  assign \new_[5103]_  = ~\new_[6919]_  | ~\new_[5276]_ ;
  assign \new_[5104]_  = ~\new_[6919]_  | ~\new_[5277]_ ;
  assign \new_[5105]_  = ~\new_[6919]_  | ~\new_[5278]_ ;
  assign \new_[5106]_  = ~\new_[6919]_  | ~\new_[5280]_ ;
  assign \new_[5107]_  = ~\new_[6745]_  | ~\new_[5279]_ ;
  assign \new_[5108]_  = ~\new_[6642]_  | ~\new_[5281]_ ;
  assign \new_[5109]_  = ~\new_[6642]_  | ~\new_[5282]_ ;
  assign \new_[5110]_  = ~\new_[6745]_  | ~\new_[5283]_ ;
  assign \new_[5111]_  = ~\new_[6745]_  | ~\new_[5285]_ ;
  assign \new_[5112]_  = ~\new_[6745]_  | ~\new_[5286]_ ;
  assign \new_[5113]_  = ~\new_[6745]_  | ~\new_[5287]_ ;
  assign \new_[5114]_  = ~\new_[5253]_ ;
  assign \new_[5115]_  = ~\new_[8307]_ ;
  assign \new_[5116]_  = \new_[8683]_  ^ \new_[8496]_ ;
  assign \new_[5117]_  = \new_[5484]_  ^ \new_[5369]_ ;
  assign \new_[5118]_  = \new_[5610]_  ^ \new_[5370]_ ;
  assign \new_[5119]_  = \new_[8682]_  ^ \new_[8527]_ ;
  assign \new_[5120]_  = \new_[8618]_  ^ \new_[5371]_ ;
  assign \new_[5121]_  = \new_[5611]_  ^ \new_[5372]_ ;
  assign \new_[5122]_  = \new_[8622]_  ^ \new_[8496]_ ;
  assign \new_[5123]_  = \new_[5485]_  ^ \new_[5373]_ ;
  assign \new_[5124]_  = \new_[5610]_  ^ \new_[5374]_ ;
  assign \new_[5125]_  = \new_[8619]_  ^ \new_[8527]_ ;
  assign \new_[5126]_  = \new_[8681]_  ^ \new_[5375]_ ;
  assign \new_[5127]_  = \new_[5611]_  ^ \new_[5376]_ ;
  assign \new_[5128]_  = \new_[5309]_  ^ \new_[5469]_ ;
  assign \new_[5129]_  = \new_[5295]_  ^ \new_[8736]_ ;
  assign \new_[5130]_  = \new_[8622]_  ^ \new_[8736]_ ;
  assign \new_[5131]_  = \new_[5311]_  ^ \new_[5476]_ ;
  assign \new_[5132]_  = \new_[5298]_  ^ \new_[8441]_ ;
  assign \new_[5133]_  = \new_[8619]_  ^ \new_[8441]_ ;
  assign \new_[5134]_  = \new_[8797]_  ^ \new_[5299]_ ;
  assign \new_[5135]_  = \new_[5301]_  ^ \new_[8758]_ ;
  assign \new_[5136]_  = \new_[8683]_  ^ \new_[8758]_ ;
  assign \new_[5137]_  = \new_[8857]_  ^ \new_[5302]_ ;
  assign \new_[5138]_  = \new_[5304]_  ^ \new_[8790]_ ;
  assign \new_[5139]_  = \new_[8682]_  ^ \new_[8790]_ ;
  assign \new_[5140]_  = \new_[8444]_  ^ \new_[5305]_ ;
  assign \new_[5141]_  = \new_[8762]_  ^ \new_[5296]_ ;
  assign \new_[5142]_  = ~\new_[5248]_ ;
  assign \new_[5143]_  = ~\new_[8401]_  | ~\new_[8805]_ ;
  assign \new_[5144]_  = ~\new_[6642]_  | ~\new_[5312]_ ;
  assign \new_[5145]_  = ~\new_[6745]_  | ~\new_[5313]_ ;
  assign \new_[5146]_  = ~\new_[6919]_  | ~\new_[5314]_ ;
  assign \new_[5147]_  = ~\new_[6919]_  | ~\new_[5315]_ ;
  assign \new_[5148]_  = ~\new_[6919]_  | ~\new_[5316]_ ;
  assign \new_[5149]_  = ~\new_[6919]_  | ~\new_[5318]_ ;
  assign \new_[5150]_  = ~\new_[6919]_  | ~\new_[5322]_ ;
  assign \new_[5151]_  = ~\new_[6919]_  | ~\new_[5323]_ ;
  assign \new_[5152]_  = ~\new_[6919]_  | ~\new_[5324]_ ;
  assign \new_[5153]_  = ~\new_[6919]_  | ~\new_[5325]_ ;
  assign \new_[5154]_  = ~\new_[6745]_  | ~\new_[5326]_ ;
  assign \new_[5155]_  = ~\new_[6642]_  | ~\new_[5317]_ ;
  assign \new_[5156]_  = ~\new_[6745]_  | ~\new_[5319]_ ;
  assign \new_[5157]_  = ~\new_[6919]_  | ~\new_[5327]_ ;
  assign \new_[5158]_  = ~\new_[6642]_  | ~\new_[5329]_ ;
  assign \new_[5159]_  = ~\new_[6919]_  | ~\new_[5337]_ ;
  assign \new_[5160]_  = ~\new_[6919]_  | ~\new_[5330]_ ;
  assign \new_[5161]_  = ~\new_[6919]_  | ~\new_[5331]_ ;
  assign \new_[5162]_  = ~\new_[6642]_  | ~\new_[5332]_ ;
  assign \new_[5163]_  = ~\new_[6919]_  | ~\new_[5333]_ ;
  assign \new_[5164]_  = ~\new_[6919]_  | ~\new_[5334]_ ;
  assign \new_[5165]_  = ~\new_[6642]_  | ~\new_[5335]_ ;
  assign \new_[5166]_  = ~\new_[6642]_  | ~\new_[5347]_ ;
  assign \new_[5167]_  = ~\new_[6642]_  | ~\new_[5336]_ ;
  assign \new_[5168]_  = ~\new_[6919]_  | ~\new_[5320]_ ;
  assign \new_[5169]_  = ~\new_[6919]_  | ~\new_[5357]_ ;
  assign \new_[5170]_  = ~\new_[6919]_  | ~\new_[5328]_ ;
  assign \new_[5171]_  = ~\new_[6642]_  | ~\new_[5339]_ ;
  assign \new_[5172]_  = ~\new_[6919]_  | ~\new_[5340]_ ;
  assign \new_[5173]_  = ~\new_[6642]_  | ~\new_[5321]_ ;
  assign \new_[5174]_  = ~\new_[6919]_  | ~\new_[5341]_ ;
  assign \new_[5175]_  = ~\new_[6919]_  | ~\new_[5343]_ ;
  assign \new_[5176]_  = ~\new_[6919]_  | ~\new_[5344]_ ;
  assign \new_[5177]_  = ~\new_[6642]_  | ~\new_[5345]_ ;
  assign \new_[5178]_  = ~\new_[6642]_  | ~\new_[5346]_ ;
  assign \new_[5179]_  = ~\new_[6642]_  | ~\new_[5348]_ ;
  assign \new_[5180]_  = ~\new_[6642]_  | ~\new_[5349]_ ;
  assign \new_[5181]_  = ~\new_[6919]_  | ~\new_[5350]_ ;
  assign \new_[5182]_  = ~\new_[6919]_  | ~\new_[5351]_ ;
  assign \new_[5183]_  = ~\new_[6642]_  | ~\new_[5352]_ ;
  assign \new_[5184]_  = ~\new_[6919]_  | ~\new_[5353]_ ;
  assign \new_[5185]_  = ~\new_[6919]_  | ~\new_[5342]_ ;
  assign \new_[5186]_  = ~\new_[6919]_  | ~\new_[5354]_ ;
  assign \new_[5187]_  = ~\new_[6919]_  | ~\new_[5355]_ ;
  assign \new_[5188]_  = ~\new_[6919]_  | ~\new_[5356]_ ;
  assign \new_[5189]_  = ~\new_[6642]_  | ~\new_[5338]_ ;
  assign \new_[5190]_  = ~\new_[6919]_  | ~\new_[5358]_ ;
  assign \new_[5191]_  = ~\new_[6642]_  | ~\new_[5359]_ ;
  assign \new_[5192]_  = ~\new_[6642]_  | ~\new_[5360]_ ;
  assign \new_[5193]_  = ~\new_[6745]_  | ~\new_[5361]_ ;
  assign \new_[5194]_  = ~\new_[6642]_  | ~\new_[5362]_ ;
  assign \new_[5195]_  = ~\new_[6642]_  | ~\new_[5363]_ ;
  assign \new_[5196]_  = ~\new_[6642]_  | ~\new_[5364]_ ;
  assign \new_[5197]_  = ~\new_[6642]_  | ~\new_[5365]_ ;
  assign \new_[5198]_  = ~\new_[6642]_  | ~\new_[5366]_ ;
  assign \new_[5199]_  = ~\new_[6642]_  | ~\new_[5367]_ ;
  assign \new_[5200]_  = ~\new_[6919]_  | ~\new_[5368]_ ;
  assign \new_[5201]_  = ~\new_[8308]_ ;
  assign \new_[5202]_  = ~\new_[5253]_ ;
  assign \new_[5203]_  = ~\new_[8727]_ ;
  assign \new_[5204]_  = \new_[6632]_  ? \new_[7624]_  : \new_[5383]_ ;
  assign \new_[5205]_  = \new_[3106]_  ? \new_[7607]_  : \new_[5410]_ ;
  assign \new_[5206]_  = \new_[6581]_  ? \new_[7607]_  : \new_[5409]_ ;
  assign \new_[5207]_  = \new_[6450]_  ? \new_[7607]_  : \new_[5387]_ ;
  assign \new_[5208]_  = \new_[6451]_  ? \new_[7624]_  : \new_[5389]_ ;
  assign \new_[5209]_  = \new_[6748]_  ? \new_[7770]_  : \new_[5386]_ ;
  assign \new_[5210]_  = \new_[3514]_  ? \new_[7770]_  : \new_[5385]_ ;
  assign \new_[5211]_  = \new_[3107]_  ? \new_[7770]_  : \new_[5388]_ ;
  assign \new_[5212]_  = \new_[3377]_  ? \new_[7770]_  : \new_[5390]_ ;
  assign \new_[5213]_  = \new_[6420]_  ? \new_[7607]_  : \new_[5391]_ ;
  assign \new_[5214]_  = \new_[6449]_  ? \new_[7770]_  : \new_[5392]_ ;
  assign \new_[5215]_  = \new_[6452]_  ? \new_[7624]_  : \new_[5393]_ ;
  assign \new_[5216]_  = \new_[2870]_  ? \new_[7624]_  : \new_[5394]_ ;
  assign \new_[5217]_  = \new_[6597]_  ? \new_[7624]_  : \new_[5404]_ ;
  assign \new_[5218]_  = \new_[6599]_  ? \new_[7624]_  : \new_[5397]_ ;
  assign \new_[5219]_  = \new_[6656]_  ? \new_[7624]_  : \new_[5396]_ ;
  assign \new_[5220]_  = \new_[6624]_  ? \new_[7624]_  : \new_[5398]_ ;
  assign \new_[5221]_  = \new_[6620]_  ? \new_[7624]_  : \new_[5400]_ ;
  assign \new_[5222]_  = \new_[6580]_  ? \new_[7770]_  : \new_[5399]_ ;
  assign \new_[5223]_  = \new_[3406]_  ? \new_[7770]_  : \new_[5384]_ ;
  assign \new_[5224]_  = \new_[6575]_  ? \new_[7770]_  : \new_[5406]_ ;
  assign \new_[5225]_  = \new_[3410]_  ? \new_[7770]_  : \new_[5395]_ ;
  assign \new_[5226]_  = \new_[6590]_  ? \new_[7624]_  : \new_[5403]_ ;
  assign \new_[5227]_  = \new_[6421]_  ? \new_[7624]_  : \new_[5405]_ ;
  assign \new_[5228]_  = \new_[6571]_  ? \new_[7624]_  : \new_[5401]_ ;
  assign \new_[5229]_  = \new_[6723]_  ? \new_[7624]_  : \new_[5407]_ ;
  assign \new_[5230]_  = \new_[3382]_  ? \new_[7624]_  : \new_[5408]_ ;
  assign \new_[5231]_  = \new_[3257]_  ? \new_[7770]_  : \new_[5411]_ ;
  assign \new_[5232]_  = \new_[6443]_  ? \new_[7624]_  : \new_[5412]_ ;
  assign \new_[5233]_  = \new_[6422]_  ? \new_[7624]_  : \new_[5413]_ ;
  assign \new_[5234]_  = \new_[6601]_  ? \new_[7624]_  : \new_[5414]_ ;
  assign \new_[5235]_  = \new_[6623]_  ? \new_[7607]_  : \new_[5402]_ ;
  assign \new_[5236]_  = \new_[6610]_  ? \new_[7624]_  : \new_[5415]_ ;
  assign \new_[5237]_  = \new_[3515]_  ? \new_[7607]_  : \new_[5416]_ ;
  assign \new_[5238]_  = \new_[6702]_  ? \new_[7607]_  : \new_[5417]_ ;
  assign \new_[5239]_  = \new_[6641]_  ? \new_[7607]_  : \new_[5382]_ ;
  assign \new_[5240]_  = \new_[5843]_  ^ \new_[5418]_ ;
  assign \new_[5241]_  = \new_[5426]_  ^ \new_[5378]_ ;
  assign \new_[5242]_  = \new_[8510]_  ^ \new_[5427]_ ;
  assign \new_[5243]_  = \new_[5427]_  ^ \new_[5428]_ ;
  assign \new_[5244]_  = \new_[8485]_  ^ \new_[8503]_ ;
  assign \new_[5245]_  = \new_[8503]_  ^ \new_[8484]_ ;
  assign \new_[5246]_  = \new_[8772]_  ^ \new_[5428]_ ;
  assign \new_[5247]_  = \new_[8504]_  ^ \new_[8484]_ ;
  assign \new_[5248]_  = (~\new_[5483]_  & ~\new_[5795]_ ) | (~\new_[5425]_  & ~\new_[5848]_ );
  assign \new_[5249]_  = ~\new_[8805]_  | ~\new_[8988]_ ;
  assign \new_[5250]_  = \new_[8754]_  ^ \new_[8637]_ ;
  assign \new_[5251]_  = \new_[8602]_  ^ \new_[8754]_ ;
  assign \new_[5252]_  = \new_[8602]_  ^ \new_[8753]_ ;
  assign \new_[5253]_  = ~\new_[8310]_ ;
  assign \new_[5254]_  = \new_[6631]_  ? \new_[7624]_  : \new_[5433]_ ;
  assign \new_[5255]_  = \new_[6594]_  ? \new_[7624]_  : \new_[5434]_ ;
  assign \new_[5256]_  = \new_[3105]_  ? \new_[7624]_  : \new_[5435]_ ;
  assign \new_[5257]_  = \new_[6432]_  ? \new_[7624]_  : \new_[5436]_ ;
  assign \new_[5258]_  = \new_[6716]_  ? \new_[7770]_  : \new_[5437]_ ;
  assign \new_[5259]_  = \new_[3443]_  ? \new_[7770]_  : \new_[5442]_ ;
  assign \new_[5260]_  = \new_[6573]_  ? \new_[7624]_  : \new_[5438]_ ;
  assign \new_[5261]_  = \new_[6630]_  ? \new_[7624]_  : \new_[5439]_ ;
  assign \new_[5262]_  = \new_[2757]_  ? \new_[7624]_  : \new_[5440]_ ;
  assign \new_[5263]_  = \new_[3109]_  ? \new_[7624]_  : \new_[5444]_ ;
  assign \new_[5264]_  = \new_[3386]_  ? \new_[7624]_  : \new_[5445]_ ;
  assign \new_[5265]_  = \new_[3863]_  ? \new_[7770]_  : \new_[5443]_ ;
  assign \new_[5266]_  = \new_[6416]_  ? \new_[7624]_  : \new_[5446]_ ;
  assign \new_[5267]_  = \new_[6572]_  ? \new_[7770]_  : \new_[5447]_ ;
  assign \new_[5268]_  = \new_[6438]_  ? \new_[7624]_  : \new_[5448]_ ;
  assign \new_[5269]_  = \new_[6666]_  ? \new_[7624]_  : \new_[5449]_ ;
  assign \new_[5270]_  = \new_[6448]_  ? \new_[7624]_  : \new_[5450]_ ;
  assign \new_[5271]_  = \new_[2934]_  ? \new_[7624]_  : \new_[5451]_ ;
  assign \new_[5272]_  = \new_[6643]_  ? \new_[7770]_  : \new_[5452]_ ;
  assign \new_[5273]_  = \new_[6625]_  ? \new_[7624]_  : \new_[5453]_ ;
  assign \new_[5274]_  = \new_[6746]_  ? \new_[7607]_  : \new_[5454]_ ;
  assign \new_[5275]_  = \new_[6639]_  ? \new_[7624]_  : \new_[5455]_ ;
  assign \new_[5276]_  = \new_[3108]_  ? \new_[7607]_  : \new_[5458]_ ;
  assign \new_[5277]_  = \new_[6663]_  ? \new_[7624]_  : \new_[5456]_ ;
  assign \new_[5278]_  = \new_[6640]_  ? \new_[7624]_  : \new_[5457]_ ;
  assign \new_[5279]_  = \new_[6424]_  ? \new_[7770]_  : \new_[5460]_ ;
  assign \new_[5280]_  = \new_[6628]_  ? \new_[7770]_  : \new_[5459]_ ;
  assign \new_[5281]_  = \new_[2758]_  ? \new_[7770]_  : \new_[5461]_ ;
  assign \new_[5282]_  = \new_[6587]_  ? \new_[7624]_  : \new_[5462]_ ;
  assign \new_[5283]_  = \new_[2755]_  ? \new_[7624]_  : \new_[5463]_ ;
  assign \new_[5284]_  = \new_[3846]_  ? \new_[7770]_  : \new_[5464]_ ;
  assign \new_[5285]_  = \new_[3409]_  ? \new_[7624]_  : \new_[5465]_ ;
  assign \new_[5286]_  = \new_[3885]_  ? \new_[7770]_  : \new_[5466]_ ;
  assign \new_[5287]_  = \new_[6574]_  ? \new_[7770]_  : \new_[5467]_ ;
  assign \new_[5288]_  = \new_[2932]_  ? \new_[7624]_  : \new_[5441]_ ;
  assign \new_[5289]_  = \new_[5421]_  ^ \new_[5428]_ ;
  assign \new_[5290]_  = \new_[5420]_  ^ \new_[8484]_ ;
  assign \new_[5291]_  = \new_[5422]_  ^ \new_[5427]_ ;
  assign \new_[5292]_  = \new_[5423]_  ^ \new_[8503]_ ;
  assign \new_[5293]_  = \\round_reg[1] ;
  assign \new_[5294]_  = \new_[8795]_  ^ \new_[8759]_ ;
  assign \new_[5295]_  = \new_[8619]_  ^ \new_[5484]_ ;
  assign \new_[5296]_  = \new_[5485]_  ^ \new_[8857]_ ;
  assign \new_[5297]_  = \new_[8833]_  ^ \new_[8793]_ ;
  assign \new_[5298]_  = \new_[8683]_  ^ \new_[8618]_ ;
  assign \new_[5299]_  = \new_[8681]_  ^ \new_[8442]_ ;
  assign \new_[5300]_  = \new_[8832]_  ^ \new_[8738]_ ;
  assign \new_[5301]_  = \new_[8682]_  ^ \new_[5485]_ ;
  assign \new_[5302]_  = \new_[5484]_  ^ \new_[8762]_ ;
  assign \new_[5303]_  = \new_[8794]_  ^ \new_[8831]_ ;
  assign \new_[5304]_  = \new_[8622]_  ^ \new_[8681]_ ;
  assign \new_[5305]_  = \new_[8618]_  ^ \new_[8791]_ ;
  assign \new_[5306]_  = \new_[5554]_  ^ \new_[5481]_ ;
  assign \new_[5307]_  = \\round_reg[2] ;
  assign \new_[5308]_  = \new_[8740]_  ^ \new_[8692]_ ;
  assign \new_[5309]_  = \new_[8741]_  ^ \new_[8692]_ ;
  assign \new_[5310]_  = \new_[8693]_  ^ \new_[8741]_ ;
  assign \new_[5311]_  = \new_[8693]_  ^ \new_[8740]_ ;
  assign \new_[5312]_  = \new_[3104]_  ? \new_[7770]_  : \new_[5538]_ ;
  assign \new_[5313]_  = \new_[2935]_  ? \new_[7624]_  : \new_[5492]_ ;
  assign \new_[5314]_  = \new_[6495]_  ? \new_[7624]_  : \new_[5493]_ ;
  assign \new_[5315]_  = \new_[6423]_  ? \new_[7770]_  : \new_[5494]_ ;
  assign \new_[5316]_  = \new_[6445]_  ? \new_[7770]_  : \new_[5495]_ ;
  assign \new_[5317]_  = \new_[6600]_  ? \new_[7624]_  : \new_[5491]_ ;
  assign \new_[5318]_  = \new_[6618]_  ? \new_[7624]_  : \new_[5496]_ ;
  assign \new_[5319]_  = \new_[3383]_  ? \new_[7770]_  : \new_[5502]_ ;
  assign \new_[5320]_  = \new_[6586]_  ? \new_[7770]_  : \new_[5533]_ ;
  assign \new_[5321]_  = \new_[6607]_  ? \new_[7624]_  : \new_[5516]_ ;
  assign \new_[5322]_  = \new_[2756]_  ? \new_[7770]_  : \new_[5497]_ ;
  assign \new_[5323]_  = \new_[6425]_  ? \new_[7770]_  : \new_[5498]_ ;
  assign \new_[5324]_  = \new_[6606]_  ? \new_[7770]_  : \new_[5500]_ ;
  assign \new_[5325]_  = \new_[6605]_  ? \new_[7770]_  : \new_[5499]_ ;
  assign \new_[5326]_  = \new_[6652]_  ? \new_[7624]_  : \new_[5501]_ ;
  assign \new_[5327]_  = \new_[6442]_  ? \new_[7624]_  : \new_[5503]_ ;
  assign \new_[5328]_  = \new_[6694]_  ? \new_[7624]_  : \new_[5515]_ ;
  assign \new_[5329]_  = \new_[3385]_  ? \new_[7770]_  : \new_[5504]_ ;
  assign \new_[5330]_  = \new_[6446]_  ? \new_[7624]_  : \new_[5505]_ ;
  assign \new_[5331]_  = \new_[6704]_  ? \new_[7624]_  : \new_[5507]_ ;
  assign \new_[5332]_  = \new_[3857]_  ? \new_[7624]_  : \new_[5506]_ ;
  assign \new_[5333]_  = \new_[6419]_  ? \new_[7624]_  : \new_[5508]_ ;
  assign \new_[5334]_  = \new_[6596]_  ? \new_[7624]_  : \new_[5509]_ ;
  assign \new_[5335]_  = \new_[6547]_  ? \new_[7624]_  : \new_[5545]_ ;
  assign \new_[5336]_  = \new_[6619]_  ? \new_[7770]_  : \new_[5511]_ ;
  assign \new_[5337]_  = \new_[6426]_  ? \new_[7770]_  : \new_[5512]_ ;
  assign \new_[5338]_  = \new_[6585]_  ? \new_[7624]_  : \new_[5531]_ ;
  assign \new_[5339]_  = \new_[6427]_  ? \new_[7624]_  : \new_[5513]_ ;
  assign \new_[5340]_  = \new_[6566]_  ? \new_[7624]_  : \new_[5514]_ ;
  assign \new_[5341]_  = \new_[6614]_  ? \new_[7770]_  : \new_[5542]_ ;
  assign \new_[5342]_  = \new_[6568]_  ? \new_[7624]_  : \new_[5524]_ ;
  assign \new_[5343]_  = \new_[6569]_  ? \new_[7624]_  : \new_[5517]_ ;
  assign \new_[5344]_  = \new_[6589]_  ? \new_[7624]_  : \new_[5519]_ ;
  assign \new_[5345]_  = \new_[6629]_  ? \new_[7770]_  : \new_[5520]_ ;
  assign \new_[5346]_  = \new_[6444]_  ? \new_[7624]_  : \new_[5521]_ ;
  assign \new_[5347]_  = \new_[6598]_  ? \new_[7770]_  : \new_[5510]_ ;
  assign \new_[5348]_  = \new_[6749]_  ? \new_[7770]_  : \new_[5522]_ ;
  assign \new_[5349]_  = \new_[6595]_  ? \new_[7770]_  : \new_[5523]_ ;
  assign \new_[5350]_  = \new_[6579]_  ? \new_[7770]_  : \new_[5527]_ ;
  assign \new_[5351]_  = \new_[6591]_  ? \new_[7624]_  : \new_[5525]_ ;
  assign \new_[5352]_  = \new_[6428]_  ? \new_[7770]_  : \new_[5526]_ ;
  assign \new_[5353]_  = \new_[6584]_  ? \new_[7624]_  : \new_[5528]_ ;
  assign \new_[5354]_  = \new_[6714]_  ? \new_[7624]_  : \new_[5529]_ ;
  assign \new_[5355]_  = \new_[6592]_  ? \new_[7770]_  : \new_[5530]_ ;
  assign \new_[5356]_  = \new_[6430]_  ? \new_[7770]_  : \new_[5518]_ ;
  assign \new_[5357]_  = \new_[6429]_  ? \new_[7770]_  : \new_[5532]_ ;
  assign \new_[5358]_  = \new_[6433]_  ? \new_[7770]_  : \new_[5534]_ ;
  assign \new_[5359]_  = \new_[6546]_  ? \new_[7624]_  : \new_[5535]_ ;
  assign \new_[5360]_  = \new_[6627]_  ? \new_[7624]_  : \new_[5536]_ ;
  assign \new_[5361]_  = \new_[6616]_  ? \new_[7607]_  : \new_[5537]_ ;
  assign \new_[5362]_  = \new_[6609]_  ? \new_[7770]_  : \new_[5539]_ ;
  assign \new_[5363]_  = \new_[6588]_  ? \new_[7624]_  : \new_[5540]_ ;
  assign \new_[5364]_  = \new_[6626]_  ? \new_[7624]_  : \new_[5541]_ ;
  assign \new_[5365]_  = \new_[6593]_  ? \new_[7770]_  : \new_[5543]_ ;
  assign \new_[5366]_  = \new_[3387]_  ? \new_[7624]_  : \new_[5544]_ ;
  assign \new_[5367]_  = \new_[3103]_  ? \new_[7770]_  : \new_[5546]_ ;
  assign \new_[5368]_  = \new_[6751]_  ? \new_[7770]_  : \new_[5547]_ ;
  assign \new_[5369]_  = \new_[8864]_  ^ \new_[5470]_ ;
  assign \new_[5370]_  = \new_[5660]_  ^ \new_[5471]_ ;
  assign \new_[5371]_  = \new_[5608]_  ^ \new_[5479]_ ;
  assign \new_[5372]_  = \new_[5662]_  ^ \new_[5473]_ ;
  assign \new_[5373]_  = \new_[8870]_  ^ \new_[5477]_ ;
  assign \new_[5374]_  = \new_[5665]_  ^ \new_[5474]_ ;
  assign \new_[5375]_  = \new_[5609]_  ^ \new_[5478]_ ;
  assign \new_[5376]_  = \new_[5663]_  ^ \new_[5475]_ ;
  assign \new_[5377]_  = \\round_reg[0] ;
  assign \new_[5378]_  = ~\new_[8808]_  | ~\new_[1227]_ ;
  assign \new_[5379]_  = \new_[5851]_  ^ \new_[5556]_ ;
  assign \new_[5380]_  = ~\new_[8457]_ ;
  assign \new_[5381]_  = ~\new_[8808]_  | ~\new_[1388]_ ;
  assign \new_[5382]_  = ~\new_[7200]_  | (~\new_[5595]_  & ~\new_[7602]_ );
  assign \new_[5383]_  = ~\new_[7300]_  | (~\new_[5561]_  & ~\new_[7584]_ );
  assign \new_[5384]_  = ~\new_[7210]_  | (~\new_[5569]_  & ~\new_[7602]_ );
  assign \new_[5385]_  = ~\new_[7292]_  | (~\new_[5571]_  & ~\new_[7602]_ );
  assign \new_[5386]_  = ~\new_[7366]_  | (~\new_[5568]_  & ~\new_[7599]_ );
  assign \new_[5387]_  = ~\new_[7208]_  | (~\new_[5565]_  & ~\new_[7602]_ );
  assign \new_[5388]_  = ~\new_[7303]_  | (~\new_[5566]_  & ~\new_[7602]_ );
  assign \new_[5389]_  = ~\new_[7353]_  | (~\new_[5567]_  & ~\new_[7602]_ );
  assign \new_[5390]_  = ~\new_[7397]_  | (~\new_[5564]_  & ~\new_[7599]_ );
  assign \new_[5391]_  = ~\new_[7237]_  | (~\new_[5586]_  & ~\new_[7602]_ );
  assign \new_[5392]_  = ~\new_[7161]_  | (~\new_[5572]_  & ~\new_[7602]_ );
  assign \new_[5393]_  = ~\new_[7282]_  | (~\new_[5573]_  & ~\new_[7602]_ );
  assign \new_[5394]_  = ~\new_[7160]_  | (~\new_[5574]_  & ~\new_[7602]_ );
  assign \new_[5395]_  = ~\new_[7315]_  | (~\new_[5570]_  & ~\new_[7602]_ );
  assign \new_[5396]_  = ~\new_[7224]_  | (~\new_[5577]_  & ~\new_[7602]_ );
  assign \new_[5397]_  = ~\new_[7241]_  | (~\new_[5575]_  & ~\new_[7602]_ );
  assign \new_[5398]_  = ~\new_[7387]_  | (~\new_[5581]_  & ~\new_[7599]_ );
  assign \new_[5399]_  = ~\new_[7229]_  | (~\new_[5583]_  & ~\new_[7599]_ );
  assign \new_[5400]_  = ~\new_[7156]_  | (~\new_[5578]_  & ~\new_[7599]_ );
  assign \new_[5401]_  = ~\new_[7320]_  | (~\new_[5582]_  & ~\new_[7602]_ );
  assign \new_[5402]_  = ~\new_[7312]_  | (~\new_[5584]_  & ~\new_[7602]_ );
  assign \new_[5403]_  = ~\new_[7310]_  | (~\new_[5579]_  & ~\new_[7602]_ );
  assign \new_[5404]_  = ~\new_[7403]_  | (~\new_[5580]_  & ~\new_[7599]_ );
  assign \new_[5405]_  = ~\new_[7219]_  | (~\new_[5576]_  & ~\new_[7599]_ );
  assign \new_[5406]_  = ~\new_[7332]_  | (~\new_[5585]_  & ~\new_[7599]_ );
  assign \new_[5407]_  = ~\new_[7386]_  | (~\new_[5588]_  & ~\new_[7599]_ );
  assign \new_[5408]_  = ~\new_[7202]_  | (~\new_[5587]_  & ~\new_[7599]_ );
  assign \new_[5409]_  = ~\new_[7230]_  | (~\new_[5563]_  & ~\new_[7599]_ );
  assign \new_[5410]_  = ~\new_[7313]_  | (~\new_[5562]_  & ~\new_[7599]_ );
  assign \new_[5411]_  = ~\new_[7174]_  | (~\new_[5589]_  & ~\new_[7599]_ );
  assign \new_[5412]_  = ~\new_[7232]_  | (~\new_[5591]_  & ~\new_[7599]_ );
  assign \new_[5413]_  = ~\new_[7227]_  | (~\new_[5590]_  & ~\new_[7602]_ );
  assign \new_[5414]_  = ~\new_[7357]_  | (~\new_[5592]_  & ~\new_[7602]_ );
  assign \new_[5415]_  = ~\new_[7305]_  | (~\new_[5593]_  & ~\new_[7599]_ );
  assign \new_[5416]_  = ~\new_[7190]_  | (~\new_[5594]_  & ~\new_[7584]_ );
  assign \new_[5417]_  = ~\new_[7329]_  | (~\new_[5596]_  & ~\new_[7602]_ );
  assign \new_[5418]_  = ~\new_[8808]_  | ~\new_[1709]_ ;
  assign \new_[5419]_  = \\round_reg[3] ;
  assign \new_[5420]_  = \new_[8869]_  ^ \new_[5609]_ ;
  assign \new_[5421]_  = \new_[8865]_  ^ \new_[8870]_ ;
  assign \new_[5422]_  = \new_[8875]_  ^ \new_[8864]_ ;
  assign \new_[5423]_  = \new_[8871]_  ^ \new_[5608]_ ;
  assign \new_[5424]_  = ~\new_[8414]_ ;
  assign \new_[5425]_  = ~\new_[5483]_ ;
  assign \new_[5426]_  = ~\new_[8592]_  | ~\new_[1709]_ ;
  assign \new_[5427]_  = \new_[8504]_  ^ \new_[8772]_ ;
  assign \new_[5428]_  = \new_[8485]_  ^ \new_[8510]_ ;
  assign \new_[5429]_  = \new_[8504]_  ^ \new_[8485]_ ;
  assign \new_[5430]_  = \new_[8772]_  ^ \new_[8510]_ ;
  assign n3555 = ~\new_[5560]_  | ~\new_[6829]_ ;
  assign n3560 = ~\new_[5559]_  | (~\new_[7565]_  & ~load_i);
  assign \new_[5433]_  = ~\new_[7330]_  | (~\new_[5622]_  & ~\new_[7584]_ );
  assign \new_[5434]_  = ~\new_[7168]_  | (~\new_[5624]_  & ~\new_[7602]_ );
  assign \new_[5435]_  = ~\new_[7306]_  | (~\new_[5623]_  & ~\new_[7602]_ );
  assign \new_[5436]_  = ~\new_[7377]_  | (~\new_[5629]_  & ~\new_[7599]_ );
  assign \new_[5437]_  = ~\new_[7209]_  | (~\new_[5630]_  & ~\new_[7599]_ );
  assign \new_[5438]_  = ~\new_[7319]_  | (~\new_[5632]_  & ~\new_[7599]_ );
  assign \new_[5439]_  = ~\new_[7385]_  | (~\new_[5634]_  & ~\new_[7599]_ );
  assign \new_[5440]_  = ~\new_[7234]_  | (~\new_[5637]_  & ~\new_[7584]_ );
  assign \new_[5441]_  = ~\new_[7287]_  | (~\new_[5628]_  & ~\new_[7602]_ );
  assign \new_[5442]_  = ~\new_[7391]_  | (~\new_[5631]_  & ~\new_[7602]_ );
  assign \new_[5443]_  = ~\new_[7267]_  | (~\new_[5642]_  & ~\new_[7602]_ );
  assign \new_[5444]_  = ~\new_[7297]_  | (~\new_[5633]_  & ~\new_[7602]_ );
  assign \new_[5445]_  = ~\new_[7356]_  | (~\new_[5625]_  & ~\new_[7599]_ );
  assign \new_[5446]_  = ~\new_[7395]_  | (~\new_[5651]_  & ~\new_[7584]_ );
  assign \new_[5447]_  = ~\new_[7350]_  | (~\new_[5635]_  & ~\new_[7599]_ );
  assign \new_[5448]_  = ~\new_[7192]_  | (~\new_[5640]_  & ~\new_[7599]_ );
  assign \new_[5449]_  = ~\new_[7383]_  | (~\new_[5653]_  & ~\new_[7599]_ );
  assign \new_[5450]_  = ~\new_[7347]_  | (~\new_[8235]_  & ~\new_[7584]_ );
  assign \new_[5451]_  = ~\new_[7341]_  | (~\new_[5636]_  & ~\new_[7599]_ );
  assign \new_[5452]_  = ~\new_[7263]_  | (~\new_[5638]_  & ~\new_[7592]_ );
  assign \new_[5453]_  = ~\new_[7182]_  | (~\new_[5639]_  & ~\new_[7602]_ );
  assign \new_[5454]_  = ~\new_[7348]_  | (~\new_[5641]_  & ~\new_[7602]_ );
  assign \new_[5455]_  = ~\new_[7187]_  | (~\new_[5643]_  & ~\new_[7602]_ );
  assign \new_[5456]_  = ~\new_[7339]_  | (~\new_[5645]_  & ~\new_[7602]_ );
  assign \new_[5457]_  = ~\new_[7349]_  | (~\new_[5627]_  & ~\new_[7602]_ );
  assign \new_[5458]_  = ~\new_[7167]_  | (~\new_[5644]_  & ~\new_[7584]_ );
  assign \new_[5459]_  = ~\new_[7373]_  | (~\new_[5646]_  & ~\new_[7602]_ );
  assign \new_[5460]_  = ~\new_[7378]_  | (~\new_[5647]_  & ~\new_[7599]_ );
  assign \new_[5461]_  = ~\new_[7351]_  | (~\new_[5649]_  & ~\new_[7599]_ );
  assign \new_[5462]_  = ~\new_[7323]_  | (~\new_[5648]_  & ~\new_[7599]_ );
  assign \new_[5463]_  = ~\new_[7193]_  | (~\new_[5650]_  & ~\new_[7599]_ );
  assign \new_[5464]_  = ~\new_[7400]_  | (~\new_[5626]_  & ~\new_[7599]_ );
  assign \new_[5465]_  = ~\new_[7151]_  | (~\new_[5652]_  & ~\new_[7599]_ );
  assign \new_[5466]_  = ~\new_[7392]_  | (~\new_[5654]_  & ~\new_[7599]_ );
  assign \new_[5467]_  = ~\new_[7390]_  | (~\new_[5655]_  & ~\new_[7584]_ );
  assign \new_[5468]_  = \new_[5660]_  ^ \new_[5665]_ ;
  assign \new_[5469]_  = \new_[8857]_  ^ \new_[8762]_ ;
  assign \new_[5470]_  = \new_[5834]_  ^ \new_[5665]_ ;
  assign \new_[5471]_  = \new_[8863]_  ^ \new_[8762]_ ;
  assign \new_[5472]_  = \new_[5663]_  ^ \new_[5662]_ ;
  assign \new_[5473]_  = \new_[8858]_  ^ \new_[8797]_ ;
  assign \new_[5474]_  = \new_[8666]_  ^ \new_[8857]_ ;
  assign \new_[5475]_  = \new_[8665]_  ^ \new_[8444]_ ;
  assign \new_[5476]_  = \new_[8444]_  ^ \new_[8797]_ ;
  assign \new_[5477]_  = \new_[5835]_  ^ \new_[5660]_ ;
  assign \new_[5478]_  = \new_[5836]_  ^ \new_[5662]_ ;
  assign \new_[5479]_  = \new_[5833]_  ^ \new_[5663]_ ;
  assign n3570 = ~\new_[5607]_  | ~\new_[6829]_ ;
  assign \new_[5481]_  = ~\new_[8952]_  | ~\new_[1254]_ ;
  assign \new_[5482]_  = ~\new_[8952]_  | ~\new_[7922]_ ;
  assign \new_[5483]_  = ~\new_[8952]_  | ~\new_[7924]_ ;
  assign \new_[5484]_  = \new_[8622]_  ^ \new_[8682]_ ;
  assign \new_[5485]_  = \new_[8683]_  ^ \new_[8619]_ ;
  assign \new_[5486]_  = \new_[8794]_  ^ \new_[8833]_ ;
  assign \new_[5487]_  = \new_[8795]_  ^ \new_[8832]_ ;
  assign \new_[5488]_  = addroundkey_start_i_reg;
  assign \new_[5489]_  = ~\new_[5555]_ ;
  assign \new_[5490]_  = ~\new_[5557]_ ;
  assign \new_[5491]_  = ~\new_[7304]_  | (~\new_[5695]_  & ~\new_[7592]_ );
  assign \new_[5492]_  = ~\new_[7321]_  | (~\new_[5673]_  & ~\new_[7592]_ );
  assign \new_[5493]_  = ~\new_[7120]_  | (~\new_[5710]_  & ~\new_[7584]_ );
  assign \new_[5494]_  = ~\new_[7172]_  | (~\new_[5674]_  & ~\new_[7592]_ );
  assign \new_[5495]_  = ~\new_[7235]_  | (~\new_[5675]_  & ~\new_[7584]_ );
  assign \new_[5496]_  = ~\new_[7296]_  | (~\new_[5676]_  & ~\new_[7592]_ );
  assign \new_[5497]_  = ~\new_[7301]_  | (~\new_[5678]_  & ~\new_[7592]_ );
  assign \new_[5498]_  = ~\new_[7365]_  | (~\new_[5679]_  & ~\new_[7592]_ );
  assign \new_[5499]_  = ~\new_[7311]_  | (~\new_[5681]_  & ~\new_[7592]_ );
  assign \new_[5500]_  = ~\new_[7178]_  | (~\new_[5694]_  & ~\new_[7592]_ );
  assign \new_[5501]_  = ~\new_[7298]_  | (~\new_[5680]_  & ~\new_[7584]_ );
  assign \new_[5502]_  = ~\new_[7338]_  | (~\new_[5682]_  & ~\new_[7584]_ );
  assign \new_[5503]_  = ~\new_[7372]_  | (~\new_[5683]_  & ~\new_[7584]_ );
  assign \new_[5504]_  = ~\new_[7398]_  | (~\new_[5684]_  & ~\new_[7592]_ );
  assign \new_[5505]_  = ~\new_[7294]_  | (~\new_[5687]_  & ~\new_[7592]_ );
  assign \new_[5506]_  = ~\new_[7299]_  | (~\new_[5688]_  & ~\new_[7592]_ );
  assign \new_[5507]_  = ~\new_[7322]_  | (~\new_[5686]_  & ~\new_[7592]_ );
  assign \new_[5508]_  = ~\new_[7216]_  | (~\new_[5726]_  & ~\new_[7592]_ );
  assign \new_[5509]_  = ~\new_[7370]_  | (~\new_[5689]_  & ~\new_[7592]_ );
  assign \new_[5510]_  = ~\new_[7333]_  | (~\new_[5691]_  & ~\new_[7584]_ );
  assign \new_[5511]_  = ~\new_[7374]_  | (~\new_[5714]_  & ~\new_[7584]_ );
  assign \new_[5512]_  = ~\new_[7231]_  | (~\new_[5685]_  & ~\new_[7592]_ );
  assign \new_[5513]_  = ~\new_[7262]_  | (~\new_[5703]_  & ~\new_[7592]_ );
  assign \new_[5514]_  = ~\new_[7254]_  | (~\new_[5698]_  & ~\new_[7592]_ );
  assign \new_[5515]_  = ~\new_[7295]_  | (~\new_[5692]_  & ~\new_[7592]_ );
  assign \new_[5516]_  = ~\new_[7251]_  | (~\new_[5697]_  & ~\new_[7592]_ );
  assign \new_[5517]_  = ~\new_[7159]_  | (~\new_[5701]_  & ~\new_[7599]_ );
  assign \new_[5518]_  = ~\new_[7170]_  | (~\new_[5709]_  & ~\new_[7592]_ );
  assign \new_[5519]_  = ~\new_[7314]_  | (~\new_[5702]_  & ~\new_[7592]_ );
  assign \new_[5520]_  = ~\new_[7327]_  | (~\new_[5704]_  & ~\new_[7592]_ );
  assign \new_[5521]_  = ~\new_[7286]_  | (~\new_[5705]_  & ~\new_[7584]_ );
  assign \new_[5522]_  = ~\new_[7203]_  | (~\new_[5706]_  & ~\new_[7592]_ );
  assign \new_[5523]_  = ~\new_[7359]_  | (~\new_[5672]_  & ~\new_[7592]_ );
  assign \new_[5524]_  = ~\new_[7236]_  | (~\new_[5700]_  & ~\new_[7602]_ );
  assign \new_[5525]_  = ~\new_[7405]_  | (~\new_[5725]_  & ~\new_[7592]_ );
  assign \new_[5526]_  = ~\new_[7284]_  | (~\new_[5708]_  & ~\new_[7592]_ );
  assign \new_[5527]_  = ~\new_[7223]_  | (~\new_[5707]_  & ~\new_[7592]_ );
  assign \new_[5528]_  = ~\new_[7271]_  | (~\new_[5677]_  & ~\new_[7584]_ );
  assign \new_[5529]_  = ~\new_[7379]_  | (~\new_[5711]_  & ~\new_[7584]_ );
  assign \new_[5530]_  = ~\new_[7361]_  | (~\new_[5712]_  & ~\new_[7584]_ );
  assign \new_[5531]_  = ~\new_[7302]_  | (~\new_[5728]_  & ~\new_[7592]_ );
  assign \new_[5532]_  = ~\new_[7228]_  | (~\new_[5693]_  & ~\new_[7592]_ );
  assign \new_[5533]_  = ~\new_[7176]_  | (~\new_[5690]_  & ~\new_[7592]_ );
  assign \new_[5534]_  = ~\new_[7404]_  | (~\new_[5713]_  & ~\new_[7592]_ );
  assign \new_[5535]_  = ~\new_[7205]_  | (~\new_[5715]_  & ~\new_[7592]_ );
  assign \new_[5536]_  = ~\new_[7364]_  | (~\new_[5716]_  & ~\new_[7592]_ );
  assign \new_[5537]_  = ~\new_[7308]_  | (~\new_[5717]_  & ~\new_[7592]_ );
  assign \new_[5538]_  = ~\new_[7175]_  | (~\new_[5727]_  & ~\new_[7592]_ );
  assign \new_[5539]_  = ~\new_[7207]_  | (~\new_[5718]_  & ~\new_[7592]_ );
  assign \new_[5540]_  = ~\new_[7290]_  | (~\new_[5719]_  & ~\new_[7584]_ );
  assign \new_[5541]_  = ~\new_[7389]_  | (~\new_[5720]_  & ~\new_[7592]_ );
  assign \new_[5542]_  = ~\new_[7214]_  | (~\new_[5699]_  & ~\new_[7592]_ );
  assign \new_[5543]_  = ~\new_[7153]_  | (~\new_[5721]_  & ~\new_[7584]_ );
  assign \new_[5544]_  = ~\new_[7169]_  | (~\new_[5722]_  & ~\new_[7584]_ );
  assign \new_[5545]_  = ~\new_[7181]_  | (~\new_[5696]_  & ~\new_[7592]_ );
  assign \new_[5546]_  = ~\new_[7291]_  | (~\new_[5724]_  & ~\new_[7592]_ );
  assign \new_[5547]_  = ~\new_[7204]_  | (~\new_[5723]_  & ~\new_[7592]_ );
  assign n3565 = ~\new_[5621]_  | (~\new_[7609]_  & ~load_i);
  assign \new_[5549]_  = \new_[5597]_ ;
  assign \new_[5550]_  = \new_[5597]_ ;
  assign \new_[5551]_  = ~\new_[5658]_ ;
  assign \new_[5552]_  = ~\new_[5658]_ ;
  assign \new_[5553]_  = ~\new_[5658]_ ;
  assign \new_[5554]_  = ~\new_[8950]_  | ~\new_[1388]_ ;
  assign \new_[5555]_  = ~\new_[7847]_  | ~\new_[8950]_ ;
  assign \new_[5556]_  = ~\new_[8950]_  | ~\new_[1254]_ ;
  assign \new_[5557]_  = ~\new_[8950]_  | ~\new_[7870]_ ;
  assign \new_[5558]_  = ~\new_[5755]_  & (~\new_[5779]_  | ~\new_[8779]_ );
  assign \new_[5559]_  = ~\new_[5955]_  | (~\new_[5762]_  & ~\new_[5914]_ );
  assign \new_[5560]_  = ~\new_[7464]_  & (~\new_[5955]_  | ~\new_[5763]_ );
  assign \new_[5561]_  = (~\new_[6235]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1249]_ );
  assign \new_[5562]_  = (~\new_[6259]_  | ~\new_[8899]_ ) & (~\new_[8911]_  | ~\new_[8053]_ );
  assign \new_[5563]_  = (~\new_[6260]_  | ~\new_[8916]_ ) & (~\new_[8911]_  | ~\new_[1200]_ );
  assign \new_[5564]_  = (~\new_[6282]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1145]_ );
  assign \new_[5565]_  = (~\new_[6262]_  | ~\new_[8910]_ ) & (~\new_[8932]_  | ~\new_[1100]_ );
  assign \new_[5566]_  = (~\new_[6264]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1384]_ );
  assign \new_[5567]_  = (~\new_[6272]_  | ~\new_[8916]_ ) & (~\new_[8898]_  | ~\new_[1101]_ );
  assign \new_[5568]_  = (~\new_[6266]_  | ~\new_[8916]_ ) & (~\new_[8929]_  | ~\new_[1201]_ );
  assign \new_[5569]_  = (~\new_[6304]_  | ~\new_[8930]_ ) & (~\new_[8907]_  | ~\new_[1113]_ );
  assign \new_[5570]_  = (~\new_[6315]_  | ~\new_[8899]_ ) & (~\new_[8929]_  | ~\new_[8026]_ );
  assign \new_[5571]_  = (~\new_[6292]_  | ~\new_[8909]_ ) & (~\new_[8922]_  | ~\new_[1136]_ );
  assign \new_[5572]_  = (~\new_[6306]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1311]_ );
  assign \new_[5573]_  = (~\new_[6307]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1383]_ );
  assign \new_[5574]_  = (~\new_[6308]_  | ~\new_[8910]_ ) & (~\new_[8922]_  | ~\new_[1217]_ );
  assign \new_[5575]_  = (~\new_[6310]_  | ~\new_[8909]_ ) & (~\new_[8922]_  | ~\new_[1241]_ );
  assign \new_[5576]_  = (~\new_[6321]_  | ~\new_[8899]_ ) & (~\new_[8932]_  | ~\new_[1191]_ );
  assign \new_[5577]_  = (~\new_[6227]_  | ~\new_[8910]_ ) & (~\new_[8932]_  | ~\new_[1458]_ );
  assign \new_[5578]_  = (~\new_[6311]_  | ~\new_[8916]_ ) & (~\new_[8908]_  | ~\new_[1190]_ );
  assign \new_[5579]_  = (~\new_[6317]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1134]_ );
  assign \new_[5580]_  = (~\new_[6322]_  | ~\new_[8899]_ ) & (~\new_[8932]_  | ~\new_[1099]_ );
  assign \new_[5581]_  = (~\new_[6312]_  | ~\new_[8916]_ ) & (~\new_[8922]_  | ~\new_[1314]_ );
  assign \new_[5582]_  = (~\new_[6324]_  | ~\new_[8930]_ ) & (~\new_[8922]_  | ~\new_[1135]_ );
  assign \new_[5583]_  = (~\new_[6319]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1197]_ );
  assign \new_[5584]_  = (~\new_[6316]_  | ~\new_[8916]_ ) & (~\new_[8914]_  | ~\new_[1196]_ );
  assign \new_[5585]_  = (~\new_[6320]_  | ~\new_[8916]_ ) & (~\new_[8911]_  | ~\new_[1198]_ );
  assign \new_[5586]_  = (~\new_[6285]_  | ~\new_[8930]_ ) & (~\new_[8907]_  | ~\new_[1457]_ );
  assign \new_[5587]_  = (~\new_[6309]_  | ~\new_[8930]_ ) & (~\new_[8922]_  | ~\new_[1096]_ );
  assign \new_[5588]_  = (~\new_[6313]_  | ~\new_[8909]_ ) & (~\new_[8908]_  | ~\new_[1243]_ );
  assign \new_[5589]_  = (~\new_[6330]_  | ~\new_[8916]_ ) & (~\new_[8911]_  | ~\new_[1312]_ );
  assign \new_[5590]_  = (~\new_[6341]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1095]_ );
  assign \new_[5591]_  = (~\new_[6343]_  | ~\new_[8930]_ ) & (~\new_[8898]_  | ~\new_[8020]_ );
  assign \new_[5592]_  = (~\new_[6345]_  | ~\new_[8910]_ ) & (~\new_[8898]_  | ~\new_[1385]_ );
  assign \new_[5593]_  = (~\new_[6347]_  | ~\new_[8916]_ ) & (~\new_[8898]_  | ~\new_[1247]_ );
  assign \new_[5594]_  = (~\new_[6349]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1112]_ );
  assign \new_[5595]_  = (~\new_[6351]_  | ~\new_[8909]_ ) & (~\new_[8908]_  | ~\new_[1192]_ );
  assign \new_[5596]_  = (~\new_[6352]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1248]_ );
  assign \new_[5597]_  = ~\new_[5658]_ ;
  assign \new_[5598]_  = (~\new_[5782]_  | ~\new_[7822]_ ) & (~\new_[5883]_  | ~\new_[8784]_ );
  assign \new_[5599]_  = \new_[6739]_  ? \new_[8992]_  : \new_[7991]_ ;
  assign \new_[5600]_  = \new_[6603]_  ? \new_[8991]_  : \new_[8109]_ ;
  assign \new_[5601]_  = \new_[6734]_  ? \new_[8991]_  : \new_[8156]_ ;
  assign \new_[5602]_  = \new_[6736]_  ? \new_[8992]_  : \new_[1089]_ ;
  assign \new_[5603]_  = \new_[6583]_  ? \new_[8991]_  : \new_[8064]_ ;
  assign \new_[5604]_  = \new_[6635]_  ? \new_[8992]_  : \new_[1119]_ ;
  assign \new_[5605]_  = \new_[6737]_  ? \new_[8991]_  : \new_[8150]_ ;
  assign \new_[5606]_  = ~\new_[5658]_ ;
  assign \new_[5607]_  = ~\new_[7428]_  & (~\new_[5955]_  | ~\new_[5785]_ );
  assign \new_[5608]_  = \new_[8875]_  ^ \new_[8869]_ ;
  assign \new_[5609]_  = \new_[8865]_  ^ \new_[8871]_ ;
  assign \new_[5610]_  = \new_[8871]_  ^ \new_[8869]_ ;
  assign \new_[5611]_  = \new_[8865]_  ^ \new_[8875]_ ;
  assign \new_[5612]_  = \\mix1_state_reg[0] ;
  assign \new_[5613]_  = ~\new_[8950]_  | ~\new_[7856]_ ;
  assign \new_[5614]_  = (~\new_[7259]_  | ~\new_[5792]_ ) & (~\new_[6706]_  | ~\new_[6636]_ );
  assign \new_[5615]_  = (~\new_[5793]_  | ~\new_[7259]_ ) & (~\new_[6700]_  | ~\new_[6636]_ );
  assign n3575 = ~\new_[5761]_  | (~\new_[6082]_  & ~\new_[5956]_ );
  assign \new_[5617]_  = ~\new_[5775]_  & (~\new_[5881]_  | ~\new_[8779]_ );
  assign \new_[5618]_  = ~\new_[5773]_  & (~\new_[5890]_  | ~\new_[8779]_ );
  assign \new_[5619]_  = ~\new_[5670]_ ;
  assign \new_[5620]_  = ~\new_[5671]_ ;
  assign \new_[5621]_  = ~\new_[5955]_  | (~\new_[5796]_  & ~\new_[5915]_ );
  assign \new_[5622]_  = (~\new_[6217]_  | ~\new_[8930]_ ) & (~\new_[8932]_  | ~\new_[1186]_ );
  assign \new_[5623]_  = (~\new_[6232]_  | ~\new_[8899]_ ) & (~\new_[8929]_  | ~\new_[8068]_ );
  assign \new_[5624]_  = (~\new_[6228]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1187]_ );
  assign \new_[5625]_  = (~\new_[6237]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1138]_ );
  assign \new_[5626]_  = (~\new_[6346]_  | ~\new_[8930]_ ) & (~\new_[8914]_  | ~\new_[1218]_ );
  assign \new_[5627]_  = (~\new_[6336]_  | ~\new_[8930]_ ) & (~\new_[8908]_  | ~\new_[1143]_ );
  assign \new_[5628]_  = (~\new_[6267]_  | ~\new_[8899]_ ) & (~\new_[8914]_  | ~\new_[1244]_ );
  assign \new_[5629]_  = (~\new_[6251]_  | ~\new_[8899]_ ) & (~\new_[8911]_  | ~\new_[1144]_ );
  assign \new_[5630]_  = (~\new_[6253]_  | ~\new_[8899]_ ) & (~\new_[8914]_  | ~\new_[1459]_ );
  assign \new_[5631]_  = (~\new_[6254]_  | ~\new_[8899]_ ) & (~\new_[8898]_  | ~\new_[1224]_ );
  assign \new_[5632]_  = (~\new_[6255]_  | ~\new_[8899]_ ) & (~\new_[8932]_  | ~\new_[1313]_ );
  assign \new_[5633]_  = (~\new_[6290]_  | ~\new_[8899]_ ) & (~\new_[8932]_  | ~\new_[1320]_ );
  assign \new_[5634]_  = (~\new_[6258]_  | ~\new_[8899]_ ) & (~\new_[8911]_  | ~\new_[1199]_ );
  assign \new_[5635]_  = (~\new_[6284]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1386]_ );
  assign \new_[5636]_  = (~\new_[6287]_  | ~\new_[8910]_ ) & (~\new_[8929]_  | ~\new_[1193]_ );
  assign \new_[5637]_  = (~\new_[6279]_  | ~\new_[8910]_ ) & (~\new_[8907]_  | ~\new_[1245]_ );
  assign \new_[5638]_  = (~\new_[6288]_  | ~\new_[8923]_ ) & (~\new_[8907]_  | ~\new_[1381]_ );
  assign \new_[5639]_  = (~\new_[6289]_  | ~\new_[8899]_ ) & (~\new_[8922]_  | ~\new_[1137]_ );
  assign \new_[5640]_  = (~\new_[6293]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1251]_ );
  assign \new_[5641]_  = (~\new_[6291]_  | ~\new_[8909]_ ) & (~\new_[8908]_  | ~\new_[1250]_ );
  assign \new_[5642]_  = (~\new_[6278]_  | ~\new_[8899]_ ) & (~\new_[8929]_  | ~\new_[1246]_ );
  assign \new_[5643]_  = (~\new_[6241]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1223]_ );
  assign \new_[5644]_  = (~\new_[6300]_  | ~\new_[8916]_ ) & (~\new_[8911]_  | ~\new_[1460]_ );
  assign \new_[5645]_  = (~\new_[6301]_  | ~\new_[8899]_ ) & (~\new_[8932]_  | ~\new_[8101]_ );
  assign \new_[5646]_  = (~\new_[6314]_  | ~\new_[8909]_ ) & (~\new_[8908]_  | ~\new_[1242]_ );
  assign \new_[5647]_  = (~\new_[6318]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1098]_ );
  assign \new_[5648]_  = (~\new_[6325]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1094]_ );
  assign \new_[5649]_  = (~\new_[6335]_  | ~\new_[8909]_ ) & (~\new_[8914]_  | ~\new_[1210]_ );
  assign \new_[5650]_  = (~\new_[6326]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1194]_ );
  assign \new_[5651]_  = (~\new_[6276]_  | ~\new_[8909]_ ) & (~\new_[8911]_  | ~\new_[1142]_ );
  assign \new_[5652]_  = (~\new_[6334]_  | ~\new_[8910]_ ) & (~\new_[8922]_  | ~\new_[1097]_ );
  assign \new_[5653]_  = (~\new_[6286]_  | ~\new_[8924]_ ) & (~\new_[8914]_  | ~\new_[1252]_ );
  assign \new_[5654]_  = (~\new_[6338]_  | ~\new_[8909]_ ) & (~\new_[8907]_  | ~\new_[1195]_ );
  assign \new_[5655]_  = (~\new_[6340]_  | ~\new_[8910]_ ) & (~\new_[8908]_  | ~\new_[1225]_ );
  assign \new_[5656]_  = ~\new_[5777]_  & (~\new_[5882]_  | ~\new_[7822]_ );
  assign \new_[5657]_  = ~\new_[5774]_  & (~\new_[5885]_  | ~\new_[8784]_ );
  assign \new_[5658]_  = ~\new_[7269]_  & ~\new_[8991]_ ;
  assign \new_[5659]_  = \\mix1_state_reg[1] ;
  assign \new_[5660]_  = \new_[5833]_  ^ \new_[5834]_ ;
  assign \new_[5661]_  = \new_[8858]_  ^ \new_[8665]_ ;
  assign \new_[5662]_  = \new_[5835]_  ^ \new_[5833]_ ;
  assign \new_[5663]_  = \new_[5834]_  ^ \new_[5836]_ ;
  assign \new_[5664]_  = \new_[8863]_  ^ \new_[8666]_ ;
  assign \new_[5665]_  = \new_[5835]_  ^ \new_[5836]_ ;
  assign \new_[5666]_  = (~\new_[5839]_  | ~\new_[7259]_ ) & (~\new_[6699]_  | ~\new_[6636]_ );
  assign \new_[5667]_  = (~\new_[5840]_  | ~\new_[7259]_ ) & (~\new_[6823]_  | ~\new_[6636]_ );
  assign \new_[5668]_  = (~\new_[5838]_  | ~\new_[7259]_ ) & (~\new_[6956]_  | ~\new_[6636]_ );
  assign \new_[5669]_  = ~\new_[8566]_ ;
  assign \new_[5670]_  = \new_[5853]_  ^ \new_[5844]_ ;
  assign \new_[5671]_  = \new_[5855]_  ^ \new_[5847]_ ;
  assign \new_[5672]_  = (~\new_[6294]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1151]_ );
  assign \new_[5673]_  = (~\new_[6229]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1207]_ );
  assign \new_[5674]_  = (~\new_[6231]_  | ~\new_[8923]_ ) & (~\new_[8932]_  | ~\new_[1147]_ );
  assign \new_[5675]_  = (~\new_[6269]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1463]_ );
  assign \new_[5676]_  = (~\new_[6236]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1322]_ );
  assign \new_[5677]_  = (~\new_[6299]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1108]_ );
  assign \new_[5678]_  = (~\new_[6238]_  | ~\new_[8924]_ ) & (~\new_[8929]_  | ~\new_[1206]_ );
  assign \new_[5679]_  = (~\new_[6239]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1216]_ );
  assign \new_[5680]_  = (~\new_[6240]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1530]_ );
  assign \new_[5681]_  = (~\new_[6242]_  | ~\new_[8923]_ ) & (~\new_[8907]_  | ~\new_[1215]_ );
  assign \new_[5682]_  = (~\new_[6243]_  | ~\new_[8924]_ ) & (~\new_[8911]_  | ~\new_[1106]_ );
  assign \new_[5683]_  = (~\new_[6244]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1115]_ );
  assign \new_[5684]_  = (~\new_[6245]_  | ~\new_[8923]_ ) & (~\new_[8898]_  | ~\new_[1107]_ );
  assign \new_[5685]_  = (~\new_[6246]_  | ~\new_[8916]_ ) & (~\new_[8898]_  | ~\new_[1114]_ );
  assign \new_[5686]_  = (~\new_[6248]_  | ~\new_[8909]_ ) & (~\new_[8929]_  | ~\new_[1315]_ );
  assign \new_[5687]_  = (~\new_[6249]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1219]_ );
  assign \new_[5688]_  = (~\new_[6250]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1208]_ );
  assign \new_[5689]_  = (~\new_[6257]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1203]_ );
  assign \new_[5690]_  = (~\new_[6268]_  | ~\new_[8923]_ ) & (~\new_[8932]_  | ~\new_[1202]_ );
  assign \new_[5691]_  = (~\new_[6302]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1150]_ );
  assign \new_[5692]_  = (~\new_[6234]_  | ~\new_[8916]_ ) & (~\new_[8898]_  | ~\new_[1105]_ );
  assign \new_[5693]_  = (~\new_[6331]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1323]_ );
  assign \new_[5694]_  = (~\new_[6233]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1103]_ );
  assign \new_[5695]_  = (~\new_[6263]_  | ~\new_[8923]_ ) & (~\new_[8914]_  | ~\new_[1221]_ );
  assign \new_[5696]_  = (~\new_[6265]_  | ~\new_[8916]_ ) & (~\new_[8907]_  | ~\new_[1204]_ );
  assign \new_[5697]_  = (~\new_[6271]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1104]_ );
  assign \new_[5698]_  = (~\new_[6273]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1117]_ );
  assign \new_[5699]_  = (~\new_[6275]_  | ~\new_[8923]_ ) & (~\new_[8932]_  | ~\new_[1222]_ );
  assign \new_[5700]_  = (~\new_[6277]_  | ~\new_[8909]_ ) & (~\new_[8908]_  | ~\new_[1226]_ );
  assign \new_[5701]_  = (~\new_[6274]_  | ~\new_[8899]_ ) & (~\new_[8929]_  | ~\new_[7939]_ );
  assign \new_[5702]_  = (~\new_[6281]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1205]_ );
  assign \new_[5703]_  = (~\new_[6270]_  | ~\new_[8916]_ ) & (~\new_[8898]_  | ~\new_[1116]_ );
  assign \new_[5704]_  = (~\new_[6283]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1209]_ );
  assign \new_[5705]_  = (~\new_[6256]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1538]_ );
  assign \new_[5706]_  = (~\new_[6261]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1237]_ );
  assign \new_[5707]_  = (~\new_[6295]_  | ~\new_[8924]_ ) & (~\new_[8929]_  | ~\new_[1464]_ );
  assign \new_[5708]_  = (~\new_[6297]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1324]_ );
  assign \new_[5709]_  = (~\new_[6298]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1240]_ );
  assign \new_[5710]_  = (~\new_[6303]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1149]_ );
  assign \new_[5711]_  = (~\new_[6339]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1109]_ );
  assign \new_[5712]_  = (~\new_[6305]_  | ~\new_[8923]_ ) & (~\new_[8914]_  | ~\new_[1238]_ );
  assign \new_[5713]_  = (~\new_[6333]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1152]_ );
  assign \new_[5714]_  = (~\new_[6247]_  | ~\new_[8923]_ ) & (~\new_[8907]_  | ~\new_[1520]_ );
  assign \new_[5715]_  = (~\new_[6323]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1521]_ );
  assign \new_[5716]_  = (~\new_[6327]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1321]_ );
  assign \new_[5717]_  = (~\new_[6328]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1211]_ );
  assign \new_[5718]_  = (~\new_[6329]_  | ~\new_[8909]_ ) & (~\new_[8932]_  | ~\new_[1212]_ );
  assign \new_[5719]_  = (~\new_[6332]_  | ~\new_[8923]_ ) & (~\new_[8929]_  | ~\new_[1110]_ );
  assign \new_[5720]_  = (~\new_[6230]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1111]_ );
  assign \new_[5721]_  = (~\new_[6337]_  | ~\new_[8924]_ ) & (~\new_[8929]_  | ~\new_[1213]_ );
  assign \new_[5722]_  = (~\new_[6344]_  | ~\new_[8916]_ ) & (~\new_[8911]_  | ~\new_[1148]_ );
  assign \new_[5723]_  = (~\new_[6350]_  | ~\new_[8923]_ ) & (~\new_[8932]_  | ~\new_[1234]_ );
  assign \new_[5724]_  = (~\new_[6348]_  | ~\new_[8916]_ ) & (~\new_[8914]_  | ~\new_[1461]_ );
  assign \new_[5725]_  = (~\new_[6296]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1214]_ );
  assign \new_[5726]_  = (~\new_[6252]_  | ~\new_[8924]_ ) & (~\new_[8907]_  | ~\new_[1102]_ );
  assign \new_[5727]_  = (~\new_[6353]_  | ~\new_[8924]_ ) & (~\new_[8898]_  | ~\new_[1319]_ );
  assign \new_[5728]_  = (~\new_[6342]_  | ~\new_[8909]_ ) & (~\new_[8898]_  | ~\new_[1220]_ );
  assign \new_[5729]_  = ~\new_[5821]_  | (~\new_[6741]_  & ~\new_[8991]_ );
  assign \new_[5730]_  = ~\new_[5817]_  | (~\new_[6608]_  & ~\new_[8992]_ );
  assign \new_[5731]_  = ~\new_[5815]_  | (~\new_[6735]_  & ~\new_[8992]_ );
  assign \new_[5732]_  = ~\new_[5819]_  | (~\new_[6742]_  & ~\new_[8991]_ );
  assign \new_[5733]_  = \new_[6898]_  ? \new_[8992]_  : \new_[8094]_ ;
  assign \new_[5734]_  = \new_[7054]_  ? \new_[8991]_  : \new_[1133]_ ;
  assign \new_[5735]_  = \new_[7047]_  ? \new_[8992]_  : \new_[1125]_ ;
  assign \new_[5736]_  = \new_[6773]_  ? \new_[8991]_  : \new_[8130]_ ;
  assign \new_[5737]_  = \new_[7061]_  ? \new_[8992]_  : \new_[1126]_ ;
  assign \new_[5738]_  = \new_[6762]_  ? \new_[8992]_  : \new_[1132]_ ;
  assign \new_[5739]_  = \new_[7041]_  ? \new_[8992]_  : \new_[1141]_ ;
  assign \new_[5740]_  = ~\new_[5816]_  | (~\new_[6924]_  & ~\new_[8992]_ );
  assign \new_[5741]_  = ~\new_[5825]_  | (~\new_[6738]_  & ~\new_[8992]_ );
  assign \new_[5742]_  = ~\new_[5818]_  | (~\new_[7055]_  & ~\new_[8992]_ );
  assign \new_[5743]_  = ~\new_[5820]_  | (~\new_[7048]_  & ~\new_[8991]_ );
  assign \new_[5744]_  = ~\new_[5822]_  | (~\new_[7039]_  & ~\new_[8991]_ );
  assign \new_[5745]_  = ~\new_[5823]_  | (~\new_[7053]_  & ~\new_[8992]_ );
  assign \new_[5746]_  = ~\new_[5824]_  | (~\new_[6743]_  & ~\new_[8992]_ );
  assign \new_[5747]_  = \new_[6899]_  ? \new_[8992]_  : \new_[8037]_ ;
  assign \new_[5748]_  = ~\new_[5826]_  | (~\new_[6744]_  & ~\new_[8992]_ );
  assign \new_[5749]_  = ~\new_[8563]_  & (~\new_[5939]_  | ~\new_[5895]_ );
  assign \new_[5750]_  = ~\new_[8563]_  & (~\new_[5897]_  | ~\new_[5891]_ );
  assign \new_[5751]_  = ~\new_[7829]_  & (~\new_[5941]_  | ~\new_[5893]_ );
  assign \new_[5752]_  = ~\new_[7829]_  & (~\new_[5902]_  | ~\new_[5829]_ );
  assign \new_[5753]_  = ~\new_[8562]_  & (~\new_[5938]_  | ~\new_[5892]_ );
  assign \new_[5754]_  = ~\new_[7829]_  & (~\new_[5901]_  | ~\new_[5831]_ );
  assign \new_[5755]_  = ~\new_[7829]_  & (~\new_[5896]_  | ~\new_[5894]_ );
  assign \new_[5756]_  = (~\new_[5906]_  | ~\new_[7259]_ ) & (~\new_[6826]_  | ~\new_[6636]_ );
  assign \new_[5757]_  = (~\new_[5905]_  | ~\new_[7259]_ ) & (~\new_[6822]_  | ~\new_[6636]_ );
  assign n3580 = ~\new_[5837]_  | ~\new_[7829]_ ;
  assign \new_[5759]_  = ~\new_[5878]_  & (~\new_[5979]_  | ~\new_[8779]_ );
  assign \new_[5760]_  = ~\new_[5876]_  & (~\new_[5976]_  | ~\new_[8779]_ );
  assign \new_[5761]_  = ~\new_[5841]_  & (~\new_[7206]_  | ~\new_[5784]_ );
  assign \new_[5762]_  = ~\new_[6919]_  & ~\new_[5850]_ ;
  assign \new_[5763]_  = (~\new_[6788]_  & ~\new_[6202]_ ) | (~\new_[6919]_  & ~\new_[5918]_ );
  assign \new_[5764]_  = \new_[5828]_  & \new_[6198]_ ;
  assign \new_[5765]_  = ~\new_[5858]_  | ~\new_[6101]_ ;
  assign \new_[5766]_  = ~\new_[5877]_  & (~\new_[5980]_  | ~\new_[8784]_ );
  assign \new_[5767]_  = ~\new_[5873]_  | (~\new_[6740]_  & ~\new_[8992]_ );
  assign \new_[5768]_  = ~\new_[5871]_  | (~\new_[7051]_  & ~\new_[8992]_ );
  assign \new_[5769]_  = ~\new_[5874]_  | (~\new_[7059]_  & ~\new_[8992]_ );
  assign \new_[5770]_  = ~\new_[5872]_  | (~\new_[7060]_  & ~\new_[8992]_ );
  assign \new_[5771]_  = (~\new_[7040]_  & ~\new_[8991]_ ) | (~\new_[2025]_  & ~\new_[8993]_ );
  assign \new_[5772]_  = ~\new_[8563]_  & (~\new_[5985]_  | ~\new_[5934]_ );
  assign \new_[5773]_  = ~\new_[8563]_  & (~\new_[5943]_  | ~\new_[5936]_ );
  assign \new_[5774]_  = ~\new_[7829]_  & (~\new_[5986]_  | ~\new_[5935]_ );
  assign \new_[5775]_  = ~\new_[8562]_  & (~\new_[5940]_  | ~\new_[5937]_ );
  assign \new_[5776]_  = ~\new_[7829]_  & (~\new_[5987]_  | ~\new_[5899]_ );
  assign \new_[5777]_  = ~\new_[7829]_  & (~\new_[5984]_  | ~\new_[5900]_ );
  assign \new_[5778]_  = \data_o[121]  ? \new_[8912]_  : \new_[8101]_ ;
  assign \new_[5779]_  = \data_o[105]  ? \new_[8934]_  : \new_[1457]_ ;
  assign \new_[5780]_  = \data_o[89]  ? \new_[8934]_  : \new_[7939]_ ;
  assign \new_[5781]_  = \data_o[65]  ? \new_[8915]_  : \new_[1463]_ ;
  assign \new_[5782]_  = \data_o[73]  ? \new_[8934]_  : \new_[1459]_ ;
  assign \new_[5783]_  = \data_o[97]  ? \new_[8899]_  : \new_[1464]_ ;
  assign \new_[5784]_  = ~state_reg;
  assign \new_[5785]_  = (~\new_[6163]_  & ~\new_[6788]_ ) | (~\new_[6919]_  & ~\new_[5951]_ );
  assign n3585 = ~\new_[8562]_  | ~\new_[7829]_  | ~\new_[5944]_ ;
  assign \new_[5787]_  = ~\new_[5927]_  & (~\new_[5977]_  | ~\new_[8779]_ );
  assign \new_[5788]_  = ~\new_[5930]_  & (~\new_[5982]_  | ~\new_[8779]_ );
  assign \new_[5789]_  = ~\new_[5933]_  & (~\new_[6042]_  | ~\new_[8779]_ );
  assign \new_[5790]_  = ~\new_[5923]_  & (~\new_[5971]_  | ~\new_[8779]_ );
  assign \new_[5791]_  = ~\new_[5924]_  & (~\new_[5981]_  | ~\new_[8779]_ );
  assign \new_[5792]_  = ~\new_[6220]_  | ~\new_[6096]_  | ~\new_[5908]_  | ~\new_[6374]_ ;
  assign \new_[5793]_  = ~\new_[6179]_  | ~\new_[6095]_  | ~\new_[5907]_  | ~\new_[6097]_ ;
  assign \new_[5794]_  = \new_[5998]_  | \new_[5913]_ ;
  assign \new_[5795]_  = ~\new_[5848]_ ;
  assign \new_[5796]_  = ~\new_[6919]_  & ~\new_[5920]_ ;
  assign \new_[5797]_  = ~\new_[5856]_ ;
  assign \new_[5798]_  = ~\new_[5928]_  & (~\new_[5945]_  | ~\new_[8558]_ );
  assign \new_[5799]_  = ~\new_[5929]_  & (~\new_[5973]_  | ~\new_[8558]_ );
  assign \new_[5800]_  = ~\new_[5932]_  & (~\new_[5992]_  | ~\new_[8784]_ );
  assign \new_[5801]_  = (~\new_[5970]_  | ~\new_[8558]_ ) & (~\new_[6040]_  | ~\new_[8784]_ );
  assign \new_[5802]_  = (~\new_[5946]_  | ~\new_[7822]_ ) & (~\new_[5972]_  | ~\new_[8784]_ );
  assign \new_[5803]_  = ~\new_[5926]_  & (~\new_[5969]_  | ~\new_[8784]_ );
  assign \new_[5804]_  = \new_[7142]_  ? \new_[8991]_  : \new_[2353]_ ;
  assign \new_[5805]_  = \new_[7140]_  ? \new_[8991]_  : \new_[2350]_ ;
  assign \new_[5806]_  = ~\new_[5922]_  | (~\new_[7042]_  & ~\new_[8992]_ );
  assign \new_[5807]_  = \new_[7149]_  ? \new_[8992]_  : \new_[2352]_ ;
  assign \new_[5808]_  = \new_[7143]_  ? \new_[8991]_  : \new_[7949]_ ;
  assign \new_[5809]_  = \new_[7112]_  ? \new_[8992]_  : \new_[2422]_ ;
  assign \new_[5810]_  = \new_[7119]_  ? \new_[8992]_  : \new_[2351]_ ;
  assign \new_[5811]_  = ~\new_[5921]_  | (~\new_[7049]_  & ~\new_[8992]_ );
  assign \new_[5812]_  = \new_[7100]_  ? \new_[8992]_  : \new_[2423]_ ;
  assign \new_[5813]_  = \new_[7046]_  ? \new_[8992]_  : \new_[2411]_ ;
  assign \new_[5814]_  = \new_[7050]_  ? \new_[8992]_  : \new_[2461]_ ;
  assign \new_[5815]_  = ~\new_[2162]_  | ~\new_[8992]_ ;
  assign \new_[5816]_  = ~\new_[2198]_  | ~\new_[8992]_ ;
  assign \new_[5817]_  = ~\new_[2069]_  | ~\new_[8992]_ ;
  assign \new_[5818]_  = ~\new_[2199]_  | ~\new_[8992]_ ;
  assign \new_[5819]_  = ~\new_[2067]_  | ~\new_[8991]_ ;
  assign \new_[5820]_  = ~\new_[2200]_  | ~\new_[8992]_ ;
  assign \new_[5821]_  = ~\new_[2068]_  | ~\new_[8991]_ ;
  assign \new_[5822]_  = ~\new_[2201]_  | ~\new_[8992]_ ;
  assign \new_[5823]_  = ~\new_[2203]_  | ~\new_[8992]_ ;
  assign \new_[5824]_  = ~\new_[2070]_  | ~\new_[8991]_ ;
  assign \new_[5825]_  = ~\new_[2202]_  | ~\new_[8992]_ ;
  assign \new_[5826]_  = ~\new_[2043]_  | ~\new_[8991]_ ;
  assign \new_[5827]_  = ~\new_[7829]_  & (~\new_[5988]_  | ~\new_[5983]_ );
  assign \new_[5828]_  = ~\new_[7269]_  | ~\new_[5965]_ ;
  assign \new_[5829]_  = ~\new_[8911]_  | ~\data_o[57] ;
  assign \new_[5830]_  = \data_o[0]  ? \new_[8924]_  : \new_[8026]_ ;
  assign \new_[5831]_  = ~\new_[8929]_  | ~\data_o[49] ;
  assign \new_[5832]_  = \new_[7092]_  ? \new_[8992]_  : \new_[8075]_ ;
  assign \new_[5833]_  = ~\new_[5964]_  | ~\new_[5948]_ ;
  assign \new_[5834]_  = ~\new_[6033]_  | ~\new_[5947]_ ;
  assign \new_[5835]_  = ~\new_[5963]_  | ~\new_[5949]_ ;
  assign \new_[5836]_  = ~\new_[5959]_  | ~\new_[5950]_ ;
  assign \new_[5837]_  = ~\new_[8713]_  | (~\new_[8710]_  & ~\new_[5612]_ );
  assign \new_[5838]_  = ~\new_[6377]_  | ~\new_[6182]_  | ~\new_[5954]_  | ~\new_[6492]_ ;
  assign \new_[5839]_  = ~\new_[6373]_  | ~\new_[6378]_  | ~\new_[5953]_  | ~\new_[6093]_ ;
  assign \new_[5840]_  = ~\new_[6280]_  | ~\new_[6183]_  | ~\new_[5952]_  | ~\new_[6094]_ ;
  assign \new_[5841]_  = ~\new_[5956]_  & ~\new_[6079]_ ;
  assign \new_[5842]_  = ~\new_[5910]_ ;
  assign \new_[5843]_  = ~\new_[9005]_  | ~\new_[1227]_ ;
  assign \new_[5844]_  = ~\new_[9005]_  | ~\new_[1709]_ ;
  assign \new_[5845]_  = ~\new_[5911]_ ;
  assign \new_[5846]_  = ~\new_[5912]_ ;
  assign \new_[5847]_  = ~\new_[9005]_  | ~\new_[1388]_ ;
  assign \new_[5848]_  = ~\new_[9005]_  | ~\new_[1592]_ ;
  assign \new_[5849]_  = ~\new_[5942]_  | ~\new_[6171]_ ;
  assign \new_[5850]_  = \new_[6030]_  ? \new_[7906]_  : \new_[7675]_ ;
  assign \new_[5851]_  = \new_[8970]_  & \new_[1388]_ ;
  assign \new_[5852]_  = ~\new_[5916]_ ;
  assign \new_[5853]_  = ~\new_[8970]_  | ~\new_[1227]_ ;
  assign \new_[5854]_  = ~\new_[5917]_ ;
  assign \new_[5855]_  = ~\new_[8970]_  | ~\new_[1254]_ ;
  assign \new_[5856]_  = ~\new_[8970]_  | ~\new_[7856]_ ;
  assign \new_[5857]_  = ~\new_[5962]_  | ~\new_[6114]_ ;
  assign \new_[5858]_  = ~\new_[7269]_  | ~\new_[5966]_ ;
  assign \new_[5859]_  = \new_[7111]_  ? \new_[8991]_  : \new_[2537]_ ;
  assign \new_[5860]_  = \new_[7095]_  ? \new_[8992]_  : \new_[2425]_ ;
  assign \new_[5861]_  = \new_[7103]_  ? \new_[8992]_  : \new_[7971]_ ;
  assign \new_[5862]_  = \new_[7148]_  ? \new_[8991]_  : \new_[7986]_ ;
  assign \new_[5863]_  = \new_[7094]_  ? \new_[8992]_  : \new_[8004]_ ;
  assign \new_[5864]_  = \new_[7045]_  ? \new_[8992]_  : \new_[2348]_ ;
  assign \new_[5865]_  = \new_[7052]_  ? \new_[8992]_  : \new_[2424]_ ;
  assign \new_[5866]_  = \new_[7141]_  ? \new_[8991]_  : \new_[7984]_ ;
  assign \new_[5867]_  = \new_[7044]_  ? \new_[8992]_  : \new_[2421]_ ;
  assign \new_[5868]_  = \new_[7144]_  ? \new_[8992]_  : \new_[2354]_ ;
  assign \new_[5869]_  = \new_[7058]_  ? \new_[8992]_  : \new_[2344]_ ;
  assign \new_[5870]_  = \new_[7037]_  ? \new_[8992]_  : \new_[2349]_ ;
  assign \new_[5871]_  = ~\new_[2132]_  | ~\new_[8992]_ ;
  assign \new_[5872]_  = ~\new_[2139]_  | ~\new_[8992]_ ;
  assign \new_[5873]_  = ~\new_[2135]_  | ~\new_[8992]_ ;
  assign \new_[5874]_  = ~\new_[2133]_  | ~\new_[8992]_ ;
  assign \new_[5875]_  = ~\new_[8563]_  & (~\new_[6128]_  | ~\new_[6046]_ );
  assign \new_[5876]_  = ~\new_[7829]_  & (~\new_[6052]_  | ~\new_[6043]_ );
  assign \new_[5877]_  = ~\new_[7902]_  & (~\new_[6051]_  | ~\new_[6044]_ );
  assign \new_[5878]_  = ~\new_[8562]_  & (~\new_[6050]_  | ~\new_[6047]_ );
  assign \new_[5879]_  = ~\new_[7902]_  & (~\new_[6129]_  | ~\new_[6048]_ );
  assign \new_[5880]_  = \data_o[113]  ? \new_[8899]_  : \new_[1530]_ ;
  assign \new_[5881]_  = \data_o[104]  ? \new_[8913]_  : \new_[1142]_ ;
  assign \new_[5882]_  = \data_o[80]  ? \new_[8930]_  : \new_[1150]_ ;
  assign \new_[5883]_  = \data_o[9]  ? \new_[8915]_  : \new_[1460]_ ;
  assign \new_[5884]_  = \data_o[17]  ? \new_[8910]_  : \new_[1461]_ ;
  assign \new_[5885]_  = \data_o[8]  ? \new_[8915]_  : \new_[1145]_ ;
  assign \new_[5886]_  = \data_o[120]  ? \new_[8931]_  : \new_[1223]_ ;
  assign \new_[5887]_  = \data_o[88]  ? \new_[8912]_  : \new_[1226]_ ;
  assign \new_[5888]_  = \data_o[96]  ? \new_[8931]_  : \new_[1151]_ ;
  assign \new_[5889]_  = \data_o[64]  ? \new_[8934]_  : \new_[1149]_ ;
  assign \new_[5890]_  = \data_o[112]  ? \new_[8930]_  : \new_[1147]_ ;
  assign \new_[5891]_  = ~\new_[8911]_  | ~\data_o[25] ;
  assign \new_[5892]_  = ~\new_[8933]_  | ~\data_o[81] ;
  assign \new_[5893]_  = ~\new_[8907]_  | ~\data_o[33] ;
  assign \new_[5894]_  = ~\new_[8898]_  | ~\data_o[41] ;
  assign \new_[5895]_  = ~\new_[8914]_  | ~\data_o[1] ;
  assign \new_[5896]_  = ~\new_[8912]_  | ~\new_[1458]_ ;
  assign \new_[5897]_  = ~\new_[8899]_  | ~\new_[8053]_ ;
  assign \new_[5898]_  = \\sub1_state_reg[0] ;
  assign \new_[5899]_  = ~\new_[8917]_  | ~\data_o[56] ;
  assign \new_[5900]_  = ~\new_[8917]_  | ~\data_o[48] ;
  assign \new_[5901]_  = ~\new_[8916]_  | ~\new_[1521]_ ;
  assign \new_[5902]_  = ~\new_[8916]_  | ~\new_[8020]_ ;
  assign \new_[5903]_  = ~\new_[6038]_  & (~\new_[6403]_  | ~\new_[8780]_ );
  assign \new_[5904]_  = ~\new_[6037]_  & (~\new_[6152]_  | ~\new_[8780]_ );
  assign \new_[5905]_  = ~\new_[6375]_  | ~\new_[6185]_  | ~\new_[5994]_  | ~\new_[6175]_ ;
  assign \new_[5906]_  = ~\new_[6381]_  | ~\new_[6379]_  | ~\new_[5995]_  | ~\new_[6181]_ ;
  assign \new_[5907]_  = ~\new_[5997]_  & ~\new_[6178]_ ;
  assign \new_[5908]_  = ~\new_[5996]_  & ~\new_[6176]_ ;
  assign n3590 = ~\new_[7585]_  | (~\new_[6081]_  & ~\new_[5784]_ );
  assign \new_[5910]_  = ~\new_[9005]_  | ~\new_[7856]_ ;
  assign \new_[5911]_  = ~\new_[9005]_  | ~\new_[1254]_ ;
  assign \new_[5912]_  = ~\new_[9005]_  | ~\new_[7924]_ ;
  assign \new_[5913]_  = ~\new_[6184]_  | ~\new_[6380]_  | ~\new_[6412]_  | ~\new_[6174]_ ;
  assign \new_[5914]_  = ~\new_[6030]_  & ~\new_[6788]_ ;
  assign \new_[5915]_  = ~\new_[6788]_  & ~\new_[6112]_ ;
  assign \new_[5916]_  = ~\new_[8971]_  | ~\new_[1592]_ ;
  assign \new_[5917]_  = ~\new_[8970]_  | ~\new_[7870]_ ;
  assign \new_[5918]_  = ~\new_[6031]_  & (~\new_[7848]_  | ~\new_[7906]_ );
  assign \new_[5919]_  = ~\new_[5989]_  & (~\new_[6219]_  | ~\new_[8784]_ );
  assign \new_[5920]_  = \new_[6112]_  ? \new_[7906]_  : \new_[7926]_ ;
  assign \new_[5921]_  = ~\new_[1456]_  | ~\new_[8992]_ ;
  assign \new_[5922]_  = ~\new_[1455]_  | ~\new_[8991]_ ;
  assign \new_[5923]_  = ~\new_[8563]_  & (~\new_[6125]_  | ~\new_[6071]_ );
  assign \new_[5924]_  = ~\new_[8563]_  & (~\new_[6131]_  | ~\new_[6120]_ );
  assign ready_o = ready_o_reg;
  assign \new_[5926]_  = ~\new_[7902]_  & (~\new_[6132]_  | ~\new_[6122]_ );
  assign \new_[5927]_  = ~\new_[7902]_  & (~\new_[6126]_  | ~\new_[6116]_ );
  assign \new_[5928]_  = ~\new_[7902]_  & (~\new_[6130]_  | ~\new_[6118]_ );
  assign \new_[5929]_  = ~\new_[7902]_  & (~\new_[6127]_  | ~\new_[6117]_ );
  assign \new_[5930]_  = ~\new_[8562]_  & (~\new_[6072]_  | ~\new_[6123]_ );
  assign \new_[5931]_  = ~\new_[8562]_  & (~\new_[6153]_  | ~\new_[6121]_ );
  assign \new_[5932]_  = ~\new_[7902]_  & (~\new_[6212]_  | ~\new_[6124]_ );
  assign \new_[5933]_  = ~\new_[8562]_  & (~\new_[6150]_  | ~\new_[6115]_ );
  assign \new_[5934]_  = ~\new_[8897]_  | ~\data_o[24] ;
  assign \new_[5935]_  = ~\new_[8917]_  | ~\data_o[40] ;
  assign \new_[5936]_  = ~\new_[8917]_  | ~\data_o[16] ;
  assign \new_[5937]_  = ~\new_[8917]_  | ~\data_o[72] ;
  assign \new_[5938]_  = ~\new_[8910]_  | ~\new_[1520]_ ;
  assign \new_[5939]_  = ~\new_[8912]_  | ~\new_[8068]_ ;
  assign \new_[5940]_  = ~\new_[8931]_  | ~\new_[1144]_ ;
  assign \new_[5941]_  = ~\new_[8912]_  | ~\new_[1538]_ ;
  assign \new_[5942]_  = ~\new_[7269]_  | ~\new_[6099]_ ;
  assign \new_[5943]_  = ~\new_[8928]_  | ~\new_[1148]_ ;
  assign \new_[5944]_  = ~\new_[5659]_  | ~\new_[8469]_  | ~\new_[8713]_ ;
  assign \new_[5945]_  = \data_o[90]  ? \new_[8946]_  : \new_[1386]_ ;
  assign \new_[5946]_  = \data_o[76]  ? \new_[8896]_  : \new_[1200]_ ;
  assign \new_[5947]_  = ~\new_[6110]_  & (~\new_[6203]_  | ~\new_[8780]_ );
  assign \new_[5948]_  = ~\new_[6106]_  & (~\new_[6206]_  | ~\new_[8780]_ );
  assign \new_[5949]_  = ~\new_[6098]_  & (~\new_[6226]_  | ~\new_[8780]_ );
  assign \new_[5950]_  = ~\new_[6187]_  & (~\new_[6205]_  | ~\new_[8780]_ );
  assign \new_[5951]_  = \new_[6163]_  ? \new_[7906]_  : \new_[7580]_ ;
  assign \new_[5952]_  = ~\new_[6078]_  & ~\new_[6222]_ ;
  assign \new_[5953]_  = ~\new_[6076]_  & ~\new_[6180]_ ;
  assign \new_[5954]_  = ~\new_[6077]_  & ~\new_[6177]_ ;
  assign \new_[5955]_  = ~\new_[6082]_  | ~\new_[6079]_ ;
  assign \new_[5956]_  = (~\new_[6418]_  | ~\new_[6919]_ ) & (~\new_[6788]_  | ~\new_[7906]_ );
  assign \new_[5957]_  = ~\new_[1096]_  | ~\new_[6092]_ ;
  assign \new_[5958]_  = ~\new_[1097]_  | ~\new_[6092]_ ;
  assign \new_[5959]_  = ~\new_[6111]_  & (~\new_[6204]_  | ~\new_[8558]_ );
  assign \new_[5960]_  = \\sub1_state_reg[3] ;
  assign \new_[5961]_  = ~\new_[6114]_  | ~\new_[6199]_ ;
  assign \new_[5962]_  = ~\new_[7269]_  | ~\new_[6100]_ ;
  assign \new_[5963]_  = ~\new_[6104]_  & (~\new_[6395]_  | ~\new_[8558]_ );
  assign \new_[5964]_  = ~\new_[6105]_  & (~\new_[6209]_  | ~\new_[8784]_ );
  assign \new_[5965]_  = ~\new_[6035]_ ;
  assign \new_[5966]_  = ~\new_[6036]_ ;
  assign \new_[5967]_  = ~\new_[7902]_  & (~\new_[6211]_  | ~\new_[6149]_ );
  assign \new_[5968]_  = ~\new_[7902]_  & (~\new_[6213]_  | ~\new_[6210]_ );
  assign \new_[5969]_  = \data_o[10]  ? \new_[8934]_  : \new_[1312]_ ;
  assign \new_[5970]_  = \data_o[66]  ? \new_[8931]_  : \new_[1322]_ ;
  assign \new_[5971]_  = \data_o[114]  ? \new_[8900]_  : \new_[1315]_ ;
  assign \new_[5972]_  = \data_o[12]  ? \new_[8918]_  : \new_[1194]_ ;
  assign \new_[5973]_  = \data_o[82]  ? \new_[8924]_  : \new_[1323]_ ;
  assign \new_[5974]_  = \data_o[84]  ? \new_[8924]_  : \new_[1220]_ ;
  assign \new_[5975]_  = \data_o[92]  ? \new_[8918]_  : \new_[1252]_ ;
  assign \new_[5976]_  = \data_o[108]  ? \new_[8912]_  : \new_[1191]_ ;
  assign \new_[5977]_  = \data_o[98]  ? \new_[8924]_  : \new_[1324]_ ;
  assign \new_[5978]_  = \data_o[124]  ? \new_[8900]_  : \new_[1242]_ ;
  assign \new_[5979]_  = \data_o[100]  ? \new_[8912]_  : \new_[1234]_ ;
  assign \new_[5980]_  = \data_o[4]  ? \new_[8924]_  : \new_[1210]_ ;
  assign \new_[5981]_  = \data_o[122]  ? \new_[8912]_  : \new_[1383]_ ;
  assign \new_[5982]_  = \data_o[106]  ? \new_[8924]_  : \new_[1311]_ ;
  assign \new_[5983]_  = ~\new_[8897]_  | ~\data_o[32] ;
  assign \new_[5984]_  = ~\new_[8931]_  | ~\new_[1152]_ ;
  assign \new_[5985]_  = ~\new_[8931]_  | ~\new_[1224]_ ;
  assign \new_[5986]_  = ~\new_[8931]_  | ~\new_[1143]_ ;
  assign \new_[5987]_  = ~\new_[8924]_  | ~\new_[1225]_ ;
  assign \new_[5988]_  = ~\new_[8931]_  | ~\new_[1209]_ ;
  assign \new_[5989]_  = ~\new_[7902]_  & (~\new_[6224]_  | ~\new_[6408]_ );
  assign \new_[5990]_  = \\sub1_state_reg[2] ;
  assign \new_[5991]_  = \\sub1_state_reg[1] ;
  assign \new_[5992]_  = \data_o[19]  ? \new_[8896]_  : \new_[1207]_ ;
  assign n3595 = ~\new_[6155]_  | (~\new_[6803]_  & ~\new_[7934]_ );
  assign \new_[5994]_  = ~\new_[6164]_  & ~\new_[6376]_ ;
  assign \new_[5995]_  = ~\new_[6165]_  & ~\new_[6369]_ ;
  assign \new_[5996]_  = ~\new_[6665]_  | ~\new_[6496]_  | ~\new_[6455]_  | ~\new_[6490]_ ;
  assign \new_[5997]_  = ~\new_[6497]_  | ~\new_[6489]_  | ~\new_[6456]_  | ~\new_[6491]_ ;
  assign \new_[5998]_  = ~\new_[6457]_  | ~\new_[6488]_  | ~\new_[6493]_  | ~\new_[6382]_ ;
  assign \new_[5999]_  = ~\new_[6168]_  | ~\new_[1211]_ ;
  assign n3600 = ~\new_[6080]_ ;
  assign \new_[6001]_  = ~\new_[1115]_  | ~\new_[6417]_ ;
  assign \new_[6002]_  = ~\new_[6454]_  | ~\new_[1094]_ ;
  assign \new_[6003]_  = ~\new_[6173]_  | ~\new_[1108]_ ;
  assign \new_[6004]_  = ~\new_[6454]_  | ~\new_[1095]_ ;
  assign \new_[6005]_  = ~\new_[1100]_  | ~\new_[6170]_ ;
  assign \new_[6006]_  = ~\new_[6434]_  | ~\new_[1105]_ ;
  assign \new_[6007]_  = ~\new_[6434]_  | ~\new_[1104]_ ;
  assign \new_[6008]_  = ~\new_[1099]_  | ~\new_[6436]_ ;
  assign \new_[6009]_  = ~\new_[6168]_  | ~\new_[1213]_ ;
  assign \new_[6010]_  = ~\new_[1098]_  | ~\new_[6436]_ ;
  assign \new_[6011]_  = ~\new_[6168]_  | ~\new_[1521]_ ;
  assign \new_[6012]_  = ~\new_[6168]_  | ~\new_[1321]_ ;
  assign \new_[6013]_  = ~\new_[1320]_  | ~\new_[6169]_ ;
  assign \new_[6014]_  = \new_[6173]_  & \new_[1209]_ ;
  assign \new_[6015]_  = ~\new_[6169]_  | ~\new_[1218]_ ;
  assign \new_[6016]_  = ~\new_[6168]_  | ~\new_[1111]_ ;
  assign \new_[6017]_  = ~\new_[6173]_  | ~\new_[1214]_ ;
  assign \new_[6018]_  = ~\new_[1210]_  | ~\new_[6169]_ ;
  assign \new_[6019]_  = ~\new_[6168]_  | ~\new_[1152]_ ;
  assign \new_[6020]_  = ~\new_[1117]_  | ~\new_[6435]_ ;
  assign \new_[6021]_  = ~\new_[6168]_  | ~\new_[1212]_ ;
  assign \new_[6022]_  = ~\new_[6168]_  | ~\new_[1110]_ ;
  assign \new_[6023]_  = ~\new_[1112]_  | ~\new_[6169]_ ;
  assign \new_[6024]_  = ~\new_[1116]_  | ~\new_[6435]_ ;
  assign \new_[6025]_  = ~\new_[1113]_  | ~\new_[6169]_ ;
  assign \new_[6026]_  = ~\new_[1114]_  | ~\new_[6417]_ ;
  assign \new_[6027]_  = ~\new_[1217]_  | ~\new_[6169]_ ;
  assign \new_[6028]_  = ~\new_[1101]_  | ~\new_[6170]_ ;
  assign \new_[6029]_  = ~\new_[6173]_  | ~\new_[1109]_ ;
  assign \new_[6030]_  = \new_[7675]_  ? \new_[7607]_  : \new_[6393]_ ;
  assign \new_[6031]_  = ~\new_[6202]_  & ~\new_[7906]_ ;
  assign \new_[6032]_  = (~\new_[6401]_  | ~\new_[8784]_ ) & (~\new_[6402]_  | ~\new_[8558]_ );
  assign \new_[6033]_  = ~\new_[6200]_  & (~\new_[6225]_  | ~\new_[8784]_ );
  assign \new_[6034]_  = ~\new_[8563]_  & (~\new_[6560]_  | ~\new_[6221]_ );
  assign \new_[6035]_  = ~\new_[8993]_  | ~\new_[7923]_ ;
  assign \new_[6036]_  = ~\new_[8993]_  | ~\new_[7928]_ ;
  assign \new_[6037]_  = ~\new_[7902]_  & (~\new_[6411]_  | ~\new_[6410]_ );
  assign \new_[6038]_  = ~\new_[8562]_  & (~\new_[6413]_  | ~\new_[6409]_ );
  assign \new_[6039]_  = \data_o[99]  ? \new_[8924]_  : \new_[1240]_ ;
  assign \new_[6040]_  = \data_o[2]  ? \new_[8918]_  : \new_[1320]_ ;
  assign \new_[6041]_  = \\sub1_state_reg[4] ;
  assign \new_[6042]_  = \data_o[115]  ? \new_[8946]_  : \new_[1203]_ ;
  assign \new_[6043]_  = ~\new_[8919]_  | ~\data_o[44] ;
  assign \new_[6044]_  = ~\new_[8914]_  | ~\data_o[36] ;
  assign \new_[6045]_  = ~\new_[8932]_  | ~\data_o[52] ;
  assign \new_[6046]_  = ~\new_[8914]_  | ~\data_o[28] ;
  assign \new_[6047]_  = ~\new_[8911]_  | ~\data_o[68] ;
  assign \new_[6048]_  = ~\new_[8897]_  | ~\data_o[60] ;
  assign \new_[6049]_  = ~\new_[8931]_  | ~\new_[1212]_ ;
  assign \new_[6050]_  = ~\new_[8924]_  | ~\new_[1215]_ ;
  assign \new_[6051]_  = ~\new_[8918]_  | ~\new_[1214]_ ;
  assign \new_[6052]_  = ~\new_[8899]_  | ~\new_[1196]_ ;
  assign \new_[6053]_  = (~\new_[7660]_  | ~\key_i[62] ) & (~\new_[7075]_  | ~\new_[8005]_ );
  assign \new_[6054]_  = (~\new_[7660]_  | ~\key_i[63] ) & (~\new_[7075]_  | ~\new_[7941]_ );
  assign \new_[6055]_  = \key_i[48]  ? \new_[7075]_  : \new_[8008]_ ;
  assign \new_[6056]_  = (~\new_[7660]_  | ~\key_i[59] ) & (~\new_[7075]_  | ~\new_[7957]_ );
  assign \new_[6057]_  = \key_i[53]  ? \new_[7075]_  : \new_[7993]_ ;
  assign \new_[6058]_  = \key_i[58]  ? \new_[7075]_  : \new_[8055]_ ;
  assign \new_[6059]_  = (~\new_[7660]_  | ~\key_i[56] ) & (~\new_[7075]_  | ~\new_[8000]_ );
  assign \new_[6060]_  = \key_i[61]  ? \new_[7075]_  : \new_[8001]_ ;
  assign \new_[6061]_  = \key_i[52]  ? \new_[7075]_  : \new_[8138]_ ;
  assign \new_[6062]_  = \key_i[32]  ? \new_[7075]_  : \new_[7973]_ ;
  assign \new_[6063]_  = \key_i[44]  ? \new_[7075]_  : \new_[1080]_ ;
  assign \new_[6064]_  = \key_i[51]  ? \new_[7075]_  : \new_[8057]_ ;
  assign \new_[6065]_  = \key_i[49]  ? \new_[7075]_  : \new_[8141]_ ;
  assign \new_[6066]_  = \key_i[60]  ? \new_[7075]_  : \new_[8028]_ ;
  assign \new_[6067]_  = \key_i[55]  ? \new_[7075]_  : \new_[8009]_ ;
  assign \new_[6068]_  = (~\new_[7660]_  | ~\key_i[57] ) & (~\new_[7075]_  | ~\new_[8124]_ );
  assign \new_[6069]_  = \key_i[54]  ? \new_[7075]_  : \new_[8122]_ ;
  assign \new_[6070]_  = (~\new_[7660]_  | ~\key_i[70] ) & (~\new_[7075]_  | ~\new_[2137]_ );
  assign \new_[6071]_  = ~\new_[8897]_  | ~\data_o[18] ;
  assign \new_[6072]_  = ~\new_[8931]_  | ~\new_[1313]_ ;
  assign \new_[6073]_  = \data_o[123]  ? \new_[8912]_  : \new_[1241]_ ;
  assign \new_[6074]_  = ~\new_[6364]_  | ~\new_[1208]_ ;
  assign n3605 = (~\new_[7605]_  & ~\new_[6808]_ ) | (~\new_[6511]_  & ~\new_[6636]_ );
  assign \new_[6076]_  = ~\new_[6657]_  | ~\new_[6648]_  | ~\new_[6498]_  | ~\new_[6487]_ ;
  assign \new_[6077]_  = ~\new_[6646]_  | ~\new_[6801]_  | ~\new_[6806]_  | ~\new_[6659]_ ;
  assign \new_[6078]_  = ~\new_[6655]_  | ~\new_[6647]_  | ~\new_[6658]_  | ~\new_[6661]_ ;
  assign \new_[6079]_  = \new_[6763]_  | \new_[5784]_ ;
  assign \new_[6080]_  = ~\new_[2426]_  | ~\new_[6763]_  | ~\new_[7884]_ ;
  assign \new_[6081]_  = \new_[6763]_  & \new_[2426]_ ;
  assign \new_[6082]_  = ~\new_[7932]_  | ~\new_[6763]_  | ~\new_[7884]_ ;
  assign \new_[6083]_  = ~\new_[6364]_  | ~\new_[1319]_ ;
  assign \new_[6084]_  = \new_[1146]_  | \new_[6355]_ ;
  assign \new_[6085]_  = ~\new_[6364]_  | ~\new_[1207]_ ;
  assign \new_[6086]_  = ~\new_[6364]_  | ~\new_[1461]_ ;
  assign \new_[6087]_  = \new_[1462]_  | \new_[6355]_ ;
  assign \new_[6088]_  = ~\new_[6364]_  | ~\new_[1206]_ ;
  assign \new_[6089]_  = ~\new_[6364]_  | ~\new_[1148]_ ;
  assign \new_[6090]_  = ~\new_[6364]_  | ~\new_[1106]_ ;
  assign \new_[6091]_  = ~\new_[6364]_  | ~\new_[1107]_ ;
  assign \new_[6092]_  = ~\new_[6356]_ ;
  assign \new_[6093]_  = ~\new_[6372]_  & (~\new_[6757]_  | ~\new_[7865]_ );
  assign \new_[6094]_  = ~\new_[6371]_  & (~\new_[6863]_  | ~\new_[7831]_ );
  assign \new_[6095]_  = ~\new_[6370]_  & (~\new_[6876]_  | ~\new_[7820]_ );
  assign \new_[6096]_  = ~\new_[6389]_  & (~\new_[6615]_  | ~\new_[7831]_ );
  assign \new_[6097]_  = ~\new_[6390]_  & (~\new_[6718]_  | ~\new_[7854]_ );
  assign \new_[6098]_  = \new_[6407]_  & \new_[8784]_ ;
  assign \new_[6099]_  = ~\new_[6197]_ ;
  assign \new_[6100]_  = ~\new_[6199]_ ;
  assign \new_[6101]_  = ~\new_[7892]_  | ~\new_[8991]_  | ~\new_[7859]_ ;
  assign \new_[6102]_  = ~\new_[7902]_  & (~\new_[6732]_  | ~\new_[6556]_ );
  assign \new_[6103]_  = ~\new_[8562]_  & (~\new_[6561]_  | ~\new_[6555]_ );
  assign \new_[6104]_  = ~\new_[7902]_  & (~\new_[6570]_  | ~\new_[6729]_ );
  assign \new_[6105]_  = ~\new_[7902]_  & (~\new_[6562]_  | ~\new_[6728]_ );
  assign \new_[6106]_  = ~\new_[6405]_  & ~\new_[8562]_ ;
  assign \new_[6107]_  = ~\new_[7902]_  & (~\new_[6557]_  | ~\new_[6554]_ );
  assign \new_[6108]_  = ~\new_[7902]_  & (~\new_[6558]_  | ~\new_[6439]_ );
  assign \new_[6109]_  = ~\new_[7902]_  & (~\new_[6559]_  | ~\new_[6441]_ );
  assign \new_[6110]_  = \new_[6400]_  & \new_[8558]_ ;
  assign \new_[6111]_  = ~\new_[7902]_  & (~\new_[6415]_  | ~\new_[6730]_ );
  assign \new_[6112]_  = \new_[6414]_  ? \new_[7662]_  : \new_[7926]_ ;
  assign \new_[6113]_  = \data_o[107]  ? \new_[8912]_  : \new_[1190]_ ;
  assign \new_[6114]_  = ~\new_[7819]_  | ~\new_[8991]_  | ~\new_[7835]_ ;
  assign \new_[6115]_  = ~\new_[8905]_  | ~\data_o[83] ;
  assign \new_[6116]_  = ~\new_[8911]_  | ~\data_o[34] ;
  assign \new_[6117]_  = ~\new_[8911]_  | ~\data_o[50] ;
  assign \new_[6118]_  = ~\new_[8914]_  | ~\data_o[58] ;
  assign \new_[6119]_  = ~\new_[8925]_  | ~\data_o[35] ;
  assign \new_[6120]_  = ~\new_[8925]_  | ~\data_o[26] ;
  assign \new_[6121]_  = ~\new_[8917]_  | ~\data_o[67] ;
  assign \new_[6122]_  = ~\new_[8911]_  | ~\data_o[42] ;
  assign \new_[6123]_  = ~\new_[8911]_  | ~\data_o[74] ;
  assign \new_[6124]_  = ~\new_[8919]_  | ~\data_o[51] ;
  assign \new_[6125]_  = ~\new_[8915]_  | ~\new_[1319]_ ;
  assign \new_[6126]_  = ~\new_[8924]_  | ~\new_[1381]_ ;
  assign \new_[6127]_  = ~\new_[8924]_  | ~\new_[1321]_ ;
  assign \new_[6128]_  = ~\new_[8904]_  | ~\new_[1245]_ ;
  assign \new_[6129]_  = ~\new_[8931]_  | ~\new_[1248]_ ;
  assign \new_[6130]_  = ~\new_[8931]_  | ~\new_[1385]_ ;
  assign \new_[6131]_  = ~\new_[8931]_  | ~\new_[1384]_ ;
  assign \new_[6132]_  = ~\new_[8915]_  | ~\new_[1314]_ ;
  assign \new_[6133]_  = (~\new_[7660]_  | ~\key_i[68] ) & (~\new_[7075]_  | ~\new_[2136]_ );
  assign \new_[6134]_  = (~\new_[7660]_  | ~\key_i[71] ) & (~\new_[7075]_  | ~\new_[2138]_ );
  assign \new_[6135]_  = \key_i[34]  ? \new_[7075]_  : \new_[7980]_ ;
  assign \new_[6136]_  = \key_i[42]  ? \new_[7075]_  : \new_[1118]_ ;
  assign \new_[6137]_  = \key_i[50]  ? \new_[7075]_  : \new_[8011]_ ;
  assign \new_[6138]_  = \key_i[33]  ? \new_[7075]_  : \new_[7968]_ ;
  assign \new_[6139]_  = \key_i[43]  ? \new_[7075]_  : \new_[1079]_ ;
  assign \new_[6140]_  = (~\new_[7660]_  | ~\key_i[69] ) & (~\new_[7075]_  | ~\new_[2095]_ );
  assign \new_[6141]_  = ~\new_[7075]_  | ~\new_[1084]_ ;
  assign \new_[6142]_  = ~\new_[7075]_  | ~\new_[1083]_ ;
  assign \new_[6143]_  = ~\new_[7075]_  | ~\new_[1082]_ ;
  assign \new_[6144]_  = ~\new_[7660]_  | ~\key_i[45] ;
  assign \new_[6145]_  = ~\new_[7660]_  | ~\key_i[47] ;
  assign \new_[6146]_  = ~\new_[7660]_  | ~\key_i[46] ;
  assign \new_[6147]_  = ~\new_[8469]_ ;
  assign \new_[6148]_  = \data_o[93]  ? \new_[8918]_  : \new_[1139]_ ;
  assign \new_[6149]_  = ~\new_[8925]_  | ~\data_o[43] ;
  assign \new_[6150]_  = ~\new_[8899]_  | ~\new_[1221]_ ;
  assign \new_[6151]_  = ~\new_[7116]_  | ~\new_[1100]_ ;
  assign \new_[6152]_  = \data_o[117]  ? \new_[8924]_  : \new_[1105]_ ;
  assign \new_[6153]_  = ~\new_[8924]_  | ~\new_[1216]_ ;
  assign n3615 = (~\new_[6668]_  & ~\new_[6636]_ ) | (~\new_[7867]_  & ~\new_[7427]_ );
  assign \new_[6155]_  = ~\new_[7116]_  | (~\new_[6636]_  & ~\new_[7934]_ );
  assign n3620 = (~\new_[6634]_  & ~\new_[6636]_ ) | (~\new_[7576]_  & ~\new_[7427]_ );
  assign n3610 = (~\new_[6578]_  & ~\new_[6636]_ ) | (~\new_[7830]_  & ~\new_[6954]_ );
  assign \new_[6158]_  = \new_[7931]_  ? \new_[9009]_  : \new_[8699]_ ;
  assign \new_[6159]_  = ~\new_[8469]_ ;
  assign \new_[6160]_  = ~\new_[8469]_ ;
  assign \new_[6161]_  = ~\new_[8469]_ ;
  assign \new_[6162]_  = ~\new_[8469]_ ;
  assign \new_[6163]_  = \new_[7580]_  ? \new_[7607]_  : \new_[6644]_ ;
  assign \new_[6164]_  = ~\new_[6789]_  | ~\new_[6800]_  | ~\new_[6664]_  | ~\new_[6662]_ ;
  assign \new_[6165]_  = ~\new_[6804]_  | ~\new_[6799]_  | ~\new_[6645]_  | ~\new_[6660]_ ;
  assign \new_[6166]_  = ~\new_[1103]_  | ~\new_[6453]_ ;
  assign \new_[6167]_  = ~\new_[1102]_  | ~\new_[6453]_ ;
  assign \new_[6168]_  = ~\new_[6354]_ ;
  assign \new_[6169]_  = ~\new_[6355]_ ;
  assign \new_[6170]_  = ~\new_[6359]_ ;
  assign \new_[6171]_  = \new_[7587]_  | \new_[8993]_ ;
  assign \new_[6172]_  = ~\new_[6364]_ ;
  assign \new_[6173]_  = ~\new_[6367]_ ;
  assign \new_[6174]_  = ~\new_[6459]_  & (~\new_[7026]_  | ~\new_[7865]_ );
  assign \new_[6175]_  = ~\new_[6458]_  & (~\new_[6830]_  | ~\new_[7854]_ );
  assign \new_[6176]_  = ~\new_[6544]_  | (~\new_[6719]_  & ~\new_[7817]_ );
  assign \new_[6177]_  = ~\new_[6545]_  | (~\new_[6875]_  & ~\new_[7817]_ );
  assign \new_[6178]_  = ~\new_[6541]_  | ~\new_[6536]_ ;
  assign \new_[6179]_  = (~\new_[6721]_  | ~\new_[7865]_ ) & (~\new_[7010]_  | ~\new_[7831]_ );
  assign \new_[6180]_  = ~\new_[6543]_  | (~\new_[6720]_  & ~\new_[7827]_ );
  assign \new_[6181]_  = ~\new_[6534]_  & (~\new_[6758]_  | ~\new_[7831]_ );
  assign \new_[6182]_  = ~\new_[6532]_  & (~\new_[6871]_  | ~\new_[7818]_ );
  assign \new_[6183]_  = ~\new_[6533]_  & (~\new_[6861]_  | ~\new_[7818]_ );
  assign \new_[6184]_  = ~\new_[6535]_  & (~\new_[6931]_  | ~\new_[7818]_ );
  assign \new_[6185]_  = ~\new_[6542]_  & (~\new_[6920]_  | ~\new_[7818]_ );
  assign \new_[6186]_  = \new_[7562]_  ? \new_[8994]_  : \new_[1981]_ ;
  assign \new_[6187]_  = \new_[6548]_  & \new_[8784]_ ;
  assign \new_[6188]_  = ~\new_[7116]_  | ~\new_[1097]_ ;
  assign \new_[6189]_  = ~\new_[7116]_  | ~\new_[1096]_ ;
  assign \new_[6190]_  = ~\new_[7116]_  | ~\new_[1099]_ ;
  assign \new_[6191]_  = ~\new_[7116]_  | ~\new_[1095]_ ;
  assign \new_[6192]_  = ~\new_[7116]_  | ~\new_[1094]_ ;
  assign \new_[6193]_  = ~\new_[7116]_  | ~\new_[1098]_ ;
  assign \new_[6194]_  = ~\new_[7116]_  | ~\new_[1101]_ ;
  assign \new_[6195]_  = \new_[6549]_  & \new_[8784]_ ;
  assign \new_[6196]_  = \new_[6550]_  & \new_[8784]_ ;
  assign \new_[6197]_  = ~\new_[8993]_  | ~\new_[7918]_ ;
  assign \new_[6198]_  = \new_[8993]_  | \new_[7923]_ ;
  assign \new_[6199]_  = ~\new_[8993]_  | ~\new_[7916]_ ;
  assign \new_[6200]_  = ~\new_[7902]_  & (~\new_[6731]_  | ~\new_[6724]_ );
  assign \new_[6201]_  = ~\new_[7902]_  & (~\new_[6750]_  | ~\new_[6613]_ );
  assign \new_[6202]_  = (~\new_[6733]_  | ~\new_[7607]_ ) & (~\new_[7848]_  | ~\new_[7662]_ );
  assign \new_[6203]_  = \new_[6900]_  | \new_[6440]_ ;
  assign \new_[6204]_  = \data_o[94]  ? \new_[8918]_  : \new_[1137]_ ;
  assign \new_[6205]_  = \data_o[126]  ? \new_[8918]_  : \new_[1135]_ ;
  assign \new_[6206]_  = \data_o[110]  ? \new_[8918]_  : \new_[1095]_ ;
  assign \new_[6207]_  = \data_o[101]  ? \new_[8904]_  : \new_[1103]_ ;
  assign \new_[6208]_  = \data_o[125]  ? \new_[8900]_  : \new_[1134]_ ;
  assign \new_[6209]_  = \data_o[14]  ? \new_[8900]_  : \new_[1097]_ ;
  assign \new_[6210]_  = ~\new_[8925]_  | ~\data_o[59] ;
  assign \new_[6211]_  = ~\new_[8924]_  | ~\new_[1197]_ ;
  assign \new_[6212]_  = ~\new_[8924]_  | ~\new_[1211]_ ;
  assign \new_[6213]_  = ~\new_[8946]_  | ~\new_[1247]_ ;
  assign \new_[6214]_  = ~\new_[8946]_  | ~\new_[1237]_ ;
  assign \new_[6215]_  = \key_i[73]  ? \new_[7075]_  : \new_[8119]_ ;
  assign \new_[6216]_  = ~\new_[7660]_  | ~\key_i[72] ;
  assign \new_[6217]_  = \data_i[61]  ? \new_[6777]_  : \new_[6631]_ ;
  assign \new_[6218]_  = \data_o[15]  ? \new_[8918]_  : \new_[1195]_ ;
  assign \new_[6219]_  = \data_o[13]  ? \new_[8918]_  : \new_[1096]_ ;
  assign \new_[6220]_  = (~\new_[6874]_  | ~\new_[7865]_ ) & (~\new_[7024]_  | ~\new_[7820]_ );
  assign \new_[6221]_  = ~\new_[8933]_  | ~\data_o[29] ;
  assign \new_[6222]_  = ~\new_[6437]_ ;
  assign \new_[6223]_  = \new_[6621]_  | \new_[6633]_ ;
  assign \new_[6224]_  = ~\new_[8946]_  | ~\new_[1098]_ ;
  assign \new_[6225]_  = \data_o[6]  ? \new_[8900]_  : \new_[1113]_ ;
  assign \new_[6226]_  = \new_[6901]_  | \new_[6725]_ ;
  assign \new_[6227]_  = \data_i[41]  ? \new_[6777]_  : \new_[6656]_ ;
  assign \new_[6228]_  = \data_i[62]  ? \new_[6795]_  : \new_[6594]_ ;
  assign \new_[6229]_  = \data_i[19]  ? \new_[6794]_  : \new_[2935]_ ;
  assign \new_[6230]_  = \data_i[54]  ? \new_[6796]_  : \new_[6626]_ ;
  assign \new_[6231]_  = \data_i[112]  ? \new_[6778]_  : \new_[6423]_ ;
  assign \new_[6232]_  = \data_i[1]  ? \new_[6778]_  : \new_[3105]_ ;
  assign \new_[6233]_  = \data_i[101]  ? \new_[6796]_  : \new_[6606]_ ;
  assign \new_[6234]_  = \data_i[117]  ? \new_[6752]_  : \new_[6694]_ ;
  assign \new_[6235]_  = \data_i[63]  ? \new_[6777]_  : \new_[6632]_ ;
  assign \new_[6236]_  = \data_i[66]  ? \new_[6752]_  : \new_[6618]_ ;
  assign \new_[6237]_  = \data_i[30]  ? \new_[6795]_  : \new_[3386]_ ;
  assign \new_[6238]_  = \data_i[20]  ? \new_[6794]_  : \new_[2756]_ ;
  assign \new_[6239]_  = \data_i[67]  ? \new_[6776]_  : \new_[6425]_ ;
  assign \new_[6240]_  = \data_i[113]  ? \new_[6794]_  : \new_[6652]_ ;
  assign \new_[6241]_  = \data_i[120]  ? \new_[6794]_  : \new_[6639]_ ;
  assign \new_[6242]_  = \data_i[68]  ? \new_[6796]_  : \new_[6605]_ ;
  assign \new_[6243]_  = \data_i[21]  ? \new_[6795]_  : \new_[3383]_ ;
  assign \new_[6244]_  = \data_i[69]  ? \new_[6752]_  : \new_[6442]_ ;
  assign \new_[6245]_  = \data_i[22]  ? \new_[6752]_  : \new_[3385]_ ;
  assign \new_[6246]_  = \data_i[70]  ? \new_[6793]_  : \new_[6426]_ ;
  assign \new_[6247]_  = \data_i[81]  ? \new_[6776]_  : \new_[6619]_ ;
  assign \new_[6248]_  = \data_i[114]  ? \new_[6776]_  : \new_[6704]_ ;
  assign \new_[6249]_  = \data_i[71]  ? \new_[6794]_  : \new_[6446]_ ;
  assign \new_[6250]_  = \data_i[23]  ? \new_[6752]_  : \new_[3857]_ ;
  assign \new_[6251]_  = \data_i[72]  ? \new_[6778]_  : \new_[6432]_ ;
  assign \new_[6252]_  = \data_i[102]  ? \new_[6793]_  : \new_[6419]_ ;
  assign \new_[6253]_  = \data_i[73]  ? \new_[6778]_  : \new_[6716]_ ;
  assign \new_[6254]_  = \data_i[24]  ? \new_[6793]_  : \new_[3443]_ ;
  assign \new_[6255]_  = \data_i[74]  ? \new_[6777]_  : \new_[6573]_ ;
  assign \new_[6256]_  = \data_i[33]  ? \new_[6776]_  : \new_[6444]_ ;
  assign \new_[6257]_  = \data_i[115]  ? \new_[6796]_  : \new_[6596]_ ;
  assign \new_[6258]_  = \data_i[75]  ? \new_[6777]_  : \new_[6630]_ ;
  assign \new_[6259]_  = \data_i[25]  ? \new_[6796]_  : \new_[3106]_ ;
  assign \new_[6260]_  = \data_i[76]  ? \new_[6793]_  : \new_[6581]_ ;
  assign \new_[6261]_  = \data_i[35]  ? \new_[6795]_  : \new_[6749]_ ;
  assign \new_[6262]_  = \data_i[77]  ? \new_[6793]_  : \new_[6450]_ ;
  assign \new_[6263]_  = \data_i[83]  ? \new_[6776]_  : \new_[6600]_ ;
  assign \new_[6264]_  = \data_i[26]  ? \new_[6776]_  : \new_[3107]_ ;
  assign \new_[6265]_  = \data_i[116]  ? \new_[6794]_  : \new_[6547]_ ;
  assign \new_[6266]_  = \data_i[79]  ? \new_[6777]_  : \new_[6748]_ ;
  assign \new_[6267]_  = \data_i[27]  ? \new_[6796]_  : \new_[2932]_ ;
  assign \new_[6268]_  = \data_i[103]  ? \new_[6795]_  : \new_[6586]_ ;
  assign \new_[6269]_  = \data_i[65]  ? \new_[6793]_  : \new_[6445]_ ;
  assign \new_[6270]_  = \data_i[85]  ? \new_[6752]_  : \new_[6427]_ ;
  assign \new_[6271]_  = \data_i[118]  ? \new_[6796]_  : \new_[6607]_ ;
  assign \new_[6272]_  = \data_i[78]  ? \new_[6795]_  : \new_[6451]_ ;
  assign \new_[6273]_  = \data_i[86]  ? \new_[6778]_  : \new_[6566]_ ;
  assign \new_[6274]_  = \data_i[89]  ? \new_[6778]_  : \new_[6569]_ ;
  assign \new_[6275]_  = \data_i[87]  ? \new_[6794]_  : \new_[6614]_ ;
  assign \new_[6276]_  = \data_i[104]  ? \new_[6777]_  : \new_[6416]_ ;
  assign \new_[6277]_  = \data_i[88]  ? \new_[6778]_  : \new_[6568]_ ;
  assign \new_[6278]_  = \data_i[31]  ? \new_[6795]_  : \new_[3863]_ ;
  assign \new_[6279]_  = \data_i[28]  ? \new_[6795]_  : \new_[2757]_ ;
  assign \new_[6280]_  = (~\new_[6768]_  | ~\new_[7854]_ ) & (~\new_[6869]_  | ~\new_[7865]_ );
  assign \new_[6281]_  = \data_i[119]  ? \new_[6776]_  : \new_[6589]_ ;
  assign \new_[6282]_  = \data_i[8]  ? \new_[6793]_  : \new_[3377]_ ;
  assign \new_[6283]_  = \data_i[32]  ? \new_[6794]_  : \new_[6629]_ ;
  assign \new_[6284]_  = \data_i[90]  ? \new_[6777]_  : \new_[6572]_ ;
  assign \new_[6285]_  = \data_i[105]  ? \new_[6777]_  : \new_[6420]_ ;
  assign \new_[6286]_  = \data_i[92]  ? \new_[6777]_  : \new_[6666]_ ;
  assign \new_[6287]_  = \data_i[11]  ? \new_[6795]_  : \new_[2934]_ ;
  assign \new_[6288]_  = \data_i[34]  ? \new_[6796]_  : \new_[6643]_ ;
  assign \new_[6289]_  = \data_i[94]  ? \new_[6777]_  : \new_[6625]_ ;
  assign \new_[6290]_  = \data_i[2]  ? \new_[6794]_  : \new_[3109]_ ;
  assign \new_[6291]_  = \data_i[95]  ? \new_[6794]_  : \new_[6746]_ ;
  assign \new_[6292]_  = \data_i[29]  ? \new_[6796]_  : \new_[3514]_ ;
  assign \new_[6293]_  = \data_i[91]  ? \new_[6793]_  : \new_[6438]_ ;
  assign \new_[6294]_  = \data_i[96]  ? \new_[6776]_  : \new_[6595]_ ;
  assign \new_[6295]_  = \data_i[97]  ? \new_[6796]_  : \new_[6579]_ ;
  assign \new_[6296]_  = \data_i[36]  ? \new_[6794]_  : \new_[6591]_ ;
  assign \new_[6297]_  = \data_i[98]  ? \new_[6794]_  : \new_[6428]_ ;
  assign \new_[6298]_  = \data_i[99]  ? \new_[6796]_  : \new_[6430]_ ;
  assign \new_[6299]_  = \data_i[37]  ? \new_[6752]_  : \new_[6584]_ ;
  assign \new_[6300]_  = \data_i[9]  ? \new_[6793]_  : \new_[3108]_ ;
  assign \new_[6301]_  = \data_i[121]  ? \new_[6776]_  : \new_[6663]_ ;
  assign \new_[6302]_  = \data_i[80]  ? \new_[6778]_  : \new_[6598]_ ;
  assign \new_[6303]_  = \data_i[64]  ? \new_[6752]_  : \new_[6495]_ ;
  assign \new_[6304]_  = \data_i[6]  ? \new_[6776]_  : \new_[3406]_ ;
  assign \new_[6305]_  = \data_i[39]  ? \new_[6794]_  : \new_[6592]_ ;
  assign \new_[6306]_  = \data_i[106]  ? \new_[6776]_  : \new_[6449]_ ;
  assign \new_[6307]_  = \data_i[122]  ? \new_[6777]_  : \new_[6452]_ ;
  assign \new_[6308]_  = \data_i[3]  ? \new_[6777]_  : \new_[2870]_ ;
  assign \new_[6309]_  = \data_i[13]  ? \new_[6752]_  : \new_[3382]_ ;
  assign \new_[6310]_  = \data_i[123]  ? \new_[6752]_  : \new_[6599]_ ;
  assign \new_[6311]_  = \data_i[107]  ? \new_[6752]_  : \new_[6620]_ ;
  assign \new_[6312]_  = \data_i[42]  ? \new_[6752]_  : \new_[6624]_ ;
  assign \new_[6313]_  = \data_i[127]  ? \new_[6795]_  : \new_[6723]_ ;
  assign \new_[6314]_  = \data_i[124]  ? \new_[6778]_  : \new_[6628]_ ;
  assign \new_[6315]_  = \data_i[0]  ? \new_[6778]_  : \new_[3410]_ ;
  assign \new_[6316]_  = \data_i[44]  ? \new_[6776]_  : \new_[6623]_ ;
  assign \new_[6317]_  = \data_i[125]  ? \new_[6793]_  : \new_[6590]_ ;
  assign \new_[6318]_  = \data_i[45]  ? \new_[6793]_  : \new_[6424]_ ;
  assign \new_[6319]_  = \data_i[43]  ? \new_[6795]_  : \new_[6580]_ ;
  assign \new_[6320]_  = \data_i[47]  ? \new_[6795]_  : \new_[6575]_ ;
  assign \new_[6321]_  = \data_i[108]  ? \new_[6778]_  : \new_[6421]_ ;
  assign \new_[6322]_  = \data_i[46]  ? \new_[6777]_  : \new_[6597]_ ;
  assign \new_[6323]_  = \data_i[49]  ? \new_[6778]_  : \new_[6546]_ ;
  assign \new_[6324]_  = \data_i[126]  ? \new_[6777]_  : \new_[6571]_ ;
  assign \new_[6325]_  = \data_i[109]  ? \new_[6777]_  : \new_[6587]_ ;
  assign \new_[6326]_  = \data_i[12]  ? \new_[6778]_  : \new_[2755]_ ;
  assign \new_[6327]_  = \data_i[50]  ? \new_[6794]_  : \new_[6627]_ ;
  assign \new_[6328]_  = \data_i[51]  ? \new_[6752]_  : \new_[6616]_ ;
  assign \new_[6329]_  = \data_i[52]  ? \new_[6752]_  : \new_[6609]_ ;
  assign \new_[6330]_  = \data_i[10]  ? \new_[6778]_  : \new_[3257]_ ;
  assign \new_[6331]_  = \data_i[82]  ? \new_[6794]_  : \new_[6429]_ ;
  assign \new_[6332]_  = \data_i[53]  ? \new_[6793]_  : \new_[6588]_ ;
  assign \new_[6333]_  = \data_i[48]  ? \new_[6796]_  : \new_[6433]_ ;
  assign \new_[6334]_  = \data_i[14]  ? \new_[6795]_  : \new_[3409]_ ;
  assign \new_[6335]_  = \data_i[4]  ? \new_[6795]_  : \new_[2758]_ ;
  assign \new_[6336]_  = \data_i[40]  ? \new_[6776]_  : \new_[6640]_ ;
  assign \new_[6337]_  = \data_i[55]  ? \new_[6796]_  : \new_[6593]_ ;
  assign \new_[6338]_  = \data_i[15]  ? \new_[6793]_  : \new_[3885]_ ;
  assign \new_[6339]_  = \data_i[38]  ? \new_[6795]_  : \new_[6714]_ ;
  assign \new_[6340]_  = \data_i[56]  ? \new_[6793]_  : \new_[6574]_ ;
  assign \new_[6341]_  = \data_i[110]  ? \new_[6796]_  : \new_[6422]_ ;
  assign \new_[6342]_  = \data_i[84]  ? \new_[6752]_  : \new_[6585]_ ;
  assign \new_[6343]_  = \data_i[57]  ? \new_[6776]_  : \new_[6443]_ ;
  assign \new_[6344]_  = \data_i[16]  ? \new_[6796]_  : \new_[3387]_ ;
  assign \new_[6345]_  = \data_i[58]  ? \new_[6795]_  : \new_[6601]_ ;
  assign \new_[6346]_  = \data_i[7]  ? \new_[6776]_  : \new_[3846]_ ;
  assign \new_[6347]_  = \data_i[59]  ? \new_[6793]_  : \new_[6610]_ ;
  assign \new_[6348]_  = \data_i[17]  ? \new_[6776]_  : \new_[3103]_ ;
  assign \new_[6349]_  = \data_i[5]  ? \new_[6778]_  : \new_[3515]_ ;
  assign \new_[6350]_  = \data_i[100]  ? \new_[6796]_  : \new_[6751]_ ;
  assign \new_[6351]_  = \data_i[111]  ? \new_[6793]_  : \new_[6641]_ ;
  assign \new_[6352]_  = \data_i[60]  ? \new_[6794]_  : \new_[6702]_ ;
  assign \new_[6353]_  = \data_i[18]  ? \new_[6752]_  : \new_[3104]_ ;
  assign \new_[6354]_  = ~\new_[6654]_  & ~\new_[7117]_ ;
  assign \new_[6355]_  = ~\new_[7117]_  & ~\new_[6650]_ ;
  assign \new_[6356]_  = ~\new_[6650]_  & ~\new_[6790]_ ;
  assign \new_[6357]_  = \new_[6651]_  | \new_[6790]_ ;
  assign \new_[6358]_  = \new_[6651]_  | \new_[6649]_ ;
  assign \new_[6359]_  = ~\new_[6649]_  & ~\new_[6650]_ ;
  assign \new_[6360]_  = ~\new_[6454]_ ;
  assign \new_[6361]_  = \new_[6654]_  | \new_[6790]_ ;
  assign \new_[6362]_  = ~\new_[6417]_ ;
  assign \new_[6363]_  = \new_[6654]_  | \new_[6649]_ ;
  assign \new_[6364]_  = \new_[7117]_  | \new_[6651]_ ;
  assign \new_[6365]_  = ~\new_[6436]_ ;
  assign \new_[6366]_  = ~\new_[6435]_ ;
  assign \new_[6367]_  = ~\new_[7117]_  & ~\new_[6653]_ ;
  assign \new_[6368]_  = ~\new_[6434]_ ;
  assign \new_[6369]_  = ~\new_[6712]_  | (~\new_[6754]_  & ~\new_[7817]_ );
  assign \new_[6370]_  = ~\new_[7817]_  & (~\new_[6889]_  | ~\new_[6887]_ );
  assign \new_[6371]_  = ~\new_[7817]_  & (~\new_[6888]_  | ~\new_[6886]_ );
  assign \new_[6372]_  = ~\new_[7817]_  & (~\new_[6892]_  | ~\new_[6884]_ );
  assign \new_[6373]_  = (~\new_[6772]_  | ~\new_[7818]_ ) & (~\new_[6865]_  | ~\new_[7832]_ );
  assign \new_[6374]_  = (~\new_[6862]_  | ~\new_[7832]_ ) & (~\new_[6870]_  | ~\new_[7818]_ );
  assign \new_[6375]_  = (~\new_[6867]_  | ~\new_[7831]_ ) & (~\new_[7022]_  | ~\new_[7865]_ );
  assign \new_[6376]_  = ~\new_[6494]_ ;
  assign \new_[6377]_  = (~\new_[6882]_  | ~\new_[7865]_ ) & (~\new_[7006]_  | ~\new_[7832]_ );
  assign \new_[6378]_  = (~\new_[6883]_  | ~\new_[7831]_ ) & (~\new_[6880]_  | ~\new_[7854]_ );
  assign \new_[6379]_  = (~\new_[6873]_  | ~\new_[7820]_ ) & (~\new_[6929]_  | ~\new_[7832]_ );
  assign \new_[6380]_  = (~\new_[6860]_  | ~\new_[7820]_ ) & (~\new_[7021]_  | ~\new_[7832]_ );
  assign \new_[6381]_  = (~\new_[6877]_  | ~\new_[7818]_ ) & (~\new_[7014]_  | ~\new_[7854]_ );
  assign \new_[6382]_  = (~\new_[6866]_  | ~\new_[7838]_ ) & (~\new_[6921]_  | ~\new_[7861]_ );
  assign \new_[6383]_  = ~\new_[6701]_  & (~\new_[1950]_  | ~\new_[8994]_ );
  assign \new_[6384]_  = \new_[6802]_  & \new_[6667]_ ;
  assign \new_[6385]_  = (~\new_[7561]_  & ~\new_[8989]_ ) | (~\new_[7961]_  & ~\new_[8996]_ );
  assign \new_[6386]_  = \new_[6814]_  & \new_[6708]_ ;
  assign \new_[6387]_  = ~\new_[6709]_  & (~\new_[1964]_  | ~\new_[8989]_ );
  assign \new_[6388]_  = \new_[6820]_  & \new_[6713]_ ;
  assign \new_[6389]_  = ~\new_[7827]_  & (~\new_[6890]_  | ~\new_[6761]_ );
  assign \new_[6390]_  = ~\new_[7827]_  & (~\new_[6767]_  | ~\new_[6885]_ );
  assign \new_[6391]_  = \new_[6717]_  & \new_[8558]_ ;
  assign \new_[6392]_  = \new_[6722]_  & \new_[7893]_ ;
  assign \new_[6393]_  = ~\new_[6715]_  & (~\new_[7648]_  | ~\new_[7921]_ );
  assign \new_[6394]_  = ~\new_[6453]_ ;
  assign \new_[6395]_  = \data_o[86]  ? \new_[8941]_  : \new_[1117]_ ;
  assign \new_[6396]_  = \new_[6576]_  | \new_[6727]_ ;
  assign \new_[6397]_  = \data_o[95]  ? \new_[8931]_  : \new_[1250]_ ;
  assign \new_[6398]_  = \data_o[5]  ? \new_[8924]_  : \new_[1112]_ ;
  assign \new_[6399]_  = \data_o[87]  ? \new_[8918]_  : \new_[1222]_ ;
  assign \new_[6400]_  = \data_o[70]  ? \new_[8896]_  : \new_[1114]_ ;
  assign \new_[6401]_  = \data_o[21]  ? \new_[8924]_  : \new_[1106]_ ;
  assign \new_[6402]_  = \data_o[85]  ? \new_[8941]_  : \new_[1116]_ ;
  assign \new_[6403]_  = \data_o[109]  ? \new_[8900]_  : \new_[1094]_ ;
  assign \new_[6404]_  = \new_[6747]_  | \new_[6726]_ ;
  assign \new_[6405]_  = (~\new_[8917]_  | ~\data_o[78] ) & (~\new_[8941]_  | ~\new_[1101]_ );
  assign \new_[6406]_  = \new_[6893]_  | \new_[6611]_ ;
  assign \new_[6407]_  = \data_o[22]  ? \new_[8896]_  : \new_[1107]_ ;
  assign \new_[6408]_  = ~\new_[8925]_  | ~\data_o[45] ;
  assign \new_[6409]_  = ~\new_[8933]_  | ~\data_o[77] ;
  assign \new_[6410]_  = ~\new_[8897]_  | ~\data_o[53] ;
  assign \new_[6411]_  = ~\new_[8918]_  | ~\new_[1110]_ ;
  assign \new_[6412]_  = (~\new_[6864]_  | ~\new_[7831]_ ) & (~\new_[6868]_  | ~\new_[7854]_ );
  assign \new_[6413]_  = ~\new_[8918]_  | ~\new_[1100]_ ;
  assign \new_[6414]_  = \new_[7926]_  ^ \new_[7648]_ ;
  assign \new_[6415]_  = ~\new_[8941]_  | ~\new_[1187]_ ;
  assign \new_[6416]_  = \\mix1_data_o_reg_reg[104] ;
  assign \new_[6417]_  = ~\new_[6949]_  | ~\new_[6791]_ ;
  assign \new_[6418]_  = ~\new_[7607]_  | ~\new_[7406]_  | ~\new_[7648]_ ;
  assign \new_[6419]_  = \\mix1_data_o_reg_reg[102] ;
  assign \new_[6420]_  = \\mix1_data_o_reg_reg[105] ;
  assign \new_[6421]_  = \\mix1_data_o_reg_reg[108] ;
  assign \new_[6422]_  = \\mix1_data_o_reg_reg[110] ;
  assign \new_[6423]_  = \\mix1_data_o_reg_reg[112] ;
  assign \new_[6424]_  = \\mix1_data_o_reg_reg[45] ;
  assign \new_[6425]_  = \\mix1_data_o_reg_reg[67] ;
  assign \new_[6426]_  = \\mix1_data_o_reg_reg[70] ;
  assign \new_[6427]_  = \\mix1_data_o_reg_reg[85] ;
  assign \new_[6428]_  = \\mix1_data_o_reg_reg[98] ;
  assign \new_[6429]_  = \\mix1_data_o_reg_reg[82] ;
  assign \new_[6430]_  = \\mix1_data_o_reg_reg[99] ;
  assign \new_[6431]_  = ~\new_[8101]_  | ~\new_[6954]_ ;
  assign \new_[6432]_  = \\mix1_data_o_reg_reg[72] ;
  assign \new_[6433]_  = \\mix1_data_o_reg_reg[48] ;
  assign \new_[6434]_  = ~\new_[6798]_  | ~\new_[6949]_ ;
  assign \new_[6435]_  = ~\new_[6792]_  | ~\new_[6949]_ ;
  assign \new_[6436]_  = ~\new_[6797]_  | ~\new_[6950]_ ;
  assign \new_[6437]_  = (~\new_[6915]_  | ~\new_[7832]_ ) & (~\new_[7016]_  | ~\new_[7820]_ );
  assign \new_[6438]_  = \\mix1_data_o_reg_reg[91] ;
  assign \new_[6439]_  = ~\new_[8897]_  | ~\data_o[37] ;
  assign \new_[6440]_  = \new_[8919]_  & \data_o[102] ;
  assign \new_[6441]_  = ~\new_[8897]_  | ~\data_o[61] ;
  assign \new_[6442]_  = \\mix1_data_o_reg_reg[69] ;
  assign \new_[6443]_  = \\mix1_data_o_reg_reg[57] ;
  assign \new_[6444]_  = \\mix1_data_o_reg_reg[33] ;
  assign \new_[6445]_  = \\mix1_data_o_reg_reg[65] ;
  assign \new_[6446]_  = \\mix1_data_o_reg_reg[71] ;
  assign \new_[6447]_  = \new_[7116]_  & \new_[1111]_ ;
  assign \new_[6448]_  = \\mix1_data_o_reg_reg[93] ;
  assign \new_[6449]_  = \\mix1_data_o_reg_reg[106] ;
  assign \new_[6450]_  = \\mix1_data_o_reg_reg[77] ;
  assign \new_[6451]_  = \\mix1_data_o_reg_reg[78] ;
  assign \new_[6452]_  = \\mix1_data_o_reg_reg[122] ;
  assign \new_[6453]_  = ~\new_[6797]_  | ~\new_[6949]_ ;
  assign \new_[6454]_  = ~\new_[6827]_  | ~\new_[6797]_ ;
  assign \new_[6455]_  = (~\new_[7036]_  | ~\new_[7836]_ ) & (~\new_[7125]_  | ~\new_[7833]_ );
  assign \new_[6456]_  = (~\new_[7017]_  | ~\new_[7836]_ ) & (~\new_[7107]_  | ~\new_[7833]_ );
  assign \new_[6457]_  = (~\new_[6934]_  | ~\new_[7833]_ ) & (~\new_[7020]_  | ~\new_[7866]_ );
  assign \new_[6458]_  = ~\new_[7817]_  & (~\new_[6912]_  | ~\new_[7030]_ );
  assign \new_[6459]_  = ~\new_[7817]_  & (~\new_[7139]_  | ~\new_[7029]_ );
  assign \new_[6460]_  = ~\new_[1137]_  | ~\new_[6954]_ ;
  assign \new_[6461]_  = ~\new_[1250]_  | ~\new_[6954]_ ;
  assign \new_[6462]_  = ~\new_[1139]_  | ~\new_[6954]_ ;
  assign \new_[6463]_  = ~\new_[1134]_  | ~\new_[6954]_ ;
  assign \new_[6464]_  = ~\new_[1241]_  | ~\new_[6954]_ ;
  assign \new_[6465]_  = ~\new_[1385]_  | ~\new_[6954]_ ;
  assign \new_[6466]_  = ~\new_[1386]_  | ~\new_[6954]_ ;
  assign \new_[6467]_  = ~\new_[1251]_  | ~\new_[6954]_ ;
  assign \new_[6468]_  = ~\new_[1224]_  | ~\new_[6954]_ ;
  assign \new_[6469]_  = ~\new_[1186]_  | ~\new_[6954]_ ;
  assign \new_[6470]_  = ~\new_[8053]_  | ~\new_[6954]_ ;
  assign \new_[6471]_  = ~\new_[1223]_  | ~\new_[6954]_ ;
  assign \new_[6472]_  = ~\new_[1135]_  | ~\new_[6954]_ ;
  assign \new_[6473]_  = ~\new_[1383]_  | ~\new_[6954]_ ;
  assign \new_[6474]_  = ~\new_[1136]_  | ~\new_[6954]_ ;
  assign \new_[6475]_  = ~\new_[1187]_  | ~\new_[6954]_ ;
  assign \new_[6476]_  = ~\new_[1246]_  | ~\new_[6954]_ ;
  assign \new_[6477]_  = ~\new_[1138]_  | ~\new_[6954]_ ;
  assign \new_[6478]_  = ~\new_[1245]_  | ~\new_[6954]_ ;
  assign \new_[6479]_  = ~\new_[1249]_  | ~\new_[6954]_ ;
  assign \new_[6480]_  = ~\new_[8020]_  | ~\new_[6954]_ ;
  assign \new_[6481]_  = ~\new_[1247]_  | ~\new_[6954]_ ;
  assign \new_[6482]_  = ~\new_[1244]_  | ~\new_[6954]_ ;
  assign \new_[6483]_  = ~\new_[1252]_  | ~\new_[6954]_ ;
  assign \new_[6484]_  = ~\new_[1248]_  | ~\new_[6954]_ ;
  assign \new_[6485]_  = ~\new_[7939]_  | ~\new_[6954]_ ;
  assign \new_[6486]_  = ~\new_[1226]_  | ~\new_[6954]_ ;
  assign \new_[6487]_  = (~\new_[6932]_  | ~\new_[7815]_ ) & (~\new_[7275]_  | ~\new_[7838]_ );
  assign \new_[6488]_  = (~\new_[7023]_  | ~\new_[7815]_ ) & (~\new_[7009]_  | ~\new_[7864]_ );
  assign \new_[6489]_  = (~\new_[7019]_  | ~\new_[7815]_ ) & (~\new_[7104]_  | ~\new_[7838]_ );
  assign \new_[6490]_  = (~\new_[7013]_  | ~\new_[7815]_ ) & (~\new_[7129]_  | ~\new_[7866]_ );
  assign \new_[6491]_  = (~\new_[7018]_  | ~\new_[7852]_ ) & (~\new_[7130]_  | ~\new_[7861]_ );
  assign \new_[6492]_  = (~\new_[7056]_  | ~\new_[7831]_ ) & (~\new_[7015]_  | ~\new_[7854]_ );
  assign \new_[6493]_  = (~\new_[7025]_  | ~\new_[7836]_ ) & (~\new_[6933]_  | ~\new_[7852]_ );
  assign \new_[6494]_  = (~\new_[7008]_  | ~\new_[7820]_ ) & (~\new_[7106]_  | ~\new_[7832]_ );
  assign \new_[6495]_  = \\mix1_data_o_reg_reg[64] ;
  assign \new_[6496]_  = (~\new_[7083]_  | ~\new_[7852]_ ) & (~\new_[7127]_  | ~\new_[7864]_ );
  assign \new_[6497]_  = (~\new_[6935]_  | ~\new_[7866]_ ) & (~\new_[7281]_  | ~\new_[7864]_ );
  assign \new_[6498]_  = (~\new_[7007]_  | ~\new_[7836]_ ) & (~\new_[7126]_  | ~\new_[7864]_ );
  assign \new_[6499]_  = (~\new_[7596]_  & ~\new_[8989]_ ) | (~\new_[8106]_  & ~\new_[8996]_ );
  assign \new_[6500]_  = (~\new_[7642]_  & ~\new_[8994]_ ) | (~\new_[7953]_  & ~\new_[8996]_ );
  assign \new_[6501]_  = (~\new_[7650]_  & ~\new_[8988]_ ) | (~\new_[8148]_  & ~\new_[8987]_ );
  assign \new_[6502]_  = (~\new_[7661]_  & ~\new_[8989]_ ) | (~\new_[8006]_  & ~\new_[8990]_ );
  assign \new_[6503]_  = (~\new_[7612]_  & ~\new_[8989]_ ) | (~\new_[8051]_  & ~\new_[8987]_ );
  assign \new_[6504]_  = (~\new_[8884]_  & ~\new_[8994]_ ) | (~\new_[8018]_  & ~\new_[8998]_ );
  assign \new_[6505]_  = \new_[7613]_  ? \new_[8994]_  : \new_[1063]_ ;
  assign \new_[6506]_  = (~\new_[7594]_  & ~\new_[8994]_ ) | (~\new_[7994]_  & ~\new_[8996]_ );
  assign \new_[6507]_  = (~\new_[7641]_  & ~\new_[8989]_ ) | (~\new_[7937]_  & ~\new_[8987]_ );
  assign \new_[6508]_  = (~\new_[7652]_  & ~\new_[8989]_ ) | (~\new_[7952]_  & ~\new_[8987]_ );
  assign \new_[6509]_  = (~\new_[7611]_  & ~\new_[8989]_ ) | (~\new_[7970]_  & ~\new_[8995]_ );
  assign \new_[6510]_  = ~\new_[7116]_  | ~\new_[1142]_ ;
  assign \new_[6511]_  = ~\new_[7116]_  | ~\new_[5960]_ ;
  assign \new_[6512]_  = ~\new_[7116]_  | ~\new_[1144]_ ;
  assign \new_[6513]_  = \new_[7116]_  & \new_[1102]_ ;
  assign \new_[6514]_  = ~\new_[7116]_  | ~\new_[1459]_ ;
  assign \new_[6515]_  = ~\new_[7116]_  | ~\new_[1460]_ ;
  assign \new_[6516]_  = \new_[7116]_  & \new_[1105]_ ;
  assign \new_[6517]_  = \new_[7116]_  & \new_[1116]_ ;
  assign \new_[6518]_  = ~\new_[7116]_  | ~\new_[1313]_ ;
  assign \new_[6519]_  = ~\new_[7116]_  | ~\new_[1200]_ ;
  assign \new_[6520]_  = ~\new_[7116]_  | ~\new_[1145]_ ;
  assign \new_[6521]_  = ~\new_[7116]_  | ~\new_[1199]_ ;
  assign \new_[6522]_  = ~\new_[6775]_  | ~\new_[7564]_ ;
  assign \new_[6523]_  = ~\new_[6831]_  | ~\new_[7564]_ ;
  assign \new_[6524]_  = ~\new_[6908]_  | ~\new_[7564]_ ;
  assign \new_[6525]_  = ~\new_[6828]_  | ~\new_[7564]_ ;
  assign \new_[6526]_  = ~\new_[6902]_  | ~\new_[7564]_ ;
  assign \new_[6527]_  = ~\new_[6779]_  | ~\new_[7564]_ ;
  assign \new_[6528]_  = ~\new_[7423]_  | ~\new_[8996]_ ;
  assign \new_[6529]_  = ~\new_[8255]_  | ~\new_[8996]_ ;
  assign \new_[6530]_  = ~\new_[8313]_  | ~\new_[8996]_ ;
  assign \new_[6531]_  = ~\new_[7475]_  | ~\new_[8996]_ ;
  assign \new_[6532]_  = ~\new_[7827]_  & (~\new_[7038]_  | ~\new_[7028]_ );
  assign \new_[6533]_  = ~\new_[7827]_  & (~\new_[7035]_  | ~\new_[7027]_ );
  assign \new_[6534]_  = ~\new_[7827]_  & (~\new_[7032]_  | ~\new_[7110]_ );
  assign \new_[6535]_  = ~\new_[7827]_  & (~\new_[6943]_  | ~\new_[7099]_ );
  assign \new_[6536]_  = ~\new_[6878]_  | ~\new_[7818]_ ;
  assign \new_[6537]_  = ~\new_[7471]_  | ~\new_[8996]_ ;
  assign \new_[6538]_  = ~\new_[8302]_  | ~\new_[8996]_ ;
  assign \new_[6539]_  = ~\new_[8244]_  | ~\new_[8995]_ ;
  assign \new_[6540]_  = ~\new_[8256]_  | ~\new_[8996]_ ;
  assign \new_[6541]_  = ~\new_[6881]_  | ~\new_[7832]_ ;
  assign \new_[6542]_  = ~\new_[7827]_  & (~\new_[7031]_  | ~\new_[7098]_ );
  assign \new_[6543]_  = ~\new_[6872]_  | ~\new_[7820]_ ;
  assign \new_[6544]_  = ~\new_[6891]_  | ~\new_[7854]_ ;
  assign \new_[6545]_  = ~\new_[6879]_  | ~\new_[7820]_ ;
  assign \new_[6546]_  = \\mix1_data_o_reg_reg[49] ;
  assign \new_[6547]_  = \\mix1_data_o_reg_reg[116] ;
  assign \new_[6548]_  = \data_o[30]  ? \new_[8900]_  : \new_[1138]_ ;
  assign \new_[6549]_  = \data_o[31]  ? \new_[8941]_  : \new_[1246]_ ;
  assign \new_[6550]_  = \data_o[23]  ? \new_[8900]_  : \new_[1208]_ ;
  assign \new_[6551]_  = \data_o[79]  ? \new_[8893]_  : \new_[1201]_ ;
  assign \new_[6552]_  = \data_o[7]  ? \new_[8941]_  : \new_[1218]_ ;
  assign \new_[6553]_  = ~\new_[1384]_  | ~\new_[6954]_ ;
  assign \new_[6554]_  = ~\new_[8897]_  | ~\data_o[55] ;
  assign \new_[6555]_  = ~\new_[8897]_  | ~\data_o[69] ;
  assign \new_[6556]_  = ~\new_[8919]_  | ~\data_o[63] ;
  assign \new_[6557]_  = ~\new_[8924]_  | ~\new_[1213]_ ;
  assign \new_[6558]_  = ~\new_[8915]_  | ~\new_[1108]_ ;
  assign \new_[6559]_  = ~\new_[8900]_  | ~\new_[1186]_ ;
  assign \new_[6560]_  = ~\new_[8915]_  | ~\new_[1136]_ ;
  assign \new_[6561]_  = ~\new_[8934]_  | ~\new_[1115]_ ;
  assign \new_[6562]_  = ~\new_[8941]_  | ~\new_[1099]_ ;
  assign \new_[6563]_  = ~\new_[1242]_  | ~\new_[6954]_ ;
  assign \new_[6564]_  = ~\new_[1243]_  | ~\new_[6954]_ ;
  assign \new_[6565]_  = ~\new_[7075]_  | ~\new_[1140]_ ;
  assign \new_[6566]_  = \\mix1_data_o_reg_reg[86] ;
  assign \new_[6567]_  = ~\new_[1225]_  | ~\new_[6954]_ ;
  assign \new_[6568]_  = \\mix1_data_o_reg_reg[88] ;
  assign \new_[6569]_  = \\mix1_data_o_reg_reg[89] ;
  assign \new_[6570]_  = ~\new_[8941]_  | ~\new_[1111]_ ;
  assign \new_[6571]_  = \\mix1_data_o_reg_reg[126] ;
  assign \new_[6572]_  = \\mix1_data_o_reg_reg[90] ;
  assign \new_[6573]_  = \\mix1_data_o_reg_reg[74] ;
  assign \new_[6574]_  = \\mix1_data_o_reg_reg[56] ;
  assign \new_[6575]_  = \\mix1_data_o_reg_reg[47] ;
  assign \new_[6576]_  = \new_[8896]_  & \new_[1202]_ ;
  assign \new_[6577]_  = \new_[7116]_  & \new_[1112]_ ;
  assign \new_[6578]_  = ~\new_[7116]_  | ~\new_[5990]_ ;
  assign \new_[6579]_  = \\mix1_data_o_reg_reg[97] ;
  assign \new_[6580]_  = \\mix1_data_o_reg_reg[43] ;
  assign \new_[6581]_  = \\mix1_data_o_reg_reg[76] ;
  assign \new_[6582]_  = \new_[7116]_  & \new_[1115]_ ;
  assign \new_[6583]_  = \key_i[36]  ? \new_[7582]_  : \new_[8064]_ ;
  assign \new_[6584]_  = \\mix1_data_o_reg_reg[37] ;
  assign \new_[6585]_  = \\mix1_data_o_reg_reg[84] ;
  assign \new_[6586]_  = \\mix1_data_o_reg_reg[103] ;
  assign \new_[6587]_  = \\mix1_data_o_reg_reg[109] ;
  assign \new_[6588]_  = \\mix1_data_o_reg_reg[53] ;
  assign \new_[6589]_  = \\mix1_data_o_reg_reg[119] ;
  assign \new_[6590]_  = \\mix1_data_o_reg_reg[125] ;
  assign \new_[6591]_  = \\mix1_data_o_reg_reg[36] ;
  assign \new_[6592]_  = \\mix1_data_o_reg_reg[39] ;
  assign \new_[6593]_  = \\mix1_data_o_reg_reg[55] ;
  assign \new_[6594]_  = \\mix1_data_o_reg_reg[62] ;
  assign \new_[6595]_  = \\mix1_data_o_reg_reg[96] ;
  assign \new_[6596]_  = \\mix1_data_o_reg_reg[115] ;
  assign \new_[6597]_  = \\mix1_data_o_reg_reg[46] ;
  assign \new_[6598]_  = \\mix1_data_o_reg_reg[80] ;
  assign \new_[6599]_  = \\mix1_data_o_reg_reg[123] ;
  assign \new_[6600]_  = \\mix1_data_o_reg_reg[83] ;
  assign \new_[6601]_  = \\mix1_data_o_reg_reg[58] ;
  assign \new_[6602]_  = (~\new_[7660]_  | ~\key_i[67] ) & (~\new_[7620]_  | ~\new_[2134]_ );
  assign \new_[6603]_  = \key_i[37]  ? \new_[7582]_  : \new_[8109]_ ;
  assign \new_[6604]_  = ~\new_[7114]_  | ~\new_[1193]_ ;
  assign \new_[6605]_  = \\mix1_data_o_reg_reg[68] ;
  assign \new_[6606]_  = \\mix1_data_o_reg_reg[101] ;
  assign \new_[6607]_  = \\mix1_data_o_reg_reg[118] ;
  assign \new_[6608]_  = (~\new_[7660]_  | ~\key_i[95] ) & (~\new_[7620]_  | ~\new_[2069]_ );
  assign \new_[6609]_  = \\mix1_data_o_reg_reg[52] ;
  assign \new_[6610]_  = \\mix1_data_o_reg_reg[59] ;
  assign \new_[6611]_  = \new_[8897]_  & \data_o[127] ;
  assign \new_[6612]_  = ~\new_[7114]_  | ~\new_[1191]_ ;
  assign \new_[6613]_  = ~\new_[8925]_  | ~\data_o[39] ;
  assign \new_[6614]_  = \\mix1_data_o_reg_reg[87] ;
  assign \new_[6615]_  = \new_[6595]_  ? \new_[8904]_  : \data_o[96] ;
  assign \new_[6616]_  = \\mix1_data_o_reg_reg[51] ;
  assign \new_[6617]_  = ~\new_[7114]_  | ~\new_[1311]_ ;
  assign \new_[6618]_  = \\mix1_data_o_reg_reg[66] ;
  assign \new_[6619]_  = \\mix1_data_o_reg_reg[81] ;
  assign \new_[6620]_  = \\mix1_data_o_reg_reg[107] ;
  assign \new_[6621]_  = \new_[8941]_  & \new_[1205]_ ;
  assign \new_[6622]_  = \new_[7116]_  & \new_[1104]_ ;
  assign \new_[6623]_  = \\mix1_data_o_reg_reg[44] ;
  assign \new_[6624]_  = \\mix1_data_o_reg_reg[42] ;
  assign \new_[6625]_  = \\mix1_data_o_reg_reg[94] ;
  assign \new_[6626]_  = \\mix1_data_o_reg_reg[54] ;
  assign \new_[6627]_  = \\mix1_data_o_reg_reg[50] ;
  assign \new_[6628]_  = \\mix1_data_o_reg_reg[124] ;
  assign \new_[6629]_  = \\mix1_data_o_reg_reg[32] ;
  assign \new_[6630]_  = \\mix1_data_o_reg_reg[75] ;
  assign \new_[6631]_  = \\mix1_data_o_reg_reg[61] ;
  assign \new_[6632]_  = \\mix1_data_o_reg_reg[63] ;
  assign \new_[6633]_  = \new_[8919]_  & \data_o[119] ;
  assign \new_[6634]_  = ~\new_[7116]_  | ~\new_[6041]_ ;
  assign \new_[6635]_  = \key_i[41]  ? \new_[7582]_  : \new_[1119]_ ;
  assign \new_[6636]_  = ~\new_[6953]_  & (~\new_[7683]_  | ~\new_[7851]_ );
  assign \new_[6637]_  = ~\new_[6755]_ ;
  assign \new_[6638]_  = ~\new_[6755]_ ;
  assign \new_[6639]_  = \\mix1_data_o_reg_reg[120] ;
  assign \new_[6640]_  = \\mix1_data_o_reg_reg[40] ;
  assign \new_[6641]_  = \\mix1_data_o_reg_reg[111] ;
  assign \new_[6642]_  = ~\new_[7115]_ ;
  assign \new_[6643]_  = \\mix1_data_o_reg_reg[34] ;
  assign \new_[6644]_  = ~\new_[6951]_  & (~\new_[7648]_  | ~\new_[7927]_ );
  assign \new_[6645]_  = (~\new_[7201]_  | ~\new_[7836]_ ) & (~\new_[7105]_  | ~\new_[7833]_ );
  assign \new_[6646]_  = (~\new_[7137]_  | ~\new_[7833]_ ) & (~\new_[7245]_  | ~\new_[7866]_ );
  assign \new_[6647]_  = (~\new_[7101]_  | ~\new_[7833]_ ) & (~\new_[7087]_  | ~\new_[7866]_ );
  assign \new_[6648]_  = (~\new_[7136]_  | ~\new_[7833]_ ) & (~\new_[7393]_  | ~\new_[7861]_ );
  assign \new_[6649]_  = ~\new_[6827]_ ;
  assign \new_[6650]_  = ~\new_[6791]_ ;
  assign \new_[6651]_  = ~\new_[6792]_ ;
  assign \new_[6652]_  = \\mix1_data_o_reg_reg[113] ;
  assign \new_[6653]_  = ~\new_[6797]_ ;
  assign \new_[6654]_  = ~\new_[6798]_ ;
  assign \new_[6655]_  = (~\new_[7134]_  | ~\new_[7815]_ ) & (~\new_[7272]_  | ~\new_[7864]_ );
  assign \new_[6656]_  = \\mix1_data_o_reg_reg[41] ;
  assign \new_[6657]_  = (~\new_[7133]_  | ~\new_[7866]_ ) & (~\new_[7085]_  | ~\new_[7852]_ );
  assign \new_[6658]_  = (~\new_[7096]_  | ~\new_[7836]_ ) & (~\new_[7246]_  | ~\new_[7852]_ );
  assign \new_[6659]_  = (~\new_[7124]_  | ~\new_[7838]_ ) & (~\new_[7248]_  | ~\new_[7861]_ );
  assign \new_[6660]_  = (~\new_[7088]_  | ~\new_[7864]_ ) & (~\new_[7279]_  | ~\new_[7852]_ );
  assign \new_[6661]_  = (~\new_[7132]_  | ~\new_[7838]_ ) & (~\new_[7268]_  | ~\new_[7861]_ );
  assign \new_[6662]_  = (~\new_[7086]_  | ~\new_[7838]_ ) & (~\new_[7217]_  | ~\new_[7861]_ );
  assign \new_[6663]_  = \\mix1_data_o_reg_reg[121] ;
  assign \new_[6664]_  = (~\new_[7093]_  | ~\new_[7836]_ ) & (~\new_[7135]_  | ~\new_[7852]_ );
  assign \new_[6665]_  = (~\new_[7128]_  | ~\new_[7861]_ ) & (~\new_[7274]_  | ~\new_[7838]_ );
  assign \new_[6666]_  = \\mix1_data_o_reg_reg[92] ;
  assign \new_[6667]_  = ~\new_[7570]_  | ~\new_[8990]_ ;
  assign \new_[6668]_  = ~\new_[7116]_  | ~\new_[5991]_ ;
  assign \new_[6669]_  = ~\new_[7114]_  | ~\new_[1198]_ ;
  assign \new_[6670]_  = \new_[7116]_  & \new_[1103]_ ;
  assign \new_[6671]_  = ~\new_[7114]_  | ~\new_[1457]_ ;
  assign \new_[6672]_  = ~\new_[7114]_  | ~\new_[1312]_ ;
  assign \new_[6673]_  = ~\new_[7114]_  | ~\new_[1192]_ ;
  assign \new_[6674]_  = ~\new_[7114]_  | ~\new_[1190]_ ;
  assign \new_[6675]_  = ~\new_[7114]_  | ~\new_[1201]_ ;
  assign \new_[6676]_  = ~\new_[7114]_  | ~\new_[1458]_ ;
  assign \new_[6677]_  = ~\new_[7114]_  | ~\new_[1195]_ ;
  assign \new_[6678]_  = ~\new_[7114]_  | ~\new_[1196]_ ;
  assign \new_[6679]_  = \new_[7116]_  & \new_[1107]_ ;
  assign \new_[6680]_  = \new_[7116]_  & \new_[1106]_ ;
  assign \new_[6681]_  = ~\new_[7114]_  | ~\new_[1314]_ ;
  assign \new_[6682]_  = ~\new_[7114]_  | ~\new_[1197]_ ;
  assign \new_[6683]_  = ~\new_[7114]_  | ~\new_[1143]_ ;
  assign \new_[6684]_  = \new_[7116]_  & \new_[1113]_ ;
  assign \new_[6685]_  = \new_[7116]_  & \new_[1109]_ ;
  assign \new_[6686]_  = \new_[7116]_  & \new_[1110]_ ;
  assign \new_[6687]_  = ~\new_[7114]_  | ~\new_[1194]_ ;
  assign \new_[6688]_  = \new_[7116]_  & \new_[1114]_ ;
  assign \new_[6689]_  = \new_[7116]_  & \new_[1108]_ ;
  assign \new_[6690]_  = \new_[7116]_  & \new_[1117]_ ;
  assign \new_[6691]_  = ~\new_[7084]_  | ~\new_[7564]_ ;
  assign \new_[6692]_  = ~\new_[7065]_  | ~\new_[7564]_ ;
  assign \new_[6693]_  = ~\new_[7067]_  | ~\new_[7564]_ ;
  assign \new_[6694]_  = \\mix1_data_o_reg_reg[117] ;
  assign \new_[6695]_  = ~\new_[6938]_  | ~\new_[7564]_ ;
  assign \new_[6696]_  = ~\new_[7079]_  | ~\new_[7564]_ ;
  assign \new_[6697]_  = ~\new_[7074]_  | ~\new_[7564]_ ;
  assign \new_[6698]_  = ~\new_[7568]_  | ~\new_[8996]_ ;
  assign \new_[6699]_  = \new_[7007]_  & \new_[7604]_ ;
  assign \new_[6700]_  = \new_[7017]_  & \new_[7604]_ ;
  assign \new_[6701]_  = \new_[7651]_  & \new_[8990]_ ;
  assign \new_[6702]_  = \\mix1_data_o_reg_reg[60] ;
  assign \new_[6703]_  = ~\new_[7259]_ ;
  assign \new_[6704]_  = \\mix1_data_o_reg_reg[114] ;
  assign \new_[6705]_  = ~\new_[8303]_  | ~\new_[8995]_ ;
  assign \new_[6706]_  = \new_[7036]_  & \new_[7604]_ ;
  assign \new_[6707]_  = ~\new_[7574]_  | ~\new_[8996]_ ;
  assign \new_[6708]_  = ~\new_[7575]_  | ~\new_[8987]_ ;
  assign \new_[6709]_  = \new_[7649]_  & \new_[8996]_ ;
  assign \new_[6710]_  = ~\new_[7610]_  | ~\new_[8996]_ ;
  assign \new_[6711]_  = \new_[8284]_  & \new_[8996]_ ;
  assign \new_[6712]_  = ~\new_[7012]_  | ~\new_[7865]_ ;
  assign \new_[6713]_  = ~\new_[7578]_  | ~\new_[8987]_ ;
  assign \new_[6714]_  = \\mix1_data_o_reg_reg[38] ;
  assign \new_[6715]_  = ~\new_[7627]_  & ~\new_[7648]_ ;
  assign \new_[6716]_  = \\mix1_data_o_reg_reg[73] ;
  assign \new_[6717]_  = \data_o[71]  ? \new_[8902]_  : \new_[1219]_ ;
  assign \new_[6718]_  = \new_[6427]_  ? \new_[8941]_  : \data_o[85] ;
  assign \new_[6719]_  = (~\new_[6574]_  | ~\new_[8945]_ ) & (~\new_[8918]_  | ~\data_o[56] );
  assign \new_[6720]_  = (~\new_[6596]_  | ~\new_[8897]_ ) & (~\new_[8893]_  | ~\data_o[115] );
  assign \new_[6721]_  = \new_[6584]_  ? \new_[8904]_  : \data_o[37] ;
  assign \new_[6722]_  = \data_o[47]  ? \new_[8902]_  : \new_[1198]_ ;
  assign \new_[6723]_  = \\mix1_data_o_reg_reg[127] ;
  assign \new_[6724]_  = ~\new_[8942]_  | ~\data_o[38] ;
  assign \new_[6725]_  = \new_[8933]_  & \data_o[118] ;
  assign \new_[6726]_  = \new_[8933]_  & \data_o[111] ;
  assign \new_[6727]_  = \new_[8933]_  & \data_o[103] ;
  assign \new_[6728]_  = ~\new_[8905]_  | ~\data_o[46] ;
  assign \new_[6729]_  = ~\new_[8919]_  | ~\data_o[54] ;
  assign \new_[6730]_  = ~\new_[8919]_  | ~\data_o[62] ;
  assign \new_[6731]_  = ~\new_[8924]_  | ~\new_[1109]_ ;
  assign \new_[6732]_  = ~\new_[8915]_  | ~\new_[1249]_ ;
  assign \new_[6733]_  = \new_[7930]_  ? \new_[7584]_  : \new_[7840]_ ;
  assign \new_[6734]_  = \key_i[38]  ? \new_[7582]_  : \new_[8156]_ ;
  assign \new_[6735]_  = (~\new_[7660]_  | ~\key_i[81] ) & (~\new_[7581]_  | ~\new_[2162]_ );
  assign \new_[6736]_  = \key_i[40]  ? \new_[7582]_  : \new_[1089]_ ;
  assign \new_[6737]_  = \key_i[39]  ? \new_[7582]_  : \new_[8150]_ ;
  assign \new_[6738]_  = (~\new_[7660]_  | ~\key_i[82] ) & (~\new_[7581]_  | ~\new_[2202]_ );
  assign \new_[6739]_  = \key_i[35]  ? \new_[7582]_  : \new_[7991]_ ;
  assign \new_[6740]_  = (~\new_[7660]_  | ~\key_i[66] ) & (~\new_[7581]_  | ~\new_[2135]_ );
  assign \new_[6741]_  = (~\new_[7660]_  | ~\key_i[94] ) & (~\new_[7620]_  | ~\new_[2068]_ );
  assign \new_[6742]_  = (~\new_[7660]_  | ~\key_i[88] ) & (~\new_[7769]_  | ~\new_[2067]_ );
  assign \new_[6743]_  = (~\new_[7660]_  | ~\key_i[89] ) & (~\new_[7769]_  | ~\new_[2070]_ );
  assign \new_[6744]_  = (~\new_[7660]_  | ~\key_i[91] ) & (~\new_[7620]_  | ~\new_[2043]_ );
  assign \new_[6745]_  = ~\new_[7115]_ ;
  assign \new_[6746]_  = \\mix1_data_o_reg_reg[95] ;
  assign \new_[6747]_  = \new_[8918]_  & \new_[1192]_ ;
  assign \new_[6748]_  = \\mix1_data_o_reg_reg[79] ;
  assign \new_[6749]_  = \\mix1_data_o_reg_reg[35] ;
  assign \new_[6750]_  = ~\new_[8946]_  | ~\new_[1238]_ ;
  assign \new_[6751]_  = \\mix1_data_o_reg_reg[100] ;
  assign \new_[6752]_  = ~\new_[7102]_ ;
  assign \new_[6753]_  = (~\new_[1234]_  | ~\new_[7632]_ ) & (~\new_[1214]_  | ~\new_[7738]_ );
  assign \new_[6754]_  = (~\new_[6702]_  | ~\new_[8919]_ ) & (~\new_[8940]_  | ~\data_o[60] );
  assign \new_[6755]_  = ~\new_[6914]_ ;
  assign \new_[6756]_  = \new_[8158]_  | \new_[8996]_ ;
  assign \new_[6757]_  = \new_[6749]_  ? \new_[8921]_  : \data_o[35] ;
  assign \new_[6758]_  = \new_[6751]_  ? \new_[8926]_  : \data_o[100] ;
  assign n3745 = ~\new_[7484]_  | ~\new_[7177]_ ;
  assign \new_[6760]_  = (~\new_[1237]_  | ~\new_[7632]_ ) & (~\new_[1240]_  | ~\new_[7738]_ );
  assign \new_[6761]_  = ~\new_[6423]_  | ~\new_[8919]_ ;
  assign \new_[6762]_  = \key_i[77]  ? \new_[7620]_  : \new_[1132]_ ;
  assign \new_[6763]_  = ~\new_[6947]_ ;
  assign \new_[6764]_  = ~\new_[6947]_ ;
  assign n3725 = ~\new_[7431]_  | ~\new_[7188]_ ;
  assign \new_[6766]_  = (~\new_[1319]_  | ~\new_[7632]_ ) & (~\new_[1323]_  | ~\new_[7738]_ );
  assign \new_[6767]_  = ~\new_[8900]_  | ~\data_o[117] ;
  assign \new_[6768]_  = \new_[6566]_  ? \new_[8946]_  : \data_o[86] ;
  assign \new_[6769]_  = \new_[8078]_  | \new_[8987]_ ;
  assign \new_[6770]_  = ~\new_[7239]_ ;
  assign \new_[6771]_  = ks1_ready_o_reg;
  assign \new_[6772]_  = \new_[6620]_  ? \new_[8918]_  : \data_o[107] ;
  assign \new_[6773]_  = \key_i[74]  ? \new_[7620]_  : \new_[8130]_ ;
  assign \new_[6774]_  = ~\new_[7239]_ ;
  assign \new_[6775]_  = \new_[1110]_  ? \new_[7632]_  : \new_[1105]_ ;
  assign \new_[6776]_  = ~\new_[7102]_ ;
  assign \new_[6777]_  = ~\new_[7102]_ ;
  assign \new_[6778]_  = ~\new_[7102]_ ;
  assign \new_[6779]_  = \new_[1102]_  ? \new_[7632]_  : \new_[1109]_ ;
  assign \new_[6780]_  = \new_[6914]_ ;
  assign n3680 = ~\new_[7516]_  | ~\new_[7108]_ ;
  assign n3675 = ~\new_[7553]_  | ~\new_[7185]_ ;
  assign n3765 = ~\new_[7433]_  | ~\new_[7184]_ ;
  assign \new_[6784]_  = ~\new_[7239]_ ;
  assign \new_[6785]_  = ~\new_[6947]_ ;
  assign \new_[6786]_  = ~\new_[6947]_ ;
  assign \new_[6787]_  = (~\new_[1207]_  | ~\new_[7632]_ ) & (~\new_[1221]_  | ~\new_[7738]_ );
  assign \new_[6788]_  = ~\new_[6919]_ ;
  assign \new_[6789]_  = (~\new_[7244]_  | ~\new_[7833]_ ) & (~\new_[7252]_  | ~\new_[7866]_ );
  assign \new_[6790]_  = ~\new_[6950]_ ;
  assign \new_[6791]_  = ~\new_[7118]_  & ~\new_[7853]_ ;
  assign \new_[6792]_  = ~\new_[7118]_  & ~\new_[7837]_ ;
  assign \new_[6793]_  = ~\new_[7102]_ ;
  assign \new_[6794]_  = ~\new_[7102]_ ;
  assign \new_[6795]_  = ~\new_[7102]_ ;
  assign \new_[6796]_  = ~\new_[7102]_ ;
  assign \new_[6797]_  = ~\new_[7131]_  & ~\new_[7853]_ ;
  assign \new_[6798]_  = ~\new_[7131]_  & ~\new_[7837]_ ;
  assign \new_[6799]_  = (~\new_[7280]_  | ~\new_[7815]_ ) & (~\new_[7256]_  | ~\new_[7838]_ );
  assign \new_[6800]_  = (~\new_[7213]_  | ~\new_[7815]_ ) & (~\new_[7273]_  | ~\new_[7864]_ );
  assign \new_[6801]_  = (~\new_[7276]_  | ~\new_[7815]_ ) & (~\new_[7277]_  | ~\new_[7864]_ );
  assign \new_[6802]_  = \new_[8058]_  | \new_[8995]_ ;
  assign \new_[6803]_  = ~\new_[7259]_ ;
  assign \new_[6804]_  = (~\new_[7222]_  | ~\new_[7866]_ ) & (~\new_[7396]_  | ~\new_[7861]_ );
  assign \new_[6805]_  = (~\new_[1521]_  | ~\new_[7632]_ ) & (~\new_[1530]_  | ~\new_[7738]_ );
  assign \new_[6806]_  = (~\new_[7278]_  | ~\new_[7836]_ ) & (~\new_[7218]_  | ~\new_[7852]_ );
  assign \new_[6807]_  = (~\new_[1321]_  | ~\new_[7632]_ ) & (~\new_[1315]_  | ~\new_[7738]_ );
  assign \new_[6808]_  = ~\new_[7259]_ ;
  assign \new_[6809]_  = ~\new_[7259]_ ;
  assign \new_[6810]_  = \new_[7936]_  | \new_[8996]_ ;
  assign \new_[6811]_  = \new_[8072]_  | \new_[8987]_ ;
  assign \new_[6812]_  = \new_[8071]_  | \new_[8990]_ ;
  assign \new_[6813]_  = \new_[7996]_  | \new_[8996]_ ;
  assign \new_[6814]_  = \new_[8034]_  | \new_[8996]_ ;
  assign \new_[6815]_  = \new_[7995]_  | \new_[8987]_ ;
  assign \new_[6816]_  = \new_[7946]_  | \new_[8996]_ ;
  assign \new_[6817]_  = \new_[8105]_  | \new_[8990]_ ;
  assign \new_[6818]_  = \new_[8103]_  | \new_[8990]_ ;
  assign \new_[6819]_  = \new_[7950]_  | \new_[8996]_ ;
  assign \new_[6820]_  = \new_[8031]_  | \new_[8996]_ ;
  assign \new_[6821]_  = \new_[8139]_  | \new_[8987]_ ;
  assign \new_[6822]_  = \new_[7093]_  & \new_[7604]_ ;
  assign \new_[6823]_  = \new_[7096]_  & \new_[7604]_ ;
  assign \new_[6824]_  = ~\new_[7259]_ ;
  assign \new_[6825]_  = ~\new_[7259]_ ;
  assign \new_[6826]_  = \new_[7201]_  & \new_[7604]_ ;
  assign \new_[6827]_  = ~\new_[7622]_  & ~\new_[7196]_ ;
  assign \new_[6828]_  = \new_[1103]_  ? \new_[7632]_  : \new_[1108]_ ;
  assign \new_[6829]_  = ~\new_[7632]_  | ~load_i | ~\new_[5784]_ ;
  assign \new_[6830]_  = \new_[6619]_  ? \new_[8894]_  : \data_o[81] ;
  assign \new_[6831]_  = \new_[1111]_  ? \new_[7632]_  : \new_[1104]_ ;
  assign \new_[6832]_  = ~\new_[7261]_ ;
  assign n3780 = ~\new_[7505]_  | ~\new_[7154]_ ;
  assign n3685 = ~\new_[7506]_  | ~\new_[7195]_ ;
  assign n3645 = ~\new_[7418]_  | ~\new_[7165]_ ;
  assign n3695 = ~\new_[7512]_  | ~\new_[7109]_ ;
  assign n3635 = ~\new_[7489]_  | ~\new_[7091]_ ;
  assign n3730 = ~\new_[7555]_  | ~\new_[7090]_ ;
  assign n3735 = ~\new_[7508]_  | ~\new_[7152]_ ;
  assign n3640 = ~\new_[7445]_  | ~\new_[7171]_ ;
  assign n3700 = ~\new_[7522]_  | ~\new_[7150]_ ;
  assign n3715 = ~\new_[7518]_  | ~\new_[7186]_ ;
  assign n3650 = ~\new_[7442]_  | ~\new_[7197]_ ;
  assign n3655 = ~\new_[7551]_  | ~\new_[7199]_ ;
  assign n3760 = ~\new_[7421]_  | ~\new_[7157]_ ;
  assign n3755 = ~\new_[7447]_  | ~\new_[7189]_ ;
  assign n3740 = ~\new_[7527]_  | ~\new_[7173]_ ;
  assign n3690 = ~\new_[7407]_  | ~\new_[7194]_ ;
  assign n3665 = ~\new_[7519]_  | ~\new_[7198]_ ;
  assign n3750 = ~\new_[7483]_  | ~\new_[7180]_ ;
  assign n3775 = ~\new_[7425]_  | ~\new_[7166]_ ;
  assign n3670 = ~\new_[7468]_  | ~\new_[7179]_ ;
  assign n3705 = ~\new_[7533]_  | ~\new_[7162]_ ;
  assign n3625 = ~\new_[7492]_  | ~\new_[7163]_ ;
  assign n3720 = ~\new_[7510]_  | ~\new_[7191]_ ;
  assign n3770 = ~\new_[7554]_  | ~\new_[7183]_ ;
  assign n3660 = ~\new_[7534]_  | ~\new_[7155]_ ;
  assign n3710 = ~\new_[7548]_  | ~\new_[7164]_ ;
  assign n3630 = ~\new_[7466]_  | ~\new_[7158]_ ;
  assign \new_[6860]_  = \new_[3863]_  ? \new_[8921]_  : \data_o[31] ;
  assign \new_[6861]_  = \new_[6422]_  ? \new_[8904]_  : \data_o[110] ;
  assign \new_[6862]_  = \new_[3377]_  ? \new_[8900]_  : \data_o[8] ;
  assign \new_[6863]_  = \new_[6419]_  ? \new_[8902]_  : \data_o[102] ;
  assign \new_[6864]_  = \new_[6586]_  ? \new_[8893]_  : \data_o[103] ;
  assign \new_[6865]_  = \new_[2934]_  ? \new_[8904]_  : \data_o[11] ;
  assign \new_[6866]_  = \new_[3846]_  ? \new_[8904]_  : \data_o[7] ;
  assign \new_[6867]_  = \new_[6579]_  ? \new_[8902]_  : \data_o[97] ;
  assign \new_[6868]_  = \new_[6614]_  ? \new_[8938]_  : \data_o[87] ;
  assign \new_[6869]_  = \new_[6714]_  ? \new_[8900]_  : \data_o[38] ;
  assign \new_[6870]_  = \new_[6416]_  ? \new_[8918]_  : \data_o[104] ;
  assign \new_[6871]_  = \new_[6449]_  ? \new_[8940]_  : \data_o[106] ;
  assign \new_[6872]_  = \new_[2932]_  ? \new_[8918]_  : \data_o[27] ;
  assign \new_[6873]_  = \new_[2757]_  ? \new_[8944]_  : \data_o[28] ;
  assign \new_[6874]_  = \new_[6629]_  ? \new_[8938]_  : \data_o[32] ;
  assign \new_[6875]_  = (~\new_[6601]_  | ~\new_[8945]_ ) & (~\new_[8893]_  | ~\data_o[58] );
  assign \new_[6876]_  = \new_[3514]_  ? \new_[8902]_  : \data_o[29] ;
  assign \new_[6877]_  = \new_[6421]_  ? \new_[8921]_  : \data_o[108] ;
  assign \new_[6878]_  = \new_[6587]_  ? \new_[8946]_  : \data_o[109] ;
  assign \new_[6879]_  = \new_[3107]_  ? \new_[8918]_  : \data_o[26] ;
  assign \new_[6880]_  = \new_[6600]_  ? \new_[8900]_  : \data_o[83] ;
  assign \new_[6881]_  = \new_[3382]_  ? \new_[8904]_  : \data_o[13] ;
  assign \new_[6882]_  = \new_[6643]_  ? \new_[8940]_  : \data_o[34] ;
  assign \new_[6883]_  = \new_[6430]_  ? \new_[8940]_  : \data_o[99] ;
  assign \new_[6884]_  = ~\new_[6610]_  | ~\new_[8925]_ ;
  assign \new_[6885]_  = ~\new_[6694]_  | ~\new_[8947]_ ;
  assign \new_[6886]_  = ~\new_[6594]_  | ~\new_[8905]_ ;
  assign \new_[6887]_  = ~\new_[6631]_  | ~\new_[8919]_ ;
  assign \new_[6888]_  = ~\new_[8900]_  | ~\data_o[62] ;
  assign \new_[6889]_  = ~\new_[8918]_  | ~\data_o[61] ;
  assign \new_[6890]_  = ~\new_[8918]_  | ~\data_o[112] ;
  assign \new_[6891]_  = \new_[6598]_  ? \new_[8893]_  : \data_o[80] ;
  assign \new_[6892]_  = ~\new_[8900]_  | ~\data_o[59] ;
  assign \new_[6893]_  = \new_[8941]_  & \new_[1243]_ ;
  assign \new_[6894]_  = \key_i[127]  ? \new_[7620]_  : \new_[2266]_ ;
  assign \new_[6895]_  = \key_i[120]  ? \new_[7620]_  : \new_[2264]_ ;
  assign \new_[6896]_  = \key_i[121]  ? \new_[7620]_  : \new_[2265]_ ;
  assign \new_[6897]_  = \key_i[122]  ? \new_[7769]_  : \new_[2273]_ ;
  assign \new_[6898]_  = \key_i[93]  ? \new_[7582]_  : \new_[8094]_ ;
  assign \new_[6899]_  = \key_i[90]  ? \new_[7582]_  : \new_[8037]_ ;
  assign \new_[6900]_  = \new_[8915]_  & \new_[1102]_ ;
  assign \new_[6901]_  = \new_[8918]_  & \new_[1104]_ ;
  assign \new_[6902]_  = \new_[1106]_  ? \new_[7632]_  : \new_[1116]_ ;
  assign \new_[6903]_  = (~\new_[1152]_  | ~\new_[7632]_ ) & (~\new_[1147]_  | ~\new_[7738]_ );
  assign \new_[6904]_  = (~\new_[1381]_  | ~\new_[7632]_ ) & (~\new_[1324]_  | ~\new_[7738]_ );
  assign \new_[6905]_  = (~\new_[1238]_  | ~\new_[7632]_ ) & (~\new_[1202]_  | ~\new_[7738]_ );
  assign \new_[6906]_  = (~\new_[1538]_  | ~\new_[7632]_ ) & (~\new_[1464]_  | ~\new_[7738]_ );
  assign \new_[6907]_  = (~\new_[1461]_  | ~\new_[7632]_ ) & (~\new_[1520]_  | ~\new_[7738]_ );
  assign \new_[6908]_  = \new_[1107]_  ? \new_[7632]_  : \new_[1117]_ ;
  assign \new_[6909]_  = (~\new_[1208]_  | ~\new_[7632]_ ) & (~\new_[1222]_  | ~\new_[7738]_ );
  assign n3915 = ~\new_[7439]_  | ~\new_[7340]_ ;
  assign \new_[6911]_  = (~\new_[1148]_  | ~\new_[7632]_ ) & (~\new_[1150]_  | ~\new_[7738]_ );
  assign \new_[6912]_  = ~\new_[8900]_  | ~\data_o[57] ;
  assign \new_[6913]_  = (~\new_[1211]_  | ~\new_[7632]_ ) & (~\new_[1203]_  | ~\new_[7738]_ );
  assign \new_[6914]_  = ~\new_[7260]_  & ~\new_[8052]_ ;
  assign \new_[6915]_  = \new_[3409]_  ? \new_[8935]_  : \data_o[14] ;
  assign n3835 = ~\new_[7528]_  | ~\new_[7382]_ ;
  assign n3940 = ~\new_[7520]_  | ~\new_[7253]_ ;
  assign \new_[6918]_  = (~\new_[1319]_  | ~\new_[7738]_ ) & (~\new_[1323]_  | ~\new_[7632]_ );
  assign \new_[6919]_  = ~\new_[7115]_ ;
  assign \new_[6920]_  = \new_[6420]_  ? \new_[8935]_  : \data_o[105] ;
  assign \new_[6921]_  = \new_[6575]_  ? \new_[8926]_  : \data_o[47] ;
  assign n4080 = ~\new_[7435]_  | ~\new_[7336]_ ;
  assign \new_[6923]_  = (~\new_[1208]_  | ~\new_[7738]_ ) & (~\new_[1222]_  | ~\new_[7569]_ );
  assign \new_[6924]_  = (~\new_[7660]_  | ~\key_i[80] ) & (~\new_[7581]_  | ~\new_[2198]_ );
  assign \new_[6925]_  = ~\new_[8343]_  | ~\new_[8119]_ ;
  assign \new_[6926]_  = (~\new_[1321]_  | ~\new_[7738]_ ) & (~\new_[1315]_  | ~\new_[7569]_ );
  assign n3930 = ~\new_[7545]_  | ~\new_[7288]_ ;
  assign \new_[6928]_  = (~\new_[1212]_  | ~\new_[7632]_ ) & (~\new_[1204]_  | ~\new_[7738]_ );
  assign \new_[6929]_  = \new_[2755]_  ? \new_[8920]_  : \data_o[12] ;
  assign n3995 = ~\new_[7517]_  | ~\new_[7220]_ ;
  assign \new_[6931]_  = \new_[6641]_  ? \new_[8938]_  : \data_o[111] ;
  assign \new_[6932]_  = \new_[2935]_  ? \new_[8944]_  : \data_o[19] ;
  assign \new_[6933]_  = \new_[6748]_  ? \new_[8918]_  : \data_o[79] ;
  assign \new_[6934]_  = \new_[6446]_  ? \new_[8918]_  : \data_o[71] ;
  assign \new_[6935]_  = \new_[6588]_  ? \new_[8904]_  : \data_o[53] ;
  assign \new_[6936]_  = ~\new_[7384]_  | ~\new_[1072]_ ;
  assign \new_[6937]_  = (~\new_[1213]_  | ~\new_[7632]_ ) & (~\new_[1205]_  | ~\new_[7738]_ );
  assign \new_[6938]_  = \new_[1107]_  ? \new_[7738]_  : \new_[1117]_ ;
  assign \new_[6939]_  = (~\new_[1538]_  | ~\new_[7738]_ ) & (~\new_[1464]_  | ~\new_[7632]_ );
  assign n4025 = ~\new_[7513]_  | ~\new_[7368]_ ;
  assign n3810 = ~\new_[7422]_  | ~\new_[7343]_ ;
  assign n3850 = ~\new_[7531]_  | ~\new_[7375]_ ;
  assign \new_[6943]_  = ~\new_[8920]_  | ~\data_o[119] ;
  assign n3830 = ~\new_[7416]_  | ~\new_[7337]_ ;
  assign n3800 = ~\new_[7515]_  | ~\new_[7258]_ ;
  assign n3925 = ~\new_[7541]_  | ~\new_[7307]_ ;
  assign \new_[6947]_  = ~\new_[7097]_ ;
  assign n4020 = ~\new_[7426]_  | ~\new_[7331]_ ;
  assign \new_[6949]_  = ~\new_[7622]_  & ~\new_[7265]_ ;
  assign \new_[6950]_  = \new_[7622]_  & \new_[7264]_ ;
  assign \new_[6951]_  = ~\new_[7648]_  & (~\new_[7640]_  | ~\new_[7488]_ );
  assign \new_[6952]_  = mix1_ready_o_reg;
  assign \new_[6953]_  = ~\new_[7239]_  & ~\new_[5784]_ ;
  assign \new_[6954]_  = ~\new_[7259]_ ;
  assign \new_[6955]_  = ~\new_[7250]_  | ~\new_[7826]_ ;
  assign \new_[6956]_  = \new_[7278]_  & \new_[7604]_ ;
  assign \new_[6957]_  = ~\new_[7250]_  | ~\new_[7688]_ ;
  assign \new_[6958]_  = ~\new_[7266]_  | ~\new_[7588]_ ;
  assign n3825 = ~\new_[7417]_  | ~\new_[7346]_ ;
  assign n3815 = ~\new_[7507]_  | ~\new_[7369]_ ;
  assign n4085 = ~\new_[7495]_  | ~\new_[7352]_ ;
  assign n4095 = ~\new_[7461]_  | ~\new_[7316]_ ;
  assign n3960 = ~\new_[7504]_  | ~\new_[7238]_ ;
  assign n4065 = ~\new_[7493]_  | ~\new_[7326]_ ;
  assign n3885 = ~\new_[7514]_  | ~\new_[7342]_ ;
  assign n4015 = ~\new_[7529]_  | ~\new_[7257]_ ;
  assign n3990 = ~\new_[7547]_  | ~\new_[7226]_ ;
  assign n3905 = ~\new_[7487]_  | ~\new_[7249]_ ;
  assign n3955 = ~\new_[7455]_  | ~\new_[7225]_ ;
  assign n3970 = ~\new_[7414]_  | ~\new_[7309]_ ;
  assign n4035 = ~\new_[7476]_  | ~\new_[7367]_ ;
  assign n4070 = ~\new_[7481]_  | ~\new_[7335]_ ;
  assign n4040 = ~\new_[7502]_  | ~\new_[7376]_ ;
  assign n4005 = ~\new_[7436]_  | ~\new_[7289]_ ;
  assign n3875 = ~\new_[7424]_  | ~\new_[7355]_ ;
  assign n3855 = ~\new_[7546]_  | ~\new_[7380]_ ;
  assign n4000 = ~\new_[7530]_  | ~\new_[7317]_ ;
  assign n3895 = ~\new_[7441]_  | ~\new_[7247]_ ;
  assign n3790 = ~\new_[7552]_  | ~\new_[7212]_ ;
  assign n4050 = ~\new_[7558]_  | ~\new_[7328]_ ;
  assign n3975 = ~\new_[7446]_  | ~\new_[7318]_ ;
  assign n3820 = ~\new_[7521]_  | ~\new_[7360]_ ;
  assign n3840 = ~\new_[7524]_  | ~\new_[7381]_ ;
  assign n3985 = ~\new_[7465]_  | ~\new_[7388]_ ;
  assign n3900 = ~\new_[7525]_  | ~\new_[7399]_ ;
  assign n3865 = ~\new_[7550]_  | ~\new_[7344]_ ;
  assign n4045 = ~\new_[7503]_  | ~\new_[7402]_ ;
  assign n4090 = ~\new_[7456]_  | ~\new_[7334]_ ;
  assign n4075 = ~\new_[7451]_  | ~\new_[7211]_ ;
  assign n3950 = ~\new_[7482]_  | ~\new_[7242]_ ;
  assign n3910 = ~\new_[7462]_  | ~\new_[7358]_ ;
  assign n4010 = ~\new_[7448]_  | ~\new_[7362]_ ;
  assign n3805 = ~\new_[7537]_  | ~\new_[7233]_ ;
  assign n4060 = ~\new_[7500]_  | ~\new_[7345]_ ;
  assign n3890 = ~\new_[7535]_  | ~\new_[7363]_ ;
  assign n3920 = ~\new_[7540]_  | ~\new_[7221]_ ;
  assign n4100 = ~\new_[7438]_  | ~\new_[7240]_ ;
  assign n3795 = ~\new_[7454]_  | ~\new_[7324]_ ;
  assign n4055 = ~\new_[7430]_  | ~\new_[7215]_ ;
  assign n3980 = ~\new_[7544]_  | ~\new_[7371]_ ;
  assign n3945 = ~\new_[7539]_  | ~\new_[7401]_ ;
  assign n3880 = ~\new_[7549]_  | ~\new_[7243]_ ;
  assign n3785 = ~\new_[7523]_  | ~\new_[7325]_ ;
  assign n3870 = ~\new_[7538]_  | ~\new_[7293]_ ;
  assign n3935 = ~\new_[7477]_  | ~\new_[7394]_ ;
  assign \new_[7006]_  = \new_[3257]_  ? \new_[8935]_  : \data_o[10] ;
  assign \new_[7007]_  = \new_[6599]_  ? \new_[8894]_  : \data_o[123] ;
  assign \new_[7008]_  = \new_[3106]_  ? \new_[8893]_  : \data_o[25] ;
  assign \new_[7009]_  = \new_[6746]_  ? \new_[8900]_  : \data_o[95] ;
  assign \new_[7010]_  = \new_[6606]_  ? \new_[8893]_  : \data_o[101] ;
  assign \new_[7011]_  = (~\new_[1207]_  | ~\new_[7738]_ ) & (~\new_[1221]_  | ~\new_[7569]_ );
  assign \new_[7012]_  = \new_[6591]_  ? \new_[8946]_  : \data_o[36] ;
  assign \new_[7013]_  = \new_[3387]_  ? \new_[8935]_  : \data_o[16] ;
  assign \new_[7014]_  = \new_[6585]_  ? \new_[8894]_  : \data_o[84] ;
  assign \new_[7015]_  = \new_[6429]_  ? \new_[8918]_  : \data_o[82] ;
  assign \new_[7016]_  = \new_[3386]_  ? \new_[8920]_  : \data_o[30] ;
  assign \new_[7017]_  = \new_[6590]_  ? \new_[8927]_  : \data_o[125] ;
  assign \new_[7018]_  = \new_[6450]_  ? \new_[8927]_  : \data_o[77] ;
  assign \new_[7019]_  = \new_[3383]_  ? \new_[8894]_  : \data_o[21] ;
  assign \new_[7020]_  = \new_[6593]_  ? \new_[8940]_  : \data_o[55] ;
  assign \new_[7021]_  = \new_[3885]_  ? \new_[8894]_  : \data_o[15] ;
  assign \new_[7022]_  = \new_[6444]_  ? \new_[8893]_  : \data_o[33] ;
  assign \new_[7023]_  = \new_[3857]_  ? \new_[8946]_  : \data_o[23] ;
  assign \new_[7024]_  = \new_[3443]_  ? \new_[8902]_  : \data_o[24] ;
  assign \new_[7025]_  = \new_[6723]_  ? \new_[8940]_  : \data_o[127] ;
  assign \new_[7026]_  = \new_[6592]_  ? \new_[8902]_  : \data_o[39] ;
  assign \new_[7027]_  = ~\new_[6607]_  | ~\new_[8925]_ ;
  assign \new_[7028]_  = ~\new_[6704]_  | ~\new_[8919]_ ;
  assign \new_[7029]_  = ~\new_[6632]_  | ~\new_[8905]_ ;
  assign \new_[7030]_  = ~\new_[6443]_  | ~\new_[8905]_ ;
  assign \new_[7031]_  = ~\new_[8900]_  | ~\data_o[113] ;
  assign \new_[7032]_  = ~\new_[8900]_  | ~\data_o[116] ;
  assign \new_[7033]_  = (~\new_[1238]_  | ~\new_[7738]_ ) & (~\new_[1202]_  | ~\new_[7632]_ );
  assign n4030 = ~\new_[7450]_  | ~\new_[7283]_ ;
  assign \new_[7035]_  = ~\new_[8918]_  | ~\data_o[118] ;
  assign \new_[7036]_  = \new_[6639]_  ? \new_[8943]_  : \data_o[120] ;
  assign \new_[7037]_  = \new_[2349]_  ? \new_[7660]_  : \key_i[98] ;
  assign \new_[7038]_  = ~\new_[8900]_  | ~\data_o[114] ;
  assign \new_[7039]_  = (~\new_[7660]_  | ~\key_i[85] ) & (~\new_[7581]_  | ~\new_[2201]_ );
  assign \new_[7040]_  = (~\new_[7660]_  | ~\key_i[92] ) & (~\new_[7582]_  | ~\new_[8151]_ );
  assign \new_[7041]_  = \key_i[79]  ? \new_[7582]_  : \new_[1141]_ ;
  assign \new_[7042]_  = (~\new_[7660]_  | ~\key_i[110] ) & (~\new_[7769]_  | ~\new_[1455]_ );
  assign n3845 = ~\new_[7444]_  | ~\new_[7354]_ ;
  assign \new_[7044]_  = \key_i[112]  ? \new_[7620]_  : \new_[2421]_ ;
  assign \new_[7045]_  = \key_i[96]  ? \new_[7620]_  : \new_[2348]_ ;
  assign \new_[7046]_  = \key_i[113]  ? \new_[7620]_  : \new_[2411]_ ;
  assign \new_[7047]_  = \key_i[76]  ? \new_[7582]_  : \new_[1125]_ ;
  assign \new_[7048]_  = (~\new_[7660]_  | ~\key_i[84] ) & (~\new_[7581]_  | ~\new_[2200]_ );
  assign \new_[7049]_  = (~\new_[7660]_  | ~\key_i[109] ) & (~\new_[7581]_  | ~\new_[1456]_ );
  assign \new_[7050]_  = \key_i[117]  ? \new_[7620]_  : \new_[2461]_ ;
  assign \new_[7051]_  = (~\new_[7660]_  | ~\key_i[64] ) & (~\new_[7581]_  | ~\new_[2132]_ );
  assign \new_[7052]_  = \key_i[114]  ? \new_[7620]_  : \new_[2424]_ ;
  assign \new_[7053]_  = (~\new_[7660]_  | ~\key_i[86] ) & (~\new_[7581]_  | ~\new_[2203]_ );
  assign \new_[7054]_  = \key_i[78]  ? \new_[7582]_  : \new_[1133]_ ;
  assign \new_[7055]_  = (~\new_[7660]_  | ~\key_i[83] ) & (~\new_[7581]_  | ~\new_[2199]_ );
  assign \new_[7056]_  = \new_[6428]_  ? \new_[8900]_  : \data_o[98] ;
  assign n3965 = ~\new_[7408]_  | ~\new_[7285]_ ;
  assign \new_[7058]_  = \key_i[97]  ? \new_[7620]_  : \new_[2344]_ ;
  assign \new_[7059]_  = (~\new_[7660]_  | ~\key_i[65] ) & (~\new_[7581]_  | ~\new_[2133]_ );
  assign \new_[7060]_  = (~\new_[7660]_  | ~\key_i[87] ) & (~\new_[7581]_  | ~\new_[2139]_ );
  assign \new_[7061]_  = \key_i[75]  ? \new_[7582]_  : \new_[1126]_ ;
  assign \new_[7062]_  = ~\new_[8343]_  | ~\new_[8130]_ ;
  assign \new_[7063]_  = (~\new_[1234]_  | ~\new_[7738]_ ) & (~\new_[1214]_  | ~\new_[7632]_ );
  assign \new_[7064]_  = (~\new_[1212]_  | ~\new_[7738]_ ) & (~\new_[1204]_  | ~\new_[7632]_ );
  assign \new_[7065]_  = \new_[1103]_  ? \new_[7738]_  : \new_[1108]_ ;
  assign n3860 = ~\new_[7413]_  | ~\new_[7255]_ ;
  assign \new_[7067]_  = \new_[1110]_  ? \new_[7738]_  : \new_[1105]_ ;
  assign \new_[7068]_  = (~\new_[1461]_  | ~\new_[7738]_ ) & (~\new_[1520]_  | ~\new_[7632]_ );
  assign \new_[7069]_  = (~\new_[1148]_  | ~\new_[7738]_ ) & (~\new_[1150]_  | ~\new_[7632]_ );
  assign \new_[7070]_  = (~\new_[1381]_  | ~\new_[7738]_ ) & (~\new_[1324]_  | ~\new_[7569]_ );
  assign \new_[7071]_  = (~\new_[1209]_  | ~\new_[7632]_ ) & (~\new_[1151]_  | ~\new_[7738]_ );
  assign \new_[7072]_  = (~\new_[1211]_  | ~\new_[7738]_ ) & (~\new_[1203]_  | ~\new_[7632]_ );
  assign \new_[7073]_  = (~\new_[1213]_  | ~\new_[7738]_ ) & (~\new_[1205]_  | ~\new_[7569]_ );
  assign \new_[7074]_  = \new_[1106]_  ? \new_[7738]_  : \new_[1116]_ ;
  assign \new_[7075]_  = ~\new_[7660]_ ;
  assign \new_[7076]_  = (~\new_[1152]_  | ~\new_[7738]_ ) & (~\new_[1147]_  | ~\new_[7632]_ );
  assign \new_[7077]_  = (~\new_[1209]_  | ~\new_[7738]_ ) & (~\new_[1151]_  | ~\new_[7569]_ );
  assign \new_[7078]_  = (~\new_[1237]_  | ~\new_[7738]_ ) & (~\new_[1240]_  | ~\new_[7569]_ );
  assign \new_[7079]_  = \new_[1111]_  ? \new_[7738]_  : \new_[1104]_ ;
  assign \new_[7080]_  = (~\new_[1206]_  | ~\new_[7738]_ ) & (~\new_[1220]_  | ~\new_[7632]_ );
  assign \new_[7081]_  = (~\new_[1206]_  | ~\new_[7632]_ ) & (~\new_[1220]_  | ~\new_[7738]_ );
  assign \new_[7082]_  = (~\new_[1521]_  | ~\new_[7738]_ ) & (~\new_[1530]_  | ~\new_[7632]_ );
  assign \new_[7083]_  = \new_[6432]_  ? \new_[8921]_  : \data_o[72] ;
  assign \new_[7084]_  = \new_[1102]_  ? \new_[7738]_  : \new_[1109]_ ;
  assign \new_[7085]_  = \new_[6630]_  ? \new_[8944]_  : \data_o[75] ;
  assign \new_[7086]_  = \new_[3105]_  ? \new_[8946]_  : \data_o[1] ;
  assign \new_[7087]_  = \new_[6626]_  ? \new_[8894]_  : \data_o[54] ;
  assign \new_[7088]_  = \new_[6666]_  ? \new_[8946]_  : \data_o[92] ;
  assign \new_[7089]_  = \key_i[126]  ? \new_[7620]_  : \new_[2271]_ ;
  assign \new_[7090]_  = ~\new_[8133]_  | ~n4110;
  assign \new_[7091]_  = ~\new_[8063]_  | ~n4110;
  assign \new_[7092]_  = \key_i[106]  ? \new_[7769]_  : \new_[8075]_ ;
  assign \new_[7093]_  = \new_[6663]_  ? \new_[8946]_  : \data_o[121] ;
  assign \new_[7094]_  = \key_i[108]  ? \new_[7620]_  : \new_[8004]_ ;
  assign \new_[7095]_  = \key_i[118]  ? \new_[7582]_  : \new_[2425]_ ;
  assign \new_[7096]_  = \new_[6571]_  ? \new_[8921]_  : \data_o[126] ;
  assign \new_[7097]_  = ~\new_[7239]_ ;
  assign \new_[7098]_  = ~\new_[6652]_  | ~\new_[8945]_ ;
  assign \new_[7099]_  = ~\new_[6589]_  | ~\new_[8925]_ ;
  assign \new_[7100]_  = \key_i[116]  ? \new_[7582]_  : \new_[2423]_ ;
  assign \new_[7101]_  = \new_[6426]_  ? \new_[8902]_  : \data_o[70] ;
  assign \new_[7102]_  = ~\new_[7488]_  | ~\new_[8237]_ ;
  assign \new_[7103]_  = \key_i[107]  ? \new_[7620]_  : \new_[7971]_ ;
  assign \new_[7104]_  = \new_[3515]_  ? \new_[8893]_  : \data_o[5] ;
  assign \new_[7105]_  = \new_[6605]_  ? \new_[8920]_  : \data_o[68] ;
  assign \new_[7106]_  = \new_[3108]_  ? \new_[8940]_  : \data_o[9] ;
  assign \new_[7107]_  = \new_[6442]_  ? \new_[8904]_  : \data_o[69] ;
  assign \new_[7108]_  = ~\new_[7998]_  | ~n4110;
  assign \new_[7109]_  = ~\new_[8030]_  | ~n4110;
  assign \new_[7110]_  = ~\new_[6547]_  | ~\new_[8939]_ ;
  assign \new_[7111]_  = \key_i[99]  ? \new_[7620]_  : \new_[2537]_ ;
  assign \new_[7112]_  = \key_i[115]  ? \new_[7582]_  : \new_[2422]_ ;
  assign \new_[7113]_  = ~\new_[7486]_  | ~\new_[1070]_ ;
  assign \new_[7114]_  = ~\new_[7261]_ ;
  assign \new_[7115]_  = ~\new_[7260]_ ;
  assign \new_[7116]_  = ~\new_[7261]_ ;
  assign \new_[7117]_  = ~\new_[7622]_  | ~\new_[7472]_ ;
  assign \new_[7118]_  = ~\new_[7491]_  | ~\new_[7467]_ ;
  assign \new_[7119]_  = \key_i[101]  ? \new_[7582]_  : \new_[2351]_ ;
  assign \new_[7120]_  = ~\new_[7603]_  | ~\new_[1149]_ ;
  assign \new_[7121]_  = ~\new_[7486]_  | ~\new_[1064]_ ;
  assign \new_[7122]_  = ~\new_[7579]_  | ~\new_[7412]_ ;
  assign \new_[7123]_  = ~\new_[7849]_  & (~\new_[8947]_  | ~\new_[2426]_ );
  assign \new_[7124]_  = \new_[3109]_  ? \new_[8893]_  : \data_o[2] ;
  assign \new_[7125]_  = \new_[6495]_  ? \new_[8940]_  : \data_o[64] ;
  assign \new_[7126]_  = \new_[6438]_  ? \new_[8946]_  : \data_o[91] ;
  assign \new_[7127]_  = \new_[6568]_  ? \new_[8893]_  : \data_o[88] ;
  assign \new_[7128]_  = \new_[6640]_  ? \new_[8940]_  : \data_o[40] ;
  assign \new_[7129]_  = \new_[6433]_  ? \new_[8893]_  : \data_o[48] ;
  assign \new_[7130]_  = \new_[6424]_  ? \new_[8946]_  : \data_o[45] ;
  assign \new_[7131]_  = ~\new_[7577]_  | ~\new_[7467]_  | ~\new_[7841]_ ;
  assign \new_[7132]_  = \new_[3406]_  ? \new_[8921]_  : \data_o[6] ;
  assign \new_[7133]_  = \new_[6616]_  ? \new_[8904]_  : \data_o[51] ;
  assign \new_[7134]_  = \new_[3385]_  ? \new_[8940]_  : \data_o[22] ;
  assign \new_[7135]_  = \new_[6716]_  ? \new_[8894]_  : \data_o[73] ;
  assign \new_[7136]_  = \new_[6425]_  ? \new_[8904]_  : \data_o[67] ;
  assign \new_[7137]_  = \new_[6618]_  ? \new_[8940]_  : \data_o[66] ;
  assign \new_[7138]_  = ~\new_[7260]_ ;
  assign \new_[7139]_  = ~\new_[8900]_  | ~\data_o[63] ;
  assign \new_[7140]_  = \key_i[100]  ? \new_[7582]_  : \new_[2350]_ ;
  assign \new_[7141]_  = \key_i[111]  ? \new_[7769]_  : \new_[7984]_ ;
  assign \new_[7142]_  = \key_i[103]  ? \new_[7582]_  : \new_[2353]_ ;
  assign \new_[7143]_  = \key_i[104]  ? \new_[7582]_  : \new_[7949]_ ;
  assign \new_[7144]_  = \key_i[119]  ? \new_[7582]_  : \new_[2354]_ ;
  assign \new_[7145]_  = \key_i[123]  ? \new_[7620]_  : \new_[2197]_ ;
  assign \new_[7146]_  = (~\new_[7660]_  | ~\key_i[124] ) & (~\new_[7620]_  | ~\new_[2131]_ );
  assign \new_[7147]_  = \key_i[125]  ? \new_[7620]_  : \new_[2196]_ ;
  assign \new_[7148]_  = \key_i[105]  ? \new_[7769]_  : \new_[7986]_ ;
  assign \new_[7149]_  = \key_i[102]  ? \new_[7582]_  : \new_[2352]_ ;
  assign \new_[7150]_  = ~\new_[8100]_  | ~n4110;
  assign \new_[7151]_  = ~\new_[7603]_  | ~\new_[1097]_ ;
  assign \new_[7152]_  = ~\new_[8019]_  | ~n4110;
  assign \new_[7153]_  = ~\new_[7603]_  | ~\new_[1213]_ ;
  assign \new_[7154]_  = ~\new_[8081]_  | ~n4110;
  assign \new_[7155]_  = ~\new_[8010]_  | ~n4110;
  assign \new_[7156]_  = ~\new_[7603]_  | ~\new_[1190]_ ;
  assign \new_[7157]_  = ~\new_[8090]_  | ~n4110;
  assign \new_[7158]_  = ~\new_[8085]_  | ~n4110;
  assign \new_[7159]_  = ~\new_[7592]_  | ~\new_[7939]_ ;
  assign \new_[7160]_  = ~\new_[7603]_  | ~\new_[1217]_ ;
  assign \new_[7161]_  = ~\new_[7592]_  | ~\new_[1311]_ ;
  assign \new_[7162]_  = ~\new_[8092]_  | ~n4110;
  assign \new_[7163]_  = ~\new_[8040]_  | ~n4110;
  assign \new_[7164]_  = ~\new_[8062]_  | ~n4110;
  assign \new_[7165]_  = ~\new_[7948]_  | ~n4110;
  assign \new_[7166]_  = ~\new_[8110]_  | ~n4110;
  assign \new_[7167]_  = ~\new_[7584]_  | ~\new_[1460]_ ;
  assign \new_[7168]_  = ~\new_[7603]_  | ~\new_[1187]_ ;
  assign \new_[7169]_  = ~\new_[7603]_  | ~\new_[1148]_ ;
  assign \new_[7170]_  = ~\new_[7603]_  | ~\new_[1240]_ ;
  assign \new_[7171]_  = ~\new_[8468]_  | ~n4110;
  assign \new_[7172]_  = ~\new_[7603]_  | ~\new_[1147]_ ;
  assign \new_[7173]_  = ~\new_[8025]_  | ~n4110;
  assign \new_[7174]_  = ~\new_[7603]_  | ~\new_[1312]_ ;
  assign \new_[7175]_  = ~\new_[7603]_  | ~\new_[1319]_ ;
  assign \new_[7176]_  = ~\new_[7603]_  | ~\new_[1202]_ ;
  assign \new_[7177]_  = ~\new_[8088]_  | ~n4110;
  assign \new_[7178]_  = ~\new_[7603]_  | ~\new_[1103]_ ;
  assign \new_[7179]_  = ~\new_[8147]_  | ~n4110;
  assign \new_[7180]_  = ~\new_[8590]_  | ~n4110;
  assign \new_[7181]_  = ~\new_[7603]_  | ~\new_[1204]_ ;
  assign \new_[7182]_  = ~\new_[7603]_  | ~\new_[1137]_ ;
  assign \new_[7183]_  = ~\new_[8136]_  | ~n4110;
  assign \new_[7184]_  = ~\new_[8478]_  | ~n4110;
  assign \new_[7185]_  = ~\new_[8102]_  | ~n4110;
  assign \new_[7186]_  = ~\new_[8016]_  | ~n4110;
  assign \new_[7187]_  = ~\new_[7603]_  | ~\new_[1223]_ ;
  assign \new_[7188]_  = ~\new_[8127]_  | ~n4110;
  assign \new_[7189]_  = ~\new_[8043]_  | ~n4110;
  assign \new_[7190]_  = ~\new_[7603]_  | ~\new_[1112]_ ;
  assign \new_[7191]_  = ~\new_[8067]_  | ~n4110;
  assign \new_[7192]_  = ~\new_[7603]_  | ~\new_[1251]_ ;
  assign \new_[7193]_  = ~\new_[7592]_  | ~\new_[1194]_ ;
  assign \new_[7194]_  = ~\new_[7992]_  | ~n4110;
  assign \new_[7195]_  = ~\new_[8070]_  | ~n4110;
  assign \new_[7196]_  = ~\new_[7264]_ ;
  assign \new_[7197]_  = ~\new_[8036]_  | ~n4110;
  assign \new_[7198]_  = ~\new_[8042]_  | ~n4110;
  assign \new_[7199]_  = ~\new_[8035]_  | ~n4110;
  assign \new_[7200]_  = ~\new_[7603]_  | ~\new_[1192]_ ;
  assign \new_[7201]_  = \new_[6628]_  ? \new_[8893]_  : \data_o[124] ;
  assign \new_[7202]_  = ~\new_[7592]_  | ~\new_[1096]_ ;
  assign \new_[7203]_  = ~\new_[7603]_  | ~\new_[1237]_ ;
  assign \new_[7204]_  = ~\new_[7603]_  | ~\new_[1234]_ ;
  assign \new_[7205]_  = ~\new_[7603]_  | ~\new_[1521]_ ;
  assign \new_[7206]_  = ~\new_[7406]_ ;
  assign \new_[7207]_  = ~\new_[7623]_  | ~\new_[1212]_ ;
  assign \new_[7208]_  = ~\new_[7603]_  | ~\new_[1100]_ ;
  assign \new_[7209]_  = ~\new_[7623]_  | ~\new_[1459]_ ;
  assign \new_[7210]_  = ~\new_[7603]_  | ~\new_[1113]_ ;
  assign \new_[7211]_  = ~\new_[7940]_  | ~n4110;
  assign \new_[7212]_  = ~\new_[8091]_  | ~n4110;
  assign \new_[7213]_  = \new_[3103]_  ? \new_[8920]_  : \data_o[17] ;
  assign \new_[7214]_  = ~\new_[7623]_  | ~\new_[1222]_ ;
  assign \new_[7215]_  = ~\new_[8002]_  | ~n4110;
  assign \new_[7216]_  = ~\new_[7623]_  | ~\new_[1102]_ ;
  assign \new_[7217]_  = \new_[6656]_  ? \new_[8920]_  : \data_o[41] ;
  assign \new_[7218]_  = \new_[6573]_  ? \new_[8904]_  : \data_o[74] ;
  assign \new_[7219]_  = ~\new_[7603]_  | ~\new_[1191]_ ;
  assign \new_[7220]_  = ~\new_[8155]_  | ~n4110;
  assign \new_[7221]_  = ~\new_[8066]_  | ~n4110;
  assign \new_[7222]_  = \new_[6609]_  ? \new_[8894]_  : \data_o[52] ;
  assign \new_[7223]_  = ~\new_[7623]_  | ~\new_[1464]_ ;
  assign \new_[7224]_  = ~\new_[7623]_  | ~\new_[1458]_ ;
  assign \new_[7225]_  = ~\new_[8126]_  | ~n4110;
  assign \new_[7226]_  = ~\new_[8463]_  | ~n4110;
  assign \new_[7227]_  = ~\new_[7603]_  | ~\new_[1095]_ ;
  assign \new_[7228]_  = ~\new_[7623]_  | ~\new_[1323]_ ;
  assign \new_[7229]_  = ~\new_[7603]_  | ~\new_[1197]_ ;
  assign \new_[7230]_  = ~\new_[7623]_  | ~\new_[1200]_ ;
  assign \new_[7231]_  = ~\new_[7623]_  | ~\new_[1114]_ ;
  assign \new_[7232]_  = ~\new_[7623]_  | ~\new_[8020]_ ;
  assign \new_[7233]_  = ~\new_[8087]_  | ~n4110;
  assign \new_[7234]_  = ~\new_[7623]_  | ~\new_[1245]_ ;
  assign \new_[7235]_  = ~\new_[7623]_  | ~\new_[1463]_ ;
  assign \new_[7236]_  = ~\new_[7623]_  | ~\new_[1226]_ ;
  assign \new_[7237]_  = ~\new_[7584]_  | ~\new_[1457]_ ;
  assign \new_[7238]_  = ~\new_[8437]_  | ~n4110;
  assign \new_[7239]_  = ~\new_[7563]_  & (~\new_[8238]_  | ~\new_[8237]_ );
  assign \new_[7240]_  = ~\new_[7960]_  | ~n4110;
  assign \new_[7241]_  = ~\new_[7623]_  | ~\new_[1241]_ ;
  assign \new_[7242]_  = ~\new_[8129]_  | ~n4110;
  assign \new_[7243]_  = ~\new_[8015]_  | ~n4110;
  assign \new_[7244]_  = \new_[6445]_  ? \new_[8894]_  : \data_o[65] ;
  assign \new_[7245]_  = \new_[6627]_  ? \new_[8894]_  : \data_o[50] ;
  assign \new_[7246]_  = \new_[6451]_  ? \new_[8904]_  : \data_o[78] ;
  assign \new_[7247]_  = ~\new_[8144]_  | ~n4110;
  assign \new_[7248]_  = \new_[6624]_  ? \new_[8920]_  : \data_o[42] ;
  assign \new_[7249]_  = ~\new_[7978]_  | ~n4110;
  assign \new_[7250]_  = ~\new_[7688]_  | ~\new_[7614]_  | ~\new_[7862]_ ;
  assign \new_[7251]_  = ~\new_[7623]_  | ~\new_[1104]_ ;
  assign \new_[7252]_  = \new_[6546]_  ? \new_[8920]_  : \data_o[49] ;
  assign \new_[7253]_  = ~\new_[8152]_  | ~n4110;
  assign \new_[7254]_  = ~\new_[7623]_  | ~\new_[1117]_ ;
  assign \new_[7255]_  = ~\new_[8114]_  | ~n4110;
  assign \new_[7256]_  = \new_[2758]_  ? \new_[8920]_  : \data_o[4] ;
  assign \new_[7257]_  = ~\new_[8112]_  | ~n4110;
  assign \new_[7258]_  = ~\new_[8054]_  | ~n4110;
  assign \new_[7259]_  = ~\new_[7427]_ ;
  assign \new_[7260]_  = ~\new_[7563]_  & (~\new_[7894]_  | ~\new_[7668]_ );
  assign \new_[7261]_  = ~\new_[7604]_ ;
  assign \new_[7262]_  = ~\new_[7623]_  | ~\new_[1116]_ ;
  assign \new_[7263]_  = ~\new_[7623]_  | ~\new_[1381]_ ;
  assign \new_[7264]_  = \new_[7577]_  & \new_[7934]_ ;
  assign \new_[7265]_  = ~\new_[7472]_ ;
  assign \new_[7266]_  = ~\new_[7412]_ ;
  assign \new_[7267]_  = ~\new_[7623]_  | ~\new_[1246]_ ;
  assign \new_[7268]_  = \new_[6597]_  ? \new_[8946]_  : \data_o[46] ;
  assign \new_[7269]_  = ~\new_[7571]_  | ~\new_[6771]_ ;
  assign \new_[7270]_  = ~\new_[7480]_ ;
  assign \new_[7271]_  = ~\new_[7623]_  | ~\new_[1108]_ ;
  assign \new_[7272]_  = \new_[6625]_  ? \new_[8902]_  : \data_o[94] ;
  assign \new_[7273]_  = \new_[6569]_  ? \new_[8920]_  : \data_o[89] ;
  assign \new_[7274]_  = \new_[3410]_  ? \new_[8943]_  : \data_o[0] ;
  assign \new_[7275]_  = \new_[2870]_  ? \new_[8893]_  : \data_o[3] ;
  assign \new_[7276]_  = \new_[3104]_  ? \new_[8902]_  : \data_o[18] ;
  assign \new_[7277]_  = \new_[6572]_  ? \new_[8893]_  : \data_o[90] ;
  assign \new_[7278]_  = \new_[6452]_  ? \new_[8935]_  : \data_o[122] ;
  assign \new_[7279]_  = \new_[6581]_  ? \new_[8920]_  : \data_o[76] ;
  assign \new_[7280]_  = \new_[2756]_  ? \new_[8902]_  : \data_o[20] ;
  assign \new_[7281]_  = \new_[6448]_  ? \new_[8894]_  : \data_o[93] ;
  assign \new_[7282]_  = ~\new_[7603]_  | ~\new_[1383]_ ;
  assign \new_[7283]_  = ~\new_[8099]_  | ~n4110;
  assign \new_[7284]_  = ~\new_[7623]_  | ~\new_[1324]_ ;
  assign \new_[7285]_  = ~\new_[8093]_  | ~n4110;
  assign \new_[7286]_  = ~\new_[7623]_  | ~\new_[1538]_ ;
  assign \new_[7287]_  = ~\new_[7603]_  | ~\new_[1244]_ ;
  assign \new_[7288]_  = ~\new_[7945]_  | ~n4110;
  assign \new_[7289]_  = ~\new_[8116]_  | ~n4110;
  assign \new_[7290]_  = ~\new_[7623]_  | ~\new_[1110]_ ;
  assign \new_[7291]_  = ~\new_[7623]_  | ~\new_[1461]_ ;
  assign \new_[7292]_  = ~\new_[7603]_  | ~\new_[1136]_ ;
  assign \new_[7293]_  = ~\new_[8132]_  | ~n4110;
  assign \new_[7294]_  = ~\new_[7623]_  | ~\new_[1219]_ ;
  assign \new_[7295]_  = ~\new_[7623]_  | ~\new_[1105]_ ;
  assign \new_[7296]_  = ~\new_[7623]_  | ~\new_[1322]_ ;
  assign \new_[7297]_  = ~\new_[7623]_  | ~\new_[1320]_ ;
  assign \new_[7298]_  = ~\new_[7623]_  | ~\new_[1530]_ ;
  assign \new_[7299]_  = ~\new_[7623]_  | ~\new_[1208]_ ;
  assign \new_[7300]_  = ~\new_[7623]_  | ~\new_[1249]_ ;
  assign \new_[7301]_  = ~\new_[7623]_  | ~\new_[1206]_ ;
  assign \new_[7302]_  = ~\new_[7584]_  | ~\new_[1220]_ ;
  assign \new_[7303]_  = ~\new_[7603]_  | ~\new_[1384]_ ;
  assign \new_[7304]_  = ~\new_[7623]_  | ~\new_[1221]_ ;
  assign \new_[7305]_  = ~\new_[7623]_  | ~\new_[1247]_ ;
  assign \new_[7306]_  = ~\new_[7623]_  | ~\new_[8068]_ ;
  assign \new_[7307]_  = ~\new_[8118]_  | ~n4110;
  assign \new_[7308]_  = ~\new_[7584]_  | ~\new_[1211]_ ;
  assign \new_[7309]_  = ~\new_[8007]_  | ~n4110;
  assign \new_[7310]_  = ~\new_[7623]_  | ~\new_[1134]_ ;
  assign \new_[7311]_  = ~\new_[7623]_  | ~\new_[1215]_ ;
  assign \new_[7312]_  = ~\new_[7623]_  | ~\new_[1196]_ ;
  assign \new_[7313]_  = ~\new_[7603]_  | ~\new_[8053]_ ;
  assign \new_[7314]_  = ~\new_[7623]_  | ~\new_[1205]_ ;
  assign \new_[7315]_  = ~\new_[7603]_  | ~\new_[8026]_ ;
  assign \new_[7316]_  = ~\new_[8143]_  | ~n4110;
  assign \new_[7317]_  = ~\new_[7972]_  | ~n4110;
  assign \new_[7318]_  = ~\new_[8082]_  | ~n4110;
  assign \new_[7319]_  = ~\new_[7623]_  | ~\new_[1313]_ ;
  assign \new_[7320]_  = ~\new_[7603]_  | ~\new_[1135]_ ;
  assign \new_[7321]_  = ~\new_[7623]_  | ~\new_[1207]_ ;
  assign \new_[7322]_  = ~\new_[7623]_  | ~\new_[1315]_ ;
  assign \new_[7323]_  = ~\new_[7603]_  | ~\new_[1094]_ ;
  assign \new_[7324]_  = ~\new_[7938]_  | ~n4110;
  assign \new_[7325]_  = ~\new_[7966]_  | ~n4110;
  assign \new_[7326]_  = ~\new_[8074]_  | ~n4110;
  assign \new_[7327]_  = ~\new_[7623]_  | ~\new_[1209]_ ;
  assign \new_[7328]_  = ~\new_[7977]_  | ~n4110;
  assign \new_[7329]_  = ~\new_[7603]_  | ~\new_[1248]_ ;
  assign \new_[7330]_  = ~\new_[7603]_  | ~\new_[1186]_ ;
  assign \new_[7331]_  = ~\new_[8145]_  | ~n4110;
  assign \new_[7332]_  = ~\new_[7623]_  | ~\new_[1198]_ ;
  assign \new_[7333]_  = ~\new_[7623]_  | ~\new_[1150]_ ;
  assign \new_[7334]_  = ~\new_[7956]_  | ~n4110;
  assign \new_[7335]_  = ~\new_[7974]_  | ~n4110;
  assign \new_[7336]_  = ~\new_[8069]_  | ~n4110;
  assign \new_[7337]_  = ~\new_[8076]_  | ~n4110;
  assign \new_[7338]_  = ~\new_[7584]_  | ~\new_[1106]_ ;
  assign \new_[7339]_  = ~\new_[7603]_  | ~\new_[8101]_ ;
  assign \new_[7340]_  = ~\new_[8032]_  | ~n4110;
  assign \new_[7341]_  = ~\new_[7603]_  | ~\new_[1193]_ ;
  assign \new_[7342]_  = ~\new_[8003]_  | ~n4110;
  assign \new_[7343]_  = ~\new_[8021]_  | ~n4110;
  assign \new_[7344]_  = ~\new_[8059]_  | ~n4110;
  assign \new_[7345]_  = ~\new_[7981]_  | ~n4110;
  assign \new_[7346]_  = ~\new_[7942]_  | ~n4110;
  assign \new_[7347]_  = ~\new_[7623]_  | ~\new_[1139]_ ;
  assign \new_[7348]_  = ~\new_[7603]_  | ~\new_[1250]_ ;
  assign \new_[7349]_  = ~\new_[7603]_  | ~\new_[1143]_ ;
  assign \new_[7350]_  = ~\new_[7603]_  | ~\new_[1386]_ ;
  assign \new_[7351]_  = ~\new_[7603]_  | ~\new_[1210]_ ;
  assign \new_[7352]_  = ~\new_[8104]_  | ~n4110;
  assign \new_[7353]_  = ~\new_[7603]_  | ~\new_[1101]_ ;
  assign \new_[7354]_  = ~\new_[7985]_  | ~n4110;
  assign \new_[7355]_  = ~\new_[8089]_  | ~n4110;
  assign \new_[7356]_  = ~\new_[7603]_  | ~\new_[1138]_ ;
  assign \new_[7357]_  = ~\new_[7623]_  | ~\new_[1385]_ ;
  assign \new_[7358]_  = ~\new_[8048]_  | ~n4110;
  assign \new_[7359]_  = ~\new_[7623]_  | ~\new_[1151]_ ;
  assign \new_[7360]_  = ~\new_[8065]_  | ~n4110;
  assign \new_[7361]_  = ~\new_[7623]_  | ~\new_[1238]_ ;
  assign \new_[7362]_  = ~\new_[8080]_  | ~n4110;
  assign \new_[7363]_  = ~\new_[7969]_  | ~n4110;
  assign \new_[7364]_  = ~\new_[7623]_  | ~\new_[1321]_ ;
  assign \new_[7365]_  = ~\new_[7623]_  | ~\new_[1216]_ ;
  assign \new_[7366]_  = ~\new_[7603]_  | ~\new_[1201]_ ;
  assign \new_[7367]_  = ~\new_[7976]_  | ~n4110;
  assign \new_[7368]_  = ~\new_[8073]_  | ~n4110;
  assign \new_[7369]_  = ~\new_[8033]_  | ~n4110;
  assign \new_[7370]_  = ~\new_[7623]_  | ~\new_[1203]_ ;
  assign \new_[7371]_  = ~\new_[8061]_  | ~n4110;
  assign \new_[7372]_  = ~\new_[7623]_  | ~\new_[1115]_ ;
  assign \new_[7373]_  = ~\new_[7603]_  | ~\new_[1242]_ ;
  assign \new_[7374]_  = ~\new_[7623]_  | ~\new_[1520]_ ;
  assign \new_[7375]_  = ~\new_[8149]_  | ~n4110;
  assign \new_[7376]_  = ~\new_[8044]_  | ~n4110;
  assign \new_[7377]_  = ~\new_[7623]_  | ~\new_[1144]_ ;
  assign \new_[7378]_  = ~\new_[7603]_  | ~\new_[1098]_ ;
  assign \new_[7379]_  = ~\new_[7623]_  | ~\new_[1109]_ ;
  assign \new_[7380]_  = ~\new_[8117]_  | ~n4110;
  assign \new_[7381]_  = ~\new_[7988]_  | ~n4110;
  assign \new_[7382]_  = ~\new_[7983]_  | ~n4110;
  assign \new_[7383]_  = ~\new_[7623]_  | ~\new_[1252]_ ;
  assign \new_[7384]_  = ~\new_[7410]_ ;
  assign \new_[7385]_  = ~\new_[7603]_  | ~\new_[1199]_ ;
  assign \new_[7386]_  = ~\new_[7603]_  | ~\new_[1243]_ ;
  assign \new_[7387]_  = ~\new_[7603]_  | ~\new_[1314]_ ;
  assign \new_[7388]_  = ~\new_[8128]_  | ~n4110;
  assign \new_[7389]_  = ~\new_[7623]_  | ~\new_[1111]_ ;
  assign \new_[7390]_  = ~\new_[7603]_  | ~\new_[1225]_ ;
  assign \new_[7391]_  = ~\new_[7623]_  | ~\new_[1224]_ ;
  assign \new_[7392]_  = ~\new_[7603]_  | ~\new_[1195]_ ;
  assign \new_[7393]_  = \new_[6580]_  ? \new_[8893]_  : \data_o[43] ;
  assign \new_[7394]_  = ~\new_[8154]_  | ~n4110;
  assign \new_[7395]_  = ~\new_[7623]_  | ~\new_[1142]_ ;
  assign \new_[7396]_  = \new_[6623]_  ? \new_[8920]_  : \data_o[44] ;
  assign \new_[7397]_  = ~\new_[7603]_  | ~\new_[1145]_ ;
  assign \new_[7398]_  = ~\new_[7623]_  | ~\new_[1107]_ ;
  assign \new_[7399]_  = ~\new_[8717]_  | ~n4110;
  assign \new_[7400]_  = ~\new_[7623]_  | ~\new_[1218]_ ;
  assign \new_[7401]_  = ~\new_[8039]_  | ~n4110;
  assign \new_[7402]_  = ~\new_[7990]_  | ~n4110;
  assign \new_[7403]_  = ~\new_[7623]_  | ~\new_[1099]_ ;
  assign \new_[7404]_  = ~\new_[7584]_  | ~\new_[1152]_ ;
  assign \new_[7405]_  = ~\new_[7623]_  | ~\new_[1214]_ ;
  assign \new_[7406]_  = ~first_round_reg_reg;
  assign \new_[7407]_  = ~\new_[7619]_  | ~\new_[6432]_ ;
  assign \new_[7408]_  = ~\new_[7619]_  | ~\new_[6623]_ ;
  assign \new_[7409]_  = ~\new_[7619]_  | ~\new_[3107]_ ;
  assign \new_[7410]_  = ~\new_[7573]_ ;
  assign \new_[7411]_  = ~\new_[7619]_  | ~\new_[3104]_ ;
  assign \new_[7412]_  = ~\new_[7600]_  | ~\new_[7658]_ ;
  assign \new_[7413]_  = ~\new_[7619]_  | ~\new_[6591]_ ;
  assign \new_[7414]_  = ~\new_[7619]_  | ~\new_[6624]_ ;
  assign \new_[7415]_  = ~\new_[7619]_  | ~\new_[2755]_ ;
  assign \new_[7416]_  = ~\new_[7619]_  | ~\new_[6585]_ ;
  assign \new_[7417]_  = ~\new_[7619]_  | ~\new_[6584]_ ;
  assign \new_[7418]_  = ~\new_[7619]_  | ~\new_[6422]_ ;
  assign \new_[7419]_  = ~\new_[7619]_  | ~\new_[3108]_ ;
  assign \new_[7420]_  = ~\new_[7619]_  | ~\new_[3846]_ ;
  assign \new_[7421]_  = ~\new_[7619]_  | ~\new_[6546]_ ;
  assign \new_[7422]_  = ~\new_[7619]_  | ~\new_[6579]_ ;
  assign \new_[7423]_  = ~\new_[7656]_  | ~\new_[7615]_ ;
  assign \new_[7424]_  = ~\new_[7619]_  | ~\new_[6594]_ ;
  assign \new_[7425]_  = ~\new_[7619]_  | ~\new_[6568]_ ;
  assign \new_[7426]_  = ~\new_[7619]_  | ~\new_[6640]_ ;
  assign \new_[7427]_  = \new_[7586]_  | \new_[7604]_ ;
  assign \new_[7428]_  = ~\new_[7901]_  & ~load_i & ~\new_[7884]_ ;
  assign \new_[7429]_  = ~\new_[7619]_  | ~\new_[3377]_ ;
  assign \new_[7430]_  = ~\new_[7619]_  | ~\new_[6694]_ ;
  assign \new_[7431]_  = ~\new_[7619]_  | ~\new_[6446]_ ;
  assign \new_[7432]_  = ~\new_[7619]_  | ~\new_[3387]_ ;
  assign \new_[7433]_  = ~\new_[7619]_  | ~\new_[6547]_ ;
  assign \new_[7434]_  = ~\new_[7619]_  | ~\new_[2870]_ ;
  assign \new_[7435]_  = ~\new_[7619]_  | ~\new_[6723]_ ;
  assign \new_[7436]_  = ~\new_[7619]_  | ~\new_[6631]_ ;
  assign \new_[7437]_  = ~\new_[7619]_  | ~\new_[3863]_ ;
  assign \new_[7438]_  = ~\new_[7619]_  | ~\new_[6751]_ ;
  assign \new_[7439]_  = ~\new_[7619]_  | ~\new_[6605]_ ;
  assign \new_[7440]_  = ~\new_[7619]_  | ~\new_[3409]_ ;
  assign \new_[7441]_  = ~\new_[7619]_  | ~\new_[6598]_ ;
  assign \new_[7442]_  = ~\new_[7619]_  | ~\new_[6423]_ ;
  assign n4105 = ~\new_[8343]_ ;
  assign \new_[7444]_  = ~\new_[7619]_  | ~\new_[6588]_ ;
  assign \new_[7445]_  = ~\new_[7619]_  | ~\new_[6421]_ ;
  assign \new_[7446]_  = ~\new_[7619]_  | ~\new_[6625]_ ;
  assign \new_[7447]_  = ~\new_[7619]_  | ~\new_[6495]_ ;
  assign \new_[7448]_  = ~\new_[7619]_  | ~\new_[6632]_ ;
  assign \new_[7449]_  = ~\new_[7619]_  | ~\new_[2934]_ ;
  assign \new_[7450]_  = ~\new_[7619]_  | ~\new_[6643]_ ;
  assign \new_[7451]_  = ~\new_[7619]_  | ~\new_[6716]_ ;
  assign \new_[7452]_  = ~\new_[7619]_  | ~\new_[3514]_ ;
  assign \new_[7453]_  = ~\new_[7619]_  | ~\new_[3383]_ ;
  assign \new_[7454]_  = ~\new_[7619]_  | ~\new_[6573]_ ;
  assign \new_[7455]_  = ~\new_[7619]_  | ~\new_[6619]_ ;
  assign \new_[7456]_  = ~\new_[7619]_  | ~\new_[6748]_ ;
  assign \new_[7457]_  = ~\new_[7619]_  | ~\new_[3385]_ ;
  assign \new_[7458]_  = ~\new_[7619]_  | ~\new_[3857]_ ;
  assign \new_[7459]_  = ~\new_[7619]_  | ~\new_[3257]_ ;
  assign \new_[7460]_  = ~\new_[7619]_  | ~\new_[3885]_ ;
  assign \new_[7461]_  = ~\new_[7619]_  | ~\new_[6749]_ ;
  assign \new_[7462]_  = ~\new_[7619]_  | ~\new_[6601]_ ;
  assign \new_[7463]_  = ~\new_[7619]_  | ~\new_[3382]_ ;
  assign \new_[7464]_  = ~\new_[7917]_  & ~load_i & ~\new_[7884]_ ;
  assign \new_[7465]_  = ~\new_[7619]_  | ~\new_[6627]_ ;
  assign \new_[7466]_  = ~\new_[7619]_  | ~\new_[6419]_ ;
  assign \new_[7467]_  = ~\new_[7593]_  & (~\new_[7751]_  | ~\new_[6041]_ );
  assign \new_[7468]_  = ~\new_[7619]_  | ~\new_[6427]_ ;
  assign \new_[7469]_  = ~\new_[7573]_ ;
  assign \new_[7470]_  = ~\new_[7573]_ ;
  assign \new_[7471]_  = ~\new_[7626]_  | ~\new_[7617]_ ;
  assign \new_[7472]_  = ~\new_[7593]_  & ~\new_[7934]_ ;
  assign \new_[7473]_  = ~\new_[7619]_  | ~\new_[2932]_ ;
  assign \new_[7474]_  = ~\new_[7619]_  | ~\new_[3105]_ ;
  assign \new_[7475]_  = ~\new_[7655]_  | ~\new_[7621]_ ;
  assign \new_[7476]_  = ~\new_[7619]_  | ~\new_[6652]_ ;
  assign \new_[7477]_  = ~\new_[7619]_  | ~\new_[6610]_ ;
  assign \new_[7478]_  = ~\new_[7619]_  | ~\new_[2757]_ ;
  assign \new_[7479]_  = ~\new_[7606]_ ;
  assign \new_[7480]_  = ~\new_[7564]_ ;
  assign \new_[7481]_  = ~\new_[7619]_  | ~\new_[6714]_ ;
  assign \new_[7482]_  = ~\new_[7619]_  | ~\new_[6618]_ ;
  assign \new_[7483]_  = ~\new_[7619]_  | ~\new_[6452]_ ;
  assign \new_[7484]_  = ~\new_[7619]_  | ~\new_[6451]_ ;
  assign \new_[7485]_  = ~\new_[7619]_  | ~\new_[3443]_ ;
  assign \new_[7486]_  = \new_[8343]_ ;
  assign \new_[7487]_  = ~\new_[7619]_  | ~\new_[6600]_ ;
  assign \new_[7488]_  = ~\new_[8881]_ ;
  assign \new_[7489]_  = ~\new_[7619]_  | ~\new_[6420]_ ;
  assign \new_[7490]_  = ~\new_[7619]_  | ~\new_[2758]_ ;
  assign \new_[7491]_  = ~\new_[7841]_  & ~\new_[7593]_ ;
  assign \new_[7492]_  = ~\new_[7619]_  | ~\new_[6416]_ ;
  assign \new_[7493]_  = ~\new_[7619]_  | ~\new_[6704]_ ;
  assign \new_[7494]_  = ~\new_[7606]_ ;
  assign \new_[7495]_  = ~\new_[7619]_  | ~\new_[6746]_ ;
  assign \new_[7496]_  = ~\new_[7566]_ ;
  assign \new_[7497]_  = ~\new_[7606]_ ;
  assign \new_[7498]_  = ~\new_[7606]_ ;
  assign \new_[7499]_  = \new_[7893]_  | \new_[8713]_ ;
  assign \new_[7500]_  = ~\new_[7619]_  | ~\new_[6702]_ ;
  assign \new_[7501]_  = ~\new_[7619]_  | ~\new_[3106]_ ;
  assign \new_[7502]_  = ~\new_[7619]_  | ~\new_[6656]_ ;
  assign \new_[7503]_  = ~\new_[7619]_  | ~\new_[6663]_ ;
  assign \new_[7504]_  = ~\new_[7619]_  | ~\new_[6620]_ ;
  assign \new_[7505]_  = ~\new_[7619]_  | ~\new_[6569]_ ;
  assign \new_[7506]_  = ~\new_[7619]_  | ~\new_[6430]_ ;
  assign \new_[7507]_  = ~\new_[7619]_  | ~\new_[6580]_ ;
  assign \new_[7508]_  = ~\new_[7619]_  | ~\new_[6449]_ ;
  assign \new_[7509]_  = ~\new_[7619]_  | ~\new_[3515]_ ;
  assign \new_[7510]_  = ~\new_[7619]_  | ~\new_[6445]_ ;
  assign \new_[7511]_  = ~\new_[7619]_  | ~\new_[3109]_ ;
  assign \new_[7512]_  = ~\new_[7619]_  | ~\new_[6433]_ ;
  assign \new_[7513]_  = ~\new_[7619]_  | ~\new_[6641]_ ;
  assign \new_[7514]_  = ~\new_[7619]_  | ~\new_[6596]_ ;
  assign \new_[7515]_  = ~\new_[7619]_  | ~\new_[6574]_ ;
  assign \new_[7516]_  = ~\new_[7619]_  | ~\new_[6429]_ ;
  assign \new_[7517]_  = ~\new_[7619]_  | ~\new_[6629]_ ;
  assign \new_[7518]_  = ~\new_[7619]_  | ~\new_[6444]_ ;
  assign \new_[7519]_  = ~\new_[7619]_  | ~\new_[6426]_ ;
  assign \new_[7520]_  = ~\new_[7619]_  | ~\new_[6614]_ ;
  assign \new_[7521]_  = ~\new_[7619]_  | ~\new_[6581]_ ;
  assign \new_[7522]_  = ~\new_[7619]_  | ~\new_[6438]_ ;
  assign \new_[7523]_  = ~\new_[7619]_  | ~\new_[6571]_ ;
  assign \new_[7524]_  = ~\new_[7619]_  | ~\new_[6587]_ ;
  assign \new_[7525]_  = ~\new_[7619]_  | ~\new_[6599]_ ;
  assign \new_[7526]_  = ~\new_[7619]_  | ~\new_[2756]_ ;
  assign \new_[7527]_  = ~\new_[7619]_  | ~\new_[6450]_ ;
  assign \new_[7528]_  = ~\new_[7619]_  | ~\new_[6586]_ ;
  assign \new_[7529]_  = ~\new_[7619]_  | ~\new_[6639]_ ;
  assign \new_[7530]_  = ~\new_[7619]_  | ~\new_[6630]_ ;
  assign \new_[7531]_  = ~\new_[7619]_  | ~\new_[6589]_ ;
  assign \new_[7532]_  = ~\new_[7619]_  | ~\new_[3406]_ ;
  assign \new_[7533]_  = ~\new_[7619]_  | ~\new_[6442]_ ;
  assign \new_[7534]_  = ~\new_[7619]_  | ~\new_[6425]_ ;
  assign \new_[7535]_  = ~\new_[7619]_  | ~\new_[6597]_ ;
  assign \new_[7536]_  = \\ks1_state_reg[1] ;
  assign \new_[7537]_  = ~\new_[7619]_  | ~\new_[6575]_ ;
  assign \new_[7538]_  = ~\new_[7619]_  | ~\new_[6593]_ ;
  assign \new_[7539]_  = ~\new_[7619]_  | ~\new_[6616]_ ;
  assign \new_[7540]_  = ~\new_[7619]_  | ~\new_[6606]_ ;
  assign \new_[7541]_  = ~\new_[7619]_  | ~\new_[6607]_ ;
  assign \new_[7542]_  = ~\new_[7619]_  | ~\new_[2935]_ ;
  assign \new_[7543]_  = ~\new_[7619]_  | ~\new_[3410]_ ;
  assign \new_[7544]_  = ~\new_[7619]_  | ~\new_[6626]_ ;
  assign \new_[7545]_  = ~\new_[7619]_  | ~\new_[6609]_ ;
  assign \new_[7546]_  = ~\new_[7619]_  | ~\new_[6590]_ ;
  assign \new_[7547]_  = ~\new_[7619]_  | ~\new_[6628]_ ;
  assign \new_[7548]_  = ~\new_[7619]_  | ~\new_[6443]_ ;
  assign \new_[7549]_  = ~\new_[7619]_  | ~\new_[6595]_ ;
  assign \new_[7550]_  = ~\new_[7619]_  | ~\new_[6592]_ ;
  assign \new_[7551]_  = ~\new_[7619]_  | ~\new_[6424]_ ;
  assign \new_[7552]_  = ~\new_[7619]_  | ~\new_[6572]_ ;
  assign \new_[7553]_  = ~\new_[7619]_  | ~\new_[6428]_ ;
  assign \new_[7554]_  = ~\new_[7619]_  | ~\new_[6566]_ ;
  assign \new_[7555]_  = ~\new_[7619]_  | ~\new_[6448]_ ;
  assign \new_[7556]_  = ~\new_[7619]_  | ~\new_[3386]_ ;
  assign \new_[7557]_  = ~\new_[7619]_  | ~\new_[3103]_ ;
  assign \new_[7558]_  = ~\new_[7619]_  | ~\new_[6666]_ ;
  assign \new_[7559]_  = ~\new_[7606]_ ;
  assign \new_[7560]_  = ~n4110;
  assign \new_[7561]_  = \new_[7958]_  ? \new_[7769]_  : \new_[7961]_ ;
  assign \new_[7562]_  = \key_i[21]  ? \new_[7769]_  : \new_[1981]_ ;
  assign \new_[7563]_  = \new_[8807]_  & decrypt_i;
  assign \new_[7564]_  = \new_[7606]_ ;
  assign \new_[7565]_  = ~\new_[5784]_  | ~\new_[7921]_ ;
  assign \new_[7566]_  = \new_[8948]_  | \new_[7905]_ ;
  assign n4115 = ~\new_[7585]_ ;
  assign \new_[7568]_  = ~\new_[7730]_  | ~\new_[7657]_ ;
  assign \new_[7569]_  = ~\new_[7738]_ ;
  assign \new_[7570]_  = ~\new_[7629]_  | ~\new_[7765]_ ;
  assign \new_[7571]_  = ~\new_[8730]_ ;
  assign \new_[7572]_  = ~sub1_ready_o_reg;
  assign \new_[7573]_  = ~\new_[8853]_ ;
  assign \new_[7574]_  = ~\new_[7729]_  | ~\new_[7628]_ ;
  assign \new_[7575]_  = ~\new_[7639]_  | ~\new_[7761]_ ;
  assign \new_[7576]_  = \new_[6041]_  ^ \new_[7752]_ ;
  assign \new_[7577]_  = ~\new_[7593]_ ;
  assign \new_[7578]_  = ~\new_[7636]_  | ~\new_[7682]_ ;
  assign \new_[7579]_  = ~\new_[7588]_ ;
  assign \new_[7580]_  = \new_[7927]_  ^ \new_[7690]_ ;
  assign \new_[7581]_  = ~\new_[7660]_ ;
  assign \new_[7582]_  = ~\new_[7660]_ ;
  assign \new_[7583]_  = ~\new_[7738]_ ;
  assign \new_[7584]_  = ~\new_[7648]_ ;
  assign \new_[7585]_  = ~load_i | ~\new_[5784]_ ;
  assign \new_[7586]_  = ~\new_[7646]_ ;
  assign \new_[7587]_  = \new_[7918]_  ^ \new_[7819]_ ;
  assign \new_[7588]_  = ~\new_[7767]_  | ~\new_[7676]_ ;
  assign \new_[7589]_  = ~\new_[7860]_  | ~\key_i[14] ;
  assign \new_[7590]_  = \new_[8098]_  ? \new_[7844]_  : \new_[8107]_ ;
  assign \new_[7591]_  = ~\new_[7874]_  | ~\key_i[22] ;
  assign \new_[7592]_  = ~\new_[7648]_ ;
  assign \new_[7593]_  = ~\new_[7751]_  & ~\new_[6041]_ ;
  assign \new_[7594]_  = \new_[8017]_  ? \new_[7845]_  : \new_[7994]_ ;
  assign \new_[7595]_  = ~\new_[7860]_  | ~\key_i[6] ;
  assign \new_[7596]_  = \new_[8084]_  ? \new_[7844]_  : \new_[8106]_ ;
  assign \new_[7597]_  = ~\new_[8343]_ ;
  assign \new_[7598]_  = ~\new_[7764]_  & (~\new_[7843]_  | ~\new_[4230]_ );
  assign \new_[7599]_  = ~\new_[7648]_ ;
  assign \new_[7600]_  = ~\new_[8949]_  | ~\new_[7905]_ ;
  assign n4110 = \new_[8784]_ ;
  assign \new_[7602]_  = ~\new_[7648]_ ;
  assign \new_[7603]_  = ~\new_[7648]_ ;
  assign \new_[7604]_  = ~\new_[7643]_ ;
  assign \new_[7605]_  = ~\new_[7833]_  & (~\new_[7880]_  | ~\new_[5960]_ );
  assign \new_[7606]_  = ~\new_[7646]_ ;
  assign \new_[7607]_  = ~\new_[7662]_ ;
  assign n4120 = \new_[7679]_  | \new_[7764]_ ;
  assign \new_[7609]_  = ~\new_[5784]_  | ~\new_[7926]_ ;
  assign \new_[7610]_  = ~\new_[7760]_  | ~\new_[7762]_ ;
  assign \new_[7611]_  = \new_[8153]_  ? \new_[7844]_  : \new_[7970]_ ;
  assign \new_[7612]_  = \new_[7999]_  ? \new_[7844]_  : \new_[8051]_ ;
  assign \new_[7613]_  = (~\new_[7844]_  & ~\new_[8123]_ ) | (~\new_[7873]_  & ~\new_[8047]_ );
  assign \new_[7614]_  = ~\new_[8422]_  & ~\new_[8853]_ ;
  assign \new_[7615]_  = ~\new_[7874]_  | ~\key_i[17] ;
  assign \new_[7616]_  = ~\new_[7874]_  | ~\key_i[20] ;
  assign \new_[7617]_  = ~\new_[7860]_  | ~\key_i[11] ;
  assign \new_[7618]_  = ~\new_[7860]_  | ~\key_i[16] ;
  assign \new_[7619]_  = ~\new_[7694]_  | ~\new_[7829]_ ;
  assign \new_[7620]_  = ~\new_[7660]_ ;
  assign \new_[7621]_  = ~\new_[7874]_  | ~\key_i[3] ;
  assign \new_[7622]_  = \new_[5960]_  ^ \new_[7891]_ ;
  assign \new_[7623]_  = ~\new_[7648]_ ;
  assign \new_[7624]_  = ~\new_[7662]_ ;
  assign \new_[7625]_  = ~\new_[7659]_ ;
  assign \new_[7626]_  = ~\new_[7844]_  | ~\new_[1061]_ ;
  assign \new_[7627]_  = ~\new_[9018]_  & (~\new_[7904]_  | ~\new_[7921]_ );
  assign \new_[7628]_  = ~\new_[7846]_  | ~\key_i[1] ;
  assign \new_[7629]_  = ~\new_[7845]_  | ~\new_[1966]_ ;
  assign n4125 = \new_[7842]_  & \new_[7872]_ ;
  assign \new_[7631]_  = ~\new_[7688]_ ;
  assign \new_[7632]_  = ~\new_[7738]_ ;
  assign \new_[7633]_  = ~\new_[7572]_  & ~\new_[1146]_ ;
  assign \new_[7634]_  = ~\new_[7844]_  | ~\new_[1978]_ ;
  assign \new_[7635]_  = ~\new_[8853]_  & ~\new_[7821]_ ;
  assign \new_[7636]_  = ~\new_[7850]_  | ~\new_[1980]_ ;
  assign \new_[7637]_  = ~\new_[7850]_  | ~\new_[1942]_ ;
  assign \new_[7638]_  = ~\new_[7572]_  & ~\new_[1540]_ ;
  assign \new_[7639]_  = ~\new_[7850]_  | ~\new_[1072]_ ;
  assign \new_[7640]_  = \new_[9018]_  | \new_[7901]_ ;
  assign \new_[7641]_  = \new_[8077]_  ? \new_[7855]_  : \new_[7937]_ ;
  assign \new_[7642]_  = \new_[7943]_  ? \new_[7855]_  : \new_[7953]_ ;
  assign \new_[7643]_  = ~\new_[7891]_  | ~\new_[7824]_ ;
  assign \new_[7644]_  = ~\new_[7572]_  & ~\new_[1558]_ ;
  assign \new_[7645]_  = ~\new_[7694]_ ;
  assign \new_[7646]_  = ~\new_[6041]_  | ~\new_[7891]_  | ~\new_[8049]_ ;
  assign \new_[7647]_  = ~\new_[7572]_  & ~\new_[1539]_ ;
  assign \new_[7648]_  = ~\new_[8052]_  | ~decrypt_i;
  assign \new_[7649]_  = (~\new_[7875]_  & ~\new_[8135]_ ) | (~\new_[7860]_  & ~\new_[7979]_ );
  assign \new_[7650]_  = \new_[8022]_  ? \new_[7875]_  : \new_[8148]_ ;
  assign \new_[7651]_  = (~\new_[7897]_  & ~\new_[8131]_ ) | (~\new_[7874]_  & ~\new_[7951]_ );
  assign \new_[7652]_  = \new_[7962]_  ? \new_[7855]_  : \new_[7952]_ ;
  assign \new_[7653]_  = ~\new_[7844]_  | ~\new_[1963]_ ;
  assign \new_[7654]_  = ~\new_[7844]_  | ~\new_[1064]_ ;
  assign \new_[7655]_  = ~\new_[7844]_  | ~\new_[1960]_ ;
  assign \new_[7656]_  = ~\new_[7844]_  | ~\new_[1977]_ ;
  assign \new_[7657]_  = ~\new_[7846]_  | ~\key_i[2] ;
  assign \new_[7658]_  = ~\new_[8698]_  | ~\new_[7889]_ ;
  assign \new_[7659]_  = ~\new_[8698]_  & ~\new_[8799]_ ;
  assign \new_[7660]_  = ~\new_[7769]_ ;
  assign \new_[7661]_  = \new_[8097]_  ? \new_[7855]_  : \new_[8006]_ ;
  assign \new_[7662]_  = ~\new_[7770]_ ;
  assign \new_[7663]_  = ~\new_[7572]_  & ~\new_[1462]_ ;
  assign \new_[7664]_  = \new_[8799]_  | \new_[7839]_ ;
  assign \new_[7665]_  = ~\new_[7572]_  & ~\new_[1541]_ ;
  assign \new_[7666]_  = \new_[7900]_  & \new_[1249]_ ;
  assign \new_[7667]_  = \new_[7906]_  & \new_[1190]_ ;
  assign \new_[7668]_  = \new_[7871]_  & \new_[8195]_ ;
  assign \new_[7669]_  = \new_[7900]_  & \new_[1210]_ ;
  assign \new_[7670]_  = \new_[7900]_  & \new_[1191]_ ;
  assign \new_[7671]_  = \new_[7900]_  & \new_[1224]_ ;
  assign \new_[7672]_  = \new_[7906]_  & \new_[1219]_ ;
  assign \new_[7673]_  = \new_[7900]_  & \new_[1192]_ ;
  assign \new_[7674]_  = \new_[7906]_  & \new_[1109]_ ;
  assign \new_[7675]_  = \new_[7921]_  ^ \new_[7887]_ ;
  assign \new_[7676]_  = ~\new_[8664]_  | ~\new_[8799]_ ;
  assign \new_[7677]_  = \new_[7906]_  & \new_[1200]_ ;
  assign \new_[7678]_  = \new_[7906]_  & \new_[1240]_ ;
  assign \new_[7679]_  = \new_[7879]_  & \new_[7881]_ ;
  assign \new_[7680]_  = \new_[7906]_  & \new_[1148]_ ;
  assign \new_[7681]_  = ~\new_[7873]_  | ~\key_i[28] ;
  assign \new_[7682]_  = ~\new_[7873]_  | ~\key_i[18] ;
  assign \new_[7683]_  = ~decrypt_i | ~\new_[8238]_  | ~\new_[2426]_ ;
  assign \new_[7684]_  = \new_[7900]_  & \new_[1099]_ ;
  assign \new_[7685]_  = \new_[7900]_  & \new_[1247]_ ;
  assign \new_[7686]_  = \new_[7900]_  & \new_[1459]_ ;
  assign \new_[7687]_  = \new_[7900]_  & \new_[1105]_ ;
  assign \new_[7688]_  = ~\new_[8329]_ ;
  assign \new_[7689]_  = \new_[7900]_  & \new_[1248]_ ;
  assign \new_[7690]_  = ~\new_[7857]_  | ~\new_[7921]_ ;
  assign \new_[7691]_  = \new_[7906]_  & \new_[1461]_ ;
  assign \new_[7692]_  = \new_[7900]_  & \new_[1095]_ ;
  assign \new_[7693]_  = \new_[7906]_  & \new_[1221]_ ;
  assign \new_[7694]_  = ~\new_[8558]_  & ~\new_[8713]_ ;
  assign \new_[7695]_  = \new_[7900]_  & \new_[1134]_ ;
  assign \new_[7696]_  = \new_[7906]_  & \new_[1216]_ ;
  assign \new_[7697]_  = \new_[7906]_  & \new_[1319]_ ;
  assign \new_[7698]_  = \new_[7906]_  & \new_[1324]_ ;
  assign \new_[7699]_  = \new_[7900]_  & \new_[1195]_ ;
  assign \new_[7700]_  = \new_[7900]_  & \new_[1137]_ ;
  assign \new_[7701]_  = \new_[7906]_  & \new_[1114]_ ;
  assign \new_[7702]_  = \new_[7906]_  & \new_[1530]_ ;
  assign \new_[7703]_  = \new_[7906]_  & \new_[1207]_ ;
  assign \new_[7704]_  = \new_[7900]_  & \new_[1101]_ ;
  assign \new_[7705]_  = \new_[7906]_  & \new_[1106]_ ;
  assign \new_[7706]_  = \new_[7900]_  & \new_[1206]_ ;
  assign \new_[7707]_  = \new_[7900]_  & \new_[1246]_ ;
  assign \new_[7708]_  = \new_[7906]_  & \new_[1204]_ ;
  assign \new_[7709]_  = \new_[7906]_  & \new_[1214]_ ;
  assign \new_[7710]_  = \new_[7906]_  & \new_[1110]_ ;
  assign \new_[7711]_  = \new_[7906]_  & \new_[1220]_ ;
  assign \new_[7712]_  = \new_[7900]_  & \new_[1201]_ ;
  assign \new_[7713]_  = \new_[7900]_  & \new_[1323]_ ;
  assign \new_[7714]_  = \new_[7906]_  & \new_[1136]_ ;
  assign \new_[7715]_  = \new_[7906]_  & \new_[1199]_ ;
  assign \new_[7716]_  = \new_[7906]_  & \new_[1520]_ ;
  assign \new_[7717]_  = \new_[7900]_  & \new_[1385]_ ;
  assign \new_[7718]_  = \new_[7906]_  & \new_[1203]_ ;
  assign \new_[7719]_  = \new_[7906]_  & \new_[1381]_ ;
  assign \new_[7720]_  = \new_[7906]_  & \new_[1151]_ ;
  assign \new_[7721]_  = \new_[7906]_  & \new_[1147]_ ;
  assign \new_[7722]_  = \new_[7906]_  & \new_[1321]_ ;
  assign \new_[7723]_  = \new_[7900]_  & \new_[1314]_ ;
  assign \new_[7724]_  = \new_[7900]_  & \new_[1244]_ ;
  assign \new_[7725]_  = \new_[7900]_  & \new_[1226]_ ;
  assign \new_[7726]_  = \new_[7900]_  & \new_[1313]_ ;
  assign \new_[7727]_  = ~\new_[7875]_  | ~\new_[1982]_ ;
  assign \new_[7728]_  = \new_[7900]_  & \new_[1211]_ ;
  assign \new_[7729]_  = ~\new_[7855]_  | ~\new_[1965]_ ;
  assign \new_[7730]_  = ~\new_[7875]_  | ~\new_[1959]_ ;
  assign \new_[7731]_  = \new_[7900]_  & \new_[1097]_ ;
  assign \new_[7732]_  = \new_[7900]_  & \new_[1193]_ ;
  assign \new_[7733]_  = \new_[7900]_  & \new_[1138]_ ;
  assign \new_[7734]_  = \new_[7900]_  & \new_[1250]_ ;
  assign \new_[7735]_  = \new_[7906]_  & \new_[1205]_ ;
  assign \new_[7736]_  = \new_[7900]_  & \new_[1187]_ ;
  assign \new_[7737]_  = \new_[7900]_  & \new_[1135]_ ;
  assign \new_[7738]_  = ~decrypt_i;
  assign \new_[7739]_  = \new_[7906]_  & \new_[1242]_ ;
  assign \new_[7740]_  = \new_[7906]_  & \new_[1222]_ ;
  assign \new_[7741]_  = \new_[7906]_  & \new_[1208]_ ;
  assign \new_[7742]_  = \new_[7906]_  & \new_[1108]_ ;
  assign \new_[7743]_  = \new_[7906]_  & \new_[1521]_ ;
  assign \new_[7744]_  = \new_[7906]_  & \new_[1117]_ ;
  assign \new_[7745]_  = \new_[7900]_  & \new_[1098]_ ;
  assign \new_[7746]_  = \new_[7900]_  & \new_[1312]_ ;
  assign \new_[7747]_  = ~\new_[8663]_ ;
  assign \new_[7748]_  = \new_[7906]_  & \new_[1322]_ ;
  assign \new_[7749]_  = \new_[7900]_  & \new_[1241]_ ;
  assign \new_[7750]_  = \new_[7900]_  & \new_[1243]_ ;
  assign \new_[7751]_  = ~\new_[7836]_ ;
  assign \new_[7752]_  = ~\new_[7838]_ ;
  assign \new_[7753]_  = \new_[7900]_  & \new_[1139]_ ;
  assign \new_[7754]_  = \new_[7900]_  & \new_[1238]_ ;
  assign \new_[7755]_  = \new_[7900]_  & \new_[1152]_ ;
  assign \new_[7756]_  = \new_[7906]_  & \new_[1094]_ ;
  assign \new_[7757]_  = \new_[7906]_  & \new_[1212]_ ;
  assign \new_[7758]_  = \new_[7900]_  & \new_[1100]_ ;
  assign \new_[7759]_  = \new_[7900]_  & \new_[1386]_ ;
  assign \new_[7760]_  = ~\new_[7855]_  | ~\new_[1062]_ ;
  assign \new_[7761]_  = ~\new_[7873]_  | ~\key_i[10] ;
  assign \new_[7762]_  = ~\new_[7873]_  | ~\key_i[12] ;
  assign \new_[7763]_  = \new_[7906]_  & \new_[1150]_ ;
  assign \new_[7764]_  = \new_[7881]_  & \new_[7925]_ ;
  assign \new_[7765]_  = ~\new_[7873]_  | ~\key_i[23] ;
  assign \new_[7766]_  = \new_[7900]_  & \new_[1144]_ ;
  assign \new_[7767]_  = \new_[8664]_  | \new_[8799]_ ;
  assign \new_[7768]_  = ~\new_[7875]_  | ~\new_[1993]_ ;
  assign \new_[7769]_  = ~\new_[7846]_ ;
  assign \new_[7770]_  = ~\new_[6952]_  | ~\new_[8237]_ ;
  assign \new_[7771]_  = \new_[7906]_  & \new_[1103]_ ;
  assign \new_[7772]_  = \new_[7900]_  & \new_[1113]_ ;
  assign \new_[7773]_  = \new_[7900]_  & \new_[1143]_ ;
  assign \new_[7774]_  = \new_[7906]_  & \new_[1194]_ ;
  assign \new_[7775]_  = \new_[7900]_  & \new_[1457]_ ;
  assign \new_[7776]_  = \new_[7900]_  & \new_[1251]_ ;
  assign \new_[7777]_  = \new_[7900]_  & \new_[1196]_ ;
  assign \new_[7778]_  = \new_[7900]_  & \new_[1145]_ ;
  assign \new_[7779]_  = \new_[7906]_  & \new_[1213]_ ;
  assign \new_[7780]_  = \new_[7906]_  & \new_[1111]_ ;
  assign \new_[7781]_  = \new_[7906]_  & \new_[1463]_ ;
  assign \new_[7782]_  = \new_[7900]_  & \new_[1197]_ ;
  assign \new_[7783]_  = \new_[7900]_  & \new_[1384]_ ;
  assign \new_[7784]_  = \new_[7906]_  & \new_[1215]_ ;
  assign \new_[7785]_  = \new_[7906]_  & \new_[1202]_ ;
  assign \new_[7786]_  = \new_[7900]_  & \new_[1225]_ ;
  assign \new_[7787]_  = \new_[7900]_  & \new_[1096]_ ;
  assign \new_[7788]_  = \new_[7906]_  & \new_[1237]_ ;
  assign \new_[7789]_  = \new_[7900]_  & \new_[1320]_ ;
  assign \new_[7790]_  = \new_[7906]_  & \new_[1234]_ ;
  assign \new_[7791]_  = \new_[7906]_  & \new_[1116]_ ;
  assign \new_[7792]_  = \new_[7906]_  & \new_[1104]_ ;
  assign \new_[7793]_  = \new_[7906]_  & \new_[1186]_ ;
  assign \new_[7794]_  = \new_[7900]_  & \new_[1245]_ ;
  assign \new_[7795]_  = \new_[7900]_  & \new_[1252]_ ;
  assign \new_[7796]_  = \new_[7900]_  & \new_[1223]_ ;
  assign \new_[7797]_  = \new_[7906]_  & \new_[1102]_ ;
  assign \new_[7798]_  = \new_[7906]_  & \new_[1149]_ ;
  assign \new_[7799]_  = \new_[7900]_  & \new_[1209]_ ;
  assign \new_[7800]_  = \new_[7906]_  & \new_[1464]_ ;
  assign \new_[7801]_  = \new_[7900]_  & \new_[1198]_ ;
  assign \new_[7802]_  = \new_[7906]_  & \new_[1538]_ ;
  assign \new_[7803]_  = \new_[7900]_  & \new_[1383]_ ;
  assign \new_[7804]_  = \new_[7906]_  & \new_[1115]_ ;
  assign \new_[7805]_  = \new_[7906]_  & \new_[1315]_ ;
  assign \new_[7806]_  = \new_[7900]_  & \new_[1458]_ ;
  assign \new_[7807]_  = \new_[7906]_  & \new_[1107]_ ;
  assign \new_[7808]_  = \new_[7906]_  & \new_[1311]_ ;
  assign \new_[7809]_  = \new_[7906]_  & \new_[1460]_ ;
  assign \new_[7810]_  = \new_[7900]_  & \new_[1142]_ ;
  assign \new_[7811]_  = \new_[7900]_  & \new_[1112]_ ;
  assign \new_[7812]_  = \new_[7900]_  & \new_[1217]_ ;
  assign \new_[7813]_  = \new_[7906]_  & \new_[1218]_ ;
  assign \new_[7814]_  = ~\new_[7858]_ ;
  assign \new_[7815]_  = ~\new_[7883]_  & ~\new_[7907]_ ;
  assign \new_[7816]_  = ~\new_[8802]_ ;
  assign \new_[7817]_  = ~\new_[7891]_  | ~\new_[5960]_ ;
  assign \new_[7818]_  = ~\new_[7895]_  & ~\new_[7898]_ ;
  assign \new_[7819]_  = \new_[7892]_  | \new_[7982]_ ;
  assign \new_[7820]_  = ~\new_[7883]_  & ~\new_[7919]_ ;
  assign \new_[7821]_  = ~\new_[7862]_ ;
  assign \new_[7822]_  = ~\new_[8562]_ ;
  assign \new_[7823]_  = \new_[7877]_  | \new_[8160]_ ;
  assign \new_[7824]_  = ~\new_[5960]_  & ~\new_[6041]_ ;
  assign \new_[7825]_  = ~\new_[8714]_ ;
  assign \new_[7826]_  = ~\new_[8422]_ ;
  assign \new_[7827]_  = \new_[7895]_  | \new_[7907]_ ;
  assign \new_[7828]_  = ~\new_[8185]_ ;
  assign \new_[7829]_  = ~\new_[7893]_ ;
  assign \new_[7830]_  = \new_[5990]_  ^ \new_[7913]_ ;
  assign \new_[7831]_  = ~\new_[7895]_  & ~\new_[7913]_ ;
  assign \new_[7832]_  = ~\new_[7883]_  & ~\new_[7898]_ ;
  assign \new_[7833]_  = ~\new_[7880]_  & ~\new_[5960]_ ;
  assign \new_[7834]_  = ~\new_[7863]_ ;
  assign \new_[7835]_  = ~\new_[7892]_  | ~\new_[7982]_ ;
  assign \new_[7836]_  = ~\new_[7895]_  & ~\new_[7919]_ ;
  assign \new_[7837]_  = ~\new_[7853]_ ;
  assign \new_[7838]_  = ~\new_[7880]_  & ~\new_[8049]_ ;
  assign \new_[7839]_  = ~\new_[8664]_ ;
  assign \new_[7840]_  = ~\new_[7887]_  | ~\new_[7904]_ ;
  assign \new_[7841]_  = ~\new_[7891]_  & (~\new_[7919]_  | ~\new_[5990]_ );
  assign \new_[7842]_  = ~\new_[7895]_  & ~\new_[7934]_ ;
  assign \new_[7843]_  = ~\new_[7881]_ ;
  assign \new_[7844]_  = ~\new_[7873]_ ;
  assign \new_[7845]_  = ~\new_[7860]_ ;
  assign \new_[7846]_  = ~\new_[7875]_ ;
  assign \new_[7847]_  = ~\new_[7886]_  & (~\new_[7924]_  | ~\new_[1592]_ );
  assign \new_[7848]_  = \new_[7917]_  ^ \new_[8125]_ ;
  assign \new_[7849]_  = ~\new_[7572]_  & ~decrypt_i;
  assign \new_[7850]_  = ~\new_[7874]_ ;
  assign \new_[7851]_  = \new_[8137]_  ? \new_[8237]_  : \new_[7932]_ ;
  assign \new_[7852]_  = ~\new_[7909]_  & ~\new_[7898]_ ;
  assign \new_[7853]_  = \new_[7919]_  & \new_[7913]_ ;
  assign \new_[7854]_  = ~\new_[7909]_  & ~\new_[7907]_ ;
  assign \new_[7855]_  = \new_[7897]_ ;
  assign \new_[7856]_  = ~\new_[7908]_  | ~\new_[7911]_ ;
  assign \new_[7857]_  = ~\new_[7887]_ ;
  assign \new_[7858]_  = \new_[7905]_  | \new_[8799]_ ;
  assign \new_[7859]_  = ~\new_[8113]_  | ~\new_[7975]_ ;
  assign \new_[7860]_  = ~\new_[7897]_ ;
  assign \new_[7861]_  = ~\new_[7915]_  & ~\new_[7898]_ ;
  assign \new_[7862]_  = ~\new_[8378]_ ;
  assign \new_[7863]_  = \new_[8689]_  | \new_[8799]_ ;
  assign \new_[7864]_  = ~\new_[7909]_  & ~\new_[7919]_ ;
  assign \new_[7865]_  = ~\new_[7915]_  & ~\new_[7913]_ ;
  assign \new_[7866]_  = ~\new_[7915]_  & ~\new_[7907]_ ;
  assign \new_[7867]_  = \new_[7898]_  & \new_[7907]_ ;
  assign \new_[7868]_  = ~\new_[7912]_  & (~\new_[8113]_  | ~\new_[8195]_ );
  assign \new_[7869]_  = \new_[7914]_  & \new_[7929]_ ;
  assign \new_[7870]_  = \new_[1387]_  ^ \new_[7922]_ ;
  assign \new_[7871]_  = ~\new_[7901]_  & ~decrypt_i;
  assign \new_[7872]_  = ~\new_[5991]_  & ~\new_[7987]_ ;
  assign \new_[7873]_  = ~\new_[7897]_ ;
  assign \new_[7874]_  = ~\new_[7897]_ ;
  assign \new_[7875]_  = \new_[7897]_ ;
  assign \new_[7876]_  = ~\new_[7910]_  & (~\new_[7975]_  | ~\new_[7963]_ );
  assign \new_[7877]_  = ~\new_[7536]_  & ~\new_[4230]_ ;
  assign \new_[7878]_  = ~\new_[5784]_ ;
  assign \new_[7879]_  = ~\new_[7536]_  & ~\new_[4362]_ ;
  assign \new_[7880]_  = ~\new_[7935]_  | ~\new_[5990]_ ;
  assign \new_[7881]_  = ~\new_[7925]_  | ~\new_[8060]_ ;
  assign \new_[7882]_  = ~\new_[5784]_ ;
  assign \new_[7883]_  = ~\new_[5990]_  | ~\new_[5960]_ ;
  assign \new_[7884]_  = ~\new_[5784]_ ;
  assign \new_[7885]_  = ~\new_[5784]_ ;
  assign \new_[7886]_  = ~\new_[7924]_  & ~\new_[1592]_ ;
  assign \new_[7887]_  = ~\new_[7926]_  | ~\new_[7930]_ ;
  assign \new_[7888]_  = ~\new_[5784]_ ;
  assign \new_[7889]_  = ~\new_[7905]_ ;
  assign \new_[7890]_  = ~\new_[7904]_ ;
  assign \new_[7891]_  = ~\new_[7919]_  & ~\new_[5990]_ ;
  assign \new_[7892]_  = ~\new_[7928]_  | ~\new_[7923]_ ;
  assign \new_[7893]_  = ~\new_[7902]_ ;
  assign \new_[7894]_  = \new_[7926]_  & \new_[8046]_ ;
  assign \new_[7895]_  = \new_[5990]_  | \new_[5960]_ ;
  assign \new_[7896]_  = ~\new_[7920]_  & (~\new_[7982]_  | ~\new_[8046]_ );
  assign \new_[7897]_  = \new_[7933]_  | \new_[3981]_ ;
  assign \new_[7898]_  = \new_[5898]_  | \new_[7965]_ ;
  assign \new_[7899]_  = \new_[4230]_  & \new_[8160]_ ;
  assign \new_[7900]_  = ~\new_[7572]_ ;
  assign \new_[7901]_  = ~\new_[7927]_ ;
  assign \new_[7902]_  = ~\new_[8108]_  | ~\new_[5659]_ ;
  assign \new_[7903]_  = ~\new_[7927]_ ;
  assign \new_[7904]_  = ~\new_[7963]_  | ~\new_[8195]_ ;
  assign \new_[7905]_  = ~\new_[1068]_ ;
  assign \new_[7906]_  = ~\new_[7572]_ ;
  assign \new_[7907]_  = ~\new_[5898]_  | ~\new_[7965]_ ;
  assign \new_[7908]_  = \new_[8086]_  | \new_[1467]_ ;
  assign \new_[7909]_  = ~\new_[5990]_  | ~\new_[8049]_ ;
  assign \new_[7910]_  = ~\new_[7975]_  & ~\new_[8125]_ ;
  assign \new_[7911]_  = ~\new_[8086]_  | ~\new_[1467]_ ;
  assign \new_[7912]_  = ~\new_[8113]_  & ~\new_[8195]_ ;
  assign \new_[7913]_  = ~\new_[7935]_ ;
  assign \new_[7914]_  = \new_[8014]_  | \new_[8196]_ ;
  assign \new_[7915]_  = \new_[5990]_  | \new_[8049]_ ;
  assign \new_[7916]_  = ~\new_[7982]_ ;
  assign \new_[7917]_  = ~\new_[7930]_ ;
  assign \new_[7918]_  = ~\new_[8014]_ ;
  assign \new_[7919]_  = \new_[5898]_  | \new_[5991]_ ;
  assign \new_[7920]_  = \new_[3996]_  & \new_[5307]_ ;
  assign \new_[7921]_  = ~\new_[8046]_ ;
  assign \new_[7922]_  = ~\new_[8086]_ ;
  assign \new_[7923]_  = ~\new_[7975]_ ;
  assign \new_[7924]_  = ~\new_[8157]_ ;
  assign \new_[7925]_  = ~\new_[4230]_  & ~\new_[4362]_ ;
  assign \new_[7926]_  = ~\new_[8125]_ ;
  assign \new_[7927]_  = ~\new_[8196]_ ;
  assign \new_[7928]_  = ~\new_[8113]_ ;
  assign \new_[7929]_  = \new_[3982]_  | \new_[5419]_ ;
  assign \new_[7930]_  = ~\new_[8195]_ ;
  assign \new_[7931]_  = ~\new_[8699]_ ;
  assign \new_[7932]_  = ~\new_[2426]_ ;
  assign \new_[7933]_  = \new_[3996]_  | \new_[3982]_ ;
  assign \new_[7934]_  = ~\new_[7944]_ ;
  assign \new_[7935]_  = \new_[5898]_  & \new_[5991]_ ;
  assign \new_[7936]_  = ~\new_[1977]_ ;
  assign \new_[7937]_  = ~\new_[1969]_ ;
  assign \new_[7938]_  = ~\new_[2771]_ ;
  assign \new_[7939]_  = ~\new_[1540]_ ;
  assign \new_[7940]_  = ~\new_[2772]_ ;
  assign \new_[7941]_  = ~\new_[2006]_ ;
  assign \new_[7942]_  = ~\new_[2867]_ ;
  assign \new_[7943]_  = ~\key_i[31] ;
  assign \new_[7944]_  = ~\new_[5898]_ ;
  assign \new_[7945]_  = ~\new_[2417]_ ;
  assign \new_[7946]_  = ~\new_[1965]_ ;
  assign \new_[7947]_  = ~\new_[1189]_ ;
  assign \new_[7948]_  = ~\new_[2653]_ ;
  assign \new_[7949]_  = ~\new_[1308]_ ;
  assign \new_[7950]_  = ~\new_[1982]_ ;
  assign \new_[7951]_  = ~\new_[1950]_ ;
  assign \new_[7952]_  = ~\new_[1955]_ ;
  assign \new_[7953]_  = ~\new_[1951]_ ;
  assign \new_[7954]_  = ~\new_[1343]_ ;
  assign \new_[7955]_  = ~\new_[1188]_ ;
  assign \new_[7956]_  = ~\new_[3376]_ ;
  assign \new_[7957]_  = ~\new_[1976]_ ;
  assign \new_[7958]_  = ~\key_i[8] ;
  assign \new_[7959]_  = ~\new_[1379]_ ;
  assign \new_[7960]_  = ~\new_[2224]_ ;
  assign \new_[7961]_  = ~\new_[1070]_ ;
  assign \new_[7962]_  = ~\key_i[26] ;
  assign \new_[7963]_  = ~\new_[5377]_ ;
  assign \new_[7964]_  = ~\key_i[23] ;
  assign \new_[7965]_  = ~\new_[5991]_ ;
  assign \new_[7966]_  = ~\new_[2630]_ ;
  assign \new_[7967]_  = ~\key_i[28] ;
  assign \new_[7968]_  = ~\new_[2027]_ ;
  assign \new_[7969]_  = ~\new_[2873]_ ;
  assign \new_[7970]_  = ~\new_[1947]_ ;
  assign \new_[7971]_  = ~\new_[1305]_ ;
  assign \new_[7972]_  = ~\new_[2549]_ ;
  assign \new_[7973]_  = ~\new_[2026]_ ;
  assign \new_[7974]_  = ~\new_[2872]_ ;
  assign \new_[7975]_  = ~\new_[2267]_ ;
  assign \new_[7976]_  = ~\new_[2540]_ ;
  assign \new_[7977]_  = ~\new_[2420]_ ;
  assign \new_[7978]_  = ~\new_[2577]_ ;
  assign \new_[7979]_  = ~\new_[1964]_ ;
  assign \new_[7980]_  = ~\new_[2028]_ ;
  assign \new_[7981]_  = ~\new_[2415]_ ;
  assign \new_[7982]_  = ~\new_[3996]_ ;
  assign \new_[7983]_  = ~\new_[2998]_ ;
  assign \new_[7984]_  = ~\new_[1378]_ ;
  assign \new_[7985]_  = ~\new_[2868]_ ;
  assign \new_[7986]_  = ~\new_[1465]_ ;
  assign \new_[7987]_  = ~\new_[6041]_ ;
  assign \new_[7988]_  = ~\new_[2659]_ ;
  assign \new_[7989]_  = ~\key_i[5] ;
  assign \new_[7990]_  = ~\new_[2542]_ ;
  assign \new_[7991]_  = ~\new_[2029]_ ;
  assign \new_[7992]_  = ~\new_[2926]_ ;
  assign \new_[7993]_  = ~\new_[2052]_ ;
  assign \new_[7994]_  = ~\new_[1065]_ ;
  assign \new_[7995]_  = ~\new_[1064]_ ;
  assign \new_[7996]_  = ~\new_[1963]_ ;
  assign \new_[7997]_  = ~\new_[1309]_ ;
  assign \new_[7998]_  = ~\new_[2774]_ ;
  assign \new_[7999]_  = ~\key_i[25] ;
  assign \new_[8000]_  = ~\new_[2009]_ ;
  assign \new_[8001]_  = ~\new_[1975]_ ;
  assign \new_[8002]_  = ~\new_[2618]_ ;
  assign \new_[8003]_  = ~\new_[2346]_ ;
  assign \new_[8004]_  = ~\new_[1306]_ ;
  assign \new_[8005]_  = ~\new_[2007]_ ;
  assign \new_[8006]_  = ~\new_[1961]_ ;
  assign \new_[8007]_  = ~\new_[2763]_ ;
  assign \new_[8008]_  = ~\new_[2051]_ ;
  assign \new_[8009]_  = ~\new_[2033]_ ;
  assign \new_[8010]_  = ~\new_[2548]_ ;
  assign \new_[8011]_  = ~\new_[2046]_ ;
  assign \new_[8012]_  = ~\new_[1317]_ ;
  assign \new_[8013]_  = ~\new_[1979]_ ;
  assign \new_[8014]_  = ~\new_[3982]_ ;
  assign \new_[8015]_  = ~\new_[2628]_ ;
  assign \new_[8016]_  = ~\new_[2761]_ ;
  assign \new_[8017]_  = ~\key_i[15] ;
  assign \new_[8018]_  = ~\new_[1962]_ ;
  assign \new_[8019]_  = ~\new_[2539]_ ;
  assign \new_[8020]_  = ~\new_[1539]_ ;
  assign \new_[8021]_  = ~\new_[2550]_ ;
  assign \new_[8022]_  = ~\key_i[9] ;
  assign \new_[8023]_  = ~\new_[1542]_ ;
  assign \new_[8024]_  = ~\new_[1715]_ ;
  assign \new_[8025]_  = ~\new_[2869]_ ;
  assign \new_[8026]_  = ~\new_[1146]_ ;
  assign \new_[8027]_  = ~\new_[1233]_ ;
  assign \new_[8028]_  = ~\new_[1958]_ ;
  assign \new_[8029]_  = ~\new_[1596]_ ;
  assign \new_[8030]_  = ~\new_[2881]_ ;
  assign \new_[8031]_  = ~\new_[1980]_ ;
  assign \new_[8032]_  = ~\new_[2416]_ ;
  assign \new_[8033]_  = ~\new_[2545]_ ;
  assign \new_[8034]_  = ~\new_[1072]_ ;
  assign \new_[8035]_  = ~\new_[2866]_ ;
  assign \new_[8036]_  = ~\new_[2627]_ ;
  assign \new_[8037]_  = ~\new_[2066]_ ;
  assign \new_[8038]_  = ~\new_[1307]_ ;
  assign \new_[8039]_  = ~\new_[2546]_ ;
  assign \new_[8040]_  = ~\new_[2626]_ ;
  assign \new_[8041]_  = ~\new_[1316]_ ;
  assign \new_[8042]_  = ~\new_[2876]_ ;
  assign \new_[8043]_  = ~\new_[2883]_ ;
  assign \new_[8044]_  = ~\new_[2764]_ ;
  assign \new_[8045]_  = ~\new_[1382]_ ;
  assign \new_[8046]_  = ~\new_[5307]_ ;
  assign \new_[8047]_  = ~\new_[1063]_ ;
  assign \new_[8048]_  = ~\new_[2768]_ ;
  assign \new_[8049]_  = ~\new_[5960]_ ;
  assign \new_[8050]_  = ~\new_[1380]_ ;
  assign \new_[8051]_  = ~\new_[1952]_ ;
  assign \new_[8052]_  = ~\new_[7572]_ ;
  assign \new_[8053]_  = ~\new_[1541]_ ;
  assign \new_[8054]_  = ~\new_[2882]_ ;
  assign \new_[8055]_  = ~\new_[2005]_ ;
  assign \new_[8056]_  = ~\new_[1253]_ ;
  assign \new_[8057]_  = ~\new_[2047]_ ;
  assign \new_[8058]_  = ~\new_[1966]_ ;
  assign \new_[8059]_  = ~\new_[3389]_ ;
  assign \new_[8060]_  = ~\new_[7536]_ ;
  assign \new_[8061]_  = ~\new_[2874]_ ;
  assign \new_[8062]_  = ~\new_[2767]_ ;
  assign \new_[8063]_  = ~\new_[2538]_ ;
  assign \new_[8064]_  = ~\new_[2030]_ ;
  assign \new_[8065]_  = ~\new_[2419]_ ;
  assign \new_[8066]_  = ~\new_[2660]_ ;
  assign \new_[8067]_  = ~\new_[2769]_ ;
  assign \new_[8068]_  = ~\new_[1462]_ ;
  assign \new_[8069]_  = ~\new_[3000]_ ;
  assign \new_[8070]_  = ~\new_[2347]_ ;
  assign \new_[8071]_  = ~\new_[1978]_ ;
  assign \new_[8072]_  = ~\new_[1960]_ ;
  assign \new_[8073]_  = ~\new_[2999]_ ;
  assign \new_[8074]_  = ~\new_[2541]_ ;
  assign \new_[8075]_  = ~\new_[1590]_ ;
  assign \new_[8076]_  = ~\new_[2418]_ ;
  assign \new_[8077]_  = ~\key_i[7] ;
  assign \new_[8078]_  = ~\new_[1062]_ ;
  assign \new_[8079]_  = ~\new_[1318]_ ;
  assign \new_[8080]_  = ~\new_[3384]_ ;
  assign \new_[8081]_  = ~\new_[2775]_ ;
  assign \new_[8082]_  = ~\new_[2879]_ ;
  assign \new_[8083]_  = ~\new_[1466]_ ;
  assign \new_[8084]_  = ~\key_i[30] ;
  assign \new_[8085]_  = ~\new_[2658]_ ;
  assign \new_[8086]_  = ~\new_[1866]_ ;
  assign \new_[8087]_  = ~\new_[3388]_ ;
  assign \new_[8088]_  = ~\new_[2877]_ ;
  assign \new_[8089]_  = ~\new_[2862]_ ;
  assign \new_[8090]_  = ~\new_[2765]_ ;
  assign \new_[8091]_  = ~\new_[2776]_ ;
  assign \new_[8092]_  = ~\new_[2864]_ ;
  assign \new_[8093]_  = ~\new_[2414]_ ;
  assign \new_[8094]_  = ~\new_[2044]_ ;
  assign \new_[8095]_  = ~\new_[1236]_ ;
  assign \new_[8096]_  = ~\new_[1375]_ ;
  assign \new_[8097]_  = ~\key_i[4] ;
  assign \new_[8098]_  = ~\key_i[27] ;
  assign \new_[8099]_  = ~\new_[2762]_ ;
  assign \new_[8100]_  = ~\new_[2552]_ ;
  assign \new_[8101]_  = ~\new_[1558]_ ;
  assign \new_[8102]_  = ~\new_[2551]_ ;
  assign \new_[8103]_  = ~\new_[1959]_ ;
  assign \new_[8104]_  = ~\new_[3513]_ ;
  assign \new_[8105]_  = ~\new_[1993]_ ;
  assign \new_[8106]_  = ~\new_[1949]_ ;
  assign \new_[8107]_  = ~\new_[1946]_ ;
  assign \new_[8108]_  = ~\new_[5612]_ ;
  assign \new_[8109]_  = ~\new_[2034]_ ;
  assign \new_[8110]_  = ~\new_[2884]_ ;
  assign \new_[8111]_  = ~\new_[1761]_ ;
  assign \new_[8112]_  = ~\new_[2617]_ ;
  assign \new_[8113]_  = ~\new_[3981]_ ;
  assign \new_[8114]_  = ~\new_[2413]_ ;
  assign \new_[8115]_  = ~\new_[5659]_ ;
  assign \new_[8116]_  = ~\new_[2861]_ ;
  assign \new_[8117]_  = ~\new_[2619]_ ;
  assign \new_[8118]_  = ~\new_[2620]_ ;
  assign \new_[8119]_  = ~\new_[1128]_ ;
  assign \new_[8120]_  = ~\new_[1239]_ ;
  assign \new_[8121]_  = ~\new_[5784]_ ;
  assign \new_[8122]_  = ~\new_[2049]_ ;
  assign \new_[8123]_  = ~\key_i[13] ;
  assign \new_[8124]_  = ~\new_[2004]_ ;
  assign \new_[8125]_  = ~\new_[5377]_ ;
  assign \new_[8126]_  = ~\new_[2773]_ ;
  assign \new_[8127]_  = ~\new_[3381]_ ;
  assign \new_[8128]_  = ~\new_[2766]_ ;
  assign \new_[8129]_  = ~\new_[2770]_ ;
  assign \new_[8130]_  = ~\new_[1127]_ ;
  assign \new_[8131]_  = ~\key_i[24] ;
  assign \new_[8132]_  = ~\new_[3378]_ ;
  assign \new_[8133]_  = ~\new_[2953]_ ;
  assign \new_[8134]_  = ~\new_[1235]_ ;
  assign \new_[8135]_  = ~\key_i[0] ;
  assign \new_[8136]_  = ~\new_[2878]_ ;
  assign \new_[8137]_  = ~\new_[6952]_ ;
  assign \new_[8138]_  = ~\new_[2048]_ ;
  assign \new_[8139]_  = ~\new_[1942]_ ;
  assign \new_[8140]_  = ~\new_[1310]_ ;
  assign \new_[8141]_  = ~\new_[2045]_ ;
  assign \new_[8142]_  = ~\new_[1591]_ ;
  assign \new_[8143]_  = ~\new_[2544]_ ;
  assign \new_[8144]_  = ~\new_[2885]_ ;
  assign \new_[8145]_  = ~\new_[2931]_ ;
  assign \new_[8146]_  = ~\key_i[10] ;
  assign \new_[8147]_  = ~\new_[2936]_ ;
  assign \new_[8148]_  = ~\new_[1076]_ ;
  assign \new_[8149]_  = ~\new_[3001]_ ;
  assign \new_[8150]_  = ~\new_[2032]_ ;
  assign \new_[8151]_  = ~\new_[2025]_ ;
  assign \new_[8152]_  = ~\new_[3519]_ ;
  assign \new_[8153]_  = ~\key_i[29] ;
  assign \new_[8154]_  = ~\new_[2547]_ ;
  assign \new_[8155]_  = ~\new_[2880]_ ;
  assign \new_[8156]_  = ~\new_[2031]_ ;
  assign \new_[8157]_  = ~\new_[1387]_ ;
  assign \new_[8158]_  = ~\new_[1061]_ ;
  assign \new_[8159]_  = ~\key_i[18] ;
  assign \new_[8160]_  = ~\new_[4362]_ ;
  assign \new_[8161]_  = ~\new_[8162]_ ;
  assign \new_[8162]_  = \new_[8404]_ ;
  assign \new_[8163]_  = ~\new_[8180]_ ;
  assign \new_[8164]_  = ~\new_[8166]_ ;
  assign \new_[8165]_  = ~\new_[8166]_ ;
  assign \new_[8166]_  = ~\new_[8580]_ ;
  assign \new_[8167]_  = ~\new_[8580]_ ;
  assign \new_[8168]_  = ~\new_[8209]_ ;
  assign \new_[8169]_  = ~\new_[8170]_ ;
  assign \new_[8170]_  = \new_[8209]_ ;
  assign \new_[8171]_  = ~\new_[8172]_ ;
  assign \new_[8172]_  = \new_[8651]_ ;
  assign \new_[8173]_  = ~n850 | ~\new_[8174]_ ;
  assign \new_[8174]_  = (~\new_[7613]_  | ~\new_[9001]_ ) & (~\new_[4789]_  | ~\new_[8966]_ );
  assign \new_[8175]_  = ~\new_[8546]_  | ~\new_[8176]_  | ~\new_[8548]_ ;
  assign \new_[8176]_  = ~\new_[8174]_ ;
  assign \new_[8177]_  = ~\new_[8583]_  | ~\new_[8337]_ ;
  assign \new_[8178]_  = ~\new_[8322]_ ;
  assign \new_[8179]_  = ~\new_[8355]_ ;
  assign \new_[8180]_  = \new_[8479]_ ;
  assign \new_[8181]_  = ~\new_[8975]_ ;
  assign \new_[8182]_  = ~\new_[8810]_  | ~\new_[1592]_ ;
  assign \new_[8183]_  = ~\new_[7863]_  & ~\new_[7659]_ ;
  assign \new_[8184]_  = ~\new_[7625]_  & ~\new_[7834]_ ;
  assign \new_[8185]_  = ~\new_[1067]_  | ~\new_[1069]_ ;
  assign \new_[8186]_  = ~\new_[8961]_  | ~\new_[4335]_ ;
  assign \new_[8187]_  = ~\new_[8964]_  | ~\new_[7103]_ ;
  assign \new_[8188]_  = ~\new_[8961]_  | ~\new_[4340]_ ;
  assign \new_[8189]_  = ~\new_[8963]_  | ~\new_[7094]_ ;
  assign \new_[8190]_  = ~\new_[8229]_  | ~\new_[8230]_ ;
  assign \new_[8191]_  = ~\new_[8725]_  & ~\new_[8553]_ ;
  assign \new_[8192]_  = ~\new_[8625]_ ;
  assign \new_[8193]_  = ~\new_[5293]_  | ~\new_[5419]_ ;
  assign \new_[8194]_  = \new_[5377]_  | \new_[5307]_ ;
  assign \new_[8195]_  = ~\new_[5293]_ ;
  assign \new_[8196]_  = ~\new_[5419]_ ;
  assign \new_[8197]_  = ~\new_[8198]_ ;
  assign \new_[8198]_  = (~\new_[5490]_  & ~\new_[5856]_ ) | (~\new_[5557]_  & ~\new_[5797]_ );
  assign \new_[8199]_  = \new_[5142]_  ? \new_[8749]_  : \new_[5248]_ ;
  assign n835 = ~\new_[8201]_  | ~\new_[8205]_ ;
  assign \new_[8201]_  = ~\new_[8843]_  | ~\new_[8202]_  | ~\new_[8203]_ ;
  assign \new_[8202]_  = \new_[8803]_  | n995;
  assign \new_[8203]_  = ~\new_[8803]_  | ~n995;
  assign \new_[8204]_  = \new_[4230]_  | \new_[8160]_ ;
  assign \new_[8205]_  = ~\new_[7486]_  | ~\new_[1076]_ ;
  assign \new_[8206]_  = ~\new_[8885]_ ;
  assign \new_[8207]_  = \new_[8163]_  ^ \new_[8411]_ ;
  assign \new_[8208]_  = \new_[8892]_  ? \new_[4361]_  : \new_[8886]_ ;
  assign \new_[8209]_  = ~\new_[8213]_  | ~\new_[8210]_  | ~\new_[8212]_ ;
  assign \new_[8210]_  = ~\new_[8191]_  | ~\new_[8211]_ ;
  assign \new_[8211]_  = ~\new_[2035]_  | ~\new_[2008]_ ;
  assign \new_[8212]_  = ~\new_[8624]_  | ~\new_[2035]_  | ~\new_[2008]_ ;
  assign \new_[8213]_  = \new_[8373]_  | \new_[4542]_ ;
  assign \new_[8214]_  = \new_[8192]_  ? \new_[8366]_  : \new_[8331]_ ;
  assign \new_[8215]_  = \new_[8216]_  ? \new_[8629]_  : \new_[8877]_ ;
  assign \new_[8216]_  = \new_[4464]_  ? \new_[8363]_  : \new_[4542]_ ;
  assign \new_[8217]_  = ~\new_[8265]_  | ~\new_[8266]_ ;
  assign \new_[8218]_  = ~\new_[1953]_  | ~\new_[1967]_ ;
  assign \new_[8219]_  = ~\new_[8434]_ ;
  assign \new_[8220]_  = \new_[8185]_  ? \new_[7664]_  : \new_[7828]_ ;
  assign \new_[8221]_  = ~\new_[8220]_ ;
  assign \new_[8222]_  = ~\new_[7122]_  | ~\new_[6958]_ ;
  assign \new_[8223]_  = ~\new_[9007]_  | ~\new_[7828]_ ;
  assign \new_[8224]_  = ~\new_[8185]_  | ~\new_[9008]_ ;
  assign \new_[8225]_  = ~\new_[8226]_ ;
  assign \new_[8226]_  = \new_[8566]_  ? \new_[8591]_  : \new_[5669]_ ;
  assign \new_[8227]_  = \new_[5845]_  ? \new_[5381]_  : \new_[5911]_ ;
  assign \new_[8228]_  = ~\new_[8229]_  | ~\new_[8230]_ ;
  assign \new_[8229]_  = ~\new_[1943]_  | ~\new_[8538]_ ;
  assign \new_[8230]_  = ~\new_[8337]_  | ~\new_[9003]_ ;
  assign \new_[8231]_  = \new_[8188]_  & \new_[8189]_ ;
  assign \new_[8232]_  = ~\new_[8434]_  & ~\new_[8655]_ ;
  assign \new_[8233]_  = ~\new_[8553]_  | ~\new_[2089]_ ;
  assign \new_[8234]_  = ~\new_[8625]_  | ~\new_[8854]_ ;
  assign \new_[8235]_  = (~\new_[8909]_  | ~\new_[8239]_ ) & (~\new_[8932]_  | ~\new_[1139]_ );
  assign \new_[8236]_  = ~\new_[8237]_  & ~\new_[8238]_ ;
  assign \new_[8237]_  = ~decrypt_i;
  assign \new_[8238]_  = ~\new_[8193]_  & ~\new_[8194]_ ;
  assign \new_[8239]_  = \data_i[93]  ? \new_[6778]_  : \new_[6448]_ ;
  assign \new_[8240]_  = \new_[8241]_  | \new_[8242]_ ;
  assign \new_[8241]_  = \new_[5253]_  & \key_i[14] ;
  assign \new_[8242]_  = ~\new_[5203]_  & (~\new_[6539]_  | ~\new_[6815]_ );
  assign \new_[8243]_  = \new_[8244]_  & \new_[9001]_ ;
  assign \new_[8244]_  = ~\new_[7589]_  | ~\new_[7654]_ ;
  assign \new_[8245]_  = ~\new_[4431]_  | ~\new_[8422]_ ;
  assign \new_[8246]_  = ~\new_[8247]_  & (~\new_[8396]_  | ~\new_[8424]_ );
  assign \new_[8247]_  = ~\new_[7688]_  & ~\new_[8278]_ ;
  assign \new_[8248]_  = ~\new_[8249]_  | ~\new_[8378]_ ;
  assign \new_[8249]_  = ~\new_[8357]_ ;
  assign \new_[8250]_  = ~\new_[8254]_  | (~\new_[8251]_  & ~\new_[8252]_ );
  assign \new_[8251]_  = ~\new_[5201]_  & (~\new_[6529]_  | ~\new_[6813]_ );
  assign \new_[8252]_  = ~\new_[8253]_  | ~\new_[8880]_ ;
  assign \new_[8253]_  = ~\new_[5253]_  | ~\key_i[6] ;
  assign \new_[8254]_  = \new_[8966]_  | \new_[8255]_ ;
  assign \new_[8255]_  = ~\new_[7595]_  | ~\new_[7653]_ ;
  assign \new_[8256]_  = ~\new_[7618]_  | ~\new_[7634]_ ;
  assign \new_[8257]_  = ~\new_[8272]_  | ~\new_[8258]_  | ~\new_[8273]_ ;
  assign \new_[8258]_  = ~\new_[8274]_ ;
  assign \new_[8259]_  = \new_[8260]_ ;
  assign \new_[8260]_  = ~\new_[8261]_  | ~\new_[8263]_ ;
  assign \new_[8261]_  = ~\new_[8262]_  | ~\new_[8373]_ ;
  assign \new_[8262]_  = ~\new_[8233]_  | ~\new_[8234]_ ;
  assign \new_[8263]_  = ~\new_[8725]_  | ~\new_[8363]_ ;
  assign \new_[8264]_  = ~\new_[8265]_  | ~\new_[8266]_ ;
  assign \new_[8265]_  = ~\new_[8218]_  | ~\new_[8219]_ ;
  assign \new_[8266]_  = ~\new_[8370]_  | ~\new_[8434]_ ;
  assign \new_[8267]_  = \new_[8186]_  & \new_[8187]_ ;
  assign \new_[8268]_  = ~\new_[8288]_  | ~\new_[8269]_  | ~\new_[8289]_ ;
  assign \new_[8269]_  = ~\new_[8290]_ ;
  assign \new_[8270]_  = ~\new_[8271]_  | ~\new_[8274]_ ;
  assign \new_[8271]_  = ~\new_[8272]_  | ~\new_[8273]_ ;
  assign \new_[8272]_  = ~\new_[1897]_  | ~\new_[3358]_ ;
  assign \new_[8273]_  = ~\new_[8228]_  | ~\new_[8231]_ ;
  assign \new_[8274]_  = \new_[8275]_  & \new_[8276]_ ;
  assign \new_[8275]_  = ~\new_[4154]_  | ~\new_[8960]_ ;
  assign \new_[8276]_  = ~\new_[8954]_  | ~\new_[7047]_ ;
  assign \new_[8277]_  = ~\new_[4893]_  | (~\new_[4794]_  & ~\new_[9001]_ );
  assign \new_[8278]_  = ~\new_[8282]_  & (~\new_[8279]_  | ~\new_[8965]_ );
  assign \new_[8279]_  = ~\new_[8281]_  | (~\new_[8280]_  & ~\new_[8307]_ );
  assign \new_[8280]_  = ~\new_[6711]_  & (~\new_[1979]_  | ~\new_[8988]_ );
  assign \new_[8281]_  = ~\new_[8307]_  | ~\key_i[19] ;
  assign \new_[8282]_  = ~\new_[8283]_  & ~\new_[8965]_ ;
  assign \new_[8283]_  = ~\new_[8284]_ ;
  assign \new_[8284]_  = (~\new_[7860]_  & ~\new_[8013]_ ) | (~\new_[7897]_  & ~\new_[8285]_ );
  assign \new_[8285]_  = ~\key_i[19] ;
  assign \new_[8286]_  = ~\new_[8287]_  | ~\new_[8290]_ ;
  assign \new_[8287]_  = ~\new_[8288]_  | ~\new_[8289]_ ;
  assign \new_[8288]_  = ~\new_[8986]_  | ~\new_[3357]_ ;
  assign \new_[8289]_  = ~\new_[8264]_  | ~\new_[8267]_ ;
  assign \new_[8290]_  = \new_[8291]_  & \new_[8292]_ ;
  assign \new_[8291]_  = ~\new_[4153]_  | ~\new_[8965]_ ;
  assign \new_[8292]_  = ~\new_[8954]_  | ~\new_[7061]_ ;
  assign \new_[8293]_  = ~\new_[8294]_ ;
  assign \new_[8294]_  = ~\new_[8295]_  | (~\new_[7747]_  & ~\new_[7816]_ );
  assign \new_[8295]_  = \new_[8663]_  | \new_[8802]_ ;
  assign \new_[8296]_  = \new_[7566]_  ? \new_[6158]_  : \new_[7496]_ ;
  assign \new_[8297]_  = ~\new_[8301]_  | (~\new_[8298]_  & ~\new_[8299]_ );
  assign \new_[8298]_  = ~\new_[5201]_  & (~\new_[6538]_  | ~\new_[6819]_ );
  assign \new_[8299]_  = ~\new_[8300]_  | ~\new_[8880]_ ;
  assign \new_[8300]_  = ~\new_[5253]_  | ~\key_i[22] ;
  assign \new_[8301]_  = \new_[8966]_  | \new_[8302]_ ;
  assign \new_[8302]_  = ~\new_[7591]_  | ~\new_[7727]_ ;
  assign \new_[8303]_  = ~\new_[7637]_  | ~\new_[7681]_ ;
  assign \new_[8304]_  = ~\new_[9001]_  & (~\new_[8305]_  | ~\new_[8309]_ );
  assign \new_[8305]_  = ~\new_[8306]_ ;
  assign \new_[8306]_  = ~\new_[8307]_  & (~\new_[6705]_  | ~\new_[6821]_ );
  assign \new_[8307]_  = ~\new_[8308]_ ;
  assign \new_[8308]_  = ~\new_[8401]_ ;
  assign \new_[8309]_  = \new_[7967]_  | \new_[8727]_ ;
  assign \new_[8310]_  = ~\new_[8882]_  | ~\new_[5488]_ ;
  assign \new_[8311]_  = ~\new_[8324]_ ;
  assign \new_[8312]_  = ~\new_[8314]_  & (~\new_[8313]_  | ~\new_[8967]_ );
  assign \new_[8313]_  = ~\new_[7616]_  | ~\new_[7768]_ ;
  assign \new_[8314]_  = ~\new_[8967]_  & (~\new_[8315]_  | ~\new_[8317]_ );
  assign \new_[8315]_  = ~\new_[8316]_ ;
  assign \new_[8316]_  = ~\new_[5201]_  & (~\new_[6530]_  | ~\new_[6817]_ );
  assign \new_[8317]_  = ~\new_[5201]_  | ~\key_i[20] ;
  assign n785 = ~\new_[8319]_  | ~\new_[8320]_ ;
  assign \new_[8319]_  = ~\new_[8321]_  | ~\new_[8843]_ ;
  assign \new_[8320]_  = ~\new_[7384]_  | ~\new_[1062]_ ;
  assign \new_[8321]_  = \new_[8178]_  ? n845 : \new_[8322]_ ;
  assign \new_[8322]_  = ~\new_[8323]_  & (~\new_[4788]_  | ~\new_[9000]_ );
  assign \new_[8323]_  = \new_[9001]_  & \new_[7610]_ ;
  assign \new_[8324]_  = ~\new_[8323]_  & (~\new_[4788]_  | ~\new_[9000]_ );
  assign \new_[8325]_  = ~\new_[8607]_ ;
  assign \new_[8326]_  = ~\new_[8327]_  | ~\new_[8328]_ ;
  assign \new_[8327]_  = ~\new_[4791]_  | ~\new_[8966]_ ;
  assign \new_[8328]_  = ~\new_[8967]_  | ~\new_[7423]_ ;
  assign \new_[8329]_  = \new_[7879]_  & \new_[4230]_ ;
  assign \new_[8330]_  = ~\new_[8326]_ ;
  assign \new_[8331]_  = ~\new_[8332]_  | (~\new_[2216]_  & ~\new_[8373]_ );
  assign \new_[8332]_  = \new_[8333]_  ? \new_[8629]_  : \new_[8334]_ ;
  assign \new_[8333]_  = \new_[8337]_  | \new_[8626]_ ;
  assign \new_[8334]_  = ~\new_[8626]_  | ~\new_[8373]_ ;
  assign \new_[8335]_  = ~\new_[8336]_  | ~\new_[8338]_ ;
  assign \new_[8336]_  = ~\new_[8337]_  & (~\new_[2090]_  | ~\new_[8553]_ );
  assign \new_[8337]_  = ~\new_[8373]_ ;
  assign \new_[8338]_  = ~\new_[8625]_  | ~\new_[8339]_ ;
  assign \new_[8339]_  = ~\new_[2302]_  | ~\new_[2301]_ ;
  assign n780 = ~\new_[8341]_  | ~\new_[8342]_ ;
  assign \new_[8341]_  = ~\new_[8354]_  | ~\new_[8852]_ ;
  assign \new_[8342]_  = ~\new_[7384]_  | ~\new_[1061]_ ;
  assign \new_[8343]_  = ~\new_[8853]_ ;
  assign \new_[8344]_  = ~\new_[8345]_  & (~\new_[8167]_  | ~\new_[8362]_ );
  assign \new_[8345]_  = ~\new_[8655]_  | ~\new_[8724]_ ;
  assign \new_[8346]_  = ~\new_[8373]_  & ~\new_[8856]_ ;
  assign \new_[8347]_  = ~\new_[8353]_  | ~\new_[8348]_  | ~\new_[8350]_ ;
  assign \new_[8348]_  = ~\new_[8383]_  | ~\new_[8349]_ ;
  assign \new_[8349]_  = ~\new_[8724]_  & ~\new_[8487]_ ;
  assign \new_[8350]_  = ~\new_[8352]_  | ~\new_[8351]_  | ~\new_[8487]_ ;
  assign \new_[8351]_  = ~\new_[8383]_ ;
  assign \new_[8352]_  = ~\new_[8724]_ ;
  assign \new_[8353]_  = ~\new_[8720]_  | ~\new_[8724]_ ;
  assign \new_[8354]_  = \new_[8179]_  ? n840 : \new_[8355]_ ;
  assign \new_[8355]_  = ~\new_[8356]_  & (~\new_[8958]_  | ~\new_[4787]_ );
  assign \new_[8356]_  = \new_[9001]_  & \new_[7471]_ ;
  assign \new_[8357]_  = ~\new_[8356]_  & (~\new_[4787]_  | ~\new_[8965]_ );
  assign \new_[8358]_  = ~\new_[4891]_  | (~\new_[4781]_  & ~\new_[9001]_ );
  assign \new_[8359]_  = ~\new_[8360]_  | ~\new_[8365]_ ;
  assign \new_[8360]_  = ~\new_[8361]_ ;
  assign \new_[8361]_  = ~\new_[8362]_  & ~\new_[8364]_ ;
  assign \new_[8362]_  = \new_[8363]_ ;
  assign \new_[8363]_  = ~\new_[3002]_  | ~\new_[3235]_ ;
  assign \new_[8364]_  = ~\new_[8580]_ ;
  assign \new_[8365]_  = ~\new_[8167]_  | ~\new_[8362]_ ;
  assign \new_[8366]_  = ~\new_[8373]_  | ~\new_[8367]_  | ~\new_[8371]_ ;
  assign \new_[8367]_  = ~\new_[8368]_  | ~\new_[8370]_ ;
  assign \new_[8368]_  = ~\new_[8369]_ ;
  assign \new_[8369]_  = \new_[8855]_  ? \new_[8973]_  : \new_[8206]_ ;
  assign \new_[8370]_  = \new_[8584]_ ;
  assign \new_[8371]_  = ~\new_[8369]_  | ~\new_[8372]_ ;
  assign \new_[8372]_  = ~\new_[8370]_ ;
  assign \new_[8373]_  = \new_[8724]_ ;
  assign \new_[8374]_  = ~\new_[8375]_  | ~\new_[8380]_  | ~\new_[8381]_  | ~\new_[8379]_ ;
  assign \new_[8375]_  = ~\new_[8376]_  | ~\new_[8378]_ ;
  assign \new_[8376]_  = ~\new_[8377]_ ;
  assign \new_[8377]_  = ~\new_[8243]_  & (~\new_[8240]_  | ~\new_[8965]_ );
  assign \new_[8378]_  = \new_[7925]_  & \new_[7536]_ ;
  assign \new_[8379]_  = ~\new_[4434]_  | ~\new_[8422]_ ;
  assign \new_[8380]_  = ~\new_[4439]_  | ~\new_[8329]_ ;
  assign \new_[8381]_  = ~\new_[8358]_  | ~\new_[8424]_ ;
  assign \new_[8382]_  = ~\new_[8376]_ ;
  assign \new_[8383]_  = ~\new_[8384]_  | ~\new_[8386]_ ;
  assign \new_[8384]_  = ~\new_[2666]_  | ~\new_[8385]_ ;
  assign \new_[8385]_  = ~\new_[3508]_  | ~\new_[4321]_ ;
  assign \new_[8386]_  = ~\new_[8387]_  | ~\new_[8388]_ ;
  assign \new_[8387]_  = ~\new_[8385]_ ;
  assign \new_[8388]_  = ~\new_[3043]_  | ~\new_[4325]_ ;
  assign \new_[8389]_  = ~\new_[8395]_  | ~\new_[8390]_  | ~\new_[8394]_ ;
  assign \new_[8390]_  = ~\new_[8391]_  & (~\new_[8326]_  | ~\new_[8329]_ );
  assign \new_[8391]_  = ~\new_[7826]_  & ~\new_[8392]_ ;
  assign \new_[8392]_  = ~\new_[8393]_  & (~\new_[4889]_  | ~\new_[9002]_ );
  assign \new_[8393]_  = \new_[9001]_  & \new_[7574]_ ;
  assign \new_[8394]_  = ~\new_[8277]_  | ~\new_[8424]_ ;
  assign \new_[8395]_  = ~\new_[8803]_  | ~\new_[8378]_ ;
  assign \new_[8396]_  = ~\new_[8400]_  | (~\new_[8397]_  & ~\new_[9001]_ );
  assign \new_[8397]_  = (~\key_i[27]  | ~\new_[5203]_ ) & (~\new_[8398]_  | ~\new_[8727]_ );
  assign \new_[8398]_  = ~\new_[8399]_  | (~\new_[8997]_  & ~\new_[7590]_ );
  assign \new_[8399]_  = \new_[8107]_  | \new_[8998]_ ;
  assign \new_[8400]_  = \new_[7590]_  | \new_[8965]_ ;
  assign \new_[8401]_  = ~\new_[8728]_ ;
  assign \new_[8402]_  = ~\new_[8403]_ ;
  assign \new_[8403]_  = \new_[4346]_  ? \new_[8954]_  : \new_[7049]_ ;
  assign \new_[8404]_  = ~\new_[8405]_  | ~\new_[8406]_ ;
  assign \new_[8405]_  = ~\new_[8359]_  | ~\new_[8232]_ ;
  assign \new_[8406]_  = ~\new_[8346]_  & (~\new_[8360]_  | ~\new_[8344]_ );
  assign n790 = ~\new_[8408]_  | ~\new_[8410]_ ;
  assign \new_[8408]_  = ~\new_[8409]_  | ~\new_[8843]_ ;
  assign \new_[8409]_  = ~\new_[8173]_  | ~\new_[8175]_ ;
  assign \new_[8410]_  = ~\new_[7384]_  | ~\new_[1063]_ ;
  assign \new_[8411]_  = ~\new_[4995]_  | ~\new_[4994]_ ;
  assign \new_[8412]_  = ~\new_[8824]_  | ~\new_[3408]_ ;
  assign \new_[8413]_  = \new_[8414]_  ? \new_[8479]_  : \new_[5424]_ ;
  assign \new_[8414]_  = ~\new_[1592]_  | ~\new_[8952]_ ;
  assign \new_[8415]_  = ~\new_[8421]_  | ~\new_[8416]_  | ~\new_[8420]_ ;
  assign \new_[8416]_  = ~\new_[8417]_  & (~\new_[8311]_  | ~\new_[8378]_ );
  assign \new_[8417]_  = ~\new_[8418]_  & ~\new_[9016]_ ;
  assign \new_[8418]_  = ~\new_[8419]_ ;
  assign \new_[8419]_  = \new_[4934]_  & \new_[7843]_ ;
  assign \new_[8420]_  = ~\new_[4437]_  | ~\new_[8329]_ ;
  assign \new_[8421]_  = ~\new_[8422]_  | ~\new_[8423]_ ;
  assign \new_[8422]_  = \new_[7899]_  & \new_[7536]_ ;
  assign \new_[8423]_  = ~\new_[4939]_  | (~\new_[4784]_  & ~\new_[9001]_ );
  assign \new_[8424]_  = ~\new_[8418]_ ;
  assign \new_[8425]_  = ~\new_[8426]_  | ~\new_[8427]_ ;
  assign \new_[8426]_  = ~\new_[8445]_  | ~\new_[8518]_ ;
  assign \new_[8427]_  = ~\new_[8706]_  | ~\new_[8446]_ ;
  assign \new_[8428]_  = ~\new_[8445]_ ;
  assign \new_[8429]_  = ~\new_[8430]_ ;
  assign \new_[8430]_  = ~\new_[2091]_  | ~\new_[2357]_ ;
  assign \new_[8431]_  = ~\new_[1971]_  | ~\new_[1957]_ ;
  assign \new_[8432]_  = ~\new_[8431]_ ;
  assign \new_[8433]_  = ~\new_[8449]_  & ~\new_[8434]_ ;
  assign \new_[8434]_  = ~\new_[8373]_ ;
  assign \new_[8435]_  = \new_[8436]_  | \new_[8438]_ ;
  assign \new_[8436]_  = ~\new_[8713]_  & (~\new_[8716]_  | ~\new_[8437]_ );
  assign \new_[8437]_  = ~\new_[2345]_ ;
  assign \new_[8438]_  = ~\new_[8439]_  & (~\new_[6162]_  | ~\new_[3864]_ );
  assign \new_[8439]_  = ~\new_[2345]_  & (~\new_[8440]_  | ~\new_[8710]_ );
  assign \new_[8440]_  = ~\new_[8716]_ ;
  assign \new_[8441]_  = \new_[8442]_  ? \new_[8831]_  : \new_[8443]_ ;
  assign \new_[8442]_  = \new_[8858]_  ^ \new_[8666]_ ;
  assign \new_[8443]_  = ~\new_[8442]_ ;
  assign \new_[8444]_  = \new_[8442]_ ;
  assign \new_[8445]_  = \new_[8446]_  ? \new_[8706]_  : \new_[8518]_ ;
  assign \new_[8446]_  = ~\new_[8518]_ ;
  assign \new_[8447]_  = ~\new_[8448]_  | ~\new_[8450]_ ;
  assign \new_[8448]_  = ~\new_[8449]_  | ~\new_[8720]_ ;
  assign \new_[8449]_  = \new_[8488]_  & \new_[8492]_ ;
  assign \new_[8450]_  = ~\new_[8723]_  | ~\new_[8487]_ ;
  assign \new_[8451]_  = (~\new_[8784]_  | ~\new_[6552]_ ) & (~\new_[6396]_  | ~\new_[8780]_ );
  assign \new_[8452]_  = ~\new_[6391]_  & ~\new_[6201]_ ;
  assign \new_[8453]_  = \new_[8454]_  ? \new_[8456]_  : \new_[8455]_ ;
  assign \new_[8454]_  = ~\new_[8455]_ ;
  assign \new_[8455]_  = (~\new_[8430]_  | ~\new_[8432]_ ) & (~\new_[8431]_  | ~\new_[8429]_ );
  assign \new_[8456]_  = ~\new_[8679]_  & (~\new_[8674]_  | ~\new_[8673]_ );
  assign \new_[8457]_  = \new_[5916]_  ? \new_[5613]_  : \new_[5852]_ ;
  assign \new_[8458]_  = \new_[5912]_  ? \new_[5482]_  : \new_[5846]_ ;
  assign \new_[8459]_  = ~\new_[8462]_  & (~\new_[8460]_  | ~\new_[8713]_ );
  assign \new_[8460]_  = ~\new_[8461]_  | (~\new_[8710]_  & ~\new_[2227]_ );
  assign \new_[8461]_  = ~\new_[6161]_  | ~\new_[3652]_ ;
  assign \new_[8462]_  = \new_[8716]_  & \new_[8463]_ ;
  assign \new_[8463]_  = ~\new_[2227]_ ;
  assign \new_[8464]_  = ~\new_[8467]_  & (~\new_[8465]_  | ~\new_[8713]_ );
  assign \new_[8465]_  = ~\new_[8466]_  | (~\new_[8710]_  & ~\new_[2225]_ );
  assign \new_[8466]_  = ~\new_[6160]_  | ~\new_[3648]_ ;
  assign \new_[8467]_  = \new_[8716]_  & \new_[8468]_ ;
  assign \new_[8468]_  = ~\new_[2225]_ ;
  assign \new_[8469]_  = ~\new_[8710]_ ;
  assign \new_[8470]_  = ~\new_[5664]_ ;
  assign \new_[8471]_  = \new_[5834]_  ^ \new_[5835]_ ;
  assign \new_[8472]_  = ~\new_[8471]_ ;
  assign \new_[8473]_  = \new_[5608]_  ^ \new_[5609]_ ;
  assign \new_[8474]_  = ~\new_[8477]_  & (~\new_[8475]_  | ~\new_[8713]_ );
  assign \new_[8475]_  = ~\new_[8476]_  | (~\new_[8710]_  & ~\new_[2226]_ );
  assign \new_[8476]_  = ~\new_[6160]_  | ~\new_[3650]_ ;
  assign \new_[8477]_  = \new_[8716]_  & \new_[8478]_ ;
  assign \new_[8478]_  = ~\new_[2226]_ ;
  assign \new_[8479]_  = \new_[8480]_  ^ \new_[8481]_ ;
  assign \new_[8480]_  = \new_[8976]_  ? \new_[8182]_  : \new_[8181]_ ;
  assign \new_[8481]_  = \new_[8482]_  ? \new_[8483]_  : \new_[8528]_ ;
  assign \new_[8482]_  = ~\new_[8528]_ ;
  assign \new_[8483]_  = ~\new_[8809]_  | ~\new_[1467]_ ;
  assign \new_[8484]_  = ~\new_[8486]_  & (~\new_[8772]_  | ~\new_[8485]_ );
  assign \new_[8485]_  = ~\new_[5760]_  | ~\new_[5802]_ ;
  assign \new_[8486]_  = ~\new_[8485]_  & ~\new_[8772]_ ;
  assign \new_[8487]_  = ~\new_[8488]_  | ~\new_[8492]_ ;
  assign \new_[8488]_  = ~\new_[8489]_  | ~\new_[8491]_ ;
  assign \new_[8489]_  = ~\new_[8490]_ ;
  assign \new_[8490]_  = ~\new_[8419]_  & (~\new_[7823]_  | ~\new_[7881]_ );
  assign \new_[8491]_  = ~\new_[8246]_  | ~\new_[8245]_  | ~\new_[8248]_ ;
  assign \new_[8492]_  = ~\new_[8493]_  | ~\new_[8490]_ ;
  assign \new_[8493]_  = ~\new_[5666]_ ;
  assign \new_[8494]_  = \new_[8495]_ ;
  assign \new_[8495]_  = ~\new_[8502]_  & (~\new_[8496]_  | ~\new_[8498]_ );
  assign \new_[8496]_  = \new_[5661]_  ? \new_[5468]_  : \new_[8497]_ ;
  assign \new_[8497]_  = ~\new_[5661]_ ;
  assign \new_[8498]_  = \new_[8499]_  ? \new_[8501]_  : \new_[8500]_ ;
  assign \new_[8499]_  = \new_[5833]_  ^ \new_[5836]_ ;
  assign \new_[8500]_  = ~\new_[8499]_ ;
  assign \new_[8501]_  = \new_[8864]_  ^ \new_[8870]_ ;
  assign \new_[8502]_  = ~\new_[8498]_  & ~\new_[8496]_ ;
  assign \new_[8503]_  = ~\new_[8511]_  & (~\new_[8504]_  | ~\new_[8510]_ );
  assign \new_[8504]_  = ~\new_[8507]_  | ~\new_[8505]_  | ~\new_[8506]_ ;
  assign \new_[8505]_  = ~\new_[5879]_ ;
  assign \new_[8506]_  = ~\new_[5875]_ ;
  assign \new_[8507]_  = \new_[8508]_  & \new_[8509]_ ;
  assign \new_[8508]_  = ~\new_[8779]_  | ~\new_[5978]_ ;
  assign \new_[8509]_  = ~\new_[5975]_  | ~\new_[8558]_ ;
  assign \new_[8510]_  = ~\new_[5766]_  | ~\new_[5759]_ ;
  assign \new_[8511]_  = ~\new_[8510]_  & ~\new_[8504]_ ;
  assign \new_[8512]_  = \new_[8513]_  ? \new_[8515]_  : \new_[8514]_ ;
  assign \new_[8513]_  = \new_[2014]_  ^ \new_[8680]_ ;
  assign \new_[8514]_  = ~\new_[8513]_ ;
  assign \new_[8515]_  = \new_[1987]_  ? \new_[1930]_  : \new_[8429]_ ;
  assign \new_[8516]_  = ~\new_[8979]_  | ~\new_[8707]_ ;
  assign \new_[8517]_  = ~\new_[2015]_  & ~\new_[8680]_ ;
  assign \new_[8518]_  = ~\new_[8673]_ ;
  assign \new_[8519]_  = ~\new_[8520]_  | ~\new_[8784]_ ;
  assign \new_[8520]_  = \data_o[27]  ? \new_[8912]_  : \new_[1244]_ ;
  assign \new_[8521]_  = ~\new_[5968]_  & (~\new_[8522]_  | ~\new_[8558]_ );
  assign \new_[8522]_  = \data_o[91]  ? \new_[8934]_  : \new_[1251]_ ;
  assign \new_[8523]_  = \new_[8524]_  ? \new_[8526]_  : \new_[8525]_ ;
  assign \new_[8524]_  = \new_[5664]_  ? \new_[5472]_  : \new_[8470]_ ;
  assign \new_[8525]_  = ~\new_[8524]_ ;
  assign \new_[8526]_  = \new_[8471]_  ? \new_[8473]_  : \new_[8472]_ ;
  assign \new_[8527]_  = \new_[8524]_ ;
  assign \new_[8528]_  = ~\new_[8569]_  | ~\new_[1866]_ ;
  assign \new_[8529]_  = ~\new_[6039]_  | ~\new_[8779]_ ;
  assign \new_[8530]_  = ~\new_[8531]_  | ~\new_[8784]_ ;
  assign \new_[8531]_  = \data_o[3]  ? \new_[8924]_  : \new_[1217]_ ;
  assign \new_[8532]_  = ~\new_[8533]_  & ~\new_[5931]_ ;
  assign \new_[8533]_  = ~\new_[7902]_  & (~\new_[6119]_  | ~\new_[6214]_ );
  assign \new_[8534]_  = ~\new_[8541]_  & (~\new_[8535]_  | ~\new_[8539]_ );
  assign \new_[8535]_  = ~\new_[8433]_  & ~\new_[8536]_ ;
  assign \new_[8536]_  = ~\new_[2665]_  | ~\new_[8537]_ ;
  assign \new_[8537]_  = \new_[8538]_  | \new_[2218]_ ;
  assign \new_[8538]_  = \new_[8373]_ ;
  assign \new_[8539]_  = ~\new_[8540]_ ;
  assign \new_[8540]_  = ~\new_[8538]_  & ~\new_[2063]_ ;
  assign \new_[8541]_  = \new_[8677]_  & \new_[8536]_ ;
  assign n850 = ~\new_[8543]_  | ~\new_[8546]_ ;
  assign \new_[8543]_  = ~\new_[8544]_  | ~n1020;
  assign \new_[8544]_  = ~\new_[3570]_  & ~\new_[3525]_ ;
  assign n1020 = ~\new_[1587]_  | ~\new_[1691]_ ;
  assign \new_[8546]_  = ~\new_[1587]_  | ~\new_[8547]_  | ~\new_[1691]_ ;
  assign \new_[8547]_  = ~\new_[8544]_ ;
  assign \new_[8548]_  = ~n1020 | ~\new_[8544]_ ;
  assign n845 = \new_[8550]_  ^ n1000;
  assign \new_[8550]_  = ~\new_[8551]_ ;
  assign \new_[8551]_  = ~\new_[2974]_  & (~\new_[3983]_  | ~\new_[6063]_ );
  assign n1000 = ~\new_[8270]_  | ~\new_[8257]_ ;
  assign \new_[8553]_  = \new_[8627]_  ? \new_[8555]_  : \new_[8626]_ ;
  assign \new_[8554]_  = ~\new_[8207]_ ;
  assign \new_[8555]_  = \new_[8556]_  & \new_[8659]_ ;
  assign \new_[8556]_  = ~\new_[8206]_  | ~\new_[4735]_ ;
  assign \new_[8557]_  = \data_o[75]  ? \new_[8904]_  : \new_[1199]_ ;
  assign \new_[8558]_  = ~\new_[5659]_  & ~\new_[8108]_ ;
  assign \new_[8559]_  = ~\new_[8560]_ ;
  assign \new_[8560]_  = ~\new_[5967]_  & (~\new_[8561]_  | ~\new_[8784]_ );
  assign \new_[8561]_  = \data_o[11]  ? \new_[8924]_  : \new_[1193]_ ;
  assign \new_[8562]_  = ~\new_[8558]_ ;
  assign \new_[8563]_  = ~\new_[8784]_ ;
  assign \new_[8564]_  = ~\new_[6102]_  & (~\new_[6406]_  | ~\new_[8780]_ );
  assign \new_[8565]_  = ~\new_[6195]_  & (~\new_[6397]_  | ~\new_[8558]_ );
  assign \new_[8566]_  = ~\new_[1709]_  | ~\new_[8567]_  | ~\new_[8568]_ ;
  assign \new_[8567]_  = \new_[8969]_  | \new_[9006]_ ;
  assign \new_[8568]_  = ~\new_[9006]_  | ~\new_[8971]_ ;
  assign \new_[8569]_  = \new_[8570]_  ? \new_[8572]_  : \new_[8571]_ ;
  assign \new_[8570]_  = ~\new_[8571]_ ;
  assign \new_[8571]_  = ~\new_[8183]_  & ~\new_[8184]_ ;
  assign \new_[8572]_  = \new_[8798]_  ? \new_[8662]_  : \new_[8573]_ ;
  assign \new_[8573]_  = ~\new_[8798]_ ;
  assign n840 = \new_[8575]_  ^ n1005;
  assign \new_[8575]_  = ~\new_[8576]_ ;
  assign \new_[8576]_  = ~\new_[2973]_  & (~\new_[3983]_  | ~\new_[6139]_ );
  assign n1005 = ~\new_[8286]_  | ~\new_[8268]_ ;
  assign \new_[8578]_  = ~\new_[8579]_  | ~\new_[8626]_ ;
  assign \new_[8579]_  = ~\new_[8580]_ ;
  assign \new_[8580]_  = ~\new_[8581]_ ;
  assign \new_[8581]_  = \new_[8582]_  ? \new_[8584]_  : \new_[8583]_ ;
  assign \new_[8582]_  = ~\new_[8583]_ ;
  assign \new_[8583]_  = \new_[8824]_  & \new_[3408]_ ;
  assign \new_[8584]_  = \new_[8197]_  ? \new_[8199]_  : \new_[8198]_ ;
  assign \new_[8585]_  = ~\new_[8626]_ ;
  assign \new_[8586]_  = ~\new_[8589]_  & (~\new_[8587]_  | ~\new_[8713]_ );
  assign \new_[8587]_  = ~\new_[8588]_  | (~\new_[8710]_  & ~\new_[2543]_ );
  assign \new_[8588]_  = ~\new_[4173]_  | ~\new_[6160]_ ;
  assign \new_[8589]_  = \new_[8716]_  & \new_[8590]_ ;
  assign \new_[8590]_  = ~\new_[2543]_ ;
  assign \new_[8591]_  = ~\new_[8592]_  | ~\new_[1227]_ ;
  assign \new_[8592]_  = \new_[8972]_  ? \new_[8951]_  : \new_[8971]_ ;
  assign \new_[8593]_  = \new_[8220]_  ? \new_[8222]_  : \new_[8221]_ ;
  assign \new_[8594]_  = ~\new_[8595]_  | ~\new_[8599]_ ;
  assign \new_[8595]_  = ~n1065;
  assign n1065 = ~\new_[8597]_  | ~\new_[8598]_ ;
  assign \new_[8597]_  = ~\new_[1742]_  | ~\new_[2997]_ ;
  assign \new_[8598]_  = ~\new_[3100]_  | ~\new_[1805]_ ;
  assign \new_[8599]_  = ~\new_[8600]_ ;
  assign \new_[8600]_  = ~\new_[3561]_  & ~\new_[2975]_ ;
  assign \new_[8601]_  = ~\new_[8605]_  & (~\new_[8637]_  | ~\new_[8602]_ );
  assign \new_[8602]_  = ~\new_[8603]_  | ~\new_[8604]_ ;
  assign \new_[8603]_  = ~\new_[5754]_  & (~\new_[5880]_  | ~\new_[8779]_ );
  assign \new_[8604]_  = ~\new_[5753]_  & (~\new_[5884]_  | ~\new_[8784]_ );
  assign \new_[8605]_  = ~\new_[8602]_  & ~\new_[8637]_ ;
  assign n995 = \new_[8325]_  ? \new_[8608]_  : \new_[8607]_ ;
  assign \new_[8607]_  = (~\new_[3862]_  | ~\new_[8958]_ ) & (~\new_[8962]_  | ~\new_[6635]_ );
  assign \new_[8608]_  = ~\new_[1811]_  | ~\new_[1851]_ ;
  assign \new_[8609]_  = ~\new_[8610]_  | ~\new_[8614]_ ;
  assign \new_[8610]_  = ~\new_[8611]_ ;
  assign \new_[8611]_  = \new_[8612]_  ? \new_[8651]_  : \new_[8613]_ ;
  assign \new_[8612]_  = ~\new_[8613]_ ;
  assign \new_[8613]_  = \new_[4347]_  ? \new_[8964]_  : \new_[7042]_ ;
  assign \new_[8614]_  = ~\new_[8615]_ ;
  assign \new_[8615]_  = (~\new_[7054]_  | ~\new_[8964]_ ) & (~\new_[4248]_  | ~\new_[8960]_ );
  assign n1610 = \new_[8612]_  ? \new_[8617]_  : \new_[8613]_ ;
  assign \new_[8617]_  = ~\new_[8652]_  | ~\new_[8658]_  | ~\new_[8656]_ ;
  assign \new_[8618]_  = \new_[8619]_  ? \new_[8622]_  : \new_[8620]_ ;
  assign \new_[8619]_  = ~\new_[8532]_  | ~\new_[8530]_  | ~\new_[8529]_ ;
  assign \new_[8620]_  = ~\new_[8621]_ ;
  assign \new_[8621]_  = ~\new_[8532]_  | ~\new_[8530]_  | ~\new_[8529]_ ;
  assign \new_[8622]_  = ~\new_[8521]_  | ~\new_[8519]_  | ~\new_[8623]_ ;
  assign \new_[8623]_  = ~\new_[6073]_  | ~\new_[8779]_ ;
  assign \new_[8624]_  = ~\new_[8625]_  & ~\new_[8725]_ ;
  assign \new_[8625]_  = \new_[8585]_  ? \new_[8628]_  : \new_[8626]_ ;
  assign \new_[8626]_  = ~\new_[8627]_ ;
  assign \new_[8627]_  = \new_[8207]_  ? \new_[8208]_  : \new_[8554]_ ;
  assign \new_[8628]_  = ~\new_[8556]_  | ~\new_[8659]_ ;
  assign \new_[8629]_  = ~\new_[8556]_  | ~\new_[8659]_ ;
  assign n820 = ~\new_[8635]_  | (~\new_[8631]_  & ~\new_[8633]_ );
  assign \new_[8631]_  = \new_[1289]_  ^ \new_[8632]_ ;
  assign \new_[8632]_  = ~\new_[1453]_ ;
  assign \new_[8633]_  = \new_[8634]_  ? \new_[1181]_  : \new_[1377]_ ;
  assign \new_[8634]_  = ~\new_[1377]_ ;
  assign \new_[8635]_  = ~\new_[8633]_  | ~\new_[8631]_ ;
  assign \new_[8636]_  = ~\new_[8641]_  & (~\new_[8637]_  | ~\new_[8753]_ );
  assign \new_[8637]_  = ~\new_[5558]_  | ~\new_[5598]_ ;
  assign \new_[8638]_  = ~\new_[5751]_  & ~\new_[5749]_ ;
  assign \new_[8639]_  = ~\new_[5783]_  | ~\new_[8779]_ ;
  assign \new_[8640]_  = ~\new_[5781]_  | ~\new_[7822]_ ;
  assign \new_[8641]_  = ~\new_[8753]_  & ~\new_[8637]_ ;
  assign \new_[8642]_  = ~\new_[8643]_  | ~\new_[8648]_ ;
  assign \new_[8643]_  = ~\new_[8644]_  | ~\new_[8646]_ ;
  assign \new_[8644]_  = ~\new_[8645]_  | ~\new_[1420]_ ;
  assign \new_[8645]_  = ~\new_[1595]_  | ~\new_[8516]_ ;
  assign \new_[8646]_  = ~\new_[8647]_ ;
  assign \new_[8647]_  = ~\new_[8514]_  & ~n1670;
  assign \new_[8648]_  = ~\new_[8647]_  | ~\new_[8645]_  | ~\new_[1420]_ ;
  assign n800 = ~\new_[8836]_  | ~\new_[8650]_ ;
  assign \new_[8650]_  = ~\new_[7486]_  | ~\new_[1065]_ ;
  assign \new_[8651]_  = ~\new_[8658]_  | ~\new_[8652]_  | ~\new_[8656]_ ;
  assign \new_[8652]_  = ~\new_[8724]_  | ~\new_[8653]_  | ~\new_[8654]_ ;
  assign \new_[8653]_  = ~\new_[8578]_  | ~\new_[1983]_ ;
  assign \new_[8654]_  = ~\new_[8655]_ ;
  assign \new_[8655]_  = \new_[8855]_  ? \new_[8974]_  : \new_[8206]_ ;
  assign \new_[8656]_  = ~\new_[8657]_  | ~\new_[8578]_  | ~\new_[1983]_ ;
  assign \new_[8657]_  = \new_[8655]_  & \new_[8373]_ ;
  assign \new_[8658]_  = \new_[8373]_  | \new_[8585]_ ;
  assign \new_[8659]_  = ~\new_[8885]_  | ~\new_[8660]_ ;
  assign \new_[8660]_  = ~\new_[8661]_ ;
  assign \new_[8661]_  = \new_[8457]_  ? \new_[8458]_  : \new_[5380]_ ;
  assign \new_[8662]_  = \new_[8948]_  ^ \new_[8663]_ ;
  assign \new_[8663]_  = ~\new_[8664]_ ;
  assign \new_[8664]_  = \new_[1068]_  & \new_[1069]_ ;
  assign \new_[8665]_  = ~\new_[8564]_  | ~\new_[8565]_ ;
  assign \new_[8666]_  = ~\new_[8669]_  | ~\new_[8667]_  | ~\new_[8668]_ ;
  assign \new_[8667]_  = ~\new_[6196]_  & ~\new_[6107]_ ;
  assign \new_[8668]_  = ~\new_[6399]_  | ~\new_[8558]_ ;
  assign \new_[8669]_  = ~\new_[6223]_  | ~\new_[8780]_ ;
  assign \new_[8670]_  = ~\new_[8666]_  & ~\new_[8665]_ ;
  assign \new_[8671]_  = (~\new_[8672]_  | ~\new_[8534]_ ) & (~\new_[8673]_  | ~\new_[8674]_ );
  assign \new_[8672]_  = ~\new_[1970]_  | ~\new_[1984]_ ;
  assign \new_[8673]_  = ~\new_[8672]_ ;
  assign \new_[8674]_  = \new_[8675]_  ^ \new_[8676]_ ;
  assign \new_[8675]_  = ~\new_[8537]_  | ~\new_[2665]_ ;
  assign \new_[8676]_  = ~\new_[8677]_ ;
  assign \new_[8677]_  = ~\new_[8539]_  | ~\new_[8678]_ ;
  assign \new_[8678]_  = ~\new_[8433]_ ;
  assign \new_[8679]_  = \new_[8534]_  & \new_[8672]_ ;
  assign \new_[8680]_  = ~\new_[8675]_ ;
  assign \new_[8681]_  = ~\new_[8686]_  & (~\new_[8682]_  | ~\new_[8683]_ );
  assign \new_[8682]_  = ~\new_[5800]_  | ~\new_[5789]_ ;
  assign \new_[8683]_  = ~\new_[8684]_  | ~\new_[8685]_ ;
  assign \new_[8684]_  = ~\new_[8557]_  | ~\new_[8558]_ ;
  assign \new_[8685]_  = ~\new_[8559]_  & (~\new_[6113]_  | ~\new_[8779]_ );
  assign \new_[8686]_  = ~\new_[8683]_  & ~\new_[8682]_ ;
  assign \new_[8687]_  = ~\new_[8688]_  | ~\new_[8689]_ ;
  assign \new_[8688]_  = ~\new_[1068]_ ;
  assign \new_[8689]_  = ~\new_[1066]_ ;
  assign \new_[8690]_  = ~\new_[1068]_  | ~\new_[1066]_ ;
  assign \new_[8691]_  = ~\new_[8697]_  & (~\new_[8692]_  | ~\new_[8693]_ );
  assign \new_[8692]_  = ~\new_[5617]_  | ~\new_[5657]_ ;
  assign \new_[8693]_  = ~\new_[8696]_  | ~\new_[8694]_  | ~\new_[8695]_ ;
  assign \new_[8694]_  = ~\new_[5827]_  & (~\new_[5830]_  | ~\new_[8784]_ );
  assign \new_[8695]_  = ~\new_[5889]_  | ~\new_[7822]_ ;
  assign \new_[8696]_  = ~\new_[5888]_  | ~\new_[8779]_ ;
  assign \new_[8697]_  = ~\new_[8693]_  & ~\new_[8692]_ ;
  assign \new_[8698]_  = ~\new_[1069]_  | ~\new_[1066]_ ;
  assign \new_[8699]_  = ~\new_[1069]_ ;
  assign \new_[8700]_  = ~\new_[1948]_  | ~\new_[8432]_ ;
  assign \new_[8701]_  = ~\new_[1937]_  | ~\new_[1944]_ ;
  assign \new_[8702]_  = \new_[8703]_  ^ \new_[8704]_ ;
  assign \new_[8703]_  = ~\new_[1941]_  | ~\new_[1848]_ ;
  assign \new_[8704]_  = ~\new_[8705]_  | ~\new_[8707]_ ;
  assign \new_[8705]_  = \new_[8706]_ ;
  assign \new_[8706]_  = ~\new_[8701]_  | ~\new_[8700]_ ;
  assign \new_[8707]_  = ~\new_[8517]_  & (~\new_[8680]_  | ~\new_[2015]_ );
  assign \new_[8708]_  = ~\new_[8715]_  & (~\new_[8709]_  | ~\new_[8713]_ );
  assign \new_[8709]_  = ~\new_[8712]_  | (~\new_[8710]_  & ~\new_[2356]_ );
  assign \new_[8710]_  = \new_[8711]_ ;
  assign \new_[8711]_  = ~\new_[7123]_  & (~\new_[7138]_  | ~\new_[8121]_ );
  assign \new_[8712]_  = ~\new_[3866]_  | ~\new_[6161]_ ;
  assign \new_[8713]_  = ~\new_[8714]_ ;
  assign \new_[8714]_  = ~\new_[8115]_  | ~\new_[8108]_ ;
  assign \new_[8715]_  = \new_[8716]_  & \new_[8717]_ ;
  assign \new_[8716]_  = ~\new_[8562]_  | ~\new_[7829]_ ;
  assign \new_[8717]_  = ~\new_[2356]_ ;
  assign \new_[8718]_  = ~\new_[8352]_  | ~\new_[8719]_  | ~\new_[8722]_ ;
  assign \new_[8719]_  = ~\new_[8720]_  | ~\new_[8721]_ ;
  assign \new_[8720]_  = ~\new_[3507]_  | ~\new_[4323]_ ;
  assign \new_[8721]_  = ~\new_[2807]_  | ~\new_[2808]_ ;
  assign \new_[8722]_  = ~\new_[2807]_  | ~\new_[8723]_  | ~\new_[2808]_ ;
  assign \new_[8723]_  = ~\new_[8720]_ ;
  assign \new_[8724]_  = ~\new_[4329]_  | ~decrypt_i;
  assign \new_[8725]_  = ~\new_[8724]_ ;
  assign \new_[8726]_  = \new_[8727]_  & \new_[8989]_ ;
  assign \new_[8727]_  = \new_[8728]_ ;
  assign \new_[8728]_  = ~\new_[8882]_  | ~\new_[5488]_ ;
  assign \new_[8729]_  = ~\new_[8730]_  | ~\new_[6771]_ ;
  assign \new_[8730]_  = ~\new_[8731]_  | ~\new_[8732]_ ;
  assign \new_[8731]_  = ~\new_[7876]_  & ~\new_[7869]_ ;
  assign \new_[8732]_  = ~\new_[7896]_  & ~\new_[7868]_ ;
  assign \new_[8733]_  = ~\new_[9014]_ ;
  assign \new_[8734]_  = ~\new_[8687]_  | ~\new_[8690]_ ;
  assign \new_[8735]_  = ~\new_[8690]_  | ~\new_[8687]_  | ~\new_[9015]_ ;
  assign \new_[8736]_  = \new_[8857]_  ? \new_[8738]_  : \new_[8737]_ ;
  assign \new_[8737]_  = ~\new_[8857]_ ;
  assign \new_[8738]_  = \new_[8833]_  ^ \new_[8795]_ ;
  assign \new_[8739]_  = ~\new_[8745]_  & (~\new_[8740]_  | ~\new_[8741]_ );
  assign \new_[8740]_  = ~\new_[5618]_  | ~\new_[5656]_ ;
  assign \new_[8741]_  = ~\new_[8744]_  | ~\new_[8742]_  | ~\new_[8743]_ ;
  assign \new_[8742]_  = ~\new_[5886]_  | ~\new_[8779]_ ;
  assign \new_[8743]_  = ~\new_[5776]_  & ~\new_[5772]_ ;
  assign \new_[8744]_  = ~\new_[5887]_  | ~\new_[7822]_ ;
  assign \new_[8745]_  = ~\new_[8741]_  & ~\new_[8740]_ ;
  assign \new_[8746]_  = ~\new_[4243]_  | ~\new_[8961]_ ;
  assign \new_[8747]_  = ~\new_[8964]_  | ~\new_[6773]_ ;
  assign \new_[8748]_  = \new_[8818]_  ? \new_[8822]_  : \new_[8821]_ ;
  assign \new_[8749]_  = \new_[8978]_  ? \new_[8829]_  : \new_[8977]_ ;
  assign \new_[8750]_  = \new_[8225]_  ? \new_[8227]_  : \new_[8226]_ ;
  assign \new_[8751]_  = \new_[8753]_  ? \new_[8754]_  : \new_[8752]_ ;
  assign \new_[8752]_  = ~\new_[8753]_ ;
  assign \new_[8753]_  = ~\new_[8640]_  | ~\new_[8639]_  | ~\new_[8638]_ ;
  assign \new_[8754]_  = ~\new_[8755]_  | ~\new_[8757]_ ;
  assign \new_[8755]_  = ~\new_[8756]_  & (~\new_[5780]_  | ~\new_[7822]_ );
  assign \new_[8756]_  = \new_[5750]_  | \new_[5752]_ ;
  assign \new_[8757]_  = ~\new_[5778]_  | ~\new_[8779]_ ;
  assign \new_[8758]_  = ~\new_[8764]_  & (~\new_[8759]_  | ~\new_[8762]_ );
  assign \new_[8759]_  = \new_[8794]_  ? \new_[8761]_  : \new_[8760]_ ;
  assign \new_[8760]_  = ~\new_[8794]_ ;
  assign \new_[8761]_  = ~\new_[5799]_  | ~\new_[5790]_ ;
  assign \new_[8762]_  = \new_[8763]_ ;
  assign \new_[8763]_  = ~\new_[8670]_  & (~\new_[8665]_  | ~\new_[8666]_ );
  assign \new_[8764]_  = ~\new_[8762]_  & ~\new_[8759]_ ;
  assign \new_[8765]_  = ~\new_[8766]_  | ~\new_[8767]_ ;
  assign \new_[8766]_  = ~\new_[8335]_  | ~\new_[8177]_ ;
  assign \new_[8767]_  = ~\new_[8768]_ ;
  assign \new_[8768]_  = \new_[8769]_  & \new_[8770]_ ;
  assign \new_[8769]_  = ~\new_[4445]_  | ~\new_[8960]_ ;
  assign \new_[8770]_  = ~\new_[8964]_  | ~\new_[7092]_ ;
  assign \new_[8771]_  = ~\new_[8768]_  | ~\new_[8335]_  | ~\new_[8177]_ ;
  assign \new_[8772]_  = ~\new_[8773]_  | ~\new_[8775]_ ;
  assign \new_[8773]_  = ~\new_[8774]_  | ~\new_[7893]_ ;
  assign \new_[8774]_  = ~\new_[6045]_  | ~\new_[6049]_ ;
  assign \new_[8775]_  = ~\new_[8776]_  & (~\new_[5974]_  | ~\new_[7822]_ );
  assign \new_[8776]_  = ~\new_[8777]_  | ~\new_[8782]_ ;
  assign \new_[8777]_  = ~\new_[8778]_  | ~\new_[8779]_ ;
  assign \new_[8778]_  = \data_o[116]  ? \new_[8912]_  : \new_[1204]_ ;
  assign \new_[8779]_  = ~\new_[8781]_ ;
  assign \new_[8780]_  = ~\new_[8781]_ ;
  assign \new_[8781]_  = ~\new_[8711]_  | ~\new_[8713]_ ;
  assign \new_[8782]_  = ~\new_[8783]_  | ~\new_[8784]_ ;
  assign \new_[8783]_  = \data_o[20]  ? \new_[8912]_  : \new_[1206]_ ;
  assign \new_[8784]_  = \new_[5612]_  & \new_[5659]_ ;
  assign \new_[8785]_  = ~\new_[8789]_  | (~\new_[8786]_  & ~\new_[8788]_ );
  assign \new_[8786]_  = ~\new_[8787]_  | ~\new_[8880]_ ;
  assign \new_[8787]_  = ~\new_[5253]_  | ~\key_i[16] ;
  assign \new_[8788]_  = ~\new_[5201]_  & (~\new_[6540]_  | ~\new_[6812]_ );
  assign \new_[8789]_  = \new_[8880]_  | \new_[8256]_ ;
  assign \new_[8790]_  = \new_[8791]_  ? \new_[8793]_  : \new_[8792]_ ;
  assign \new_[8791]_  = \new_[8665]_  ^ \new_[8863]_ ;
  assign \new_[8792]_  = ~\new_[8791]_ ;
  assign \new_[8793]_  = ~\new_[8796]_  & (~\new_[8794]_  | ~\new_[8795]_ );
  assign \new_[8794]_  = ~\new_[5798]_  | ~\new_[5791]_ ;
  assign \new_[8795]_  = ~\new_[5801]_  | ~\new_[5787]_ ;
  assign \new_[8796]_  = ~\new_[8795]_  & ~\new_[8794]_ ;
  assign \new_[8797]_  = \new_[8791]_ ;
  assign \new_[8798]_  = \new_[8799]_  ^ \new_[8800]_ ;
  assign \new_[8799]_  = ~\new_[1067]_ ;
  assign \new_[8800]_  = \new_[8801]_ ;
  assign \new_[8801]_  = ~\new_[1068]_  | ~\new_[1066]_ ;
  assign \new_[8802]_  = ~\new_[8800]_ ;
  assign \new_[8803]_  = ~\new_[8806]_  | (~\new_[8804]_  & ~\new_[9001]_ );
  assign \new_[8804]_  = ~\new_[4945]_  & (~\new_[6501]_  | ~\new_[5115]_ );
  assign \new_[8805]_  = ~\new_[8881]_  | ~\new_[5488]_ ;
  assign \new_[8806]_  = \new_[7650]_  | \new_[9002]_ ;
  assign \new_[8807]_  = ~\new_[8882]_ ;
  assign \new_[8808]_  = ~\new_[8814]_  & (~\new_[8953]_  | ~\new_[8950]_ );
  assign \new_[8809]_  = \new_[8293]_  ? \new_[8296]_  : \new_[8294]_ ;
  assign \new_[8810]_  = \new_[8811]_  ? \new_[8813]_  : \new_[8812]_ ;
  assign \new_[8811]_  = (~\new_[7814]_  & ~\new_[7863]_ ) | (~\new_[7834]_  & ~\new_[7858]_ );
  assign \new_[8812]_  = ~\new_[8811]_ ;
  assign \new_[8813]_  = ~\new_[8223]_  | ~\new_[8224]_ ;
  assign \new_[8814]_  = ~\new_[8953]_  & ~\new_[8950]_ ;
  assign \new_[8815]_  = ~\new_[8816]_  | ~\new_[8820]_ ;
  assign \new_[8816]_  = ~\new_[8819]_  & (~\new_[8817]_  | ~\new_[8765]_ );
  assign \new_[8817]_  = \new_[8771]_  & \new_[8818]_ ;
  assign \new_[8818]_  = ~\new_[8746]_  | ~\new_[8747]_ ;
  assign \new_[8819]_  = ~\new_[2972]_  & (~\new_[3983]_  | ~\new_[6136]_ );
  assign \new_[8820]_  = ~\new_[8821]_  | ~\new_[8822]_ ;
  assign \new_[8821]_  = ~\new_[8818]_ ;
  assign \new_[8822]_  = ~\new_[8765]_  | ~\new_[8771]_ ;
  assign \new_[8823]_  = \new_[8821]_  ^ \new_[9004]_ ;
  assign \new_[8824]_  = ~\new_[8825]_  | ~\new_[8828]_ ;
  assign \new_[8825]_  = ~\new_[8891]_ ;
  assign \new_[8826]_  = (~\new_[5842]_  & ~\new_[5917]_ ) | (~\new_[5910]_  & ~\new_[5854]_ );
  assign \new_[8827]_  = \new_[5555]_  ? \new_[8413]_  : \new_[5489]_ ;
  assign \new_[8828]_  = \new_[4827]_  ? \new_[8750]_  : \new_[8661]_ ;
  assign \new_[8829]_  = \new_[8890]_  ? \new_[8830]_  : \new_[8826]_ ;
  assign \new_[8830]_  = \new_[5555]_  ? \new_[8413]_  : \new_[5489]_ ;
  assign \new_[8831]_  = ~\new_[8834]_  & (~\new_[8832]_  | ~\new_[8833]_ );
  assign \new_[8832]_  = ~\new_[5790]_  | ~\new_[5799]_ ;
  assign \new_[8833]_  = ~\new_[5788]_  | ~\new_[5803]_ ;
  assign \new_[8834]_  = ~\new_[8835]_  & ~\new_[8832]_ ;
  assign \new_[8835]_  = ~\new_[5788]_  | ~\new_[5803]_ ;
  assign \new_[8836]_  = ~\new_[8843]_  | ~\new_[8837]_  | ~\new_[8841]_ ;
  assign \new_[8837]_  = ~n860 | ~\new_[8839]_ ;
  assign n860 = ~\new_[1299]_  | ~\new_[8594]_ ;
  assign \new_[8839]_  = \new_[8840]_ ;
  assign \new_[8840]_  = ~\new_[5075]_  | (~\new_[4790]_  & ~\new_[8967]_ );
  assign \new_[8841]_  = ~\new_[8594]_  | ~\new_[8842]_  | ~\new_[1299]_ ;
  assign \new_[8842]_  = ~\new_[8839]_ ;
  assign \new_[8843]_  = \new_[8853]_ ;
  assign \new_[8844]_  = ~\new_[8852]_  | ~\new_[8845]_  | ~\new_[8849]_ ;
  assign \new_[8845]_  = ~n865 | ~\new_[8847]_ ;
  assign n865 = ~\new_[1358]_  | ~\new_[1300]_ ;
  assign \new_[8847]_  = ~\new_[8848]_  | (~\new_[4786]_  & ~\new_[8964]_ );
  assign \new_[8848]_  = \new_[7561]_  | \new_[8966]_ ;
  assign \new_[8849]_  = ~\new_[8850]_  | ~\new_[1300]_ ;
  assign \new_[8850]_  = \new_[1358]_  & \new_[8851]_ ;
  assign \new_[8851]_  = ~\new_[8847]_ ;
  assign \new_[8852]_  = \new_[8853]_ ;
  assign \new_[8853]_  = ~\new_[7536]_  & ~\new_[8204]_ ;
  assign \new_[8854]_  = \new_[8877]_  ? \new_[8855]_  : \new_[8216]_ ;
  assign \new_[8855]_  = \new_[8885]_ ;
  assign \new_[8856]_  = ~\new_[8855]_ ;
  assign \new_[8857]_  = \new_[8858]_  ? \new_[8863]_  : \new_[8862]_ ;
  assign \new_[8858]_  = ~\new_[8861]_  | ~\new_[8859]_  | ~\new_[8860]_ ;
  assign \new_[8859]_  = ~\new_[6218]_  | ~\new_[8784]_ ;
  assign \new_[8860]_  = ~\new_[6404]_  | ~\new_[8780]_ ;
  assign \new_[8861]_  = ~\new_[6392]_  & (~\new_[6551]_  | ~\new_[8558]_ );
  assign \new_[8862]_  = ~\new_[8858]_ ;
  assign \new_[8863]_  = ~\new_[8451]_  | ~\new_[8452]_ ;
  assign \new_[8864]_  = \new_[8865]_  ^ \new_[8869]_ ;
  assign \new_[8865]_  = ~\new_[8868]_  | ~\new_[8866]_  | ~\new_[8867]_ ;
  assign \new_[8866]_  = ~\new_[6207]_  | ~\new_[8780]_ ;
  assign \new_[8867]_  = ~\new_[6108]_  & ~\new_[6103]_ ;
  assign \new_[8868]_  = ~\new_[6398]_  | ~\new_[8784]_ ;
  assign \new_[8869]_  = ~\new_[5919]_  | ~\new_[5903]_ ;
  assign \new_[8870]_  = \new_[8871]_  ^ \new_[8875]_ ;
  assign \new_[8871]_  = ~\new_[8874]_  | ~\new_[8872]_  | ~\new_[8873]_ ;
  assign \new_[8872]_  = ~\new_[6148]_  | ~\new_[8558]_ ;
  assign \new_[8873]_  = ~\new_[6208]_  | ~\new_[8780]_ ;
  assign \new_[8874]_  = ~\new_[6034]_  & ~\new_[6109]_ ;
  assign \new_[8875]_  = ~\new_[6032]_  | ~\new_[5904]_ ;
  assign \new_[8876]_  = \new_[8216]_  ? \new_[9003]_  : \new_[8877]_ ;
  assign \new_[8877]_  = \new_[4542]_  ? \new_[8363]_  : \new_[4464]_ ;
  assign \new_[8878]_  = ~\new_[8879]_  | ~\new_[8883]_ ;
  assign \new_[8879]_  = ~\new_[8966]_  | ~\new_[4942]_  | ~\new_[4941]_ ;
  assign \new_[8880]_  = ~\new_[8881]_  | ~\new_[5488]_ ;
  assign \new_[8881]_  = ~\new_[8882]_ ;
  assign \new_[8882]_  = ~\new_[7903]_  | ~\new_[9019]_ ;
  assign \new_[8883]_  = ~\new_[8884]_  | ~\new_[8967]_ ;
  assign \new_[8884]_  = \new_[7989]_  ? \new_[7875]_  : \new_[8018]_ ;
  assign \new_[8885]_  = \new_[8886]_  ^ \new_[8888]_ ;
  assign \new_[8886]_  = (~\new_[5241]_  & ~\new_[5620]_ ) | (~\new_[8887]_  & ~\new_[5671]_ );
  assign \new_[8887]_  = ~\new_[5241]_ ;
  assign \new_[8888]_  = ~\new_[8889]_ ;
  assign \new_[8889]_  = \new_[8826]_  ? \new_[8827]_  : \new_[8890]_ ;
  assign \new_[8890]_  = ~\new_[8826]_ ;
  assign \new_[8891]_  = \new_[8826]_  ? \new_[8827]_  : \new_[8890]_ ;
  assign \new_[8892]_  = ~\new_[8886]_ ;
  assign \new_[8893]_  = ~\new_[8905]_ ;
  assign \new_[8894]_  = ~\new_[8895]_ ;
  assign \new_[8895]_  = ~\new_[8906]_ ;
  assign \new_[8896]_  = ~\new_[8897]_ ;
  assign \new_[8897]_  = ~\new_[8900]_ ;
  assign \new_[8898]_  = ~\new_[8899]_ ;
  assign \new_[8899]_  = \new_[8900]_ ;
  assign \new_[8900]_  = ~\new_[8901]_ ;
  assign \new_[8901]_  = ~\new_[8902]_ ;
  assign \new_[8902]_  = ~\new_[8903]_ ;
  assign \new_[8903]_  = ~\new_[8906]_ ;
  assign \new_[8904]_  = ~\new_[8905]_ ;
  assign \new_[8905]_  = ~\new_[8906]_ ;
  assign \new_[8906]_  = ~\new_[8236]_ ;
  assign \new_[8907]_  = ~\new_[8912]_ ;
  assign \new_[8908]_  = \new_[8911]_ ;
  assign \new_[8909]_  = ~\new_[8911]_ ;
  assign \new_[8910]_  = ~\new_[8911]_ ;
  assign \new_[8911]_  = ~\new_[8912]_ ;
  assign \new_[8912]_  = \new_[8915]_ ;
  assign \new_[8913]_  = ~\new_[8914]_ ;
  assign \new_[8914]_  = ~\new_[8915]_ ;
  assign \new_[8915]_  = \new_[8920]_ ;
  assign \new_[8916]_  = ~\new_[8917]_ ;
  assign \new_[8917]_  = ~\new_[8918]_ ;
  assign \new_[8918]_  = ~\new_[8919]_ ;
  assign \new_[8919]_  = ~\new_[8920]_ ;
  assign \new_[8920]_  = ~\new_[8937]_ ;
  assign \new_[8921]_  = \new_[8920]_ ;
  assign \new_[8922]_  = ~\new_[8924]_ ;
  assign \new_[8923]_  = ~\new_[8922]_ ;
  assign \new_[8924]_  = ~\new_[8925]_ ;
  assign \new_[8925]_  = ~\new_[8927]_ ;
  assign \new_[8926]_  = \new_[8927]_ ;
  assign \new_[8927]_  = ~\new_[8936]_ ;
  assign \new_[8928]_  = ~\new_[8929]_ ;
  assign \new_[8929]_  = \new_[8933]_ ;
  assign \new_[8930]_  = ~\new_[8932]_ ;
  assign \new_[8931]_  = ~\new_[8933]_ ;
  assign \new_[8932]_  = \new_[8933]_ ;
  assign \new_[8933]_  = ~\new_[8934]_ ;
  assign \new_[8934]_  = \new_[8935]_ ;
  assign \new_[8935]_  = ~\new_[8936]_ ;
  assign \new_[8936]_  = ~\new_[8920]_ ;
  assign \new_[8937]_  = \new_[8236]_ ;
  assign \new_[8938]_  = ~\new_[8939]_ ;
  assign \new_[8939]_  = ~\new_[8940]_ ;
  assign \new_[8940]_  = ~\new_[8947]_ ;
  assign \new_[8941]_  = ~\new_[8942]_ ;
  assign \new_[8942]_  = \new_[8947]_ ;
  assign \new_[8943]_  = ~\new_[8947]_ ;
  assign \new_[8944]_  = ~\new_[8947]_ ;
  assign \new_[8945]_  = ~\new_[8946]_ ;
  assign \new_[8946]_  = ~\new_[8947]_ ;
  assign \new_[8947]_  = \new_[8236]_ ;
  assign \new_[8948]_  = ~\new_[8949]_ ;
  assign \new_[8949]_  = ~\new_[8698]_ ;
  assign \new_[8950]_  = ~\new_[8951]_ ;
  assign \new_[8951]_  = ~\new_[8810]_ ;
  assign \new_[8952]_  = \new_[8953]_ ;
  assign \new_[8953]_  = \new_[8809]_ ;
  assign \new_[8954]_  = ~\new_[8961]_ ;
  assign \new_[8955]_  = ~\new_[8959]_ ;
  assign \new_[8956]_  = ~\new_[8959]_ ;
  assign \new_[8957]_  = \new_[8958]_ ;
  assign \new_[8958]_  = ~\new_[8959]_ ;
  assign \new_[8959]_  = ~\new_[8960]_ ;
  assign \new_[8960]_  = ~\new_[8963]_ ;
  assign \new_[8961]_  = ~\new_[8964]_ ;
  assign \new_[8962]_  = ~\new_[8961]_ ;
  assign \new_[8963]_  = \new_[8964]_ ;
  assign \new_[8964]_  = ~\new_[8965]_ ;
  assign \new_[8965]_  = ~\new_[8967]_ ;
  assign \new_[8966]_  = ~\new_[8967]_ ;
  assign \new_[8967]_  = ~\new_[8880]_ ;
  assign \new_[8968]_  = \new_[8392]_ ;
  assign \new_[8969]_  = ~\new_[8972]_ ;
  assign \new_[8970]_  = \new_[8971]_ ;
  assign \new_[8971]_  = ~\new_[8972]_ ;
  assign \new_[8972]_  = ~\new_[8593]_ ;
  assign \new_[8973]_  = \new_[8411]_  ? \new_[8412]_  : \new_[4729]_ ;
  assign \new_[8974]_  = \new_[8411]_  ? \new_[8412]_  : \new_[4729]_ ;
  assign \new_[8975]_  = ~\new_[1387]_  | ~\new_[8593]_ ;
  assign \new_[8976]_  = ~\new_[1387]_  | ~\new_[8593]_ ;
  assign \new_[8977]_  = ~\new_[8978]_ ;
  assign \new_[8978]_  = \new_[8750]_ ;
  assign \new_[8979]_  = ~\new_[8983]_ ;
  assign n1600 = \new_[8981]_ ;
  assign \new_[8981]_  = ~\new_[8982]_ ;
  assign \new_[8982]_  = ~\new_[8979]_ ;
  assign \new_[8983]_  = ~\new_[8671]_ ;
  assign \new_[8984]_  = ~\new_[8985]_ ;
  assign \new_[8985]_  = \new_[8986]_ ;
  assign \new_[8986]_  = ~\new_[8217]_ ;
  assign \new_[8987]_  = ~\new_[8988]_ ;
  assign \new_[8988]_  = \new_[8999]_ ;
  assign \new_[8989]_  = ~\new_[8990]_ ;
  assign \new_[8990]_  = \new_[8998]_ ;
  assign \new_[8991]_  = ~\new_[8993]_ ;
  assign \new_[8992]_  = ~\new_[8993]_ ;
  assign \new_[8993]_  = \new_[8995]_ ;
  assign \new_[8994]_  = ~\new_[8995]_ ;
  assign \new_[8995]_  = \new_[8998]_ ;
  assign \new_[8996]_  = ~\new_[8997]_ ;
  assign \new_[8997]_  = ~\new_[8998]_ ;
  assign \new_[8998]_  = ~\new_[8999]_ ;
  assign \new_[8999]_  = ~\new_[8729]_ ;
  assign \new_[9000]_  = ~\new_[9001]_ ;
  assign \new_[9001]_  = ~\new_[9002]_ ;
  assign \new_[9002]_  = \new_[8805]_ ;
  assign \new_[9003]_  = \new_[8973]_ ;
  assign \new_[9004]_  = \new_[8822]_ ;
  assign \new_[9005]_  = \new_[9006]_ ;
  assign \new_[9006]_  = \new_[8569]_ ;
  assign \new_[9007]_  = ~\new_[9008]_ ;
  assign \new_[9008]_  = ~\new_[9010]_  | ~\new_[8735]_ ;
  assign \new_[9009]_  = ~\new_[9011]_  | ~\new_[8735]_ ;
  assign \new_[9010]_  = ~\new_[8734]_  | ~\new_[8733]_ ;
  assign \new_[9011]_  = ~\new_[8734]_  | ~\new_[8733]_ ;
  assign n1615 = \new_[8402]_  ? \new_[8404]_  : \new_[8403]_ ;
  assign \new_[9013]_  = \new_[8402]_  ? \new_[8404]_  : \new_[8403]_ ;
  assign \new_[9014]_  = ~\new_[8801]_  | ~\new_[1067]_ ;
  assign \new_[9015]_  = ~\new_[8801]_  | ~\new_[1067]_ ;
  assign \new_[9016]_  = ~\new_[8304]_  & (~\new_[9001]_  | ~\new_[8303]_ );
  assign \new_[9017]_  = ~\new_[8304]_  & (~\new_[9001]_  | ~\new_[8303]_ );
  assign \new_[9018]_  = \new_[7890]_  & \new_[8046]_ ;
  assign \new_[9019]_  = \new_[7890]_  & \new_[8046]_ ;
  always @ (posedge clock) begin
    \\ks1_key_reg_reg[11]  <= n780;
    \\ks1_key_reg_reg[12]  <= n785;
    \\ks1_key_reg_reg[13]  <= n790;
    \\ks1_key_reg_reg[14]  <= n795;
    \\ks1_key_reg_reg[15]  <= n800;
    \\sbox1_to_invert_reg[1]  <= n805;
    \\sbox1_to_invert_reg[3]  <= n810;
    \\sbox1_to_invert_reg[2]  <= n815;
    \\sbox1_to_invert_reg[0]  <= n820;
    \\ks1_key_reg_reg[8]  <= n825;
    \\ks1_key_reg_reg[10]  <= n830;
    \\ks1_key_reg_reg[9]  <= n835;
    \\ks1_key_reg_reg[43]  <= n840;
    \\ks1_key_reg_reg[44]  <= n845;
    \\ks1_key_reg_reg[45]  <= n850;
    \\ks1_key_reg_reg[46]  <= n855;
    \\ks1_key_reg_reg[47]  <= n860;
    \\ks1_key_reg_reg[40]  <= n865;
    \\sub1_data_reg_reg[109]  <= n870;
    \\sub1_data_reg_reg[110]  <= n875;
    \\sub1_data_reg_reg[13]  <= n880;
    \\sub1_data_reg_reg[14]  <= n885;
    \\sub1_data_reg_reg[45]  <= n890;
    \\sub1_data_reg_reg[46]  <= n895;
    \\sub1_data_reg_reg[77]  <= n900;
    \\sub1_data_reg_reg[78]  <= n905;
    \\sub1_data_reg_reg[102]  <= n910;
    \\sub1_data_reg_reg[101]  <= n915;
    \\sub1_data_reg_reg[118]  <= n920;
    \\sub1_data_reg_reg[117]  <= n925;
    \\sub1_data_reg_reg[21]  <= n930;
    \\sub1_data_reg_reg[22]  <= n935;
    \\sub1_data_reg_reg[37]  <= n940;
    \\sub1_data_reg_reg[38]  <= n945;
    \\sub1_data_reg_reg[53]  <= n950;
    \\sub1_data_reg_reg[54]  <= n955;
    \\sub1_data_reg_reg[5]  <= n960;
    \\sub1_data_reg_reg[6]  <= n965;
    \\sub1_data_reg_reg[70]  <= n970;
    \\sub1_data_reg_reg[69]  <= n975;
    \\sub1_data_reg_reg[85]  <= n980;
    \\sub1_data_reg_reg[86]  <= n985;
    \\ks1_key_reg_reg[42]  <= n990;
    \\ks1_key_reg_reg[41]  <= n995;
    \\ks1_key_reg_reg[76]  <= n1000;
    \\ks1_key_reg_reg[75]  <= n1005;
    \\ks1_key_reg_reg[74]  <= n1010;
    \\ks1_key_reg_reg[73]  <= n1015;
    \\ks1_key_reg_reg[77]  <= n1020;
    \\ks1_key_reg_reg[78]  <= n1025;
    \\sub1_data_reg_reg[125]  <= n1030;
    \\sub1_data_reg_reg[126]  <= n1035;
    \\sub1_data_reg_reg[29]  <= n1040;
    \\sub1_data_reg_reg[94]  <= n1045;
    \\sub1_data_reg_reg[30]  <= n1050;
    \\sub1_data_reg_reg[93]  <= n1055;
    \\ks1_key_reg_reg[72]  <= n1060;
    \\ks1_key_reg_reg[79]  <= n1065;
    \\sub1_data_reg_reg[104]  <= n1070;
    \\sub1_data_reg_reg[40]  <= n1075;
    \\sub1_data_reg_reg[72]  <= n1080;
    \\sub1_data_reg_reg[8]  <= n1085;
    \\sub1_data_reg_reg[0]  <= n1090;
    \\sub1_data_reg_reg[112]  <= n1095;
    \\sub1_data_reg_reg[16]  <= n1100;
    \\sub1_data_reg_reg[64]  <= n1105;
    \\sub1_data_reg_reg[80]  <= n1110;
    \\sub1_data_reg_reg[96]  <= n1115;
    \\sub1_data_reg_reg[48]  <= n1120;
    \\sub1_data_reg_reg[61]  <= n1125;
    \\sub1_data_reg_reg[62]  <= n1130;
    \\ks1_col_reg[21]  <= n1135;
    \\ks1_col_reg[22]  <= n1140;
    \\sub1_data_reg_reg[107]  <= n1145;
    \\sub1_data_reg_reg[108]  <= n1150;
    \\sub1_data_reg_reg[111]  <= n1155;
    \\sub1_data_reg_reg[11]  <= n1160;
    \\sub1_data_reg_reg[12]  <= n1165;
    \\sub1_data_reg_reg[15]  <= n1170;
    \\sub1_data_reg_reg[44]  <= n1175;
    \\sub1_data_reg_reg[43]  <= n1180;
    \\sub1_data_reg_reg[47]  <= n1185;
    \\sub1_data_reg_reg[75]  <= n1190;
    \\sub1_data_reg_reg[76]  <= n1195;
    \\sub1_data_reg_reg[79]  <= n1200;
    \\sub1_data_reg_reg[103]  <= n1205;
    \\sub1_data_reg_reg[115]  <= n1210;
    \\sub1_data_reg_reg[116]  <= n1215;
    \\sub1_data_reg_reg[119]  <= n1220;
    \\sub1_data_reg_reg[20]  <= n1225;
    \\sub1_data_reg_reg[19]  <= n1230;
    \\sub1_data_reg_reg[23]  <= n1235;
    \\sub1_data_reg_reg[32]  <= n1240;
    \\sub1_data_reg_reg[4]  <= n1245;
    \\sub1_data_reg_reg[51]  <= n1250;
    \\sub1_data_reg_reg[52]  <= n1255;
    \\sub1_data_reg_reg[55]  <= n1260;
    \\sub1_data_reg_reg[36]  <= n1265;
    \\sub1_data_reg_reg[68]  <= n1270;
    \\sub1_data_reg_reg[67]  <= n1275;
    \\sub1_data_reg_reg[3]  <= n1280;
    \\sub1_data_reg_reg[7]  <= n1285;
    \\sub1_data_reg_reg[71]  <= n1290;
    \\sub1_data_reg_reg[84]  <= n1295;
    \\sub1_data_reg_reg[83]  <= n1300;
    \\sub1_data_reg_reg[87]  <= n1305;
    \\sub1_data_reg_reg[120]  <= n1310;
    \\sub1_data_reg_reg[24]  <= n1315;
    \\sub1_data_reg_reg[56]  <= n1320;
    \\sub1_data_reg_reg[88]  <= n1325;
    \\sbox1_alph_reg[2]  <= n1330;
    \\ks1_col_reg[30]  <= n1335;
    \\sub1_data_reg_reg[100]  <= n1340;
    \\ks1_col_reg[6]  <= n1345;
    \\ks1_col_reg[5]  <= n1350;
    \\sub1_data_reg_reg[35]  <= n1355;
    \\sub1_data_reg_reg[39]  <= n1360;
    \\ks1_col_reg[29]  <= n1365;
    \\sub1_data_reg_reg[99]  <= n1370;
    \\sub1_data_reg_reg[123]  <= n1375;
    \\sub1_data_reg_reg[124]  <= n1380;
    \\sub1_data_reg_reg[127]  <= n1385;
    \\sub1_data_reg_reg[27]  <= n1390;
    \\sub1_data_reg_reg[28]  <= n1395;
    \\sub1_data_reg_reg[31]  <= n1400;
    \\sub1_data_reg_reg[59]  <= n1405;
    \\sub1_data_reg_reg[60]  <= n1410;
    \\sub1_data_reg_reg[63]  <= n1415;
    \\sub1_data_reg_reg[95]  <= n1420;
    \\sub1_data_reg_reg[91]  <= n1425;
    \\sub1_data_reg_reg[92]  <= n1430;
    \\ks1_col_reg[16]  <= n1435;
    \\sbox1_alph_reg[0]  <= n1440;
    \\ks1_key_reg_reg[107]  <= n1445;
    \\ks1_key_reg_reg[108]  <= n1450;
    \\ks1_col_reg[20]  <= n1455;
    \\ks1_key_reg_reg[104]  <= n1460;
    \\ks1_col_reg[23]  <= n1465;
    \\ks1_col_reg[19]  <= n1470;
    \\sub1_data_reg_reg[106]  <= n1475;
    \\sub1_data_reg_reg[10]  <= n1480;
    \\sub1_data_reg_reg[74]  <= n1485;
    \\sub1_data_reg_reg[42]  <= n1490;
    \\sub1_data_reg_reg[114]  <= n1495;
    \\ks1_col_reg[24]  <= n1500;
    \\ks1_col_reg[3]  <= n1505;
    \\ks1_col_reg[4]  <= n1510;
    \\sub1_data_reg_reg[18]  <= n1515;
    \\sub1_data_reg_reg[2]  <= n1520;
    \\sub1_data_reg_reg[50]  <= n1525;
    \\sub1_data_reg_reg[66]  <= n1530;
    \\sub1_data_reg_reg[82]  <= n1535;
    \\sub1_data_reg_reg[98]  <= n1540;
    \\ks1_col_reg[0]  <= n1545;
    \\ks1_col_reg[28]  <= n1550;
    \\ks1_key_reg_reg[111]  <= n1555;
    \\ks1_col_reg[27]  <= n1560;
    \\ks1_col_reg[31]  <= n1565;
    \\sub1_data_reg_reg[34]  <= n1570;
    \\ks1_col_reg[7]  <= n1575;
    \\sub1_data_reg_reg[122]  <= n1580;
    \\sub1_data_reg_reg[26]  <= n1585;
    \\sub1_data_reg_reg[58]  <= n1590;
    \\sub1_data_reg_reg[90]  <= n1595;
    \\sbox1_ah_reg_reg[2]  <= n1600;
    \\sbox1_alph_reg[1]  <= n1605;
    \\ks1_key_reg_reg[110]  <= n1610;
    \\ks1_key_reg_reg[109]  <= n1615;
    \\sub1_data_reg_reg[105]  <= n1620;
    \\sub1_data_reg_reg[41]  <= n1625;
    \\sub1_data_reg_reg[73]  <= n1630;
    \\sub1_data_reg_reg[9]  <= n1635;
    \\sub1_data_reg_reg[17]  <= n1640;
    \\sub1_data_reg_reg[1]  <= n1645;
    \\sub1_data_reg_reg[65]  <= n1650;
    \\sub1_data_reg_reg[97]  <= n1655;
    \\ks1_key_reg_reg[105]  <= n1660;
    \\ks1_col_reg[18]  <= n1665;
    \\sbox1_ah_reg_reg[0]  <= n1670;
    \\sub1_data_reg_reg[81]  <= n1675;
    \\sub1_data_reg_reg[49]  <= n1680;
    \\sub1_data_reg_reg[113]  <= n1685;
    \\sub1_data_reg_reg[33]  <= n1690;
    \\sub1_data_reg_reg[57]  <= n1695;
    \\sub1_data_reg_reg[89]  <= n1700;
    \\sub1_data_reg_reg[25]  <= n1705;
    \\ks1_col_reg[26]  <= n1710;
    \\sub1_data_reg_reg[121]  <= n1715;
    \\ks1_key_reg_reg[106]  <= n1720;
    \\ks1_col_reg[2]  <= n1725;
    \\sbox1_ah_reg_reg[1]  <= n1730;
    \\ks1_col_reg[17]  <= n1735;
    \\sbox1_alph_reg[3]  <= n1740;
    \\ks1_col_reg[25]  <= n1745;
    \\ks1_col_reg[1]  <= n1750;
    \\sbox1_ah_reg_reg[3]  <= n1755;
    \\ks1_key_reg_reg[28]  <= n1760;
    \\ks1_key_reg_reg[27]  <= n1765;
    \\ks1_key_reg_reg[29]  <= n1770;
    \\ks1_key_reg_reg[30]  <= n1775;
    \\ks1_key_reg_reg[24]  <= n1780;
    \\ks1_key_reg_reg[31]  <= n1785;
    \\ks1_key_reg_reg[25]  <= n1790;
    \\ks1_key_reg_reg[26]  <= n1795;
    \\ks1_key_reg_reg[60]  <= n1800;
    \\ks1_key_reg_reg[2]  <= n1805;
    \\ks1_key_reg_reg[3]  <= n1810;
    \\ks1_key_reg_reg[4]  <= n1815;
    \\ks1_key_reg_reg[5]  <= n1820;
    \\ks1_key_reg_reg[6]  <= n1825;
    \\ks1_key_reg_reg[0]  <= n1830;
    \\ks1_key_reg_reg[1]  <= n1835;
    \\ks1_key_reg_reg[23]  <= n1840;
    \\ks1_key_reg_reg[7]  <= n1845;
    \\ks1_key_reg_reg[61]  <= n1850;
    \\ks1_key_reg_reg[59]  <= n1855;
    \\ks1_key_reg_reg[17]  <= n1860;
    \\ks1_key_reg_reg[16]  <= n1865;
    \\ks1_key_reg_reg[19]  <= n1870;
    \\ks1_key_reg_reg[18]  <= n1875;
    \\ks1_key_reg_reg[21]  <= n1880;
    \\ks1_key_reg_reg[22]  <= n1885;
    \\ks1_key_reg_reg[20]  <= n1890;
    \\ks1_key_reg_reg[57]  <= n1895;
    \\ks1_key_reg_reg[58]  <= n1900;
    \\ks1_key_reg_reg[63]  <= n1905;
    \\ks1_key_reg_reg[62]  <= n1910;
    \\ks1_key_reg_reg[56]  <= n1915;
    \\ks1_key_reg_reg[92]  <= n1920;
    \\ks1_key_reg_reg[32]  <= n1925;
    \\ks1_key_reg_reg[33]  <= n1930;
    \\ks1_key_reg_reg[34]  <= n1935;
    \\ks1_key_reg_reg[35]  <= n1940;
    \\ks1_key_reg_reg[36]  <= n1945;
    \\ks1_key_reg_reg[38]  <= n1950;
    \\ks1_key_reg_reg[39]  <= n1955;
    \\ks1_key_reg_reg[55]  <= n1960;
    \\ks1_key_reg_reg[37]  <= n1965;
    \\ks1_key_reg_reg[91]  <= n1970;
    \\ks1_key_reg_reg[93]  <= n1975;
    \\ks1_key_reg_reg[49]  <= n1980;
    \\ks1_key_reg_reg[50]  <= n1985;
    \\ks1_key_reg_reg[51]  <= n1990;
    \\ks1_key_reg_reg[52]  <= n1995;
    \\ks1_key_reg_reg[54]  <= n2000;
    \\ks1_key_reg_reg[48]  <= n2005;
    \\ks1_key_reg_reg[53]  <= n2010;
    \\ks1_key_reg_reg[90]  <= n2015;
    \\ks1_key_reg_reg[88]  <= n2020;
    \\ks1_key_reg_reg[94]  <= n2025;
    \\ks1_key_reg_reg[95]  <= n2030;
    \\ks1_key_reg_reg[89]  <= n2035;
    \\ks1_key_reg_reg[69]  <= n2040;
    \\addroundkey_data_reg_reg[60]  <= n2045;
    \\addroundkey_data_reg_reg[111]  <= n2050;
    \\addroundkey_data_reg_reg[63]  <= n2055;
    \\addroundkey_data_reg_reg[6]  <= n2060;
    \\addroundkey_data_reg_reg[76]  <= n2065;
    \\addroundkey_data_reg_reg[25]  <= n2070;
    \\addroundkey_data_reg_reg[77]  <= n2075;
    \\addroundkey_data_reg_reg[78]  <= n2080;
    \\addroundkey_data_reg_reg[79]  <= n2085;
    \\addroundkey_data_reg_reg[26]  <= n2090;
    \\addroundkey_data_reg_reg[29]  <= n2095;
    \\addroundkey_data_reg_reg[8]  <= n2100;
    \\addroundkey_data_reg_reg[105]  <= n2105;
    \\addroundkey_data_reg_reg[0]  <= n2110;
    \\addroundkey_data_reg_reg[106]  <= n2115;
    \\addroundkey_data_reg_reg[107]  <= n2120;
    \\addroundkey_data_reg_reg[122]  <= n2125;
    \\addroundkey_data_reg_reg[3]  <= n2130;
    \\addroundkey_data_reg_reg[41]  <= n2135;
    \\addroundkey_data_reg_reg[123]  <= n2140;
    \\addroundkey_data_reg_reg[42]  <= n2145;
    \\addroundkey_data_reg_reg[43]  <= n2150;
    \\addroundkey_data_reg_reg[44]  <= n2155;
    \\addroundkey_data_reg_reg[108]  <= n2160;
    \\addroundkey_data_reg_reg[125]  <= n2165;
    \\addroundkey_data_reg_reg[46]  <= n2170;
    \\addroundkey_data_reg_reg[47]  <= n2175;
    \\addroundkey_data_reg_reg[126]  <= n2180;
    \\addroundkey_data_reg_reg[127]  <= n2185;
    \\addroundkey_data_reg_reg[10]  <= n2190;
    \\addroundkey_data_reg_reg[13]  <= n2195;
    \\addroundkey_data_reg_reg[110]  <= n2200;
    \\addroundkey_data_reg_reg[58]  <= n2205;
    \\addroundkey_data_reg_reg[57]  <= n2210;
    \\addroundkey_data_reg_reg[59]  <= n2215;
    \\ks1_key_reg_reg[124]  <= n2220;
    \\ks1_key_reg_reg[64]  <= n2225;
    \\ks1_key_reg_reg[65]  <= n2230;
    \\ks1_key_reg_reg[67]  <= n2235;
    \\ks1_key_reg_reg[66]  <= n2240;
    \\ks1_key_reg_reg[68]  <= n2245;
    \\ks1_key_reg_reg[70]  <= n2250;
    \\ks1_key_reg_reg[71]  <= n2255;
    \\ks1_key_reg_reg[87]  <= n2260;
    \\addroundkey_data_reg_reg[5]  <= n2265;
    \\ks1_key_reg_reg[81]  <= n2270;
    \\addroundkey_data_reg_reg[40]  <= n2275;
    \\addroundkey_data_reg_reg[124]  <= n2280;
    \\addroundkey_data_reg_reg[61]  <= n2285;
    \\addroundkey_data_reg_reg[62]  <= n2290;
    \\addroundkey_data_reg_reg[1]  <= n2295;
    \\addroundkey_data_reg_reg[73]  <= n2300;
    \\addroundkey_data_reg_reg[74]  <= n2305;
    \\addroundkey_data_reg_reg[24]  <= n2310;
    \\addroundkey_data_reg_reg[72]  <= n2315;
    \\addroundkey_data_reg_reg[7]  <= n2320;
    \\addroundkey_data_reg_reg[28]  <= n2325;
    \\addroundkey_data_reg_reg[104]  <= n2330;
    \\addroundkey_data_reg_reg[30]  <= n2335;
    \\addroundkey_data_reg_reg[2]  <= n2340;
    \\addroundkey_data_reg_reg[31]  <= n2345;
    \\addroundkey_data_reg_reg[90]  <= n2350;
    \\addroundkey_data_reg_reg[91]  <= n2355;
    \\addroundkey_data_reg_reg[92]  <= n2360;
    \\addroundkey_data_reg_reg[34]  <= n2365;
    \\addroundkey_data_reg_reg[93]  <= n2370;
    \\addroundkey_data_reg_reg[11]  <= n2375;
    \\addroundkey_data_reg_reg[94]  <= n2380;
    \\addroundkey_data_reg_reg[95]  <= n2385;
    \\addroundkey_data_reg_reg[120]  <= n2390;
    \\addroundkey_data_reg_reg[9]  <= n2395;
    \\addroundkey_data_reg_reg[121]  <= n2400;
    \\addroundkey_data_reg_reg[45]  <= n2405;
    \\addroundkey_data_reg_reg[4]  <= n2410;
    \\addroundkey_data_reg_reg[12]  <= n2415;
    \\addroundkey_data_reg_reg[109]  <= n2420;
    \\addroundkey_data_reg_reg[14]  <= n2425;
    \\addroundkey_data_reg_reg[56]  <= n2430;
    \\addroundkey_data_reg_reg[15]  <= n2435;
    \\ks1_key_reg_reg[125]  <= n2440;
    \\ks1_key_reg_reg[123]  <= n2445;
    \\ks1_key_reg_reg[80]  <= n2450;
    \\ks1_key_reg_reg[83]  <= n2455;
    \\ks1_key_reg_reg[84]  <= n2460;
    \\ks1_key_reg_reg[85]  <= n2465;
    \\ks1_key_reg_reg[82]  <= n2470;
    \\ks1_key_reg_reg[86]  <= n2475;
    \\addroundkey_data_reg_reg[27]  <= n2480;
    \\addroundkey_data_reg_reg[75]  <= n2485;
    \\addroundkey_data_reg_reg[100]  <= n2490;
    \\addroundkey_data_reg_reg[33]  <= n2495;
    \\addroundkey_data_reg_reg[103]  <= n2500;
    \\addroundkey_data_reg_reg[98]  <= n2505;
    \\addroundkey_data_reg_reg[35]  <= n2510;
    \\mix1_data_reg_reg[100]  <= n2515;
    \\mix1_data_reg_reg[108]  <= n2520;
    \\mix1_data_reg_reg[116]  <= n2525;
    \\mix1_data_reg_reg[124]  <= n2530;
    \\addroundkey_data_reg_reg[101]  <= n2535;
    \\addroundkey_data_reg_reg[112]  <= n2540;
    \\addroundkey_data_reg_reg[64]  <= n2545;
    \\addroundkey_data_reg_reg[65]  <= n2550;
    \\addroundkey_data_reg_reg[20]  <= n2555;
    \\addroundkey_data_reg_reg[66]  <= n2560;
    \\addroundkey_data_reg_reg[67]  <= n2565;
    \\addroundkey_data_reg_reg[21]  <= n2570;
    \\addroundkey_data_reg_reg[69]  <= n2575;
    \\addroundkey_data_reg_reg[22]  <= n2580;
    \\addroundkey_data_reg_reg[70]  <= n2585;
    \\addroundkey_data_reg_reg[102]  <= n2590;
    \\addroundkey_data_reg_reg[23]  <= n2595;
    \\addroundkey_data_reg_reg[115]  <= n2600;
    \\addroundkey_data_reg_reg[116]  <= n2605;
    \\addroundkey_data_reg_reg[80]  <= n2610;
    \\addroundkey_data_reg_reg[81]  <= n2615;
    \\addroundkey_data_reg_reg[83]  <= n2620;
    \\addroundkey_data_reg_reg[85]  <= n2625;
    \\addroundkey_data_reg_reg[86]  <= n2630;
    \\addroundkey_data_reg_reg[84]  <= n2635;
    \\addroundkey_data_reg_reg[87]  <= n2640;
    \\addroundkey_data_reg_reg[88]  <= n2645;
    \\addroundkey_data_reg_reg[32]  <= n2650;
    \\addroundkey_data_reg_reg[119]  <= n2655;
    \\addroundkey_data_reg_reg[96]  <= n2660;
    \\addroundkey_data_reg_reg[97]  <= n2665;
    \\addroundkey_data_reg_reg[36]  <= n2670;
    \\addroundkey_data_reg_reg[99]  <= n2675;
    \\addroundkey_data_reg_reg[37]  <= n2680;
    \\addroundkey_data_reg_reg[38]  <= n2685;
    \\addroundkey_data_reg_reg[39]  <= n2690;
    \\addroundkey_data_reg_reg[49]  <= n2695;
    \\addroundkey_data_reg_reg[52]  <= n2700;
    \\addroundkey_data_reg_reg[55]  <= n2705;
    \\addroundkey_data_reg_reg[17]  <= n2710;
    \\ks1_key_reg_reg[120]  <= n2715;
    \\ks1_key_reg_reg[121]  <= n2720;
    \\ks1_key_reg_reg[127]  <= n2725;
    \\addroundkey_round_reg[0]  <= n2730;
    \\addroundkey_data_reg_reg[118]  <= n2735;
    \\addroundkey_data_reg_reg[89]  <= n2740;
    \\addroundkey_data_reg_reg[117]  <= n2745;
    \\ks1_key_reg_reg[126]  <= n2750;
    \\addroundkey_data_reg_reg[82]  <= n2755;
    \\ks1_key_reg_reg[122]  <= n2760;
    \\addroundkey_data_reg_reg[114]  <= n2765;
    \\addroundkey_data_reg_reg[54]  <= n2770;
    \\addroundkey_data_reg_reg[71]  <= n2775;
    \\addroundkey_data_reg_reg[16]  <= n2780;
    \\addroundkey_data_reg_reg[68]  <= n2785;
    \\addroundkey_data_reg_reg[53]  <= n2790;
    \\addroundkey_data_reg_reg[113]  <= n2795;
    \\addroundkey_data_reg_reg[19]  <= n2800;
    \\addroundkey_data_reg_reg[51]  <= n2805;
    \\addroundkey_data_reg_reg[50]  <= n2810;
    \\addroundkey_data_reg_reg[18]  <= n2815;
    \\addroundkey_data_reg_reg[48]  <= n2820;
    \\ks1_key_reg_reg[97]  <= n2825;
    \\mix1_data_reg_reg[107]  <= n2830;
    \\mix1_data_reg_reg[115]  <= n2835;
    \\mix1_data_reg_reg[99]  <= n2840;
    \\ks1_key_reg_reg[96]  <= n2845;
    \\ks1_key_reg_reg[98]  <= n2850;
    \\ks1_key_reg_reg[100]  <= n2855;
    \\ks1_key_reg_reg[101]  <= n2860;
    \\ks1_key_reg_reg[102]  <= n2865;
    \\ks1_key_reg_reg[103]  <= n2870;
    \\ks1_key_reg_reg[119]  <= n2875;
    \\mix1_data_reg_reg[123]  <= n2880;
    \\ks1_key_reg_reg[113]  <= n2885;
    \\mix1_data_reg_reg[36]  <= n2890;
    \\mix1_data_reg_reg[44]  <= n2895;
    \\mix1_data_reg_reg[60]  <= n2900;
    \\mix1_data_reg_reg[68]  <= n2905;
    \\mix1_data_reg_reg[52]  <= n2910;
    \\mix1_data_reg_reg[84]  <= n2915;
    \\mix1_data_reg_reg[76]  <= n2920;
    \\mix1_data_reg_reg[92]  <= n2925;
    \\ks1_key_reg_reg[112]  <= n2930;
    \\ks1_key_reg_reg[115]  <= n2935;
    \\ks1_key_reg_reg[116]  <= n2940;
    \\ks1_key_reg_reg[114]  <= n2945;
    \\ks1_key_reg_reg[118]  <= n2950;
    addroundkey_ready_o_reg <= n2955;
    \\ks1_key_reg_reg[117]  <= n2960;
    \\ks1_key_reg_reg[99]  <= n2965;
    \\mix1_data_reg_reg[105]  <= n2970;
    \\mix1_data_reg_reg[106]  <= n2975;
    \\mix1_data_reg_reg[113]  <= n2980;
    \\mix1_data_reg_reg[114]  <= n2985;
    \\mix1_data_reg_reg[121]  <= n2990;
    \\mix1_data_reg_reg[122]  <= n2995;
    \\mix1_data_reg_reg[35]  <= n3000;
    \\mix1_data_reg_reg[43]  <= n3005;
    \\mix1_data_reg_reg[51]  <= n3010;
    \\mix1_data_reg_reg[59]  <= n3015;
    \\mix1_data_reg_reg[67]  <= n3020;
    \\mix1_data_reg_reg[75]  <= n3025;
    \\mix1_data_reg_reg[97]  <= n3030;
    \\mix1_data_reg_reg[98]  <= n3035;
    \\mix1_data_reg_reg[91]  <= n3040;
    \\mix1_data_reg_reg[83]  <= n3045;
    \\mix1_data_reg_reg[120]  <= n3050;
    \\mix1_data_reg_reg[117]  <= n3055;
    \\mix1_data_reg_reg[125]  <= n3060;
    \\mix1_data_reg_reg[118]  <= n3065;
    \\mix1_data_reg_reg[104]  <= n3070;
    \\mix1_data_reg_reg[112]  <= n3075;
    \\mix1_data_reg_reg[96]  <= n3080;
    \\mix1_data_reg_reg[126]  <= n3085;
    \\mix1_data_reg_reg[110]  <= n3090;
    \\mix1_data_reg_reg[102]  <= n3095;
    \\mix1_data_reg_reg[109]  <= n3100;
    \\mix1_data_reg_reg[101]  <= n3105;
    \\mix1_data_o_reg_reg[12]  <= n3110;
    \\mix1_data_o_reg_reg[20]  <= n3115;
    \\mix1_data_o_reg_reg[28]  <= n3120;
    \\mix1_data_o_reg_reg[4]  <= n3125;
    \\mix1_data_reg_reg[33]  <= n3130;
    \\mix1_data_reg_reg[34]  <= n3135;
    \\mix1_data_reg_reg[42]  <= n3140;
    \\mix1_data_reg_reg[41]  <= n3145;
    \\mix1_data_reg_reg[49]  <= n3150;
    \\mix1_data_reg_reg[50]  <= n3155;
    \\mix1_data_reg_reg[57]  <= n3160;
    \\mix1_data_reg_reg[58]  <= n3165;
    \\mix1_data_reg_reg[65]  <= n3170;
    \\mix1_data_reg_reg[66]  <= n3175;
    \\mix1_data_reg_reg[74]  <= n3180;
    \\mix1_data_reg_reg[73]  <= n3185;
    \\mix1_data_reg_reg[81]  <= n3190;
    \\mix1_data_reg_reg[82]  <= n3195;
    \\mix1_data_reg_reg[89]  <= n3200;
    \\mix1_data_reg_reg[90]  <= n3205;
    \\mix1_data_reg_reg[61]  <= n3210;
    \\mix1_data_reg_reg[62]  <= n3215;
    \\mix1_data_reg_reg[69]  <= n3220;
    \\mix1_data_reg_reg[45]  <= n3225;
    \\mix1_data_reg_reg[37]  <= n3230;
    \\mix1_data_reg_reg[53]  <= n3235;
    \\mix1_data_reg_reg[77]  <= n3240;
    \\mix1_data_o_reg_reg[3]  <= n3245;
    \\mix1_data_reg_reg[38]  <= n3250;
    \\mix1_data_reg_reg[46]  <= n3255;
    \\mix1_data_reg_reg[54]  <= n3260;
    \\mix1_data_reg_reg[70]  <= n3265;
    \\mix1_data_reg_reg[78]  <= n3270;
    \\mix1_data_reg_reg[86]  <= n3275;
    \\mix1_data_reg_reg[94]  <= n3280;
    \\mix1_data_reg_reg[32]  <= n3285;
    \\mix1_data_reg_reg[48]  <= n3290;
    \\mix1_data_reg_reg[56]  <= n3295;
    \\mix1_data_reg_reg[64]  <= n3300;
    \\mix1_data_reg_reg[88]  <= n3305;
    \\mix1_data_reg_reg[80]  <= n3310;
    \\mix1_data_reg_reg[72]  <= n3315;
    \\mix1_data_reg_reg[40]  <= n3320;
    \\mix1_data_o_reg_reg[27]  <= n3325;
    \\mix1_data_o_reg_reg[11]  <= n3330;
    \\mix1_data_o_reg_reg[19]  <= n3335;
    \\mix1_data_reg_reg[85]  <= n3340;
    \\mix1_data_reg_reg[93]  <= n3345;
    \\mix1_data_reg_reg[103]  <= n3350;
    \\mix1_data_reg_reg[111]  <= n3355;
    \\mix1_data_reg_reg[127]  <= n3360;
    \\mix1_data_reg_reg[119]  <= n3365;
    \\mix1_data_o_reg_reg[17]  <= n3370;
    \\mix1_data_o_reg_reg[18]  <= n3375;
    \\mix1_data_o_reg_reg[1]  <= n3380;
    \\mix1_data_o_reg_reg[25]  <= n3385;
    \\mix1_data_o_reg_reg[26]  <= n3390;
    \\mix1_data_o_reg_reg[9]  <= n3395;
    \\mix1_data_o_reg_reg[2]  <= n3400;
    \\mix1_data_o_reg_reg[10]  <= n3405;
    \\mix1_data_reg_reg[79]  <= n3410;
    \\mix1_data_o_reg_reg[8]  <= n3415;
    \\mix1_data_reg_reg[55]  <= n3420;
    \\mix1_data_reg_reg[71]  <= n3425;
    \\mix1_data_o_reg_reg[13]  <= n3430;
    \\mix1_data_o_reg_reg[21]  <= n3435;
    \\mix1_data_reg_reg[63]  <= n3440;
    \\mix1_data_o_reg_reg[22]  <= n3445;
    \\mix1_data_o_reg_reg[30]  <= n3450;
    \\mix1_data_o_reg_reg[16]  <= n3455;
    \\mix1_data_reg_reg[47]  <= n3460;
    \\mix1_data_reg_reg[39]  <= n3465;
    \\mix1_data_o_reg_reg[6]  <= n3470;
    \\mix1_data_o_reg_reg[14]  <= n3475;
    \\mix1_data_o_reg_reg[0]  <= n3480;
    \\mix1_data_o_reg_reg[24]  <= n3485;
    \\mix1_data_reg_reg[95]  <= n3490;
    \\mix1_data_o_reg_reg[29]  <= n3495;
    \\mix1_data_o_reg_reg[5]  <= n3500;
    \\mix1_data_reg_reg[87]  <= n3505;
    \\mix1_data_o_reg_reg[7]  <= n3510;
    \\mix1_data_o_reg_reg[23]  <= n3515;
    \\mix1_data_o_reg_reg[31]  <= n3520;
    \\mix1_data_o_reg_reg[15]  <= n3525;
    \\addroundkey_round_reg[1]  <= n3530;
    \\addroundkey_round_reg[3]  <= n3535;
    \\addroundkey_round_reg[2]  <= n3540;
    \\ks1_state_reg[0]  <= n3545;
    \\ks1_state_reg[2]  <= n3550;
    \\round_reg[1]  <= n3555;
    \\round_reg[2]  <= n3560;
    \\round_reg[0]  <= n3565;
    \\round_reg[3]  <= n3570;
    addroundkey_start_i_reg <= n3575;
    \\mix1_state_reg[0]  <= n3580;
    \\mix1_state_reg[1]  <= n3585;
    state_reg <= n3590;
    \\sub1_state_reg[0]  <= n3595;
    ready_o_reg <= n3600;
    \\sub1_state_reg[3]  <= n3605;
    \\sub1_state_reg[2]  <= n3610;
    \\sub1_state_reg[1]  <= n3615;
    \\sub1_state_reg[4]  <= n3620;
    \\mix1_data_o_reg_reg[104]  <= n3625;
    \\mix1_data_o_reg_reg[102]  <= n3630;
    \\mix1_data_o_reg_reg[105]  <= n3635;
    \\mix1_data_o_reg_reg[108]  <= n3640;
    \\mix1_data_o_reg_reg[110]  <= n3645;
    \\mix1_data_o_reg_reg[112]  <= n3650;
    \\mix1_data_o_reg_reg[45]  <= n3655;
    \\mix1_data_o_reg_reg[67]  <= n3660;
    \\mix1_data_o_reg_reg[70]  <= n3665;
    \\mix1_data_o_reg_reg[85]  <= n3670;
    \\mix1_data_o_reg_reg[98]  <= n3675;
    \\mix1_data_o_reg_reg[82]  <= n3680;
    \\mix1_data_o_reg_reg[99]  <= n3685;
    \\mix1_data_o_reg_reg[72]  <= n3690;
    \\mix1_data_o_reg_reg[48]  <= n3695;
    \\mix1_data_o_reg_reg[91]  <= n3700;
    \\mix1_data_o_reg_reg[69]  <= n3705;
    \\mix1_data_o_reg_reg[57]  <= n3710;
    \\mix1_data_o_reg_reg[33]  <= n3715;
    \\mix1_data_o_reg_reg[65]  <= n3720;
    \\mix1_data_o_reg_reg[71]  <= n3725;
    \\mix1_data_o_reg_reg[93]  <= n3730;
    \\mix1_data_o_reg_reg[106]  <= n3735;
    \\mix1_data_o_reg_reg[77]  <= n3740;
    \\mix1_data_o_reg_reg[78]  <= n3745;
    \\mix1_data_o_reg_reg[122]  <= n3750;
    \\mix1_data_o_reg_reg[64]  <= n3755;
    \\mix1_data_o_reg_reg[49]  <= n3760;
    \\mix1_data_o_reg_reg[116]  <= n3765;
    \\mix1_data_o_reg_reg[86]  <= n3770;
    \\mix1_data_o_reg_reg[88]  <= n3775;
    \\mix1_data_o_reg_reg[89]  <= n3780;
    \\mix1_data_o_reg_reg[126]  <= n3785;
    \\mix1_data_o_reg_reg[90]  <= n3790;
    \\mix1_data_o_reg_reg[74]  <= n3795;
    \\mix1_data_o_reg_reg[56]  <= n3800;
    \\mix1_data_o_reg_reg[47]  <= n3805;
    \\mix1_data_o_reg_reg[97]  <= n3810;
    \\mix1_data_o_reg_reg[43]  <= n3815;
    \\mix1_data_o_reg_reg[76]  <= n3820;
    \\mix1_data_o_reg_reg[37]  <= n3825;
    \\mix1_data_o_reg_reg[84]  <= n3830;
    \\mix1_data_o_reg_reg[103]  <= n3835;
    \\mix1_data_o_reg_reg[109]  <= n3840;
    \\mix1_data_o_reg_reg[53]  <= n3845;
    \\mix1_data_o_reg_reg[119]  <= n3850;
    \\mix1_data_o_reg_reg[125]  <= n3855;
    \\mix1_data_o_reg_reg[36]  <= n3860;
    \\mix1_data_o_reg_reg[39]  <= n3865;
    \\mix1_data_o_reg_reg[55]  <= n3870;
    \\mix1_data_o_reg_reg[62]  <= n3875;
    \\mix1_data_o_reg_reg[96]  <= n3880;
    \\mix1_data_o_reg_reg[115]  <= n3885;
    \\mix1_data_o_reg_reg[46]  <= n3890;
    \\mix1_data_o_reg_reg[80]  <= n3895;
    \\mix1_data_o_reg_reg[123]  <= n3900;
    \\mix1_data_o_reg_reg[83]  <= n3905;
    \\mix1_data_o_reg_reg[58]  <= n3910;
    \\mix1_data_o_reg_reg[68]  <= n3915;
    \\mix1_data_o_reg_reg[101]  <= n3920;
    \\mix1_data_o_reg_reg[118]  <= n3925;
    \\mix1_data_o_reg_reg[52]  <= n3930;
    \\mix1_data_o_reg_reg[59]  <= n3935;
    \\mix1_data_o_reg_reg[87]  <= n3940;
    \\mix1_data_o_reg_reg[51]  <= n3945;
    \\mix1_data_o_reg_reg[66]  <= n3950;
    \\mix1_data_o_reg_reg[81]  <= n3955;
    \\mix1_data_o_reg_reg[107]  <= n3960;
    \\mix1_data_o_reg_reg[44]  <= n3965;
    \\mix1_data_o_reg_reg[42]  <= n3970;
    \\mix1_data_o_reg_reg[94]  <= n3975;
    \\mix1_data_o_reg_reg[54]  <= n3980;
    \\mix1_data_o_reg_reg[50]  <= n3985;
    \\mix1_data_o_reg_reg[124]  <= n3990;
    \\mix1_data_o_reg_reg[32]  <= n3995;
    \\mix1_data_o_reg_reg[75]  <= n4000;
    \\mix1_data_o_reg_reg[61]  <= n4005;
    \\mix1_data_o_reg_reg[63]  <= n4010;
    \\mix1_data_o_reg_reg[120]  <= n4015;
    \\mix1_data_o_reg_reg[40]  <= n4020;
    \\mix1_data_o_reg_reg[111]  <= n4025;
    \\mix1_data_o_reg_reg[34]  <= n4030;
    \\mix1_data_o_reg_reg[113]  <= n4035;
    \\mix1_data_o_reg_reg[41]  <= n4040;
    \\mix1_data_o_reg_reg[121]  <= n4045;
    \\mix1_data_o_reg_reg[92]  <= n4050;
    \\mix1_data_o_reg_reg[117]  <= n4055;
    \\mix1_data_o_reg_reg[60]  <= n4060;
    \\mix1_data_o_reg_reg[114]  <= n4065;
    \\mix1_data_o_reg_reg[38]  <= n4070;
    \\mix1_data_o_reg_reg[73]  <= n4075;
    \\mix1_data_o_reg_reg[127]  <= n4080;
    \\mix1_data_o_reg_reg[95]  <= n4085;
    \\mix1_data_o_reg_reg[79]  <= n4090;
    \\mix1_data_o_reg_reg[35]  <= n4095;
    \\mix1_data_o_reg_reg[100]  <= n4100;
    ks1_ready_o_reg <= n4105;
    mix1_ready_o_reg <= n4110;
    first_round_reg_reg <= n4115;
    \\ks1_state_reg[1]  <= n4120;
    sub1_ready_o_reg <= n4125;
  end
  initial begin
    \\ks1_key_reg_reg[11]  <= 1'b0;
    \\ks1_key_reg_reg[12]  <= 1'b0;
    \\ks1_key_reg_reg[13]  <= 1'b0;
    \\ks1_key_reg_reg[14]  <= 1'b0;
    \\ks1_key_reg_reg[15]  <= 1'b0;
    \\sbox1_to_invert_reg[1]  <= 1'b0;
    \\sbox1_to_invert_reg[3]  <= 1'b0;
    \\sbox1_to_invert_reg[2]  <= 1'b0;
    \\sbox1_to_invert_reg[0]  <= 1'b0;
    \\ks1_key_reg_reg[8]  <= 1'b0;
    \\ks1_key_reg_reg[10]  <= 1'b0;
    \\ks1_key_reg_reg[9]  <= 1'b0;
    \\ks1_key_reg_reg[43]  <= 1'b0;
    \\ks1_key_reg_reg[44]  <= 1'b0;
    \\ks1_key_reg_reg[45]  <= 1'b0;
    \\ks1_key_reg_reg[46]  <= 1'b0;
    \\ks1_key_reg_reg[47]  <= 1'b0;
    \\ks1_key_reg_reg[40]  <= 1'b0;
    \\sub1_data_reg_reg[109]  <= 1'b0;
    \\sub1_data_reg_reg[110]  <= 1'b0;
    \\sub1_data_reg_reg[13]  <= 1'b0;
    \\sub1_data_reg_reg[14]  <= 1'b0;
    \\sub1_data_reg_reg[45]  <= 1'b0;
    \\sub1_data_reg_reg[46]  <= 1'b0;
    \\sub1_data_reg_reg[77]  <= 1'b0;
    \\sub1_data_reg_reg[78]  <= 1'b0;
    \\sub1_data_reg_reg[102]  <= 1'b0;
    \\sub1_data_reg_reg[101]  <= 1'b0;
    \\sub1_data_reg_reg[118]  <= 1'b0;
    \\sub1_data_reg_reg[117]  <= 1'b0;
    \\sub1_data_reg_reg[21]  <= 1'b0;
    \\sub1_data_reg_reg[22]  <= 1'b0;
    \\sub1_data_reg_reg[37]  <= 1'b0;
    \\sub1_data_reg_reg[38]  <= 1'b0;
    \\sub1_data_reg_reg[53]  <= 1'b0;
    \\sub1_data_reg_reg[54]  <= 1'b0;
    \\sub1_data_reg_reg[5]  <= 1'b0;
    \\sub1_data_reg_reg[6]  <= 1'b0;
    \\sub1_data_reg_reg[70]  <= 1'b0;
    \\sub1_data_reg_reg[69]  <= 1'b0;
    \\sub1_data_reg_reg[85]  <= 1'b0;
    \\sub1_data_reg_reg[86]  <= 1'b0;
    \\ks1_key_reg_reg[42]  <= 1'b0;
    \\ks1_key_reg_reg[41]  <= 1'b0;
    \\ks1_key_reg_reg[76]  <= 1'b0;
    \\ks1_key_reg_reg[75]  <= 1'b0;
    \\ks1_key_reg_reg[74]  <= 1'b0;
    \\ks1_key_reg_reg[73]  <= 1'b0;
    \\ks1_key_reg_reg[77]  <= 1'b0;
    \\ks1_key_reg_reg[78]  <= 1'b0;
    \\sub1_data_reg_reg[125]  <= 1'b0;
    \\sub1_data_reg_reg[126]  <= 1'b0;
    \\sub1_data_reg_reg[29]  <= 1'b0;
    \\sub1_data_reg_reg[94]  <= 1'b0;
    \\sub1_data_reg_reg[30]  <= 1'b0;
    \\sub1_data_reg_reg[93]  <= 1'b0;
    \\ks1_key_reg_reg[72]  <= 1'b0;
    \\ks1_key_reg_reg[79]  <= 1'b0;
    \\sub1_data_reg_reg[104]  <= 1'b0;
    \\sub1_data_reg_reg[40]  <= 1'b0;
    \\sub1_data_reg_reg[72]  <= 1'b0;
    \\sub1_data_reg_reg[8]  <= 1'b0;
    \\sub1_data_reg_reg[0]  <= 1'b0;
    \\sub1_data_reg_reg[112]  <= 1'b0;
    \\sub1_data_reg_reg[16]  <= 1'b0;
    \\sub1_data_reg_reg[64]  <= 1'b0;
    \\sub1_data_reg_reg[80]  <= 1'b0;
    \\sub1_data_reg_reg[96]  <= 1'b0;
    \\sub1_data_reg_reg[48]  <= 1'b0;
    \\sub1_data_reg_reg[61]  <= 1'b0;
    \\sub1_data_reg_reg[62]  <= 1'b0;
    \\ks1_col_reg[21]  <= 1'b0;
    \\ks1_col_reg[22]  <= 1'b0;
    \\sub1_data_reg_reg[107]  <= 1'b0;
    \\sub1_data_reg_reg[108]  <= 1'b0;
    \\sub1_data_reg_reg[111]  <= 1'b0;
    \\sub1_data_reg_reg[11]  <= 1'b0;
    \\sub1_data_reg_reg[12]  <= 1'b0;
    \\sub1_data_reg_reg[15]  <= 1'b0;
    \\sub1_data_reg_reg[44]  <= 1'b0;
    \\sub1_data_reg_reg[43]  <= 1'b0;
    \\sub1_data_reg_reg[47]  <= 1'b0;
    \\sub1_data_reg_reg[75]  <= 1'b0;
    \\sub1_data_reg_reg[76]  <= 1'b0;
    \\sub1_data_reg_reg[79]  <= 1'b0;
    \\sub1_data_reg_reg[103]  <= 1'b0;
    \\sub1_data_reg_reg[115]  <= 1'b0;
    \\sub1_data_reg_reg[116]  <= 1'b0;
    \\sub1_data_reg_reg[119]  <= 1'b0;
    \\sub1_data_reg_reg[20]  <= 1'b0;
    \\sub1_data_reg_reg[19]  <= 1'b0;
    \\sub1_data_reg_reg[23]  <= 1'b0;
    \\sub1_data_reg_reg[32]  <= 1'b0;
    \\sub1_data_reg_reg[4]  <= 1'b0;
    \\sub1_data_reg_reg[51]  <= 1'b0;
    \\sub1_data_reg_reg[52]  <= 1'b0;
    \\sub1_data_reg_reg[55]  <= 1'b0;
    \\sub1_data_reg_reg[36]  <= 1'b0;
    \\sub1_data_reg_reg[68]  <= 1'b0;
    \\sub1_data_reg_reg[67]  <= 1'b0;
    \\sub1_data_reg_reg[3]  <= 1'b0;
    \\sub1_data_reg_reg[7]  <= 1'b0;
    \\sub1_data_reg_reg[71]  <= 1'b0;
    \\sub1_data_reg_reg[84]  <= 1'b0;
    \\sub1_data_reg_reg[83]  <= 1'b0;
    \\sub1_data_reg_reg[87]  <= 1'b0;
    \\sub1_data_reg_reg[120]  <= 1'b0;
    \\sub1_data_reg_reg[24]  <= 1'b0;
    \\sub1_data_reg_reg[56]  <= 1'b0;
    \\sub1_data_reg_reg[88]  <= 1'b0;
    \\sbox1_alph_reg[2]  <= 1'b0;
    \\ks1_col_reg[30]  <= 1'b0;
    \\sub1_data_reg_reg[100]  <= 1'b0;
    \\ks1_col_reg[6]  <= 1'b0;
    \\ks1_col_reg[5]  <= 1'b0;
    \\sub1_data_reg_reg[35]  <= 1'b0;
    \\sub1_data_reg_reg[39]  <= 1'b0;
    \\ks1_col_reg[29]  <= 1'b0;
    \\sub1_data_reg_reg[99]  <= 1'b0;
    \\sub1_data_reg_reg[123]  <= 1'b0;
    \\sub1_data_reg_reg[124]  <= 1'b0;
    \\sub1_data_reg_reg[127]  <= 1'b0;
    \\sub1_data_reg_reg[27]  <= 1'b0;
    \\sub1_data_reg_reg[28]  <= 1'b0;
    \\sub1_data_reg_reg[31]  <= 1'b0;
    \\sub1_data_reg_reg[59]  <= 1'b0;
    \\sub1_data_reg_reg[60]  <= 1'b0;
    \\sub1_data_reg_reg[63]  <= 1'b0;
    \\sub1_data_reg_reg[95]  <= 1'b0;
    \\sub1_data_reg_reg[91]  <= 1'b0;
    \\sub1_data_reg_reg[92]  <= 1'b0;
    \\ks1_col_reg[16]  <= 1'b0;
    \\sbox1_alph_reg[0]  <= 1'b0;
    \\ks1_key_reg_reg[107]  <= 1'b0;
    \\ks1_key_reg_reg[108]  <= 1'b0;
    \\ks1_col_reg[20]  <= 1'b0;
    \\ks1_key_reg_reg[104]  <= 1'b0;
    \\ks1_col_reg[23]  <= 1'b0;
    \\ks1_col_reg[19]  <= 1'b0;
    \\sub1_data_reg_reg[106]  <= 1'b0;
    \\sub1_data_reg_reg[10]  <= 1'b0;
    \\sub1_data_reg_reg[74]  <= 1'b0;
    \\sub1_data_reg_reg[42]  <= 1'b0;
    \\sub1_data_reg_reg[114]  <= 1'b0;
    \\ks1_col_reg[24]  <= 1'b0;
    \\ks1_col_reg[3]  <= 1'b0;
    \\ks1_col_reg[4]  <= 1'b0;
    \\sub1_data_reg_reg[18]  <= 1'b0;
    \\sub1_data_reg_reg[2]  <= 1'b0;
    \\sub1_data_reg_reg[50]  <= 1'b0;
    \\sub1_data_reg_reg[66]  <= 1'b0;
    \\sub1_data_reg_reg[82]  <= 1'b0;
    \\sub1_data_reg_reg[98]  <= 1'b0;
    \\ks1_col_reg[0]  <= 1'b0;
    \\ks1_col_reg[28]  <= 1'b0;
    \\ks1_key_reg_reg[111]  <= 1'b0;
    \\ks1_col_reg[27]  <= 1'b0;
    \\ks1_col_reg[31]  <= 1'b0;
    \\sub1_data_reg_reg[34]  <= 1'b0;
    \\ks1_col_reg[7]  <= 1'b0;
    \\sub1_data_reg_reg[122]  <= 1'b0;
    \\sub1_data_reg_reg[26]  <= 1'b0;
    \\sub1_data_reg_reg[58]  <= 1'b0;
    \\sub1_data_reg_reg[90]  <= 1'b0;
    \\sbox1_ah_reg_reg[2]  <= 1'b0;
    \\sbox1_alph_reg[1]  <= 1'b0;
    \\ks1_key_reg_reg[110]  <= 1'b0;
    \\ks1_key_reg_reg[109]  <= 1'b0;
    \\sub1_data_reg_reg[105]  <= 1'b0;
    \\sub1_data_reg_reg[41]  <= 1'b0;
    \\sub1_data_reg_reg[73]  <= 1'b0;
    \\sub1_data_reg_reg[9]  <= 1'b0;
    \\sub1_data_reg_reg[17]  <= 1'b0;
    \\sub1_data_reg_reg[1]  <= 1'b0;
    \\sub1_data_reg_reg[65]  <= 1'b0;
    \\sub1_data_reg_reg[97]  <= 1'b0;
    \\ks1_key_reg_reg[105]  <= 1'b0;
    \\ks1_col_reg[18]  <= 1'b0;
    \\sbox1_ah_reg_reg[0]  <= 1'b0;
    \\sub1_data_reg_reg[81]  <= 1'b0;
    \\sub1_data_reg_reg[49]  <= 1'b0;
    \\sub1_data_reg_reg[113]  <= 1'b0;
    \\sub1_data_reg_reg[33]  <= 1'b0;
    \\sub1_data_reg_reg[57]  <= 1'b0;
    \\sub1_data_reg_reg[89]  <= 1'b0;
    \\sub1_data_reg_reg[25]  <= 1'b0;
    \\ks1_col_reg[26]  <= 1'b0;
    \\sub1_data_reg_reg[121]  <= 1'b0;
    \\ks1_key_reg_reg[106]  <= 1'b0;
    \\ks1_col_reg[2]  <= 1'b0;
    \\sbox1_ah_reg_reg[1]  <= 1'b0;
    \\ks1_col_reg[17]  <= 1'b0;
    \\sbox1_alph_reg[3]  <= 1'b0;
    \\ks1_col_reg[25]  <= 1'b0;
    \\ks1_col_reg[1]  <= 1'b0;
    \\sbox1_ah_reg_reg[3]  <= 1'b0;
    \\ks1_key_reg_reg[28]  <= 1'b0;
    \\ks1_key_reg_reg[27]  <= 1'b0;
    \\ks1_key_reg_reg[29]  <= 1'b0;
    \\ks1_key_reg_reg[30]  <= 1'b0;
    \\ks1_key_reg_reg[24]  <= 1'b0;
    \\ks1_key_reg_reg[31]  <= 1'b0;
    \\ks1_key_reg_reg[25]  <= 1'b0;
    \\ks1_key_reg_reg[26]  <= 1'b0;
    \\ks1_key_reg_reg[60]  <= 1'b0;
    \\ks1_key_reg_reg[2]  <= 1'b0;
    \\ks1_key_reg_reg[3]  <= 1'b0;
    \\ks1_key_reg_reg[4]  <= 1'b0;
    \\ks1_key_reg_reg[5]  <= 1'b0;
    \\ks1_key_reg_reg[6]  <= 1'b0;
    \\ks1_key_reg_reg[0]  <= 1'b0;
    \\ks1_key_reg_reg[1]  <= 1'b0;
    \\ks1_key_reg_reg[23]  <= 1'b0;
    \\ks1_key_reg_reg[7]  <= 1'b0;
    \\ks1_key_reg_reg[61]  <= 1'b0;
    \\ks1_key_reg_reg[59]  <= 1'b0;
    \\ks1_key_reg_reg[17]  <= 1'b0;
    \\ks1_key_reg_reg[16]  <= 1'b0;
    \\ks1_key_reg_reg[19]  <= 1'b0;
    \\ks1_key_reg_reg[18]  <= 1'b0;
    \\ks1_key_reg_reg[21]  <= 1'b0;
    \\ks1_key_reg_reg[22]  <= 1'b0;
    \\ks1_key_reg_reg[20]  <= 1'b0;
    \\ks1_key_reg_reg[57]  <= 1'b0;
    \\ks1_key_reg_reg[58]  <= 1'b0;
    \\ks1_key_reg_reg[63]  <= 1'b0;
    \\ks1_key_reg_reg[62]  <= 1'b0;
    \\ks1_key_reg_reg[56]  <= 1'b0;
    \\ks1_key_reg_reg[92]  <= 1'b0;
    \\ks1_key_reg_reg[32]  <= 1'b0;
    \\ks1_key_reg_reg[33]  <= 1'b0;
    \\ks1_key_reg_reg[34]  <= 1'b0;
    \\ks1_key_reg_reg[35]  <= 1'b0;
    \\ks1_key_reg_reg[36]  <= 1'b0;
    \\ks1_key_reg_reg[38]  <= 1'b0;
    \\ks1_key_reg_reg[39]  <= 1'b0;
    \\ks1_key_reg_reg[55]  <= 1'b0;
    \\ks1_key_reg_reg[37]  <= 1'b0;
    \\ks1_key_reg_reg[91]  <= 1'b0;
    \\ks1_key_reg_reg[93]  <= 1'b0;
    \\ks1_key_reg_reg[49]  <= 1'b0;
    \\ks1_key_reg_reg[50]  <= 1'b0;
    \\ks1_key_reg_reg[51]  <= 1'b0;
    \\ks1_key_reg_reg[52]  <= 1'b0;
    \\ks1_key_reg_reg[54]  <= 1'b0;
    \\ks1_key_reg_reg[48]  <= 1'b0;
    \\ks1_key_reg_reg[53]  <= 1'b0;
    \\ks1_key_reg_reg[90]  <= 1'b0;
    \\ks1_key_reg_reg[88]  <= 1'b0;
    \\ks1_key_reg_reg[94]  <= 1'b0;
    \\ks1_key_reg_reg[95]  <= 1'b0;
    \\ks1_key_reg_reg[89]  <= 1'b0;
    \\ks1_key_reg_reg[69]  <= 1'b0;
    \\addroundkey_data_reg_reg[60]  <= 1'b0;
    \\addroundkey_data_reg_reg[111]  <= 1'b0;
    \\addroundkey_data_reg_reg[63]  <= 1'b0;
    \\addroundkey_data_reg_reg[6]  <= 1'b0;
    \\addroundkey_data_reg_reg[76]  <= 1'b0;
    \\addroundkey_data_reg_reg[25]  <= 1'b0;
    \\addroundkey_data_reg_reg[77]  <= 1'b0;
    \\addroundkey_data_reg_reg[78]  <= 1'b0;
    \\addroundkey_data_reg_reg[79]  <= 1'b0;
    \\addroundkey_data_reg_reg[26]  <= 1'b0;
    \\addroundkey_data_reg_reg[29]  <= 1'b0;
    \\addroundkey_data_reg_reg[8]  <= 1'b0;
    \\addroundkey_data_reg_reg[105]  <= 1'b0;
    \\addroundkey_data_reg_reg[0]  <= 1'b0;
    \\addroundkey_data_reg_reg[106]  <= 1'b0;
    \\addroundkey_data_reg_reg[107]  <= 1'b0;
    \\addroundkey_data_reg_reg[122]  <= 1'b0;
    \\addroundkey_data_reg_reg[3]  <= 1'b0;
    \\addroundkey_data_reg_reg[41]  <= 1'b0;
    \\addroundkey_data_reg_reg[123]  <= 1'b0;
    \\addroundkey_data_reg_reg[42]  <= 1'b0;
    \\addroundkey_data_reg_reg[43]  <= 1'b0;
    \\addroundkey_data_reg_reg[44]  <= 1'b0;
    \\addroundkey_data_reg_reg[108]  <= 1'b0;
    \\addroundkey_data_reg_reg[125]  <= 1'b0;
    \\addroundkey_data_reg_reg[46]  <= 1'b0;
    \\addroundkey_data_reg_reg[47]  <= 1'b0;
    \\addroundkey_data_reg_reg[126]  <= 1'b0;
    \\addroundkey_data_reg_reg[127]  <= 1'b0;
    \\addroundkey_data_reg_reg[10]  <= 1'b0;
    \\addroundkey_data_reg_reg[13]  <= 1'b0;
    \\addroundkey_data_reg_reg[110]  <= 1'b0;
    \\addroundkey_data_reg_reg[58]  <= 1'b0;
    \\addroundkey_data_reg_reg[57]  <= 1'b0;
    \\addroundkey_data_reg_reg[59]  <= 1'b0;
    \\ks1_key_reg_reg[124]  <= 1'b0;
    \\ks1_key_reg_reg[64]  <= 1'b0;
    \\ks1_key_reg_reg[65]  <= 1'b0;
    \\ks1_key_reg_reg[67]  <= 1'b0;
    \\ks1_key_reg_reg[66]  <= 1'b0;
    \\ks1_key_reg_reg[68]  <= 1'b0;
    \\ks1_key_reg_reg[70]  <= 1'b0;
    \\ks1_key_reg_reg[71]  <= 1'b0;
    \\ks1_key_reg_reg[87]  <= 1'b0;
    \\addroundkey_data_reg_reg[5]  <= 1'b0;
    \\ks1_key_reg_reg[81]  <= 1'b0;
    \\addroundkey_data_reg_reg[40]  <= 1'b0;
    \\addroundkey_data_reg_reg[124]  <= 1'b0;
    \\addroundkey_data_reg_reg[61]  <= 1'b0;
    \\addroundkey_data_reg_reg[62]  <= 1'b0;
    \\addroundkey_data_reg_reg[1]  <= 1'b0;
    \\addroundkey_data_reg_reg[73]  <= 1'b0;
    \\addroundkey_data_reg_reg[74]  <= 1'b0;
    \\addroundkey_data_reg_reg[24]  <= 1'b0;
    \\addroundkey_data_reg_reg[72]  <= 1'b0;
    \\addroundkey_data_reg_reg[7]  <= 1'b0;
    \\addroundkey_data_reg_reg[28]  <= 1'b0;
    \\addroundkey_data_reg_reg[104]  <= 1'b0;
    \\addroundkey_data_reg_reg[30]  <= 1'b0;
    \\addroundkey_data_reg_reg[2]  <= 1'b0;
    \\addroundkey_data_reg_reg[31]  <= 1'b0;
    \\addroundkey_data_reg_reg[90]  <= 1'b0;
    \\addroundkey_data_reg_reg[91]  <= 1'b0;
    \\addroundkey_data_reg_reg[92]  <= 1'b0;
    \\addroundkey_data_reg_reg[34]  <= 1'b0;
    \\addroundkey_data_reg_reg[93]  <= 1'b0;
    \\addroundkey_data_reg_reg[11]  <= 1'b0;
    \\addroundkey_data_reg_reg[94]  <= 1'b0;
    \\addroundkey_data_reg_reg[95]  <= 1'b0;
    \\addroundkey_data_reg_reg[120]  <= 1'b0;
    \\addroundkey_data_reg_reg[9]  <= 1'b0;
    \\addroundkey_data_reg_reg[121]  <= 1'b0;
    \\addroundkey_data_reg_reg[45]  <= 1'b0;
    \\addroundkey_data_reg_reg[4]  <= 1'b0;
    \\addroundkey_data_reg_reg[12]  <= 1'b0;
    \\addroundkey_data_reg_reg[109]  <= 1'b0;
    \\addroundkey_data_reg_reg[14]  <= 1'b0;
    \\addroundkey_data_reg_reg[56]  <= 1'b0;
    \\addroundkey_data_reg_reg[15]  <= 1'b0;
    \\ks1_key_reg_reg[125]  <= 1'b0;
    \\ks1_key_reg_reg[123]  <= 1'b0;
    \\ks1_key_reg_reg[80]  <= 1'b0;
    \\ks1_key_reg_reg[83]  <= 1'b0;
    \\ks1_key_reg_reg[84]  <= 1'b0;
    \\ks1_key_reg_reg[85]  <= 1'b0;
    \\ks1_key_reg_reg[82]  <= 1'b0;
    \\ks1_key_reg_reg[86]  <= 1'b0;
    \\addroundkey_data_reg_reg[27]  <= 1'b0;
    \\addroundkey_data_reg_reg[75]  <= 1'b0;
    \\addroundkey_data_reg_reg[100]  <= 1'b0;
    \\addroundkey_data_reg_reg[33]  <= 1'b0;
    \\addroundkey_data_reg_reg[103]  <= 1'b0;
    \\addroundkey_data_reg_reg[98]  <= 1'b0;
    \\addroundkey_data_reg_reg[35]  <= 1'b0;
    \\mix1_data_reg_reg[100]  <= 1'b0;
    \\mix1_data_reg_reg[108]  <= 1'b0;
    \\mix1_data_reg_reg[116]  <= 1'b0;
    \\mix1_data_reg_reg[124]  <= 1'b0;
    \\addroundkey_data_reg_reg[101]  <= 1'b0;
    \\addroundkey_data_reg_reg[112]  <= 1'b0;
    \\addroundkey_data_reg_reg[64]  <= 1'b0;
    \\addroundkey_data_reg_reg[65]  <= 1'b0;
    \\addroundkey_data_reg_reg[20]  <= 1'b0;
    \\addroundkey_data_reg_reg[66]  <= 1'b0;
    \\addroundkey_data_reg_reg[67]  <= 1'b0;
    \\addroundkey_data_reg_reg[21]  <= 1'b0;
    \\addroundkey_data_reg_reg[69]  <= 1'b0;
    \\addroundkey_data_reg_reg[22]  <= 1'b0;
    \\addroundkey_data_reg_reg[70]  <= 1'b0;
    \\addroundkey_data_reg_reg[102]  <= 1'b0;
    \\addroundkey_data_reg_reg[23]  <= 1'b0;
    \\addroundkey_data_reg_reg[115]  <= 1'b0;
    \\addroundkey_data_reg_reg[116]  <= 1'b0;
    \\addroundkey_data_reg_reg[80]  <= 1'b0;
    \\addroundkey_data_reg_reg[81]  <= 1'b0;
    \\addroundkey_data_reg_reg[83]  <= 1'b0;
    \\addroundkey_data_reg_reg[85]  <= 1'b0;
    \\addroundkey_data_reg_reg[86]  <= 1'b0;
    \\addroundkey_data_reg_reg[84]  <= 1'b0;
    \\addroundkey_data_reg_reg[87]  <= 1'b0;
    \\addroundkey_data_reg_reg[88]  <= 1'b0;
    \\addroundkey_data_reg_reg[32]  <= 1'b0;
    \\addroundkey_data_reg_reg[119]  <= 1'b0;
    \\addroundkey_data_reg_reg[96]  <= 1'b0;
    \\addroundkey_data_reg_reg[97]  <= 1'b0;
    \\addroundkey_data_reg_reg[36]  <= 1'b0;
    \\addroundkey_data_reg_reg[99]  <= 1'b0;
    \\addroundkey_data_reg_reg[37]  <= 1'b0;
    \\addroundkey_data_reg_reg[38]  <= 1'b0;
    \\addroundkey_data_reg_reg[39]  <= 1'b0;
    \\addroundkey_data_reg_reg[49]  <= 1'b0;
    \\addroundkey_data_reg_reg[52]  <= 1'b0;
    \\addroundkey_data_reg_reg[55]  <= 1'b0;
    \\addroundkey_data_reg_reg[17]  <= 1'b0;
    \\ks1_key_reg_reg[120]  <= 1'b0;
    \\ks1_key_reg_reg[121]  <= 1'b0;
    \\ks1_key_reg_reg[127]  <= 1'b0;
    \\addroundkey_round_reg[0]  <= 1'b0;
    \\addroundkey_data_reg_reg[118]  <= 1'b0;
    \\addroundkey_data_reg_reg[89]  <= 1'b0;
    \\addroundkey_data_reg_reg[117]  <= 1'b0;
    \\ks1_key_reg_reg[126]  <= 1'b0;
    \\addroundkey_data_reg_reg[82]  <= 1'b0;
    \\ks1_key_reg_reg[122]  <= 1'b0;
    \\addroundkey_data_reg_reg[114]  <= 1'b0;
    \\addroundkey_data_reg_reg[54]  <= 1'b0;
    \\addroundkey_data_reg_reg[71]  <= 1'b0;
    \\addroundkey_data_reg_reg[16]  <= 1'b0;
    \\addroundkey_data_reg_reg[68]  <= 1'b0;
    \\addroundkey_data_reg_reg[53]  <= 1'b0;
    \\addroundkey_data_reg_reg[113]  <= 1'b0;
    \\addroundkey_data_reg_reg[19]  <= 1'b0;
    \\addroundkey_data_reg_reg[51]  <= 1'b0;
    \\addroundkey_data_reg_reg[50]  <= 1'b0;
    \\addroundkey_data_reg_reg[18]  <= 1'b0;
    \\addroundkey_data_reg_reg[48]  <= 1'b0;
    \\ks1_key_reg_reg[97]  <= 1'b0;
    \\mix1_data_reg_reg[107]  <= 1'b0;
    \\mix1_data_reg_reg[115]  <= 1'b0;
    \\mix1_data_reg_reg[99]  <= 1'b0;
    \\ks1_key_reg_reg[96]  <= 1'b0;
    \\ks1_key_reg_reg[98]  <= 1'b0;
    \\ks1_key_reg_reg[100]  <= 1'b0;
    \\ks1_key_reg_reg[101]  <= 1'b0;
    \\ks1_key_reg_reg[102]  <= 1'b0;
    \\ks1_key_reg_reg[103]  <= 1'b0;
    \\ks1_key_reg_reg[119]  <= 1'b0;
    \\mix1_data_reg_reg[123]  <= 1'b0;
    \\ks1_key_reg_reg[113]  <= 1'b0;
    \\mix1_data_reg_reg[36]  <= 1'b0;
    \\mix1_data_reg_reg[44]  <= 1'b0;
    \\mix1_data_reg_reg[60]  <= 1'b0;
    \\mix1_data_reg_reg[68]  <= 1'b0;
    \\mix1_data_reg_reg[52]  <= 1'b0;
    \\mix1_data_reg_reg[84]  <= 1'b0;
    \\mix1_data_reg_reg[76]  <= 1'b0;
    \\mix1_data_reg_reg[92]  <= 1'b0;
    \\ks1_key_reg_reg[112]  <= 1'b0;
    \\ks1_key_reg_reg[115]  <= 1'b0;
    \\ks1_key_reg_reg[116]  <= 1'b0;
    \\ks1_key_reg_reg[114]  <= 1'b0;
    \\ks1_key_reg_reg[118]  <= 1'b0;
    addroundkey_ready_o_reg <= 1'b0;
    \\ks1_key_reg_reg[117]  <= 1'b0;
    \\ks1_key_reg_reg[99]  <= 1'b0;
    \\mix1_data_reg_reg[105]  <= 1'b0;
    \\mix1_data_reg_reg[106]  <= 1'b0;
    \\mix1_data_reg_reg[113]  <= 1'b0;
    \\mix1_data_reg_reg[114]  <= 1'b0;
    \\mix1_data_reg_reg[121]  <= 1'b0;
    \\mix1_data_reg_reg[122]  <= 1'b0;
    \\mix1_data_reg_reg[35]  <= 1'b0;
    \\mix1_data_reg_reg[43]  <= 1'b0;
    \\mix1_data_reg_reg[51]  <= 1'b0;
    \\mix1_data_reg_reg[59]  <= 1'b0;
    \\mix1_data_reg_reg[67]  <= 1'b0;
    \\mix1_data_reg_reg[75]  <= 1'b0;
    \\mix1_data_reg_reg[97]  <= 1'b0;
    \\mix1_data_reg_reg[98]  <= 1'b0;
    \\mix1_data_reg_reg[91]  <= 1'b0;
    \\mix1_data_reg_reg[83]  <= 1'b0;
    \\mix1_data_reg_reg[120]  <= 1'b0;
    \\mix1_data_reg_reg[117]  <= 1'b0;
    \\mix1_data_reg_reg[125]  <= 1'b0;
    \\mix1_data_reg_reg[118]  <= 1'b0;
    \\mix1_data_reg_reg[104]  <= 1'b0;
    \\mix1_data_reg_reg[112]  <= 1'b0;
    \\mix1_data_reg_reg[96]  <= 1'b0;
    \\mix1_data_reg_reg[126]  <= 1'b0;
    \\mix1_data_reg_reg[110]  <= 1'b0;
    \\mix1_data_reg_reg[102]  <= 1'b0;
    \\mix1_data_reg_reg[109]  <= 1'b0;
    \\mix1_data_reg_reg[101]  <= 1'b0;
    \\mix1_data_o_reg_reg[12]  <= 1'b0;
    \\mix1_data_o_reg_reg[20]  <= 1'b0;
    \\mix1_data_o_reg_reg[28]  <= 1'b0;
    \\mix1_data_o_reg_reg[4]  <= 1'b0;
    \\mix1_data_reg_reg[33]  <= 1'b0;
    \\mix1_data_reg_reg[34]  <= 1'b0;
    \\mix1_data_reg_reg[42]  <= 1'b0;
    \\mix1_data_reg_reg[41]  <= 1'b0;
    \\mix1_data_reg_reg[49]  <= 1'b0;
    \\mix1_data_reg_reg[50]  <= 1'b0;
    \\mix1_data_reg_reg[57]  <= 1'b0;
    \\mix1_data_reg_reg[58]  <= 1'b0;
    \\mix1_data_reg_reg[65]  <= 1'b0;
    \\mix1_data_reg_reg[66]  <= 1'b0;
    \\mix1_data_reg_reg[74]  <= 1'b0;
    \\mix1_data_reg_reg[73]  <= 1'b0;
    \\mix1_data_reg_reg[81]  <= 1'b0;
    \\mix1_data_reg_reg[82]  <= 1'b0;
    \\mix1_data_reg_reg[89]  <= 1'b0;
    \\mix1_data_reg_reg[90]  <= 1'b0;
    \\mix1_data_reg_reg[61]  <= 1'b0;
    \\mix1_data_reg_reg[62]  <= 1'b0;
    \\mix1_data_reg_reg[69]  <= 1'b0;
    \\mix1_data_reg_reg[45]  <= 1'b0;
    \\mix1_data_reg_reg[37]  <= 1'b0;
    \\mix1_data_reg_reg[53]  <= 1'b0;
    \\mix1_data_reg_reg[77]  <= 1'b0;
    \\mix1_data_o_reg_reg[3]  <= 1'b0;
    \\mix1_data_reg_reg[38]  <= 1'b0;
    \\mix1_data_reg_reg[46]  <= 1'b0;
    \\mix1_data_reg_reg[54]  <= 1'b0;
    \\mix1_data_reg_reg[70]  <= 1'b0;
    \\mix1_data_reg_reg[78]  <= 1'b0;
    \\mix1_data_reg_reg[86]  <= 1'b0;
    \\mix1_data_reg_reg[94]  <= 1'b0;
    \\mix1_data_reg_reg[32]  <= 1'b0;
    \\mix1_data_reg_reg[48]  <= 1'b0;
    \\mix1_data_reg_reg[56]  <= 1'b0;
    \\mix1_data_reg_reg[64]  <= 1'b0;
    \\mix1_data_reg_reg[88]  <= 1'b0;
    \\mix1_data_reg_reg[80]  <= 1'b0;
    \\mix1_data_reg_reg[72]  <= 1'b0;
    \\mix1_data_reg_reg[40]  <= 1'b0;
    \\mix1_data_o_reg_reg[27]  <= 1'b0;
    \\mix1_data_o_reg_reg[11]  <= 1'b0;
    \\mix1_data_o_reg_reg[19]  <= 1'b0;
    \\mix1_data_reg_reg[85]  <= 1'b0;
    \\mix1_data_reg_reg[93]  <= 1'b0;
    \\mix1_data_reg_reg[103]  <= 1'b0;
    \\mix1_data_reg_reg[111]  <= 1'b0;
    \\mix1_data_reg_reg[127]  <= 1'b0;
    \\mix1_data_reg_reg[119]  <= 1'b0;
    \\mix1_data_o_reg_reg[17]  <= 1'b0;
    \\mix1_data_o_reg_reg[18]  <= 1'b0;
    \\mix1_data_o_reg_reg[1]  <= 1'b0;
    \\mix1_data_o_reg_reg[25]  <= 1'b0;
    \\mix1_data_o_reg_reg[26]  <= 1'b0;
    \\mix1_data_o_reg_reg[9]  <= 1'b0;
    \\mix1_data_o_reg_reg[2]  <= 1'b0;
    \\mix1_data_o_reg_reg[10]  <= 1'b0;
    \\mix1_data_reg_reg[79]  <= 1'b0;
    \\mix1_data_o_reg_reg[8]  <= 1'b0;
    \\mix1_data_reg_reg[55]  <= 1'b0;
    \\mix1_data_reg_reg[71]  <= 1'b0;
    \\mix1_data_o_reg_reg[13]  <= 1'b0;
    \\mix1_data_o_reg_reg[21]  <= 1'b0;
    \\mix1_data_reg_reg[63]  <= 1'b0;
    \\mix1_data_o_reg_reg[22]  <= 1'b0;
    \\mix1_data_o_reg_reg[30]  <= 1'b0;
    \\mix1_data_o_reg_reg[16]  <= 1'b0;
    \\mix1_data_reg_reg[47]  <= 1'b0;
    \\mix1_data_reg_reg[39]  <= 1'b0;
    \\mix1_data_o_reg_reg[6]  <= 1'b0;
    \\mix1_data_o_reg_reg[14]  <= 1'b0;
    \\mix1_data_o_reg_reg[0]  <= 1'b0;
    \\mix1_data_o_reg_reg[24]  <= 1'b0;
    \\mix1_data_reg_reg[95]  <= 1'b0;
    \\mix1_data_o_reg_reg[29]  <= 1'b0;
    \\mix1_data_o_reg_reg[5]  <= 1'b0;
    \\mix1_data_reg_reg[87]  <= 1'b0;
    \\mix1_data_o_reg_reg[7]  <= 1'b0;
    \\mix1_data_o_reg_reg[23]  <= 1'b0;
    \\mix1_data_o_reg_reg[31]  <= 1'b0;
    \\mix1_data_o_reg_reg[15]  <= 1'b0;
    \\addroundkey_round_reg[1]  <= 1'b0;
    \\addroundkey_round_reg[3]  <= 1'b0;
    \\addroundkey_round_reg[2]  <= 1'b0;
    \\ks1_state_reg[0]  <= 1'b0;
    \\ks1_state_reg[2]  <= 1'b0;
    \\round_reg[1]  <= 1'b0;
    \\round_reg[2]  <= 1'b0;
    \\round_reg[0]  <= 1'b0;
    \\round_reg[3]  <= 1'b0;
    addroundkey_start_i_reg <= 1'b0;
    \\mix1_state_reg[0]  <= 1'b0;
    \\mix1_state_reg[1]  <= 1'b0;
    state_reg <= 1'b0;
    \\sub1_state_reg[0]  <= 1'b0;
    ready_o_reg <= 1'b0;
    \\sub1_state_reg[3]  <= 1'b0;
    \\sub1_state_reg[2]  <= 1'b0;
    \\sub1_state_reg[1]  <= 1'b0;
    \\sub1_state_reg[4]  <= 1'b0;
    \\mix1_data_o_reg_reg[104]  <= 1'b0;
    \\mix1_data_o_reg_reg[102]  <= 1'b0;
    \\mix1_data_o_reg_reg[105]  <= 1'b0;
    \\mix1_data_o_reg_reg[108]  <= 1'b0;
    \\mix1_data_o_reg_reg[110]  <= 1'b0;
    \\mix1_data_o_reg_reg[112]  <= 1'b0;
    \\mix1_data_o_reg_reg[45]  <= 1'b0;
    \\mix1_data_o_reg_reg[67]  <= 1'b0;
    \\mix1_data_o_reg_reg[70]  <= 1'b0;
    \\mix1_data_o_reg_reg[85]  <= 1'b0;
    \\mix1_data_o_reg_reg[98]  <= 1'b0;
    \\mix1_data_o_reg_reg[82]  <= 1'b0;
    \\mix1_data_o_reg_reg[99]  <= 1'b0;
    \\mix1_data_o_reg_reg[72]  <= 1'b0;
    \\mix1_data_o_reg_reg[48]  <= 1'b0;
    \\mix1_data_o_reg_reg[91]  <= 1'b0;
    \\mix1_data_o_reg_reg[69]  <= 1'b0;
    \\mix1_data_o_reg_reg[57]  <= 1'b0;
    \\mix1_data_o_reg_reg[33]  <= 1'b0;
    \\mix1_data_o_reg_reg[65]  <= 1'b0;
    \\mix1_data_o_reg_reg[71]  <= 1'b0;
    \\mix1_data_o_reg_reg[93]  <= 1'b0;
    \\mix1_data_o_reg_reg[106]  <= 1'b0;
    \\mix1_data_o_reg_reg[77]  <= 1'b0;
    \\mix1_data_o_reg_reg[78]  <= 1'b0;
    \\mix1_data_o_reg_reg[122]  <= 1'b0;
    \\mix1_data_o_reg_reg[64]  <= 1'b0;
    \\mix1_data_o_reg_reg[49]  <= 1'b0;
    \\mix1_data_o_reg_reg[116]  <= 1'b0;
    \\mix1_data_o_reg_reg[86]  <= 1'b0;
    \\mix1_data_o_reg_reg[88]  <= 1'b0;
    \\mix1_data_o_reg_reg[89]  <= 1'b0;
    \\mix1_data_o_reg_reg[126]  <= 1'b0;
    \\mix1_data_o_reg_reg[90]  <= 1'b0;
    \\mix1_data_o_reg_reg[74]  <= 1'b0;
    \\mix1_data_o_reg_reg[56]  <= 1'b0;
    \\mix1_data_o_reg_reg[47]  <= 1'b0;
    \\mix1_data_o_reg_reg[97]  <= 1'b0;
    \\mix1_data_o_reg_reg[43]  <= 1'b0;
    \\mix1_data_o_reg_reg[76]  <= 1'b0;
    \\mix1_data_o_reg_reg[37]  <= 1'b0;
    \\mix1_data_o_reg_reg[84]  <= 1'b0;
    \\mix1_data_o_reg_reg[103]  <= 1'b0;
    \\mix1_data_o_reg_reg[109]  <= 1'b0;
    \\mix1_data_o_reg_reg[53]  <= 1'b0;
    \\mix1_data_o_reg_reg[119]  <= 1'b0;
    \\mix1_data_o_reg_reg[125]  <= 1'b0;
    \\mix1_data_o_reg_reg[36]  <= 1'b0;
    \\mix1_data_o_reg_reg[39]  <= 1'b0;
    \\mix1_data_o_reg_reg[55]  <= 1'b0;
    \\mix1_data_o_reg_reg[62]  <= 1'b0;
    \\mix1_data_o_reg_reg[96]  <= 1'b0;
    \\mix1_data_o_reg_reg[115]  <= 1'b0;
    \\mix1_data_o_reg_reg[46]  <= 1'b0;
    \\mix1_data_o_reg_reg[80]  <= 1'b0;
    \\mix1_data_o_reg_reg[123]  <= 1'b0;
    \\mix1_data_o_reg_reg[83]  <= 1'b0;
    \\mix1_data_o_reg_reg[58]  <= 1'b0;
    \\mix1_data_o_reg_reg[68]  <= 1'b0;
    \\mix1_data_o_reg_reg[101]  <= 1'b0;
    \\mix1_data_o_reg_reg[118]  <= 1'b0;
    \\mix1_data_o_reg_reg[52]  <= 1'b0;
    \\mix1_data_o_reg_reg[59]  <= 1'b0;
    \\mix1_data_o_reg_reg[87]  <= 1'b0;
    \\mix1_data_o_reg_reg[51]  <= 1'b0;
    \\mix1_data_o_reg_reg[66]  <= 1'b0;
    \\mix1_data_o_reg_reg[81]  <= 1'b0;
    \\mix1_data_o_reg_reg[107]  <= 1'b0;
    \\mix1_data_o_reg_reg[44]  <= 1'b0;
    \\mix1_data_o_reg_reg[42]  <= 1'b0;
    \\mix1_data_o_reg_reg[94]  <= 1'b0;
    \\mix1_data_o_reg_reg[54]  <= 1'b0;
    \\mix1_data_o_reg_reg[50]  <= 1'b0;
    \\mix1_data_o_reg_reg[124]  <= 1'b0;
    \\mix1_data_o_reg_reg[32]  <= 1'b0;
    \\mix1_data_o_reg_reg[75]  <= 1'b0;
    \\mix1_data_o_reg_reg[61]  <= 1'b0;
    \\mix1_data_o_reg_reg[63]  <= 1'b0;
    \\mix1_data_o_reg_reg[120]  <= 1'b0;
    \\mix1_data_o_reg_reg[40]  <= 1'b0;
    \\mix1_data_o_reg_reg[111]  <= 1'b0;
    \\mix1_data_o_reg_reg[34]  <= 1'b0;
    \\mix1_data_o_reg_reg[113]  <= 1'b0;
    \\mix1_data_o_reg_reg[41]  <= 1'b0;
    \\mix1_data_o_reg_reg[121]  <= 1'b0;
    \\mix1_data_o_reg_reg[92]  <= 1'b0;
    \\mix1_data_o_reg_reg[117]  <= 1'b0;
    \\mix1_data_o_reg_reg[60]  <= 1'b0;
    \\mix1_data_o_reg_reg[114]  <= 1'b0;
    \\mix1_data_o_reg_reg[38]  <= 1'b0;
    \\mix1_data_o_reg_reg[73]  <= 1'b0;
    \\mix1_data_o_reg_reg[127]  <= 1'b0;
    \\mix1_data_o_reg_reg[95]  <= 1'b0;
    \\mix1_data_o_reg_reg[79]  <= 1'b0;
    \\mix1_data_o_reg_reg[35]  <= 1'b0;
    \\mix1_data_o_reg_reg[100]  <= 1'b0;
    ks1_ready_o_reg <= 1'b0;
    mix1_ready_o_reg <= 1'b0;
    first_round_reg_reg <= 1'b0;
    \\ks1_state_reg[1]  <= 1'b0;
    sub1_ready_o_reg <= 1'b0;
  end
endmodule


