// Benchmark "testing" written by ABC on Thu Oct  8 22:16:31 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A73  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A73;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1014]_ , \new_[1015]_ ,
    \new_[1018]_ , \new_[1021]_ , \new_[1022]_ , \new_[1023]_ ,
    \new_[1026]_ , \new_[1029]_ , \new_[1030]_ , \new_[1033]_ ,
    \new_[1036]_ , \new_[1037]_ , \new_[1038]_ , \new_[1039]_ ,
    \new_[1042]_ , \new_[1045]_ , \new_[1046]_ , \new_[1049]_ ,
    \new_[1052]_ , \new_[1053]_ , \new_[1054]_ , \new_[1057]_ ,
    \new_[1060]_ , \new_[1061]_ , \new_[1064]_ , \new_[1067]_ ,
    \new_[1068]_ , \new_[1069]_ , \new_[1070]_ , \new_[1071]_ ,
    \new_[1074]_ , \new_[1077]_ , \new_[1078]_ , \new_[1081]_ ,
    \new_[1084]_ , \new_[1085]_ , \new_[1086]_ , \new_[1089]_ ,
    \new_[1092]_ , \new_[1093]_ , \new_[1096]_ , \new_[1099]_ ,
    \new_[1100]_ , \new_[1101]_ , \new_[1102]_ , \new_[1105]_ ,
    \new_[1108]_ , \new_[1109]_ , \new_[1112]_ , \new_[1115]_ ,
    \new_[1116]_ , \new_[1117]_ , \new_[1120]_ , \new_[1123]_ ,
    \new_[1124]_ , \new_[1127]_ , \new_[1130]_ , \new_[1131]_ ,
    \new_[1132]_ , \new_[1133]_ , \new_[1134]_ , \new_[1135]_ ,
    \new_[1139]_ , \new_[1140]_ , \new_[1143]_ , \new_[1146]_ ,
    \new_[1147]_ , \new_[1148]_ , \new_[1151]_ , \new_[1154]_ ,
    \new_[1155]_ , \new_[1158]_ , \new_[1161]_ , \new_[1162]_ ,
    \new_[1163]_ , \new_[1164]_ , \new_[1167]_ , \new_[1170]_ ,
    \new_[1171]_ , \new_[1174]_ , \new_[1177]_ , \new_[1178]_ ,
    \new_[1179]_ , \new_[1182]_ , \new_[1185]_ , \new_[1186]_ ,
    \new_[1189]_ , \new_[1192]_ , \new_[1193]_ , \new_[1194]_ ,
    \new_[1195]_ , \new_[1196]_ , \new_[1199]_ , \new_[1202]_ ,
    \new_[1203]_ , \new_[1206]_ , \new_[1209]_ , \new_[1210]_ ,
    \new_[1211]_ , \new_[1214]_ , \new_[1217]_ , \new_[1218]_ ,
    \new_[1221]_ , \new_[1224]_ , \new_[1225]_ , \new_[1226]_ ,
    \new_[1227]_ , \new_[1230]_ , \new_[1233]_ , \new_[1234]_ ,
    \new_[1237]_ , \new_[1240]_ , \new_[1241]_ , \new_[1242]_ ,
    \new_[1245]_ , \new_[1248]_ , \new_[1249]_ , \new_[1252]_ ,
    \new_[1255]_ , \new_[1256]_ , \new_[1257]_ , \new_[1258]_ ,
    \new_[1259]_ , \new_[1260]_ , \new_[1261]_ , \new_[1265]_ ,
    \new_[1266]_ , \new_[1269]_ , \new_[1272]_ , \new_[1273]_ ,
    \new_[1274]_ , \new_[1277]_ , \new_[1280]_ , \new_[1281]_ ,
    \new_[1284]_ , \new_[1287]_ , \new_[1288]_ , \new_[1289]_ ,
    \new_[1290]_ , \new_[1293]_ , \new_[1296]_ , \new_[1297]_ ,
    \new_[1300]_ , \new_[1303]_ , \new_[1304]_ , \new_[1305]_ ,
    \new_[1308]_ , \new_[1311]_ , \new_[1312]_ , \new_[1315]_ ,
    \new_[1318]_ , \new_[1319]_ , \new_[1320]_ , \new_[1321]_ ,
    \new_[1322]_ , \new_[1325]_ , \new_[1328]_ , \new_[1329]_ ,
    \new_[1332]_ , \new_[1335]_ , \new_[1336]_ , \new_[1337]_ ,
    \new_[1340]_ , \new_[1343]_ , \new_[1344]_ , \new_[1347]_ ,
    \new_[1350]_ , \new_[1351]_ , \new_[1352]_ , \new_[1353]_ ,
    \new_[1356]_ , \new_[1359]_ , \new_[1360]_ , \new_[1363]_ ,
    \new_[1366]_ , \new_[1367]_ , \new_[1368]_ , \new_[1371]_ ,
    \new_[1374]_ , \new_[1375]_ , \new_[1378]_ , \new_[1381]_ ,
    \new_[1382]_ , \new_[1383]_ , \new_[1384]_ , \new_[1385]_ ,
    \new_[1386]_ , \new_[1390]_ , \new_[1391]_ , \new_[1394]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1402]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1409]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1418]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1425]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1433]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1440]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1450]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1457]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1465]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1472]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1481]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1488]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1496]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1503]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1517]_ , \new_[1518]_ , \new_[1521]_ ,
    \new_[1524]_ , \new_[1525]_ , \new_[1526]_ , \new_[1529]_ ,
    \new_[1532]_ , \new_[1533]_ , \new_[1536]_ , \new_[1539]_ ,
    \new_[1540]_ , \new_[1541]_ , \new_[1542]_ , \new_[1545]_ ,
    \new_[1548]_ , \new_[1549]_ , \new_[1552]_ , \new_[1555]_ ,
    \new_[1556]_ , \new_[1557]_ , \new_[1560]_ , \new_[1563]_ ,
    \new_[1564]_ , \new_[1567]_ , \new_[1570]_ , \new_[1571]_ ,
    \new_[1572]_ , \new_[1573]_ , \new_[1574]_ , \new_[1577]_ ,
    \new_[1580]_ , \new_[1581]_ , \new_[1584]_ , \new_[1587]_ ,
    \new_[1588]_ , \new_[1589]_ , \new_[1592]_ , \new_[1595]_ ,
    \new_[1596]_ , \new_[1599]_ , \new_[1602]_ , \new_[1603]_ ,
    \new_[1604]_ , \new_[1605]_ , \new_[1608]_ , \new_[1611]_ ,
    \new_[1612]_ , \new_[1615]_ , \new_[1618]_ , \new_[1619]_ ,
    \new_[1620]_ , \new_[1623]_ , \new_[1626]_ , \new_[1627]_ ,
    \new_[1630]_ , \new_[1633]_ , \new_[1634]_ , \new_[1635]_ ,
    \new_[1636]_ , \new_[1637]_ , \new_[1638]_ , \new_[1642]_ ,
    \new_[1643]_ , \new_[1646]_ , \new_[1649]_ , \new_[1650]_ ,
    \new_[1651]_ , \new_[1654]_ , \new_[1657]_ , \new_[1658]_ ,
    \new_[1661]_ , \new_[1664]_ , \new_[1665]_ , \new_[1666]_ ,
    \new_[1667]_ , \new_[1670]_ , \new_[1673]_ , \new_[1674]_ ,
    \new_[1677]_ , \new_[1680]_ , \new_[1681]_ , \new_[1682]_ ,
    \new_[1685]_ , \new_[1688]_ , \new_[1689]_ , \new_[1692]_ ,
    \new_[1695]_ , \new_[1696]_ , \new_[1697]_ , \new_[1698]_ ,
    \new_[1699]_ , \new_[1702]_ , \new_[1705]_ , \new_[1706]_ ,
    \new_[1709]_ , \new_[1712]_ , \new_[1713]_ , \new_[1714]_ ,
    \new_[1717]_ , \new_[1720]_ , \new_[1721]_ , \new_[1724]_ ,
    \new_[1727]_ , \new_[1728]_ , \new_[1729]_ , \new_[1730]_ ,
    \new_[1733]_ , \new_[1736]_ , \new_[1737]_ , \new_[1740]_ ,
    \new_[1743]_ , \new_[1744]_ , \new_[1745]_ , \new_[1748]_ ,
    \new_[1751]_ , \new_[1752]_ , \new_[1755]_ , \new_[1758]_ ,
    \new_[1759]_ , \new_[1760]_ , \new_[1761]_ , \new_[1762]_ ,
    \new_[1763]_ , \new_[1764]_ , \new_[1768]_ , \new_[1769]_ ,
    \new_[1772]_ , \new_[1775]_ , \new_[1776]_ , \new_[1777]_ ,
    \new_[1780]_ , \new_[1783]_ , \new_[1784]_ , \new_[1787]_ ,
    \new_[1790]_ , \new_[1791]_ , \new_[1792]_ , \new_[1793]_ ,
    \new_[1796]_ , \new_[1799]_ , \new_[1800]_ , \new_[1803]_ ,
    \new_[1806]_ , \new_[1807]_ , \new_[1808]_ , \new_[1811]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1818]_ , \new_[1821]_ ,
    \new_[1822]_ , \new_[1823]_ , \new_[1824]_ , \new_[1825]_ ,
    \new_[1828]_ , \new_[1831]_ , \new_[1832]_ , \new_[1835]_ ,
    \new_[1838]_ , \new_[1839]_ , \new_[1840]_ , \new_[1843]_ ,
    \new_[1846]_ , \new_[1847]_ , \new_[1850]_ , \new_[1853]_ ,
    \new_[1854]_ , \new_[1855]_ , \new_[1856]_ , \new_[1859]_ ,
    \new_[1862]_ , \new_[1863]_ , \new_[1866]_ , \new_[1869]_ ,
    \new_[1870]_ , \new_[1871]_ , \new_[1874]_ , \new_[1877]_ ,
    \new_[1878]_ , \new_[1881]_ , \new_[1884]_ , \new_[1885]_ ,
    \new_[1886]_ , \new_[1887]_ , \new_[1888]_ , \new_[1889]_ ,
    \new_[1892]_ , \new_[1895]_ , \new_[1896]_ , \new_[1899]_ ,
    \new_[1902]_ , \new_[1903]_ , \new_[1904]_ , \new_[1907]_ ,
    \new_[1910]_ , \new_[1911]_ , \new_[1914]_ , \new_[1917]_ ,
    \new_[1918]_ , \new_[1919]_ , \new_[1920]_ , \new_[1923]_ ,
    \new_[1926]_ , \new_[1927]_ , \new_[1930]_ , \new_[1933]_ ,
    \new_[1934]_ , \new_[1935]_ , \new_[1938]_ , \new_[1941]_ ,
    \new_[1942]_ , \new_[1945]_ , \new_[1948]_ , \new_[1949]_ ,
    \new_[1950]_ , \new_[1951]_ , \new_[1952]_ , \new_[1955]_ ,
    \new_[1958]_ , \new_[1959]_ , \new_[1962]_ , \new_[1965]_ ,
    \new_[1966]_ , \new_[1967]_ , \new_[1970]_ , \new_[1973]_ ,
    \new_[1974]_ , \new_[1977]_ , \new_[1980]_ , \new_[1981]_ ,
    \new_[1982]_ , \new_[1983]_ , \new_[1986]_ , \new_[1989]_ ,
    \new_[1990]_ , \new_[1993]_ , \new_[1996]_ , \new_[1997]_ ,
    \new_[1998]_ , \new_[2001]_ , \new_[2004]_ , \new_[2005]_ ,
    \new_[2008]_ , \new_[2011]_ , \new_[2012]_ , \new_[2013]_ ,
    \new_[2014]_ , \new_[2015]_ , \new_[2016]_ , \new_[2017]_ ,
    \new_[2018]_ , \new_[2019]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2027]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2035]_ , \new_[2038]_ , \new_[2039]_ , \new_[2042]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2051]_ , \new_[2054]_ , \new_[2055]_ , \new_[2058]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2066]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2073]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2083]_ , \new_[2086]_ , \new_[2087]_ , \new_[2090]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2098]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2105]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2114]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2121]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2129]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2136]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2148]_ , \new_[2149]_ , \new_[2152]_ , \new_[2155]_ ,
    \new_[2156]_ , \new_[2157]_ , \new_[2160]_ , \new_[2163]_ ,
    \new_[2164]_ , \new_[2167]_ , \new_[2170]_ , \new_[2171]_ ,
    \new_[2172]_ , \new_[2173]_ , \new_[2176]_ , \new_[2179]_ ,
    \new_[2180]_ , \new_[2183]_ , \new_[2186]_ , \new_[2187]_ ,
    \new_[2188]_ , \new_[2191]_ , \new_[2194]_ , \new_[2195]_ ,
    \new_[2198]_ , \new_[2201]_ , \new_[2202]_ , \new_[2203]_ ,
    \new_[2204]_ , \new_[2205]_ , \new_[2208]_ , \new_[2211]_ ,
    \new_[2212]_ , \new_[2215]_ , \new_[2218]_ , \new_[2219]_ ,
    \new_[2220]_ , \new_[2223]_ , \new_[2226]_ , \new_[2227]_ ,
    \new_[2230]_ , \new_[2233]_ , \new_[2234]_ , \new_[2235]_ ,
    \new_[2236]_ , \new_[2239]_ , \new_[2242]_ , \new_[2243]_ ,
    \new_[2246]_ , \new_[2249]_ , \new_[2250]_ , \new_[2251]_ ,
    \new_[2254]_ , \new_[2257]_ , \new_[2258]_ , \new_[2261]_ ,
    \new_[2264]_ , \new_[2265]_ , \new_[2266]_ , \new_[2267]_ ,
    \new_[2268]_ , \new_[2269]_ , \new_[2270]_ , \new_[2274]_ ,
    \new_[2275]_ , \new_[2278]_ , \new_[2281]_ , \new_[2282]_ ,
    \new_[2283]_ , \new_[2286]_ , \new_[2289]_ , \new_[2290]_ ,
    \new_[2293]_ , \new_[2296]_ , \new_[2297]_ , \new_[2298]_ ,
    \new_[2299]_ , \new_[2302]_ , \new_[2305]_ , \new_[2306]_ ,
    \new_[2309]_ , \new_[2312]_ , \new_[2313]_ , \new_[2314]_ ,
    \new_[2317]_ , \new_[2320]_ , \new_[2321]_ , \new_[2324]_ ,
    \new_[2327]_ , \new_[2328]_ , \new_[2329]_ , \new_[2330]_ ,
    \new_[2331]_ , \new_[2334]_ , \new_[2337]_ , \new_[2338]_ ,
    \new_[2341]_ , \new_[2344]_ , \new_[2345]_ , \new_[2346]_ ,
    \new_[2349]_ , \new_[2352]_ , \new_[2353]_ , \new_[2356]_ ,
    \new_[2359]_ , \new_[2360]_ , \new_[2361]_ , \new_[2362]_ ,
    \new_[2365]_ , \new_[2368]_ , \new_[2369]_ , \new_[2372]_ ,
    \new_[2375]_ , \new_[2376]_ , \new_[2377]_ , \new_[2380]_ ,
    \new_[2383]_ , \new_[2384]_ , \new_[2387]_ , \new_[2390]_ ,
    \new_[2391]_ , \new_[2392]_ , \new_[2393]_ , \new_[2394]_ ,
    \new_[2395]_ , \new_[2399]_ , \new_[2400]_ , \new_[2403]_ ,
    \new_[2406]_ , \new_[2407]_ , \new_[2408]_ , \new_[2411]_ ,
    \new_[2414]_ , \new_[2415]_ , \new_[2418]_ , \new_[2421]_ ,
    \new_[2422]_ , \new_[2423]_ , \new_[2424]_ , \new_[2427]_ ,
    \new_[2430]_ , \new_[2431]_ , \new_[2434]_ , \new_[2437]_ ,
    \new_[2438]_ , \new_[2439]_ , \new_[2442]_ , \new_[2445]_ ,
    \new_[2446]_ , \new_[2449]_ , \new_[2452]_ , \new_[2453]_ ,
    \new_[2454]_ , \new_[2455]_ , \new_[2456]_ , \new_[2459]_ ,
    \new_[2462]_ , \new_[2463]_ , \new_[2466]_ , \new_[2469]_ ,
    \new_[2470]_ , \new_[2471]_ , \new_[2474]_ , \new_[2477]_ ,
    \new_[2478]_ , \new_[2481]_ , \new_[2484]_ , \new_[2485]_ ,
    \new_[2486]_ , \new_[2487]_ , \new_[2490]_ , \new_[2493]_ ,
    \new_[2494]_ , \new_[2497]_ , \new_[2500]_ , \new_[2501]_ ,
    \new_[2502]_ , \new_[2505]_ , \new_[2508]_ , \new_[2509]_ ,
    \new_[2512]_ , \new_[2515]_ , \new_[2516]_ , \new_[2517]_ ,
    \new_[2518]_ , \new_[2519]_ , \new_[2520]_ , \new_[2521]_ ,
    \new_[2522]_ , \new_[2526]_ , \new_[2527]_ , \new_[2530]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2538]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2545]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2554]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2561]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2569]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2576]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2586]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2593]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2601]_ , \new_[2604]_ ,
    \new_[2605]_ , \new_[2608]_ , \new_[2611]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2614]_ , \new_[2617]_ , \new_[2620]_ ,
    \new_[2621]_ , \new_[2624]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2632]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2639]_ , \new_[2642]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2646]_ , \new_[2647]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2655]_ , \new_[2658]_ , \new_[2659]_ ,
    \new_[2660]_ , \new_[2663]_ , \new_[2666]_ , \new_[2667]_ ,
    \new_[2670]_ , \new_[2673]_ , \new_[2674]_ , \new_[2675]_ ,
    \new_[2676]_ , \new_[2679]_ , \new_[2682]_ , \new_[2683]_ ,
    \new_[2686]_ , \new_[2689]_ , \new_[2690]_ , \new_[2691]_ ,
    \new_[2694]_ , \new_[2697]_ , \new_[2698]_ , \new_[2701]_ ,
    \new_[2704]_ , \new_[2705]_ , \new_[2706]_ , \new_[2707]_ ,
    \new_[2708]_ , \new_[2711]_ , \new_[2714]_ , \new_[2715]_ ,
    \new_[2718]_ , \new_[2721]_ , \new_[2722]_ , \new_[2723]_ ,
    \new_[2726]_ , \new_[2729]_ , \new_[2730]_ , \new_[2733]_ ,
    \new_[2736]_ , \new_[2737]_ , \new_[2738]_ , \new_[2739]_ ,
    \new_[2742]_ , \new_[2745]_ , \new_[2746]_ , \new_[2749]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2757]_ ,
    \new_[2760]_ , \new_[2761]_ , \new_[2764]_ , \new_[2767]_ ,
    \new_[2768]_ , \new_[2769]_ , \new_[2770]_ , \new_[2771]_ ,
    \new_[2772]_ , \new_[2773]_ , \new_[2777]_ , \new_[2778]_ ,
    \new_[2781]_ , \new_[2784]_ , \new_[2785]_ , \new_[2786]_ ,
    \new_[2789]_ , \new_[2792]_ , \new_[2793]_ , \new_[2796]_ ,
    \new_[2799]_ , \new_[2800]_ , \new_[2801]_ , \new_[2802]_ ,
    \new_[2805]_ , \new_[2808]_ , \new_[2809]_ , \new_[2812]_ ,
    \new_[2815]_ , \new_[2816]_ , \new_[2817]_ , \new_[2820]_ ,
    \new_[2823]_ , \new_[2824]_ , \new_[2827]_ , \new_[2830]_ ,
    \new_[2831]_ , \new_[2832]_ , \new_[2833]_ , \new_[2834]_ ,
    \new_[2837]_ , \new_[2840]_ , \new_[2841]_ , \new_[2844]_ ,
    \new_[2847]_ , \new_[2848]_ , \new_[2849]_ , \new_[2852]_ ,
    \new_[2855]_ , \new_[2856]_ , \new_[2859]_ , \new_[2862]_ ,
    \new_[2863]_ , \new_[2864]_ , \new_[2865]_ , \new_[2868]_ ,
    \new_[2871]_ , \new_[2872]_ , \new_[2875]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2880]_ , \new_[2883]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2890]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2896]_ , \new_[2897]_ , \new_[2898]_ ,
    \new_[2901]_ , \new_[2904]_ , \new_[2905]_ , \new_[2908]_ ,
    \new_[2911]_ , \new_[2912]_ , \new_[2913]_ , \new_[2916]_ ,
    \new_[2919]_ , \new_[2920]_ , \new_[2923]_ , \new_[2926]_ ,
    \new_[2927]_ , \new_[2928]_ , \new_[2929]_ , \new_[2932]_ ,
    \new_[2935]_ , \new_[2936]_ , \new_[2939]_ , \new_[2942]_ ,
    \new_[2943]_ , \new_[2944]_ , \new_[2947]_ , \new_[2950]_ ,
    \new_[2951]_ , \new_[2954]_ , \new_[2957]_ , \new_[2958]_ ,
    \new_[2959]_ , \new_[2960]_ , \new_[2961]_ , \new_[2964]_ ,
    \new_[2967]_ , \new_[2968]_ , \new_[2971]_ , \new_[2974]_ ,
    \new_[2975]_ , \new_[2976]_ , \new_[2979]_ , \new_[2982]_ ,
    \new_[2983]_ , \new_[2986]_ , \new_[2989]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2992]_ , \new_[2995]_ , \new_[2998]_ ,
    \new_[2999]_ , \new_[3002]_ , \new_[3005]_ , \new_[3006]_ ,
    \new_[3007]_ , \new_[3010]_ , \new_[3013]_ , \new_[3014]_ ,
    \new_[3017]_ , \new_[3020]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3024]_ , \new_[3025]_ , \new_[3026]_ ,
    \new_[3027]_ , \new_[3028]_ , \new_[3036]_ , \new_[3040]_ ,
    \new_[3044]_ , \new_[3048]_ , \new_[3052]_ , \new_[3056]_ ,
    \new_[3060]_ , \new_[3064]_ , \new_[3067]_ , \new_[3070]_ ,
    \new_[3073]_ , \new_[3076]_ , \new_[3079]_ , \new_[3082]_ ,
    \new_[3085]_ , \new_[3088]_ , \new_[3091]_ , \new_[3094]_ ,
    \new_[3097]_ , \new_[3100]_ , \new_[3103]_ , \new_[3106]_ ,
    \new_[3109]_ , \new_[3112]_ , \new_[3115]_ , \new_[3118]_ ,
    \new_[3121]_ , \new_[3124]_ , \new_[3127]_ , \new_[3130]_ ,
    \new_[3133]_ , \new_[3136]_ , \new_[3139]_ , \new_[3142]_ ,
    \new_[3145]_ , \new_[3148]_ , \new_[3151]_ , \new_[3154]_ ,
    \new_[3157]_ , \new_[3160]_ , \new_[3163]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3171]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3179]_ , \new_[3183]_ , \new_[3184]_ , \new_[3187]_ ,
    \new_[3191]_ , \new_[3192]_ , \new_[3195]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3203]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3211]_ , \new_[3215]_ , \new_[3216]_ , \new_[3219]_ ,
    \new_[3223]_ , \new_[3224]_ , \new_[3227]_ , \new_[3231]_ ,
    \new_[3232]_ , \new_[3235]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3243]_ , \new_[3247]_ , \new_[3248]_ , \new_[3251]_ ,
    \new_[3255]_ , \new_[3256]_ , \new_[3259]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3267]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3275]_ , \new_[3279]_ , \new_[3280]_ , \new_[3283]_ ,
    \new_[3287]_ , \new_[3288]_ , \new_[3292]_ , \new_[3293]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3302]_ , \new_[3303]_ ,
    \new_[3307]_ , \new_[3308]_ , \new_[3312]_ , \new_[3313]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3327]_ , \new_[3328]_ , \new_[3332]_ , \new_[3333]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3342]_ , \new_[3343]_ ,
    \new_[3347]_ , \new_[3348]_ , \new_[3352]_ , \new_[3353]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3362]_ , \new_[3363]_ ,
    \new_[3367]_ , \new_[3368]_ , \new_[3372]_ , \new_[3373]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3382]_ , \new_[3383]_ ,
    \new_[3387]_ , \new_[3388]_ , \new_[3392]_ , \new_[3393]_ ,
    \new_[3396]_ , \new_[3399]_ , \new_[3400]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3408]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3416]_ , \new_[3417]_ , \new_[3420]_ , \new_[3423]_ ,
    \new_[3424]_ , \new_[3428]_ , \new_[3429]_ , \new_[3432]_ ,
    \new_[3435]_ , \new_[3436]_ , \new_[3440]_ , \new_[3441]_ ,
    \new_[3444]_ , \new_[3447]_ , \new_[3448]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3456]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3464]_ , \new_[3465]_ , \new_[3468]_ , \new_[3471]_ ,
    \new_[3472]_ , \new_[3476]_ , \new_[3477]_ , \new_[3480]_ ,
    \new_[3483]_ , \new_[3484]_ , \new_[3488]_ , \new_[3489]_ ,
    \new_[3492]_ , \new_[3495]_ , \new_[3496]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3504]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3512]_ , \new_[3513]_ , \new_[3516]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3524]_ , \new_[3525]_ , \new_[3528]_ ,
    \new_[3531]_ , \new_[3532]_ , \new_[3536]_ , \new_[3537]_ ,
    \new_[3540]_ , \new_[3543]_ , \new_[3544]_ , \new_[3547]_ ,
    \new_[3550]_ , \new_[3551]_ , \new_[3554]_ , \new_[3557]_ ,
    \new_[3558]_ , \new_[3561]_ , \new_[3564]_ , \new_[3565]_ ,
    \new_[3568]_ , \new_[3571]_ , \new_[3572]_ , \new_[3575]_ ,
    \new_[3578]_ , \new_[3579]_ , \new_[3582]_ , \new_[3585]_ ,
    \new_[3586]_ , \new_[3589]_ , \new_[3592]_ , \new_[3593]_ ,
    \new_[3596]_ , \new_[3599]_ , \new_[3600]_ , \new_[3603]_ ,
    \new_[3606]_ , \new_[3607]_ , \new_[3610]_ , \new_[3613]_ ,
    \new_[3614]_ , \new_[3617]_ , \new_[3620]_ , \new_[3621]_ ,
    \new_[3624]_ , \new_[3627]_ , \new_[3628]_ , \new_[3631]_ ,
    \new_[3634]_ , \new_[3635]_ , \new_[3638]_ , \new_[3641]_ ,
    \new_[3642]_ , \new_[3645]_ , \new_[3648]_ , \new_[3649]_ ,
    \new_[3652]_ , \new_[3655]_ , \new_[3656]_ , \new_[3659]_ ,
    \new_[3662]_ , \new_[3663]_ , \new_[3666]_ , \new_[3669]_ ,
    \new_[3670]_ , \new_[3673]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3680]_ , \new_[3683]_ , \new_[3684]_ , \new_[3687]_ ,
    \new_[3690]_ , \new_[3691]_ , \new_[3694]_ , \new_[3697]_ ,
    \new_[3698]_ , \new_[3701]_ , \new_[3704]_ , \new_[3705]_ ,
    \new_[3708]_ , \new_[3711]_ , \new_[3712]_ , \new_[3715]_ ,
    \new_[3718]_ , \new_[3719]_ , \new_[3722]_ , \new_[3725]_ ,
    \new_[3726]_ , \new_[3729]_ , \new_[3732]_ , \new_[3733]_ ,
    \new_[3736]_ , \new_[3739]_ , \new_[3740]_ , \new_[3743]_ ,
    \new_[3746]_ , \new_[3747]_ , \new_[3750]_ , \new_[3753]_ ,
    \new_[3754]_ , \new_[3757]_ , \new_[3760]_ , \new_[3761]_ ,
    \new_[3764]_ , \new_[3767]_ , \new_[3768]_ , \new_[3771]_ ,
    \new_[3774]_ , \new_[3775]_ , \new_[3778]_ , \new_[3781]_ ,
    \new_[3782]_ , \new_[3785]_ , \new_[3788]_ , \new_[3789]_ ,
    \new_[3792]_ , \new_[3795]_ , \new_[3796]_ , \new_[3799]_ ,
    \new_[3802]_ , \new_[3803]_ , \new_[3806]_ , \new_[3809]_ ,
    \new_[3810]_ , \new_[3813]_ , \new_[3816]_ , \new_[3817]_ ,
    \new_[3820]_ , \new_[3823]_ , \new_[3824]_ , \new_[3827]_ ,
    \new_[3830]_ , \new_[3831]_ , \new_[3834]_ , \new_[3837]_ ,
    \new_[3838]_ , \new_[3841]_ , \new_[3844]_ , \new_[3845]_ ,
    \new_[3848]_ , \new_[3851]_ , \new_[3852]_ , \new_[3855]_ ,
    \new_[3858]_ , \new_[3859]_ , \new_[3862]_ , \new_[3865]_ ,
    \new_[3866]_ , \new_[3869]_ , \new_[3872]_ , \new_[3873]_ ,
    \new_[3876]_ , \new_[3879]_ , \new_[3880]_ , \new_[3883]_ ,
    \new_[3886]_ , \new_[3887]_ , \new_[3890]_ , \new_[3893]_ ,
    \new_[3894]_ , \new_[3897]_ , \new_[3900]_ , \new_[3901]_ ,
    \new_[3904]_ , \new_[3907]_ , \new_[3908]_ , \new_[3911]_ ,
    \new_[3914]_ , \new_[3915]_ , \new_[3918]_ , \new_[3921]_ ,
    \new_[3922]_ , \new_[3925]_ , \new_[3928]_ , \new_[3929]_ ,
    \new_[3932]_ , \new_[3935]_ , \new_[3936]_ , \new_[3939]_ ,
    \new_[3942]_ , \new_[3943]_ , \new_[3946]_ , \new_[3949]_ ,
    \new_[3950]_ , \new_[3953]_ , \new_[3956]_ , \new_[3957]_ ,
    \new_[3960]_ , \new_[3963]_ , \new_[3964]_ , \new_[3967]_ ,
    \new_[3970]_ , \new_[3971]_ , \new_[3974]_ , \new_[3977]_ ,
    \new_[3978]_ , \new_[3981]_ , \new_[3984]_ , \new_[3985]_ ,
    \new_[3988]_ , \new_[3991]_ , \new_[3992]_ , \new_[3995]_ ,
    \new_[3998]_ , \new_[3999]_ , \new_[4002]_ , \new_[4005]_ ,
    \new_[4006]_ , \new_[4009]_ , \new_[4012]_ , \new_[4013]_ ,
    \new_[4016]_ , \new_[4019]_ , \new_[4020]_ , \new_[4023]_ ,
    \new_[4026]_ , \new_[4027]_ , \new_[4030]_ , \new_[4033]_ ,
    \new_[4034]_ , \new_[4037]_ , \new_[4040]_ , \new_[4041]_ ,
    \new_[4044]_ , \new_[4047]_ , \new_[4048]_ , \new_[4051]_ ,
    \new_[4054]_ , \new_[4055]_ , \new_[4058]_ , \new_[4061]_ ,
    \new_[4062]_ , \new_[4065]_ , \new_[4068]_ , \new_[4069]_ ,
    \new_[4072]_ , \new_[4075]_ , \new_[4076]_ , \new_[4079]_ ,
    \new_[4082]_ , \new_[4083]_ , \new_[4086]_ , \new_[4089]_ ,
    \new_[4090]_ , \new_[4093]_ , \new_[4096]_ , \new_[4097]_ ,
    \new_[4100]_ , \new_[4103]_ , \new_[4104]_ , \new_[4107]_ ,
    \new_[4110]_ , \new_[4111]_ , \new_[4114]_ , \new_[4117]_ ,
    \new_[4118]_ , \new_[4121]_ , \new_[4124]_ , \new_[4125]_ ,
    \new_[4128]_ , \new_[4131]_ , \new_[4132]_ , \new_[4135]_ ,
    \new_[4138]_ , \new_[4139]_ , \new_[4142]_ , \new_[4145]_ ,
    \new_[4146]_ , \new_[4149]_ , \new_[4152]_ , \new_[4153]_ ,
    \new_[4156]_ , \new_[4159]_ , \new_[4160]_ , \new_[4163]_ ,
    \new_[4166]_ , \new_[4167]_ , \new_[4170]_ , \new_[4173]_ ,
    \new_[4174]_ , \new_[4177]_ , \new_[4180]_ , \new_[4181]_ ,
    \new_[4184]_ , \new_[4187]_ , \new_[4188]_ , \new_[4191]_ ,
    \new_[4194]_ , \new_[4195]_ , \new_[4198]_ , \new_[4201]_ ,
    \new_[4202]_ , \new_[4205]_ , \new_[4208]_ , \new_[4209]_ ,
    \new_[4212]_ , \new_[4215]_ , \new_[4216]_ , \new_[4219]_ ,
    \new_[4222]_ , \new_[4223]_ , \new_[4226]_ , \new_[4229]_ ,
    \new_[4230]_ , \new_[4233]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4240]_ , \new_[4243]_ , \new_[4244]_ , \new_[4247]_ ,
    \new_[4250]_ , \new_[4251]_ , \new_[4254]_ , \new_[4258]_ ,
    \new_[4259]_ , \new_[4260]_ , \new_[4263]_ , \new_[4266]_ ,
    \new_[4267]_ , \new_[4270]_ , \new_[4274]_ , \new_[4275]_ ,
    \new_[4276]_ , \new_[4279]_ , \new_[4282]_ , \new_[4283]_ ,
    \new_[4286]_ , \new_[4290]_ , \new_[4291]_ , \new_[4292]_ ,
    \new_[4295]_ , \new_[4298]_ , \new_[4299]_ , \new_[4302]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4311]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4318]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4327]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4334]_ , \new_[4338]_ , \new_[4339]_ ,
    \new_[4340]_ , \new_[4343]_ , \new_[4346]_ , \new_[4347]_ ,
    \new_[4350]_ , \new_[4354]_ , \new_[4355]_ , \new_[4356]_ ,
    \new_[4359]_ , \new_[4362]_ , \new_[4363]_ , \new_[4366]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4372]_ , \new_[4375]_ ,
    \new_[4378]_ , \new_[4379]_ , \new_[4382]_ , \new_[4386]_ ,
    \new_[4387]_ , \new_[4388]_ , \new_[4391]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4398]_ , \new_[4402]_ , \new_[4403]_ ,
    \new_[4404]_ , \new_[4407]_ , \new_[4410]_ , \new_[4411]_ ,
    \new_[4414]_ , \new_[4418]_ , \new_[4419]_ , \new_[4420]_ ,
    \new_[4423]_ , \new_[4426]_ , \new_[4427]_ , \new_[4430]_ ,
    \new_[4434]_ , \new_[4435]_ , \new_[4436]_ , \new_[4439]_ ,
    \new_[4442]_ , \new_[4443]_ , \new_[4446]_ , \new_[4450]_ ,
    \new_[4451]_ , \new_[4452]_ , \new_[4455]_ , \new_[4458]_ ,
    \new_[4459]_ , \new_[4462]_ , \new_[4466]_ , \new_[4467]_ ,
    \new_[4468]_ , \new_[4471]_ , \new_[4474]_ , \new_[4475]_ ,
    \new_[4478]_ , \new_[4482]_ , \new_[4483]_ , \new_[4484]_ ,
    \new_[4487]_ , \new_[4490]_ , \new_[4491]_ , \new_[4494]_ ,
    \new_[4498]_ , \new_[4499]_ , \new_[4500]_ , \new_[4503]_ ,
    \new_[4506]_ , \new_[4507]_ , \new_[4510]_ , \new_[4514]_ ,
    \new_[4515]_ , \new_[4516]_ , \new_[4519]_ , \new_[4522]_ ,
    \new_[4523]_ , \new_[4526]_ , \new_[4530]_ , \new_[4531]_ ,
    \new_[4532]_ , \new_[4535]_ , \new_[4538]_ , \new_[4539]_ ,
    \new_[4542]_ , \new_[4546]_ , \new_[4547]_ , \new_[4548]_ ,
    \new_[4551]_ , \new_[4554]_ , \new_[4555]_ , \new_[4558]_ ,
    \new_[4562]_ , \new_[4563]_ , \new_[4564]_ , \new_[4567]_ ,
    \new_[4570]_ , \new_[4571]_ , \new_[4574]_ , \new_[4578]_ ,
    \new_[4579]_ , \new_[4580]_ , \new_[4583]_ , \new_[4586]_ ,
    \new_[4587]_ , \new_[4590]_ , \new_[4594]_ , \new_[4595]_ ,
    \new_[4596]_ , \new_[4599]_ , \new_[4602]_ , \new_[4603]_ ,
    \new_[4606]_ , \new_[4610]_ , \new_[4611]_ , \new_[4612]_ ,
    \new_[4615]_ , \new_[4618]_ , \new_[4619]_ , \new_[4622]_ ,
    \new_[4626]_ , \new_[4627]_ , \new_[4628]_ , \new_[4631]_ ,
    \new_[4634]_ , \new_[4635]_ , \new_[4638]_ , \new_[4642]_ ,
    \new_[4643]_ , \new_[4644]_ , \new_[4647]_ , \new_[4650]_ ,
    \new_[4651]_ , \new_[4654]_ , \new_[4658]_ , \new_[4659]_ ,
    \new_[4660]_ , \new_[4663]_ , \new_[4666]_ , \new_[4667]_ ,
    \new_[4670]_ , \new_[4674]_ , \new_[4675]_ , \new_[4676]_ ,
    \new_[4679]_ , \new_[4682]_ , \new_[4683]_ , \new_[4686]_ ,
    \new_[4690]_ , \new_[4691]_ , \new_[4692]_ , \new_[4695]_ ,
    \new_[4698]_ , \new_[4699]_ , \new_[4702]_ , \new_[4706]_ ,
    \new_[4707]_ , \new_[4708]_ , \new_[4711]_ , \new_[4714]_ ,
    \new_[4715]_ , \new_[4718]_ , \new_[4722]_ , \new_[4723]_ ,
    \new_[4724]_ , \new_[4727]_ , \new_[4730]_ , \new_[4731]_ ,
    \new_[4734]_ , \new_[4738]_ , \new_[4739]_ , \new_[4740]_ ,
    \new_[4743]_ , \new_[4746]_ , \new_[4747]_ , \new_[4750]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4759]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4766]_ , \new_[4770]_ ,
    \new_[4771]_ , \new_[4772]_ , \new_[4775]_ , \new_[4778]_ ,
    \new_[4779]_ , \new_[4782]_ , \new_[4786]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4791]_ , \new_[4794]_ , \new_[4795]_ ,
    \new_[4798]_ , \new_[4802]_ , \new_[4803]_ , \new_[4804]_ ,
    \new_[4807]_ , \new_[4810]_ , \new_[4811]_ , \new_[4814]_ ,
    \new_[4818]_ , \new_[4819]_ , \new_[4820]_ , \new_[4823]_ ,
    \new_[4826]_ , \new_[4827]_ , \new_[4830]_ , \new_[4834]_ ,
    \new_[4835]_ , \new_[4836]_ , \new_[4839]_ , \new_[4842]_ ,
    \new_[4843]_ , \new_[4846]_ , \new_[4850]_ , \new_[4851]_ ,
    \new_[4852]_ , \new_[4855]_ , \new_[4858]_ , \new_[4859]_ ,
    \new_[4862]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4871]_ , \new_[4874]_ , \new_[4875]_ , \new_[4878]_ ,
    \new_[4882]_ , \new_[4883]_ , \new_[4884]_ , \new_[4887]_ ,
    \new_[4890]_ , \new_[4891]_ , \new_[4894]_ , \new_[4898]_ ,
    \new_[4899]_ , \new_[4900]_ , \new_[4903]_ , \new_[4906]_ ,
    \new_[4907]_ , \new_[4910]_ , \new_[4914]_ , \new_[4915]_ ,
    \new_[4916]_ , \new_[4919]_ , \new_[4922]_ , \new_[4923]_ ,
    \new_[4926]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4935]_ , \new_[4938]_ , \new_[4939]_ , \new_[4942]_ ,
    \new_[4946]_ , \new_[4947]_ , \new_[4948]_ , \new_[4951]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4958]_ , \new_[4962]_ ,
    \new_[4963]_ , \new_[4964]_ , \new_[4967]_ , \new_[4970]_ ,
    \new_[4971]_ , \new_[4974]_ , \new_[4978]_ , \new_[4979]_ ,
    \new_[4980]_ , \new_[4983]_ , \new_[4986]_ , \new_[4987]_ ,
    \new_[4990]_ , \new_[4994]_ , \new_[4995]_ , \new_[4996]_ ,
    \new_[4999]_ , \new_[5002]_ , \new_[5003]_ , \new_[5006]_ ,
    \new_[5010]_ , \new_[5011]_ , \new_[5012]_ , \new_[5015]_ ,
    \new_[5018]_ , \new_[5019]_ , \new_[5022]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5031]_ , \new_[5034]_ ,
    \new_[5035]_ , \new_[5038]_ , \new_[5042]_ , \new_[5043]_ ,
    \new_[5044]_ , \new_[5047]_ , \new_[5050]_ , \new_[5051]_ ,
    \new_[5054]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5063]_ , \new_[5066]_ , \new_[5067]_ , \new_[5070]_ ,
    \new_[5074]_ , \new_[5075]_ , \new_[5076]_ , \new_[5079]_ ,
    \new_[5082]_ , \new_[5083]_ , \new_[5086]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5095]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5102]_ , \new_[5106]_ , \new_[5107]_ ,
    \new_[5108]_ , \new_[5111]_ , \new_[5114]_ , \new_[5115]_ ,
    \new_[5118]_ , \new_[5122]_ , \new_[5123]_ , \new_[5124]_ ,
    \new_[5127]_ , \new_[5130]_ , \new_[5131]_ , \new_[5134]_ ,
    \new_[5138]_ , \new_[5139]_ , \new_[5140]_ , \new_[5143]_ ,
    \new_[5146]_ , \new_[5147]_ , \new_[5150]_ , \new_[5154]_ ,
    \new_[5155]_ , \new_[5156]_ , \new_[5159]_ , \new_[5162]_ ,
    \new_[5163]_ , \new_[5166]_ , \new_[5170]_ , \new_[5171]_ ,
    \new_[5172]_ , \new_[5175]_ , \new_[5178]_ , \new_[5179]_ ,
    \new_[5182]_ , \new_[5186]_ , \new_[5187]_ , \new_[5188]_ ,
    \new_[5191]_ , \new_[5194]_ , \new_[5195]_ , \new_[5198]_ ,
    \new_[5202]_ , \new_[5203]_ , \new_[5204]_ , \new_[5207]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5214]_ , \new_[5218]_ ,
    \new_[5219]_ , \new_[5220]_ , \new_[5223]_ , \new_[5226]_ ,
    \new_[5227]_ , \new_[5230]_ , \new_[5234]_ , \new_[5235]_ ,
    \new_[5236]_ , \new_[5239]_ , \new_[5242]_ , \new_[5243]_ ,
    \new_[5246]_ , \new_[5250]_ , \new_[5251]_ , \new_[5252]_ ,
    \new_[5255]_ , \new_[5258]_ , \new_[5259]_ , \new_[5262]_ ,
    \new_[5266]_ , \new_[5267]_ , \new_[5268]_ , \new_[5271]_ ,
    \new_[5274]_ , \new_[5275]_ , \new_[5278]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5287]_ , \new_[5290]_ ,
    \new_[5291]_ , \new_[5294]_ , \new_[5298]_ , \new_[5299]_ ,
    \new_[5300]_ , \new_[5303]_ , \new_[5306]_ , \new_[5307]_ ,
    \new_[5310]_ , \new_[5314]_ , \new_[5315]_ , \new_[5316]_ ,
    \new_[5319]_ , \new_[5322]_ , \new_[5323]_ , \new_[5326]_ ,
    \new_[5330]_ , \new_[5331]_ , \new_[5332]_ , \new_[5335]_ ,
    \new_[5338]_ , \new_[5339]_ , \new_[5342]_ , \new_[5346]_ ,
    \new_[5347]_ , \new_[5348]_ , \new_[5351]_ , \new_[5354]_ ,
    \new_[5355]_ , \new_[5358]_ , \new_[5362]_ , \new_[5363]_ ,
    \new_[5364]_ , \new_[5367]_ , \new_[5370]_ , \new_[5371]_ ,
    \new_[5374]_ , \new_[5378]_ , \new_[5379]_ , \new_[5380]_ ,
    \new_[5383]_ , \new_[5386]_ , \new_[5387]_ , \new_[5390]_ ,
    \new_[5394]_ , \new_[5395]_ , \new_[5396]_ , \new_[5399]_ ,
    \new_[5402]_ , \new_[5403]_ , \new_[5406]_ , \new_[5410]_ ,
    \new_[5411]_ , \new_[5412]_ , \new_[5415]_ , \new_[5418]_ ,
    \new_[5419]_ , \new_[5422]_ , \new_[5426]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5431]_ , \new_[5434]_ , \new_[5435]_ ,
    \new_[5438]_ , \new_[5442]_ , \new_[5443]_ , \new_[5444]_ ,
    \new_[5447]_ , \new_[5450]_ , \new_[5451]_ , \new_[5454]_ ,
    \new_[5458]_ , \new_[5459]_ , \new_[5460]_ , \new_[5463]_ ,
    \new_[5466]_ , \new_[5467]_ , \new_[5470]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5476]_ , \new_[5479]_ , \new_[5482]_ ,
    \new_[5483]_ , \new_[5486]_ , \new_[5490]_ , \new_[5491]_ ,
    \new_[5492]_ , \new_[5495]_ , \new_[5498]_ , \new_[5499]_ ,
    \new_[5502]_ , \new_[5506]_ , \new_[5507]_ , \new_[5508]_ ,
    \new_[5511]_ , \new_[5514]_ , \new_[5515]_ , \new_[5518]_ ,
    \new_[5522]_ , \new_[5523]_ , \new_[5524]_ , \new_[5527]_ ,
    \new_[5530]_ , \new_[5531]_ , \new_[5534]_ , \new_[5538]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5543]_ , \new_[5546]_ ,
    \new_[5547]_ , \new_[5550]_ , \new_[5554]_ , \new_[5555]_ ,
    \new_[5556]_ , \new_[5559]_ , \new_[5562]_ , \new_[5563]_ ,
    \new_[5566]_ , \new_[5570]_ , \new_[5571]_ , \new_[5572]_ ,
    \new_[5575]_ , \new_[5578]_ , \new_[5579]_ , \new_[5582]_ ,
    \new_[5586]_ , \new_[5587]_ , \new_[5588]_ , \new_[5591]_ ,
    \new_[5594]_ , \new_[5595]_ , \new_[5598]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5607]_ , \new_[5610]_ ,
    \new_[5611]_ , \new_[5614]_ , \new_[5618]_ , \new_[5619]_ ,
    \new_[5620]_ , \new_[5623]_ , \new_[5626]_ , \new_[5627]_ ,
    \new_[5630]_ , \new_[5634]_ , \new_[5635]_ , \new_[5636]_ ,
    \new_[5639]_ , \new_[5642]_ , \new_[5643]_ , \new_[5646]_ ,
    \new_[5650]_ , \new_[5651]_ , \new_[5652]_ , \new_[5655]_ ,
    \new_[5658]_ , \new_[5659]_ , \new_[5662]_ , \new_[5666]_ ,
    \new_[5667]_ , \new_[5668]_ , \new_[5671]_ , \new_[5674]_ ,
    \new_[5675]_ , \new_[5678]_ , \new_[5682]_ , \new_[5683]_ ,
    \new_[5684]_ , \new_[5687]_ , \new_[5690]_ , \new_[5691]_ ,
    \new_[5694]_ , \new_[5698]_ , \new_[5699]_ , \new_[5700]_ ,
    \new_[5703]_ , \new_[5706]_ , \new_[5707]_ , \new_[5710]_ ,
    \new_[5714]_ , \new_[5715]_ , \new_[5716]_ , \new_[5719]_ ,
    \new_[5722]_ , \new_[5723]_ , \new_[5726]_ , \new_[5730]_ ,
    \new_[5731]_ , \new_[5732]_ , \new_[5735]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5742]_ , \new_[5746]_ , \new_[5747]_ ,
    \new_[5748]_ , \new_[5751]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5758]_ , \new_[5762]_ , \new_[5763]_ , \new_[5764]_ ,
    \new_[5767]_ , \new_[5770]_ , \new_[5771]_ , \new_[5774]_ ,
    \new_[5778]_ , \new_[5779]_ , \new_[5780]_ , \new_[5783]_ ,
    \new_[5786]_ , \new_[5787]_ , \new_[5790]_ , \new_[5794]_ ,
    \new_[5795]_ , \new_[5796]_ , \new_[5799]_ , \new_[5802]_ ,
    \new_[5803]_ , \new_[5806]_ , \new_[5810]_ , \new_[5811]_ ,
    \new_[5812]_ , \new_[5815]_ , \new_[5818]_ , \new_[5819]_ ,
    \new_[5822]_ , \new_[5826]_ , \new_[5827]_ , \new_[5828]_ ,
    \new_[5831]_ , \new_[5834]_ , \new_[5835]_ , \new_[5838]_ ,
    \new_[5842]_ , \new_[5843]_ , \new_[5844]_ , \new_[5847]_ ,
    \new_[5850]_ , \new_[5851]_ , \new_[5854]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5863]_ , \new_[5866]_ ,
    \new_[5867]_ , \new_[5870]_ , \new_[5874]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5879]_ , \new_[5882]_ , \new_[5883]_ ,
    \new_[5886]_ , \new_[5890]_ , \new_[5891]_ , \new_[5892]_ ,
    \new_[5895]_ , \new_[5898]_ , \new_[5899]_ , \new_[5902]_ ,
    \new_[5906]_ , \new_[5907]_ , \new_[5908]_ , \new_[5911]_ ,
    \new_[5914]_ , \new_[5915]_ , \new_[5918]_ , \new_[5922]_ ,
    \new_[5923]_ , \new_[5924]_ , \new_[5927]_ , \new_[5930]_ ,
    \new_[5931]_ , \new_[5934]_ , \new_[5938]_ , \new_[5939]_ ,
    \new_[5940]_ , \new_[5943]_ , \new_[5946]_ , \new_[5947]_ ,
    \new_[5950]_ , \new_[5954]_ , \new_[5955]_ , \new_[5956]_ ,
    \new_[5959]_ , \new_[5962]_ , \new_[5963]_ , \new_[5966]_ ,
    \new_[5970]_ , \new_[5971]_ , \new_[5972]_ , \new_[5975]_ ,
    \new_[5978]_ , \new_[5979]_ , \new_[5982]_ , \new_[5986]_ ,
    \new_[5987]_ , \new_[5988]_ , \new_[5991]_ , \new_[5994]_ ,
    \new_[5995]_ , \new_[5998]_ , \new_[6002]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6007]_ , \new_[6010]_ , \new_[6011]_ ,
    \new_[6014]_ , \new_[6018]_ , \new_[6019]_ , \new_[6020]_ ,
    \new_[6023]_ , \new_[6026]_ , \new_[6027]_ , \new_[6030]_ ,
    \new_[6034]_ , \new_[6035]_ , \new_[6036]_ , \new_[6039]_ ,
    \new_[6042]_ , \new_[6043]_ , \new_[6046]_ , \new_[6050]_ ,
    \new_[6051]_ , \new_[6052]_ , \new_[6055]_ , \new_[6058]_ ,
    \new_[6059]_ , \new_[6062]_ , \new_[6066]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6071]_ , \new_[6074]_ , \new_[6075]_ ,
    \new_[6078]_ , \new_[6082]_ , \new_[6083]_ , \new_[6084]_ ,
    \new_[6087]_ , \new_[6090]_ , \new_[6091]_ , \new_[6094]_ ,
    \new_[6098]_ , \new_[6099]_ , \new_[6100]_ , \new_[6103]_ ,
    \new_[6106]_ , \new_[6107]_ , \new_[6110]_ , \new_[6114]_ ,
    \new_[6115]_ , \new_[6116]_ , \new_[6119]_ , \new_[6122]_ ,
    \new_[6123]_ , \new_[6126]_ , \new_[6130]_ , \new_[6131]_ ,
    \new_[6132]_ , \new_[6135]_ , \new_[6138]_ , \new_[6139]_ ,
    \new_[6142]_ , \new_[6146]_ , \new_[6147]_ , \new_[6148]_ ,
    \new_[6151]_ , \new_[6154]_ , \new_[6155]_ , \new_[6158]_ ,
    \new_[6162]_ , \new_[6163]_ , \new_[6164]_ , \new_[6167]_ ,
    \new_[6170]_ , \new_[6171]_ , \new_[6174]_ , \new_[6178]_ ,
    \new_[6179]_ , \new_[6180]_ , \new_[6183]_ , \new_[6186]_ ,
    \new_[6187]_ , \new_[6190]_ , \new_[6194]_ , \new_[6195]_ ,
    \new_[6196]_ , \new_[6199]_ , \new_[6203]_ , \new_[6204]_ ,
    \new_[6205]_ , \new_[6208]_ , \new_[6212]_ , \new_[6213]_ ,
    \new_[6214]_ , \new_[6217]_ , \new_[6221]_ , \new_[6222]_ ,
    \new_[6223]_ , \new_[6226]_ , \new_[6230]_ , \new_[6231]_ ,
    \new_[6232]_ , \new_[6235]_ , \new_[6239]_ , \new_[6240]_ ,
    \new_[6241]_ , \new_[6244]_ , \new_[6248]_ , \new_[6249]_ ,
    \new_[6250]_ , \new_[6253]_ , \new_[6257]_ , \new_[6258]_ ,
    \new_[6259]_ , \new_[6262]_ , \new_[6266]_ , \new_[6267]_ ,
    \new_[6268]_ , \new_[6271]_ , \new_[6275]_ , \new_[6276]_ ,
    \new_[6277]_ , \new_[6280]_ , \new_[6284]_ , \new_[6285]_ ,
    \new_[6286]_ , \new_[6289]_ , \new_[6293]_ , \new_[6294]_ ,
    \new_[6295]_ , \new_[6298]_ , \new_[6302]_ , \new_[6303]_ ,
    \new_[6304]_ , \new_[6307]_ , \new_[6311]_ , \new_[6312]_ ,
    \new_[6313]_ , \new_[6316]_ , \new_[6320]_ , \new_[6321]_ ,
    \new_[6322]_ , \new_[6325]_ , \new_[6329]_ , \new_[6330]_ ,
    \new_[6331]_ , \new_[6334]_ , \new_[6338]_ , \new_[6339]_ ,
    \new_[6340]_ , \new_[6343]_ , \new_[6347]_ , \new_[6348]_ ,
    \new_[6349]_ , \new_[6352]_ , \new_[6356]_ , \new_[6357]_ ,
    \new_[6358]_ , \new_[6361]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6367]_ , \new_[6370]_ , \new_[6374]_ , \new_[6375]_ ,
    \new_[6376]_ , \new_[6379]_ , \new_[6383]_ , \new_[6384]_ ,
    \new_[6385]_ , \new_[6388]_ , \new_[6392]_ , \new_[6393]_ ,
    \new_[6394]_ , \new_[6397]_ , \new_[6401]_ , \new_[6402]_ ,
    \new_[6403]_ , \new_[6406]_ , \new_[6410]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6415]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6421]_ , \new_[6424]_ , \new_[6428]_ , \new_[6429]_ ,
    \new_[6430]_ , \new_[6433]_ , \new_[6437]_ , \new_[6438]_ ,
    \new_[6439]_ , \new_[6442]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6451]_ , \new_[6455]_ , \new_[6456]_ ,
    \new_[6457]_ , \new_[6460]_ , \new_[6464]_ , \new_[6465]_ ,
    \new_[6466]_ , \new_[6469]_ , \new_[6473]_ , \new_[6474]_ ,
    \new_[6475]_ , \new_[6478]_ , \new_[6482]_ , \new_[6483]_ ,
    \new_[6484]_ , \new_[6487]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6493]_ , \new_[6496]_ , \new_[6500]_ , \new_[6501]_ ,
    \new_[6502]_ , \new_[6505]_ , \new_[6509]_ , \new_[6510]_ ,
    \new_[6511]_ , \new_[6514]_ , \new_[6518]_ , \new_[6519]_ ,
    \new_[6520]_ , \new_[6523]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6532]_ , \new_[6536]_ , \new_[6537]_ ,
    \new_[6538]_ , \new_[6541]_ , \new_[6545]_ , \new_[6546]_ ,
    \new_[6547]_ , \new_[6550]_ , \new_[6554]_ , \new_[6555]_ ,
    \new_[6556]_ , \new_[6559]_ , \new_[6563]_ , \new_[6564]_ ,
    \new_[6565]_ , \new_[6568]_ , \new_[6572]_ , \new_[6573]_ ,
    \new_[6574]_ , \new_[6577]_ , \new_[6581]_ , \new_[6582]_ ,
    \new_[6583]_ , \new_[6586]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6592]_ , \new_[6595]_ , \new_[6599]_ , \new_[6600]_ ,
    \new_[6601]_ , \new_[6604]_ , \new_[6608]_ , \new_[6609]_ ,
    \new_[6610]_ , \new_[6613]_ , \new_[6617]_ , \new_[6618]_ ,
    \new_[6619]_ , \new_[6622]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6628]_ , \new_[6631]_ , \new_[6635]_ , \new_[6636]_ ,
    \new_[6637]_ , \new_[6640]_ , \new_[6644]_ , \new_[6645]_ ,
    \new_[6646]_ , \new_[6649]_ , \new_[6653]_ , \new_[6654]_ ,
    \new_[6655]_ , \new_[6658]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6664]_ , \new_[6667]_ , \new_[6671]_ , \new_[6672]_ ,
    \new_[6673]_ , \new_[6676]_ , \new_[6680]_ , \new_[6681]_ ,
    \new_[6682]_ , \new_[6685]_ , \new_[6689]_ , \new_[6690]_ ,
    \new_[6691]_ , \new_[6694]_ , \new_[6698]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6703]_ , \new_[6707]_ , \new_[6708]_ ,
    \new_[6709]_ , \new_[6712]_ , \new_[6716]_ , \new_[6717]_ ,
    \new_[6718]_ , \new_[6721]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6727]_ , \new_[6730]_ , \new_[6734]_ , \new_[6735]_ ,
    \new_[6736]_ , \new_[6739]_ , \new_[6743]_ , \new_[6744]_ ,
    \new_[6745]_ , \new_[6748]_ , \new_[6752]_ , \new_[6753]_ ,
    \new_[6754]_ , \new_[6757]_ , \new_[6761]_ , \new_[6762]_ ,
    \new_[6763]_ , \new_[6766]_ , \new_[6770]_ , \new_[6771]_ ,
    \new_[6772]_ , \new_[6775]_ , \new_[6779]_ , \new_[6780]_ ,
    \new_[6781]_ , \new_[6784]_ , \new_[6788]_ , \new_[6789]_ ,
    \new_[6790]_ , \new_[6793]_ , \new_[6797]_ , \new_[6798]_ ,
    \new_[6799]_ , \new_[6802]_ , \new_[6806]_ , \new_[6807]_ ,
    \new_[6808]_ , \new_[6811]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6817]_ , \new_[6820]_ , \new_[6824]_ , \new_[6825]_ ,
    \new_[6826]_ , \new_[6829]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6835]_ , \new_[6838]_ , \new_[6842]_ , \new_[6843]_ ,
    \new_[6844]_ , \new_[6847]_ , \new_[6851]_ , \new_[6852]_ ,
    \new_[6853]_ , \new_[6856]_ , \new_[6860]_ , \new_[6861]_ ,
    \new_[6862]_ , \new_[6865]_ , \new_[6869]_ , \new_[6870]_ ,
    \new_[6871]_ , \new_[6874]_ , \new_[6878]_ , \new_[6879]_ ,
    \new_[6880]_ , \new_[6883]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6889]_ , \new_[6892]_ , \new_[6896]_ , \new_[6897]_ ,
    \new_[6898]_ , \new_[6901]_ , \new_[6905]_ , \new_[6906]_ ,
    \new_[6907]_ , \new_[6910]_ , \new_[6914]_ , \new_[6915]_ ,
    \new_[6916]_ , \new_[6919]_ , \new_[6923]_ , \new_[6924]_ ,
    \new_[6925]_ , \new_[6928]_ , \new_[6932]_ , \new_[6933]_ ,
    \new_[6934]_ , \new_[6937]_ , \new_[6941]_ , \new_[6942]_ ,
    \new_[6943]_ , \new_[6946]_ , \new_[6950]_ , \new_[6951]_ ,
    \new_[6952]_ , \new_[6955]_ , \new_[6959]_ , \new_[6960]_ ,
    \new_[6961]_ , \new_[6964]_ , \new_[6968]_ , \new_[6969]_ ,
    \new_[6970]_ , \new_[6973]_ , \new_[6977]_ , \new_[6978]_ ,
    \new_[6979]_ , \new_[6982]_ , \new_[6986]_ , \new_[6987]_ ,
    \new_[6988]_ , \new_[6991]_ , \new_[6995]_ , \new_[6996]_ ,
    \new_[6997]_ , \new_[7000]_ , \new_[7004]_ , \new_[7005]_ ,
    \new_[7006]_ , \new_[7009]_ , \new_[7013]_ , \new_[7014]_ ,
    \new_[7015]_ , \new_[7018]_ , \new_[7022]_ , \new_[7023]_ ,
    \new_[7024]_ , \new_[7027]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7033]_ , \new_[7036]_ , \new_[7040]_ , \new_[7041]_ ,
    \new_[7042]_ , \new_[7045]_ , \new_[7049]_ , \new_[7050]_ ,
    \new_[7051]_ , \new_[7054]_ , \new_[7058]_ , \new_[7059]_ ,
    \new_[7060]_ , \new_[7063]_ , \new_[7067]_ , \new_[7068]_ ,
    \new_[7069]_ , \new_[7072]_ , \new_[7076]_ , \new_[7077]_ ,
    \new_[7078]_ , \new_[7081]_ , \new_[7085]_ , \new_[7086]_ ,
    \new_[7087]_ , \new_[7090]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7096]_ , \new_[7099]_ , \new_[7103]_ , \new_[7104]_ ,
    \new_[7105]_ , \new_[7108]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7114]_ , \new_[7117]_ , \new_[7121]_ , \new_[7122]_ ,
    \new_[7123]_ , \new_[7126]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7132]_ , \new_[7135]_ , \new_[7139]_ , \new_[7140]_ ,
    \new_[7141]_ , \new_[7144]_ , \new_[7148]_ , \new_[7149]_ ,
    \new_[7150]_ , \new_[7153]_ , \new_[7157]_ , \new_[7158]_ ,
    \new_[7159]_ , \new_[7162]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7171]_ , \new_[7175]_ , \new_[7176]_ ,
    \new_[7177]_ , \new_[7180]_ , \new_[7184]_ , \new_[7185]_ ,
    \new_[7186]_ , \new_[7189]_ , \new_[7193]_ , \new_[7194]_ ,
    \new_[7195]_ , \new_[7198]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7207]_ , \new_[7211]_ , \new_[7212]_ ,
    \new_[7213]_ , \new_[7216]_ , \new_[7220]_ , \new_[7221]_ ,
    \new_[7222]_ , \new_[7225]_ , \new_[7229]_ , \new_[7230]_ ,
    \new_[7231]_ , \new_[7234]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7243]_ , \new_[7247]_ , \new_[7248]_ ,
    \new_[7249]_ , \new_[7252]_ , \new_[7256]_ , \new_[7257]_ ,
    \new_[7258]_ , \new_[7261]_ , \new_[7265]_ , \new_[7266]_ ,
    \new_[7267]_ , \new_[7270]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7276]_ , \new_[7279]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7288]_ , \new_[7292]_ , \new_[7293]_ ,
    \new_[7294]_ , \new_[7297]_ , \new_[7301]_ , \new_[7302]_ ,
    \new_[7303]_ , \new_[7306]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7312]_ , \new_[7315]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7321]_ , \new_[7324]_ , \new_[7328]_ , \new_[7329]_ ,
    \new_[7330]_ , \new_[7333]_ , \new_[7337]_ , \new_[7338]_ ,
    \new_[7339]_ , \new_[7342]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7348]_ , \new_[7351]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7357]_ , \new_[7360]_ , \new_[7364]_ , \new_[7365]_ ,
    \new_[7366]_ , \new_[7369]_ , \new_[7373]_ , \new_[7374]_ ,
    \new_[7375]_ , \new_[7378]_ , \new_[7382]_ , \new_[7383]_ ,
    \new_[7384]_ , \new_[7387]_ , \new_[7391]_ , \new_[7392]_ ,
    \new_[7393]_ , \new_[7396]_ , \new_[7400]_ , \new_[7401]_ ,
    \new_[7402]_ , \new_[7405]_ , \new_[7409]_ , \new_[7410]_ ,
    \new_[7411]_ , \new_[7414]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7423]_ , \new_[7427]_ , \new_[7428]_ ,
    \new_[7429]_ , \new_[7432]_ , \new_[7436]_ , \new_[7437]_ ,
    \new_[7438]_ , \new_[7441]_ , \new_[7445]_ , \new_[7446]_ ,
    \new_[7447]_ , \new_[7450]_ , \new_[7454]_ , \new_[7455]_ ,
    \new_[7456]_ , \new_[7459]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7465]_ , \new_[7468]_ , \new_[7472]_ , \new_[7473]_ ,
    \new_[7474]_ , \new_[7477]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7483]_ , \new_[7486]_ , \new_[7490]_ , \new_[7491]_ ,
    \new_[7492]_ , \new_[7495]_ , \new_[7499]_ , \new_[7500]_ ,
    \new_[7501]_ , \new_[7504]_ , \new_[7508]_ , \new_[7509]_ ,
    \new_[7510]_ , \new_[7513]_ , \new_[7517]_ , \new_[7518]_ ,
    \new_[7519]_ , \new_[7522]_ , \new_[7526]_ , \new_[7527]_ ,
    \new_[7528]_ , \new_[7531]_ , \new_[7535]_ , \new_[7536]_ ,
    \new_[7537]_ , \new_[7540]_ , \new_[7544]_ , \new_[7545]_ ,
    \new_[7546]_ , \new_[7549]_ , \new_[7553]_ , \new_[7554]_ ,
    \new_[7555]_ , \new_[7558]_ , \new_[7562]_ , \new_[7563]_ ,
    \new_[7564]_ , \new_[7567]_ , \new_[7571]_ , \new_[7572]_ ,
    \new_[7573]_ , \new_[7576]_ , \new_[7580]_ , \new_[7581]_ ,
    \new_[7582]_ , \new_[7585]_ , \new_[7589]_ , \new_[7590]_ ,
    \new_[7591]_ , \new_[7594]_ , \new_[7598]_ , \new_[7599]_ ,
    \new_[7600]_ , \new_[7603]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7609]_ , \new_[7612]_ , \new_[7616]_ , \new_[7617]_ ,
    \new_[7618]_ , \new_[7621]_ , \new_[7625]_ , \new_[7626]_ ,
    \new_[7627]_ , \new_[7630]_ , \new_[7634]_ , \new_[7635]_ ,
    \new_[7636]_ , \new_[7639]_ , \new_[7643]_ , \new_[7644]_ ,
    \new_[7645]_ , \new_[7648]_ , \new_[7652]_ , \new_[7653]_ ,
    \new_[7654]_ , \new_[7657]_ , \new_[7661]_ , \new_[7662]_ ,
    \new_[7663]_ , \new_[7666]_ , \new_[7670]_ , \new_[7671]_ ,
    \new_[7672]_ , \new_[7675]_ , \new_[7679]_ , \new_[7680]_ ,
    \new_[7681]_ , \new_[7684]_ , \new_[7688]_ , \new_[7689]_ ,
    \new_[7690]_ , \new_[7693]_ , \new_[7697]_ , \new_[7698]_ ,
    \new_[7699]_ , \new_[7702]_ , \new_[7706]_ , \new_[7707]_ ,
    \new_[7708]_ , \new_[7711]_ , \new_[7715]_ , \new_[7716]_ ,
    \new_[7717]_ , \new_[7720]_ , \new_[7724]_ , \new_[7725]_ ,
    \new_[7726]_ , \new_[7729]_ , \new_[7733]_ , \new_[7734]_ ,
    \new_[7735]_ , \new_[7738]_ , \new_[7742]_ , \new_[7743]_ ,
    \new_[7744]_ , \new_[7747]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7756]_ , \new_[7760]_ , \new_[7761]_ ,
    \new_[7762]_ , \new_[7765]_ , \new_[7769]_ , \new_[7770]_ ,
    \new_[7771]_ , \new_[7774]_ , \new_[7778]_ , \new_[7779]_ ,
    \new_[7780]_ , \new_[7783]_ , \new_[7787]_ , \new_[7788]_ ,
    \new_[7789]_ , \new_[7792]_ , \new_[7796]_ , \new_[7797]_ ,
    \new_[7798]_ , \new_[7801]_ , \new_[7805]_ , \new_[7806]_ ,
    \new_[7807]_ , \new_[7810]_ , \new_[7814]_ , \new_[7815]_ ,
    \new_[7816]_ , \new_[7819]_ , \new_[7823]_ , \new_[7824]_ ,
    \new_[7825]_ , \new_[7828]_ , \new_[7832]_ , \new_[7833]_ ,
    \new_[7834]_ , \new_[7837]_ , \new_[7841]_ , \new_[7842]_ ,
    \new_[7843]_ , \new_[7846]_ , \new_[7850]_ , \new_[7851]_ ,
    \new_[7852]_ , \new_[7855]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7861]_ , \new_[7864]_ , \new_[7868]_ , \new_[7869]_ ,
    \new_[7870]_ , \new_[7873]_ , \new_[7877]_ , \new_[7878]_ ,
    \new_[7879]_ , \new_[7882]_ , \new_[7886]_ , \new_[7887]_ ,
    \new_[7888]_ , \new_[7891]_ , \new_[7895]_ , \new_[7896]_ ,
    \new_[7897]_ , \new_[7900]_ , \new_[7904]_ , \new_[7905]_ ,
    \new_[7906]_ , \new_[7909]_ , \new_[7913]_ , \new_[7914]_ ,
    \new_[7915]_ , \new_[7918]_ , \new_[7922]_ , \new_[7923]_ ,
    \new_[7924]_ , \new_[7927]_ , \new_[7931]_ , \new_[7932]_ ,
    \new_[7933]_ , \new_[7936]_ , \new_[7940]_ , \new_[7941]_ ,
    \new_[7942]_ , \new_[7945]_ , \new_[7949]_ , \new_[7950]_ ,
    \new_[7951]_ , \new_[7954]_ , \new_[7958]_ , \new_[7959]_ ,
    \new_[7960]_ , \new_[7963]_ , \new_[7967]_ , \new_[7968]_ ,
    \new_[7969]_ , \new_[7972]_ , \new_[7976]_ , \new_[7977]_ ,
    \new_[7978]_ , \new_[7981]_ , \new_[7985]_ , \new_[7986]_ ,
    \new_[7987]_ , \new_[7990]_ , \new_[7994]_ , \new_[7995]_ ,
    \new_[7996]_ , \new_[7999]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8005]_ , \new_[8008]_ , \new_[8012]_ , \new_[8013]_ ,
    \new_[8014]_ , \new_[8017]_ , \new_[8021]_ , \new_[8022]_ ,
    \new_[8023]_ , \new_[8026]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8032]_ , \new_[8035]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8041]_ , \new_[8044]_ , \new_[8048]_ , \new_[8049]_ ,
    \new_[8050]_ , \new_[8053]_ , \new_[8057]_ , \new_[8058]_ ,
    \new_[8059]_ , \new_[8062]_ , \new_[8066]_ , \new_[8067]_ ,
    \new_[8068]_ , \new_[8071]_ , \new_[8075]_ , \new_[8076]_ ,
    \new_[8077]_ , \new_[8080]_ , \new_[8084]_ , \new_[8085]_ ,
    \new_[8086]_ , \new_[8089]_ , \new_[8093]_ , \new_[8094]_ ,
    \new_[8095]_ , \new_[8098]_ , \new_[8102]_ , \new_[8103]_ ,
    \new_[8104]_ , \new_[8107]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8113]_ , \new_[8116]_ , \new_[8120]_ , \new_[8121]_ ,
    \new_[8122]_ , \new_[8125]_ , \new_[8129]_ , \new_[8130]_ ,
    \new_[8131]_ , \new_[8134]_ , \new_[8138]_ , \new_[8139]_ ,
    \new_[8140]_ , \new_[8143]_ , \new_[8147]_ , \new_[8148]_ ,
    \new_[8149]_ , \new_[8152]_ , \new_[8156]_ , \new_[8157]_ ,
    \new_[8158]_ , \new_[8161]_ , \new_[8165]_ , \new_[8166]_ ,
    \new_[8167]_ , \new_[8170]_ , \new_[8174]_ , \new_[8175]_ ,
    \new_[8176]_ , \new_[8179]_ , \new_[8183]_ , \new_[8184]_ ,
    \new_[8185]_ , \new_[8188]_ , \new_[8192]_ , \new_[8193]_ ,
    \new_[8194]_ , \new_[8197]_ , \new_[8201]_ , \new_[8202]_ ,
    \new_[8203]_ , \new_[8206]_ , \new_[8210]_ , \new_[8211]_ ,
    \new_[8212]_ , \new_[8215]_ , \new_[8219]_ , \new_[8220]_ ,
    \new_[8221]_ , \new_[8224]_ , \new_[8228]_ , \new_[8229]_ ,
    \new_[8230]_ , \new_[8233]_ , \new_[8237]_ , \new_[8238]_ ,
    \new_[8239]_ , \new_[8242]_ , \new_[8246]_ , \new_[8247]_ ,
    \new_[8248]_ , \new_[8251]_ , \new_[8255]_ , \new_[8256]_ ,
    \new_[8257]_ , \new_[8260]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8266]_ , \new_[8269]_ , \new_[8273]_ , \new_[8274]_ ,
    \new_[8275]_ , \new_[8278]_ , \new_[8282]_ , \new_[8283]_ ,
    \new_[8284]_ , \new_[8287]_ , \new_[8291]_ , \new_[8292]_ ,
    \new_[8293]_ , \new_[8296]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8302]_ , \new_[8305]_ , \new_[8309]_ , \new_[8310]_ ,
    \new_[8311]_ , \new_[8314]_ , \new_[8318]_ , \new_[8319]_ ,
    \new_[8320]_ , \new_[8323]_ , \new_[8327]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8332]_ , \new_[8336]_ , \new_[8337]_ ,
    \new_[8338]_ , \new_[8341]_ , \new_[8345]_ , \new_[8346]_ ,
    \new_[8347]_ , \new_[8350]_ , \new_[8354]_ , \new_[8355]_ ,
    \new_[8356]_ , \new_[8359]_ , \new_[8363]_ , \new_[8364]_ ,
    \new_[8365]_ , \new_[8368]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8377]_ , \new_[8381]_ , \new_[8382]_ ,
    \new_[8383]_ , \new_[8386]_ , \new_[8390]_ , \new_[8391]_ ,
    \new_[8392]_ , \new_[8395]_ , \new_[8399]_ , \new_[8400]_ ,
    \new_[8401]_ , \new_[8404]_ , \new_[8408]_ , \new_[8409]_ ,
    \new_[8410]_ , \new_[8413]_ , \new_[8417]_ , \new_[8418]_ ,
    \new_[8419]_ , \new_[8422]_ , \new_[8426]_ , \new_[8427]_ ,
    \new_[8428]_ , \new_[8431]_ , \new_[8435]_ , \new_[8436]_ ,
    \new_[8437]_ , \new_[8440]_ , \new_[8444]_ , \new_[8445]_ ,
    \new_[8446]_ , \new_[8449]_ , \new_[8453]_ , \new_[8454]_ ,
    \new_[8455]_ , \new_[8458]_ , \new_[8462]_ , \new_[8463]_ ,
    \new_[8464]_ , \new_[8467]_ , \new_[8471]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8476]_ , \new_[8480]_ , \new_[8481]_ ,
    \new_[8482]_ , \new_[8485]_ , \new_[8489]_ , \new_[8490]_ ,
    \new_[8491]_ , \new_[8494]_ , \new_[8498]_ , \new_[8499]_ ,
    \new_[8500]_ , \new_[8503]_ , \new_[8507]_ , \new_[8508]_ ,
    \new_[8509]_ , \new_[8512]_ , \new_[8516]_ , \new_[8517]_ ,
    \new_[8518]_ , \new_[8521]_ , \new_[8525]_ , \new_[8526]_ ,
    \new_[8527]_ , \new_[8530]_ , \new_[8534]_ , \new_[8535]_ ,
    \new_[8536]_ , \new_[8539]_ , \new_[8543]_ , \new_[8544]_ ,
    \new_[8545]_ , \new_[8548]_ , \new_[8552]_ , \new_[8553]_ ,
    \new_[8554]_ , \new_[8557]_ , \new_[8561]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8566]_ , \new_[8570]_ , \new_[8571]_ ,
    \new_[8572]_ , \new_[8575]_ , \new_[8579]_ , \new_[8580]_ ,
    \new_[8581]_ , \new_[8584]_ , \new_[8588]_ , \new_[8589]_ ,
    \new_[8590]_ , \new_[8593]_ , \new_[8597]_ , \new_[8598]_ ,
    \new_[8599]_ , \new_[8602]_ , \new_[8606]_ , \new_[8607]_ ,
    \new_[8608]_ , \new_[8611]_ , \new_[8615]_ , \new_[8616]_ ,
    \new_[8617]_ , \new_[8620]_ , \new_[8624]_ , \new_[8625]_ ,
    \new_[8626]_ , \new_[8629]_ , \new_[8633]_ , \new_[8634]_ ,
    \new_[8635]_ , \new_[8638]_ , \new_[8642]_ , \new_[8643]_ ,
    \new_[8644]_ , \new_[8647]_ , \new_[8651]_ , \new_[8652]_ ,
    \new_[8653]_ , \new_[8656]_ , \new_[8660]_ , \new_[8661]_ ,
    \new_[8662]_ , \new_[8665]_ , \new_[8669]_ , \new_[8670]_ ,
    \new_[8671]_ , \new_[8674]_ , \new_[8678]_ , \new_[8679]_ ,
    \new_[8680]_ , \new_[8683]_ , \new_[8687]_ , \new_[8688]_ ,
    \new_[8689]_ , \new_[8692]_ , \new_[8696]_ , \new_[8697]_ ,
    \new_[8698]_ , \new_[8701]_ , \new_[8705]_ , \new_[8706]_ ,
    \new_[8707]_ , \new_[8710]_ , \new_[8714]_ , \new_[8715]_ ,
    \new_[8716]_ , \new_[8719]_ , \new_[8723]_ , \new_[8724]_ ,
    \new_[8725]_ , \new_[8728]_ , \new_[8732]_ , \new_[8733]_ ,
    \new_[8734]_ , \new_[8737]_ , \new_[8741]_ , \new_[8742]_ ,
    \new_[8743]_ , \new_[8746]_ , \new_[8750]_ , \new_[8751]_ ,
    \new_[8752]_ , \new_[8755]_ , \new_[8759]_ , \new_[8760]_ ,
    \new_[8761]_ , \new_[8764]_ , \new_[8768]_ , \new_[8769]_ ,
    \new_[8770]_ , \new_[8773]_ , \new_[8777]_ , \new_[8778]_ ,
    \new_[8779]_ , \new_[8782]_ , \new_[8786]_ , \new_[8787]_ ,
    \new_[8788]_ , \new_[8791]_ , \new_[8795]_ , \new_[8796]_ ,
    \new_[8797]_ , \new_[8800]_ , \new_[8804]_ , \new_[8805]_ ,
    \new_[8806]_ , \new_[8809]_ , \new_[8813]_ , \new_[8814]_ ,
    \new_[8815]_ , \new_[8818]_ , \new_[8822]_ , \new_[8823]_ ,
    \new_[8824]_ , \new_[8827]_ , \new_[8831]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8836]_ , \new_[8840]_ , \new_[8841]_ ,
    \new_[8842]_ , \new_[8845]_ , \new_[8849]_ , \new_[8850]_ ,
    \new_[8851]_ , \new_[8854]_ , \new_[8858]_ , \new_[8859]_ ,
    \new_[8860]_ , \new_[8863]_ , \new_[8867]_ , \new_[8868]_ ,
    \new_[8869]_ , \new_[8872]_ , \new_[8876]_ , \new_[8877]_ ,
    \new_[8878]_ , \new_[8881]_ , \new_[8885]_ , \new_[8886]_ ,
    \new_[8887]_ , \new_[8890]_ , \new_[8894]_ , \new_[8895]_ ,
    \new_[8896]_ , \new_[8899]_ , \new_[8903]_ , \new_[8904]_ ,
    \new_[8905]_ , \new_[8908]_ , \new_[8912]_ , \new_[8913]_ ,
    \new_[8914]_ , \new_[8917]_ , \new_[8921]_ , \new_[8922]_ ,
    \new_[8923]_ , \new_[8926]_ , \new_[8930]_ , \new_[8931]_ ,
    \new_[8932]_ , \new_[8935]_ , \new_[8939]_ , \new_[8940]_ ,
    \new_[8941]_ , \new_[8944]_ , \new_[8948]_ , \new_[8949]_ ,
    \new_[8950]_ , \new_[8953]_ , \new_[8957]_ , \new_[8958]_ ,
    \new_[8959]_ , \new_[8962]_ , \new_[8966]_ , \new_[8967]_ ,
    \new_[8968]_ , \new_[8971]_ , \new_[8975]_ , \new_[8976]_ ,
    \new_[8977]_ , \new_[8980]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8986]_ , \new_[8989]_ , \new_[8993]_ , \new_[8994]_ ,
    \new_[8995]_ , \new_[8998]_ , \new_[9002]_ , \new_[9003]_ ,
    \new_[9004]_ , \new_[9007]_ , \new_[9011]_ , \new_[9012]_ ,
    \new_[9013]_ , \new_[9016]_ , \new_[9020]_ , \new_[9021]_ ,
    \new_[9022]_ , \new_[9025]_ , \new_[9029]_ , \new_[9030]_ ,
    \new_[9031]_ , \new_[9034]_ , \new_[9038]_ , \new_[9039]_ ,
    \new_[9040]_ , \new_[9043]_ , \new_[9047]_ , \new_[9048]_ ,
    \new_[9049]_ , \new_[9052]_ , \new_[9056]_ , \new_[9057]_ ,
    \new_[9058]_ , \new_[9061]_ , \new_[9065]_ , \new_[9066]_ ,
    \new_[9067]_ , \new_[9070]_ , \new_[9074]_ , \new_[9075]_ ,
    \new_[9076]_ , \new_[9079]_ , \new_[9083]_ , \new_[9084]_ ,
    \new_[9085]_ , \new_[9088]_ , \new_[9092]_ , \new_[9093]_ ,
    \new_[9094]_ , \new_[9097]_ , \new_[9101]_ , \new_[9102]_ ,
    \new_[9103]_ , \new_[9106]_ , \new_[9110]_ , \new_[9111]_ ,
    \new_[9112]_ , \new_[9115]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9121]_ , \new_[9124]_ , \new_[9128]_ , \new_[9129]_ ,
    \new_[9130]_ , \new_[9133]_ , \new_[9137]_ , \new_[9138]_ ,
    \new_[9139]_ , \new_[9142]_ , \new_[9146]_ , \new_[9147]_ ,
    \new_[9148]_ , \new_[9151]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9160]_ , \new_[9164]_ , \new_[9165]_ ,
    \new_[9166]_ , \new_[9169]_ , \new_[9173]_ , \new_[9174]_ ,
    \new_[9175]_ , \new_[9178]_ , \new_[9182]_ , \new_[9183]_ ,
    \new_[9184]_ , \new_[9187]_ , \new_[9191]_ , \new_[9192]_ ,
    \new_[9193]_ , \new_[9196]_ , \new_[9200]_ , \new_[9201]_ ,
    \new_[9202]_ , \new_[9205]_ , \new_[9209]_ , \new_[9210]_ ,
    \new_[9211]_ , \new_[9214]_ , \new_[9218]_ , \new_[9219]_ ,
    \new_[9220]_ , \new_[9223]_ , \new_[9227]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9232]_ , \new_[9236]_ , \new_[9237]_ ,
    \new_[9238]_ , \new_[9241]_ , \new_[9245]_ , \new_[9246]_ ,
    \new_[9247]_ , \new_[9250]_ , \new_[9254]_ , \new_[9255]_ ,
    \new_[9256]_ , \new_[9259]_ , \new_[9263]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9268]_ , \new_[9272]_ , \new_[9273]_ ,
    \new_[9274]_ , \new_[9277]_ , \new_[9281]_ , \new_[9282]_ ,
    \new_[9283]_ , \new_[9286]_ , \new_[9290]_ , \new_[9291]_ ,
    \new_[9292]_ , \new_[9295]_ , \new_[9299]_ , \new_[9300]_ ,
    \new_[9301]_ , \new_[9304]_ , \new_[9308]_ , \new_[9309]_ ,
    \new_[9310]_ , \new_[9313]_ , \new_[9317]_ , \new_[9318]_ ,
    \new_[9319]_ , \new_[9322]_ , \new_[9326]_ , \new_[9327]_ ,
    \new_[9328]_ , \new_[9331]_ , \new_[9335]_ , \new_[9336]_ ,
    \new_[9337]_ , \new_[9340]_ , \new_[9344]_ , \new_[9345]_ ,
    \new_[9346]_ , \new_[9349]_ , \new_[9353]_ , \new_[9354]_ ,
    \new_[9355]_ , \new_[9358]_ , \new_[9362]_ , \new_[9363]_ ,
    \new_[9364]_ , \new_[9367]_ , \new_[9371]_ , \new_[9372]_ ,
    \new_[9373]_ , \new_[9376]_ , \new_[9380]_ , \new_[9381]_ ,
    \new_[9382]_ , \new_[9385]_ , \new_[9389]_ , \new_[9390]_ ,
    \new_[9391]_ , \new_[9394]_ , \new_[9398]_ , \new_[9399]_ ,
    \new_[9400]_ , \new_[9403]_ , \new_[9407]_ , \new_[9408]_ ,
    \new_[9409]_ , \new_[9412]_ , \new_[9416]_ , \new_[9417]_ ,
    \new_[9418]_ , \new_[9421]_ , \new_[9425]_ , \new_[9426]_ ,
    \new_[9427]_ , \new_[9430]_ , \new_[9434]_ , \new_[9435]_ ,
    \new_[9436]_ , \new_[9439]_ , \new_[9443]_ , \new_[9444]_ ,
    \new_[9445]_ , \new_[9448]_ , \new_[9452]_ , \new_[9453]_ ,
    \new_[9454]_ , \new_[9457]_ , \new_[9461]_ , \new_[9462]_ ,
    \new_[9463]_ , \new_[9466]_ , \new_[9470]_ , \new_[9471]_ ,
    \new_[9472]_ , \new_[9475]_ , \new_[9479]_ , \new_[9480]_ ,
    \new_[9481]_ , \new_[9484]_ , \new_[9488]_ , \new_[9489]_ ,
    \new_[9490]_ , \new_[9493]_ , \new_[9497]_ , \new_[9498]_ ,
    \new_[9499]_ , \new_[9502]_ , \new_[9506]_ , \new_[9507]_ ,
    \new_[9508]_ , \new_[9511]_ , \new_[9515]_ , \new_[9516]_ ,
    \new_[9517]_ , \new_[9520]_ , \new_[9524]_ , \new_[9525]_ ,
    \new_[9526]_ , \new_[9529]_ , \new_[9533]_ , \new_[9534]_ ,
    \new_[9535]_ , \new_[9538]_ , \new_[9542]_ , \new_[9543]_ ,
    \new_[9544]_ , \new_[9547]_ , \new_[9551]_ , \new_[9552]_ ,
    \new_[9553]_ , \new_[9556]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9562]_ , \new_[9565]_ , \new_[9569]_ , \new_[9570]_ ,
    \new_[9571]_ , \new_[9574]_ , \new_[9578]_ , \new_[9579]_ ,
    \new_[9580]_ , \new_[9583]_ , \new_[9587]_ , \new_[9588]_ ,
    \new_[9589]_ , \new_[9592]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9598]_ , \new_[9601]_ , \new_[9605]_ , \new_[9606]_ ,
    \new_[9607]_ , \new_[9610]_ , \new_[9614]_ , \new_[9615]_ ,
    \new_[9616]_ , \new_[9619]_ , \new_[9623]_ , \new_[9624]_ ,
    \new_[9625]_ , \new_[9628]_ , \new_[9632]_ , \new_[9633]_ ,
    \new_[9634]_ , \new_[9637]_ , \new_[9641]_ , \new_[9642]_ ,
    \new_[9643]_ , \new_[9646]_ , \new_[9650]_ , \new_[9651]_ ,
    \new_[9652]_ , \new_[9655]_ , \new_[9659]_ , \new_[9660]_ ,
    \new_[9661]_ , \new_[9664]_ , \new_[9668]_ , \new_[9669]_ ,
    \new_[9670]_ , \new_[9673]_ , \new_[9677]_ , \new_[9678]_ ,
    \new_[9679]_ , \new_[9682]_ , \new_[9686]_ , \new_[9687]_ ,
    \new_[9688]_ , \new_[9691]_ , \new_[9695]_ , \new_[9696]_ ,
    \new_[9697]_ , \new_[9700]_ , \new_[9704]_ , \new_[9705]_ ,
    \new_[9706]_ , \new_[9709]_ , \new_[9713]_ , \new_[9714]_ ,
    \new_[9715]_ , \new_[9718]_ , \new_[9722]_ , \new_[9723]_ ,
    \new_[9724]_ , \new_[9727]_ , \new_[9731]_ , \new_[9732]_ ,
    \new_[9733]_ , \new_[9736]_ , \new_[9740]_ , \new_[9741]_ ,
    \new_[9742]_ , \new_[9745]_ , \new_[9749]_ , \new_[9750]_ ,
    \new_[9751]_ , \new_[9754]_ , \new_[9758]_ , \new_[9759]_ ,
    \new_[9760]_ , \new_[9763]_ , \new_[9767]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9772]_ , \new_[9776]_ , \new_[9777]_ ,
    \new_[9778]_ , \new_[9781]_ , \new_[9785]_ , \new_[9786]_ ,
    \new_[9787]_ , \new_[9790]_ , \new_[9794]_ , \new_[9795]_ ,
    \new_[9796]_ , \new_[9799]_ , \new_[9803]_ , \new_[9804]_ ,
    \new_[9805]_ , \new_[9808]_ , \new_[9812]_ , \new_[9813]_ ,
    \new_[9814]_ , \new_[9817]_ , \new_[9821]_ , \new_[9822]_ ,
    \new_[9823]_ , \new_[9826]_ , \new_[9830]_ , \new_[9831]_ ,
    \new_[9832]_ , \new_[9835]_ , \new_[9839]_ , \new_[9840]_ ,
    \new_[9841]_ , \new_[9844]_ , \new_[9848]_ , \new_[9849]_ ,
    \new_[9850]_ , \new_[9853]_ , \new_[9857]_ , \new_[9858]_ ,
    \new_[9859]_ , \new_[9862]_ , \new_[9866]_ , \new_[9867]_ ,
    \new_[9868]_ , \new_[9871]_ , \new_[9875]_ , \new_[9876]_ ,
    \new_[9877]_ , \new_[9880]_ , \new_[9884]_ , \new_[9885]_ ,
    \new_[9886]_ , \new_[9889]_ , \new_[9893]_ , \new_[9894]_ ,
    \new_[9895]_ , \new_[9898]_ , \new_[9902]_ , \new_[9903]_ ,
    \new_[9904]_ , \new_[9907]_ , \new_[9911]_ , \new_[9912]_ ,
    \new_[9913]_ , \new_[9916]_ , \new_[9920]_ , \new_[9921]_ ,
    \new_[9922]_ , \new_[9925]_ , \new_[9929]_ , \new_[9930]_ ,
    \new_[9931]_ , \new_[9934]_ , \new_[9938]_ , \new_[9939]_ ,
    \new_[9940]_ , \new_[9943]_ , \new_[9947]_ , \new_[9948]_ ,
    \new_[9949]_ , \new_[9952]_ , \new_[9956]_ , \new_[9957]_ ,
    \new_[9958]_ , \new_[9961]_ , \new_[9965]_ , \new_[9966]_ ,
    \new_[9967]_ , \new_[9970]_ , \new_[9974]_ , \new_[9975]_ ,
    \new_[9976]_ , \new_[9979]_ , \new_[9983]_ , \new_[9984]_ ,
    \new_[9985]_ , \new_[9989]_ , \new_[9990]_ , \new_[9994]_ ,
    \new_[9995]_ , \new_[9996]_ , \new_[9999]_ , \new_[10003]_ ,
    \new_[10004]_ , \new_[10005]_ , \new_[10009]_ , \new_[10010]_ ,
    \new_[10014]_ , \new_[10015]_ , \new_[10016]_ , \new_[10019]_ ,
    \new_[10023]_ , \new_[10024]_ , \new_[10025]_ , \new_[10029]_ ,
    \new_[10030]_ , \new_[10034]_ , \new_[10035]_ , \new_[10036]_ ,
    \new_[10039]_ , \new_[10043]_ , \new_[10044]_ , \new_[10045]_ ,
    \new_[10049]_ , \new_[10050]_ , \new_[10054]_ , \new_[10055]_ ,
    \new_[10056]_ , \new_[10059]_ , \new_[10063]_ , \new_[10064]_ ,
    \new_[10065]_ , \new_[10069]_ , \new_[10070]_ , \new_[10074]_ ,
    \new_[10075]_ , \new_[10076]_ , \new_[10079]_ , \new_[10083]_ ,
    \new_[10084]_ , \new_[10085]_ , \new_[10089]_ , \new_[10090]_ ,
    \new_[10094]_ , \new_[10095]_ , \new_[10096]_ , \new_[10099]_ ,
    \new_[10103]_ , \new_[10104]_ , \new_[10105]_ , \new_[10109]_ ,
    \new_[10110]_ , \new_[10114]_ , \new_[10115]_ , \new_[10116]_ ,
    \new_[10119]_ , \new_[10123]_ , \new_[10124]_ , \new_[10125]_ ,
    \new_[10129]_ , \new_[10130]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10136]_ , \new_[10139]_ , \new_[10143]_ , \new_[10144]_ ,
    \new_[10145]_ , \new_[10149]_ , \new_[10150]_ , \new_[10154]_ ,
    \new_[10155]_ , \new_[10156]_ , \new_[10159]_ , \new_[10163]_ ,
    \new_[10164]_ , \new_[10165]_ , \new_[10169]_ , \new_[10170]_ ,
    \new_[10174]_ , \new_[10175]_ , \new_[10176]_ , \new_[10179]_ ,
    \new_[10183]_ , \new_[10184]_ , \new_[10185]_ , \new_[10189]_ ,
    \new_[10190]_ , \new_[10194]_ , \new_[10195]_ , \new_[10196]_ ,
    \new_[10199]_ , \new_[10203]_ , \new_[10204]_ , \new_[10205]_ ,
    \new_[10209]_ , \new_[10210]_ , \new_[10214]_ , \new_[10215]_ ,
    \new_[10216]_ , \new_[10219]_ , \new_[10223]_ , \new_[10224]_ ,
    \new_[10225]_ , \new_[10229]_ , \new_[10230]_ , \new_[10234]_ ,
    \new_[10235]_ , \new_[10236]_ , \new_[10239]_ , \new_[10243]_ ,
    \new_[10244]_ , \new_[10245]_ , \new_[10249]_ , \new_[10250]_ ,
    \new_[10254]_ , \new_[10255]_ , \new_[10256]_ , \new_[10259]_ ,
    \new_[10263]_ , \new_[10264]_ , \new_[10265]_ , \new_[10269]_ ,
    \new_[10270]_ , \new_[10274]_ , \new_[10275]_ , \new_[10276]_ ,
    \new_[10279]_ , \new_[10283]_ , \new_[10284]_ , \new_[10285]_ ,
    \new_[10289]_ , \new_[10290]_ , \new_[10294]_ , \new_[10295]_ ,
    \new_[10296]_ , \new_[10299]_ , \new_[10303]_ , \new_[10304]_ ,
    \new_[10305]_ , \new_[10309]_ , \new_[10310]_ , \new_[10314]_ ,
    \new_[10315]_ , \new_[10316]_ , \new_[10319]_ , \new_[10323]_ ,
    \new_[10324]_ , \new_[10325]_ , \new_[10329]_ , \new_[10330]_ ,
    \new_[10334]_ , \new_[10335]_ , \new_[10336]_ , \new_[10339]_ ,
    \new_[10343]_ , \new_[10344]_ , \new_[10345]_ , \new_[10349]_ ,
    \new_[10350]_ , \new_[10354]_ , \new_[10355]_ , \new_[10356]_ ,
    \new_[10359]_ , \new_[10363]_ , \new_[10364]_ , \new_[10365]_ ,
    \new_[10369]_ , \new_[10370]_ , \new_[10374]_ , \new_[10375]_ ,
    \new_[10376]_ , \new_[10379]_ , \new_[10383]_ , \new_[10384]_ ,
    \new_[10385]_ , \new_[10389]_ , \new_[10390]_ , \new_[10394]_ ,
    \new_[10395]_ , \new_[10396]_ , \new_[10399]_ , \new_[10403]_ ,
    \new_[10404]_ , \new_[10405]_ , \new_[10409]_ , \new_[10410]_ ,
    \new_[10414]_ , \new_[10415]_ , \new_[10416]_ , \new_[10419]_ ,
    \new_[10423]_ , \new_[10424]_ , \new_[10425]_ , \new_[10429]_ ,
    \new_[10430]_ , \new_[10434]_ , \new_[10435]_ , \new_[10436]_ ,
    \new_[10439]_ , \new_[10443]_ , \new_[10444]_ , \new_[10445]_ ,
    \new_[10449]_ , \new_[10450]_ , \new_[10454]_ , \new_[10455]_ ,
    \new_[10456]_ , \new_[10459]_ , \new_[10463]_ , \new_[10464]_ ,
    \new_[10465]_ , \new_[10469]_ , \new_[10470]_ , \new_[10474]_ ,
    \new_[10475]_ , \new_[10476]_ , \new_[10479]_ , \new_[10483]_ ,
    \new_[10484]_ , \new_[10485]_ , \new_[10489]_ , \new_[10490]_ ,
    \new_[10494]_ , \new_[10495]_ , \new_[10496]_ , \new_[10499]_ ,
    \new_[10503]_ , \new_[10504]_ , \new_[10505]_ , \new_[10509]_ ,
    \new_[10510]_ , \new_[10514]_ , \new_[10515]_ , \new_[10516]_ ,
    \new_[10519]_ , \new_[10523]_ , \new_[10524]_ , \new_[10525]_ ,
    \new_[10529]_ , \new_[10530]_ , \new_[10534]_ , \new_[10535]_ ,
    \new_[10536]_ , \new_[10539]_ , \new_[10543]_ , \new_[10544]_ ,
    \new_[10545]_ , \new_[10549]_ , \new_[10550]_ , \new_[10554]_ ,
    \new_[10555]_ , \new_[10556]_ , \new_[10559]_ , \new_[10563]_ ,
    \new_[10564]_ , \new_[10565]_ , \new_[10569]_ , \new_[10570]_ ,
    \new_[10574]_ , \new_[10575]_ , \new_[10576]_ , \new_[10579]_ ,
    \new_[10583]_ , \new_[10584]_ , \new_[10585]_ , \new_[10589]_ ,
    \new_[10590]_ , \new_[10594]_ , \new_[10595]_ , \new_[10596]_ ,
    \new_[10599]_ , \new_[10603]_ , \new_[10604]_ , \new_[10605]_ ,
    \new_[10609]_ , \new_[10610]_ , \new_[10614]_ , \new_[10615]_ ,
    \new_[10616]_ , \new_[10619]_ , \new_[10623]_ , \new_[10624]_ ,
    \new_[10625]_ , \new_[10629]_ , \new_[10630]_ , \new_[10634]_ ,
    \new_[10635]_ , \new_[10636]_ , \new_[10639]_ , \new_[10643]_ ,
    \new_[10644]_ , \new_[10645]_ , \new_[10649]_ , \new_[10650]_ ,
    \new_[10654]_ , \new_[10655]_ , \new_[10656]_ , \new_[10659]_ ,
    \new_[10663]_ , \new_[10664]_ , \new_[10665]_ , \new_[10669]_ ,
    \new_[10670]_ , \new_[10674]_ , \new_[10675]_ , \new_[10676]_ ,
    \new_[10679]_ , \new_[10683]_ , \new_[10684]_ , \new_[10685]_ ,
    \new_[10689]_ , \new_[10690]_ , \new_[10694]_ , \new_[10695]_ ,
    \new_[10696]_ , \new_[10699]_ , \new_[10703]_ , \new_[10704]_ ,
    \new_[10705]_ , \new_[10709]_ , \new_[10710]_ , \new_[10714]_ ,
    \new_[10715]_ , \new_[10716]_ , \new_[10719]_ , \new_[10723]_ ,
    \new_[10724]_ , \new_[10725]_ , \new_[10729]_ , \new_[10730]_ ,
    \new_[10734]_ , \new_[10735]_ , \new_[10736]_ , \new_[10739]_ ,
    \new_[10743]_ , \new_[10744]_ , \new_[10745]_ , \new_[10749]_ ,
    \new_[10750]_ , \new_[10754]_ , \new_[10755]_ , \new_[10756]_ ,
    \new_[10759]_ , \new_[10763]_ , \new_[10764]_ , \new_[10765]_ ,
    \new_[10769]_ , \new_[10770]_ , \new_[10774]_ , \new_[10775]_ ,
    \new_[10776]_ , \new_[10779]_ , \new_[10783]_ , \new_[10784]_ ,
    \new_[10785]_ , \new_[10789]_ , \new_[10790]_ , \new_[10794]_ ,
    \new_[10795]_ , \new_[10796]_ , \new_[10799]_ , \new_[10803]_ ,
    \new_[10804]_ , \new_[10805]_ , \new_[10809]_ , \new_[10810]_ ,
    \new_[10814]_ , \new_[10815]_ , \new_[10816]_ , \new_[10819]_ ,
    \new_[10823]_ , \new_[10824]_ , \new_[10825]_ , \new_[10829]_ ,
    \new_[10830]_ , \new_[10834]_ , \new_[10835]_ , \new_[10836]_ ,
    \new_[10839]_ , \new_[10843]_ , \new_[10844]_ , \new_[10845]_ ,
    \new_[10849]_ , \new_[10850]_ , \new_[10854]_ , \new_[10855]_ ,
    \new_[10856]_ , \new_[10859]_ , \new_[10863]_ , \new_[10864]_ ,
    \new_[10865]_ , \new_[10869]_ , \new_[10870]_ , \new_[10874]_ ,
    \new_[10875]_ , \new_[10876]_ , \new_[10879]_ , \new_[10883]_ ,
    \new_[10884]_ , \new_[10885]_ , \new_[10889]_ , \new_[10890]_ ,
    \new_[10894]_ , \new_[10895]_ , \new_[10896]_ , \new_[10899]_ ,
    \new_[10903]_ , \new_[10904]_ , \new_[10905]_ , \new_[10909]_ ,
    \new_[10910]_ , \new_[10914]_ , \new_[10915]_ , \new_[10916]_ ,
    \new_[10919]_ , \new_[10923]_ , \new_[10924]_ , \new_[10925]_ ,
    \new_[10929]_ , \new_[10930]_ , \new_[10934]_ , \new_[10935]_ ,
    \new_[10936]_ , \new_[10939]_ , \new_[10943]_ , \new_[10944]_ ,
    \new_[10945]_ , \new_[10949]_ , \new_[10950]_ , \new_[10954]_ ,
    \new_[10955]_ , \new_[10956]_ , \new_[10959]_ , \new_[10963]_ ,
    \new_[10964]_ , \new_[10965]_ , \new_[10969]_ , \new_[10970]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10976]_ , \new_[10979]_ ,
    \new_[10983]_ , \new_[10984]_ , \new_[10985]_ , \new_[10989]_ ,
    \new_[10990]_ , \new_[10994]_ , \new_[10995]_ , \new_[10996]_ ,
    \new_[10999]_ , \new_[11003]_ , \new_[11004]_ , \new_[11005]_ ,
    \new_[11009]_ , \new_[11010]_ , \new_[11014]_ , \new_[11015]_ ,
    \new_[11016]_ , \new_[11019]_ , \new_[11023]_ , \new_[11024]_ ,
    \new_[11025]_ , \new_[11029]_ , \new_[11030]_ , \new_[11034]_ ,
    \new_[11035]_ , \new_[11036]_ , \new_[11039]_ , \new_[11043]_ ,
    \new_[11044]_ , \new_[11045]_ , \new_[11049]_ , \new_[11050]_ ,
    \new_[11054]_ , \new_[11055]_ , \new_[11056]_ , \new_[11059]_ ,
    \new_[11063]_ , \new_[11064]_ , \new_[11065]_ , \new_[11069]_ ,
    \new_[11070]_ , \new_[11074]_ , \new_[11075]_ , \new_[11076]_ ,
    \new_[11079]_ , \new_[11083]_ , \new_[11084]_ , \new_[11085]_ ,
    \new_[11089]_ , \new_[11090]_ , \new_[11094]_ , \new_[11095]_ ,
    \new_[11096]_ , \new_[11099]_ , \new_[11103]_ , \new_[11104]_ ,
    \new_[11105]_ , \new_[11109]_ , \new_[11110]_ , \new_[11114]_ ,
    \new_[11115]_ , \new_[11116]_ , \new_[11119]_ , \new_[11123]_ ,
    \new_[11124]_ , \new_[11125]_ , \new_[11129]_ , \new_[11130]_ ,
    \new_[11134]_ , \new_[11135]_ , \new_[11136]_ , \new_[11139]_ ,
    \new_[11143]_ , \new_[11144]_ , \new_[11145]_ , \new_[11149]_ ,
    \new_[11150]_ , \new_[11154]_ , \new_[11155]_ , \new_[11156]_ ,
    \new_[11159]_ , \new_[11163]_ , \new_[11164]_ , \new_[11165]_ ,
    \new_[11169]_ , \new_[11170]_ , \new_[11174]_ , \new_[11175]_ ,
    \new_[11176]_ , \new_[11179]_ , \new_[11183]_ , \new_[11184]_ ,
    \new_[11185]_ , \new_[11189]_ , \new_[11190]_ , \new_[11194]_ ,
    \new_[11195]_ , \new_[11196]_ , \new_[11199]_ , \new_[11203]_ ,
    \new_[11204]_ , \new_[11205]_ , \new_[11209]_ , \new_[11210]_ ,
    \new_[11214]_ , \new_[11215]_ , \new_[11216]_ , \new_[11219]_ ,
    \new_[11223]_ , \new_[11224]_ , \new_[11225]_ , \new_[11229]_ ,
    \new_[11230]_ , \new_[11234]_ , \new_[11235]_ , \new_[11236]_ ,
    \new_[11239]_ , \new_[11243]_ , \new_[11244]_ , \new_[11245]_ ,
    \new_[11249]_ , \new_[11250]_ , \new_[11254]_ , \new_[11255]_ ,
    \new_[11256]_ , \new_[11259]_ , \new_[11263]_ , \new_[11264]_ ,
    \new_[11265]_ , \new_[11269]_ , \new_[11270]_ , \new_[11274]_ ,
    \new_[11275]_ , \new_[11276]_ , \new_[11279]_ , \new_[11283]_ ,
    \new_[11284]_ , \new_[11285]_ , \new_[11289]_ , \new_[11290]_ ,
    \new_[11294]_ , \new_[11295]_ , \new_[11296]_ , \new_[11299]_ ,
    \new_[11303]_ , \new_[11304]_ , \new_[11305]_ , \new_[11309]_ ,
    \new_[11310]_ , \new_[11314]_ , \new_[11315]_ , \new_[11316]_ ,
    \new_[11319]_ , \new_[11323]_ , \new_[11324]_ , \new_[11325]_ ,
    \new_[11329]_ , \new_[11330]_ , \new_[11334]_ , \new_[11335]_ ,
    \new_[11336]_ , \new_[11339]_ , \new_[11343]_ , \new_[11344]_ ,
    \new_[11345]_ , \new_[11349]_ , \new_[11350]_ , \new_[11354]_ ,
    \new_[11355]_ , \new_[11356]_ , \new_[11359]_ , \new_[11363]_ ,
    \new_[11364]_ , \new_[11365]_ , \new_[11369]_ , \new_[11370]_ ,
    \new_[11374]_ , \new_[11375]_ , \new_[11376]_ , \new_[11379]_ ,
    \new_[11383]_ , \new_[11384]_ , \new_[11385]_ , \new_[11389]_ ,
    \new_[11390]_ , \new_[11394]_ , \new_[11395]_ , \new_[11396]_ ,
    \new_[11399]_ , \new_[11403]_ , \new_[11404]_ , \new_[11405]_ ,
    \new_[11409]_ , \new_[11410]_ , \new_[11414]_ , \new_[11415]_ ,
    \new_[11416]_ , \new_[11419]_ , \new_[11423]_ , \new_[11424]_ ,
    \new_[11425]_ , \new_[11429]_ , \new_[11430]_ , \new_[11434]_ ,
    \new_[11435]_ , \new_[11436]_ , \new_[11439]_ , \new_[11443]_ ,
    \new_[11444]_ , \new_[11445]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11454]_ , \new_[11455]_ , \new_[11456]_ , \new_[11459]_ ,
    \new_[11463]_ , \new_[11464]_ , \new_[11465]_ , \new_[11469]_ ,
    \new_[11470]_ , \new_[11474]_ , \new_[11475]_ , \new_[11476]_ ,
    \new_[11479]_ , \new_[11483]_ , \new_[11484]_ , \new_[11485]_ ,
    \new_[11489]_ , \new_[11490]_ , \new_[11494]_ , \new_[11495]_ ,
    \new_[11496]_ , \new_[11499]_ , \new_[11503]_ , \new_[11504]_ ,
    \new_[11505]_ , \new_[11509]_ , \new_[11510]_ , \new_[11514]_ ,
    \new_[11515]_ , \new_[11516]_ , \new_[11519]_ , \new_[11523]_ ,
    \new_[11524]_ , \new_[11525]_ , \new_[11529]_ , \new_[11530]_ ,
    \new_[11534]_ , \new_[11535]_ , \new_[11536]_ , \new_[11539]_ ,
    \new_[11543]_ , \new_[11544]_ , \new_[11545]_ , \new_[11549]_ ,
    \new_[11550]_ , \new_[11554]_ , \new_[11555]_ , \new_[11556]_ ,
    \new_[11559]_ , \new_[11563]_ , \new_[11564]_ , \new_[11565]_ ,
    \new_[11569]_ , \new_[11570]_ , \new_[11574]_ , \new_[11575]_ ,
    \new_[11576]_ , \new_[11579]_ , \new_[11583]_ , \new_[11584]_ ,
    \new_[11585]_ , \new_[11589]_ , \new_[11590]_ , \new_[11594]_ ,
    \new_[11595]_ , \new_[11596]_ , \new_[11599]_ , \new_[11603]_ ,
    \new_[11604]_ , \new_[11605]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11614]_ , \new_[11615]_ , \new_[11616]_ , \new_[11619]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11625]_ , \new_[11629]_ ,
    \new_[11630]_ , \new_[11634]_ , \new_[11635]_ , \new_[11636]_ ,
    \new_[11639]_ , \new_[11643]_ , \new_[11644]_ , \new_[11645]_ ,
    \new_[11649]_ , \new_[11650]_ , \new_[11654]_ , \new_[11655]_ ,
    \new_[11656]_ , \new_[11659]_ , \new_[11663]_ , \new_[11664]_ ,
    \new_[11665]_ , \new_[11669]_ , \new_[11670]_ , \new_[11674]_ ,
    \new_[11675]_ , \new_[11676]_ , \new_[11679]_ , \new_[11683]_ ,
    \new_[11684]_ , \new_[11685]_ , \new_[11689]_ , \new_[11690]_ ,
    \new_[11694]_ , \new_[11695]_ , \new_[11696]_ , \new_[11699]_ ,
    \new_[11703]_ , \new_[11704]_ , \new_[11705]_ , \new_[11709]_ ,
    \new_[11710]_ , \new_[11714]_ , \new_[11715]_ , \new_[11716]_ ,
    \new_[11719]_ , \new_[11723]_ , \new_[11724]_ , \new_[11725]_ ,
    \new_[11729]_ , \new_[11730]_ , \new_[11734]_ , \new_[11735]_ ,
    \new_[11736]_ , \new_[11739]_ , \new_[11743]_ , \new_[11744]_ ,
    \new_[11745]_ , \new_[11749]_ , \new_[11750]_ , \new_[11754]_ ,
    \new_[11755]_ , \new_[11756]_ , \new_[11759]_ , \new_[11763]_ ,
    \new_[11764]_ , \new_[11765]_ , \new_[11769]_ , \new_[11770]_ ,
    \new_[11774]_ , \new_[11775]_ , \new_[11776]_ , \new_[11779]_ ,
    \new_[11783]_ , \new_[11784]_ , \new_[11785]_ , \new_[11789]_ ,
    \new_[11790]_ , \new_[11794]_ , \new_[11795]_ , \new_[11796]_ ,
    \new_[11799]_ , \new_[11803]_ , \new_[11804]_ , \new_[11805]_ ,
    \new_[11809]_ , \new_[11810]_ , \new_[11814]_ , \new_[11815]_ ,
    \new_[11816]_ , \new_[11819]_ , \new_[11823]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11829]_ , \new_[11830]_ , \new_[11834]_ ,
    \new_[11835]_ , \new_[11836]_ , \new_[11839]_ , \new_[11843]_ ,
    \new_[11844]_ , \new_[11845]_ , \new_[11849]_ , \new_[11850]_ ,
    \new_[11854]_ , \new_[11855]_ , \new_[11856]_ , \new_[11859]_ ,
    \new_[11863]_ , \new_[11864]_ , \new_[11865]_ , \new_[11869]_ ,
    \new_[11870]_ , \new_[11874]_ , \new_[11875]_ , \new_[11876]_ ,
    \new_[11879]_ , \new_[11883]_ , \new_[11884]_ , \new_[11885]_ ,
    \new_[11889]_ , \new_[11890]_ , \new_[11894]_ , \new_[11895]_ ,
    \new_[11896]_ , \new_[11899]_ , \new_[11903]_ , \new_[11904]_ ,
    \new_[11905]_ , \new_[11909]_ , \new_[11910]_ , \new_[11914]_ ,
    \new_[11915]_ , \new_[11916]_ , \new_[11919]_ , \new_[11923]_ ,
    \new_[11924]_ , \new_[11925]_ , \new_[11929]_ , \new_[11930]_ ,
    \new_[11934]_ , \new_[11935]_ , \new_[11936]_ , \new_[11939]_ ,
    \new_[11943]_ , \new_[11944]_ , \new_[11945]_ , \new_[11949]_ ,
    \new_[11950]_ , \new_[11954]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11959]_ , \new_[11963]_ , \new_[11964]_ , \new_[11965]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11974]_ , \new_[11975]_ ,
    \new_[11976]_ , \new_[11979]_ , \new_[11983]_ , \new_[11984]_ ,
    \new_[11985]_ , \new_[11989]_ , \new_[11990]_ , \new_[11994]_ ,
    \new_[11995]_ , \new_[11996]_ , \new_[11999]_ , \new_[12003]_ ,
    \new_[12004]_ , \new_[12005]_ , \new_[12009]_ , \new_[12010]_ ,
    \new_[12014]_ , \new_[12015]_ , \new_[12016]_ , \new_[12019]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12025]_ , \new_[12029]_ ,
    \new_[12030]_ , \new_[12034]_ , \new_[12035]_ , \new_[12036]_ ,
    \new_[12039]_ , \new_[12043]_ , \new_[12044]_ , \new_[12045]_ ,
    \new_[12049]_ , \new_[12050]_ , \new_[12054]_ , \new_[12055]_ ,
    \new_[12056]_ , \new_[12059]_ , \new_[12063]_ , \new_[12064]_ ,
    \new_[12065]_ , \new_[12069]_ , \new_[12070]_ , \new_[12074]_ ,
    \new_[12075]_ , \new_[12076]_ , \new_[12079]_ , \new_[12083]_ ,
    \new_[12084]_ , \new_[12085]_ , \new_[12089]_ , \new_[12090]_ ,
    \new_[12094]_ , \new_[12095]_ , \new_[12096]_ , \new_[12099]_ ,
    \new_[12103]_ , \new_[12104]_ , \new_[12105]_ , \new_[12109]_ ,
    \new_[12110]_ , \new_[12114]_ , \new_[12115]_ , \new_[12116]_ ,
    \new_[12119]_ , \new_[12123]_ , \new_[12124]_ , \new_[12125]_ ,
    \new_[12129]_ , \new_[12130]_ , \new_[12134]_ , \new_[12135]_ ,
    \new_[12136]_ , \new_[12139]_ , \new_[12143]_ , \new_[12144]_ ,
    \new_[12145]_ , \new_[12149]_ , \new_[12150]_ , \new_[12154]_ ,
    \new_[12155]_ , \new_[12156]_ , \new_[12159]_ , \new_[12163]_ ,
    \new_[12164]_ , \new_[12165]_ , \new_[12169]_ , \new_[12170]_ ,
    \new_[12174]_ , \new_[12175]_ , \new_[12176]_ , \new_[12179]_ ,
    \new_[12183]_ , \new_[12184]_ , \new_[12185]_ , \new_[12189]_ ,
    \new_[12190]_ , \new_[12194]_ , \new_[12195]_ , \new_[12196]_ ,
    \new_[12199]_ , \new_[12203]_ , \new_[12204]_ , \new_[12205]_ ,
    \new_[12209]_ , \new_[12210]_ , \new_[12214]_ , \new_[12215]_ ,
    \new_[12216]_ , \new_[12219]_ , \new_[12223]_ , \new_[12224]_ ,
    \new_[12225]_ , \new_[12229]_ , \new_[12230]_ , \new_[12234]_ ,
    \new_[12235]_ , \new_[12236]_ , \new_[12239]_ , \new_[12243]_ ,
    \new_[12244]_ , \new_[12245]_ , \new_[12249]_ , \new_[12250]_ ,
    \new_[12254]_ , \new_[12255]_ , \new_[12256]_ , \new_[12259]_ ,
    \new_[12263]_ , \new_[12264]_ , \new_[12265]_ , \new_[12269]_ ,
    \new_[12270]_ , \new_[12274]_ , \new_[12275]_ , \new_[12276]_ ,
    \new_[12279]_ , \new_[12283]_ , \new_[12284]_ , \new_[12285]_ ,
    \new_[12289]_ , \new_[12290]_ , \new_[12294]_ , \new_[12295]_ ,
    \new_[12296]_ , \new_[12299]_ , \new_[12303]_ , \new_[12304]_ ,
    \new_[12305]_ , \new_[12309]_ , \new_[12310]_ , \new_[12314]_ ,
    \new_[12315]_ , \new_[12316]_ , \new_[12319]_ , \new_[12323]_ ,
    \new_[12324]_ , \new_[12325]_ , \new_[12329]_ , \new_[12330]_ ,
    \new_[12334]_ , \new_[12335]_ , \new_[12336]_ , \new_[12339]_ ,
    \new_[12343]_ , \new_[12344]_ , \new_[12345]_ , \new_[12349]_ ,
    \new_[12350]_ , \new_[12354]_ , \new_[12355]_ , \new_[12356]_ ,
    \new_[12359]_ , \new_[12363]_ , \new_[12364]_ , \new_[12365]_ ,
    \new_[12369]_ , \new_[12370]_ , \new_[12374]_ , \new_[12375]_ ,
    \new_[12376]_ , \new_[12379]_ , \new_[12383]_ , \new_[12384]_ ,
    \new_[12385]_ , \new_[12389]_ , \new_[12390]_ , \new_[12394]_ ,
    \new_[12395]_ , \new_[12396]_ , \new_[12399]_ , \new_[12403]_ ,
    \new_[12404]_ , \new_[12405]_ , \new_[12409]_ , \new_[12410]_ ,
    \new_[12414]_ , \new_[12415]_ , \new_[12416]_ , \new_[12419]_ ,
    \new_[12423]_ , \new_[12424]_ , \new_[12425]_ , \new_[12429]_ ,
    \new_[12430]_ , \new_[12434]_ , \new_[12435]_ , \new_[12436]_ ,
    \new_[12439]_ , \new_[12443]_ , \new_[12444]_ , \new_[12445]_ ,
    \new_[12449]_ , \new_[12450]_ , \new_[12454]_ , \new_[12455]_ ,
    \new_[12456]_ , \new_[12459]_ , \new_[12463]_ , \new_[12464]_ ,
    \new_[12465]_ , \new_[12469]_ , \new_[12470]_ , \new_[12474]_ ,
    \new_[12475]_ , \new_[12476]_ , \new_[12479]_ , \new_[12483]_ ,
    \new_[12484]_ , \new_[12485]_ , \new_[12489]_ , \new_[12490]_ ,
    \new_[12494]_ , \new_[12495]_ , \new_[12496]_ , \new_[12499]_ ,
    \new_[12503]_ , \new_[12504]_ , \new_[12505]_ , \new_[12509]_ ,
    \new_[12510]_ , \new_[12514]_ , \new_[12515]_ , \new_[12516]_ ,
    \new_[12519]_ , \new_[12523]_ , \new_[12524]_ , \new_[12525]_ ,
    \new_[12529]_ , \new_[12530]_ , \new_[12534]_ , \new_[12535]_ ,
    \new_[12536]_ , \new_[12539]_ , \new_[12543]_ , \new_[12544]_ ,
    \new_[12545]_ , \new_[12549]_ , \new_[12550]_ , \new_[12554]_ ,
    \new_[12555]_ , \new_[12556]_ , \new_[12559]_ , \new_[12563]_ ,
    \new_[12564]_ , \new_[12565]_ , \new_[12569]_ , \new_[12570]_ ,
    \new_[12574]_ , \new_[12575]_ , \new_[12576]_ , \new_[12579]_ ,
    \new_[12583]_ , \new_[12584]_ , \new_[12585]_ , \new_[12589]_ ,
    \new_[12590]_ , \new_[12594]_ , \new_[12595]_ , \new_[12596]_ ,
    \new_[12599]_ , \new_[12603]_ , \new_[12604]_ , \new_[12605]_ ,
    \new_[12609]_ , \new_[12610]_ , \new_[12614]_ , \new_[12615]_ ,
    \new_[12616]_ , \new_[12619]_ , \new_[12623]_ , \new_[12624]_ ,
    \new_[12625]_ , \new_[12629]_ , \new_[12630]_ , \new_[12634]_ ,
    \new_[12635]_ , \new_[12636]_ , \new_[12639]_ , \new_[12643]_ ,
    \new_[12644]_ , \new_[12645]_ , \new_[12649]_ , \new_[12650]_ ,
    \new_[12654]_ , \new_[12655]_ , \new_[12656]_ , \new_[12659]_ ,
    \new_[12663]_ , \new_[12664]_ , \new_[12665]_ , \new_[12669]_ ,
    \new_[12670]_ , \new_[12674]_ , \new_[12675]_ , \new_[12676]_ ,
    \new_[12679]_ , \new_[12683]_ , \new_[12684]_ , \new_[12685]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12694]_ , \new_[12695]_ ,
    \new_[12696]_ , \new_[12699]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12705]_ , \new_[12709]_ , \new_[12710]_ , \new_[12714]_ ,
    \new_[12715]_ , \new_[12716]_ , \new_[12719]_ , \new_[12723]_ ,
    \new_[12724]_ , \new_[12725]_ , \new_[12729]_ , \new_[12730]_ ,
    \new_[12734]_ , \new_[12735]_ , \new_[12736]_ , \new_[12739]_ ,
    \new_[12743]_ , \new_[12744]_ , \new_[12745]_ , \new_[12749]_ ,
    \new_[12750]_ , \new_[12754]_ , \new_[12755]_ , \new_[12756]_ ,
    \new_[12759]_ , \new_[12763]_ , \new_[12764]_ , \new_[12765]_ ,
    \new_[12769]_ , \new_[12770]_ , \new_[12774]_ , \new_[12775]_ ,
    \new_[12776]_ , \new_[12779]_ , \new_[12783]_ , \new_[12784]_ ,
    \new_[12785]_ , \new_[12789]_ , \new_[12790]_ , \new_[12794]_ ,
    \new_[12795]_ , \new_[12796]_ , \new_[12799]_ , \new_[12803]_ ,
    \new_[12804]_ , \new_[12805]_ , \new_[12809]_ , \new_[12810]_ ,
    \new_[12814]_ , \new_[12815]_ , \new_[12816]_ , \new_[12819]_ ,
    \new_[12823]_ , \new_[12824]_ , \new_[12825]_ , \new_[12829]_ ,
    \new_[12830]_ , \new_[12834]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12839]_ , \new_[12843]_ , \new_[12844]_ , \new_[12845]_ ,
    \new_[12849]_ , \new_[12850]_ , \new_[12854]_ , \new_[12855]_ ,
    \new_[12856]_ , \new_[12859]_ , \new_[12863]_ , \new_[12864]_ ,
    \new_[12865]_ , \new_[12869]_ , \new_[12870]_ , \new_[12874]_ ,
    \new_[12875]_ , \new_[12876]_ , \new_[12879]_ , \new_[12883]_ ,
    \new_[12884]_ , \new_[12885]_ , \new_[12889]_ , \new_[12890]_ ,
    \new_[12894]_ , \new_[12895]_ , \new_[12896]_ , \new_[12899]_ ,
    \new_[12903]_ , \new_[12904]_ , \new_[12905]_ , \new_[12909]_ ,
    \new_[12910]_ , \new_[12914]_ , \new_[12915]_ , \new_[12916]_ ,
    \new_[12919]_ , \new_[12923]_ , \new_[12924]_ , \new_[12925]_ ,
    \new_[12929]_ , \new_[12930]_ , \new_[12934]_ , \new_[12935]_ ,
    \new_[12936]_ , \new_[12939]_ , \new_[12943]_ , \new_[12944]_ ,
    \new_[12945]_ , \new_[12949]_ , \new_[12950]_ , \new_[12954]_ ,
    \new_[12955]_ , \new_[12956]_ , \new_[12959]_ , \new_[12963]_ ,
    \new_[12964]_ , \new_[12965]_ , \new_[12969]_ , \new_[12970]_ ,
    \new_[12974]_ , \new_[12975]_ , \new_[12976]_ , \new_[12979]_ ,
    \new_[12983]_ , \new_[12984]_ , \new_[12985]_ , \new_[12989]_ ,
    \new_[12990]_ , \new_[12994]_ , \new_[12995]_ , \new_[12996]_ ,
    \new_[12999]_ , \new_[13003]_ , \new_[13004]_ , \new_[13005]_ ,
    \new_[13009]_ , \new_[13010]_ , \new_[13014]_ , \new_[13015]_ ,
    \new_[13016]_ , \new_[13019]_ , \new_[13023]_ , \new_[13024]_ ,
    \new_[13025]_ , \new_[13029]_ , \new_[13030]_ , \new_[13034]_ ,
    \new_[13035]_ , \new_[13036]_ , \new_[13039]_ , \new_[13043]_ ,
    \new_[13044]_ , \new_[13045]_ , \new_[13049]_ , \new_[13050]_ ,
    \new_[13054]_ , \new_[13055]_ , \new_[13056]_ , \new_[13059]_ ,
    \new_[13063]_ , \new_[13064]_ , \new_[13065]_ , \new_[13069]_ ,
    \new_[13070]_ , \new_[13074]_ , \new_[13075]_ , \new_[13076]_ ,
    \new_[13079]_ , \new_[13083]_ , \new_[13084]_ , \new_[13085]_ ,
    \new_[13089]_ , \new_[13090]_ , \new_[13094]_ , \new_[13095]_ ,
    \new_[13096]_ , \new_[13099]_ , \new_[13103]_ , \new_[13104]_ ,
    \new_[13105]_ , \new_[13109]_ , \new_[13110]_ , \new_[13114]_ ,
    \new_[13115]_ , \new_[13116]_ , \new_[13119]_ , \new_[13123]_ ,
    \new_[13124]_ , \new_[13125]_ , \new_[13129]_ , \new_[13130]_ ,
    \new_[13134]_ , \new_[13135]_ , \new_[13136]_ , \new_[13139]_ ,
    \new_[13143]_ , \new_[13144]_ , \new_[13145]_ , \new_[13149]_ ,
    \new_[13150]_ , \new_[13154]_ , \new_[13155]_ , \new_[13156]_ ,
    \new_[13159]_ , \new_[13163]_ , \new_[13164]_ , \new_[13165]_ ,
    \new_[13169]_ , \new_[13170]_ , \new_[13174]_ , \new_[13175]_ ,
    \new_[13176]_ , \new_[13179]_ , \new_[13183]_ , \new_[13184]_ ,
    \new_[13185]_ , \new_[13189]_ , \new_[13190]_ , \new_[13194]_ ,
    \new_[13195]_ , \new_[13196]_ , \new_[13199]_ , \new_[13203]_ ,
    \new_[13204]_ , \new_[13205]_ , \new_[13209]_ , \new_[13210]_ ,
    \new_[13214]_ , \new_[13215]_ , \new_[13216]_ , \new_[13219]_ ,
    \new_[13223]_ , \new_[13224]_ , \new_[13225]_ , \new_[13229]_ ,
    \new_[13230]_ , \new_[13234]_ , \new_[13235]_ , \new_[13236]_ ,
    \new_[13239]_ , \new_[13243]_ , \new_[13244]_ , \new_[13245]_ ,
    \new_[13249]_ , \new_[13250]_ , \new_[13254]_ , \new_[13255]_ ,
    \new_[13256]_ , \new_[13259]_ , \new_[13263]_ , \new_[13264]_ ,
    \new_[13265]_ , \new_[13269]_ , \new_[13270]_ , \new_[13274]_ ,
    \new_[13275]_ , \new_[13276]_ , \new_[13279]_ , \new_[13283]_ ,
    \new_[13284]_ , \new_[13285]_ , \new_[13289]_ , \new_[13290]_ ,
    \new_[13294]_ , \new_[13295]_ , \new_[13296]_ , \new_[13299]_ ,
    \new_[13303]_ , \new_[13304]_ , \new_[13305]_ , \new_[13309]_ ,
    \new_[13310]_ , \new_[13314]_ , \new_[13315]_ , \new_[13316]_ ,
    \new_[13319]_ , \new_[13323]_ , \new_[13324]_ , \new_[13325]_ ,
    \new_[13329]_ , \new_[13330]_ , \new_[13334]_ , \new_[13335]_ ,
    \new_[13336]_ , \new_[13339]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13345]_ , \new_[13349]_ , \new_[13350]_ , \new_[13354]_ ,
    \new_[13355]_ , \new_[13356]_ , \new_[13359]_ , \new_[13363]_ ,
    \new_[13364]_ , \new_[13365]_ , \new_[13369]_ , \new_[13370]_ ,
    \new_[13374]_ , \new_[13375]_ , \new_[13376]_ , \new_[13379]_ ,
    \new_[13383]_ , \new_[13384]_ , \new_[13385]_ , \new_[13389]_ ,
    \new_[13390]_ , \new_[13394]_ , \new_[13395]_ , \new_[13396]_ ,
    \new_[13399]_ , \new_[13403]_ , \new_[13404]_ , \new_[13405]_ ,
    \new_[13409]_ , \new_[13410]_ , \new_[13414]_ , \new_[13415]_ ,
    \new_[13416]_ , \new_[13419]_ , \new_[13423]_ , \new_[13424]_ ,
    \new_[13425]_ , \new_[13429]_ , \new_[13430]_ , \new_[13434]_ ,
    \new_[13435]_ , \new_[13436]_ , \new_[13439]_ , \new_[13443]_ ,
    \new_[13444]_ , \new_[13445]_ , \new_[13449]_ , \new_[13450]_ ,
    \new_[13454]_ , \new_[13455]_ , \new_[13456]_ , \new_[13459]_ ,
    \new_[13463]_ , \new_[13464]_ , \new_[13465]_ , \new_[13469]_ ,
    \new_[13470]_ , \new_[13474]_ , \new_[13475]_ , \new_[13476]_ ,
    \new_[13479]_ , \new_[13483]_ , \new_[13484]_ , \new_[13485]_ ,
    \new_[13489]_ , \new_[13490]_ , \new_[13494]_ , \new_[13495]_ ,
    \new_[13496]_ , \new_[13499]_ , \new_[13503]_ , \new_[13504]_ ,
    \new_[13505]_ , \new_[13509]_ , \new_[13510]_ , \new_[13514]_ ,
    \new_[13515]_ , \new_[13516]_ , \new_[13519]_ , \new_[13523]_ ,
    \new_[13524]_ , \new_[13525]_ , \new_[13529]_ , \new_[13530]_ ,
    \new_[13534]_ , \new_[13535]_ , \new_[13536]_ , \new_[13539]_ ,
    \new_[13543]_ , \new_[13544]_ , \new_[13545]_ , \new_[13549]_ ,
    \new_[13550]_ , \new_[13554]_ , \new_[13555]_ , \new_[13556]_ ,
    \new_[13559]_ , \new_[13563]_ , \new_[13564]_ , \new_[13565]_ ,
    \new_[13569]_ , \new_[13570]_ , \new_[13574]_ , \new_[13575]_ ,
    \new_[13576]_ , \new_[13579]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13589]_ , \new_[13590]_ , \new_[13594]_ ,
    \new_[13595]_ , \new_[13596]_ , \new_[13599]_ , \new_[13603]_ ,
    \new_[13604]_ , \new_[13605]_ , \new_[13609]_ , \new_[13610]_ ,
    \new_[13614]_ , \new_[13615]_ , \new_[13616]_ , \new_[13619]_ ,
    \new_[13623]_ , \new_[13624]_ , \new_[13625]_ , \new_[13629]_ ,
    \new_[13630]_ , \new_[13634]_ , \new_[13635]_ , \new_[13636]_ ,
    \new_[13639]_ , \new_[13643]_ , \new_[13644]_ , \new_[13645]_ ,
    \new_[13649]_ , \new_[13650]_ , \new_[13654]_ , \new_[13655]_ ,
    \new_[13656]_ , \new_[13659]_ , \new_[13663]_ , \new_[13664]_ ,
    \new_[13665]_ , \new_[13669]_ , \new_[13670]_ , \new_[13674]_ ,
    \new_[13675]_ , \new_[13676]_ , \new_[13679]_ , \new_[13683]_ ,
    \new_[13684]_ , \new_[13685]_ , \new_[13689]_ , \new_[13690]_ ,
    \new_[13694]_ , \new_[13695]_ , \new_[13696]_ , \new_[13699]_ ,
    \new_[13703]_ , \new_[13704]_ , \new_[13705]_ , \new_[13709]_ ,
    \new_[13710]_ , \new_[13714]_ , \new_[13715]_ , \new_[13716]_ ,
    \new_[13719]_ , \new_[13723]_ , \new_[13724]_ , \new_[13725]_ ,
    \new_[13729]_ , \new_[13730]_ , \new_[13734]_ , \new_[13735]_ ,
    \new_[13736]_ , \new_[13739]_ , \new_[13743]_ , \new_[13744]_ ,
    \new_[13745]_ , \new_[13749]_ , \new_[13750]_ , \new_[13754]_ ,
    \new_[13755]_ , \new_[13756]_ , \new_[13759]_ , \new_[13763]_ ,
    \new_[13764]_ , \new_[13765]_ , \new_[13769]_ , \new_[13770]_ ,
    \new_[13774]_ , \new_[13775]_ , \new_[13776]_ , \new_[13779]_ ,
    \new_[13783]_ , \new_[13784]_ , \new_[13785]_ , \new_[13789]_ ,
    \new_[13790]_ , \new_[13794]_ , \new_[13795]_ , \new_[13796]_ ,
    \new_[13799]_ , \new_[13803]_ , \new_[13804]_ , \new_[13805]_ ,
    \new_[13809]_ , \new_[13810]_ , \new_[13814]_ , \new_[13815]_ ,
    \new_[13816]_ , \new_[13819]_ , \new_[13823]_ , \new_[13824]_ ,
    \new_[13825]_ , \new_[13829]_ , \new_[13830]_ , \new_[13834]_ ,
    \new_[13835]_ , \new_[13836]_ , \new_[13839]_ , \new_[13843]_ ,
    \new_[13844]_ , \new_[13845]_ , \new_[13849]_ , \new_[13850]_ ,
    \new_[13854]_ , \new_[13855]_ , \new_[13856]_ , \new_[13859]_ ,
    \new_[13863]_ , \new_[13864]_ , \new_[13865]_ , \new_[13869]_ ,
    \new_[13870]_ , \new_[13874]_ , \new_[13875]_ , \new_[13876]_ ,
    \new_[13879]_ , \new_[13883]_ , \new_[13884]_ , \new_[13885]_ ,
    \new_[13889]_ , \new_[13890]_ , \new_[13894]_ , \new_[13895]_ ,
    \new_[13896]_ , \new_[13899]_ , \new_[13903]_ , \new_[13904]_ ,
    \new_[13905]_ , \new_[13909]_ , \new_[13910]_ , \new_[13914]_ ,
    \new_[13915]_ , \new_[13916]_ , \new_[13919]_ , \new_[13923]_ ,
    \new_[13924]_ , \new_[13925]_ , \new_[13929]_ , \new_[13930]_ ,
    \new_[13934]_ , \new_[13935]_ , \new_[13936]_ , \new_[13939]_ ,
    \new_[13943]_ , \new_[13944]_ , \new_[13945]_ , \new_[13949]_ ,
    \new_[13950]_ , \new_[13954]_ , \new_[13955]_ , \new_[13956]_ ,
    \new_[13959]_ , \new_[13963]_ , \new_[13964]_ , \new_[13965]_ ,
    \new_[13969]_ , \new_[13970]_ , \new_[13974]_ , \new_[13975]_ ,
    \new_[13976]_ , \new_[13979]_ , \new_[13983]_ , \new_[13984]_ ,
    \new_[13985]_ , \new_[13989]_ , \new_[13990]_ , \new_[13994]_ ,
    \new_[13995]_ , \new_[13996]_ , \new_[13999]_ , \new_[14003]_ ,
    \new_[14004]_ , \new_[14005]_ , \new_[14009]_ , \new_[14010]_ ,
    \new_[14014]_ , \new_[14015]_ , \new_[14016]_ , \new_[14019]_ ,
    \new_[14023]_ , \new_[14024]_ , \new_[14025]_ , \new_[14029]_ ,
    \new_[14030]_ , \new_[14034]_ , \new_[14035]_ , \new_[14036]_ ,
    \new_[14039]_ , \new_[14043]_ , \new_[14044]_ , \new_[14045]_ ,
    \new_[14049]_ , \new_[14050]_ , \new_[14054]_ , \new_[14055]_ ,
    \new_[14056]_ , \new_[14059]_ , \new_[14063]_ , \new_[14064]_ ,
    \new_[14065]_ , \new_[14069]_ , \new_[14070]_ , \new_[14074]_ ,
    \new_[14075]_ , \new_[14076]_ , \new_[14079]_ , \new_[14083]_ ,
    \new_[14084]_ , \new_[14085]_ , \new_[14089]_ , \new_[14090]_ ,
    \new_[14094]_ , \new_[14095]_ , \new_[14096]_ , \new_[14099]_ ,
    \new_[14103]_ , \new_[14104]_ , \new_[14105]_ , \new_[14109]_ ,
    \new_[14110]_ , \new_[14114]_ , \new_[14115]_ , \new_[14116]_ ,
    \new_[14119]_ , \new_[14123]_ , \new_[14124]_ , \new_[14125]_ ,
    \new_[14129]_ , \new_[14130]_ , \new_[14134]_ , \new_[14135]_ ,
    \new_[14136]_ , \new_[14139]_ , \new_[14143]_ , \new_[14144]_ ,
    \new_[14145]_ , \new_[14149]_ , \new_[14150]_ , \new_[14154]_ ,
    \new_[14155]_ , \new_[14156]_ , \new_[14159]_ , \new_[14163]_ ,
    \new_[14164]_ , \new_[14165]_ , \new_[14169]_ , \new_[14170]_ ,
    \new_[14174]_ , \new_[14175]_ , \new_[14176]_ , \new_[14179]_ ,
    \new_[14183]_ , \new_[14184]_ , \new_[14185]_ , \new_[14189]_ ,
    \new_[14190]_ , \new_[14194]_ , \new_[14195]_ , \new_[14196]_ ,
    \new_[14199]_ , \new_[14203]_ , \new_[14204]_ , \new_[14205]_ ,
    \new_[14209]_ , \new_[14210]_ , \new_[14214]_ , \new_[14215]_ ,
    \new_[14216]_ , \new_[14219]_ , \new_[14223]_ , \new_[14224]_ ,
    \new_[14225]_ , \new_[14229]_ , \new_[14230]_ , \new_[14234]_ ,
    \new_[14235]_ , \new_[14236]_ , \new_[14239]_ , \new_[14243]_ ,
    \new_[14244]_ , \new_[14245]_ , \new_[14249]_ , \new_[14250]_ ,
    \new_[14254]_ , \new_[14255]_ , \new_[14256]_ , \new_[14259]_ ,
    \new_[14263]_ , \new_[14264]_ , \new_[14265]_ , \new_[14269]_ ,
    \new_[14270]_ , \new_[14274]_ , \new_[14275]_ , \new_[14276]_ ,
    \new_[14279]_ , \new_[14283]_ , \new_[14284]_ , \new_[14285]_ ,
    \new_[14289]_ , \new_[14290]_ , \new_[14294]_ , \new_[14295]_ ,
    \new_[14296]_ , \new_[14299]_ , \new_[14303]_ , \new_[14304]_ ,
    \new_[14305]_ , \new_[14309]_ , \new_[14310]_ , \new_[14314]_ ,
    \new_[14315]_ , \new_[14316]_ , \new_[14319]_ , \new_[14323]_ ,
    \new_[14324]_ , \new_[14325]_ , \new_[14329]_ , \new_[14330]_ ,
    \new_[14334]_ , \new_[14335]_ , \new_[14336]_ , \new_[14339]_ ,
    \new_[14343]_ , \new_[14344]_ , \new_[14345]_ , \new_[14349]_ ,
    \new_[14350]_ , \new_[14354]_ , \new_[14355]_ , \new_[14356]_ ,
    \new_[14359]_ , \new_[14363]_ , \new_[14364]_ , \new_[14365]_ ,
    \new_[14369]_ , \new_[14370]_ , \new_[14374]_ , \new_[14375]_ ,
    \new_[14376]_ , \new_[14379]_ , \new_[14383]_ , \new_[14384]_ ,
    \new_[14385]_ , \new_[14389]_ , \new_[14390]_ , \new_[14394]_ ,
    \new_[14395]_ , \new_[14396]_ , \new_[14399]_ , \new_[14403]_ ,
    \new_[14404]_ , \new_[14405]_ , \new_[14409]_ , \new_[14410]_ ,
    \new_[14414]_ , \new_[14415]_ , \new_[14416]_ , \new_[14419]_ ,
    \new_[14423]_ , \new_[14424]_ , \new_[14425]_ , \new_[14429]_ ,
    \new_[14430]_ , \new_[14434]_ , \new_[14435]_ , \new_[14436]_ ,
    \new_[14439]_ , \new_[14443]_ , \new_[14444]_ , \new_[14445]_ ,
    \new_[14449]_ , \new_[14450]_ , \new_[14454]_ , \new_[14455]_ ,
    \new_[14456]_ , \new_[14459]_ , \new_[14463]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14469]_ , \new_[14470]_ , \new_[14474]_ ,
    \new_[14475]_ , \new_[14476]_ , \new_[14479]_ , \new_[14483]_ ,
    \new_[14484]_ , \new_[14485]_ , \new_[14489]_ , \new_[14490]_ ,
    \new_[14494]_ , \new_[14495]_ , \new_[14496]_ , \new_[14499]_ ,
    \new_[14503]_ , \new_[14504]_ , \new_[14505]_ , \new_[14509]_ ,
    \new_[14510]_ , \new_[14514]_ , \new_[14515]_ , \new_[14516]_ ,
    \new_[14519]_ , \new_[14523]_ , \new_[14524]_ , \new_[14525]_ ,
    \new_[14529]_ , \new_[14530]_ , \new_[14534]_ , \new_[14535]_ ,
    \new_[14536]_ , \new_[14539]_ , \new_[14543]_ , \new_[14544]_ ,
    \new_[14545]_ , \new_[14549]_ , \new_[14550]_ , \new_[14554]_ ,
    \new_[14555]_ , \new_[14556]_ , \new_[14559]_ , \new_[14563]_ ,
    \new_[14564]_ , \new_[14565]_ , \new_[14569]_ , \new_[14570]_ ,
    \new_[14574]_ , \new_[14575]_ , \new_[14576]_ , \new_[14579]_ ,
    \new_[14583]_ , \new_[14584]_ , \new_[14585]_ , \new_[14589]_ ,
    \new_[14590]_ , \new_[14594]_ , \new_[14595]_ , \new_[14596]_ ,
    \new_[14599]_ , \new_[14603]_ , \new_[14604]_ , \new_[14605]_ ,
    \new_[14609]_ , \new_[14610]_ , \new_[14614]_ , \new_[14615]_ ,
    \new_[14616]_ , \new_[14619]_ , \new_[14623]_ , \new_[14624]_ ,
    \new_[14625]_ , \new_[14629]_ , \new_[14630]_ , \new_[14634]_ ,
    \new_[14635]_ , \new_[14636]_ , \new_[14639]_ , \new_[14643]_ ,
    \new_[14644]_ , \new_[14645]_ , \new_[14649]_ , \new_[14650]_ ,
    \new_[14654]_ , \new_[14655]_ , \new_[14656]_ , \new_[14659]_ ,
    \new_[14663]_ , \new_[14664]_ , \new_[14665]_ , \new_[14669]_ ,
    \new_[14670]_ , \new_[14674]_ , \new_[14675]_ , \new_[14676]_ ,
    \new_[14679]_ , \new_[14683]_ , \new_[14684]_ , \new_[14685]_ ,
    \new_[14689]_ , \new_[14690]_ , \new_[14694]_ , \new_[14695]_ ,
    \new_[14696]_ , \new_[14699]_ , \new_[14703]_ , \new_[14704]_ ,
    \new_[14705]_ , \new_[14709]_ , \new_[14710]_ , \new_[14714]_ ,
    \new_[14715]_ , \new_[14716]_ , \new_[14719]_ , \new_[14723]_ ,
    \new_[14724]_ , \new_[14725]_ , \new_[14729]_ , \new_[14730]_ ,
    \new_[14734]_ , \new_[14735]_ , \new_[14736]_ , \new_[14739]_ ,
    \new_[14743]_ , \new_[14744]_ , \new_[14745]_ , \new_[14749]_ ,
    \new_[14750]_ , \new_[14754]_ , \new_[14755]_ , \new_[14756]_ ,
    \new_[14759]_ , \new_[14763]_ , \new_[14764]_ , \new_[14765]_ ,
    \new_[14769]_ , \new_[14770]_ , \new_[14774]_ , \new_[14775]_ ,
    \new_[14776]_ , \new_[14779]_ , \new_[14783]_ , \new_[14784]_ ,
    \new_[14785]_ , \new_[14789]_ , \new_[14790]_ , \new_[14794]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14799]_ , \new_[14803]_ ,
    \new_[14804]_ , \new_[14805]_ , \new_[14809]_ , \new_[14810]_ ,
    \new_[14814]_ , \new_[14815]_ , \new_[14816]_ , \new_[14819]_ ,
    \new_[14823]_ , \new_[14824]_ , \new_[14825]_ , \new_[14829]_ ,
    \new_[14830]_ , \new_[14834]_ , \new_[14835]_ , \new_[14836]_ ,
    \new_[14839]_ , \new_[14843]_ , \new_[14844]_ , \new_[14845]_ ,
    \new_[14849]_ , \new_[14850]_ , \new_[14854]_ , \new_[14855]_ ,
    \new_[14856]_ , \new_[14859]_ , \new_[14863]_ , \new_[14864]_ ,
    \new_[14865]_ , \new_[14869]_ , \new_[14870]_ , \new_[14874]_ ,
    \new_[14875]_ , \new_[14876]_ , \new_[14879]_ , \new_[14883]_ ,
    \new_[14884]_ , \new_[14885]_ , \new_[14889]_ , \new_[14890]_ ,
    \new_[14894]_ , \new_[14895]_ , \new_[14896]_ , \new_[14899]_ ,
    \new_[14903]_ , \new_[14904]_ , \new_[14905]_ , \new_[14909]_ ,
    \new_[14910]_ , \new_[14914]_ , \new_[14915]_ , \new_[14916]_ ,
    \new_[14919]_ , \new_[14923]_ , \new_[14924]_ , \new_[14925]_ ,
    \new_[14929]_ , \new_[14930]_ , \new_[14934]_ , \new_[14935]_ ,
    \new_[14936]_ , \new_[14940]_ , \new_[14941]_ , \new_[14945]_ ,
    \new_[14946]_ , \new_[14947]_ , \new_[14951]_ , \new_[14952]_ ,
    \new_[14956]_ , \new_[14957]_ , \new_[14958]_ , \new_[14962]_ ,
    \new_[14963]_ , \new_[14967]_ , \new_[14968]_ , \new_[14969]_ ,
    \new_[14973]_ , \new_[14974]_ , \new_[14978]_ , \new_[14979]_ ,
    \new_[14980]_ , \new_[14984]_ , \new_[14985]_ , \new_[14989]_ ,
    \new_[14990]_ , \new_[14991]_ , \new_[14995]_ , \new_[14996]_ ,
    \new_[15000]_ , \new_[15001]_ , \new_[15002]_ , \new_[15006]_ ,
    \new_[15007]_ , \new_[15011]_ , \new_[15012]_ , \new_[15013]_ ,
    \new_[15017]_ , \new_[15018]_ , \new_[15022]_ , \new_[15023]_ ,
    \new_[15024]_ , \new_[15028]_ , \new_[15029]_ , \new_[15033]_ ,
    \new_[15034]_ , \new_[15035]_ , \new_[15039]_ , \new_[15040]_ ,
    \new_[15044]_ , \new_[15045]_ , \new_[15046]_ , \new_[15050]_ ,
    \new_[15051]_ , \new_[15055]_ , \new_[15056]_ , \new_[15057]_ ,
    \new_[15061]_ , \new_[15062]_ , \new_[15066]_ , \new_[15067]_ ,
    \new_[15068]_ , \new_[15072]_ , \new_[15073]_ , \new_[15077]_ ,
    \new_[15078]_ , \new_[15079]_ , \new_[15083]_ , \new_[15084]_ ,
    \new_[15088]_ , \new_[15089]_ , \new_[15090]_ , \new_[15094]_ ,
    \new_[15095]_ , \new_[15099]_ , \new_[15100]_ , \new_[15101]_ ,
    \new_[15105]_ , \new_[15106]_ , \new_[15110]_ , \new_[15111]_ ,
    \new_[15112]_ , \new_[15116]_ , \new_[15117]_ , \new_[15121]_ ,
    \new_[15122]_ , \new_[15123]_ , \new_[15127]_ , \new_[15128]_ ,
    \new_[15132]_ , \new_[15133]_ , \new_[15134]_ , \new_[15138]_ ,
    \new_[15139]_ , \new_[15143]_ , \new_[15144]_ , \new_[15145]_ ,
    \new_[15149]_ , \new_[15150]_ , \new_[15154]_ , \new_[15155]_ ,
    \new_[15156]_ , \new_[15160]_ , \new_[15161]_ , \new_[15165]_ ,
    \new_[15166]_ , \new_[15167]_ , \new_[15171]_ , \new_[15172]_ ,
    \new_[15176]_ , \new_[15177]_ , \new_[15178]_ , \new_[15182]_ ,
    \new_[15183]_ , \new_[15187]_ , \new_[15188]_ , \new_[15189]_ ,
    \new_[15193]_ , \new_[15194]_ , \new_[15198]_ , \new_[15199]_ ,
    \new_[15200]_ , \new_[15204]_ , \new_[15205]_ , \new_[15209]_ ,
    \new_[15210]_ , \new_[15211]_ , \new_[15215]_ , \new_[15216]_ ,
    \new_[15220]_ , \new_[15221]_ , \new_[15222]_ , \new_[15226]_ ,
    \new_[15227]_ , \new_[15231]_ , \new_[15232]_ , \new_[15233]_ ,
    \new_[15237]_ , \new_[15238]_ , \new_[15242]_ , \new_[15243]_ ,
    \new_[15244]_ , \new_[15248]_ , \new_[15249]_ , \new_[15253]_ ,
    \new_[15254]_ , \new_[15255]_ , \new_[15259]_ , \new_[15260]_ ,
    \new_[15264]_ , \new_[15265]_ , \new_[15266]_ , \new_[15270]_ ,
    \new_[15271]_ , \new_[15275]_ , \new_[15276]_ , \new_[15277]_ ,
    \new_[15281]_ , \new_[15282]_ , \new_[15286]_ , \new_[15287]_ ,
    \new_[15288]_ , \new_[15292]_ , \new_[15293]_ , \new_[15297]_ ,
    \new_[15298]_ , \new_[15299]_ , \new_[15303]_ , \new_[15304]_ ,
    \new_[15308]_ , \new_[15309]_ , \new_[15310]_ , \new_[15314]_ ,
    \new_[15315]_ , \new_[15319]_ , \new_[15320]_ , \new_[15321]_ ,
    \new_[15325]_ , \new_[15326]_ , \new_[15330]_ , \new_[15331]_ ,
    \new_[15332]_ , \new_[15336]_ , \new_[15337]_ , \new_[15341]_ ,
    \new_[15342]_ , \new_[15343]_ , \new_[15347]_ , \new_[15348]_ ,
    \new_[15352]_ , \new_[15353]_ , \new_[15354]_ , \new_[15358]_ ,
    \new_[15359]_ , \new_[15363]_ , \new_[15364]_ , \new_[15365]_ ,
    \new_[15369]_ , \new_[15370]_ , \new_[15374]_ , \new_[15375]_ ,
    \new_[15376]_ , \new_[15380]_ , \new_[15381]_ , \new_[15385]_ ,
    \new_[15386]_ , \new_[15387]_ , \new_[15391]_ , \new_[15392]_ ,
    \new_[15396]_ , \new_[15397]_ , \new_[15398]_ , \new_[15402]_ ,
    \new_[15403]_ , \new_[15407]_ , \new_[15408]_ , \new_[15409]_ ,
    \new_[15413]_ , \new_[15414]_ , \new_[15418]_ , \new_[15419]_ ,
    \new_[15420]_ , \new_[15424]_ , \new_[15425]_ , \new_[15429]_ ,
    \new_[15430]_ , \new_[15431]_ , \new_[15435]_ , \new_[15436]_ ,
    \new_[15440]_ , \new_[15441]_ , \new_[15442]_ , \new_[15446]_ ,
    \new_[15447]_ , \new_[15451]_ , \new_[15452]_ , \new_[15453]_ ,
    \new_[15457]_ , \new_[15458]_ , \new_[15462]_ , \new_[15463]_ ,
    \new_[15464]_ , \new_[15468]_ , \new_[15469]_ , \new_[15473]_ ,
    \new_[15474]_ , \new_[15475]_ , \new_[15479]_ , \new_[15480]_ ,
    \new_[15484]_ , \new_[15485]_ , \new_[15486]_ , \new_[15490]_ ,
    \new_[15491]_ , \new_[15495]_ , \new_[15496]_ , \new_[15497]_ ,
    \new_[15501]_ , \new_[15502]_ , \new_[15506]_ , \new_[15507]_ ,
    \new_[15508]_ , \new_[15512]_ , \new_[15513]_ , \new_[15517]_ ,
    \new_[15518]_ , \new_[15519]_ , \new_[15523]_ , \new_[15524]_ ,
    \new_[15528]_ , \new_[15529]_ , \new_[15530]_ , \new_[15534]_ ,
    \new_[15535]_ , \new_[15539]_ , \new_[15540]_ , \new_[15541]_ ,
    \new_[15545]_ , \new_[15546]_ , \new_[15550]_ , \new_[15551]_ ,
    \new_[15552]_ , \new_[15556]_ , \new_[15557]_ , \new_[15561]_ ,
    \new_[15562]_ , \new_[15563]_ , \new_[15567]_ , \new_[15568]_ ,
    \new_[15572]_ , \new_[15573]_ , \new_[15574]_ , \new_[15578]_ ,
    \new_[15579]_ , \new_[15583]_ , \new_[15584]_ , \new_[15585]_ ,
    \new_[15589]_ , \new_[15590]_ , \new_[15594]_ , \new_[15595]_ ,
    \new_[15596]_ , \new_[15600]_ , \new_[15601]_ , \new_[15605]_ ,
    \new_[15606]_ , \new_[15607]_ , \new_[15611]_ , \new_[15612]_ ,
    \new_[15616]_ , \new_[15617]_ , \new_[15618]_ , \new_[15622]_ ,
    \new_[15623]_ , \new_[15627]_ , \new_[15628]_ , \new_[15629]_ ,
    \new_[15633]_ , \new_[15634]_ , \new_[15638]_ , \new_[15639]_ ,
    \new_[15640]_ , \new_[15644]_ , \new_[15645]_ , \new_[15649]_ ,
    \new_[15650]_ , \new_[15651]_ , \new_[15655]_ , \new_[15656]_ ,
    \new_[15660]_ , \new_[15661]_ , \new_[15662]_ , \new_[15666]_ ,
    \new_[15667]_ , \new_[15671]_ , \new_[15672]_ , \new_[15673]_ ,
    \new_[15677]_ , \new_[15678]_ , \new_[15682]_ , \new_[15683]_ ,
    \new_[15684]_ , \new_[15688]_ , \new_[15689]_ , \new_[15693]_ ,
    \new_[15694]_ , \new_[15695]_ , \new_[15699]_ , \new_[15700]_ ,
    \new_[15704]_ , \new_[15705]_ , \new_[15706]_ , \new_[15710]_ ,
    \new_[15711]_ , \new_[15715]_ , \new_[15716]_ , \new_[15717]_ ,
    \new_[15721]_ , \new_[15722]_ , \new_[15726]_ , \new_[15727]_ ,
    \new_[15728]_ , \new_[15732]_ , \new_[15733]_ , \new_[15737]_ ,
    \new_[15738]_ , \new_[15739]_ , \new_[15743]_ , \new_[15744]_ ,
    \new_[15748]_ , \new_[15749]_ , \new_[15750]_ , \new_[15754]_ ,
    \new_[15755]_ , \new_[15759]_ , \new_[15760]_ , \new_[15761]_ ,
    \new_[15765]_ , \new_[15766]_ , \new_[15770]_ , \new_[15771]_ ,
    \new_[15772]_ , \new_[15776]_ , \new_[15777]_ , \new_[15781]_ ,
    \new_[15782]_ , \new_[15783]_ , \new_[15787]_ , \new_[15788]_ ,
    \new_[15792]_ , \new_[15793]_ , \new_[15794]_ , \new_[15798]_ ,
    \new_[15799]_ , \new_[15803]_ , \new_[15804]_ , \new_[15805]_ ,
    \new_[15809]_ , \new_[15810]_ , \new_[15814]_ , \new_[15815]_ ,
    \new_[15816]_ , \new_[15820]_ , \new_[15821]_ , \new_[15825]_ ,
    \new_[15826]_ , \new_[15827]_ , \new_[15831]_ , \new_[15832]_ ,
    \new_[15836]_ , \new_[15837]_ , \new_[15838]_ , \new_[15842]_ ,
    \new_[15843]_ , \new_[15847]_ , \new_[15848]_ , \new_[15849]_ ,
    \new_[15853]_ , \new_[15854]_ , \new_[15858]_ , \new_[15859]_ ,
    \new_[15860]_ , \new_[15864]_ , \new_[15865]_ , \new_[15869]_ ,
    \new_[15870]_ , \new_[15871]_ , \new_[15875]_ , \new_[15876]_ ,
    \new_[15880]_ , \new_[15881]_ , \new_[15882]_ , \new_[15886]_ ,
    \new_[15887]_ , \new_[15891]_ , \new_[15892]_ , \new_[15893]_ ,
    \new_[15897]_ , \new_[15898]_ , \new_[15902]_ , \new_[15903]_ ,
    \new_[15904]_ , \new_[15908]_ , \new_[15909]_ , \new_[15913]_ ,
    \new_[15914]_ , \new_[15915]_ , \new_[15919]_ , \new_[15920]_ ,
    \new_[15924]_ , \new_[15925]_ , \new_[15926]_ , \new_[15930]_ ,
    \new_[15931]_ , \new_[15935]_ , \new_[15936]_ , \new_[15937]_ ,
    \new_[15941]_ , \new_[15942]_ , \new_[15946]_ , \new_[15947]_ ,
    \new_[15948]_ , \new_[15952]_ , \new_[15953]_ , \new_[15957]_ ,
    \new_[15958]_ , \new_[15959]_ , \new_[15963]_ , \new_[15964]_ ,
    \new_[15968]_ , \new_[15969]_ , \new_[15970]_ , \new_[15974]_ ,
    \new_[15975]_ , \new_[15979]_ , \new_[15980]_ , \new_[15981]_ ,
    \new_[15985]_ , \new_[15986]_ , \new_[15990]_ , \new_[15991]_ ,
    \new_[15992]_ , \new_[15996]_ , \new_[15997]_ , \new_[16001]_ ,
    \new_[16002]_ , \new_[16003]_ , \new_[16007]_ , \new_[16008]_ ,
    \new_[16012]_ , \new_[16013]_ , \new_[16014]_ , \new_[16018]_ ,
    \new_[16019]_ , \new_[16023]_ , \new_[16024]_ , \new_[16025]_ ,
    \new_[16029]_ , \new_[16030]_ , \new_[16034]_ , \new_[16035]_ ,
    \new_[16036]_ , \new_[16040]_ , \new_[16041]_ , \new_[16045]_ ,
    \new_[16046]_ , \new_[16047]_ , \new_[16051]_ , \new_[16052]_ ,
    \new_[16056]_ , \new_[16057]_ , \new_[16058]_ , \new_[16062]_ ,
    \new_[16063]_ , \new_[16067]_ , \new_[16068]_ , \new_[16069]_ ,
    \new_[16073]_ , \new_[16074]_ , \new_[16078]_ , \new_[16079]_ ,
    \new_[16080]_ , \new_[16084]_ , \new_[16085]_ , \new_[16089]_ ,
    \new_[16090]_ , \new_[16091]_ , \new_[16095]_ , \new_[16096]_ ,
    \new_[16100]_ , \new_[16101]_ , \new_[16102]_ , \new_[16106]_ ,
    \new_[16107]_ , \new_[16111]_ , \new_[16112]_ , \new_[16113]_ ,
    \new_[16117]_ , \new_[16118]_ , \new_[16122]_ , \new_[16123]_ ,
    \new_[16124]_ , \new_[16128]_ , \new_[16129]_ , \new_[16133]_ ,
    \new_[16134]_ , \new_[16135]_ , \new_[16139]_ , \new_[16140]_ ,
    \new_[16144]_ , \new_[16145]_ , \new_[16146]_ , \new_[16150]_ ,
    \new_[16151]_ , \new_[16155]_ , \new_[16156]_ , \new_[16157]_ ,
    \new_[16161]_ , \new_[16162]_ , \new_[16166]_ , \new_[16167]_ ,
    \new_[16168]_ , \new_[16172]_ , \new_[16173]_ , \new_[16177]_ ,
    \new_[16178]_ , \new_[16179]_ , \new_[16183]_ , \new_[16184]_ ,
    \new_[16188]_ , \new_[16189]_ , \new_[16190]_ , \new_[16194]_ ,
    \new_[16195]_ , \new_[16199]_ , \new_[16200]_ , \new_[16201]_ ,
    \new_[16205]_ , \new_[16206]_ , \new_[16210]_ , \new_[16211]_ ,
    \new_[16212]_ , \new_[16216]_ , \new_[16217]_ , \new_[16221]_ ,
    \new_[16222]_ , \new_[16223]_ , \new_[16227]_ , \new_[16228]_ ,
    \new_[16232]_ , \new_[16233]_ , \new_[16234]_ , \new_[16238]_ ,
    \new_[16239]_ , \new_[16243]_ , \new_[16244]_ , \new_[16245]_ ,
    \new_[16249]_ , \new_[16250]_ , \new_[16254]_ , \new_[16255]_ ,
    \new_[16256]_ , \new_[16260]_ , \new_[16261]_ , \new_[16265]_ ,
    \new_[16266]_ , \new_[16267]_ , \new_[16271]_ , \new_[16272]_ ,
    \new_[16276]_ , \new_[16277]_ , \new_[16278]_ , \new_[16282]_ ,
    \new_[16283]_ , \new_[16287]_ , \new_[16288]_ , \new_[16289]_ ,
    \new_[16293]_ , \new_[16294]_ , \new_[16298]_ , \new_[16299]_ ,
    \new_[16300]_ , \new_[16304]_ , \new_[16305]_ , \new_[16309]_ ,
    \new_[16310]_ , \new_[16311]_ , \new_[16315]_ , \new_[16316]_ ,
    \new_[16320]_ , \new_[16321]_ , \new_[16322]_ , \new_[16326]_ ,
    \new_[16327]_ , \new_[16331]_ , \new_[16332]_ , \new_[16333]_ ,
    \new_[16337]_ , \new_[16338]_ , \new_[16342]_ , \new_[16343]_ ,
    \new_[16344]_ , \new_[16348]_ , \new_[16349]_ , \new_[16353]_ ,
    \new_[16354]_ , \new_[16355]_ , \new_[16359]_ , \new_[16360]_ ,
    \new_[16364]_ , \new_[16365]_ , \new_[16366]_ , \new_[16370]_ ,
    \new_[16371]_ , \new_[16375]_ , \new_[16376]_ , \new_[16377]_ ,
    \new_[16381]_ , \new_[16382]_ , \new_[16386]_ , \new_[16387]_ ,
    \new_[16388]_ , \new_[16392]_ , \new_[16393]_ , \new_[16397]_ ,
    \new_[16398]_ , \new_[16399]_ , \new_[16403]_ , \new_[16404]_ ,
    \new_[16408]_ , \new_[16409]_ , \new_[16410]_ , \new_[16414]_ ,
    \new_[16415]_ , \new_[16419]_ , \new_[16420]_ , \new_[16421]_ ,
    \new_[16425]_ , \new_[16426]_ , \new_[16430]_ , \new_[16431]_ ,
    \new_[16432]_ , \new_[16436]_ , \new_[16437]_ , \new_[16441]_ ,
    \new_[16442]_ , \new_[16443]_ , \new_[16447]_ , \new_[16448]_ ,
    \new_[16452]_ , \new_[16453]_ , \new_[16454]_ , \new_[16458]_ ,
    \new_[16459]_ , \new_[16463]_ , \new_[16464]_ , \new_[16465]_ ,
    \new_[16469]_ , \new_[16470]_ , \new_[16474]_ , \new_[16475]_ ,
    \new_[16476]_ , \new_[16480]_ , \new_[16481]_ , \new_[16485]_ ,
    \new_[16486]_ , \new_[16487]_ , \new_[16491]_ , \new_[16492]_ ,
    \new_[16496]_ , \new_[16497]_ , \new_[16498]_ , \new_[16502]_ ,
    \new_[16503]_ , \new_[16507]_ , \new_[16508]_ , \new_[16509]_ ,
    \new_[16513]_ , \new_[16514]_ , \new_[16518]_ , \new_[16519]_ ,
    \new_[16520]_ , \new_[16524]_ , \new_[16525]_ , \new_[16529]_ ,
    \new_[16530]_ , \new_[16531]_ , \new_[16535]_ , \new_[16536]_ ,
    \new_[16540]_ , \new_[16541]_ , \new_[16542]_ , \new_[16546]_ ,
    \new_[16547]_ , \new_[16551]_ , \new_[16552]_ , \new_[16553]_ ,
    \new_[16557]_ , \new_[16558]_ , \new_[16562]_ , \new_[16563]_ ,
    \new_[16564]_ , \new_[16568]_ , \new_[16569]_ , \new_[16573]_ ,
    \new_[16574]_ , \new_[16575]_ , \new_[16579]_ , \new_[16580]_ ,
    \new_[16584]_ , \new_[16585]_ , \new_[16586]_ , \new_[16590]_ ,
    \new_[16591]_ , \new_[16595]_ , \new_[16596]_ , \new_[16597]_ ,
    \new_[16601]_ , \new_[16602]_ , \new_[16606]_ , \new_[16607]_ ,
    \new_[16608]_ , \new_[16612]_ , \new_[16613]_ , \new_[16617]_ ,
    \new_[16618]_ , \new_[16619]_ , \new_[16623]_ , \new_[16624]_ ,
    \new_[16628]_ , \new_[16629]_ , \new_[16630]_ , \new_[16634]_ ,
    \new_[16635]_ , \new_[16639]_ , \new_[16640]_ , \new_[16641]_ ,
    \new_[16645]_ , \new_[16646]_ , \new_[16650]_ , \new_[16651]_ ,
    \new_[16652]_ , \new_[16656]_ , \new_[16657]_ , \new_[16661]_ ,
    \new_[16662]_ , \new_[16663]_ , \new_[16667]_ , \new_[16668]_ ,
    \new_[16672]_ , \new_[16673]_ , \new_[16674]_ , \new_[16678]_ ,
    \new_[16679]_ , \new_[16683]_ , \new_[16684]_ , \new_[16685]_ ,
    \new_[16689]_ , \new_[16690]_ , \new_[16694]_ , \new_[16695]_ ,
    \new_[16696]_ , \new_[16700]_ , \new_[16701]_ , \new_[16705]_ ,
    \new_[16706]_ , \new_[16707]_ , \new_[16711]_ , \new_[16712]_ ,
    \new_[16716]_ , \new_[16717]_ , \new_[16718]_ , \new_[16722]_ ,
    \new_[16723]_ , \new_[16727]_ , \new_[16728]_ , \new_[16729]_ ,
    \new_[16733]_ , \new_[16734]_ , \new_[16738]_ , \new_[16739]_ ,
    \new_[16740]_ , \new_[16744]_ , \new_[16745]_ , \new_[16749]_ ,
    \new_[16750]_ , \new_[16751]_ , \new_[16755]_ , \new_[16756]_ ,
    \new_[16760]_ , \new_[16761]_ , \new_[16762]_ , \new_[16766]_ ,
    \new_[16767]_ , \new_[16771]_ , \new_[16772]_ , \new_[16773]_ ,
    \new_[16777]_ , \new_[16778]_ , \new_[16782]_ , \new_[16783]_ ,
    \new_[16784]_ , \new_[16788]_ , \new_[16789]_ , \new_[16793]_ ,
    \new_[16794]_ , \new_[16795]_ , \new_[16799]_ , \new_[16800]_ ,
    \new_[16804]_ , \new_[16805]_ , \new_[16806]_ , \new_[16810]_ ,
    \new_[16811]_ , \new_[16815]_ , \new_[16816]_ , \new_[16817]_ ,
    \new_[16821]_ , \new_[16822]_ , \new_[16826]_ , \new_[16827]_ ,
    \new_[16828]_ , \new_[16832]_ , \new_[16833]_ , \new_[16837]_ ,
    \new_[16838]_ , \new_[16839]_ , \new_[16843]_ , \new_[16844]_ ,
    \new_[16848]_ , \new_[16849]_ , \new_[16850]_ , \new_[16854]_ ,
    \new_[16855]_ , \new_[16859]_ , \new_[16860]_ , \new_[16861]_ ,
    \new_[16865]_ , \new_[16866]_ , \new_[16870]_ , \new_[16871]_ ,
    \new_[16872]_ , \new_[16876]_ , \new_[16877]_ , \new_[16881]_ ,
    \new_[16882]_ , \new_[16883]_ , \new_[16887]_ , \new_[16888]_ ,
    \new_[16892]_ , \new_[16893]_ , \new_[16894]_ , \new_[16898]_ ,
    \new_[16899]_ , \new_[16903]_ , \new_[16904]_ , \new_[16905]_ ,
    \new_[16909]_ , \new_[16910]_ , \new_[16914]_ , \new_[16915]_ ,
    \new_[16916]_ , \new_[16920]_ , \new_[16921]_ , \new_[16925]_ ,
    \new_[16926]_ , \new_[16927]_ , \new_[16931]_ , \new_[16932]_ ,
    \new_[16936]_ , \new_[16937]_ , \new_[16938]_ , \new_[16942]_ ,
    \new_[16943]_ , \new_[16947]_ , \new_[16948]_ , \new_[16949]_ ,
    \new_[16953]_ , \new_[16954]_ , \new_[16958]_ , \new_[16959]_ ,
    \new_[16960]_ , \new_[16964]_ , \new_[16965]_ , \new_[16969]_ ,
    \new_[16970]_ , \new_[16971]_ , \new_[16975]_ , \new_[16976]_ ,
    \new_[16980]_ , \new_[16981]_ , \new_[16982]_ , \new_[16986]_ ,
    \new_[16987]_ , \new_[16991]_ , \new_[16992]_ , \new_[16993]_ ,
    \new_[16997]_ , \new_[16998]_ , \new_[17002]_ , \new_[17003]_ ,
    \new_[17004]_ , \new_[17008]_ , \new_[17009]_ , \new_[17013]_ ,
    \new_[17014]_ , \new_[17015]_ , \new_[17019]_ , \new_[17020]_ ,
    \new_[17024]_ , \new_[17025]_ , \new_[17026]_ , \new_[17030]_ ,
    \new_[17031]_ , \new_[17035]_ , \new_[17036]_ , \new_[17037]_ ,
    \new_[17041]_ , \new_[17042]_ , \new_[17046]_ , \new_[17047]_ ,
    \new_[17048]_ , \new_[17052]_ , \new_[17053]_ , \new_[17057]_ ,
    \new_[17058]_ , \new_[17059]_ , \new_[17063]_ , \new_[17064]_ ,
    \new_[17068]_ , \new_[17069]_ , \new_[17070]_ , \new_[17074]_ ,
    \new_[17075]_ , \new_[17079]_ , \new_[17080]_ , \new_[17081]_ ,
    \new_[17085]_ , \new_[17086]_ , \new_[17090]_ , \new_[17091]_ ,
    \new_[17092]_ , \new_[17096]_ , \new_[17097]_ , \new_[17101]_ ,
    \new_[17102]_ , \new_[17103]_ , \new_[17107]_ , \new_[17108]_ ,
    \new_[17112]_ , \new_[17113]_ , \new_[17114]_ , \new_[17118]_ ,
    \new_[17119]_ , \new_[17123]_ , \new_[17124]_ , \new_[17125]_ ,
    \new_[17129]_ , \new_[17130]_ , \new_[17134]_ , \new_[17135]_ ,
    \new_[17136]_ , \new_[17140]_ , \new_[17141]_ , \new_[17145]_ ,
    \new_[17146]_ , \new_[17147]_ , \new_[17151]_ , \new_[17152]_ ,
    \new_[17156]_ , \new_[17157]_ , \new_[17158]_ , \new_[17162]_ ,
    \new_[17163]_ , \new_[17167]_ , \new_[17168]_ , \new_[17169]_ ,
    \new_[17173]_ , \new_[17174]_ , \new_[17178]_ , \new_[17179]_ ,
    \new_[17180]_ , \new_[17184]_ , \new_[17185]_ , \new_[17189]_ ,
    \new_[17190]_ , \new_[17191]_ , \new_[17195]_ , \new_[17196]_ ,
    \new_[17200]_ , \new_[17201]_ , \new_[17202]_ , \new_[17206]_ ,
    \new_[17207]_ , \new_[17211]_ , \new_[17212]_ , \new_[17213]_ ,
    \new_[17217]_ , \new_[17218]_ , \new_[17222]_ , \new_[17223]_ ,
    \new_[17224]_ , \new_[17228]_ , \new_[17229]_ , \new_[17233]_ ,
    \new_[17234]_ , \new_[17235]_ , \new_[17239]_ , \new_[17240]_ ,
    \new_[17244]_ , \new_[17245]_ , \new_[17246]_ , \new_[17250]_ ,
    \new_[17251]_ , \new_[17255]_ , \new_[17256]_ , \new_[17257]_ ,
    \new_[17261]_ , \new_[17262]_ , \new_[17266]_ , \new_[17267]_ ,
    \new_[17268]_ , \new_[17272]_ , \new_[17273]_ , \new_[17277]_ ,
    \new_[17278]_ , \new_[17279]_ , \new_[17283]_ , \new_[17284]_ ,
    \new_[17288]_ , \new_[17289]_ , \new_[17290]_ , \new_[17294]_ ,
    \new_[17295]_ , \new_[17299]_ , \new_[17300]_ , \new_[17301]_ ,
    \new_[17305]_ , \new_[17306]_ , \new_[17310]_ , \new_[17311]_ ,
    \new_[17312]_ , \new_[17316]_ , \new_[17317]_ , \new_[17321]_ ,
    \new_[17322]_ , \new_[17323]_ , \new_[17327]_ , \new_[17328]_ ,
    \new_[17332]_ , \new_[17333]_ , \new_[17334]_ , \new_[17338]_ ,
    \new_[17339]_ , \new_[17343]_ , \new_[17344]_ , \new_[17345]_ ,
    \new_[17349]_ , \new_[17350]_ , \new_[17354]_ , \new_[17355]_ ,
    \new_[17356]_ , \new_[17360]_ , \new_[17361]_ , \new_[17365]_ ,
    \new_[17366]_ , \new_[17367]_ , \new_[17371]_ , \new_[17372]_ ,
    \new_[17376]_ , \new_[17377]_ , \new_[17378]_ , \new_[17382]_ ,
    \new_[17383]_ , \new_[17387]_ , \new_[17388]_ , \new_[17389]_ ,
    \new_[17393]_ , \new_[17394]_ , \new_[17398]_ , \new_[17399]_ ,
    \new_[17400]_ , \new_[17404]_ , \new_[17405]_ , \new_[17409]_ ,
    \new_[17410]_ , \new_[17411]_ , \new_[17415]_ , \new_[17416]_ ,
    \new_[17420]_ , \new_[17421]_ , \new_[17422]_ , \new_[17426]_ ,
    \new_[17427]_ , \new_[17431]_ , \new_[17432]_ , \new_[17433]_ ,
    \new_[17437]_ , \new_[17438]_ , \new_[17442]_ , \new_[17443]_ ,
    \new_[17444]_ , \new_[17448]_ , \new_[17449]_ , \new_[17453]_ ,
    \new_[17454]_ , \new_[17455]_ , \new_[17459]_ , \new_[17460]_ ,
    \new_[17464]_ , \new_[17465]_ , \new_[17466]_ , \new_[17470]_ ,
    \new_[17471]_ , \new_[17475]_ , \new_[17476]_ , \new_[17477]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17486]_ , \new_[17487]_ ,
    \new_[17488]_ , \new_[17492]_ , \new_[17493]_ , \new_[17497]_ ,
    \new_[17498]_ , \new_[17499]_ , \new_[17503]_ , \new_[17504]_ ,
    \new_[17508]_ , \new_[17509]_ , \new_[17510]_ , \new_[17514]_ ,
    \new_[17515]_ , \new_[17519]_ , \new_[17520]_ , \new_[17521]_ ,
    \new_[17525]_ , \new_[17526]_ , \new_[17530]_ , \new_[17531]_ ,
    \new_[17532]_ , \new_[17536]_ , \new_[17537]_ , \new_[17541]_ ,
    \new_[17542]_ , \new_[17543]_ , \new_[17547]_ , \new_[17548]_ ,
    \new_[17552]_ , \new_[17553]_ , \new_[17554]_ , \new_[17558]_ ,
    \new_[17559]_ , \new_[17563]_ , \new_[17564]_ , \new_[17565]_ ,
    \new_[17569]_ , \new_[17570]_ , \new_[17574]_ , \new_[17575]_ ,
    \new_[17576]_ , \new_[17580]_ , \new_[17581]_ , \new_[17585]_ ,
    \new_[17586]_ , \new_[17587]_ , \new_[17591]_ , \new_[17592]_ ,
    \new_[17596]_ , \new_[17597]_ , \new_[17598]_ , \new_[17602]_ ,
    \new_[17603]_ , \new_[17607]_ , \new_[17608]_ , \new_[17609]_ ,
    \new_[17613]_ , \new_[17614]_ , \new_[17618]_ , \new_[17619]_ ,
    \new_[17620]_ , \new_[17624]_ , \new_[17625]_ , \new_[17629]_ ,
    \new_[17630]_ , \new_[17631]_ , \new_[17635]_ , \new_[17636]_ ,
    \new_[17640]_ , \new_[17641]_ , \new_[17642]_ , \new_[17646]_ ,
    \new_[17647]_ , \new_[17651]_ , \new_[17652]_ , \new_[17653]_ ,
    \new_[17657]_ , \new_[17658]_ , \new_[17662]_ , \new_[17663]_ ,
    \new_[17664]_ , \new_[17668]_ , \new_[17669]_ , \new_[17673]_ ,
    \new_[17674]_ , \new_[17675]_ , \new_[17679]_ , \new_[17680]_ ,
    \new_[17684]_ , \new_[17685]_ , \new_[17686]_ , \new_[17690]_ ,
    \new_[17691]_ , \new_[17695]_ , \new_[17696]_ , \new_[17697]_ ,
    \new_[17701]_ , \new_[17702]_ , \new_[17706]_ , \new_[17707]_ ,
    \new_[17708]_ , \new_[17712]_ , \new_[17713]_ , \new_[17717]_ ,
    \new_[17718]_ , \new_[17719]_ , \new_[17723]_ , \new_[17724]_ ,
    \new_[17728]_ , \new_[17729]_ , \new_[17730]_ , \new_[17734]_ ,
    \new_[17735]_ , \new_[17739]_ , \new_[17740]_ , \new_[17741]_ ,
    \new_[17745]_ , \new_[17746]_ , \new_[17750]_ , \new_[17751]_ ,
    \new_[17752]_ , \new_[17756]_ , \new_[17757]_ , \new_[17761]_ ,
    \new_[17762]_ , \new_[17763]_ , \new_[17767]_ , \new_[17768]_ ,
    \new_[17772]_ , \new_[17773]_ , \new_[17774]_ , \new_[17778]_ ,
    \new_[17779]_ , \new_[17783]_ , \new_[17784]_ , \new_[17785]_ ,
    \new_[17789]_ , \new_[17790]_ , \new_[17794]_ , \new_[17795]_ ,
    \new_[17796]_ , \new_[17800]_ , \new_[17801]_ , \new_[17805]_ ,
    \new_[17806]_ , \new_[17807]_ , \new_[17811]_ , \new_[17812]_ ,
    \new_[17816]_ , \new_[17817]_ , \new_[17818]_ , \new_[17822]_ ,
    \new_[17823]_ , \new_[17827]_ , \new_[17828]_ , \new_[17829]_ ,
    \new_[17833]_ , \new_[17834]_ , \new_[17838]_ , \new_[17839]_ ,
    \new_[17840]_ , \new_[17844]_ , \new_[17845]_ , \new_[17849]_ ,
    \new_[17850]_ , \new_[17851]_ , \new_[17855]_ , \new_[17856]_ ,
    \new_[17860]_ , \new_[17861]_ , \new_[17862]_ , \new_[17866]_ ,
    \new_[17867]_ , \new_[17871]_ , \new_[17872]_ , \new_[17873]_ ,
    \new_[17877]_ , \new_[17878]_ , \new_[17882]_ , \new_[17883]_ ,
    \new_[17884]_ , \new_[17888]_ , \new_[17889]_ , \new_[17893]_ ,
    \new_[17894]_ , \new_[17895]_ , \new_[17899]_ , \new_[17900]_ ,
    \new_[17904]_ , \new_[17905]_ , \new_[17906]_ , \new_[17910]_ ,
    \new_[17911]_ , \new_[17915]_ , \new_[17916]_ , \new_[17917]_ ,
    \new_[17921]_ , \new_[17922]_ , \new_[17926]_ , \new_[17927]_ ,
    \new_[17928]_ , \new_[17932]_ , \new_[17933]_ , \new_[17937]_ ,
    \new_[17938]_ , \new_[17939]_ , \new_[17943]_ , \new_[17944]_ ,
    \new_[17948]_ , \new_[17949]_ , \new_[17950]_ , \new_[17954]_ ,
    \new_[17955]_ , \new_[17959]_ , \new_[17960]_ , \new_[17961]_ ,
    \new_[17965]_ , \new_[17966]_ , \new_[17970]_ , \new_[17971]_ ,
    \new_[17972]_ , \new_[17976]_ , \new_[17977]_ , \new_[17981]_ ,
    \new_[17982]_ , \new_[17983]_ , \new_[17987]_ , \new_[17988]_ ,
    \new_[17992]_ , \new_[17993]_ , \new_[17994]_ , \new_[17998]_ ,
    \new_[17999]_ , \new_[18003]_ , \new_[18004]_ , \new_[18005]_ ,
    \new_[18009]_ , \new_[18010]_ , \new_[18014]_ , \new_[18015]_ ,
    \new_[18016]_ , \new_[18020]_ , \new_[18021]_ , \new_[18025]_ ,
    \new_[18026]_ , \new_[18027]_ , \new_[18031]_ , \new_[18032]_ ,
    \new_[18036]_ , \new_[18037]_ , \new_[18038]_ , \new_[18042]_ ,
    \new_[18043]_ , \new_[18047]_ , \new_[18048]_ , \new_[18049]_ ,
    \new_[18053]_ , \new_[18054]_ , \new_[18058]_ , \new_[18059]_ ,
    \new_[18060]_ , \new_[18064]_ , \new_[18065]_ , \new_[18069]_ ,
    \new_[18070]_ , \new_[18071]_ , \new_[18075]_ , \new_[18076]_ ,
    \new_[18080]_ , \new_[18081]_ , \new_[18082]_ , \new_[18086]_ ,
    \new_[18087]_ , \new_[18091]_ , \new_[18092]_ , \new_[18093]_ ,
    \new_[18097]_ , \new_[18098]_ , \new_[18102]_ , \new_[18103]_ ,
    \new_[18104]_ , \new_[18108]_ , \new_[18109]_ , \new_[18113]_ ,
    \new_[18114]_ , \new_[18115]_ , \new_[18119]_ , \new_[18120]_ ,
    \new_[18124]_ , \new_[18125]_ , \new_[18126]_ , \new_[18130]_ ,
    \new_[18131]_ , \new_[18135]_ , \new_[18136]_ , \new_[18137]_ ,
    \new_[18141]_ , \new_[18142]_ , \new_[18146]_ , \new_[18147]_ ,
    \new_[18148]_ , \new_[18152]_ , \new_[18153]_ , \new_[18157]_ ,
    \new_[18158]_ , \new_[18159]_ , \new_[18163]_ , \new_[18164]_ ,
    \new_[18168]_ , \new_[18169]_ , \new_[18170]_ , \new_[18174]_ ,
    \new_[18175]_ , \new_[18179]_ , \new_[18180]_ , \new_[18181]_ ,
    \new_[18185]_ , \new_[18186]_ , \new_[18190]_ , \new_[18191]_ ,
    \new_[18192]_ , \new_[18196]_ , \new_[18197]_ , \new_[18201]_ ,
    \new_[18202]_ , \new_[18203]_ , \new_[18207]_ , \new_[18208]_ ,
    \new_[18212]_ , \new_[18213]_ , \new_[18214]_ , \new_[18218]_ ,
    \new_[18219]_ , \new_[18223]_ , \new_[18224]_ , \new_[18225]_ ,
    \new_[18229]_ , \new_[18230]_ , \new_[18234]_ , \new_[18235]_ ,
    \new_[18236]_ , \new_[18240]_ , \new_[18241]_ , \new_[18245]_ ,
    \new_[18246]_ , \new_[18247]_ , \new_[18251]_ , \new_[18252]_ ,
    \new_[18256]_ , \new_[18257]_ , \new_[18258]_ , \new_[18262]_ ,
    \new_[18263]_ , \new_[18267]_ , \new_[18268]_ , \new_[18269]_ ,
    \new_[18273]_ , \new_[18274]_ , \new_[18278]_ , \new_[18279]_ ,
    \new_[18280]_ , \new_[18284]_ , \new_[18285]_ , \new_[18289]_ ,
    \new_[18290]_ , \new_[18291]_ , \new_[18295]_ , \new_[18296]_ ,
    \new_[18300]_ , \new_[18301]_ , \new_[18302]_ , \new_[18306]_ ,
    \new_[18307]_ , \new_[18311]_ , \new_[18312]_ , \new_[18313]_ ,
    \new_[18317]_ , \new_[18318]_ , \new_[18322]_ , \new_[18323]_ ,
    \new_[18324]_ , \new_[18328]_ , \new_[18329]_ , \new_[18333]_ ,
    \new_[18334]_ , \new_[18335]_ , \new_[18339]_ , \new_[18340]_ ,
    \new_[18344]_ , \new_[18345]_ , \new_[18346]_ , \new_[18350]_ ,
    \new_[18351]_ , \new_[18355]_ , \new_[18356]_ , \new_[18357]_ ,
    \new_[18361]_ , \new_[18362]_ , \new_[18366]_ , \new_[18367]_ ,
    \new_[18368]_ , \new_[18372]_ , \new_[18373]_ , \new_[18377]_ ,
    \new_[18378]_ , \new_[18379]_ , \new_[18383]_ , \new_[18384]_ ,
    \new_[18388]_ , \new_[18389]_ , \new_[18390]_ , \new_[18394]_ ,
    \new_[18395]_ , \new_[18399]_ , \new_[18400]_ , \new_[18401]_ ,
    \new_[18405]_ , \new_[18406]_ , \new_[18410]_ , \new_[18411]_ ,
    \new_[18412]_ , \new_[18416]_ , \new_[18417]_ , \new_[18421]_ ,
    \new_[18422]_ , \new_[18423]_ , \new_[18427]_ , \new_[18428]_ ,
    \new_[18432]_ , \new_[18433]_ , \new_[18434]_ , \new_[18438]_ ,
    \new_[18439]_ , \new_[18443]_ , \new_[18444]_ , \new_[18445]_ ,
    \new_[18449]_ , \new_[18450]_ , \new_[18454]_ , \new_[18455]_ ,
    \new_[18456]_ , \new_[18460]_ , \new_[18461]_ , \new_[18465]_ ,
    \new_[18466]_ , \new_[18467]_ , \new_[18471]_ , \new_[18472]_ ,
    \new_[18476]_ , \new_[18477]_ , \new_[18478]_ , \new_[18482]_ ,
    \new_[18483]_ , \new_[18487]_ , \new_[18488]_ , \new_[18489]_ ,
    \new_[18493]_ , \new_[18494]_ , \new_[18498]_ , \new_[18499]_ ,
    \new_[18500]_ , \new_[18504]_ , \new_[18505]_ , \new_[18509]_ ,
    \new_[18510]_ , \new_[18511]_ , \new_[18515]_ , \new_[18516]_ ,
    \new_[18520]_ , \new_[18521]_ , \new_[18522]_ , \new_[18526]_ ,
    \new_[18527]_ , \new_[18531]_ , \new_[18532]_ , \new_[18533]_ ,
    \new_[18537]_ , \new_[18538]_ , \new_[18542]_ , \new_[18543]_ ,
    \new_[18544]_ , \new_[18548]_ , \new_[18549]_ , \new_[18553]_ ,
    \new_[18554]_ , \new_[18555]_ , \new_[18559]_ , \new_[18560]_ ,
    \new_[18564]_ , \new_[18565]_ , \new_[18566]_ , \new_[18570]_ ,
    \new_[18571]_ , \new_[18575]_ , \new_[18576]_ , \new_[18577]_ ,
    \new_[18581]_ , \new_[18582]_ , \new_[18586]_ , \new_[18587]_ ,
    \new_[18588]_ , \new_[18592]_ , \new_[18593]_ , \new_[18597]_ ,
    \new_[18598]_ , \new_[18599]_ , \new_[18603]_ , \new_[18604]_ ,
    \new_[18608]_ , \new_[18609]_ , \new_[18610]_ , \new_[18614]_ ,
    \new_[18615]_ , \new_[18619]_ , \new_[18620]_ , \new_[18621]_ ,
    \new_[18625]_ , \new_[18626]_ , \new_[18630]_ , \new_[18631]_ ,
    \new_[18632]_ , \new_[18636]_ , \new_[18637]_ , \new_[18641]_ ,
    \new_[18642]_ , \new_[18643]_ , \new_[18647]_ , \new_[18648]_ ,
    \new_[18652]_ , \new_[18653]_ , \new_[18654]_ , \new_[18658]_ ,
    \new_[18659]_ , \new_[18663]_ , \new_[18664]_ , \new_[18665]_ ,
    \new_[18669]_ , \new_[18670]_ , \new_[18674]_ , \new_[18675]_ ,
    \new_[18676]_ , \new_[18680]_ , \new_[18681]_ , \new_[18685]_ ,
    \new_[18686]_ , \new_[18687]_ , \new_[18691]_ , \new_[18692]_ ,
    \new_[18696]_ , \new_[18697]_ , \new_[18698]_ , \new_[18702]_ ,
    \new_[18703]_ , \new_[18707]_ , \new_[18708]_ , \new_[18709]_ ,
    \new_[18713]_ , \new_[18714]_ , \new_[18718]_ , \new_[18719]_ ,
    \new_[18720]_ , \new_[18724]_ , \new_[18725]_ , \new_[18729]_ ,
    \new_[18730]_ , \new_[18731]_ , \new_[18735]_ , \new_[18736]_ ,
    \new_[18740]_ , \new_[18741]_ , \new_[18742]_ , \new_[18746]_ ,
    \new_[18747]_ , \new_[18751]_ , \new_[18752]_ , \new_[18753]_ ,
    \new_[18757]_ , \new_[18758]_ , \new_[18762]_ , \new_[18763]_ ,
    \new_[18764]_ , \new_[18768]_ , \new_[18769]_ , \new_[18773]_ ,
    \new_[18774]_ , \new_[18775]_ , \new_[18779]_ , \new_[18780]_ ,
    \new_[18784]_ , \new_[18785]_ , \new_[18786]_ , \new_[18790]_ ,
    \new_[18791]_ , \new_[18795]_ , \new_[18796]_ , \new_[18797]_ ,
    \new_[18801]_ , \new_[18802]_ , \new_[18806]_ , \new_[18807]_ ,
    \new_[18808]_ , \new_[18812]_ , \new_[18813]_ , \new_[18817]_ ,
    \new_[18818]_ , \new_[18819]_ , \new_[18823]_ , \new_[18824]_ ,
    \new_[18828]_ , \new_[18829]_ , \new_[18830]_ , \new_[18834]_ ,
    \new_[18835]_ , \new_[18839]_ , \new_[18840]_ , \new_[18841]_ ,
    \new_[18845]_ , \new_[18846]_ , \new_[18850]_ , \new_[18851]_ ,
    \new_[18852]_ , \new_[18856]_ , \new_[18857]_ , \new_[18861]_ ,
    \new_[18862]_ , \new_[18863]_ , \new_[18867]_ , \new_[18868]_ ,
    \new_[18872]_ , \new_[18873]_ , \new_[18874]_ , \new_[18878]_ ,
    \new_[18879]_ , \new_[18883]_ , \new_[18884]_ , \new_[18885]_ ,
    \new_[18889]_ , \new_[18890]_ , \new_[18894]_ , \new_[18895]_ ,
    \new_[18896]_ , \new_[18900]_ , \new_[18901]_ , \new_[18905]_ ,
    \new_[18906]_ , \new_[18907]_ , \new_[18911]_ , \new_[18912]_ ,
    \new_[18916]_ , \new_[18917]_ , \new_[18918]_ , \new_[18922]_ ,
    \new_[18923]_ , \new_[18927]_ , \new_[18928]_ , \new_[18929]_ ,
    \new_[18933]_ , \new_[18934]_ , \new_[18938]_ , \new_[18939]_ ,
    \new_[18940]_ , \new_[18944]_ , \new_[18945]_ , \new_[18949]_ ,
    \new_[18950]_ , \new_[18951]_ , \new_[18955]_ , \new_[18956]_ ,
    \new_[18960]_ , \new_[18961]_ , \new_[18962]_ , \new_[18966]_ ,
    \new_[18967]_ , \new_[18971]_ , \new_[18972]_ , \new_[18973]_ ,
    \new_[18977]_ , \new_[18978]_ , \new_[18982]_ , \new_[18983]_ ,
    \new_[18984]_ , \new_[18988]_ , \new_[18989]_ , \new_[18993]_ ,
    \new_[18994]_ , \new_[18995]_ , \new_[18999]_ , \new_[19000]_ ,
    \new_[19004]_ , \new_[19005]_ , \new_[19006]_ , \new_[19010]_ ,
    \new_[19011]_ , \new_[19015]_ , \new_[19016]_ , \new_[19017]_ ,
    \new_[19021]_ , \new_[19022]_ , \new_[19026]_ , \new_[19027]_ ,
    \new_[19028]_ , \new_[19032]_ , \new_[19033]_ , \new_[19037]_ ,
    \new_[19038]_ , \new_[19039]_ , \new_[19043]_ , \new_[19044]_ ,
    \new_[19048]_ , \new_[19049]_ , \new_[19050]_ , \new_[19054]_ ,
    \new_[19055]_ , \new_[19059]_ , \new_[19060]_ , \new_[19061]_ ,
    \new_[19065]_ , \new_[19066]_ , \new_[19070]_ , \new_[19071]_ ,
    \new_[19072]_ , \new_[19076]_ , \new_[19077]_ , \new_[19081]_ ,
    \new_[19082]_ , \new_[19083]_ , \new_[19087]_ , \new_[19088]_ ,
    \new_[19092]_ , \new_[19093]_ , \new_[19094]_ , \new_[19098]_ ,
    \new_[19099]_ , \new_[19103]_ , \new_[19104]_ , \new_[19105]_ ,
    \new_[19109]_ , \new_[19110]_ , \new_[19114]_ , \new_[19115]_ ,
    \new_[19116]_ , \new_[19120]_ , \new_[19121]_ , \new_[19125]_ ,
    \new_[19126]_ , \new_[19127]_ , \new_[19131]_ , \new_[19132]_ ,
    \new_[19136]_ , \new_[19137]_ , \new_[19138]_ , \new_[19142]_ ,
    \new_[19143]_ , \new_[19147]_ , \new_[19148]_ , \new_[19149]_ ,
    \new_[19153]_ , \new_[19154]_ , \new_[19158]_ , \new_[19159]_ ,
    \new_[19160]_ , \new_[19164]_ , \new_[19165]_ , \new_[19169]_ ,
    \new_[19170]_ , \new_[19171]_ , \new_[19175]_ , \new_[19176]_ ,
    \new_[19180]_ , \new_[19181]_ , \new_[19182]_ , \new_[19186]_ ,
    \new_[19187]_ , \new_[19191]_ , \new_[19192]_ , \new_[19193]_ ,
    \new_[19197]_ , \new_[19198]_ , \new_[19202]_ , \new_[19203]_ ,
    \new_[19204]_ , \new_[19208]_ , \new_[19209]_ , \new_[19213]_ ,
    \new_[19214]_ , \new_[19215]_ , \new_[19219]_ , \new_[19220]_ ,
    \new_[19224]_ , \new_[19225]_ , \new_[19226]_ , \new_[19230]_ ,
    \new_[19231]_ , \new_[19235]_ , \new_[19236]_ , \new_[19237]_ ,
    \new_[19241]_ , \new_[19242]_ , \new_[19246]_ , \new_[19247]_ ,
    \new_[19248]_ , \new_[19252]_ , \new_[19253]_ , \new_[19257]_ ,
    \new_[19258]_ , \new_[19259]_ , \new_[19263]_ , \new_[19264]_ ,
    \new_[19268]_ , \new_[19269]_ , \new_[19270]_ , \new_[19274]_ ,
    \new_[19275]_ , \new_[19279]_ , \new_[19280]_ , \new_[19281]_ ,
    \new_[19285]_ , \new_[19286]_ , \new_[19290]_ , \new_[19291]_ ,
    \new_[19292]_ , \new_[19296]_ , \new_[19297]_ , \new_[19301]_ ,
    \new_[19302]_ , \new_[19303]_ , \new_[19307]_ , \new_[19308]_ ,
    \new_[19311]_ , \new_[19314]_ , \new_[19315]_ , \new_[19316]_ ,
    \new_[19320]_ , \new_[19321]_ , \new_[19325]_ , \new_[19326]_ ,
    \new_[19327]_ , \new_[19331]_ , \new_[19332]_ , \new_[19335]_ ,
    \new_[19338]_ , \new_[19339]_ , \new_[19340]_ , \new_[19344]_ ,
    \new_[19345]_ , \new_[19349]_ , \new_[19350]_ , \new_[19351]_ ,
    \new_[19355]_ , \new_[19356]_ , \new_[19359]_ , \new_[19362]_ ,
    \new_[19363]_ , \new_[19364]_ , \new_[19368]_ , \new_[19369]_ ,
    \new_[19373]_ , \new_[19374]_ , \new_[19375]_ , \new_[19379]_ ,
    \new_[19380]_ , \new_[19383]_ , \new_[19386]_ , \new_[19387]_ ,
    \new_[19388]_ , \new_[19392]_ , \new_[19393]_ , \new_[19397]_ ,
    \new_[19398]_ , \new_[19399]_ , \new_[19403]_ , \new_[19404]_ ,
    \new_[19407]_ , \new_[19410]_ , \new_[19411]_ , \new_[19412]_ ,
    \new_[19416]_ , \new_[19417]_ , \new_[19421]_ , \new_[19422]_ ,
    \new_[19423]_ , \new_[19427]_ , \new_[19428]_ , \new_[19431]_ ,
    \new_[19434]_ , \new_[19435]_ , \new_[19436]_ , \new_[19440]_ ,
    \new_[19441]_ , \new_[19445]_ , \new_[19446]_ , \new_[19447]_ ,
    \new_[19451]_ , \new_[19452]_ , \new_[19455]_ , \new_[19458]_ ,
    \new_[19459]_ , \new_[19460]_ , \new_[19464]_ , \new_[19465]_ ,
    \new_[19469]_ , \new_[19470]_ , \new_[19471]_ , \new_[19475]_ ,
    \new_[19476]_ , \new_[19479]_ , \new_[19482]_ , \new_[19483]_ ,
    \new_[19484]_ , \new_[19488]_ , \new_[19489]_ , \new_[19493]_ ,
    \new_[19494]_ , \new_[19495]_ , \new_[19499]_ , \new_[19500]_ ,
    \new_[19503]_ , \new_[19506]_ , \new_[19507]_ , \new_[19508]_ ,
    \new_[19512]_ , \new_[19513]_ , \new_[19517]_ , \new_[19518]_ ,
    \new_[19519]_ , \new_[19523]_ , \new_[19524]_ , \new_[19527]_ ,
    \new_[19530]_ , \new_[19531]_ , \new_[19532]_ , \new_[19536]_ ,
    \new_[19537]_ , \new_[19541]_ , \new_[19542]_ , \new_[19543]_ ,
    \new_[19547]_ , \new_[19548]_ , \new_[19551]_ , \new_[19554]_ ,
    \new_[19555]_ , \new_[19556]_ , \new_[19560]_ , \new_[19561]_ ,
    \new_[19565]_ , \new_[19566]_ , \new_[19567]_ , \new_[19571]_ ,
    \new_[19572]_ , \new_[19575]_ , \new_[19578]_ , \new_[19579]_ ,
    \new_[19580]_ , \new_[19584]_ , \new_[19585]_ , \new_[19589]_ ,
    \new_[19590]_ , \new_[19591]_ , \new_[19595]_ , \new_[19596]_ ,
    \new_[19599]_ , \new_[19602]_ , \new_[19603]_ , \new_[19604]_ ,
    \new_[19608]_ , \new_[19609]_ , \new_[19613]_ , \new_[19614]_ ,
    \new_[19615]_ , \new_[19619]_ , \new_[19620]_ , \new_[19623]_ ,
    \new_[19626]_ , \new_[19627]_ , \new_[19628]_ , \new_[19632]_ ,
    \new_[19633]_ , \new_[19637]_ , \new_[19638]_ , \new_[19639]_ ,
    \new_[19643]_ , \new_[19644]_ , \new_[19647]_ , \new_[19650]_ ,
    \new_[19651]_ , \new_[19652]_ , \new_[19656]_ , \new_[19657]_ ,
    \new_[19661]_ , \new_[19662]_ , \new_[19663]_ , \new_[19667]_ ,
    \new_[19668]_ , \new_[19671]_ , \new_[19674]_ , \new_[19675]_ ,
    \new_[19676]_ , \new_[19680]_ , \new_[19681]_ , \new_[19685]_ ,
    \new_[19686]_ , \new_[19687]_ , \new_[19691]_ , \new_[19692]_ ,
    \new_[19695]_ , \new_[19698]_ , \new_[19699]_ , \new_[19700]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19709]_ , \new_[19710]_ ,
    \new_[19711]_ , \new_[19715]_ , \new_[19716]_ , \new_[19719]_ ,
    \new_[19722]_ , \new_[19723]_ , \new_[19724]_ , \new_[19728]_ ,
    \new_[19729]_ , \new_[19733]_ , \new_[19734]_ , \new_[19735]_ ,
    \new_[19739]_ , \new_[19740]_ , \new_[19743]_ , \new_[19746]_ ,
    \new_[19747]_ , \new_[19748]_ , \new_[19752]_ , \new_[19753]_ ,
    \new_[19757]_ , \new_[19758]_ , \new_[19759]_ , \new_[19763]_ ,
    \new_[19764]_ , \new_[19767]_ , \new_[19770]_ , \new_[19771]_ ,
    \new_[19772]_ , \new_[19776]_ , \new_[19777]_ , \new_[19781]_ ,
    \new_[19782]_ , \new_[19783]_ , \new_[19787]_ , \new_[19788]_ ,
    \new_[19791]_ , \new_[19794]_ , \new_[19795]_ , \new_[19796]_ ,
    \new_[19800]_ , \new_[19801]_ , \new_[19805]_ , \new_[19806]_ ,
    \new_[19807]_ , \new_[19811]_ , \new_[19812]_ , \new_[19815]_ ,
    \new_[19818]_ , \new_[19819]_ , \new_[19820]_ , \new_[19824]_ ,
    \new_[19825]_ , \new_[19829]_ , \new_[19830]_ , \new_[19831]_ ,
    \new_[19835]_ , \new_[19836]_ , \new_[19839]_ , \new_[19842]_ ,
    \new_[19843]_ , \new_[19844]_ , \new_[19848]_ , \new_[19849]_ ,
    \new_[19853]_ , \new_[19854]_ , \new_[19855]_ , \new_[19859]_ ,
    \new_[19860]_ , \new_[19863]_ , \new_[19866]_ , \new_[19867]_ ,
    \new_[19868]_ , \new_[19872]_ , \new_[19873]_ , \new_[19877]_ ,
    \new_[19878]_ , \new_[19879]_ , \new_[19883]_ , \new_[19884]_ ,
    \new_[19887]_ , \new_[19890]_ , \new_[19891]_ , \new_[19892]_ ,
    \new_[19896]_ , \new_[19897]_ , \new_[19901]_ , \new_[19902]_ ,
    \new_[19903]_ , \new_[19907]_ , \new_[19908]_ , \new_[19911]_ ,
    \new_[19914]_ , \new_[19915]_ , \new_[19916]_ , \new_[19920]_ ,
    \new_[19921]_ , \new_[19925]_ , \new_[19926]_ , \new_[19927]_ ,
    \new_[19931]_ , \new_[19932]_ , \new_[19935]_ , \new_[19938]_ ,
    \new_[19939]_ , \new_[19940]_ , \new_[19944]_ , \new_[19945]_ ,
    \new_[19949]_ , \new_[19950]_ , \new_[19951]_ , \new_[19955]_ ,
    \new_[19956]_ , \new_[19959]_ , \new_[19962]_ , \new_[19963]_ ,
    \new_[19964]_ , \new_[19968]_ , \new_[19969]_ , \new_[19973]_ ,
    \new_[19974]_ , \new_[19975]_ , \new_[19979]_ , \new_[19980]_ ,
    \new_[19983]_ , \new_[19986]_ , \new_[19987]_ , \new_[19988]_ ,
    \new_[19992]_ , \new_[19993]_ , \new_[19997]_ , \new_[19998]_ ,
    \new_[19999]_ , \new_[20003]_ , \new_[20004]_ , \new_[20007]_ ,
    \new_[20010]_ , \new_[20011]_ , \new_[20012]_ , \new_[20016]_ ,
    \new_[20017]_ , \new_[20021]_ , \new_[20022]_ , \new_[20023]_ ,
    \new_[20027]_ , \new_[20028]_ , \new_[20031]_ , \new_[20034]_ ,
    \new_[20035]_ , \new_[20036]_ , \new_[20040]_ , \new_[20041]_ ,
    \new_[20045]_ , \new_[20046]_ , \new_[20047]_ , \new_[20051]_ ,
    \new_[20052]_ , \new_[20055]_ , \new_[20058]_ , \new_[20059]_ ,
    \new_[20060]_ , \new_[20064]_ , \new_[20065]_ , \new_[20069]_ ,
    \new_[20070]_ , \new_[20071]_ , \new_[20075]_ , \new_[20076]_ ,
    \new_[20079]_ , \new_[20082]_ , \new_[20083]_ , \new_[20084]_ ,
    \new_[20088]_ , \new_[20089]_ , \new_[20093]_ , \new_[20094]_ ,
    \new_[20095]_ , \new_[20099]_ , \new_[20100]_ , \new_[20103]_ ,
    \new_[20106]_ , \new_[20107]_ , \new_[20108]_ , \new_[20112]_ ,
    \new_[20113]_ , \new_[20117]_ , \new_[20118]_ , \new_[20119]_ ,
    \new_[20123]_ , \new_[20124]_ , \new_[20127]_ , \new_[20130]_ ,
    \new_[20131]_ , \new_[20132]_ , \new_[20136]_ , \new_[20137]_ ,
    \new_[20141]_ , \new_[20142]_ , \new_[20143]_ , \new_[20147]_ ,
    \new_[20148]_ , \new_[20151]_ , \new_[20154]_ , \new_[20155]_ ,
    \new_[20156]_ , \new_[20160]_ , \new_[20161]_ , \new_[20165]_ ,
    \new_[20166]_ , \new_[20167]_ , \new_[20171]_ , \new_[20172]_ ,
    \new_[20175]_ , \new_[20178]_ , \new_[20179]_ , \new_[20180]_ ,
    \new_[20184]_ , \new_[20185]_ , \new_[20189]_ , \new_[20190]_ ,
    \new_[20191]_ , \new_[20195]_ , \new_[20196]_ , \new_[20199]_ ,
    \new_[20202]_ , \new_[20203]_ , \new_[20204]_ , \new_[20208]_ ,
    \new_[20209]_ , \new_[20213]_ , \new_[20214]_ , \new_[20215]_ ,
    \new_[20219]_ , \new_[20220]_ , \new_[20223]_ , \new_[20226]_ ,
    \new_[20227]_ , \new_[20228]_ , \new_[20232]_ , \new_[20233]_ ,
    \new_[20237]_ , \new_[20238]_ , \new_[20239]_ , \new_[20243]_ ,
    \new_[20244]_ , \new_[20247]_ , \new_[20250]_ , \new_[20251]_ ,
    \new_[20252]_ , \new_[20256]_ , \new_[20257]_ , \new_[20261]_ ,
    \new_[20262]_ , \new_[20263]_ , \new_[20267]_ , \new_[20268]_ ,
    \new_[20271]_ , \new_[20274]_ , \new_[20275]_ , \new_[20276]_ ,
    \new_[20280]_ , \new_[20281]_ , \new_[20285]_ , \new_[20286]_ ,
    \new_[20287]_ , \new_[20291]_ , \new_[20292]_ , \new_[20295]_ ,
    \new_[20298]_ , \new_[20299]_ , \new_[20300]_ , \new_[20304]_ ,
    \new_[20305]_ , \new_[20309]_ , \new_[20310]_ , \new_[20311]_ ,
    \new_[20315]_ , \new_[20316]_ , \new_[20319]_ , \new_[20322]_ ,
    \new_[20323]_ , \new_[20324]_ , \new_[20328]_ , \new_[20329]_ ,
    \new_[20333]_ , \new_[20334]_ , \new_[20335]_ , \new_[20339]_ ,
    \new_[20340]_ , \new_[20343]_ , \new_[20346]_ , \new_[20347]_ ,
    \new_[20348]_ , \new_[20352]_ , \new_[20353]_ , \new_[20357]_ ,
    \new_[20358]_ , \new_[20359]_ , \new_[20363]_ , \new_[20364]_ ,
    \new_[20367]_ , \new_[20370]_ , \new_[20371]_ , \new_[20372]_ ,
    \new_[20376]_ , \new_[20377]_ , \new_[20381]_ , \new_[20382]_ ,
    \new_[20383]_ , \new_[20387]_ , \new_[20388]_ , \new_[20391]_ ,
    \new_[20394]_ , \new_[20395]_ , \new_[20396]_ , \new_[20400]_ ,
    \new_[20401]_ , \new_[20405]_ , \new_[20406]_ , \new_[20407]_ ,
    \new_[20411]_ , \new_[20412]_ , \new_[20415]_ , \new_[20418]_ ,
    \new_[20419]_ , \new_[20420]_ , \new_[20424]_ , \new_[20425]_ ,
    \new_[20429]_ , \new_[20430]_ , \new_[20431]_ , \new_[20435]_ ,
    \new_[20436]_ , \new_[20439]_ , \new_[20442]_ , \new_[20443]_ ,
    \new_[20444]_ , \new_[20448]_ , \new_[20449]_ , \new_[20453]_ ,
    \new_[20454]_ , \new_[20455]_ , \new_[20459]_ , \new_[20460]_ ,
    \new_[20463]_ , \new_[20466]_ , \new_[20467]_ , \new_[20468]_ ,
    \new_[20472]_ , \new_[20473]_ , \new_[20477]_ , \new_[20478]_ ,
    \new_[20479]_ , \new_[20483]_ , \new_[20484]_ , \new_[20487]_ ,
    \new_[20490]_ , \new_[20491]_ , \new_[20492]_ , \new_[20496]_ ,
    \new_[20497]_ , \new_[20501]_ , \new_[20502]_ , \new_[20503]_ ,
    \new_[20507]_ , \new_[20508]_ , \new_[20511]_ , \new_[20514]_ ,
    \new_[20515]_ , \new_[20516]_ , \new_[20520]_ , \new_[20521]_ ,
    \new_[20525]_ , \new_[20526]_ , \new_[20527]_ , \new_[20531]_ ,
    \new_[20532]_ , \new_[20535]_ , \new_[20538]_ , \new_[20539]_ ,
    \new_[20540]_ , \new_[20544]_ , \new_[20545]_ , \new_[20549]_ ,
    \new_[20550]_ , \new_[20551]_ , \new_[20555]_ , \new_[20556]_ ,
    \new_[20559]_ , \new_[20562]_ , \new_[20563]_ , \new_[20564]_ ,
    \new_[20568]_ , \new_[20569]_ , \new_[20573]_ , \new_[20574]_ ,
    \new_[20575]_ , \new_[20579]_ , \new_[20580]_ , \new_[20583]_ ,
    \new_[20586]_ , \new_[20587]_ , \new_[20588]_ , \new_[20592]_ ,
    \new_[20593]_ , \new_[20597]_ , \new_[20598]_ , \new_[20599]_ ,
    \new_[20603]_ , \new_[20604]_ , \new_[20607]_ , \new_[20610]_ ,
    \new_[20611]_ , \new_[20612]_ , \new_[20616]_ , \new_[20617]_ ,
    \new_[20621]_ , \new_[20622]_ , \new_[20623]_ , \new_[20627]_ ,
    \new_[20628]_ , \new_[20631]_ , \new_[20634]_ , \new_[20635]_ ,
    \new_[20636]_ , \new_[20640]_ , \new_[20641]_ , \new_[20645]_ ,
    \new_[20646]_ , \new_[20647]_ , \new_[20651]_ , \new_[20652]_ ,
    \new_[20655]_ , \new_[20658]_ , \new_[20659]_ , \new_[20660]_ ,
    \new_[20664]_ , \new_[20665]_ , \new_[20669]_ , \new_[20670]_ ,
    \new_[20671]_ , \new_[20675]_ , \new_[20676]_ , \new_[20679]_ ,
    \new_[20682]_ , \new_[20683]_ , \new_[20684]_ , \new_[20688]_ ,
    \new_[20689]_ , \new_[20693]_ , \new_[20694]_ , \new_[20695]_ ,
    \new_[20699]_ , \new_[20700]_ , \new_[20703]_ , \new_[20706]_ ,
    \new_[20707]_ , \new_[20708]_ , \new_[20712]_ , \new_[20713]_ ,
    \new_[20717]_ , \new_[20718]_ , \new_[20719]_ , \new_[20723]_ ,
    \new_[20724]_ , \new_[20727]_ , \new_[20730]_ , \new_[20731]_ ,
    \new_[20732]_ , \new_[20736]_ , \new_[20737]_ , \new_[20741]_ ,
    \new_[20742]_ , \new_[20743]_ , \new_[20747]_ , \new_[20748]_ ,
    \new_[20751]_ , \new_[20754]_ , \new_[20755]_ , \new_[20756]_ ,
    \new_[20760]_ , \new_[20761]_ , \new_[20765]_ , \new_[20766]_ ,
    \new_[20767]_ , \new_[20771]_ , \new_[20772]_ , \new_[20775]_ ,
    \new_[20778]_ , \new_[20779]_ , \new_[20780]_ , \new_[20784]_ ,
    \new_[20785]_ , \new_[20789]_ , \new_[20790]_ , \new_[20791]_ ,
    \new_[20795]_ , \new_[20796]_ , \new_[20799]_ , \new_[20802]_ ,
    \new_[20803]_ , \new_[20804]_ , \new_[20808]_ , \new_[20809]_ ,
    \new_[20813]_ , \new_[20814]_ , \new_[20815]_ , \new_[20819]_ ,
    \new_[20820]_ , \new_[20823]_ , \new_[20826]_ , \new_[20827]_ ,
    \new_[20828]_ , \new_[20832]_ , \new_[20833]_ , \new_[20837]_ ,
    \new_[20838]_ , \new_[20839]_ , \new_[20843]_ , \new_[20844]_ ,
    \new_[20847]_ , \new_[20850]_ , \new_[20851]_ , \new_[20852]_ ,
    \new_[20856]_ , \new_[20857]_ , \new_[20861]_ , \new_[20862]_ ,
    \new_[20863]_ , \new_[20867]_ , \new_[20868]_ , \new_[20871]_ ,
    \new_[20874]_ , \new_[20875]_ , \new_[20876]_ , \new_[20880]_ ,
    \new_[20881]_ , \new_[20885]_ , \new_[20886]_ , \new_[20887]_ ,
    \new_[20891]_ , \new_[20892]_ , \new_[20895]_ , \new_[20898]_ ,
    \new_[20899]_ , \new_[20900]_ , \new_[20904]_ , \new_[20905]_ ,
    \new_[20909]_ , \new_[20910]_ , \new_[20911]_ , \new_[20915]_ ,
    \new_[20916]_ , \new_[20919]_ , \new_[20922]_ , \new_[20923]_ ,
    \new_[20924]_ , \new_[20928]_ , \new_[20929]_ , \new_[20933]_ ,
    \new_[20934]_ , \new_[20935]_ , \new_[20939]_ , \new_[20940]_ ,
    \new_[20943]_ , \new_[20946]_ , \new_[20947]_ , \new_[20948]_ ,
    \new_[20952]_ , \new_[20953]_ , \new_[20957]_ , \new_[20958]_ ,
    \new_[20959]_ , \new_[20963]_ , \new_[20964]_ , \new_[20967]_ ,
    \new_[20970]_ , \new_[20971]_ , \new_[20972]_ , \new_[20976]_ ,
    \new_[20977]_ , \new_[20981]_ , \new_[20982]_ , \new_[20983]_ ,
    \new_[20987]_ , \new_[20988]_ , \new_[20991]_ , \new_[20994]_ ,
    \new_[20995]_ , \new_[20996]_ , \new_[21000]_ , \new_[21001]_ ,
    \new_[21005]_ , \new_[21006]_ , \new_[21007]_ , \new_[21011]_ ,
    \new_[21012]_ , \new_[21015]_ , \new_[21018]_ , \new_[21019]_ ,
    \new_[21020]_ , \new_[21024]_ , \new_[21025]_ , \new_[21029]_ ,
    \new_[21030]_ , \new_[21031]_ , \new_[21035]_ , \new_[21036]_ ,
    \new_[21039]_ , \new_[21042]_ , \new_[21043]_ , \new_[21044]_ ,
    \new_[21048]_ , \new_[21049]_ , \new_[21053]_ , \new_[21054]_ ,
    \new_[21055]_ , \new_[21059]_ , \new_[21060]_ , \new_[21063]_ ,
    \new_[21066]_ , \new_[21067]_ , \new_[21068]_ , \new_[21072]_ ,
    \new_[21073]_ , \new_[21077]_ , \new_[21078]_ , \new_[21079]_ ,
    \new_[21083]_ , \new_[21084]_ , \new_[21087]_ , \new_[21090]_ ,
    \new_[21091]_ , \new_[21092]_ , \new_[21096]_ , \new_[21097]_ ,
    \new_[21101]_ , \new_[21102]_ , \new_[21103]_ , \new_[21107]_ ,
    \new_[21108]_ , \new_[21111]_ , \new_[21114]_ , \new_[21115]_ ,
    \new_[21116]_ , \new_[21120]_ , \new_[21121]_ , \new_[21125]_ ,
    \new_[21126]_ , \new_[21127]_ , \new_[21131]_ , \new_[21132]_ ,
    \new_[21135]_ , \new_[21138]_ , \new_[21139]_ , \new_[21140]_ ,
    \new_[21144]_ , \new_[21145]_ , \new_[21149]_ , \new_[21150]_ ,
    \new_[21151]_ , \new_[21155]_ , \new_[21156]_ , \new_[21159]_ ,
    \new_[21162]_ , \new_[21163]_ , \new_[21164]_ , \new_[21168]_ ,
    \new_[21169]_ , \new_[21173]_ , \new_[21174]_ , \new_[21175]_ ,
    \new_[21179]_ , \new_[21180]_ , \new_[21183]_ , \new_[21186]_ ,
    \new_[21187]_ , \new_[21188]_ , \new_[21192]_ , \new_[21193]_ ,
    \new_[21197]_ , \new_[21198]_ , \new_[21199]_ , \new_[21203]_ ,
    \new_[21204]_ , \new_[21207]_ , \new_[21210]_ , \new_[21211]_ ,
    \new_[21212]_ , \new_[21216]_ , \new_[21217]_ , \new_[21221]_ ,
    \new_[21222]_ , \new_[21223]_ , \new_[21227]_ , \new_[21228]_ ,
    \new_[21231]_ , \new_[21234]_ , \new_[21235]_ , \new_[21236]_ ,
    \new_[21240]_ , \new_[21241]_ , \new_[21245]_ , \new_[21246]_ ,
    \new_[21247]_ , \new_[21251]_ , \new_[21252]_ , \new_[21255]_ ,
    \new_[21258]_ , \new_[21259]_ , \new_[21260]_ , \new_[21264]_ ,
    \new_[21265]_ , \new_[21269]_ , \new_[21270]_ , \new_[21271]_ ,
    \new_[21275]_ , \new_[21276]_ , \new_[21279]_ , \new_[21282]_ ,
    \new_[21283]_ , \new_[21284]_ , \new_[21288]_ , \new_[21289]_ ,
    \new_[21293]_ , \new_[21294]_ , \new_[21295]_ , \new_[21299]_ ,
    \new_[21300]_ , \new_[21303]_ , \new_[21306]_ , \new_[21307]_ ,
    \new_[21308]_ , \new_[21312]_ , \new_[21313]_ , \new_[21317]_ ,
    \new_[21318]_ , \new_[21319]_ , \new_[21323]_ , \new_[21324]_ ,
    \new_[21327]_ , \new_[21330]_ , \new_[21331]_ , \new_[21332]_ ,
    \new_[21336]_ , \new_[21337]_ , \new_[21341]_ , \new_[21342]_ ,
    \new_[21343]_ , \new_[21347]_ , \new_[21348]_ , \new_[21351]_ ,
    \new_[21354]_ , \new_[21355]_ , \new_[21356]_ , \new_[21360]_ ,
    \new_[21361]_ , \new_[21365]_ , \new_[21366]_ , \new_[21367]_ ,
    \new_[21371]_ , \new_[21372]_ , \new_[21375]_ , \new_[21378]_ ,
    \new_[21379]_ , \new_[21380]_ , \new_[21384]_ , \new_[21385]_ ,
    \new_[21389]_ , \new_[21390]_ , \new_[21391]_ , \new_[21395]_ ,
    \new_[21396]_ , \new_[21399]_ , \new_[21402]_ , \new_[21403]_ ,
    \new_[21404]_ , \new_[21408]_ , \new_[21409]_ , \new_[21413]_ ,
    \new_[21414]_ , \new_[21415]_ , \new_[21419]_ , \new_[21420]_ ,
    \new_[21423]_ , \new_[21426]_ , \new_[21427]_ , \new_[21428]_ ,
    \new_[21432]_ , \new_[21433]_ , \new_[21437]_ , \new_[21438]_ ,
    \new_[21439]_ , \new_[21443]_ , \new_[21444]_ , \new_[21447]_ ,
    \new_[21450]_ , \new_[21451]_ , \new_[21452]_ , \new_[21456]_ ,
    \new_[21457]_ , \new_[21461]_ , \new_[21462]_ , \new_[21463]_ ,
    \new_[21467]_ , \new_[21468]_ , \new_[21471]_ , \new_[21474]_ ,
    \new_[21475]_ , \new_[21476]_ , \new_[21480]_ , \new_[21481]_ ,
    \new_[21485]_ , \new_[21486]_ , \new_[21487]_ , \new_[21491]_ ,
    \new_[21492]_ , \new_[21495]_ , \new_[21498]_ , \new_[21499]_ ,
    \new_[21500]_ , \new_[21504]_ , \new_[21505]_ , \new_[21509]_ ,
    \new_[21510]_ , \new_[21511]_ , \new_[21515]_ , \new_[21516]_ ,
    \new_[21519]_ , \new_[21522]_ , \new_[21523]_ , \new_[21524]_ ,
    \new_[21528]_ , \new_[21529]_ , \new_[21532]_ , \new_[21535]_ ,
    \new_[21536]_ , \new_[21537]_ , \new_[21541]_ , \new_[21542]_ ,
    \new_[21545]_ , \new_[21548]_ , \new_[21549]_ , \new_[21550]_ ,
    \new_[21554]_ , \new_[21555]_ , \new_[21558]_ , \new_[21561]_ ,
    \new_[21562]_ , \new_[21563]_ , \new_[21567]_ , \new_[21568]_ ,
    \new_[21571]_ , \new_[21574]_ , \new_[21575]_ , \new_[21576]_ ,
    \new_[21580]_ , \new_[21581]_ , \new_[21584]_ , \new_[21587]_ ,
    \new_[21588]_ , \new_[21589]_ , \new_[21593]_ , \new_[21594]_ ,
    \new_[21597]_ , \new_[21600]_ , \new_[21601]_ , \new_[21602]_ ,
    \new_[21606]_ , \new_[21607]_ , \new_[21610]_ , \new_[21613]_ ,
    \new_[21614]_ , \new_[21615]_ , \new_[21619]_ , \new_[21620]_ ,
    \new_[21623]_ , \new_[21626]_ , \new_[21627]_ , \new_[21628]_ ,
    \new_[21632]_ , \new_[21633]_ , \new_[21636]_ , \new_[21639]_ ,
    \new_[21640]_ , \new_[21641]_ , \new_[21645]_ , \new_[21646]_ ,
    \new_[21649]_ , \new_[21652]_ , \new_[21653]_ , \new_[21654]_ ,
    \new_[21658]_ , \new_[21659]_ , \new_[21662]_ , \new_[21665]_ ,
    \new_[21666]_ , \new_[21667]_ , \new_[21671]_ , \new_[21672]_ ,
    \new_[21675]_ , \new_[21678]_ , \new_[21679]_ , \new_[21680]_ ,
    \new_[21684]_ , \new_[21685]_ , \new_[21688]_ , \new_[21691]_ ,
    \new_[21692]_ , \new_[21693]_ , \new_[21697]_ , \new_[21698]_ ,
    \new_[21701]_ , \new_[21704]_ , \new_[21705]_ , \new_[21706]_ ,
    \new_[21710]_ , \new_[21711]_ , \new_[21714]_ , \new_[21717]_ ,
    \new_[21718]_ , \new_[21719]_ , \new_[21723]_ , \new_[21724]_ ,
    \new_[21727]_ , \new_[21730]_ , \new_[21731]_ , \new_[21732]_ ,
    \new_[21736]_ , \new_[21737]_ , \new_[21740]_ , \new_[21743]_ ,
    \new_[21744]_ , \new_[21745]_ , \new_[21749]_ , \new_[21750]_ ,
    \new_[21753]_ , \new_[21756]_ , \new_[21757]_ , \new_[21758]_ ,
    \new_[21762]_ , \new_[21763]_ , \new_[21766]_ , \new_[21769]_ ,
    \new_[21770]_ , \new_[21771]_ , \new_[21775]_ , \new_[21776]_ ,
    \new_[21779]_ , \new_[21782]_ , \new_[21783]_ , \new_[21784]_ ,
    \new_[21788]_ , \new_[21789]_ , \new_[21792]_ , \new_[21795]_ ,
    \new_[21796]_ , \new_[21797]_ , \new_[21801]_ , \new_[21802]_ ,
    \new_[21805]_ , \new_[21808]_ , \new_[21809]_ , \new_[21810]_ ,
    \new_[21814]_ , \new_[21815]_ , \new_[21818]_ , \new_[21821]_ ,
    \new_[21822]_ , \new_[21823]_ , \new_[21827]_ , \new_[21828]_ ,
    \new_[21831]_ , \new_[21834]_ , \new_[21835]_ , \new_[21836]_ ,
    \new_[21840]_ , \new_[21841]_ , \new_[21844]_ , \new_[21847]_ ,
    \new_[21848]_ , \new_[21849]_ , \new_[21853]_ , \new_[21854]_ ,
    \new_[21857]_ , \new_[21860]_ , \new_[21861]_ , \new_[21862]_ ,
    \new_[21866]_ , \new_[21867]_ , \new_[21870]_ , \new_[21873]_ ,
    \new_[21874]_ , \new_[21875]_ , \new_[21879]_ , \new_[21880]_ ,
    \new_[21883]_ , \new_[21886]_ , \new_[21887]_ , \new_[21888]_ ,
    \new_[21892]_ , \new_[21893]_ , \new_[21896]_ , \new_[21899]_ ,
    \new_[21900]_ , \new_[21901]_ , \new_[21905]_ , \new_[21906]_ ,
    \new_[21909]_ , \new_[21912]_ , \new_[21913]_ , \new_[21914]_ ,
    \new_[21918]_ , \new_[21919]_ , \new_[21922]_ , \new_[21925]_ ,
    \new_[21926]_ , \new_[21927]_ , \new_[21931]_ , \new_[21932]_ ,
    \new_[21935]_ , \new_[21938]_ , \new_[21939]_ , \new_[21940]_ ,
    \new_[21944]_ , \new_[21945]_ , \new_[21948]_ , \new_[21951]_ ,
    \new_[21952]_ , \new_[21953]_ , \new_[21957]_ , \new_[21958]_ ,
    \new_[21961]_ , \new_[21964]_ , \new_[21965]_ , \new_[21966]_ ,
    \new_[21970]_ , \new_[21971]_ , \new_[21974]_ , \new_[21977]_ ,
    \new_[21978]_ , \new_[21979]_ , \new_[21983]_ , \new_[21984]_ ,
    \new_[21987]_ , \new_[21990]_ , \new_[21991]_ , \new_[21992]_ ,
    \new_[21996]_ , \new_[21997]_ , \new_[22000]_ , \new_[22003]_ ,
    \new_[22004]_ , \new_[22005]_ , \new_[22009]_ , \new_[22010]_ ,
    \new_[22013]_ , \new_[22016]_ , \new_[22017]_ , \new_[22018]_ ,
    \new_[22022]_ , \new_[22023]_ , \new_[22026]_ , \new_[22029]_ ,
    \new_[22030]_ , \new_[22031]_ , \new_[22035]_ , \new_[22036]_ ,
    \new_[22039]_ , \new_[22042]_ , \new_[22043]_ , \new_[22044]_ ,
    \new_[22048]_ , \new_[22049]_ , \new_[22052]_ , \new_[22055]_ ,
    \new_[22056]_ , \new_[22057]_ , \new_[22061]_ , \new_[22062]_ ,
    \new_[22065]_ , \new_[22068]_ , \new_[22069]_ , \new_[22070]_ ,
    \new_[22074]_ , \new_[22075]_ , \new_[22078]_ , \new_[22081]_ ,
    \new_[22082]_ , \new_[22083]_ , \new_[22087]_ , \new_[22088]_ ,
    \new_[22091]_ , \new_[22094]_ , \new_[22095]_ , \new_[22096]_ ,
    \new_[22100]_ , \new_[22101]_ , \new_[22104]_ , \new_[22107]_ ,
    \new_[22108]_ , \new_[22109]_ , \new_[22112]_ , \new_[22115]_ ,
    \new_[22116]_ , \new_[22119]_ , \new_[22122]_ , \new_[22123]_ ,
    \new_[22124]_ , \new_[22128]_ , \new_[22129]_ , \new_[22132]_ ,
    \new_[22135]_ , \new_[22136]_ , \new_[22137]_ , \new_[22140]_ ,
    \new_[22143]_ , \new_[22144]_ , \new_[22147]_ , \new_[22150]_ ,
    \new_[22151]_ , \new_[22152]_ ;
  assign A73 = \new_[3028]_  | \new_[2019]_ ;
  assign \new_[1]_  = \new_[22152]_  & \new_[22137]_ ;
  assign \new_[2]_  = \new_[22124]_  & \new_[22109]_ ;
  assign \new_[3]_  = \new_[22096]_  & \new_[22083]_ ;
  assign \new_[4]_  = \new_[22070]_  & \new_[22057]_ ;
  assign \new_[5]_  = \new_[22044]_  & \new_[22031]_ ;
  assign \new_[6]_  = \new_[22018]_  & \new_[22005]_ ;
  assign \new_[7]_  = \new_[21992]_  & \new_[21979]_ ;
  assign \new_[8]_  = \new_[21966]_  & \new_[21953]_ ;
  assign \new_[9]_  = \new_[21940]_  & \new_[21927]_ ;
  assign \new_[10]_  = \new_[21914]_  & \new_[21901]_ ;
  assign \new_[11]_  = \new_[21888]_  & \new_[21875]_ ;
  assign \new_[12]_  = \new_[21862]_  & \new_[21849]_ ;
  assign \new_[13]_  = \new_[21836]_  & \new_[21823]_ ;
  assign \new_[14]_  = \new_[21810]_  & \new_[21797]_ ;
  assign \new_[15]_  = \new_[21784]_  & \new_[21771]_ ;
  assign \new_[16]_  = \new_[21758]_  & \new_[21745]_ ;
  assign \new_[17]_  = \new_[21732]_  & \new_[21719]_ ;
  assign \new_[18]_  = \new_[21706]_  & \new_[21693]_ ;
  assign \new_[19]_  = \new_[21680]_  & \new_[21667]_ ;
  assign \new_[20]_  = \new_[21654]_  & \new_[21641]_ ;
  assign \new_[21]_  = \new_[21628]_  & \new_[21615]_ ;
  assign \new_[22]_  = \new_[21602]_  & \new_[21589]_ ;
  assign \new_[23]_  = \new_[21576]_  & \new_[21563]_ ;
  assign \new_[24]_  = \new_[21550]_  & \new_[21537]_ ;
  assign \new_[25]_  = \new_[21524]_  & \new_[21511]_ ;
  assign \new_[26]_  = \new_[21500]_  & \new_[21487]_ ;
  assign \new_[27]_  = \new_[21476]_  & \new_[21463]_ ;
  assign \new_[28]_  = \new_[21452]_  & \new_[21439]_ ;
  assign \new_[29]_  = \new_[21428]_  & \new_[21415]_ ;
  assign \new_[30]_  = \new_[21404]_  & \new_[21391]_ ;
  assign \new_[31]_  = \new_[21380]_  & \new_[21367]_ ;
  assign \new_[32]_  = \new_[21356]_  & \new_[21343]_ ;
  assign \new_[33]_  = \new_[21332]_  & \new_[21319]_ ;
  assign \new_[34]_  = \new_[21308]_  & \new_[21295]_ ;
  assign \new_[35]_  = \new_[21284]_  & \new_[21271]_ ;
  assign \new_[36]_  = \new_[21260]_  & \new_[21247]_ ;
  assign \new_[37]_  = \new_[21236]_  & \new_[21223]_ ;
  assign \new_[38]_  = \new_[21212]_  & \new_[21199]_ ;
  assign \new_[39]_  = \new_[21188]_  & \new_[21175]_ ;
  assign \new_[40]_  = \new_[21164]_  & \new_[21151]_ ;
  assign \new_[41]_  = \new_[21140]_  & \new_[21127]_ ;
  assign \new_[42]_  = \new_[21116]_  & \new_[21103]_ ;
  assign \new_[43]_  = \new_[21092]_  & \new_[21079]_ ;
  assign \new_[44]_  = \new_[21068]_  & \new_[21055]_ ;
  assign \new_[45]_  = \new_[21044]_  & \new_[21031]_ ;
  assign \new_[46]_  = \new_[21020]_  & \new_[21007]_ ;
  assign \new_[47]_  = \new_[20996]_  & \new_[20983]_ ;
  assign \new_[48]_  = \new_[20972]_  & \new_[20959]_ ;
  assign \new_[49]_  = \new_[20948]_  & \new_[20935]_ ;
  assign \new_[50]_  = \new_[20924]_  & \new_[20911]_ ;
  assign \new_[51]_  = \new_[20900]_  & \new_[20887]_ ;
  assign \new_[52]_  = \new_[20876]_  & \new_[20863]_ ;
  assign \new_[53]_  = \new_[20852]_  & \new_[20839]_ ;
  assign \new_[54]_  = \new_[20828]_  & \new_[20815]_ ;
  assign \new_[55]_  = \new_[20804]_  & \new_[20791]_ ;
  assign \new_[56]_  = \new_[20780]_  & \new_[20767]_ ;
  assign \new_[57]_  = \new_[20756]_  & \new_[20743]_ ;
  assign \new_[58]_  = \new_[20732]_  & \new_[20719]_ ;
  assign \new_[59]_  = \new_[20708]_  & \new_[20695]_ ;
  assign \new_[60]_  = \new_[20684]_  & \new_[20671]_ ;
  assign \new_[61]_  = \new_[20660]_  & \new_[20647]_ ;
  assign \new_[62]_  = \new_[20636]_  & \new_[20623]_ ;
  assign \new_[63]_  = \new_[20612]_  & \new_[20599]_ ;
  assign \new_[64]_  = \new_[20588]_  & \new_[20575]_ ;
  assign \new_[65]_  = \new_[20564]_  & \new_[20551]_ ;
  assign \new_[66]_  = \new_[20540]_  & \new_[20527]_ ;
  assign \new_[67]_  = \new_[20516]_  & \new_[20503]_ ;
  assign \new_[68]_  = \new_[20492]_  & \new_[20479]_ ;
  assign \new_[69]_  = \new_[20468]_  & \new_[20455]_ ;
  assign \new_[70]_  = \new_[20444]_  & \new_[20431]_ ;
  assign \new_[71]_  = \new_[20420]_  & \new_[20407]_ ;
  assign \new_[72]_  = \new_[20396]_  & \new_[20383]_ ;
  assign \new_[73]_  = \new_[20372]_  & \new_[20359]_ ;
  assign \new_[74]_  = \new_[20348]_  & \new_[20335]_ ;
  assign \new_[75]_  = \new_[20324]_  & \new_[20311]_ ;
  assign \new_[76]_  = \new_[20300]_  & \new_[20287]_ ;
  assign \new_[77]_  = \new_[20276]_  & \new_[20263]_ ;
  assign \new_[78]_  = \new_[20252]_  & \new_[20239]_ ;
  assign \new_[79]_  = \new_[20228]_  & \new_[20215]_ ;
  assign \new_[80]_  = \new_[20204]_  & \new_[20191]_ ;
  assign \new_[81]_  = \new_[20180]_  & \new_[20167]_ ;
  assign \new_[82]_  = \new_[20156]_  & \new_[20143]_ ;
  assign \new_[83]_  = \new_[20132]_  & \new_[20119]_ ;
  assign \new_[84]_  = \new_[20108]_  & \new_[20095]_ ;
  assign \new_[85]_  = \new_[20084]_  & \new_[20071]_ ;
  assign \new_[86]_  = \new_[20060]_  & \new_[20047]_ ;
  assign \new_[87]_  = \new_[20036]_  & \new_[20023]_ ;
  assign \new_[88]_  = \new_[20012]_  & \new_[19999]_ ;
  assign \new_[89]_  = \new_[19988]_  & \new_[19975]_ ;
  assign \new_[90]_  = \new_[19964]_  & \new_[19951]_ ;
  assign \new_[91]_  = \new_[19940]_  & \new_[19927]_ ;
  assign \new_[92]_  = \new_[19916]_  & \new_[19903]_ ;
  assign \new_[93]_  = \new_[19892]_  & \new_[19879]_ ;
  assign \new_[94]_  = \new_[19868]_  & \new_[19855]_ ;
  assign \new_[95]_  = \new_[19844]_  & \new_[19831]_ ;
  assign \new_[96]_  = \new_[19820]_  & \new_[19807]_ ;
  assign \new_[97]_  = \new_[19796]_  & \new_[19783]_ ;
  assign \new_[98]_  = \new_[19772]_  & \new_[19759]_ ;
  assign \new_[99]_  = \new_[19748]_  & \new_[19735]_ ;
  assign \new_[100]_  = \new_[19724]_  & \new_[19711]_ ;
  assign \new_[101]_  = \new_[19700]_  & \new_[19687]_ ;
  assign \new_[102]_  = \new_[19676]_  & \new_[19663]_ ;
  assign \new_[103]_  = \new_[19652]_  & \new_[19639]_ ;
  assign \new_[104]_  = \new_[19628]_  & \new_[19615]_ ;
  assign \new_[105]_  = \new_[19604]_  & \new_[19591]_ ;
  assign \new_[106]_  = \new_[19580]_  & \new_[19567]_ ;
  assign \new_[107]_  = \new_[19556]_  & \new_[19543]_ ;
  assign \new_[108]_  = \new_[19532]_  & \new_[19519]_ ;
  assign \new_[109]_  = \new_[19508]_  & \new_[19495]_ ;
  assign \new_[110]_  = \new_[19484]_  & \new_[19471]_ ;
  assign \new_[111]_  = \new_[19460]_  & \new_[19447]_ ;
  assign \new_[112]_  = \new_[19436]_  & \new_[19423]_ ;
  assign \new_[113]_  = \new_[19412]_  & \new_[19399]_ ;
  assign \new_[114]_  = \new_[19388]_  & \new_[19375]_ ;
  assign \new_[115]_  = \new_[19364]_  & \new_[19351]_ ;
  assign \new_[116]_  = \new_[19340]_  & \new_[19327]_ ;
  assign \new_[117]_  = \new_[19316]_  & \new_[19303]_ ;
  assign \new_[118]_  = \new_[19292]_  & \new_[19281]_ ;
  assign \new_[119]_  = \new_[19270]_  & \new_[19259]_ ;
  assign \new_[120]_  = \new_[19248]_  & \new_[19237]_ ;
  assign \new_[121]_  = \new_[19226]_  & \new_[19215]_ ;
  assign \new_[122]_  = \new_[19204]_  & \new_[19193]_ ;
  assign \new_[123]_  = \new_[19182]_  & \new_[19171]_ ;
  assign \new_[124]_  = \new_[19160]_  & \new_[19149]_ ;
  assign \new_[125]_  = \new_[19138]_  & \new_[19127]_ ;
  assign \new_[126]_  = \new_[19116]_  & \new_[19105]_ ;
  assign \new_[127]_  = \new_[19094]_  & \new_[19083]_ ;
  assign \new_[128]_  = \new_[19072]_  & \new_[19061]_ ;
  assign \new_[129]_  = \new_[19050]_  & \new_[19039]_ ;
  assign \new_[130]_  = \new_[19028]_  & \new_[19017]_ ;
  assign \new_[131]_  = \new_[19006]_  & \new_[18995]_ ;
  assign \new_[132]_  = \new_[18984]_  & \new_[18973]_ ;
  assign \new_[133]_  = \new_[18962]_  & \new_[18951]_ ;
  assign \new_[134]_  = \new_[18940]_  & \new_[18929]_ ;
  assign \new_[135]_  = \new_[18918]_  & \new_[18907]_ ;
  assign \new_[136]_  = \new_[18896]_  & \new_[18885]_ ;
  assign \new_[137]_  = \new_[18874]_  & \new_[18863]_ ;
  assign \new_[138]_  = \new_[18852]_  & \new_[18841]_ ;
  assign \new_[139]_  = \new_[18830]_  & \new_[18819]_ ;
  assign \new_[140]_  = \new_[18808]_  & \new_[18797]_ ;
  assign \new_[141]_  = \new_[18786]_  & \new_[18775]_ ;
  assign \new_[142]_  = \new_[18764]_  & \new_[18753]_ ;
  assign \new_[143]_  = \new_[18742]_  & \new_[18731]_ ;
  assign \new_[144]_  = \new_[18720]_  & \new_[18709]_ ;
  assign \new_[145]_  = \new_[18698]_  & \new_[18687]_ ;
  assign \new_[146]_  = \new_[18676]_  & \new_[18665]_ ;
  assign \new_[147]_  = \new_[18654]_  & \new_[18643]_ ;
  assign \new_[148]_  = \new_[18632]_  & \new_[18621]_ ;
  assign \new_[149]_  = \new_[18610]_  & \new_[18599]_ ;
  assign \new_[150]_  = \new_[18588]_  & \new_[18577]_ ;
  assign \new_[151]_  = \new_[18566]_  & \new_[18555]_ ;
  assign \new_[152]_  = \new_[18544]_  & \new_[18533]_ ;
  assign \new_[153]_  = \new_[18522]_  & \new_[18511]_ ;
  assign \new_[154]_  = \new_[18500]_  & \new_[18489]_ ;
  assign \new_[155]_  = \new_[18478]_  & \new_[18467]_ ;
  assign \new_[156]_  = \new_[18456]_  & \new_[18445]_ ;
  assign \new_[157]_  = \new_[18434]_  & \new_[18423]_ ;
  assign \new_[158]_  = \new_[18412]_  & \new_[18401]_ ;
  assign \new_[159]_  = \new_[18390]_  & \new_[18379]_ ;
  assign \new_[160]_  = \new_[18368]_  & \new_[18357]_ ;
  assign \new_[161]_  = \new_[18346]_  & \new_[18335]_ ;
  assign \new_[162]_  = \new_[18324]_  & \new_[18313]_ ;
  assign \new_[163]_  = \new_[18302]_  & \new_[18291]_ ;
  assign \new_[164]_  = \new_[18280]_  & \new_[18269]_ ;
  assign \new_[165]_  = \new_[18258]_  & \new_[18247]_ ;
  assign \new_[166]_  = \new_[18236]_  & \new_[18225]_ ;
  assign \new_[167]_  = \new_[18214]_  & \new_[18203]_ ;
  assign \new_[168]_  = \new_[18192]_  & \new_[18181]_ ;
  assign \new_[169]_  = \new_[18170]_  & \new_[18159]_ ;
  assign \new_[170]_  = \new_[18148]_  & \new_[18137]_ ;
  assign \new_[171]_  = \new_[18126]_  & \new_[18115]_ ;
  assign \new_[172]_  = \new_[18104]_  & \new_[18093]_ ;
  assign \new_[173]_  = \new_[18082]_  & \new_[18071]_ ;
  assign \new_[174]_  = \new_[18060]_  & \new_[18049]_ ;
  assign \new_[175]_  = \new_[18038]_  & \new_[18027]_ ;
  assign \new_[176]_  = \new_[18016]_  & \new_[18005]_ ;
  assign \new_[177]_  = \new_[17994]_  & \new_[17983]_ ;
  assign \new_[178]_  = \new_[17972]_  & \new_[17961]_ ;
  assign \new_[179]_  = \new_[17950]_  & \new_[17939]_ ;
  assign \new_[180]_  = \new_[17928]_  & \new_[17917]_ ;
  assign \new_[181]_  = \new_[17906]_  & \new_[17895]_ ;
  assign \new_[182]_  = \new_[17884]_  & \new_[17873]_ ;
  assign \new_[183]_  = \new_[17862]_  & \new_[17851]_ ;
  assign \new_[184]_  = \new_[17840]_  & \new_[17829]_ ;
  assign \new_[185]_  = \new_[17818]_  & \new_[17807]_ ;
  assign \new_[186]_  = \new_[17796]_  & \new_[17785]_ ;
  assign \new_[187]_  = \new_[17774]_  & \new_[17763]_ ;
  assign \new_[188]_  = \new_[17752]_  & \new_[17741]_ ;
  assign \new_[189]_  = \new_[17730]_  & \new_[17719]_ ;
  assign \new_[190]_  = \new_[17708]_  & \new_[17697]_ ;
  assign \new_[191]_  = \new_[17686]_  & \new_[17675]_ ;
  assign \new_[192]_  = \new_[17664]_  & \new_[17653]_ ;
  assign \new_[193]_  = \new_[17642]_  & \new_[17631]_ ;
  assign \new_[194]_  = \new_[17620]_  & \new_[17609]_ ;
  assign \new_[195]_  = \new_[17598]_  & \new_[17587]_ ;
  assign \new_[196]_  = \new_[17576]_  & \new_[17565]_ ;
  assign \new_[197]_  = \new_[17554]_  & \new_[17543]_ ;
  assign \new_[198]_  = \new_[17532]_  & \new_[17521]_ ;
  assign \new_[199]_  = \new_[17510]_  & \new_[17499]_ ;
  assign \new_[200]_  = \new_[17488]_  & \new_[17477]_ ;
  assign \new_[201]_  = \new_[17466]_  & \new_[17455]_ ;
  assign \new_[202]_  = \new_[17444]_  & \new_[17433]_ ;
  assign \new_[203]_  = \new_[17422]_  & \new_[17411]_ ;
  assign \new_[204]_  = \new_[17400]_  & \new_[17389]_ ;
  assign \new_[205]_  = \new_[17378]_  & \new_[17367]_ ;
  assign \new_[206]_  = \new_[17356]_  & \new_[17345]_ ;
  assign \new_[207]_  = \new_[17334]_  & \new_[17323]_ ;
  assign \new_[208]_  = \new_[17312]_  & \new_[17301]_ ;
  assign \new_[209]_  = \new_[17290]_  & \new_[17279]_ ;
  assign \new_[210]_  = \new_[17268]_  & \new_[17257]_ ;
  assign \new_[211]_  = \new_[17246]_  & \new_[17235]_ ;
  assign \new_[212]_  = \new_[17224]_  & \new_[17213]_ ;
  assign \new_[213]_  = \new_[17202]_  & \new_[17191]_ ;
  assign \new_[214]_  = \new_[17180]_  & \new_[17169]_ ;
  assign \new_[215]_  = \new_[17158]_  & \new_[17147]_ ;
  assign \new_[216]_  = \new_[17136]_  & \new_[17125]_ ;
  assign \new_[217]_  = \new_[17114]_  & \new_[17103]_ ;
  assign \new_[218]_  = \new_[17092]_  & \new_[17081]_ ;
  assign \new_[219]_  = \new_[17070]_  & \new_[17059]_ ;
  assign \new_[220]_  = \new_[17048]_  & \new_[17037]_ ;
  assign \new_[221]_  = \new_[17026]_  & \new_[17015]_ ;
  assign \new_[222]_  = \new_[17004]_  & \new_[16993]_ ;
  assign \new_[223]_  = \new_[16982]_  & \new_[16971]_ ;
  assign \new_[224]_  = \new_[16960]_  & \new_[16949]_ ;
  assign \new_[225]_  = \new_[16938]_  & \new_[16927]_ ;
  assign \new_[226]_  = \new_[16916]_  & \new_[16905]_ ;
  assign \new_[227]_  = \new_[16894]_  & \new_[16883]_ ;
  assign \new_[228]_  = \new_[16872]_  & \new_[16861]_ ;
  assign \new_[229]_  = \new_[16850]_  & \new_[16839]_ ;
  assign \new_[230]_  = \new_[16828]_  & \new_[16817]_ ;
  assign \new_[231]_  = \new_[16806]_  & \new_[16795]_ ;
  assign \new_[232]_  = \new_[16784]_  & \new_[16773]_ ;
  assign \new_[233]_  = \new_[16762]_  & \new_[16751]_ ;
  assign \new_[234]_  = \new_[16740]_  & \new_[16729]_ ;
  assign \new_[235]_  = \new_[16718]_  & \new_[16707]_ ;
  assign \new_[236]_  = \new_[16696]_  & \new_[16685]_ ;
  assign \new_[237]_  = \new_[16674]_  & \new_[16663]_ ;
  assign \new_[238]_  = \new_[16652]_  & \new_[16641]_ ;
  assign \new_[239]_  = \new_[16630]_  & \new_[16619]_ ;
  assign \new_[240]_  = \new_[16608]_  & \new_[16597]_ ;
  assign \new_[241]_  = \new_[16586]_  & \new_[16575]_ ;
  assign \new_[242]_  = \new_[16564]_  & \new_[16553]_ ;
  assign \new_[243]_  = \new_[16542]_  & \new_[16531]_ ;
  assign \new_[244]_  = \new_[16520]_  & \new_[16509]_ ;
  assign \new_[245]_  = \new_[16498]_  & \new_[16487]_ ;
  assign \new_[246]_  = \new_[16476]_  & \new_[16465]_ ;
  assign \new_[247]_  = \new_[16454]_  & \new_[16443]_ ;
  assign \new_[248]_  = \new_[16432]_  & \new_[16421]_ ;
  assign \new_[249]_  = \new_[16410]_  & \new_[16399]_ ;
  assign \new_[250]_  = \new_[16388]_  & \new_[16377]_ ;
  assign \new_[251]_  = \new_[16366]_  & \new_[16355]_ ;
  assign \new_[252]_  = \new_[16344]_  & \new_[16333]_ ;
  assign \new_[253]_  = \new_[16322]_  & \new_[16311]_ ;
  assign \new_[254]_  = \new_[16300]_  & \new_[16289]_ ;
  assign \new_[255]_  = \new_[16278]_  & \new_[16267]_ ;
  assign \new_[256]_  = \new_[16256]_  & \new_[16245]_ ;
  assign \new_[257]_  = \new_[16234]_  & \new_[16223]_ ;
  assign \new_[258]_  = \new_[16212]_  & \new_[16201]_ ;
  assign \new_[259]_  = \new_[16190]_  & \new_[16179]_ ;
  assign \new_[260]_  = \new_[16168]_  & \new_[16157]_ ;
  assign \new_[261]_  = \new_[16146]_  & \new_[16135]_ ;
  assign \new_[262]_  = \new_[16124]_  & \new_[16113]_ ;
  assign \new_[263]_  = \new_[16102]_  & \new_[16091]_ ;
  assign \new_[264]_  = \new_[16080]_  & \new_[16069]_ ;
  assign \new_[265]_  = \new_[16058]_  & \new_[16047]_ ;
  assign \new_[266]_  = \new_[16036]_  & \new_[16025]_ ;
  assign \new_[267]_  = \new_[16014]_  & \new_[16003]_ ;
  assign \new_[268]_  = \new_[15992]_  & \new_[15981]_ ;
  assign \new_[269]_  = \new_[15970]_  & \new_[15959]_ ;
  assign \new_[270]_  = \new_[15948]_  & \new_[15937]_ ;
  assign \new_[271]_  = \new_[15926]_  & \new_[15915]_ ;
  assign \new_[272]_  = \new_[15904]_  & \new_[15893]_ ;
  assign \new_[273]_  = \new_[15882]_  & \new_[15871]_ ;
  assign \new_[274]_  = \new_[15860]_  & \new_[15849]_ ;
  assign \new_[275]_  = \new_[15838]_  & \new_[15827]_ ;
  assign \new_[276]_  = \new_[15816]_  & \new_[15805]_ ;
  assign \new_[277]_  = \new_[15794]_  & \new_[15783]_ ;
  assign \new_[278]_  = \new_[15772]_  & \new_[15761]_ ;
  assign \new_[279]_  = \new_[15750]_  & \new_[15739]_ ;
  assign \new_[280]_  = \new_[15728]_  & \new_[15717]_ ;
  assign \new_[281]_  = \new_[15706]_  & \new_[15695]_ ;
  assign \new_[282]_  = \new_[15684]_  & \new_[15673]_ ;
  assign \new_[283]_  = \new_[15662]_  & \new_[15651]_ ;
  assign \new_[284]_  = \new_[15640]_  & \new_[15629]_ ;
  assign \new_[285]_  = \new_[15618]_  & \new_[15607]_ ;
  assign \new_[286]_  = \new_[15596]_  & \new_[15585]_ ;
  assign \new_[287]_  = \new_[15574]_  & \new_[15563]_ ;
  assign \new_[288]_  = \new_[15552]_  & \new_[15541]_ ;
  assign \new_[289]_  = \new_[15530]_  & \new_[15519]_ ;
  assign \new_[290]_  = \new_[15508]_  & \new_[15497]_ ;
  assign \new_[291]_  = \new_[15486]_  & \new_[15475]_ ;
  assign \new_[292]_  = \new_[15464]_  & \new_[15453]_ ;
  assign \new_[293]_  = \new_[15442]_  & \new_[15431]_ ;
  assign \new_[294]_  = \new_[15420]_  & \new_[15409]_ ;
  assign \new_[295]_  = \new_[15398]_  & \new_[15387]_ ;
  assign \new_[296]_  = \new_[15376]_  & \new_[15365]_ ;
  assign \new_[297]_  = \new_[15354]_  & \new_[15343]_ ;
  assign \new_[298]_  = \new_[15332]_  & \new_[15321]_ ;
  assign \new_[299]_  = \new_[15310]_  & \new_[15299]_ ;
  assign \new_[300]_  = \new_[15288]_  & \new_[15277]_ ;
  assign \new_[301]_  = \new_[15266]_  & \new_[15255]_ ;
  assign \new_[302]_  = \new_[15244]_  & \new_[15233]_ ;
  assign \new_[303]_  = \new_[15222]_  & \new_[15211]_ ;
  assign \new_[304]_  = \new_[15200]_  & \new_[15189]_ ;
  assign \new_[305]_  = \new_[15178]_  & \new_[15167]_ ;
  assign \new_[306]_  = \new_[15156]_  & \new_[15145]_ ;
  assign \new_[307]_  = \new_[15134]_  & \new_[15123]_ ;
  assign \new_[308]_  = \new_[15112]_  & \new_[15101]_ ;
  assign \new_[309]_  = \new_[15090]_  & \new_[15079]_ ;
  assign \new_[310]_  = \new_[15068]_  & \new_[15057]_ ;
  assign \new_[311]_  = \new_[15046]_  & \new_[15035]_ ;
  assign \new_[312]_  = \new_[15024]_  & \new_[15013]_ ;
  assign \new_[313]_  = \new_[15002]_  & \new_[14991]_ ;
  assign \new_[314]_  = \new_[14980]_  & \new_[14969]_ ;
  assign \new_[315]_  = \new_[14958]_  & \new_[14947]_ ;
  assign \new_[316]_  = \new_[14936]_  & \new_[14925]_ ;
  assign \new_[317]_  = \new_[14916]_  & \new_[14905]_ ;
  assign \new_[318]_  = \new_[14896]_  & \new_[14885]_ ;
  assign \new_[319]_  = \new_[14876]_  & \new_[14865]_ ;
  assign \new_[320]_  = \new_[14856]_  & \new_[14845]_ ;
  assign \new_[321]_  = \new_[14836]_  & \new_[14825]_ ;
  assign \new_[322]_  = \new_[14816]_  & \new_[14805]_ ;
  assign \new_[323]_  = \new_[14796]_  & \new_[14785]_ ;
  assign \new_[324]_  = \new_[14776]_  & \new_[14765]_ ;
  assign \new_[325]_  = \new_[14756]_  & \new_[14745]_ ;
  assign \new_[326]_  = \new_[14736]_  & \new_[14725]_ ;
  assign \new_[327]_  = \new_[14716]_  & \new_[14705]_ ;
  assign \new_[328]_  = \new_[14696]_  & \new_[14685]_ ;
  assign \new_[329]_  = \new_[14676]_  & \new_[14665]_ ;
  assign \new_[330]_  = \new_[14656]_  & \new_[14645]_ ;
  assign \new_[331]_  = \new_[14636]_  & \new_[14625]_ ;
  assign \new_[332]_  = \new_[14616]_  & \new_[14605]_ ;
  assign \new_[333]_  = \new_[14596]_  & \new_[14585]_ ;
  assign \new_[334]_  = \new_[14576]_  & \new_[14565]_ ;
  assign \new_[335]_  = \new_[14556]_  & \new_[14545]_ ;
  assign \new_[336]_  = \new_[14536]_  & \new_[14525]_ ;
  assign \new_[337]_  = \new_[14516]_  & \new_[14505]_ ;
  assign \new_[338]_  = \new_[14496]_  & \new_[14485]_ ;
  assign \new_[339]_  = \new_[14476]_  & \new_[14465]_ ;
  assign \new_[340]_  = \new_[14456]_  & \new_[14445]_ ;
  assign \new_[341]_  = \new_[14436]_  & \new_[14425]_ ;
  assign \new_[342]_  = \new_[14416]_  & \new_[14405]_ ;
  assign \new_[343]_  = \new_[14396]_  & \new_[14385]_ ;
  assign \new_[344]_  = \new_[14376]_  & \new_[14365]_ ;
  assign \new_[345]_  = \new_[14356]_  & \new_[14345]_ ;
  assign \new_[346]_  = \new_[14336]_  & \new_[14325]_ ;
  assign \new_[347]_  = \new_[14316]_  & \new_[14305]_ ;
  assign \new_[348]_  = \new_[14296]_  & \new_[14285]_ ;
  assign \new_[349]_  = \new_[14276]_  & \new_[14265]_ ;
  assign \new_[350]_  = \new_[14256]_  & \new_[14245]_ ;
  assign \new_[351]_  = \new_[14236]_  & \new_[14225]_ ;
  assign \new_[352]_  = \new_[14216]_  & \new_[14205]_ ;
  assign \new_[353]_  = \new_[14196]_  & \new_[14185]_ ;
  assign \new_[354]_  = \new_[14176]_  & \new_[14165]_ ;
  assign \new_[355]_  = \new_[14156]_  & \new_[14145]_ ;
  assign \new_[356]_  = \new_[14136]_  & \new_[14125]_ ;
  assign \new_[357]_  = \new_[14116]_  & \new_[14105]_ ;
  assign \new_[358]_  = \new_[14096]_  & \new_[14085]_ ;
  assign \new_[359]_  = \new_[14076]_  & \new_[14065]_ ;
  assign \new_[360]_  = \new_[14056]_  & \new_[14045]_ ;
  assign \new_[361]_  = \new_[14036]_  & \new_[14025]_ ;
  assign \new_[362]_  = \new_[14016]_  & \new_[14005]_ ;
  assign \new_[363]_  = \new_[13996]_  & \new_[13985]_ ;
  assign \new_[364]_  = \new_[13976]_  & \new_[13965]_ ;
  assign \new_[365]_  = \new_[13956]_  & \new_[13945]_ ;
  assign \new_[366]_  = \new_[13936]_  & \new_[13925]_ ;
  assign \new_[367]_  = \new_[13916]_  & \new_[13905]_ ;
  assign \new_[368]_  = \new_[13896]_  & \new_[13885]_ ;
  assign \new_[369]_  = \new_[13876]_  & \new_[13865]_ ;
  assign \new_[370]_  = \new_[13856]_  & \new_[13845]_ ;
  assign \new_[371]_  = \new_[13836]_  & \new_[13825]_ ;
  assign \new_[372]_  = \new_[13816]_  & \new_[13805]_ ;
  assign \new_[373]_  = \new_[13796]_  & \new_[13785]_ ;
  assign \new_[374]_  = \new_[13776]_  & \new_[13765]_ ;
  assign \new_[375]_  = \new_[13756]_  & \new_[13745]_ ;
  assign \new_[376]_  = \new_[13736]_  & \new_[13725]_ ;
  assign \new_[377]_  = \new_[13716]_  & \new_[13705]_ ;
  assign \new_[378]_  = \new_[13696]_  & \new_[13685]_ ;
  assign \new_[379]_  = \new_[13676]_  & \new_[13665]_ ;
  assign \new_[380]_  = \new_[13656]_  & \new_[13645]_ ;
  assign \new_[381]_  = \new_[13636]_  & \new_[13625]_ ;
  assign \new_[382]_  = \new_[13616]_  & \new_[13605]_ ;
  assign \new_[383]_  = \new_[13596]_  & \new_[13585]_ ;
  assign \new_[384]_  = \new_[13576]_  & \new_[13565]_ ;
  assign \new_[385]_  = \new_[13556]_  & \new_[13545]_ ;
  assign \new_[386]_  = \new_[13536]_  & \new_[13525]_ ;
  assign \new_[387]_  = \new_[13516]_  & \new_[13505]_ ;
  assign \new_[388]_  = \new_[13496]_  & \new_[13485]_ ;
  assign \new_[389]_  = \new_[13476]_  & \new_[13465]_ ;
  assign \new_[390]_  = \new_[13456]_  & \new_[13445]_ ;
  assign \new_[391]_  = \new_[13436]_  & \new_[13425]_ ;
  assign \new_[392]_  = \new_[13416]_  & \new_[13405]_ ;
  assign \new_[393]_  = \new_[13396]_  & \new_[13385]_ ;
  assign \new_[394]_  = \new_[13376]_  & \new_[13365]_ ;
  assign \new_[395]_  = \new_[13356]_  & \new_[13345]_ ;
  assign \new_[396]_  = \new_[13336]_  & \new_[13325]_ ;
  assign \new_[397]_  = \new_[13316]_  & \new_[13305]_ ;
  assign \new_[398]_  = \new_[13296]_  & \new_[13285]_ ;
  assign \new_[399]_  = \new_[13276]_  & \new_[13265]_ ;
  assign \new_[400]_  = \new_[13256]_  & \new_[13245]_ ;
  assign \new_[401]_  = \new_[13236]_  & \new_[13225]_ ;
  assign \new_[402]_  = \new_[13216]_  & \new_[13205]_ ;
  assign \new_[403]_  = \new_[13196]_  & \new_[13185]_ ;
  assign \new_[404]_  = \new_[13176]_  & \new_[13165]_ ;
  assign \new_[405]_  = \new_[13156]_  & \new_[13145]_ ;
  assign \new_[406]_  = \new_[13136]_  & \new_[13125]_ ;
  assign \new_[407]_  = \new_[13116]_  & \new_[13105]_ ;
  assign \new_[408]_  = \new_[13096]_  & \new_[13085]_ ;
  assign \new_[409]_  = \new_[13076]_  & \new_[13065]_ ;
  assign \new_[410]_  = \new_[13056]_  & \new_[13045]_ ;
  assign \new_[411]_  = \new_[13036]_  & \new_[13025]_ ;
  assign \new_[412]_  = \new_[13016]_  & \new_[13005]_ ;
  assign \new_[413]_  = \new_[12996]_  & \new_[12985]_ ;
  assign \new_[414]_  = \new_[12976]_  & \new_[12965]_ ;
  assign \new_[415]_  = \new_[12956]_  & \new_[12945]_ ;
  assign \new_[416]_  = \new_[12936]_  & \new_[12925]_ ;
  assign \new_[417]_  = \new_[12916]_  & \new_[12905]_ ;
  assign \new_[418]_  = \new_[12896]_  & \new_[12885]_ ;
  assign \new_[419]_  = \new_[12876]_  & \new_[12865]_ ;
  assign \new_[420]_  = \new_[12856]_  & \new_[12845]_ ;
  assign \new_[421]_  = \new_[12836]_  & \new_[12825]_ ;
  assign \new_[422]_  = \new_[12816]_  & \new_[12805]_ ;
  assign \new_[423]_  = \new_[12796]_  & \new_[12785]_ ;
  assign \new_[424]_  = \new_[12776]_  & \new_[12765]_ ;
  assign \new_[425]_  = \new_[12756]_  & \new_[12745]_ ;
  assign \new_[426]_  = \new_[12736]_  & \new_[12725]_ ;
  assign \new_[427]_  = \new_[12716]_  & \new_[12705]_ ;
  assign \new_[428]_  = \new_[12696]_  & \new_[12685]_ ;
  assign \new_[429]_  = \new_[12676]_  & \new_[12665]_ ;
  assign \new_[430]_  = \new_[12656]_  & \new_[12645]_ ;
  assign \new_[431]_  = \new_[12636]_  & \new_[12625]_ ;
  assign \new_[432]_  = \new_[12616]_  & \new_[12605]_ ;
  assign \new_[433]_  = \new_[12596]_  & \new_[12585]_ ;
  assign \new_[434]_  = \new_[12576]_  & \new_[12565]_ ;
  assign \new_[435]_  = \new_[12556]_  & \new_[12545]_ ;
  assign \new_[436]_  = \new_[12536]_  & \new_[12525]_ ;
  assign \new_[437]_  = \new_[12516]_  & \new_[12505]_ ;
  assign \new_[438]_  = \new_[12496]_  & \new_[12485]_ ;
  assign \new_[439]_  = \new_[12476]_  & \new_[12465]_ ;
  assign \new_[440]_  = \new_[12456]_  & \new_[12445]_ ;
  assign \new_[441]_  = \new_[12436]_  & \new_[12425]_ ;
  assign \new_[442]_  = \new_[12416]_  & \new_[12405]_ ;
  assign \new_[443]_  = \new_[12396]_  & \new_[12385]_ ;
  assign \new_[444]_  = \new_[12376]_  & \new_[12365]_ ;
  assign \new_[445]_  = \new_[12356]_  & \new_[12345]_ ;
  assign \new_[446]_  = \new_[12336]_  & \new_[12325]_ ;
  assign \new_[447]_  = \new_[12316]_  & \new_[12305]_ ;
  assign \new_[448]_  = \new_[12296]_  & \new_[12285]_ ;
  assign \new_[449]_  = \new_[12276]_  & \new_[12265]_ ;
  assign \new_[450]_  = \new_[12256]_  & \new_[12245]_ ;
  assign \new_[451]_  = \new_[12236]_  & \new_[12225]_ ;
  assign \new_[452]_  = \new_[12216]_  & \new_[12205]_ ;
  assign \new_[453]_  = \new_[12196]_  & \new_[12185]_ ;
  assign \new_[454]_  = \new_[12176]_  & \new_[12165]_ ;
  assign \new_[455]_  = \new_[12156]_  & \new_[12145]_ ;
  assign \new_[456]_  = \new_[12136]_  & \new_[12125]_ ;
  assign \new_[457]_  = \new_[12116]_  & \new_[12105]_ ;
  assign \new_[458]_  = \new_[12096]_  & \new_[12085]_ ;
  assign \new_[459]_  = \new_[12076]_  & \new_[12065]_ ;
  assign \new_[460]_  = \new_[12056]_  & \new_[12045]_ ;
  assign \new_[461]_  = \new_[12036]_  & \new_[12025]_ ;
  assign \new_[462]_  = \new_[12016]_  & \new_[12005]_ ;
  assign \new_[463]_  = \new_[11996]_  & \new_[11985]_ ;
  assign \new_[464]_  = \new_[11976]_  & \new_[11965]_ ;
  assign \new_[465]_  = \new_[11956]_  & \new_[11945]_ ;
  assign \new_[466]_  = \new_[11936]_  & \new_[11925]_ ;
  assign \new_[467]_  = \new_[11916]_  & \new_[11905]_ ;
  assign \new_[468]_  = \new_[11896]_  & \new_[11885]_ ;
  assign \new_[469]_  = \new_[11876]_  & \new_[11865]_ ;
  assign \new_[470]_  = \new_[11856]_  & \new_[11845]_ ;
  assign \new_[471]_  = \new_[11836]_  & \new_[11825]_ ;
  assign \new_[472]_  = \new_[11816]_  & \new_[11805]_ ;
  assign \new_[473]_  = \new_[11796]_  & \new_[11785]_ ;
  assign \new_[474]_  = \new_[11776]_  & \new_[11765]_ ;
  assign \new_[475]_  = \new_[11756]_  & \new_[11745]_ ;
  assign \new_[476]_  = \new_[11736]_  & \new_[11725]_ ;
  assign \new_[477]_  = \new_[11716]_  & \new_[11705]_ ;
  assign \new_[478]_  = \new_[11696]_  & \new_[11685]_ ;
  assign \new_[479]_  = \new_[11676]_  & \new_[11665]_ ;
  assign \new_[480]_  = \new_[11656]_  & \new_[11645]_ ;
  assign \new_[481]_  = \new_[11636]_  & \new_[11625]_ ;
  assign \new_[482]_  = \new_[11616]_  & \new_[11605]_ ;
  assign \new_[483]_  = \new_[11596]_  & \new_[11585]_ ;
  assign \new_[484]_  = \new_[11576]_  & \new_[11565]_ ;
  assign \new_[485]_  = \new_[11556]_  & \new_[11545]_ ;
  assign \new_[486]_  = \new_[11536]_  & \new_[11525]_ ;
  assign \new_[487]_  = \new_[11516]_  & \new_[11505]_ ;
  assign \new_[488]_  = \new_[11496]_  & \new_[11485]_ ;
  assign \new_[489]_  = \new_[11476]_  & \new_[11465]_ ;
  assign \new_[490]_  = \new_[11456]_  & \new_[11445]_ ;
  assign \new_[491]_  = \new_[11436]_  & \new_[11425]_ ;
  assign \new_[492]_  = \new_[11416]_  & \new_[11405]_ ;
  assign \new_[493]_  = \new_[11396]_  & \new_[11385]_ ;
  assign \new_[494]_  = \new_[11376]_  & \new_[11365]_ ;
  assign \new_[495]_  = \new_[11356]_  & \new_[11345]_ ;
  assign \new_[496]_  = \new_[11336]_  & \new_[11325]_ ;
  assign \new_[497]_  = \new_[11316]_  & \new_[11305]_ ;
  assign \new_[498]_  = \new_[11296]_  & \new_[11285]_ ;
  assign \new_[499]_  = \new_[11276]_  & \new_[11265]_ ;
  assign \new_[500]_  = \new_[11256]_  & \new_[11245]_ ;
  assign \new_[501]_  = \new_[11236]_  & \new_[11225]_ ;
  assign \new_[502]_  = \new_[11216]_  & \new_[11205]_ ;
  assign \new_[503]_  = \new_[11196]_  & \new_[11185]_ ;
  assign \new_[504]_  = \new_[11176]_  & \new_[11165]_ ;
  assign \new_[505]_  = \new_[11156]_  & \new_[11145]_ ;
  assign \new_[506]_  = \new_[11136]_  & \new_[11125]_ ;
  assign \new_[507]_  = \new_[11116]_  & \new_[11105]_ ;
  assign \new_[508]_  = \new_[11096]_  & \new_[11085]_ ;
  assign \new_[509]_  = \new_[11076]_  & \new_[11065]_ ;
  assign \new_[510]_  = \new_[11056]_  & \new_[11045]_ ;
  assign \new_[511]_  = \new_[11036]_  & \new_[11025]_ ;
  assign \new_[512]_  = \new_[11016]_  & \new_[11005]_ ;
  assign \new_[513]_  = \new_[10996]_  & \new_[10985]_ ;
  assign \new_[514]_  = \new_[10976]_  & \new_[10965]_ ;
  assign \new_[515]_  = \new_[10956]_  & \new_[10945]_ ;
  assign \new_[516]_  = \new_[10936]_  & \new_[10925]_ ;
  assign \new_[517]_  = \new_[10916]_  & \new_[10905]_ ;
  assign \new_[518]_  = \new_[10896]_  & \new_[10885]_ ;
  assign \new_[519]_  = \new_[10876]_  & \new_[10865]_ ;
  assign \new_[520]_  = \new_[10856]_  & \new_[10845]_ ;
  assign \new_[521]_  = \new_[10836]_  & \new_[10825]_ ;
  assign \new_[522]_  = \new_[10816]_  & \new_[10805]_ ;
  assign \new_[523]_  = \new_[10796]_  & \new_[10785]_ ;
  assign \new_[524]_  = \new_[10776]_  & \new_[10765]_ ;
  assign \new_[525]_  = \new_[10756]_  & \new_[10745]_ ;
  assign \new_[526]_  = \new_[10736]_  & \new_[10725]_ ;
  assign \new_[527]_  = \new_[10716]_  & \new_[10705]_ ;
  assign \new_[528]_  = \new_[10696]_  & \new_[10685]_ ;
  assign \new_[529]_  = \new_[10676]_  & \new_[10665]_ ;
  assign \new_[530]_  = \new_[10656]_  & \new_[10645]_ ;
  assign \new_[531]_  = \new_[10636]_  & \new_[10625]_ ;
  assign \new_[532]_  = \new_[10616]_  & \new_[10605]_ ;
  assign \new_[533]_  = \new_[10596]_  & \new_[10585]_ ;
  assign \new_[534]_  = \new_[10576]_  & \new_[10565]_ ;
  assign \new_[535]_  = \new_[10556]_  & \new_[10545]_ ;
  assign \new_[536]_  = \new_[10536]_  & \new_[10525]_ ;
  assign \new_[537]_  = \new_[10516]_  & \new_[10505]_ ;
  assign \new_[538]_  = \new_[10496]_  & \new_[10485]_ ;
  assign \new_[539]_  = \new_[10476]_  & \new_[10465]_ ;
  assign \new_[540]_  = \new_[10456]_  & \new_[10445]_ ;
  assign \new_[541]_  = \new_[10436]_  & \new_[10425]_ ;
  assign \new_[542]_  = \new_[10416]_  & \new_[10405]_ ;
  assign \new_[543]_  = \new_[10396]_  & \new_[10385]_ ;
  assign \new_[544]_  = \new_[10376]_  & \new_[10365]_ ;
  assign \new_[545]_  = \new_[10356]_  & \new_[10345]_ ;
  assign \new_[546]_  = \new_[10336]_  & \new_[10325]_ ;
  assign \new_[547]_  = \new_[10316]_  & \new_[10305]_ ;
  assign \new_[548]_  = \new_[10296]_  & \new_[10285]_ ;
  assign \new_[549]_  = \new_[10276]_  & \new_[10265]_ ;
  assign \new_[550]_  = \new_[10256]_  & \new_[10245]_ ;
  assign \new_[551]_  = \new_[10236]_  & \new_[10225]_ ;
  assign \new_[552]_  = \new_[10216]_  & \new_[10205]_ ;
  assign \new_[553]_  = \new_[10196]_  & \new_[10185]_ ;
  assign \new_[554]_  = \new_[10176]_  & \new_[10165]_ ;
  assign \new_[555]_  = \new_[10156]_  & \new_[10145]_ ;
  assign \new_[556]_  = \new_[10136]_  & \new_[10125]_ ;
  assign \new_[557]_  = \new_[10116]_  & \new_[10105]_ ;
  assign \new_[558]_  = \new_[10096]_  & \new_[10085]_ ;
  assign \new_[559]_  = \new_[10076]_  & \new_[10065]_ ;
  assign \new_[560]_  = \new_[10056]_  & \new_[10045]_ ;
  assign \new_[561]_  = \new_[10036]_  & \new_[10025]_ ;
  assign \new_[562]_  = \new_[10016]_  & \new_[10005]_ ;
  assign \new_[563]_  = \new_[9996]_  & \new_[9985]_ ;
  assign \new_[564]_  = \new_[9976]_  & \new_[9967]_ ;
  assign \new_[565]_  = \new_[9958]_  & \new_[9949]_ ;
  assign \new_[566]_  = \new_[9940]_  & \new_[9931]_ ;
  assign \new_[567]_  = \new_[9922]_  & \new_[9913]_ ;
  assign \new_[568]_  = \new_[9904]_  & \new_[9895]_ ;
  assign \new_[569]_  = \new_[9886]_  & \new_[9877]_ ;
  assign \new_[570]_  = \new_[9868]_  & \new_[9859]_ ;
  assign \new_[571]_  = \new_[9850]_  & \new_[9841]_ ;
  assign \new_[572]_  = \new_[9832]_  & \new_[9823]_ ;
  assign \new_[573]_  = \new_[9814]_  & \new_[9805]_ ;
  assign \new_[574]_  = \new_[9796]_  & \new_[9787]_ ;
  assign \new_[575]_  = \new_[9778]_  & \new_[9769]_ ;
  assign \new_[576]_  = \new_[9760]_  & \new_[9751]_ ;
  assign \new_[577]_  = \new_[9742]_  & \new_[9733]_ ;
  assign \new_[578]_  = \new_[9724]_  & \new_[9715]_ ;
  assign \new_[579]_  = \new_[9706]_  & \new_[9697]_ ;
  assign \new_[580]_  = \new_[9688]_  & \new_[9679]_ ;
  assign \new_[581]_  = \new_[9670]_  & \new_[9661]_ ;
  assign \new_[582]_  = \new_[9652]_  & \new_[9643]_ ;
  assign \new_[583]_  = \new_[9634]_  & \new_[9625]_ ;
  assign \new_[584]_  = \new_[9616]_  & \new_[9607]_ ;
  assign \new_[585]_  = \new_[9598]_  & \new_[9589]_ ;
  assign \new_[586]_  = \new_[9580]_  & \new_[9571]_ ;
  assign \new_[587]_  = \new_[9562]_  & \new_[9553]_ ;
  assign \new_[588]_  = \new_[9544]_  & \new_[9535]_ ;
  assign \new_[589]_  = \new_[9526]_  & \new_[9517]_ ;
  assign \new_[590]_  = \new_[9508]_  & \new_[9499]_ ;
  assign \new_[591]_  = \new_[9490]_  & \new_[9481]_ ;
  assign \new_[592]_  = \new_[9472]_  & \new_[9463]_ ;
  assign \new_[593]_  = \new_[9454]_  & \new_[9445]_ ;
  assign \new_[594]_  = \new_[9436]_  & \new_[9427]_ ;
  assign \new_[595]_  = \new_[9418]_  & \new_[9409]_ ;
  assign \new_[596]_  = \new_[9400]_  & \new_[9391]_ ;
  assign \new_[597]_  = \new_[9382]_  & \new_[9373]_ ;
  assign \new_[598]_  = \new_[9364]_  & \new_[9355]_ ;
  assign \new_[599]_  = \new_[9346]_  & \new_[9337]_ ;
  assign \new_[600]_  = \new_[9328]_  & \new_[9319]_ ;
  assign \new_[601]_  = \new_[9310]_  & \new_[9301]_ ;
  assign \new_[602]_  = \new_[9292]_  & \new_[9283]_ ;
  assign \new_[603]_  = \new_[9274]_  & \new_[9265]_ ;
  assign \new_[604]_  = \new_[9256]_  & \new_[9247]_ ;
  assign \new_[605]_  = \new_[9238]_  & \new_[9229]_ ;
  assign \new_[606]_  = \new_[9220]_  & \new_[9211]_ ;
  assign \new_[607]_  = \new_[9202]_  & \new_[9193]_ ;
  assign \new_[608]_  = \new_[9184]_  & \new_[9175]_ ;
  assign \new_[609]_  = \new_[9166]_  & \new_[9157]_ ;
  assign \new_[610]_  = \new_[9148]_  & \new_[9139]_ ;
  assign \new_[611]_  = \new_[9130]_  & \new_[9121]_ ;
  assign \new_[612]_  = \new_[9112]_  & \new_[9103]_ ;
  assign \new_[613]_  = \new_[9094]_  & \new_[9085]_ ;
  assign \new_[614]_  = \new_[9076]_  & \new_[9067]_ ;
  assign \new_[615]_  = \new_[9058]_  & \new_[9049]_ ;
  assign \new_[616]_  = \new_[9040]_  & \new_[9031]_ ;
  assign \new_[617]_  = \new_[9022]_  & \new_[9013]_ ;
  assign \new_[618]_  = \new_[9004]_  & \new_[8995]_ ;
  assign \new_[619]_  = \new_[8986]_  & \new_[8977]_ ;
  assign \new_[620]_  = \new_[8968]_  & \new_[8959]_ ;
  assign \new_[621]_  = \new_[8950]_  & \new_[8941]_ ;
  assign \new_[622]_  = \new_[8932]_  & \new_[8923]_ ;
  assign \new_[623]_  = \new_[8914]_  & \new_[8905]_ ;
  assign \new_[624]_  = \new_[8896]_  & \new_[8887]_ ;
  assign \new_[625]_  = \new_[8878]_  & \new_[8869]_ ;
  assign \new_[626]_  = \new_[8860]_  & \new_[8851]_ ;
  assign \new_[627]_  = \new_[8842]_  & \new_[8833]_ ;
  assign \new_[628]_  = \new_[8824]_  & \new_[8815]_ ;
  assign \new_[629]_  = \new_[8806]_  & \new_[8797]_ ;
  assign \new_[630]_  = \new_[8788]_  & \new_[8779]_ ;
  assign \new_[631]_  = \new_[8770]_  & \new_[8761]_ ;
  assign \new_[632]_  = \new_[8752]_  & \new_[8743]_ ;
  assign \new_[633]_  = \new_[8734]_  & \new_[8725]_ ;
  assign \new_[634]_  = \new_[8716]_  & \new_[8707]_ ;
  assign \new_[635]_  = \new_[8698]_  & \new_[8689]_ ;
  assign \new_[636]_  = \new_[8680]_  & \new_[8671]_ ;
  assign \new_[637]_  = \new_[8662]_  & \new_[8653]_ ;
  assign \new_[638]_  = \new_[8644]_  & \new_[8635]_ ;
  assign \new_[639]_  = \new_[8626]_  & \new_[8617]_ ;
  assign \new_[640]_  = \new_[8608]_  & \new_[8599]_ ;
  assign \new_[641]_  = \new_[8590]_  & \new_[8581]_ ;
  assign \new_[642]_  = \new_[8572]_  & \new_[8563]_ ;
  assign \new_[643]_  = \new_[8554]_  & \new_[8545]_ ;
  assign \new_[644]_  = \new_[8536]_  & \new_[8527]_ ;
  assign \new_[645]_  = \new_[8518]_  & \new_[8509]_ ;
  assign \new_[646]_  = \new_[8500]_  & \new_[8491]_ ;
  assign \new_[647]_  = \new_[8482]_  & \new_[8473]_ ;
  assign \new_[648]_  = \new_[8464]_  & \new_[8455]_ ;
  assign \new_[649]_  = \new_[8446]_  & \new_[8437]_ ;
  assign \new_[650]_  = \new_[8428]_  & \new_[8419]_ ;
  assign \new_[651]_  = \new_[8410]_  & \new_[8401]_ ;
  assign \new_[652]_  = \new_[8392]_  & \new_[8383]_ ;
  assign \new_[653]_  = \new_[8374]_  & \new_[8365]_ ;
  assign \new_[654]_  = \new_[8356]_  & \new_[8347]_ ;
  assign \new_[655]_  = \new_[8338]_  & \new_[8329]_ ;
  assign \new_[656]_  = \new_[8320]_  & \new_[8311]_ ;
  assign \new_[657]_  = \new_[8302]_  & \new_[8293]_ ;
  assign \new_[658]_  = \new_[8284]_  & \new_[8275]_ ;
  assign \new_[659]_  = \new_[8266]_  & \new_[8257]_ ;
  assign \new_[660]_  = \new_[8248]_  & \new_[8239]_ ;
  assign \new_[661]_  = \new_[8230]_  & \new_[8221]_ ;
  assign \new_[662]_  = \new_[8212]_  & \new_[8203]_ ;
  assign \new_[663]_  = \new_[8194]_  & \new_[8185]_ ;
  assign \new_[664]_  = \new_[8176]_  & \new_[8167]_ ;
  assign \new_[665]_  = \new_[8158]_  & \new_[8149]_ ;
  assign \new_[666]_  = \new_[8140]_  & \new_[8131]_ ;
  assign \new_[667]_  = \new_[8122]_  & \new_[8113]_ ;
  assign \new_[668]_  = \new_[8104]_  & \new_[8095]_ ;
  assign \new_[669]_  = \new_[8086]_  & \new_[8077]_ ;
  assign \new_[670]_  = \new_[8068]_  & \new_[8059]_ ;
  assign \new_[671]_  = \new_[8050]_  & \new_[8041]_ ;
  assign \new_[672]_  = \new_[8032]_  & \new_[8023]_ ;
  assign \new_[673]_  = \new_[8014]_  & \new_[8005]_ ;
  assign \new_[674]_  = \new_[7996]_  & \new_[7987]_ ;
  assign \new_[675]_  = \new_[7978]_  & \new_[7969]_ ;
  assign \new_[676]_  = \new_[7960]_  & \new_[7951]_ ;
  assign \new_[677]_  = \new_[7942]_  & \new_[7933]_ ;
  assign \new_[678]_  = \new_[7924]_  & \new_[7915]_ ;
  assign \new_[679]_  = \new_[7906]_  & \new_[7897]_ ;
  assign \new_[680]_  = \new_[7888]_  & \new_[7879]_ ;
  assign \new_[681]_  = \new_[7870]_  & \new_[7861]_ ;
  assign \new_[682]_  = \new_[7852]_  & \new_[7843]_ ;
  assign \new_[683]_  = \new_[7834]_  & \new_[7825]_ ;
  assign \new_[684]_  = \new_[7816]_  & \new_[7807]_ ;
  assign \new_[685]_  = \new_[7798]_  & \new_[7789]_ ;
  assign \new_[686]_  = \new_[7780]_  & \new_[7771]_ ;
  assign \new_[687]_  = \new_[7762]_  & \new_[7753]_ ;
  assign \new_[688]_  = \new_[7744]_  & \new_[7735]_ ;
  assign \new_[689]_  = \new_[7726]_  & \new_[7717]_ ;
  assign \new_[690]_  = \new_[7708]_  & \new_[7699]_ ;
  assign \new_[691]_  = \new_[7690]_  & \new_[7681]_ ;
  assign \new_[692]_  = \new_[7672]_  & \new_[7663]_ ;
  assign \new_[693]_  = \new_[7654]_  & \new_[7645]_ ;
  assign \new_[694]_  = \new_[7636]_  & \new_[7627]_ ;
  assign \new_[695]_  = \new_[7618]_  & \new_[7609]_ ;
  assign \new_[696]_  = \new_[7600]_  & \new_[7591]_ ;
  assign \new_[697]_  = \new_[7582]_  & \new_[7573]_ ;
  assign \new_[698]_  = \new_[7564]_  & \new_[7555]_ ;
  assign \new_[699]_  = \new_[7546]_  & \new_[7537]_ ;
  assign \new_[700]_  = \new_[7528]_  & \new_[7519]_ ;
  assign \new_[701]_  = \new_[7510]_  & \new_[7501]_ ;
  assign \new_[702]_  = \new_[7492]_  & \new_[7483]_ ;
  assign \new_[703]_  = \new_[7474]_  & \new_[7465]_ ;
  assign \new_[704]_  = \new_[7456]_  & \new_[7447]_ ;
  assign \new_[705]_  = \new_[7438]_  & \new_[7429]_ ;
  assign \new_[706]_  = \new_[7420]_  & \new_[7411]_ ;
  assign \new_[707]_  = \new_[7402]_  & \new_[7393]_ ;
  assign \new_[708]_  = \new_[7384]_  & \new_[7375]_ ;
  assign \new_[709]_  = \new_[7366]_  & \new_[7357]_ ;
  assign \new_[710]_  = \new_[7348]_  & \new_[7339]_ ;
  assign \new_[711]_  = \new_[7330]_  & \new_[7321]_ ;
  assign \new_[712]_  = \new_[7312]_  & \new_[7303]_ ;
  assign \new_[713]_  = \new_[7294]_  & \new_[7285]_ ;
  assign \new_[714]_  = \new_[7276]_  & \new_[7267]_ ;
  assign \new_[715]_  = \new_[7258]_  & \new_[7249]_ ;
  assign \new_[716]_  = \new_[7240]_  & \new_[7231]_ ;
  assign \new_[717]_  = \new_[7222]_  & \new_[7213]_ ;
  assign \new_[718]_  = \new_[7204]_  & \new_[7195]_ ;
  assign \new_[719]_  = \new_[7186]_  & \new_[7177]_ ;
  assign \new_[720]_  = \new_[7168]_  & \new_[7159]_ ;
  assign \new_[721]_  = \new_[7150]_  & \new_[7141]_ ;
  assign \new_[722]_  = \new_[7132]_  & \new_[7123]_ ;
  assign \new_[723]_  = \new_[7114]_  & \new_[7105]_ ;
  assign \new_[724]_  = \new_[7096]_  & \new_[7087]_ ;
  assign \new_[725]_  = \new_[7078]_  & \new_[7069]_ ;
  assign \new_[726]_  = \new_[7060]_  & \new_[7051]_ ;
  assign \new_[727]_  = \new_[7042]_  & \new_[7033]_ ;
  assign \new_[728]_  = \new_[7024]_  & \new_[7015]_ ;
  assign \new_[729]_  = \new_[7006]_  & \new_[6997]_ ;
  assign \new_[730]_  = \new_[6988]_  & \new_[6979]_ ;
  assign \new_[731]_  = \new_[6970]_  & \new_[6961]_ ;
  assign \new_[732]_  = \new_[6952]_  & \new_[6943]_ ;
  assign \new_[733]_  = \new_[6934]_  & \new_[6925]_ ;
  assign \new_[734]_  = \new_[6916]_  & \new_[6907]_ ;
  assign \new_[735]_  = \new_[6898]_  & \new_[6889]_ ;
  assign \new_[736]_  = \new_[6880]_  & \new_[6871]_ ;
  assign \new_[737]_  = \new_[6862]_  & \new_[6853]_ ;
  assign \new_[738]_  = \new_[6844]_  & \new_[6835]_ ;
  assign \new_[739]_  = \new_[6826]_  & \new_[6817]_ ;
  assign \new_[740]_  = \new_[6808]_  & \new_[6799]_ ;
  assign \new_[741]_  = \new_[6790]_  & \new_[6781]_ ;
  assign \new_[742]_  = \new_[6772]_  & \new_[6763]_ ;
  assign \new_[743]_  = \new_[6754]_  & \new_[6745]_ ;
  assign \new_[744]_  = \new_[6736]_  & \new_[6727]_ ;
  assign \new_[745]_  = \new_[6718]_  & \new_[6709]_ ;
  assign \new_[746]_  = \new_[6700]_  & \new_[6691]_ ;
  assign \new_[747]_  = \new_[6682]_  & \new_[6673]_ ;
  assign \new_[748]_  = \new_[6664]_  & \new_[6655]_ ;
  assign \new_[749]_  = \new_[6646]_  & \new_[6637]_ ;
  assign \new_[750]_  = \new_[6628]_  & \new_[6619]_ ;
  assign \new_[751]_  = \new_[6610]_  & \new_[6601]_ ;
  assign \new_[752]_  = \new_[6592]_  & \new_[6583]_ ;
  assign \new_[753]_  = \new_[6574]_  & \new_[6565]_ ;
  assign \new_[754]_  = \new_[6556]_  & \new_[6547]_ ;
  assign \new_[755]_  = \new_[6538]_  & \new_[6529]_ ;
  assign \new_[756]_  = \new_[6520]_  & \new_[6511]_ ;
  assign \new_[757]_  = \new_[6502]_  & \new_[6493]_ ;
  assign \new_[758]_  = \new_[6484]_  & \new_[6475]_ ;
  assign \new_[759]_  = \new_[6466]_  & \new_[6457]_ ;
  assign \new_[760]_  = \new_[6448]_  & \new_[6439]_ ;
  assign \new_[761]_  = \new_[6430]_  & \new_[6421]_ ;
  assign \new_[762]_  = \new_[6412]_  & \new_[6403]_ ;
  assign \new_[763]_  = \new_[6394]_  & \new_[6385]_ ;
  assign \new_[764]_  = \new_[6376]_  & \new_[6367]_ ;
  assign \new_[765]_  = \new_[6358]_  & \new_[6349]_ ;
  assign \new_[766]_  = \new_[6340]_  & \new_[6331]_ ;
  assign \new_[767]_  = \new_[6322]_  & \new_[6313]_ ;
  assign \new_[768]_  = \new_[6304]_  & \new_[6295]_ ;
  assign \new_[769]_  = \new_[6286]_  & \new_[6277]_ ;
  assign \new_[770]_  = \new_[6268]_  & \new_[6259]_ ;
  assign \new_[771]_  = \new_[6250]_  & \new_[6241]_ ;
  assign \new_[772]_  = \new_[6232]_  & \new_[6223]_ ;
  assign \new_[773]_  = \new_[6214]_  & \new_[6205]_ ;
  assign \new_[774]_  = \new_[6196]_  & \new_[6187]_ ;
  assign \new_[775]_  = \new_[6180]_  & \new_[6171]_ ;
  assign \new_[776]_  = \new_[6164]_  & \new_[6155]_ ;
  assign \new_[777]_  = \new_[6148]_  & \new_[6139]_ ;
  assign \new_[778]_  = \new_[6132]_  & \new_[6123]_ ;
  assign \new_[779]_  = \new_[6116]_  & \new_[6107]_ ;
  assign \new_[780]_  = \new_[6100]_  & \new_[6091]_ ;
  assign \new_[781]_  = \new_[6084]_  & \new_[6075]_ ;
  assign \new_[782]_  = \new_[6068]_  & \new_[6059]_ ;
  assign \new_[783]_  = \new_[6052]_  & \new_[6043]_ ;
  assign \new_[784]_  = \new_[6036]_  & \new_[6027]_ ;
  assign \new_[785]_  = \new_[6020]_  & \new_[6011]_ ;
  assign \new_[786]_  = \new_[6004]_  & \new_[5995]_ ;
  assign \new_[787]_  = \new_[5988]_  & \new_[5979]_ ;
  assign \new_[788]_  = \new_[5972]_  & \new_[5963]_ ;
  assign \new_[789]_  = \new_[5956]_  & \new_[5947]_ ;
  assign \new_[790]_  = \new_[5940]_  & \new_[5931]_ ;
  assign \new_[791]_  = \new_[5924]_  & \new_[5915]_ ;
  assign \new_[792]_  = \new_[5908]_  & \new_[5899]_ ;
  assign \new_[793]_  = \new_[5892]_  & \new_[5883]_ ;
  assign \new_[794]_  = \new_[5876]_  & \new_[5867]_ ;
  assign \new_[795]_  = \new_[5860]_  & \new_[5851]_ ;
  assign \new_[796]_  = \new_[5844]_  & \new_[5835]_ ;
  assign \new_[797]_  = \new_[5828]_  & \new_[5819]_ ;
  assign \new_[798]_  = \new_[5812]_  & \new_[5803]_ ;
  assign \new_[799]_  = \new_[5796]_  & \new_[5787]_ ;
  assign \new_[800]_  = \new_[5780]_  & \new_[5771]_ ;
  assign \new_[801]_  = \new_[5764]_  & \new_[5755]_ ;
  assign \new_[802]_  = \new_[5748]_  & \new_[5739]_ ;
  assign \new_[803]_  = \new_[5732]_  & \new_[5723]_ ;
  assign \new_[804]_  = \new_[5716]_  & \new_[5707]_ ;
  assign \new_[805]_  = \new_[5700]_  & \new_[5691]_ ;
  assign \new_[806]_  = \new_[5684]_  & \new_[5675]_ ;
  assign \new_[807]_  = \new_[5668]_  & \new_[5659]_ ;
  assign \new_[808]_  = \new_[5652]_  & \new_[5643]_ ;
  assign \new_[809]_  = \new_[5636]_  & \new_[5627]_ ;
  assign \new_[810]_  = \new_[5620]_  & \new_[5611]_ ;
  assign \new_[811]_  = \new_[5604]_  & \new_[5595]_ ;
  assign \new_[812]_  = \new_[5588]_  & \new_[5579]_ ;
  assign \new_[813]_  = \new_[5572]_  & \new_[5563]_ ;
  assign \new_[814]_  = \new_[5556]_  & \new_[5547]_ ;
  assign \new_[815]_  = \new_[5540]_  & \new_[5531]_ ;
  assign \new_[816]_  = \new_[5524]_  & \new_[5515]_ ;
  assign \new_[817]_  = \new_[5508]_  & \new_[5499]_ ;
  assign \new_[818]_  = \new_[5492]_  & \new_[5483]_ ;
  assign \new_[819]_  = \new_[5476]_  & \new_[5467]_ ;
  assign \new_[820]_  = \new_[5460]_  & \new_[5451]_ ;
  assign \new_[821]_  = \new_[5444]_  & \new_[5435]_ ;
  assign \new_[822]_  = \new_[5428]_  & \new_[5419]_ ;
  assign \new_[823]_  = \new_[5412]_  & \new_[5403]_ ;
  assign \new_[824]_  = \new_[5396]_  & \new_[5387]_ ;
  assign \new_[825]_  = \new_[5380]_  & \new_[5371]_ ;
  assign \new_[826]_  = \new_[5364]_  & \new_[5355]_ ;
  assign \new_[827]_  = \new_[5348]_  & \new_[5339]_ ;
  assign \new_[828]_  = \new_[5332]_  & \new_[5323]_ ;
  assign \new_[829]_  = \new_[5316]_  & \new_[5307]_ ;
  assign \new_[830]_  = \new_[5300]_  & \new_[5291]_ ;
  assign \new_[831]_  = \new_[5284]_  & \new_[5275]_ ;
  assign \new_[832]_  = \new_[5268]_  & \new_[5259]_ ;
  assign \new_[833]_  = \new_[5252]_  & \new_[5243]_ ;
  assign \new_[834]_  = \new_[5236]_  & \new_[5227]_ ;
  assign \new_[835]_  = \new_[5220]_  & \new_[5211]_ ;
  assign \new_[836]_  = \new_[5204]_  & \new_[5195]_ ;
  assign \new_[837]_  = \new_[5188]_  & \new_[5179]_ ;
  assign \new_[838]_  = \new_[5172]_  & \new_[5163]_ ;
  assign \new_[839]_  = \new_[5156]_  & \new_[5147]_ ;
  assign \new_[840]_  = \new_[5140]_  & \new_[5131]_ ;
  assign \new_[841]_  = \new_[5124]_  & \new_[5115]_ ;
  assign \new_[842]_  = \new_[5108]_  & \new_[5099]_ ;
  assign \new_[843]_  = \new_[5092]_  & \new_[5083]_ ;
  assign \new_[844]_  = \new_[5076]_  & \new_[5067]_ ;
  assign \new_[845]_  = \new_[5060]_  & \new_[5051]_ ;
  assign \new_[846]_  = \new_[5044]_  & \new_[5035]_ ;
  assign \new_[847]_  = \new_[5028]_  & \new_[5019]_ ;
  assign \new_[848]_  = \new_[5012]_  & \new_[5003]_ ;
  assign \new_[849]_  = \new_[4996]_  & \new_[4987]_ ;
  assign \new_[850]_  = \new_[4980]_  & \new_[4971]_ ;
  assign \new_[851]_  = \new_[4964]_  & \new_[4955]_ ;
  assign \new_[852]_  = \new_[4948]_  & \new_[4939]_ ;
  assign \new_[853]_  = \new_[4932]_  & \new_[4923]_ ;
  assign \new_[854]_  = \new_[4916]_  & \new_[4907]_ ;
  assign \new_[855]_  = \new_[4900]_  & \new_[4891]_ ;
  assign \new_[856]_  = \new_[4884]_  & \new_[4875]_ ;
  assign \new_[857]_  = \new_[4868]_  & \new_[4859]_ ;
  assign \new_[858]_  = \new_[4852]_  & \new_[4843]_ ;
  assign \new_[859]_  = \new_[4836]_  & \new_[4827]_ ;
  assign \new_[860]_  = \new_[4820]_  & \new_[4811]_ ;
  assign \new_[861]_  = \new_[4804]_  & \new_[4795]_ ;
  assign \new_[862]_  = \new_[4788]_  & \new_[4779]_ ;
  assign \new_[863]_  = \new_[4772]_  & \new_[4763]_ ;
  assign \new_[864]_  = \new_[4756]_  & \new_[4747]_ ;
  assign \new_[865]_  = \new_[4740]_  & \new_[4731]_ ;
  assign \new_[866]_  = \new_[4724]_  & \new_[4715]_ ;
  assign \new_[867]_  = \new_[4708]_  & \new_[4699]_ ;
  assign \new_[868]_  = \new_[4692]_  & \new_[4683]_ ;
  assign \new_[869]_  = \new_[4676]_  & \new_[4667]_ ;
  assign \new_[870]_  = \new_[4660]_  & \new_[4651]_ ;
  assign \new_[871]_  = \new_[4644]_  & \new_[4635]_ ;
  assign \new_[872]_  = \new_[4628]_  & \new_[4619]_ ;
  assign \new_[873]_  = \new_[4612]_  & \new_[4603]_ ;
  assign \new_[874]_  = \new_[4596]_  & \new_[4587]_ ;
  assign \new_[875]_  = \new_[4580]_  & \new_[4571]_ ;
  assign \new_[876]_  = \new_[4564]_  & \new_[4555]_ ;
  assign \new_[877]_  = \new_[4548]_  & \new_[4539]_ ;
  assign \new_[878]_  = \new_[4532]_  & \new_[4523]_ ;
  assign \new_[879]_  = \new_[4516]_  & \new_[4507]_ ;
  assign \new_[880]_  = \new_[4500]_  & \new_[4491]_ ;
  assign \new_[881]_  = \new_[4484]_  & \new_[4475]_ ;
  assign \new_[882]_  = \new_[4468]_  & \new_[4459]_ ;
  assign \new_[883]_  = \new_[4452]_  & \new_[4443]_ ;
  assign \new_[884]_  = \new_[4436]_  & \new_[4427]_ ;
  assign \new_[885]_  = \new_[4420]_  & \new_[4411]_ ;
  assign \new_[886]_  = \new_[4404]_  & \new_[4395]_ ;
  assign \new_[887]_  = \new_[4388]_  & \new_[4379]_ ;
  assign \new_[888]_  = \new_[4372]_  & \new_[4363]_ ;
  assign \new_[889]_  = \new_[4356]_  & \new_[4347]_ ;
  assign \new_[890]_  = \new_[4340]_  & \new_[4331]_ ;
  assign \new_[891]_  = \new_[4324]_  & \new_[4315]_ ;
  assign \new_[892]_  = \new_[4308]_  & \new_[4299]_ ;
  assign \new_[893]_  = \new_[4292]_  & \new_[4283]_ ;
  assign \new_[894]_  = \new_[4276]_  & \new_[4267]_ ;
  assign \new_[895]_  = \new_[4260]_  & \new_[4251]_ ;
  assign \new_[896]_  = \new_[4244]_  & \new_[4237]_ ;
  assign \new_[897]_  = \new_[4230]_  & \new_[4223]_ ;
  assign \new_[898]_  = \new_[4216]_  & \new_[4209]_ ;
  assign \new_[899]_  = \new_[4202]_  & \new_[4195]_ ;
  assign \new_[900]_  = \new_[4188]_  & \new_[4181]_ ;
  assign \new_[901]_  = \new_[4174]_  & \new_[4167]_ ;
  assign \new_[902]_  = \new_[4160]_  & \new_[4153]_ ;
  assign \new_[903]_  = \new_[4146]_  & \new_[4139]_ ;
  assign \new_[904]_  = \new_[4132]_  & \new_[4125]_ ;
  assign \new_[905]_  = \new_[4118]_  & \new_[4111]_ ;
  assign \new_[906]_  = \new_[4104]_  & \new_[4097]_ ;
  assign \new_[907]_  = \new_[4090]_  & \new_[4083]_ ;
  assign \new_[908]_  = \new_[4076]_  & \new_[4069]_ ;
  assign \new_[909]_  = \new_[4062]_  & \new_[4055]_ ;
  assign \new_[910]_  = \new_[4048]_  & \new_[4041]_ ;
  assign \new_[911]_  = \new_[4034]_  & \new_[4027]_ ;
  assign \new_[912]_  = \new_[4020]_  & \new_[4013]_ ;
  assign \new_[913]_  = \new_[4006]_  & \new_[3999]_ ;
  assign \new_[914]_  = \new_[3992]_  & \new_[3985]_ ;
  assign \new_[915]_  = \new_[3978]_  & \new_[3971]_ ;
  assign \new_[916]_  = \new_[3964]_  & \new_[3957]_ ;
  assign \new_[917]_  = \new_[3950]_  & \new_[3943]_ ;
  assign \new_[918]_  = \new_[3936]_  & \new_[3929]_ ;
  assign \new_[919]_  = \new_[3922]_  & \new_[3915]_ ;
  assign \new_[920]_  = \new_[3908]_  & \new_[3901]_ ;
  assign \new_[921]_  = \new_[3894]_  & \new_[3887]_ ;
  assign \new_[922]_  = \new_[3880]_  & \new_[3873]_ ;
  assign \new_[923]_  = \new_[3866]_  & \new_[3859]_ ;
  assign \new_[924]_  = \new_[3852]_  & \new_[3845]_ ;
  assign \new_[925]_  = \new_[3838]_  & \new_[3831]_ ;
  assign \new_[926]_  = \new_[3824]_  & \new_[3817]_ ;
  assign \new_[927]_  = \new_[3810]_  & \new_[3803]_ ;
  assign \new_[928]_  = \new_[3796]_  & \new_[3789]_ ;
  assign \new_[929]_  = \new_[3782]_  & \new_[3775]_ ;
  assign \new_[930]_  = \new_[3768]_  & \new_[3761]_ ;
  assign \new_[931]_  = \new_[3754]_  & \new_[3747]_ ;
  assign \new_[932]_  = \new_[3740]_  & \new_[3733]_ ;
  assign \new_[933]_  = \new_[3726]_  & \new_[3719]_ ;
  assign \new_[934]_  = \new_[3712]_  & \new_[3705]_ ;
  assign \new_[935]_  = \new_[3698]_  & \new_[3691]_ ;
  assign \new_[936]_  = \new_[3684]_  & \new_[3677]_ ;
  assign \new_[937]_  = \new_[3670]_  & \new_[3663]_ ;
  assign \new_[938]_  = \new_[3656]_  & \new_[3649]_ ;
  assign \new_[939]_  = \new_[3642]_  & \new_[3635]_ ;
  assign \new_[940]_  = \new_[3628]_  & \new_[3621]_ ;
  assign \new_[941]_  = \new_[3614]_  & \new_[3607]_ ;
  assign \new_[942]_  = \new_[3600]_  & \new_[3593]_ ;
  assign \new_[943]_  = \new_[3586]_  & \new_[3579]_ ;
  assign \new_[944]_  = \new_[3572]_  & \new_[3565]_ ;
  assign \new_[945]_  = \new_[3558]_  & \new_[3551]_ ;
  assign \new_[946]_  = \new_[3544]_  & \new_[3537]_ ;
  assign \new_[947]_  = \new_[3532]_  & \new_[3525]_ ;
  assign \new_[948]_  = \new_[3520]_  & \new_[3513]_ ;
  assign \new_[949]_  = \new_[3508]_  & \new_[3501]_ ;
  assign \new_[950]_  = \new_[3496]_  & \new_[3489]_ ;
  assign \new_[951]_  = \new_[3484]_  & \new_[3477]_ ;
  assign \new_[952]_  = \new_[3472]_  & \new_[3465]_ ;
  assign \new_[953]_  = \new_[3460]_  & \new_[3453]_ ;
  assign \new_[954]_  = \new_[3448]_  & \new_[3441]_ ;
  assign \new_[955]_  = \new_[3436]_  & \new_[3429]_ ;
  assign \new_[956]_  = \new_[3424]_  & \new_[3417]_ ;
  assign \new_[957]_  = \new_[3412]_  & \new_[3405]_ ;
  assign \new_[958]_  = \new_[3400]_  & \new_[3393]_ ;
  assign \new_[959]_  = \new_[3388]_  & \new_[3383]_ ;
  assign \new_[960]_  = \new_[3378]_  & \new_[3373]_ ;
  assign \new_[961]_  = \new_[3368]_  & \new_[3363]_ ;
  assign \new_[962]_  = \new_[3358]_  & \new_[3353]_ ;
  assign \new_[963]_  = \new_[3348]_  & \new_[3343]_ ;
  assign \new_[964]_  = \new_[3338]_  & \new_[3333]_ ;
  assign \new_[965]_  = \new_[3328]_  & \new_[3323]_ ;
  assign \new_[966]_  = \new_[3318]_  & \new_[3313]_ ;
  assign \new_[967]_  = \new_[3308]_  & \new_[3303]_ ;
  assign \new_[968]_  = \new_[3298]_  & \new_[3293]_ ;
  assign \new_[969]_  = \new_[3288]_  & \new_[3283]_ ;
  assign \new_[970]_  = \new_[3280]_  & \new_[3275]_ ;
  assign \new_[971]_  = \new_[3272]_  & \new_[3267]_ ;
  assign \new_[972]_  = \new_[3264]_  & \new_[3259]_ ;
  assign \new_[973]_  = \new_[3256]_  & \new_[3251]_ ;
  assign \new_[974]_  = \new_[3248]_  & \new_[3243]_ ;
  assign \new_[975]_  = \new_[3240]_  & \new_[3235]_ ;
  assign \new_[976]_  = \new_[3232]_  & \new_[3227]_ ;
  assign \new_[977]_  = \new_[3224]_  & \new_[3219]_ ;
  assign \new_[978]_  = \new_[3216]_  & \new_[3211]_ ;
  assign \new_[979]_  = \new_[3208]_  & \new_[3203]_ ;
  assign \new_[980]_  = \new_[3200]_  & \new_[3195]_ ;
  assign \new_[981]_  = \new_[3192]_  & \new_[3187]_ ;
  assign \new_[982]_  = \new_[3184]_  & \new_[3179]_ ;
  assign \new_[983]_  = \new_[3176]_  & \new_[3171]_ ;
  assign \new_[984]_  = \new_[3168]_  & \new_[3163]_ ;
  assign \new_[985]_  = \new_[3160]_  & \new_[3157]_ ;
  assign \new_[986]_  = \new_[3154]_  & \new_[3151]_ ;
  assign \new_[987]_  = \new_[3148]_  & \new_[3145]_ ;
  assign \new_[988]_  = \new_[3142]_  & \new_[3139]_ ;
  assign \new_[989]_  = \new_[3136]_  & \new_[3133]_ ;
  assign \new_[990]_  = \new_[3130]_  & \new_[3127]_ ;
  assign \new_[991]_  = \new_[3124]_  & \new_[3121]_ ;
  assign \new_[992]_  = \new_[3118]_  & \new_[3115]_ ;
  assign \new_[993]_  = \new_[3112]_  & \new_[3109]_ ;
  assign \new_[994]_  = \new_[3106]_  & \new_[3103]_ ;
  assign \new_[995]_  = \new_[3100]_  & \new_[3097]_ ;
  assign \new_[996]_  = \new_[3094]_  & \new_[3091]_ ;
  assign \new_[997]_  = \new_[3088]_  & \new_[3085]_ ;
  assign \new_[998]_  = \new_[3082]_  & \new_[3079]_ ;
  assign \new_[999]_  = \new_[3076]_  & \new_[3073]_ ;
  assign \new_[1000]_  = \new_[3070]_  & \new_[3067]_ ;
  assign \new_[1001]_  = A169 & \new_[3064]_ ;
  assign \new_[1002]_  = A169 & \new_[3060]_ ;
  assign \new_[1003]_  = A168 & \new_[3056]_ ;
  assign \new_[1004]_  = A168 & \new_[3052]_ ;
  assign \new_[1005]_  = A200 & \new_[3048]_ ;
  assign \new_[1006]_  = A199 & \new_[3044]_ ;
  assign \new_[1007]_  = A202 & \new_[3040]_ ;
  assign \new_[1008]_  = A202 & \new_[3036]_ ;
  assign \new_[1009]_  = A235 & A169;
  assign \new_[1010]_  = A235 & A202;
  assign \new_[1014]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[1015]_  = \new_[1010]_  | \new_[1014]_ ;
  assign \new_[1018]_  = \new_[1006]_  | \new_[1007]_ ;
  assign \new_[1021]_  = \new_[1004]_  | \new_[1005]_ ;
  assign \new_[1022]_  = \new_[1021]_  | \new_[1018]_ ;
  assign \new_[1023]_  = \new_[1022]_  | \new_[1015]_ ;
  assign \new_[1026]_  = \new_[1002]_  | \new_[1003]_ ;
  assign \new_[1029]_  = \new_[1000]_  | \new_[1001]_ ;
  assign \new_[1030]_  = \new_[1029]_  | \new_[1026]_ ;
  assign \new_[1033]_  = \new_[998]_  | \new_[999]_ ;
  assign \new_[1036]_  = \new_[996]_  | \new_[997]_ ;
  assign \new_[1037]_  = \new_[1036]_  | \new_[1033]_ ;
  assign \new_[1038]_  = \new_[1037]_  | \new_[1030]_ ;
  assign \new_[1039]_  = \new_[1038]_  | \new_[1023]_ ;
  assign \new_[1042]_  = \new_[994]_  | \new_[995]_ ;
  assign \new_[1045]_  = \new_[992]_  | \new_[993]_ ;
  assign \new_[1046]_  = \new_[1045]_  | \new_[1042]_ ;
  assign \new_[1049]_  = \new_[990]_  | \new_[991]_ ;
  assign \new_[1052]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[1053]_  = \new_[1052]_  | \new_[1049]_ ;
  assign \new_[1054]_  = \new_[1053]_  | \new_[1046]_ ;
  assign \new_[1057]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[1060]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[1061]_  = \new_[1060]_  | \new_[1057]_ ;
  assign \new_[1064]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[1067]_  = \new_[980]_  | \new_[981]_ ;
  assign \new_[1068]_  = \new_[1067]_  | \new_[1064]_ ;
  assign \new_[1069]_  = \new_[1068]_  | \new_[1061]_ ;
  assign \new_[1070]_  = \new_[1069]_  | \new_[1054]_ ;
  assign \new_[1071]_  = \new_[1070]_  | \new_[1039]_ ;
  assign \new_[1074]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[1077]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[1078]_  = \new_[1077]_  | \new_[1074]_ ;
  assign \new_[1081]_  = \new_[974]_  | \new_[975]_ ;
  assign \new_[1084]_  = \new_[972]_  | \new_[973]_ ;
  assign \new_[1085]_  = \new_[1084]_  | \new_[1081]_ ;
  assign \new_[1086]_  = \new_[1085]_  | \new_[1078]_ ;
  assign \new_[1089]_  = \new_[970]_  | \new_[971]_ ;
  assign \new_[1092]_  = \new_[968]_  | \new_[969]_ ;
  assign \new_[1093]_  = \new_[1092]_  | \new_[1089]_ ;
  assign \new_[1096]_  = \new_[966]_  | \new_[967]_ ;
  assign \new_[1099]_  = \new_[964]_  | \new_[965]_ ;
  assign \new_[1100]_  = \new_[1099]_  | \new_[1096]_ ;
  assign \new_[1101]_  = \new_[1100]_  | \new_[1093]_ ;
  assign \new_[1102]_  = \new_[1101]_  | \new_[1086]_ ;
  assign \new_[1105]_  = \new_[962]_  | \new_[963]_ ;
  assign \new_[1108]_  = \new_[960]_  | \new_[961]_ ;
  assign \new_[1109]_  = \new_[1108]_  | \new_[1105]_ ;
  assign \new_[1112]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[1115]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[1116]_  = \new_[1115]_  | \new_[1112]_ ;
  assign \new_[1117]_  = \new_[1116]_  | \new_[1109]_ ;
  assign \new_[1120]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[1123]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[1124]_  = \new_[1123]_  | \new_[1120]_ ;
  assign \new_[1127]_  = \new_[950]_  | \new_[951]_ ;
  assign \new_[1130]_  = \new_[948]_  | \new_[949]_ ;
  assign \new_[1131]_  = \new_[1130]_  | \new_[1127]_ ;
  assign \new_[1132]_  = \new_[1131]_  | \new_[1124]_ ;
  assign \new_[1133]_  = \new_[1132]_  | \new_[1117]_ ;
  assign \new_[1134]_  = \new_[1133]_  | \new_[1102]_ ;
  assign \new_[1135]_  = \new_[1134]_  | \new_[1071]_ ;
  assign \new_[1139]_  = \new_[945]_  | \new_[946]_ ;
  assign \new_[1140]_  = \new_[947]_  | \new_[1139]_ ;
  assign \new_[1143]_  = \new_[943]_  | \new_[944]_ ;
  assign \new_[1146]_  = \new_[941]_  | \new_[942]_ ;
  assign \new_[1147]_  = \new_[1146]_  | \new_[1143]_ ;
  assign \new_[1148]_  = \new_[1147]_  | \new_[1140]_ ;
  assign \new_[1151]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[1154]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[1155]_  = \new_[1154]_  | \new_[1151]_ ;
  assign \new_[1158]_  = \new_[935]_  | \new_[936]_ ;
  assign \new_[1161]_  = \new_[933]_  | \new_[934]_ ;
  assign \new_[1162]_  = \new_[1161]_  | \new_[1158]_ ;
  assign \new_[1163]_  = \new_[1162]_  | \new_[1155]_ ;
  assign \new_[1164]_  = \new_[1163]_  | \new_[1148]_ ;
  assign \new_[1167]_  = \new_[931]_  | \new_[932]_ ;
  assign \new_[1170]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[1171]_  = \new_[1170]_  | \new_[1167]_ ;
  assign \new_[1174]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[1177]_  = \new_[925]_  | \new_[926]_ ;
  assign \new_[1178]_  = \new_[1177]_  | \new_[1174]_ ;
  assign \new_[1179]_  = \new_[1178]_  | \new_[1171]_ ;
  assign \new_[1182]_  = \new_[923]_  | \new_[924]_ ;
  assign \new_[1185]_  = \new_[921]_  | \new_[922]_ ;
  assign \new_[1186]_  = \new_[1185]_  | \new_[1182]_ ;
  assign \new_[1189]_  = \new_[919]_  | \new_[920]_ ;
  assign \new_[1192]_  = \new_[917]_  | \new_[918]_ ;
  assign \new_[1193]_  = \new_[1192]_  | \new_[1189]_ ;
  assign \new_[1194]_  = \new_[1193]_  | \new_[1186]_ ;
  assign \new_[1195]_  = \new_[1194]_  | \new_[1179]_ ;
  assign \new_[1196]_  = \new_[1195]_  | \new_[1164]_ ;
  assign \new_[1199]_  = \new_[915]_  | \new_[916]_ ;
  assign \new_[1202]_  = \new_[913]_  | \new_[914]_ ;
  assign \new_[1203]_  = \new_[1202]_  | \new_[1199]_ ;
  assign \new_[1206]_  = \new_[911]_  | \new_[912]_ ;
  assign \new_[1209]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[1210]_  = \new_[1209]_  | \new_[1206]_ ;
  assign \new_[1211]_  = \new_[1210]_  | \new_[1203]_ ;
  assign \new_[1214]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[1217]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[1218]_  = \new_[1217]_  | \new_[1214]_ ;
  assign \new_[1221]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[1224]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[1225]_  = \new_[1224]_  | \new_[1221]_ ;
  assign \new_[1226]_  = \new_[1225]_  | \new_[1218]_ ;
  assign \new_[1227]_  = \new_[1226]_  | \new_[1211]_ ;
  assign \new_[1230]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[1233]_  = \new_[897]_  | \new_[898]_ ;
  assign \new_[1234]_  = \new_[1233]_  | \new_[1230]_ ;
  assign \new_[1237]_  = \new_[895]_  | \new_[896]_ ;
  assign \new_[1240]_  = \new_[893]_  | \new_[894]_ ;
  assign \new_[1241]_  = \new_[1240]_  | \new_[1237]_ ;
  assign \new_[1242]_  = \new_[1241]_  | \new_[1234]_ ;
  assign \new_[1245]_  = \new_[891]_  | \new_[892]_ ;
  assign \new_[1248]_  = \new_[889]_  | \new_[890]_ ;
  assign \new_[1249]_  = \new_[1248]_  | \new_[1245]_ ;
  assign \new_[1252]_  = \new_[887]_  | \new_[888]_ ;
  assign \new_[1255]_  = \new_[885]_  | \new_[886]_ ;
  assign \new_[1256]_  = \new_[1255]_  | \new_[1252]_ ;
  assign \new_[1257]_  = \new_[1256]_  | \new_[1249]_ ;
  assign \new_[1258]_  = \new_[1257]_  | \new_[1242]_ ;
  assign \new_[1259]_  = \new_[1258]_  | \new_[1227]_ ;
  assign \new_[1260]_  = \new_[1259]_  | \new_[1196]_ ;
  assign \new_[1261]_  = \new_[1260]_  | \new_[1135]_ ;
  assign \new_[1265]_  = \new_[882]_  | \new_[883]_ ;
  assign \new_[1266]_  = \new_[884]_  | \new_[1265]_ ;
  assign \new_[1269]_  = \new_[880]_  | \new_[881]_ ;
  assign \new_[1272]_  = \new_[878]_  | \new_[879]_ ;
  assign \new_[1273]_  = \new_[1272]_  | \new_[1269]_ ;
  assign \new_[1274]_  = \new_[1273]_  | \new_[1266]_ ;
  assign \new_[1277]_  = \new_[876]_  | \new_[877]_ ;
  assign \new_[1280]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[1281]_  = \new_[1280]_  | \new_[1277]_ ;
  assign \new_[1284]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[1287]_  = \new_[870]_  | \new_[871]_ ;
  assign \new_[1288]_  = \new_[1287]_  | \new_[1284]_ ;
  assign \new_[1289]_  = \new_[1288]_  | \new_[1281]_ ;
  assign \new_[1290]_  = \new_[1289]_  | \new_[1274]_ ;
  assign \new_[1293]_  = \new_[868]_  | \new_[869]_ ;
  assign \new_[1296]_  = \new_[866]_  | \new_[867]_ ;
  assign \new_[1297]_  = \new_[1296]_  | \new_[1293]_ ;
  assign \new_[1300]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[1303]_  = \new_[862]_  | \new_[863]_ ;
  assign \new_[1304]_  = \new_[1303]_  | \new_[1300]_ ;
  assign \new_[1305]_  = \new_[1304]_  | \new_[1297]_ ;
  assign \new_[1308]_  = \new_[860]_  | \new_[861]_ ;
  assign \new_[1311]_  = \new_[858]_  | \new_[859]_ ;
  assign \new_[1312]_  = \new_[1311]_  | \new_[1308]_ ;
  assign \new_[1315]_  = \new_[856]_  | \new_[857]_ ;
  assign \new_[1318]_  = \new_[854]_  | \new_[855]_ ;
  assign \new_[1319]_  = \new_[1318]_  | \new_[1315]_ ;
  assign \new_[1320]_  = \new_[1319]_  | \new_[1312]_ ;
  assign \new_[1321]_  = \new_[1320]_  | \new_[1305]_ ;
  assign \new_[1322]_  = \new_[1321]_  | \new_[1290]_ ;
  assign \new_[1325]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[1328]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[1329]_  = \new_[1328]_  | \new_[1325]_ ;
  assign \new_[1332]_  = \new_[848]_  | \new_[849]_ ;
  assign \new_[1335]_  = \new_[846]_  | \new_[847]_ ;
  assign \new_[1336]_  = \new_[1335]_  | \new_[1332]_ ;
  assign \new_[1337]_  = \new_[1336]_  | \new_[1329]_ ;
  assign \new_[1340]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[1343]_  = \new_[842]_  | \new_[843]_ ;
  assign \new_[1344]_  = \new_[1343]_  | \new_[1340]_ ;
  assign \new_[1347]_  = \new_[840]_  | \new_[841]_ ;
  assign \new_[1350]_  = \new_[838]_  | \new_[839]_ ;
  assign \new_[1351]_  = \new_[1350]_  | \new_[1347]_ ;
  assign \new_[1352]_  = \new_[1351]_  | \new_[1344]_ ;
  assign \new_[1353]_  = \new_[1352]_  | \new_[1337]_ ;
  assign \new_[1356]_  = \new_[836]_  | \new_[837]_ ;
  assign \new_[1359]_  = \new_[834]_  | \new_[835]_ ;
  assign \new_[1360]_  = \new_[1359]_  | \new_[1356]_ ;
  assign \new_[1363]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[1366]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[1367]_  = \new_[1366]_  | \new_[1363]_ ;
  assign \new_[1368]_  = \new_[1367]_  | \new_[1360]_ ;
  assign \new_[1371]_  = \new_[828]_  | \new_[829]_ ;
  assign \new_[1374]_  = \new_[826]_  | \new_[827]_ ;
  assign \new_[1375]_  = \new_[1374]_  | \new_[1371]_ ;
  assign \new_[1378]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[1381]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[1382]_  = \new_[1381]_  | \new_[1378]_ ;
  assign \new_[1383]_  = \new_[1382]_  | \new_[1375]_ ;
  assign \new_[1384]_  = \new_[1383]_  | \new_[1368]_ ;
  assign \new_[1385]_  = \new_[1384]_  | \new_[1353]_ ;
  assign \new_[1386]_  = \new_[1385]_  | \new_[1322]_ ;
  assign \new_[1390]_  = \new_[819]_  | \new_[820]_ ;
  assign \new_[1391]_  = \new_[821]_  | \new_[1390]_ ;
  assign \new_[1394]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[1397]_  = \new_[815]_  | \new_[816]_ ;
  assign \new_[1398]_  = \new_[1397]_  | \new_[1394]_ ;
  assign \new_[1399]_  = \new_[1398]_  | \new_[1391]_ ;
  assign \new_[1402]_  = \new_[813]_  | \new_[814]_ ;
  assign \new_[1405]_  = \new_[811]_  | \new_[812]_ ;
  assign \new_[1406]_  = \new_[1405]_  | \new_[1402]_ ;
  assign \new_[1409]_  = \new_[809]_  | \new_[810]_ ;
  assign \new_[1412]_  = \new_[807]_  | \new_[808]_ ;
  assign \new_[1413]_  = \new_[1412]_  | \new_[1409]_ ;
  assign \new_[1414]_  = \new_[1413]_  | \new_[1406]_ ;
  assign \new_[1415]_  = \new_[1414]_  | \new_[1399]_ ;
  assign \new_[1418]_  = \new_[805]_  | \new_[806]_ ;
  assign \new_[1421]_  = \new_[803]_  | \new_[804]_ ;
  assign \new_[1422]_  = \new_[1421]_  | \new_[1418]_ ;
  assign \new_[1425]_  = \new_[801]_  | \new_[802]_ ;
  assign \new_[1428]_  = \new_[799]_  | \new_[800]_ ;
  assign \new_[1429]_  = \new_[1428]_  | \new_[1425]_ ;
  assign \new_[1430]_  = \new_[1429]_  | \new_[1422]_ ;
  assign \new_[1433]_  = \new_[797]_  | \new_[798]_ ;
  assign \new_[1436]_  = \new_[795]_  | \new_[796]_ ;
  assign \new_[1437]_  = \new_[1436]_  | \new_[1433]_ ;
  assign \new_[1440]_  = \new_[793]_  | \new_[794]_ ;
  assign \new_[1443]_  = \new_[791]_  | \new_[792]_ ;
  assign \new_[1444]_  = \new_[1443]_  | \new_[1440]_ ;
  assign \new_[1445]_  = \new_[1444]_  | \new_[1437]_ ;
  assign \new_[1446]_  = \new_[1445]_  | \new_[1430]_ ;
  assign \new_[1447]_  = \new_[1446]_  | \new_[1415]_ ;
  assign \new_[1450]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[1453]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[1454]_  = \new_[1453]_  | \new_[1450]_ ;
  assign \new_[1457]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[1460]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[1461]_  = \new_[1460]_  | \new_[1457]_ ;
  assign \new_[1462]_  = \new_[1461]_  | \new_[1454]_ ;
  assign \new_[1465]_  = \new_[781]_  | \new_[782]_ ;
  assign \new_[1468]_  = \new_[779]_  | \new_[780]_ ;
  assign \new_[1469]_  = \new_[1468]_  | \new_[1465]_ ;
  assign \new_[1472]_  = \new_[777]_  | \new_[778]_ ;
  assign \new_[1475]_  = \new_[775]_  | \new_[776]_ ;
  assign \new_[1476]_  = \new_[1475]_  | \new_[1472]_ ;
  assign \new_[1477]_  = \new_[1476]_  | \new_[1469]_ ;
  assign \new_[1478]_  = \new_[1477]_  | \new_[1462]_ ;
  assign \new_[1481]_  = \new_[773]_  | \new_[774]_ ;
  assign \new_[1484]_  = \new_[771]_  | \new_[772]_ ;
  assign \new_[1485]_  = \new_[1484]_  | \new_[1481]_ ;
  assign \new_[1488]_  = \new_[769]_  | \new_[770]_ ;
  assign \new_[1491]_  = \new_[767]_  | \new_[768]_ ;
  assign \new_[1492]_  = \new_[1491]_  | \new_[1488]_ ;
  assign \new_[1493]_  = \new_[1492]_  | \new_[1485]_ ;
  assign \new_[1496]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[1499]_  = \new_[763]_  | \new_[764]_ ;
  assign \new_[1500]_  = \new_[1499]_  | \new_[1496]_ ;
  assign \new_[1503]_  = \new_[761]_  | \new_[762]_ ;
  assign \new_[1506]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[1507]_  = \new_[1506]_  | \new_[1503]_ ;
  assign \new_[1508]_  = \new_[1507]_  | \new_[1500]_ ;
  assign \new_[1509]_  = \new_[1508]_  | \new_[1493]_ ;
  assign \new_[1510]_  = \new_[1509]_  | \new_[1478]_ ;
  assign \new_[1511]_  = \new_[1510]_  | \new_[1447]_ ;
  assign \new_[1512]_  = \new_[1511]_  | \new_[1386]_ ;
  assign \new_[1513]_  = \new_[1512]_  | \new_[1261]_ ;
  assign \new_[1517]_  = \new_[756]_  | \new_[757]_ ;
  assign \new_[1518]_  = \new_[758]_  | \new_[1517]_ ;
  assign \new_[1521]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[1524]_  = \new_[752]_  | \new_[753]_ ;
  assign \new_[1525]_  = \new_[1524]_  | \new_[1521]_ ;
  assign \new_[1526]_  = \new_[1525]_  | \new_[1518]_ ;
  assign \new_[1529]_  = \new_[750]_  | \new_[751]_ ;
  assign \new_[1532]_  = \new_[748]_  | \new_[749]_ ;
  assign \new_[1533]_  = \new_[1532]_  | \new_[1529]_ ;
  assign \new_[1536]_  = \new_[746]_  | \new_[747]_ ;
  assign \new_[1539]_  = \new_[744]_  | \new_[745]_ ;
  assign \new_[1540]_  = \new_[1539]_  | \new_[1536]_ ;
  assign \new_[1541]_  = \new_[1540]_  | \new_[1533]_ ;
  assign \new_[1542]_  = \new_[1541]_  | \new_[1526]_ ;
  assign \new_[1545]_  = \new_[742]_  | \new_[743]_ ;
  assign \new_[1548]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[1549]_  = \new_[1548]_  | \new_[1545]_ ;
  assign \new_[1552]_  = \new_[738]_  | \new_[739]_ ;
  assign \new_[1555]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[1556]_  = \new_[1555]_  | \new_[1552]_ ;
  assign \new_[1557]_  = \new_[1556]_  | \new_[1549]_ ;
  assign \new_[1560]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[1563]_  = \new_[732]_  | \new_[733]_ ;
  assign \new_[1564]_  = \new_[1563]_  | \new_[1560]_ ;
  assign \new_[1567]_  = \new_[730]_  | \new_[731]_ ;
  assign \new_[1570]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[1571]_  = \new_[1570]_  | \new_[1567]_ ;
  assign \new_[1572]_  = \new_[1571]_  | \new_[1564]_ ;
  assign \new_[1573]_  = \new_[1572]_  | \new_[1557]_ ;
  assign \new_[1574]_  = \new_[1573]_  | \new_[1542]_ ;
  assign \new_[1577]_  = \new_[726]_  | \new_[727]_ ;
  assign \new_[1580]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[1581]_  = \new_[1580]_  | \new_[1577]_ ;
  assign \new_[1584]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[1587]_  = \new_[720]_  | \new_[721]_ ;
  assign \new_[1588]_  = \new_[1587]_  | \new_[1584]_ ;
  assign \new_[1589]_  = \new_[1588]_  | \new_[1581]_ ;
  assign \new_[1592]_  = \new_[718]_  | \new_[719]_ ;
  assign \new_[1595]_  = \new_[716]_  | \new_[717]_ ;
  assign \new_[1596]_  = \new_[1595]_  | \new_[1592]_ ;
  assign \new_[1599]_  = \new_[714]_  | \new_[715]_ ;
  assign \new_[1602]_  = \new_[712]_  | \new_[713]_ ;
  assign \new_[1603]_  = \new_[1602]_  | \new_[1599]_ ;
  assign \new_[1604]_  = \new_[1603]_  | \new_[1596]_ ;
  assign \new_[1605]_  = \new_[1604]_  | \new_[1589]_ ;
  assign \new_[1608]_  = \new_[710]_  | \new_[711]_ ;
  assign \new_[1611]_  = \new_[708]_  | \new_[709]_ ;
  assign \new_[1612]_  = \new_[1611]_  | \new_[1608]_ ;
  assign \new_[1615]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[1618]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[1619]_  = \new_[1618]_  | \new_[1615]_ ;
  assign \new_[1620]_  = \new_[1619]_  | \new_[1612]_ ;
  assign \new_[1623]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[1626]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[1627]_  = \new_[1626]_  | \new_[1623]_ ;
  assign \new_[1630]_  = \new_[698]_  | \new_[699]_ ;
  assign \new_[1633]_  = \new_[696]_  | \new_[697]_ ;
  assign \new_[1634]_  = \new_[1633]_  | \new_[1630]_ ;
  assign \new_[1635]_  = \new_[1634]_  | \new_[1627]_ ;
  assign \new_[1636]_  = \new_[1635]_  | \new_[1620]_ ;
  assign \new_[1637]_  = \new_[1636]_  | \new_[1605]_ ;
  assign \new_[1638]_  = \new_[1637]_  | \new_[1574]_ ;
  assign \new_[1642]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[1643]_  = \new_[695]_  | \new_[1642]_ ;
  assign \new_[1646]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[1649]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[1650]_  = \new_[1649]_  | \new_[1646]_ ;
  assign \new_[1651]_  = \new_[1650]_  | \new_[1643]_ ;
  assign \new_[1654]_  = \new_[687]_  | \new_[688]_ ;
  assign \new_[1657]_  = \new_[685]_  | \new_[686]_ ;
  assign \new_[1658]_  = \new_[1657]_  | \new_[1654]_ ;
  assign \new_[1661]_  = \new_[683]_  | \new_[684]_ ;
  assign \new_[1664]_  = \new_[681]_  | \new_[682]_ ;
  assign \new_[1665]_  = \new_[1664]_  | \new_[1661]_ ;
  assign \new_[1666]_  = \new_[1665]_  | \new_[1658]_ ;
  assign \new_[1667]_  = \new_[1666]_  | \new_[1651]_ ;
  assign \new_[1670]_  = \new_[679]_  | \new_[680]_ ;
  assign \new_[1673]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[1674]_  = \new_[1673]_  | \new_[1670]_ ;
  assign \new_[1677]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[1680]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[1681]_  = \new_[1680]_  | \new_[1677]_ ;
  assign \new_[1682]_  = \new_[1681]_  | \new_[1674]_ ;
  assign \new_[1685]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[1688]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[1689]_  = \new_[1688]_  | \new_[1685]_ ;
  assign \new_[1692]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[1695]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[1696]_  = \new_[1695]_  | \new_[1692]_ ;
  assign \new_[1697]_  = \new_[1696]_  | \new_[1689]_ ;
  assign \new_[1698]_  = \new_[1697]_  | \new_[1682]_ ;
  assign \new_[1699]_  = \new_[1698]_  | \new_[1667]_ ;
  assign \new_[1702]_  = \new_[663]_  | \new_[664]_ ;
  assign \new_[1705]_  = \new_[661]_  | \new_[662]_ ;
  assign \new_[1706]_  = \new_[1705]_  | \new_[1702]_ ;
  assign \new_[1709]_  = \new_[659]_  | \new_[660]_ ;
  assign \new_[1712]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[1713]_  = \new_[1712]_  | \new_[1709]_ ;
  assign \new_[1714]_  = \new_[1713]_  | \new_[1706]_ ;
  assign \new_[1717]_  = \new_[655]_  | \new_[656]_ ;
  assign \new_[1720]_  = \new_[653]_  | \new_[654]_ ;
  assign \new_[1721]_  = \new_[1720]_  | \new_[1717]_ ;
  assign \new_[1724]_  = \new_[651]_  | \new_[652]_ ;
  assign \new_[1727]_  = \new_[649]_  | \new_[650]_ ;
  assign \new_[1728]_  = \new_[1727]_  | \new_[1724]_ ;
  assign \new_[1729]_  = \new_[1728]_  | \new_[1721]_ ;
  assign \new_[1730]_  = \new_[1729]_  | \new_[1714]_ ;
  assign \new_[1733]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[1736]_  = \new_[645]_  | \new_[646]_ ;
  assign \new_[1737]_  = \new_[1736]_  | \new_[1733]_ ;
  assign \new_[1740]_  = \new_[643]_  | \new_[644]_ ;
  assign \new_[1743]_  = \new_[641]_  | \new_[642]_ ;
  assign \new_[1744]_  = \new_[1743]_  | \new_[1740]_ ;
  assign \new_[1745]_  = \new_[1744]_  | \new_[1737]_ ;
  assign \new_[1748]_  = \new_[639]_  | \new_[640]_ ;
  assign \new_[1751]_  = \new_[637]_  | \new_[638]_ ;
  assign \new_[1752]_  = \new_[1751]_  | \new_[1748]_ ;
  assign \new_[1755]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[1758]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[1759]_  = \new_[1758]_  | \new_[1755]_ ;
  assign \new_[1760]_  = \new_[1759]_  | \new_[1752]_ ;
  assign \new_[1761]_  = \new_[1760]_  | \new_[1745]_ ;
  assign \new_[1762]_  = \new_[1761]_  | \new_[1730]_ ;
  assign \new_[1763]_  = \new_[1762]_  | \new_[1699]_ ;
  assign \new_[1764]_  = \new_[1763]_  | \new_[1638]_ ;
  assign \new_[1768]_  = \new_[630]_  | \new_[631]_ ;
  assign \new_[1769]_  = \new_[632]_  | \new_[1768]_ ;
  assign \new_[1772]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[1775]_  = \new_[626]_  | \new_[627]_ ;
  assign \new_[1776]_  = \new_[1775]_  | \new_[1772]_ ;
  assign \new_[1777]_  = \new_[1776]_  | \new_[1769]_ ;
  assign \new_[1780]_  = \new_[624]_  | \new_[625]_ ;
  assign \new_[1783]_  = \new_[622]_  | \new_[623]_ ;
  assign \new_[1784]_  = \new_[1783]_  | \new_[1780]_ ;
  assign \new_[1787]_  = \new_[620]_  | \new_[621]_ ;
  assign \new_[1790]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[1791]_  = \new_[1790]_  | \new_[1787]_ ;
  assign \new_[1792]_  = \new_[1791]_  | \new_[1784]_ ;
  assign \new_[1793]_  = \new_[1792]_  | \new_[1777]_ ;
  assign \new_[1796]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[1799]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[1800]_  = \new_[1799]_  | \new_[1796]_ ;
  assign \new_[1803]_  = \new_[612]_  | \new_[613]_ ;
  assign \new_[1806]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[1807]_  = \new_[1806]_  | \new_[1803]_ ;
  assign \new_[1808]_  = \new_[1807]_  | \new_[1800]_ ;
  assign \new_[1811]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[1814]_  = \new_[606]_  | \new_[607]_ ;
  assign \new_[1815]_  = \new_[1814]_  | \new_[1811]_ ;
  assign \new_[1818]_  = \new_[604]_  | \new_[605]_ ;
  assign \new_[1821]_  = \new_[602]_  | \new_[603]_ ;
  assign \new_[1822]_  = \new_[1821]_  | \new_[1818]_ ;
  assign \new_[1823]_  = \new_[1822]_  | \new_[1815]_ ;
  assign \new_[1824]_  = \new_[1823]_  | \new_[1808]_ ;
  assign \new_[1825]_  = \new_[1824]_  | \new_[1793]_ ;
  assign \new_[1828]_  = \new_[600]_  | \new_[601]_ ;
  assign \new_[1831]_  = \new_[598]_  | \new_[599]_ ;
  assign \new_[1832]_  = \new_[1831]_  | \new_[1828]_ ;
  assign \new_[1835]_  = \new_[596]_  | \new_[597]_ ;
  assign \new_[1838]_  = \new_[594]_  | \new_[595]_ ;
  assign \new_[1839]_  = \new_[1838]_  | \new_[1835]_ ;
  assign \new_[1840]_  = \new_[1839]_  | \new_[1832]_ ;
  assign \new_[1843]_  = \new_[592]_  | \new_[593]_ ;
  assign \new_[1846]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[1847]_  = \new_[1846]_  | \new_[1843]_ ;
  assign \new_[1850]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[1853]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[1854]_  = \new_[1853]_  | \new_[1850]_ ;
  assign \new_[1855]_  = \new_[1854]_  | \new_[1847]_ ;
  assign \new_[1856]_  = \new_[1855]_  | \new_[1840]_ ;
  assign \new_[1859]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[1862]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[1863]_  = \new_[1862]_  | \new_[1859]_ ;
  assign \new_[1866]_  = \new_[580]_  | \new_[581]_ ;
  assign \new_[1869]_  = \new_[578]_  | \new_[579]_ ;
  assign \new_[1870]_  = \new_[1869]_  | \new_[1866]_ ;
  assign \new_[1871]_  = \new_[1870]_  | \new_[1863]_ ;
  assign \new_[1874]_  = \new_[576]_  | \new_[577]_ ;
  assign \new_[1877]_  = \new_[574]_  | \new_[575]_ ;
  assign \new_[1878]_  = \new_[1877]_  | \new_[1874]_ ;
  assign \new_[1881]_  = \new_[572]_  | \new_[573]_ ;
  assign \new_[1884]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[1885]_  = \new_[1884]_  | \new_[1881]_ ;
  assign \new_[1886]_  = \new_[1885]_  | \new_[1878]_ ;
  assign \new_[1887]_  = \new_[1886]_  | \new_[1871]_ ;
  assign \new_[1888]_  = \new_[1887]_  | \new_[1856]_ ;
  assign \new_[1889]_  = \new_[1888]_  | \new_[1825]_ ;
  assign \new_[1892]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[1895]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[1896]_  = \new_[1895]_  | \new_[1892]_ ;
  assign \new_[1899]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[1902]_  = \new_[562]_  | \new_[563]_ ;
  assign \new_[1903]_  = \new_[1902]_  | \new_[1899]_ ;
  assign \new_[1904]_  = \new_[1903]_  | \new_[1896]_ ;
  assign \new_[1907]_  = \new_[560]_  | \new_[561]_ ;
  assign \new_[1910]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[1911]_  = \new_[1910]_  | \new_[1907]_ ;
  assign \new_[1914]_  = \new_[556]_  | \new_[557]_ ;
  assign \new_[1917]_  = \new_[554]_  | \new_[555]_ ;
  assign \new_[1918]_  = \new_[1917]_  | \new_[1914]_ ;
  assign \new_[1919]_  = \new_[1918]_  | \new_[1911]_ ;
  assign \new_[1920]_  = \new_[1919]_  | \new_[1904]_ ;
  assign \new_[1923]_  = \new_[552]_  | \new_[553]_ ;
  assign \new_[1926]_  = \new_[550]_  | \new_[551]_ ;
  assign \new_[1927]_  = \new_[1926]_  | \new_[1923]_ ;
  assign \new_[1930]_  = \new_[548]_  | \new_[549]_ ;
  assign \new_[1933]_  = \new_[546]_  | \new_[547]_ ;
  assign \new_[1934]_  = \new_[1933]_  | \new_[1930]_ ;
  assign \new_[1935]_  = \new_[1934]_  | \new_[1927]_ ;
  assign \new_[1938]_  = \new_[544]_  | \new_[545]_ ;
  assign \new_[1941]_  = \new_[542]_  | \new_[543]_ ;
  assign \new_[1942]_  = \new_[1941]_  | \new_[1938]_ ;
  assign \new_[1945]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[1948]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[1949]_  = \new_[1948]_  | \new_[1945]_ ;
  assign \new_[1950]_  = \new_[1949]_  | \new_[1942]_ ;
  assign \new_[1951]_  = \new_[1950]_  | \new_[1935]_ ;
  assign \new_[1952]_  = \new_[1951]_  | \new_[1920]_ ;
  assign \new_[1955]_  = \new_[536]_  | \new_[537]_ ;
  assign \new_[1958]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[1959]_  = \new_[1958]_  | \new_[1955]_ ;
  assign \new_[1962]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[1965]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[1966]_  = \new_[1965]_  | \new_[1962]_ ;
  assign \new_[1967]_  = \new_[1966]_  | \new_[1959]_ ;
  assign \new_[1970]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[1973]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[1974]_  = \new_[1973]_  | \new_[1970]_ ;
  assign \new_[1977]_  = \new_[524]_  | \new_[525]_ ;
  assign \new_[1980]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[1981]_  = \new_[1980]_  | \new_[1977]_ ;
  assign \new_[1982]_  = \new_[1981]_  | \new_[1974]_ ;
  assign \new_[1983]_  = \new_[1982]_  | \new_[1967]_ ;
  assign \new_[1986]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[1989]_  = \new_[518]_  | \new_[519]_ ;
  assign \new_[1990]_  = \new_[1989]_  | \new_[1986]_ ;
  assign \new_[1993]_  = \new_[516]_  | \new_[517]_ ;
  assign \new_[1996]_  = \new_[514]_  | \new_[515]_ ;
  assign \new_[1997]_  = \new_[1996]_  | \new_[1993]_ ;
  assign \new_[1998]_  = \new_[1997]_  | \new_[1990]_ ;
  assign \new_[2001]_  = \new_[512]_  | \new_[513]_ ;
  assign \new_[2004]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[2005]_  = \new_[2004]_  | \new_[2001]_ ;
  assign \new_[2008]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[2011]_  = \new_[506]_  | \new_[507]_ ;
  assign \new_[2012]_  = \new_[2011]_  | \new_[2008]_ ;
  assign \new_[2013]_  = \new_[2012]_  | \new_[2005]_ ;
  assign \new_[2014]_  = \new_[2013]_  | \new_[1998]_ ;
  assign \new_[2015]_  = \new_[2014]_  | \new_[1983]_ ;
  assign \new_[2016]_  = \new_[2015]_  | \new_[1952]_ ;
  assign \new_[2017]_  = \new_[2016]_  | \new_[1889]_ ;
  assign \new_[2018]_  = \new_[2017]_  | \new_[1764]_ ;
  assign \new_[2019]_  = \new_[2018]_  | \new_[1513]_ ;
  assign \new_[2023]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[2024]_  = \new_[505]_  | \new_[2023]_ ;
  assign \new_[2027]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[2030]_  = \new_[499]_  | \new_[500]_ ;
  assign \new_[2031]_  = \new_[2030]_  | \new_[2027]_ ;
  assign \new_[2032]_  = \new_[2031]_  | \new_[2024]_ ;
  assign \new_[2035]_  = \new_[497]_  | \new_[498]_ ;
  assign \new_[2038]_  = \new_[495]_  | \new_[496]_ ;
  assign \new_[2039]_  = \new_[2038]_  | \new_[2035]_ ;
  assign \new_[2042]_  = \new_[493]_  | \new_[494]_ ;
  assign \new_[2045]_  = \new_[491]_  | \new_[492]_ ;
  assign \new_[2046]_  = \new_[2045]_  | \new_[2042]_ ;
  assign \new_[2047]_  = \new_[2046]_  | \new_[2039]_ ;
  assign \new_[2048]_  = \new_[2047]_  | \new_[2032]_ ;
  assign \new_[2051]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[2054]_  = \new_[487]_  | \new_[488]_ ;
  assign \new_[2055]_  = \new_[2054]_  | \new_[2051]_ ;
  assign \new_[2058]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[2061]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[2062]_  = \new_[2061]_  | \new_[2058]_ ;
  assign \new_[2063]_  = \new_[2062]_  | \new_[2055]_ ;
  assign \new_[2066]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[2069]_  = \new_[479]_  | \new_[480]_ ;
  assign \new_[2070]_  = \new_[2069]_  | \new_[2066]_ ;
  assign \new_[2073]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[2076]_  = \new_[475]_  | \new_[476]_ ;
  assign \new_[2077]_  = \new_[2076]_  | \new_[2073]_ ;
  assign \new_[2078]_  = \new_[2077]_  | \new_[2070]_ ;
  assign \new_[2079]_  = \new_[2078]_  | \new_[2063]_ ;
  assign \new_[2080]_  = \new_[2079]_  | \new_[2048]_ ;
  assign \new_[2083]_  = \new_[473]_  | \new_[474]_ ;
  assign \new_[2086]_  = \new_[471]_  | \new_[472]_ ;
  assign \new_[2087]_  = \new_[2086]_  | \new_[2083]_ ;
  assign \new_[2090]_  = \new_[469]_  | \new_[470]_ ;
  assign \new_[2093]_  = \new_[467]_  | \new_[468]_ ;
  assign \new_[2094]_  = \new_[2093]_  | \new_[2090]_ ;
  assign \new_[2095]_  = \new_[2094]_  | \new_[2087]_ ;
  assign \new_[2098]_  = \new_[465]_  | \new_[466]_ ;
  assign \new_[2101]_  = \new_[463]_  | \new_[464]_ ;
  assign \new_[2102]_  = \new_[2101]_  | \new_[2098]_ ;
  assign \new_[2105]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[2108]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[2109]_  = \new_[2108]_  | \new_[2105]_ ;
  assign \new_[2110]_  = \new_[2109]_  | \new_[2102]_ ;
  assign \new_[2111]_  = \new_[2110]_  | \new_[2095]_ ;
  assign \new_[2114]_  = \new_[457]_  | \new_[458]_ ;
  assign \new_[2117]_  = \new_[455]_  | \new_[456]_ ;
  assign \new_[2118]_  = \new_[2117]_  | \new_[2114]_ ;
  assign \new_[2121]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[2124]_  = \new_[451]_  | \new_[452]_ ;
  assign \new_[2125]_  = \new_[2124]_  | \new_[2121]_ ;
  assign \new_[2126]_  = \new_[2125]_  | \new_[2118]_ ;
  assign \new_[2129]_  = \new_[449]_  | \new_[450]_ ;
  assign \new_[2132]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[2133]_  = \new_[2132]_  | \new_[2129]_ ;
  assign \new_[2136]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[2139]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[2140]_  = \new_[2139]_  | \new_[2136]_ ;
  assign \new_[2141]_  = \new_[2140]_  | \new_[2133]_ ;
  assign \new_[2142]_  = \new_[2141]_  | \new_[2126]_ ;
  assign \new_[2143]_  = \new_[2142]_  | \new_[2111]_ ;
  assign \new_[2144]_  = \new_[2143]_  | \new_[2080]_ ;
  assign \new_[2148]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[2149]_  = \new_[442]_  | \new_[2148]_ ;
  assign \new_[2152]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[2155]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[2156]_  = \new_[2155]_  | \new_[2152]_ ;
  assign \new_[2157]_  = \new_[2156]_  | \new_[2149]_ ;
  assign \new_[2160]_  = \new_[434]_  | \new_[435]_ ;
  assign \new_[2163]_  = \new_[432]_  | \new_[433]_ ;
  assign \new_[2164]_  = \new_[2163]_  | \new_[2160]_ ;
  assign \new_[2167]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[2170]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[2171]_  = \new_[2170]_  | \new_[2167]_ ;
  assign \new_[2172]_  = \new_[2171]_  | \new_[2164]_ ;
  assign \new_[2173]_  = \new_[2172]_  | \new_[2157]_ ;
  assign \new_[2176]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[2179]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[2180]_  = \new_[2179]_  | \new_[2176]_ ;
  assign \new_[2183]_  = \new_[422]_  | \new_[423]_ ;
  assign \new_[2186]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[2187]_  = \new_[2186]_  | \new_[2183]_ ;
  assign \new_[2188]_  = \new_[2187]_  | \new_[2180]_ ;
  assign \new_[2191]_  = \new_[418]_  | \new_[419]_ ;
  assign \new_[2194]_  = \new_[416]_  | \new_[417]_ ;
  assign \new_[2195]_  = \new_[2194]_  | \new_[2191]_ ;
  assign \new_[2198]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[2201]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[2202]_  = \new_[2201]_  | \new_[2198]_ ;
  assign \new_[2203]_  = \new_[2202]_  | \new_[2195]_ ;
  assign \new_[2204]_  = \new_[2203]_  | \new_[2188]_ ;
  assign \new_[2205]_  = \new_[2204]_  | \new_[2173]_ ;
  assign \new_[2208]_  = \new_[410]_  | \new_[411]_ ;
  assign \new_[2211]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[2212]_  = \new_[2211]_  | \new_[2208]_ ;
  assign \new_[2215]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[2218]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[2219]_  = \new_[2218]_  | \new_[2215]_ ;
  assign \new_[2220]_  = \new_[2219]_  | \new_[2212]_ ;
  assign \new_[2223]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[2226]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[2227]_  = \new_[2226]_  | \new_[2223]_ ;
  assign \new_[2230]_  = \new_[398]_  | \new_[399]_ ;
  assign \new_[2233]_  = \new_[396]_  | \new_[397]_ ;
  assign \new_[2234]_  = \new_[2233]_  | \new_[2230]_ ;
  assign \new_[2235]_  = \new_[2234]_  | \new_[2227]_ ;
  assign \new_[2236]_  = \new_[2235]_  | \new_[2220]_ ;
  assign \new_[2239]_  = \new_[394]_  | \new_[395]_ ;
  assign \new_[2242]_  = \new_[392]_  | \new_[393]_ ;
  assign \new_[2243]_  = \new_[2242]_  | \new_[2239]_ ;
  assign \new_[2246]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[2249]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[2250]_  = \new_[2249]_  | \new_[2246]_ ;
  assign \new_[2251]_  = \new_[2250]_  | \new_[2243]_ ;
  assign \new_[2254]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[2257]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[2258]_  = \new_[2257]_  | \new_[2254]_ ;
  assign \new_[2261]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[2264]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[2265]_  = \new_[2264]_  | \new_[2261]_ ;
  assign \new_[2266]_  = \new_[2265]_  | \new_[2258]_ ;
  assign \new_[2267]_  = \new_[2266]_  | \new_[2251]_ ;
  assign \new_[2268]_  = \new_[2267]_  | \new_[2236]_ ;
  assign \new_[2269]_  = \new_[2268]_  | \new_[2205]_ ;
  assign \new_[2270]_  = \new_[2269]_  | \new_[2144]_ ;
  assign \new_[2274]_  = \new_[377]_  | \new_[378]_ ;
  assign \new_[2275]_  = \new_[379]_  | \new_[2274]_ ;
  assign \new_[2278]_  = \new_[375]_  | \new_[376]_ ;
  assign \new_[2281]_  = \new_[373]_  | \new_[374]_ ;
  assign \new_[2282]_  = \new_[2281]_  | \new_[2278]_ ;
  assign \new_[2283]_  = \new_[2282]_  | \new_[2275]_ ;
  assign \new_[2286]_  = \new_[371]_  | \new_[372]_ ;
  assign \new_[2289]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[2290]_  = \new_[2289]_  | \new_[2286]_ ;
  assign \new_[2293]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[2296]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[2297]_  = \new_[2296]_  | \new_[2293]_ ;
  assign \new_[2298]_  = \new_[2297]_  | \new_[2290]_ ;
  assign \new_[2299]_  = \new_[2298]_  | \new_[2283]_ ;
  assign \new_[2302]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[2305]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[2306]_  = \new_[2305]_  | \new_[2302]_ ;
  assign \new_[2309]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[2312]_  = \new_[357]_  | \new_[358]_ ;
  assign \new_[2313]_  = \new_[2312]_  | \new_[2309]_ ;
  assign \new_[2314]_  = \new_[2313]_  | \new_[2306]_ ;
  assign \new_[2317]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[2320]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[2321]_  = \new_[2320]_  | \new_[2317]_ ;
  assign \new_[2324]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[2327]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[2328]_  = \new_[2327]_  | \new_[2324]_ ;
  assign \new_[2329]_  = \new_[2328]_  | \new_[2321]_ ;
  assign \new_[2330]_  = \new_[2329]_  | \new_[2314]_ ;
  assign \new_[2331]_  = \new_[2330]_  | \new_[2299]_ ;
  assign \new_[2334]_  = \new_[347]_  | \new_[348]_ ;
  assign \new_[2337]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[2338]_  = \new_[2337]_  | \new_[2334]_ ;
  assign \new_[2341]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[2344]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[2345]_  = \new_[2344]_  | \new_[2341]_ ;
  assign \new_[2346]_  = \new_[2345]_  | \new_[2338]_ ;
  assign \new_[2349]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[2352]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[2353]_  = \new_[2352]_  | \new_[2349]_ ;
  assign \new_[2356]_  = \new_[335]_  | \new_[336]_ ;
  assign \new_[2359]_  = \new_[333]_  | \new_[334]_ ;
  assign \new_[2360]_  = \new_[2359]_  | \new_[2356]_ ;
  assign \new_[2361]_  = \new_[2360]_  | \new_[2353]_ ;
  assign \new_[2362]_  = \new_[2361]_  | \new_[2346]_ ;
  assign \new_[2365]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[2368]_  = \new_[329]_  | \new_[330]_ ;
  assign \new_[2369]_  = \new_[2368]_  | \new_[2365]_ ;
  assign \new_[2372]_  = \new_[327]_  | \new_[328]_ ;
  assign \new_[2375]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[2376]_  = \new_[2375]_  | \new_[2372]_ ;
  assign \new_[2377]_  = \new_[2376]_  | \new_[2369]_ ;
  assign \new_[2380]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[2383]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[2384]_  = \new_[2383]_  | \new_[2380]_ ;
  assign \new_[2387]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[2390]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[2391]_  = \new_[2390]_  | \new_[2387]_ ;
  assign \new_[2392]_  = \new_[2391]_  | \new_[2384]_ ;
  assign \new_[2393]_  = \new_[2392]_  | \new_[2377]_ ;
  assign \new_[2394]_  = \new_[2393]_  | \new_[2362]_ ;
  assign \new_[2395]_  = \new_[2394]_  | \new_[2331]_ ;
  assign \new_[2399]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[2400]_  = \new_[316]_  | \new_[2399]_ ;
  assign \new_[2403]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[2406]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[2407]_  = \new_[2406]_  | \new_[2403]_ ;
  assign \new_[2408]_  = \new_[2407]_  | \new_[2400]_ ;
  assign \new_[2411]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[2414]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[2415]_  = \new_[2414]_  | \new_[2411]_ ;
  assign \new_[2418]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[2421]_  = \new_[302]_  | \new_[303]_ ;
  assign \new_[2422]_  = \new_[2421]_  | \new_[2418]_ ;
  assign \new_[2423]_  = \new_[2422]_  | \new_[2415]_ ;
  assign \new_[2424]_  = \new_[2423]_  | \new_[2408]_ ;
  assign \new_[2427]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[2430]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[2431]_  = \new_[2430]_  | \new_[2427]_ ;
  assign \new_[2434]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[2437]_  = \new_[294]_  | \new_[295]_ ;
  assign \new_[2438]_  = \new_[2437]_  | \new_[2434]_ ;
  assign \new_[2439]_  = \new_[2438]_  | \new_[2431]_ ;
  assign \new_[2442]_  = \new_[292]_  | \new_[293]_ ;
  assign \new_[2445]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[2446]_  = \new_[2445]_  | \new_[2442]_ ;
  assign \new_[2449]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[2452]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[2453]_  = \new_[2452]_  | \new_[2449]_ ;
  assign \new_[2454]_  = \new_[2453]_  | \new_[2446]_ ;
  assign \new_[2455]_  = \new_[2454]_  | \new_[2439]_ ;
  assign \new_[2456]_  = \new_[2455]_  | \new_[2424]_ ;
  assign \new_[2459]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[2462]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[2463]_  = \new_[2462]_  | \new_[2459]_ ;
  assign \new_[2466]_  = \new_[280]_  | \new_[281]_ ;
  assign \new_[2469]_  = \new_[278]_  | \new_[279]_ ;
  assign \new_[2470]_  = \new_[2469]_  | \new_[2466]_ ;
  assign \new_[2471]_  = \new_[2470]_  | \new_[2463]_ ;
  assign \new_[2474]_  = \new_[276]_  | \new_[277]_ ;
  assign \new_[2477]_  = \new_[274]_  | \new_[275]_ ;
  assign \new_[2478]_  = \new_[2477]_  | \new_[2474]_ ;
  assign \new_[2481]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[2484]_  = \new_[270]_  | \new_[271]_ ;
  assign \new_[2485]_  = \new_[2484]_  | \new_[2481]_ ;
  assign \new_[2486]_  = \new_[2485]_  | \new_[2478]_ ;
  assign \new_[2487]_  = \new_[2486]_  | \new_[2471]_ ;
  assign \new_[2490]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[2493]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[2494]_  = \new_[2493]_  | \new_[2490]_ ;
  assign \new_[2497]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[2500]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[2501]_  = \new_[2500]_  | \new_[2497]_ ;
  assign \new_[2502]_  = \new_[2501]_  | \new_[2494]_ ;
  assign \new_[2505]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[2508]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[2509]_  = \new_[2508]_  | \new_[2505]_ ;
  assign \new_[2512]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[2515]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[2516]_  = \new_[2515]_  | \new_[2512]_ ;
  assign \new_[2517]_  = \new_[2516]_  | \new_[2509]_ ;
  assign \new_[2518]_  = \new_[2517]_  | \new_[2502]_ ;
  assign \new_[2519]_  = \new_[2518]_  | \new_[2487]_ ;
  assign \new_[2520]_  = \new_[2519]_  | \new_[2456]_ ;
  assign \new_[2521]_  = \new_[2520]_  | \new_[2395]_ ;
  assign \new_[2522]_  = \new_[2521]_  | \new_[2270]_ ;
  assign \new_[2526]_  = \new_[251]_  | \new_[252]_ ;
  assign \new_[2527]_  = \new_[253]_  | \new_[2526]_ ;
  assign \new_[2530]_  = \new_[249]_  | \new_[250]_ ;
  assign \new_[2533]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[2534]_  = \new_[2533]_  | \new_[2530]_ ;
  assign \new_[2535]_  = \new_[2534]_  | \new_[2527]_ ;
  assign \new_[2538]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[2541]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[2542]_  = \new_[2541]_  | \new_[2538]_ ;
  assign \new_[2545]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[2548]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[2549]_  = \new_[2548]_  | \new_[2545]_ ;
  assign \new_[2550]_  = \new_[2549]_  | \new_[2542]_ ;
  assign \new_[2551]_  = \new_[2550]_  | \new_[2535]_ ;
  assign \new_[2554]_  = \new_[237]_  | \new_[238]_ ;
  assign \new_[2557]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[2558]_  = \new_[2557]_  | \new_[2554]_ ;
  assign \new_[2561]_  = \new_[233]_  | \new_[234]_ ;
  assign \new_[2564]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[2565]_  = \new_[2564]_  | \new_[2561]_ ;
  assign \new_[2566]_  = \new_[2565]_  | \new_[2558]_ ;
  assign \new_[2569]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[2572]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[2573]_  = \new_[2572]_  | \new_[2569]_ ;
  assign \new_[2576]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[2579]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[2580]_  = \new_[2579]_  | \new_[2576]_ ;
  assign \new_[2581]_  = \new_[2580]_  | \new_[2573]_ ;
  assign \new_[2582]_  = \new_[2581]_  | \new_[2566]_ ;
  assign \new_[2583]_  = \new_[2582]_  | \new_[2551]_ ;
  assign \new_[2586]_  = \new_[221]_  | \new_[222]_ ;
  assign \new_[2589]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[2590]_  = \new_[2589]_  | \new_[2586]_ ;
  assign \new_[2593]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[2596]_  = \new_[215]_  | \new_[216]_ ;
  assign \new_[2597]_  = \new_[2596]_  | \new_[2593]_ ;
  assign \new_[2598]_  = \new_[2597]_  | \new_[2590]_ ;
  assign \new_[2601]_  = \new_[213]_  | \new_[214]_ ;
  assign \new_[2604]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[2605]_  = \new_[2604]_  | \new_[2601]_ ;
  assign \new_[2608]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[2611]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[2612]_  = \new_[2611]_  | \new_[2608]_ ;
  assign \new_[2613]_  = \new_[2612]_  | \new_[2605]_ ;
  assign \new_[2614]_  = \new_[2613]_  | \new_[2598]_ ;
  assign \new_[2617]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[2620]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[2621]_  = \new_[2620]_  | \new_[2617]_ ;
  assign \new_[2624]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[2627]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[2628]_  = \new_[2627]_  | \new_[2624]_ ;
  assign \new_[2629]_  = \new_[2628]_  | \new_[2621]_ ;
  assign \new_[2632]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[2635]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[2636]_  = \new_[2635]_  | \new_[2632]_ ;
  assign \new_[2639]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[2642]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[2643]_  = \new_[2642]_  | \new_[2639]_ ;
  assign \new_[2644]_  = \new_[2643]_  | \new_[2636]_ ;
  assign \new_[2645]_  = \new_[2644]_  | \new_[2629]_ ;
  assign \new_[2646]_  = \new_[2645]_  | \new_[2614]_ ;
  assign \new_[2647]_  = \new_[2646]_  | \new_[2583]_ ;
  assign \new_[2651]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[2652]_  = \new_[190]_  | \new_[2651]_ ;
  assign \new_[2655]_  = \new_[186]_  | \new_[187]_ ;
  assign \new_[2658]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[2659]_  = \new_[2658]_  | \new_[2655]_ ;
  assign \new_[2660]_  = \new_[2659]_  | \new_[2652]_ ;
  assign \new_[2663]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[2666]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[2667]_  = \new_[2666]_  | \new_[2663]_ ;
  assign \new_[2670]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[2673]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[2674]_  = \new_[2673]_  | \new_[2670]_ ;
  assign \new_[2675]_  = \new_[2674]_  | \new_[2667]_ ;
  assign \new_[2676]_  = \new_[2675]_  | \new_[2660]_ ;
  assign \new_[2679]_  = \new_[174]_  | \new_[175]_ ;
  assign \new_[2682]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[2683]_  = \new_[2682]_  | \new_[2679]_ ;
  assign \new_[2686]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[2689]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[2690]_  = \new_[2689]_  | \new_[2686]_ ;
  assign \new_[2691]_  = \new_[2690]_  | \new_[2683]_ ;
  assign \new_[2694]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[2697]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[2698]_  = \new_[2697]_  | \new_[2694]_ ;
  assign \new_[2701]_  = \new_[162]_  | \new_[163]_ ;
  assign \new_[2704]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[2705]_  = \new_[2704]_  | \new_[2701]_ ;
  assign \new_[2706]_  = \new_[2705]_  | \new_[2698]_ ;
  assign \new_[2707]_  = \new_[2706]_  | \new_[2691]_ ;
  assign \new_[2708]_  = \new_[2707]_  | \new_[2676]_ ;
  assign \new_[2711]_  = \new_[158]_  | \new_[159]_ ;
  assign \new_[2714]_  = \new_[156]_  | \new_[157]_ ;
  assign \new_[2715]_  = \new_[2714]_  | \new_[2711]_ ;
  assign \new_[2718]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[2721]_  = \new_[152]_  | \new_[153]_ ;
  assign \new_[2722]_  = \new_[2721]_  | \new_[2718]_ ;
  assign \new_[2723]_  = \new_[2722]_  | \new_[2715]_ ;
  assign \new_[2726]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[2729]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[2730]_  = \new_[2729]_  | \new_[2726]_ ;
  assign \new_[2733]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[2736]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[2737]_  = \new_[2736]_  | \new_[2733]_ ;
  assign \new_[2738]_  = \new_[2737]_  | \new_[2730]_ ;
  assign \new_[2739]_  = \new_[2738]_  | \new_[2723]_ ;
  assign \new_[2742]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[2745]_  = \new_[140]_  | \new_[141]_ ;
  assign \new_[2746]_  = \new_[2745]_  | \new_[2742]_ ;
  assign \new_[2749]_  = \new_[138]_  | \new_[139]_ ;
  assign \new_[2752]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[2753]_  = \new_[2752]_  | \new_[2749]_ ;
  assign \new_[2754]_  = \new_[2753]_  | \new_[2746]_ ;
  assign \new_[2757]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[2760]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[2761]_  = \new_[2760]_  | \new_[2757]_ ;
  assign \new_[2764]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[2767]_  = \new_[128]_  | \new_[129]_ ;
  assign \new_[2768]_  = \new_[2767]_  | \new_[2764]_ ;
  assign \new_[2769]_  = \new_[2768]_  | \new_[2761]_ ;
  assign \new_[2770]_  = \new_[2769]_  | \new_[2754]_ ;
  assign \new_[2771]_  = \new_[2770]_  | \new_[2739]_ ;
  assign \new_[2772]_  = \new_[2771]_  | \new_[2708]_ ;
  assign \new_[2773]_  = \new_[2772]_  | \new_[2647]_ ;
  assign \new_[2777]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[2778]_  = \new_[127]_  | \new_[2777]_ ;
  assign \new_[2781]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[2784]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[2785]_  = \new_[2784]_  | \new_[2781]_ ;
  assign \new_[2786]_  = \new_[2785]_  | \new_[2778]_ ;
  assign \new_[2789]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[2792]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[2793]_  = \new_[2792]_  | \new_[2789]_ ;
  assign \new_[2796]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[2799]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[2800]_  = \new_[2799]_  | \new_[2796]_ ;
  assign \new_[2801]_  = \new_[2800]_  | \new_[2793]_ ;
  assign \new_[2802]_  = \new_[2801]_  | \new_[2786]_ ;
  assign \new_[2805]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[2808]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[2809]_  = \new_[2808]_  | \new_[2805]_ ;
  assign \new_[2812]_  = \new_[107]_  | \new_[108]_ ;
  assign \new_[2815]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[2816]_  = \new_[2815]_  | \new_[2812]_ ;
  assign \new_[2817]_  = \new_[2816]_  | \new_[2809]_ ;
  assign \new_[2820]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[2823]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[2824]_  = \new_[2823]_  | \new_[2820]_ ;
  assign \new_[2827]_  = \new_[99]_  | \new_[100]_ ;
  assign \new_[2830]_  = \new_[97]_  | \new_[98]_ ;
  assign \new_[2831]_  = \new_[2830]_  | \new_[2827]_ ;
  assign \new_[2832]_  = \new_[2831]_  | \new_[2824]_ ;
  assign \new_[2833]_  = \new_[2832]_  | \new_[2817]_ ;
  assign \new_[2834]_  = \new_[2833]_  | \new_[2802]_ ;
  assign \new_[2837]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[2840]_  = \new_[93]_  | \new_[94]_ ;
  assign \new_[2841]_  = \new_[2840]_  | \new_[2837]_ ;
  assign \new_[2844]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[2847]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[2848]_  = \new_[2847]_  | \new_[2844]_ ;
  assign \new_[2849]_  = \new_[2848]_  | \new_[2841]_ ;
  assign \new_[2852]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[2855]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[2856]_  = \new_[2855]_  | \new_[2852]_ ;
  assign \new_[2859]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[2862]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[2863]_  = \new_[2862]_  | \new_[2859]_ ;
  assign \new_[2864]_  = \new_[2863]_  | \new_[2856]_ ;
  assign \new_[2865]_  = \new_[2864]_  | \new_[2849]_ ;
  assign \new_[2868]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[2871]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[2872]_  = \new_[2871]_  | \new_[2868]_ ;
  assign \new_[2875]_  = \new_[75]_  | \new_[76]_ ;
  assign \new_[2878]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[2879]_  = \new_[2878]_  | \new_[2875]_ ;
  assign \new_[2880]_  = \new_[2879]_  | \new_[2872]_ ;
  assign \new_[2883]_  = \new_[71]_  | \new_[72]_ ;
  assign \new_[2886]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[2887]_  = \new_[2886]_  | \new_[2883]_ ;
  assign \new_[2890]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[2893]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[2894]_  = \new_[2893]_  | \new_[2890]_ ;
  assign \new_[2895]_  = \new_[2894]_  | \new_[2887]_ ;
  assign \new_[2896]_  = \new_[2895]_  | \new_[2880]_ ;
  assign \new_[2897]_  = \new_[2896]_  | \new_[2865]_ ;
  assign \new_[2898]_  = \new_[2897]_  | \new_[2834]_ ;
  assign \new_[2901]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[2904]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[2905]_  = \new_[2904]_  | \new_[2901]_ ;
  assign \new_[2908]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[2911]_  = \new_[57]_  | \new_[58]_ ;
  assign \new_[2912]_  = \new_[2911]_  | \new_[2908]_ ;
  assign \new_[2913]_  = \new_[2912]_  | \new_[2905]_ ;
  assign \new_[2916]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[2919]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[2920]_  = \new_[2919]_  | \new_[2916]_ ;
  assign \new_[2923]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[2926]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[2927]_  = \new_[2926]_  | \new_[2923]_ ;
  assign \new_[2928]_  = \new_[2927]_  | \new_[2920]_ ;
  assign \new_[2929]_  = \new_[2928]_  | \new_[2913]_ ;
  assign \new_[2932]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[2935]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[2936]_  = \new_[2935]_  | \new_[2932]_ ;
  assign \new_[2939]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[2942]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[2943]_  = \new_[2942]_  | \new_[2939]_ ;
  assign \new_[2944]_  = \new_[2943]_  | \new_[2936]_ ;
  assign \new_[2947]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[2950]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[2951]_  = \new_[2950]_  | \new_[2947]_ ;
  assign \new_[2954]_  = \new_[35]_  | \new_[36]_ ;
  assign \new_[2957]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[2958]_  = \new_[2957]_  | \new_[2954]_ ;
  assign \new_[2959]_  = \new_[2958]_  | \new_[2951]_ ;
  assign \new_[2960]_  = \new_[2959]_  | \new_[2944]_ ;
  assign \new_[2961]_  = \new_[2960]_  | \new_[2929]_ ;
  assign \new_[2964]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[2967]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[2968]_  = \new_[2967]_  | \new_[2964]_ ;
  assign \new_[2971]_  = \new_[27]_  | \new_[28]_ ;
  assign \new_[2974]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[2975]_  = \new_[2974]_  | \new_[2971]_ ;
  assign \new_[2976]_  = \new_[2975]_  | \new_[2968]_ ;
  assign \new_[2979]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[2982]_  = \new_[21]_  | \new_[22]_ ;
  assign \new_[2983]_  = \new_[2982]_  | \new_[2979]_ ;
  assign \new_[2986]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[2989]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[2990]_  = \new_[2989]_  | \new_[2986]_ ;
  assign \new_[2991]_  = \new_[2990]_  | \new_[2983]_ ;
  assign \new_[2992]_  = \new_[2991]_  | \new_[2976]_ ;
  assign \new_[2995]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[2998]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[2999]_  = \new_[2998]_  | \new_[2995]_ ;
  assign \new_[3002]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[3005]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[3006]_  = \new_[3005]_  | \new_[3002]_ ;
  assign \new_[3007]_  = \new_[3006]_  | \new_[2999]_ ;
  assign \new_[3010]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[3013]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[3014]_  = \new_[3013]_  | \new_[3010]_ ;
  assign \new_[3017]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[3020]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[3021]_  = \new_[3020]_  | \new_[3017]_ ;
  assign \new_[3022]_  = \new_[3021]_  | \new_[3014]_ ;
  assign \new_[3023]_  = \new_[3022]_  | \new_[3007]_ ;
  assign \new_[3024]_  = \new_[3023]_  | \new_[2992]_ ;
  assign \new_[3025]_  = \new_[3024]_  | \new_[2961]_ ;
  assign \new_[3026]_  = \new_[3025]_  | \new_[2898]_ ;
  assign \new_[3027]_  = \new_[3026]_  | \new_[2773]_ ;
  assign \new_[3028]_  = \new_[3027]_  | \new_[2522]_ ;
  assign \new_[3036]_  = A234 & A232;
  assign \new_[3040]_  = A234 & A233;
  assign \new_[3044]_  = A235 & A201;
  assign \new_[3048]_  = A235 & A201;
  assign \new_[3052]_  = A235 & A166;
  assign \new_[3056]_  = A235 & A167;
  assign \new_[3060]_  = A234 & A232;
  assign \new_[3064]_  = A234 & A233;
  assign \new_[3067]_  = ~A232 & A202;
  assign \new_[3070]_  = A236 & A233;
  assign \new_[3073]_  = A232 & A202;
  assign \new_[3076]_  = A236 & ~A233;
  assign \new_[3079]_  = A201 & A199;
  assign \new_[3082]_  = A234 & A232;
  assign \new_[3085]_  = A201 & A199;
  assign \new_[3088]_  = A234 & A233;
  assign \new_[3091]_  = A201 & A200;
  assign \new_[3094]_  = A234 & A232;
  assign \new_[3097]_  = A201 & A200;
  assign \new_[3100]_  = A234 & A233;
  assign \new_[3103]_  = A200 & ~A199;
  assign \new_[3106]_  = A235 & A203;
  assign \new_[3109]_  = ~A200 & A199;
  assign \new_[3112]_  = A235 & A203;
  assign \new_[3115]_  = A166 & A168;
  assign \new_[3118]_  = A234 & A232;
  assign \new_[3121]_  = A166 & A168;
  assign \new_[3124]_  = A234 & A233;
  assign \new_[3127]_  = A167 & A168;
  assign \new_[3130]_  = A234 & A232;
  assign \new_[3133]_  = A167 & A168;
  assign \new_[3136]_  = A234 & A233;
  assign \new_[3139]_  = A167 & A170;
  assign \new_[3142]_  = A235 & ~A166;
  assign \new_[3145]_  = ~A167 & A170;
  assign \new_[3148]_  = A235 & A166;
  assign \new_[3151]_  = ~A232 & A169;
  assign \new_[3154]_  = A236 & A233;
  assign \new_[3157]_  = A232 & A169;
  assign \new_[3160]_  = A236 & ~A233;
  assign \new_[3163]_  = A201 & A199;
  assign \new_[3167]_  = A236 & A233;
  assign \new_[3168]_  = ~A232 & \new_[3167]_ ;
  assign \new_[3171]_  = A201 & A199;
  assign \new_[3175]_  = A236 & ~A233;
  assign \new_[3176]_  = A232 & \new_[3175]_ ;
  assign \new_[3179]_  = A201 & A200;
  assign \new_[3183]_  = A236 & A233;
  assign \new_[3184]_  = ~A232 & \new_[3183]_ ;
  assign \new_[3187]_  = A201 & A200;
  assign \new_[3191]_  = A236 & ~A233;
  assign \new_[3192]_  = A232 & \new_[3191]_ ;
  assign \new_[3195]_  = A200 & ~A199;
  assign \new_[3199]_  = A234 & A232;
  assign \new_[3200]_  = A203 & \new_[3199]_ ;
  assign \new_[3203]_  = A200 & ~A199;
  assign \new_[3207]_  = A234 & A233;
  assign \new_[3208]_  = A203 & \new_[3207]_ ;
  assign \new_[3211]_  = ~A200 & A199;
  assign \new_[3215]_  = A234 & A232;
  assign \new_[3216]_  = A203 & \new_[3215]_ ;
  assign \new_[3219]_  = ~A200 & A199;
  assign \new_[3223]_  = A234 & A233;
  assign \new_[3224]_  = A203 & \new_[3223]_ ;
  assign \new_[3227]_  = A166 & A168;
  assign \new_[3231]_  = A236 & A233;
  assign \new_[3232]_  = ~A232 & \new_[3231]_ ;
  assign \new_[3235]_  = A166 & A168;
  assign \new_[3239]_  = A236 & ~A233;
  assign \new_[3240]_  = A232 & \new_[3239]_ ;
  assign \new_[3243]_  = A167 & A168;
  assign \new_[3247]_  = A236 & A233;
  assign \new_[3248]_  = ~A232 & \new_[3247]_ ;
  assign \new_[3251]_  = A167 & A168;
  assign \new_[3255]_  = A236 & ~A233;
  assign \new_[3256]_  = A232 & \new_[3255]_ ;
  assign \new_[3259]_  = A167 & A170;
  assign \new_[3263]_  = A234 & A232;
  assign \new_[3264]_  = ~A166 & \new_[3263]_ ;
  assign \new_[3267]_  = A167 & A170;
  assign \new_[3271]_  = A234 & A233;
  assign \new_[3272]_  = ~A166 & \new_[3271]_ ;
  assign \new_[3275]_  = ~A167 & A170;
  assign \new_[3279]_  = A234 & A232;
  assign \new_[3280]_  = A166 & \new_[3279]_ ;
  assign \new_[3283]_  = ~A167 & A170;
  assign \new_[3287]_  = A234 & A233;
  assign \new_[3288]_  = A166 & \new_[3287]_ ;
  assign \new_[3292]_  = A203 & A200;
  assign \new_[3293]_  = ~A199 & \new_[3292]_ ;
  assign \new_[3297]_  = A236 & A233;
  assign \new_[3298]_  = ~A232 & \new_[3297]_ ;
  assign \new_[3302]_  = A203 & A200;
  assign \new_[3303]_  = ~A199 & \new_[3302]_ ;
  assign \new_[3307]_  = A236 & ~A233;
  assign \new_[3308]_  = A232 & \new_[3307]_ ;
  assign \new_[3312]_  = A203 & ~A200;
  assign \new_[3313]_  = A199 & \new_[3312]_ ;
  assign \new_[3317]_  = A236 & A233;
  assign \new_[3318]_  = ~A232 & \new_[3317]_ ;
  assign \new_[3322]_  = A203 & ~A200;
  assign \new_[3323]_  = A199 & \new_[3322]_ ;
  assign \new_[3327]_  = A236 & ~A233;
  assign \new_[3328]_  = A232 & \new_[3327]_ ;
  assign \new_[3332]_  = ~A166 & A167;
  assign \new_[3333]_  = A170 & \new_[3332]_ ;
  assign \new_[3337]_  = A236 & A233;
  assign \new_[3338]_  = ~A232 & \new_[3337]_ ;
  assign \new_[3342]_  = ~A166 & A167;
  assign \new_[3343]_  = A170 & \new_[3342]_ ;
  assign \new_[3347]_  = A236 & ~A233;
  assign \new_[3348]_  = A232 & \new_[3347]_ ;
  assign \new_[3352]_  = A166 & ~A167;
  assign \new_[3353]_  = A170 & \new_[3352]_ ;
  assign \new_[3357]_  = A236 & A233;
  assign \new_[3358]_  = ~A232 & \new_[3357]_ ;
  assign \new_[3362]_  = A166 & ~A167;
  assign \new_[3363]_  = A170 & \new_[3362]_ ;
  assign \new_[3367]_  = A236 & ~A233;
  assign \new_[3368]_  = A232 & \new_[3367]_ ;
  assign \new_[3372]_  = A268 & A202;
  assign \new_[3373]_  = A169 & \new_[3372]_ ;
  assign \new_[3377]_  = ~A302 & ~A301;
  assign \new_[3378]_  = ~A300 & \new_[3377]_ ;
  assign \new_[3382]_  = A268 & A202;
  assign \new_[3383]_  = A169 & \new_[3382]_ ;
  assign \new_[3387]_  = ~A301 & ~A299;
  assign \new_[3388]_  = ~A298 & \new_[3387]_ ;
  assign \new_[3392]_  = A202 & A166;
  assign \new_[3393]_  = A168 & \new_[3392]_ ;
  assign \new_[3396]_  = ~A300 & A268;
  assign \new_[3399]_  = ~A302 & ~A301;
  assign \new_[3400]_  = \new_[3399]_  & \new_[3396]_ ;
  assign \new_[3404]_  = A202 & A166;
  assign \new_[3405]_  = A168 & \new_[3404]_ ;
  assign \new_[3408]_  = ~A298 & A268;
  assign \new_[3411]_  = ~A301 & ~A299;
  assign \new_[3412]_  = \new_[3411]_  & \new_[3408]_ ;
  assign \new_[3416]_  = A202 & A167;
  assign \new_[3417]_  = A168 & \new_[3416]_ ;
  assign \new_[3420]_  = ~A300 & A268;
  assign \new_[3423]_  = ~A302 & ~A301;
  assign \new_[3424]_  = \new_[3423]_  & \new_[3420]_ ;
  assign \new_[3428]_  = A202 & A167;
  assign \new_[3429]_  = A168 & \new_[3428]_ ;
  assign \new_[3432]_  = ~A298 & A268;
  assign \new_[3435]_  = ~A301 & ~A299;
  assign \new_[3436]_  = \new_[3435]_  & \new_[3432]_ ;
  assign \new_[3440]_  = A268 & A202;
  assign \new_[3441]_  = A169 & \new_[3440]_ ;
  assign \new_[3444]_  = A299 & A298;
  assign \new_[3447]_  = ~A301 & ~A300;
  assign \new_[3448]_  = \new_[3447]_  & \new_[3444]_ ;
  assign \new_[3452]_  = A265 & A202;
  assign \new_[3453]_  = A169 & \new_[3452]_ ;
  assign \new_[3456]_  = ~A300 & A267;
  assign \new_[3459]_  = ~A302 & ~A301;
  assign \new_[3460]_  = \new_[3459]_  & \new_[3456]_ ;
  assign \new_[3464]_  = A265 & A202;
  assign \new_[3465]_  = A169 & \new_[3464]_ ;
  assign \new_[3468]_  = ~A298 & A267;
  assign \new_[3471]_  = ~A301 & ~A299;
  assign \new_[3472]_  = \new_[3471]_  & \new_[3468]_ ;
  assign \new_[3476]_  = A266 & A202;
  assign \new_[3477]_  = A169 & \new_[3476]_ ;
  assign \new_[3480]_  = ~A300 & A267;
  assign \new_[3483]_  = ~A302 & ~A301;
  assign \new_[3484]_  = \new_[3483]_  & \new_[3480]_ ;
  assign \new_[3488]_  = A266 & A202;
  assign \new_[3489]_  = A169 & \new_[3488]_ ;
  assign \new_[3492]_  = ~A298 & A267;
  assign \new_[3495]_  = ~A301 & ~A299;
  assign \new_[3496]_  = \new_[3495]_  & \new_[3492]_ ;
  assign \new_[3500]_  = A201 & A199;
  assign \new_[3501]_  = A169 & \new_[3500]_ ;
  assign \new_[3504]_  = ~A300 & A268;
  assign \new_[3507]_  = ~A302 & ~A301;
  assign \new_[3508]_  = \new_[3507]_  & \new_[3504]_ ;
  assign \new_[3512]_  = A201 & A199;
  assign \new_[3513]_  = A169 & \new_[3512]_ ;
  assign \new_[3516]_  = ~A298 & A268;
  assign \new_[3519]_  = ~A301 & ~A299;
  assign \new_[3520]_  = \new_[3519]_  & \new_[3516]_ ;
  assign \new_[3524]_  = A201 & A200;
  assign \new_[3525]_  = A169 & \new_[3524]_ ;
  assign \new_[3528]_  = ~A300 & A268;
  assign \new_[3531]_  = ~A302 & ~A301;
  assign \new_[3532]_  = \new_[3531]_  & \new_[3528]_ ;
  assign \new_[3536]_  = A201 & A200;
  assign \new_[3537]_  = A169 & \new_[3536]_ ;
  assign \new_[3540]_  = ~A298 & A268;
  assign \new_[3543]_  = ~A301 & ~A299;
  assign \new_[3544]_  = \new_[3543]_  & \new_[3540]_ ;
  assign \new_[3547]_  = A166 & A168;
  assign \new_[3550]_  = A268 & A202;
  assign \new_[3551]_  = \new_[3550]_  & \new_[3547]_ ;
  assign \new_[3554]_  = A299 & A298;
  assign \new_[3557]_  = ~A301 & ~A300;
  assign \new_[3558]_  = \new_[3557]_  & \new_[3554]_ ;
  assign \new_[3561]_  = A166 & A168;
  assign \new_[3564]_  = A265 & A202;
  assign \new_[3565]_  = \new_[3564]_  & \new_[3561]_ ;
  assign \new_[3568]_  = ~A300 & A267;
  assign \new_[3571]_  = ~A302 & ~A301;
  assign \new_[3572]_  = \new_[3571]_  & \new_[3568]_ ;
  assign \new_[3575]_  = A166 & A168;
  assign \new_[3578]_  = A265 & A202;
  assign \new_[3579]_  = \new_[3578]_  & \new_[3575]_ ;
  assign \new_[3582]_  = ~A298 & A267;
  assign \new_[3585]_  = ~A301 & ~A299;
  assign \new_[3586]_  = \new_[3585]_  & \new_[3582]_ ;
  assign \new_[3589]_  = A166 & A168;
  assign \new_[3592]_  = A266 & A202;
  assign \new_[3593]_  = \new_[3592]_  & \new_[3589]_ ;
  assign \new_[3596]_  = ~A300 & A267;
  assign \new_[3599]_  = ~A302 & ~A301;
  assign \new_[3600]_  = \new_[3599]_  & \new_[3596]_ ;
  assign \new_[3603]_  = A166 & A168;
  assign \new_[3606]_  = A266 & A202;
  assign \new_[3607]_  = \new_[3606]_  & \new_[3603]_ ;
  assign \new_[3610]_  = ~A298 & A267;
  assign \new_[3613]_  = ~A301 & ~A299;
  assign \new_[3614]_  = \new_[3613]_  & \new_[3610]_ ;
  assign \new_[3617]_  = A166 & A168;
  assign \new_[3620]_  = A201 & A199;
  assign \new_[3621]_  = \new_[3620]_  & \new_[3617]_ ;
  assign \new_[3624]_  = ~A300 & A268;
  assign \new_[3627]_  = ~A302 & ~A301;
  assign \new_[3628]_  = \new_[3627]_  & \new_[3624]_ ;
  assign \new_[3631]_  = A166 & A168;
  assign \new_[3634]_  = A201 & A199;
  assign \new_[3635]_  = \new_[3634]_  & \new_[3631]_ ;
  assign \new_[3638]_  = ~A298 & A268;
  assign \new_[3641]_  = ~A301 & ~A299;
  assign \new_[3642]_  = \new_[3641]_  & \new_[3638]_ ;
  assign \new_[3645]_  = A166 & A168;
  assign \new_[3648]_  = A201 & A200;
  assign \new_[3649]_  = \new_[3648]_  & \new_[3645]_ ;
  assign \new_[3652]_  = ~A300 & A268;
  assign \new_[3655]_  = ~A302 & ~A301;
  assign \new_[3656]_  = \new_[3655]_  & \new_[3652]_ ;
  assign \new_[3659]_  = A166 & A168;
  assign \new_[3662]_  = A201 & A200;
  assign \new_[3663]_  = \new_[3662]_  & \new_[3659]_ ;
  assign \new_[3666]_  = ~A298 & A268;
  assign \new_[3669]_  = ~A301 & ~A299;
  assign \new_[3670]_  = \new_[3669]_  & \new_[3666]_ ;
  assign \new_[3673]_  = A167 & A168;
  assign \new_[3676]_  = A268 & A202;
  assign \new_[3677]_  = \new_[3676]_  & \new_[3673]_ ;
  assign \new_[3680]_  = A299 & A298;
  assign \new_[3683]_  = ~A301 & ~A300;
  assign \new_[3684]_  = \new_[3683]_  & \new_[3680]_ ;
  assign \new_[3687]_  = A167 & A168;
  assign \new_[3690]_  = A265 & A202;
  assign \new_[3691]_  = \new_[3690]_  & \new_[3687]_ ;
  assign \new_[3694]_  = ~A300 & A267;
  assign \new_[3697]_  = ~A302 & ~A301;
  assign \new_[3698]_  = \new_[3697]_  & \new_[3694]_ ;
  assign \new_[3701]_  = A167 & A168;
  assign \new_[3704]_  = A265 & A202;
  assign \new_[3705]_  = \new_[3704]_  & \new_[3701]_ ;
  assign \new_[3708]_  = ~A298 & A267;
  assign \new_[3711]_  = ~A301 & ~A299;
  assign \new_[3712]_  = \new_[3711]_  & \new_[3708]_ ;
  assign \new_[3715]_  = A167 & A168;
  assign \new_[3718]_  = A266 & A202;
  assign \new_[3719]_  = \new_[3718]_  & \new_[3715]_ ;
  assign \new_[3722]_  = ~A300 & A267;
  assign \new_[3725]_  = ~A302 & ~A301;
  assign \new_[3726]_  = \new_[3725]_  & \new_[3722]_ ;
  assign \new_[3729]_  = A167 & A168;
  assign \new_[3732]_  = A266 & A202;
  assign \new_[3733]_  = \new_[3732]_  & \new_[3729]_ ;
  assign \new_[3736]_  = ~A298 & A267;
  assign \new_[3739]_  = ~A301 & ~A299;
  assign \new_[3740]_  = \new_[3739]_  & \new_[3736]_ ;
  assign \new_[3743]_  = A167 & A168;
  assign \new_[3746]_  = A201 & A199;
  assign \new_[3747]_  = \new_[3746]_  & \new_[3743]_ ;
  assign \new_[3750]_  = ~A300 & A268;
  assign \new_[3753]_  = ~A302 & ~A301;
  assign \new_[3754]_  = \new_[3753]_  & \new_[3750]_ ;
  assign \new_[3757]_  = A167 & A168;
  assign \new_[3760]_  = A201 & A199;
  assign \new_[3761]_  = \new_[3760]_  & \new_[3757]_ ;
  assign \new_[3764]_  = ~A298 & A268;
  assign \new_[3767]_  = ~A301 & ~A299;
  assign \new_[3768]_  = \new_[3767]_  & \new_[3764]_ ;
  assign \new_[3771]_  = A167 & A168;
  assign \new_[3774]_  = A201 & A200;
  assign \new_[3775]_  = \new_[3774]_  & \new_[3771]_ ;
  assign \new_[3778]_  = ~A300 & A268;
  assign \new_[3781]_  = ~A302 & ~A301;
  assign \new_[3782]_  = \new_[3781]_  & \new_[3778]_ ;
  assign \new_[3785]_  = A167 & A168;
  assign \new_[3788]_  = A201 & A200;
  assign \new_[3789]_  = \new_[3788]_  & \new_[3785]_ ;
  assign \new_[3792]_  = ~A298 & A268;
  assign \new_[3795]_  = ~A301 & ~A299;
  assign \new_[3796]_  = \new_[3795]_  & \new_[3792]_ ;
  assign \new_[3799]_  = A167 & A170;
  assign \new_[3802]_  = A202 & ~A166;
  assign \new_[3803]_  = \new_[3802]_  & \new_[3799]_ ;
  assign \new_[3806]_  = ~A300 & A268;
  assign \new_[3809]_  = ~A302 & ~A301;
  assign \new_[3810]_  = \new_[3809]_  & \new_[3806]_ ;
  assign \new_[3813]_  = A167 & A170;
  assign \new_[3816]_  = A202 & ~A166;
  assign \new_[3817]_  = \new_[3816]_  & \new_[3813]_ ;
  assign \new_[3820]_  = ~A298 & A268;
  assign \new_[3823]_  = ~A301 & ~A299;
  assign \new_[3824]_  = \new_[3823]_  & \new_[3820]_ ;
  assign \new_[3827]_  = ~A167 & A170;
  assign \new_[3830]_  = A202 & A166;
  assign \new_[3831]_  = \new_[3830]_  & \new_[3827]_ ;
  assign \new_[3834]_  = ~A300 & A268;
  assign \new_[3837]_  = ~A302 & ~A301;
  assign \new_[3838]_  = \new_[3837]_  & \new_[3834]_ ;
  assign \new_[3841]_  = ~A167 & A170;
  assign \new_[3844]_  = A202 & A166;
  assign \new_[3845]_  = \new_[3844]_  & \new_[3841]_ ;
  assign \new_[3848]_  = ~A298 & A268;
  assign \new_[3851]_  = ~A301 & ~A299;
  assign \new_[3852]_  = \new_[3851]_  & \new_[3848]_ ;
  assign \new_[3855]_  = A202 & A169;
  assign \new_[3858]_  = A267 & A265;
  assign \new_[3859]_  = \new_[3858]_  & \new_[3855]_ ;
  assign \new_[3862]_  = A299 & A298;
  assign \new_[3865]_  = ~A301 & ~A300;
  assign \new_[3866]_  = \new_[3865]_  & \new_[3862]_ ;
  assign \new_[3869]_  = A202 & A169;
  assign \new_[3872]_  = A267 & A266;
  assign \new_[3873]_  = \new_[3872]_  & \new_[3869]_ ;
  assign \new_[3876]_  = A299 & A298;
  assign \new_[3879]_  = ~A301 & ~A300;
  assign \new_[3880]_  = \new_[3879]_  & \new_[3876]_ ;
  assign \new_[3883]_  = A202 & A169;
  assign \new_[3886]_  = A266 & ~A265;
  assign \new_[3887]_  = \new_[3886]_  & \new_[3883]_ ;
  assign \new_[3890]_  = ~A300 & A269;
  assign \new_[3893]_  = ~A302 & ~A301;
  assign \new_[3894]_  = \new_[3893]_  & \new_[3890]_ ;
  assign \new_[3897]_  = A202 & A169;
  assign \new_[3900]_  = A266 & ~A265;
  assign \new_[3901]_  = \new_[3900]_  & \new_[3897]_ ;
  assign \new_[3904]_  = ~A298 & A269;
  assign \new_[3907]_  = ~A301 & ~A299;
  assign \new_[3908]_  = \new_[3907]_  & \new_[3904]_ ;
  assign \new_[3911]_  = A202 & A169;
  assign \new_[3914]_  = ~A266 & A265;
  assign \new_[3915]_  = \new_[3914]_  & \new_[3911]_ ;
  assign \new_[3918]_  = ~A300 & A269;
  assign \new_[3921]_  = ~A302 & ~A301;
  assign \new_[3922]_  = \new_[3921]_  & \new_[3918]_ ;
  assign \new_[3925]_  = A202 & A169;
  assign \new_[3928]_  = ~A266 & A265;
  assign \new_[3929]_  = \new_[3928]_  & \new_[3925]_ ;
  assign \new_[3932]_  = ~A298 & A269;
  assign \new_[3935]_  = ~A301 & ~A299;
  assign \new_[3936]_  = \new_[3935]_  & \new_[3932]_ ;
  assign \new_[3939]_  = ~A201 & A169;
  assign \new_[3942]_  = ~A203 & ~A202;
  assign \new_[3943]_  = \new_[3942]_  & \new_[3939]_ ;
  assign \new_[3946]_  = ~A268 & ~A267;
  assign \new_[3949]_  = A301 & ~A269;
  assign \new_[3950]_  = \new_[3949]_  & \new_[3946]_ ;
  assign \new_[3953]_  = ~A201 & A169;
  assign \new_[3956]_  = ~A203 & ~A202;
  assign \new_[3957]_  = \new_[3956]_  & \new_[3953]_ ;
  assign \new_[3960]_  = ~A266 & ~A265;
  assign \new_[3963]_  = A301 & ~A268;
  assign \new_[3964]_  = \new_[3963]_  & \new_[3960]_ ;
  assign \new_[3967]_  = A199 & A169;
  assign \new_[3970]_  = A268 & A201;
  assign \new_[3971]_  = \new_[3970]_  & \new_[3967]_ ;
  assign \new_[3974]_  = A299 & A298;
  assign \new_[3977]_  = ~A301 & ~A300;
  assign \new_[3978]_  = \new_[3977]_  & \new_[3974]_ ;
  assign \new_[3981]_  = A199 & A169;
  assign \new_[3984]_  = A265 & A201;
  assign \new_[3985]_  = \new_[3984]_  & \new_[3981]_ ;
  assign \new_[3988]_  = ~A300 & A267;
  assign \new_[3991]_  = ~A302 & ~A301;
  assign \new_[3992]_  = \new_[3991]_  & \new_[3988]_ ;
  assign \new_[3995]_  = A199 & A169;
  assign \new_[3998]_  = A265 & A201;
  assign \new_[3999]_  = \new_[3998]_  & \new_[3995]_ ;
  assign \new_[4002]_  = ~A298 & A267;
  assign \new_[4005]_  = ~A301 & ~A299;
  assign \new_[4006]_  = \new_[4005]_  & \new_[4002]_ ;
  assign \new_[4009]_  = A199 & A169;
  assign \new_[4012]_  = A266 & A201;
  assign \new_[4013]_  = \new_[4012]_  & \new_[4009]_ ;
  assign \new_[4016]_  = ~A300 & A267;
  assign \new_[4019]_  = ~A302 & ~A301;
  assign \new_[4020]_  = \new_[4019]_  & \new_[4016]_ ;
  assign \new_[4023]_  = A199 & A169;
  assign \new_[4026]_  = A266 & A201;
  assign \new_[4027]_  = \new_[4026]_  & \new_[4023]_ ;
  assign \new_[4030]_  = ~A298 & A267;
  assign \new_[4033]_  = ~A301 & ~A299;
  assign \new_[4034]_  = \new_[4033]_  & \new_[4030]_ ;
  assign \new_[4037]_  = A200 & A169;
  assign \new_[4040]_  = A268 & A201;
  assign \new_[4041]_  = \new_[4040]_  & \new_[4037]_ ;
  assign \new_[4044]_  = A299 & A298;
  assign \new_[4047]_  = ~A301 & ~A300;
  assign \new_[4048]_  = \new_[4047]_  & \new_[4044]_ ;
  assign \new_[4051]_  = A200 & A169;
  assign \new_[4054]_  = A265 & A201;
  assign \new_[4055]_  = \new_[4054]_  & \new_[4051]_ ;
  assign \new_[4058]_  = ~A300 & A267;
  assign \new_[4061]_  = ~A302 & ~A301;
  assign \new_[4062]_  = \new_[4061]_  & \new_[4058]_ ;
  assign \new_[4065]_  = A200 & A169;
  assign \new_[4068]_  = A265 & A201;
  assign \new_[4069]_  = \new_[4068]_  & \new_[4065]_ ;
  assign \new_[4072]_  = ~A298 & A267;
  assign \new_[4075]_  = ~A301 & ~A299;
  assign \new_[4076]_  = \new_[4075]_  & \new_[4072]_ ;
  assign \new_[4079]_  = A200 & A169;
  assign \new_[4082]_  = A266 & A201;
  assign \new_[4083]_  = \new_[4082]_  & \new_[4079]_ ;
  assign \new_[4086]_  = ~A300 & A267;
  assign \new_[4089]_  = ~A302 & ~A301;
  assign \new_[4090]_  = \new_[4089]_  & \new_[4086]_ ;
  assign \new_[4093]_  = A200 & A169;
  assign \new_[4096]_  = A266 & A201;
  assign \new_[4097]_  = \new_[4096]_  & \new_[4093]_ ;
  assign \new_[4100]_  = ~A298 & A267;
  assign \new_[4103]_  = ~A301 & ~A299;
  assign \new_[4104]_  = \new_[4103]_  & \new_[4100]_ ;
  assign \new_[4107]_  = ~A199 & A169;
  assign \new_[4110]_  = A203 & A200;
  assign \new_[4111]_  = \new_[4110]_  & \new_[4107]_ ;
  assign \new_[4114]_  = ~A300 & A268;
  assign \new_[4117]_  = ~A302 & ~A301;
  assign \new_[4118]_  = \new_[4117]_  & \new_[4114]_ ;
  assign \new_[4121]_  = ~A199 & A169;
  assign \new_[4124]_  = A203 & A200;
  assign \new_[4125]_  = \new_[4124]_  & \new_[4121]_ ;
  assign \new_[4128]_  = ~A298 & A268;
  assign \new_[4131]_  = ~A301 & ~A299;
  assign \new_[4132]_  = \new_[4131]_  & \new_[4128]_ ;
  assign \new_[4135]_  = A199 & A169;
  assign \new_[4138]_  = A203 & ~A200;
  assign \new_[4139]_  = \new_[4138]_  & \new_[4135]_ ;
  assign \new_[4142]_  = ~A300 & A268;
  assign \new_[4145]_  = ~A302 & ~A301;
  assign \new_[4146]_  = \new_[4145]_  & \new_[4142]_ ;
  assign \new_[4149]_  = A199 & A169;
  assign \new_[4152]_  = A203 & ~A200;
  assign \new_[4153]_  = \new_[4152]_  & \new_[4149]_ ;
  assign \new_[4156]_  = ~A298 & A268;
  assign \new_[4159]_  = ~A301 & ~A299;
  assign \new_[4160]_  = \new_[4159]_  & \new_[4156]_ ;
  assign \new_[4163]_  = ~A199 & A169;
  assign \new_[4166]_  = ~A202 & ~A200;
  assign \new_[4167]_  = \new_[4166]_  & \new_[4163]_ ;
  assign \new_[4170]_  = ~A268 & ~A267;
  assign \new_[4173]_  = A301 & ~A269;
  assign \new_[4174]_  = \new_[4173]_  & \new_[4170]_ ;
  assign \new_[4177]_  = ~A199 & A169;
  assign \new_[4180]_  = ~A202 & ~A200;
  assign \new_[4181]_  = \new_[4180]_  & \new_[4177]_ ;
  assign \new_[4184]_  = ~A266 & ~A265;
  assign \new_[4187]_  = A301 & ~A268;
  assign \new_[4188]_  = \new_[4187]_  & \new_[4184]_ ;
  assign \new_[4191]_  = ~A167 & ~A169;
  assign \new_[4194]_  = A202 & ~A166;
  assign \new_[4195]_  = \new_[4194]_  & \new_[4191]_ ;
  assign \new_[4198]_  = ~A268 & ~A267;
  assign \new_[4201]_  = A301 & ~A269;
  assign \new_[4202]_  = \new_[4201]_  & \new_[4198]_ ;
  assign \new_[4205]_  = ~A167 & ~A169;
  assign \new_[4208]_  = A202 & ~A166;
  assign \new_[4209]_  = \new_[4208]_  & \new_[4205]_ ;
  assign \new_[4212]_  = ~A266 & ~A265;
  assign \new_[4215]_  = A301 & ~A268;
  assign \new_[4216]_  = \new_[4215]_  & \new_[4212]_ ;
  assign \new_[4219]_  = ~A169 & ~A170;
  assign \new_[4222]_  = A202 & ~A168;
  assign \new_[4223]_  = \new_[4222]_  & \new_[4219]_ ;
  assign \new_[4226]_  = ~A268 & ~A267;
  assign \new_[4229]_  = A301 & ~A269;
  assign \new_[4230]_  = \new_[4229]_  & \new_[4226]_ ;
  assign \new_[4233]_  = ~A169 & ~A170;
  assign \new_[4236]_  = A202 & ~A168;
  assign \new_[4237]_  = \new_[4236]_  & \new_[4233]_ ;
  assign \new_[4240]_  = ~A266 & ~A265;
  assign \new_[4243]_  = A301 & ~A268;
  assign \new_[4244]_  = \new_[4243]_  & \new_[4240]_ ;
  assign \new_[4247]_  = A166 & A168;
  assign \new_[4250]_  = A265 & A202;
  assign \new_[4251]_  = \new_[4250]_  & \new_[4247]_ ;
  assign \new_[4254]_  = A298 & A267;
  assign \new_[4258]_  = ~A301 & ~A300;
  assign \new_[4259]_  = A299 & \new_[4258]_ ;
  assign \new_[4260]_  = \new_[4259]_  & \new_[4254]_ ;
  assign \new_[4263]_  = A166 & A168;
  assign \new_[4266]_  = A266 & A202;
  assign \new_[4267]_  = \new_[4266]_  & \new_[4263]_ ;
  assign \new_[4270]_  = A298 & A267;
  assign \new_[4274]_  = ~A301 & ~A300;
  assign \new_[4275]_  = A299 & \new_[4274]_ ;
  assign \new_[4276]_  = \new_[4275]_  & \new_[4270]_ ;
  assign \new_[4279]_  = A166 & A168;
  assign \new_[4282]_  = ~A265 & A202;
  assign \new_[4283]_  = \new_[4282]_  & \new_[4279]_ ;
  assign \new_[4286]_  = A269 & A266;
  assign \new_[4290]_  = ~A302 & ~A301;
  assign \new_[4291]_  = ~A300 & \new_[4290]_ ;
  assign \new_[4292]_  = \new_[4291]_  & \new_[4286]_ ;
  assign \new_[4295]_  = A166 & A168;
  assign \new_[4298]_  = ~A265 & A202;
  assign \new_[4299]_  = \new_[4298]_  & \new_[4295]_ ;
  assign \new_[4302]_  = A269 & A266;
  assign \new_[4306]_  = ~A301 & ~A299;
  assign \new_[4307]_  = ~A298 & \new_[4306]_ ;
  assign \new_[4308]_  = \new_[4307]_  & \new_[4302]_ ;
  assign \new_[4311]_  = A166 & A168;
  assign \new_[4314]_  = A265 & A202;
  assign \new_[4315]_  = \new_[4314]_  & \new_[4311]_ ;
  assign \new_[4318]_  = A269 & ~A266;
  assign \new_[4322]_  = ~A302 & ~A301;
  assign \new_[4323]_  = ~A300 & \new_[4322]_ ;
  assign \new_[4324]_  = \new_[4323]_  & \new_[4318]_ ;
  assign \new_[4327]_  = A166 & A168;
  assign \new_[4330]_  = A265 & A202;
  assign \new_[4331]_  = \new_[4330]_  & \new_[4327]_ ;
  assign \new_[4334]_  = A269 & ~A266;
  assign \new_[4338]_  = ~A301 & ~A299;
  assign \new_[4339]_  = ~A298 & \new_[4338]_ ;
  assign \new_[4340]_  = \new_[4339]_  & \new_[4334]_ ;
  assign \new_[4343]_  = A166 & A168;
  assign \new_[4346]_  = ~A202 & ~A201;
  assign \new_[4347]_  = \new_[4346]_  & \new_[4343]_ ;
  assign \new_[4350]_  = ~A267 & ~A203;
  assign \new_[4354]_  = A301 & ~A269;
  assign \new_[4355]_  = ~A268 & \new_[4354]_ ;
  assign \new_[4356]_  = \new_[4355]_  & \new_[4350]_ ;
  assign \new_[4359]_  = A166 & A168;
  assign \new_[4362]_  = ~A202 & ~A201;
  assign \new_[4363]_  = \new_[4362]_  & \new_[4359]_ ;
  assign \new_[4366]_  = ~A265 & ~A203;
  assign \new_[4370]_  = A301 & ~A268;
  assign \new_[4371]_  = ~A266 & \new_[4370]_ ;
  assign \new_[4372]_  = \new_[4371]_  & \new_[4366]_ ;
  assign \new_[4375]_  = A166 & A168;
  assign \new_[4378]_  = A201 & A199;
  assign \new_[4379]_  = \new_[4378]_  & \new_[4375]_ ;
  assign \new_[4382]_  = A298 & A268;
  assign \new_[4386]_  = ~A301 & ~A300;
  assign \new_[4387]_  = A299 & \new_[4386]_ ;
  assign \new_[4388]_  = \new_[4387]_  & \new_[4382]_ ;
  assign \new_[4391]_  = A166 & A168;
  assign \new_[4394]_  = A201 & A199;
  assign \new_[4395]_  = \new_[4394]_  & \new_[4391]_ ;
  assign \new_[4398]_  = A267 & A265;
  assign \new_[4402]_  = ~A302 & ~A301;
  assign \new_[4403]_  = ~A300 & \new_[4402]_ ;
  assign \new_[4404]_  = \new_[4403]_  & \new_[4398]_ ;
  assign \new_[4407]_  = A166 & A168;
  assign \new_[4410]_  = A201 & A199;
  assign \new_[4411]_  = \new_[4410]_  & \new_[4407]_ ;
  assign \new_[4414]_  = A267 & A265;
  assign \new_[4418]_  = ~A301 & ~A299;
  assign \new_[4419]_  = ~A298 & \new_[4418]_ ;
  assign \new_[4420]_  = \new_[4419]_  & \new_[4414]_ ;
  assign \new_[4423]_  = A166 & A168;
  assign \new_[4426]_  = A201 & A199;
  assign \new_[4427]_  = \new_[4426]_  & \new_[4423]_ ;
  assign \new_[4430]_  = A267 & A266;
  assign \new_[4434]_  = ~A302 & ~A301;
  assign \new_[4435]_  = ~A300 & \new_[4434]_ ;
  assign \new_[4436]_  = \new_[4435]_  & \new_[4430]_ ;
  assign \new_[4439]_  = A166 & A168;
  assign \new_[4442]_  = A201 & A199;
  assign \new_[4443]_  = \new_[4442]_  & \new_[4439]_ ;
  assign \new_[4446]_  = A267 & A266;
  assign \new_[4450]_  = ~A301 & ~A299;
  assign \new_[4451]_  = ~A298 & \new_[4450]_ ;
  assign \new_[4452]_  = \new_[4451]_  & \new_[4446]_ ;
  assign \new_[4455]_  = A166 & A168;
  assign \new_[4458]_  = A201 & A200;
  assign \new_[4459]_  = \new_[4458]_  & \new_[4455]_ ;
  assign \new_[4462]_  = A298 & A268;
  assign \new_[4466]_  = ~A301 & ~A300;
  assign \new_[4467]_  = A299 & \new_[4466]_ ;
  assign \new_[4468]_  = \new_[4467]_  & \new_[4462]_ ;
  assign \new_[4471]_  = A166 & A168;
  assign \new_[4474]_  = A201 & A200;
  assign \new_[4475]_  = \new_[4474]_  & \new_[4471]_ ;
  assign \new_[4478]_  = A267 & A265;
  assign \new_[4482]_  = ~A302 & ~A301;
  assign \new_[4483]_  = ~A300 & \new_[4482]_ ;
  assign \new_[4484]_  = \new_[4483]_  & \new_[4478]_ ;
  assign \new_[4487]_  = A166 & A168;
  assign \new_[4490]_  = A201 & A200;
  assign \new_[4491]_  = \new_[4490]_  & \new_[4487]_ ;
  assign \new_[4494]_  = A267 & A265;
  assign \new_[4498]_  = ~A301 & ~A299;
  assign \new_[4499]_  = ~A298 & \new_[4498]_ ;
  assign \new_[4500]_  = \new_[4499]_  & \new_[4494]_ ;
  assign \new_[4503]_  = A166 & A168;
  assign \new_[4506]_  = A201 & A200;
  assign \new_[4507]_  = \new_[4506]_  & \new_[4503]_ ;
  assign \new_[4510]_  = A267 & A266;
  assign \new_[4514]_  = ~A302 & ~A301;
  assign \new_[4515]_  = ~A300 & \new_[4514]_ ;
  assign \new_[4516]_  = \new_[4515]_  & \new_[4510]_ ;
  assign \new_[4519]_  = A166 & A168;
  assign \new_[4522]_  = A201 & A200;
  assign \new_[4523]_  = \new_[4522]_  & \new_[4519]_ ;
  assign \new_[4526]_  = A267 & A266;
  assign \new_[4530]_  = ~A301 & ~A299;
  assign \new_[4531]_  = ~A298 & \new_[4530]_ ;
  assign \new_[4532]_  = \new_[4531]_  & \new_[4526]_ ;
  assign \new_[4535]_  = A166 & A168;
  assign \new_[4538]_  = A200 & ~A199;
  assign \new_[4539]_  = \new_[4538]_  & \new_[4535]_ ;
  assign \new_[4542]_  = A268 & A203;
  assign \new_[4546]_  = ~A302 & ~A301;
  assign \new_[4547]_  = ~A300 & \new_[4546]_ ;
  assign \new_[4548]_  = \new_[4547]_  & \new_[4542]_ ;
  assign \new_[4551]_  = A166 & A168;
  assign \new_[4554]_  = A200 & ~A199;
  assign \new_[4555]_  = \new_[4554]_  & \new_[4551]_ ;
  assign \new_[4558]_  = A268 & A203;
  assign \new_[4562]_  = ~A301 & ~A299;
  assign \new_[4563]_  = ~A298 & \new_[4562]_ ;
  assign \new_[4564]_  = \new_[4563]_  & \new_[4558]_ ;
  assign \new_[4567]_  = A166 & A168;
  assign \new_[4570]_  = ~A200 & A199;
  assign \new_[4571]_  = \new_[4570]_  & \new_[4567]_ ;
  assign \new_[4574]_  = A268 & A203;
  assign \new_[4578]_  = ~A302 & ~A301;
  assign \new_[4579]_  = ~A300 & \new_[4578]_ ;
  assign \new_[4580]_  = \new_[4579]_  & \new_[4574]_ ;
  assign \new_[4583]_  = A166 & A168;
  assign \new_[4586]_  = ~A200 & A199;
  assign \new_[4587]_  = \new_[4586]_  & \new_[4583]_ ;
  assign \new_[4590]_  = A268 & A203;
  assign \new_[4594]_  = ~A301 & ~A299;
  assign \new_[4595]_  = ~A298 & \new_[4594]_ ;
  assign \new_[4596]_  = \new_[4595]_  & \new_[4590]_ ;
  assign \new_[4599]_  = A166 & A168;
  assign \new_[4602]_  = ~A200 & ~A199;
  assign \new_[4603]_  = \new_[4602]_  & \new_[4599]_ ;
  assign \new_[4606]_  = ~A267 & ~A202;
  assign \new_[4610]_  = A301 & ~A269;
  assign \new_[4611]_  = ~A268 & \new_[4610]_ ;
  assign \new_[4612]_  = \new_[4611]_  & \new_[4606]_ ;
  assign \new_[4615]_  = A166 & A168;
  assign \new_[4618]_  = ~A200 & ~A199;
  assign \new_[4619]_  = \new_[4618]_  & \new_[4615]_ ;
  assign \new_[4622]_  = ~A265 & ~A202;
  assign \new_[4626]_  = A301 & ~A268;
  assign \new_[4627]_  = ~A266 & \new_[4626]_ ;
  assign \new_[4628]_  = \new_[4627]_  & \new_[4622]_ ;
  assign \new_[4631]_  = A167 & A168;
  assign \new_[4634]_  = A265 & A202;
  assign \new_[4635]_  = \new_[4634]_  & \new_[4631]_ ;
  assign \new_[4638]_  = A298 & A267;
  assign \new_[4642]_  = ~A301 & ~A300;
  assign \new_[4643]_  = A299 & \new_[4642]_ ;
  assign \new_[4644]_  = \new_[4643]_  & \new_[4638]_ ;
  assign \new_[4647]_  = A167 & A168;
  assign \new_[4650]_  = A266 & A202;
  assign \new_[4651]_  = \new_[4650]_  & \new_[4647]_ ;
  assign \new_[4654]_  = A298 & A267;
  assign \new_[4658]_  = ~A301 & ~A300;
  assign \new_[4659]_  = A299 & \new_[4658]_ ;
  assign \new_[4660]_  = \new_[4659]_  & \new_[4654]_ ;
  assign \new_[4663]_  = A167 & A168;
  assign \new_[4666]_  = ~A265 & A202;
  assign \new_[4667]_  = \new_[4666]_  & \new_[4663]_ ;
  assign \new_[4670]_  = A269 & A266;
  assign \new_[4674]_  = ~A302 & ~A301;
  assign \new_[4675]_  = ~A300 & \new_[4674]_ ;
  assign \new_[4676]_  = \new_[4675]_  & \new_[4670]_ ;
  assign \new_[4679]_  = A167 & A168;
  assign \new_[4682]_  = ~A265 & A202;
  assign \new_[4683]_  = \new_[4682]_  & \new_[4679]_ ;
  assign \new_[4686]_  = A269 & A266;
  assign \new_[4690]_  = ~A301 & ~A299;
  assign \new_[4691]_  = ~A298 & \new_[4690]_ ;
  assign \new_[4692]_  = \new_[4691]_  & \new_[4686]_ ;
  assign \new_[4695]_  = A167 & A168;
  assign \new_[4698]_  = A265 & A202;
  assign \new_[4699]_  = \new_[4698]_  & \new_[4695]_ ;
  assign \new_[4702]_  = A269 & ~A266;
  assign \new_[4706]_  = ~A302 & ~A301;
  assign \new_[4707]_  = ~A300 & \new_[4706]_ ;
  assign \new_[4708]_  = \new_[4707]_  & \new_[4702]_ ;
  assign \new_[4711]_  = A167 & A168;
  assign \new_[4714]_  = A265 & A202;
  assign \new_[4715]_  = \new_[4714]_  & \new_[4711]_ ;
  assign \new_[4718]_  = A269 & ~A266;
  assign \new_[4722]_  = ~A301 & ~A299;
  assign \new_[4723]_  = ~A298 & \new_[4722]_ ;
  assign \new_[4724]_  = \new_[4723]_  & \new_[4718]_ ;
  assign \new_[4727]_  = A167 & A168;
  assign \new_[4730]_  = ~A202 & ~A201;
  assign \new_[4731]_  = \new_[4730]_  & \new_[4727]_ ;
  assign \new_[4734]_  = ~A267 & ~A203;
  assign \new_[4738]_  = A301 & ~A269;
  assign \new_[4739]_  = ~A268 & \new_[4738]_ ;
  assign \new_[4740]_  = \new_[4739]_  & \new_[4734]_ ;
  assign \new_[4743]_  = A167 & A168;
  assign \new_[4746]_  = ~A202 & ~A201;
  assign \new_[4747]_  = \new_[4746]_  & \new_[4743]_ ;
  assign \new_[4750]_  = ~A265 & ~A203;
  assign \new_[4754]_  = A301 & ~A268;
  assign \new_[4755]_  = ~A266 & \new_[4754]_ ;
  assign \new_[4756]_  = \new_[4755]_  & \new_[4750]_ ;
  assign \new_[4759]_  = A167 & A168;
  assign \new_[4762]_  = A201 & A199;
  assign \new_[4763]_  = \new_[4762]_  & \new_[4759]_ ;
  assign \new_[4766]_  = A298 & A268;
  assign \new_[4770]_  = ~A301 & ~A300;
  assign \new_[4771]_  = A299 & \new_[4770]_ ;
  assign \new_[4772]_  = \new_[4771]_  & \new_[4766]_ ;
  assign \new_[4775]_  = A167 & A168;
  assign \new_[4778]_  = A201 & A199;
  assign \new_[4779]_  = \new_[4778]_  & \new_[4775]_ ;
  assign \new_[4782]_  = A267 & A265;
  assign \new_[4786]_  = ~A302 & ~A301;
  assign \new_[4787]_  = ~A300 & \new_[4786]_ ;
  assign \new_[4788]_  = \new_[4787]_  & \new_[4782]_ ;
  assign \new_[4791]_  = A167 & A168;
  assign \new_[4794]_  = A201 & A199;
  assign \new_[4795]_  = \new_[4794]_  & \new_[4791]_ ;
  assign \new_[4798]_  = A267 & A265;
  assign \new_[4802]_  = ~A301 & ~A299;
  assign \new_[4803]_  = ~A298 & \new_[4802]_ ;
  assign \new_[4804]_  = \new_[4803]_  & \new_[4798]_ ;
  assign \new_[4807]_  = A167 & A168;
  assign \new_[4810]_  = A201 & A199;
  assign \new_[4811]_  = \new_[4810]_  & \new_[4807]_ ;
  assign \new_[4814]_  = A267 & A266;
  assign \new_[4818]_  = ~A302 & ~A301;
  assign \new_[4819]_  = ~A300 & \new_[4818]_ ;
  assign \new_[4820]_  = \new_[4819]_  & \new_[4814]_ ;
  assign \new_[4823]_  = A167 & A168;
  assign \new_[4826]_  = A201 & A199;
  assign \new_[4827]_  = \new_[4826]_  & \new_[4823]_ ;
  assign \new_[4830]_  = A267 & A266;
  assign \new_[4834]_  = ~A301 & ~A299;
  assign \new_[4835]_  = ~A298 & \new_[4834]_ ;
  assign \new_[4836]_  = \new_[4835]_  & \new_[4830]_ ;
  assign \new_[4839]_  = A167 & A168;
  assign \new_[4842]_  = A201 & A200;
  assign \new_[4843]_  = \new_[4842]_  & \new_[4839]_ ;
  assign \new_[4846]_  = A298 & A268;
  assign \new_[4850]_  = ~A301 & ~A300;
  assign \new_[4851]_  = A299 & \new_[4850]_ ;
  assign \new_[4852]_  = \new_[4851]_  & \new_[4846]_ ;
  assign \new_[4855]_  = A167 & A168;
  assign \new_[4858]_  = A201 & A200;
  assign \new_[4859]_  = \new_[4858]_  & \new_[4855]_ ;
  assign \new_[4862]_  = A267 & A265;
  assign \new_[4866]_  = ~A302 & ~A301;
  assign \new_[4867]_  = ~A300 & \new_[4866]_ ;
  assign \new_[4868]_  = \new_[4867]_  & \new_[4862]_ ;
  assign \new_[4871]_  = A167 & A168;
  assign \new_[4874]_  = A201 & A200;
  assign \new_[4875]_  = \new_[4874]_  & \new_[4871]_ ;
  assign \new_[4878]_  = A267 & A265;
  assign \new_[4882]_  = ~A301 & ~A299;
  assign \new_[4883]_  = ~A298 & \new_[4882]_ ;
  assign \new_[4884]_  = \new_[4883]_  & \new_[4878]_ ;
  assign \new_[4887]_  = A167 & A168;
  assign \new_[4890]_  = A201 & A200;
  assign \new_[4891]_  = \new_[4890]_  & \new_[4887]_ ;
  assign \new_[4894]_  = A267 & A266;
  assign \new_[4898]_  = ~A302 & ~A301;
  assign \new_[4899]_  = ~A300 & \new_[4898]_ ;
  assign \new_[4900]_  = \new_[4899]_  & \new_[4894]_ ;
  assign \new_[4903]_  = A167 & A168;
  assign \new_[4906]_  = A201 & A200;
  assign \new_[4907]_  = \new_[4906]_  & \new_[4903]_ ;
  assign \new_[4910]_  = A267 & A266;
  assign \new_[4914]_  = ~A301 & ~A299;
  assign \new_[4915]_  = ~A298 & \new_[4914]_ ;
  assign \new_[4916]_  = \new_[4915]_  & \new_[4910]_ ;
  assign \new_[4919]_  = A167 & A168;
  assign \new_[4922]_  = A200 & ~A199;
  assign \new_[4923]_  = \new_[4922]_  & \new_[4919]_ ;
  assign \new_[4926]_  = A268 & A203;
  assign \new_[4930]_  = ~A302 & ~A301;
  assign \new_[4931]_  = ~A300 & \new_[4930]_ ;
  assign \new_[4932]_  = \new_[4931]_  & \new_[4926]_ ;
  assign \new_[4935]_  = A167 & A168;
  assign \new_[4938]_  = A200 & ~A199;
  assign \new_[4939]_  = \new_[4938]_  & \new_[4935]_ ;
  assign \new_[4942]_  = A268 & A203;
  assign \new_[4946]_  = ~A301 & ~A299;
  assign \new_[4947]_  = ~A298 & \new_[4946]_ ;
  assign \new_[4948]_  = \new_[4947]_  & \new_[4942]_ ;
  assign \new_[4951]_  = A167 & A168;
  assign \new_[4954]_  = ~A200 & A199;
  assign \new_[4955]_  = \new_[4954]_  & \new_[4951]_ ;
  assign \new_[4958]_  = A268 & A203;
  assign \new_[4962]_  = ~A302 & ~A301;
  assign \new_[4963]_  = ~A300 & \new_[4962]_ ;
  assign \new_[4964]_  = \new_[4963]_  & \new_[4958]_ ;
  assign \new_[4967]_  = A167 & A168;
  assign \new_[4970]_  = ~A200 & A199;
  assign \new_[4971]_  = \new_[4970]_  & \new_[4967]_ ;
  assign \new_[4974]_  = A268 & A203;
  assign \new_[4978]_  = ~A301 & ~A299;
  assign \new_[4979]_  = ~A298 & \new_[4978]_ ;
  assign \new_[4980]_  = \new_[4979]_  & \new_[4974]_ ;
  assign \new_[4983]_  = A167 & A168;
  assign \new_[4986]_  = ~A200 & ~A199;
  assign \new_[4987]_  = \new_[4986]_  & \new_[4983]_ ;
  assign \new_[4990]_  = ~A267 & ~A202;
  assign \new_[4994]_  = A301 & ~A269;
  assign \new_[4995]_  = ~A268 & \new_[4994]_ ;
  assign \new_[4996]_  = \new_[4995]_  & \new_[4990]_ ;
  assign \new_[4999]_  = A167 & A168;
  assign \new_[5002]_  = ~A200 & ~A199;
  assign \new_[5003]_  = \new_[5002]_  & \new_[4999]_ ;
  assign \new_[5006]_  = ~A265 & ~A202;
  assign \new_[5010]_  = A301 & ~A268;
  assign \new_[5011]_  = ~A266 & \new_[5010]_ ;
  assign \new_[5012]_  = \new_[5011]_  & \new_[5006]_ ;
  assign \new_[5015]_  = A167 & A170;
  assign \new_[5018]_  = A202 & ~A166;
  assign \new_[5019]_  = \new_[5018]_  & \new_[5015]_ ;
  assign \new_[5022]_  = A298 & A268;
  assign \new_[5026]_  = ~A301 & ~A300;
  assign \new_[5027]_  = A299 & \new_[5026]_ ;
  assign \new_[5028]_  = \new_[5027]_  & \new_[5022]_ ;
  assign \new_[5031]_  = A167 & A170;
  assign \new_[5034]_  = A202 & ~A166;
  assign \new_[5035]_  = \new_[5034]_  & \new_[5031]_ ;
  assign \new_[5038]_  = A267 & A265;
  assign \new_[5042]_  = ~A302 & ~A301;
  assign \new_[5043]_  = ~A300 & \new_[5042]_ ;
  assign \new_[5044]_  = \new_[5043]_  & \new_[5038]_ ;
  assign \new_[5047]_  = A167 & A170;
  assign \new_[5050]_  = A202 & ~A166;
  assign \new_[5051]_  = \new_[5050]_  & \new_[5047]_ ;
  assign \new_[5054]_  = A267 & A265;
  assign \new_[5058]_  = ~A301 & ~A299;
  assign \new_[5059]_  = ~A298 & \new_[5058]_ ;
  assign \new_[5060]_  = \new_[5059]_  & \new_[5054]_ ;
  assign \new_[5063]_  = A167 & A170;
  assign \new_[5066]_  = A202 & ~A166;
  assign \new_[5067]_  = \new_[5066]_  & \new_[5063]_ ;
  assign \new_[5070]_  = A267 & A266;
  assign \new_[5074]_  = ~A302 & ~A301;
  assign \new_[5075]_  = ~A300 & \new_[5074]_ ;
  assign \new_[5076]_  = \new_[5075]_  & \new_[5070]_ ;
  assign \new_[5079]_  = A167 & A170;
  assign \new_[5082]_  = A202 & ~A166;
  assign \new_[5083]_  = \new_[5082]_  & \new_[5079]_ ;
  assign \new_[5086]_  = A267 & A266;
  assign \new_[5090]_  = ~A301 & ~A299;
  assign \new_[5091]_  = ~A298 & \new_[5090]_ ;
  assign \new_[5092]_  = \new_[5091]_  & \new_[5086]_ ;
  assign \new_[5095]_  = A167 & A170;
  assign \new_[5098]_  = A199 & ~A166;
  assign \new_[5099]_  = \new_[5098]_  & \new_[5095]_ ;
  assign \new_[5102]_  = A268 & A201;
  assign \new_[5106]_  = ~A302 & ~A301;
  assign \new_[5107]_  = ~A300 & \new_[5106]_ ;
  assign \new_[5108]_  = \new_[5107]_  & \new_[5102]_ ;
  assign \new_[5111]_  = A167 & A170;
  assign \new_[5114]_  = A199 & ~A166;
  assign \new_[5115]_  = \new_[5114]_  & \new_[5111]_ ;
  assign \new_[5118]_  = A268 & A201;
  assign \new_[5122]_  = ~A301 & ~A299;
  assign \new_[5123]_  = ~A298 & \new_[5122]_ ;
  assign \new_[5124]_  = \new_[5123]_  & \new_[5118]_ ;
  assign \new_[5127]_  = A167 & A170;
  assign \new_[5130]_  = A200 & ~A166;
  assign \new_[5131]_  = \new_[5130]_  & \new_[5127]_ ;
  assign \new_[5134]_  = A268 & A201;
  assign \new_[5138]_  = ~A302 & ~A301;
  assign \new_[5139]_  = ~A300 & \new_[5138]_ ;
  assign \new_[5140]_  = \new_[5139]_  & \new_[5134]_ ;
  assign \new_[5143]_  = A167 & A170;
  assign \new_[5146]_  = A200 & ~A166;
  assign \new_[5147]_  = \new_[5146]_  & \new_[5143]_ ;
  assign \new_[5150]_  = A268 & A201;
  assign \new_[5154]_  = ~A301 & ~A299;
  assign \new_[5155]_  = ~A298 & \new_[5154]_ ;
  assign \new_[5156]_  = \new_[5155]_  & \new_[5150]_ ;
  assign \new_[5159]_  = ~A167 & A170;
  assign \new_[5162]_  = A202 & A166;
  assign \new_[5163]_  = \new_[5162]_  & \new_[5159]_ ;
  assign \new_[5166]_  = A298 & A268;
  assign \new_[5170]_  = ~A301 & ~A300;
  assign \new_[5171]_  = A299 & \new_[5170]_ ;
  assign \new_[5172]_  = \new_[5171]_  & \new_[5166]_ ;
  assign \new_[5175]_  = ~A167 & A170;
  assign \new_[5178]_  = A202 & A166;
  assign \new_[5179]_  = \new_[5178]_  & \new_[5175]_ ;
  assign \new_[5182]_  = A267 & A265;
  assign \new_[5186]_  = ~A302 & ~A301;
  assign \new_[5187]_  = ~A300 & \new_[5186]_ ;
  assign \new_[5188]_  = \new_[5187]_  & \new_[5182]_ ;
  assign \new_[5191]_  = ~A167 & A170;
  assign \new_[5194]_  = A202 & A166;
  assign \new_[5195]_  = \new_[5194]_  & \new_[5191]_ ;
  assign \new_[5198]_  = A267 & A265;
  assign \new_[5202]_  = ~A301 & ~A299;
  assign \new_[5203]_  = ~A298 & \new_[5202]_ ;
  assign \new_[5204]_  = \new_[5203]_  & \new_[5198]_ ;
  assign \new_[5207]_  = ~A167 & A170;
  assign \new_[5210]_  = A202 & A166;
  assign \new_[5211]_  = \new_[5210]_  & \new_[5207]_ ;
  assign \new_[5214]_  = A267 & A266;
  assign \new_[5218]_  = ~A302 & ~A301;
  assign \new_[5219]_  = ~A300 & \new_[5218]_ ;
  assign \new_[5220]_  = \new_[5219]_  & \new_[5214]_ ;
  assign \new_[5223]_  = ~A167 & A170;
  assign \new_[5226]_  = A202 & A166;
  assign \new_[5227]_  = \new_[5226]_  & \new_[5223]_ ;
  assign \new_[5230]_  = A267 & A266;
  assign \new_[5234]_  = ~A301 & ~A299;
  assign \new_[5235]_  = ~A298 & \new_[5234]_ ;
  assign \new_[5236]_  = \new_[5235]_  & \new_[5230]_ ;
  assign \new_[5239]_  = ~A167 & A170;
  assign \new_[5242]_  = A199 & A166;
  assign \new_[5243]_  = \new_[5242]_  & \new_[5239]_ ;
  assign \new_[5246]_  = A268 & A201;
  assign \new_[5250]_  = ~A302 & ~A301;
  assign \new_[5251]_  = ~A300 & \new_[5250]_ ;
  assign \new_[5252]_  = \new_[5251]_  & \new_[5246]_ ;
  assign \new_[5255]_  = ~A167 & A170;
  assign \new_[5258]_  = A199 & A166;
  assign \new_[5259]_  = \new_[5258]_  & \new_[5255]_ ;
  assign \new_[5262]_  = A268 & A201;
  assign \new_[5266]_  = ~A301 & ~A299;
  assign \new_[5267]_  = ~A298 & \new_[5266]_ ;
  assign \new_[5268]_  = \new_[5267]_  & \new_[5262]_ ;
  assign \new_[5271]_  = ~A167 & A170;
  assign \new_[5274]_  = A200 & A166;
  assign \new_[5275]_  = \new_[5274]_  & \new_[5271]_ ;
  assign \new_[5278]_  = A268 & A201;
  assign \new_[5282]_  = ~A302 & ~A301;
  assign \new_[5283]_  = ~A300 & \new_[5282]_ ;
  assign \new_[5284]_  = \new_[5283]_  & \new_[5278]_ ;
  assign \new_[5287]_  = ~A167 & A170;
  assign \new_[5290]_  = A200 & A166;
  assign \new_[5291]_  = \new_[5290]_  & \new_[5287]_ ;
  assign \new_[5294]_  = A268 & A201;
  assign \new_[5298]_  = ~A301 & ~A299;
  assign \new_[5299]_  = ~A298 & \new_[5298]_ ;
  assign \new_[5300]_  = \new_[5299]_  & \new_[5294]_ ;
  assign \new_[5303]_  = A202 & A169;
  assign \new_[5306]_  = A266 & ~A265;
  assign \new_[5307]_  = \new_[5306]_  & \new_[5303]_ ;
  assign \new_[5310]_  = A298 & A269;
  assign \new_[5314]_  = ~A301 & ~A300;
  assign \new_[5315]_  = A299 & \new_[5314]_ ;
  assign \new_[5316]_  = \new_[5315]_  & \new_[5310]_ ;
  assign \new_[5319]_  = A202 & A169;
  assign \new_[5322]_  = ~A266 & A265;
  assign \new_[5323]_  = \new_[5322]_  & \new_[5319]_ ;
  assign \new_[5326]_  = A298 & A269;
  assign \new_[5330]_  = ~A301 & ~A300;
  assign \new_[5331]_  = A299 & \new_[5330]_ ;
  assign \new_[5332]_  = \new_[5331]_  & \new_[5326]_ ;
  assign \new_[5335]_  = ~A201 & A169;
  assign \new_[5338]_  = ~A203 & ~A202;
  assign \new_[5339]_  = \new_[5338]_  & \new_[5335]_ ;
  assign \new_[5342]_  = ~A268 & ~A267;
  assign \new_[5346]_  = A300 & A299;
  assign \new_[5347]_  = ~A269 & \new_[5346]_ ;
  assign \new_[5348]_  = \new_[5347]_  & \new_[5342]_ ;
  assign \new_[5351]_  = ~A201 & A169;
  assign \new_[5354]_  = ~A203 & ~A202;
  assign \new_[5355]_  = \new_[5354]_  & \new_[5351]_ ;
  assign \new_[5358]_  = ~A268 & ~A267;
  assign \new_[5362]_  = A300 & A298;
  assign \new_[5363]_  = ~A269 & \new_[5362]_ ;
  assign \new_[5364]_  = \new_[5363]_  & \new_[5358]_ ;
  assign \new_[5367]_  = ~A201 & A169;
  assign \new_[5370]_  = ~A203 & ~A202;
  assign \new_[5371]_  = \new_[5370]_  & \new_[5367]_ ;
  assign \new_[5374]_  = A266 & A265;
  assign \new_[5378]_  = A301 & ~A268;
  assign \new_[5379]_  = ~A267 & \new_[5378]_ ;
  assign \new_[5380]_  = \new_[5379]_  & \new_[5374]_ ;
  assign \new_[5383]_  = ~A201 & A169;
  assign \new_[5386]_  = ~A203 & ~A202;
  assign \new_[5387]_  = \new_[5386]_  & \new_[5383]_ ;
  assign \new_[5390]_  = ~A266 & ~A265;
  assign \new_[5394]_  = A300 & A299;
  assign \new_[5395]_  = ~A268 & \new_[5394]_ ;
  assign \new_[5396]_  = \new_[5395]_  & \new_[5390]_ ;
  assign \new_[5399]_  = ~A201 & A169;
  assign \new_[5402]_  = ~A203 & ~A202;
  assign \new_[5403]_  = \new_[5402]_  & \new_[5399]_ ;
  assign \new_[5406]_  = ~A266 & ~A265;
  assign \new_[5410]_  = A300 & A298;
  assign \new_[5411]_  = ~A268 & \new_[5410]_ ;
  assign \new_[5412]_  = \new_[5411]_  & \new_[5406]_ ;
  assign \new_[5415]_  = A199 & A169;
  assign \new_[5418]_  = A265 & A201;
  assign \new_[5419]_  = \new_[5418]_  & \new_[5415]_ ;
  assign \new_[5422]_  = A298 & A267;
  assign \new_[5426]_  = ~A301 & ~A300;
  assign \new_[5427]_  = A299 & \new_[5426]_ ;
  assign \new_[5428]_  = \new_[5427]_  & \new_[5422]_ ;
  assign \new_[5431]_  = A199 & A169;
  assign \new_[5434]_  = A266 & A201;
  assign \new_[5435]_  = \new_[5434]_  & \new_[5431]_ ;
  assign \new_[5438]_  = A298 & A267;
  assign \new_[5442]_  = ~A301 & ~A300;
  assign \new_[5443]_  = A299 & \new_[5442]_ ;
  assign \new_[5444]_  = \new_[5443]_  & \new_[5438]_ ;
  assign \new_[5447]_  = A199 & A169;
  assign \new_[5450]_  = ~A265 & A201;
  assign \new_[5451]_  = \new_[5450]_  & \new_[5447]_ ;
  assign \new_[5454]_  = A269 & A266;
  assign \new_[5458]_  = ~A302 & ~A301;
  assign \new_[5459]_  = ~A300 & \new_[5458]_ ;
  assign \new_[5460]_  = \new_[5459]_  & \new_[5454]_ ;
  assign \new_[5463]_  = A199 & A169;
  assign \new_[5466]_  = ~A265 & A201;
  assign \new_[5467]_  = \new_[5466]_  & \new_[5463]_ ;
  assign \new_[5470]_  = A269 & A266;
  assign \new_[5474]_  = ~A301 & ~A299;
  assign \new_[5475]_  = ~A298 & \new_[5474]_ ;
  assign \new_[5476]_  = \new_[5475]_  & \new_[5470]_ ;
  assign \new_[5479]_  = A199 & A169;
  assign \new_[5482]_  = A265 & A201;
  assign \new_[5483]_  = \new_[5482]_  & \new_[5479]_ ;
  assign \new_[5486]_  = A269 & ~A266;
  assign \new_[5490]_  = ~A302 & ~A301;
  assign \new_[5491]_  = ~A300 & \new_[5490]_ ;
  assign \new_[5492]_  = \new_[5491]_  & \new_[5486]_ ;
  assign \new_[5495]_  = A199 & A169;
  assign \new_[5498]_  = A265 & A201;
  assign \new_[5499]_  = \new_[5498]_  & \new_[5495]_ ;
  assign \new_[5502]_  = A269 & ~A266;
  assign \new_[5506]_  = ~A301 & ~A299;
  assign \new_[5507]_  = ~A298 & \new_[5506]_ ;
  assign \new_[5508]_  = \new_[5507]_  & \new_[5502]_ ;
  assign \new_[5511]_  = A200 & A169;
  assign \new_[5514]_  = A265 & A201;
  assign \new_[5515]_  = \new_[5514]_  & \new_[5511]_ ;
  assign \new_[5518]_  = A298 & A267;
  assign \new_[5522]_  = ~A301 & ~A300;
  assign \new_[5523]_  = A299 & \new_[5522]_ ;
  assign \new_[5524]_  = \new_[5523]_  & \new_[5518]_ ;
  assign \new_[5527]_  = A200 & A169;
  assign \new_[5530]_  = A266 & A201;
  assign \new_[5531]_  = \new_[5530]_  & \new_[5527]_ ;
  assign \new_[5534]_  = A298 & A267;
  assign \new_[5538]_  = ~A301 & ~A300;
  assign \new_[5539]_  = A299 & \new_[5538]_ ;
  assign \new_[5540]_  = \new_[5539]_  & \new_[5534]_ ;
  assign \new_[5543]_  = A200 & A169;
  assign \new_[5546]_  = ~A265 & A201;
  assign \new_[5547]_  = \new_[5546]_  & \new_[5543]_ ;
  assign \new_[5550]_  = A269 & A266;
  assign \new_[5554]_  = ~A302 & ~A301;
  assign \new_[5555]_  = ~A300 & \new_[5554]_ ;
  assign \new_[5556]_  = \new_[5555]_  & \new_[5550]_ ;
  assign \new_[5559]_  = A200 & A169;
  assign \new_[5562]_  = ~A265 & A201;
  assign \new_[5563]_  = \new_[5562]_  & \new_[5559]_ ;
  assign \new_[5566]_  = A269 & A266;
  assign \new_[5570]_  = ~A301 & ~A299;
  assign \new_[5571]_  = ~A298 & \new_[5570]_ ;
  assign \new_[5572]_  = \new_[5571]_  & \new_[5566]_ ;
  assign \new_[5575]_  = A200 & A169;
  assign \new_[5578]_  = A265 & A201;
  assign \new_[5579]_  = \new_[5578]_  & \new_[5575]_ ;
  assign \new_[5582]_  = A269 & ~A266;
  assign \new_[5586]_  = ~A302 & ~A301;
  assign \new_[5587]_  = ~A300 & \new_[5586]_ ;
  assign \new_[5588]_  = \new_[5587]_  & \new_[5582]_ ;
  assign \new_[5591]_  = A200 & A169;
  assign \new_[5594]_  = A265 & A201;
  assign \new_[5595]_  = \new_[5594]_  & \new_[5591]_ ;
  assign \new_[5598]_  = A269 & ~A266;
  assign \new_[5602]_  = ~A301 & ~A299;
  assign \new_[5603]_  = ~A298 & \new_[5602]_ ;
  assign \new_[5604]_  = \new_[5603]_  & \new_[5598]_ ;
  assign \new_[5607]_  = A199 & A169;
  assign \new_[5610]_  = ~A201 & A200;
  assign \new_[5611]_  = \new_[5610]_  & \new_[5607]_ ;
  assign \new_[5614]_  = ~A267 & ~A202;
  assign \new_[5618]_  = A301 & ~A269;
  assign \new_[5619]_  = ~A268 & \new_[5618]_ ;
  assign \new_[5620]_  = \new_[5619]_  & \new_[5614]_ ;
  assign \new_[5623]_  = A199 & A169;
  assign \new_[5626]_  = ~A201 & A200;
  assign \new_[5627]_  = \new_[5626]_  & \new_[5623]_ ;
  assign \new_[5630]_  = ~A265 & ~A202;
  assign \new_[5634]_  = A301 & ~A268;
  assign \new_[5635]_  = ~A266 & \new_[5634]_ ;
  assign \new_[5636]_  = \new_[5635]_  & \new_[5630]_ ;
  assign \new_[5639]_  = ~A199 & A169;
  assign \new_[5642]_  = A203 & A200;
  assign \new_[5643]_  = \new_[5642]_  & \new_[5639]_ ;
  assign \new_[5646]_  = A298 & A268;
  assign \new_[5650]_  = ~A301 & ~A300;
  assign \new_[5651]_  = A299 & \new_[5650]_ ;
  assign \new_[5652]_  = \new_[5651]_  & \new_[5646]_ ;
  assign \new_[5655]_  = ~A199 & A169;
  assign \new_[5658]_  = A203 & A200;
  assign \new_[5659]_  = \new_[5658]_  & \new_[5655]_ ;
  assign \new_[5662]_  = A267 & A265;
  assign \new_[5666]_  = ~A302 & ~A301;
  assign \new_[5667]_  = ~A300 & \new_[5666]_ ;
  assign \new_[5668]_  = \new_[5667]_  & \new_[5662]_ ;
  assign \new_[5671]_  = ~A199 & A169;
  assign \new_[5674]_  = A203 & A200;
  assign \new_[5675]_  = \new_[5674]_  & \new_[5671]_ ;
  assign \new_[5678]_  = A267 & A265;
  assign \new_[5682]_  = ~A301 & ~A299;
  assign \new_[5683]_  = ~A298 & \new_[5682]_ ;
  assign \new_[5684]_  = \new_[5683]_  & \new_[5678]_ ;
  assign \new_[5687]_  = ~A199 & A169;
  assign \new_[5690]_  = A203 & A200;
  assign \new_[5691]_  = \new_[5690]_  & \new_[5687]_ ;
  assign \new_[5694]_  = A267 & A266;
  assign \new_[5698]_  = ~A302 & ~A301;
  assign \new_[5699]_  = ~A300 & \new_[5698]_ ;
  assign \new_[5700]_  = \new_[5699]_  & \new_[5694]_ ;
  assign \new_[5703]_  = ~A199 & A169;
  assign \new_[5706]_  = A203 & A200;
  assign \new_[5707]_  = \new_[5706]_  & \new_[5703]_ ;
  assign \new_[5710]_  = A267 & A266;
  assign \new_[5714]_  = ~A301 & ~A299;
  assign \new_[5715]_  = ~A298 & \new_[5714]_ ;
  assign \new_[5716]_  = \new_[5715]_  & \new_[5710]_ ;
  assign \new_[5719]_  = A199 & A169;
  assign \new_[5722]_  = A203 & ~A200;
  assign \new_[5723]_  = \new_[5722]_  & \new_[5719]_ ;
  assign \new_[5726]_  = A298 & A268;
  assign \new_[5730]_  = ~A301 & ~A300;
  assign \new_[5731]_  = A299 & \new_[5730]_ ;
  assign \new_[5732]_  = \new_[5731]_  & \new_[5726]_ ;
  assign \new_[5735]_  = A199 & A169;
  assign \new_[5738]_  = A203 & ~A200;
  assign \new_[5739]_  = \new_[5738]_  & \new_[5735]_ ;
  assign \new_[5742]_  = A267 & A265;
  assign \new_[5746]_  = ~A302 & ~A301;
  assign \new_[5747]_  = ~A300 & \new_[5746]_ ;
  assign \new_[5748]_  = \new_[5747]_  & \new_[5742]_ ;
  assign \new_[5751]_  = A199 & A169;
  assign \new_[5754]_  = A203 & ~A200;
  assign \new_[5755]_  = \new_[5754]_  & \new_[5751]_ ;
  assign \new_[5758]_  = A267 & A265;
  assign \new_[5762]_  = ~A301 & ~A299;
  assign \new_[5763]_  = ~A298 & \new_[5762]_ ;
  assign \new_[5764]_  = \new_[5763]_  & \new_[5758]_ ;
  assign \new_[5767]_  = A199 & A169;
  assign \new_[5770]_  = A203 & ~A200;
  assign \new_[5771]_  = \new_[5770]_  & \new_[5767]_ ;
  assign \new_[5774]_  = A267 & A266;
  assign \new_[5778]_  = ~A302 & ~A301;
  assign \new_[5779]_  = ~A300 & \new_[5778]_ ;
  assign \new_[5780]_  = \new_[5779]_  & \new_[5774]_ ;
  assign \new_[5783]_  = A199 & A169;
  assign \new_[5786]_  = A203 & ~A200;
  assign \new_[5787]_  = \new_[5786]_  & \new_[5783]_ ;
  assign \new_[5790]_  = A267 & A266;
  assign \new_[5794]_  = ~A301 & ~A299;
  assign \new_[5795]_  = ~A298 & \new_[5794]_ ;
  assign \new_[5796]_  = \new_[5795]_  & \new_[5790]_ ;
  assign \new_[5799]_  = ~A199 & A169;
  assign \new_[5802]_  = ~A202 & ~A200;
  assign \new_[5803]_  = \new_[5802]_  & \new_[5799]_ ;
  assign \new_[5806]_  = ~A268 & ~A267;
  assign \new_[5810]_  = A300 & A299;
  assign \new_[5811]_  = ~A269 & \new_[5810]_ ;
  assign \new_[5812]_  = \new_[5811]_  & \new_[5806]_ ;
  assign \new_[5815]_  = ~A199 & A169;
  assign \new_[5818]_  = ~A202 & ~A200;
  assign \new_[5819]_  = \new_[5818]_  & \new_[5815]_ ;
  assign \new_[5822]_  = ~A268 & ~A267;
  assign \new_[5826]_  = A300 & A298;
  assign \new_[5827]_  = ~A269 & \new_[5826]_ ;
  assign \new_[5828]_  = \new_[5827]_  & \new_[5822]_ ;
  assign \new_[5831]_  = ~A199 & A169;
  assign \new_[5834]_  = ~A202 & ~A200;
  assign \new_[5835]_  = \new_[5834]_  & \new_[5831]_ ;
  assign \new_[5838]_  = A266 & A265;
  assign \new_[5842]_  = A301 & ~A268;
  assign \new_[5843]_  = ~A267 & \new_[5842]_ ;
  assign \new_[5844]_  = \new_[5843]_  & \new_[5838]_ ;
  assign \new_[5847]_  = ~A199 & A169;
  assign \new_[5850]_  = ~A202 & ~A200;
  assign \new_[5851]_  = \new_[5850]_  & \new_[5847]_ ;
  assign \new_[5854]_  = ~A266 & ~A265;
  assign \new_[5858]_  = A300 & A299;
  assign \new_[5859]_  = ~A268 & \new_[5858]_ ;
  assign \new_[5860]_  = \new_[5859]_  & \new_[5854]_ ;
  assign \new_[5863]_  = ~A199 & A169;
  assign \new_[5866]_  = ~A202 & ~A200;
  assign \new_[5867]_  = \new_[5866]_  & \new_[5863]_ ;
  assign \new_[5870]_  = ~A266 & ~A265;
  assign \new_[5874]_  = A300 & A298;
  assign \new_[5875]_  = ~A268 & \new_[5874]_ ;
  assign \new_[5876]_  = \new_[5875]_  & \new_[5870]_ ;
  assign \new_[5879]_  = ~A167 & ~A169;
  assign \new_[5882]_  = A202 & ~A166;
  assign \new_[5883]_  = \new_[5882]_  & \new_[5879]_ ;
  assign \new_[5886]_  = ~A268 & ~A267;
  assign \new_[5890]_  = A300 & A299;
  assign \new_[5891]_  = ~A269 & \new_[5890]_ ;
  assign \new_[5892]_  = \new_[5891]_  & \new_[5886]_ ;
  assign \new_[5895]_  = ~A167 & ~A169;
  assign \new_[5898]_  = A202 & ~A166;
  assign \new_[5899]_  = \new_[5898]_  & \new_[5895]_ ;
  assign \new_[5902]_  = ~A268 & ~A267;
  assign \new_[5906]_  = A300 & A298;
  assign \new_[5907]_  = ~A269 & \new_[5906]_ ;
  assign \new_[5908]_  = \new_[5907]_  & \new_[5902]_ ;
  assign \new_[5911]_  = ~A167 & ~A169;
  assign \new_[5914]_  = A202 & ~A166;
  assign \new_[5915]_  = \new_[5914]_  & \new_[5911]_ ;
  assign \new_[5918]_  = A266 & A265;
  assign \new_[5922]_  = A301 & ~A268;
  assign \new_[5923]_  = ~A267 & \new_[5922]_ ;
  assign \new_[5924]_  = \new_[5923]_  & \new_[5918]_ ;
  assign \new_[5927]_  = ~A167 & ~A169;
  assign \new_[5930]_  = A202 & ~A166;
  assign \new_[5931]_  = \new_[5930]_  & \new_[5927]_ ;
  assign \new_[5934]_  = ~A266 & ~A265;
  assign \new_[5938]_  = A300 & A299;
  assign \new_[5939]_  = ~A268 & \new_[5938]_ ;
  assign \new_[5940]_  = \new_[5939]_  & \new_[5934]_ ;
  assign \new_[5943]_  = ~A167 & ~A169;
  assign \new_[5946]_  = A202 & ~A166;
  assign \new_[5947]_  = \new_[5946]_  & \new_[5943]_ ;
  assign \new_[5950]_  = ~A266 & ~A265;
  assign \new_[5954]_  = A300 & A298;
  assign \new_[5955]_  = ~A268 & \new_[5954]_ ;
  assign \new_[5956]_  = \new_[5955]_  & \new_[5950]_ ;
  assign \new_[5959]_  = ~A167 & ~A169;
  assign \new_[5962]_  = A199 & ~A166;
  assign \new_[5963]_  = \new_[5962]_  & \new_[5959]_ ;
  assign \new_[5966]_  = ~A267 & A201;
  assign \new_[5970]_  = A301 & ~A269;
  assign \new_[5971]_  = ~A268 & \new_[5970]_ ;
  assign \new_[5972]_  = \new_[5971]_  & \new_[5966]_ ;
  assign \new_[5975]_  = ~A167 & ~A169;
  assign \new_[5978]_  = A199 & ~A166;
  assign \new_[5979]_  = \new_[5978]_  & \new_[5975]_ ;
  assign \new_[5982]_  = ~A265 & A201;
  assign \new_[5986]_  = A301 & ~A268;
  assign \new_[5987]_  = ~A266 & \new_[5986]_ ;
  assign \new_[5988]_  = \new_[5987]_  & \new_[5982]_ ;
  assign \new_[5991]_  = ~A167 & ~A169;
  assign \new_[5994]_  = A200 & ~A166;
  assign \new_[5995]_  = \new_[5994]_  & \new_[5991]_ ;
  assign \new_[5998]_  = ~A267 & A201;
  assign \new_[6002]_  = A301 & ~A269;
  assign \new_[6003]_  = ~A268 & \new_[6002]_ ;
  assign \new_[6004]_  = \new_[6003]_  & \new_[5998]_ ;
  assign \new_[6007]_  = ~A167 & ~A169;
  assign \new_[6010]_  = A200 & ~A166;
  assign \new_[6011]_  = \new_[6010]_  & \new_[6007]_ ;
  assign \new_[6014]_  = ~A265 & A201;
  assign \new_[6018]_  = A301 & ~A268;
  assign \new_[6019]_  = ~A266 & \new_[6018]_ ;
  assign \new_[6020]_  = \new_[6019]_  & \new_[6014]_ ;
  assign \new_[6023]_  = ~A168 & ~A169;
  assign \new_[6026]_  = A166 & A167;
  assign \new_[6027]_  = \new_[6026]_  & \new_[6023]_ ;
  assign \new_[6030]_  = ~A267 & A202;
  assign \new_[6034]_  = A301 & ~A269;
  assign \new_[6035]_  = ~A268 & \new_[6034]_ ;
  assign \new_[6036]_  = \new_[6035]_  & \new_[6030]_ ;
  assign \new_[6039]_  = ~A168 & ~A169;
  assign \new_[6042]_  = A166 & A167;
  assign \new_[6043]_  = \new_[6042]_  & \new_[6039]_ ;
  assign \new_[6046]_  = ~A265 & A202;
  assign \new_[6050]_  = A301 & ~A268;
  assign \new_[6051]_  = ~A266 & \new_[6050]_ ;
  assign \new_[6052]_  = \new_[6051]_  & \new_[6046]_ ;
  assign \new_[6055]_  = ~A169 & ~A170;
  assign \new_[6058]_  = A202 & ~A168;
  assign \new_[6059]_  = \new_[6058]_  & \new_[6055]_ ;
  assign \new_[6062]_  = ~A268 & ~A267;
  assign \new_[6066]_  = A300 & A299;
  assign \new_[6067]_  = ~A269 & \new_[6066]_ ;
  assign \new_[6068]_  = \new_[6067]_  & \new_[6062]_ ;
  assign \new_[6071]_  = ~A169 & ~A170;
  assign \new_[6074]_  = A202 & ~A168;
  assign \new_[6075]_  = \new_[6074]_  & \new_[6071]_ ;
  assign \new_[6078]_  = ~A268 & ~A267;
  assign \new_[6082]_  = A300 & A298;
  assign \new_[6083]_  = ~A269 & \new_[6082]_ ;
  assign \new_[6084]_  = \new_[6083]_  & \new_[6078]_ ;
  assign \new_[6087]_  = ~A169 & ~A170;
  assign \new_[6090]_  = A202 & ~A168;
  assign \new_[6091]_  = \new_[6090]_  & \new_[6087]_ ;
  assign \new_[6094]_  = A266 & A265;
  assign \new_[6098]_  = A301 & ~A268;
  assign \new_[6099]_  = ~A267 & \new_[6098]_ ;
  assign \new_[6100]_  = \new_[6099]_  & \new_[6094]_ ;
  assign \new_[6103]_  = ~A169 & ~A170;
  assign \new_[6106]_  = A202 & ~A168;
  assign \new_[6107]_  = \new_[6106]_  & \new_[6103]_ ;
  assign \new_[6110]_  = ~A266 & ~A265;
  assign \new_[6114]_  = A300 & A299;
  assign \new_[6115]_  = ~A268 & \new_[6114]_ ;
  assign \new_[6116]_  = \new_[6115]_  & \new_[6110]_ ;
  assign \new_[6119]_  = ~A169 & ~A170;
  assign \new_[6122]_  = A202 & ~A168;
  assign \new_[6123]_  = \new_[6122]_  & \new_[6119]_ ;
  assign \new_[6126]_  = ~A266 & ~A265;
  assign \new_[6130]_  = A300 & A298;
  assign \new_[6131]_  = ~A268 & \new_[6130]_ ;
  assign \new_[6132]_  = \new_[6131]_  & \new_[6126]_ ;
  assign \new_[6135]_  = ~A169 & ~A170;
  assign \new_[6138]_  = A199 & ~A168;
  assign \new_[6139]_  = \new_[6138]_  & \new_[6135]_ ;
  assign \new_[6142]_  = ~A267 & A201;
  assign \new_[6146]_  = A301 & ~A269;
  assign \new_[6147]_  = ~A268 & \new_[6146]_ ;
  assign \new_[6148]_  = \new_[6147]_  & \new_[6142]_ ;
  assign \new_[6151]_  = ~A169 & ~A170;
  assign \new_[6154]_  = A199 & ~A168;
  assign \new_[6155]_  = \new_[6154]_  & \new_[6151]_ ;
  assign \new_[6158]_  = ~A265 & A201;
  assign \new_[6162]_  = A301 & ~A268;
  assign \new_[6163]_  = ~A266 & \new_[6162]_ ;
  assign \new_[6164]_  = \new_[6163]_  & \new_[6158]_ ;
  assign \new_[6167]_  = ~A169 & ~A170;
  assign \new_[6170]_  = A200 & ~A168;
  assign \new_[6171]_  = \new_[6170]_  & \new_[6167]_ ;
  assign \new_[6174]_  = ~A267 & A201;
  assign \new_[6178]_  = A301 & ~A269;
  assign \new_[6179]_  = ~A268 & \new_[6178]_ ;
  assign \new_[6180]_  = \new_[6179]_  & \new_[6174]_ ;
  assign \new_[6183]_  = ~A169 & ~A170;
  assign \new_[6186]_  = A200 & ~A168;
  assign \new_[6187]_  = \new_[6186]_  & \new_[6183]_ ;
  assign \new_[6190]_  = ~A265 & A201;
  assign \new_[6194]_  = A301 & ~A268;
  assign \new_[6195]_  = ~A266 & \new_[6194]_ ;
  assign \new_[6196]_  = \new_[6195]_  & \new_[6190]_ ;
  assign \new_[6199]_  = A166 & A168;
  assign \new_[6203]_  = A266 & ~A265;
  assign \new_[6204]_  = A202 & \new_[6203]_ ;
  assign \new_[6205]_  = \new_[6204]_  & \new_[6199]_ ;
  assign \new_[6208]_  = A298 & A269;
  assign \new_[6212]_  = ~A301 & ~A300;
  assign \new_[6213]_  = A299 & \new_[6212]_ ;
  assign \new_[6214]_  = \new_[6213]_  & \new_[6208]_ ;
  assign \new_[6217]_  = A166 & A168;
  assign \new_[6221]_  = ~A266 & A265;
  assign \new_[6222]_  = A202 & \new_[6221]_ ;
  assign \new_[6223]_  = \new_[6222]_  & \new_[6217]_ ;
  assign \new_[6226]_  = A298 & A269;
  assign \new_[6230]_  = ~A301 & ~A300;
  assign \new_[6231]_  = A299 & \new_[6230]_ ;
  assign \new_[6232]_  = \new_[6231]_  & \new_[6226]_ ;
  assign \new_[6235]_  = A166 & A168;
  assign \new_[6239]_  = ~A203 & ~A202;
  assign \new_[6240]_  = ~A201 & \new_[6239]_ ;
  assign \new_[6241]_  = \new_[6240]_  & \new_[6235]_ ;
  assign \new_[6244]_  = ~A268 & ~A267;
  assign \new_[6248]_  = A300 & A299;
  assign \new_[6249]_  = ~A269 & \new_[6248]_ ;
  assign \new_[6250]_  = \new_[6249]_  & \new_[6244]_ ;
  assign \new_[6253]_  = A166 & A168;
  assign \new_[6257]_  = ~A203 & ~A202;
  assign \new_[6258]_  = ~A201 & \new_[6257]_ ;
  assign \new_[6259]_  = \new_[6258]_  & \new_[6253]_ ;
  assign \new_[6262]_  = ~A268 & ~A267;
  assign \new_[6266]_  = A300 & A298;
  assign \new_[6267]_  = ~A269 & \new_[6266]_ ;
  assign \new_[6268]_  = \new_[6267]_  & \new_[6262]_ ;
  assign \new_[6271]_  = A166 & A168;
  assign \new_[6275]_  = ~A203 & ~A202;
  assign \new_[6276]_  = ~A201 & \new_[6275]_ ;
  assign \new_[6277]_  = \new_[6276]_  & \new_[6271]_ ;
  assign \new_[6280]_  = A266 & A265;
  assign \new_[6284]_  = A301 & ~A268;
  assign \new_[6285]_  = ~A267 & \new_[6284]_ ;
  assign \new_[6286]_  = \new_[6285]_  & \new_[6280]_ ;
  assign \new_[6289]_  = A166 & A168;
  assign \new_[6293]_  = ~A203 & ~A202;
  assign \new_[6294]_  = ~A201 & \new_[6293]_ ;
  assign \new_[6295]_  = \new_[6294]_  & \new_[6289]_ ;
  assign \new_[6298]_  = ~A266 & ~A265;
  assign \new_[6302]_  = A300 & A299;
  assign \new_[6303]_  = ~A268 & \new_[6302]_ ;
  assign \new_[6304]_  = \new_[6303]_  & \new_[6298]_ ;
  assign \new_[6307]_  = A166 & A168;
  assign \new_[6311]_  = ~A203 & ~A202;
  assign \new_[6312]_  = ~A201 & \new_[6311]_ ;
  assign \new_[6313]_  = \new_[6312]_  & \new_[6307]_ ;
  assign \new_[6316]_  = ~A266 & ~A265;
  assign \new_[6320]_  = A300 & A298;
  assign \new_[6321]_  = ~A268 & \new_[6320]_ ;
  assign \new_[6322]_  = \new_[6321]_  & \new_[6316]_ ;
  assign \new_[6325]_  = A166 & A168;
  assign \new_[6329]_  = A265 & A201;
  assign \new_[6330]_  = A199 & \new_[6329]_ ;
  assign \new_[6331]_  = \new_[6330]_  & \new_[6325]_ ;
  assign \new_[6334]_  = A298 & A267;
  assign \new_[6338]_  = ~A301 & ~A300;
  assign \new_[6339]_  = A299 & \new_[6338]_ ;
  assign \new_[6340]_  = \new_[6339]_  & \new_[6334]_ ;
  assign \new_[6343]_  = A166 & A168;
  assign \new_[6347]_  = A266 & A201;
  assign \new_[6348]_  = A199 & \new_[6347]_ ;
  assign \new_[6349]_  = \new_[6348]_  & \new_[6343]_ ;
  assign \new_[6352]_  = A298 & A267;
  assign \new_[6356]_  = ~A301 & ~A300;
  assign \new_[6357]_  = A299 & \new_[6356]_ ;
  assign \new_[6358]_  = \new_[6357]_  & \new_[6352]_ ;
  assign \new_[6361]_  = A166 & A168;
  assign \new_[6365]_  = ~A265 & A201;
  assign \new_[6366]_  = A199 & \new_[6365]_ ;
  assign \new_[6367]_  = \new_[6366]_  & \new_[6361]_ ;
  assign \new_[6370]_  = A269 & A266;
  assign \new_[6374]_  = ~A302 & ~A301;
  assign \new_[6375]_  = ~A300 & \new_[6374]_ ;
  assign \new_[6376]_  = \new_[6375]_  & \new_[6370]_ ;
  assign \new_[6379]_  = A166 & A168;
  assign \new_[6383]_  = ~A265 & A201;
  assign \new_[6384]_  = A199 & \new_[6383]_ ;
  assign \new_[6385]_  = \new_[6384]_  & \new_[6379]_ ;
  assign \new_[6388]_  = A269 & A266;
  assign \new_[6392]_  = ~A301 & ~A299;
  assign \new_[6393]_  = ~A298 & \new_[6392]_ ;
  assign \new_[6394]_  = \new_[6393]_  & \new_[6388]_ ;
  assign \new_[6397]_  = A166 & A168;
  assign \new_[6401]_  = A265 & A201;
  assign \new_[6402]_  = A199 & \new_[6401]_ ;
  assign \new_[6403]_  = \new_[6402]_  & \new_[6397]_ ;
  assign \new_[6406]_  = A269 & ~A266;
  assign \new_[6410]_  = ~A302 & ~A301;
  assign \new_[6411]_  = ~A300 & \new_[6410]_ ;
  assign \new_[6412]_  = \new_[6411]_  & \new_[6406]_ ;
  assign \new_[6415]_  = A166 & A168;
  assign \new_[6419]_  = A265 & A201;
  assign \new_[6420]_  = A199 & \new_[6419]_ ;
  assign \new_[6421]_  = \new_[6420]_  & \new_[6415]_ ;
  assign \new_[6424]_  = A269 & ~A266;
  assign \new_[6428]_  = ~A301 & ~A299;
  assign \new_[6429]_  = ~A298 & \new_[6428]_ ;
  assign \new_[6430]_  = \new_[6429]_  & \new_[6424]_ ;
  assign \new_[6433]_  = A166 & A168;
  assign \new_[6437]_  = A265 & A201;
  assign \new_[6438]_  = A200 & \new_[6437]_ ;
  assign \new_[6439]_  = \new_[6438]_  & \new_[6433]_ ;
  assign \new_[6442]_  = A298 & A267;
  assign \new_[6446]_  = ~A301 & ~A300;
  assign \new_[6447]_  = A299 & \new_[6446]_ ;
  assign \new_[6448]_  = \new_[6447]_  & \new_[6442]_ ;
  assign \new_[6451]_  = A166 & A168;
  assign \new_[6455]_  = A266 & A201;
  assign \new_[6456]_  = A200 & \new_[6455]_ ;
  assign \new_[6457]_  = \new_[6456]_  & \new_[6451]_ ;
  assign \new_[6460]_  = A298 & A267;
  assign \new_[6464]_  = ~A301 & ~A300;
  assign \new_[6465]_  = A299 & \new_[6464]_ ;
  assign \new_[6466]_  = \new_[6465]_  & \new_[6460]_ ;
  assign \new_[6469]_  = A166 & A168;
  assign \new_[6473]_  = ~A265 & A201;
  assign \new_[6474]_  = A200 & \new_[6473]_ ;
  assign \new_[6475]_  = \new_[6474]_  & \new_[6469]_ ;
  assign \new_[6478]_  = A269 & A266;
  assign \new_[6482]_  = ~A302 & ~A301;
  assign \new_[6483]_  = ~A300 & \new_[6482]_ ;
  assign \new_[6484]_  = \new_[6483]_  & \new_[6478]_ ;
  assign \new_[6487]_  = A166 & A168;
  assign \new_[6491]_  = ~A265 & A201;
  assign \new_[6492]_  = A200 & \new_[6491]_ ;
  assign \new_[6493]_  = \new_[6492]_  & \new_[6487]_ ;
  assign \new_[6496]_  = A269 & A266;
  assign \new_[6500]_  = ~A301 & ~A299;
  assign \new_[6501]_  = ~A298 & \new_[6500]_ ;
  assign \new_[6502]_  = \new_[6501]_  & \new_[6496]_ ;
  assign \new_[6505]_  = A166 & A168;
  assign \new_[6509]_  = A265 & A201;
  assign \new_[6510]_  = A200 & \new_[6509]_ ;
  assign \new_[6511]_  = \new_[6510]_  & \new_[6505]_ ;
  assign \new_[6514]_  = A269 & ~A266;
  assign \new_[6518]_  = ~A302 & ~A301;
  assign \new_[6519]_  = ~A300 & \new_[6518]_ ;
  assign \new_[6520]_  = \new_[6519]_  & \new_[6514]_ ;
  assign \new_[6523]_  = A166 & A168;
  assign \new_[6527]_  = A265 & A201;
  assign \new_[6528]_  = A200 & \new_[6527]_ ;
  assign \new_[6529]_  = \new_[6528]_  & \new_[6523]_ ;
  assign \new_[6532]_  = A269 & ~A266;
  assign \new_[6536]_  = ~A301 & ~A299;
  assign \new_[6537]_  = ~A298 & \new_[6536]_ ;
  assign \new_[6538]_  = \new_[6537]_  & \new_[6532]_ ;
  assign \new_[6541]_  = A166 & A168;
  assign \new_[6545]_  = ~A201 & A200;
  assign \new_[6546]_  = A199 & \new_[6545]_ ;
  assign \new_[6547]_  = \new_[6546]_  & \new_[6541]_ ;
  assign \new_[6550]_  = ~A267 & ~A202;
  assign \new_[6554]_  = A301 & ~A269;
  assign \new_[6555]_  = ~A268 & \new_[6554]_ ;
  assign \new_[6556]_  = \new_[6555]_  & \new_[6550]_ ;
  assign \new_[6559]_  = A166 & A168;
  assign \new_[6563]_  = ~A201 & A200;
  assign \new_[6564]_  = A199 & \new_[6563]_ ;
  assign \new_[6565]_  = \new_[6564]_  & \new_[6559]_ ;
  assign \new_[6568]_  = ~A265 & ~A202;
  assign \new_[6572]_  = A301 & ~A268;
  assign \new_[6573]_  = ~A266 & \new_[6572]_ ;
  assign \new_[6574]_  = \new_[6573]_  & \new_[6568]_ ;
  assign \new_[6577]_  = A166 & A168;
  assign \new_[6581]_  = A203 & A200;
  assign \new_[6582]_  = ~A199 & \new_[6581]_ ;
  assign \new_[6583]_  = \new_[6582]_  & \new_[6577]_ ;
  assign \new_[6586]_  = A298 & A268;
  assign \new_[6590]_  = ~A301 & ~A300;
  assign \new_[6591]_  = A299 & \new_[6590]_ ;
  assign \new_[6592]_  = \new_[6591]_  & \new_[6586]_ ;
  assign \new_[6595]_  = A166 & A168;
  assign \new_[6599]_  = A203 & A200;
  assign \new_[6600]_  = ~A199 & \new_[6599]_ ;
  assign \new_[6601]_  = \new_[6600]_  & \new_[6595]_ ;
  assign \new_[6604]_  = A267 & A265;
  assign \new_[6608]_  = ~A302 & ~A301;
  assign \new_[6609]_  = ~A300 & \new_[6608]_ ;
  assign \new_[6610]_  = \new_[6609]_  & \new_[6604]_ ;
  assign \new_[6613]_  = A166 & A168;
  assign \new_[6617]_  = A203 & A200;
  assign \new_[6618]_  = ~A199 & \new_[6617]_ ;
  assign \new_[6619]_  = \new_[6618]_  & \new_[6613]_ ;
  assign \new_[6622]_  = A267 & A265;
  assign \new_[6626]_  = ~A301 & ~A299;
  assign \new_[6627]_  = ~A298 & \new_[6626]_ ;
  assign \new_[6628]_  = \new_[6627]_  & \new_[6622]_ ;
  assign \new_[6631]_  = A166 & A168;
  assign \new_[6635]_  = A203 & A200;
  assign \new_[6636]_  = ~A199 & \new_[6635]_ ;
  assign \new_[6637]_  = \new_[6636]_  & \new_[6631]_ ;
  assign \new_[6640]_  = A267 & A266;
  assign \new_[6644]_  = ~A302 & ~A301;
  assign \new_[6645]_  = ~A300 & \new_[6644]_ ;
  assign \new_[6646]_  = \new_[6645]_  & \new_[6640]_ ;
  assign \new_[6649]_  = A166 & A168;
  assign \new_[6653]_  = A203 & A200;
  assign \new_[6654]_  = ~A199 & \new_[6653]_ ;
  assign \new_[6655]_  = \new_[6654]_  & \new_[6649]_ ;
  assign \new_[6658]_  = A267 & A266;
  assign \new_[6662]_  = ~A301 & ~A299;
  assign \new_[6663]_  = ~A298 & \new_[6662]_ ;
  assign \new_[6664]_  = \new_[6663]_  & \new_[6658]_ ;
  assign \new_[6667]_  = A166 & A168;
  assign \new_[6671]_  = A203 & ~A200;
  assign \new_[6672]_  = A199 & \new_[6671]_ ;
  assign \new_[6673]_  = \new_[6672]_  & \new_[6667]_ ;
  assign \new_[6676]_  = A298 & A268;
  assign \new_[6680]_  = ~A301 & ~A300;
  assign \new_[6681]_  = A299 & \new_[6680]_ ;
  assign \new_[6682]_  = \new_[6681]_  & \new_[6676]_ ;
  assign \new_[6685]_  = A166 & A168;
  assign \new_[6689]_  = A203 & ~A200;
  assign \new_[6690]_  = A199 & \new_[6689]_ ;
  assign \new_[6691]_  = \new_[6690]_  & \new_[6685]_ ;
  assign \new_[6694]_  = A267 & A265;
  assign \new_[6698]_  = ~A302 & ~A301;
  assign \new_[6699]_  = ~A300 & \new_[6698]_ ;
  assign \new_[6700]_  = \new_[6699]_  & \new_[6694]_ ;
  assign \new_[6703]_  = A166 & A168;
  assign \new_[6707]_  = A203 & ~A200;
  assign \new_[6708]_  = A199 & \new_[6707]_ ;
  assign \new_[6709]_  = \new_[6708]_  & \new_[6703]_ ;
  assign \new_[6712]_  = A267 & A265;
  assign \new_[6716]_  = ~A301 & ~A299;
  assign \new_[6717]_  = ~A298 & \new_[6716]_ ;
  assign \new_[6718]_  = \new_[6717]_  & \new_[6712]_ ;
  assign \new_[6721]_  = A166 & A168;
  assign \new_[6725]_  = A203 & ~A200;
  assign \new_[6726]_  = A199 & \new_[6725]_ ;
  assign \new_[6727]_  = \new_[6726]_  & \new_[6721]_ ;
  assign \new_[6730]_  = A267 & A266;
  assign \new_[6734]_  = ~A302 & ~A301;
  assign \new_[6735]_  = ~A300 & \new_[6734]_ ;
  assign \new_[6736]_  = \new_[6735]_  & \new_[6730]_ ;
  assign \new_[6739]_  = A166 & A168;
  assign \new_[6743]_  = A203 & ~A200;
  assign \new_[6744]_  = A199 & \new_[6743]_ ;
  assign \new_[6745]_  = \new_[6744]_  & \new_[6739]_ ;
  assign \new_[6748]_  = A267 & A266;
  assign \new_[6752]_  = ~A301 & ~A299;
  assign \new_[6753]_  = ~A298 & \new_[6752]_ ;
  assign \new_[6754]_  = \new_[6753]_  & \new_[6748]_ ;
  assign \new_[6757]_  = A166 & A168;
  assign \new_[6761]_  = ~A202 & ~A200;
  assign \new_[6762]_  = ~A199 & \new_[6761]_ ;
  assign \new_[6763]_  = \new_[6762]_  & \new_[6757]_ ;
  assign \new_[6766]_  = ~A268 & ~A267;
  assign \new_[6770]_  = A300 & A299;
  assign \new_[6771]_  = ~A269 & \new_[6770]_ ;
  assign \new_[6772]_  = \new_[6771]_  & \new_[6766]_ ;
  assign \new_[6775]_  = A166 & A168;
  assign \new_[6779]_  = ~A202 & ~A200;
  assign \new_[6780]_  = ~A199 & \new_[6779]_ ;
  assign \new_[6781]_  = \new_[6780]_  & \new_[6775]_ ;
  assign \new_[6784]_  = ~A268 & ~A267;
  assign \new_[6788]_  = A300 & A298;
  assign \new_[6789]_  = ~A269 & \new_[6788]_ ;
  assign \new_[6790]_  = \new_[6789]_  & \new_[6784]_ ;
  assign \new_[6793]_  = A166 & A168;
  assign \new_[6797]_  = ~A202 & ~A200;
  assign \new_[6798]_  = ~A199 & \new_[6797]_ ;
  assign \new_[6799]_  = \new_[6798]_  & \new_[6793]_ ;
  assign \new_[6802]_  = A266 & A265;
  assign \new_[6806]_  = A301 & ~A268;
  assign \new_[6807]_  = ~A267 & \new_[6806]_ ;
  assign \new_[6808]_  = \new_[6807]_  & \new_[6802]_ ;
  assign \new_[6811]_  = A166 & A168;
  assign \new_[6815]_  = ~A202 & ~A200;
  assign \new_[6816]_  = ~A199 & \new_[6815]_ ;
  assign \new_[6817]_  = \new_[6816]_  & \new_[6811]_ ;
  assign \new_[6820]_  = ~A266 & ~A265;
  assign \new_[6824]_  = A300 & A299;
  assign \new_[6825]_  = ~A268 & \new_[6824]_ ;
  assign \new_[6826]_  = \new_[6825]_  & \new_[6820]_ ;
  assign \new_[6829]_  = A166 & A168;
  assign \new_[6833]_  = ~A202 & ~A200;
  assign \new_[6834]_  = ~A199 & \new_[6833]_ ;
  assign \new_[6835]_  = \new_[6834]_  & \new_[6829]_ ;
  assign \new_[6838]_  = ~A266 & ~A265;
  assign \new_[6842]_  = A300 & A298;
  assign \new_[6843]_  = ~A268 & \new_[6842]_ ;
  assign \new_[6844]_  = \new_[6843]_  & \new_[6838]_ ;
  assign \new_[6847]_  = A167 & A168;
  assign \new_[6851]_  = A266 & ~A265;
  assign \new_[6852]_  = A202 & \new_[6851]_ ;
  assign \new_[6853]_  = \new_[6852]_  & \new_[6847]_ ;
  assign \new_[6856]_  = A298 & A269;
  assign \new_[6860]_  = ~A301 & ~A300;
  assign \new_[6861]_  = A299 & \new_[6860]_ ;
  assign \new_[6862]_  = \new_[6861]_  & \new_[6856]_ ;
  assign \new_[6865]_  = A167 & A168;
  assign \new_[6869]_  = ~A266 & A265;
  assign \new_[6870]_  = A202 & \new_[6869]_ ;
  assign \new_[6871]_  = \new_[6870]_  & \new_[6865]_ ;
  assign \new_[6874]_  = A298 & A269;
  assign \new_[6878]_  = ~A301 & ~A300;
  assign \new_[6879]_  = A299 & \new_[6878]_ ;
  assign \new_[6880]_  = \new_[6879]_  & \new_[6874]_ ;
  assign \new_[6883]_  = A167 & A168;
  assign \new_[6887]_  = ~A203 & ~A202;
  assign \new_[6888]_  = ~A201 & \new_[6887]_ ;
  assign \new_[6889]_  = \new_[6888]_  & \new_[6883]_ ;
  assign \new_[6892]_  = ~A268 & ~A267;
  assign \new_[6896]_  = A300 & A299;
  assign \new_[6897]_  = ~A269 & \new_[6896]_ ;
  assign \new_[6898]_  = \new_[6897]_  & \new_[6892]_ ;
  assign \new_[6901]_  = A167 & A168;
  assign \new_[6905]_  = ~A203 & ~A202;
  assign \new_[6906]_  = ~A201 & \new_[6905]_ ;
  assign \new_[6907]_  = \new_[6906]_  & \new_[6901]_ ;
  assign \new_[6910]_  = ~A268 & ~A267;
  assign \new_[6914]_  = A300 & A298;
  assign \new_[6915]_  = ~A269 & \new_[6914]_ ;
  assign \new_[6916]_  = \new_[6915]_  & \new_[6910]_ ;
  assign \new_[6919]_  = A167 & A168;
  assign \new_[6923]_  = ~A203 & ~A202;
  assign \new_[6924]_  = ~A201 & \new_[6923]_ ;
  assign \new_[6925]_  = \new_[6924]_  & \new_[6919]_ ;
  assign \new_[6928]_  = A266 & A265;
  assign \new_[6932]_  = A301 & ~A268;
  assign \new_[6933]_  = ~A267 & \new_[6932]_ ;
  assign \new_[6934]_  = \new_[6933]_  & \new_[6928]_ ;
  assign \new_[6937]_  = A167 & A168;
  assign \new_[6941]_  = ~A203 & ~A202;
  assign \new_[6942]_  = ~A201 & \new_[6941]_ ;
  assign \new_[6943]_  = \new_[6942]_  & \new_[6937]_ ;
  assign \new_[6946]_  = ~A266 & ~A265;
  assign \new_[6950]_  = A300 & A299;
  assign \new_[6951]_  = ~A268 & \new_[6950]_ ;
  assign \new_[6952]_  = \new_[6951]_  & \new_[6946]_ ;
  assign \new_[6955]_  = A167 & A168;
  assign \new_[6959]_  = ~A203 & ~A202;
  assign \new_[6960]_  = ~A201 & \new_[6959]_ ;
  assign \new_[6961]_  = \new_[6960]_  & \new_[6955]_ ;
  assign \new_[6964]_  = ~A266 & ~A265;
  assign \new_[6968]_  = A300 & A298;
  assign \new_[6969]_  = ~A268 & \new_[6968]_ ;
  assign \new_[6970]_  = \new_[6969]_  & \new_[6964]_ ;
  assign \new_[6973]_  = A167 & A168;
  assign \new_[6977]_  = A265 & A201;
  assign \new_[6978]_  = A199 & \new_[6977]_ ;
  assign \new_[6979]_  = \new_[6978]_  & \new_[6973]_ ;
  assign \new_[6982]_  = A298 & A267;
  assign \new_[6986]_  = ~A301 & ~A300;
  assign \new_[6987]_  = A299 & \new_[6986]_ ;
  assign \new_[6988]_  = \new_[6987]_  & \new_[6982]_ ;
  assign \new_[6991]_  = A167 & A168;
  assign \new_[6995]_  = A266 & A201;
  assign \new_[6996]_  = A199 & \new_[6995]_ ;
  assign \new_[6997]_  = \new_[6996]_  & \new_[6991]_ ;
  assign \new_[7000]_  = A298 & A267;
  assign \new_[7004]_  = ~A301 & ~A300;
  assign \new_[7005]_  = A299 & \new_[7004]_ ;
  assign \new_[7006]_  = \new_[7005]_  & \new_[7000]_ ;
  assign \new_[7009]_  = A167 & A168;
  assign \new_[7013]_  = ~A265 & A201;
  assign \new_[7014]_  = A199 & \new_[7013]_ ;
  assign \new_[7015]_  = \new_[7014]_  & \new_[7009]_ ;
  assign \new_[7018]_  = A269 & A266;
  assign \new_[7022]_  = ~A302 & ~A301;
  assign \new_[7023]_  = ~A300 & \new_[7022]_ ;
  assign \new_[7024]_  = \new_[7023]_  & \new_[7018]_ ;
  assign \new_[7027]_  = A167 & A168;
  assign \new_[7031]_  = ~A265 & A201;
  assign \new_[7032]_  = A199 & \new_[7031]_ ;
  assign \new_[7033]_  = \new_[7032]_  & \new_[7027]_ ;
  assign \new_[7036]_  = A269 & A266;
  assign \new_[7040]_  = ~A301 & ~A299;
  assign \new_[7041]_  = ~A298 & \new_[7040]_ ;
  assign \new_[7042]_  = \new_[7041]_  & \new_[7036]_ ;
  assign \new_[7045]_  = A167 & A168;
  assign \new_[7049]_  = A265 & A201;
  assign \new_[7050]_  = A199 & \new_[7049]_ ;
  assign \new_[7051]_  = \new_[7050]_  & \new_[7045]_ ;
  assign \new_[7054]_  = A269 & ~A266;
  assign \new_[7058]_  = ~A302 & ~A301;
  assign \new_[7059]_  = ~A300 & \new_[7058]_ ;
  assign \new_[7060]_  = \new_[7059]_  & \new_[7054]_ ;
  assign \new_[7063]_  = A167 & A168;
  assign \new_[7067]_  = A265 & A201;
  assign \new_[7068]_  = A199 & \new_[7067]_ ;
  assign \new_[7069]_  = \new_[7068]_  & \new_[7063]_ ;
  assign \new_[7072]_  = A269 & ~A266;
  assign \new_[7076]_  = ~A301 & ~A299;
  assign \new_[7077]_  = ~A298 & \new_[7076]_ ;
  assign \new_[7078]_  = \new_[7077]_  & \new_[7072]_ ;
  assign \new_[7081]_  = A167 & A168;
  assign \new_[7085]_  = A265 & A201;
  assign \new_[7086]_  = A200 & \new_[7085]_ ;
  assign \new_[7087]_  = \new_[7086]_  & \new_[7081]_ ;
  assign \new_[7090]_  = A298 & A267;
  assign \new_[7094]_  = ~A301 & ~A300;
  assign \new_[7095]_  = A299 & \new_[7094]_ ;
  assign \new_[7096]_  = \new_[7095]_  & \new_[7090]_ ;
  assign \new_[7099]_  = A167 & A168;
  assign \new_[7103]_  = A266 & A201;
  assign \new_[7104]_  = A200 & \new_[7103]_ ;
  assign \new_[7105]_  = \new_[7104]_  & \new_[7099]_ ;
  assign \new_[7108]_  = A298 & A267;
  assign \new_[7112]_  = ~A301 & ~A300;
  assign \new_[7113]_  = A299 & \new_[7112]_ ;
  assign \new_[7114]_  = \new_[7113]_  & \new_[7108]_ ;
  assign \new_[7117]_  = A167 & A168;
  assign \new_[7121]_  = ~A265 & A201;
  assign \new_[7122]_  = A200 & \new_[7121]_ ;
  assign \new_[7123]_  = \new_[7122]_  & \new_[7117]_ ;
  assign \new_[7126]_  = A269 & A266;
  assign \new_[7130]_  = ~A302 & ~A301;
  assign \new_[7131]_  = ~A300 & \new_[7130]_ ;
  assign \new_[7132]_  = \new_[7131]_  & \new_[7126]_ ;
  assign \new_[7135]_  = A167 & A168;
  assign \new_[7139]_  = ~A265 & A201;
  assign \new_[7140]_  = A200 & \new_[7139]_ ;
  assign \new_[7141]_  = \new_[7140]_  & \new_[7135]_ ;
  assign \new_[7144]_  = A269 & A266;
  assign \new_[7148]_  = ~A301 & ~A299;
  assign \new_[7149]_  = ~A298 & \new_[7148]_ ;
  assign \new_[7150]_  = \new_[7149]_  & \new_[7144]_ ;
  assign \new_[7153]_  = A167 & A168;
  assign \new_[7157]_  = A265 & A201;
  assign \new_[7158]_  = A200 & \new_[7157]_ ;
  assign \new_[7159]_  = \new_[7158]_  & \new_[7153]_ ;
  assign \new_[7162]_  = A269 & ~A266;
  assign \new_[7166]_  = ~A302 & ~A301;
  assign \new_[7167]_  = ~A300 & \new_[7166]_ ;
  assign \new_[7168]_  = \new_[7167]_  & \new_[7162]_ ;
  assign \new_[7171]_  = A167 & A168;
  assign \new_[7175]_  = A265 & A201;
  assign \new_[7176]_  = A200 & \new_[7175]_ ;
  assign \new_[7177]_  = \new_[7176]_  & \new_[7171]_ ;
  assign \new_[7180]_  = A269 & ~A266;
  assign \new_[7184]_  = ~A301 & ~A299;
  assign \new_[7185]_  = ~A298 & \new_[7184]_ ;
  assign \new_[7186]_  = \new_[7185]_  & \new_[7180]_ ;
  assign \new_[7189]_  = A167 & A168;
  assign \new_[7193]_  = ~A201 & A200;
  assign \new_[7194]_  = A199 & \new_[7193]_ ;
  assign \new_[7195]_  = \new_[7194]_  & \new_[7189]_ ;
  assign \new_[7198]_  = ~A267 & ~A202;
  assign \new_[7202]_  = A301 & ~A269;
  assign \new_[7203]_  = ~A268 & \new_[7202]_ ;
  assign \new_[7204]_  = \new_[7203]_  & \new_[7198]_ ;
  assign \new_[7207]_  = A167 & A168;
  assign \new_[7211]_  = ~A201 & A200;
  assign \new_[7212]_  = A199 & \new_[7211]_ ;
  assign \new_[7213]_  = \new_[7212]_  & \new_[7207]_ ;
  assign \new_[7216]_  = ~A265 & ~A202;
  assign \new_[7220]_  = A301 & ~A268;
  assign \new_[7221]_  = ~A266 & \new_[7220]_ ;
  assign \new_[7222]_  = \new_[7221]_  & \new_[7216]_ ;
  assign \new_[7225]_  = A167 & A168;
  assign \new_[7229]_  = A203 & A200;
  assign \new_[7230]_  = ~A199 & \new_[7229]_ ;
  assign \new_[7231]_  = \new_[7230]_  & \new_[7225]_ ;
  assign \new_[7234]_  = A298 & A268;
  assign \new_[7238]_  = ~A301 & ~A300;
  assign \new_[7239]_  = A299 & \new_[7238]_ ;
  assign \new_[7240]_  = \new_[7239]_  & \new_[7234]_ ;
  assign \new_[7243]_  = A167 & A168;
  assign \new_[7247]_  = A203 & A200;
  assign \new_[7248]_  = ~A199 & \new_[7247]_ ;
  assign \new_[7249]_  = \new_[7248]_  & \new_[7243]_ ;
  assign \new_[7252]_  = A267 & A265;
  assign \new_[7256]_  = ~A302 & ~A301;
  assign \new_[7257]_  = ~A300 & \new_[7256]_ ;
  assign \new_[7258]_  = \new_[7257]_  & \new_[7252]_ ;
  assign \new_[7261]_  = A167 & A168;
  assign \new_[7265]_  = A203 & A200;
  assign \new_[7266]_  = ~A199 & \new_[7265]_ ;
  assign \new_[7267]_  = \new_[7266]_  & \new_[7261]_ ;
  assign \new_[7270]_  = A267 & A265;
  assign \new_[7274]_  = ~A301 & ~A299;
  assign \new_[7275]_  = ~A298 & \new_[7274]_ ;
  assign \new_[7276]_  = \new_[7275]_  & \new_[7270]_ ;
  assign \new_[7279]_  = A167 & A168;
  assign \new_[7283]_  = A203 & A200;
  assign \new_[7284]_  = ~A199 & \new_[7283]_ ;
  assign \new_[7285]_  = \new_[7284]_  & \new_[7279]_ ;
  assign \new_[7288]_  = A267 & A266;
  assign \new_[7292]_  = ~A302 & ~A301;
  assign \new_[7293]_  = ~A300 & \new_[7292]_ ;
  assign \new_[7294]_  = \new_[7293]_  & \new_[7288]_ ;
  assign \new_[7297]_  = A167 & A168;
  assign \new_[7301]_  = A203 & A200;
  assign \new_[7302]_  = ~A199 & \new_[7301]_ ;
  assign \new_[7303]_  = \new_[7302]_  & \new_[7297]_ ;
  assign \new_[7306]_  = A267 & A266;
  assign \new_[7310]_  = ~A301 & ~A299;
  assign \new_[7311]_  = ~A298 & \new_[7310]_ ;
  assign \new_[7312]_  = \new_[7311]_  & \new_[7306]_ ;
  assign \new_[7315]_  = A167 & A168;
  assign \new_[7319]_  = A203 & ~A200;
  assign \new_[7320]_  = A199 & \new_[7319]_ ;
  assign \new_[7321]_  = \new_[7320]_  & \new_[7315]_ ;
  assign \new_[7324]_  = A298 & A268;
  assign \new_[7328]_  = ~A301 & ~A300;
  assign \new_[7329]_  = A299 & \new_[7328]_ ;
  assign \new_[7330]_  = \new_[7329]_  & \new_[7324]_ ;
  assign \new_[7333]_  = A167 & A168;
  assign \new_[7337]_  = A203 & ~A200;
  assign \new_[7338]_  = A199 & \new_[7337]_ ;
  assign \new_[7339]_  = \new_[7338]_  & \new_[7333]_ ;
  assign \new_[7342]_  = A267 & A265;
  assign \new_[7346]_  = ~A302 & ~A301;
  assign \new_[7347]_  = ~A300 & \new_[7346]_ ;
  assign \new_[7348]_  = \new_[7347]_  & \new_[7342]_ ;
  assign \new_[7351]_  = A167 & A168;
  assign \new_[7355]_  = A203 & ~A200;
  assign \new_[7356]_  = A199 & \new_[7355]_ ;
  assign \new_[7357]_  = \new_[7356]_  & \new_[7351]_ ;
  assign \new_[7360]_  = A267 & A265;
  assign \new_[7364]_  = ~A301 & ~A299;
  assign \new_[7365]_  = ~A298 & \new_[7364]_ ;
  assign \new_[7366]_  = \new_[7365]_  & \new_[7360]_ ;
  assign \new_[7369]_  = A167 & A168;
  assign \new_[7373]_  = A203 & ~A200;
  assign \new_[7374]_  = A199 & \new_[7373]_ ;
  assign \new_[7375]_  = \new_[7374]_  & \new_[7369]_ ;
  assign \new_[7378]_  = A267 & A266;
  assign \new_[7382]_  = ~A302 & ~A301;
  assign \new_[7383]_  = ~A300 & \new_[7382]_ ;
  assign \new_[7384]_  = \new_[7383]_  & \new_[7378]_ ;
  assign \new_[7387]_  = A167 & A168;
  assign \new_[7391]_  = A203 & ~A200;
  assign \new_[7392]_  = A199 & \new_[7391]_ ;
  assign \new_[7393]_  = \new_[7392]_  & \new_[7387]_ ;
  assign \new_[7396]_  = A267 & A266;
  assign \new_[7400]_  = ~A301 & ~A299;
  assign \new_[7401]_  = ~A298 & \new_[7400]_ ;
  assign \new_[7402]_  = \new_[7401]_  & \new_[7396]_ ;
  assign \new_[7405]_  = A167 & A168;
  assign \new_[7409]_  = ~A202 & ~A200;
  assign \new_[7410]_  = ~A199 & \new_[7409]_ ;
  assign \new_[7411]_  = \new_[7410]_  & \new_[7405]_ ;
  assign \new_[7414]_  = ~A268 & ~A267;
  assign \new_[7418]_  = A300 & A299;
  assign \new_[7419]_  = ~A269 & \new_[7418]_ ;
  assign \new_[7420]_  = \new_[7419]_  & \new_[7414]_ ;
  assign \new_[7423]_  = A167 & A168;
  assign \new_[7427]_  = ~A202 & ~A200;
  assign \new_[7428]_  = ~A199 & \new_[7427]_ ;
  assign \new_[7429]_  = \new_[7428]_  & \new_[7423]_ ;
  assign \new_[7432]_  = ~A268 & ~A267;
  assign \new_[7436]_  = A300 & A298;
  assign \new_[7437]_  = ~A269 & \new_[7436]_ ;
  assign \new_[7438]_  = \new_[7437]_  & \new_[7432]_ ;
  assign \new_[7441]_  = A167 & A168;
  assign \new_[7445]_  = ~A202 & ~A200;
  assign \new_[7446]_  = ~A199 & \new_[7445]_ ;
  assign \new_[7447]_  = \new_[7446]_  & \new_[7441]_ ;
  assign \new_[7450]_  = A266 & A265;
  assign \new_[7454]_  = A301 & ~A268;
  assign \new_[7455]_  = ~A267 & \new_[7454]_ ;
  assign \new_[7456]_  = \new_[7455]_  & \new_[7450]_ ;
  assign \new_[7459]_  = A167 & A168;
  assign \new_[7463]_  = ~A202 & ~A200;
  assign \new_[7464]_  = ~A199 & \new_[7463]_ ;
  assign \new_[7465]_  = \new_[7464]_  & \new_[7459]_ ;
  assign \new_[7468]_  = ~A266 & ~A265;
  assign \new_[7472]_  = A300 & A299;
  assign \new_[7473]_  = ~A268 & \new_[7472]_ ;
  assign \new_[7474]_  = \new_[7473]_  & \new_[7468]_ ;
  assign \new_[7477]_  = A167 & A168;
  assign \new_[7481]_  = ~A202 & ~A200;
  assign \new_[7482]_  = ~A199 & \new_[7481]_ ;
  assign \new_[7483]_  = \new_[7482]_  & \new_[7477]_ ;
  assign \new_[7486]_  = ~A266 & ~A265;
  assign \new_[7490]_  = A300 & A298;
  assign \new_[7491]_  = ~A268 & \new_[7490]_ ;
  assign \new_[7492]_  = \new_[7491]_  & \new_[7486]_ ;
  assign \new_[7495]_  = A167 & A170;
  assign \new_[7499]_  = A265 & A202;
  assign \new_[7500]_  = ~A166 & \new_[7499]_ ;
  assign \new_[7501]_  = \new_[7500]_  & \new_[7495]_ ;
  assign \new_[7504]_  = A298 & A267;
  assign \new_[7508]_  = ~A301 & ~A300;
  assign \new_[7509]_  = A299 & \new_[7508]_ ;
  assign \new_[7510]_  = \new_[7509]_  & \new_[7504]_ ;
  assign \new_[7513]_  = A167 & A170;
  assign \new_[7517]_  = A266 & A202;
  assign \new_[7518]_  = ~A166 & \new_[7517]_ ;
  assign \new_[7519]_  = \new_[7518]_  & \new_[7513]_ ;
  assign \new_[7522]_  = A298 & A267;
  assign \new_[7526]_  = ~A301 & ~A300;
  assign \new_[7527]_  = A299 & \new_[7526]_ ;
  assign \new_[7528]_  = \new_[7527]_  & \new_[7522]_ ;
  assign \new_[7531]_  = A167 & A170;
  assign \new_[7535]_  = ~A265 & A202;
  assign \new_[7536]_  = ~A166 & \new_[7535]_ ;
  assign \new_[7537]_  = \new_[7536]_  & \new_[7531]_ ;
  assign \new_[7540]_  = A269 & A266;
  assign \new_[7544]_  = ~A302 & ~A301;
  assign \new_[7545]_  = ~A300 & \new_[7544]_ ;
  assign \new_[7546]_  = \new_[7545]_  & \new_[7540]_ ;
  assign \new_[7549]_  = A167 & A170;
  assign \new_[7553]_  = ~A265 & A202;
  assign \new_[7554]_  = ~A166 & \new_[7553]_ ;
  assign \new_[7555]_  = \new_[7554]_  & \new_[7549]_ ;
  assign \new_[7558]_  = A269 & A266;
  assign \new_[7562]_  = ~A301 & ~A299;
  assign \new_[7563]_  = ~A298 & \new_[7562]_ ;
  assign \new_[7564]_  = \new_[7563]_  & \new_[7558]_ ;
  assign \new_[7567]_  = A167 & A170;
  assign \new_[7571]_  = A265 & A202;
  assign \new_[7572]_  = ~A166 & \new_[7571]_ ;
  assign \new_[7573]_  = \new_[7572]_  & \new_[7567]_ ;
  assign \new_[7576]_  = A269 & ~A266;
  assign \new_[7580]_  = ~A302 & ~A301;
  assign \new_[7581]_  = ~A300 & \new_[7580]_ ;
  assign \new_[7582]_  = \new_[7581]_  & \new_[7576]_ ;
  assign \new_[7585]_  = A167 & A170;
  assign \new_[7589]_  = A265 & A202;
  assign \new_[7590]_  = ~A166 & \new_[7589]_ ;
  assign \new_[7591]_  = \new_[7590]_  & \new_[7585]_ ;
  assign \new_[7594]_  = A269 & ~A266;
  assign \new_[7598]_  = ~A301 & ~A299;
  assign \new_[7599]_  = ~A298 & \new_[7598]_ ;
  assign \new_[7600]_  = \new_[7599]_  & \new_[7594]_ ;
  assign \new_[7603]_  = A167 & A170;
  assign \new_[7607]_  = ~A202 & ~A201;
  assign \new_[7608]_  = ~A166 & \new_[7607]_ ;
  assign \new_[7609]_  = \new_[7608]_  & \new_[7603]_ ;
  assign \new_[7612]_  = ~A267 & ~A203;
  assign \new_[7616]_  = A301 & ~A269;
  assign \new_[7617]_  = ~A268 & \new_[7616]_ ;
  assign \new_[7618]_  = \new_[7617]_  & \new_[7612]_ ;
  assign \new_[7621]_  = A167 & A170;
  assign \new_[7625]_  = ~A202 & ~A201;
  assign \new_[7626]_  = ~A166 & \new_[7625]_ ;
  assign \new_[7627]_  = \new_[7626]_  & \new_[7621]_ ;
  assign \new_[7630]_  = ~A265 & ~A203;
  assign \new_[7634]_  = A301 & ~A268;
  assign \new_[7635]_  = ~A266 & \new_[7634]_ ;
  assign \new_[7636]_  = \new_[7635]_  & \new_[7630]_ ;
  assign \new_[7639]_  = A167 & A170;
  assign \new_[7643]_  = A201 & A199;
  assign \new_[7644]_  = ~A166 & \new_[7643]_ ;
  assign \new_[7645]_  = \new_[7644]_  & \new_[7639]_ ;
  assign \new_[7648]_  = A298 & A268;
  assign \new_[7652]_  = ~A301 & ~A300;
  assign \new_[7653]_  = A299 & \new_[7652]_ ;
  assign \new_[7654]_  = \new_[7653]_  & \new_[7648]_ ;
  assign \new_[7657]_  = A167 & A170;
  assign \new_[7661]_  = A201 & A199;
  assign \new_[7662]_  = ~A166 & \new_[7661]_ ;
  assign \new_[7663]_  = \new_[7662]_  & \new_[7657]_ ;
  assign \new_[7666]_  = A267 & A265;
  assign \new_[7670]_  = ~A302 & ~A301;
  assign \new_[7671]_  = ~A300 & \new_[7670]_ ;
  assign \new_[7672]_  = \new_[7671]_  & \new_[7666]_ ;
  assign \new_[7675]_  = A167 & A170;
  assign \new_[7679]_  = A201 & A199;
  assign \new_[7680]_  = ~A166 & \new_[7679]_ ;
  assign \new_[7681]_  = \new_[7680]_  & \new_[7675]_ ;
  assign \new_[7684]_  = A267 & A265;
  assign \new_[7688]_  = ~A301 & ~A299;
  assign \new_[7689]_  = ~A298 & \new_[7688]_ ;
  assign \new_[7690]_  = \new_[7689]_  & \new_[7684]_ ;
  assign \new_[7693]_  = A167 & A170;
  assign \new_[7697]_  = A201 & A199;
  assign \new_[7698]_  = ~A166 & \new_[7697]_ ;
  assign \new_[7699]_  = \new_[7698]_  & \new_[7693]_ ;
  assign \new_[7702]_  = A267 & A266;
  assign \new_[7706]_  = ~A302 & ~A301;
  assign \new_[7707]_  = ~A300 & \new_[7706]_ ;
  assign \new_[7708]_  = \new_[7707]_  & \new_[7702]_ ;
  assign \new_[7711]_  = A167 & A170;
  assign \new_[7715]_  = A201 & A199;
  assign \new_[7716]_  = ~A166 & \new_[7715]_ ;
  assign \new_[7717]_  = \new_[7716]_  & \new_[7711]_ ;
  assign \new_[7720]_  = A267 & A266;
  assign \new_[7724]_  = ~A301 & ~A299;
  assign \new_[7725]_  = ~A298 & \new_[7724]_ ;
  assign \new_[7726]_  = \new_[7725]_  & \new_[7720]_ ;
  assign \new_[7729]_  = A167 & A170;
  assign \new_[7733]_  = A201 & A200;
  assign \new_[7734]_  = ~A166 & \new_[7733]_ ;
  assign \new_[7735]_  = \new_[7734]_  & \new_[7729]_ ;
  assign \new_[7738]_  = A298 & A268;
  assign \new_[7742]_  = ~A301 & ~A300;
  assign \new_[7743]_  = A299 & \new_[7742]_ ;
  assign \new_[7744]_  = \new_[7743]_  & \new_[7738]_ ;
  assign \new_[7747]_  = A167 & A170;
  assign \new_[7751]_  = A201 & A200;
  assign \new_[7752]_  = ~A166 & \new_[7751]_ ;
  assign \new_[7753]_  = \new_[7752]_  & \new_[7747]_ ;
  assign \new_[7756]_  = A267 & A265;
  assign \new_[7760]_  = ~A302 & ~A301;
  assign \new_[7761]_  = ~A300 & \new_[7760]_ ;
  assign \new_[7762]_  = \new_[7761]_  & \new_[7756]_ ;
  assign \new_[7765]_  = A167 & A170;
  assign \new_[7769]_  = A201 & A200;
  assign \new_[7770]_  = ~A166 & \new_[7769]_ ;
  assign \new_[7771]_  = \new_[7770]_  & \new_[7765]_ ;
  assign \new_[7774]_  = A267 & A265;
  assign \new_[7778]_  = ~A301 & ~A299;
  assign \new_[7779]_  = ~A298 & \new_[7778]_ ;
  assign \new_[7780]_  = \new_[7779]_  & \new_[7774]_ ;
  assign \new_[7783]_  = A167 & A170;
  assign \new_[7787]_  = A201 & A200;
  assign \new_[7788]_  = ~A166 & \new_[7787]_ ;
  assign \new_[7789]_  = \new_[7788]_  & \new_[7783]_ ;
  assign \new_[7792]_  = A267 & A266;
  assign \new_[7796]_  = ~A302 & ~A301;
  assign \new_[7797]_  = ~A300 & \new_[7796]_ ;
  assign \new_[7798]_  = \new_[7797]_  & \new_[7792]_ ;
  assign \new_[7801]_  = A167 & A170;
  assign \new_[7805]_  = A201 & A200;
  assign \new_[7806]_  = ~A166 & \new_[7805]_ ;
  assign \new_[7807]_  = \new_[7806]_  & \new_[7801]_ ;
  assign \new_[7810]_  = A267 & A266;
  assign \new_[7814]_  = ~A301 & ~A299;
  assign \new_[7815]_  = ~A298 & \new_[7814]_ ;
  assign \new_[7816]_  = \new_[7815]_  & \new_[7810]_ ;
  assign \new_[7819]_  = A167 & A170;
  assign \new_[7823]_  = A200 & ~A199;
  assign \new_[7824]_  = ~A166 & \new_[7823]_ ;
  assign \new_[7825]_  = \new_[7824]_  & \new_[7819]_ ;
  assign \new_[7828]_  = A268 & A203;
  assign \new_[7832]_  = ~A302 & ~A301;
  assign \new_[7833]_  = ~A300 & \new_[7832]_ ;
  assign \new_[7834]_  = \new_[7833]_  & \new_[7828]_ ;
  assign \new_[7837]_  = A167 & A170;
  assign \new_[7841]_  = A200 & ~A199;
  assign \new_[7842]_  = ~A166 & \new_[7841]_ ;
  assign \new_[7843]_  = \new_[7842]_  & \new_[7837]_ ;
  assign \new_[7846]_  = A268 & A203;
  assign \new_[7850]_  = ~A301 & ~A299;
  assign \new_[7851]_  = ~A298 & \new_[7850]_ ;
  assign \new_[7852]_  = \new_[7851]_  & \new_[7846]_ ;
  assign \new_[7855]_  = A167 & A170;
  assign \new_[7859]_  = ~A200 & A199;
  assign \new_[7860]_  = ~A166 & \new_[7859]_ ;
  assign \new_[7861]_  = \new_[7860]_  & \new_[7855]_ ;
  assign \new_[7864]_  = A268 & A203;
  assign \new_[7868]_  = ~A302 & ~A301;
  assign \new_[7869]_  = ~A300 & \new_[7868]_ ;
  assign \new_[7870]_  = \new_[7869]_  & \new_[7864]_ ;
  assign \new_[7873]_  = A167 & A170;
  assign \new_[7877]_  = ~A200 & A199;
  assign \new_[7878]_  = ~A166 & \new_[7877]_ ;
  assign \new_[7879]_  = \new_[7878]_  & \new_[7873]_ ;
  assign \new_[7882]_  = A268 & A203;
  assign \new_[7886]_  = ~A301 & ~A299;
  assign \new_[7887]_  = ~A298 & \new_[7886]_ ;
  assign \new_[7888]_  = \new_[7887]_  & \new_[7882]_ ;
  assign \new_[7891]_  = A167 & A170;
  assign \new_[7895]_  = ~A200 & ~A199;
  assign \new_[7896]_  = ~A166 & \new_[7895]_ ;
  assign \new_[7897]_  = \new_[7896]_  & \new_[7891]_ ;
  assign \new_[7900]_  = ~A267 & ~A202;
  assign \new_[7904]_  = A301 & ~A269;
  assign \new_[7905]_  = ~A268 & \new_[7904]_ ;
  assign \new_[7906]_  = \new_[7905]_  & \new_[7900]_ ;
  assign \new_[7909]_  = A167 & A170;
  assign \new_[7913]_  = ~A200 & ~A199;
  assign \new_[7914]_  = ~A166 & \new_[7913]_ ;
  assign \new_[7915]_  = \new_[7914]_  & \new_[7909]_ ;
  assign \new_[7918]_  = ~A265 & ~A202;
  assign \new_[7922]_  = A301 & ~A268;
  assign \new_[7923]_  = ~A266 & \new_[7922]_ ;
  assign \new_[7924]_  = \new_[7923]_  & \new_[7918]_ ;
  assign \new_[7927]_  = ~A167 & A170;
  assign \new_[7931]_  = A265 & A202;
  assign \new_[7932]_  = A166 & \new_[7931]_ ;
  assign \new_[7933]_  = \new_[7932]_  & \new_[7927]_ ;
  assign \new_[7936]_  = A298 & A267;
  assign \new_[7940]_  = ~A301 & ~A300;
  assign \new_[7941]_  = A299 & \new_[7940]_ ;
  assign \new_[7942]_  = \new_[7941]_  & \new_[7936]_ ;
  assign \new_[7945]_  = ~A167 & A170;
  assign \new_[7949]_  = A266 & A202;
  assign \new_[7950]_  = A166 & \new_[7949]_ ;
  assign \new_[7951]_  = \new_[7950]_  & \new_[7945]_ ;
  assign \new_[7954]_  = A298 & A267;
  assign \new_[7958]_  = ~A301 & ~A300;
  assign \new_[7959]_  = A299 & \new_[7958]_ ;
  assign \new_[7960]_  = \new_[7959]_  & \new_[7954]_ ;
  assign \new_[7963]_  = ~A167 & A170;
  assign \new_[7967]_  = ~A265 & A202;
  assign \new_[7968]_  = A166 & \new_[7967]_ ;
  assign \new_[7969]_  = \new_[7968]_  & \new_[7963]_ ;
  assign \new_[7972]_  = A269 & A266;
  assign \new_[7976]_  = ~A302 & ~A301;
  assign \new_[7977]_  = ~A300 & \new_[7976]_ ;
  assign \new_[7978]_  = \new_[7977]_  & \new_[7972]_ ;
  assign \new_[7981]_  = ~A167 & A170;
  assign \new_[7985]_  = ~A265 & A202;
  assign \new_[7986]_  = A166 & \new_[7985]_ ;
  assign \new_[7987]_  = \new_[7986]_  & \new_[7981]_ ;
  assign \new_[7990]_  = A269 & A266;
  assign \new_[7994]_  = ~A301 & ~A299;
  assign \new_[7995]_  = ~A298 & \new_[7994]_ ;
  assign \new_[7996]_  = \new_[7995]_  & \new_[7990]_ ;
  assign \new_[7999]_  = ~A167 & A170;
  assign \new_[8003]_  = A265 & A202;
  assign \new_[8004]_  = A166 & \new_[8003]_ ;
  assign \new_[8005]_  = \new_[8004]_  & \new_[7999]_ ;
  assign \new_[8008]_  = A269 & ~A266;
  assign \new_[8012]_  = ~A302 & ~A301;
  assign \new_[8013]_  = ~A300 & \new_[8012]_ ;
  assign \new_[8014]_  = \new_[8013]_  & \new_[8008]_ ;
  assign \new_[8017]_  = ~A167 & A170;
  assign \new_[8021]_  = A265 & A202;
  assign \new_[8022]_  = A166 & \new_[8021]_ ;
  assign \new_[8023]_  = \new_[8022]_  & \new_[8017]_ ;
  assign \new_[8026]_  = A269 & ~A266;
  assign \new_[8030]_  = ~A301 & ~A299;
  assign \new_[8031]_  = ~A298 & \new_[8030]_ ;
  assign \new_[8032]_  = \new_[8031]_  & \new_[8026]_ ;
  assign \new_[8035]_  = ~A167 & A170;
  assign \new_[8039]_  = ~A202 & ~A201;
  assign \new_[8040]_  = A166 & \new_[8039]_ ;
  assign \new_[8041]_  = \new_[8040]_  & \new_[8035]_ ;
  assign \new_[8044]_  = ~A267 & ~A203;
  assign \new_[8048]_  = A301 & ~A269;
  assign \new_[8049]_  = ~A268 & \new_[8048]_ ;
  assign \new_[8050]_  = \new_[8049]_  & \new_[8044]_ ;
  assign \new_[8053]_  = ~A167 & A170;
  assign \new_[8057]_  = ~A202 & ~A201;
  assign \new_[8058]_  = A166 & \new_[8057]_ ;
  assign \new_[8059]_  = \new_[8058]_  & \new_[8053]_ ;
  assign \new_[8062]_  = ~A265 & ~A203;
  assign \new_[8066]_  = A301 & ~A268;
  assign \new_[8067]_  = ~A266 & \new_[8066]_ ;
  assign \new_[8068]_  = \new_[8067]_  & \new_[8062]_ ;
  assign \new_[8071]_  = ~A167 & A170;
  assign \new_[8075]_  = A201 & A199;
  assign \new_[8076]_  = A166 & \new_[8075]_ ;
  assign \new_[8077]_  = \new_[8076]_  & \new_[8071]_ ;
  assign \new_[8080]_  = A298 & A268;
  assign \new_[8084]_  = ~A301 & ~A300;
  assign \new_[8085]_  = A299 & \new_[8084]_ ;
  assign \new_[8086]_  = \new_[8085]_  & \new_[8080]_ ;
  assign \new_[8089]_  = ~A167 & A170;
  assign \new_[8093]_  = A201 & A199;
  assign \new_[8094]_  = A166 & \new_[8093]_ ;
  assign \new_[8095]_  = \new_[8094]_  & \new_[8089]_ ;
  assign \new_[8098]_  = A267 & A265;
  assign \new_[8102]_  = ~A302 & ~A301;
  assign \new_[8103]_  = ~A300 & \new_[8102]_ ;
  assign \new_[8104]_  = \new_[8103]_  & \new_[8098]_ ;
  assign \new_[8107]_  = ~A167 & A170;
  assign \new_[8111]_  = A201 & A199;
  assign \new_[8112]_  = A166 & \new_[8111]_ ;
  assign \new_[8113]_  = \new_[8112]_  & \new_[8107]_ ;
  assign \new_[8116]_  = A267 & A265;
  assign \new_[8120]_  = ~A301 & ~A299;
  assign \new_[8121]_  = ~A298 & \new_[8120]_ ;
  assign \new_[8122]_  = \new_[8121]_  & \new_[8116]_ ;
  assign \new_[8125]_  = ~A167 & A170;
  assign \new_[8129]_  = A201 & A199;
  assign \new_[8130]_  = A166 & \new_[8129]_ ;
  assign \new_[8131]_  = \new_[8130]_  & \new_[8125]_ ;
  assign \new_[8134]_  = A267 & A266;
  assign \new_[8138]_  = ~A302 & ~A301;
  assign \new_[8139]_  = ~A300 & \new_[8138]_ ;
  assign \new_[8140]_  = \new_[8139]_  & \new_[8134]_ ;
  assign \new_[8143]_  = ~A167 & A170;
  assign \new_[8147]_  = A201 & A199;
  assign \new_[8148]_  = A166 & \new_[8147]_ ;
  assign \new_[8149]_  = \new_[8148]_  & \new_[8143]_ ;
  assign \new_[8152]_  = A267 & A266;
  assign \new_[8156]_  = ~A301 & ~A299;
  assign \new_[8157]_  = ~A298 & \new_[8156]_ ;
  assign \new_[8158]_  = \new_[8157]_  & \new_[8152]_ ;
  assign \new_[8161]_  = ~A167 & A170;
  assign \new_[8165]_  = A201 & A200;
  assign \new_[8166]_  = A166 & \new_[8165]_ ;
  assign \new_[8167]_  = \new_[8166]_  & \new_[8161]_ ;
  assign \new_[8170]_  = A298 & A268;
  assign \new_[8174]_  = ~A301 & ~A300;
  assign \new_[8175]_  = A299 & \new_[8174]_ ;
  assign \new_[8176]_  = \new_[8175]_  & \new_[8170]_ ;
  assign \new_[8179]_  = ~A167 & A170;
  assign \new_[8183]_  = A201 & A200;
  assign \new_[8184]_  = A166 & \new_[8183]_ ;
  assign \new_[8185]_  = \new_[8184]_  & \new_[8179]_ ;
  assign \new_[8188]_  = A267 & A265;
  assign \new_[8192]_  = ~A302 & ~A301;
  assign \new_[8193]_  = ~A300 & \new_[8192]_ ;
  assign \new_[8194]_  = \new_[8193]_  & \new_[8188]_ ;
  assign \new_[8197]_  = ~A167 & A170;
  assign \new_[8201]_  = A201 & A200;
  assign \new_[8202]_  = A166 & \new_[8201]_ ;
  assign \new_[8203]_  = \new_[8202]_  & \new_[8197]_ ;
  assign \new_[8206]_  = A267 & A265;
  assign \new_[8210]_  = ~A301 & ~A299;
  assign \new_[8211]_  = ~A298 & \new_[8210]_ ;
  assign \new_[8212]_  = \new_[8211]_  & \new_[8206]_ ;
  assign \new_[8215]_  = ~A167 & A170;
  assign \new_[8219]_  = A201 & A200;
  assign \new_[8220]_  = A166 & \new_[8219]_ ;
  assign \new_[8221]_  = \new_[8220]_  & \new_[8215]_ ;
  assign \new_[8224]_  = A267 & A266;
  assign \new_[8228]_  = ~A302 & ~A301;
  assign \new_[8229]_  = ~A300 & \new_[8228]_ ;
  assign \new_[8230]_  = \new_[8229]_  & \new_[8224]_ ;
  assign \new_[8233]_  = ~A167 & A170;
  assign \new_[8237]_  = A201 & A200;
  assign \new_[8238]_  = A166 & \new_[8237]_ ;
  assign \new_[8239]_  = \new_[8238]_  & \new_[8233]_ ;
  assign \new_[8242]_  = A267 & A266;
  assign \new_[8246]_  = ~A301 & ~A299;
  assign \new_[8247]_  = ~A298 & \new_[8246]_ ;
  assign \new_[8248]_  = \new_[8247]_  & \new_[8242]_ ;
  assign \new_[8251]_  = ~A167 & A170;
  assign \new_[8255]_  = A200 & ~A199;
  assign \new_[8256]_  = A166 & \new_[8255]_ ;
  assign \new_[8257]_  = \new_[8256]_  & \new_[8251]_ ;
  assign \new_[8260]_  = A268 & A203;
  assign \new_[8264]_  = ~A302 & ~A301;
  assign \new_[8265]_  = ~A300 & \new_[8264]_ ;
  assign \new_[8266]_  = \new_[8265]_  & \new_[8260]_ ;
  assign \new_[8269]_  = ~A167 & A170;
  assign \new_[8273]_  = A200 & ~A199;
  assign \new_[8274]_  = A166 & \new_[8273]_ ;
  assign \new_[8275]_  = \new_[8274]_  & \new_[8269]_ ;
  assign \new_[8278]_  = A268 & A203;
  assign \new_[8282]_  = ~A301 & ~A299;
  assign \new_[8283]_  = ~A298 & \new_[8282]_ ;
  assign \new_[8284]_  = \new_[8283]_  & \new_[8278]_ ;
  assign \new_[8287]_  = ~A167 & A170;
  assign \new_[8291]_  = ~A200 & A199;
  assign \new_[8292]_  = A166 & \new_[8291]_ ;
  assign \new_[8293]_  = \new_[8292]_  & \new_[8287]_ ;
  assign \new_[8296]_  = A268 & A203;
  assign \new_[8300]_  = ~A302 & ~A301;
  assign \new_[8301]_  = ~A300 & \new_[8300]_ ;
  assign \new_[8302]_  = \new_[8301]_  & \new_[8296]_ ;
  assign \new_[8305]_  = ~A167 & A170;
  assign \new_[8309]_  = ~A200 & A199;
  assign \new_[8310]_  = A166 & \new_[8309]_ ;
  assign \new_[8311]_  = \new_[8310]_  & \new_[8305]_ ;
  assign \new_[8314]_  = A268 & A203;
  assign \new_[8318]_  = ~A301 & ~A299;
  assign \new_[8319]_  = ~A298 & \new_[8318]_ ;
  assign \new_[8320]_  = \new_[8319]_  & \new_[8314]_ ;
  assign \new_[8323]_  = ~A167 & A170;
  assign \new_[8327]_  = ~A200 & ~A199;
  assign \new_[8328]_  = A166 & \new_[8327]_ ;
  assign \new_[8329]_  = \new_[8328]_  & \new_[8323]_ ;
  assign \new_[8332]_  = ~A267 & ~A202;
  assign \new_[8336]_  = A301 & ~A269;
  assign \new_[8337]_  = ~A268 & \new_[8336]_ ;
  assign \new_[8338]_  = \new_[8337]_  & \new_[8332]_ ;
  assign \new_[8341]_  = ~A167 & A170;
  assign \new_[8345]_  = ~A200 & ~A199;
  assign \new_[8346]_  = A166 & \new_[8345]_ ;
  assign \new_[8347]_  = \new_[8346]_  & \new_[8341]_ ;
  assign \new_[8350]_  = ~A265 & ~A202;
  assign \new_[8354]_  = A301 & ~A268;
  assign \new_[8355]_  = ~A266 & \new_[8354]_ ;
  assign \new_[8356]_  = \new_[8355]_  & \new_[8350]_ ;
  assign \new_[8359]_  = ~A201 & A169;
  assign \new_[8363]_  = ~A267 & ~A203;
  assign \new_[8364]_  = ~A202 & \new_[8363]_ ;
  assign \new_[8365]_  = \new_[8364]_  & \new_[8359]_ ;
  assign \new_[8368]_  = ~A269 & ~A268;
  assign \new_[8372]_  = A302 & ~A299;
  assign \new_[8373]_  = A298 & \new_[8372]_ ;
  assign \new_[8374]_  = \new_[8373]_  & \new_[8368]_ ;
  assign \new_[8377]_  = ~A201 & A169;
  assign \new_[8381]_  = ~A267 & ~A203;
  assign \new_[8382]_  = ~A202 & \new_[8381]_ ;
  assign \new_[8383]_  = \new_[8382]_  & \new_[8377]_ ;
  assign \new_[8386]_  = ~A269 & ~A268;
  assign \new_[8390]_  = A302 & A299;
  assign \new_[8391]_  = ~A298 & \new_[8390]_ ;
  assign \new_[8392]_  = \new_[8391]_  & \new_[8386]_ ;
  assign \new_[8395]_  = ~A201 & A169;
  assign \new_[8399]_  = A265 & ~A203;
  assign \new_[8400]_  = ~A202 & \new_[8399]_ ;
  assign \new_[8401]_  = \new_[8400]_  & \new_[8395]_ ;
  assign \new_[8404]_  = ~A267 & A266;
  assign \new_[8408]_  = A300 & A299;
  assign \new_[8409]_  = ~A268 & \new_[8408]_ ;
  assign \new_[8410]_  = \new_[8409]_  & \new_[8404]_ ;
  assign \new_[8413]_  = ~A201 & A169;
  assign \new_[8417]_  = A265 & ~A203;
  assign \new_[8418]_  = ~A202 & \new_[8417]_ ;
  assign \new_[8419]_  = \new_[8418]_  & \new_[8413]_ ;
  assign \new_[8422]_  = ~A267 & A266;
  assign \new_[8426]_  = A300 & A298;
  assign \new_[8427]_  = ~A268 & \new_[8426]_ ;
  assign \new_[8428]_  = \new_[8427]_  & \new_[8422]_ ;
  assign \new_[8431]_  = ~A201 & A169;
  assign \new_[8435]_  = ~A265 & ~A203;
  assign \new_[8436]_  = ~A202 & \new_[8435]_ ;
  assign \new_[8437]_  = \new_[8436]_  & \new_[8431]_ ;
  assign \new_[8440]_  = ~A268 & ~A266;
  assign \new_[8444]_  = A302 & ~A299;
  assign \new_[8445]_  = A298 & \new_[8444]_ ;
  assign \new_[8446]_  = \new_[8445]_  & \new_[8440]_ ;
  assign \new_[8449]_  = ~A201 & A169;
  assign \new_[8453]_  = ~A265 & ~A203;
  assign \new_[8454]_  = ~A202 & \new_[8453]_ ;
  assign \new_[8455]_  = \new_[8454]_  & \new_[8449]_ ;
  assign \new_[8458]_  = ~A268 & ~A266;
  assign \new_[8462]_  = A302 & A299;
  assign \new_[8463]_  = ~A298 & \new_[8462]_ ;
  assign \new_[8464]_  = \new_[8463]_  & \new_[8458]_ ;
  assign \new_[8467]_  = A199 & A169;
  assign \new_[8471]_  = A266 & ~A265;
  assign \new_[8472]_  = A201 & \new_[8471]_ ;
  assign \new_[8473]_  = \new_[8472]_  & \new_[8467]_ ;
  assign \new_[8476]_  = A298 & A269;
  assign \new_[8480]_  = ~A301 & ~A300;
  assign \new_[8481]_  = A299 & \new_[8480]_ ;
  assign \new_[8482]_  = \new_[8481]_  & \new_[8476]_ ;
  assign \new_[8485]_  = A199 & A169;
  assign \new_[8489]_  = ~A266 & A265;
  assign \new_[8490]_  = A201 & \new_[8489]_ ;
  assign \new_[8491]_  = \new_[8490]_  & \new_[8485]_ ;
  assign \new_[8494]_  = A298 & A269;
  assign \new_[8498]_  = ~A301 & ~A300;
  assign \new_[8499]_  = A299 & \new_[8498]_ ;
  assign \new_[8500]_  = \new_[8499]_  & \new_[8494]_ ;
  assign \new_[8503]_  = A200 & A169;
  assign \new_[8507]_  = A266 & ~A265;
  assign \new_[8508]_  = A201 & \new_[8507]_ ;
  assign \new_[8509]_  = \new_[8508]_  & \new_[8503]_ ;
  assign \new_[8512]_  = A298 & A269;
  assign \new_[8516]_  = ~A301 & ~A300;
  assign \new_[8517]_  = A299 & \new_[8516]_ ;
  assign \new_[8518]_  = \new_[8517]_  & \new_[8512]_ ;
  assign \new_[8521]_  = A200 & A169;
  assign \new_[8525]_  = ~A266 & A265;
  assign \new_[8526]_  = A201 & \new_[8525]_ ;
  assign \new_[8527]_  = \new_[8526]_  & \new_[8521]_ ;
  assign \new_[8530]_  = A298 & A269;
  assign \new_[8534]_  = ~A301 & ~A300;
  assign \new_[8535]_  = A299 & \new_[8534]_ ;
  assign \new_[8536]_  = \new_[8535]_  & \new_[8530]_ ;
  assign \new_[8539]_  = A199 & A169;
  assign \new_[8543]_  = ~A202 & ~A201;
  assign \new_[8544]_  = A200 & \new_[8543]_ ;
  assign \new_[8545]_  = \new_[8544]_  & \new_[8539]_ ;
  assign \new_[8548]_  = ~A268 & ~A267;
  assign \new_[8552]_  = A300 & A299;
  assign \new_[8553]_  = ~A269 & \new_[8552]_ ;
  assign \new_[8554]_  = \new_[8553]_  & \new_[8548]_ ;
  assign \new_[8557]_  = A199 & A169;
  assign \new_[8561]_  = ~A202 & ~A201;
  assign \new_[8562]_  = A200 & \new_[8561]_ ;
  assign \new_[8563]_  = \new_[8562]_  & \new_[8557]_ ;
  assign \new_[8566]_  = ~A268 & ~A267;
  assign \new_[8570]_  = A300 & A298;
  assign \new_[8571]_  = ~A269 & \new_[8570]_ ;
  assign \new_[8572]_  = \new_[8571]_  & \new_[8566]_ ;
  assign \new_[8575]_  = A199 & A169;
  assign \new_[8579]_  = ~A202 & ~A201;
  assign \new_[8580]_  = A200 & \new_[8579]_ ;
  assign \new_[8581]_  = \new_[8580]_  & \new_[8575]_ ;
  assign \new_[8584]_  = A266 & A265;
  assign \new_[8588]_  = A301 & ~A268;
  assign \new_[8589]_  = ~A267 & \new_[8588]_ ;
  assign \new_[8590]_  = \new_[8589]_  & \new_[8584]_ ;
  assign \new_[8593]_  = A199 & A169;
  assign \new_[8597]_  = ~A202 & ~A201;
  assign \new_[8598]_  = A200 & \new_[8597]_ ;
  assign \new_[8599]_  = \new_[8598]_  & \new_[8593]_ ;
  assign \new_[8602]_  = ~A266 & ~A265;
  assign \new_[8606]_  = A300 & A299;
  assign \new_[8607]_  = ~A268 & \new_[8606]_ ;
  assign \new_[8608]_  = \new_[8607]_  & \new_[8602]_ ;
  assign \new_[8611]_  = A199 & A169;
  assign \new_[8615]_  = ~A202 & ~A201;
  assign \new_[8616]_  = A200 & \new_[8615]_ ;
  assign \new_[8617]_  = \new_[8616]_  & \new_[8611]_ ;
  assign \new_[8620]_  = ~A266 & ~A265;
  assign \new_[8624]_  = A300 & A298;
  assign \new_[8625]_  = ~A268 & \new_[8624]_ ;
  assign \new_[8626]_  = \new_[8625]_  & \new_[8620]_ ;
  assign \new_[8629]_  = ~A199 & A169;
  assign \new_[8633]_  = A265 & A203;
  assign \new_[8634]_  = A200 & \new_[8633]_ ;
  assign \new_[8635]_  = \new_[8634]_  & \new_[8629]_ ;
  assign \new_[8638]_  = A298 & A267;
  assign \new_[8642]_  = ~A301 & ~A300;
  assign \new_[8643]_  = A299 & \new_[8642]_ ;
  assign \new_[8644]_  = \new_[8643]_  & \new_[8638]_ ;
  assign \new_[8647]_  = ~A199 & A169;
  assign \new_[8651]_  = A266 & A203;
  assign \new_[8652]_  = A200 & \new_[8651]_ ;
  assign \new_[8653]_  = \new_[8652]_  & \new_[8647]_ ;
  assign \new_[8656]_  = A298 & A267;
  assign \new_[8660]_  = ~A301 & ~A300;
  assign \new_[8661]_  = A299 & \new_[8660]_ ;
  assign \new_[8662]_  = \new_[8661]_  & \new_[8656]_ ;
  assign \new_[8665]_  = ~A199 & A169;
  assign \new_[8669]_  = ~A265 & A203;
  assign \new_[8670]_  = A200 & \new_[8669]_ ;
  assign \new_[8671]_  = \new_[8670]_  & \new_[8665]_ ;
  assign \new_[8674]_  = A269 & A266;
  assign \new_[8678]_  = ~A302 & ~A301;
  assign \new_[8679]_  = ~A300 & \new_[8678]_ ;
  assign \new_[8680]_  = \new_[8679]_  & \new_[8674]_ ;
  assign \new_[8683]_  = ~A199 & A169;
  assign \new_[8687]_  = ~A265 & A203;
  assign \new_[8688]_  = A200 & \new_[8687]_ ;
  assign \new_[8689]_  = \new_[8688]_  & \new_[8683]_ ;
  assign \new_[8692]_  = A269 & A266;
  assign \new_[8696]_  = ~A301 & ~A299;
  assign \new_[8697]_  = ~A298 & \new_[8696]_ ;
  assign \new_[8698]_  = \new_[8697]_  & \new_[8692]_ ;
  assign \new_[8701]_  = ~A199 & A169;
  assign \new_[8705]_  = A265 & A203;
  assign \new_[8706]_  = A200 & \new_[8705]_ ;
  assign \new_[8707]_  = \new_[8706]_  & \new_[8701]_ ;
  assign \new_[8710]_  = A269 & ~A266;
  assign \new_[8714]_  = ~A302 & ~A301;
  assign \new_[8715]_  = ~A300 & \new_[8714]_ ;
  assign \new_[8716]_  = \new_[8715]_  & \new_[8710]_ ;
  assign \new_[8719]_  = ~A199 & A169;
  assign \new_[8723]_  = A265 & A203;
  assign \new_[8724]_  = A200 & \new_[8723]_ ;
  assign \new_[8725]_  = \new_[8724]_  & \new_[8719]_ ;
  assign \new_[8728]_  = A269 & ~A266;
  assign \new_[8732]_  = ~A301 & ~A299;
  assign \new_[8733]_  = ~A298 & \new_[8732]_ ;
  assign \new_[8734]_  = \new_[8733]_  & \new_[8728]_ ;
  assign \new_[8737]_  = A199 & A169;
  assign \new_[8741]_  = A265 & A203;
  assign \new_[8742]_  = ~A200 & \new_[8741]_ ;
  assign \new_[8743]_  = \new_[8742]_  & \new_[8737]_ ;
  assign \new_[8746]_  = A298 & A267;
  assign \new_[8750]_  = ~A301 & ~A300;
  assign \new_[8751]_  = A299 & \new_[8750]_ ;
  assign \new_[8752]_  = \new_[8751]_  & \new_[8746]_ ;
  assign \new_[8755]_  = A199 & A169;
  assign \new_[8759]_  = A266 & A203;
  assign \new_[8760]_  = ~A200 & \new_[8759]_ ;
  assign \new_[8761]_  = \new_[8760]_  & \new_[8755]_ ;
  assign \new_[8764]_  = A298 & A267;
  assign \new_[8768]_  = ~A301 & ~A300;
  assign \new_[8769]_  = A299 & \new_[8768]_ ;
  assign \new_[8770]_  = \new_[8769]_  & \new_[8764]_ ;
  assign \new_[8773]_  = A199 & A169;
  assign \new_[8777]_  = ~A265 & A203;
  assign \new_[8778]_  = ~A200 & \new_[8777]_ ;
  assign \new_[8779]_  = \new_[8778]_  & \new_[8773]_ ;
  assign \new_[8782]_  = A269 & A266;
  assign \new_[8786]_  = ~A302 & ~A301;
  assign \new_[8787]_  = ~A300 & \new_[8786]_ ;
  assign \new_[8788]_  = \new_[8787]_  & \new_[8782]_ ;
  assign \new_[8791]_  = A199 & A169;
  assign \new_[8795]_  = ~A265 & A203;
  assign \new_[8796]_  = ~A200 & \new_[8795]_ ;
  assign \new_[8797]_  = \new_[8796]_  & \new_[8791]_ ;
  assign \new_[8800]_  = A269 & A266;
  assign \new_[8804]_  = ~A301 & ~A299;
  assign \new_[8805]_  = ~A298 & \new_[8804]_ ;
  assign \new_[8806]_  = \new_[8805]_  & \new_[8800]_ ;
  assign \new_[8809]_  = A199 & A169;
  assign \new_[8813]_  = A265 & A203;
  assign \new_[8814]_  = ~A200 & \new_[8813]_ ;
  assign \new_[8815]_  = \new_[8814]_  & \new_[8809]_ ;
  assign \new_[8818]_  = A269 & ~A266;
  assign \new_[8822]_  = ~A302 & ~A301;
  assign \new_[8823]_  = ~A300 & \new_[8822]_ ;
  assign \new_[8824]_  = \new_[8823]_  & \new_[8818]_ ;
  assign \new_[8827]_  = A199 & A169;
  assign \new_[8831]_  = A265 & A203;
  assign \new_[8832]_  = ~A200 & \new_[8831]_ ;
  assign \new_[8833]_  = \new_[8832]_  & \new_[8827]_ ;
  assign \new_[8836]_  = A269 & ~A266;
  assign \new_[8840]_  = ~A301 & ~A299;
  assign \new_[8841]_  = ~A298 & \new_[8840]_ ;
  assign \new_[8842]_  = \new_[8841]_  & \new_[8836]_ ;
  assign \new_[8845]_  = ~A199 & A169;
  assign \new_[8849]_  = ~A267 & ~A202;
  assign \new_[8850]_  = ~A200 & \new_[8849]_ ;
  assign \new_[8851]_  = \new_[8850]_  & \new_[8845]_ ;
  assign \new_[8854]_  = ~A269 & ~A268;
  assign \new_[8858]_  = A302 & ~A299;
  assign \new_[8859]_  = A298 & \new_[8858]_ ;
  assign \new_[8860]_  = \new_[8859]_  & \new_[8854]_ ;
  assign \new_[8863]_  = ~A199 & A169;
  assign \new_[8867]_  = ~A267 & ~A202;
  assign \new_[8868]_  = ~A200 & \new_[8867]_ ;
  assign \new_[8869]_  = \new_[8868]_  & \new_[8863]_ ;
  assign \new_[8872]_  = ~A269 & ~A268;
  assign \new_[8876]_  = A302 & A299;
  assign \new_[8877]_  = ~A298 & \new_[8876]_ ;
  assign \new_[8878]_  = \new_[8877]_  & \new_[8872]_ ;
  assign \new_[8881]_  = ~A199 & A169;
  assign \new_[8885]_  = A265 & ~A202;
  assign \new_[8886]_  = ~A200 & \new_[8885]_ ;
  assign \new_[8887]_  = \new_[8886]_  & \new_[8881]_ ;
  assign \new_[8890]_  = ~A267 & A266;
  assign \new_[8894]_  = A300 & A299;
  assign \new_[8895]_  = ~A268 & \new_[8894]_ ;
  assign \new_[8896]_  = \new_[8895]_  & \new_[8890]_ ;
  assign \new_[8899]_  = ~A199 & A169;
  assign \new_[8903]_  = A265 & ~A202;
  assign \new_[8904]_  = ~A200 & \new_[8903]_ ;
  assign \new_[8905]_  = \new_[8904]_  & \new_[8899]_ ;
  assign \new_[8908]_  = ~A267 & A266;
  assign \new_[8912]_  = A300 & A298;
  assign \new_[8913]_  = ~A268 & \new_[8912]_ ;
  assign \new_[8914]_  = \new_[8913]_  & \new_[8908]_ ;
  assign \new_[8917]_  = ~A199 & A169;
  assign \new_[8921]_  = ~A265 & ~A202;
  assign \new_[8922]_  = ~A200 & \new_[8921]_ ;
  assign \new_[8923]_  = \new_[8922]_  & \new_[8917]_ ;
  assign \new_[8926]_  = ~A268 & ~A266;
  assign \new_[8930]_  = A302 & ~A299;
  assign \new_[8931]_  = A298 & \new_[8930]_ ;
  assign \new_[8932]_  = \new_[8931]_  & \new_[8926]_ ;
  assign \new_[8935]_  = ~A199 & A169;
  assign \new_[8939]_  = ~A265 & ~A202;
  assign \new_[8940]_  = ~A200 & \new_[8939]_ ;
  assign \new_[8941]_  = \new_[8940]_  & \new_[8935]_ ;
  assign \new_[8944]_  = ~A268 & ~A266;
  assign \new_[8948]_  = A302 & A299;
  assign \new_[8949]_  = ~A298 & \new_[8948]_ ;
  assign \new_[8950]_  = \new_[8949]_  & \new_[8944]_ ;
  assign \new_[8953]_  = ~A167 & ~A169;
  assign \new_[8957]_  = ~A267 & A202;
  assign \new_[8958]_  = ~A166 & \new_[8957]_ ;
  assign \new_[8959]_  = \new_[8958]_  & \new_[8953]_ ;
  assign \new_[8962]_  = ~A269 & ~A268;
  assign \new_[8966]_  = A302 & ~A299;
  assign \new_[8967]_  = A298 & \new_[8966]_ ;
  assign \new_[8968]_  = \new_[8967]_  & \new_[8962]_ ;
  assign \new_[8971]_  = ~A167 & ~A169;
  assign \new_[8975]_  = ~A267 & A202;
  assign \new_[8976]_  = ~A166 & \new_[8975]_ ;
  assign \new_[8977]_  = \new_[8976]_  & \new_[8971]_ ;
  assign \new_[8980]_  = ~A269 & ~A268;
  assign \new_[8984]_  = A302 & A299;
  assign \new_[8985]_  = ~A298 & \new_[8984]_ ;
  assign \new_[8986]_  = \new_[8985]_  & \new_[8980]_ ;
  assign \new_[8989]_  = ~A167 & ~A169;
  assign \new_[8993]_  = A265 & A202;
  assign \new_[8994]_  = ~A166 & \new_[8993]_ ;
  assign \new_[8995]_  = \new_[8994]_  & \new_[8989]_ ;
  assign \new_[8998]_  = ~A267 & A266;
  assign \new_[9002]_  = A300 & A299;
  assign \new_[9003]_  = ~A268 & \new_[9002]_ ;
  assign \new_[9004]_  = \new_[9003]_  & \new_[8998]_ ;
  assign \new_[9007]_  = ~A167 & ~A169;
  assign \new_[9011]_  = A265 & A202;
  assign \new_[9012]_  = ~A166 & \new_[9011]_ ;
  assign \new_[9013]_  = \new_[9012]_  & \new_[9007]_ ;
  assign \new_[9016]_  = ~A267 & A266;
  assign \new_[9020]_  = A300 & A298;
  assign \new_[9021]_  = ~A268 & \new_[9020]_ ;
  assign \new_[9022]_  = \new_[9021]_  & \new_[9016]_ ;
  assign \new_[9025]_  = ~A167 & ~A169;
  assign \new_[9029]_  = ~A265 & A202;
  assign \new_[9030]_  = ~A166 & \new_[9029]_ ;
  assign \new_[9031]_  = \new_[9030]_  & \new_[9025]_ ;
  assign \new_[9034]_  = ~A268 & ~A266;
  assign \new_[9038]_  = A302 & ~A299;
  assign \new_[9039]_  = A298 & \new_[9038]_ ;
  assign \new_[9040]_  = \new_[9039]_  & \new_[9034]_ ;
  assign \new_[9043]_  = ~A167 & ~A169;
  assign \new_[9047]_  = ~A265 & A202;
  assign \new_[9048]_  = ~A166 & \new_[9047]_ ;
  assign \new_[9049]_  = \new_[9048]_  & \new_[9043]_ ;
  assign \new_[9052]_  = ~A268 & ~A266;
  assign \new_[9056]_  = A302 & A299;
  assign \new_[9057]_  = ~A298 & \new_[9056]_ ;
  assign \new_[9058]_  = \new_[9057]_  & \new_[9052]_ ;
  assign \new_[9061]_  = ~A167 & ~A169;
  assign \new_[9065]_  = ~A202 & ~A201;
  assign \new_[9066]_  = ~A166 & \new_[9065]_ ;
  assign \new_[9067]_  = \new_[9066]_  & \new_[9061]_ ;
  assign \new_[9070]_  = A268 & ~A203;
  assign \new_[9074]_  = ~A302 & ~A301;
  assign \new_[9075]_  = ~A300 & \new_[9074]_ ;
  assign \new_[9076]_  = \new_[9075]_  & \new_[9070]_ ;
  assign \new_[9079]_  = ~A167 & ~A169;
  assign \new_[9083]_  = ~A202 & ~A201;
  assign \new_[9084]_  = ~A166 & \new_[9083]_ ;
  assign \new_[9085]_  = \new_[9084]_  & \new_[9079]_ ;
  assign \new_[9088]_  = A268 & ~A203;
  assign \new_[9092]_  = ~A301 & ~A299;
  assign \new_[9093]_  = ~A298 & \new_[9092]_ ;
  assign \new_[9094]_  = \new_[9093]_  & \new_[9088]_ ;
  assign \new_[9097]_  = ~A167 & ~A169;
  assign \new_[9101]_  = A201 & A199;
  assign \new_[9102]_  = ~A166 & \new_[9101]_ ;
  assign \new_[9103]_  = \new_[9102]_  & \new_[9097]_ ;
  assign \new_[9106]_  = ~A268 & ~A267;
  assign \new_[9110]_  = A300 & A299;
  assign \new_[9111]_  = ~A269 & \new_[9110]_ ;
  assign \new_[9112]_  = \new_[9111]_  & \new_[9106]_ ;
  assign \new_[9115]_  = ~A167 & ~A169;
  assign \new_[9119]_  = A201 & A199;
  assign \new_[9120]_  = ~A166 & \new_[9119]_ ;
  assign \new_[9121]_  = \new_[9120]_  & \new_[9115]_ ;
  assign \new_[9124]_  = ~A268 & ~A267;
  assign \new_[9128]_  = A300 & A298;
  assign \new_[9129]_  = ~A269 & \new_[9128]_ ;
  assign \new_[9130]_  = \new_[9129]_  & \new_[9124]_ ;
  assign \new_[9133]_  = ~A167 & ~A169;
  assign \new_[9137]_  = A201 & A199;
  assign \new_[9138]_  = ~A166 & \new_[9137]_ ;
  assign \new_[9139]_  = \new_[9138]_  & \new_[9133]_ ;
  assign \new_[9142]_  = A266 & A265;
  assign \new_[9146]_  = A301 & ~A268;
  assign \new_[9147]_  = ~A267 & \new_[9146]_ ;
  assign \new_[9148]_  = \new_[9147]_  & \new_[9142]_ ;
  assign \new_[9151]_  = ~A167 & ~A169;
  assign \new_[9155]_  = A201 & A199;
  assign \new_[9156]_  = ~A166 & \new_[9155]_ ;
  assign \new_[9157]_  = \new_[9156]_  & \new_[9151]_ ;
  assign \new_[9160]_  = ~A266 & ~A265;
  assign \new_[9164]_  = A300 & A299;
  assign \new_[9165]_  = ~A268 & \new_[9164]_ ;
  assign \new_[9166]_  = \new_[9165]_  & \new_[9160]_ ;
  assign \new_[9169]_  = ~A167 & ~A169;
  assign \new_[9173]_  = A201 & A199;
  assign \new_[9174]_  = ~A166 & \new_[9173]_ ;
  assign \new_[9175]_  = \new_[9174]_  & \new_[9169]_ ;
  assign \new_[9178]_  = ~A266 & ~A265;
  assign \new_[9182]_  = A300 & A298;
  assign \new_[9183]_  = ~A268 & \new_[9182]_ ;
  assign \new_[9184]_  = \new_[9183]_  & \new_[9178]_ ;
  assign \new_[9187]_  = ~A167 & ~A169;
  assign \new_[9191]_  = A201 & A200;
  assign \new_[9192]_  = ~A166 & \new_[9191]_ ;
  assign \new_[9193]_  = \new_[9192]_  & \new_[9187]_ ;
  assign \new_[9196]_  = ~A268 & ~A267;
  assign \new_[9200]_  = A300 & A299;
  assign \new_[9201]_  = ~A269 & \new_[9200]_ ;
  assign \new_[9202]_  = \new_[9201]_  & \new_[9196]_ ;
  assign \new_[9205]_  = ~A167 & ~A169;
  assign \new_[9209]_  = A201 & A200;
  assign \new_[9210]_  = ~A166 & \new_[9209]_ ;
  assign \new_[9211]_  = \new_[9210]_  & \new_[9205]_ ;
  assign \new_[9214]_  = ~A268 & ~A267;
  assign \new_[9218]_  = A300 & A298;
  assign \new_[9219]_  = ~A269 & \new_[9218]_ ;
  assign \new_[9220]_  = \new_[9219]_  & \new_[9214]_ ;
  assign \new_[9223]_  = ~A167 & ~A169;
  assign \new_[9227]_  = A201 & A200;
  assign \new_[9228]_  = ~A166 & \new_[9227]_ ;
  assign \new_[9229]_  = \new_[9228]_  & \new_[9223]_ ;
  assign \new_[9232]_  = A266 & A265;
  assign \new_[9236]_  = A301 & ~A268;
  assign \new_[9237]_  = ~A267 & \new_[9236]_ ;
  assign \new_[9238]_  = \new_[9237]_  & \new_[9232]_ ;
  assign \new_[9241]_  = ~A167 & ~A169;
  assign \new_[9245]_  = A201 & A200;
  assign \new_[9246]_  = ~A166 & \new_[9245]_ ;
  assign \new_[9247]_  = \new_[9246]_  & \new_[9241]_ ;
  assign \new_[9250]_  = ~A266 & ~A265;
  assign \new_[9254]_  = A300 & A299;
  assign \new_[9255]_  = ~A268 & \new_[9254]_ ;
  assign \new_[9256]_  = \new_[9255]_  & \new_[9250]_ ;
  assign \new_[9259]_  = ~A167 & ~A169;
  assign \new_[9263]_  = A201 & A200;
  assign \new_[9264]_  = ~A166 & \new_[9263]_ ;
  assign \new_[9265]_  = \new_[9264]_  & \new_[9259]_ ;
  assign \new_[9268]_  = ~A266 & ~A265;
  assign \new_[9272]_  = A300 & A298;
  assign \new_[9273]_  = ~A268 & \new_[9272]_ ;
  assign \new_[9274]_  = \new_[9273]_  & \new_[9268]_ ;
  assign \new_[9277]_  = ~A167 & ~A169;
  assign \new_[9281]_  = A200 & ~A199;
  assign \new_[9282]_  = ~A166 & \new_[9281]_ ;
  assign \new_[9283]_  = \new_[9282]_  & \new_[9277]_ ;
  assign \new_[9286]_  = ~A267 & A203;
  assign \new_[9290]_  = A301 & ~A269;
  assign \new_[9291]_  = ~A268 & \new_[9290]_ ;
  assign \new_[9292]_  = \new_[9291]_  & \new_[9286]_ ;
  assign \new_[9295]_  = ~A167 & ~A169;
  assign \new_[9299]_  = A200 & ~A199;
  assign \new_[9300]_  = ~A166 & \new_[9299]_ ;
  assign \new_[9301]_  = \new_[9300]_  & \new_[9295]_ ;
  assign \new_[9304]_  = ~A265 & A203;
  assign \new_[9308]_  = A301 & ~A268;
  assign \new_[9309]_  = ~A266 & \new_[9308]_ ;
  assign \new_[9310]_  = \new_[9309]_  & \new_[9304]_ ;
  assign \new_[9313]_  = ~A167 & ~A169;
  assign \new_[9317]_  = ~A200 & A199;
  assign \new_[9318]_  = ~A166 & \new_[9317]_ ;
  assign \new_[9319]_  = \new_[9318]_  & \new_[9313]_ ;
  assign \new_[9322]_  = ~A267 & A203;
  assign \new_[9326]_  = A301 & ~A269;
  assign \new_[9327]_  = ~A268 & \new_[9326]_ ;
  assign \new_[9328]_  = \new_[9327]_  & \new_[9322]_ ;
  assign \new_[9331]_  = ~A167 & ~A169;
  assign \new_[9335]_  = ~A200 & A199;
  assign \new_[9336]_  = ~A166 & \new_[9335]_ ;
  assign \new_[9337]_  = \new_[9336]_  & \new_[9331]_ ;
  assign \new_[9340]_  = ~A265 & A203;
  assign \new_[9344]_  = A301 & ~A268;
  assign \new_[9345]_  = ~A266 & \new_[9344]_ ;
  assign \new_[9346]_  = \new_[9345]_  & \new_[9340]_ ;
  assign \new_[9349]_  = ~A167 & ~A169;
  assign \new_[9353]_  = ~A200 & ~A199;
  assign \new_[9354]_  = ~A166 & \new_[9353]_ ;
  assign \new_[9355]_  = \new_[9354]_  & \new_[9349]_ ;
  assign \new_[9358]_  = A268 & ~A202;
  assign \new_[9362]_  = ~A302 & ~A301;
  assign \new_[9363]_  = ~A300 & \new_[9362]_ ;
  assign \new_[9364]_  = \new_[9363]_  & \new_[9358]_ ;
  assign \new_[9367]_  = ~A167 & ~A169;
  assign \new_[9371]_  = ~A200 & ~A199;
  assign \new_[9372]_  = ~A166 & \new_[9371]_ ;
  assign \new_[9373]_  = \new_[9372]_  & \new_[9367]_ ;
  assign \new_[9376]_  = A268 & ~A202;
  assign \new_[9380]_  = ~A301 & ~A299;
  assign \new_[9381]_  = ~A298 & \new_[9380]_ ;
  assign \new_[9382]_  = \new_[9381]_  & \new_[9376]_ ;
  assign \new_[9385]_  = ~A168 & ~A169;
  assign \new_[9389]_  = A202 & A166;
  assign \new_[9390]_  = A167 & \new_[9389]_ ;
  assign \new_[9391]_  = \new_[9390]_  & \new_[9385]_ ;
  assign \new_[9394]_  = ~A268 & ~A267;
  assign \new_[9398]_  = A300 & A299;
  assign \new_[9399]_  = ~A269 & \new_[9398]_ ;
  assign \new_[9400]_  = \new_[9399]_  & \new_[9394]_ ;
  assign \new_[9403]_  = ~A168 & ~A169;
  assign \new_[9407]_  = A202 & A166;
  assign \new_[9408]_  = A167 & \new_[9407]_ ;
  assign \new_[9409]_  = \new_[9408]_  & \new_[9403]_ ;
  assign \new_[9412]_  = ~A268 & ~A267;
  assign \new_[9416]_  = A300 & A298;
  assign \new_[9417]_  = ~A269 & \new_[9416]_ ;
  assign \new_[9418]_  = \new_[9417]_  & \new_[9412]_ ;
  assign \new_[9421]_  = ~A168 & ~A169;
  assign \new_[9425]_  = A202 & A166;
  assign \new_[9426]_  = A167 & \new_[9425]_ ;
  assign \new_[9427]_  = \new_[9426]_  & \new_[9421]_ ;
  assign \new_[9430]_  = A266 & A265;
  assign \new_[9434]_  = A301 & ~A268;
  assign \new_[9435]_  = ~A267 & \new_[9434]_ ;
  assign \new_[9436]_  = \new_[9435]_  & \new_[9430]_ ;
  assign \new_[9439]_  = ~A168 & ~A169;
  assign \new_[9443]_  = A202 & A166;
  assign \new_[9444]_  = A167 & \new_[9443]_ ;
  assign \new_[9445]_  = \new_[9444]_  & \new_[9439]_ ;
  assign \new_[9448]_  = ~A266 & ~A265;
  assign \new_[9452]_  = A300 & A299;
  assign \new_[9453]_  = ~A268 & \new_[9452]_ ;
  assign \new_[9454]_  = \new_[9453]_  & \new_[9448]_ ;
  assign \new_[9457]_  = ~A168 & ~A169;
  assign \new_[9461]_  = A202 & A166;
  assign \new_[9462]_  = A167 & \new_[9461]_ ;
  assign \new_[9463]_  = \new_[9462]_  & \new_[9457]_ ;
  assign \new_[9466]_  = ~A266 & ~A265;
  assign \new_[9470]_  = A300 & A298;
  assign \new_[9471]_  = ~A268 & \new_[9470]_ ;
  assign \new_[9472]_  = \new_[9471]_  & \new_[9466]_ ;
  assign \new_[9475]_  = ~A168 & ~A169;
  assign \new_[9479]_  = A199 & A166;
  assign \new_[9480]_  = A167 & \new_[9479]_ ;
  assign \new_[9481]_  = \new_[9480]_  & \new_[9475]_ ;
  assign \new_[9484]_  = ~A267 & A201;
  assign \new_[9488]_  = A301 & ~A269;
  assign \new_[9489]_  = ~A268 & \new_[9488]_ ;
  assign \new_[9490]_  = \new_[9489]_  & \new_[9484]_ ;
  assign \new_[9493]_  = ~A168 & ~A169;
  assign \new_[9497]_  = A199 & A166;
  assign \new_[9498]_  = A167 & \new_[9497]_ ;
  assign \new_[9499]_  = \new_[9498]_  & \new_[9493]_ ;
  assign \new_[9502]_  = ~A265 & A201;
  assign \new_[9506]_  = A301 & ~A268;
  assign \new_[9507]_  = ~A266 & \new_[9506]_ ;
  assign \new_[9508]_  = \new_[9507]_  & \new_[9502]_ ;
  assign \new_[9511]_  = ~A168 & ~A169;
  assign \new_[9515]_  = A200 & A166;
  assign \new_[9516]_  = A167 & \new_[9515]_ ;
  assign \new_[9517]_  = \new_[9516]_  & \new_[9511]_ ;
  assign \new_[9520]_  = ~A267 & A201;
  assign \new_[9524]_  = A301 & ~A269;
  assign \new_[9525]_  = ~A268 & \new_[9524]_ ;
  assign \new_[9526]_  = \new_[9525]_  & \new_[9520]_ ;
  assign \new_[9529]_  = ~A168 & ~A169;
  assign \new_[9533]_  = A200 & A166;
  assign \new_[9534]_  = A167 & \new_[9533]_ ;
  assign \new_[9535]_  = \new_[9534]_  & \new_[9529]_ ;
  assign \new_[9538]_  = ~A265 & A201;
  assign \new_[9542]_  = A301 & ~A268;
  assign \new_[9543]_  = ~A266 & \new_[9542]_ ;
  assign \new_[9544]_  = \new_[9543]_  & \new_[9538]_ ;
  assign \new_[9547]_  = ~A169 & ~A170;
  assign \new_[9551]_  = ~A267 & A202;
  assign \new_[9552]_  = ~A168 & \new_[9551]_ ;
  assign \new_[9553]_  = \new_[9552]_  & \new_[9547]_ ;
  assign \new_[9556]_  = ~A269 & ~A268;
  assign \new_[9560]_  = A302 & ~A299;
  assign \new_[9561]_  = A298 & \new_[9560]_ ;
  assign \new_[9562]_  = \new_[9561]_  & \new_[9556]_ ;
  assign \new_[9565]_  = ~A169 & ~A170;
  assign \new_[9569]_  = ~A267 & A202;
  assign \new_[9570]_  = ~A168 & \new_[9569]_ ;
  assign \new_[9571]_  = \new_[9570]_  & \new_[9565]_ ;
  assign \new_[9574]_  = ~A269 & ~A268;
  assign \new_[9578]_  = A302 & A299;
  assign \new_[9579]_  = ~A298 & \new_[9578]_ ;
  assign \new_[9580]_  = \new_[9579]_  & \new_[9574]_ ;
  assign \new_[9583]_  = ~A169 & ~A170;
  assign \new_[9587]_  = A265 & A202;
  assign \new_[9588]_  = ~A168 & \new_[9587]_ ;
  assign \new_[9589]_  = \new_[9588]_  & \new_[9583]_ ;
  assign \new_[9592]_  = ~A267 & A266;
  assign \new_[9596]_  = A300 & A299;
  assign \new_[9597]_  = ~A268 & \new_[9596]_ ;
  assign \new_[9598]_  = \new_[9597]_  & \new_[9592]_ ;
  assign \new_[9601]_  = ~A169 & ~A170;
  assign \new_[9605]_  = A265 & A202;
  assign \new_[9606]_  = ~A168 & \new_[9605]_ ;
  assign \new_[9607]_  = \new_[9606]_  & \new_[9601]_ ;
  assign \new_[9610]_  = ~A267 & A266;
  assign \new_[9614]_  = A300 & A298;
  assign \new_[9615]_  = ~A268 & \new_[9614]_ ;
  assign \new_[9616]_  = \new_[9615]_  & \new_[9610]_ ;
  assign \new_[9619]_  = ~A169 & ~A170;
  assign \new_[9623]_  = ~A265 & A202;
  assign \new_[9624]_  = ~A168 & \new_[9623]_ ;
  assign \new_[9625]_  = \new_[9624]_  & \new_[9619]_ ;
  assign \new_[9628]_  = ~A268 & ~A266;
  assign \new_[9632]_  = A302 & ~A299;
  assign \new_[9633]_  = A298 & \new_[9632]_ ;
  assign \new_[9634]_  = \new_[9633]_  & \new_[9628]_ ;
  assign \new_[9637]_  = ~A169 & ~A170;
  assign \new_[9641]_  = ~A265 & A202;
  assign \new_[9642]_  = ~A168 & \new_[9641]_ ;
  assign \new_[9643]_  = \new_[9642]_  & \new_[9637]_ ;
  assign \new_[9646]_  = ~A268 & ~A266;
  assign \new_[9650]_  = A302 & A299;
  assign \new_[9651]_  = ~A298 & \new_[9650]_ ;
  assign \new_[9652]_  = \new_[9651]_  & \new_[9646]_ ;
  assign \new_[9655]_  = ~A169 & ~A170;
  assign \new_[9659]_  = ~A202 & ~A201;
  assign \new_[9660]_  = ~A168 & \new_[9659]_ ;
  assign \new_[9661]_  = \new_[9660]_  & \new_[9655]_ ;
  assign \new_[9664]_  = A268 & ~A203;
  assign \new_[9668]_  = ~A302 & ~A301;
  assign \new_[9669]_  = ~A300 & \new_[9668]_ ;
  assign \new_[9670]_  = \new_[9669]_  & \new_[9664]_ ;
  assign \new_[9673]_  = ~A169 & ~A170;
  assign \new_[9677]_  = ~A202 & ~A201;
  assign \new_[9678]_  = ~A168 & \new_[9677]_ ;
  assign \new_[9679]_  = \new_[9678]_  & \new_[9673]_ ;
  assign \new_[9682]_  = A268 & ~A203;
  assign \new_[9686]_  = ~A301 & ~A299;
  assign \new_[9687]_  = ~A298 & \new_[9686]_ ;
  assign \new_[9688]_  = \new_[9687]_  & \new_[9682]_ ;
  assign \new_[9691]_  = ~A169 & ~A170;
  assign \new_[9695]_  = A201 & A199;
  assign \new_[9696]_  = ~A168 & \new_[9695]_ ;
  assign \new_[9697]_  = \new_[9696]_  & \new_[9691]_ ;
  assign \new_[9700]_  = ~A268 & ~A267;
  assign \new_[9704]_  = A300 & A299;
  assign \new_[9705]_  = ~A269 & \new_[9704]_ ;
  assign \new_[9706]_  = \new_[9705]_  & \new_[9700]_ ;
  assign \new_[9709]_  = ~A169 & ~A170;
  assign \new_[9713]_  = A201 & A199;
  assign \new_[9714]_  = ~A168 & \new_[9713]_ ;
  assign \new_[9715]_  = \new_[9714]_  & \new_[9709]_ ;
  assign \new_[9718]_  = ~A268 & ~A267;
  assign \new_[9722]_  = A300 & A298;
  assign \new_[9723]_  = ~A269 & \new_[9722]_ ;
  assign \new_[9724]_  = \new_[9723]_  & \new_[9718]_ ;
  assign \new_[9727]_  = ~A169 & ~A170;
  assign \new_[9731]_  = A201 & A199;
  assign \new_[9732]_  = ~A168 & \new_[9731]_ ;
  assign \new_[9733]_  = \new_[9732]_  & \new_[9727]_ ;
  assign \new_[9736]_  = A266 & A265;
  assign \new_[9740]_  = A301 & ~A268;
  assign \new_[9741]_  = ~A267 & \new_[9740]_ ;
  assign \new_[9742]_  = \new_[9741]_  & \new_[9736]_ ;
  assign \new_[9745]_  = ~A169 & ~A170;
  assign \new_[9749]_  = A201 & A199;
  assign \new_[9750]_  = ~A168 & \new_[9749]_ ;
  assign \new_[9751]_  = \new_[9750]_  & \new_[9745]_ ;
  assign \new_[9754]_  = ~A266 & ~A265;
  assign \new_[9758]_  = A300 & A299;
  assign \new_[9759]_  = ~A268 & \new_[9758]_ ;
  assign \new_[9760]_  = \new_[9759]_  & \new_[9754]_ ;
  assign \new_[9763]_  = ~A169 & ~A170;
  assign \new_[9767]_  = A201 & A199;
  assign \new_[9768]_  = ~A168 & \new_[9767]_ ;
  assign \new_[9769]_  = \new_[9768]_  & \new_[9763]_ ;
  assign \new_[9772]_  = ~A266 & ~A265;
  assign \new_[9776]_  = A300 & A298;
  assign \new_[9777]_  = ~A268 & \new_[9776]_ ;
  assign \new_[9778]_  = \new_[9777]_  & \new_[9772]_ ;
  assign \new_[9781]_  = ~A169 & ~A170;
  assign \new_[9785]_  = A201 & A200;
  assign \new_[9786]_  = ~A168 & \new_[9785]_ ;
  assign \new_[9787]_  = \new_[9786]_  & \new_[9781]_ ;
  assign \new_[9790]_  = ~A268 & ~A267;
  assign \new_[9794]_  = A300 & A299;
  assign \new_[9795]_  = ~A269 & \new_[9794]_ ;
  assign \new_[9796]_  = \new_[9795]_  & \new_[9790]_ ;
  assign \new_[9799]_  = ~A169 & ~A170;
  assign \new_[9803]_  = A201 & A200;
  assign \new_[9804]_  = ~A168 & \new_[9803]_ ;
  assign \new_[9805]_  = \new_[9804]_  & \new_[9799]_ ;
  assign \new_[9808]_  = ~A268 & ~A267;
  assign \new_[9812]_  = A300 & A298;
  assign \new_[9813]_  = ~A269 & \new_[9812]_ ;
  assign \new_[9814]_  = \new_[9813]_  & \new_[9808]_ ;
  assign \new_[9817]_  = ~A169 & ~A170;
  assign \new_[9821]_  = A201 & A200;
  assign \new_[9822]_  = ~A168 & \new_[9821]_ ;
  assign \new_[9823]_  = \new_[9822]_  & \new_[9817]_ ;
  assign \new_[9826]_  = A266 & A265;
  assign \new_[9830]_  = A301 & ~A268;
  assign \new_[9831]_  = ~A267 & \new_[9830]_ ;
  assign \new_[9832]_  = \new_[9831]_  & \new_[9826]_ ;
  assign \new_[9835]_  = ~A169 & ~A170;
  assign \new_[9839]_  = A201 & A200;
  assign \new_[9840]_  = ~A168 & \new_[9839]_ ;
  assign \new_[9841]_  = \new_[9840]_  & \new_[9835]_ ;
  assign \new_[9844]_  = ~A266 & ~A265;
  assign \new_[9848]_  = A300 & A299;
  assign \new_[9849]_  = ~A268 & \new_[9848]_ ;
  assign \new_[9850]_  = \new_[9849]_  & \new_[9844]_ ;
  assign \new_[9853]_  = ~A169 & ~A170;
  assign \new_[9857]_  = A201 & A200;
  assign \new_[9858]_  = ~A168 & \new_[9857]_ ;
  assign \new_[9859]_  = \new_[9858]_  & \new_[9853]_ ;
  assign \new_[9862]_  = ~A266 & ~A265;
  assign \new_[9866]_  = A300 & A298;
  assign \new_[9867]_  = ~A268 & \new_[9866]_ ;
  assign \new_[9868]_  = \new_[9867]_  & \new_[9862]_ ;
  assign \new_[9871]_  = ~A169 & ~A170;
  assign \new_[9875]_  = A200 & ~A199;
  assign \new_[9876]_  = ~A168 & \new_[9875]_ ;
  assign \new_[9877]_  = \new_[9876]_  & \new_[9871]_ ;
  assign \new_[9880]_  = ~A267 & A203;
  assign \new_[9884]_  = A301 & ~A269;
  assign \new_[9885]_  = ~A268 & \new_[9884]_ ;
  assign \new_[9886]_  = \new_[9885]_  & \new_[9880]_ ;
  assign \new_[9889]_  = ~A169 & ~A170;
  assign \new_[9893]_  = A200 & ~A199;
  assign \new_[9894]_  = ~A168 & \new_[9893]_ ;
  assign \new_[9895]_  = \new_[9894]_  & \new_[9889]_ ;
  assign \new_[9898]_  = ~A265 & A203;
  assign \new_[9902]_  = A301 & ~A268;
  assign \new_[9903]_  = ~A266 & \new_[9902]_ ;
  assign \new_[9904]_  = \new_[9903]_  & \new_[9898]_ ;
  assign \new_[9907]_  = ~A169 & ~A170;
  assign \new_[9911]_  = ~A200 & A199;
  assign \new_[9912]_  = ~A168 & \new_[9911]_ ;
  assign \new_[9913]_  = \new_[9912]_  & \new_[9907]_ ;
  assign \new_[9916]_  = ~A267 & A203;
  assign \new_[9920]_  = A301 & ~A269;
  assign \new_[9921]_  = ~A268 & \new_[9920]_ ;
  assign \new_[9922]_  = \new_[9921]_  & \new_[9916]_ ;
  assign \new_[9925]_  = ~A169 & ~A170;
  assign \new_[9929]_  = ~A200 & A199;
  assign \new_[9930]_  = ~A168 & \new_[9929]_ ;
  assign \new_[9931]_  = \new_[9930]_  & \new_[9925]_ ;
  assign \new_[9934]_  = ~A265 & A203;
  assign \new_[9938]_  = A301 & ~A268;
  assign \new_[9939]_  = ~A266 & \new_[9938]_ ;
  assign \new_[9940]_  = \new_[9939]_  & \new_[9934]_ ;
  assign \new_[9943]_  = ~A169 & ~A170;
  assign \new_[9947]_  = ~A200 & ~A199;
  assign \new_[9948]_  = ~A168 & \new_[9947]_ ;
  assign \new_[9949]_  = \new_[9948]_  & \new_[9943]_ ;
  assign \new_[9952]_  = A268 & ~A202;
  assign \new_[9956]_  = ~A302 & ~A301;
  assign \new_[9957]_  = ~A300 & \new_[9956]_ ;
  assign \new_[9958]_  = \new_[9957]_  & \new_[9952]_ ;
  assign \new_[9961]_  = ~A169 & ~A170;
  assign \new_[9965]_  = ~A200 & ~A199;
  assign \new_[9966]_  = ~A168 & \new_[9965]_ ;
  assign \new_[9967]_  = \new_[9966]_  & \new_[9961]_ ;
  assign \new_[9970]_  = A268 & ~A202;
  assign \new_[9974]_  = ~A301 & ~A299;
  assign \new_[9975]_  = ~A298 & \new_[9974]_ ;
  assign \new_[9976]_  = \new_[9975]_  & \new_[9970]_ ;
  assign \new_[9979]_  = A166 & A168;
  assign \new_[9983]_  = ~A203 & ~A202;
  assign \new_[9984]_  = ~A201 & \new_[9983]_ ;
  assign \new_[9985]_  = \new_[9984]_  & \new_[9979]_ ;
  assign \new_[9989]_  = ~A269 & ~A268;
  assign \new_[9990]_  = ~A267 & \new_[9989]_ ;
  assign \new_[9994]_  = A302 & ~A299;
  assign \new_[9995]_  = A298 & \new_[9994]_ ;
  assign \new_[9996]_  = \new_[9995]_  & \new_[9990]_ ;
  assign \new_[9999]_  = A166 & A168;
  assign \new_[10003]_  = ~A203 & ~A202;
  assign \new_[10004]_  = ~A201 & \new_[10003]_ ;
  assign \new_[10005]_  = \new_[10004]_  & \new_[9999]_ ;
  assign \new_[10009]_  = ~A269 & ~A268;
  assign \new_[10010]_  = ~A267 & \new_[10009]_ ;
  assign \new_[10014]_  = A302 & A299;
  assign \new_[10015]_  = ~A298 & \new_[10014]_ ;
  assign \new_[10016]_  = \new_[10015]_  & \new_[10010]_ ;
  assign \new_[10019]_  = A166 & A168;
  assign \new_[10023]_  = ~A203 & ~A202;
  assign \new_[10024]_  = ~A201 & \new_[10023]_ ;
  assign \new_[10025]_  = \new_[10024]_  & \new_[10019]_ ;
  assign \new_[10029]_  = ~A267 & A266;
  assign \new_[10030]_  = A265 & \new_[10029]_ ;
  assign \new_[10034]_  = A300 & A299;
  assign \new_[10035]_  = ~A268 & \new_[10034]_ ;
  assign \new_[10036]_  = \new_[10035]_  & \new_[10030]_ ;
  assign \new_[10039]_  = A166 & A168;
  assign \new_[10043]_  = ~A203 & ~A202;
  assign \new_[10044]_  = ~A201 & \new_[10043]_ ;
  assign \new_[10045]_  = \new_[10044]_  & \new_[10039]_ ;
  assign \new_[10049]_  = ~A267 & A266;
  assign \new_[10050]_  = A265 & \new_[10049]_ ;
  assign \new_[10054]_  = A300 & A298;
  assign \new_[10055]_  = ~A268 & \new_[10054]_ ;
  assign \new_[10056]_  = \new_[10055]_  & \new_[10050]_ ;
  assign \new_[10059]_  = A166 & A168;
  assign \new_[10063]_  = ~A203 & ~A202;
  assign \new_[10064]_  = ~A201 & \new_[10063]_ ;
  assign \new_[10065]_  = \new_[10064]_  & \new_[10059]_ ;
  assign \new_[10069]_  = ~A268 & ~A266;
  assign \new_[10070]_  = ~A265 & \new_[10069]_ ;
  assign \new_[10074]_  = A302 & ~A299;
  assign \new_[10075]_  = A298 & \new_[10074]_ ;
  assign \new_[10076]_  = \new_[10075]_  & \new_[10070]_ ;
  assign \new_[10079]_  = A166 & A168;
  assign \new_[10083]_  = ~A203 & ~A202;
  assign \new_[10084]_  = ~A201 & \new_[10083]_ ;
  assign \new_[10085]_  = \new_[10084]_  & \new_[10079]_ ;
  assign \new_[10089]_  = ~A268 & ~A266;
  assign \new_[10090]_  = ~A265 & \new_[10089]_ ;
  assign \new_[10094]_  = A302 & A299;
  assign \new_[10095]_  = ~A298 & \new_[10094]_ ;
  assign \new_[10096]_  = \new_[10095]_  & \new_[10090]_ ;
  assign \new_[10099]_  = A166 & A168;
  assign \new_[10103]_  = ~A265 & A201;
  assign \new_[10104]_  = A199 & \new_[10103]_ ;
  assign \new_[10105]_  = \new_[10104]_  & \new_[10099]_ ;
  assign \new_[10109]_  = A298 & A269;
  assign \new_[10110]_  = A266 & \new_[10109]_ ;
  assign \new_[10114]_  = ~A301 & ~A300;
  assign \new_[10115]_  = A299 & \new_[10114]_ ;
  assign \new_[10116]_  = \new_[10115]_  & \new_[10110]_ ;
  assign \new_[10119]_  = A166 & A168;
  assign \new_[10123]_  = A265 & A201;
  assign \new_[10124]_  = A199 & \new_[10123]_ ;
  assign \new_[10125]_  = \new_[10124]_  & \new_[10119]_ ;
  assign \new_[10129]_  = A298 & A269;
  assign \new_[10130]_  = ~A266 & \new_[10129]_ ;
  assign \new_[10134]_  = ~A301 & ~A300;
  assign \new_[10135]_  = A299 & \new_[10134]_ ;
  assign \new_[10136]_  = \new_[10135]_  & \new_[10130]_ ;
  assign \new_[10139]_  = A166 & A168;
  assign \new_[10143]_  = ~A265 & A201;
  assign \new_[10144]_  = A200 & \new_[10143]_ ;
  assign \new_[10145]_  = \new_[10144]_  & \new_[10139]_ ;
  assign \new_[10149]_  = A298 & A269;
  assign \new_[10150]_  = A266 & \new_[10149]_ ;
  assign \new_[10154]_  = ~A301 & ~A300;
  assign \new_[10155]_  = A299 & \new_[10154]_ ;
  assign \new_[10156]_  = \new_[10155]_  & \new_[10150]_ ;
  assign \new_[10159]_  = A166 & A168;
  assign \new_[10163]_  = A265 & A201;
  assign \new_[10164]_  = A200 & \new_[10163]_ ;
  assign \new_[10165]_  = \new_[10164]_  & \new_[10159]_ ;
  assign \new_[10169]_  = A298 & A269;
  assign \new_[10170]_  = ~A266 & \new_[10169]_ ;
  assign \new_[10174]_  = ~A301 & ~A300;
  assign \new_[10175]_  = A299 & \new_[10174]_ ;
  assign \new_[10176]_  = \new_[10175]_  & \new_[10170]_ ;
  assign \new_[10179]_  = A166 & A168;
  assign \new_[10183]_  = ~A201 & A200;
  assign \new_[10184]_  = A199 & \new_[10183]_ ;
  assign \new_[10185]_  = \new_[10184]_  & \new_[10179]_ ;
  assign \new_[10189]_  = ~A268 & ~A267;
  assign \new_[10190]_  = ~A202 & \new_[10189]_ ;
  assign \new_[10194]_  = A300 & A299;
  assign \new_[10195]_  = ~A269 & \new_[10194]_ ;
  assign \new_[10196]_  = \new_[10195]_  & \new_[10190]_ ;
  assign \new_[10199]_  = A166 & A168;
  assign \new_[10203]_  = ~A201 & A200;
  assign \new_[10204]_  = A199 & \new_[10203]_ ;
  assign \new_[10205]_  = \new_[10204]_  & \new_[10199]_ ;
  assign \new_[10209]_  = ~A268 & ~A267;
  assign \new_[10210]_  = ~A202 & \new_[10209]_ ;
  assign \new_[10214]_  = A300 & A298;
  assign \new_[10215]_  = ~A269 & \new_[10214]_ ;
  assign \new_[10216]_  = \new_[10215]_  & \new_[10210]_ ;
  assign \new_[10219]_  = A166 & A168;
  assign \new_[10223]_  = ~A201 & A200;
  assign \new_[10224]_  = A199 & \new_[10223]_ ;
  assign \new_[10225]_  = \new_[10224]_  & \new_[10219]_ ;
  assign \new_[10229]_  = A266 & A265;
  assign \new_[10230]_  = ~A202 & \new_[10229]_ ;
  assign \new_[10234]_  = A301 & ~A268;
  assign \new_[10235]_  = ~A267 & \new_[10234]_ ;
  assign \new_[10236]_  = \new_[10235]_  & \new_[10230]_ ;
  assign \new_[10239]_  = A166 & A168;
  assign \new_[10243]_  = ~A201 & A200;
  assign \new_[10244]_  = A199 & \new_[10243]_ ;
  assign \new_[10245]_  = \new_[10244]_  & \new_[10239]_ ;
  assign \new_[10249]_  = ~A266 & ~A265;
  assign \new_[10250]_  = ~A202 & \new_[10249]_ ;
  assign \new_[10254]_  = A300 & A299;
  assign \new_[10255]_  = ~A268 & \new_[10254]_ ;
  assign \new_[10256]_  = \new_[10255]_  & \new_[10250]_ ;
  assign \new_[10259]_  = A166 & A168;
  assign \new_[10263]_  = ~A201 & A200;
  assign \new_[10264]_  = A199 & \new_[10263]_ ;
  assign \new_[10265]_  = \new_[10264]_  & \new_[10259]_ ;
  assign \new_[10269]_  = ~A266 & ~A265;
  assign \new_[10270]_  = ~A202 & \new_[10269]_ ;
  assign \new_[10274]_  = A300 & A298;
  assign \new_[10275]_  = ~A268 & \new_[10274]_ ;
  assign \new_[10276]_  = \new_[10275]_  & \new_[10270]_ ;
  assign \new_[10279]_  = A166 & A168;
  assign \new_[10283]_  = A203 & A200;
  assign \new_[10284]_  = ~A199 & \new_[10283]_ ;
  assign \new_[10285]_  = \new_[10284]_  & \new_[10279]_ ;
  assign \new_[10289]_  = A298 & A267;
  assign \new_[10290]_  = A265 & \new_[10289]_ ;
  assign \new_[10294]_  = ~A301 & ~A300;
  assign \new_[10295]_  = A299 & \new_[10294]_ ;
  assign \new_[10296]_  = \new_[10295]_  & \new_[10290]_ ;
  assign \new_[10299]_  = A166 & A168;
  assign \new_[10303]_  = A203 & A200;
  assign \new_[10304]_  = ~A199 & \new_[10303]_ ;
  assign \new_[10305]_  = \new_[10304]_  & \new_[10299]_ ;
  assign \new_[10309]_  = A298 & A267;
  assign \new_[10310]_  = A266 & \new_[10309]_ ;
  assign \new_[10314]_  = ~A301 & ~A300;
  assign \new_[10315]_  = A299 & \new_[10314]_ ;
  assign \new_[10316]_  = \new_[10315]_  & \new_[10310]_ ;
  assign \new_[10319]_  = A166 & A168;
  assign \new_[10323]_  = A203 & A200;
  assign \new_[10324]_  = ~A199 & \new_[10323]_ ;
  assign \new_[10325]_  = \new_[10324]_  & \new_[10319]_ ;
  assign \new_[10329]_  = A269 & A266;
  assign \new_[10330]_  = ~A265 & \new_[10329]_ ;
  assign \new_[10334]_  = ~A302 & ~A301;
  assign \new_[10335]_  = ~A300 & \new_[10334]_ ;
  assign \new_[10336]_  = \new_[10335]_  & \new_[10330]_ ;
  assign \new_[10339]_  = A166 & A168;
  assign \new_[10343]_  = A203 & A200;
  assign \new_[10344]_  = ~A199 & \new_[10343]_ ;
  assign \new_[10345]_  = \new_[10344]_  & \new_[10339]_ ;
  assign \new_[10349]_  = A269 & A266;
  assign \new_[10350]_  = ~A265 & \new_[10349]_ ;
  assign \new_[10354]_  = ~A301 & ~A299;
  assign \new_[10355]_  = ~A298 & \new_[10354]_ ;
  assign \new_[10356]_  = \new_[10355]_  & \new_[10350]_ ;
  assign \new_[10359]_  = A166 & A168;
  assign \new_[10363]_  = A203 & A200;
  assign \new_[10364]_  = ~A199 & \new_[10363]_ ;
  assign \new_[10365]_  = \new_[10364]_  & \new_[10359]_ ;
  assign \new_[10369]_  = A269 & ~A266;
  assign \new_[10370]_  = A265 & \new_[10369]_ ;
  assign \new_[10374]_  = ~A302 & ~A301;
  assign \new_[10375]_  = ~A300 & \new_[10374]_ ;
  assign \new_[10376]_  = \new_[10375]_  & \new_[10370]_ ;
  assign \new_[10379]_  = A166 & A168;
  assign \new_[10383]_  = A203 & A200;
  assign \new_[10384]_  = ~A199 & \new_[10383]_ ;
  assign \new_[10385]_  = \new_[10384]_  & \new_[10379]_ ;
  assign \new_[10389]_  = A269 & ~A266;
  assign \new_[10390]_  = A265 & \new_[10389]_ ;
  assign \new_[10394]_  = ~A301 & ~A299;
  assign \new_[10395]_  = ~A298 & \new_[10394]_ ;
  assign \new_[10396]_  = \new_[10395]_  & \new_[10390]_ ;
  assign \new_[10399]_  = A166 & A168;
  assign \new_[10403]_  = A203 & ~A200;
  assign \new_[10404]_  = A199 & \new_[10403]_ ;
  assign \new_[10405]_  = \new_[10404]_  & \new_[10399]_ ;
  assign \new_[10409]_  = A298 & A267;
  assign \new_[10410]_  = A265 & \new_[10409]_ ;
  assign \new_[10414]_  = ~A301 & ~A300;
  assign \new_[10415]_  = A299 & \new_[10414]_ ;
  assign \new_[10416]_  = \new_[10415]_  & \new_[10410]_ ;
  assign \new_[10419]_  = A166 & A168;
  assign \new_[10423]_  = A203 & ~A200;
  assign \new_[10424]_  = A199 & \new_[10423]_ ;
  assign \new_[10425]_  = \new_[10424]_  & \new_[10419]_ ;
  assign \new_[10429]_  = A298 & A267;
  assign \new_[10430]_  = A266 & \new_[10429]_ ;
  assign \new_[10434]_  = ~A301 & ~A300;
  assign \new_[10435]_  = A299 & \new_[10434]_ ;
  assign \new_[10436]_  = \new_[10435]_  & \new_[10430]_ ;
  assign \new_[10439]_  = A166 & A168;
  assign \new_[10443]_  = A203 & ~A200;
  assign \new_[10444]_  = A199 & \new_[10443]_ ;
  assign \new_[10445]_  = \new_[10444]_  & \new_[10439]_ ;
  assign \new_[10449]_  = A269 & A266;
  assign \new_[10450]_  = ~A265 & \new_[10449]_ ;
  assign \new_[10454]_  = ~A302 & ~A301;
  assign \new_[10455]_  = ~A300 & \new_[10454]_ ;
  assign \new_[10456]_  = \new_[10455]_  & \new_[10450]_ ;
  assign \new_[10459]_  = A166 & A168;
  assign \new_[10463]_  = A203 & ~A200;
  assign \new_[10464]_  = A199 & \new_[10463]_ ;
  assign \new_[10465]_  = \new_[10464]_  & \new_[10459]_ ;
  assign \new_[10469]_  = A269 & A266;
  assign \new_[10470]_  = ~A265 & \new_[10469]_ ;
  assign \new_[10474]_  = ~A301 & ~A299;
  assign \new_[10475]_  = ~A298 & \new_[10474]_ ;
  assign \new_[10476]_  = \new_[10475]_  & \new_[10470]_ ;
  assign \new_[10479]_  = A166 & A168;
  assign \new_[10483]_  = A203 & ~A200;
  assign \new_[10484]_  = A199 & \new_[10483]_ ;
  assign \new_[10485]_  = \new_[10484]_  & \new_[10479]_ ;
  assign \new_[10489]_  = A269 & ~A266;
  assign \new_[10490]_  = A265 & \new_[10489]_ ;
  assign \new_[10494]_  = ~A302 & ~A301;
  assign \new_[10495]_  = ~A300 & \new_[10494]_ ;
  assign \new_[10496]_  = \new_[10495]_  & \new_[10490]_ ;
  assign \new_[10499]_  = A166 & A168;
  assign \new_[10503]_  = A203 & ~A200;
  assign \new_[10504]_  = A199 & \new_[10503]_ ;
  assign \new_[10505]_  = \new_[10504]_  & \new_[10499]_ ;
  assign \new_[10509]_  = A269 & ~A266;
  assign \new_[10510]_  = A265 & \new_[10509]_ ;
  assign \new_[10514]_  = ~A301 & ~A299;
  assign \new_[10515]_  = ~A298 & \new_[10514]_ ;
  assign \new_[10516]_  = \new_[10515]_  & \new_[10510]_ ;
  assign \new_[10519]_  = A166 & A168;
  assign \new_[10523]_  = ~A202 & ~A200;
  assign \new_[10524]_  = ~A199 & \new_[10523]_ ;
  assign \new_[10525]_  = \new_[10524]_  & \new_[10519]_ ;
  assign \new_[10529]_  = ~A269 & ~A268;
  assign \new_[10530]_  = ~A267 & \new_[10529]_ ;
  assign \new_[10534]_  = A302 & ~A299;
  assign \new_[10535]_  = A298 & \new_[10534]_ ;
  assign \new_[10536]_  = \new_[10535]_  & \new_[10530]_ ;
  assign \new_[10539]_  = A166 & A168;
  assign \new_[10543]_  = ~A202 & ~A200;
  assign \new_[10544]_  = ~A199 & \new_[10543]_ ;
  assign \new_[10545]_  = \new_[10544]_  & \new_[10539]_ ;
  assign \new_[10549]_  = ~A269 & ~A268;
  assign \new_[10550]_  = ~A267 & \new_[10549]_ ;
  assign \new_[10554]_  = A302 & A299;
  assign \new_[10555]_  = ~A298 & \new_[10554]_ ;
  assign \new_[10556]_  = \new_[10555]_  & \new_[10550]_ ;
  assign \new_[10559]_  = A166 & A168;
  assign \new_[10563]_  = ~A202 & ~A200;
  assign \new_[10564]_  = ~A199 & \new_[10563]_ ;
  assign \new_[10565]_  = \new_[10564]_  & \new_[10559]_ ;
  assign \new_[10569]_  = ~A267 & A266;
  assign \new_[10570]_  = A265 & \new_[10569]_ ;
  assign \new_[10574]_  = A300 & A299;
  assign \new_[10575]_  = ~A268 & \new_[10574]_ ;
  assign \new_[10576]_  = \new_[10575]_  & \new_[10570]_ ;
  assign \new_[10579]_  = A166 & A168;
  assign \new_[10583]_  = ~A202 & ~A200;
  assign \new_[10584]_  = ~A199 & \new_[10583]_ ;
  assign \new_[10585]_  = \new_[10584]_  & \new_[10579]_ ;
  assign \new_[10589]_  = ~A267 & A266;
  assign \new_[10590]_  = A265 & \new_[10589]_ ;
  assign \new_[10594]_  = A300 & A298;
  assign \new_[10595]_  = ~A268 & \new_[10594]_ ;
  assign \new_[10596]_  = \new_[10595]_  & \new_[10590]_ ;
  assign \new_[10599]_  = A166 & A168;
  assign \new_[10603]_  = ~A202 & ~A200;
  assign \new_[10604]_  = ~A199 & \new_[10603]_ ;
  assign \new_[10605]_  = \new_[10604]_  & \new_[10599]_ ;
  assign \new_[10609]_  = ~A268 & ~A266;
  assign \new_[10610]_  = ~A265 & \new_[10609]_ ;
  assign \new_[10614]_  = A302 & ~A299;
  assign \new_[10615]_  = A298 & \new_[10614]_ ;
  assign \new_[10616]_  = \new_[10615]_  & \new_[10610]_ ;
  assign \new_[10619]_  = A166 & A168;
  assign \new_[10623]_  = ~A202 & ~A200;
  assign \new_[10624]_  = ~A199 & \new_[10623]_ ;
  assign \new_[10625]_  = \new_[10624]_  & \new_[10619]_ ;
  assign \new_[10629]_  = ~A268 & ~A266;
  assign \new_[10630]_  = ~A265 & \new_[10629]_ ;
  assign \new_[10634]_  = A302 & A299;
  assign \new_[10635]_  = ~A298 & \new_[10634]_ ;
  assign \new_[10636]_  = \new_[10635]_  & \new_[10630]_ ;
  assign \new_[10639]_  = A167 & A168;
  assign \new_[10643]_  = ~A203 & ~A202;
  assign \new_[10644]_  = ~A201 & \new_[10643]_ ;
  assign \new_[10645]_  = \new_[10644]_  & \new_[10639]_ ;
  assign \new_[10649]_  = ~A269 & ~A268;
  assign \new_[10650]_  = ~A267 & \new_[10649]_ ;
  assign \new_[10654]_  = A302 & ~A299;
  assign \new_[10655]_  = A298 & \new_[10654]_ ;
  assign \new_[10656]_  = \new_[10655]_  & \new_[10650]_ ;
  assign \new_[10659]_  = A167 & A168;
  assign \new_[10663]_  = ~A203 & ~A202;
  assign \new_[10664]_  = ~A201 & \new_[10663]_ ;
  assign \new_[10665]_  = \new_[10664]_  & \new_[10659]_ ;
  assign \new_[10669]_  = ~A269 & ~A268;
  assign \new_[10670]_  = ~A267 & \new_[10669]_ ;
  assign \new_[10674]_  = A302 & A299;
  assign \new_[10675]_  = ~A298 & \new_[10674]_ ;
  assign \new_[10676]_  = \new_[10675]_  & \new_[10670]_ ;
  assign \new_[10679]_  = A167 & A168;
  assign \new_[10683]_  = ~A203 & ~A202;
  assign \new_[10684]_  = ~A201 & \new_[10683]_ ;
  assign \new_[10685]_  = \new_[10684]_  & \new_[10679]_ ;
  assign \new_[10689]_  = ~A267 & A266;
  assign \new_[10690]_  = A265 & \new_[10689]_ ;
  assign \new_[10694]_  = A300 & A299;
  assign \new_[10695]_  = ~A268 & \new_[10694]_ ;
  assign \new_[10696]_  = \new_[10695]_  & \new_[10690]_ ;
  assign \new_[10699]_  = A167 & A168;
  assign \new_[10703]_  = ~A203 & ~A202;
  assign \new_[10704]_  = ~A201 & \new_[10703]_ ;
  assign \new_[10705]_  = \new_[10704]_  & \new_[10699]_ ;
  assign \new_[10709]_  = ~A267 & A266;
  assign \new_[10710]_  = A265 & \new_[10709]_ ;
  assign \new_[10714]_  = A300 & A298;
  assign \new_[10715]_  = ~A268 & \new_[10714]_ ;
  assign \new_[10716]_  = \new_[10715]_  & \new_[10710]_ ;
  assign \new_[10719]_  = A167 & A168;
  assign \new_[10723]_  = ~A203 & ~A202;
  assign \new_[10724]_  = ~A201 & \new_[10723]_ ;
  assign \new_[10725]_  = \new_[10724]_  & \new_[10719]_ ;
  assign \new_[10729]_  = ~A268 & ~A266;
  assign \new_[10730]_  = ~A265 & \new_[10729]_ ;
  assign \new_[10734]_  = A302 & ~A299;
  assign \new_[10735]_  = A298 & \new_[10734]_ ;
  assign \new_[10736]_  = \new_[10735]_  & \new_[10730]_ ;
  assign \new_[10739]_  = A167 & A168;
  assign \new_[10743]_  = ~A203 & ~A202;
  assign \new_[10744]_  = ~A201 & \new_[10743]_ ;
  assign \new_[10745]_  = \new_[10744]_  & \new_[10739]_ ;
  assign \new_[10749]_  = ~A268 & ~A266;
  assign \new_[10750]_  = ~A265 & \new_[10749]_ ;
  assign \new_[10754]_  = A302 & A299;
  assign \new_[10755]_  = ~A298 & \new_[10754]_ ;
  assign \new_[10756]_  = \new_[10755]_  & \new_[10750]_ ;
  assign \new_[10759]_  = A167 & A168;
  assign \new_[10763]_  = ~A265 & A201;
  assign \new_[10764]_  = A199 & \new_[10763]_ ;
  assign \new_[10765]_  = \new_[10764]_  & \new_[10759]_ ;
  assign \new_[10769]_  = A298 & A269;
  assign \new_[10770]_  = A266 & \new_[10769]_ ;
  assign \new_[10774]_  = ~A301 & ~A300;
  assign \new_[10775]_  = A299 & \new_[10774]_ ;
  assign \new_[10776]_  = \new_[10775]_  & \new_[10770]_ ;
  assign \new_[10779]_  = A167 & A168;
  assign \new_[10783]_  = A265 & A201;
  assign \new_[10784]_  = A199 & \new_[10783]_ ;
  assign \new_[10785]_  = \new_[10784]_  & \new_[10779]_ ;
  assign \new_[10789]_  = A298 & A269;
  assign \new_[10790]_  = ~A266 & \new_[10789]_ ;
  assign \new_[10794]_  = ~A301 & ~A300;
  assign \new_[10795]_  = A299 & \new_[10794]_ ;
  assign \new_[10796]_  = \new_[10795]_  & \new_[10790]_ ;
  assign \new_[10799]_  = A167 & A168;
  assign \new_[10803]_  = ~A265 & A201;
  assign \new_[10804]_  = A200 & \new_[10803]_ ;
  assign \new_[10805]_  = \new_[10804]_  & \new_[10799]_ ;
  assign \new_[10809]_  = A298 & A269;
  assign \new_[10810]_  = A266 & \new_[10809]_ ;
  assign \new_[10814]_  = ~A301 & ~A300;
  assign \new_[10815]_  = A299 & \new_[10814]_ ;
  assign \new_[10816]_  = \new_[10815]_  & \new_[10810]_ ;
  assign \new_[10819]_  = A167 & A168;
  assign \new_[10823]_  = A265 & A201;
  assign \new_[10824]_  = A200 & \new_[10823]_ ;
  assign \new_[10825]_  = \new_[10824]_  & \new_[10819]_ ;
  assign \new_[10829]_  = A298 & A269;
  assign \new_[10830]_  = ~A266 & \new_[10829]_ ;
  assign \new_[10834]_  = ~A301 & ~A300;
  assign \new_[10835]_  = A299 & \new_[10834]_ ;
  assign \new_[10836]_  = \new_[10835]_  & \new_[10830]_ ;
  assign \new_[10839]_  = A167 & A168;
  assign \new_[10843]_  = ~A201 & A200;
  assign \new_[10844]_  = A199 & \new_[10843]_ ;
  assign \new_[10845]_  = \new_[10844]_  & \new_[10839]_ ;
  assign \new_[10849]_  = ~A268 & ~A267;
  assign \new_[10850]_  = ~A202 & \new_[10849]_ ;
  assign \new_[10854]_  = A300 & A299;
  assign \new_[10855]_  = ~A269 & \new_[10854]_ ;
  assign \new_[10856]_  = \new_[10855]_  & \new_[10850]_ ;
  assign \new_[10859]_  = A167 & A168;
  assign \new_[10863]_  = ~A201 & A200;
  assign \new_[10864]_  = A199 & \new_[10863]_ ;
  assign \new_[10865]_  = \new_[10864]_  & \new_[10859]_ ;
  assign \new_[10869]_  = ~A268 & ~A267;
  assign \new_[10870]_  = ~A202 & \new_[10869]_ ;
  assign \new_[10874]_  = A300 & A298;
  assign \new_[10875]_  = ~A269 & \new_[10874]_ ;
  assign \new_[10876]_  = \new_[10875]_  & \new_[10870]_ ;
  assign \new_[10879]_  = A167 & A168;
  assign \new_[10883]_  = ~A201 & A200;
  assign \new_[10884]_  = A199 & \new_[10883]_ ;
  assign \new_[10885]_  = \new_[10884]_  & \new_[10879]_ ;
  assign \new_[10889]_  = A266 & A265;
  assign \new_[10890]_  = ~A202 & \new_[10889]_ ;
  assign \new_[10894]_  = A301 & ~A268;
  assign \new_[10895]_  = ~A267 & \new_[10894]_ ;
  assign \new_[10896]_  = \new_[10895]_  & \new_[10890]_ ;
  assign \new_[10899]_  = A167 & A168;
  assign \new_[10903]_  = ~A201 & A200;
  assign \new_[10904]_  = A199 & \new_[10903]_ ;
  assign \new_[10905]_  = \new_[10904]_  & \new_[10899]_ ;
  assign \new_[10909]_  = ~A266 & ~A265;
  assign \new_[10910]_  = ~A202 & \new_[10909]_ ;
  assign \new_[10914]_  = A300 & A299;
  assign \new_[10915]_  = ~A268 & \new_[10914]_ ;
  assign \new_[10916]_  = \new_[10915]_  & \new_[10910]_ ;
  assign \new_[10919]_  = A167 & A168;
  assign \new_[10923]_  = ~A201 & A200;
  assign \new_[10924]_  = A199 & \new_[10923]_ ;
  assign \new_[10925]_  = \new_[10924]_  & \new_[10919]_ ;
  assign \new_[10929]_  = ~A266 & ~A265;
  assign \new_[10930]_  = ~A202 & \new_[10929]_ ;
  assign \new_[10934]_  = A300 & A298;
  assign \new_[10935]_  = ~A268 & \new_[10934]_ ;
  assign \new_[10936]_  = \new_[10935]_  & \new_[10930]_ ;
  assign \new_[10939]_  = A167 & A168;
  assign \new_[10943]_  = A203 & A200;
  assign \new_[10944]_  = ~A199 & \new_[10943]_ ;
  assign \new_[10945]_  = \new_[10944]_  & \new_[10939]_ ;
  assign \new_[10949]_  = A298 & A267;
  assign \new_[10950]_  = A265 & \new_[10949]_ ;
  assign \new_[10954]_  = ~A301 & ~A300;
  assign \new_[10955]_  = A299 & \new_[10954]_ ;
  assign \new_[10956]_  = \new_[10955]_  & \new_[10950]_ ;
  assign \new_[10959]_  = A167 & A168;
  assign \new_[10963]_  = A203 & A200;
  assign \new_[10964]_  = ~A199 & \new_[10963]_ ;
  assign \new_[10965]_  = \new_[10964]_  & \new_[10959]_ ;
  assign \new_[10969]_  = A298 & A267;
  assign \new_[10970]_  = A266 & \new_[10969]_ ;
  assign \new_[10974]_  = ~A301 & ~A300;
  assign \new_[10975]_  = A299 & \new_[10974]_ ;
  assign \new_[10976]_  = \new_[10975]_  & \new_[10970]_ ;
  assign \new_[10979]_  = A167 & A168;
  assign \new_[10983]_  = A203 & A200;
  assign \new_[10984]_  = ~A199 & \new_[10983]_ ;
  assign \new_[10985]_  = \new_[10984]_  & \new_[10979]_ ;
  assign \new_[10989]_  = A269 & A266;
  assign \new_[10990]_  = ~A265 & \new_[10989]_ ;
  assign \new_[10994]_  = ~A302 & ~A301;
  assign \new_[10995]_  = ~A300 & \new_[10994]_ ;
  assign \new_[10996]_  = \new_[10995]_  & \new_[10990]_ ;
  assign \new_[10999]_  = A167 & A168;
  assign \new_[11003]_  = A203 & A200;
  assign \new_[11004]_  = ~A199 & \new_[11003]_ ;
  assign \new_[11005]_  = \new_[11004]_  & \new_[10999]_ ;
  assign \new_[11009]_  = A269 & A266;
  assign \new_[11010]_  = ~A265 & \new_[11009]_ ;
  assign \new_[11014]_  = ~A301 & ~A299;
  assign \new_[11015]_  = ~A298 & \new_[11014]_ ;
  assign \new_[11016]_  = \new_[11015]_  & \new_[11010]_ ;
  assign \new_[11019]_  = A167 & A168;
  assign \new_[11023]_  = A203 & A200;
  assign \new_[11024]_  = ~A199 & \new_[11023]_ ;
  assign \new_[11025]_  = \new_[11024]_  & \new_[11019]_ ;
  assign \new_[11029]_  = A269 & ~A266;
  assign \new_[11030]_  = A265 & \new_[11029]_ ;
  assign \new_[11034]_  = ~A302 & ~A301;
  assign \new_[11035]_  = ~A300 & \new_[11034]_ ;
  assign \new_[11036]_  = \new_[11035]_  & \new_[11030]_ ;
  assign \new_[11039]_  = A167 & A168;
  assign \new_[11043]_  = A203 & A200;
  assign \new_[11044]_  = ~A199 & \new_[11043]_ ;
  assign \new_[11045]_  = \new_[11044]_  & \new_[11039]_ ;
  assign \new_[11049]_  = A269 & ~A266;
  assign \new_[11050]_  = A265 & \new_[11049]_ ;
  assign \new_[11054]_  = ~A301 & ~A299;
  assign \new_[11055]_  = ~A298 & \new_[11054]_ ;
  assign \new_[11056]_  = \new_[11055]_  & \new_[11050]_ ;
  assign \new_[11059]_  = A167 & A168;
  assign \new_[11063]_  = A203 & ~A200;
  assign \new_[11064]_  = A199 & \new_[11063]_ ;
  assign \new_[11065]_  = \new_[11064]_  & \new_[11059]_ ;
  assign \new_[11069]_  = A298 & A267;
  assign \new_[11070]_  = A265 & \new_[11069]_ ;
  assign \new_[11074]_  = ~A301 & ~A300;
  assign \new_[11075]_  = A299 & \new_[11074]_ ;
  assign \new_[11076]_  = \new_[11075]_  & \new_[11070]_ ;
  assign \new_[11079]_  = A167 & A168;
  assign \new_[11083]_  = A203 & ~A200;
  assign \new_[11084]_  = A199 & \new_[11083]_ ;
  assign \new_[11085]_  = \new_[11084]_  & \new_[11079]_ ;
  assign \new_[11089]_  = A298 & A267;
  assign \new_[11090]_  = A266 & \new_[11089]_ ;
  assign \new_[11094]_  = ~A301 & ~A300;
  assign \new_[11095]_  = A299 & \new_[11094]_ ;
  assign \new_[11096]_  = \new_[11095]_  & \new_[11090]_ ;
  assign \new_[11099]_  = A167 & A168;
  assign \new_[11103]_  = A203 & ~A200;
  assign \new_[11104]_  = A199 & \new_[11103]_ ;
  assign \new_[11105]_  = \new_[11104]_  & \new_[11099]_ ;
  assign \new_[11109]_  = A269 & A266;
  assign \new_[11110]_  = ~A265 & \new_[11109]_ ;
  assign \new_[11114]_  = ~A302 & ~A301;
  assign \new_[11115]_  = ~A300 & \new_[11114]_ ;
  assign \new_[11116]_  = \new_[11115]_  & \new_[11110]_ ;
  assign \new_[11119]_  = A167 & A168;
  assign \new_[11123]_  = A203 & ~A200;
  assign \new_[11124]_  = A199 & \new_[11123]_ ;
  assign \new_[11125]_  = \new_[11124]_  & \new_[11119]_ ;
  assign \new_[11129]_  = A269 & A266;
  assign \new_[11130]_  = ~A265 & \new_[11129]_ ;
  assign \new_[11134]_  = ~A301 & ~A299;
  assign \new_[11135]_  = ~A298 & \new_[11134]_ ;
  assign \new_[11136]_  = \new_[11135]_  & \new_[11130]_ ;
  assign \new_[11139]_  = A167 & A168;
  assign \new_[11143]_  = A203 & ~A200;
  assign \new_[11144]_  = A199 & \new_[11143]_ ;
  assign \new_[11145]_  = \new_[11144]_  & \new_[11139]_ ;
  assign \new_[11149]_  = A269 & ~A266;
  assign \new_[11150]_  = A265 & \new_[11149]_ ;
  assign \new_[11154]_  = ~A302 & ~A301;
  assign \new_[11155]_  = ~A300 & \new_[11154]_ ;
  assign \new_[11156]_  = \new_[11155]_  & \new_[11150]_ ;
  assign \new_[11159]_  = A167 & A168;
  assign \new_[11163]_  = A203 & ~A200;
  assign \new_[11164]_  = A199 & \new_[11163]_ ;
  assign \new_[11165]_  = \new_[11164]_  & \new_[11159]_ ;
  assign \new_[11169]_  = A269 & ~A266;
  assign \new_[11170]_  = A265 & \new_[11169]_ ;
  assign \new_[11174]_  = ~A301 & ~A299;
  assign \new_[11175]_  = ~A298 & \new_[11174]_ ;
  assign \new_[11176]_  = \new_[11175]_  & \new_[11170]_ ;
  assign \new_[11179]_  = A167 & A168;
  assign \new_[11183]_  = ~A202 & ~A200;
  assign \new_[11184]_  = ~A199 & \new_[11183]_ ;
  assign \new_[11185]_  = \new_[11184]_  & \new_[11179]_ ;
  assign \new_[11189]_  = ~A269 & ~A268;
  assign \new_[11190]_  = ~A267 & \new_[11189]_ ;
  assign \new_[11194]_  = A302 & ~A299;
  assign \new_[11195]_  = A298 & \new_[11194]_ ;
  assign \new_[11196]_  = \new_[11195]_  & \new_[11190]_ ;
  assign \new_[11199]_  = A167 & A168;
  assign \new_[11203]_  = ~A202 & ~A200;
  assign \new_[11204]_  = ~A199 & \new_[11203]_ ;
  assign \new_[11205]_  = \new_[11204]_  & \new_[11199]_ ;
  assign \new_[11209]_  = ~A269 & ~A268;
  assign \new_[11210]_  = ~A267 & \new_[11209]_ ;
  assign \new_[11214]_  = A302 & A299;
  assign \new_[11215]_  = ~A298 & \new_[11214]_ ;
  assign \new_[11216]_  = \new_[11215]_  & \new_[11210]_ ;
  assign \new_[11219]_  = A167 & A168;
  assign \new_[11223]_  = ~A202 & ~A200;
  assign \new_[11224]_  = ~A199 & \new_[11223]_ ;
  assign \new_[11225]_  = \new_[11224]_  & \new_[11219]_ ;
  assign \new_[11229]_  = ~A267 & A266;
  assign \new_[11230]_  = A265 & \new_[11229]_ ;
  assign \new_[11234]_  = A300 & A299;
  assign \new_[11235]_  = ~A268 & \new_[11234]_ ;
  assign \new_[11236]_  = \new_[11235]_  & \new_[11230]_ ;
  assign \new_[11239]_  = A167 & A168;
  assign \new_[11243]_  = ~A202 & ~A200;
  assign \new_[11244]_  = ~A199 & \new_[11243]_ ;
  assign \new_[11245]_  = \new_[11244]_  & \new_[11239]_ ;
  assign \new_[11249]_  = ~A267 & A266;
  assign \new_[11250]_  = A265 & \new_[11249]_ ;
  assign \new_[11254]_  = A300 & A298;
  assign \new_[11255]_  = ~A268 & \new_[11254]_ ;
  assign \new_[11256]_  = \new_[11255]_  & \new_[11250]_ ;
  assign \new_[11259]_  = A167 & A168;
  assign \new_[11263]_  = ~A202 & ~A200;
  assign \new_[11264]_  = ~A199 & \new_[11263]_ ;
  assign \new_[11265]_  = \new_[11264]_  & \new_[11259]_ ;
  assign \new_[11269]_  = ~A268 & ~A266;
  assign \new_[11270]_  = ~A265 & \new_[11269]_ ;
  assign \new_[11274]_  = A302 & ~A299;
  assign \new_[11275]_  = A298 & \new_[11274]_ ;
  assign \new_[11276]_  = \new_[11275]_  & \new_[11270]_ ;
  assign \new_[11279]_  = A167 & A168;
  assign \new_[11283]_  = ~A202 & ~A200;
  assign \new_[11284]_  = ~A199 & \new_[11283]_ ;
  assign \new_[11285]_  = \new_[11284]_  & \new_[11279]_ ;
  assign \new_[11289]_  = ~A268 & ~A266;
  assign \new_[11290]_  = ~A265 & \new_[11289]_ ;
  assign \new_[11294]_  = A302 & A299;
  assign \new_[11295]_  = ~A298 & \new_[11294]_ ;
  assign \new_[11296]_  = \new_[11295]_  & \new_[11290]_ ;
  assign \new_[11299]_  = A167 & A170;
  assign \new_[11303]_  = ~A265 & A202;
  assign \new_[11304]_  = ~A166 & \new_[11303]_ ;
  assign \new_[11305]_  = \new_[11304]_  & \new_[11299]_ ;
  assign \new_[11309]_  = A298 & A269;
  assign \new_[11310]_  = A266 & \new_[11309]_ ;
  assign \new_[11314]_  = ~A301 & ~A300;
  assign \new_[11315]_  = A299 & \new_[11314]_ ;
  assign \new_[11316]_  = \new_[11315]_  & \new_[11310]_ ;
  assign \new_[11319]_  = A167 & A170;
  assign \new_[11323]_  = A265 & A202;
  assign \new_[11324]_  = ~A166 & \new_[11323]_ ;
  assign \new_[11325]_  = \new_[11324]_  & \new_[11319]_ ;
  assign \new_[11329]_  = A298 & A269;
  assign \new_[11330]_  = ~A266 & \new_[11329]_ ;
  assign \new_[11334]_  = ~A301 & ~A300;
  assign \new_[11335]_  = A299 & \new_[11334]_ ;
  assign \new_[11336]_  = \new_[11335]_  & \new_[11330]_ ;
  assign \new_[11339]_  = A167 & A170;
  assign \new_[11343]_  = ~A202 & ~A201;
  assign \new_[11344]_  = ~A166 & \new_[11343]_ ;
  assign \new_[11345]_  = \new_[11344]_  & \new_[11339]_ ;
  assign \new_[11349]_  = ~A268 & ~A267;
  assign \new_[11350]_  = ~A203 & \new_[11349]_ ;
  assign \new_[11354]_  = A300 & A299;
  assign \new_[11355]_  = ~A269 & \new_[11354]_ ;
  assign \new_[11356]_  = \new_[11355]_  & \new_[11350]_ ;
  assign \new_[11359]_  = A167 & A170;
  assign \new_[11363]_  = ~A202 & ~A201;
  assign \new_[11364]_  = ~A166 & \new_[11363]_ ;
  assign \new_[11365]_  = \new_[11364]_  & \new_[11359]_ ;
  assign \new_[11369]_  = ~A268 & ~A267;
  assign \new_[11370]_  = ~A203 & \new_[11369]_ ;
  assign \new_[11374]_  = A300 & A298;
  assign \new_[11375]_  = ~A269 & \new_[11374]_ ;
  assign \new_[11376]_  = \new_[11375]_  & \new_[11370]_ ;
  assign \new_[11379]_  = A167 & A170;
  assign \new_[11383]_  = ~A202 & ~A201;
  assign \new_[11384]_  = ~A166 & \new_[11383]_ ;
  assign \new_[11385]_  = \new_[11384]_  & \new_[11379]_ ;
  assign \new_[11389]_  = A266 & A265;
  assign \new_[11390]_  = ~A203 & \new_[11389]_ ;
  assign \new_[11394]_  = A301 & ~A268;
  assign \new_[11395]_  = ~A267 & \new_[11394]_ ;
  assign \new_[11396]_  = \new_[11395]_  & \new_[11390]_ ;
  assign \new_[11399]_  = A167 & A170;
  assign \new_[11403]_  = ~A202 & ~A201;
  assign \new_[11404]_  = ~A166 & \new_[11403]_ ;
  assign \new_[11405]_  = \new_[11404]_  & \new_[11399]_ ;
  assign \new_[11409]_  = ~A266 & ~A265;
  assign \new_[11410]_  = ~A203 & \new_[11409]_ ;
  assign \new_[11414]_  = A300 & A299;
  assign \new_[11415]_  = ~A268 & \new_[11414]_ ;
  assign \new_[11416]_  = \new_[11415]_  & \new_[11410]_ ;
  assign \new_[11419]_  = A167 & A170;
  assign \new_[11423]_  = ~A202 & ~A201;
  assign \new_[11424]_  = ~A166 & \new_[11423]_ ;
  assign \new_[11425]_  = \new_[11424]_  & \new_[11419]_ ;
  assign \new_[11429]_  = ~A266 & ~A265;
  assign \new_[11430]_  = ~A203 & \new_[11429]_ ;
  assign \new_[11434]_  = A300 & A298;
  assign \new_[11435]_  = ~A268 & \new_[11434]_ ;
  assign \new_[11436]_  = \new_[11435]_  & \new_[11430]_ ;
  assign \new_[11439]_  = A167 & A170;
  assign \new_[11443]_  = A201 & A199;
  assign \new_[11444]_  = ~A166 & \new_[11443]_ ;
  assign \new_[11445]_  = \new_[11444]_  & \new_[11439]_ ;
  assign \new_[11449]_  = A298 & A267;
  assign \new_[11450]_  = A265 & \new_[11449]_ ;
  assign \new_[11454]_  = ~A301 & ~A300;
  assign \new_[11455]_  = A299 & \new_[11454]_ ;
  assign \new_[11456]_  = \new_[11455]_  & \new_[11450]_ ;
  assign \new_[11459]_  = A167 & A170;
  assign \new_[11463]_  = A201 & A199;
  assign \new_[11464]_  = ~A166 & \new_[11463]_ ;
  assign \new_[11465]_  = \new_[11464]_  & \new_[11459]_ ;
  assign \new_[11469]_  = A298 & A267;
  assign \new_[11470]_  = A266 & \new_[11469]_ ;
  assign \new_[11474]_  = ~A301 & ~A300;
  assign \new_[11475]_  = A299 & \new_[11474]_ ;
  assign \new_[11476]_  = \new_[11475]_  & \new_[11470]_ ;
  assign \new_[11479]_  = A167 & A170;
  assign \new_[11483]_  = A201 & A199;
  assign \new_[11484]_  = ~A166 & \new_[11483]_ ;
  assign \new_[11485]_  = \new_[11484]_  & \new_[11479]_ ;
  assign \new_[11489]_  = A269 & A266;
  assign \new_[11490]_  = ~A265 & \new_[11489]_ ;
  assign \new_[11494]_  = ~A302 & ~A301;
  assign \new_[11495]_  = ~A300 & \new_[11494]_ ;
  assign \new_[11496]_  = \new_[11495]_  & \new_[11490]_ ;
  assign \new_[11499]_  = A167 & A170;
  assign \new_[11503]_  = A201 & A199;
  assign \new_[11504]_  = ~A166 & \new_[11503]_ ;
  assign \new_[11505]_  = \new_[11504]_  & \new_[11499]_ ;
  assign \new_[11509]_  = A269 & A266;
  assign \new_[11510]_  = ~A265 & \new_[11509]_ ;
  assign \new_[11514]_  = ~A301 & ~A299;
  assign \new_[11515]_  = ~A298 & \new_[11514]_ ;
  assign \new_[11516]_  = \new_[11515]_  & \new_[11510]_ ;
  assign \new_[11519]_  = A167 & A170;
  assign \new_[11523]_  = A201 & A199;
  assign \new_[11524]_  = ~A166 & \new_[11523]_ ;
  assign \new_[11525]_  = \new_[11524]_  & \new_[11519]_ ;
  assign \new_[11529]_  = A269 & ~A266;
  assign \new_[11530]_  = A265 & \new_[11529]_ ;
  assign \new_[11534]_  = ~A302 & ~A301;
  assign \new_[11535]_  = ~A300 & \new_[11534]_ ;
  assign \new_[11536]_  = \new_[11535]_  & \new_[11530]_ ;
  assign \new_[11539]_  = A167 & A170;
  assign \new_[11543]_  = A201 & A199;
  assign \new_[11544]_  = ~A166 & \new_[11543]_ ;
  assign \new_[11545]_  = \new_[11544]_  & \new_[11539]_ ;
  assign \new_[11549]_  = A269 & ~A266;
  assign \new_[11550]_  = A265 & \new_[11549]_ ;
  assign \new_[11554]_  = ~A301 & ~A299;
  assign \new_[11555]_  = ~A298 & \new_[11554]_ ;
  assign \new_[11556]_  = \new_[11555]_  & \new_[11550]_ ;
  assign \new_[11559]_  = A167 & A170;
  assign \new_[11563]_  = A201 & A200;
  assign \new_[11564]_  = ~A166 & \new_[11563]_ ;
  assign \new_[11565]_  = \new_[11564]_  & \new_[11559]_ ;
  assign \new_[11569]_  = A298 & A267;
  assign \new_[11570]_  = A265 & \new_[11569]_ ;
  assign \new_[11574]_  = ~A301 & ~A300;
  assign \new_[11575]_  = A299 & \new_[11574]_ ;
  assign \new_[11576]_  = \new_[11575]_  & \new_[11570]_ ;
  assign \new_[11579]_  = A167 & A170;
  assign \new_[11583]_  = A201 & A200;
  assign \new_[11584]_  = ~A166 & \new_[11583]_ ;
  assign \new_[11585]_  = \new_[11584]_  & \new_[11579]_ ;
  assign \new_[11589]_  = A298 & A267;
  assign \new_[11590]_  = A266 & \new_[11589]_ ;
  assign \new_[11594]_  = ~A301 & ~A300;
  assign \new_[11595]_  = A299 & \new_[11594]_ ;
  assign \new_[11596]_  = \new_[11595]_  & \new_[11590]_ ;
  assign \new_[11599]_  = A167 & A170;
  assign \new_[11603]_  = A201 & A200;
  assign \new_[11604]_  = ~A166 & \new_[11603]_ ;
  assign \new_[11605]_  = \new_[11604]_  & \new_[11599]_ ;
  assign \new_[11609]_  = A269 & A266;
  assign \new_[11610]_  = ~A265 & \new_[11609]_ ;
  assign \new_[11614]_  = ~A302 & ~A301;
  assign \new_[11615]_  = ~A300 & \new_[11614]_ ;
  assign \new_[11616]_  = \new_[11615]_  & \new_[11610]_ ;
  assign \new_[11619]_  = A167 & A170;
  assign \new_[11623]_  = A201 & A200;
  assign \new_[11624]_  = ~A166 & \new_[11623]_ ;
  assign \new_[11625]_  = \new_[11624]_  & \new_[11619]_ ;
  assign \new_[11629]_  = A269 & A266;
  assign \new_[11630]_  = ~A265 & \new_[11629]_ ;
  assign \new_[11634]_  = ~A301 & ~A299;
  assign \new_[11635]_  = ~A298 & \new_[11634]_ ;
  assign \new_[11636]_  = \new_[11635]_  & \new_[11630]_ ;
  assign \new_[11639]_  = A167 & A170;
  assign \new_[11643]_  = A201 & A200;
  assign \new_[11644]_  = ~A166 & \new_[11643]_ ;
  assign \new_[11645]_  = \new_[11644]_  & \new_[11639]_ ;
  assign \new_[11649]_  = A269 & ~A266;
  assign \new_[11650]_  = A265 & \new_[11649]_ ;
  assign \new_[11654]_  = ~A302 & ~A301;
  assign \new_[11655]_  = ~A300 & \new_[11654]_ ;
  assign \new_[11656]_  = \new_[11655]_  & \new_[11650]_ ;
  assign \new_[11659]_  = A167 & A170;
  assign \new_[11663]_  = A201 & A200;
  assign \new_[11664]_  = ~A166 & \new_[11663]_ ;
  assign \new_[11665]_  = \new_[11664]_  & \new_[11659]_ ;
  assign \new_[11669]_  = A269 & ~A266;
  assign \new_[11670]_  = A265 & \new_[11669]_ ;
  assign \new_[11674]_  = ~A301 & ~A299;
  assign \new_[11675]_  = ~A298 & \new_[11674]_ ;
  assign \new_[11676]_  = \new_[11675]_  & \new_[11670]_ ;
  assign \new_[11679]_  = A167 & A170;
  assign \new_[11683]_  = A200 & A199;
  assign \new_[11684]_  = ~A166 & \new_[11683]_ ;
  assign \new_[11685]_  = \new_[11684]_  & \new_[11679]_ ;
  assign \new_[11689]_  = ~A267 & ~A202;
  assign \new_[11690]_  = ~A201 & \new_[11689]_ ;
  assign \new_[11694]_  = A301 & ~A269;
  assign \new_[11695]_  = ~A268 & \new_[11694]_ ;
  assign \new_[11696]_  = \new_[11695]_  & \new_[11690]_ ;
  assign \new_[11699]_  = A167 & A170;
  assign \new_[11703]_  = A200 & A199;
  assign \new_[11704]_  = ~A166 & \new_[11703]_ ;
  assign \new_[11705]_  = \new_[11704]_  & \new_[11699]_ ;
  assign \new_[11709]_  = ~A265 & ~A202;
  assign \new_[11710]_  = ~A201 & \new_[11709]_ ;
  assign \new_[11714]_  = A301 & ~A268;
  assign \new_[11715]_  = ~A266 & \new_[11714]_ ;
  assign \new_[11716]_  = \new_[11715]_  & \new_[11710]_ ;
  assign \new_[11719]_  = A167 & A170;
  assign \new_[11723]_  = A200 & ~A199;
  assign \new_[11724]_  = ~A166 & \new_[11723]_ ;
  assign \new_[11725]_  = \new_[11724]_  & \new_[11719]_ ;
  assign \new_[11729]_  = A298 & A268;
  assign \new_[11730]_  = A203 & \new_[11729]_ ;
  assign \new_[11734]_  = ~A301 & ~A300;
  assign \new_[11735]_  = A299 & \new_[11734]_ ;
  assign \new_[11736]_  = \new_[11735]_  & \new_[11730]_ ;
  assign \new_[11739]_  = A167 & A170;
  assign \new_[11743]_  = A200 & ~A199;
  assign \new_[11744]_  = ~A166 & \new_[11743]_ ;
  assign \new_[11745]_  = \new_[11744]_  & \new_[11739]_ ;
  assign \new_[11749]_  = A267 & A265;
  assign \new_[11750]_  = A203 & \new_[11749]_ ;
  assign \new_[11754]_  = ~A302 & ~A301;
  assign \new_[11755]_  = ~A300 & \new_[11754]_ ;
  assign \new_[11756]_  = \new_[11755]_  & \new_[11750]_ ;
  assign \new_[11759]_  = A167 & A170;
  assign \new_[11763]_  = A200 & ~A199;
  assign \new_[11764]_  = ~A166 & \new_[11763]_ ;
  assign \new_[11765]_  = \new_[11764]_  & \new_[11759]_ ;
  assign \new_[11769]_  = A267 & A265;
  assign \new_[11770]_  = A203 & \new_[11769]_ ;
  assign \new_[11774]_  = ~A301 & ~A299;
  assign \new_[11775]_  = ~A298 & \new_[11774]_ ;
  assign \new_[11776]_  = \new_[11775]_  & \new_[11770]_ ;
  assign \new_[11779]_  = A167 & A170;
  assign \new_[11783]_  = A200 & ~A199;
  assign \new_[11784]_  = ~A166 & \new_[11783]_ ;
  assign \new_[11785]_  = \new_[11784]_  & \new_[11779]_ ;
  assign \new_[11789]_  = A267 & A266;
  assign \new_[11790]_  = A203 & \new_[11789]_ ;
  assign \new_[11794]_  = ~A302 & ~A301;
  assign \new_[11795]_  = ~A300 & \new_[11794]_ ;
  assign \new_[11796]_  = \new_[11795]_  & \new_[11790]_ ;
  assign \new_[11799]_  = A167 & A170;
  assign \new_[11803]_  = A200 & ~A199;
  assign \new_[11804]_  = ~A166 & \new_[11803]_ ;
  assign \new_[11805]_  = \new_[11804]_  & \new_[11799]_ ;
  assign \new_[11809]_  = A267 & A266;
  assign \new_[11810]_  = A203 & \new_[11809]_ ;
  assign \new_[11814]_  = ~A301 & ~A299;
  assign \new_[11815]_  = ~A298 & \new_[11814]_ ;
  assign \new_[11816]_  = \new_[11815]_  & \new_[11810]_ ;
  assign \new_[11819]_  = A167 & A170;
  assign \new_[11823]_  = ~A200 & A199;
  assign \new_[11824]_  = ~A166 & \new_[11823]_ ;
  assign \new_[11825]_  = \new_[11824]_  & \new_[11819]_ ;
  assign \new_[11829]_  = A298 & A268;
  assign \new_[11830]_  = A203 & \new_[11829]_ ;
  assign \new_[11834]_  = ~A301 & ~A300;
  assign \new_[11835]_  = A299 & \new_[11834]_ ;
  assign \new_[11836]_  = \new_[11835]_  & \new_[11830]_ ;
  assign \new_[11839]_  = A167 & A170;
  assign \new_[11843]_  = ~A200 & A199;
  assign \new_[11844]_  = ~A166 & \new_[11843]_ ;
  assign \new_[11845]_  = \new_[11844]_  & \new_[11839]_ ;
  assign \new_[11849]_  = A267 & A265;
  assign \new_[11850]_  = A203 & \new_[11849]_ ;
  assign \new_[11854]_  = ~A302 & ~A301;
  assign \new_[11855]_  = ~A300 & \new_[11854]_ ;
  assign \new_[11856]_  = \new_[11855]_  & \new_[11850]_ ;
  assign \new_[11859]_  = A167 & A170;
  assign \new_[11863]_  = ~A200 & A199;
  assign \new_[11864]_  = ~A166 & \new_[11863]_ ;
  assign \new_[11865]_  = \new_[11864]_  & \new_[11859]_ ;
  assign \new_[11869]_  = A267 & A265;
  assign \new_[11870]_  = A203 & \new_[11869]_ ;
  assign \new_[11874]_  = ~A301 & ~A299;
  assign \new_[11875]_  = ~A298 & \new_[11874]_ ;
  assign \new_[11876]_  = \new_[11875]_  & \new_[11870]_ ;
  assign \new_[11879]_  = A167 & A170;
  assign \new_[11883]_  = ~A200 & A199;
  assign \new_[11884]_  = ~A166 & \new_[11883]_ ;
  assign \new_[11885]_  = \new_[11884]_  & \new_[11879]_ ;
  assign \new_[11889]_  = A267 & A266;
  assign \new_[11890]_  = A203 & \new_[11889]_ ;
  assign \new_[11894]_  = ~A302 & ~A301;
  assign \new_[11895]_  = ~A300 & \new_[11894]_ ;
  assign \new_[11896]_  = \new_[11895]_  & \new_[11890]_ ;
  assign \new_[11899]_  = A167 & A170;
  assign \new_[11903]_  = ~A200 & A199;
  assign \new_[11904]_  = ~A166 & \new_[11903]_ ;
  assign \new_[11905]_  = \new_[11904]_  & \new_[11899]_ ;
  assign \new_[11909]_  = A267 & A266;
  assign \new_[11910]_  = A203 & \new_[11909]_ ;
  assign \new_[11914]_  = ~A301 & ~A299;
  assign \new_[11915]_  = ~A298 & \new_[11914]_ ;
  assign \new_[11916]_  = \new_[11915]_  & \new_[11910]_ ;
  assign \new_[11919]_  = A167 & A170;
  assign \new_[11923]_  = ~A200 & ~A199;
  assign \new_[11924]_  = ~A166 & \new_[11923]_ ;
  assign \new_[11925]_  = \new_[11924]_  & \new_[11919]_ ;
  assign \new_[11929]_  = ~A268 & ~A267;
  assign \new_[11930]_  = ~A202 & \new_[11929]_ ;
  assign \new_[11934]_  = A300 & A299;
  assign \new_[11935]_  = ~A269 & \new_[11934]_ ;
  assign \new_[11936]_  = \new_[11935]_  & \new_[11930]_ ;
  assign \new_[11939]_  = A167 & A170;
  assign \new_[11943]_  = ~A200 & ~A199;
  assign \new_[11944]_  = ~A166 & \new_[11943]_ ;
  assign \new_[11945]_  = \new_[11944]_  & \new_[11939]_ ;
  assign \new_[11949]_  = ~A268 & ~A267;
  assign \new_[11950]_  = ~A202 & \new_[11949]_ ;
  assign \new_[11954]_  = A300 & A298;
  assign \new_[11955]_  = ~A269 & \new_[11954]_ ;
  assign \new_[11956]_  = \new_[11955]_  & \new_[11950]_ ;
  assign \new_[11959]_  = A167 & A170;
  assign \new_[11963]_  = ~A200 & ~A199;
  assign \new_[11964]_  = ~A166 & \new_[11963]_ ;
  assign \new_[11965]_  = \new_[11964]_  & \new_[11959]_ ;
  assign \new_[11969]_  = A266 & A265;
  assign \new_[11970]_  = ~A202 & \new_[11969]_ ;
  assign \new_[11974]_  = A301 & ~A268;
  assign \new_[11975]_  = ~A267 & \new_[11974]_ ;
  assign \new_[11976]_  = \new_[11975]_  & \new_[11970]_ ;
  assign \new_[11979]_  = A167 & A170;
  assign \new_[11983]_  = ~A200 & ~A199;
  assign \new_[11984]_  = ~A166 & \new_[11983]_ ;
  assign \new_[11985]_  = \new_[11984]_  & \new_[11979]_ ;
  assign \new_[11989]_  = ~A266 & ~A265;
  assign \new_[11990]_  = ~A202 & \new_[11989]_ ;
  assign \new_[11994]_  = A300 & A299;
  assign \new_[11995]_  = ~A268 & \new_[11994]_ ;
  assign \new_[11996]_  = \new_[11995]_  & \new_[11990]_ ;
  assign \new_[11999]_  = A167 & A170;
  assign \new_[12003]_  = ~A200 & ~A199;
  assign \new_[12004]_  = ~A166 & \new_[12003]_ ;
  assign \new_[12005]_  = \new_[12004]_  & \new_[11999]_ ;
  assign \new_[12009]_  = ~A266 & ~A265;
  assign \new_[12010]_  = ~A202 & \new_[12009]_ ;
  assign \new_[12014]_  = A300 & A298;
  assign \new_[12015]_  = ~A268 & \new_[12014]_ ;
  assign \new_[12016]_  = \new_[12015]_  & \new_[12010]_ ;
  assign \new_[12019]_  = ~A167 & A170;
  assign \new_[12023]_  = ~A265 & A202;
  assign \new_[12024]_  = A166 & \new_[12023]_ ;
  assign \new_[12025]_  = \new_[12024]_  & \new_[12019]_ ;
  assign \new_[12029]_  = A298 & A269;
  assign \new_[12030]_  = A266 & \new_[12029]_ ;
  assign \new_[12034]_  = ~A301 & ~A300;
  assign \new_[12035]_  = A299 & \new_[12034]_ ;
  assign \new_[12036]_  = \new_[12035]_  & \new_[12030]_ ;
  assign \new_[12039]_  = ~A167 & A170;
  assign \new_[12043]_  = A265 & A202;
  assign \new_[12044]_  = A166 & \new_[12043]_ ;
  assign \new_[12045]_  = \new_[12044]_  & \new_[12039]_ ;
  assign \new_[12049]_  = A298 & A269;
  assign \new_[12050]_  = ~A266 & \new_[12049]_ ;
  assign \new_[12054]_  = ~A301 & ~A300;
  assign \new_[12055]_  = A299 & \new_[12054]_ ;
  assign \new_[12056]_  = \new_[12055]_  & \new_[12050]_ ;
  assign \new_[12059]_  = ~A167 & A170;
  assign \new_[12063]_  = ~A202 & ~A201;
  assign \new_[12064]_  = A166 & \new_[12063]_ ;
  assign \new_[12065]_  = \new_[12064]_  & \new_[12059]_ ;
  assign \new_[12069]_  = ~A268 & ~A267;
  assign \new_[12070]_  = ~A203 & \new_[12069]_ ;
  assign \new_[12074]_  = A300 & A299;
  assign \new_[12075]_  = ~A269 & \new_[12074]_ ;
  assign \new_[12076]_  = \new_[12075]_  & \new_[12070]_ ;
  assign \new_[12079]_  = ~A167 & A170;
  assign \new_[12083]_  = ~A202 & ~A201;
  assign \new_[12084]_  = A166 & \new_[12083]_ ;
  assign \new_[12085]_  = \new_[12084]_  & \new_[12079]_ ;
  assign \new_[12089]_  = ~A268 & ~A267;
  assign \new_[12090]_  = ~A203 & \new_[12089]_ ;
  assign \new_[12094]_  = A300 & A298;
  assign \new_[12095]_  = ~A269 & \new_[12094]_ ;
  assign \new_[12096]_  = \new_[12095]_  & \new_[12090]_ ;
  assign \new_[12099]_  = ~A167 & A170;
  assign \new_[12103]_  = ~A202 & ~A201;
  assign \new_[12104]_  = A166 & \new_[12103]_ ;
  assign \new_[12105]_  = \new_[12104]_  & \new_[12099]_ ;
  assign \new_[12109]_  = A266 & A265;
  assign \new_[12110]_  = ~A203 & \new_[12109]_ ;
  assign \new_[12114]_  = A301 & ~A268;
  assign \new_[12115]_  = ~A267 & \new_[12114]_ ;
  assign \new_[12116]_  = \new_[12115]_  & \new_[12110]_ ;
  assign \new_[12119]_  = ~A167 & A170;
  assign \new_[12123]_  = ~A202 & ~A201;
  assign \new_[12124]_  = A166 & \new_[12123]_ ;
  assign \new_[12125]_  = \new_[12124]_  & \new_[12119]_ ;
  assign \new_[12129]_  = ~A266 & ~A265;
  assign \new_[12130]_  = ~A203 & \new_[12129]_ ;
  assign \new_[12134]_  = A300 & A299;
  assign \new_[12135]_  = ~A268 & \new_[12134]_ ;
  assign \new_[12136]_  = \new_[12135]_  & \new_[12130]_ ;
  assign \new_[12139]_  = ~A167 & A170;
  assign \new_[12143]_  = ~A202 & ~A201;
  assign \new_[12144]_  = A166 & \new_[12143]_ ;
  assign \new_[12145]_  = \new_[12144]_  & \new_[12139]_ ;
  assign \new_[12149]_  = ~A266 & ~A265;
  assign \new_[12150]_  = ~A203 & \new_[12149]_ ;
  assign \new_[12154]_  = A300 & A298;
  assign \new_[12155]_  = ~A268 & \new_[12154]_ ;
  assign \new_[12156]_  = \new_[12155]_  & \new_[12150]_ ;
  assign \new_[12159]_  = ~A167 & A170;
  assign \new_[12163]_  = A201 & A199;
  assign \new_[12164]_  = A166 & \new_[12163]_ ;
  assign \new_[12165]_  = \new_[12164]_  & \new_[12159]_ ;
  assign \new_[12169]_  = A298 & A267;
  assign \new_[12170]_  = A265 & \new_[12169]_ ;
  assign \new_[12174]_  = ~A301 & ~A300;
  assign \new_[12175]_  = A299 & \new_[12174]_ ;
  assign \new_[12176]_  = \new_[12175]_  & \new_[12170]_ ;
  assign \new_[12179]_  = ~A167 & A170;
  assign \new_[12183]_  = A201 & A199;
  assign \new_[12184]_  = A166 & \new_[12183]_ ;
  assign \new_[12185]_  = \new_[12184]_  & \new_[12179]_ ;
  assign \new_[12189]_  = A298 & A267;
  assign \new_[12190]_  = A266 & \new_[12189]_ ;
  assign \new_[12194]_  = ~A301 & ~A300;
  assign \new_[12195]_  = A299 & \new_[12194]_ ;
  assign \new_[12196]_  = \new_[12195]_  & \new_[12190]_ ;
  assign \new_[12199]_  = ~A167 & A170;
  assign \new_[12203]_  = A201 & A199;
  assign \new_[12204]_  = A166 & \new_[12203]_ ;
  assign \new_[12205]_  = \new_[12204]_  & \new_[12199]_ ;
  assign \new_[12209]_  = A269 & A266;
  assign \new_[12210]_  = ~A265 & \new_[12209]_ ;
  assign \new_[12214]_  = ~A302 & ~A301;
  assign \new_[12215]_  = ~A300 & \new_[12214]_ ;
  assign \new_[12216]_  = \new_[12215]_  & \new_[12210]_ ;
  assign \new_[12219]_  = ~A167 & A170;
  assign \new_[12223]_  = A201 & A199;
  assign \new_[12224]_  = A166 & \new_[12223]_ ;
  assign \new_[12225]_  = \new_[12224]_  & \new_[12219]_ ;
  assign \new_[12229]_  = A269 & A266;
  assign \new_[12230]_  = ~A265 & \new_[12229]_ ;
  assign \new_[12234]_  = ~A301 & ~A299;
  assign \new_[12235]_  = ~A298 & \new_[12234]_ ;
  assign \new_[12236]_  = \new_[12235]_  & \new_[12230]_ ;
  assign \new_[12239]_  = ~A167 & A170;
  assign \new_[12243]_  = A201 & A199;
  assign \new_[12244]_  = A166 & \new_[12243]_ ;
  assign \new_[12245]_  = \new_[12244]_  & \new_[12239]_ ;
  assign \new_[12249]_  = A269 & ~A266;
  assign \new_[12250]_  = A265 & \new_[12249]_ ;
  assign \new_[12254]_  = ~A302 & ~A301;
  assign \new_[12255]_  = ~A300 & \new_[12254]_ ;
  assign \new_[12256]_  = \new_[12255]_  & \new_[12250]_ ;
  assign \new_[12259]_  = ~A167 & A170;
  assign \new_[12263]_  = A201 & A199;
  assign \new_[12264]_  = A166 & \new_[12263]_ ;
  assign \new_[12265]_  = \new_[12264]_  & \new_[12259]_ ;
  assign \new_[12269]_  = A269 & ~A266;
  assign \new_[12270]_  = A265 & \new_[12269]_ ;
  assign \new_[12274]_  = ~A301 & ~A299;
  assign \new_[12275]_  = ~A298 & \new_[12274]_ ;
  assign \new_[12276]_  = \new_[12275]_  & \new_[12270]_ ;
  assign \new_[12279]_  = ~A167 & A170;
  assign \new_[12283]_  = A201 & A200;
  assign \new_[12284]_  = A166 & \new_[12283]_ ;
  assign \new_[12285]_  = \new_[12284]_  & \new_[12279]_ ;
  assign \new_[12289]_  = A298 & A267;
  assign \new_[12290]_  = A265 & \new_[12289]_ ;
  assign \new_[12294]_  = ~A301 & ~A300;
  assign \new_[12295]_  = A299 & \new_[12294]_ ;
  assign \new_[12296]_  = \new_[12295]_  & \new_[12290]_ ;
  assign \new_[12299]_  = ~A167 & A170;
  assign \new_[12303]_  = A201 & A200;
  assign \new_[12304]_  = A166 & \new_[12303]_ ;
  assign \new_[12305]_  = \new_[12304]_  & \new_[12299]_ ;
  assign \new_[12309]_  = A298 & A267;
  assign \new_[12310]_  = A266 & \new_[12309]_ ;
  assign \new_[12314]_  = ~A301 & ~A300;
  assign \new_[12315]_  = A299 & \new_[12314]_ ;
  assign \new_[12316]_  = \new_[12315]_  & \new_[12310]_ ;
  assign \new_[12319]_  = ~A167 & A170;
  assign \new_[12323]_  = A201 & A200;
  assign \new_[12324]_  = A166 & \new_[12323]_ ;
  assign \new_[12325]_  = \new_[12324]_  & \new_[12319]_ ;
  assign \new_[12329]_  = A269 & A266;
  assign \new_[12330]_  = ~A265 & \new_[12329]_ ;
  assign \new_[12334]_  = ~A302 & ~A301;
  assign \new_[12335]_  = ~A300 & \new_[12334]_ ;
  assign \new_[12336]_  = \new_[12335]_  & \new_[12330]_ ;
  assign \new_[12339]_  = ~A167 & A170;
  assign \new_[12343]_  = A201 & A200;
  assign \new_[12344]_  = A166 & \new_[12343]_ ;
  assign \new_[12345]_  = \new_[12344]_  & \new_[12339]_ ;
  assign \new_[12349]_  = A269 & A266;
  assign \new_[12350]_  = ~A265 & \new_[12349]_ ;
  assign \new_[12354]_  = ~A301 & ~A299;
  assign \new_[12355]_  = ~A298 & \new_[12354]_ ;
  assign \new_[12356]_  = \new_[12355]_  & \new_[12350]_ ;
  assign \new_[12359]_  = ~A167 & A170;
  assign \new_[12363]_  = A201 & A200;
  assign \new_[12364]_  = A166 & \new_[12363]_ ;
  assign \new_[12365]_  = \new_[12364]_  & \new_[12359]_ ;
  assign \new_[12369]_  = A269 & ~A266;
  assign \new_[12370]_  = A265 & \new_[12369]_ ;
  assign \new_[12374]_  = ~A302 & ~A301;
  assign \new_[12375]_  = ~A300 & \new_[12374]_ ;
  assign \new_[12376]_  = \new_[12375]_  & \new_[12370]_ ;
  assign \new_[12379]_  = ~A167 & A170;
  assign \new_[12383]_  = A201 & A200;
  assign \new_[12384]_  = A166 & \new_[12383]_ ;
  assign \new_[12385]_  = \new_[12384]_  & \new_[12379]_ ;
  assign \new_[12389]_  = A269 & ~A266;
  assign \new_[12390]_  = A265 & \new_[12389]_ ;
  assign \new_[12394]_  = ~A301 & ~A299;
  assign \new_[12395]_  = ~A298 & \new_[12394]_ ;
  assign \new_[12396]_  = \new_[12395]_  & \new_[12390]_ ;
  assign \new_[12399]_  = ~A167 & A170;
  assign \new_[12403]_  = A200 & A199;
  assign \new_[12404]_  = A166 & \new_[12403]_ ;
  assign \new_[12405]_  = \new_[12404]_  & \new_[12399]_ ;
  assign \new_[12409]_  = ~A267 & ~A202;
  assign \new_[12410]_  = ~A201 & \new_[12409]_ ;
  assign \new_[12414]_  = A301 & ~A269;
  assign \new_[12415]_  = ~A268 & \new_[12414]_ ;
  assign \new_[12416]_  = \new_[12415]_  & \new_[12410]_ ;
  assign \new_[12419]_  = ~A167 & A170;
  assign \new_[12423]_  = A200 & A199;
  assign \new_[12424]_  = A166 & \new_[12423]_ ;
  assign \new_[12425]_  = \new_[12424]_  & \new_[12419]_ ;
  assign \new_[12429]_  = ~A265 & ~A202;
  assign \new_[12430]_  = ~A201 & \new_[12429]_ ;
  assign \new_[12434]_  = A301 & ~A268;
  assign \new_[12435]_  = ~A266 & \new_[12434]_ ;
  assign \new_[12436]_  = \new_[12435]_  & \new_[12430]_ ;
  assign \new_[12439]_  = ~A167 & A170;
  assign \new_[12443]_  = A200 & ~A199;
  assign \new_[12444]_  = A166 & \new_[12443]_ ;
  assign \new_[12445]_  = \new_[12444]_  & \new_[12439]_ ;
  assign \new_[12449]_  = A298 & A268;
  assign \new_[12450]_  = A203 & \new_[12449]_ ;
  assign \new_[12454]_  = ~A301 & ~A300;
  assign \new_[12455]_  = A299 & \new_[12454]_ ;
  assign \new_[12456]_  = \new_[12455]_  & \new_[12450]_ ;
  assign \new_[12459]_  = ~A167 & A170;
  assign \new_[12463]_  = A200 & ~A199;
  assign \new_[12464]_  = A166 & \new_[12463]_ ;
  assign \new_[12465]_  = \new_[12464]_  & \new_[12459]_ ;
  assign \new_[12469]_  = A267 & A265;
  assign \new_[12470]_  = A203 & \new_[12469]_ ;
  assign \new_[12474]_  = ~A302 & ~A301;
  assign \new_[12475]_  = ~A300 & \new_[12474]_ ;
  assign \new_[12476]_  = \new_[12475]_  & \new_[12470]_ ;
  assign \new_[12479]_  = ~A167 & A170;
  assign \new_[12483]_  = A200 & ~A199;
  assign \new_[12484]_  = A166 & \new_[12483]_ ;
  assign \new_[12485]_  = \new_[12484]_  & \new_[12479]_ ;
  assign \new_[12489]_  = A267 & A265;
  assign \new_[12490]_  = A203 & \new_[12489]_ ;
  assign \new_[12494]_  = ~A301 & ~A299;
  assign \new_[12495]_  = ~A298 & \new_[12494]_ ;
  assign \new_[12496]_  = \new_[12495]_  & \new_[12490]_ ;
  assign \new_[12499]_  = ~A167 & A170;
  assign \new_[12503]_  = A200 & ~A199;
  assign \new_[12504]_  = A166 & \new_[12503]_ ;
  assign \new_[12505]_  = \new_[12504]_  & \new_[12499]_ ;
  assign \new_[12509]_  = A267 & A266;
  assign \new_[12510]_  = A203 & \new_[12509]_ ;
  assign \new_[12514]_  = ~A302 & ~A301;
  assign \new_[12515]_  = ~A300 & \new_[12514]_ ;
  assign \new_[12516]_  = \new_[12515]_  & \new_[12510]_ ;
  assign \new_[12519]_  = ~A167 & A170;
  assign \new_[12523]_  = A200 & ~A199;
  assign \new_[12524]_  = A166 & \new_[12523]_ ;
  assign \new_[12525]_  = \new_[12524]_  & \new_[12519]_ ;
  assign \new_[12529]_  = A267 & A266;
  assign \new_[12530]_  = A203 & \new_[12529]_ ;
  assign \new_[12534]_  = ~A301 & ~A299;
  assign \new_[12535]_  = ~A298 & \new_[12534]_ ;
  assign \new_[12536]_  = \new_[12535]_  & \new_[12530]_ ;
  assign \new_[12539]_  = ~A167 & A170;
  assign \new_[12543]_  = ~A200 & A199;
  assign \new_[12544]_  = A166 & \new_[12543]_ ;
  assign \new_[12545]_  = \new_[12544]_  & \new_[12539]_ ;
  assign \new_[12549]_  = A298 & A268;
  assign \new_[12550]_  = A203 & \new_[12549]_ ;
  assign \new_[12554]_  = ~A301 & ~A300;
  assign \new_[12555]_  = A299 & \new_[12554]_ ;
  assign \new_[12556]_  = \new_[12555]_  & \new_[12550]_ ;
  assign \new_[12559]_  = ~A167 & A170;
  assign \new_[12563]_  = ~A200 & A199;
  assign \new_[12564]_  = A166 & \new_[12563]_ ;
  assign \new_[12565]_  = \new_[12564]_  & \new_[12559]_ ;
  assign \new_[12569]_  = A267 & A265;
  assign \new_[12570]_  = A203 & \new_[12569]_ ;
  assign \new_[12574]_  = ~A302 & ~A301;
  assign \new_[12575]_  = ~A300 & \new_[12574]_ ;
  assign \new_[12576]_  = \new_[12575]_  & \new_[12570]_ ;
  assign \new_[12579]_  = ~A167 & A170;
  assign \new_[12583]_  = ~A200 & A199;
  assign \new_[12584]_  = A166 & \new_[12583]_ ;
  assign \new_[12585]_  = \new_[12584]_  & \new_[12579]_ ;
  assign \new_[12589]_  = A267 & A265;
  assign \new_[12590]_  = A203 & \new_[12589]_ ;
  assign \new_[12594]_  = ~A301 & ~A299;
  assign \new_[12595]_  = ~A298 & \new_[12594]_ ;
  assign \new_[12596]_  = \new_[12595]_  & \new_[12590]_ ;
  assign \new_[12599]_  = ~A167 & A170;
  assign \new_[12603]_  = ~A200 & A199;
  assign \new_[12604]_  = A166 & \new_[12603]_ ;
  assign \new_[12605]_  = \new_[12604]_  & \new_[12599]_ ;
  assign \new_[12609]_  = A267 & A266;
  assign \new_[12610]_  = A203 & \new_[12609]_ ;
  assign \new_[12614]_  = ~A302 & ~A301;
  assign \new_[12615]_  = ~A300 & \new_[12614]_ ;
  assign \new_[12616]_  = \new_[12615]_  & \new_[12610]_ ;
  assign \new_[12619]_  = ~A167 & A170;
  assign \new_[12623]_  = ~A200 & A199;
  assign \new_[12624]_  = A166 & \new_[12623]_ ;
  assign \new_[12625]_  = \new_[12624]_  & \new_[12619]_ ;
  assign \new_[12629]_  = A267 & A266;
  assign \new_[12630]_  = A203 & \new_[12629]_ ;
  assign \new_[12634]_  = ~A301 & ~A299;
  assign \new_[12635]_  = ~A298 & \new_[12634]_ ;
  assign \new_[12636]_  = \new_[12635]_  & \new_[12630]_ ;
  assign \new_[12639]_  = ~A167 & A170;
  assign \new_[12643]_  = ~A200 & ~A199;
  assign \new_[12644]_  = A166 & \new_[12643]_ ;
  assign \new_[12645]_  = \new_[12644]_  & \new_[12639]_ ;
  assign \new_[12649]_  = ~A268 & ~A267;
  assign \new_[12650]_  = ~A202 & \new_[12649]_ ;
  assign \new_[12654]_  = A300 & A299;
  assign \new_[12655]_  = ~A269 & \new_[12654]_ ;
  assign \new_[12656]_  = \new_[12655]_  & \new_[12650]_ ;
  assign \new_[12659]_  = ~A167 & A170;
  assign \new_[12663]_  = ~A200 & ~A199;
  assign \new_[12664]_  = A166 & \new_[12663]_ ;
  assign \new_[12665]_  = \new_[12664]_  & \new_[12659]_ ;
  assign \new_[12669]_  = ~A268 & ~A267;
  assign \new_[12670]_  = ~A202 & \new_[12669]_ ;
  assign \new_[12674]_  = A300 & A298;
  assign \new_[12675]_  = ~A269 & \new_[12674]_ ;
  assign \new_[12676]_  = \new_[12675]_  & \new_[12670]_ ;
  assign \new_[12679]_  = ~A167 & A170;
  assign \new_[12683]_  = ~A200 & ~A199;
  assign \new_[12684]_  = A166 & \new_[12683]_ ;
  assign \new_[12685]_  = \new_[12684]_  & \new_[12679]_ ;
  assign \new_[12689]_  = A266 & A265;
  assign \new_[12690]_  = ~A202 & \new_[12689]_ ;
  assign \new_[12694]_  = A301 & ~A268;
  assign \new_[12695]_  = ~A267 & \new_[12694]_ ;
  assign \new_[12696]_  = \new_[12695]_  & \new_[12690]_ ;
  assign \new_[12699]_  = ~A167 & A170;
  assign \new_[12703]_  = ~A200 & ~A199;
  assign \new_[12704]_  = A166 & \new_[12703]_ ;
  assign \new_[12705]_  = \new_[12704]_  & \new_[12699]_ ;
  assign \new_[12709]_  = ~A266 & ~A265;
  assign \new_[12710]_  = ~A202 & \new_[12709]_ ;
  assign \new_[12714]_  = A300 & A299;
  assign \new_[12715]_  = ~A268 & \new_[12714]_ ;
  assign \new_[12716]_  = \new_[12715]_  & \new_[12710]_ ;
  assign \new_[12719]_  = ~A167 & A170;
  assign \new_[12723]_  = ~A200 & ~A199;
  assign \new_[12724]_  = A166 & \new_[12723]_ ;
  assign \new_[12725]_  = \new_[12724]_  & \new_[12719]_ ;
  assign \new_[12729]_  = ~A266 & ~A265;
  assign \new_[12730]_  = ~A202 & \new_[12729]_ ;
  assign \new_[12734]_  = A300 & A298;
  assign \new_[12735]_  = ~A268 & \new_[12734]_ ;
  assign \new_[12736]_  = \new_[12735]_  & \new_[12730]_ ;
  assign \new_[12739]_  = ~A201 & A169;
  assign \new_[12743]_  = A265 & ~A203;
  assign \new_[12744]_  = ~A202 & \new_[12743]_ ;
  assign \new_[12745]_  = \new_[12744]_  & \new_[12739]_ ;
  assign \new_[12749]_  = ~A268 & ~A267;
  assign \new_[12750]_  = A266 & \new_[12749]_ ;
  assign \new_[12754]_  = A302 & ~A299;
  assign \new_[12755]_  = A298 & \new_[12754]_ ;
  assign \new_[12756]_  = \new_[12755]_  & \new_[12750]_ ;
  assign \new_[12759]_  = ~A201 & A169;
  assign \new_[12763]_  = A265 & ~A203;
  assign \new_[12764]_  = ~A202 & \new_[12763]_ ;
  assign \new_[12765]_  = \new_[12764]_  & \new_[12759]_ ;
  assign \new_[12769]_  = ~A268 & ~A267;
  assign \new_[12770]_  = A266 & \new_[12769]_ ;
  assign \new_[12774]_  = A302 & A299;
  assign \new_[12775]_  = ~A298 & \new_[12774]_ ;
  assign \new_[12776]_  = \new_[12775]_  & \new_[12770]_ ;
  assign \new_[12779]_  = A199 & A169;
  assign \new_[12783]_  = ~A202 & ~A201;
  assign \new_[12784]_  = A200 & \new_[12783]_ ;
  assign \new_[12785]_  = \new_[12784]_  & \new_[12779]_ ;
  assign \new_[12789]_  = ~A269 & ~A268;
  assign \new_[12790]_  = ~A267 & \new_[12789]_ ;
  assign \new_[12794]_  = A302 & ~A299;
  assign \new_[12795]_  = A298 & \new_[12794]_ ;
  assign \new_[12796]_  = \new_[12795]_  & \new_[12790]_ ;
  assign \new_[12799]_  = A199 & A169;
  assign \new_[12803]_  = ~A202 & ~A201;
  assign \new_[12804]_  = A200 & \new_[12803]_ ;
  assign \new_[12805]_  = \new_[12804]_  & \new_[12799]_ ;
  assign \new_[12809]_  = ~A269 & ~A268;
  assign \new_[12810]_  = ~A267 & \new_[12809]_ ;
  assign \new_[12814]_  = A302 & A299;
  assign \new_[12815]_  = ~A298 & \new_[12814]_ ;
  assign \new_[12816]_  = \new_[12815]_  & \new_[12810]_ ;
  assign \new_[12819]_  = A199 & A169;
  assign \new_[12823]_  = ~A202 & ~A201;
  assign \new_[12824]_  = A200 & \new_[12823]_ ;
  assign \new_[12825]_  = \new_[12824]_  & \new_[12819]_ ;
  assign \new_[12829]_  = ~A267 & A266;
  assign \new_[12830]_  = A265 & \new_[12829]_ ;
  assign \new_[12834]_  = A300 & A299;
  assign \new_[12835]_  = ~A268 & \new_[12834]_ ;
  assign \new_[12836]_  = \new_[12835]_  & \new_[12830]_ ;
  assign \new_[12839]_  = A199 & A169;
  assign \new_[12843]_  = ~A202 & ~A201;
  assign \new_[12844]_  = A200 & \new_[12843]_ ;
  assign \new_[12845]_  = \new_[12844]_  & \new_[12839]_ ;
  assign \new_[12849]_  = ~A267 & A266;
  assign \new_[12850]_  = A265 & \new_[12849]_ ;
  assign \new_[12854]_  = A300 & A298;
  assign \new_[12855]_  = ~A268 & \new_[12854]_ ;
  assign \new_[12856]_  = \new_[12855]_  & \new_[12850]_ ;
  assign \new_[12859]_  = A199 & A169;
  assign \new_[12863]_  = ~A202 & ~A201;
  assign \new_[12864]_  = A200 & \new_[12863]_ ;
  assign \new_[12865]_  = \new_[12864]_  & \new_[12859]_ ;
  assign \new_[12869]_  = ~A268 & ~A266;
  assign \new_[12870]_  = ~A265 & \new_[12869]_ ;
  assign \new_[12874]_  = A302 & ~A299;
  assign \new_[12875]_  = A298 & \new_[12874]_ ;
  assign \new_[12876]_  = \new_[12875]_  & \new_[12870]_ ;
  assign \new_[12879]_  = A199 & A169;
  assign \new_[12883]_  = ~A202 & ~A201;
  assign \new_[12884]_  = A200 & \new_[12883]_ ;
  assign \new_[12885]_  = \new_[12884]_  & \new_[12879]_ ;
  assign \new_[12889]_  = ~A268 & ~A266;
  assign \new_[12890]_  = ~A265 & \new_[12889]_ ;
  assign \new_[12894]_  = A302 & A299;
  assign \new_[12895]_  = ~A298 & \new_[12894]_ ;
  assign \new_[12896]_  = \new_[12895]_  & \new_[12890]_ ;
  assign \new_[12899]_  = ~A199 & A169;
  assign \new_[12903]_  = ~A265 & A203;
  assign \new_[12904]_  = A200 & \new_[12903]_ ;
  assign \new_[12905]_  = \new_[12904]_  & \new_[12899]_ ;
  assign \new_[12909]_  = A298 & A269;
  assign \new_[12910]_  = A266 & \new_[12909]_ ;
  assign \new_[12914]_  = ~A301 & ~A300;
  assign \new_[12915]_  = A299 & \new_[12914]_ ;
  assign \new_[12916]_  = \new_[12915]_  & \new_[12910]_ ;
  assign \new_[12919]_  = ~A199 & A169;
  assign \new_[12923]_  = A265 & A203;
  assign \new_[12924]_  = A200 & \new_[12923]_ ;
  assign \new_[12925]_  = \new_[12924]_  & \new_[12919]_ ;
  assign \new_[12929]_  = A298 & A269;
  assign \new_[12930]_  = ~A266 & \new_[12929]_ ;
  assign \new_[12934]_  = ~A301 & ~A300;
  assign \new_[12935]_  = A299 & \new_[12934]_ ;
  assign \new_[12936]_  = \new_[12935]_  & \new_[12930]_ ;
  assign \new_[12939]_  = A199 & A169;
  assign \new_[12943]_  = ~A265 & A203;
  assign \new_[12944]_  = ~A200 & \new_[12943]_ ;
  assign \new_[12945]_  = \new_[12944]_  & \new_[12939]_ ;
  assign \new_[12949]_  = A298 & A269;
  assign \new_[12950]_  = A266 & \new_[12949]_ ;
  assign \new_[12954]_  = ~A301 & ~A300;
  assign \new_[12955]_  = A299 & \new_[12954]_ ;
  assign \new_[12956]_  = \new_[12955]_  & \new_[12950]_ ;
  assign \new_[12959]_  = A199 & A169;
  assign \new_[12963]_  = A265 & A203;
  assign \new_[12964]_  = ~A200 & \new_[12963]_ ;
  assign \new_[12965]_  = \new_[12964]_  & \new_[12959]_ ;
  assign \new_[12969]_  = A298 & A269;
  assign \new_[12970]_  = ~A266 & \new_[12969]_ ;
  assign \new_[12974]_  = ~A301 & ~A300;
  assign \new_[12975]_  = A299 & \new_[12974]_ ;
  assign \new_[12976]_  = \new_[12975]_  & \new_[12970]_ ;
  assign \new_[12979]_  = ~A199 & A169;
  assign \new_[12983]_  = A265 & ~A202;
  assign \new_[12984]_  = ~A200 & \new_[12983]_ ;
  assign \new_[12985]_  = \new_[12984]_  & \new_[12979]_ ;
  assign \new_[12989]_  = ~A268 & ~A267;
  assign \new_[12990]_  = A266 & \new_[12989]_ ;
  assign \new_[12994]_  = A302 & ~A299;
  assign \new_[12995]_  = A298 & \new_[12994]_ ;
  assign \new_[12996]_  = \new_[12995]_  & \new_[12990]_ ;
  assign \new_[12999]_  = ~A199 & A169;
  assign \new_[13003]_  = A265 & ~A202;
  assign \new_[13004]_  = ~A200 & \new_[13003]_ ;
  assign \new_[13005]_  = \new_[13004]_  & \new_[12999]_ ;
  assign \new_[13009]_  = ~A268 & ~A267;
  assign \new_[13010]_  = A266 & \new_[13009]_ ;
  assign \new_[13014]_  = A302 & A299;
  assign \new_[13015]_  = ~A298 & \new_[13014]_ ;
  assign \new_[13016]_  = \new_[13015]_  & \new_[13010]_ ;
  assign \new_[13019]_  = ~A167 & ~A169;
  assign \new_[13023]_  = A265 & A202;
  assign \new_[13024]_  = ~A166 & \new_[13023]_ ;
  assign \new_[13025]_  = \new_[13024]_  & \new_[13019]_ ;
  assign \new_[13029]_  = ~A268 & ~A267;
  assign \new_[13030]_  = A266 & \new_[13029]_ ;
  assign \new_[13034]_  = A302 & ~A299;
  assign \new_[13035]_  = A298 & \new_[13034]_ ;
  assign \new_[13036]_  = \new_[13035]_  & \new_[13030]_ ;
  assign \new_[13039]_  = ~A167 & ~A169;
  assign \new_[13043]_  = A265 & A202;
  assign \new_[13044]_  = ~A166 & \new_[13043]_ ;
  assign \new_[13045]_  = \new_[13044]_  & \new_[13039]_ ;
  assign \new_[13049]_  = ~A268 & ~A267;
  assign \new_[13050]_  = A266 & \new_[13049]_ ;
  assign \new_[13054]_  = A302 & A299;
  assign \new_[13055]_  = ~A298 & \new_[13054]_ ;
  assign \new_[13056]_  = \new_[13055]_  & \new_[13050]_ ;
  assign \new_[13059]_  = ~A167 & ~A169;
  assign \new_[13063]_  = ~A202 & ~A201;
  assign \new_[13064]_  = ~A166 & \new_[13063]_ ;
  assign \new_[13065]_  = \new_[13064]_  & \new_[13059]_ ;
  assign \new_[13069]_  = A298 & A268;
  assign \new_[13070]_  = ~A203 & \new_[13069]_ ;
  assign \new_[13074]_  = ~A301 & ~A300;
  assign \new_[13075]_  = A299 & \new_[13074]_ ;
  assign \new_[13076]_  = \new_[13075]_  & \new_[13070]_ ;
  assign \new_[13079]_  = ~A167 & ~A169;
  assign \new_[13083]_  = ~A202 & ~A201;
  assign \new_[13084]_  = ~A166 & \new_[13083]_ ;
  assign \new_[13085]_  = \new_[13084]_  & \new_[13079]_ ;
  assign \new_[13089]_  = A267 & A265;
  assign \new_[13090]_  = ~A203 & \new_[13089]_ ;
  assign \new_[13094]_  = ~A302 & ~A301;
  assign \new_[13095]_  = ~A300 & \new_[13094]_ ;
  assign \new_[13096]_  = \new_[13095]_  & \new_[13090]_ ;
  assign \new_[13099]_  = ~A167 & ~A169;
  assign \new_[13103]_  = ~A202 & ~A201;
  assign \new_[13104]_  = ~A166 & \new_[13103]_ ;
  assign \new_[13105]_  = \new_[13104]_  & \new_[13099]_ ;
  assign \new_[13109]_  = A267 & A265;
  assign \new_[13110]_  = ~A203 & \new_[13109]_ ;
  assign \new_[13114]_  = ~A301 & ~A299;
  assign \new_[13115]_  = ~A298 & \new_[13114]_ ;
  assign \new_[13116]_  = \new_[13115]_  & \new_[13110]_ ;
  assign \new_[13119]_  = ~A167 & ~A169;
  assign \new_[13123]_  = ~A202 & ~A201;
  assign \new_[13124]_  = ~A166 & \new_[13123]_ ;
  assign \new_[13125]_  = \new_[13124]_  & \new_[13119]_ ;
  assign \new_[13129]_  = A267 & A266;
  assign \new_[13130]_  = ~A203 & \new_[13129]_ ;
  assign \new_[13134]_  = ~A302 & ~A301;
  assign \new_[13135]_  = ~A300 & \new_[13134]_ ;
  assign \new_[13136]_  = \new_[13135]_  & \new_[13130]_ ;
  assign \new_[13139]_  = ~A167 & ~A169;
  assign \new_[13143]_  = ~A202 & ~A201;
  assign \new_[13144]_  = ~A166 & \new_[13143]_ ;
  assign \new_[13145]_  = \new_[13144]_  & \new_[13139]_ ;
  assign \new_[13149]_  = A267 & A266;
  assign \new_[13150]_  = ~A203 & \new_[13149]_ ;
  assign \new_[13154]_  = ~A301 & ~A299;
  assign \new_[13155]_  = ~A298 & \new_[13154]_ ;
  assign \new_[13156]_  = \new_[13155]_  & \new_[13150]_ ;
  assign \new_[13159]_  = ~A167 & ~A169;
  assign \new_[13163]_  = A201 & A199;
  assign \new_[13164]_  = ~A166 & \new_[13163]_ ;
  assign \new_[13165]_  = \new_[13164]_  & \new_[13159]_ ;
  assign \new_[13169]_  = ~A269 & ~A268;
  assign \new_[13170]_  = ~A267 & \new_[13169]_ ;
  assign \new_[13174]_  = A302 & ~A299;
  assign \new_[13175]_  = A298 & \new_[13174]_ ;
  assign \new_[13176]_  = \new_[13175]_  & \new_[13170]_ ;
  assign \new_[13179]_  = ~A167 & ~A169;
  assign \new_[13183]_  = A201 & A199;
  assign \new_[13184]_  = ~A166 & \new_[13183]_ ;
  assign \new_[13185]_  = \new_[13184]_  & \new_[13179]_ ;
  assign \new_[13189]_  = ~A269 & ~A268;
  assign \new_[13190]_  = ~A267 & \new_[13189]_ ;
  assign \new_[13194]_  = A302 & A299;
  assign \new_[13195]_  = ~A298 & \new_[13194]_ ;
  assign \new_[13196]_  = \new_[13195]_  & \new_[13190]_ ;
  assign \new_[13199]_  = ~A167 & ~A169;
  assign \new_[13203]_  = A201 & A199;
  assign \new_[13204]_  = ~A166 & \new_[13203]_ ;
  assign \new_[13205]_  = \new_[13204]_  & \new_[13199]_ ;
  assign \new_[13209]_  = ~A267 & A266;
  assign \new_[13210]_  = A265 & \new_[13209]_ ;
  assign \new_[13214]_  = A300 & A299;
  assign \new_[13215]_  = ~A268 & \new_[13214]_ ;
  assign \new_[13216]_  = \new_[13215]_  & \new_[13210]_ ;
  assign \new_[13219]_  = ~A167 & ~A169;
  assign \new_[13223]_  = A201 & A199;
  assign \new_[13224]_  = ~A166 & \new_[13223]_ ;
  assign \new_[13225]_  = \new_[13224]_  & \new_[13219]_ ;
  assign \new_[13229]_  = ~A267 & A266;
  assign \new_[13230]_  = A265 & \new_[13229]_ ;
  assign \new_[13234]_  = A300 & A298;
  assign \new_[13235]_  = ~A268 & \new_[13234]_ ;
  assign \new_[13236]_  = \new_[13235]_  & \new_[13230]_ ;
  assign \new_[13239]_  = ~A167 & ~A169;
  assign \new_[13243]_  = A201 & A199;
  assign \new_[13244]_  = ~A166 & \new_[13243]_ ;
  assign \new_[13245]_  = \new_[13244]_  & \new_[13239]_ ;
  assign \new_[13249]_  = ~A268 & ~A266;
  assign \new_[13250]_  = ~A265 & \new_[13249]_ ;
  assign \new_[13254]_  = A302 & ~A299;
  assign \new_[13255]_  = A298 & \new_[13254]_ ;
  assign \new_[13256]_  = \new_[13255]_  & \new_[13250]_ ;
  assign \new_[13259]_  = ~A167 & ~A169;
  assign \new_[13263]_  = A201 & A199;
  assign \new_[13264]_  = ~A166 & \new_[13263]_ ;
  assign \new_[13265]_  = \new_[13264]_  & \new_[13259]_ ;
  assign \new_[13269]_  = ~A268 & ~A266;
  assign \new_[13270]_  = ~A265 & \new_[13269]_ ;
  assign \new_[13274]_  = A302 & A299;
  assign \new_[13275]_  = ~A298 & \new_[13274]_ ;
  assign \new_[13276]_  = \new_[13275]_  & \new_[13270]_ ;
  assign \new_[13279]_  = ~A167 & ~A169;
  assign \new_[13283]_  = A201 & A200;
  assign \new_[13284]_  = ~A166 & \new_[13283]_ ;
  assign \new_[13285]_  = \new_[13284]_  & \new_[13279]_ ;
  assign \new_[13289]_  = ~A269 & ~A268;
  assign \new_[13290]_  = ~A267 & \new_[13289]_ ;
  assign \new_[13294]_  = A302 & ~A299;
  assign \new_[13295]_  = A298 & \new_[13294]_ ;
  assign \new_[13296]_  = \new_[13295]_  & \new_[13290]_ ;
  assign \new_[13299]_  = ~A167 & ~A169;
  assign \new_[13303]_  = A201 & A200;
  assign \new_[13304]_  = ~A166 & \new_[13303]_ ;
  assign \new_[13305]_  = \new_[13304]_  & \new_[13299]_ ;
  assign \new_[13309]_  = ~A269 & ~A268;
  assign \new_[13310]_  = ~A267 & \new_[13309]_ ;
  assign \new_[13314]_  = A302 & A299;
  assign \new_[13315]_  = ~A298 & \new_[13314]_ ;
  assign \new_[13316]_  = \new_[13315]_  & \new_[13310]_ ;
  assign \new_[13319]_  = ~A167 & ~A169;
  assign \new_[13323]_  = A201 & A200;
  assign \new_[13324]_  = ~A166 & \new_[13323]_ ;
  assign \new_[13325]_  = \new_[13324]_  & \new_[13319]_ ;
  assign \new_[13329]_  = ~A267 & A266;
  assign \new_[13330]_  = A265 & \new_[13329]_ ;
  assign \new_[13334]_  = A300 & A299;
  assign \new_[13335]_  = ~A268 & \new_[13334]_ ;
  assign \new_[13336]_  = \new_[13335]_  & \new_[13330]_ ;
  assign \new_[13339]_  = ~A167 & ~A169;
  assign \new_[13343]_  = A201 & A200;
  assign \new_[13344]_  = ~A166 & \new_[13343]_ ;
  assign \new_[13345]_  = \new_[13344]_  & \new_[13339]_ ;
  assign \new_[13349]_  = ~A267 & A266;
  assign \new_[13350]_  = A265 & \new_[13349]_ ;
  assign \new_[13354]_  = A300 & A298;
  assign \new_[13355]_  = ~A268 & \new_[13354]_ ;
  assign \new_[13356]_  = \new_[13355]_  & \new_[13350]_ ;
  assign \new_[13359]_  = ~A167 & ~A169;
  assign \new_[13363]_  = A201 & A200;
  assign \new_[13364]_  = ~A166 & \new_[13363]_ ;
  assign \new_[13365]_  = \new_[13364]_  & \new_[13359]_ ;
  assign \new_[13369]_  = ~A268 & ~A266;
  assign \new_[13370]_  = ~A265 & \new_[13369]_ ;
  assign \new_[13374]_  = A302 & ~A299;
  assign \new_[13375]_  = A298 & \new_[13374]_ ;
  assign \new_[13376]_  = \new_[13375]_  & \new_[13370]_ ;
  assign \new_[13379]_  = ~A167 & ~A169;
  assign \new_[13383]_  = A201 & A200;
  assign \new_[13384]_  = ~A166 & \new_[13383]_ ;
  assign \new_[13385]_  = \new_[13384]_  & \new_[13379]_ ;
  assign \new_[13389]_  = ~A268 & ~A266;
  assign \new_[13390]_  = ~A265 & \new_[13389]_ ;
  assign \new_[13394]_  = A302 & A299;
  assign \new_[13395]_  = ~A298 & \new_[13394]_ ;
  assign \new_[13396]_  = \new_[13395]_  & \new_[13390]_ ;
  assign \new_[13399]_  = ~A167 & ~A169;
  assign \new_[13403]_  = A200 & A199;
  assign \new_[13404]_  = ~A166 & \new_[13403]_ ;
  assign \new_[13405]_  = \new_[13404]_  & \new_[13399]_ ;
  assign \new_[13409]_  = A268 & ~A202;
  assign \new_[13410]_  = ~A201 & \new_[13409]_ ;
  assign \new_[13414]_  = ~A302 & ~A301;
  assign \new_[13415]_  = ~A300 & \new_[13414]_ ;
  assign \new_[13416]_  = \new_[13415]_  & \new_[13410]_ ;
  assign \new_[13419]_  = ~A167 & ~A169;
  assign \new_[13423]_  = A200 & A199;
  assign \new_[13424]_  = ~A166 & \new_[13423]_ ;
  assign \new_[13425]_  = \new_[13424]_  & \new_[13419]_ ;
  assign \new_[13429]_  = A268 & ~A202;
  assign \new_[13430]_  = ~A201 & \new_[13429]_ ;
  assign \new_[13434]_  = ~A301 & ~A299;
  assign \new_[13435]_  = ~A298 & \new_[13434]_ ;
  assign \new_[13436]_  = \new_[13435]_  & \new_[13430]_ ;
  assign \new_[13439]_  = ~A167 & ~A169;
  assign \new_[13443]_  = A200 & ~A199;
  assign \new_[13444]_  = ~A166 & \new_[13443]_ ;
  assign \new_[13445]_  = \new_[13444]_  & \new_[13439]_ ;
  assign \new_[13449]_  = ~A268 & ~A267;
  assign \new_[13450]_  = A203 & \new_[13449]_ ;
  assign \new_[13454]_  = A300 & A299;
  assign \new_[13455]_  = ~A269 & \new_[13454]_ ;
  assign \new_[13456]_  = \new_[13455]_  & \new_[13450]_ ;
  assign \new_[13459]_  = ~A167 & ~A169;
  assign \new_[13463]_  = A200 & ~A199;
  assign \new_[13464]_  = ~A166 & \new_[13463]_ ;
  assign \new_[13465]_  = \new_[13464]_  & \new_[13459]_ ;
  assign \new_[13469]_  = ~A268 & ~A267;
  assign \new_[13470]_  = A203 & \new_[13469]_ ;
  assign \new_[13474]_  = A300 & A298;
  assign \new_[13475]_  = ~A269 & \new_[13474]_ ;
  assign \new_[13476]_  = \new_[13475]_  & \new_[13470]_ ;
  assign \new_[13479]_  = ~A167 & ~A169;
  assign \new_[13483]_  = A200 & ~A199;
  assign \new_[13484]_  = ~A166 & \new_[13483]_ ;
  assign \new_[13485]_  = \new_[13484]_  & \new_[13479]_ ;
  assign \new_[13489]_  = A266 & A265;
  assign \new_[13490]_  = A203 & \new_[13489]_ ;
  assign \new_[13494]_  = A301 & ~A268;
  assign \new_[13495]_  = ~A267 & \new_[13494]_ ;
  assign \new_[13496]_  = \new_[13495]_  & \new_[13490]_ ;
  assign \new_[13499]_  = ~A167 & ~A169;
  assign \new_[13503]_  = A200 & ~A199;
  assign \new_[13504]_  = ~A166 & \new_[13503]_ ;
  assign \new_[13505]_  = \new_[13504]_  & \new_[13499]_ ;
  assign \new_[13509]_  = ~A266 & ~A265;
  assign \new_[13510]_  = A203 & \new_[13509]_ ;
  assign \new_[13514]_  = A300 & A299;
  assign \new_[13515]_  = ~A268 & \new_[13514]_ ;
  assign \new_[13516]_  = \new_[13515]_  & \new_[13510]_ ;
  assign \new_[13519]_  = ~A167 & ~A169;
  assign \new_[13523]_  = A200 & ~A199;
  assign \new_[13524]_  = ~A166 & \new_[13523]_ ;
  assign \new_[13525]_  = \new_[13524]_  & \new_[13519]_ ;
  assign \new_[13529]_  = ~A266 & ~A265;
  assign \new_[13530]_  = A203 & \new_[13529]_ ;
  assign \new_[13534]_  = A300 & A298;
  assign \new_[13535]_  = ~A268 & \new_[13534]_ ;
  assign \new_[13536]_  = \new_[13535]_  & \new_[13530]_ ;
  assign \new_[13539]_  = ~A167 & ~A169;
  assign \new_[13543]_  = ~A200 & A199;
  assign \new_[13544]_  = ~A166 & \new_[13543]_ ;
  assign \new_[13545]_  = \new_[13544]_  & \new_[13539]_ ;
  assign \new_[13549]_  = ~A268 & ~A267;
  assign \new_[13550]_  = A203 & \new_[13549]_ ;
  assign \new_[13554]_  = A300 & A299;
  assign \new_[13555]_  = ~A269 & \new_[13554]_ ;
  assign \new_[13556]_  = \new_[13555]_  & \new_[13550]_ ;
  assign \new_[13559]_  = ~A167 & ~A169;
  assign \new_[13563]_  = ~A200 & A199;
  assign \new_[13564]_  = ~A166 & \new_[13563]_ ;
  assign \new_[13565]_  = \new_[13564]_  & \new_[13559]_ ;
  assign \new_[13569]_  = ~A268 & ~A267;
  assign \new_[13570]_  = A203 & \new_[13569]_ ;
  assign \new_[13574]_  = A300 & A298;
  assign \new_[13575]_  = ~A269 & \new_[13574]_ ;
  assign \new_[13576]_  = \new_[13575]_  & \new_[13570]_ ;
  assign \new_[13579]_  = ~A167 & ~A169;
  assign \new_[13583]_  = ~A200 & A199;
  assign \new_[13584]_  = ~A166 & \new_[13583]_ ;
  assign \new_[13585]_  = \new_[13584]_  & \new_[13579]_ ;
  assign \new_[13589]_  = A266 & A265;
  assign \new_[13590]_  = A203 & \new_[13589]_ ;
  assign \new_[13594]_  = A301 & ~A268;
  assign \new_[13595]_  = ~A267 & \new_[13594]_ ;
  assign \new_[13596]_  = \new_[13595]_  & \new_[13590]_ ;
  assign \new_[13599]_  = ~A167 & ~A169;
  assign \new_[13603]_  = ~A200 & A199;
  assign \new_[13604]_  = ~A166 & \new_[13603]_ ;
  assign \new_[13605]_  = \new_[13604]_  & \new_[13599]_ ;
  assign \new_[13609]_  = ~A266 & ~A265;
  assign \new_[13610]_  = A203 & \new_[13609]_ ;
  assign \new_[13614]_  = A300 & A299;
  assign \new_[13615]_  = ~A268 & \new_[13614]_ ;
  assign \new_[13616]_  = \new_[13615]_  & \new_[13610]_ ;
  assign \new_[13619]_  = ~A167 & ~A169;
  assign \new_[13623]_  = ~A200 & A199;
  assign \new_[13624]_  = ~A166 & \new_[13623]_ ;
  assign \new_[13625]_  = \new_[13624]_  & \new_[13619]_ ;
  assign \new_[13629]_  = ~A266 & ~A265;
  assign \new_[13630]_  = A203 & \new_[13629]_ ;
  assign \new_[13634]_  = A300 & A298;
  assign \new_[13635]_  = ~A268 & \new_[13634]_ ;
  assign \new_[13636]_  = \new_[13635]_  & \new_[13630]_ ;
  assign \new_[13639]_  = ~A167 & ~A169;
  assign \new_[13643]_  = ~A200 & ~A199;
  assign \new_[13644]_  = ~A166 & \new_[13643]_ ;
  assign \new_[13645]_  = \new_[13644]_  & \new_[13639]_ ;
  assign \new_[13649]_  = A298 & A268;
  assign \new_[13650]_  = ~A202 & \new_[13649]_ ;
  assign \new_[13654]_  = ~A301 & ~A300;
  assign \new_[13655]_  = A299 & \new_[13654]_ ;
  assign \new_[13656]_  = \new_[13655]_  & \new_[13650]_ ;
  assign \new_[13659]_  = ~A167 & ~A169;
  assign \new_[13663]_  = ~A200 & ~A199;
  assign \new_[13664]_  = ~A166 & \new_[13663]_ ;
  assign \new_[13665]_  = \new_[13664]_  & \new_[13659]_ ;
  assign \new_[13669]_  = A267 & A265;
  assign \new_[13670]_  = ~A202 & \new_[13669]_ ;
  assign \new_[13674]_  = ~A302 & ~A301;
  assign \new_[13675]_  = ~A300 & \new_[13674]_ ;
  assign \new_[13676]_  = \new_[13675]_  & \new_[13670]_ ;
  assign \new_[13679]_  = ~A167 & ~A169;
  assign \new_[13683]_  = ~A200 & ~A199;
  assign \new_[13684]_  = ~A166 & \new_[13683]_ ;
  assign \new_[13685]_  = \new_[13684]_  & \new_[13679]_ ;
  assign \new_[13689]_  = A267 & A265;
  assign \new_[13690]_  = ~A202 & \new_[13689]_ ;
  assign \new_[13694]_  = ~A301 & ~A299;
  assign \new_[13695]_  = ~A298 & \new_[13694]_ ;
  assign \new_[13696]_  = \new_[13695]_  & \new_[13690]_ ;
  assign \new_[13699]_  = ~A167 & ~A169;
  assign \new_[13703]_  = ~A200 & ~A199;
  assign \new_[13704]_  = ~A166 & \new_[13703]_ ;
  assign \new_[13705]_  = \new_[13704]_  & \new_[13699]_ ;
  assign \new_[13709]_  = A267 & A266;
  assign \new_[13710]_  = ~A202 & \new_[13709]_ ;
  assign \new_[13714]_  = ~A302 & ~A301;
  assign \new_[13715]_  = ~A300 & \new_[13714]_ ;
  assign \new_[13716]_  = \new_[13715]_  & \new_[13710]_ ;
  assign \new_[13719]_  = ~A167 & ~A169;
  assign \new_[13723]_  = ~A200 & ~A199;
  assign \new_[13724]_  = ~A166 & \new_[13723]_ ;
  assign \new_[13725]_  = \new_[13724]_  & \new_[13719]_ ;
  assign \new_[13729]_  = A267 & A266;
  assign \new_[13730]_  = ~A202 & \new_[13729]_ ;
  assign \new_[13734]_  = ~A301 & ~A299;
  assign \new_[13735]_  = ~A298 & \new_[13734]_ ;
  assign \new_[13736]_  = \new_[13735]_  & \new_[13730]_ ;
  assign \new_[13739]_  = ~A168 & ~A169;
  assign \new_[13743]_  = A202 & A166;
  assign \new_[13744]_  = A167 & \new_[13743]_ ;
  assign \new_[13745]_  = \new_[13744]_  & \new_[13739]_ ;
  assign \new_[13749]_  = ~A269 & ~A268;
  assign \new_[13750]_  = ~A267 & \new_[13749]_ ;
  assign \new_[13754]_  = A302 & ~A299;
  assign \new_[13755]_  = A298 & \new_[13754]_ ;
  assign \new_[13756]_  = \new_[13755]_  & \new_[13750]_ ;
  assign \new_[13759]_  = ~A168 & ~A169;
  assign \new_[13763]_  = A202 & A166;
  assign \new_[13764]_  = A167 & \new_[13763]_ ;
  assign \new_[13765]_  = \new_[13764]_  & \new_[13759]_ ;
  assign \new_[13769]_  = ~A269 & ~A268;
  assign \new_[13770]_  = ~A267 & \new_[13769]_ ;
  assign \new_[13774]_  = A302 & A299;
  assign \new_[13775]_  = ~A298 & \new_[13774]_ ;
  assign \new_[13776]_  = \new_[13775]_  & \new_[13770]_ ;
  assign \new_[13779]_  = ~A168 & ~A169;
  assign \new_[13783]_  = A202 & A166;
  assign \new_[13784]_  = A167 & \new_[13783]_ ;
  assign \new_[13785]_  = \new_[13784]_  & \new_[13779]_ ;
  assign \new_[13789]_  = ~A267 & A266;
  assign \new_[13790]_  = A265 & \new_[13789]_ ;
  assign \new_[13794]_  = A300 & A299;
  assign \new_[13795]_  = ~A268 & \new_[13794]_ ;
  assign \new_[13796]_  = \new_[13795]_  & \new_[13790]_ ;
  assign \new_[13799]_  = ~A168 & ~A169;
  assign \new_[13803]_  = A202 & A166;
  assign \new_[13804]_  = A167 & \new_[13803]_ ;
  assign \new_[13805]_  = \new_[13804]_  & \new_[13799]_ ;
  assign \new_[13809]_  = ~A267 & A266;
  assign \new_[13810]_  = A265 & \new_[13809]_ ;
  assign \new_[13814]_  = A300 & A298;
  assign \new_[13815]_  = ~A268 & \new_[13814]_ ;
  assign \new_[13816]_  = \new_[13815]_  & \new_[13810]_ ;
  assign \new_[13819]_  = ~A168 & ~A169;
  assign \new_[13823]_  = A202 & A166;
  assign \new_[13824]_  = A167 & \new_[13823]_ ;
  assign \new_[13825]_  = \new_[13824]_  & \new_[13819]_ ;
  assign \new_[13829]_  = ~A268 & ~A266;
  assign \new_[13830]_  = ~A265 & \new_[13829]_ ;
  assign \new_[13834]_  = A302 & ~A299;
  assign \new_[13835]_  = A298 & \new_[13834]_ ;
  assign \new_[13836]_  = \new_[13835]_  & \new_[13830]_ ;
  assign \new_[13839]_  = ~A168 & ~A169;
  assign \new_[13843]_  = A202 & A166;
  assign \new_[13844]_  = A167 & \new_[13843]_ ;
  assign \new_[13845]_  = \new_[13844]_  & \new_[13839]_ ;
  assign \new_[13849]_  = ~A268 & ~A266;
  assign \new_[13850]_  = ~A265 & \new_[13849]_ ;
  assign \new_[13854]_  = A302 & A299;
  assign \new_[13855]_  = ~A298 & \new_[13854]_ ;
  assign \new_[13856]_  = \new_[13855]_  & \new_[13850]_ ;
  assign \new_[13859]_  = ~A168 & ~A169;
  assign \new_[13863]_  = ~A201 & A166;
  assign \new_[13864]_  = A167 & \new_[13863]_ ;
  assign \new_[13865]_  = \new_[13864]_  & \new_[13859]_ ;
  assign \new_[13869]_  = A268 & ~A203;
  assign \new_[13870]_  = ~A202 & \new_[13869]_ ;
  assign \new_[13874]_  = ~A302 & ~A301;
  assign \new_[13875]_  = ~A300 & \new_[13874]_ ;
  assign \new_[13876]_  = \new_[13875]_  & \new_[13870]_ ;
  assign \new_[13879]_  = ~A168 & ~A169;
  assign \new_[13883]_  = ~A201 & A166;
  assign \new_[13884]_  = A167 & \new_[13883]_ ;
  assign \new_[13885]_  = \new_[13884]_  & \new_[13879]_ ;
  assign \new_[13889]_  = A268 & ~A203;
  assign \new_[13890]_  = ~A202 & \new_[13889]_ ;
  assign \new_[13894]_  = ~A301 & ~A299;
  assign \new_[13895]_  = ~A298 & \new_[13894]_ ;
  assign \new_[13896]_  = \new_[13895]_  & \new_[13890]_ ;
  assign \new_[13899]_  = ~A168 & ~A169;
  assign \new_[13903]_  = A199 & A166;
  assign \new_[13904]_  = A167 & \new_[13903]_ ;
  assign \new_[13905]_  = \new_[13904]_  & \new_[13899]_ ;
  assign \new_[13909]_  = ~A268 & ~A267;
  assign \new_[13910]_  = A201 & \new_[13909]_ ;
  assign \new_[13914]_  = A300 & A299;
  assign \new_[13915]_  = ~A269 & \new_[13914]_ ;
  assign \new_[13916]_  = \new_[13915]_  & \new_[13910]_ ;
  assign \new_[13919]_  = ~A168 & ~A169;
  assign \new_[13923]_  = A199 & A166;
  assign \new_[13924]_  = A167 & \new_[13923]_ ;
  assign \new_[13925]_  = \new_[13924]_  & \new_[13919]_ ;
  assign \new_[13929]_  = ~A268 & ~A267;
  assign \new_[13930]_  = A201 & \new_[13929]_ ;
  assign \new_[13934]_  = A300 & A298;
  assign \new_[13935]_  = ~A269 & \new_[13934]_ ;
  assign \new_[13936]_  = \new_[13935]_  & \new_[13930]_ ;
  assign \new_[13939]_  = ~A168 & ~A169;
  assign \new_[13943]_  = A199 & A166;
  assign \new_[13944]_  = A167 & \new_[13943]_ ;
  assign \new_[13945]_  = \new_[13944]_  & \new_[13939]_ ;
  assign \new_[13949]_  = A266 & A265;
  assign \new_[13950]_  = A201 & \new_[13949]_ ;
  assign \new_[13954]_  = A301 & ~A268;
  assign \new_[13955]_  = ~A267 & \new_[13954]_ ;
  assign \new_[13956]_  = \new_[13955]_  & \new_[13950]_ ;
  assign \new_[13959]_  = ~A168 & ~A169;
  assign \new_[13963]_  = A199 & A166;
  assign \new_[13964]_  = A167 & \new_[13963]_ ;
  assign \new_[13965]_  = \new_[13964]_  & \new_[13959]_ ;
  assign \new_[13969]_  = ~A266 & ~A265;
  assign \new_[13970]_  = A201 & \new_[13969]_ ;
  assign \new_[13974]_  = A300 & A299;
  assign \new_[13975]_  = ~A268 & \new_[13974]_ ;
  assign \new_[13976]_  = \new_[13975]_  & \new_[13970]_ ;
  assign \new_[13979]_  = ~A168 & ~A169;
  assign \new_[13983]_  = A199 & A166;
  assign \new_[13984]_  = A167 & \new_[13983]_ ;
  assign \new_[13985]_  = \new_[13984]_  & \new_[13979]_ ;
  assign \new_[13989]_  = ~A266 & ~A265;
  assign \new_[13990]_  = A201 & \new_[13989]_ ;
  assign \new_[13994]_  = A300 & A298;
  assign \new_[13995]_  = ~A268 & \new_[13994]_ ;
  assign \new_[13996]_  = \new_[13995]_  & \new_[13990]_ ;
  assign \new_[13999]_  = ~A168 & ~A169;
  assign \new_[14003]_  = A200 & A166;
  assign \new_[14004]_  = A167 & \new_[14003]_ ;
  assign \new_[14005]_  = \new_[14004]_  & \new_[13999]_ ;
  assign \new_[14009]_  = ~A268 & ~A267;
  assign \new_[14010]_  = A201 & \new_[14009]_ ;
  assign \new_[14014]_  = A300 & A299;
  assign \new_[14015]_  = ~A269 & \new_[14014]_ ;
  assign \new_[14016]_  = \new_[14015]_  & \new_[14010]_ ;
  assign \new_[14019]_  = ~A168 & ~A169;
  assign \new_[14023]_  = A200 & A166;
  assign \new_[14024]_  = A167 & \new_[14023]_ ;
  assign \new_[14025]_  = \new_[14024]_  & \new_[14019]_ ;
  assign \new_[14029]_  = ~A268 & ~A267;
  assign \new_[14030]_  = A201 & \new_[14029]_ ;
  assign \new_[14034]_  = A300 & A298;
  assign \new_[14035]_  = ~A269 & \new_[14034]_ ;
  assign \new_[14036]_  = \new_[14035]_  & \new_[14030]_ ;
  assign \new_[14039]_  = ~A168 & ~A169;
  assign \new_[14043]_  = A200 & A166;
  assign \new_[14044]_  = A167 & \new_[14043]_ ;
  assign \new_[14045]_  = \new_[14044]_  & \new_[14039]_ ;
  assign \new_[14049]_  = A266 & A265;
  assign \new_[14050]_  = A201 & \new_[14049]_ ;
  assign \new_[14054]_  = A301 & ~A268;
  assign \new_[14055]_  = ~A267 & \new_[14054]_ ;
  assign \new_[14056]_  = \new_[14055]_  & \new_[14050]_ ;
  assign \new_[14059]_  = ~A168 & ~A169;
  assign \new_[14063]_  = A200 & A166;
  assign \new_[14064]_  = A167 & \new_[14063]_ ;
  assign \new_[14065]_  = \new_[14064]_  & \new_[14059]_ ;
  assign \new_[14069]_  = ~A266 & ~A265;
  assign \new_[14070]_  = A201 & \new_[14069]_ ;
  assign \new_[14074]_  = A300 & A299;
  assign \new_[14075]_  = ~A268 & \new_[14074]_ ;
  assign \new_[14076]_  = \new_[14075]_  & \new_[14070]_ ;
  assign \new_[14079]_  = ~A168 & ~A169;
  assign \new_[14083]_  = A200 & A166;
  assign \new_[14084]_  = A167 & \new_[14083]_ ;
  assign \new_[14085]_  = \new_[14084]_  & \new_[14079]_ ;
  assign \new_[14089]_  = ~A266 & ~A265;
  assign \new_[14090]_  = A201 & \new_[14089]_ ;
  assign \new_[14094]_  = A300 & A298;
  assign \new_[14095]_  = ~A268 & \new_[14094]_ ;
  assign \new_[14096]_  = \new_[14095]_  & \new_[14090]_ ;
  assign \new_[14099]_  = ~A168 & ~A169;
  assign \new_[14103]_  = ~A199 & A166;
  assign \new_[14104]_  = A167 & \new_[14103]_ ;
  assign \new_[14105]_  = \new_[14104]_  & \new_[14099]_ ;
  assign \new_[14109]_  = ~A267 & A203;
  assign \new_[14110]_  = A200 & \new_[14109]_ ;
  assign \new_[14114]_  = A301 & ~A269;
  assign \new_[14115]_  = ~A268 & \new_[14114]_ ;
  assign \new_[14116]_  = \new_[14115]_  & \new_[14110]_ ;
  assign \new_[14119]_  = ~A168 & ~A169;
  assign \new_[14123]_  = ~A199 & A166;
  assign \new_[14124]_  = A167 & \new_[14123]_ ;
  assign \new_[14125]_  = \new_[14124]_  & \new_[14119]_ ;
  assign \new_[14129]_  = ~A265 & A203;
  assign \new_[14130]_  = A200 & \new_[14129]_ ;
  assign \new_[14134]_  = A301 & ~A268;
  assign \new_[14135]_  = ~A266 & \new_[14134]_ ;
  assign \new_[14136]_  = \new_[14135]_  & \new_[14130]_ ;
  assign \new_[14139]_  = ~A168 & ~A169;
  assign \new_[14143]_  = A199 & A166;
  assign \new_[14144]_  = A167 & \new_[14143]_ ;
  assign \new_[14145]_  = \new_[14144]_  & \new_[14139]_ ;
  assign \new_[14149]_  = ~A267 & A203;
  assign \new_[14150]_  = ~A200 & \new_[14149]_ ;
  assign \new_[14154]_  = A301 & ~A269;
  assign \new_[14155]_  = ~A268 & \new_[14154]_ ;
  assign \new_[14156]_  = \new_[14155]_  & \new_[14150]_ ;
  assign \new_[14159]_  = ~A168 & ~A169;
  assign \new_[14163]_  = A199 & A166;
  assign \new_[14164]_  = A167 & \new_[14163]_ ;
  assign \new_[14165]_  = \new_[14164]_  & \new_[14159]_ ;
  assign \new_[14169]_  = ~A265 & A203;
  assign \new_[14170]_  = ~A200 & \new_[14169]_ ;
  assign \new_[14174]_  = A301 & ~A268;
  assign \new_[14175]_  = ~A266 & \new_[14174]_ ;
  assign \new_[14176]_  = \new_[14175]_  & \new_[14170]_ ;
  assign \new_[14179]_  = ~A168 & ~A169;
  assign \new_[14183]_  = ~A199 & A166;
  assign \new_[14184]_  = A167 & \new_[14183]_ ;
  assign \new_[14185]_  = \new_[14184]_  & \new_[14179]_ ;
  assign \new_[14189]_  = A268 & ~A202;
  assign \new_[14190]_  = ~A200 & \new_[14189]_ ;
  assign \new_[14194]_  = ~A302 & ~A301;
  assign \new_[14195]_  = ~A300 & \new_[14194]_ ;
  assign \new_[14196]_  = \new_[14195]_  & \new_[14190]_ ;
  assign \new_[14199]_  = ~A168 & ~A169;
  assign \new_[14203]_  = ~A199 & A166;
  assign \new_[14204]_  = A167 & \new_[14203]_ ;
  assign \new_[14205]_  = \new_[14204]_  & \new_[14199]_ ;
  assign \new_[14209]_  = A268 & ~A202;
  assign \new_[14210]_  = ~A200 & \new_[14209]_ ;
  assign \new_[14214]_  = ~A301 & ~A299;
  assign \new_[14215]_  = ~A298 & \new_[14214]_ ;
  assign \new_[14216]_  = \new_[14215]_  & \new_[14210]_ ;
  assign \new_[14219]_  = ~A169 & ~A170;
  assign \new_[14223]_  = A265 & A202;
  assign \new_[14224]_  = ~A168 & \new_[14223]_ ;
  assign \new_[14225]_  = \new_[14224]_  & \new_[14219]_ ;
  assign \new_[14229]_  = ~A268 & ~A267;
  assign \new_[14230]_  = A266 & \new_[14229]_ ;
  assign \new_[14234]_  = A302 & ~A299;
  assign \new_[14235]_  = A298 & \new_[14234]_ ;
  assign \new_[14236]_  = \new_[14235]_  & \new_[14230]_ ;
  assign \new_[14239]_  = ~A169 & ~A170;
  assign \new_[14243]_  = A265 & A202;
  assign \new_[14244]_  = ~A168 & \new_[14243]_ ;
  assign \new_[14245]_  = \new_[14244]_  & \new_[14239]_ ;
  assign \new_[14249]_  = ~A268 & ~A267;
  assign \new_[14250]_  = A266 & \new_[14249]_ ;
  assign \new_[14254]_  = A302 & A299;
  assign \new_[14255]_  = ~A298 & \new_[14254]_ ;
  assign \new_[14256]_  = \new_[14255]_  & \new_[14250]_ ;
  assign \new_[14259]_  = ~A169 & ~A170;
  assign \new_[14263]_  = ~A202 & ~A201;
  assign \new_[14264]_  = ~A168 & \new_[14263]_ ;
  assign \new_[14265]_  = \new_[14264]_  & \new_[14259]_ ;
  assign \new_[14269]_  = A298 & A268;
  assign \new_[14270]_  = ~A203 & \new_[14269]_ ;
  assign \new_[14274]_  = ~A301 & ~A300;
  assign \new_[14275]_  = A299 & \new_[14274]_ ;
  assign \new_[14276]_  = \new_[14275]_  & \new_[14270]_ ;
  assign \new_[14279]_  = ~A169 & ~A170;
  assign \new_[14283]_  = ~A202 & ~A201;
  assign \new_[14284]_  = ~A168 & \new_[14283]_ ;
  assign \new_[14285]_  = \new_[14284]_  & \new_[14279]_ ;
  assign \new_[14289]_  = A267 & A265;
  assign \new_[14290]_  = ~A203 & \new_[14289]_ ;
  assign \new_[14294]_  = ~A302 & ~A301;
  assign \new_[14295]_  = ~A300 & \new_[14294]_ ;
  assign \new_[14296]_  = \new_[14295]_  & \new_[14290]_ ;
  assign \new_[14299]_  = ~A169 & ~A170;
  assign \new_[14303]_  = ~A202 & ~A201;
  assign \new_[14304]_  = ~A168 & \new_[14303]_ ;
  assign \new_[14305]_  = \new_[14304]_  & \new_[14299]_ ;
  assign \new_[14309]_  = A267 & A265;
  assign \new_[14310]_  = ~A203 & \new_[14309]_ ;
  assign \new_[14314]_  = ~A301 & ~A299;
  assign \new_[14315]_  = ~A298 & \new_[14314]_ ;
  assign \new_[14316]_  = \new_[14315]_  & \new_[14310]_ ;
  assign \new_[14319]_  = ~A169 & ~A170;
  assign \new_[14323]_  = ~A202 & ~A201;
  assign \new_[14324]_  = ~A168 & \new_[14323]_ ;
  assign \new_[14325]_  = \new_[14324]_  & \new_[14319]_ ;
  assign \new_[14329]_  = A267 & A266;
  assign \new_[14330]_  = ~A203 & \new_[14329]_ ;
  assign \new_[14334]_  = ~A302 & ~A301;
  assign \new_[14335]_  = ~A300 & \new_[14334]_ ;
  assign \new_[14336]_  = \new_[14335]_  & \new_[14330]_ ;
  assign \new_[14339]_  = ~A169 & ~A170;
  assign \new_[14343]_  = ~A202 & ~A201;
  assign \new_[14344]_  = ~A168 & \new_[14343]_ ;
  assign \new_[14345]_  = \new_[14344]_  & \new_[14339]_ ;
  assign \new_[14349]_  = A267 & A266;
  assign \new_[14350]_  = ~A203 & \new_[14349]_ ;
  assign \new_[14354]_  = ~A301 & ~A299;
  assign \new_[14355]_  = ~A298 & \new_[14354]_ ;
  assign \new_[14356]_  = \new_[14355]_  & \new_[14350]_ ;
  assign \new_[14359]_  = ~A169 & ~A170;
  assign \new_[14363]_  = A201 & A199;
  assign \new_[14364]_  = ~A168 & \new_[14363]_ ;
  assign \new_[14365]_  = \new_[14364]_  & \new_[14359]_ ;
  assign \new_[14369]_  = ~A269 & ~A268;
  assign \new_[14370]_  = ~A267 & \new_[14369]_ ;
  assign \new_[14374]_  = A302 & ~A299;
  assign \new_[14375]_  = A298 & \new_[14374]_ ;
  assign \new_[14376]_  = \new_[14375]_  & \new_[14370]_ ;
  assign \new_[14379]_  = ~A169 & ~A170;
  assign \new_[14383]_  = A201 & A199;
  assign \new_[14384]_  = ~A168 & \new_[14383]_ ;
  assign \new_[14385]_  = \new_[14384]_  & \new_[14379]_ ;
  assign \new_[14389]_  = ~A269 & ~A268;
  assign \new_[14390]_  = ~A267 & \new_[14389]_ ;
  assign \new_[14394]_  = A302 & A299;
  assign \new_[14395]_  = ~A298 & \new_[14394]_ ;
  assign \new_[14396]_  = \new_[14395]_  & \new_[14390]_ ;
  assign \new_[14399]_  = ~A169 & ~A170;
  assign \new_[14403]_  = A201 & A199;
  assign \new_[14404]_  = ~A168 & \new_[14403]_ ;
  assign \new_[14405]_  = \new_[14404]_  & \new_[14399]_ ;
  assign \new_[14409]_  = ~A267 & A266;
  assign \new_[14410]_  = A265 & \new_[14409]_ ;
  assign \new_[14414]_  = A300 & A299;
  assign \new_[14415]_  = ~A268 & \new_[14414]_ ;
  assign \new_[14416]_  = \new_[14415]_  & \new_[14410]_ ;
  assign \new_[14419]_  = ~A169 & ~A170;
  assign \new_[14423]_  = A201 & A199;
  assign \new_[14424]_  = ~A168 & \new_[14423]_ ;
  assign \new_[14425]_  = \new_[14424]_  & \new_[14419]_ ;
  assign \new_[14429]_  = ~A267 & A266;
  assign \new_[14430]_  = A265 & \new_[14429]_ ;
  assign \new_[14434]_  = A300 & A298;
  assign \new_[14435]_  = ~A268 & \new_[14434]_ ;
  assign \new_[14436]_  = \new_[14435]_  & \new_[14430]_ ;
  assign \new_[14439]_  = ~A169 & ~A170;
  assign \new_[14443]_  = A201 & A199;
  assign \new_[14444]_  = ~A168 & \new_[14443]_ ;
  assign \new_[14445]_  = \new_[14444]_  & \new_[14439]_ ;
  assign \new_[14449]_  = ~A268 & ~A266;
  assign \new_[14450]_  = ~A265 & \new_[14449]_ ;
  assign \new_[14454]_  = A302 & ~A299;
  assign \new_[14455]_  = A298 & \new_[14454]_ ;
  assign \new_[14456]_  = \new_[14455]_  & \new_[14450]_ ;
  assign \new_[14459]_  = ~A169 & ~A170;
  assign \new_[14463]_  = A201 & A199;
  assign \new_[14464]_  = ~A168 & \new_[14463]_ ;
  assign \new_[14465]_  = \new_[14464]_  & \new_[14459]_ ;
  assign \new_[14469]_  = ~A268 & ~A266;
  assign \new_[14470]_  = ~A265 & \new_[14469]_ ;
  assign \new_[14474]_  = A302 & A299;
  assign \new_[14475]_  = ~A298 & \new_[14474]_ ;
  assign \new_[14476]_  = \new_[14475]_  & \new_[14470]_ ;
  assign \new_[14479]_  = ~A169 & ~A170;
  assign \new_[14483]_  = A201 & A200;
  assign \new_[14484]_  = ~A168 & \new_[14483]_ ;
  assign \new_[14485]_  = \new_[14484]_  & \new_[14479]_ ;
  assign \new_[14489]_  = ~A269 & ~A268;
  assign \new_[14490]_  = ~A267 & \new_[14489]_ ;
  assign \new_[14494]_  = A302 & ~A299;
  assign \new_[14495]_  = A298 & \new_[14494]_ ;
  assign \new_[14496]_  = \new_[14495]_  & \new_[14490]_ ;
  assign \new_[14499]_  = ~A169 & ~A170;
  assign \new_[14503]_  = A201 & A200;
  assign \new_[14504]_  = ~A168 & \new_[14503]_ ;
  assign \new_[14505]_  = \new_[14504]_  & \new_[14499]_ ;
  assign \new_[14509]_  = ~A269 & ~A268;
  assign \new_[14510]_  = ~A267 & \new_[14509]_ ;
  assign \new_[14514]_  = A302 & A299;
  assign \new_[14515]_  = ~A298 & \new_[14514]_ ;
  assign \new_[14516]_  = \new_[14515]_  & \new_[14510]_ ;
  assign \new_[14519]_  = ~A169 & ~A170;
  assign \new_[14523]_  = A201 & A200;
  assign \new_[14524]_  = ~A168 & \new_[14523]_ ;
  assign \new_[14525]_  = \new_[14524]_  & \new_[14519]_ ;
  assign \new_[14529]_  = ~A267 & A266;
  assign \new_[14530]_  = A265 & \new_[14529]_ ;
  assign \new_[14534]_  = A300 & A299;
  assign \new_[14535]_  = ~A268 & \new_[14534]_ ;
  assign \new_[14536]_  = \new_[14535]_  & \new_[14530]_ ;
  assign \new_[14539]_  = ~A169 & ~A170;
  assign \new_[14543]_  = A201 & A200;
  assign \new_[14544]_  = ~A168 & \new_[14543]_ ;
  assign \new_[14545]_  = \new_[14544]_  & \new_[14539]_ ;
  assign \new_[14549]_  = ~A267 & A266;
  assign \new_[14550]_  = A265 & \new_[14549]_ ;
  assign \new_[14554]_  = A300 & A298;
  assign \new_[14555]_  = ~A268 & \new_[14554]_ ;
  assign \new_[14556]_  = \new_[14555]_  & \new_[14550]_ ;
  assign \new_[14559]_  = ~A169 & ~A170;
  assign \new_[14563]_  = A201 & A200;
  assign \new_[14564]_  = ~A168 & \new_[14563]_ ;
  assign \new_[14565]_  = \new_[14564]_  & \new_[14559]_ ;
  assign \new_[14569]_  = ~A268 & ~A266;
  assign \new_[14570]_  = ~A265 & \new_[14569]_ ;
  assign \new_[14574]_  = A302 & ~A299;
  assign \new_[14575]_  = A298 & \new_[14574]_ ;
  assign \new_[14576]_  = \new_[14575]_  & \new_[14570]_ ;
  assign \new_[14579]_  = ~A169 & ~A170;
  assign \new_[14583]_  = A201 & A200;
  assign \new_[14584]_  = ~A168 & \new_[14583]_ ;
  assign \new_[14585]_  = \new_[14584]_  & \new_[14579]_ ;
  assign \new_[14589]_  = ~A268 & ~A266;
  assign \new_[14590]_  = ~A265 & \new_[14589]_ ;
  assign \new_[14594]_  = A302 & A299;
  assign \new_[14595]_  = ~A298 & \new_[14594]_ ;
  assign \new_[14596]_  = \new_[14595]_  & \new_[14590]_ ;
  assign \new_[14599]_  = ~A169 & ~A170;
  assign \new_[14603]_  = A200 & A199;
  assign \new_[14604]_  = ~A168 & \new_[14603]_ ;
  assign \new_[14605]_  = \new_[14604]_  & \new_[14599]_ ;
  assign \new_[14609]_  = A268 & ~A202;
  assign \new_[14610]_  = ~A201 & \new_[14609]_ ;
  assign \new_[14614]_  = ~A302 & ~A301;
  assign \new_[14615]_  = ~A300 & \new_[14614]_ ;
  assign \new_[14616]_  = \new_[14615]_  & \new_[14610]_ ;
  assign \new_[14619]_  = ~A169 & ~A170;
  assign \new_[14623]_  = A200 & A199;
  assign \new_[14624]_  = ~A168 & \new_[14623]_ ;
  assign \new_[14625]_  = \new_[14624]_  & \new_[14619]_ ;
  assign \new_[14629]_  = A268 & ~A202;
  assign \new_[14630]_  = ~A201 & \new_[14629]_ ;
  assign \new_[14634]_  = ~A301 & ~A299;
  assign \new_[14635]_  = ~A298 & \new_[14634]_ ;
  assign \new_[14636]_  = \new_[14635]_  & \new_[14630]_ ;
  assign \new_[14639]_  = ~A169 & ~A170;
  assign \new_[14643]_  = A200 & ~A199;
  assign \new_[14644]_  = ~A168 & \new_[14643]_ ;
  assign \new_[14645]_  = \new_[14644]_  & \new_[14639]_ ;
  assign \new_[14649]_  = ~A268 & ~A267;
  assign \new_[14650]_  = A203 & \new_[14649]_ ;
  assign \new_[14654]_  = A300 & A299;
  assign \new_[14655]_  = ~A269 & \new_[14654]_ ;
  assign \new_[14656]_  = \new_[14655]_  & \new_[14650]_ ;
  assign \new_[14659]_  = ~A169 & ~A170;
  assign \new_[14663]_  = A200 & ~A199;
  assign \new_[14664]_  = ~A168 & \new_[14663]_ ;
  assign \new_[14665]_  = \new_[14664]_  & \new_[14659]_ ;
  assign \new_[14669]_  = ~A268 & ~A267;
  assign \new_[14670]_  = A203 & \new_[14669]_ ;
  assign \new_[14674]_  = A300 & A298;
  assign \new_[14675]_  = ~A269 & \new_[14674]_ ;
  assign \new_[14676]_  = \new_[14675]_  & \new_[14670]_ ;
  assign \new_[14679]_  = ~A169 & ~A170;
  assign \new_[14683]_  = A200 & ~A199;
  assign \new_[14684]_  = ~A168 & \new_[14683]_ ;
  assign \new_[14685]_  = \new_[14684]_  & \new_[14679]_ ;
  assign \new_[14689]_  = A266 & A265;
  assign \new_[14690]_  = A203 & \new_[14689]_ ;
  assign \new_[14694]_  = A301 & ~A268;
  assign \new_[14695]_  = ~A267 & \new_[14694]_ ;
  assign \new_[14696]_  = \new_[14695]_  & \new_[14690]_ ;
  assign \new_[14699]_  = ~A169 & ~A170;
  assign \new_[14703]_  = A200 & ~A199;
  assign \new_[14704]_  = ~A168 & \new_[14703]_ ;
  assign \new_[14705]_  = \new_[14704]_  & \new_[14699]_ ;
  assign \new_[14709]_  = ~A266 & ~A265;
  assign \new_[14710]_  = A203 & \new_[14709]_ ;
  assign \new_[14714]_  = A300 & A299;
  assign \new_[14715]_  = ~A268 & \new_[14714]_ ;
  assign \new_[14716]_  = \new_[14715]_  & \new_[14710]_ ;
  assign \new_[14719]_  = ~A169 & ~A170;
  assign \new_[14723]_  = A200 & ~A199;
  assign \new_[14724]_  = ~A168 & \new_[14723]_ ;
  assign \new_[14725]_  = \new_[14724]_  & \new_[14719]_ ;
  assign \new_[14729]_  = ~A266 & ~A265;
  assign \new_[14730]_  = A203 & \new_[14729]_ ;
  assign \new_[14734]_  = A300 & A298;
  assign \new_[14735]_  = ~A268 & \new_[14734]_ ;
  assign \new_[14736]_  = \new_[14735]_  & \new_[14730]_ ;
  assign \new_[14739]_  = ~A169 & ~A170;
  assign \new_[14743]_  = ~A200 & A199;
  assign \new_[14744]_  = ~A168 & \new_[14743]_ ;
  assign \new_[14745]_  = \new_[14744]_  & \new_[14739]_ ;
  assign \new_[14749]_  = ~A268 & ~A267;
  assign \new_[14750]_  = A203 & \new_[14749]_ ;
  assign \new_[14754]_  = A300 & A299;
  assign \new_[14755]_  = ~A269 & \new_[14754]_ ;
  assign \new_[14756]_  = \new_[14755]_  & \new_[14750]_ ;
  assign \new_[14759]_  = ~A169 & ~A170;
  assign \new_[14763]_  = ~A200 & A199;
  assign \new_[14764]_  = ~A168 & \new_[14763]_ ;
  assign \new_[14765]_  = \new_[14764]_  & \new_[14759]_ ;
  assign \new_[14769]_  = ~A268 & ~A267;
  assign \new_[14770]_  = A203 & \new_[14769]_ ;
  assign \new_[14774]_  = A300 & A298;
  assign \new_[14775]_  = ~A269 & \new_[14774]_ ;
  assign \new_[14776]_  = \new_[14775]_  & \new_[14770]_ ;
  assign \new_[14779]_  = ~A169 & ~A170;
  assign \new_[14783]_  = ~A200 & A199;
  assign \new_[14784]_  = ~A168 & \new_[14783]_ ;
  assign \new_[14785]_  = \new_[14784]_  & \new_[14779]_ ;
  assign \new_[14789]_  = A266 & A265;
  assign \new_[14790]_  = A203 & \new_[14789]_ ;
  assign \new_[14794]_  = A301 & ~A268;
  assign \new_[14795]_  = ~A267 & \new_[14794]_ ;
  assign \new_[14796]_  = \new_[14795]_  & \new_[14790]_ ;
  assign \new_[14799]_  = ~A169 & ~A170;
  assign \new_[14803]_  = ~A200 & A199;
  assign \new_[14804]_  = ~A168 & \new_[14803]_ ;
  assign \new_[14805]_  = \new_[14804]_  & \new_[14799]_ ;
  assign \new_[14809]_  = ~A266 & ~A265;
  assign \new_[14810]_  = A203 & \new_[14809]_ ;
  assign \new_[14814]_  = A300 & A299;
  assign \new_[14815]_  = ~A268 & \new_[14814]_ ;
  assign \new_[14816]_  = \new_[14815]_  & \new_[14810]_ ;
  assign \new_[14819]_  = ~A169 & ~A170;
  assign \new_[14823]_  = ~A200 & A199;
  assign \new_[14824]_  = ~A168 & \new_[14823]_ ;
  assign \new_[14825]_  = \new_[14824]_  & \new_[14819]_ ;
  assign \new_[14829]_  = ~A266 & ~A265;
  assign \new_[14830]_  = A203 & \new_[14829]_ ;
  assign \new_[14834]_  = A300 & A298;
  assign \new_[14835]_  = ~A268 & \new_[14834]_ ;
  assign \new_[14836]_  = \new_[14835]_  & \new_[14830]_ ;
  assign \new_[14839]_  = ~A169 & ~A170;
  assign \new_[14843]_  = ~A200 & ~A199;
  assign \new_[14844]_  = ~A168 & \new_[14843]_ ;
  assign \new_[14845]_  = \new_[14844]_  & \new_[14839]_ ;
  assign \new_[14849]_  = A298 & A268;
  assign \new_[14850]_  = ~A202 & \new_[14849]_ ;
  assign \new_[14854]_  = ~A301 & ~A300;
  assign \new_[14855]_  = A299 & \new_[14854]_ ;
  assign \new_[14856]_  = \new_[14855]_  & \new_[14850]_ ;
  assign \new_[14859]_  = ~A169 & ~A170;
  assign \new_[14863]_  = ~A200 & ~A199;
  assign \new_[14864]_  = ~A168 & \new_[14863]_ ;
  assign \new_[14865]_  = \new_[14864]_  & \new_[14859]_ ;
  assign \new_[14869]_  = A267 & A265;
  assign \new_[14870]_  = ~A202 & \new_[14869]_ ;
  assign \new_[14874]_  = ~A302 & ~A301;
  assign \new_[14875]_  = ~A300 & \new_[14874]_ ;
  assign \new_[14876]_  = \new_[14875]_  & \new_[14870]_ ;
  assign \new_[14879]_  = ~A169 & ~A170;
  assign \new_[14883]_  = ~A200 & ~A199;
  assign \new_[14884]_  = ~A168 & \new_[14883]_ ;
  assign \new_[14885]_  = \new_[14884]_  & \new_[14879]_ ;
  assign \new_[14889]_  = A267 & A265;
  assign \new_[14890]_  = ~A202 & \new_[14889]_ ;
  assign \new_[14894]_  = ~A301 & ~A299;
  assign \new_[14895]_  = ~A298 & \new_[14894]_ ;
  assign \new_[14896]_  = \new_[14895]_  & \new_[14890]_ ;
  assign \new_[14899]_  = ~A169 & ~A170;
  assign \new_[14903]_  = ~A200 & ~A199;
  assign \new_[14904]_  = ~A168 & \new_[14903]_ ;
  assign \new_[14905]_  = \new_[14904]_  & \new_[14899]_ ;
  assign \new_[14909]_  = A267 & A266;
  assign \new_[14910]_  = ~A202 & \new_[14909]_ ;
  assign \new_[14914]_  = ~A302 & ~A301;
  assign \new_[14915]_  = ~A300 & \new_[14914]_ ;
  assign \new_[14916]_  = \new_[14915]_  & \new_[14910]_ ;
  assign \new_[14919]_  = ~A169 & ~A170;
  assign \new_[14923]_  = ~A200 & ~A199;
  assign \new_[14924]_  = ~A168 & \new_[14923]_ ;
  assign \new_[14925]_  = \new_[14924]_  & \new_[14919]_ ;
  assign \new_[14929]_  = A267 & A266;
  assign \new_[14930]_  = ~A202 & \new_[14929]_ ;
  assign \new_[14934]_  = ~A301 & ~A299;
  assign \new_[14935]_  = ~A298 & \new_[14934]_ ;
  assign \new_[14936]_  = \new_[14935]_  & \new_[14930]_ ;
  assign \new_[14940]_  = ~A201 & A166;
  assign \new_[14941]_  = A168 & \new_[14940]_ ;
  assign \new_[14945]_  = A265 & ~A203;
  assign \new_[14946]_  = ~A202 & \new_[14945]_ ;
  assign \new_[14947]_  = \new_[14946]_  & \new_[14941]_ ;
  assign \new_[14951]_  = ~A268 & ~A267;
  assign \new_[14952]_  = A266 & \new_[14951]_ ;
  assign \new_[14956]_  = A302 & ~A299;
  assign \new_[14957]_  = A298 & \new_[14956]_ ;
  assign \new_[14958]_  = \new_[14957]_  & \new_[14952]_ ;
  assign \new_[14962]_  = ~A201 & A166;
  assign \new_[14963]_  = A168 & \new_[14962]_ ;
  assign \new_[14967]_  = A265 & ~A203;
  assign \new_[14968]_  = ~A202 & \new_[14967]_ ;
  assign \new_[14969]_  = \new_[14968]_  & \new_[14963]_ ;
  assign \new_[14973]_  = ~A268 & ~A267;
  assign \new_[14974]_  = A266 & \new_[14973]_ ;
  assign \new_[14978]_  = A302 & A299;
  assign \new_[14979]_  = ~A298 & \new_[14978]_ ;
  assign \new_[14980]_  = \new_[14979]_  & \new_[14974]_ ;
  assign \new_[14984]_  = A199 & A166;
  assign \new_[14985]_  = A168 & \new_[14984]_ ;
  assign \new_[14989]_  = ~A202 & ~A201;
  assign \new_[14990]_  = A200 & \new_[14989]_ ;
  assign \new_[14991]_  = \new_[14990]_  & \new_[14985]_ ;
  assign \new_[14995]_  = ~A269 & ~A268;
  assign \new_[14996]_  = ~A267 & \new_[14995]_ ;
  assign \new_[15000]_  = A302 & ~A299;
  assign \new_[15001]_  = A298 & \new_[15000]_ ;
  assign \new_[15002]_  = \new_[15001]_  & \new_[14996]_ ;
  assign \new_[15006]_  = A199 & A166;
  assign \new_[15007]_  = A168 & \new_[15006]_ ;
  assign \new_[15011]_  = ~A202 & ~A201;
  assign \new_[15012]_  = A200 & \new_[15011]_ ;
  assign \new_[15013]_  = \new_[15012]_  & \new_[15007]_ ;
  assign \new_[15017]_  = ~A269 & ~A268;
  assign \new_[15018]_  = ~A267 & \new_[15017]_ ;
  assign \new_[15022]_  = A302 & A299;
  assign \new_[15023]_  = ~A298 & \new_[15022]_ ;
  assign \new_[15024]_  = \new_[15023]_  & \new_[15018]_ ;
  assign \new_[15028]_  = A199 & A166;
  assign \new_[15029]_  = A168 & \new_[15028]_ ;
  assign \new_[15033]_  = ~A202 & ~A201;
  assign \new_[15034]_  = A200 & \new_[15033]_ ;
  assign \new_[15035]_  = \new_[15034]_  & \new_[15029]_ ;
  assign \new_[15039]_  = ~A267 & A266;
  assign \new_[15040]_  = A265 & \new_[15039]_ ;
  assign \new_[15044]_  = A300 & A299;
  assign \new_[15045]_  = ~A268 & \new_[15044]_ ;
  assign \new_[15046]_  = \new_[15045]_  & \new_[15040]_ ;
  assign \new_[15050]_  = A199 & A166;
  assign \new_[15051]_  = A168 & \new_[15050]_ ;
  assign \new_[15055]_  = ~A202 & ~A201;
  assign \new_[15056]_  = A200 & \new_[15055]_ ;
  assign \new_[15057]_  = \new_[15056]_  & \new_[15051]_ ;
  assign \new_[15061]_  = ~A267 & A266;
  assign \new_[15062]_  = A265 & \new_[15061]_ ;
  assign \new_[15066]_  = A300 & A298;
  assign \new_[15067]_  = ~A268 & \new_[15066]_ ;
  assign \new_[15068]_  = \new_[15067]_  & \new_[15062]_ ;
  assign \new_[15072]_  = A199 & A166;
  assign \new_[15073]_  = A168 & \new_[15072]_ ;
  assign \new_[15077]_  = ~A202 & ~A201;
  assign \new_[15078]_  = A200 & \new_[15077]_ ;
  assign \new_[15079]_  = \new_[15078]_  & \new_[15073]_ ;
  assign \new_[15083]_  = ~A268 & ~A266;
  assign \new_[15084]_  = ~A265 & \new_[15083]_ ;
  assign \new_[15088]_  = A302 & ~A299;
  assign \new_[15089]_  = A298 & \new_[15088]_ ;
  assign \new_[15090]_  = \new_[15089]_  & \new_[15084]_ ;
  assign \new_[15094]_  = A199 & A166;
  assign \new_[15095]_  = A168 & \new_[15094]_ ;
  assign \new_[15099]_  = ~A202 & ~A201;
  assign \new_[15100]_  = A200 & \new_[15099]_ ;
  assign \new_[15101]_  = \new_[15100]_  & \new_[15095]_ ;
  assign \new_[15105]_  = ~A268 & ~A266;
  assign \new_[15106]_  = ~A265 & \new_[15105]_ ;
  assign \new_[15110]_  = A302 & A299;
  assign \new_[15111]_  = ~A298 & \new_[15110]_ ;
  assign \new_[15112]_  = \new_[15111]_  & \new_[15106]_ ;
  assign \new_[15116]_  = ~A199 & A166;
  assign \new_[15117]_  = A168 & \new_[15116]_ ;
  assign \new_[15121]_  = ~A265 & A203;
  assign \new_[15122]_  = A200 & \new_[15121]_ ;
  assign \new_[15123]_  = \new_[15122]_  & \new_[15117]_ ;
  assign \new_[15127]_  = A298 & A269;
  assign \new_[15128]_  = A266 & \new_[15127]_ ;
  assign \new_[15132]_  = ~A301 & ~A300;
  assign \new_[15133]_  = A299 & \new_[15132]_ ;
  assign \new_[15134]_  = \new_[15133]_  & \new_[15128]_ ;
  assign \new_[15138]_  = ~A199 & A166;
  assign \new_[15139]_  = A168 & \new_[15138]_ ;
  assign \new_[15143]_  = A265 & A203;
  assign \new_[15144]_  = A200 & \new_[15143]_ ;
  assign \new_[15145]_  = \new_[15144]_  & \new_[15139]_ ;
  assign \new_[15149]_  = A298 & A269;
  assign \new_[15150]_  = ~A266 & \new_[15149]_ ;
  assign \new_[15154]_  = ~A301 & ~A300;
  assign \new_[15155]_  = A299 & \new_[15154]_ ;
  assign \new_[15156]_  = \new_[15155]_  & \new_[15150]_ ;
  assign \new_[15160]_  = A199 & A166;
  assign \new_[15161]_  = A168 & \new_[15160]_ ;
  assign \new_[15165]_  = ~A265 & A203;
  assign \new_[15166]_  = ~A200 & \new_[15165]_ ;
  assign \new_[15167]_  = \new_[15166]_  & \new_[15161]_ ;
  assign \new_[15171]_  = A298 & A269;
  assign \new_[15172]_  = A266 & \new_[15171]_ ;
  assign \new_[15176]_  = ~A301 & ~A300;
  assign \new_[15177]_  = A299 & \new_[15176]_ ;
  assign \new_[15178]_  = \new_[15177]_  & \new_[15172]_ ;
  assign \new_[15182]_  = A199 & A166;
  assign \new_[15183]_  = A168 & \new_[15182]_ ;
  assign \new_[15187]_  = A265 & A203;
  assign \new_[15188]_  = ~A200 & \new_[15187]_ ;
  assign \new_[15189]_  = \new_[15188]_  & \new_[15183]_ ;
  assign \new_[15193]_  = A298 & A269;
  assign \new_[15194]_  = ~A266 & \new_[15193]_ ;
  assign \new_[15198]_  = ~A301 & ~A300;
  assign \new_[15199]_  = A299 & \new_[15198]_ ;
  assign \new_[15200]_  = \new_[15199]_  & \new_[15194]_ ;
  assign \new_[15204]_  = ~A199 & A166;
  assign \new_[15205]_  = A168 & \new_[15204]_ ;
  assign \new_[15209]_  = A265 & ~A202;
  assign \new_[15210]_  = ~A200 & \new_[15209]_ ;
  assign \new_[15211]_  = \new_[15210]_  & \new_[15205]_ ;
  assign \new_[15215]_  = ~A268 & ~A267;
  assign \new_[15216]_  = A266 & \new_[15215]_ ;
  assign \new_[15220]_  = A302 & ~A299;
  assign \new_[15221]_  = A298 & \new_[15220]_ ;
  assign \new_[15222]_  = \new_[15221]_  & \new_[15216]_ ;
  assign \new_[15226]_  = ~A199 & A166;
  assign \new_[15227]_  = A168 & \new_[15226]_ ;
  assign \new_[15231]_  = A265 & ~A202;
  assign \new_[15232]_  = ~A200 & \new_[15231]_ ;
  assign \new_[15233]_  = \new_[15232]_  & \new_[15227]_ ;
  assign \new_[15237]_  = ~A268 & ~A267;
  assign \new_[15238]_  = A266 & \new_[15237]_ ;
  assign \new_[15242]_  = A302 & A299;
  assign \new_[15243]_  = ~A298 & \new_[15242]_ ;
  assign \new_[15244]_  = \new_[15243]_  & \new_[15238]_ ;
  assign \new_[15248]_  = ~A201 & A167;
  assign \new_[15249]_  = A168 & \new_[15248]_ ;
  assign \new_[15253]_  = A265 & ~A203;
  assign \new_[15254]_  = ~A202 & \new_[15253]_ ;
  assign \new_[15255]_  = \new_[15254]_  & \new_[15249]_ ;
  assign \new_[15259]_  = ~A268 & ~A267;
  assign \new_[15260]_  = A266 & \new_[15259]_ ;
  assign \new_[15264]_  = A302 & ~A299;
  assign \new_[15265]_  = A298 & \new_[15264]_ ;
  assign \new_[15266]_  = \new_[15265]_  & \new_[15260]_ ;
  assign \new_[15270]_  = ~A201 & A167;
  assign \new_[15271]_  = A168 & \new_[15270]_ ;
  assign \new_[15275]_  = A265 & ~A203;
  assign \new_[15276]_  = ~A202 & \new_[15275]_ ;
  assign \new_[15277]_  = \new_[15276]_  & \new_[15271]_ ;
  assign \new_[15281]_  = ~A268 & ~A267;
  assign \new_[15282]_  = A266 & \new_[15281]_ ;
  assign \new_[15286]_  = A302 & A299;
  assign \new_[15287]_  = ~A298 & \new_[15286]_ ;
  assign \new_[15288]_  = \new_[15287]_  & \new_[15282]_ ;
  assign \new_[15292]_  = A199 & A167;
  assign \new_[15293]_  = A168 & \new_[15292]_ ;
  assign \new_[15297]_  = ~A202 & ~A201;
  assign \new_[15298]_  = A200 & \new_[15297]_ ;
  assign \new_[15299]_  = \new_[15298]_  & \new_[15293]_ ;
  assign \new_[15303]_  = ~A269 & ~A268;
  assign \new_[15304]_  = ~A267 & \new_[15303]_ ;
  assign \new_[15308]_  = A302 & ~A299;
  assign \new_[15309]_  = A298 & \new_[15308]_ ;
  assign \new_[15310]_  = \new_[15309]_  & \new_[15304]_ ;
  assign \new_[15314]_  = A199 & A167;
  assign \new_[15315]_  = A168 & \new_[15314]_ ;
  assign \new_[15319]_  = ~A202 & ~A201;
  assign \new_[15320]_  = A200 & \new_[15319]_ ;
  assign \new_[15321]_  = \new_[15320]_  & \new_[15315]_ ;
  assign \new_[15325]_  = ~A269 & ~A268;
  assign \new_[15326]_  = ~A267 & \new_[15325]_ ;
  assign \new_[15330]_  = A302 & A299;
  assign \new_[15331]_  = ~A298 & \new_[15330]_ ;
  assign \new_[15332]_  = \new_[15331]_  & \new_[15326]_ ;
  assign \new_[15336]_  = A199 & A167;
  assign \new_[15337]_  = A168 & \new_[15336]_ ;
  assign \new_[15341]_  = ~A202 & ~A201;
  assign \new_[15342]_  = A200 & \new_[15341]_ ;
  assign \new_[15343]_  = \new_[15342]_  & \new_[15337]_ ;
  assign \new_[15347]_  = ~A267 & A266;
  assign \new_[15348]_  = A265 & \new_[15347]_ ;
  assign \new_[15352]_  = A300 & A299;
  assign \new_[15353]_  = ~A268 & \new_[15352]_ ;
  assign \new_[15354]_  = \new_[15353]_  & \new_[15348]_ ;
  assign \new_[15358]_  = A199 & A167;
  assign \new_[15359]_  = A168 & \new_[15358]_ ;
  assign \new_[15363]_  = ~A202 & ~A201;
  assign \new_[15364]_  = A200 & \new_[15363]_ ;
  assign \new_[15365]_  = \new_[15364]_  & \new_[15359]_ ;
  assign \new_[15369]_  = ~A267 & A266;
  assign \new_[15370]_  = A265 & \new_[15369]_ ;
  assign \new_[15374]_  = A300 & A298;
  assign \new_[15375]_  = ~A268 & \new_[15374]_ ;
  assign \new_[15376]_  = \new_[15375]_  & \new_[15370]_ ;
  assign \new_[15380]_  = A199 & A167;
  assign \new_[15381]_  = A168 & \new_[15380]_ ;
  assign \new_[15385]_  = ~A202 & ~A201;
  assign \new_[15386]_  = A200 & \new_[15385]_ ;
  assign \new_[15387]_  = \new_[15386]_  & \new_[15381]_ ;
  assign \new_[15391]_  = ~A268 & ~A266;
  assign \new_[15392]_  = ~A265 & \new_[15391]_ ;
  assign \new_[15396]_  = A302 & ~A299;
  assign \new_[15397]_  = A298 & \new_[15396]_ ;
  assign \new_[15398]_  = \new_[15397]_  & \new_[15392]_ ;
  assign \new_[15402]_  = A199 & A167;
  assign \new_[15403]_  = A168 & \new_[15402]_ ;
  assign \new_[15407]_  = ~A202 & ~A201;
  assign \new_[15408]_  = A200 & \new_[15407]_ ;
  assign \new_[15409]_  = \new_[15408]_  & \new_[15403]_ ;
  assign \new_[15413]_  = ~A268 & ~A266;
  assign \new_[15414]_  = ~A265 & \new_[15413]_ ;
  assign \new_[15418]_  = A302 & A299;
  assign \new_[15419]_  = ~A298 & \new_[15418]_ ;
  assign \new_[15420]_  = \new_[15419]_  & \new_[15414]_ ;
  assign \new_[15424]_  = ~A199 & A167;
  assign \new_[15425]_  = A168 & \new_[15424]_ ;
  assign \new_[15429]_  = ~A265 & A203;
  assign \new_[15430]_  = A200 & \new_[15429]_ ;
  assign \new_[15431]_  = \new_[15430]_  & \new_[15425]_ ;
  assign \new_[15435]_  = A298 & A269;
  assign \new_[15436]_  = A266 & \new_[15435]_ ;
  assign \new_[15440]_  = ~A301 & ~A300;
  assign \new_[15441]_  = A299 & \new_[15440]_ ;
  assign \new_[15442]_  = \new_[15441]_  & \new_[15436]_ ;
  assign \new_[15446]_  = ~A199 & A167;
  assign \new_[15447]_  = A168 & \new_[15446]_ ;
  assign \new_[15451]_  = A265 & A203;
  assign \new_[15452]_  = A200 & \new_[15451]_ ;
  assign \new_[15453]_  = \new_[15452]_  & \new_[15447]_ ;
  assign \new_[15457]_  = A298 & A269;
  assign \new_[15458]_  = ~A266 & \new_[15457]_ ;
  assign \new_[15462]_  = ~A301 & ~A300;
  assign \new_[15463]_  = A299 & \new_[15462]_ ;
  assign \new_[15464]_  = \new_[15463]_  & \new_[15458]_ ;
  assign \new_[15468]_  = A199 & A167;
  assign \new_[15469]_  = A168 & \new_[15468]_ ;
  assign \new_[15473]_  = ~A265 & A203;
  assign \new_[15474]_  = ~A200 & \new_[15473]_ ;
  assign \new_[15475]_  = \new_[15474]_  & \new_[15469]_ ;
  assign \new_[15479]_  = A298 & A269;
  assign \new_[15480]_  = A266 & \new_[15479]_ ;
  assign \new_[15484]_  = ~A301 & ~A300;
  assign \new_[15485]_  = A299 & \new_[15484]_ ;
  assign \new_[15486]_  = \new_[15485]_  & \new_[15480]_ ;
  assign \new_[15490]_  = A199 & A167;
  assign \new_[15491]_  = A168 & \new_[15490]_ ;
  assign \new_[15495]_  = A265 & A203;
  assign \new_[15496]_  = ~A200 & \new_[15495]_ ;
  assign \new_[15497]_  = \new_[15496]_  & \new_[15491]_ ;
  assign \new_[15501]_  = A298 & A269;
  assign \new_[15502]_  = ~A266 & \new_[15501]_ ;
  assign \new_[15506]_  = ~A301 & ~A300;
  assign \new_[15507]_  = A299 & \new_[15506]_ ;
  assign \new_[15508]_  = \new_[15507]_  & \new_[15502]_ ;
  assign \new_[15512]_  = ~A199 & A167;
  assign \new_[15513]_  = A168 & \new_[15512]_ ;
  assign \new_[15517]_  = A265 & ~A202;
  assign \new_[15518]_  = ~A200 & \new_[15517]_ ;
  assign \new_[15519]_  = \new_[15518]_  & \new_[15513]_ ;
  assign \new_[15523]_  = ~A268 & ~A267;
  assign \new_[15524]_  = A266 & \new_[15523]_ ;
  assign \new_[15528]_  = A302 & ~A299;
  assign \new_[15529]_  = A298 & \new_[15528]_ ;
  assign \new_[15530]_  = \new_[15529]_  & \new_[15524]_ ;
  assign \new_[15534]_  = ~A199 & A167;
  assign \new_[15535]_  = A168 & \new_[15534]_ ;
  assign \new_[15539]_  = A265 & ~A202;
  assign \new_[15540]_  = ~A200 & \new_[15539]_ ;
  assign \new_[15541]_  = \new_[15540]_  & \new_[15535]_ ;
  assign \new_[15545]_  = ~A268 & ~A267;
  assign \new_[15546]_  = A266 & \new_[15545]_ ;
  assign \new_[15550]_  = A302 & A299;
  assign \new_[15551]_  = ~A298 & \new_[15550]_ ;
  assign \new_[15552]_  = \new_[15551]_  & \new_[15546]_ ;
  assign \new_[15556]_  = ~A166 & A167;
  assign \new_[15557]_  = A170 & \new_[15556]_ ;
  assign \new_[15561]_  = ~A203 & ~A202;
  assign \new_[15562]_  = ~A201 & \new_[15561]_ ;
  assign \new_[15563]_  = \new_[15562]_  & \new_[15557]_ ;
  assign \new_[15567]_  = ~A269 & ~A268;
  assign \new_[15568]_  = ~A267 & \new_[15567]_ ;
  assign \new_[15572]_  = A302 & ~A299;
  assign \new_[15573]_  = A298 & \new_[15572]_ ;
  assign \new_[15574]_  = \new_[15573]_  & \new_[15568]_ ;
  assign \new_[15578]_  = ~A166 & A167;
  assign \new_[15579]_  = A170 & \new_[15578]_ ;
  assign \new_[15583]_  = ~A203 & ~A202;
  assign \new_[15584]_  = ~A201 & \new_[15583]_ ;
  assign \new_[15585]_  = \new_[15584]_  & \new_[15579]_ ;
  assign \new_[15589]_  = ~A269 & ~A268;
  assign \new_[15590]_  = ~A267 & \new_[15589]_ ;
  assign \new_[15594]_  = A302 & A299;
  assign \new_[15595]_  = ~A298 & \new_[15594]_ ;
  assign \new_[15596]_  = \new_[15595]_  & \new_[15590]_ ;
  assign \new_[15600]_  = ~A166 & A167;
  assign \new_[15601]_  = A170 & \new_[15600]_ ;
  assign \new_[15605]_  = ~A203 & ~A202;
  assign \new_[15606]_  = ~A201 & \new_[15605]_ ;
  assign \new_[15607]_  = \new_[15606]_  & \new_[15601]_ ;
  assign \new_[15611]_  = ~A267 & A266;
  assign \new_[15612]_  = A265 & \new_[15611]_ ;
  assign \new_[15616]_  = A300 & A299;
  assign \new_[15617]_  = ~A268 & \new_[15616]_ ;
  assign \new_[15618]_  = \new_[15617]_  & \new_[15612]_ ;
  assign \new_[15622]_  = ~A166 & A167;
  assign \new_[15623]_  = A170 & \new_[15622]_ ;
  assign \new_[15627]_  = ~A203 & ~A202;
  assign \new_[15628]_  = ~A201 & \new_[15627]_ ;
  assign \new_[15629]_  = \new_[15628]_  & \new_[15623]_ ;
  assign \new_[15633]_  = ~A267 & A266;
  assign \new_[15634]_  = A265 & \new_[15633]_ ;
  assign \new_[15638]_  = A300 & A298;
  assign \new_[15639]_  = ~A268 & \new_[15638]_ ;
  assign \new_[15640]_  = \new_[15639]_  & \new_[15634]_ ;
  assign \new_[15644]_  = ~A166 & A167;
  assign \new_[15645]_  = A170 & \new_[15644]_ ;
  assign \new_[15649]_  = ~A203 & ~A202;
  assign \new_[15650]_  = ~A201 & \new_[15649]_ ;
  assign \new_[15651]_  = \new_[15650]_  & \new_[15645]_ ;
  assign \new_[15655]_  = ~A268 & ~A266;
  assign \new_[15656]_  = ~A265 & \new_[15655]_ ;
  assign \new_[15660]_  = A302 & ~A299;
  assign \new_[15661]_  = A298 & \new_[15660]_ ;
  assign \new_[15662]_  = \new_[15661]_  & \new_[15656]_ ;
  assign \new_[15666]_  = ~A166 & A167;
  assign \new_[15667]_  = A170 & \new_[15666]_ ;
  assign \new_[15671]_  = ~A203 & ~A202;
  assign \new_[15672]_  = ~A201 & \new_[15671]_ ;
  assign \new_[15673]_  = \new_[15672]_  & \new_[15667]_ ;
  assign \new_[15677]_  = ~A268 & ~A266;
  assign \new_[15678]_  = ~A265 & \new_[15677]_ ;
  assign \new_[15682]_  = A302 & A299;
  assign \new_[15683]_  = ~A298 & \new_[15682]_ ;
  assign \new_[15684]_  = \new_[15683]_  & \new_[15678]_ ;
  assign \new_[15688]_  = ~A166 & A167;
  assign \new_[15689]_  = A170 & \new_[15688]_ ;
  assign \new_[15693]_  = ~A265 & A201;
  assign \new_[15694]_  = A199 & \new_[15693]_ ;
  assign \new_[15695]_  = \new_[15694]_  & \new_[15689]_ ;
  assign \new_[15699]_  = A298 & A269;
  assign \new_[15700]_  = A266 & \new_[15699]_ ;
  assign \new_[15704]_  = ~A301 & ~A300;
  assign \new_[15705]_  = A299 & \new_[15704]_ ;
  assign \new_[15706]_  = \new_[15705]_  & \new_[15700]_ ;
  assign \new_[15710]_  = ~A166 & A167;
  assign \new_[15711]_  = A170 & \new_[15710]_ ;
  assign \new_[15715]_  = A265 & A201;
  assign \new_[15716]_  = A199 & \new_[15715]_ ;
  assign \new_[15717]_  = \new_[15716]_  & \new_[15711]_ ;
  assign \new_[15721]_  = A298 & A269;
  assign \new_[15722]_  = ~A266 & \new_[15721]_ ;
  assign \new_[15726]_  = ~A301 & ~A300;
  assign \new_[15727]_  = A299 & \new_[15726]_ ;
  assign \new_[15728]_  = \new_[15727]_  & \new_[15722]_ ;
  assign \new_[15732]_  = ~A166 & A167;
  assign \new_[15733]_  = A170 & \new_[15732]_ ;
  assign \new_[15737]_  = ~A265 & A201;
  assign \new_[15738]_  = A200 & \new_[15737]_ ;
  assign \new_[15739]_  = \new_[15738]_  & \new_[15733]_ ;
  assign \new_[15743]_  = A298 & A269;
  assign \new_[15744]_  = A266 & \new_[15743]_ ;
  assign \new_[15748]_  = ~A301 & ~A300;
  assign \new_[15749]_  = A299 & \new_[15748]_ ;
  assign \new_[15750]_  = \new_[15749]_  & \new_[15744]_ ;
  assign \new_[15754]_  = ~A166 & A167;
  assign \new_[15755]_  = A170 & \new_[15754]_ ;
  assign \new_[15759]_  = A265 & A201;
  assign \new_[15760]_  = A200 & \new_[15759]_ ;
  assign \new_[15761]_  = \new_[15760]_  & \new_[15755]_ ;
  assign \new_[15765]_  = A298 & A269;
  assign \new_[15766]_  = ~A266 & \new_[15765]_ ;
  assign \new_[15770]_  = ~A301 & ~A300;
  assign \new_[15771]_  = A299 & \new_[15770]_ ;
  assign \new_[15772]_  = \new_[15771]_  & \new_[15766]_ ;
  assign \new_[15776]_  = ~A166 & A167;
  assign \new_[15777]_  = A170 & \new_[15776]_ ;
  assign \new_[15781]_  = ~A201 & A200;
  assign \new_[15782]_  = A199 & \new_[15781]_ ;
  assign \new_[15783]_  = \new_[15782]_  & \new_[15777]_ ;
  assign \new_[15787]_  = ~A268 & ~A267;
  assign \new_[15788]_  = ~A202 & \new_[15787]_ ;
  assign \new_[15792]_  = A300 & A299;
  assign \new_[15793]_  = ~A269 & \new_[15792]_ ;
  assign \new_[15794]_  = \new_[15793]_  & \new_[15788]_ ;
  assign \new_[15798]_  = ~A166 & A167;
  assign \new_[15799]_  = A170 & \new_[15798]_ ;
  assign \new_[15803]_  = ~A201 & A200;
  assign \new_[15804]_  = A199 & \new_[15803]_ ;
  assign \new_[15805]_  = \new_[15804]_  & \new_[15799]_ ;
  assign \new_[15809]_  = ~A268 & ~A267;
  assign \new_[15810]_  = ~A202 & \new_[15809]_ ;
  assign \new_[15814]_  = A300 & A298;
  assign \new_[15815]_  = ~A269 & \new_[15814]_ ;
  assign \new_[15816]_  = \new_[15815]_  & \new_[15810]_ ;
  assign \new_[15820]_  = ~A166 & A167;
  assign \new_[15821]_  = A170 & \new_[15820]_ ;
  assign \new_[15825]_  = ~A201 & A200;
  assign \new_[15826]_  = A199 & \new_[15825]_ ;
  assign \new_[15827]_  = \new_[15826]_  & \new_[15821]_ ;
  assign \new_[15831]_  = A266 & A265;
  assign \new_[15832]_  = ~A202 & \new_[15831]_ ;
  assign \new_[15836]_  = A301 & ~A268;
  assign \new_[15837]_  = ~A267 & \new_[15836]_ ;
  assign \new_[15838]_  = \new_[15837]_  & \new_[15832]_ ;
  assign \new_[15842]_  = ~A166 & A167;
  assign \new_[15843]_  = A170 & \new_[15842]_ ;
  assign \new_[15847]_  = ~A201 & A200;
  assign \new_[15848]_  = A199 & \new_[15847]_ ;
  assign \new_[15849]_  = \new_[15848]_  & \new_[15843]_ ;
  assign \new_[15853]_  = ~A266 & ~A265;
  assign \new_[15854]_  = ~A202 & \new_[15853]_ ;
  assign \new_[15858]_  = A300 & A299;
  assign \new_[15859]_  = ~A268 & \new_[15858]_ ;
  assign \new_[15860]_  = \new_[15859]_  & \new_[15854]_ ;
  assign \new_[15864]_  = ~A166 & A167;
  assign \new_[15865]_  = A170 & \new_[15864]_ ;
  assign \new_[15869]_  = ~A201 & A200;
  assign \new_[15870]_  = A199 & \new_[15869]_ ;
  assign \new_[15871]_  = \new_[15870]_  & \new_[15865]_ ;
  assign \new_[15875]_  = ~A266 & ~A265;
  assign \new_[15876]_  = ~A202 & \new_[15875]_ ;
  assign \new_[15880]_  = A300 & A298;
  assign \new_[15881]_  = ~A268 & \new_[15880]_ ;
  assign \new_[15882]_  = \new_[15881]_  & \new_[15876]_ ;
  assign \new_[15886]_  = ~A166 & A167;
  assign \new_[15887]_  = A170 & \new_[15886]_ ;
  assign \new_[15891]_  = A203 & A200;
  assign \new_[15892]_  = ~A199 & \new_[15891]_ ;
  assign \new_[15893]_  = \new_[15892]_  & \new_[15887]_ ;
  assign \new_[15897]_  = A298 & A267;
  assign \new_[15898]_  = A265 & \new_[15897]_ ;
  assign \new_[15902]_  = ~A301 & ~A300;
  assign \new_[15903]_  = A299 & \new_[15902]_ ;
  assign \new_[15904]_  = \new_[15903]_  & \new_[15898]_ ;
  assign \new_[15908]_  = ~A166 & A167;
  assign \new_[15909]_  = A170 & \new_[15908]_ ;
  assign \new_[15913]_  = A203 & A200;
  assign \new_[15914]_  = ~A199 & \new_[15913]_ ;
  assign \new_[15915]_  = \new_[15914]_  & \new_[15909]_ ;
  assign \new_[15919]_  = A298 & A267;
  assign \new_[15920]_  = A266 & \new_[15919]_ ;
  assign \new_[15924]_  = ~A301 & ~A300;
  assign \new_[15925]_  = A299 & \new_[15924]_ ;
  assign \new_[15926]_  = \new_[15925]_  & \new_[15920]_ ;
  assign \new_[15930]_  = ~A166 & A167;
  assign \new_[15931]_  = A170 & \new_[15930]_ ;
  assign \new_[15935]_  = A203 & A200;
  assign \new_[15936]_  = ~A199 & \new_[15935]_ ;
  assign \new_[15937]_  = \new_[15936]_  & \new_[15931]_ ;
  assign \new_[15941]_  = A269 & A266;
  assign \new_[15942]_  = ~A265 & \new_[15941]_ ;
  assign \new_[15946]_  = ~A302 & ~A301;
  assign \new_[15947]_  = ~A300 & \new_[15946]_ ;
  assign \new_[15948]_  = \new_[15947]_  & \new_[15942]_ ;
  assign \new_[15952]_  = ~A166 & A167;
  assign \new_[15953]_  = A170 & \new_[15952]_ ;
  assign \new_[15957]_  = A203 & A200;
  assign \new_[15958]_  = ~A199 & \new_[15957]_ ;
  assign \new_[15959]_  = \new_[15958]_  & \new_[15953]_ ;
  assign \new_[15963]_  = A269 & A266;
  assign \new_[15964]_  = ~A265 & \new_[15963]_ ;
  assign \new_[15968]_  = ~A301 & ~A299;
  assign \new_[15969]_  = ~A298 & \new_[15968]_ ;
  assign \new_[15970]_  = \new_[15969]_  & \new_[15964]_ ;
  assign \new_[15974]_  = ~A166 & A167;
  assign \new_[15975]_  = A170 & \new_[15974]_ ;
  assign \new_[15979]_  = A203 & A200;
  assign \new_[15980]_  = ~A199 & \new_[15979]_ ;
  assign \new_[15981]_  = \new_[15980]_  & \new_[15975]_ ;
  assign \new_[15985]_  = A269 & ~A266;
  assign \new_[15986]_  = A265 & \new_[15985]_ ;
  assign \new_[15990]_  = ~A302 & ~A301;
  assign \new_[15991]_  = ~A300 & \new_[15990]_ ;
  assign \new_[15992]_  = \new_[15991]_  & \new_[15986]_ ;
  assign \new_[15996]_  = ~A166 & A167;
  assign \new_[15997]_  = A170 & \new_[15996]_ ;
  assign \new_[16001]_  = A203 & A200;
  assign \new_[16002]_  = ~A199 & \new_[16001]_ ;
  assign \new_[16003]_  = \new_[16002]_  & \new_[15997]_ ;
  assign \new_[16007]_  = A269 & ~A266;
  assign \new_[16008]_  = A265 & \new_[16007]_ ;
  assign \new_[16012]_  = ~A301 & ~A299;
  assign \new_[16013]_  = ~A298 & \new_[16012]_ ;
  assign \new_[16014]_  = \new_[16013]_  & \new_[16008]_ ;
  assign \new_[16018]_  = ~A166 & A167;
  assign \new_[16019]_  = A170 & \new_[16018]_ ;
  assign \new_[16023]_  = A203 & ~A200;
  assign \new_[16024]_  = A199 & \new_[16023]_ ;
  assign \new_[16025]_  = \new_[16024]_  & \new_[16019]_ ;
  assign \new_[16029]_  = A298 & A267;
  assign \new_[16030]_  = A265 & \new_[16029]_ ;
  assign \new_[16034]_  = ~A301 & ~A300;
  assign \new_[16035]_  = A299 & \new_[16034]_ ;
  assign \new_[16036]_  = \new_[16035]_  & \new_[16030]_ ;
  assign \new_[16040]_  = ~A166 & A167;
  assign \new_[16041]_  = A170 & \new_[16040]_ ;
  assign \new_[16045]_  = A203 & ~A200;
  assign \new_[16046]_  = A199 & \new_[16045]_ ;
  assign \new_[16047]_  = \new_[16046]_  & \new_[16041]_ ;
  assign \new_[16051]_  = A298 & A267;
  assign \new_[16052]_  = A266 & \new_[16051]_ ;
  assign \new_[16056]_  = ~A301 & ~A300;
  assign \new_[16057]_  = A299 & \new_[16056]_ ;
  assign \new_[16058]_  = \new_[16057]_  & \new_[16052]_ ;
  assign \new_[16062]_  = ~A166 & A167;
  assign \new_[16063]_  = A170 & \new_[16062]_ ;
  assign \new_[16067]_  = A203 & ~A200;
  assign \new_[16068]_  = A199 & \new_[16067]_ ;
  assign \new_[16069]_  = \new_[16068]_  & \new_[16063]_ ;
  assign \new_[16073]_  = A269 & A266;
  assign \new_[16074]_  = ~A265 & \new_[16073]_ ;
  assign \new_[16078]_  = ~A302 & ~A301;
  assign \new_[16079]_  = ~A300 & \new_[16078]_ ;
  assign \new_[16080]_  = \new_[16079]_  & \new_[16074]_ ;
  assign \new_[16084]_  = ~A166 & A167;
  assign \new_[16085]_  = A170 & \new_[16084]_ ;
  assign \new_[16089]_  = A203 & ~A200;
  assign \new_[16090]_  = A199 & \new_[16089]_ ;
  assign \new_[16091]_  = \new_[16090]_  & \new_[16085]_ ;
  assign \new_[16095]_  = A269 & A266;
  assign \new_[16096]_  = ~A265 & \new_[16095]_ ;
  assign \new_[16100]_  = ~A301 & ~A299;
  assign \new_[16101]_  = ~A298 & \new_[16100]_ ;
  assign \new_[16102]_  = \new_[16101]_  & \new_[16096]_ ;
  assign \new_[16106]_  = ~A166 & A167;
  assign \new_[16107]_  = A170 & \new_[16106]_ ;
  assign \new_[16111]_  = A203 & ~A200;
  assign \new_[16112]_  = A199 & \new_[16111]_ ;
  assign \new_[16113]_  = \new_[16112]_  & \new_[16107]_ ;
  assign \new_[16117]_  = A269 & ~A266;
  assign \new_[16118]_  = A265 & \new_[16117]_ ;
  assign \new_[16122]_  = ~A302 & ~A301;
  assign \new_[16123]_  = ~A300 & \new_[16122]_ ;
  assign \new_[16124]_  = \new_[16123]_  & \new_[16118]_ ;
  assign \new_[16128]_  = ~A166 & A167;
  assign \new_[16129]_  = A170 & \new_[16128]_ ;
  assign \new_[16133]_  = A203 & ~A200;
  assign \new_[16134]_  = A199 & \new_[16133]_ ;
  assign \new_[16135]_  = \new_[16134]_  & \new_[16129]_ ;
  assign \new_[16139]_  = A269 & ~A266;
  assign \new_[16140]_  = A265 & \new_[16139]_ ;
  assign \new_[16144]_  = ~A301 & ~A299;
  assign \new_[16145]_  = ~A298 & \new_[16144]_ ;
  assign \new_[16146]_  = \new_[16145]_  & \new_[16140]_ ;
  assign \new_[16150]_  = ~A166 & A167;
  assign \new_[16151]_  = A170 & \new_[16150]_ ;
  assign \new_[16155]_  = ~A202 & ~A200;
  assign \new_[16156]_  = ~A199 & \new_[16155]_ ;
  assign \new_[16157]_  = \new_[16156]_  & \new_[16151]_ ;
  assign \new_[16161]_  = ~A269 & ~A268;
  assign \new_[16162]_  = ~A267 & \new_[16161]_ ;
  assign \new_[16166]_  = A302 & ~A299;
  assign \new_[16167]_  = A298 & \new_[16166]_ ;
  assign \new_[16168]_  = \new_[16167]_  & \new_[16162]_ ;
  assign \new_[16172]_  = ~A166 & A167;
  assign \new_[16173]_  = A170 & \new_[16172]_ ;
  assign \new_[16177]_  = ~A202 & ~A200;
  assign \new_[16178]_  = ~A199 & \new_[16177]_ ;
  assign \new_[16179]_  = \new_[16178]_  & \new_[16173]_ ;
  assign \new_[16183]_  = ~A269 & ~A268;
  assign \new_[16184]_  = ~A267 & \new_[16183]_ ;
  assign \new_[16188]_  = A302 & A299;
  assign \new_[16189]_  = ~A298 & \new_[16188]_ ;
  assign \new_[16190]_  = \new_[16189]_  & \new_[16184]_ ;
  assign \new_[16194]_  = ~A166 & A167;
  assign \new_[16195]_  = A170 & \new_[16194]_ ;
  assign \new_[16199]_  = ~A202 & ~A200;
  assign \new_[16200]_  = ~A199 & \new_[16199]_ ;
  assign \new_[16201]_  = \new_[16200]_  & \new_[16195]_ ;
  assign \new_[16205]_  = ~A267 & A266;
  assign \new_[16206]_  = A265 & \new_[16205]_ ;
  assign \new_[16210]_  = A300 & A299;
  assign \new_[16211]_  = ~A268 & \new_[16210]_ ;
  assign \new_[16212]_  = \new_[16211]_  & \new_[16206]_ ;
  assign \new_[16216]_  = ~A166 & A167;
  assign \new_[16217]_  = A170 & \new_[16216]_ ;
  assign \new_[16221]_  = ~A202 & ~A200;
  assign \new_[16222]_  = ~A199 & \new_[16221]_ ;
  assign \new_[16223]_  = \new_[16222]_  & \new_[16217]_ ;
  assign \new_[16227]_  = ~A267 & A266;
  assign \new_[16228]_  = A265 & \new_[16227]_ ;
  assign \new_[16232]_  = A300 & A298;
  assign \new_[16233]_  = ~A268 & \new_[16232]_ ;
  assign \new_[16234]_  = \new_[16233]_  & \new_[16228]_ ;
  assign \new_[16238]_  = ~A166 & A167;
  assign \new_[16239]_  = A170 & \new_[16238]_ ;
  assign \new_[16243]_  = ~A202 & ~A200;
  assign \new_[16244]_  = ~A199 & \new_[16243]_ ;
  assign \new_[16245]_  = \new_[16244]_  & \new_[16239]_ ;
  assign \new_[16249]_  = ~A268 & ~A266;
  assign \new_[16250]_  = ~A265 & \new_[16249]_ ;
  assign \new_[16254]_  = A302 & ~A299;
  assign \new_[16255]_  = A298 & \new_[16254]_ ;
  assign \new_[16256]_  = \new_[16255]_  & \new_[16250]_ ;
  assign \new_[16260]_  = ~A166 & A167;
  assign \new_[16261]_  = A170 & \new_[16260]_ ;
  assign \new_[16265]_  = ~A202 & ~A200;
  assign \new_[16266]_  = ~A199 & \new_[16265]_ ;
  assign \new_[16267]_  = \new_[16266]_  & \new_[16261]_ ;
  assign \new_[16271]_  = ~A268 & ~A266;
  assign \new_[16272]_  = ~A265 & \new_[16271]_ ;
  assign \new_[16276]_  = A302 & A299;
  assign \new_[16277]_  = ~A298 & \new_[16276]_ ;
  assign \new_[16278]_  = \new_[16277]_  & \new_[16272]_ ;
  assign \new_[16282]_  = A166 & ~A167;
  assign \new_[16283]_  = A170 & \new_[16282]_ ;
  assign \new_[16287]_  = ~A203 & ~A202;
  assign \new_[16288]_  = ~A201 & \new_[16287]_ ;
  assign \new_[16289]_  = \new_[16288]_  & \new_[16283]_ ;
  assign \new_[16293]_  = ~A269 & ~A268;
  assign \new_[16294]_  = ~A267 & \new_[16293]_ ;
  assign \new_[16298]_  = A302 & ~A299;
  assign \new_[16299]_  = A298 & \new_[16298]_ ;
  assign \new_[16300]_  = \new_[16299]_  & \new_[16294]_ ;
  assign \new_[16304]_  = A166 & ~A167;
  assign \new_[16305]_  = A170 & \new_[16304]_ ;
  assign \new_[16309]_  = ~A203 & ~A202;
  assign \new_[16310]_  = ~A201 & \new_[16309]_ ;
  assign \new_[16311]_  = \new_[16310]_  & \new_[16305]_ ;
  assign \new_[16315]_  = ~A269 & ~A268;
  assign \new_[16316]_  = ~A267 & \new_[16315]_ ;
  assign \new_[16320]_  = A302 & A299;
  assign \new_[16321]_  = ~A298 & \new_[16320]_ ;
  assign \new_[16322]_  = \new_[16321]_  & \new_[16316]_ ;
  assign \new_[16326]_  = A166 & ~A167;
  assign \new_[16327]_  = A170 & \new_[16326]_ ;
  assign \new_[16331]_  = ~A203 & ~A202;
  assign \new_[16332]_  = ~A201 & \new_[16331]_ ;
  assign \new_[16333]_  = \new_[16332]_  & \new_[16327]_ ;
  assign \new_[16337]_  = ~A267 & A266;
  assign \new_[16338]_  = A265 & \new_[16337]_ ;
  assign \new_[16342]_  = A300 & A299;
  assign \new_[16343]_  = ~A268 & \new_[16342]_ ;
  assign \new_[16344]_  = \new_[16343]_  & \new_[16338]_ ;
  assign \new_[16348]_  = A166 & ~A167;
  assign \new_[16349]_  = A170 & \new_[16348]_ ;
  assign \new_[16353]_  = ~A203 & ~A202;
  assign \new_[16354]_  = ~A201 & \new_[16353]_ ;
  assign \new_[16355]_  = \new_[16354]_  & \new_[16349]_ ;
  assign \new_[16359]_  = ~A267 & A266;
  assign \new_[16360]_  = A265 & \new_[16359]_ ;
  assign \new_[16364]_  = A300 & A298;
  assign \new_[16365]_  = ~A268 & \new_[16364]_ ;
  assign \new_[16366]_  = \new_[16365]_  & \new_[16360]_ ;
  assign \new_[16370]_  = A166 & ~A167;
  assign \new_[16371]_  = A170 & \new_[16370]_ ;
  assign \new_[16375]_  = ~A203 & ~A202;
  assign \new_[16376]_  = ~A201 & \new_[16375]_ ;
  assign \new_[16377]_  = \new_[16376]_  & \new_[16371]_ ;
  assign \new_[16381]_  = ~A268 & ~A266;
  assign \new_[16382]_  = ~A265 & \new_[16381]_ ;
  assign \new_[16386]_  = A302 & ~A299;
  assign \new_[16387]_  = A298 & \new_[16386]_ ;
  assign \new_[16388]_  = \new_[16387]_  & \new_[16382]_ ;
  assign \new_[16392]_  = A166 & ~A167;
  assign \new_[16393]_  = A170 & \new_[16392]_ ;
  assign \new_[16397]_  = ~A203 & ~A202;
  assign \new_[16398]_  = ~A201 & \new_[16397]_ ;
  assign \new_[16399]_  = \new_[16398]_  & \new_[16393]_ ;
  assign \new_[16403]_  = ~A268 & ~A266;
  assign \new_[16404]_  = ~A265 & \new_[16403]_ ;
  assign \new_[16408]_  = A302 & A299;
  assign \new_[16409]_  = ~A298 & \new_[16408]_ ;
  assign \new_[16410]_  = \new_[16409]_  & \new_[16404]_ ;
  assign \new_[16414]_  = A166 & ~A167;
  assign \new_[16415]_  = A170 & \new_[16414]_ ;
  assign \new_[16419]_  = ~A265 & A201;
  assign \new_[16420]_  = A199 & \new_[16419]_ ;
  assign \new_[16421]_  = \new_[16420]_  & \new_[16415]_ ;
  assign \new_[16425]_  = A298 & A269;
  assign \new_[16426]_  = A266 & \new_[16425]_ ;
  assign \new_[16430]_  = ~A301 & ~A300;
  assign \new_[16431]_  = A299 & \new_[16430]_ ;
  assign \new_[16432]_  = \new_[16431]_  & \new_[16426]_ ;
  assign \new_[16436]_  = A166 & ~A167;
  assign \new_[16437]_  = A170 & \new_[16436]_ ;
  assign \new_[16441]_  = A265 & A201;
  assign \new_[16442]_  = A199 & \new_[16441]_ ;
  assign \new_[16443]_  = \new_[16442]_  & \new_[16437]_ ;
  assign \new_[16447]_  = A298 & A269;
  assign \new_[16448]_  = ~A266 & \new_[16447]_ ;
  assign \new_[16452]_  = ~A301 & ~A300;
  assign \new_[16453]_  = A299 & \new_[16452]_ ;
  assign \new_[16454]_  = \new_[16453]_  & \new_[16448]_ ;
  assign \new_[16458]_  = A166 & ~A167;
  assign \new_[16459]_  = A170 & \new_[16458]_ ;
  assign \new_[16463]_  = ~A265 & A201;
  assign \new_[16464]_  = A200 & \new_[16463]_ ;
  assign \new_[16465]_  = \new_[16464]_  & \new_[16459]_ ;
  assign \new_[16469]_  = A298 & A269;
  assign \new_[16470]_  = A266 & \new_[16469]_ ;
  assign \new_[16474]_  = ~A301 & ~A300;
  assign \new_[16475]_  = A299 & \new_[16474]_ ;
  assign \new_[16476]_  = \new_[16475]_  & \new_[16470]_ ;
  assign \new_[16480]_  = A166 & ~A167;
  assign \new_[16481]_  = A170 & \new_[16480]_ ;
  assign \new_[16485]_  = A265 & A201;
  assign \new_[16486]_  = A200 & \new_[16485]_ ;
  assign \new_[16487]_  = \new_[16486]_  & \new_[16481]_ ;
  assign \new_[16491]_  = A298 & A269;
  assign \new_[16492]_  = ~A266 & \new_[16491]_ ;
  assign \new_[16496]_  = ~A301 & ~A300;
  assign \new_[16497]_  = A299 & \new_[16496]_ ;
  assign \new_[16498]_  = \new_[16497]_  & \new_[16492]_ ;
  assign \new_[16502]_  = A166 & ~A167;
  assign \new_[16503]_  = A170 & \new_[16502]_ ;
  assign \new_[16507]_  = ~A201 & A200;
  assign \new_[16508]_  = A199 & \new_[16507]_ ;
  assign \new_[16509]_  = \new_[16508]_  & \new_[16503]_ ;
  assign \new_[16513]_  = ~A268 & ~A267;
  assign \new_[16514]_  = ~A202 & \new_[16513]_ ;
  assign \new_[16518]_  = A300 & A299;
  assign \new_[16519]_  = ~A269 & \new_[16518]_ ;
  assign \new_[16520]_  = \new_[16519]_  & \new_[16514]_ ;
  assign \new_[16524]_  = A166 & ~A167;
  assign \new_[16525]_  = A170 & \new_[16524]_ ;
  assign \new_[16529]_  = ~A201 & A200;
  assign \new_[16530]_  = A199 & \new_[16529]_ ;
  assign \new_[16531]_  = \new_[16530]_  & \new_[16525]_ ;
  assign \new_[16535]_  = ~A268 & ~A267;
  assign \new_[16536]_  = ~A202 & \new_[16535]_ ;
  assign \new_[16540]_  = A300 & A298;
  assign \new_[16541]_  = ~A269 & \new_[16540]_ ;
  assign \new_[16542]_  = \new_[16541]_  & \new_[16536]_ ;
  assign \new_[16546]_  = A166 & ~A167;
  assign \new_[16547]_  = A170 & \new_[16546]_ ;
  assign \new_[16551]_  = ~A201 & A200;
  assign \new_[16552]_  = A199 & \new_[16551]_ ;
  assign \new_[16553]_  = \new_[16552]_  & \new_[16547]_ ;
  assign \new_[16557]_  = A266 & A265;
  assign \new_[16558]_  = ~A202 & \new_[16557]_ ;
  assign \new_[16562]_  = A301 & ~A268;
  assign \new_[16563]_  = ~A267 & \new_[16562]_ ;
  assign \new_[16564]_  = \new_[16563]_  & \new_[16558]_ ;
  assign \new_[16568]_  = A166 & ~A167;
  assign \new_[16569]_  = A170 & \new_[16568]_ ;
  assign \new_[16573]_  = ~A201 & A200;
  assign \new_[16574]_  = A199 & \new_[16573]_ ;
  assign \new_[16575]_  = \new_[16574]_  & \new_[16569]_ ;
  assign \new_[16579]_  = ~A266 & ~A265;
  assign \new_[16580]_  = ~A202 & \new_[16579]_ ;
  assign \new_[16584]_  = A300 & A299;
  assign \new_[16585]_  = ~A268 & \new_[16584]_ ;
  assign \new_[16586]_  = \new_[16585]_  & \new_[16580]_ ;
  assign \new_[16590]_  = A166 & ~A167;
  assign \new_[16591]_  = A170 & \new_[16590]_ ;
  assign \new_[16595]_  = ~A201 & A200;
  assign \new_[16596]_  = A199 & \new_[16595]_ ;
  assign \new_[16597]_  = \new_[16596]_  & \new_[16591]_ ;
  assign \new_[16601]_  = ~A266 & ~A265;
  assign \new_[16602]_  = ~A202 & \new_[16601]_ ;
  assign \new_[16606]_  = A300 & A298;
  assign \new_[16607]_  = ~A268 & \new_[16606]_ ;
  assign \new_[16608]_  = \new_[16607]_  & \new_[16602]_ ;
  assign \new_[16612]_  = A166 & ~A167;
  assign \new_[16613]_  = A170 & \new_[16612]_ ;
  assign \new_[16617]_  = A203 & A200;
  assign \new_[16618]_  = ~A199 & \new_[16617]_ ;
  assign \new_[16619]_  = \new_[16618]_  & \new_[16613]_ ;
  assign \new_[16623]_  = A298 & A267;
  assign \new_[16624]_  = A265 & \new_[16623]_ ;
  assign \new_[16628]_  = ~A301 & ~A300;
  assign \new_[16629]_  = A299 & \new_[16628]_ ;
  assign \new_[16630]_  = \new_[16629]_  & \new_[16624]_ ;
  assign \new_[16634]_  = A166 & ~A167;
  assign \new_[16635]_  = A170 & \new_[16634]_ ;
  assign \new_[16639]_  = A203 & A200;
  assign \new_[16640]_  = ~A199 & \new_[16639]_ ;
  assign \new_[16641]_  = \new_[16640]_  & \new_[16635]_ ;
  assign \new_[16645]_  = A298 & A267;
  assign \new_[16646]_  = A266 & \new_[16645]_ ;
  assign \new_[16650]_  = ~A301 & ~A300;
  assign \new_[16651]_  = A299 & \new_[16650]_ ;
  assign \new_[16652]_  = \new_[16651]_  & \new_[16646]_ ;
  assign \new_[16656]_  = A166 & ~A167;
  assign \new_[16657]_  = A170 & \new_[16656]_ ;
  assign \new_[16661]_  = A203 & A200;
  assign \new_[16662]_  = ~A199 & \new_[16661]_ ;
  assign \new_[16663]_  = \new_[16662]_  & \new_[16657]_ ;
  assign \new_[16667]_  = A269 & A266;
  assign \new_[16668]_  = ~A265 & \new_[16667]_ ;
  assign \new_[16672]_  = ~A302 & ~A301;
  assign \new_[16673]_  = ~A300 & \new_[16672]_ ;
  assign \new_[16674]_  = \new_[16673]_  & \new_[16668]_ ;
  assign \new_[16678]_  = A166 & ~A167;
  assign \new_[16679]_  = A170 & \new_[16678]_ ;
  assign \new_[16683]_  = A203 & A200;
  assign \new_[16684]_  = ~A199 & \new_[16683]_ ;
  assign \new_[16685]_  = \new_[16684]_  & \new_[16679]_ ;
  assign \new_[16689]_  = A269 & A266;
  assign \new_[16690]_  = ~A265 & \new_[16689]_ ;
  assign \new_[16694]_  = ~A301 & ~A299;
  assign \new_[16695]_  = ~A298 & \new_[16694]_ ;
  assign \new_[16696]_  = \new_[16695]_  & \new_[16690]_ ;
  assign \new_[16700]_  = A166 & ~A167;
  assign \new_[16701]_  = A170 & \new_[16700]_ ;
  assign \new_[16705]_  = A203 & A200;
  assign \new_[16706]_  = ~A199 & \new_[16705]_ ;
  assign \new_[16707]_  = \new_[16706]_  & \new_[16701]_ ;
  assign \new_[16711]_  = A269 & ~A266;
  assign \new_[16712]_  = A265 & \new_[16711]_ ;
  assign \new_[16716]_  = ~A302 & ~A301;
  assign \new_[16717]_  = ~A300 & \new_[16716]_ ;
  assign \new_[16718]_  = \new_[16717]_  & \new_[16712]_ ;
  assign \new_[16722]_  = A166 & ~A167;
  assign \new_[16723]_  = A170 & \new_[16722]_ ;
  assign \new_[16727]_  = A203 & A200;
  assign \new_[16728]_  = ~A199 & \new_[16727]_ ;
  assign \new_[16729]_  = \new_[16728]_  & \new_[16723]_ ;
  assign \new_[16733]_  = A269 & ~A266;
  assign \new_[16734]_  = A265 & \new_[16733]_ ;
  assign \new_[16738]_  = ~A301 & ~A299;
  assign \new_[16739]_  = ~A298 & \new_[16738]_ ;
  assign \new_[16740]_  = \new_[16739]_  & \new_[16734]_ ;
  assign \new_[16744]_  = A166 & ~A167;
  assign \new_[16745]_  = A170 & \new_[16744]_ ;
  assign \new_[16749]_  = A203 & ~A200;
  assign \new_[16750]_  = A199 & \new_[16749]_ ;
  assign \new_[16751]_  = \new_[16750]_  & \new_[16745]_ ;
  assign \new_[16755]_  = A298 & A267;
  assign \new_[16756]_  = A265 & \new_[16755]_ ;
  assign \new_[16760]_  = ~A301 & ~A300;
  assign \new_[16761]_  = A299 & \new_[16760]_ ;
  assign \new_[16762]_  = \new_[16761]_  & \new_[16756]_ ;
  assign \new_[16766]_  = A166 & ~A167;
  assign \new_[16767]_  = A170 & \new_[16766]_ ;
  assign \new_[16771]_  = A203 & ~A200;
  assign \new_[16772]_  = A199 & \new_[16771]_ ;
  assign \new_[16773]_  = \new_[16772]_  & \new_[16767]_ ;
  assign \new_[16777]_  = A298 & A267;
  assign \new_[16778]_  = A266 & \new_[16777]_ ;
  assign \new_[16782]_  = ~A301 & ~A300;
  assign \new_[16783]_  = A299 & \new_[16782]_ ;
  assign \new_[16784]_  = \new_[16783]_  & \new_[16778]_ ;
  assign \new_[16788]_  = A166 & ~A167;
  assign \new_[16789]_  = A170 & \new_[16788]_ ;
  assign \new_[16793]_  = A203 & ~A200;
  assign \new_[16794]_  = A199 & \new_[16793]_ ;
  assign \new_[16795]_  = \new_[16794]_  & \new_[16789]_ ;
  assign \new_[16799]_  = A269 & A266;
  assign \new_[16800]_  = ~A265 & \new_[16799]_ ;
  assign \new_[16804]_  = ~A302 & ~A301;
  assign \new_[16805]_  = ~A300 & \new_[16804]_ ;
  assign \new_[16806]_  = \new_[16805]_  & \new_[16800]_ ;
  assign \new_[16810]_  = A166 & ~A167;
  assign \new_[16811]_  = A170 & \new_[16810]_ ;
  assign \new_[16815]_  = A203 & ~A200;
  assign \new_[16816]_  = A199 & \new_[16815]_ ;
  assign \new_[16817]_  = \new_[16816]_  & \new_[16811]_ ;
  assign \new_[16821]_  = A269 & A266;
  assign \new_[16822]_  = ~A265 & \new_[16821]_ ;
  assign \new_[16826]_  = ~A301 & ~A299;
  assign \new_[16827]_  = ~A298 & \new_[16826]_ ;
  assign \new_[16828]_  = \new_[16827]_  & \new_[16822]_ ;
  assign \new_[16832]_  = A166 & ~A167;
  assign \new_[16833]_  = A170 & \new_[16832]_ ;
  assign \new_[16837]_  = A203 & ~A200;
  assign \new_[16838]_  = A199 & \new_[16837]_ ;
  assign \new_[16839]_  = \new_[16838]_  & \new_[16833]_ ;
  assign \new_[16843]_  = A269 & ~A266;
  assign \new_[16844]_  = A265 & \new_[16843]_ ;
  assign \new_[16848]_  = ~A302 & ~A301;
  assign \new_[16849]_  = ~A300 & \new_[16848]_ ;
  assign \new_[16850]_  = \new_[16849]_  & \new_[16844]_ ;
  assign \new_[16854]_  = A166 & ~A167;
  assign \new_[16855]_  = A170 & \new_[16854]_ ;
  assign \new_[16859]_  = A203 & ~A200;
  assign \new_[16860]_  = A199 & \new_[16859]_ ;
  assign \new_[16861]_  = \new_[16860]_  & \new_[16855]_ ;
  assign \new_[16865]_  = A269 & ~A266;
  assign \new_[16866]_  = A265 & \new_[16865]_ ;
  assign \new_[16870]_  = ~A301 & ~A299;
  assign \new_[16871]_  = ~A298 & \new_[16870]_ ;
  assign \new_[16872]_  = \new_[16871]_  & \new_[16866]_ ;
  assign \new_[16876]_  = A166 & ~A167;
  assign \new_[16877]_  = A170 & \new_[16876]_ ;
  assign \new_[16881]_  = ~A202 & ~A200;
  assign \new_[16882]_  = ~A199 & \new_[16881]_ ;
  assign \new_[16883]_  = \new_[16882]_  & \new_[16877]_ ;
  assign \new_[16887]_  = ~A269 & ~A268;
  assign \new_[16888]_  = ~A267 & \new_[16887]_ ;
  assign \new_[16892]_  = A302 & ~A299;
  assign \new_[16893]_  = A298 & \new_[16892]_ ;
  assign \new_[16894]_  = \new_[16893]_  & \new_[16888]_ ;
  assign \new_[16898]_  = A166 & ~A167;
  assign \new_[16899]_  = A170 & \new_[16898]_ ;
  assign \new_[16903]_  = ~A202 & ~A200;
  assign \new_[16904]_  = ~A199 & \new_[16903]_ ;
  assign \new_[16905]_  = \new_[16904]_  & \new_[16899]_ ;
  assign \new_[16909]_  = ~A269 & ~A268;
  assign \new_[16910]_  = ~A267 & \new_[16909]_ ;
  assign \new_[16914]_  = A302 & A299;
  assign \new_[16915]_  = ~A298 & \new_[16914]_ ;
  assign \new_[16916]_  = \new_[16915]_  & \new_[16910]_ ;
  assign \new_[16920]_  = A166 & ~A167;
  assign \new_[16921]_  = A170 & \new_[16920]_ ;
  assign \new_[16925]_  = ~A202 & ~A200;
  assign \new_[16926]_  = ~A199 & \new_[16925]_ ;
  assign \new_[16927]_  = \new_[16926]_  & \new_[16921]_ ;
  assign \new_[16931]_  = ~A267 & A266;
  assign \new_[16932]_  = A265 & \new_[16931]_ ;
  assign \new_[16936]_  = A300 & A299;
  assign \new_[16937]_  = ~A268 & \new_[16936]_ ;
  assign \new_[16938]_  = \new_[16937]_  & \new_[16932]_ ;
  assign \new_[16942]_  = A166 & ~A167;
  assign \new_[16943]_  = A170 & \new_[16942]_ ;
  assign \new_[16947]_  = ~A202 & ~A200;
  assign \new_[16948]_  = ~A199 & \new_[16947]_ ;
  assign \new_[16949]_  = \new_[16948]_  & \new_[16943]_ ;
  assign \new_[16953]_  = ~A267 & A266;
  assign \new_[16954]_  = A265 & \new_[16953]_ ;
  assign \new_[16958]_  = A300 & A298;
  assign \new_[16959]_  = ~A268 & \new_[16958]_ ;
  assign \new_[16960]_  = \new_[16959]_  & \new_[16954]_ ;
  assign \new_[16964]_  = A166 & ~A167;
  assign \new_[16965]_  = A170 & \new_[16964]_ ;
  assign \new_[16969]_  = ~A202 & ~A200;
  assign \new_[16970]_  = ~A199 & \new_[16969]_ ;
  assign \new_[16971]_  = \new_[16970]_  & \new_[16965]_ ;
  assign \new_[16975]_  = ~A268 & ~A266;
  assign \new_[16976]_  = ~A265 & \new_[16975]_ ;
  assign \new_[16980]_  = A302 & ~A299;
  assign \new_[16981]_  = A298 & \new_[16980]_ ;
  assign \new_[16982]_  = \new_[16981]_  & \new_[16976]_ ;
  assign \new_[16986]_  = A166 & ~A167;
  assign \new_[16987]_  = A170 & \new_[16986]_ ;
  assign \new_[16991]_  = ~A202 & ~A200;
  assign \new_[16992]_  = ~A199 & \new_[16991]_ ;
  assign \new_[16993]_  = \new_[16992]_  & \new_[16987]_ ;
  assign \new_[16997]_  = ~A268 & ~A266;
  assign \new_[16998]_  = ~A265 & \new_[16997]_ ;
  assign \new_[17002]_  = A302 & A299;
  assign \new_[17003]_  = ~A298 & \new_[17002]_ ;
  assign \new_[17004]_  = \new_[17003]_  & \new_[16998]_ ;
  assign \new_[17008]_  = A200 & A199;
  assign \new_[17009]_  = A169 & \new_[17008]_ ;
  assign \new_[17013]_  = A265 & ~A202;
  assign \new_[17014]_  = ~A201 & \new_[17013]_ ;
  assign \new_[17015]_  = \new_[17014]_  & \new_[17009]_ ;
  assign \new_[17019]_  = ~A268 & ~A267;
  assign \new_[17020]_  = A266 & \new_[17019]_ ;
  assign \new_[17024]_  = A302 & ~A299;
  assign \new_[17025]_  = A298 & \new_[17024]_ ;
  assign \new_[17026]_  = \new_[17025]_  & \new_[17020]_ ;
  assign \new_[17030]_  = A200 & A199;
  assign \new_[17031]_  = A169 & \new_[17030]_ ;
  assign \new_[17035]_  = A265 & ~A202;
  assign \new_[17036]_  = ~A201 & \new_[17035]_ ;
  assign \new_[17037]_  = \new_[17036]_  & \new_[17031]_ ;
  assign \new_[17041]_  = ~A268 & ~A267;
  assign \new_[17042]_  = A266 & \new_[17041]_ ;
  assign \new_[17046]_  = A302 & A299;
  assign \new_[17047]_  = ~A298 & \new_[17046]_ ;
  assign \new_[17048]_  = \new_[17047]_  & \new_[17042]_ ;
  assign \new_[17052]_  = ~A166 & ~A167;
  assign \new_[17053]_  = ~A169 & \new_[17052]_ ;
  assign \new_[17057]_  = ~A203 & ~A202;
  assign \new_[17058]_  = ~A201 & \new_[17057]_ ;
  assign \new_[17059]_  = \new_[17058]_  & \new_[17053]_ ;
  assign \new_[17063]_  = A298 & A267;
  assign \new_[17064]_  = A265 & \new_[17063]_ ;
  assign \new_[17068]_  = ~A301 & ~A300;
  assign \new_[17069]_  = A299 & \new_[17068]_ ;
  assign \new_[17070]_  = \new_[17069]_  & \new_[17064]_ ;
  assign \new_[17074]_  = ~A166 & ~A167;
  assign \new_[17075]_  = ~A169 & \new_[17074]_ ;
  assign \new_[17079]_  = ~A203 & ~A202;
  assign \new_[17080]_  = ~A201 & \new_[17079]_ ;
  assign \new_[17081]_  = \new_[17080]_  & \new_[17075]_ ;
  assign \new_[17085]_  = A298 & A267;
  assign \new_[17086]_  = A266 & \new_[17085]_ ;
  assign \new_[17090]_  = ~A301 & ~A300;
  assign \new_[17091]_  = A299 & \new_[17090]_ ;
  assign \new_[17092]_  = \new_[17091]_  & \new_[17086]_ ;
  assign \new_[17096]_  = ~A166 & ~A167;
  assign \new_[17097]_  = ~A169 & \new_[17096]_ ;
  assign \new_[17101]_  = ~A203 & ~A202;
  assign \new_[17102]_  = ~A201 & \new_[17101]_ ;
  assign \new_[17103]_  = \new_[17102]_  & \new_[17097]_ ;
  assign \new_[17107]_  = A269 & A266;
  assign \new_[17108]_  = ~A265 & \new_[17107]_ ;
  assign \new_[17112]_  = ~A302 & ~A301;
  assign \new_[17113]_  = ~A300 & \new_[17112]_ ;
  assign \new_[17114]_  = \new_[17113]_  & \new_[17108]_ ;
  assign \new_[17118]_  = ~A166 & ~A167;
  assign \new_[17119]_  = ~A169 & \new_[17118]_ ;
  assign \new_[17123]_  = ~A203 & ~A202;
  assign \new_[17124]_  = ~A201 & \new_[17123]_ ;
  assign \new_[17125]_  = \new_[17124]_  & \new_[17119]_ ;
  assign \new_[17129]_  = A269 & A266;
  assign \new_[17130]_  = ~A265 & \new_[17129]_ ;
  assign \new_[17134]_  = ~A301 & ~A299;
  assign \new_[17135]_  = ~A298 & \new_[17134]_ ;
  assign \new_[17136]_  = \new_[17135]_  & \new_[17130]_ ;
  assign \new_[17140]_  = ~A166 & ~A167;
  assign \new_[17141]_  = ~A169 & \new_[17140]_ ;
  assign \new_[17145]_  = ~A203 & ~A202;
  assign \new_[17146]_  = ~A201 & \new_[17145]_ ;
  assign \new_[17147]_  = \new_[17146]_  & \new_[17141]_ ;
  assign \new_[17151]_  = A269 & ~A266;
  assign \new_[17152]_  = A265 & \new_[17151]_ ;
  assign \new_[17156]_  = ~A302 & ~A301;
  assign \new_[17157]_  = ~A300 & \new_[17156]_ ;
  assign \new_[17158]_  = \new_[17157]_  & \new_[17152]_ ;
  assign \new_[17162]_  = ~A166 & ~A167;
  assign \new_[17163]_  = ~A169 & \new_[17162]_ ;
  assign \new_[17167]_  = ~A203 & ~A202;
  assign \new_[17168]_  = ~A201 & \new_[17167]_ ;
  assign \new_[17169]_  = \new_[17168]_  & \new_[17163]_ ;
  assign \new_[17173]_  = A269 & ~A266;
  assign \new_[17174]_  = A265 & \new_[17173]_ ;
  assign \new_[17178]_  = ~A301 & ~A299;
  assign \new_[17179]_  = ~A298 & \new_[17178]_ ;
  assign \new_[17180]_  = \new_[17179]_  & \new_[17174]_ ;
  assign \new_[17184]_  = ~A166 & ~A167;
  assign \new_[17185]_  = ~A169 & \new_[17184]_ ;
  assign \new_[17189]_  = A265 & A201;
  assign \new_[17190]_  = A199 & \new_[17189]_ ;
  assign \new_[17191]_  = \new_[17190]_  & \new_[17185]_ ;
  assign \new_[17195]_  = ~A268 & ~A267;
  assign \new_[17196]_  = A266 & \new_[17195]_ ;
  assign \new_[17200]_  = A302 & ~A299;
  assign \new_[17201]_  = A298 & \new_[17200]_ ;
  assign \new_[17202]_  = \new_[17201]_  & \new_[17196]_ ;
  assign \new_[17206]_  = ~A166 & ~A167;
  assign \new_[17207]_  = ~A169 & \new_[17206]_ ;
  assign \new_[17211]_  = A265 & A201;
  assign \new_[17212]_  = A199 & \new_[17211]_ ;
  assign \new_[17213]_  = \new_[17212]_  & \new_[17207]_ ;
  assign \new_[17217]_  = ~A268 & ~A267;
  assign \new_[17218]_  = A266 & \new_[17217]_ ;
  assign \new_[17222]_  = A302 & A299;
  assign \new_[17223]_  = ~A298 & \new_[17222]_ ;
  assign \new_[17224]_  = \new_[17223]_  & \new_[17218]_ ;
  assign \new_[17228]_  = ~A166 & ~A167;
  assign \new_[17229]_  = ~A169 & \new_[17228]_ ;
  assign \new_[17233]_  = A265 & A201;
  assign \new_[17234]_  = A200 & \new_[17233]_ ;
  assign \new_[17235]_  = \new_[17234]_  & \new_[17229]_ ;
  assign \new_[17239]_  = ~A268 & ~A267;
  assign \new_[17240]_  = A266 & \new_[17239]_ ;
  assign \new_[17244]_  = A302 & ~A299;
  assign \new_[17245]_  = A298 & \new_[17244]_ ;
  assign \new_[17246]_  = \new_[17245]_  & \new_[17240]_ ;
  assign \new_[17250]_  = ~A166 & ~A167;
  assign \new_[17251]_  = ~A169 & \new_[17250]_ ;
  assign \new_[17255]_  = A265 & A201;
  assign \new_[17256]_  = A200 & \new_[17255]_ ;
  assign \new_[17257]_  = \new_[17256]_  & \new_[17251]_ ;
  assign \new_[17261]_  = ~A268 & ~A267;
  assign \new_[17262]_  = A266 & \new_[17261]_ ;
  assign \new_[17266]_  = A302 & A299;
  assign \new_[17267]_  = ~A298 & \new_[17266]_ ;
  assign \new_[17268]_  = \new_[17267]_  & \new_[17262]_ ;
  assign \new_[17272]_  = ~A166 & ~A167;
  assign \new_[17273]_  = ~A169 & \new_[17272]_ ;
  assign \new_[17277]_  = ~A201 & A200;
  assign \new_[17278]_  = A199 & \new_[17277]_ ;
  assign \new_[17279]_  = \new_[17278]_  & \new_[17273]_ ;
  assign \new_[17283]_  = A298 & A268;
  assign \new_[17284]_  = ~A202 & \new_[17283]_ ;
  assign \new_[17288]_  = ~A301 & ~A300;
  assign \new_[17289]_  = A299 & \new_[17288]_ ;
  assign \new_[17290]_  = \new_[17289]_  & \new_[17284]_ ;
  assign \new_[17294]_  = ~A166 & ~A167;
  assign \new_[17295]_  = ~A169 & \new_[17294]_ ;
  assign \new_[17299]_  = ~A201 & A200;
  assign \new_[17300]_  = A199 & \new_[17299]_ ;
  assign \new_[17301]_  = \new_[17300]_  & \new_[17295]_ ;
  assign \new_[17305]_  = A267 & A265;
  assign \new_[17306]_  = ~A202 & \new_[17305]_ ;
  assign \new_[17310]_  = ~A302 & ~A301;
  assign \new_[17311]_  = ~A300 & \new_[17310]_ ;
  assign \new_[17312]_  = \new_[17311]_  & \new_[17306]_ ;
  assign \new_[17316]_  = ~A166 & ~A167;
  assign \new_[17317]_  = ~A169 & \new_[17316]_ ;
  assign \new_[17321]_  = ~A201 & A200;
  assign \new_[17322]_  = A199 & \new_[17321]_ ;
  assign \new_[17323]_  = \new_[17322]_  & \new_[17317]_ ;
  assign \new_[17327]_  = A267 & A265;
  assign \new_[17328]_  = ~A202 & \new_[17327]_ ;
  assign \new_[17332]_  = ~A301 & ~A299;
  assign \new_[17333]_  = ~A298 & \new_[17332]_ ;
  assign \new_[17334]_  = \new_[17333]_  & \new_[17328]_ ;
  assign \new_[17338]_  = ~A166 & ~A167;
  assign \new_[17339]_  = ~A169 & \new_[17338]_ ;
  assign \new_[17343]_  = ~A201 & A200;
  assign \new_[17344]_  = A199 & \new_[17343]_ ;
  assign \new_[17345]_  = \new_[17344]_  & \new_[17339]_ ;
  assign \new_[17349]_  = A267 & A266;
  assign \new_[17350]_  = ~A202 & \new_[17349]_ ;
  assign \new_[17354]_  = ~A302 & ~A301;
  assign \new_[17355]_  = ~A300 & \new_[17354]_ ;
  assign \new_[17356]_  = \new_[17355]_  & \new_[17350]_ ;
  assign \new_[17360]_  = ~A166 & ~A167;
  assign \new_[17361]_  = ~A169 & \new_[17360]_ ;
  assign \new_[17365]_  = ~A201 & A200;
  assign \new_[17366]_  = A199 & \new_[17365]_ ;
  assign \new_[17367]_  = \new_[17366]_  & \new_[17361]_ ;
  assign \new_[17371]_  = A267 & A266;
  assign \new_[17372]_  = ~A202 & \new_[17371]_ ;
  assign \new_[17376]_  = ~A301 & ~A299;
  assign \new_[17377]_  = ~A298 & \new_[17376]_ ;
  assign \new_[17378]_  = \new_[17377]_  & \new_[17372]_ ;
  assign \new_[17382]_  = ~A166 & ~A167;
  assign \new_[17383]_  = ~A169 & \new_[17382]_ ;
  assign \new_[17387]_  = A203 & A200;
  assign \new_[17388]_  = ~A199 & \new_[17387]_ ;
  assign \new_[17389]_  = \new_[17388]_  & \new_[17383]_ ;
  assign \new_[17393]_  = ~A269 & ~A268;
  assign \new_[17394]_  = ~A267 & \new_[17393]_ ;
  assign \new_[17398]_  = A302 & ~A299;
  assign \new_[17399]_  = A298 & \new_[17398]_ ;
  assign \new_[17400]_  = \new_[17399]_  & \new_[17394]_ ;
  assign \new_[17404]_  = ~A166 & ~A167;
  assign \new_[17405]_  = ~A169 & \new_[17404]_ ;
  assign \new_[17409]_  = A203 & A200;
  assign \new_[17410]_  = ~A199 & \new_[17409]_ ;
  assign \new_[17411]_  = \new_[17410]_  & \new_[17405]_ ;
  assign \new_[17415]_  = ~A269 & ~A268;
  assign \new_[17416]_  = ~A267 & \new_[17415]_ ;
  assign \new_[17420]_  = A302 & A299;
  assign \new_[17421]_  = ~A298 & \new_[17420]_ ;
  assign \new_[17422]_  = \new_[17421]_  & \new_[17416]_ ;
  assign \new_[17426]_  = ~A166 & ~A167;
  assign \new_[17427]_  = ~A169 & \new_[17426]_ ;
  assign \new_[17431]_  = A203 & A200;
  assign \new_[17432]_  = ~A199 & \new_[17431]_ ;
  assign \new_[17433]_  = \new_[17432]_  & \new_[17427]_ ;
  assign \new_[17437]_  = ~A267 & A266;
  assign \new_[17438]_  = A265 & \new_[17437]_ ;
  assign \new_[17442]_  = A300 & A299;
  assign \new_[17443]_  = ~A268 & \new_[17442]_ ;
  assign \new_[17444]_  = \new_[17443]_  & \new_[17438]_ ;
  assign \new_[17448]_  = ~A166 & ~A167;
  assign \new_[17449]_  = ~A169 & \new_[17448]_ ;
  assign \new_[17453]_  = A203 & A200;
  assign \new_[17454]_  = ~A199 & \new_[17453]_ ;
  assign \new_[17455]_  = \new_[17454]_  & \new_[17449]_ ;
  assign \new_[17459]_  = ~A267 & A266;
  assign \new_[17460]_  = A265 & \new_[17459]_ ;
  assign \new_[17464]_  = A300 & A298;
  assign \new_[17465]_  = ~A268 & \new_[17464]_ ;
  assign \new_[17466]_  = \new_[17465]_  & \new_[17460]_ ;
  assign \new_[17470]_  = ~A166 & ~A167;
  assign \new_[17471]_  = ~A169 & \new_[17470]_ ;
  assign \new_[17475]_  = A203 & A200;
  assign \new_[17476]_  = ~A199 & \new_[17475]_ ;
  assign \new_[17477]_  = \new_[17476]_  & \new_[17471]_ ;
  assign \new_[17481]_  = ~A268 & ~A266;
  assign \new_[17482]_  = ~A265 & \new_[17481]_ ;
  assign \new_[17486]_  = A302 & ~A299;
  assign \new_[17487]_  = A298 & \new_[17486]_ ;
  assign \new_[17488]_  = \new_[17487]_  & \new_[17482]_ ;
  assign \new_[17492]_  = ~A166 & ~A167;
  assign \new_[17493]_  = ~A169 & \new_[17492]_ ;
  assign \new_[17497]_  = A203 & A200;
  assign \new_[17498]_  = ~A199 & \new_[17497]_ ;
  assign \new_[17499]_  = \new_[17498]_  & \new_[17493]_ ;
  assign \new_[17503]_  = ~A268 & ~A266;
  assign \new_[17504]_  = ~A265 & \new_[17503]_ ;
  assign \new_[17508]_  = A302 & A299;
  assign \new_[17509]_  = ~A298 & \new_[17508]_ ;
  assign \new_[17510]_  = \new_[17509]_  & \new_[17504]_ ;
  assign \new_[17514]_  = ~A166 & ~A167;
  assign \new_[17515]_  = ~A169 & \new_[17514]_ ;
  assign \new_[17519]_  = A203 & ~A200;
  assign \new_[17520]_  = A199 & \new_[17519]_ ;
  assign \new_[17521]_  = \new_[17520]_  & \new_[17515]_ ;
  assign \new_[17525]_  = ~A269 & ~A268;
  assign \new_[17526]_  = ~A267 & \new_[17525]_ ;
  assign \new_[17530]_  = A302 & ~A299;
  assign \new_[17531]_  = A298 & \new_[17530]_ ;
  assign \new_[17532]_  = \new_[17531]_  & \new_[17526]_ ;
  assign \new_[17536]_  = ~A166 & ~A167;
  assign \new_[17537]_  = ~A169 & \new_[17536]_ ;
  assign \new_[17541]_  = A203 & ~A200;
  assign \new_[17542]_  = A199 & \new_[17541]_ ;
  assign \new_[17543]_  = \new_[17542]_  & \new_[17537]_ ;
  assign \new_[17547]_  = ~A269 & ~A268;
  assign \new_[17548]_  = ~A267 & \new_[17547]_ ;
  assign \new_[17552]_  = A302 & A299;
  assign \new_[17553]_  = ~A298 & \new_[17552]_ ;
  assign \new_[17554]_  = \new_[17553]_  & \new_[17548]_ ;
  assign \new_[17558]_  = ~A166 & ~A167;
  assign \new_[17559]_  = ~A169 & \new_[17558]_ ;
  assign \new_[17563]_  = A203 & ~A200;
  assign \new_[17564]_  = A199 & \new_[17563]_ ;
  assign \new_[17565]_  = \new_[17564]_  & \new_[17559]_ ;
  assign \new_[17569]_  = ~A267 & A266;
  assign \new_[17570]_  = A265 & \new_[17569]_ ;
  assign \new_[17574]_  = A300 & A299;
  assign \new_[17575]_  = ~A268 & \new_[17574]_ ;
  assign \new_[17576]_  = \new_[17575]_  & \new_[17570]_ ;
  assign \new_[17580]_  = ~A166 & ~A167;
  assign \new_[17581]_  = ~A169 & \new_[17580]_ ;
  assign \new_[17585]_  = A203 & ~A200;
  assign \new_[17586]_  = A199 & \new_[17585]_ ;
  assign \new_[17587]_  = \new_[17586]_  & \new_[17581]_ ;
  assign \new_[17591]_  = ~A267 & A266;
  assign \new_[17592]_  = A265 & \new_[17591]_ ;
  assign \new_[17596]_  = A300 & A298;
  assign \new_[17597]_  = ~A268 & \new_[17596]_ ;
  assign \new_[17598]_  = \new_[17597]_  & \new_[17592]_ ;
  assign \new_[17602]_  = ~A166 & ~A167;
  assign \new_[17603]_  = ~A169 & \new_[17602]_ ;
  assign \new_[17607]_  = A203 & ~A200;
  assign \new_[17608]_  = A199 & \new_[17607]_ ;
  assign \new_[17609]_  = \new_[17608]_  & \new_[17603]_ ;
  assign \new_[17613]_  = ~A268 & ~A266;
  assign \new_[17614]_  = ~A265 & \new_[17613]_ ;
  assign \new_[17618]_  = A302 & ~A299;
  assign \new_[17619]_  = A298 & \new_[17618]_ ;
  assign \new_[17620]_  = \new_[17619]_  & \new_[17614]_ ;
  assign \new_[17624]_  = ~A166 & ~A167;
  assign \new_[17625]_  = ~A169 & \new_[17624]_ ;
  assign \new_[17629]_  = A203 & ~A200;
  assign \new_[17630]_  = A199 & \new_[17629]_ ;
  assign \new_[17631]_  = \new_[17630]_  & \new_[17625]_ ;
  assign \new_[17635]_  = ~A268 & ~A266;
  assign \new_[17636]_  = ~A265 & \new_[17635]_ ;
  assign \new_[17640]_  = A302 & A299;
  assign \new_[17641]_  = ~A298 & \new_[17640]_ ;
  assign \new_[17642]_  = \new_[17641]_  & \new_[17636]_ ;
  assign \new_[17646]_  = ~A166 & ~A167;
  assign \new_[17647]_  = ~A169 & \new_[17646]_ ;
  assign \new_[17651]_  = ~A202 & ~A200;
  assign \new_[17652]_  = ~A199 & \new_[17651]_ ;
  assign \new_[17653]_  = \new_[17652]_  & \new_[17647]_ ;
  assign \new_[17657]_  = A298 & A267;
  assign \new_[17658]_  = A265 & \new_[17657]_ ;
  assign \new_[17662]_  = ~A301 & ~A300;
  assign \new_[17663]_  = A299 & \new_[17662]_ ;
  assign \new_[17664]_  = \new_[17663]_  & \new_[17658]_ ;
  assign \new_[17668]_  = ~A166 & ~A167;
  assign \new_[17669]_  = ~A169 & \new_[17668]_ ;
  assign \new_[17673]_  = ~A202 & ~A200;
  assign \new_[17674]_  = ~A199 & \new_[17673]_ ;
  assign \new_[17675]_  = \new_[17674]_  & \new_[17669]_ ;
  assign \new_[17679]_  = A298 & A267;
  assign \new_[17680]_  = A266 & \new_[17679]_ ;
  assign \new_[17684]_  = ~A301 & ~A300;
  assign \new_[17685]_  = A299 & \new_[17684]_ ;
  assign \new_[17686]_  = \new_[17685]_  & \new_[17680]_ ;
  assign \new_[17690]_  = ~A166 & ~A167;
  assign \new_[17691]_  = ~A169 & \new_[17690]_ ;
  assign \new_[17695]_  = ~A202 & ~A200;
  assign \new_[17696]_  = ~A199 & \new_[17695]_ ;
  assign \new_[17697]_  = \new_[17696]_  & \new_[17691]_ ;
  assign \new_[17701]_  = A269 & A266;
  assign \new_[17702]_  = ~A265 & \new_[17701]_ ;
  assign \new_[17706]_  = ~A302 & ~A301;
  assign \new_[17707]_  = ~A300 & \new_[17706]_ ;
  assign \new_[17708]_  = \new_[17707]_  & \new_[17702]_ ;
  assign \new_[17712]_  = ~A166 & ~A167;
  assign \new_[17713]_  = ~A169 & \new_[17712]_ ;
  assign \new_[17717]_  = ~A202 & ~A200;
  assign \new_[17718]_  = ~A199 & \new_[17717]_ ;
  assign \new_[17719]_  = \new_[17718]_  & \new_[17713]_ ;
  assign \new_[17723]_  = A269 & A266;
  assign \new_[17724]_  = ~A265 & \new_[17723]_ ;
  assign \new_[17728]_  = ~A301 & ~A299;
  assign \new_[17729]_  = ~A298 & \new_[17728]_ ;
  assign \new_[17730]_  = \new_[17729]_  & \new_[17724]_ ;
  assign \new_[17734]_  = ~A166 & ~A167;
  assign \new_[17735]_  = ~A169 & \new_[17734]_ ;
  assign \new_[17739]_  = ~A202 & ~A200;
  assign \new_[17740]_  = ~A199 & \new_[17739]_ ;
  assign \new_[17741]_  = \new_[17740]_  & \new_[17735]_ ;
  assign \new_[17745]_  = A269 & ~A266;
  assign \new_[17746]_  = A265 & \new_[17745]_ ;
  assign \new_[17750]_  = ~A302 & ~A301;
  assign \new_[17751]_  = ~A300 & \new_[17750]_ ;
  assign \new_[17752]_  = \new_[17751]_  & \new_[17746]_ ;
  assign \new_[17756]_  = ~A166 & ~A167;
  assign \new_[17757]_  = ~A169 & \new_[17756]_ ;
  assign \new_[17761]_  = ~A202 & ~A200;
  assign \new_[17762]_  = ~A199 & \new_[17761]_ ;
  assign \new_[17763]_  = \new_[17762]_  & \new_[17757]_ ;
  assign \new_[17767]_  = A269 & ~A266;
  assign \new_[17768]_  = A265 & \new_[17767]_ ;
  assign \new_[17772]_  = ~A301 & ~A299;
  assign \new_[17773]_  = ~A298 & \new_[17772]_ ;
  assign \new_[17774]_  = \new_[17773]_  & \new_[17768]_ ;
  assign \new_[17778]_  = A167 & ~A168;
  assign \new_[17779]_  = ~A169 & \new_[17778]_ ;
  assign \new_[17783]_  = A265 & A202;
  assign \new_[17784]_  = A166 & \new_[17783]_ ;
  assign \new_[17785]_  = \new_[17784]_  & \new_[17779]_ ;
  assign \new_[17789]_  = ~A268 & ~A267;
  assign \new_[17790]_  = A266 & \new_[17789]_ ;
  assign \new_[17794]_  = A302 & ~A299;
  assign \new_[17795]_  = A298 & \new_[17794]_ ;
  assign \new_[17796]_  = \new_[17795]_  & \new_[17790]_ ;
  assign \new_[17800]_  = A167 & ~A168;
  assign \new_[17801]_  = ~A169 & \new_[17800]_ ;
  assign \new_[17805]_  = A265 & A202;
  assign \new_[17806]_  = A166 & \new_[17805]_ ;
  assign \new_[17807]_  = \new_[17806]_  & \new_[17801]_ ;
  assign \new_[17811]_  = ~A268 & ~A267;
  assign \new_[17812]_  = A266 & \new_[17811]_ ;
  assign \new_[17816]_  = A302 & A299;
  assign \new_[17817]_  = ~A298 & \new_[17816]_ ;
  assign \new_[17818]_  = \new_[17817]_  & \new_[17812]_ ;
  assign \new_[17822]_  = A167 & ~A168;
  assign \new_[17823]_  = ~A169 & \new_[17822]_ ;
  assign \new_[17827]_  = ~A202 & ~A201;
  assign \new_[17828]_  = A166 & \new_[17827]_ ;
  assign \new_[17829]_  = \new_[17828]_  & \new_[17823]_ ;
  assign \new_[17833]_  = A298 & A268;
  assign \new_[17834]_  = ~A203 & \new_[17833]_ ;
  assign \new_[17838]_  = ~A301 & ~A300;
  assign \new_[17839]_  = A299 & \new_[17838]_ ;
  assign \new_[17840]_  = \new_[17839]_  & \new_[17834]_ ;
  assign \new_[17844]_  = A167 & ~A168;
  assign \new_[17845]_  = ~A169 & \new_[17844]_ ;
  assign \new_[17849]_  = ~A202 & ~A201;
  assign \new_[17850]_  = A166 & \new_[17849]_ ;
  assign \new_[17851]_  = \new_[17850]_  & \new_[17845]_ ;
  assign \new_[17855]_  = A267 & A265;
  assign \new_[17856]_  = ~A203 & \new_[17855]_ ;
  assign \new_[17860]_  = ~A302 & ~A301;
  assign \new_[17861]_  = ~A300 & \new_[17860]_ ;
  assign \new_[17862]_  = \new_[17861]_  & \new_[17856]_ ;
  assign \new_[17866]_  = A167 & ~A168;
  assign \new_[17867]_  = ~A169 & \new_[17866]_ ;
  assign \new_[17871]_  = ~A202 & ~A201;
  assign \new_[17872]_  = A166 & \new_[17871]_ ;
  assign \new_[17873]_  = \new_[17872]_  & \new_[17867]_ ;
  assign \new_[17877]_  = A267 & A265;
  assign \new_[17878]_  = ~A203 & \new_[17877]_ ;
  assign \new_[17882]_  = ~A301 & ~A299;
  assign \new_[17883]_  = ~A298 & \new_[17882]_ ;
  assign \new_[17884]_  = \new_[17883]_  & \new_[17878]_ ;
  assign \new_[17888]_  = A167 & ~A168;
  assign \new_[17889]_  = ~A169 & \new_[17888]_ ;
  assign \new_[17893]_  = ~A202 & ~A201;
  assign \new_[17894]_  = A166 & \new_[17893]_ ;
  assign \new_[17895]_  = \new_[17894]_  & \new_[17889]_ ;
  assign \new_[17899]_  = A267 & A266;
  assign \new_[17900]_  = ~A203 & \new_[17899]_ ;
  assign \new_[17904]_  = ~A302 & ~A301;
  assign \new_[17905]_  = ~A300 & \new_[17904]_ ;
  assign \new_[17906]_  = \new_[17905]_  & \new_[17900]_ ;
  assign \new_[17910]_  = A167 & ~A168;
  assign \new_[17911]_  = ~A169 & \new_[17910]_ ;
  assign \new_[17915]_  = ~A202 & ~A201;
  assign \new_[17916]_  = A166 & \new_[17915]_ ;
  assign \new_[17917]_  = \new_[17916]_  & \new_[17911]_ ;
  assign \new_[17921]_  = A267 & A266;
  assign \new_[17922]_  = ~A203 & \new_[17921]_ ;
  assign \new_[17926]_  = ~A301 & ~A299;
  assign \new_[17927]_  = ~A298 & \new_[17926]_ ;
  assign \new_[17928]_  = \new_[17927]_  & \new_[17922]_ ;
  assign \new_[17932]_  = A167 & ~A168;
  assign \new_[17933]_  = ~A169 & \new_[17932]_ ;
  assign \new_[17937]_  = A201 & A199;
  assign \new_[17938]_  = A166 & \new_[17937]_ ;
  assign \new_[17939]_  = \new_[17938]_  & \new_[17933]_ ;
  assign \new_[17943]_  = ~A269 & ~A268;
  assign \new_[17944]_  = ~A267 & \new_[17943]_ ;
  assign \new_[17948]_  = A302 & ~A299;
  assign \new_[17949]_  = A298 & \new_[17948]_ ;
  assign \new_[17950]_  = \new_[17949]_  & \new_[17944]_ ;
  assign \new_[17954]_  = A167 & ~A168;
  assign \new_[17955]_  = ~A169 & \new_[17954]_ ;
  assign \new_[17959]_  = A201 & A199;
  assign \new_[17960]_  = A166 & \new_[17959]_ ;
  assign \new_[17961]_  = \new_[17960]_  & \new_[17955]_ ;
  assign \new_[17965]_  = ~A269 & ~A268;
  assign \new_[17966]_  = ~A267 & \new_[17965]_ ;
  assign \new_[17970]_  = A302 & A299;
  assign \new_[17971]_  = ~A298 & \new_[17970]_ ;
  assign \new_[17972]_  = \new_[17971]_  & \new_[17966]_ ;
  assign \new_[17976]_  = A167 & ~A168;
  assign \new_[17977]_  = ~A169 & \new_[17976]_ ;
  assign \new_[17981]_  = A201 & A199;
  assign \new_[17982]_  = A166 & \new_[17981]_ ;
  assign \new_[17983]_  = \new_[17982]_  & \new_[17977]_ ;
  assign \new_[17987]_  = ~A267 & A266;
  assign \new_[17988]_  = A265 & \new_[17987]_ ;
  assign \new_[17992]_  = A300 & A299;
  assign \new_[17993]_  = ~A268 & \new_[17992]_ ;
  assign \new_[17994]_  = \new_[17993]_  & \new_[17988]_ ;
  assign \new_[17998]_  = A167 & ~A168;
  assign \new_[17999]_  = ~A169 & \new_[17998]_ ;
  assign \new_[18003]_  = A201 & A199;
  assign \new_[18004]_  = A166 & \new_[18003]_ ;
  assign \new_[18005]_  = \new_[18004]_  & \new_[17999]_ ;
  assign \new_[18009]_  = ~A267 & A266;
  assign \new_[18010]_  = A265 & \new_[18009]_ ;
  assign \new_[18014]_  = A300 & A298;
  assign \new_[18015]_  = ~A268 & \new_[18014]_ ;
  assign \new_[18016]_  = \new_[18015]_  & \new_[18010]_ ;
  assign \new_[18020]_  = A167 & ~A168;
  assign \new_[18021]_  = ~A169 & \new_[18020]_ ;
  assign \new_[18025]_  = A201 & A199;
  assign \new_[18026]_  = A166 & \new_[18025]_ ;
  assign \new_[18027]_  = \new_[18026]_  & \new_[18021]_ ;
  assign \new_[18031]_  = ~A268 & ~A266;
  assign \new_[18032]_  = ~A265 & \new_[18031]_ ;
  assign \new_[18036]_  = A302 & ~A299;
  assign \new_[18037]_  = A298 & \new_[18036]_ ;
  assign \new_[18038]_  = \new_[18037]_  & \new_[18032]_ ;
  assign \new_[18042]_  = A167 & ~A168;
  assign \new_[18043]_  = ~A169 & \new_[18042]_ ;
  assign \new_[18047]_  = A201 & A199;
  assign \new_[18048]_  = A166 & \new_[18047]_ ;
  assign \new_[18049]_  = \new_[18048]_  & \new_[18043]_ ;
  assign \new_[18053]_  = ~A268 & ~A266;
  assign \new_[18054]_  = ~A265 & \new_[18053]_ ;
  assign \new_[18058]_  = A302 & A299;
  assign \new_[18059]_  = ~A298 & \new_[18058]_ ;
  assign \new_[18060]_  = \new_[18059]_  & \new_[18054]_ ;
  assign \new_[18064]_  = A167 & ~A168;
  assign \new_[18065]_  = ~A169 & \new_[18064]_ ;
  assign \new_[18069]_  = A201 & A200;
  assign \new_[18070]_  = A166 & \new_[18069]_ ;
  assign \new_[18071]_  = \new_[18070]_  & \new_[18065]_ ;
  assign \new_[18075]_  = ~A269 & ~A268;
  assign \new_[18076]_  = ~A267 & \new_[18075]_ ;
  assign \new_[18080]_  = A302 & ~A299;
  assign \new_[18081]_  = A298 & \new_[18080]_ ;
  assign \new_[18082]_  = \new_[18081]_  & \new_[18076]_ ;
  assign \new_[18086]_  = A167 & ~A168;
  assign \new_[18087]_  = ~A169 & \new_[18086]_ ;
  assign \new_[18091]_  = A201 & A200;
  assign \new_[18092]_  = A166 & \new_[18091]_ ;
  assign \new_[18093]_  = \new_[18092]_  & \new_[18087]_ ;
  assign \new_[18097]_  = ~A269 & ~A268;
  assign \new_[18098]_  = ~A267 & \new_[18097]_ ;
  assign \new_[18102]_  = A302 & A299;
  assign \new_[18103]_  = ~A298 & \new_[18102]_ ;
  assign \new_[18104]_  = \new_[18103]_  & \new_[18098]_ ;
  assign \new_[18108]_  = A167 & ~A168;
  assign \new_[18109]_  = ~A169 & \new_[18108]_ ;
  assign \new_[18113]_  = A201 & A200;
  assign \new_[18114]_  = A166 & \new_[18113]_ ;
  assign \new_[18115]_  = \new_[18114]_  & \new_[18109]_ ;
  assign \new_[18119]_  = ~A267 & A266;
  assign \new_[18120]_  = A265 & \new_[18119]_ ;
  assign \new_[18124]_  = A300 & A299;
  assign \new_[18125]_  = ~A268 & \new_[18124]_ ;
  assign \new_[18126]_  = \new_[18125]_  & \new_[18120]_ ;
  assign \new_[18130]_  = A167 & ~A168;
  assign \new_[18131]_  = ~A169 & \new_[18130]_ ;
  assign \new_[18135]_  = A201 & A200;
  assign \new_[18136]_  = A166 & \new_[18135]_ ;
  assign \new_[18137]_  = \new_[18136]_  & \new_[18131]_ ;
  assign \new_[18141]_  = ~A267 & A266;
  assign \new_[18142]_  = A265 & \new_[18141]_ ;
  assign \new_[18146]_  = A300 & A298;
  assign \new_[18147]_  = ~A268 & \new_[18146]_ ;
  assign \new_[18148]_  = \new_[18147]_  & \new_[18142]_ ;
  assign \new_[18152]_  = A167 & ~A168;
  assign \new_[18153]_  = ~A169 & \new_[18152]_ ;
  assign \new_[18157]_  = A201 & A200;
  assign \new_[18158]_  = A166 & \new_[18157]_ ;
  assign \new_[18159]_  = \new_[18158]_  & \new_[18153]_ ;
  assign \new_[18163]_  = ~A268 & ~A266;
  assign \new_[18164]_  = ~A265 & \new_[18163]_ ;
  assign \new_[18168]_  = A302 & ~A299;
  assign \new_[18169]_  = A298 & \new_[18168]_ ;
  assign \new_[18170]_  = \new_[18169]_  & \new_[18164]_ ;
  assign \new_[18174]_  = A167 & ~A168;
  assign \new_[18175]_  = ~A169 & \new_[18174]_ ;
  assign \new_[18179]_  = A201 & A200;
  assign \new_[18180]_  = A166 & \new_[18179]_ ;
  assign \new_[18181]_  = \new_[18180]_  & \new_[18175]_ ;
  assign \new_[18185]_  = ~A268 & ~A266;
  assign \new_[18186]_  = ~A265 & \new_[18185]_ ;
  assign \new_[18190]_  = A302 & A299;
  assign \new_[18191]_  = ~A298 & \new_[18190]_ ;
  assign \new_[18192]_  = \new_[18191]_  & \new_[18186]_ ;
  assign \new_[18196]_  = A167 & ~A168;
  assign \new_[18197]_  = ~A169 & \new_[18196]_ ;
  assign \new_[18201]_  = A200 & A199;
  assign \new_[18202]_  = A166 & \new_[18201]_ ;
  assign \new_[18203]_  = \new_[18202]_  & \new_[18197]_ ;
  assign \new_[18207]_  = A268 & ~A202;
  assign \new_[18208]_  = ~A201 & \new_[18207]_ ;
  assign \new_[18212]_  = ~A302 & ~A301;
  assign \new_[18213]_  = ~A300 & \new_[18212]_ ;
  assign \new_[18214]_  = \new_[18213]_  & \new_[18208]_ ;
  assign \new_[18218]_  = A167 & ~A168;
  assign \new_[18219]_  = ~A169 & \new_[18218]_ ;
  assign \new_[18223]_  = A200 & A199;
  assign \new_[18224]_  = A166 & \new_[18223]_ ;
  assign \new_[18225]_  = \new_[18224]_  & \new_[18219]_ ;
  assign \new_[18229]_  = A268 & ~A202;
  assign \new_[18230]_  = ~A201 & \new_[18229]_ ;
  assign \new_[18234]_  = ~A301 & ~A299;
  assign \new_[18235]_  = ~A298 & \new_[18234]_ ;
  assign \new_[18236]_  = \new_[18235]_  & \new_[18230]_ ;
  assign \new_[18240]_  = A167 & ~A168;
  assign \new_[18241]_  = ~A169 & \new_[18240]_ ;
  assign \new_[18245]_  = A200 & ~A199;
  assign \new_[18246]_  = A166 & \new_[18245]_ ;
  assign \new_[18247]_  = \new_[18246]_  & \new_[18241]_ ;
  assign \new_[18251]_  = ~A268 & ~A267;
  assign \new_[18252]_  = A203 & \new_[18251]_ ;
  assign \new_[18256]_  = A300 & A299;
  assign \new_[18257]_  = ~A269 & \new_[18256]_ ;
  assign \new_[18258]_  = \new_[18257]_  & \new_[18252]_ ;
  assign \new_[18262]_  = A167 & ~A168;
  assign \new_[18263]_  = ~A169 & \new_[18262]_ ;
  assign \new_[18267]_  = A200 & ~A199;
  assign \new_[18268]_  = A166 & \new_[18267]_ ;
  assign \new_[18269]_  = \new_[18268]_  & \new_[18263]_ ;
  assign \new_[18273]_  = ~A268 & ~A267;
  assign \new_[18274]_  = A203 & \new_[18273]_ ;
  assign \new_[18278]_  = A300 & A298;
  assign \new_[18279]_  = ~A269 & \new_[18278]_ ;
  assign \new_[18280]_  = \new_[18279]_  & \new_[18274]_ ;
  assign \new_[18284]_  = A167 & ~A168;
  assign \new_[18285]_  = ~A169 & \new_[18284]_ ;
  assign \new_[18289]_  = A200 & ~A199;
  assign \new_[18290]_  = A166 & \new_[18289]_ ;
  assign \new_[18291]_  = \new_[18290]_  & \new_[18285]_ ;
  assign \new_[18295]_  = A266 & A265;
  assign \new_[18296]_  = A203 & \new_[18295]_ ;
  assign \new_[18300]_  = A301 & ~A268;
  assign \new_[18301]_  = ~A267 & \new_[18300]_ ;
  assign \new_[18302]_  = \new_[18301]_  & \new_[18296]_ ;
  assign \new_[18306]_  = A167 & ~A168;
  assign \new_[18307]_  = ~A169 & \new_[18306]_ ;
  assign \new_[18311]_  = A200 & ~A199;
  assign \new_[18312]_  = A166 & \new_[18311]_ ;
  assign \new_[18313]_  = \new_[18312]_  & \new_[18307]_ ;
  assign \new_[18317]_  = ~A266 & ~A265;
  assign \new_[18318]_  = A203 & \new_[18317]_ ;
  assign \new_[18322]_  = A300 & A299;
  assign \new_[18323]_  = ~A268 & \new_[18322]_ ;
  assign \new_[18324]_  = \new_[18323]_  & \new_[18318]_ ;
  assign \new_[18328]_  = A167 & ~A168;
  assign \new_[18329]_  = ~A169 & \new_[18328]_ ;
  assign \new_[18333]_  = A200 & ~A199;
  assign \new_[18334]_  = A166 & \new_[18333]_ ;
  assign \new_[18335]_  = \new_[18334]_  & \new_[18329]_ ;
  assign \new_[18339]_  = ~A266 & ~A265;
  assign \new_[18340]_  = A203 & \new_[18339]_ ;
  assign \new_[18344]_  = A300 & A298;
  assign \new_[18345]_  = ~A268 & \new_[18344]_ ;
  assign \new_[18346]_  = \new_[18345]_  & \new_[18340]_ ;
  assign \new_[18350]_  = A167 & ~A168;
  assign \new_[18351]_  = ~A169 & \new_[18350]_ ;
  assign \new_[18355]_  = ~A200 & A199;
  assign \new_[18356]_  = A166 & \new_[18355]_ ;
  assign \new_[18357]_  = \new_[18356]_  & \new_[18351]_ ;
  assign \new_[18361]_  = ~A268 & ~A267;
  assign \new_[18362]_  = A203 & \new_[18361]_ ;
  assign \new_[18366]_  = A300 & A299;
  assign \new_[18367]_  = ~A269 & \new_[18366]_ ;
  assign \new_[18368]_  = \new_[18367]_  & \new_[18362]_ ;
  assign \new_[18372]_  = A167 & ~A168;
  assign \new_[18373]_  = ~A169 & \new_[18372]_ ;
  assign \new_[18377]_  = ~A200 & A199;
  assign \new_[18378]_  = A166 & \new_[18377]_ ;
  assign \new_[18379]_  = \new_[18378]_  & \new_[18373]_ ;
  assign \new_[18383]_  = ~A268 & ~A267;
  assign \new_[18384]_  = A203 & \new_[18383]_ ;
  assign \new_[18388]_  = A300 & A298;
  assign \new_[18389]_  = ~A269 & \new_[18388]_ ;
  assign \new_[18390]_  = \new_[18389]_  & \new_[18384]_ ;
  assign \new_[18394]_  = A167 & ~A168;
  assign \new_[18395]_  = ~A169 & \new_[18394]_ ;
  assign \new_[18399]_  = ~A200 & A199;
  assign \new_[18400]_  = A166 & \new_[18399]_ ;
  assign \new_[18401]_  = \new_[18400]_  & \new_[18395]_ ;
  assign \new_[18405]_  = A266 & A265;
  assign \new_[18406]_  = A203 & \new_[18405]_ ;
  assign \new_[18410]_  = A301 & ~A268;
  assign \new_[18411]_  = ~A267 & \new_[18410]_ ;
  assign \new_[18412]_  = \new_[18411]_  & \new_[18406]_ ;
  assign \new_[18416]_  = A167 & ~A168;
  assign \new_[18417]_  = ~A169 & \new_[18416]_ ;
  assign \new_[18421]_  = ~A200 & A199;
  assign \new_[18422]_  = A166 & \new_[18421]_ ;
  assign \new_[18423]_  = \new_[18422]_  & \new_[18417]_ ;
  assign \new_[18427]_  = ~A266 & ~A265;
  assign \new_[18428]_  = A203 & \new_[18427]_ ;
  assign \new_[18432]_  = A300 & A299;
  assign \new_[18433]_  = ~A268 & \new_[18432]_ ;
  assign \new_[18434]_  = \new_[18433]_  & \new_[18428]_ ;
  assign \new_[18438]_  = A167 & ~A168;
  assign \new_[18439]_  = ~A169 & \new_[18438]_ ;
  assign \new_[18443]_  = ~A200 & A199;
  assign \new_[18444]_  = A166 & \new_[18443]_ ;
  assign \new_[18445]_  = \new_[18444]_  & \new_[18439]_ ;
  assign \new_[18449]_  = ~A266 & ~A265;
  assign \new_[18450]_  = A203 & \new_[18449]_ ;
  assign \new_[18454]_  = A300 & A298;
  assign \new_[18455]_  = ~A268 & \new_[18454]_ ;
  assign \new_[18456]_  = \new_[18455]_  & \new_[18450]_ ;
  assign \new_[18460]_  = A167 & ~A168;
  assign \new_[18461]_  = ~A169 & \new_[18460]_ ;
  assign \new_[18465]_  = ~A200 & ~A199;
  assign \new_[18466]_  = A166 & \new_[18465]_ ;
  assign \new_[18467]_  = \new_[18466]_  & \new_[18461]_ ;
  assign \new_[18471]_  = A298 & A268;
  assign \new_[18472]_  = ~A202 & \new_[18471]_ ;
  assign \new_[18476]_  = ~A301 & ~A300;
  assign \new_[18477]_  = A299 & \new_[18476]_ ;
  assign \new_[18478]_  = \new_[18477]_  & \new_[18472]_ ;
  assign \new_[18482]_  = A167 & ~A168;
  assign \new_[18483]_  = ~A169 & \new_[18482]_ ;
  assign \new_[18487]_  = ~A200 & ~A199;
  assign \new_[18488]_  = A166 & \new_[18487]_ ;
  assign \new_[18489]_  = \new_[18488]_  & \new_[18483]_ ;
  assign \new_[18493]_  = A267 & A265;
  assign \new_[18494]_  = ~A202 & \new_[18493]_ ;
  assign \new_[18498]_  = ~A302 & ~A301;
  assign \new_[18499]_  = ~A300 & \new_[18498]_ ;
  assign \new_[18500]_  = \new_[18499]_  & \new_[18494]_ ;
  assign \new_[18504]_  = A167 & ~A168;
  assign \new_[18505]_  = ~A169 & \new_[18504]_ ;
  assign \new_[18509]_  = ~A200 & ~A199;
  assign \new_[18510]_  = A166 & \new_[18509]_ ;
  assign \new_[18511]_  = \new_[18510]_  & \new_[18505]_ ;
  assign \new_[18515]_  = A267 & A265;
  assign \new_[18516]_  = ~A202 & \new_[18515]_ ;
  assign \new_[18520]_  = ~A301 & ~A299;
  assign \new_[18521]_  = ~A298 & \new_[18520]_ ;
  assign \new_[18522]_  = \new_[18521]_  & \new_[18516]_ ;
  assign \new_[18526]_  = A167 & ~A168;
  assign \new_[18527]_  = ~A169 & \new_[18526]_ ;
  assign \new_[18531]_  = ~A200 & ~A199;
  assign \new_[18532]_  = A166 & \new_[18531]_ ;
  assign \new_[18533]_  = \new_[18532]_  & \new_[18527]_ ;
  assign \new_[18537]_  = A267 & A266;
  assign \new_[18538]_  = ~A202 & \new_[18537]_ ;
  assign \new_[18542]_  = ~A302 & ~A301;
  assign \new_[18543]_  = ~A300 & \new_[18542]_ ;
  assign \new_[18544]_  = \new_[18543]_  & \new_[18538]_ ;
  assign \new_[18548]_  = A167 & ~A168;
  assign \new_[18549]_  = ~A169 & \new_[18548]_ ;
  assign \new_[18553]_  = ~A200 & ~A199;
  assign \new_[18554]_  = A166 & \new_[18553]_ ;
  assign \new_[18555]_  = \new_[18554]_  & \new_[18549]_ ;
  assign \new_[18559]_  = A267 & A266;
  assign \new_[18560]_  = ~A202 & \new_[18559]_ ;
  assign \new_[18564]_  = ~A301 & ~A299;
  assign \new_[18565]_  = ~A298 & \new_[18564]_ ;
  assign \new_[18566]_  = \new_[18565]_  & \new_[18560]_ ;
  assign \new_[18570]_  = ~A168 & ~A169;
  assign \new_[18571]_  = ~A170 & \new_[18570]_ ;
  assign \new_[18575]_  = ~A203 & ~A202;
  assign \new_[18576]_  = ~A201 & \new_[18575]_ ;
  assign \new_[18577]_  = \new_[18576]_  & \new_[18571]_ ;
  assign \new_[18581]_  = A298 & A267;
  assign \new_[18582]_  = A265 & \new_[18581]_ ;
  assign \new_[18586]_  = ~A301 & ~A300;
  assign \new_[18587]_  = A299 & \new_[18586]_ ;
  assign \new_[18588]_  = \new_[18587]_  & \new_[18582]_ ;
  assign \new_[18592]_  = ~A168 & ~A169;
  assign \new_[18593]_  = ~A170 & \new_[18592]_ ;
  assign \new_[18597]_  = ~A203 & ~A202;
  assign \new_[18598]_  = ~A201 & \new_[18597]_ ;
  assign \new_[18599]_  = \new_[18598]_  & \new_[18593]_ ;
  assign \new_[18603]_  = A298 & A267;
  assign \new_[18604]_  = A266 & \new_[18603]_ ;
  assign \new_[18608]_  = ~A301 & ~A300;
  assign \new_[18609]_  = A299 & \new_[18608]_ ;
  assign \new_[18610]_  = \new_[18609]_  & \new_[18604]_ ;
  assign \new_[18614]_  = ~A168 & ~A169;
  assign \new_[18615]_  = ~A170 & \new_[18614]_ ;
  assign \new_[18619]_  = ~A203 & ~A202;
  assign \new_[18620]_  = ~A201 & \new_[18619]_ ;
  assign \new_[18621]_  = \new_[18620]_  & \new_[18615]_ ;
  assign \new_[18625]_  = A269 & A266;
  assign \new_[18626]_  = ~A265 & \new_[18625]_ ;
  assign \new_[18630]_  = ~A302 & ~A301;
  assign \new_[18631]_  = ~A300 & \new_[18630]_ ;
  assign \new_[18632]_  = \new_[18631]_  & \new_[18626]_ ;
  assign \new_[18636]_  = ~A168 & ~A169;
  assign \new_[18637]_  = ~A170 & \new_[18636]_ ;
  assign \new_[18641]_  = ~A203 & ~A202;
  assign \new_[18642]_  = ~A201 & \new_[18641]_ ;
  assign \new_[18643]_  = \new_[18642]_  & \new_[18637]_ ;
  assign \new_[18647]_  = A269 & A266;
  assign \new_[18648]_  = ~A265 & \new_[18647]_ ;
  assign \new_[18652]_  = ~A301 & ~A299;
  assign \new_[18653]_  = ~A298 & \new_[18652]_ ;
  assign \new_[18654]_  = \new_[18653]_  & \new_[18648]_ ;
  assign \new_[18658]_  = ~A168 & ~A169;
  assign \new_[18659]_  = ~A170 & \new_[18658]_ ;
  assign \new_[18663]_  = ~A203 & ~A202;
  assign \new_[18664]_  = ~A201 & \new_[18663]_ ;
  assign \new_[18665]_  = \new_[18664]_  & \new_[18659]_ ;
  assign \new_[18669]_  = A269 & ~A266;
  assign \new_[18670]_  = A265 & \new_[18669]_ ;
  assign \new_[18674]_  = ~A302 & ~A301;
  assign \new_[18675]_  = ~A300 & \new_[18674]_ ;
  assign \new_[18676]_  = \new_[18675]_  & \new_[18670]_ ;
  assign \new_[18680]_  = ~A168 & ~A169;
  assign \new_[18681]_  = ~A170 & \new_[18680]_ ;
  assign \new_[18685]_  = ~A203 & ~A202;
  assign \new_[18686]_  = ~A201 & \new_[18685]_ ;
  assign \new_[18687]_  = \new_[18686]_  & \new_[18681]_ ;
  assign \new_[18691]_  = A269 & ~A266;
  assign \new_[18692]_  = A265 & \new_[18691]_ ;
  assign \new_[18696]_  = ~A301 & ~A299;
  assign \new_[18697]_  = ~A298 & \new_[18696]_ ;
  assign \new_[18698]_  = \new_[18697]_  & \new_[18692]_ ;
  assign \new_[18702]_  = ~A168 & ~A169;
  assign \new_[18703]_  = ~A170 & \new_[18702]_ ;
  assign \new_[18707]_  = A265 & A201;
  assign \new_[18708]_  = A199 & \new_[18707]_ ;
  assign \new_[18709]_  = \new_[18708]_  & \new_[18703]_ ;
  assign \new_[18713]_  = ~A268 & ~A267;
  assign \new_[18714]_  = A266 & \new_[18713]_ ;
  assign \new_[18718]_  = A302 & ~A299;
  assign \new_[18719]_  = A298 & \new_[18718]_ ;
  assign \new_[18720]_  = \new_[18719]_  & \new_[18714]_ ;
  assign \new_[18724]_  = ~A168 & ~A169;
  assign \new_[18725]_  = ~A170 & \new_[18724]_ ;
  assign \new_[18729]_  = A265 & A201;
  assign \new_[18730]_  = A199 & \new_[18729]_ ;
  assign \new_[18731]_  = \new_[18730]_  & \new_[18725]_ ;
  assign \new_[18735]_  = ~A268 & ~A267;
  assign \new_[18736]_  = A266 & \new_[18735]_ ;
  assign \new_[18740]_  = A302 & A299;
  assign \new_[18741]_  = ~A298 & \new_[18740]_ ;
  assign \new_[18742]_  = \new_[18741]_  & \new_[18736]_ ;
  assign \new_[18746]_  = ~A168 & ~A169;
  assign \new_[18747]_  = ~A170 & \new_[18746]_ ;
  assign \new_[18751]_  = A265 & A201;
  assign \new_[18752]_  = A200 & \new_[18751]_ ;
  assign \new_[18753]_  = \new_[18752]_  & \new_[18747]_ ;
  assign \new_[18757]_  = ~A268 & ~A267;
  assign \new_[18758]_  = A266 & \new_[18757]_ ;
  assign \new_[18762]_  = A302 & ~A299;
  assign \new_[18763]_  = A298 & \new_[18762]_ ;
  assign \new_[18764]_  = \new_[18763]_  & \new_[18758]_ ;
  assign \new_[18768]_  = ~A168 & ~A169;
  assign \new_[18769]_  = ~A170 & \new_[18768]_ ;
  assign \new_[18773]_  = A265 & A201;
  assign \new_[18774]_  = A200 & \new_[18773]_ ;
  assign \new_[18775]_  = \new_[18774]_  & \new_[18769]_ ;
  assign \new_[18779]_  = ~A268 & ~A267;
  assign \new_[18780]_  = A266 & \new_[18779]_ ;
  assign \new_[18784]_  = A302 & A299;
  assign \new_[18785]_  = ~A298 & \new_[18784]_ ;
  assign \new_[18786]_  = \new_[18785]_  & \new_[18780]_ ;
  assign \new_[18790]_  = ~A168 & ~A169;
  assign \new_[18791]_  = ~A170 & \new_[18790]_ ;
  assign \new_[18795]_  = ~A201 & A200;
  assign \new_[18796]_  = A199 & \new_[18795]_ ;
  assign \new_[18797]_  = \new_[18796]_  & \new_[18791]_ ;
  assign \new_[18801]_  = A298 & A268;
  assign \new_[18802]_  = ~A202 & \new_[18801]_ ;
  assign \new_[18806]_  = ~A301 & ~A300;
  assign \new_[18807]_  = A299 & \new_[18806]_ ;
  assign \new_[18808]_  = \new_[18807]_  & \new_[18802]_ ;
  assign \new_[18812]_  = ~A168 & ~A169;
  assign \new_[18813]_  = ~A170 & \new_[18812]_ ;
  assign \new_[18817]_  = ~A201 & A200;
  assign \new_[18818]_  = A199 & \new_[18817]_ ;
  assign \new_[18819]_  = \new_[18818]_  & \new_[18813]_ ;
  assign \new_[18823]_  = A267 & A265;
  assign \new_[18824]_  = ~A202 & \new_[18823]_ ;
  assign \new_[18828]_  = ~A302 & ~A301;
  assign \new_[18829]_  = ~A300 & \new_[18828]_ ;
  assign \new_[18830]_  = \new_[18829]_  & \new_[18824]_ ;
  assign \new_[18834]_  = ~A168 & ~A169;
  assign \new_[18835]_  = ~A170 & \new_[18834]_ ;
  assign \new_[18839]_  = ~A201 & A200;
  assign \new_[18840]_  = A199 & \new_[18839]_ ;
  assign \new_[18841]_  = \new_[18840]_  & \new_[18835]_ ;
  assign \new_[18845]_  = A267 & A265;
  assign \new_[18846]_  = ~A202 & \new_[18845]_ ;
  assign \new_[18850]_  = ~A301 & ~A299;
  assign \new_[18851]_  = ~A298 & \new_[18850]_ ;
  assign \new_[18852]_  = \new_[18851]_  & \new_[18846]_ ;
  assign \new_[18856]_  = ~A168 & ~A169;
  assign \new_[18857]_  = ~A170 & \new_[18856]_ ;
  assign \new_[18861]_  = ~A201 & A200;
  assign \new_[18862]_  = A199 & \new_[18861]_ ;
  assign \new_[18863]_  = \new_[18862]_  & \new_[18857]_ ;
  assign \new_[18867]_  = A267 & A266;
  assign \new_[18868]_  = ~A202 & \new_[18867]_ ;
  assign \new_[18872]_  = ~A302 & ~A301;
  assign \new_[18873]_  = ~A300 & \new_[18872]_ ;
  assign \new_[18874]_  = \new_[18873]_  & \new_[18868]_ ;
  assign \new_[18878]_  = ~A168 & ~A169;
  assign \new_[18879]_  = ~A170 & \new_[18878]_ ;
  assign \new_[18883]_  = ~A201 & A200;
  assign \new_[18884]_  = A199 & \new_[18883]_ ;
  assign \new_[18885]_  = \new_[18884]_  & \new_[18879]_ ;
  assign \new_[18889]_  = A267 & A266;
  assign \new_[18890]_  = ~A202 & \new_[18889]_ ;
  assign \new_[18894]_  = ~A301 & ~A299;
  assign \new_[18895]_  = ~A298 & \new_[18894]_ ;
  assign \new_[18896]_  = \new_[18895]_  & \new_[18890]_ ;
  assign \new_[18900]_  = ~A168 & ~A169;
  assign \new_[18901]_  = ~A170 & \new_[18900]_ ;
  assign \new_[18905]_  = A203 & A200;
  assign \new_[18906]_  = ~A199 & \new_[18905]_ ;
  assign \new_[18907]_  = \new_[18906]_  & \new_[18901]_ ;
  assign \new_[18911]_  = ~A269 & ~A268;
  assign \new_[18912]_  = ~A267 & \new_[18911]_ ;
  assign \new_[18916]_  = A302 & ~A299;
  assign \new_[18917]_  = A298 & \new_[18916]_ ;
  assign \new_[18918]_  = \new_[18917]_  & \new_[18912]_ ;
  assign \new_[18922]_  = ~A168 & ~A169;
  assign \new_[18923]_  = ~A170 & \new_[18922]_ ;
  assign \new_[18927]_  = A203 & A200;
  assign \new_[18928]_  = ~A199 & \new_[18927]_ ;
  assign \new_[18929]_  = \new_[18928]_  & \new_[18923]_ ;
  assign \new_[18933]_  = ~A269 & ~A268;
  assign \new_[18934]_  = ~A267 & \new_[18933]_ ;
  assign \new_[18938]_  = A302 & A299;
  assign \new_[18939]_  = ~A298 & \new_[18938]_ ;
  assign \new_[18940]_  = \new_[18939]_  & \new_[18934]_ ;
  assign \new_[18944]_  = ~A168 & ~A169;
  assign \new_[18945]_  = ~A170 & \new_[18944]_ ;
  assign \new_[18949]_  = A203 & A200;
  assign \new_[18950]_  = ~A199 & \new_[18949]_ ;
  assign \new_[18951]_  = \new_[18950]_  & \new_[18945]_ ;
  assign \new_[18955]_  = ~A267 & A266;
  assign \new_[18956]_  = A265 & \new_[18955]_ ;
  assign \new_[18960]_  = A300 & A299;
  assign \new_[18961]_  = ~A268 & \new_[18960]_ ;
  assign \new_[18962]_  = \new_[18961]_  & \new_[18956]_ ;
  assign \new_[18966]_  = ~A168 & ~A169;
  assign \new_[18967]_  = ~A170 & \new_[18966]_ ;
  assign \new_[18971]_  = A203 & A200;
  assign \new_[18972]_  = ~A199 & \new_[18971]_ ;
  assign \new_[18973]_  = \new_[18972]_  & \new_[18967]_ ;
  assign \new_[18977]_  = ~A267 & A266;
  assign \new_[18978]_  = A265 & \new_[18977]_ ;
  assign \new_[18982]_  = A300 & A298;
  assign \new_[18983]_  = ~A268 & \new_[18982]_ ;
  assign \new_[18984]_  = \new_[18983]_  & \new_[18978]_ ;
  assign \new_[18988]_  = ~A168 & ~A169;
  assign \new_[18989]_  = ~A170 & \new_[18988]_ ;
  assign \new_[18993]_  = A203 & A200;
  assign \new_[18994]_  = ~A199 & \new_[18993]_ ;
  assign \new_[18995]_  = \new_[18994]_  & \new_[18989]_ ;
  assign \new_[18999]_  = ~A268 & ~A266;
  assign \new_[19000]_  = ~A265 & \new_[18999]_ ;
  assign \new_[19004]_  = A302 & ~A299;
  assign \new_[19005]_  = A298 & \new_[19004]_ ;
  assign \new_[19006]_  = \new_[19005]_  & \new_[19000]_ ;
  assign \new_[19010]_  = ~A168 & ~A169;
  assign \new_[19011]_  = ~A170 & \new_[19010]_ ;
  assign \new_[19015]_  = A203 & A200;
  assign \new_[19016]_  = ~A199 & \new_[19015]_ ;
  assign \new_[19017]_  = \new_[19016]_  & \new_[19011]_ ;
  assign \new_[19021]_  = ~A268 & ~A266;
  assign \new_[19022]_  = ~A265 & \new_[19021]_ ;
  assign \new_[19026]_  = A302 & A299;
  assign \new_[19027]_  = ~A298 & \new_[19026]_ ;
  assign \new_[19028]_  = \new_[19027]_  & \new_[19022]_ ;
  assign \new_[19032]_  = ~A168 & ~A169;
  assign \new_[19033]_  = ~A170 & \new_[19032]_ ;
  assign \new_[19037]_  = A203 & ~A200;
  assign \new_[19038]_  = A199 & \new_[19037]_ ;
  assign \new_[19039]_  = \new_[19038]_  & \new_[19033]_ ;
  assign \new_[19043]_  = ~A269 & ~A268;
  assign \new_[19044]_  = ~A267 & \new_[19043]_ ;
  assign \new_[19048]_  = A302 & ~A299;
  assign \new_[19049]_  = A298 & \new_[19048]_ ;
  assign \new_[19050]_  = \new_[19049]_  & \new_[19044]_ ;
  assign \new_[19054]_  = ~A168 & ~A169;
  assign \new_[19055]_  = ~A170 & \new_[19054]_ ;
  assign \new_[19059]_  = A203 & ~A200;
  assign \new_[19060]_  = A199 & \new_[19059]_ ;
  assign \new_[19061]_  = \new_[19060]_  & \new_[19055]_ ;
  assign \new_[19065]_  = ~A269 & ~A268;
  assign \new_[19066]_  = ~A267 & \new_[19065]_ ;
  assign \new_[19070]_  = A302 & A299;
  assign \new_[19071]_  = ~A298 & \new_[19070]_ ;
  assign \new_[19072]_  = \new_[19071]_  & \new_[19066]_ ;
  assign \new_[19076]_  = ~A168 & ~A169;
  assign \new_[19077]_  = ~A170 & \new_[19076]_ ;
  assign \new_[19081]_  = A203 & ~A200;
  assign \new_[19082]_  = A199 & \new_[19081]_ ;
  assign \new_[19083]_  = \new_[19082]_  & \new_[19077]_ ;
  assign \new_[19087]_  = ~A267 & A266;
  assign \new_[19088]_  = A265 & \new_[19087]_ ;
  assign \new_[19092]_  = A300 & A299;
  assign \new_[19093]_  = ~A268 & \new_[19092]_ ;
  assign \new_[19094]_  = \new_[19093]_  & \new_[19088]_ ;
  assign \new_[19098]_  = ~A168 & ~A169;
  assign \new_[19099]_  = ~A170 & \new_[19098]_ ;
  assign \new_[19103]_  = A203 & ~A200;
  assign \new_[19104]_  = A199 & \new_[19103]_ ;
  assign \new_[19105]_  = \new_[19104]_  & \new_[19099]_ ;
  assign \new_[19109]_  = ~A267 & A266;
  assign \new_[19110]_  = A265 & \new_[19109]_ ;
  assign \new_[19114]_  = A300 & A298;
  assign \new_[19115]_  = ~A268 & \new_[19114]_ ;
  assign \new_[19116]_  = \new_[19115]_  & \new_[19110]_ ;
  assign \new_[19120]_  = ~A168 & ~A169;
  assign \new_[19121]_  = ~A170 & \new_[19120]_ ;
  assign \new_[19125]_  = A203 & ~A200;
  assign \new_[19126]_  = A199 & \new_[19125]_ ;
  assign \new_[19127]_  = \new_[19126]_  & \new_[19121]_ ;
  assign \new_[19131]_  = ~A268 & ~A266;
  assign \new_[19132]_  = ~A265 & \new_[19131]_ ;
  assign \new_[19136]_  = A302 & ~A299;
  assign \new_[19137]_  = A298 & \new_[19136]_ ;
  assign \new_[19138]_  = \new_[19137]_  & \new_[19132]_ ;
  assign \new_[19142]_  = ~A168 & ~A169;
  assign \new_[19143]_  = ~A170 & \new_[19142]_ ;
  assign \new_[19147]_  = A203 & ~A200;
  assign \new_[19148]_  = A199 & \new_[19147]_ ;
  assign \new_[19149]_  = \new_[19148]_  & \new_[19143]_ ;
  assign \new_[19153]_  = ~A268 & ~A266;
  assign \new_[19154]_  = ~A265 & \new_[19153]_ ;
  assign \new_[19158]_  = A302 & A299;
  assign \new_[19159]_  = ~A298 & \new_[19158]_ ;
  assign \new_[19160]_  = \new_[19159]_  & \new_[19154]_ ;
  assign \new_[19164]_  = ~A168 & ~A169;
  assign \new_[19165]_  = ~A170 & \new_[19164]_ ;
  assign \new_[19169]_  = ~A202 & ~A200;
  assign \new_[19170]_  = ~A199 & \new_[19169]_ ;
  assign \new_[19171]_  = \new_[19170]_  & \new_[19165]_ ;
  assign \new_[19175]_  = A298 & A267;
  assign \new_[19176]_  = A265 & \new_[19175]_ ;
  assign \new_[19180]_  = ~A301 & ~A300;
  assign \new_[19181]_  = A299 & \new_[19180]_ ;
  assign \new_[19182]_  = \new_[19181]_  & \new_[19176]_ ;
  assign \new_[19186]_  = ~A168 & ~A169;
  assign \new_[19187]_  = ~A170 & \new_[19186]_ ;
  assign \new_[19191]_  = ~A202 & ~A200;
  assign \new_[19192]_  = ~A199 & \new_[19191]_ ;
  assign \new_[19193]_  = \new_[19192]_  & \new_[19187]_ ;
  assign \new_[19197]_  = A298 & A267;
  assign \new_[19198]_  = A266 & \new_[19197]_ ;
  assign \new_[19202]_  = ~A301 & ~A300;
  assign \new_[19203]_  = A299 & \new_[19202]_ ;
  assign \new_[19204]_  = \new_[19203]_  & \new_[19198]_ ;
  assign \new_[19208]_  = ~A168 & ~A169;
  assign \new_[19209]_  = ~A170 & \new_[19208]_ ;
  assign \new_[19213]_  = ~A202 & ~A200;
  assign \new_[19214]_  = ~A199 & \new_[19213]_ ;
  assign \new_[19215]_  = \new_[19214]_  & \new_[19209]_ ;
  assign \new_[19219]_  = A269 & A266;
  assign \new_[19220]_  = ~A265 & \new_[19219]_ ;
  assign \new_[19224]_  = ~A302 & ~A301;
  assign \new_[19225]_  = ~A300 & \new_[19224]_ ;
  assign \new_[19226]_  = \new_[19225]_  & \new_[19220]_ ;
  assign \new_[19230]_  = ~A168 & ~A169;
  assign \new_[19231]_  = ~A170 & \new_[19230]_ ;
  assign \new_[19235]_  = ~A202 & ~A200;
  assign \new_[19236]_  = ~A199 & \new_[19235]_ ;
  assign \new_[19237]_  = \new_[19236]_  & \new_[19231]_ ;
  assign \new_[19241]_  = A269 & A266;
  assign \new_[19242]_  = ~A265 & \new_[19241]_ ;
  assign \new_[19246]_  = ~A301 & ~A299;
  assign \new_[19247]_  = ~A298 & \new_[19246]_ ;
  assign \new_[19248]_  = \new_[19247]_  & \new_[19242]_ ;
  assign \new_[19252]_  = ~A168 & ~A169;
  assign \new_[19253]_  = ~A170 & \new_[19252]_ ;
  assign \new_[19257]_  = ~A202 & ~A200;
  assign \new_[19258]_  = ~A199 & \new_[19257]_ ;
  assign \new_[19259]_  = \new_[19258]_  & \new_[19253]_ ;
  assign \new_[19263]_  = A269 & ~A266;
  assign \new_[19264]_  = A265 & \new_[19263]_ ;
  assign \new_[19268]_  = ~A302 & ~A301;
  assign \new_[19269]_  = ~A300 & \new_[19268]_ ;
  assign \new_[19270]_  = \new_[19269]_  & \new_[19264]_ ;
  assign \new_[19274]_  = ~A168 & ~A169;
  assign \new_[19275]_  = ~A170 & \new_[19274]_ ;
  assign \new_[19279]_  = ~A202 & ~A200;
  assign \new_[19280]_  = ~A199 & \new_[19279]_ ;
  assign \new_[19281]_  = \new_[19280]_  & \new_[19275]_ ;
  assign \new_[19285]_  = A269 & ~A266;
  assign \new_[19286]_  = A265 & \new_[19285]_ ;
  assign \new_[19290]_  = ~A301 & ~A299;
  assign \new_[19291]_  = ~A298 & \new_[19290]_ ;
  assign \new_[19292]_  = \new_[19291]_  & \new_[19286]_ ;
  assign \new_[19296]_  = A199 & A166;
  assign \new_[19297]_  = A168 & \new_[19296]_ ;
  assign \new_[19301]_  = ~A202 & ~A201;
  assign \new_[19302]_  = A200 & \new_[19301]_ ;
  assign \new_[19303]_  = \new_[19302]_  & \new_[19297]_ ;
  assign \new_[19307]_  = ~A267 & A266;
  assign \new_[19308]_  = A265 & \new_[19307]_ ;
  assign \new_[19311]_  = A298 & ~A268;
  assign \new_[19314]_  = A302 & ~A299;
  assign \new_[19315]_  = \new_[19314]_  & \new_[19311]_ ;
  assign \new_[19316]_  = \new_[19315]_  & \new_[19308]_ ;
  assign \new_[19320]_  = A199 & A166;
  assign \new_[19321]_  = A168 & \new_[19320]_ ;
  assign \new_[19325]_  = ~A202 & ~A201;
  assign \new_[19326]_  = A200 & \new_[19325]_ ;
  assign \new_[19327]_  = \new_[19326]_  & \new_[19321]_ ;
  assign \new_[19331]_  = ~A267 & A266;
  assign \new_[19332]_  = A265 & \new_[19331]_ ;
  assign \new_[19335]_  = ~A298 & ~A268;
  assign \new_[19338]_  = A302 & A299;
  assign \new_[19339]_  = \new_[19338]_  & \new_[19335]_ ;
  assign \new_[19340]_  = \new_[19339]_  & \new_[19332]_ ;
  assign \new_[19344]_  = A199 & A167;
  assign \new_[19345]_  = A168 & \new_[19344]_ ;
  assign \new_[19349]_  = ~A202 & ~A201;
  assign \new_[19350]_  = A200 & \new_[19349]_ ;
  assign \new_[19351]_  = \new_[19350]_  & \new_[19345]_ ;
  assign \new_[19355]_  = ~A267 & A266;
  assign \new_[19356]_  = A265 & \new_[19355]_ ;
  assign \new_[19359]_  = A298 & ~A268;
  assign \new_[19362]_  = A302 & ~A299;
  assign \new_[19363]_  = \new_[19362]_  & \new_[19359]_ ;
  assign \new_[19364]_  = \new_[19363]_  & \new_[19356]_ ;
  assign \new_[19368]_  = A199 & A167;
  assign \new_[19369]_  = A168 & \new_[19368]_ ;
  assign \new_[19373]_  = ~A202 & ~A201;
  assign \new_[19374]_  = A200 & \new_[19373]_ ;
  assign \new_[19375]_  = \new_[19374]_  & \new_[19369]_ ;
  assign \new_[19379]_  = ~A267 & A266;
  assign \new_[19380]_  = A265 & \new_[19379]_ ;
  assign \new_[19383]_  = ~A298 & ~A268;
  assign \new_[19386]_  = A302 & A299;
  assign \new_[19387]_  = \new_[19386]_  & \new_[19383]_ ;
  assign \new_[19388]_  = \new_[19387]_  & \new_[19380]_ ;
  assign \new_[19392]_  = ~A166 & A167;
  assign \new_[19393]_  = A170 & \new_[19392]_ ;
  assign \new_[19397]_  = ~A203 & ~A202;
  assign \new_[19398]_  = ~A201 & \new_[19397]_ ;
  assign \new_[19399]_  = \new_[19398]_  & \new_[19393]_ ;
  assign \new_[19403]_  = ~A267 & A266;
  assign \new_[19404]_  = A265 & \new_[19403]_ ;
  assign \new_[19407]_  = A298 & ~A268;
  assign \new_[19410]_  = A302 & ~A299;
  assign \new_[19411]_  = \new_[19410]_  & \new_[19407]_ ;
  assign \new_[19412]_  = \new_[19411]_  & \new_[19404]_ ;
  assign \new_[19416]_  = ~A166 & A167;
  assign \new_[19417]_  = A170 & \new_[19416]_ ;
  assign \new_[19421]_  = ~A203 & ~A202;
  assign \new_[19422]_  = ~A201 & \new_[19421]_ ;
  assign \new_[19423]_  = \new_[19422]_  & \new_[19417]_ ;
  assign \new_[19427]_  = ~A267 & A266;
  assign \new_[19428]_  = A265 & \new_[19427]_ ;
  assign \new_[19431]_  = ~A298 & ~A268;
  assign \new_[19434]_  = A302 & A299;
  assign \new_[19435]_  = \new_[19434]_  & \new_[19431]_ ;
  assign \new_[19436]_  = \new_[19435]_  & \new_[19428]_ ;
  assign \new_[19440]_  = ~A166 & A167;
  assign \new_[19441]_  = A170 & \new_[19440]_ ;
  assign \new_[19445]_  = ~A201 & A200;
  assign \new_[19446]_  = A199 & \new_[19445]_ ;
  assign \new_[19447]_  = \new_[19446]_  & \new_[19441]_ ;
  assign \new_[19451]_  = ~A268 & ~A267;
  assign \new_[19452]_  = ~A202 & \new_[19451]_ ;
  assign \new_[19455]_  = A298 & ~A269;
  assign \new_[19458]_  = A302 & ~A299;
  assign \new_[19459]_  = \new_[19458]_  & \new_[19455]_ ;
  assign \new_[19460]_  = \new_[19459]_  & \new_[19452]_ ;
  assign \new_[19464]_  = ~A166 & A167;
  assign \new_[19465]_  = A170 & \new_[19464]_ ;
  assign \new_[19469]_  = ~A201 & A200;
  assign \new_[19470]_  = A199 & \new_[19469]_ ;
  assign \new_[19471]_  = \new_[19470]_  & \new_[19465]_ ;
  assign \new_[19475]_  = ~A268 & ~A267;
  assign \new_[19476]_  = ~A202 & \new_[19475]_ ;
  assign \new_[19479]_  = ~A298 & ~A269;
  assign \new_[19482]_  = A302 & A299;
  assign \new_[19483]_  = \new_[19482]_  & \new_[19479]_ ;
  assign \new_[19484]_  = \new_[19483]_  & \new_[19476]_ ;
  assign \new_[19488]_  = ~A166 & A167;
  assign \new_[19489]_  = A170 & \new_[19488]_ ;
  assign \new_[19493]_  = ~A201 & A200;
  assign \new_[19494]_  = A199 & \new_[19493]_ ;
  assign \new_[19495]_  = \new_[19494]_  & \new_[19489]_ ;
  assign \new_[19499]_  = A266 & A265;
  assign \new_[19500]_  = ~A202 & \new_[19499]_ ;
  assign \new_[19503]_  = ~A268 & ~A267;
  assign \new_[19506]_  = A300 & A299;
  assign \new_[19507]_  = \new_[19506]_  & \new_[19503]_ ;
  assign \new_[19508]_  = \new_[19507]_  & \new_[19500]_ ;
  assign \new_[19512]_  = ~A166 & A167;
  assign \new_[19513]_  = A170 & \new_[19512]_ ;
  assign \new_[19517]_  = ~A201 & A200;
  assign \new_[19518]_  = A199 & \new_[19517]_ ;
  assign \new_[19519]_  = \new_[19518]_  & \new_[19513]_ ;
  assign \new_[19523]_  = A266 & A265;
  assign \new_[19524]_  = ~A202 & \new_[19523]_ ;
  assign \new_[19527]_  = ~A268 & ~A267;
  assign \new_[19530]_  = A300 & A298;
  assign \new_[19531]_  = \new_[19530]_  & \new_[19527]_ ;
  assign \new_[19532]_  = \new_[19531]_  & \new_[19524]_ ;
  assign \new_[19536]_  = ~A166 & A167;
  assign \new_[19537]_  = A170 & \new_[19536]_ ;
  assign \new_[19541]_  = ~A201 & A200;
  assign \new_[19542]_  = A199 & \new_[19541]_ ;
  assign \new_[19543]_  = \new_[19542]_  & \new_[19537]_ ;
  assign \new_[19547]_  = ~A266 & ~A265;
  assign \new_[19548]_  = ~A202 & \new_[19547]_ ;
  assign \new_[19551]_  = A298 & ~A268;
  assign \new_[19554]_  = A302 & ~A299;
  assign \new_[19555]_  = \new_[19554]_  & \new_[19551]_ ;
  assign \new_[19556]_  = \new_[19555]_  & \new_[19548]_ ;
  assign \new_[19560]_  = ~A166 & A167;
  assign \new_[19561]_  = A170 & \new_[19560]_ ;
  assign \new_[19565]_  = ~A201 & A200;
  assign \new_[19566]_  = A199 & \new_[19565]_ ;
  assign \new_[19567]_  = \new_[19566]_  & \new_[19561]_ ;
  assign \new_[19571]_  = ~A266 & ~A265;
  assign \new_[19572]_  = ~A202 & \new_[19571]_ ;
  assign \new_[19575]_  = ~A298 & ~A268;
  assign \new_[19578]_  = A302 & A299;
  assign \new_[19579]_  = \new_[19578]_  & \new_[19575]_ ;
  assign \new_[19580]_  = \new_[19579]_  & \new_[19572]_ ;
  assign \new_[19584]_  = ~A166 & A167;
  assign \new_[19585]_  = A170 & \new_[19584]_ ;
  assign \new_[19589]_  = A203 & A200;
  assign \new_[19590]_  = ~A199 & \new_[19589]_ ;
  assign \new_[19591]_  = \new_[19590]_  & \new_[19585]_ ;
  assign \new_[19595]_  = A269 & A266;
  assign \new_[19596]_  = ~A265 & \new_[19595]_ ;
  assign \new_[19599]_  = A299 & A298;
  assign \new_[19602]_  = ~A301 & ~A300;
  assign \new_[19603]_  = \new_[19602]_  & \new_[19599]_ ;
  assign \new_[19604]_  = \new_[19603]_  & \new_[19596]_ ;
  assign \new_[19608]_  = ~A166 & A167;
  assign \new_[19609]_  = A170 & \new_[19608]_ ;
  assign \new_[19613]_  = A203 & A200;
  assign \new_[19614]_  = ~A199 & \new_[19613]_ ;
  assign \new_[19615]_  = \new_[19614]_  & \new_[19609]_ ;
  assign \new_[19619]_  = A269 & ~A266;
  assign \new_[19620]_  = A265 & \new_[19619]_ ;
  assign \new_[19623]_  = A299 & A298;
  assign \new_[19626]_  = ~A301 & ~A300;
  assign \new_[19627]_  = \new_[19626]_  & \new_[19623]_ ;
  assign \new_[19628]_  = \new_[19627]_  & \new_[19620]_ ;
  assign \new_[19632]_  = ~A166 & A167;
  assign \new_[19633]_  = A170 & \new_[19632]_ ;
  assign \new_[19637]_  = A203 & ~A200;
  assign \new_[19638]_  = A199 & \new_[19637]_ ;
  assign \new_[19639]_  = \new_[19638]_  & \new_[19633]_ ;
  assign \new_[19643]_  = A269 & A266;
  assign \new_[19644]_  = ~A265 & \new_[19643]_ ;
  assign \new_[19647]_  = A299 & A298;
  assign \new_[19650]_  = ~A301 & ~A300;
  assign \new_[19651]_  = \new_[19650]_  & \new_[19647]_ ;
  assign \new_[19652]_  = \new_[19651]_  & \new_[19644]_ ;
  assign \new_[19656]_  = ~A166 & A167;
  assign \new_[19657]_  = A170 & \new_[19656]_ ;
  assign \new_[19661]_  = A203 & ~A200;
  assign \new_[19662]_  = A199 & \new_[19661]_ ;
  assign \new_[19663]_  = \new_[19662]_  & \new_[19657]_ ;
  assign \new_[19667]_  = A269 & ~A266;
  assign \new_[19668]_  = A265 & \new_[19667]_ ;
  assign \new_[19671]_  = A299 & A298;
  assign \new_[19674]_  = ~A301 & ~A300;
  assign \new_[19675]_  = \new_[19674]_  & \new_[19671]_ ;
  assign \new_[19676]_  = \new_[19675]_  & \new_[19668]_ ;
  assign \new_[19680]_  = ~A166 & A167;
  assign \new_[19681]_  = A170 & \new_[19680]_ ;
  assign \new_[19685]_  = ~A202 & ~A200;
  assign \new_[19686]_  = ~A199 & \new_[19685]_ ;
  assign \new_[19687]_  = \new_[19686]_  & \new_[19681]_ ;
  assign \new_[19691]_  = ~A267 & A266;
  assign \new_[19692]_  = A265 & \new_[19691]_ ;
  assign \new_[19695]_  = A298 & ~A268;
  assign \new_[19698]_  = A302 & ~A299;
  assign \new_[19699]_  = \new_[19698]_  & \new_[19695]_ ;
  assign \new_[19700]_  = \new_[19699]_  & \new_[19692]_ ;
  assign \new_[19704]_  = ~A166 & A167;
  assign \new_[19705]_  = A170 & \new_[19704]_ ;
  assign \new_[19709]_  = ~A202 & ~A200;
  assign \new_[19710]_  = ~A199 & \new_[19709]_ ;
  assign \new_[19711]_  = \new_[19710]_  & \new_[19705]_ ;
  assign \new_[19715]_  = ~A267 & A266;
  assign \new_[19716]_  = A265 & \new_[19715]_ ;
  assign \new_[19719]_  = ~A298 & ~A268;
  assign \new_[19722]_  = A302 & A299;
  assign \new_[19723]_  = \new_[19722]_  & \new_[19719]_ ;
  assign \new_[19724]_  = \new_[19723]_  & \new_[19716]_ ;
  assign \new_[19728]_  = A166 & ~A167;
  assign \new_[19729]_  = A170 & \new_[19728]_ ;
  assign \new_[19733]_  = ~A203 & ~A202;
  assign \new_[19734]_  = ~A201 & \new_[19733]_ ;
  assign \new_[19735]_  = \new_[19734]_  & \new_[19729]_ ;
  assign \new_[19739]_  = ~A267 & A266;
  assign \new_[19740]_  = A265 & \new_[19739]_ ;
  assign \new_[19743]_  = A298 & ~A268;
  assign \new_[19746]_  = A302 & ~A299;
  assign \new_[19747]_  = \new_[19746]_  & \new_[19743]_ ;
  assign \new_[19748]_  = \new_[19747]_  & \new_[19740]_ ;
  assign \new_[19752]_  = A166 & ~A167;
  assign \new_[19753]_  = A170 & \new_[19752]_ ;
  assign \new_[19757]_  = ~A203 & ~A202;
  assign \new_[19758]_  = ~A201 & \new_[19757]_ ;
  assign \new_[19759]_  = \new_[19758]_  & \new_[19753]_ ;
  assign \new_[19763]_  = ~A267 & A266;
  assign \new_[19764]_  = A265 & \new_[19763]_ ;
  assign \new_[19767]_  = ~A298 & ~A268;
  assign \new_[19770]_  = A302 & A299;
  assign \new_[19771]_  = \new_[19770]_  & \new_[19767]_ ;
  assign \new_[19772]_  = \new_[19771]_  & \new_[19764]_ ;
  assign \new_[19776]_  = A166 & ~A167;
  assign \new_[19777]_  = A170 & \new_[19776]_ ;
  assign \new_[19781]_  = ~A201 & A200;
  assign \new_[19782]_  = A199 & \new_[19781]_ ;
  assign \new_[19783]_  = \new_[19782]_  & \new_[19777]_ ;
  assign \new_[19787]_  = ~A268 & ~A267;
  assign \new_[19788]_  = ~A202 & \new_[19787]_ ;
  assign \new_[19791]_  = A298 & ~A269;
  assign \new_[19794]_  = A302 & ~A299;
  assign \new_[19795]_  = \new_[19794]_  & \new_[19791]_ ;
  assign \new_[19796]_  = \new_[19795]_  & \new_[19788]_ ;
  assign \new_[19800]_  = A166 & ~A167;
  assign \new_[19801]_  = A170 & \new_[19800]_ ;
  assign \new_[19805]_  = ~A201 & A200;
  assign \new_[19806]_  = A199 & \new_[19805]_ ;
  assign \new_[19807]_  = \new_[19806]_  & \new_[19801]_ ;
  assign \new_[19811]_  = ~A268 & ~A267;
  assign \new_[19812]_  = ~A202 & \new_[19811]_ ;
  assign \new_[19815]_  = ~A298 & ~A269;
  assign \new_[19818]_  = A302 & A299;
  assign \new_[19819]_  = \new_[19818]_  & \new_[19815]_ ;
  assign \new_[19820]_  = \new_[19819]_  & \new_[19812]_ ;
  assign \new_[19824]_  = A166 & ~A167;
  assign \new_[19825]_  = A170 & \new_[19824]_ ;
  assign \new_[19829]_  = ~A201 & A200;
  assign \new_[19830]_  = A199 & \new_[19829]_ ;
  assign \new_[19831]_  = \new_[19830]_  & \new_[19825]_ ;
  assign \new_[19835]_  = A266 & A265;
  assign \new_[19836]_  = ~A202 & \new_[19835]_ ;
  assign \new_[19839]_  = ~A268 & ~A267;
  assign \new_[19842]_  = A300 & A299;
  assign \new_[19843]_  = \new_[19842]_  & \new_[19839]_ ;
  assign \new_[19844]_  = \new_[19843]_  & \new_[19836]_ ;
  assign \new_[19848]_  = A166 & ~A167;
  assign \new_[19849]_  = A170 & \new_[19848]_ ;
  assign \new_[19853]_  = ~A201 & A200;
  assign \new_[19854]_  = A199 & \new_[19853]_ ;
  assign \new_[19855]_  = \new_[19854]_  & \new_[19849]_ ;
  assign \new_[19859]_  = A266 & A265;
  assign \new_[19860]_  = ~A202 & \new_[19859]_ ;
  assign \new_[19863]_  = ~A268 & ~A267;
  assign \new_[19866]_  = A300 & A298;
  assign \new_[19867]_  = \new_[19866]_  & \new_[19863]_ ;
  assign \new_[19868]_  = \new_[19867]_  & \new_[19860]_ ;
  assign \new_[19872]_  = A166 & ~A167;
  assign \new_[19873]_  = A170 & \new_[19872]_ ;
  assign \new_[19877]_  = ~A201 & A200;
  assign \new_[19878]_  = A199 & \new_[19877]_ ;
  assign \new_[19879]_  = \new_[19878]_  & \new_[19873]_ ;
  assign \new_[19883]_  = ~A266 & ~A265;
  assign \new_[19884]_  = ~A202 & \new_[19883]_ ;
  assign \new_[19887]_  = A298 & ~A268;
  assign \new_[19890]_  = A302 & ~A299;
  assign \new_[19891]_  = \new_[19890]_  & \new_[19887]_ ;
  assign \new_[19892]_  = \new_[19891]_  & \new_[19884]_ ;
  assign \new_[19896]_  = A166 & ~A167;
  assign \new_[19897]_  = A170 & \new_[19896]_ ;
  assign \new_[19901]_  = ~A201 & A200;
  assign \new_[19902]_  = A199 & \new_[19901]_ ;
  assign \new_[19903]_  = \new_[19902]_  & \new_[19897]_ ;
  assign \new_[19907]_  = ~A266 & ~A265;
  assign \new_[19908]_  = ~A202 & \new_[19907]_ ;
  assign \new_[19911]_  = ~A298 & ~A268;
  assign \new_[19914]_  = A302 & A299;
  assign \new_[19915]_  = \new_[19914]_  & \new_[19911]_ ;
  assign \new_[19916]_  = \new_[19915]_  & \new_[19908]_ ;
  assign \new_[19920]_  = A166 & ~A167;
  assign \new_[19921]_  = A170 & \new_[19920]_ ;
  assign \new_[19925]_  = A203 & A200;
  assign \new_[19926]_  = ~A199 & \new_[19925]_ ;
  assign \new_[19927]_  = \new_[19926]_  & \new_[19921]_ ;
  assign \new_[19931]_  = A269 & A266;
  assign \new_[19932]_  = ~A265 & \new_[19931]_ ;
  assign \new_[19935]_  = A299 & A298;
  assign \new_[19938]_  = ~A301 & ~A300;
  assign \new_[19939]_  = \new_[19938]_  & \new_[19935]_ ;
  assign \new_[19940]_  = \new_[19939]_  & \new_[19932]_ ;
  assign \new_[19944]_  = A166 & ~A167;
  assign \new_[19945]_  = A170 & \new_[19944]_ ;
  assign \new_[19949]_  = A203 & A200;
  assign \new_[19950]_  = ~A199 & \new_[19949]_ ;
  assign \new_[19951]_  = \new_[19950]_  & \new_[19945]_ ;
  assign \new_[19955]_  = A269 & ~A266;
  assign \new_[19956]_  = A265 & \new_[19955]_ ;
  assign \new_[19959]_  = A299 & A298;
  assign \new_[19962]_  = ~A301 & ~A300;
  assign \new_[19963]_  = \new_[19962]_  & \new_[19959]_ ;
  assign \new_[19964]_  = \new_[19963]_  & \new_[19956]_ ;
  assign \new_[19968]_  = A166 & ~A167;
  assign \new_[19969]_  = A170 & \new_[19968]_ ;
  assign \new_[19973]_  = A203 & ~A200;
  assign \new_[19974]_  = A199 & \new_[19973]_ ;
  assign \new_[19975]_  = \new_[19974]_  & \new_[19969]_ ;
  assign \new_[19979]_  = A269 & A266;
  assign \new_[19980]_  = ~A265 & \new_[19979]_ ;
  assign \new_[19983]_  = A299 & A298;
  assign \new_[19986]_  = ~A301 & ~A300;
  assign \new_[19987]_  = \new_[19986]_  & \new_[19983]_ ;
  assign \new_[19988]_  = \new_[19987]_  & \new_[19980]_ ;
  assign \new_[19992]_  = A166 & ~A167;
  assign \new_[19993]_  = A170 & \new_[19992]_ ;
  assign \new_[19997]_  = A203 & ~A200;
  assign \new_[19998]_  = A199 & \new_[19997]_ ;
  assign \new_[19999]_  = \new_[19998]_  & \new_[19993]_ ;
  assign \new_[20003]_  = A269 & ~A266;
  assign \new_[20004]_  = A265 & \new_[20003]_ ;
  assign \new_[20007]_  = A299 & A298;
  assign \new_[20010]_  = ~A301 & ~A300;
  assign \new_[20011]_  = \new_[20010]_  & \new_[20007]_ ;
  assign \new_[20012]_  = \new_[20011]_  & \new_[20004]_ ;
  assign \new_[20016]_  = A166 & ~A167;
  assign \new_[20017]_  = A170 & \new_[20016]_ ;
  assign \new_[20021]_  = ~A202 & ~A200;
  assign \new_[20022]_  = ~A199 & \new_[20021]_ ;
  assign \new_[20023]_  = \new_[20022]_  & \new_[20017]_ ;
  assign \new_[20027]_  = ~A267 & A266;
  assign \new_[20028]_  = A265 & \new_[20027]_ ;
  assign \new_[20031]_  = A298 & ~A268;
  assign \new_[20034]_  = A302 & ~A299;
  assign \new_[20035]_  = \new_[20034]_  & \new_[20031]_ ;
  assign \new_[20036]_  = \new_[20035]_  & \new_[20028]_ ;
  assign \new_[20040]_  = A166 & ~A167;
  assign \new_[20041]_  = A170 & \new_[20040]_ ;
  assign \new_[20045]_  = ~A202 & ~A200;
  assign \new_[20046]_  = ~A199 & \new_[20045]_ ;
  assign \new_[20047]_  = \new_[20046]_  & \new_[20041]_ ;
  assign \new_[20051]_  = ~A267 & A266;
  assign \new_[20052]_  = A265 & \new_[20051]_ ;
  assign \new_[20055]_  = ~A298 & ~A268;
  assign \new_[20058]_  = A302 & A299;
  assign \new_[20059]_  = \new_[20058]_  & \new_[20055]_ ;
  assign \new_[20060]_  = \new_[20059]_  & \new_[20052]_ ;
  assign \new_[20064]_  = ~A166 & ~A167;
  assign \new_[20065]_  = ~A169 & \new_[20064]_ ;
  assign \new_[20069]_  = ~A203 & ~A202;
  assign \new_[20070]_  = ~A201 & \new_[20069]_ ;
  assign \new_[20071]_  = \new_[20070]_  & \new_[20065]_ ;
  assign \new_[20075]_  = A269 & A266;
  assign \new_[20076]_  = ~A265 & \new_[20075]_ ;
  assign \new_[20079]_  = A299 & A298;
  assign \new_[20082]_  = ~A301 & ~A300;
  assign \new_[20083]_  = \new_[20082]_  & \new_[20079]_ ;
  assign \new_[20084]_  = \new_[20083]_  & \new_[20076]_ ;
  assign \new_[20088]_  = ~A166 & ~A167;
  assign \new_[20089]_  = ~A169 & \new_[20088]_ ;
  assign \new_[20093]_  = ~A203 & ~A202;
  assign \new_[20094]_  = ~A201 & \new_[20093]_ ;
  assign \new_[20095]_  = \new_[20094]_  & \new_[20089]_ ;
  assign \new_[20099]_  = A269 & ~A266;
  assign \new_[20100]_  = A265 & \new_[20099]_ ;
  assign \new_[20103]_  = A299 & A298;
  assign \new_[20106]_  = ~A301 & ~A300;
  assign \new_[20107]_  = \new_[20106]_  & \new_[20103]_ ;
  assign \new_[20108]_  = \new_[20107]_  & \new_[20100]_ ;
  assign \new_[20112]_  = ~A166 & ~A167;
  assign \new_[20113]_  = ~A169 & \new_[20112]_ ;
  assign \new_[20117]_  = ~A201 & A200;
  assign \new_[20118]_  = A199 & \new_[20117]_ ;
  assign \new_[20119]_  = \new_[20118]_  & \new_[20113]_ ;
  assign \new_[20123]_  = A267 & A265;
  assign \new_[20124]_  = ~A202 & \new_[20123]_ ;
  assign \new_[20127]_  = A299 & A298;
  assign \new_[20130]_  = ~A301 & ~A300;
  assign \new_[20131]_  = \new_[20130]_  & \new_[20127]_ ;
  assign \new_[20132]_  = \new_[20131]_  & \new_[20124]_ ;
  assign \new_[20136]_  = ~A166 & ~A167;
  assign \new_[20137]_  = ~A169 & \new_[20136]_ ;
  assign \new_[20141]_  = ~A201 & A200;
  assign \new_[20142]_  = A199 & \new_[20141]_ ;
  assign \new_[20143]_  = \new_[20142]_  & \new_[20137]_ ;
  assign \new_[20147]_  = A267 & A266;
  assign \new_[20148]_  = ~A202 & \new_[20147]_ ;
  assign \new_[20151]_  = A299 & A298;
  assign \new_[20154]_  = ~A301 & ~A300;
  assign \new_[20155]_  = \new_[20154]_  & \new_[20151]_ ;
  assign \new_[20156]_  = \new_[20155]_  & \new_[20148]_ ;
  assign \new_[20160]_  = ~A166 & ~A167;
  assign \new_[20161]_  = ~A169 & \new_[20160]_ ;
  assign \new_[20165]_  = ~A201 & A200;
  assign \new_[20166]_  = A199 & \new_[20165]_ ;
  assign \new_[20167]_  = \new_[20166]_  & \new_[20161]_ ;
  assign \new_[20171]_  = A266 & ~A265;
  assign \new_[20172]_  = ~A202 & \new_[20171]_ ;
  assign \new_[20175]_  = ~A300 & A269;
  assign \new_[20178]_  = ~A302 & ~A301;
  assign \new_[20179]_  = \new_[20178]_  & \new_[20175]_ ;
  assign \new_[20180]_  = \new_[20179]_  & \new_[20172]_ ;
  assign \new_[20184]_  = ~A166 & ~A167;
  assign \new_[20185]_  = ~A169 & \new_[20184]_ ;
  assign \new_[20189]_  = ~A201 & A200;
  assign \new_[20190]_  = A199 & \new_[20189]_ ;
  assign \new_[20191]_  = \new_[20190]_  & \new_[20185]_ ;
  assign \new_[20195]_  = A266 & ~A265;
  assign \new_[20196]_  = ~A202 & \new_[20195]_ ;
  assign \new_[20199]_  = ~A298 & A269;
  assign \new_[20202]_  = ~A301 & ~A299;
  assign \new_[20203]_  = \new_[20202]_  & \new_[20199]_ ;
  assign \new_[20204]_  = \new_[20203]_  & \new_[20196]_ ;
  assign \new_[20208]_  = ~A166 & ~A167;
  assign \new_[20209]_  = ~A169 & \new_[20208]_ ;
  assign \new_[20213]_  = ~A201 & A200;
  assign \new_[20214]_  = A199 & \new_[20213]_ ;
  assign \new_[20215]_  = \new_[20214]_  & \new_[20209]_ ;
  assign \new_[20219]_  = ~A266 & A265;
  assign \new_[20220]_  = ~A202 & \new_[20219]_ ;
  assign \new_[20223]_  = ~A300 & A269;
  assign \new_[20226]_  = ~A302 & ~A301;
  assign \new_[20227]_  = \new_[20226]_  & \new_[20223]_ ;
  assign \new_[20228]_  = \new_[20227]_  & \new_[20220]_ ;
  assign \new_[20232]_  = ~A166 & ~A167;
  assign \new_[20233]_  = ~A169 & \new_[20232]_ ;
  assign \new_[20237]_  = ~A201 & A200;
  assign \new_[20238]_  = A199 & \new_[20237]_ ;
  assign \new_[20239]_  = \new_[20238]_  & \new_[20233]_ ;
  assign \new_[20243]_  = ~A266 & A265;
  assign \new_[20244]_  = ~A202 & \new_[20243]_ ;
  assign \new_[20247]_  = ~A298 & A269;
  assign \new_[20250]_  = ~A301 & ~A299;
  assign \new_[20251]_  = \new_[20250]_  & \new_[20247]_ ;
  assign \new_[20252]_  = \new_[20251]_  & \new_[20244]_ ;
  assign \new_[20256]_  = ~A166 & ~A167;
  assign \new_[20257]_  = ~A169 & \new_[20256]_ ;
  assign \new_[20261]_  = A203 & A200;
  assign \new_[20262]_  = ~A199 & \new_[20261]_ ;
  assign \new_[20263]_  = \new_[20262]_  & \new_[20257]_ ;
  assign \new_[20267]_  = ~A267 & A266;
  assign \new_[20268]_  = A265 & \new_[20267]_ ;
  assign \new_[20271]_  = A298 & ~A268;
  assign \new_[20274]_  = A302 & ~A299;
  assign \new_[20275]_  = \new_[20274]_  & \new_[20271]_ ;
  assign \new_[20276]_  = \new_[20275]_  & \new_[20268]_ ;
  assign \new_[20280]_  = ~A166 & ~A167;
  assign \new_[20281]_  = ~A169 & \new_[20280]_ ;
  assign \new_[20285]_  = A203 & A200;
  assign \new_[20286]_  = ~A199 & \new_[20285]_ ;
  assign \new_[20287]_  = \new_[20286]_  & \new_[20281]_ ;
  assign \new_[20291]_  = ~A267 & A266;
  assign \new_[20292]_  = A265 & \new_[20291]_ ;
  assign \new_[20295]_  = ~A298 & ~A268;
  assign \new_[20298]_  = A302 & A299;
  assign \new_[20299]_  = \new_[20298]_  & \new_[20295]_ ;
  assign \new_[20300]_  = \new_[20299]_  & \new_[20292]_ ;
  assign \new_[20304]_  = ~A166 & ~A167;
  assign \new_[20305]_  = ~A169 & \new_[20304]_ ;
  assign \new_[20309]_  = A203 & ~A200;
  assign \new_[20310]_  = A199 & \new_[20309]_ ;
  assign \new_[20311]_  = \new_[20310]_  & \new_[20305]_ ;
  assign \new_[20315]_  = ~A267 & A266;
  assign \new_[20316]_  = A265 & \new_[20315]_ ;
  assign \new_[20319]_  = A298 & ~A268;
  assign \new_[20322]_  = A302 & ~A299;
  assign \new_[20323]_  = \new_[20322]_  & \new_[20319]_ ;
  assign \new_[20324]_  = \new_[20323]_  & \new_[20316]_ ;
  assign \new_[20328]_  = ~A166 & ~A167;
  assign \new_[20329]_  = ~A169 & \new_[20328]_ ;
  assign \new_[20333]_  = A203 & ~A200;
  assign \new_[20334]_  = A199 & \new_[20333]_ ;
  assign \new_[20335]_  = \new_[20334]_  & \new_[20329]_ ;
  assign \new_[20339]_  = ~A267 & A266;
  assign \new_[20340]_  = A265 & \new_[20339]_ ;
  assign \new_[20343]_  = ~A298 & ~A268;
  assign \new_[20346]_  = A302 & A299;
  assign \new_[20347]_  = \new_[20346]_  & \new_[20343]_ ;
  assign \new_[20348]_  = \new_[20347]_  & \new_[20340]_ ;
  assign \new_[20352]_  = ~A166 & ~A167;
  assign \new_[20353]_  = ~A169 & \new_[20352]_ ;
  assign \new_[20357]_  = ~A202 & ~A200;
  assign \new_[20358]_  = ~A199 & \new_[20357]_ ;
  assign \new_[20359]_  = \new_[20358]_  & \new_[20353]_ ;
  assign \new_[20363]_  = A269 & A266;
  assign \new_[20364]_  = ~A265 & \new_[20363]_ ;
  assign \new_[20367]_  = A299 & A298;
  assign \new_[20370]_  = ~A301 & ~A300;
  assign \new_[20371]_  = \new_[20370]_  & \new_[20367]_ ;
  assign \new_[20372]_  = \new_[20371]_  & \new_[20364]_ ;
  assign \new_[20376]_  = ~A166 & ~A167;
  assign \new_[20377]_  = ~A169 & \new_[20376]_ ;
  assign \new_[20381]_  = ~A202 & ~A200;
  assign \new_[20382]_  = ~A199 & \new_[20381]_ ;
  assign \new_[20383]_  = \new_[20382]_  & \new_[20377]_ ;
  assign \new_[20387]_  = A269 & ~A266;
  assign \new_[20388]_  = A265 & \new_[20387]_ ;
  assign \new_[20391]_  = A299 & A298;
  assign \new_[20394]_  = ~A301 & ~A300;
  assign \new_[20395]_  = \new_[20394]_  & \new_[20391]_ ;
  assign \new_[20396]_  = \new_[20395]_  & \new_[20388]_ ;
  assign \new_[20400]_  = A167 & ~A168;
  assign \new_[20401]_  = ~A169 & \new_[20400]_ ;
  assign \new_[20405]_  = ~A202 & ~A201;
  assign \new_[20406]_  = A166 & \new_[20405]_ ;
  assign \new_[20407]_  = \new_[20406]_  & \new_[20401]_ ;
  assign \new_[20411]_  = A267 & A265;
  assign \new_[20412]_  = ~A203 & \new_[20411]_ ;
  assign \new_[20415]_  = A299 & A298;
  assign \new_[20418]_  = ~A301 & ~A300;
  assign \new_[20419]_  = \new_[20418]_  & \new_[20415]_ ;
  assign \new_[20420]_  = \new_[20419]_  & \new_[20412]_ ;
  assign \new_[20424]_  = A167 & ~A168;
  assign \new_[20425]_  = ~A169 & \new_[20424]_ ;
  assign \new_[20429]_  = ~A202 & ~A201;
  assign \new_[20430]_  = A166 & \new_[20429]_ ;
  assign \new_[20431]_  = \new_[20430]_  & \new_[20425]_ ;
  assign \new_[20435]_  = A267 & A266;
  assign \new_[20436]_  = ~A203 & \new_[20435]_ ;
  assign \new_[20439]_  = A299 & A298;
  assign \new_[20442]_  = ~A301 & ~A300;
  assign \new_[20443]_  = \new_[20442]_  & \new_[20439]_ ;
  assign \new_[20444]_  = \new_[20443]_  & \new_[20436]_ ;
  assign \new_[20448]_  = A167 & ~A168;
  assign \new_[20449]_  = ~A169 & \new_[20448]_ ;
  assign \new_[20453]_  = ~A202 & ~A201;
  assign \new_[20454]_  = A166 & \new_[20453]_ ;
  assign \new_[20455]_  = \new_[20454]_  & \new_[20449]_ ;
  assign \new_[20459]_  = A266 & ~A265;
  assign \new_[20460]_  = ~A203 & \new_[20459]_ ;
  assign \new_[20463]_  = ~A300 & A269;
  assign \new_[20466]_  = ~A302 & ~A301;
  assign \new_[20467]_  = \new_[20466]_  & \new_[20463]_ ;
  assign \new_[20468]_  = \new_[20467]_  & \new_[20460]_ ;
  assign \new_[20472]_  = A167 & ~A168;
  assign \new_[20473]_  = ~A169 & \new_[20472]_ ;
  assign \new_[20477]_  = ~A202 & ~A201;
  assign \new_[20478]_  = A166 & \new_[20477]_ ;
  assign \new_[20479]_  = \new_[20478]_  & \new_[20473]_ ;
  assign \new_[20483]_  = A266 & ~A265;
  assign \new_[20484]_  = ~A203 & \new_[20483]_ ;
  assign \new_[20487]_  = ~A298 & A269;
  assign \new_[20490]_  = ~A301 & ~A299;
  assign \new_[20491]_  = \new_[20490]_  & \new_[20487]_ ;
  assign \new_[20492]_  = \new_[20491]_  & \new_[20484]_ ;
  assign \new_[20496]_  = A167 & ~A168;
  assign \new_[20497]_  = ~A169 & \new_[20496]_ ;
  assign \new_[20501]_  = ~A202 & ~A201;
  assign \new_[20502]_  = A166 & \new_[20501]_ ;
  assign \new_[20503]_  = \new_[20502]_  & \new_[20497]_ ;
  assign \new_[20507]_  = ~A266 & A265;
  assign \new_[20508]_  = ~A203 & \new_[20507]_ ;
  assign \new_[20511]_  = ~A300 & A269;
  assign \new_[20514]_  = ~A302 & ~A301;
  assign \new_[20515]_  = \new_[20514]_  & \new_[20511]_ ;
  assign \new_[20516]_  = \new_[20515]_  & \new_[20508]_ ;
  assign \new_[20520]_  = A167 & ~A168;
  assign \new_[20521]_  = ~A169 & \new_[20520]_ ;
  assign \new_[20525]_  = ~A202 & ~A201;
  assign \new_[20526]_  = A166 & \new_[20525]_ ;
  assign \new_[20527]_  = \new_[20526]_  & \new_[20521]_ ;
  assign \new_[20531]_  = ~A266 & A265;
  assign \new_[20532]_  = ~A203 & \new_[20531]_ ;
  assign \new_[20535]_  = ~A298 & A269;
  assign \new_[20538]_  = ~A301 & ~A299;
  assign \new_[20539]_  = \new_[20538]_  & \new_[20535]_ ;
  assign \new_[20540]_  = \new_[20539]_  & \new_[20532]_ ;
  assign \new_[20544]_  = A167 & ~A168;
  assign \new_[20545]_  = ~A169 & \new_[20544]_ ;
  assign \new_[20549]_  = A201 & A199;
  assign \new_[20550]_  = A166 & \new_[20549]_ ;
  assign \new_[20551]_  = \new_[20550]_  & \new_[20545]_ ;
  assign \new_[20555]_  = ~A267 & A266;
  assign \new_[20556]_  = A265 & \new_[20555]_ ;
  assign \new_[20559]_  = A298 & ~A268;
  assign \new_[20562]_  = A302 & ~A299;
  assign \new_[20563]_  = \new_[20562]_  & \new_[20559]_ ;
  assign \new_[20564]_  = \new_[20563]_  & \new_[20556]_ ;
  assign \new_[20568]_  = A167 & ~A168;
  assign \new_[20569]_  = ~A169 & \new_[20568]_ ;
  assign \new_[20573]_  = A201 & A199;
  assign \new_[20574]_  = A166 & \new_[20573]_ ;
  assign \new_[20575]_  = \new_[20574]_  & \new_[20569]_ ;
  assign \new_[20579]_  = ~A267 & A266;
  assign \new_[20580]_  = A265 & \new_[20579]_ ;
  assign \new_[20583]_  = ~A298 & ~A268;
  assign \new_[20586]_  = A302 & A299;
  assign \new_[20587]_  = \new_[20586]_  & \new_[20583]_ ;
  assign \new_[20588]_  = \new_[20587]_  & \new_[20580]_ ;
  assign \new_[20592]_  = A167 & ~A168;
  assign \new_[20593]_  = ~A169 & \new_[20592]_ ;
  assign \new_[20597]_  = A201 & A200;
  assign \new_[20598]_  = A166 & \new_[20597]_ ;
  assign \new_[20599]_  = \new_[20598]_  & \new_[20593]_ ;
  assign \new_[20603]_  = ~A267 & A266;
  assign \new_[20604]_  = A265 & \new_[20603]_ ;
  assign \new_[20607]_  = A298 & ~A268;
  assign \new_[20610]_  = A302 & ~A299;
  assign \new_[20611]_  = \new_[20610]_  & \new_[20607]_ ;
  assign \new_[20612]_  = \new_[20611]_  & \new_[20604]_ ;
  assign \new_[20616]_  = A167 & ~A168;
  assign \new_[20617]_  = ~A169 & \new_[20616]_ ;
  assign \new_[20621]_  = A201 & A200;
  assign \new_[20622]_  = A166 & \new_[20621]_ ;
  assign \new_[20623]_  = \new_[20622]_  & \new_[20617]_ ;
  assign \new_[20627]_  = ~A267 & A266;
  assign \new_[20628]_  = A265 & \new_[20627]_ ;
  assign \new_[20631]_  = ~A298 & ~A268;
  assign \new_[20634]_  = A302 & A299;
  assign \new_[20635]_  = \new_[20634]_  & \new_[20631]_ ;
  assign \new_[20636]_  = \new_[20635]_  & \new_[20628]_ ;
  assign \new_[20640]_  = A167 & ~A168;
  assign \new_[20641]_  = ~A169 & \new_[20640]_ ;
  assign \new_[20645]_  = A200 & A199;
  assign \new_[20646]_  = A166 & \new_[20645]_ ;
  assign \new_[20647]_  = \new_[20646]_  & \new_[20641]_ ;
  assign \new_[20651]_  = A268 & ~A202;
  assign \new_[20652]_  = ~A201 & \new_[20651]_ ;
  assign \new_[20655]_  = A299 & A298;
  assign \new_[20658]_  = ~A301 & ~A300;
  assign \new_[20659]_  = \new_[20658]_  & \new_[20655]_ ;
  assign \new_[20660]_  = \new_[20659]_  & \new_[20652]_ ;
  assign \new_[20664]_  = A167 & ~A168;
  assign \new_[20665]_  = ~A169 & \new_[20664]_ ;
  assign \new_[20669]_  = A200 & A199;
  assign \new_[20670]_  = A166 & \new_[20669]_ ;
  assign \new_[20671]_  = \new_[20670]_  & \new_[20665]_ ;
  assign \new_[20675]_  = A265 & ~A202;
  assign \new_[20676]_  = ~A201 & \new_[20675]_ ;
  assign \new_[20679]_  = ~A300 & A267;
  assign \new_[20682]_  = ~A302 & ~A301;
  assign \new_[20683]_  = \new_[20682]_  & \new_[20679]_ ;
  assign \new_[20684]_  = \new_[20683]_  & \new_[20676]_ ;
  assign \new_[20688]_  = A167 & ~A168;
  assign \new_[20689]_  = ~A169 & \new_[20688]_ ;
  assign \new_[20693]_  = A200 & A199;
  assign \new_[20694]_  = A166 & \new_[20693]_ ;
  assign \new_[20695]_  = \new_[20694]_  & \new_[20689]_ ;
  assign \new_[20699]_  = A265 & ~A202;
  assign \new_[20700]_  = ~A201 & \new_[20699]_ ;
  assign \new_[20703]_  = ~A298 & A267;
  assign \new_[20706]_  = ~A301 & ~A299;
  assign \new_[20707]_  = \new_[20706]_  & \new_[20703]_ ;
  assign \new_[20708]_  = \new_[20707]_  & \new_[20700]_ ;
  assign \new_[20712]_  = A167 & ~A168;
  assign \new_[20713]_  = ~A169 & \new_[20712]_ ;
  assign \new_[20717]_  = A200 & A199;
  assign \new_[20718]_  = A166 & \new_[20717]_ ;
  assign \new_[20719]_  = \new_[20718]_  & \new_[20713]_ ;
  assign \new_[20723]_  = A266 & ~A202;
  assign \new_[20724]_  = ~A201 & \new_[20723]_ ;
  assign \new_[20727]_  = ~A300 & A267;
  assign \new_[20730]_  = ~A302 & ~A301;
  assign \new_[20731]_  = \new_[20730]_  & \new_[20727]_ ;
  assign \new_[20732]_  = \new_[20731]_  & \new_[20724]_ ;
  assign \new_[20736]_  = A167 & ~A168;
  assign \new_[20737]_  = ~A169 & \new_[20736]_ ;
  assign \new_[20741]_  = A200 & A199;
  assign \new_[20742]_  = A166 & \new_[20741]_ ;
  assign \new_[20743]_  = \new_[20742]_  & \new_[20737]_ ;
  assign \new_[20747]_  = A266 & ~A202;
  assign \new_[20748]_  = ~A201 & \new_[20747]_ ;
  assign \new_[20751]_  = ~A298 & A267;
  assign \new_[20754]_  = ~A301 & ~A299;
  assign \new_[20755]_  = \new_[20754]_  & \new_[20751]_ ;
  assign \new_[20756]_  = \new_[20755]_  & \new_[20748]_ ;
  assign \new_[20760]_  = A167 & ~A168;
  assign \new_[20761]_  = ~A169 & \new_[20760]_ ;
  assign \new_[20765]_  = A200 & ~A199;
  assign \new_[20766]_  = A166 & \new_[20765]_ ;
  assign \new_[20767]_  = \new_[20766]_  & \new_[20761]_ ;
  assign \new_[20771]_  = ~A268 & ~A267;
  assign \new_[20772]_  = A203 & \new_[20771]_ ;
  assign \new_[20775]_  = A298 & ~A269;
  assign \new_[20778]_  = A302 & ~A299;
  assign \new_[20779]_  = \new_[20778]_  & \new_[20775]_ ;
  assign \new_[20780]_  = \new_[20779]_  & \new_[20772]_ ;
  assign \new_[20784]_  = A167 & ~A168;
  assign \new_[20785]_  = ~A169 & \new_[20784]_ ;
  assign \new_[20789]_  = A200 & ~A199;
  assign \new_[20790]_  = A166 & \new_[20789]_ ;
  assign \new_[20791]_  = \new_[20790]_  & \new_[20785]_ ;
  assign \new_[20795]_  = ~A268 & ~A267;
  assign \new_[20796]_  = A203 & \new_[20795]_ ;
  assign \new_[20799]_  = ~A298 & ~A269;
  assign \new_[20802]_  = A302 & A299;
  assign \new_[20803]_  = \new_[20802]_  & \new_[20799]_ ;
  assign \new_[20804]_  = \new_[20803]_  & \new_[20796]_ ;
  assign \new_[20808]_  = A167 & ~A168;
  assign \new_[20809]_  = ~A169 & \new_[20808]_ ;
  assign \new_[20813]_  = A200 & ~A199;
  assign \new_[20814]_  = A166 & \new_[20813]_ ;
  assign \new_[20815]_  = \new_[20814]_  & \new_[20809]_ ;
  assign \new_[20819]_  = A266 & A265;
  assign \new_[20820]_  = A203 & \new_[20819]_ ;
  assign \new_[20823]_  = ~A268 & ~A267;
  assign \new_[20826]_  = A300 & A299;
  assign \new_[20827]_  = \new_[20826]_  & \new_[20823]_ ;
  assign \new_[20828]_  = \new_[20827]_  & \new_[20820]_ ;
  assign \new_[20832]_  = A167 & ~A168;
  assign \new_[20833]_  = ~A169 & \new_[20832]_ ;
  assign \new_[20837]_  = A200 & ~A199;
  assign \new_[20838]_  = A166 & \new_[20837]_ ;
  assign \new_[20839]_  = \new_[20838]_  & \new_[20833]_ ;
  assign \new_[20843]_  = A266 & A265;
  assign \new_[20844]_  = A203 & \new_[20843]_ ;
  assign \new_[20847]_  = ~A268 & ~A267;
  assign \new_[20850]_  = A300 & A298;
  assign \new_[20851]_  = \new_[20850]_  & \new_[20847]_ ;
  assign \new_[20852]_  = \new_[20851]_  & \new_[20844]_ ;
  assign \new_[20856]_  = A167 & ~A168;
  assign \new_[20857]_  = ~A169 & \new_[20856]_ ;
  assign \new_[20861]_  = A200 & ~A199;
  assign \new_[20862]_  = A166 & \new_[20861]_ ;
  assign \new_[20863]_  = \new_[20862]_  & \new_[20857]_ ;
  assign \new_[20867]_  = ~A266 & ~A265;
  assign \new_[20868]_  = A203 & \new_[20867]_ ;
  assign \new_[20871]_  = A298 & ~A268;
  assign \new_[20874]_  = A302 & ~A299;
  assign \new_[20875]_  = \new_[20874]_  & \new_[20871]_ ;
  assign \new_[20876]_  = \new_[20875]_  & \new_[20868]_ ;
  assign \new_[20880]_  = A167 & ~A168;
  assign \new_[20881]_  = ~A169 & \new_[20880]_ ;
  assign \new_[20885]_  = A200 & ~A199;
  assign \new_[20886]_  = A166 & \new_[20885]_ ;
  assign \new_[20887]_  = \new_[20886]_  & \new_[20881]_ ;
  assign \new_[20891]_  = ~A266 & ~A265;
  assign \new_[20892]_  = A203 & \new_[20891]_ ;
  assign \new_[20895]_  = ~A298 & ~A268;
  assign \new_[20898]_  = A302 & A299;
  assign \new_[20899]_  = \new_[20898]_  & \new_[20895]_ ;
  assign \new_[20900]_  = \new_[20899]_  & \new_[20892]_ ;
  assign \new_[20904]_  = A167 & ~A168;
  assign \new_[20905]_  = ~A169 & \new_[20904]_ ;
  assign \new_[20909]_  = ~A200 & A199;
  assign \new_[20910]_  = A166 & \new_[20909]_ ;
  assign \new_[20911]_  = \new_[20910]_  & \new_[20905]_ ;
  assign \new_[20915]_  = ~A268 & ~A267;
  assign \new_[20916]_  = A203 & \new_[20915]_ ;
  assign \new_[20919]_  = A298 & ~A269;
  assign \new_[20922]_  = A302 & ~A299;
  assign \new_[20923]_  = \new_[20922]_  & \new_[20919]_ ;
  assign \new_[20924]_  = \new_[20923]_  & \new_[20916]_ ;
  assign \new_[20928]_  = A167 & ~A168;
  assign \new_[20929]_  = ~A169 & \new_[20928]_ ;
  assign \new_[20933]_  = ~A200 & A199;
  assign \new_[20934]_  = A166 & \new_[20933]_ ;
  assign \new_[20935]_  = \new_[20934]_  & \new_[20929]_ ;
  assign \new_[20939]_  = ~A268 & ~A267;
  assign \new_[20940]_  = A203 & \new_[20939]_ ;
  assign \new_[20943]_  = ~A298 & ~A269;
  assign \new_[20946]_  = A302 & A299;
  assign \new_[20947]_  = \new_[20946]_  & \new_[20943]_ ;
  assign \new_[20948]_  = \new_[20947]_  & \new_[20940]_ ;
  assign \new_[20952]_  = A167 & ~A168;
  assign \new_[20953]_  = ~A169 & \new_[20952]_ ;
  assign \new_[20957]_  = ~A200 & A199;
  assign \new_[20958]_  = A166 & \new_[20957]_ ;
  assign \new_[20959]_  = \new_[20958]_  & \new_[20953]_ ;
  assign \new_[20963]_  = A266 & A265;
  assign \new_[20964]_  = A203 & \new_[20963]_ ;
  assign \new_[20967]_  = ~A268 & ~A267;
  assign \new_[20970]_  = A300 & A299;
  assign \new_[20971]_  = \new_[20970]_  & \new_[20967]_ ;
  assign \new_[20972]_  = \new_[20971]_  & \new_[20964]_ ;
  assign \new_[20976]_  = A167 & ~A168;
  assign \new_[20977]_  = ~A169 & \new_[20976]_ ;
  assign \new_[20981]_  = ~A200 & A199;
  assign \new_[20982]_  = A166 & \new_[20981]_ ;
  assign \new_[20983]_  = \new_[20982]_  & \new_[20977]_ ;
  assign \new_[20987]_  = A266 & A265;
  assign \new_[20988]_  = A203 & \new_[20987]_ ;
  assign \new_[20991]_  = ~A268 & ~A267;
  assign \new_[20994]_  = A300 & A298;
  assign \new_[20995]_  = \new_[20994]_  & \new_[20991]_ ;
  assign \new_[20996]_  = \new_[20995]_  & \new_[20988]_ ;
  assign \new_[21000]_  = A167 & ~A168;
  assign \new_[21001]_  = ~A169 & \new_[21000]_ ;
  assign \new_[21005]_  = ~A200 & A199;
  assign \new_[21006]_  = A166 & \new_[21005]_ ;
  assign \new_[21007]_  = \new_[21006]_  & \new_[21001]_ ;
  assign \new_[21011]_  = ~A266 & ~A265;
  assign \new_[21012]_  = A203 & \new_[21011]_ ;
  assign \new_[21015]_  = A298 & ~A268;
  assign \new_[21018]_  = A302 & ~A299;
  assign \new_[21019]_  = \new_[21018]_  & \new_[21015]_ ;
  assign \new_[21020]_  = \new_[21019]_  & \new_[21012]_ ;
  assign \new_[21024]_  = A167 & ~A168;
  assign \new_[21025]_  = ~A169 & \new_[21024]_ ;
  assign \new_[21029]_  = ~A200 & A199;
  assign \new_[21030]_  = A166 & \new_[21029]_ ;
  assign \new_[21031]_  = \new_[21030]_  & \new_[21025]_ ;
  assign \new_[21035]_  = ~A266 & ~A265;
  assign \new_[21036]_  = A203 & \new_[21035]_ ;
  assign \new_[21039]_  = ~A298 & ~A268;
  assign \new_[21042]_  = A302 & A299;
  assign \new_[21043]_  = \new_[21042]_  & \new_[21039]_ ;
  assign \new_[21044]_  = \new_[21043]_  & \new_[21036]_ ;
  assign \new_[21048]_  = A167 & ~A168;
  assign \new_[21049]_  = ~A169 & \new_[21048]_ ;
  assign \new_[21053]_  = ~A200 & ~A199;
  assign \new_[21054]_  = A166 & \new_[21053]_ ;
  assign \new_[21055]_  = \new_[21054]_  & \new_[21049]_ ;
  assign \new_[21059]_  = A267 & A265;
  assign \new_[21060]_  = ~A202 & \new_[21059]_ ;
  assign \new_[21063]_  = A299 & A298;
  assign \new_[21066]_  = ~A301 & ~A300;
  assign \new_[21067]_  = \new_[21066]_  & \new_[21063]_ ;
  assign \new_[21068]_  = \new_[21067]_  & \new_[21060]_ ;
  assign \new_[21072]_  = A167 & ~A168;
  assign \new_[21073]_  = ~A169 & \new_[21072]_ ;
  assign \new_[21077]_  = ~A200 & ~A199;
  assign \new_[21078]_  = A166 & \new_[21077]_ ;
  assign \new_[21079]_  = \new_[21078]_  & \new_[21073]_ ;
  assign \new_[21083]_  = A267 & A266;
  assign \new_[21084]_  = ~A202 & \new_[21083]_ ;
  assign \new_[21087]_  = A299 & A298;
  assign \new_[21090]_  = ~A301 & ~A300;
  assign \new_[21091]_  = \new_[21090]_  & \new_[21087]_ ;
  assign \new_[21092]_  = \new_[21091]_  & \new_[21084]_ ;
  assign \new_[21096]_  = A167 & ~A168;
  assign \new_[21097]_  = ~A169 & \new_[21096]_ ;
  assign \new_[21101]_  = ~A200 & ~A199;
  assign \new_[21102]_  = A166 & \new_[21101]_ ;
  assign \new_[21103]_  = \new_[21102]_  & \new_[21097]_ ;
  assign \new_[21107]_  = A266 & ~A265;
  assign \new_[21108]_  = ~A202 & \new_[21107]_ ;
  assign \new_[21111]_  = ~A300 & A269;
  assign \new_[21114]_  = ~A302 & ~A301;
  assign \new_[21115]_  = \new_[21114]_  & \new_[21111]_ ;
  assign \new_[21116]_  = \new_[21115]_  & \new_[21108]_ ;
  assign \new_[21120]_  = A167 & ~A168;
  assign \new_[21121]_  = ~A169 & \new_[21120]_ ;
  assign \new_[21125]_  = ~A200 & ~A199;
  assign \new_[21126]_  = A166 & \new_[21125]_ ;
  assign \new_[21127]_  = \new_[21126]_  & \new_[21121]_ ;
  assign \new_[21131]_  = A266 & ~A265;
  assign \new_[21132]_  = ~A202 & \new_[21131]_ ;
  assign \new_[21135]_  = ~A298 & A269;
  assign \new_[21138]_  = ~A301 & ~A299;
  assign \new_[21139]_  = \new_[21138]_  & \new_[21135]_ ;
  assign \new_[21140]_  = \new_[21139]_  & \new_[21132]_ ;
  assign \new_[21144]_  = A167 & ~A168;
  assign \new_[21145]_  = ~A169 & \new_[21144]_ ;
  assign \new_[21149]_  = ~A200 & ~A199;
  assign \new_[21150]_  = A166 & \new_[21149]_ ;
  assign \new_[21151]_  = \new_[21150]_  & \new_[21145]_ ;
  assign \new_[21155]_  = ~A266 & A265;
  assign \new_[21156]_  = ~A202 & \new_[21155]_ ;
  assign \new_[21159]_  = ~A300 & A269;
  assign \new_[21162]_  = ~A302 & ~A301;
  assign \new_[21163]_  = \new_[21162]_  & \new_[21159]_ ;
  assign \new_[21164]_  = \new_[21163]_  & \new_[21156]_ ;
  assign \new_[21168]_  = A167 & ~A168;
  assign \new_[21169]_  = ~A169 & \new_[21168]_ ;
  assign \new_[21173]_  = ~A200 & ~A199;
  assign \new_[21174]_  = A166 & \new_[21173]_ ;
  assign \new_[21175]_  = \new_[21174]_  & \new_[21169]_ ;
  assign \new_[21179]_  = ~A266 & A265;
  assign \new_[21180]_  = ~A202 & \new_[21179]_ ;
  assign \new_[21183]_  = ~A298 & A269;
  assign \new_[21186]_  = ~A301 & ~A299;
  assign \new_[21187]_  = \new_[21186]_  & \new_[21183]_ ;
  assign \new_[21188]_  = \new_[21187]_  & \new_[21180]_ ;
  assign \new_[21192]_  = ~A168 & ~A169;
  assign \new_[21193]_  = ~A170 & \new_[21192]_ ;
  assign \new_[21197]_  = ~A203 & ~A202;
  assign \new_[21198]_  = ~A201 & \new_[21197]_ ;
  assign \new_[21199]_  = \new_[21198]_  & \new_[21193]_ ;
  assign \new_[21203]_  = A269 & A266;
  assign \new_[21204]_  = ~A265 & \new_[21203]_ ;
  assign \new_[21207]_  = A299 & A298;
  assign \new_[21210]_  = ~A301 & ~A300;
  assign \new_[21211]_  = \new_[21210]_  & \new_[21207]_ ;
  assign \new_[21212]_  = \new_[21211]_  & \new_[21204]_ ;
  assign \new_[21216]_  = ~A168 & ~A169;
  assign \new_[21217]_  = ~A170 & \new_[21216]_ ;
  assign \new_[21221]_  = ~A203 & ~A202;
  assign \new_[21222]_  = ~A201 & \new_[21221]_ ;
  assign \new_[21223]_  = \new_[21222]_  & \new_[21217]_ ;
  assign \new_[21227]_  = A269 & ~A266;
  assign \new_[21228]_  = A265 & \new_[21227]_ ;
  assign \new_[21231]_  = A299 & A298;
  assign \new_[21234]_  = ~A301 & ~A300;
  assign \new_[21235]_  = \new_[21234]_  & \new_[21231]_ ;
  assign \new_[21236]_  = \new_[21235]_  & \new_[21228]_ ;
  assign \new_[21240]_  = ~A168 & ~A169;
  assign \new_[21241]_  = ~A170 & \new_[21240]_ ;
  assign \new_[21245]_  = ~A201 & A200;
  assign \new_[21246]_  = A199 & \new_[21245]_ ;
  assign \new_[21247]_  = \new_[21246]_  & \new_[21241]_ ;
  assign \new_[21251]_  = A267 & A265;
  assign \new_[21252]_  = ~A202 & \new_[21251]_ ;
  assign \new_[21255]_  = A299 & A298;
  assign \new_[21258]_  = ~A301 & ~A300;
  assign \new_[21259]_  = \new_[21258]_  & \new_[21255]_ ;
  assign \new_[21260]_  = \new_[21259]_  & \new_[21252]_ ;
  assign \new_[21264]_  = ~A168 & ~A169;
  assign \new_[21265]_  = ~A170 & \new_[21264]_ ;
  assign \new_[21269]_  = ~A201 & A200;
  assign \new_[21270]_  = A199 & \new_[21269]_ ;
  assign \new_[21271]_  = \new_[21270]_  & \new_[21265]_ ;
  assign \new_[21275]_  = A267 & A266;
  assign \new_[21276]_  = ~A202 & \new_[21275]_ ;
  assign \new_[21279]_  = A299 & A298;
  assign \new_[21282]_  = ~A301 & ~A300;
  assign \new_[21283]_  = \new_[21282]_  & \new_[21279]_ ;
  assign \new_[21284]_  = \new_[21283]_  & \new_[21276]_ ;
  assign \new_[21288]_  = ~A168 & ~A169;
  assign \new_[21289]_  = ~A170 & \new_[21288]_ ;
  assign \new_[21293]_  = ~A201 & A200;
  assign \new_[21294]_  = A199 & \new_[21293]_ ;
  assign \new_[21295]_  = \new_[21294]_  & \new_[21289]_ ;
  assign \new_[21299]_  = A266 & ~A265;
  assign \new_[21300]_  = ~A202 & \new_[21299]_ ;
  assign \new_[21303]_  = ~A300 & A269;
  assign \new_[21306]_  = ~A302 & ~A301;
  assign \new_[21307]_  = \new_[21306]_  & \new_[21303]_ ;
  assign \new_[21308]_  = \new_[21307]_  & \new_[21300]_ ;
  assign \new_[21312]_  = ~A168 & ~A169;
  assign \new_[21313]_  = ~A170 & \new_[21312]_ ;
  assign \new_[21317]_  = ~A201 & A200;
  assign \new_[21318]_  = A199 & \new_[21317]_ ;
  assign \new_[21319]_  = \new_[21318]_  & \new_[21313]_ ;
  assign \new_[21323]_  = A266 & ~A265;
  assign \new_[21324]_  = ~A202 & \new_[21323]_ ;
  assign \new_[21327]_  = ~A298 & A269;
  assign \new_[21330]_  = ~A301 & ~A299;
  assign \new_[21331]_  = \new_[21330]_  & \new_[21327]_ ;
  assign \new_[21332]_  = \new_[21331]_  & \new_[21324]_ ;
  assign \new_[21336]_  = ~A168 & ~A169;
  assign \new_[21337]_  = ~A170 & \new_[21336]_ ;
  assign \new_[21341]_  = ~A201 & A200;
  assign \new_[21342]_  = A199 & \new_[21341]_ ;
  assign \new_[21343]_  = \new_[21342]_  & \new_[21337]_ ;
  assign \new_[21347]_  = ~A266 & A265;
  assign \new_[21348]_  = ~A202 & \new_[21347]_ ;
  assign \new_[21351]_  = ~A300 & A269;
  assign \new_[21354]_  = ~A302 & ~A301;
  assign \new_[21355]_  = \new_[21354]_  & \new_[21351]_ ;
  assign \new_[21356]_  = \new_[21355]_  & \new_[21348]_ ;
  assign \new_[21360]_  = ~A168 & ~A169;
  assign \new_[21361]_  = ~A170 & \new_[21360]_ ;
  assign \new_[21365]_  = ~A201 & A200;
  assign \new_[21366]_  = A199 & \new_[21365]_ ;
  assign \new_[21367]_  = \new_[21366]_  & \new_[21361]_ ;
  assign \new_[21371]_  = ~A266 & A265;
  assign \new_[21372]_  = ~A202 & \new_[21371]_ ;
  assign \new_[21375]_  = ~A298 & A269;
  assign \new_[21378]_  = ~A301 & ~A299;
  assign \new_[21379]_  = \new_[21378]_  & \new_[21375]_ ;
  assign \new_[21380]_  = \new_[21379]_  & \new_[21372]_ ;
  assign \new_[21384]_  = ~A168 & ~A169;
  assign \new_[21385]_  = ~A170 & \new_[21384]_ ;
  assign \new_[21389]_  = A203 & A200;
  assign \new_[21390]_  = ~A199 & \new_[21389]_ ;
  assign \new_[21391]_  = \new_[21390]_  & \new_[21385]_ ;
  assign \new_[21395]_  = ~A267 & A266;
  assign \new_[21396]_  = A265 & \new_[21395]_ ;
  assign \new_[21399]_  = A298 & ~A268;
  assign \new_[21402]_  = A302 & ~A299;
  assign \new_[21403]_  = \new_[21402]_  & \new_[21399]_ ;
  assign \new_[21404]_  = \new_[21403]_  & \new_[21396]_ ;
  assign \new_[21408]_  = ~A168 & ~A169;
  assign \new_[21409]_  = ~A170 & \new_[21408]_ ;
  assign \new_[21413]_  = A203 & A200;
  assign \new_[21414]_  = ~A199 & \new_[21413]_ ;
  assign \new_[21415]_  = \new_[21414]_  & \new_[21409]_ ;
  assign \new_[21419]_  = ~A267 & A266;
  assign \new_[21420]_  = A265 & \new_[21419]_ ;
  assign \new_[21423]_  = ~A298 & ~A268;
  assign \new_[21426]_  = A302 & A299;
  assign \new_[21427]_  = \new_[21426]_  & \new_[21423]_ ;
  assign \new_[21428]_  = \new_[21427]_  & \new_[21420]_ ;
  assign \new_[21432]_  = ~A168 & ~A169;
  assign \new_[21433]_  = ~A170 & \new_[21432]_ ;
  assign \new_[21437]_  = A203 & ~A200;
  assign \new_[21438]_  = A199 & \new_[21437]_ ;
  assign \new_[21439]_  = \new_[21438]_  & \new_[21433]_ ;
  assign \new_[21443]_  = ~A267 & A266;
  assign \new_[21444]_  = A265 & \new_[21443]_ ;
  assign \new_[21447]_  = A298 & ~A268;
  assign \new_[21450]_  = A302 & ~A299;
  assign \new_[21451]_  = \new_[21450]_  & \new_[21447]_ ;
  assign \new_[21452]_  = \new_[21451]_  & \new_[21444]_ ;
  assign \new_[21456]_  = ~A168 & ~A169;
  assign \new_[21457]_  = ~A170 & \new_[21456]_ ;
  assign \new_[21461]_  = A203 & ~A200;
  assign \new_[21462]_  = A199 & \new_[21461]_ ;
  assign \new_[21463]_  = \new_[21462]_  & \new_[21457]_ ;
  assign \new_[21467]_  = ~A267 & A266;
  assign \new_[21468]_  = A265 & \new_[21467]_ ;
  assign \new_[21471]_  = ~A298 & ~A268;
  assign \new_[21474]_  = A302 & A299;
  assign \new_[21475]_  = \new_[21474]_  & \new_[21471]_ ;
  assign \new_[21476]_  = \new_[21475]_  & \new_[21468]_ ;
  assign \new_[21480]_  = ~A168 & ~A169;
  assign \new_[21481]_  = ~A170 & \new_[21480]_ ;
  assign \new_[21485]_  = ~A202 & ~A200;
  assign \new_[21486]_  = ~A199 & \new_[21485]_ ;
  assign \new_[21487]_  = \new_[21486]_  & \new_[21481]_ ;
  assign \new_[21491]_  = A269 & A266;
  assign \new_[21492]_  = ~A265 & \new_[21491]_ ;
  assign \new_[21495]_  = A299 & A298;
  assign \new_[21498]_  = ~A301 & ~A300;
  assign \new_[21499]_  = \new_[21498]_  & \new_[21495]_ ;
  assign \new_[21500]_  = \new_[21499]_  & \new_[21492]_ ;
  assign \new_[21504]_  = ~A168 & ~A169;
  assign \new_[21505]_  = ~A170 & \new_[21504]_ ;
  assign \new_[21509]_  = ~A202 & ~A200;
  assign \new_[21510]_  = ~A199 & \new_[21509]_ ;
  assign \new_[21511]_  = \new_[21510]_  & \new_[21505]_ ;
  assign \new_[21515]_  = A269 & ~A266;
  assign \new_[21516]_  = A265 & \new_[21515]_ ;
  assign \new_[21519]_  = A299 & A298;
  assign \new_[21522]_  = ~A301 & ~A300;
  assign \new_[21523]_  = \new_[21522]_  & \new_[21519]_ ;
  assign \new_[21524]_  = \new_[21523]_  & \new_[21516]_ ;
  assign \new_[21528]_  = ~A166 & A167;
  assign \new_[21529]_  = A170 & \new_[21528]_ ;
  assign \new_[21532]_  = A200 & A199;
  assign \new_[21535]_  = ~A202 & ~A201;
  assign \new_[21536]_  = \new_[21535]_  & \new_[21532]_ ;
  assign \new_[21537]_  = \new_[21536]_  & \new_[21529]_ ;
  assign \new_[21541]_  = ~A267 & A266;
  assign \new_[21542]_  = A265 & \new_[21541]_ ;
  assign \new_[21545]_  = A298 & ~A268;
  assign \new_[21548]_  = A302 & ~A299;
  assign \new_[21549]_  = \new_[21548]_  & \new_[21545]_ ;
  assign \new_[21550]_  = \new_[21549]_  & \new_[21542]_ ;
  assign \new_[21554]_  = ~A166 & A167;
  assign \new_[21555]_  = A170 & \new_[21554]_ ;
  assign \new_[21558]_  = A200 & A199;
  assign \new_[21561]_  = ~A202 & ~A201;
  assign \new_[21562]_  = \new_[21561]_  & \new_[21558]_ ;
  assign \new_[21563]_  = \new_[21562]_  & \new_[21555]_ ;
  assign \new_[21567]_  = ~A267 & A266;
  assign \new_[21568]_  = A265 & \new_[21567]_ ;
  assign \new_[21571]_  = ~A298 & ~A268;
  assign \new_[21574]_  = A302 & A299;
  assign \new_[21575]_  = \new_[21574]_  & \new_[21571]_ ;
  assign \new_[21576]_  = \new_[21575]_  & \new_[21568]_ ;
  assign \new_[21580]_  = A166 & ~A167;
  assign \new_[21581]_  = A170 & \new_[21580]_ ;
  assign \new_[21584]_  = A200 & A199;
  assign \new_[21587]_  = ~A202 & ~A201;
  assign \new_[21588]_  = \new_[21587]_  & \new_[21584]_ ;
  assign \new_[21589]_  = \new_[21588]_  & \new_[21581]_ ;
  assign \new_[21593]_  = ~A267 & A266;
  assign \new_[21594]_  = A265 & \new_[21593]_ ;
  assign \new_[21597]_  = A298 & ~A268;
  assign \new_[21600]_  = A302 & ~A299;
  assign \new_[21601]_  = \new_[21600]_  & \new_[21597]_ ;
  assign \new_[21602]_  = \new_[21601]_  & \new_[21594]_ ;
  assign \new_[21606]_  = A166 & ~A167;
  assign \new_[21607]_  = A170 & \new_[21606]_ ;
  assign \new_[21610]_  = A200 & A199;
  assign \new_[21613]_  = ~A202 & ~A201;
  assign \new_[21614]_  = \new_[21613]_  & \new_[21610]_ ;
  assign \new_[21615]_  = \new_[21614]_  & \new_[21607]_ ;
  assign \new_[21619]_  = ~A267 & A266;
  assign \new_[21620]_  = A265 & \new_[21619]_ ;
  assign \new_[21623]_  = ~A298 & ~A268;
  assign \new_[21626]_  = A302 & A299;
  assign \new_[21627]_  = \new_[21626]_  & \new_[21623]_ ;
  assign \new_[21628]_  = \new_[21627]_  & \new_[21620]_ ;
  assign \new_[21632]_  = ~A166 & ~A167;
  assign \new_[21633]_  = ~A169 & \new_[21632]_ ;
  assign \new_[21636]_  = A200 & A199;
  assign \new_[21639]_  = ~A202 & ~A201;
  assign \new_[21640]_  = \new_[21639]_  & \new_[21636]_ ;
  assign \new_[21641]_  = \new_[21640]_  & \new_[21633]_ ;
  assign \new_[21645]_  = A269 & A266;
  assign \new_[21646]_  = ~A265 & \new_[21645]_ ;
  assign \new_[21649]_  = A299 & A298;
  assign \new_[21652]_  = ~A301 & ~A300;
  assign \new_[21653]_  = \new_[21652]_  & \new_[21649]_ ;
  assign \new_[21654]_  = \new_[21653]_  & \new_[21646]_ ;
  assign \new_[21658]_  = ~A166 & ~A167;
  assign \new_[21659]_  = ~A169 & \new_[21658]_ ;
  assign \new_[21662]_  = A200 & A199;
  assign \new_[21665]_  = ~A202 & ~A201;
  assign \new_[21666]_  = \new_[21665]_  & \new_[21662]_ ;
  assign \new_[21667]_  = \new_[21666]_  & \new_[21659]_ ;
  assign \new_[21671]_  = A269 & ~A266;
  assign \new_[21672]_  = A265 & \new_[21671]_ ;
  assign \new_[21675]_  = A299 & A298;
  assign \new_[21678]_  = ~A301 & ~A300;
  assign \new_[21679]_  = \new_[21678]_  & \new_[21675]_ ;
  assign \new_[21680]_  = \new_[21679]_  & \new_[21672]_ ;
  assign \new_[21684]_  = A167 & ~A168;
  assign \new_[21685]_  = ~A169 & \new_[21684]_ ;
  assign \new_[21688]_  = ~A201 & A166;
  assign \new_[21691]_  = ~A203 & ~A202;
  assign \new_[21692]_  = \new_[21691]_  & \new_[21688]_ ;
  assign \new_[21693]_  = \new_[21692]_  & \new_[21685]_ ;
  assign \new_[21697]_  = A269 & A266;
  assign \new_[21698]_  = ~A265 & \new_[21697]_ ;
  assign \new_[21701]_  = A299 & A298;
  assign \new_[21704]_  = ~A301 & ~A300;
  assign \new_[21705]_  = \new_[21704]_  & \new_[21701]_ ;
  assign \new_[21706]_  = \new_[21705]_  & \new_[21698]_ ;
  assign \new_[21710]_  = A167 & ~A168;
  assign \new_[21711]_  = ~A169 & \new_[21710]_ ;
  assign \new_[21714]_  = ~A201 & A166;
  assign \new_[21717]_  = ~A203 & ~A202;
  assign \new_[21718]_  = \new_[21717]_  & \new_[21714]_ ;
  assign \new_[21719]_  = \new_[21718]_  & \new_[21711]_ ;
  assign \new_[21723]_  = A269 & ~A266;
  assign \new_[21724]_  = A265 & \new_[21723]_ ;
  assign \new_[21727]_  = A299 & A298;
  assign \new_[21730]_  = ~A301 & ~A300;
  assign \new_[21731]_  = \new_[21730]_  & \new_[21727]_ ;
  assign \new_[21732]_  = \new_[21731]_  & \new_[21724]_ ;
  assign \new_[21736]_  = A167 & ~A168;
  assign \new_[21737]_  = ~A169 & \new_[21736]_ ;
  assign \new_[21740]_  = A199 & A166;
  assign \new_[21743]_  = ~A201 & A200;
  assign \new_[21744]_  = \new_[21743]_  & \new_[21740]_ ;
  assign \new_[21745]_  = \new_[21744]_  & \new_[21737]_ ;
  assign \new_[21749]_  = A267 & A265;
  assign \new_[21750]_  = ~A202 & \new_[21749]_ ;
  assign \new_[21753]_  = A299 & A298;
  assign \new_[21756]_  = ~A301 & ~A300;
  assign \new_[21757]_  = \new_[21756]_  & \new_[21753]_ ;
  assign \new_[21758]_  = \new_[21757]_  & \new_[21750]_ ;
  assign \new_[21762]_  = A167 & ~A168;
  assign \new_[21763]_  = ~A169 & \new_[21762]_ ;
  assign \new_[21766]_  = A199 & A166;
  assign \new_[21769]_  = ~A201 & A200;
  assign \new_[21770]_  = \new_[21769]_  & \new_[21766]_ ;
  assign \new_[21771]_  = \new_[21770]_  & \new_[21763]_ ;
  assign \new_[21775]_  = A267 & A266;
  assign \new_[21776]_  = ~A202 & \new_[21775]_ ;
  assign \new_[21779]_  = A299 & A298;
  assign \new_[21782]_  = ~A301 & ~A300;
  assign \new_[21783]_  = \new_[21782]_  & \new_[21779]_ ;
  assign \new_[21784]_  = \new_[21783]_  & \new_[21776]_ ;
  assign \new_[21788]_  = A167 & ~A168;
  assign \new_[21789]_  = ~A169 & \new_[21788]_ ;
  assign \new_[21792]_  = A199 & A166;
  assign \new_[21795]_  = ~A201 & A200;
  assign \new_[21796]_  = \new_[21795]_  & \new_[21792]_ ;
  assign \new_[21797]_  = \new_[21796]_  & \new_[21789]_ ;
  assign \new_[21801]_  = A266 & ~A265;
  assign \new_[21802]_  = ~A202 & \new_[21801]_ ;
  assign \new_[21805]_  = ~A300 & A269;
  assign \new_[21808]_  = ~A302 & ~A301;
  assign \new_[21809]_  = \new_[21808]_  & \new_[21805]_ ;
  assign \new_[21810]_  = \new_[21809]_  & \new_[21802]_ ;
  assign \new_[21814]_  = A167 & ~A168;
  assign \new_[21815]_  = ~A169 & \new_[21814]_ ;
  assign \new_[21818]_  = A199 & A166;
  assign \new_[21821]_  = ~A201 & A200;
  assign \new_[21822]_  = \new_[21821]_  & \new_[21818]_ ;
  assign \new_[21823]_  = \new_[21822]_  & \new_[21815]_ ;
  assign \new_[21827]_  = A266 & ~A265;
  assign \new_[21828]_  = ~A202 & \new_[21827]_ ;
  assign \new_[21831]_  = ~A298 & A269;
  assign \new_[21834]_  = ~A301 & ~A299;
  assign \new_[21835]_  = \new_[21834]_  & \new_[21831]_ ;
  assign \new_[21836]_  = \new_[21835]_  & \new_[21828]_ ;
  assign \new_[21840]_  = A167 & ~A168;
  assign \new_[21841]_  = ~A169 & \new_[21840]_ ;
  assign \new_[21844]_  = A199 & A166;
  assign \new_[21847]_  = ~A201 & A200;
  assign \new_[21848]_  = \new_[21847]_  & \new_[21844]_ ;
  assign \new_[21849]_  = \new_[21848]_  & \new_[21841]_ ;
  assign \new_[21853]_  = ~A266 & A265;
  assign \new_[21854]_  = ~A202 & \new_[21853]_ ;
  assign \new_[21857]_  = ~A300 & A269;
  assign \new_[21860]_  = ~A302 & ~A301;
  assign \new_[21861]_  = \new_[21860]_  & \new_[21857]_ ;
  assign \new_[21862]_  = \new_[21861]_  & \new_[21854]_ ;
  assign \new_[21866]_  = A167 & ~A168;
  assign \new_[21867]_  = ~A169 & \new_[21866]_ ;
  assign \new_[21870]_  = A199 & A166;
  assign \new_[21873]_  = ~A201 & A200;
  assign \new_[21874]_  = \new_[21873]_  & \new_[21870]_ ;
  assign \new_[21875]_  = \new_[21874]_  & \new_[21867]_ ;
  assign \new_[21879]_  = ~A266 & A265;
  assign \new_[21880]_  = ~A202 & \new_[21879]_ ;
  assign \new_[21883]_  = ~A298 & A269;
  assign \new_[21886]_  = ~A301 & ~A299;
  assign \new_[21887]_  = \new_[21886]_  & \new_[21883]_ ;
  assign \new_[21888]_  = \new_[21887]_  & \new_[21880]_ ;
  assign \new_[21892]_  = A167 & ~A168;
  assign \new_[21893]_  = ~A169 & \new_[21892]_ ;
  assign \new_[21896]_  = ~A199 & A166;
  assign \new_[21899]_  = A203 & A200;
  assign \new_[21900]_  = \new_[21899]_  & \new_[21896]_ ;
  assign \new_[21901]_  = \new_[21900]_  & \new_[21893]_ ;
  assign \new_[21905]_  = ~A267 & A266;
  assign \new_[21906]_  = A265 & \new_[21905]_ ;
  assign \new_[21909]_  = A298 & ~A268;
  assign \new_[21912]_  = A302 & ~A299;
  assign \new_[21913]_  = \new_[21912]_  & \new_[21909]_ ;
  assign \new_[21914]_  = \new_[21913]_  & \new_[21906]_ ;
  assign \new_[21918]_  = A167 & ~A168;
  assign \new_[21919]_  = ~A169 & \new_[21918]_ ;
  assign \new_[21922]_  = ~A199 & A166;
  assign \new_[21925]_  = A203 & A200;
  assign \new_[21926]_  = \new_[21925]_  & \new_[21922]_ ;
  assign \new_[21927]_  = \new_[21926]_  & \new_[21919]_ ;
  assign \new_[21931]_  = ~A267 & A266;
  assign \new_[21932]_  = A265 & \new_[21931]_ ;
  assign \new_[21935]_  = ~A298 & ~A268;
  assign \new_[21938]_  = A302 & A299;
  assign \new_[21939]_  = \new_[21938]_  & \new_[21935]_ ;
  assign \new_[21940]_  = \new_[21939]_  & \new_[21932]_ ;
  assign \new_[21944]_  = A167 & ~A168;
  assign \new_[21945]_  = ~A169 & \new_[21944]_ ;
  assign \new_[21948]_  = A199 & A166;
  assign \new_[21951]_  = A203 & ~A200;
  assign \new_[21952]_  = \new_[21951]_  & \new_[21948]_ ;
  assign \new_[21953]_  = \new_[21952]_  & \new_[21945]_ ;
  assign \new_[21957]_  = ~A267 & A266;
  assign \new_[21958]_  = A265 & \new_[21957]_ ;
  assign \new_[21961]_  = A298 & ~A268;
  assign \new_[21964]_  = A302 & ~A299;
  assign \new_[21965]_  = \new_[21964]_  & \new_[21961]_ ;
  assign \new_[21966]_  = \new_[21965]_  & \new_[21958]_ ;
  assign \new_[21970]_  = A167 & ~A168;
  assign \new_[21971]_  = ~A169 & \new_[21970]_ ;
  assign \new_[21974]_  = A199 & A166;
  assign \new_[21977]_  = A203 & ~A200;
  assign \new_[21978]_  = \new_[21977]_  & \new_[21974]_ ;
  assign \new_[21979]_  = \new_[21978]_  & \new_[21971]_ ;
  assign \new_[21983]_  = ~A267 & A266;
  assign \new_[21984]_  = A265 & \new_[21983]_ ;
  assign \new_[21987]_  = ~A298 & ~A268;
  assign \new_[21990]_  = A302 & A299;
  assign \new_[21991]_  = \new_[21990]_  & \new_[21987]_ ;
  assign \new_[21992]_  = \new_[21991]_  & \new_[21984]_ ;
  assign \new_[21996]_  = A167 & ~A168;
  assign \new_[21997]_  = ~A169 & \new_[21996]_ ;
  assign \new_[22000]_  = ~A199 & A166;
  assign \new_[22003]_  = ~A202 & ~A200;
  assign \new_[22004]_  = \new_[22003]_  & \new_[22000]_ ;
  assign \new_[22005]_  = \new_[22004]_  & \new_[21997]_ ;
  assign \new_[22009]_  = A269 & A266;
  assign \new_[22010]_  = ~A265 & \new_[22009]_ ;
  assign \new_[22013]_  = A299 & A298;
  assign \new_[22016]_  = ~A301 & ~A300;
  assign \new_[22017]_  = \new_[22016]_  & \new_[22013]_ ;
  assign \new_[22018]_  = \new_[22017]_  & \new_[22010]_ ;
  assign \new_[22022]_  = A167 & ~A168;
  assign \new_[22023]_  = ~A169 & \new_[22022]_ ;
  assign \new_[22026]_  = ~A199 & A166;
  assign \new_[22029]_  = ~A202 & ~A200;
  assign \new_[22030]_  = \new_[22029]_  & \new_[22026]_ ;
  assign \new_[22031]_  = \new_[22030]_  & \new_[22023]_ ;
  assign \new_[22035]_  = A269 & ~A266;
  assign \new_[22036]_  = A265 & \new_[22035]_ ;
  assign \new_[22039]_  = A299 & A298;
  assign \new_[22042]_  = ~A301 & ~A300;
  assign \new_[22043]_  = \new_[22042]_  & \new_[22039]_ ;
  assign \new_[22044]_  = \new_[22043]_  & \new_[22036]_ ;
  assign \new_[22048]_  = ~A168 & ~A169;
  assign \new_[22049]_  = ~A170 & \new_[22048]_ ;
  assign \new_[22052]_  = A200 & A199;
  assign \new_[22055]_  = ~A202 & ~A201;
  assign \new_[22056]_  = \new_[22055]_  & \new_[22052]_ ;
  assign \new_[22057]_  = \new_[22056]_  & \new_[22049]_ ;
  assign \new_[22061]_  = A269 & A266;
  assign \new_[22062]_  = ~A265 & \new_[22061]_ ;
  assign \new_[22065]_  = A299 & A298;
  assign \new_[22068]_  = ~A301 & ~A300;
  assign \new_[22069]_  = \new_[22068]_  & \new_[22065]_ ;
  assign \new_[22070]_  = \new_[22069]_  & \new_[22062]_ ;
  assign \new_[22074]_  = ~A168 & ~A169;
  assign \new_[22075]_  = ~A170 & \new_[22074]_ ;
  assign \new_[22078]_  = A200 & A199;
  assign \new_[22081]_  = ~A202 & ~A201;
  assign \new_[22082]_  = \new_[22081]_  & \new_[22078]_ ;
  assign \new_[22083]_  = \new_[22082]_  & \new_[22075]_ ;
  assign \new_[22087]_  = A269 & ~A266;
  assign \new_[22088]_  = A265 & \new_[22087]_ ;
  assign \new_[22091]_  = A299 & A298;
  assign \new_[22094]_  = ~A301 & ~A300;
  assign \new_[22095]_  = \new_[22094]_  & \new_[22091]_ ;
  assign \new_[22096]_  = \new_[22095]_  & \new_[22088]_ ;
  assign \new_[22100]_  = A167 & ~A168;
  assign \new_[22101]_  = ~A169 & \new_[22100]_ ;
  assign \new_[22104]_  = A199 & A166;
  assign \new_[22107]_  = ~A201 & A200;
  assign \new_[22108]_  = \new_[22107]_  & \new_[22104]_ ;
  assign \new_[22109]_  = \new_[22108]_  & \new_[22101]_ ;
  assign \new_[22112]_  = ~A265 & ~A202;
  assign \new_[22115]_  = A269 & A266;
  assign \new_[22116]_  = \new_[22115]_  & \new_[22112]_ ;
  assign \new_[22119]_  = A299 & A298;
  assign \new_[22122]_  = ~A301 & ~A300;
  assign \new_[22123]_  = \new_[22122]_  & \new_[22119]_ ;
  assign \new_[22124]_  = \new_[22123]_  & \new_[22116]_ ;
  assign \new_[22128]_  = A167 & ~A168;
  assign \new_[22129]_  = ~A169 & \new_[22128]_ ;
  assign \new_[22132]_  = A199 & A166;
  assign \new_[22135]_  = ~A201 & A200;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22132]_ ;
  assign \new_[22137]_  = \new_[22136]_  & \new_[22129]_ ;
  assign \new_[22140]_  = A265 & ~A202;
  assign \new_[22143]_  = A269 & ~A266;
  assign \new_[22144]_  = \new_[22143]_  & \new_[22140]_ ;
  assign \new_[22147]_  = A299 & A298;
  assign \new_[22150]_  = ~A301 & ~A300;
  assign \new_[22151]_  = \new_[22150]_  & \new_[22147]_ ;
  assign \new_[22152]_  = \new_[22151]_  & \new_[22144]_ ;
endmodule


