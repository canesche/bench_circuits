// Benchmark "testing" written by ABC on Thu Oct  8 22:17:00 2020

module testing ( 
    B9278, B9277, B9276, B9275, B9274, B9245, B9244, B9243, B9242, B9241,
    B9212, B9211, B9210, B9209, B9208, B9179, B9178, B9177, B9176, B9175,
    B9146, B9145, B9144, B9143, B9142, B9113, B9112, B9111, B9110, B9109,
    B9080, B9079, B9078, B9077, B9076, B9047, B9046, B9045, B9044, B9043,
    B9014, B9013, B9012, B9011, B9010, B8981, B8980, B8979, B8978, B8977,
    B8948, B8947, B8946, B8945, B8944, B8915, B8914, B8913, B8912, B8911,
    B8882, B8881, B8880, B8879, B8878, B8849, B8848, B8847, B8846, B8845,
    B8816, B8815, B8814, B8813, B8812, B8783, B8782, B8781, B8780, B8779,
    B8750, B8749, B8748, B8747, B8746, B8717, B8716, B8715, B8714, B8713,
    B8684, B8683, B8682, B8681, B8680, B8651, B8650, B8649, B8648, B8647,
    B8618, B8617, B8616, B8615, B8614, B8585, B8584, B8583, B8582, B8581,
    B8552, B8551, B8550, B8549, B8548, B8519, B8518, B8517, B8516, B8515,
    B8486, B8485, B8484, B8483, B8482, B8453, B8452, B8451, B8450, B8449,
    B8420, B8419, B8418, B8417, B8416, B8387, B8386, B8385, B8384, B8383,
    B8354, B8353, B8352, B8351, B8350, B8321, B8320, B8319, B8318, B8317,
    B8288, B8287, B8286, B8285, B8284, B8255, B8254, B8253, B8252, B8251,
    B8222, B8221, B8220, B8219, B8218, B8189, B8188, B8187, B8186, B8185,
    B8156, B8155, B8154, B8153, B8152, B8123, B8122, B8121, B8120, B8119,
    B8090, B8089, B8088, B8087, B8086, B8057, B8056, B8055, B8054, B8053,
    B8024, B8023, B8022, B8021, B8020, B7991, B7990, B7989, B7988, B7987,
    B7958, B7957, B7956, B7955, B7954, B7925, B7924, B7923, B7922, B7921,
    B7892, B7891, B7890, B7889, B7888, B7859, B7858, B7857, B7856, B7855,
    B7826, B7825, B7824, B7823, B7822, B7793, B7792, B7791, B7790, B7789,
    B7760, B7759, B7758, B7757, B7756, B7727, B7726, B7725, B7724, B7723,
    B7694, B7693, B7692, B7691, B7690, B7661, B7660, B7659, B7658, B7657,
    B7628, B7627, B7626, B7625, B7624, B7595, B7594, B7593, B7592, B7591,
    B7562, B7561, B7560, B7559, B7558, B7529, B7528, B7527, B7526, B7525,
    B7496, B7495, B7494, B7493, B7492, B7463, B7462, B7461, B7460, B7459,
    B7430, B7429, B7428, B7427, B7426, B7397, B7396, B7395, B7394, B7393,
    B7364, B7363, B7362, B7361, B7360, B7331, B7330, B7329, B7328, B7327,
    B7298, B7297, B7296, B7295, B7294, B7265, B7264, B7263, B7262, B7261,
    B7232, B7231, B7230, B7229, B7228, B7199, B7198, B7197, B7196, B7195,
    B7166, B7165, B7164, B7163, B7162, B7133, B7132, B7131, B7130, B7129,
    B7100, B7099, B7098, B7097, B7096, B7067, B7066, B7065, B7064, B7063,
    B7034, B7033, B7032, B7031, B7030, B7001, B7000, B6999, B6998, B6997,
    B6968, B6967, B6966, B6965, B6964, B6935, B6934, B6933, B6932, B6931,
    B6902, B6901, B6900, B6899, B6898, B6869, B6868, B6867, B6866, B6865,
    B6836, B6835, B6834, B6833, B6832, B6803, B6802, B6801, B6800, B6799,
    B6770, B6769, B6768, B6767, B6766, B6737, B6736, B6735, B6734, B6733,
    B6704, B6703, B6702, B6701, B6700, B6671, B6670, B6669, B6668, B6667,
    B6638, B6637, B6636, B6635, B6634, B6605, B6604, B6603, B6602, B6601,
    B6572, B6571, B6570, B6569, B6568, B6539, B6538, B6537, B6536, B6535,
    B6506, B6505, B6504, B6503, B6502, B6473, B6472, B6471, B6470, B6469,
    B6440, B6439, B6438, B6437, B6436, B6407, B6406, B6405, B6404, B6403,
    B6374, B6373, B6372, B6371, B6370, B6341, B6340, B6339, B6338, B6337,
    B6308, B6307, B6306, B6305, B6304, B6275, B6274, B6273, B6272, B6271,
    B6242, B6241, B6240, B6239, B6238, B6209, B6208, B6207, B6206, B6205,
    B6176, B6175, B6174, B6173, B6172, B6143, B6142, B6141, B6140, B6139,
    B6110, B6109, B6108, B6107, B6106, B6077, B6076, B6075, B6074, B6073,
    B6044, B6043, B6042, B6041, B6040, B6011, B6010, B6009, B6008, B6007,
    B5978, B5977, B5976, B5975, B5974, B5945, B5944, B5943, B5942, B5941,
    B5912, B5911, B5910, B5909, B5908, B5879, B5878, B5877, B5876, B5875,
    B5846, B5845, B5844, B5843, B5842, B5813, B5812, B5811, B5810, B5809,
    B5780, B5779, B5778, B5777, B5776, B5747, B5746, B5745, B5744, B5743,
    B5714, B5713, B5712, B5711, B5710, B5681, B5680, B5679, B5678, B5677,
    B5648, B5647, B5646, B5645, B5644, B5615, B5614, B5613, B5612, B5611,
    B5582, B5581, B5580, B5579, B5578, B5549, B5548, B5547, B5546, B5545,
    B5516, B5515, B5514, B5513, B5512, B5483, B5482, B5481, B5480, B5479,
    B5450, B5449, B5448, B5447, B5446, B5417, B5416, B5415, B5414, B5413,
    B5384, B5383, B5382, B5381, B5380, B5351, B5350, B5349, B5348, B5347,
    B5318, B5317, B5316, B5315, B5314, B5285, B5284, B5283, B5282, B5281,
    B5252, B5251, B5250, B5249, B5248, B5219, B5218, B5217, B5216, B5215,
    B5182, B5183, B5184, B5185, B5186,
    A6907, A6906, A6905, A6904, A6903, A6874, A6873, A6872, A6871, A6870,
    A6841, A6840, A6839, A6838, A6837, A6808, A6807, A6806, A6805, A6804,
    A6775, A6774, A6773, A6772, A6771, A6742, A6741, A6740, A6739, A6738,
    A6709, A6708, A6707, A6706, A6705, A6676, A6675, A6674, A6673, A6672,
    A6643, A6642, A6641, A6640, A6639, A6610, A6609, A6608, A6607, A6606,
    A6577, A6576, A6575, A6574, A6573, A6544, A6543, A6542, A6541, A6540,
    A6511, A6510, A6509, A6508, A6507, A6478, A6477, A6476, A6475, A6474,
    A6445, A6444, A6443, A6442, A6441, A6412, A6411, A6410, A6409, A6408,
    A6379, A6378, A6377, A6376, A6375, A6346, A6345, A6344, A6343, A6342,
    A6313, A6312, A6311, A6310, A6309, A6280, A6279, A6278, A6277, A6276,
    A6247, A6246, A6245, A6244, A6243, A6214, A6213, A6212, A6211, A6210,
    A6181, A6180, A6179, A6178, A6177, A6148, A6147, A6146, A6145, A6144,
    A6115, A6114, A6113, A6112, A6111, A6082, A6081, A6080, A6079, A6078,
    A6049, A6048, A6047, A6046, A6045, A6016, A6015, A6014, A6013, A6012,
    A5983, A5982, A5981, A5980, A5979, A5950, A5949, A5948, A5947, A5946,
    A5917, A5916, A5915, A5914, A5913, A5884, A5883, A5882, A5881, A5880,
    A5851, A5850, A5849, A5848, A5847, A5818, A5817, A5816, A5815, A5814,
    A5785, A5784, A5783, A5782, A5781, A5752, A5751, A5750, A5749, A5748,
    A5719, A5718, A5717, A5716, A5715, A5686, A5685, A5684, A5683, A5682,
    A5653, A5652, A5651, A5650, A5649, A5620, A5619, A5618, A5617, A5616,
    A5587, A5586, A5585, A5584, A5583, A5554, A5553, A5552, A5551, A5550,
    A5521, A5520, A5519, A5518, A5517, A5488, A5487, A5486, A5485, A5484,
    A5455, A5454, A5453, A5452, A5451, A5422, A5421, A5420, A5419, A5418,
    A5389, A5388, A5387, A5386, A5385, A5356, A5355, A5354, A5353, A5352,
    A5323, A5322, A5321, A5320, A5319, A5290, A5289, A5288, A5287, A5286,
    A5257, A5256, A5255, A5254, A5253, A5224, A5223, A5222, A5221, A5220,
    A5191, A5190, A5189, A5188, A5187, A5158, A5157, A5156, A5155, A5154,
    A5125, A5124, A5123, A5122, A5121, A5092, A5091, A5090, A5089, A5088,
    A5059, A5058, A5057, A5056, A5055, A5026, A5025, A5024, A5023, A5022,
    A4993, A4992, A4991, A4990, A4989, A4960, A4959, A4958, A4957, A4956,
    A4927, A4926, A4925, A4924, A4923, A4894, A4893, A4892, A4891, A4890,
    A4861, A4860, A4859, A4858, A4857, A4828, A4827, A4826, A4825, A4824,
    A4795, A4794, A4793, A4792, A4791, A4762, A4761, A4760, A4759, A4758,
    A4729, A4728, A4727, A4726, A4725, A4696, A4695, A4694, A4693, A4692,
    A4663, A4662, A4661, A4660, A4659, A4630, A4629, A4628, A4627, A4626,
    A4597, A4596, A4595, A4594, A4593, A4564, A4563, A4562, A4561, A4560,
    A4531, A4530, A4529, A4528, A4527, A4498, A4497, A4496, A4495, A4494,
    A4465, A4464, A4463, A4462, A4461, A4432, A4431, A4430, A4429, A4428,
    A4399, A4398, A4397, A4396, A4395, A4366, A4365, A4364, A4363, A4362,
    A4333, A4332, A4331, A4330, A4329, A4300, A4299, A4298, A4297, A4296,
    A4267, A4266, A4265, A4264, A4263, A4234, A4233, A4232, A4231, A4230,
    A4201, A4200, A4199, A4198, A4197, A4168, A4167, A4166, A4165, A4164,
    A4135, A4134, A4133, A4132, A4131, A4102, A4101, A4100, A4099, A4098,
    A4069, A4068, A4067, A4066, A4065, A4036, A4035, A4034, A4033, A4032,
    A4003, A4002, A4001, A4000, A3999, A3970, A3969, A3968, A3967, A3966,
    A3937, A3936, A3935, A3934, A3933, A3904, A3903, A3902, A3901, A3900,
    A3871, A3870, A3869, A3868, A3867, A3838, A3837, A3836, A3835, A3834,
    A3805, A3804, A3803, A3802, A3801, A3772, A3771, A3770, A3769, A3768,
    A3739, A3738, A3737, A3736, A3735, A3706, A3705, A3704, A3703, A3702,
    A3673, A3672, A3671, A3670, A3669, A3640, A3639, A3638, A3637, A3636,
    A3607, A3606, A3605, A3604, A3603, A3574, A3573, A3572, A3571, A3570,
    A3541, A3540, A3539, A3538, A3537, A3508, A3507, A3506, A3505, A3504,
    A3475, A3474, A3473, A3472, A3471, A3442, A3441, A3440, A3439, A3438,
    A3409, A3408, A3407, A3406, A3405, A3376, A3375, A3374, A3373, A3372,
    A3343, A3342, A3341, A3340, A3339, A3310, A3309, A3308, A3307, A3306,
    A3277, A3276, A3275, A3274, A3273, A3244, A3243, A3242, A3241, A3240,
    A3211, A3210, A3209, A3208, A3207, A3178, A3177, A3176, A3175, A3174,
    A3145, A3144, A3143, A3142, A3141, A3112, A3111, A3110, A3109, A3108,
    A3079, A3078, A3077, A3076, A3075, A3046, A3045, A3044, A3043, A3042,
    A3013, A3012, A3011, A3010, A3009, A2980, A2979, A2978, A2977, A2976,
    A2947, A2946, A2945, A2944, A2943, A2914, A2913, A2912, A2911, A2910,
    A2881, A2880, A2879, A2878, A2877, A2848, A2847, A2846, A2845, A2844,
    A2811, A2812, A2813, A2814, A2815  );
  input  B9278, B9277, B9276, B9275, B9274, B9245, B9244, B9243, B9242,
    B9241, B9212, B9211, B9210, B9209, B9208, B9179, B9178, B9177, B9176,
    B9175, B9146, B9145, B9144, B9143, B9142, B9113, B9112, B9111, B9110,
    B9109, B9080, B9079, B9078, B9077, B9076, B9047, B9046, B9045, B9044,
    B9043, B9014, B9013, B9012, B9011, B9010, B8981, B8980, B8979, B8978,
    B8977, B8948, B8947, B8946, B8945, B8944, B8915, B8914, B8913, B8912,
    B8911, B8882, B8881, B8880, B8879, B8878, B8849, B8848, B8847, B8846,
    B8845, B8816, B8815, B8814, B8813, B8812, B8783, B8782, B8781, B8780,
    B8779, B8750, B8749, B8748, B8747, B8746, B8717, B8716, B8715, B8714,
    B8713, B8684, B8683, B8682, B8681, B8680, B8651, B8650, B8649, B8648,
    B8647, B8618, B8617, B8616, B8615, B8614, B8585, B8584, B8583, B8582,
    B8581, B8552, B8551, B8550, B8549, B8548, B8519, B8518, B8517, B8516,
    B8515, B8486, B8485, B8484, B8483, B8482, B8453, B8452, B8451, B8450,
    B8449, B8420, B8419, B8418, B8417, B8416, B8387, B8386, B8385, B8384,
    B8383, B8354, B8353, B8352, B8351, B8350, B8321, B8320, B8319, B8318,
    B8317, B8288, B8287, B8286, B8285, B8284, B8255, B8254, B8253, B8252,
    B8251, B8222, B8221, B8220, B8219, B8218, B8189, B8188, B8187, B8186,
    B8185, B8156, B8155, B8154, B8153, B8152, B8123, B8122, B8121, B8120,
    B8119, B8090, B8089, B8088, B8087, B8086, B8057, B8056, B8055, B8054,
    B8053, B8024, B8023, B8022, B8021, B8020, B7991, B7990, B7989, B7988,
    B7987, B7958, B7957, B7956, B7955, B7954, B7925, B7924, B7923, B7922,
    B7921, B7892, B7891, B7890, B7889, B7888, B7859, B7858, B7857, B7856,
    B7855, B7826, B7825, B7824, B7823, B7822, B7793, B7792, B7791, B7790,
    B7789, B7760, B7759, B7758, B7757, B7756, B7727, B7726, B7725, B7724,
    B7723, B7694, B7693, B7692, B7691, B7690, B7661, B7660, B7659, B7658,
    B7657, B7628, B7627, B7626, B7625, B7624, B7595, B7594, B7593, B7592,
    B7591, B7562, B7561, B7560, B7559, B7558, B7529, B7528, B7527, B7526,
    B7525, B7496, B7495, B7494, B7493, B7492, B7463, B7462, B7461, B7460,
    B7459, B7430, B7429, B7428, B7427, B7426, B7397, B7396, B7395, B7394,
    B7393, B7364, B7363, B7362, B7361, B7360, B7331, B7330, B7329, B7328,
    B7327, B7298, B7297, B7296, B7295, B7294, B7265, B7264, B7263, B7262,
    B7261, B7232, B7231, B7230, B7229, B7228, B7199, B7198, B7197, B7196,
    B7195, B7166, B7165, B7164, B7163, B7162, B7133, B7132, B7131, B7130,
    B7129, B7100, B7099, B7098, B7097, B7096, B7067, B7066, B7065, B7064,
    B7063, B7034, B7033, B7032, B7031, B7030, B7001, B7000, B6999, B6998,
    B6997, B6968, B6967, B6966, B6965, B6964, B6935, B6934, B6933, B6932,
    B6931, B6902, B6901, B6900, B6899, B6898, B6869, B6868, B6867, B6866,
    B6865, B6836, B6835, B6834, B6833, B6832, B6803, B6802, B6801, B6800,
    B6799, B6770, B6769, B6768, B6767, B6766, B6737, B6736, B6735, B6734,
    B6733, B6704, B6703, B6702, B6701, B6700, B6671, B6670, B6669, B6668,
    B6667, B6638, B6637, B6636, B6635, B6634, B6605, B6604, B6603, B6602,
    B6601, B6572, B6571, B6570, B6569, B6568, B6539, B6538, B6537, B6536,
    B6535, B6506, B6505, B6504, B6503, B6502, B6473, B6472, B6471, B6470,
    B6469, B6440, B6439, B6438, B6437, B6436, B6407, B6406, B6405, B6404,
    B6403, B6374, B6373, B6372, B6371, B6370, B6341, B6340, B6339, B6338,
    B6337, B6308, B6307, B6306, B6305, B6304, B6275, B6274, B6273, B6272,
    B6271, B6242, B6241, B6240, B6239, B6238, B6209, B6208, B6207, B6206,
    B6205, B6176, B6175, B6174, B6173, B6172, B6143, B6142, B6141, B6140,
    B6139, B6110, B6109, B6108, B6107, B6106, B6077, B6076, B6075, B6074,
    B6073, B6044, B6043, B6042, B6041, B6040, B6011, B6010, B6009, B6008,
    B6007, B5978, B5977, B5976, B5975, B5974, B5945, B5944, B5943, B5942,
    B5941, B5912, B5911, B5910, B5909, B5908, B5879, B5878, B5877, B5876,
    B5875, B5846, B5845, B5844, B5843, B5842, B5813, B5812, B5811, B5810,
    B5809, B5780, B5779, B5778, B5777, B5776, B5747, B5746, B5745, B5744,
    B5743, B5714, B5713, B5712, B5711, B5710, B5681, B5680, B5679, B5678,
    B5677, B5648, B5647, B5646, B5645, B5644, B5615, B5614, B5613, B5612,
    B5611, B5582, B5581, B5580, B5579, B5578, B5549, B5548, B5547, B5546,
    B5545, B5516, B5515, B5514, B5513, B5512, B5483, B5482, B5481, B5480,
    B5479, B5450, B5449, B5448, B5447, B5446, B5417, B5416, B5415, B5414,
    B5413, B5384, B5383, B5382, B5381, B5380, B5351, B5350, B5349, B5348,
    B5347, B5318, B5317, B5316, B5315, B5314, B5285, B5284, B5283, B5282,
    B5281, B5252, B5251, B5250, B5249, B5248, B5219, B5218, B5217, B5216,
    B5215, B5182, B5183, B5184, B5185, B5186;
  output A6907, A6906, A6905, A6904, A6903, A6874, A6873, A6872, A6871, A6870,
    A6841, A6840, A6839, A6838, A6837, A6808, A6807, A6806, A6805, A6804,
    A6775, A6774, A6773, A6772, A6771, A6742, A6741, A6740, A6739, A6738,
    A6709, A6708, A6707, A6706, A6705, A6676, A6675, A6674, A6673, A6672,
    A6643, A6642, A6641, A6640, A6639, A6610, A6609, A6608, A6607, A6606,
    A6577, A6576, A6575, A6574, A6573, A6544, A6543, A6542, A6541, A6540,
    A6511, A6510, A6509, A6508, A6507, A6478, A6477, A6476, A6475, A6474,
    A6445, A6444, A6443, A6442, A6441, A6412, A6411, A6410, A6409, A6408,
    A6379, A6378, A6377, A6376, A6375, A6346, A6345, A6344, A6343, A6342,
    A6313, A6312, A6311, A6310, A6309, A6280, A6279, A6278, A6277, A6276,
    A6247, A6246, A6245, A6244, A6243, A6214, A6213, A6212, A6211, A6210,
    A6181, A6180, A6179, A6178, A6177, A6148, A6147, A6146, A6145, A6144,
    A6115, A6114, A6113, A6112, A6111, A6082, A6081, A6080, A6079, A6078,
    A6049, A6048, A6047, A6046, A6045, A6016, A6015, A6014, A6013, A6012,
    A5983, A5982, A5981, A5980, A5979, A5950, A5949, A5948, A5947, A5946,
    A5917, A5916, A5915, A5914, A5913, A5884, A5883, A5882, A5881, A5880,
    A5851, A5850, A5849, A5848, A5847, A5818, A5817, A5816, A5815, A5814,
    A5785, A5784, A5783, A5782, A5781, A5752, A5751, A5750, A5749, A5748,
    A5719, A5718, A5717, A5716, A5715, A5686, A5685, A5684, A5683, A5682,
    A5653, A5652, A5651, A5650, A5649, A5620, A5619, A5618, A5617, A5616,
    A5587, A5586, A5585, A5584, A5583, A5554, A5553, A5552, A5551, A5550,
    A5521, A5520, A5519, A5518, A5517, A5488, A5487, A5486, A5485, A5484,
    A5455, A5454, A5453, A5452, A5451, A5422, A5421, A5420, A5419, A5418,
    A5389, A5388, A5387, A5386, A5385, A5356, A5355, A5354, A5353, A5352,
    A5323, A5322, A5321, A5320, A5319, A5290, A5289, A5288, A5287, A5286,
    A5257, A5256, A5255, A5254, A5253, A5224, A5223, A5222, A5221, A5220,
    A5191, A5190, A5189, A5188, A5187, A5158, A5157, A5156, A5155, A5154,
    A5125, A5124, A5123, A5122, A5121, A5092, A5091, A5090, A5089, A5088,
    A5059, A5058, A5057, A5056, A5055, A5026, A5025, A5024, A5023, A5022,
    A4993, A4992, A4991, A4990, A4989, A4960, A4959, A4958, A4957, A4956,
    A4927, A4926, A4925, A4924, A4923, A4894, A4893, A4892, A4891, A4890,
    A4861, A4860, A4859, A4858, A4857, A4828, A4827, A4826, A4825, A4824,
    A4795, A4794, A4793, A4792, A4791, A4762, A4761, A4760, A4759, A4758,
    A4729, A4728, A4727, A4726, A4725, A4696, A4695, A4694, A4693, A4692,
    A4663, A4662, A4661, A4660, A4659, A4630, A4629, A4628, A4627, A4626,
    A4597, A4596, A4595, A4594, A4593, A4564, A4563, A4562, A4561, A4560,
    A4531, A4530, A4529, A4528, A4527, A4498, A4497, A4496, A4495, A4494,
    A4465, A4464, A4463, A4462, A4461, A4432, A4431, A4430, A4429, A4428,
    A4399, A4398, A4397, A4396, A4395, A4366, A4365, A4364, A4363, A4362,
    A4333, A4332, A4331, A4330, A4329, A4300, A4299, A4298, A4297, A4296,
    A4267, A4266, A4265, A4264, A4263, A4234, A4233, A4232, A4231, A4230,
    A4201, A4200, A4199, A4198, A4197, A4168, A4167, A4166, A4165, A4164,
    A4135, A4134, A4133, A4132, A4131, A4102, A4101, A4100, A4099, A4098,
    A4069, A4068, A4067, A4066, A4065, A4036, A4035, A4034, A4033, A4032,
    A4003, A4002, A4001, A4000, A3999, A3970, A3969, A3968, A3967, A3966,
    A3937, A3936, A3935, A3934, A3933, A3904, A3903, A3902, A3901, A3900,
    A3871, A3870, A3869, A3868, A3867, A3838, A3837, A3836, A3835, A3834,
    A3805, A3804, A3803, A3802, A3801, A3772, A3771, A3770, A3769, A3768,
    A3739, A3738, A3737, A3736, A3735, A3706, A3705, A3704, A3703, A3702,
    A3673, A3672, A3671, A3670, A3669, A3640, A3639, A3638, A3637, A3636,
    A3607, A3606, A3605, A3604, A3603, A3574, A3573, A3572, A3571, A3570,
    A3541, A3540, A3539, A3538, A3537, A3508, A3507, A3506, A3505, A3504,
    A3475, A3474, A3473, A3472, A3471, A3442, A3441, A3440, A3439, A3438,
    A3409, A3408, A3407, A3406, A3405, A3376, A3375, A3374, A3373, A3372,
    A3343, A3342, A3341, A3340, A3339, A3310, A3309, A3308, A3307, A3306,
    A3277, A3276, A3275, A3274, A3273, A3244, A3243, A3242, A3241, A3240,
    A3211, A3210, A3209, A3208, A3207, A3178, A3177, A3176, A3175, A3174,
    A3145, A3144, A3143, A3142, A3141, A3112, A3111, A3110, A3109, A3108,
    A3079, A3078, A3077, A3076, A3075, A3046, A3045, A3044, A3043, A3042,
    A3013, A3012, A3011, A3010, A3009, A2980, A2979, A2978, A2977, A2976,
    A2947, A2946, A2945, A2944, A2943, A2914, A2913, A2912, A2911, A2910,
    A2881, A2880, A2879, A2878, A2877, A2848, A2847, A2846, A2845, A2844,
    A2811, A2812, A2813, A2814, A2815;
  wire new_B5214_, new_B5213_, new_B5212_, new_B5211_, new_B5210_,
    new_B5209_, new_B5208_, new_B5207_, new_B5206_, new_B5205_, new_B5204_,
    new_B5203_, new_B5202_, new_B5201_, new_B5200_, new_B5199_, new_B5198_,
    new_B5197_, new_B5196_, new_B5195_, new_B5194_, new_B5193_, new_B5192_,
    new_B5191_, new_B5190_, new_B5189_, new_B5188_, new_B5187_, new_B5220_,
    new_B5221_, new_B5222_, new_B5223_, new_B5224_, new_B5225_, new_B5226_,
    new_B5227_, new_B5228_, new_B5229_, new_B5230_, new_B5231_, new_B5232_,
    new_B5233_, new_B5234_, new_B5235_, new_B5236_, new_B5237_, new_B5238_,
    new_B5239_, new_B5240_, new_B5241_, new_B5242_, new_B5243_, new_B5244_,
    new_B5245_, new_B5246_, new_B5247_, new_B5253_, new_B5254_, new_B5255_,
    new_B5256_, new_B5257_, new_B5258_, new_B5259_, new_B5260_, new_B5261_,
    new_B5262_, new_B5263_, new_B5264_, new_B5265_, new_B5266_, new_B5267_,
    new_B5268_, new_B5269_, new_B5270_, new_B5271_, new_B5272_, new_B5273_,
    new_B5274_, new_B5275_, new_B5276_, new_B5277_, new_B5278_, new_B5279_,
    new_B5280_, new_B5286_, new_B5287_, new_B5288_, new_B5289_, new_B5290_,
    new_B5291_, new_B5292_, new_B5293_, new_B5294_, new_B5295_, new_B5296_,
    new_B5297_, new_B5298_, new_B5299_, new_B5300_, new_B5301_, new_B5302_,
    new_B5303_, new_B5304_, new_B5305_, new_B5306_, new_B5307_, new_B5308_,
    new_B5309_, new_B5310_, new_B5311_, new_B5312_, new_B5313_, new_B5319_,
    new_B5320_, new_B5321_, new_B5322_, new_B5323_, new_B5324_, new_B5325_,
    new_B5326_, new_B5327_, new_B5328_, new_B5329_, new_B5330_, new_B5331_,
    new_B5332_, new_B5333_, new_B5334_, new_B5335_, new_B5336_, new_B5337_,
    new_B5338_, new_B5339_, new_B5340_, new_B5341_, new_B5342_, new_B5343_,
    new_B5344_, new_B5345_, new_B5346_, new_B5352_, new_B5353_, new_B5354_,
    new_B5355_, new_B5356_, new_B5357_, new_B5358_, new_B5359_, new_B5360_,
    new_B5361_, new_B5362_, new_B5363_, new_B5364_, new_B5365_, new_B5366_,
    new_B5367_, new_B5368_, new_B5369_, new_B5370_, new_B5371_, new_B5372_,
    new_B5373_, new_B5374_, new_B5375_, new_B5376_, new_B5377_, new_B5378_,
    new_B5379_, new_B5385_, new_B5386_, new_B5387_, new_B5388_, new_B5389_,
    new_B5390_, new_B5391_, new_B5392_, new_B5393_, new_B5394_, new_B5395_,
    new_B5396_, new_B5397_, new_B5398_, new_B5399_, new_B5400_, new_B5401_,
    new_B5402_, new_B5403_, new_B5404_, new_B5405_, new_B5406_, new_B5407_,
    new_B5408_, new_B5409_, new_B5410_, new_B5411_, new_B5412_, new_B5418_,
    new_B5419_, new_B5420_, new_B5421_, new_B5422_, new_B5423_, new_B5424_,
    new_B5425_, new_B5426_, new_B5427_, new_B5428_, new_B5429_, new_B5430_,
    new_B5431_, new_B5432_, new_B5433_, new_B5434_, new_B5435_, new_B5436_,
    new_B5437_, new_B5438_, new_B5439_, new_B5440_, new_B5441_, new_B5442_,
    new_B5443_, new_B5444_, new_B5445_, new_B5451_, new_B5452_, new_B5453_,
    new_B5454_, new_B5455_, new_B5456_, new_B5457_, new_B5458_, new_B5459_,
    new_B5460_, new_B5461_, new_B5462_, new_B5463_, new_B5464_, new_B5465_,
    new_B5466_, new_B5467_, new_B5468_, new_B5469_, new_B5470_, new_B5471_,
    new_B5472_, new_B5473_, new_B5474_, new_B5475_, new_B5476_, new_B5477_,
    new_B5478_, new_B5484_, new_B5485_, new_B5486_, new_B5487_, new_B5488_,
    new_B5489_, new_B5490_, new_B5491_, new_B5492_, new_B5493_, new_B5494_,
    new_B5495_, new_B5496_, new_B5497_, new_B5498_, new_B5499_, new_B5500_,
    new_B5501_, new_B5502_, new_B5503_, new_B5504_, new_B5505_, new_B5506_,
    new_B5507_, new_B5508_, new_B5509_, new_B5510_, new_B5511_, new_B5517_,
    new_B5518_, new_B5519_, new_B5520_, new_B5521_, new_B5522_, new_B5523_,
    new_B5524_, new_B5525_, new_B5526_, new_B5527_, new_B5528_, new_B5529_,
    new_B5530_, new_B5531_, new_B5532_, new_B5533_, new_B5534_, new_B5535_,
    new_B5536_, new_B5537_, new_B5538_, new_B5539_, new_B5540_, new_B5541_,
    new_B5542_, new_B5543_, new_B5544_, new_B5550_, new_B5551_, new_B5552_,
    new_B5553_, new_B5554_, new_B5555_, new_B5556_, new_B5557_, new_B5558_,
    new_B5559_, new_B5560_, new_B5561_, new_B5562_, new_B5563_, new_B5564_,
    new_B5565_, new_B5566_, new_B5567_, new_B5568_, new_B5569_, new_B5570_,
    new_B5571_, new_B5572_, new_B5573_, new_B5574_, new_B5575_, new_B5576_,
    new_B5577_, new_B5583_, new_B5584_, new_B5585_, new_B5586_, new_B5587_,
    new_B5588_, new_B5589_, new_B5590_, new_B5591_, new_B5592_, new_B5593_,
    new_B5594_, new_B5595_, new_B5596_, new_B5597_, new_B5598_, new_B5599_,
    new_B5600_, new_B5601_, new_B5602_, new_B5603_, new_B5604_, new_B5605_,
    new_B5606_, new_B5607_, new_B5608_, new_B5609_, new_B5610_, new_B5616_,
    new_B5617_, new_B5618_, new_B5619_, new_B5620_, new_B5621_, new_B5622_,
    new_B5623_, new_B5624_, new_B5625_, new_B5626_, new_B5627_, new_B5628_,
    new_B5629_, new_B5630_, new_B5631_, new_B5632_, new_B5633_, new_B5634_,
    new_B5635_, new_B5636_, new_B5637_, new_B5638_, new_B5639_, new_B5640_,
    new_B5641_, new_B5642_, new_B5643_, new_B5649_, new_B5650_, new_B5651_,
    new_B5652_, new_B5653_, new_B5654_, new_B5655_, new_B5656_, new_B5657_,
    new_B5658_, new_B5659_, new_B5660_, new_B5661_, new_B5662_, new_B5663_,
    new_B5664_, new_B5665_, new_B5666_, new_B5667_, new_B5668_, new_B5669_,
    new_B5670_, new_B5671_, new_B5672_, new_B5673_, new_B5674_, new_B5675_,
    new_B5676_, new_B5682_, new_B5683_, new_B5684_, new_B5685_, new_B5686_,
    new_B5687_, new_B5688_, new_B5689_, new_B5690_, new_B5691_, new_B5692_,
    new_B5693_, new_B5694_, new_B5695_, new_B5696_, new_B5697_, new_B5698_,
    new_B5699_, new_B5700_, new_B5701_, new_B5702_, new_B5703_, new_B5704_,
    new_B5705_, new_B5706_, new_B5707_, new_B5708_, new_B5709_, new_B5715_,
    new_B5716_, new_B5717_, new_B5718_, new_B5719_, new_B5720_, new_B5721_,
    new_B5722_, new_B5723_, new_B5724_, new_B5725_, new_B5726_, new_B5727_,
    new_B5728_, new_B5729_, new_B5730_, new_B5731_, new_B5732_, new_B5733_,
    new_B5734_, new_B5735_, new_B5736_, new_B5737_, new_B5738_, new_B5739_,
    new_B5740_, new_B5741_, new_B5742_, new_B5748_, new_B5749_, new_B5750_,
    new_B5751_, new_B5752_, new_B5753_, new_B5754_, new_B5755_, new_B5756_,
    new_B5757_, new_B5758_, new_B5759_, new_B5760_, new_B5761_, new_B5762_,
    new_B5763_, new_B5764_, new_B5765_, new_B5766_, new_B5767_, new_B5768_,
    new_B5769_, new_B5770_, new_B5771_, new_B5772_, new_B5773_, new_B5774_,
    new_B5775_, new_B5781_, new_B5782_, new_B5783_, new_B5784_, new_B5785_,
    new_B5786_, new_B5787_, new_B5788_, new_B5789_, new_B5790_, new_B5791_,
    new_B5792_, new_B5793_, new_B5794_, new_B5795_, new_B5796_, new_B5797_,
    new_B5798_, new_B5799_, new_B5800_, new_B5801_, new_B5802_, new_B5803_,
    new_B5804_, new_B5805_, new_B5806_, new_B5807_, new_B5808_, new_B5814_,
    new_B5815_, new_B5816_, new_B5817_, new_B5818_, new_B5819_, new_B5820_,
    new_B5821_, new_B5822_, new_B5823_, new_B5824_, new_B5825_, new_B5826_,
    new_B5827_, new_B5828_, new_B5829_, new_B5830_, new_B5831_, new_B5832_,
    new_B5833_, new_B5834_, new_B5835_, new_B5836_, new_B5837_, new_B5838_,
    new_B5839_, new_B5840_, new_B5841_, new_B5847_, new_B5848_, new_B5849_,
    new_B5850_, new_B5851_, new_B5852_, new_B5853_, new_B5854_, new_B5855_,
    new_B5856_, new_B5857_, new_B5858_, new_B5859_, new_B5860_, new_B5861_,
    new_B5862_, new_B5863_, new_B5864_, new_B5865_, new_B5866_, new_B5867_,
    new_B5868_, new_B5869_, new_B5870_, new_B5871_, new_B5872_, new_B5873_,
    new_B5874_, new_B5880_, new_B5881_, new_B5882_, new_B5883_, new_B5884_,
    new_B5885_, new_B5886_, new_B5887_, new_B5888_, new_B5889_, new_B5890_,
    new_B5891_, new_B5892_, new_B5893_, new_B5894_, new_B5895_, new_B5896_,
    new_B5897_, new_B5898_, new_B5899_, new_B5900_, new_B5901_, new_B5902_,
    new_B5903_, new_B5904_, new_B5905_, new_B5906_, new_B5907_, new_B5913_,
    new_B5914_, new_B5915_, new_B5916_, new_B5917_, new_B5918_, new_B5919_,
    new_B5920_, new_B5921_, new_B5922_, new_B5923_, new_B5924_, new_B5925_,
    new_B5926_, new_B5927_, new_B5928_, new_B5929_, new_B5930_, new_B5931_,
    new_B5932_, new_B5933_, new_B5934_, new_B5935_, new_B5936_, new_B5937_,
    new_B5938_, new_B5939_, new_B5940_, new_B5946_, new_B5947_, new_B5948_,
    new_B5949_, new_B5950_, new_B5951_, new_B5952_, new_B5953_, new_B5954_,
    new_B5955_, new_B5956_, new_B5957_, new_B5958_, new_B5959_, new_B5960_,
    new_B5961_, new_B5962_, new_B5963_, new_B5964_, new_B5965_, new_B5966_,
    new_B5967_, new_B5968_, new_B5969_, new_B5970_, new_B5971_, new_B5972_,
    new_B5973_, new_B5979_, new_B5980_, new_B5981_, new_B5982_, new_B5983_,
    new_B5984_, new_B5985_, new_B5986_, new_B5987_, new_B5988_, new_B5989_,
    new_B5990_, new_B5991_, new_B5992_, new_B5993_, new_B5994_, new_B5995_,
    new_B5996_, new_B5997_, new_B5998_, new_B5999_, new_B6000_, new_B6001_,
    new_B6002_, new_B6003_, new_B6004_, new_B6005_, new_B6006_, new_B6012_,
    new_B6013_, new_B6014_, new_B6015_, new_B6016_, new_B6017_, new_B6018_,
    new_B6019_, new_B6020_, new_B6021_, new_B6022_, new_B6023_, new_B6024_,
    new_B6025_, new_B6026_, new_B6027_, new_B6028_, new_B6029_, new_B6030_,
    new_B6031_, new_B6032_, new_B6033_, new_B6034_, new_B6035_, new_B6036_,
    new_B6037_, new_B6038_, new_B6039_, new_B6045_, new_B6046_, new_B6047_,
    new_B6048_, new_B6049_, new_B6050_, new_B6051_, new_B6052_, new_B6053_,
    new_B6054_, new_B6055_, new_B6056_, new_B6057_, new_B6058_, new_B6059_,
    new_B6060_, new_B6061_, new_B6062_, new_B6063_, new_B6064_, new_B6065_,
    new_B6066_, new_B6067_, new_B6068_, new_B6069_, new_B6070_, new_B6071_,
    new_B6072_, new_B6078_, new_B6079_, new_B6080_, new_B6081_, new_B6082_,
    new_B6083_, new_B6084_, new_B6085_, new_B6086_, new_B6087_, new_B6088_,
    new_B6089_, new_B6090_, new_B6091_, new_B6092_, new_B6093_, new_B6094_,
    new_B6095_, new_B6096_, new_B6097_, new_B6098_, new_B6099_, new_B6100_,
    new_B6101_, new_B6102_, new_B6103_, new_B6104_, new_B6105_, new_B6111_,
    new_B6112_, new_B6113_, new_B6114_, new_B6115_, new_B6116_, new_B6117_,
    new_B6118_, new_B6119_, new_B6120_, new_B6121_, new_B6122_, new_B6123_,
    new_B6124_, new_B6125_, new_B6126_, new_B6127_, new_B6128_, new_B6129_,
    new_B6130_, new_B6131_, new_B6132_, new_B6133_, new_B6134_, new_B6135_,
    new_B6136_, new_B6137_, new_B6138_, new_B6144_, new_B6145_, new_B6146_,
    new_B6147_, new_B6148_, new_B6149_, new_B6150_, new_B6151_, new_B6152_,
    new_B6153_, new_B6154_, new_B6155_, new_B6156_, new_B6157_, new_B6158_,
    new_B6159_, new_B6160_, new_B6161_, new_B6162_, new_B6163_, new_B6164_,
    new_B6165_, new_B6166_, new_B6167_, new_B6168_, new_B6169_, new_B6170_,
    new_B6171_, new_B6177_, new_B6178_, new_B6179_, new_B6180_, new_B6181_,
    new_B6182_, new_B6183_, new_B6184_, new_B6185_, new_B6186_, new_B6187_,
    new_B6188_, new_B6189_, new_B6190_, new_B6191_, new_B6192_, new_B6193_,
    new_B6194_, new_B6195_, new_B6196_, new_B6197_, new_B6198_, new_B6199_,
    new_B6200_, new_B6201_, new_B6202_, new_B6203_, new_B6204_, new_B6210_,
    new_B6211_, new_B6212_, new_B6213_, new_B6214_, new_B6215_, new_B6216_,
    new_B6217_, new_B6218_, new_B6219_, new_B6220_, new_B6221_, new_B6222_,
    new_B6223_, new_B6224_, new_B6225_, new_B6226_, new_B6227_, new_B6228_,
    new_B6229_, new_B6230_, new_B6231_, new_B6232_, new_B6233_, new_B6234_,
    new_B6235_, new_B6236_, new_B6237_, new_B6243_, new_B6244_, new_B6245_,
    new_B6246_, new_B6247_, new_B6248_, new_B6249_, new_B6250_, new_B6251_,
    new_B6252_, new_B6253_, new_B6254_, new_B6255_, new_B6256_, new_B6257_,
    new_B6258_, new_B6259_, new_B6260_, new_B6261_, new_B6262_, new_B6263_,
    new_B6264_, new_B6265_, new_B6266_, new_B6267_, new_B6268_, new_B6269_,
    new_B6270_, new_B6276_, new_B6277_, new_B6278_, new_B6279_, new_B6280_,
    new_B6281_, new_B6282_, new_B6283_, new_B6284_, new_B6285_, new_B6286_,
    new_B6287_, new_B6288_, new_B6289_, new_B6290_, new_B6291_, new_B6292_,
    new_B6293_, new_B6294_, new_B6295_, new_B6296_, new_B6297_, new_B6298_,
    new_B6299_, new_B6300_, new_B6301_, new_B6302_, new_B6303_, new_B6309_,
    new_B6310_, new_B6311_, new_B6312_, new_B6313_, new_B6314_, new_B6315_,
    new_B6316_, new_B6317_, new_B6318_, new_B6319_, new_B6320_, new_B6321_,
    new_B6322_, new_B6323_, new_B6324_, new_B6325_, new_B6326_, new_B6327_,
    new_B6328_, new_B6329_, new_B6330_, new_B6331_, new_B6332_, new_B6333_,
    new_B6334_, new_B6335_, new_B6336_, new_B6342_, new_B6343_, new_B6344_,
    new_B6345_, new_B6346_, new_B6347_, new_B6348_, new_B6349_, new_B6350_,
    new_B6351_, new_B6352_, new_B6353_, new_B6354_, new_B6355_, new_B6356_,
    new_B6357_, new_B6358_, new_B6359_, new_B6360_, new_B6361_, new_B6362_,
    new_B6363_, new_B6364_, new_B6365_, new_B6366_, new_B6367_, new_B6368_,
    new_B6369_, new_B6375_, new_B6376_, new_B6377_, new_B6378_, new_B6379_,
    new_B6380_, new_B6381_, new_B6382_, new_B6383_, new_B6384_, new_B6385_,
    new_B6386_, new_B6387_, new_B6388_, new_B6389_, new_B6390_, new_B6391_,
    new_B6392_, new_B6393_, new_B6394_, new_B6395_, new_B6396_, new_B6397_,
    new_B6398_, new_B6399_, new_B6400_, new_B6401_, new_B6402_, new_B6408_,
    new_B6409_, new_B6410_, new_B6411_, new_B6412_, new_B6413_, new_B6414_,
    new_B6415_, new_B6416_, new_B6417_, new_B6418_, new_B6419_, new_B6420_,
    new_B6421_, new_B6422_, new_B6423_, new_B6424_, new_B6425_, new_B6426_,
    new_B6427_, new_B6428_, new_B6429_, new_B6430_, new_B6431_, new_B6432_,
    new_B6433_, new_B6434_, new_B6435_, new_B6441_, new_B6442_, new_B6443_,
    new_B6444_, new_B6445_, new_B6446_, new_B6447_, new_B6448_, new_B6449_,
    new_B6450_, new_B6451_, new_B6452_, new_B6453_, new_B6454_, new_B6455_,
    new_B6456_, new_B6457_, new_B6458_, new_B6459_, new_B6460_, new_B6461_,
    new_B6462_, new_B6463_, new_B6464_, new_B6465_, new_B6466_, new_B6467_,
    new_B6468_, new_B6474_, new_B6475_, new_B6476_, new_B6477_, new_B6478_,
    new_B6479_, new_B6480_, new_B6481_, new_B6482_, new_B6483_, new_B6484_,
    new_B6485_, new_B6486_, new_B6487_, new_B6488_, new_B6489_, new_B6490_,
    new_B6491_, new_B6492_, new_B6493_, new_B6494_, new_B6495_, new_B6496_,
    new_B6497_, new_B6498_, new_B6499_, new_B6500_, new_B6501_, new_B6507_,
    new_B6508_, new_B6509_, new_B6510_, new_B6511_, new_B6512_, new_B6513_,
    new_B6514_, new_B6515_, new_B6516_, new_B6517_, new_B6518_, new_B6519_,
    new_B6520_, new_B6521_, new_B6522_, new_B6523_, new_B6524_, new_B6525_,
    new_B6526_, new_B6527_, new_B6528_, new_B6529_, new_B6530_, new_B6531_,
    new_B6532_, new_B6533_, new_B6534_, new_B6540_, new_B6541_, new_B6542_,
    new_B6543_, new_B6544_, new_B6545_, new_B6546_, new_B6547_, new_B6548_,
    new_B6549_, new_B6550_, new_B6551_, new_B6552_, new_B6553_, new_B6554_,
    new_B6555_, new_B6556_, new_B6557_, new_B6558_, new_B6559_, new_B6560_,
    new_B6561_, new_B6562_, new_B6563_, new_B6564_, new_B6565_, new_B6566_,
    new_B6567_, new_B6573_, new_B6574_, new_B6575_, new_B6576_, new_B6577_,
    new_B6578_, new_B6579_, new_B6580_, new_B6581_, new_B6582_, new_B6583_,
    new_B6584_, new_B6585_, new_B6586_, new_B6587_, new_B6588_, new_B6589_,
    new_B6590_, new_B6591_, new_B6592_, new_B6593_, new_B6594_, new_B6595_,
    new_B6596_, new_B6597_, new_B6598_, new_B6599_, new_B6600_, new_B6606_,
    new_B6607_, new_B6608_, new_B6609_, new_B6610_, new_B6611_, new_B6612_,
    new_B6613_, new_B6614_, new_B6615_, new_B6616_, new_B6617_, new_B6618_,
    new_B6619_, new_B6620_, new_B6621_, new_B6622_, new_B6623_, new_B6624_,
    new_B6625_, new_B6626_, new_B6627_, new_B6628_, new_B6629_, new_B6630_,
    new_B6631_, new_B6632_, new_B6633_, new_B6639_, new_B6640_, new_B6641_,
    new_B6642_, new_B6643_, new_B6644_, new_B6645_, new_B6646_, new_B6647_,
    new_B6648_, new_B6649_, new_B6650_, new_B6651_, new_B6652_, new_B6653_,
    new_B6654_, new_B6655_, new_B6656_, new_B6657_, new_B6658_, new_B6659_,
    new_B6660_, new_B6661_, new_B6662_, new_B6663_, new_B6664_, new_B6665_,
    new_B6666_, new_B6672_, new_B6673_, new_B6674_, new_B6675_, new_B6676_,
    new_B6677_, new_B6678_, new_B6679_, new_B6680_, new_B6681_, new_B6682_,
    new_B6683_, new_B6684_, new_B6685_, new_B6686_, new_B6687_, new_B6688_,
    new_B6689_, new_B6690_, new_B6691_, new_B6692_, new_B6693_, new_B6694_,
    new_B6695_, new_B6696_, new_B6697_, new_B6698_, new_B6699_, new_B6705_,
    new_B6706_, new_B6707_, new_B6708_, new_B6709_, new_B6710_, new_B6711_,
    new_B6712_, new_B6713_, new_B6714_, new_B6715_, new_B6716_, new_B6717_,
    new_B6718_, new_B6719_, new_B6720_, new_B6721_, new_B6722_, new_B6723_,
    new_B6724_, new_B6725_, new_B6726_, new_B6727_, new_B6728_, new_B6729_,
    new_B6730_, new_B6731_, new_B6732_, new_B6738_, new_B6739_, new_B6740_,
    new_B6741_, new_B6742_, new_B6743_, new_B6744_, new_B6745_, new_B6746_,
    new_B6747_, new_B6748_, new_B6749_, new_B6750_, new_B6751_, new_B6752_,
    new_B6753_, new_B6754_, new_B6755_, new_B6756_, new_B6757_, new_B6758_,
    new_B6759_, new_B6760_, new_B6761_, new_B6762_, new_B6763_, new_B6764_,
    new_B6765_, new_B6771_, new_B6772_, new_B6773_, new_B6774_, new_B6775_,
    new_B6776_, new_B6777_, new_B6778_, new_B6779_, new_B6780_, new_B6781_,
    new_B6782_, new_B6783_, new_B6784_, new_B6785_, new_B6786_, new_B6787_,
    new_B6788_, new_B6789_, new_B6790_, new_B6791_, new_B6792_, new_B6793_,
    new_B6794_, new_B6795_, new_B6796_, new_B6797_, new_B6798_, new_B6804_,
    new_B6805_, new_B6806_, new_B6807_, new_B6808_, new_B6809_, new_B6810_,
    new_B6811_, new_B6812_, new_B6813_, new_B6814_, new_B6815_, new_B6816_,
    new_B6817_, new_B6818_, new_B6819_, new_B6820_, new_B6821_, new_B6822_,
    new_B6823_, new_B6824_, new_B6825_, new_B6826_, new_B6827_, new_B6828_,
    new_B6829_, new_B6830_, new_B6831_, new_B6837_, new_B6838_, new_B6839_,
    new_B6840_, new_B6841_, new_B6842_, new_B6843_, new_B6844_, new_B6845_,
    new_B6846_, new_B6847_, new_B6848_, new_B6849_, new_B6850_, new_B6851_,
    new_B6852_, new_B6853_, new_B6854_, new_B6855_, new_B6856_, new_B6857_,
    new_B6858_, new_B6859_, new_B6860_, new_B6861_, new_B6862_, new_B6863_,
    new_B6864_, new_B6870_, new_B6871_, new_B6872_, new_B6873_, new_B6874_,
    new_B6875_, new_B6876_, new_B6877_, new_B6878_, new_B6879_, new_B6880_,
    new_B6881_, new_B6882_, new_B6883_, new_B6884_, new_B6885_, new_B6886_,
    new_B6887_, new_B6888_, new_B6889_, new_B6890_, new_B6891_, new_B6892_,
    new_B6893_, new_B6894_, new_B6895_, new_B6896_, new_B6897_, new_B6903_,
    new_B6904_, new_B6905_, new_B6906_, new_B6907_, new_B6908_, new_B6909_,
    new_B6910_, new_B6911_, new_B6912_, new_B6913_, new_B6914_, new_B6915_,
    new_B6916_, new_B6917_, new_B6918_, new_B6919_, new_B6920_, new_B6921_,
    new_B6922_, new_B6923_, new_B6924_, new_B6925_, new_B6926_, new_B6927_,
    new_B6928_, new_B6929_, new_B6930_, new_B6936_, new_B6937_, new_B6938_,
    new_B6939_, new_B6940_, new_B6941_, new_B6942_, new_B6943_, new_B6944_,
    new_B6945_, new_B6946_, new_B6947_, new_B6948_, new_B6949_, new_B6950_,
    new_B6951_, new_B6952_, new_B6953_, new_B6954_, new_B6955_, new_B6956_,
    new_B6957_, new_B6958_, new_B6959_, new_B6960_, new_B6961_, new_B6962_,
    new_B6963_, new_B6969_, new_B6970_, new_B6971_, new_B6972_, new_B6973_,
    new_B6974_, new_B6975_, new_B6976_, new_B6977_, new_B6978_, new_B6979_,
    new_B6980_, new_B6981_, new_B6982_, new_B6983_, new_B6984_, new_B6985_,
    new_B6986_, new_B6987_, new_B6988_, new_B6989_, new_B6990_, new_B6991_,
    new_B6992_, new_B6993_, new_B6994_, new_B6995_, new_B6996_, new_B7002_,
    new_B7003_, new_B7004_, new_B7005_, new_B7006_, new_B7007_, new_B7008_,
    new_B7009_, new_B7010_, new_B7011_, new_B7012_, new_B7013_, new_B7014_,
    new_B7015_, new_B7016_, new_B7017_, new_B7018_, new_B7019_, new_B7020_,
    new_B7021_, new_B7022_, new_B7023_, new_B7024_, new_B7025_, new_B7026_,
    new_B7027_, new_B7028_, new_B7029_, new_B7035_, new_B7036_, new_B7037_,
    new_B7038_, new_B7039_, new_B7040_, new_B7041_, new_B7042_, new_B7043_,
    new_B7044_, new_B7045_, new_B7046_, new_B7047_, new_B7048_, new_B7049_,
    new_B7050_, new_B7051_, new_B7052_, new_B7053_, new_B7054_, new_B7055_,
    new_B7056_, new_B7057_, new_B7058_, new_B7059_, new_B7060_, new_B7061_,
    new_B7062_, new_B7068_, new_B7069_, new_B7070_, new_B7071_, new_B7072_,
    new_B7073_, new_B7074_, new_B7075_, new_B7076_, new_B7077_, new_B7078_,
    new_B7079_, new_B7080_, new_B7081_, new_B7082_, new_B7083_, new_B7084_,
    new_B7085_, new_B7086_, new_B7087_, new_B7088_, new_B7089_, new_B7090_,
    new_B7091_, new_B7092_, new_B7093_, new_B7094_, new_B7095_, new_B7101_,
    new_B7102_, new_B7103_, new_B7104_, new_B7105_, new_B7106_, new_B7107_,
    new_B7108_, new_B7109_, new_B7110_, new_B7111_, new_B7112_, new_B7113_,
    new_B7114_, new_B7115_, new_B7116_, new_B7117_, new_B7118_, new_B7119_,
    new_B7120_, new_B7121_, new_B7122_, new_B7123_, new_B7124_, new_B7125_,
    new_B7126_, new_B7127_, new_B7128_, new_B7134_, new_B7135_, new_B7136_,
    new_B7137_, new_B7138_, new_B7139_, new_B7140_, new_B7141_, new_B7142_,
    new_B7143_, new_B7144_, new_B7145_, new_B7146_, new_B7147_, new_B7148_,
    new_B7149_, new_B7150_, new_B7151_, new_B7152_, new_B7153_, new_B7154_,
    new_B7155_, new_B7156_, new_B7157_, new_B7158_, new_B7159_, new_B7160_,
    new_B7161_, new_B7167_, new_B7168_, new_B7169_, new_B7170_, new_B7171_,
    new_B7172_, new_B7173_, new_B7174_, new_B7175_, new_B7176_, new_B7177_,
    new_B7178_, new_B7179_, new_B7180_, new_B7181_, new_B7182_, new_B7183_,
    new_B7184_, new_B7185_, new_B7186_, new_B7187_, new_B7188_, new_B7189_,
    new_B7190_, new_B7191_, new_B7192_, new_B7193_, new_B7194_, new_B7200_,
    new_B7201_, new_B7202_, new_B7203_, new_B7204_, new_B7205_, new_B7206_,
    new_B7207_, new_B7208_, new_B7209_, new_B7210_, new_B7211_, new_B7212_,
    new_B7213_, new_B7214_, new_B7215_, new_B7216_, new_B7217_, new_B7218_,
    new_B7219_, new_B7220_, new_B7221_, new_B7222_, new_B7223_, new_B7224_,
    new_B7225_, new_B7226_, new_B7227_, new_B7233_, new_B7234_, new_B7235_,
    new_B7236_, new_B7237_, new_B7238_, new_B7239_, new_B7240_, new_B7241_,
    new_B7242_, new_B7243_, new_B7244_, new_B7245_, new_B7246_, new_B7247_,
    new_B7248_, new_B7249_, new_B7250_, new_B7251_, new_B7252_, new_B7253_,
    new_B7254_, new_B7255_, new_B7256_, new_B7257_, new_B7258_, new_B7259_,
    new_B7260_, new_B7266_, new_B7267_, new_B7268_, new_B7269_, new_B7270_,
    new_B7271_, new_B7272_, new_B7273_, new_B7274_, new_B7275_, new_B7276_,
    new_B7277_, new_B7278_, new_B7279_, new_B7280_, new_B7281_, new_B7282_,
    new_B7283_, new_B7284_, new_B7285_, new_B7286_, new_B7287_, new_B7288_,
    new_B7289_, new_B7290_, new_B7291_, new_B7292_, new_B7293_, new_B7299_,
    new_B7300_, new_B7301_, new_B7302_, new_B7303_, new_B7304_, new_B7305_,
    new_B7306_, new_B7307_, new_B7308_, new_B7309_, new_B7310_, new_B7311_,
    new_B7312_, new_B7313_, new_B7314_, new_B7315_, new_B7316_, new_B7317_,
    new_B7318_, new_B7319_, new_B7320_, new_B7321_, new_B7322_, new_B7323_,
    new_B7324_, new_B7325_, new_B7326_, new_B7332_, new_B7333_, new_B7334_,
    new_B7335_, new_B7336_, new_B7337_, new_B7338_, new_B7339_, new_B7340_,
    new_B7341_, new_B7342_, new_B7343_, new_B7344_, new_B7345_, new_B7346_,
    new_B7347_, new_B7348_, new_B7349_, new_B7350_, new_B7351_, new_B7352_,
    new_B7353_, new_B7354_, new_B7355_, new_B7356_, new_B7357_, new_B7358_,
    new_B7359_, new_B7365_, new_B7366_, new_B7367_, new_B7368_, new_B7369_,
    new_B7370_, new_B7371_, new_B7372_, new_B7373_, new_B7374_, new_B7375_,
    new_B7376_, new_B7377_, new_B7378_, new_B7379_, new_B7380_, new_B7381_,
    new_B7382_, new_B7383_, new_B7384_, new_B7385_, new_B7386_, new_B7387_,
    new_B7388_, new_B7389_, new_B7390_, new_B7391_, new_B7392_, new_B7398_,
    new_B7399_, new_B7400_, new_B7401_, new_B7402_, new_B7403_, new_B7404_,
    new_B7405_, new_B7406_, new_B7407_, new_B7408_, new_B7409_, new_B7410_,
    new_B7411_, new_B7412_, new_B7413_, new_B7414_, new_B7415_, new_B7416_,
    new_B7417_, new_B7418_, new_B7419_, new_B7420_, new_B7421_, new_B7422_,
    new_B7423_, new_B7424_, new_B7425_, new_B7431_, new_B7432_, new_B7433_,
    new_B7434_, new_B7435_, new_B7436_, new_B7437_, new_B7438_, new_B7439_,
    new_B7440_, new_B7441_, new_B7442_, new_B7443_, new_B7444_, new_B7445_,
    new_B7446_, new_B7447_, new_B7448_, new_B7449_, new_B7450_, new_B7451_,
    new_B7452_, new_B7453_, new_B7454_, new_B7455_, new_B7456_, new_B7457_,
    new_B7458_, new_B7464_, new_B7465_, new_B7466_, new_B7467_, new_B7468_,
    new_B7469_, new_B7470_, new_B7471_, new_B7472_, new_B7473_, new_B7474_,
    new_B7475_, new_B7476_, new_B7477_, new_B7478_, new_B7479_, new_B7480_,
    new_B7481_, new_B7482_, new_B7483_, new_B7484_, new_B7485_, new_B7486_,
    new_B7487_, new_B7488_, new_B7489_, new_B7490_, new_B7491_, new_B7497_,
    new_B7498_, new_B7499_, new_B7500_, new_B7501_, new_B7502_, new_B7503_,
    new_B7504_, new_B7505_, new_B7506_, new_B7507_, new_B7508_, new_B7509_,
    new_B7510_, new_B7511_, new_B7512_, new_B7513_, new_B7514_, new_B7515_,
    new_B7516_, new_B7517_, new_B7518_, new_B7519_, new_B7520_, new_B7521_,
    new_B7522_, new_B7523_, new_B7524_, new_B7530_, new_B7531_, new_B7532_,
    new_B7533_, new_B7534_, new_B7535_, new_B7536_, new_B7537_, new_B7538_,
    new_B7539_, new_B7540_, new_B7541_, new_B7542_, new_B7543_, new_B7544_,
    new_B7545_, new_B7546_, new_B7547_, new_B7548_, new_B7549_, new_B7550_,
    new_B7551_, new_B7552_, new_B7553_, new_B7554_, new_B7555_, new_B7556_,
    new_B7557_, new_B7563_, new_B7564_, new_B7565_, new_B7566_, new_B7567_,
    new_B7568_, new_B7569_, new_B7570_, new_B7571_, new_B7572_, new_B7573_,
    new_B7574_, new_B7575_, new_B7576_, new_B7577_, new_B7578_, new_B7579_,
    new_B7580_, new_B7581_, new_B7582_, new_B7583_, new_B7584_, new_B7585_,
    new_B7586_, new_B7587_, new_B7588_, new_B7589_, new_B7590_, new_B7596_,
    new_B7597_, new_B7598_, new_B7599_, new_B7600_, new_B7601_, new_B7602_,
    new_B7603_, new_B7604_, new_B7605_, new_B7606_, new_B7607_, new_B7608_,
    new_B7609_, new_B7610_, new_B7611_, new_B7612_, new_B7613_, new_B7614_,
    new_B7615_, new_B7616_, new_B7617_, new_B7618_, new_B7619_, new_B7620_,
    new_B7621_, new_B7622_, new_B7623_, new_B7629_, new_B7630_, new_B7631_,
    new_B7632_, new_B7633_, new_B7634_, new_B7635_, new_B7636_, new_B7637_,
    new_B7638_, new_B7639_, new_B7640_, new_B7641_, new_B7642_, new_B7643_,
    new_B7644_, new_B7645_, new_B7646_, new_B7647_, new_B7648_, new_B7649_,
    new_B7650_, new_B7651_, new_B7652_, new_B7653_, new_B7654_, new_B7655_,
    new_B7656_, new_B7662_, new_B7663_, new_B7664_, new_B7665_, new_B7666_,
    new_B7667_, new_B7668_, new_B7669_, new_B7670_, new_B7671_, new_B7672_,
    new_B7673_, new_B7674_, new_B7675_, new_B7676_, new_B7677_, new_B7678_,
    new_B7679_, new_B7680_, new_B7681_, new_B7682_, new_B7683_, new_B7684_,
    new_B7685_, new_B7686_, new_B7687_, new_B7688_, new_B7689_, new_B7695_,
    new_B7696_, new_B7697_, new_B7698_, new_B7699_, new_B7700_, new_B7701_,
    new_B7702_, new_B7703_, new_B7704_, new_B7705_, new_B7706_, new_B7707_,
    new_B7708_, new_B7709_, new_B7710_, new_B7711_, new_B7712_, new_B7713_,
    new_B7714_, new_B7715_, new_B7716_, new_B7717_, new_B7718_, new_B7719_,
    new_B7720_, new_B7721_, new_B7722_, new_B7728_, new_B7729_, new_B7730_,
    new_B7731_, new_B7732_, new_B7733_, new_B7734_, new_B7735_, new_B7736_,
    new_B7737_, new_B7738_, new_B7739_, new_B7740_, new_B7741_, new_B7742_,
    new_B7743_, new_B7744_, new_B7745_, new_B7746_, new_B7747_, new_B7748_,
    new_B7749_, new_B7750_, new_B7751_, new_B7752_, new_B7753_, new_B7754_,
    new_B7755_, new_B7761_, new_B7762_, new_B7763_, new_B7764_, new_B7765_,
    new_B7766_, new_B7767_, new_B7768_, new_B7769_, new_B7770_, new_B7771_,
    new_B7772_, new_B7773_, new_B7774_, new_B7775_, new_B7776_, new_B7777_,
    new_B7778_, new_B7779_, new_B7780_, new_B7781_, new_B7782_, new_B7783_,
    new_B7784_, new_B7785_, new_B7786_, new_B7787_, new_B7788_, new_B7794_,
    new_B7795_, new_B7796_, new_B7797_, new_B7798_, new_B7799_, new_B7800_,
    new_B7801_, new_B7802_, new_B7803_, new_B7804_, new_B7805_, new_B7806_,
    new_B7807_, new_B7808_, new_B7809_, new_B7810_, new_B7811_, new_B7812_,
    new_B7813_, new_B7814_, new_B7815_, new_B7816_, new_B7817_, new_B7818_,
    new_B7819_, new_B7820_, new_B7821_, new_B7827_, new_B7828_, new_B7829_,
    new_B7830_, new_B7831_, new_B7832_, new_B7833_, new_B7834_, new_B7835_,
    new_B7836_, new_B7837_, new_B7838_, new_B7839_, new_B7840_, new_B7841_,
    new_B7842_, new_B7843_, new_B7844_, new_B7845_, new_B7846_, new_B7847_,
    new_B7848_, new_B7849_, new_B7850_, new_B7851_, new_B7852_, new_B7853_,
    new_B7854_, new_B7860_, new_B7861_, new_B7862_, new_B7863_, new_B7864_,
    new_B7865_, new_B7866_, new_B7867_, new_B7868_, new_B7869_, new_B7870_,
    new_B7871_, new_B7872_, new_B7873_, new_B7874_, new_B7875_, new_B7876_,
    new_B7877_, new_B7878_, new_B7879_, new_B7880_, new_B7881_, new_B7882_,
    new_B7883_, new_B7884_, new_B7885_, new_B7886_, new_B7887_, new_B7893_,
    new_B7894_, new_B7895_, new_B7896_, new_B7897_, new_B7898_, new_B7899_,
    new_B7900_, new_B7901_, new_B7902_, new_B7903_, new_B7904_, new_B7905_,
    new_B7906_, new_B7907_, new_B7908_, new_B7909_, new_B7910_, new_B7911_,
    new_B7912_, new_B7913_, new_B7914_, new_B7915_, new_B7916_, new_B7917_,
    new_B7918_, new_B7919_, new_B7920_, new_B7926_, new_B7927_, new_B7928_,
    new_B7929_, new_B7930_, new_B7931_, new_B7932_, new_B7933_, new_B7934_,
    new_B7935_, new_B7936_, new_B7937_, new_B7938_, new_B7939_, new_B7940_,
    new_B7941_, new_B7942_, new_B7943_, new_B7944_, new_B7945_, new_B7946_,
    new_B7947_, new_B7948_, new_B7949_, new_B7950_, new_B7951_, new_B7952_,
    new_B7953_, new_B7959_, new_B7960_, new_B7961_, new_B7962_, new_B7963_,
    new_B7964_, new_B7965_, new_B7966_, new_B7967_, new_B7968_, new_B7969_,
    new_B7970_, new_B7971_, new_B7972_, new_B7973_, new_B7974_, new_B7975_,
    new_B7976_, new_B7977_, new_B7978_, new_B7979_, new_B7980_, new_B7981_,
    new_B7982_, new_B7983_, new_B7984_, new_B7985_, new_B7986_, new_B7992_,
    new_B7993_, new_B7994_, new_B7995_, new_B7996_, new_B7997_, new_B7998_,
    new_B7999_, new_B8000_, new_B8001_, new_B8002_, new_B8003_, new_B8004_,
    new_B8005_, new_B8006_, new_B8007_, new_B8008_, new_B8009_, new_B8010_,
    new_B8011_, new_B8012_, new_B8013_, new_B8014_, new_B8015_, new_B8016_,
    new_B8017_, new_B8018_, new_B8019_, new_B8025_, new_B8026_, new_B8027_,
    new_B8028_, new_B8029_, new_B8030_, new_B8031_, new_B8032_, new_B8033_,
    new_B8034_, new_B8035_, new_B8036_, new_B8037_, new_B8038_, new_B8039_,
    new_B8040_, new_B8041_, new_B8042_, new_B8043_, new_B8044_, new_B8045_,
    new_B8046_, new_B8047_, new_B8048_, new_B8049_, new_B8050_, new_B8051_,
    new_B8052_, new_B8058_, new_B8059_, new_B8060_, new_B8061_, new_B8062_,
    new_B8063_, new_B8064_, new_B8065_, new_B8066_, new_B8067_, new_B8068_,
    new_B8069_, new_B8070_, new_B8071_, new_B8072_, new_B8073_, new_B8074_,
    new_B8075_, new_B8076_, new_B8077_, new_B8078_, new_B8079_, new_B8080_,
    new_B8081_, new_B8082_, new_B8083_, new_B8084_, new_B8085_, new_B8091_,
    new_B8092_, new_B8093_, new_B8094_, new_B8095_, new_B8096_, new_B8097_,
    new_B8098_, new_B8099_, new_B8100_, new_B8101_, new_B8102_, new_B8103_,
    new_B8104_, new_B8105_, new_B8106_, new_B8107_, new_B8108_, new_B8109_,
    new_B8110_, new_B8111_, new_B8112_, new_B8113_, new_B8114_, new_B8115_,
    new_B8116_, new_B8117_, new_B8118_, new_B8124_, new_B8125_, new_B8126_,
    new_B8127_, new_B8128_, new_B8129_, new_B8130_, new_B8131_, new_B8132_,
    new_B8133_, new_B8134_, new_B8135_, new_B8136_, new_B8137_, new_B8138_,
    new_B8139_, new_B8140_, new_B8141_, new_B8142_, new_B8143_, new_B8144_,
    new_B8145_, new_B8146_, new_B8147_, new_B8148_, new_B8149_, new_B8150_,
    new_B8151_, new_B8157_, new_B8158_, new_B8159_, new_B8160_, new_B8161_,
    new_B8162_, new_B8163_, new_B8164_, new_B8165_, new_B8166_, new_B8167_,
    new_B8168_, new_B8169_, new_B8170_, new_B8171_, new_B8172_, new_B8173_,
    new_B8174_, new_B8175_, new_B8176_, new_B8177_, new_B8178_, new_B8179_,
    new_B8180_, new_B8181_, new_B8182_, new_B8183_, new_B8184_, new_B8190_,
    new_B8191_, new_B8192_, new_B8193_, new_B8194_, new_B8195_, new_B8196_,
    new_B8197_, new_B8198_, new_B8199_, new_B8200_, new_B8201_, new_B8202_,
    new_B8203_, new_B8204_, new_B8205_, new_B8206_, new_B8207_, new_B8208_,
    new_B8209_, new_B8210_, new_B8211_, new_B8212_, new_B8213_, new_B8214_,
    new_B8215_, new_B8216_, new_B8217_, new_B8223_, new_B8224_, new_B8225_,
    new_B8226_, new_B8227_, new_B8228_, new_B8229_, new_B8230_, new_B8231_,
    new_B8232_, new_B8233_, new_B8234_, new_B8235_, new_B8236_, new_B8237_,
    new_B8238_, new_B8239_, new_B8240_, new_B8241_, new_B8242_, new_B8243_,
    new_B8244_, new_B8245_, new_B8246_, new_B8247_, new_B8248_, new_B8249_,
    new_B8250_, new_B8256_, new_B8257_, new_B8258_, new_B8259_, new_B8260_,
    new_B8261_, new_B8262_, new_B8263_, new_B8264_, new_B8265_, new_B8266_,
    new_B8267_, new_B8268_, new_B8269_, new_B8270_, new_B8271_, new_B8272_,
    new_B8273_, new_B8274_, new_B8275_, new_B8276_, new_B8277_, new_B8278_,
    new_B8279_, new_B8280_, new_B8281_, new_B8282_, new_B8283_, new_B8289_,
    new_B8290_, new_B8291_, new_B8292_, new_B8293_, new_B8294_, new_B8295_,
    new_B8296_, new_B8297_, new_B8298_, new_B8299_, new_B8300_, new_B8301_,
    new_B8302_, new_B8303_, new_B8304_, new_B8305_, new_B8306_, new_B8307_,
    new_B8308_, new_B8309_, new_B8310_, new_B8311_, new_B8312_, new_B8313_,
    new_B8314_, new_B8315_, new_B8316_, new_B8322_, new_B8323_, new_B8324_,
    new_B8325_, new_B8326_, new_B8327_, new_B8328_, new_B8329_, new_B8330_,
    new_B8331_, new_B8332_, new_B8333_, new_B8334_, new_B8335_, new_B8336_,
    new_B8337_, new_B8338_, new_B8339_, new_B8340_, new_B8341_, new_B8342_,
    new_B8343_, new_B8344_, new_B8345_, new_B8346_, new_B8347_, new_B8348_,
    new_B8349_, new_B8355_, new_B8356_, new_B8357_, new_B8358_, new_B8359_,
    new_B8360_, new_B8361_, new_B8362_, new_B8363_, new_B8364_, new_B8365_,
    new_B8366_, new_B8367_, new_B8368_, new_B8369_, new_B8370_, new_B8371_,
    new_B8372_, new_B8373_, new_B8374_, new_B8375_, new_B8376_, new_B8377_,
    new_B8378_, new_B8379_, new_B8380_, new_B8381_, new_B8382_, new_B8388_,
    new_B8389_, new_B8390_, new_B8391_, new_B8392_, new_B8393_, new_B8394_,
    new_B8395_, new_B8396_, new_B8397_, new_B8398_, new_B8399_, new_B8400_,
    new_B8401_, new_B8402_, new_B8403_, new_B8404_, new_B8405_, new_B8406_,
    new_B8407_, new_B8408_, new_B8409_, new_B8410_, new_B8411_, new_B8412_,
    new_B8413_, new_B8414_, new_B8415_, new_B8421_, new_B8422_, new_B8423_,
    new_B8424_, new_B8425_, new_B8426_, new_B8427_, new_B8428_, new_B8429_,
    new_B8430_, new_B8431_, new_B8432_, new_B8433_, new_B8434_, new_B8435_,
    new_B8436_, new_B8437_, new_B8438_, new_B8439_, new_B8440_, new_B8441_,
    new_B8442_, new_B8443_, new_B8444_, new_B8445_, new_B8446_, new_B8447_,
    new_B8448_, new_B8454_, new_B8455_, new_B8456_, new_B8457_, new_B8458_,
    new_B8459_, new_B8460_, new_B8461_, new_B8462_, new_B8463_, new_B8464_,
    new_B8465_, new_B8466_, new_B8467_, new_B8468_, new_B8469_, new_B8470_,
    new_B8471_, new_B8472_, new_B8473_, new_B8474_, new_B8475_, new_B8476_,
    new_B8477_, new_B8478_, new_B8479_, new_B8480_, new_B8481_, new_B8487_,
    new_B8488_, new_B8489_, new_B8490_, new_B8491_, new_B8492_, new_B8493_,
    new_B8494_, new_B8495_, new_B8496_, new_B8497_, new_B8498_, new_B8499_,
    new_B8500_, new_B8501_, new_B8502_, new_B8503_, new_B8504_, new_B8505_,
    new_B8506_, new_B8507_, new_B8508_, new_B8509_, new_B8510_, new_B8511_,
    new_B8512_, new_B8513_, new_B8514_, new_B8520_, new_B8521_, new_B8522_,
    new_B8523_, new_B8524_, new_B8525_, new_B8526_, new_B8527_, new_B8528_,
    new_B8529_, new_B8530_, new_B8531_, new_B8532_, new_B8533_, new_B8534_,
    new_B8535_, new_B8536_, new_B8537_, new_B8538_, new_B8539_, new_B8540_,
    new_B8541_, new_B8542_, new_B8543_, new_B8544_, new_B8545_, new_B8546_,
    new_B8547_, new_B8553_, new_B8554_, new_B8555_, new_B8556_, new_B8557_,
    new_B8558_, new_B8559_, new_B8560_, new_B8561_, new_B8562_, new_B8563_,
    new_B8564_, new_B8565_, new_B8566_, new_B8567_, new_B8568_, new_B8569_,
    new_B8570_, new_B8571_, new_B8572_, new_B8573_, new_B8574_, new_B8575_,
    new_B8576_, new_B8577_, new_B8578_, new_B8579_, new_B8580_, new_B8586_,
    new_B8587_, new_B8588_, new_B8589_, new_B8590_, new_B8591_, new_B8592_,
    new_B8593_, new_B8594_, new_B8595_, new_B8596_, new_B8597_, new_B8598_,
    new_B8599_, new_B8600_, new_B8601_, new_B8602_, new_B8603_, new_B8604_,
    new_B8605_, new_B8606_, new_B8607_, new_B8608_, new_B8609_, new_B8610_,
    new_B8611_, new_B8612_, new_B8613_, new_B8619_, new_B8620_, new_B8621_,
    new_B8622_, new_B8623_, new_B8624_, new_B8625_, new_B8626_, new_B8627_,
    new_B8628_, new_B8629_, new_B8630_, new_B8631_, new_B8632_, new_B8633_,
    new_B8634_, new_B8635_, new_B8636_, new_B8637_, new_B8638_, new_B8639_,
    new_B8640_, new_B8641_, new_B8642_, new_B8643_, new_B8644_, new_B8645_,
    new_B8646_, new_B8652_, new_B8653_, new_B8654_, new_B8655_, new_B8656_,
    new_B8657_, new_B8658_, new_B8659_, new_B8660_, new_B8661_, new_B8662_,
    new_B8663_, new_B8664_, new_B8665_, new_B8666_, new_B8667_, new_B8668_,
    new_B8669_, new_B8670_, new_B8671_, new_B8672_, new_B8673_, new_B8674_,
    new_B8675_, new_B8676_, new_B8677_, new_B8678_, new_B8679_, new_B8685_,
    new_B8686_, new_B8687_, new_B8688_, new_B8689_, new_B8690_, new_B8691_,
    new_B8692_, new_B8693_, new_B8694_, new_B8695_, new_B8696_, new_B8697_,
    new_B8698_, new_B8699_, new_B8700_, new_B8701_, new_B8702_, new_B8703_,
    new_B8704_, new_B8705_, new_B8706_, new_B8707_, new_B8708_, new_B8709_,
    new_B8710_, new_B8711_, new_B8712_, new_B8718_, new_B8719_, new_B8720_,
    new_B8721_, new_B8722_, new_B8723_, new_B8724_, new_B8725_, new_B8726_,
    new_B8727_, new_B8728_, new_B8729_, new_B8730_, new_B8731_, new_B8732_,
    new_B8733_, new_B8734_, new_B8735_, new_B8736_, new_B8737_, new_B8738_,
    new_B8739_, new_B8740_, new_B8741_, new_B8742_, new_B8743_, new_B8744_,
    new_B8745_, new_B8751_, new_B8752_, new_B8753_, new_B8754_, new_B8755_,
    new_B8756_, new_B8757_, new_B8758_, new_B8759_, new_B8760_, new_B8761_,
    new_B8762_, new_B8763_, new_B8764_, new_B8765_, new_B8766_, new_B8767_,
    new_B8768_, new_B8769_, new_B8770_, new_B8771_, new_B8772_, new_B8773_,
    new_B8774_, new_B8775_, new_B8776_, new_B8777_, new_B8778_, new_B8784_,
    new_B8785_, new_B8786_, new_B8787_, new_B8788_, new_B8789_, new_B8790_,
    new_B8791_, new_B8792_, new_B8793_, new_B8794_, new_B8795_, new_B8796_,
    new_B8797_, new_B8798_, new_B8799_, new_B8800_, new_B8801_, new_B8802_,
    new_B8803_, new_B8804_, new_B8805_, new_B8806_, new_B8807_, new_B8808_,
    new_B8809_, new_B8810_, new_B8811_, new_B8817_, new_B8818_, new_B8819_,
    new_B8820_, new_B8821_, new_B8822_, new_B8823_, new_B8824_, new_B8825_,
    new_B8826_, new_B8827_, new_B8828_, new_B8829_, new_B8830_, new_B8831_,
    new_B8832_, new_B8833_, new_B8834_, new_B8835_, new_B8836_, new_B8837_,
    new_B8838_, new_B8839_, new_B8840_, new_B8841_, new_B8842_, new_B8843_,
    new_B8844_, new_B8850_, new_B8851_, new_B8852_, new_B8853_, new_B8854_,
    new_B8855_, new_B8856_, new_B8857_, new_B8858_, new_B8859_, new_B8860_,
    new_B8861_, new_B8862_, new_B8863_, new_B8864_, new_B8865_, new_B8866_,
    new_B8867_, new_B8868_, new_B8869_, new_B8870_, new_B8871_, new_B8872_,
    new_B8873_, new_B8874_, new_B8875_, new_B8876_, new_B8877_, new_B8883_,
    new_B8884_, new_B8885_, new_B8886_, new_B8887_, new_B8888_, new_B8889_,
    new_B8890_, new_B8891_, new_B8892_, new_B8893_, new_B8894_, new_B8895_,
    new_B8896_, new_B8897_, new_B8898_, new_B8899_, new_B8900_, new_B8901_,
    new_B8902_, new_B8903_, new_B8904_, new_B8905_, new_B8906_, new_B8907_,
    new_B8908_, new_B8909_, new_B8910_, new_B8916_, new_B8917_, new_B8918_,
    new_B8919_, new_B8920_, new_B8921_, new_B8922_, new_B8923_, new_B8924_,
    new_B8925_, new_B8926_, new_B8927_, new_B8928_, new_B8929_, new_B8930_,
    new_B8931_, new_B8932_, new_B8933_, new_B8934_, new_B8935_, new_B8936_,
    new_B8937_, new_B8938_, new_B8939_, new_B8940_, new_B8941_, new_B8942_,
    new_B8943_, new_B8949_, new_B8950_, new_B8951_, new_B8952_, new_B8953_,
    new_B8954_, new_B8955_, new_B8956_, new_B8957_, new_B8958_, new_B8959_,
    new_B8960_, new_B8961_, new_B8962_, new_B8963_, new_B8964_, new_B8965_,
    new_B8966_, new_B8967_, new_B8968_, new_B8969_, new_B8970_, new_B8971_,
    new_B8972_, new_B8973_, new_B8974_, new_B8975_, new_B8976_, new_B8982_,
    new_B8983_, new_B8984_, new_B8985_, new_B8986_, new_B8987_, new_B8988_,
    new_B8989_, new_B8990_, new_B8991_, new_B8992_, new_B8993_, new_B8994_,
    new_B8995_, new_B8996_, new_B8997_, new_B8998_, new_B8999_, new_B9000_,
    new_B9001_, new_B9002_, new_B9003_, new_B9004_, new_B9005_, new_B9006_,
    new_B9007_, new_B9008_, new_B9009_, new_B9015_, new_B9016_, new_B9017_,
    new_B9018_, new_B9019_, new_B9020_, new_B9021_, new_B9022_, new_B9023_,
    new_B9024_, new_B9025_, new_B9026_, new_B9027_, new_B9028_, new_B9029_,
    new_B9030_, new_B9031_, new_B9032_, new_B9033_, new_B9034_, new_B9035_,
    new_B9036_, new_B9037_, new_B9038_, new_B9039_, new_B9040_, new_B9041_,
    new_B9042_, new_B9048_, new_B9049_, new_B9050_, new_B9051_, new_B9052_,
    new_B9053_, new_B9054_, new_B9055_, new_B9056_, new_B9057_, new_B9058_,
    new_B9059_, new_B9060_, new_B9061_, new_B9062_, new_B9063_, new_B9064_,
    new_B9065_, new_B9066_, new_B9067_, new_B9068_, new_B9069_, new_B9070_,
    new_B9071_, new_B9072_, new_B9073_, new_B9074_, new_B9075_, new_B9081_,
    new_B9082_, new_B9083_, new_B9084_, new_B9085_, new_B9086_, new_B9087_,
    new_B9088_, new_B9089_, new_B9090_, new_B9091_, new_B9092_, new_B9093_,
    new_B9094_, new_B9095_, new_B9096_, new_B9097_, new_B9098_, new_B9099_,
    new_B9100_, new_B9101_, new_B9102_, new_B9103_, new_B9104_, new_B9105_,
    new_B9106_, new_B9107_, new_B9108_, new_B9114_, new_B9115_, new_B9116_,
    new_B9117_, new_B9118_, new_B9119_, new_B9120_, new_B9121_, new_B9122_,
    new_B9123_, new_B9124_, new_B9125_, new_B9126_, new_B9127_, new_B9128_,
    new_B9129_, new_B9130_, new_B9131_, new_B9132_, new_B9133_, new_B9134_,
    new_B9135_, new_B9136_, new_B9137_, new_B9138_, new_B9139_, new_B9140_,
    new_B9141_, new_B9147_, new_B9148_, new_B9149_, new_B9150_, new_B9151_,
    new_B9152_, new_B9153_, new_B9154_, new_B9155_, new_B9156_, new_B9157_,
    new_B9158_, new_B9159_, new_B9160_, new_B9161_, new_B9162_, new_B9163_,
    new_B9164_, new_B9165_, new_B9166_, new_B9167_, new_B9168_, new_B9169_,
    new_B9170_, new_B9171_, new_B9172_, new_B9173_, new_B9174_, new_B9180_,
    new_B9181_, new_B9182_, new_B9183_, new_B9184_, new_B9185_, new_B9186_,
    new_B9187_, new_B9188_, new_B9189_, new_B9190_, new_B9191_, new_B9192_,
    new_B9193_, new_B9194_, new_B9195_, new_B9196_, new_B9197_, new_B9198_,
    new_B9199_, new_B9200_, new_B9201_, new_B9202_, new_B9203_, new_B9204_,
    new_B9205_, new_B9206_, new_B9207_, new_B9213_, new_B9214_, new_B9215_,
    new_B9216_, new_B9217_, new_B9218_, new_B9219_, new_B9220_, new_B9221_,
    new_B9222_, new_B9223_, new_B9224_, new_B9225_, new_B9226_, new_B9227_,
    new_B9228_, new_B9229_, new_B9230_, new_B9231_, new_B9232_, new_B9233_,
    new_B9234_, new_B9235_, new_B9236_, new_B9237_, new_B9238_, new_B9239_,
    new_B9240_, new_B9246_, new_B9247_, new_B9248_, new_B9249_, new_B9250_,
    new_B9251_, new_B9252_, new_B9253_, new_B9254_, new_B9255_, new_B9256_,
    new_B9257_, new_B9258_, new_B9259_, new_B9260_, new_B9261_, new_B9262_,
    new_B9263_, new_B9264_, new_B9265_, new_B9266_, new_B9267_, new_B9268_,
    new_B9269_, new_B9270_, new_B9271_, new_B9272_, new_B9273_, new_B9279_,
    new_B9280_, new_B9281_, new_B9282_, new_B9283_, new_B9284_, new_B9285_,
    new_B9286_, new_B9287_, new_B9288_, new_B9289_, new_B9290_, new_B9291_,
    new_B9292_, new_B9293_, new_B9294_, new_B9295_, new_B9296_, new_B9297_,
    new_B9298_, new_B9299_, new_B9300_, new_B9301_, new_B9302_, new_B9303_,
    new_B9304_, new_B9305_, new_B9306_, new_B1089_, new_B1088_, new_B1087_,
    new_B1086_, new_B1085_, new_B1084_, new_B1083_, new_B1082_, new_B1081_,
    new_B1080_, new_B1079_, new_B1078_, new_B1077_, new_B1076_, new_B1075_,
    new_B1074_, new_B1073_, new_B1072_, new_B1071_, new_B1070_, new_B1069_,
    new_B1068_, new_B1067_, new_B1066_, new_B1065_, new_B1064_, new_B1063_,
    new_B1062_, new_B1061_, new_B1060_, new_B1059_, new_B1058_, new_B1057_,
    new_B1090_, new_B1091_, new_B1092_, new_B1093_, new_B1094_, new_B1095_,
    new_B1096_, new_B1097_, new_B1098_, new_B1099_, new_B1100_, new_B1101_,
    new_B1102_, new_B1103_, new_B1104_, new_B1105_, new_B1106_, new_B1107_,
    new_B1108_, new_B1109_, new_B1110_, new_B1111_, new_B1112_, new_B1113_,
    new_B1114_, new_B1115_, new_B1116_, new_B1117_, new_B1118_, new_B1119_,
    new_B1120_, new_B1121_, new_B1122_, new_B1123_, new_B1124_, new_B1125_,
    new_B1126_, new_B1127_, new_B1128_, new_B1129_, new_B1130_, new_B1131_,
    new_B1132_, new_B1133_, new_B1134_, new_B1135_, new_B1136_, new_B1137_,
    new_B1138_, new_B1139_, new_B1140_, new_B1141_, new_B1142_, new_B1143_,
    new_B1144_, new_B1145_, new_B1146_, new_B1147_, new_B1148_, new_B1149_,
    new_B1150_, new_B1151_, new_B1152_, new_B1153_, new_B1154_, new_B1155_,
    new_B1156_, new_B1157_, new_B1158_, new_B1159_, new_B1160_, new_B1161_,
    new_B1162_, new_B1163_, new_B1164_, new_B1165_, new_B1166_, new_B1167_,
    new_B1168_, new_B1169_, new_B1170_, new_B1171_, new_B1172_, new_B1173_,
    new_B1174_, new_B1175_, new_B1176_, new_B1177_, new_B1178_, new_B1179_,
    new_B1180_, new_B1181_, new_B1182_, new_B1183_, new_B1184_, new_B1185_,
    new_B1186_, new_B1187_, new_B1188_, new_B1189_, new_B1190_, new_B1191_,
    new_B1192_, new_B1193_, new_B1194_, new_B1195_, new_B1196_, new_B1197_,
    new_B1198_, new_B1199_, new_B1200_, new_B1201_, new_B1202_, new_B1203_,
    new_B1204_, new_B1205_, new_B1206_, new_B1207_, new_B1208_, new_B1209_,
    new_B1210_, new_B1211_, new_B1212_, new_B1213_, new_B1214_, new_B1215_,
    new_B1216_, new_B1217_, new_B1218_, new_B1219_, new_B1220_, new_B1221_,
    new_B1222_, new_B1223_, new_B1224_, new_B1225_, new_B1226_, new_B1227_,
    new_B1228_, new_B1229_, new_B1230_, new_B1231_, new_B1232_, new_B1233_,
    new_B1234_, new_B1235_, new_B1236_, new_B1237_, new_B1238_, new_B1239_,
    new_B1240_, new_B1241_, new_B1242_, new_B1243_, new_B1244_, new_B1245_,
    new_B1246_, new_B1247_, new_B1248_, new_B1249_, new_B1250_, new_B1251_,
    new_B1252_, new_B1253_, new_B1254_, new_B1255_, new_B1256_, new_B1257_,
    new_B1258_, new_B1259_, new_B1260_, new_B1261_, new_B1262_, new_B1263_,
    new_B1264_, new_B1265_, new_B1266_, new_B1267_, new_B1268_, new_B1269_,
    new_B1270_, new_B1271_, new_B1272_, new_B1273_, new_B1274_, new_B1275_,
    new_B1276_, new_B1277_, new_B1278_, new_B1279_, new_B1280_, new_B1281_,
    new_B1282_, new_B1283_, new_B1284_, new_B1285_, new_B1286_, new_B1287_,
    new_B1288_, new_B1289_, new_B1290_, new_B1291_, new_B1292_, new_B1293_,
    new_B1294_, new_B1295_, new_B1296_, new_B1297_, new_B1298_, new_B1299_,
    new_B1300_, new_B1301_, new_B1302_, new_B1303_, new_B1304_, new_B1305_,
    new_B1306_, new_B1307_, new_B1308_, new_B1309_, new_B1310_, new_B1311_,
    new_B1312_, new_B1313_, new_B1314_, new_B1315_, new_B1316_, new_B1317_,
    new_B1318_, new_B1319_, new_B1320_, new_B1321_, new_B1322_, new_B1323_,
    new_B1324_, new_B1325_, new_B1326_, new_B1327_, new_B1328_, new_B1329_,
    new_B1330_, new_B1331_, new_B1332_, new_B1333_, new_B1334_, new_B1335_,
    new_B1336_, new_B1337_, new_B1338_, new_B1339_, new_B1340_, new_B1341_,
    new_B1342_, new_B1343_, new_B1344_, new_B1345_, new_B1346_, new_B1347_,
    new_B1348_, new_B1349_, new_B1350_, new_B1351_, new_B1352_, new_B1353_,
    new_B1354_, new_B1355_, new_B1356_, new_B1357_, new_B1358_, new_B1359_,
    new_B1360_, new_B1361_, new_B1362_, new_B1363_, new_B1364_, new_B1365_,
    new_B1366_, new_B1367_, new_B1368_, new_B1369_, new_B1370_, new_B1371_,
    new_B1372_, new_B1373_, new_B1374_, new_B1375_, new_B1376_, new_B1377_,
    new_B1378_, new_B1379_, new_B1380_, new_B1381_, new_B1382_, new_B1383_,
    new_B1384_, new_B1385_, new_B1386_, new_B1387_, new_B1388_, new_B1389_,
    new_B1390_, new_B1391_, new_B1392_, new_B1393_, new_B1394_, new_B1395_,
    new_B1396_, new_B1397_, new_B1398_, new_B1399_, new_B1400_, new_B1401_,
    new_B1402_, new_B1403_, new_B1404_, new_B1405_, new_B1406_, new_B1407_,
    new_B1408_, new_B1409_, new_B1410_, new_B1411_, new_B1412_, new_B1413_,
    new_B1414_, new_B1415_, new_B1416_, new_B1417_, new_B1418_, new_B1419_,
    new_B1420_, new_B1421_, new_B1422_, new_B1423_, new_B1424_, new_B1425_,
    new_B1426_, new_B1427_, new_B1428_, new_B1429_, new_B1430_, new_B1431_,
    new_B1432_, new_B1433_, new_B1434_, new_B1435_, new_B1436_, new_B1437_,
    new_B1438_, new_B1439_, new_B1440_, new_B1441_, new_B1442_, new_B1443_,
    new_B1444_, new_B1445_, new_B1446_, new_B1447_, new_B1448_, new_B1449_,
    new_B1450_, new_B1451_, new_B1452_, new_B1453_, new_B1454_, new_B1455_,
    new_B1456_, new_B1457_, new_B1458_, new_B1459_, new_B1460_, new_B1461_,
    new_B1462_, new_B1463_, new_B1464_, new_B1465_, new_B1466_, new_B1467_,
    new_B1468_, new_B1469_, new_B1470_, new_B1471_, new_B1472_, new_B1473_,
    new_B1474_, new_B1475_, new_B1476_, new_B1477_, new_B1478_, new_B1479_,
    new_B1480_, new_B1481_, new_B1482_, new_B1483_, new_B1484_, new_B1485_,
    new_B1486_, new_B1487_, new_B1488_, new_B1489_, new_B1490_, new_B1491_,
    new_B1492_, new_B1493_, new_B1494_, new_B1495_, new_B1496_, new_B1497_,
    new_B1498_, new_B1499_, new_B1500_, new_B1501_, new_B1502_, new_B1503_,
    new_B1504_, new_B1505_, new_B1506_, new_B1507_, new_B1508_, new_B1509_,
    new_B1510_, new_B1511_, new_B1512_, new_B1513_, new_B1514_, new_B1515_,
    new_B1516_, new_B1517_, new_B1518_, new_B1519_, new_B1520_, new_B1521_,
    new_B1522_, new_B1523_, new_B1524_, new_B1525_, new_B1526_, new_B1527_,
    new_B1528_, new_B1529_, new_B1530_, new_B1531_, new_B1532_, new_B1533_,
    new_B1534_, new_B1535_, new_B1536_, new_B1537_, new_B1538_, new_B1539_,
    new_B1540_, new_B1541_, new_B1542_, new_B1543_, new_B1544_, new_B1545_,
    new_B1546_, new_B1547_, new_B1548_, new_B1549_, new_B1550_, new_B1551_,
    new_B1552_, new_B1553_, new_B1554_, new_B1555_, new_B1556_, new_B1557_,
    new_B1558_, new_B1559_, new_B1560_, new_B1561_, new_B1562_, new_B1563_,
    new_B1564_, new_B1565_, new_B1566_, new_B1567_, new_B1568_, new_B1569_,
    new_B1570_, new_B1571_, new_B1572_, new_B1573_, new_B1574_, new_B1575_,
    new_B1576_, new_B1577_, new_B1578_, new_B1579_, new_B1580_, new_B1581_,
    new_B1582_, new_B1583_, new_B1584_, new_B1585_, new_B1586_, new_B1587_,
    new_B1588_, new_B1589_, new_B1590_, new_B1591_, new_B1592_, new_B1593_,
    new_B1594_, new_B1595_, new_B1596_, new_B1597_, new_B1598_, new_B1599_,
    new_B1600_, new_B1601_, new_B1602_, new_B1603_, new_B1604_, new_B1605_,
    new_B1606_, new_B1607_, new_B1608_, new_B1609_, new_B1610_, new_B1611_,
    new_B1612_, new_B1613_, new_B1614_, new_B1615_, new_B1616_, new_B1617_,
    new_B1618_, new_B1619_, new_B1620_, new_B1621_, new_B1622_, new_B1623_,
    new_B1624_, new_B1625_, new_B1626_, new_B1627_, new_B1628_, new_B1629_,
    new_B1630_, new_B1631_, new_B1632_, new_B1633_, new_B1634_, new_B1635_,
    new_B1636_, new_B1637_, new_B1638_, new_B1639_, new_B1640_, new_B1641_,
    new_B1642_, new_B1643_, new_B1644_, new_B1645_, new_B1646_, new_B1647_,
    new_B1648_, new_B1649_, new_B1650_, new_B1651_, new_B1652_, new_B1653_,
    new_B1654_, new_B1655_, new_B1656_, new_B1657_, new_B1658_, new_B1659_,
    new_B1660_, new_B1661_, new_B1662_, new_B1663_, new_B1664_, new_B1665_,
    new_B1666_, new_B1667_, new_B1668_, new_B1669_, new_B1670_, new_B1671_,
    new_B1672_, new_B1673_, new_B1674_, new_B1675_, new_B1676_, new_B1677_,
    new_B1678_, new_B1679_, new_B1680_, new_B1681_, new_B1682_, new_B1683_,
    new_B1684_, new_B1685_, new_B1686_, new_B1687_, new_B1688_, new_B1689_,
    new_B1690_, new_B1691_, new_B1692_, new_B1693_, new_B1694_, new_B1695_,
    new_B1696_, new_B1697_, new_B1698_, new_B1699_, new_B1700_, new_B1701_,
    new_B1702_, new_B1703_, new_B1704_, new_B1705_, new_B1706_, new_B1707_,
    new_B1708_, new_B1709_, new_B1710_, new_B1711_, new_B1712_, new_B1713_,
    new_B1714_, new_B1715_, new_B1716_, new_B1717_, new_B1718_, new_B1719_,
    new_B1720_, new_B1721_, new_B1722_, new_B1723_, new_B1724_, new_B1725_,
    new_B1726_, new_B1727_, new_B1728_, new_B1729_, new_B1730_, new_B1731_,
    new_B1732_, new_B1733_, new_B1734_, new_B1735_, new_B1736_, new_B1737_,
    new_B1738_, new_B1739_, new_B1740_, new_B1741_, new_B1742_, new_B1743_,
    new_B1744_, new_B1745_, new_B1746_, new_B1747_, new_B1748_, new_B1749_,
    new_B1750_, new_B1751_, new_B1752_, new_B1753_, new_B1754_, new_B1755_,
    new_B1756_, new_B1757_, new_B1758_, new_B1759_, new_B1760_, new_B1761_,
    new_B1762_, new_B1763_, new_B1764_, new_B1765_, new_B1766_, new_B1767_,
    new_B1768_, new_B1769_, new_B1770_, new_B1771_, new_B1772_, new_B1773_,
    new_B1774_, new_B1775_, new_B1776_, new_B1777_, new_B1778_, new_B1779_,
    new_B1780_, new_B1781_, new_B1782_, new_B1783_, new_B1784_, new_B1785_,
    new_B1786_, new_B1787_, new_B1788_, new_B1789_, new_B1790_, new_B1791_,
    new_B1792_, new_B1793_, new_B1794_, new_B1795_, new_B1796_, new_B1797_,
    new_B1798_, new_B1799_, new_B1800_, new_B1801_, new_B1802_, new_B1803_,
    new_B1804_, new_B1805_, new_B1806_, new_B1807_, new_B1808_, new_B1809_,
    new_B1810_, new_B1811_, new_B1812_, new_B1813_, new_B1814_, new_B1815_,
    new_B1816_, new_B1817_, new_B1818_, new_B1819_, new_B1820_, new_B1821_,
    new_B1822_, new_B1823_, new_B1824_, new_B1825_, new_B1826_, new_B1827_,
    new_B1828_, new_B1829_, new_B1830_, new_B1831_, new_B1832_, new_B1833_,
    new_B1834_, new_B1835_, new_B1836_, new_B1837_, new_B1838_, new_B1839_,
    new_B1840_, new_B1841_, new_B1842_, new_B1843_, new_B1844_, new_B1845_,
    new_B1846_, new_B1847_, new_B1848_, new_B1849_, new_B1850_, new_B1851_,
    new_B1852_, new_B1853_, new_B1854_, new_B1855_, new_B1856_, new_B1857_,
    new_B1858_, new_B1859_, new_B1860_, new_B1861_, new_B1862_, new_B1863_,
    new_B1864_, new_B1865_, new_B1866_, new_B1867_, new_B1868_, new_B1869_,
    new_B1870_, new_B1871_, new_B1872_, new_B1873_, new_B1874_, new_B1875_,
    new_B1876_, new_B1877_, new_B1878_, new_B1879_, new_B1880_, new_B1881_,
    new_B1882_, new_B1883_, new_B1884_, new_B1885_, new_B1886_, new_B1887_,
    new_B1888_, new_B1889_, new_B1890_, new_B1891_, new_B1892_, new_B1893_,
    new_B1894_, new_B1895_, new_B1896_, new_B1897_, new_B1898_, new_B1899_,
    new_B1900_, new_B1901_, new_B1902_, new_B1903_, new_B1904_, new_B1905_,
    new_B1906_, new_B1907_, new_B1908_, new_B1909_, new_B1910_, new_B1911_,
    new_B1912_, new_B1913_, new_B1914_, new_B1915_, new_B1916_, new_B1917_,
    new_B1918_, new_B1919_, new_B1920_, new_B1921_, new_B1922_, new_B1923_,
    new_B1924_, new_B1925_, new_B1926_, new_B1927_, new_B1928_, new_B1929_,
    new_B1930_, new_B1931_, new_B1932_, new_B1933_, new_B1934_, new_B1935_,
    new_B1936_, new_B1937_, new_B1938_, new_B1939_, new_B1940_, new_B1941_,
    new_B1942_, new_B1943_, new_B1944_, new_B1945_, new_B1946_, new_B1947_,
    new_B1948_, new_B1949_, new_B1950_, new_B1951_, new_B1952_, new_B1953_,
    new_B1954_, new_B1955_, new_B1956_, new_B1957_, new_B1958_, new_B1959_,
    new_B1960_, new_B1961_, new_B1962_, new_B1963_, new_B1964_, new_B1965_,
    new_B1966_, new_B1967_, new_B1968_, new_B1969_, new_B1970_, new_B1971_,
    new_B1972_, new_B1973_, new_B1974_, new_B1975_, new_B1976_, new_B1977_,
    new_B1978_, new_B1979_, new_B1980_, new_B1981_, new_B1982_, new_B1983_,
    new_B1984_, new_B1985_, new_B1986_, new_B1987_, new_B1988_, new_B1989_,
    new_B1990_, new_B1991_, new_B1992_, new_B1993_, new_B1994_, new_B1995_,
    new_B1996_, new_B1997_, new_B1998_, new_B1999_, new_B2000_, new_B2001_,
    new_B2002_, new_B2003_, new_B2004_, new_B2005_, new_B2006_, new_B2007_,
    new_B2008_, new_B2009_, new_B2010_, new_B2011_, new_B2012_, new_B2013_,
    new_B2014_, new_B2015_, new_B2016_, new_B2017_, new_B2018_, new_B2019_,
    new_B2020_, new_B2021_, new_B2022_, new_B2023_, new_B2024_, new_B2025_,
    new_B2026_, new_B2027_, new_B2028_, new_B2029_, new_B2030_, new_B2031_,
    new_B2032_, new_B2033_, new_B2034_, new_B2035_, new_B2036_, new_B2037_,
    new_B2038_, new_B2039_, new_B2040_, new_B2041_, new_B2042_, new_B2043_,
    new_B2044_, new_B2045_, new_B2046_, new_B2047_, new_B2048_, new_B2049_,
    new_B2050_, new_B2051_, new_B2052_, new_B2053_, new_B2054_, new_B2055_,
    new_B2056_, new_B2057_, new_B2058_, new_B2059_, new_B2060_, new_B2061_,
    new_B2062_, new_B2063_, new_B2064_, new_B2065_, new_B2066_, new_B2067_,
    new_B2068_, new_B2069_, new_B2070_, new_B2071_, new_B2072_, new_B2073_,
    new_B2074_, new_B2075_, new_B2076_, new_B2077_, new_B2078_, new_B2079_,
    new_B2080_, new_B2081_, new_B2082_, new_B2083_, new_B2084_, new_B2085_,
    new_B2086_, new_B2087_, new_B2088_, new_B2089_, new_B2090_, new_B2091_,
    new_B2092_, new_B2093_, new_B2094_, new_B2095_, new_B2096_, new_B2097_,
    new_B2098_, new_B2099_, new_B2100_, new_B2101_, new_B2102_, new_B2103_,
    new_B2104_, new_B2105_, new_B2106_, new_B2107_, new_B2108_, new_B2109_,
    new_B2110_, new_B2111_, new_B2112_, new_B2113_, new_B2114_, new_B2115_,
    new_B2116_, new_B2117_, new_B2118_, new_B2119_, new_B2120_, new_B2121_,
    new_B2122_, new_B2123_, new_B2124_, new_B2125_, new_B2126_, new_B2127_,
    new_B2128_, new_B2129_, new_B2130_, new_B2131_, new_B2132_, new_B2133_,
    new_B2134_, new_B2135_, new_B2136_, new_B2137_, new_B2138_, new_B2139_,
    new_B2140_, new_B2141_, new_B2142_, new_B2143_, new_B2144_, new_B2145_,
    new_B2146_, new_B2147_, new_B2148_, new_B2149_, new_B2150_, new_B2151_,
    new_B2152_, new_B2153_, new_B2154_, new_B2155_, new_B2156_, new_B2157_,
    new_B2158_, new_B2159_, new_B2160_, new_B2161_, new_B2162_, new_B2163_,
    new_B2164_, new_B2165_, new_B2166_, new_B2167_, new_B2168_, new_B2169_,
    new_B2170_, new_B2171_, new_B2172_, new_B2173_, new_B2174_, new_B2175_,
    new_B2176_, new_B2177_, new_B2178_, new_B2179_, new_B2180_, new_B2181_,
    new_B2182_, new_B2183_, new_B2184_, new_B2185_, new_B2186_, new_B2187_,
    new_B2188_, new_B2189_, new_B2190_, new_B2191_, new_B2192_, new_B2193_,
    new_B2194_, new_B2195_, new_B2196_, new_B2197_, new_B2198_, new_B2199_,
    new_B2200_, new_B2201_, new_B2202_, new_B2203_, new_B2204_, new_B2205_,
    new_B2206_, new_B2207_, new_B2208_, new_B2209_, new_B2210_, new_B2211_,
    new_B2212_, new_B2213_, new_B2214_, new_B2215_, new_B2216_, new_B2217_,
    new_B2218_, new_B2219_, new_B2220_, new_B2221_, new_B2222_, new_B2223_,
    new_B2224_, new_B2225_, new_B2226_, new_B2227_, new_B2228_, new_B2229_,
    new_B2230_, new_B2231_, new_B2232_, new_B2233_, new_B2234_, new_B2235_,
    new_B2236_, new_B2237_, new_B2238_, new_B2239_, new_B2240_, new_B2241_,
    new_B2242_, new_B2243_, new_B2244_, new_B2245_, new_B2246_, new_B2247_,
    new_B2248_, new_B2249_, new_B2250_, new_B2251_, new_B2252_, new_B2253_,
    new_B2254_, new_B2255_, new_B2256_, new_B2257_, new_B2258_, new_B2259_,
    new_B2260_, new_B2261_, new_B2262_, new_B2263_, new_B2264_, new_B2265_,
    new_B2266_, new_B2267_, new_B2268_, new_B2269_, new_B2270_, new_B2271_,
    new_B2272_, new_B2273_, new_B2274_, new_B2275_, new_B2276_, new_B2277_,
    new_B2278_, new_B2279_, new_B2280_, new_B2281_, new_B2282_, new_B2283_,
    new_B2284_, new_B2285_, new_B2286_, new_B2287_, new_B2288_, new_B2289_,
    new_B2290_, new_B2291_, new_B2292_, new_B2293_, new_B2294_, new_B2295_,
    new_B2296_, new_B2297_, new_B2298_, new_B2299_, new_B2300_, new_B2301_,
    new_B2302_, new_B2303_, new_B2304_, new_B2305_, new_B2306_, new_B2307_,
    new_B2308_, new_B2309_, new_B2310_, new_B2311_, new_B2312_, new_B2313_,
    new_B2314_, new_B2315_, new_B2316_, new_B2317_, new_B2318_, new_B2319_,
    new_B2320_, new_B2321_, new_B2322_, new_B2323_, new_B2324_, new_B2325_,
    new_B2326_, new_B2327_, new_B2328_, new_B2329_, new_B2330_, new_B2331_,
    new_B2332_, new_B2333_, new_B2334_, new_B2335_, new_B2336_, new_B2337_,
    new_B2338_, new_B2339_, new_B2340_, new_B2341_, new_B2342_, new_B2343_,
    new_B2344_, new_B2345_, new_B2346_, new_B2347_, new_B2348_, new_B2349_,
    new_B2350_, new_B2351_, new_B2352_, new_B2353_, new_B2354_, new_B2355_,
    new_B2356_, new_B2357_, new_B2358_, new_B2359_, new_B2360_, new_B2361_,
    new_B2362_, new_B2363_, new_B2364_, new_B2365_, new_B2366_, new_B2367_,
    new_B2368_, new_B2369_, new_B2370_, new_B2371_, new_B2372_, new_B2373_,
    new_B2374_, new_B2375_, new_B2376_, new_B2377_, new_B2378_, new_B2379_,
    new_B2380_, new_B2381_, new_B2382_, new_B2383_, new_B2384_, new_B2385_,
    new_B2386_, new_B2387_, new_B2388_, new_B2389_, new_B2390_, new_B2391_,
    new_B2392_, new_B2393_, new_B2394_, new_B2395_, new_B2396_, new_B2397_,
    new_B2398_, new_B2399_, new_B2400_, new_B2401_, new_B2402_, new_B2403_,
    new_B2404_, new_B2405_, new_B2406_, new_B2407_, new_B2408_, new_B2409_,
    new_B2410_, new_B2411_, new_B2412_, new_B2413_, new_B2414_, new_B2415_,
    new_B2416_, new_B2417_, new_B2418_, new_B2419_, new_B2420_, new_B2421_,
    new_B2422_, new_B2423_, new_B2424_, new_B2425_, new_B2426_, new_B2427_,
    new_B2428_, new_B2429_, new_B2430_, new_B2431_, new_B2432_, new_B2433_,
    new_B2434_, new_B2435_, new_B2436_, new_B2437_, new_B2438_, new_B2439_,
    new_B2440_, new_B2441_, new_B2442_, new_B2443_, new_B2444_, new_B2445_,
    new_B2446_, new_B2447_, new_B2448_, new_B2449_, new_B2450_, new_B2451_,
    new_B2452_, new_B2453_, new_B2454_, new_B2455_, new_B2456_, new_B2457_,
    new_B2458_, new_B2459_, new_B2460_, new_B2461_, new_B2462_, new_B2463_,
    new_B2464_, new_B2465_, new_B2466_, new_B2467_, new_B2468_, new_B2469_,
    new_B2470_, new_B2471_, new_B2472_, new_B2473_, new_B2474_, new_B2475_,
    new_B2476_, new_B2477_, new_B2478_, new_B2479_, new_B2480_, new_B2481_,
    new_B2482_, new_B2483_, new_B2484_, new_B2485_, new_B2486_, new_B2487_,
    new_B2488_, new_B2489_, new_B2490_, new_B2491_, new_B2492_, new_B2493_,
    new_B2494_, new_B2495_, new_B2496_, new_B2497_, new_B2498_, new_B2499_,
    new_B2500_, new_B2501_, new_B2502_, new_B2503_, new_B2504_, new_B2505_,
    new_B2506_, new_B2507_, new_B2508_, new_B2509_, new_B2510_, new_B2511_,
    new_B2512_, new_B2513_, new_B2514_, new_B2515_, new_B2516_, new_B2517_,
    new_B2518_, new_B2519_, new_B2520_, new_B2521_, new_B2522_, new_B2523_,
    new_B2524_, new_B2525_, new_B2526_, new_B2527_, new_B2528_, new_B2529_,
    new_B2530_, new_B2531_, new_B2532_, new_B2533_, new_B2534_, new_B2535_,
    new_B2536_, new_B2537_, new_B2538_, new_B2539_, new_B2540_, new_B2541_,
    new_B2542_, new_B2543_, new_B2544_, new_B2545_, new_B2546_, new_B2547_,
    new_B2548_, new_B2549_, new_B2550_, new_B2551_, new_B2552_, new_B2553_,
    new_B2554_, new_B2555_, new_B2556_, new_B2557_, new_B2558_, new_B2559_,
    new_B2560_, new_B2561_, new_B2562_, new_B2563_, new_B2564_, new_B2565_,
    new_B2566_, new_B2567_, new_B2568_, new_B2569_, new_B2570_, new_B2571_,
    new_B2572_, new_B2573_, new_B2574_, new_B2575_, new_B2576_, new_B2577_,
    new_B2578_, new_B2579_, new_B2580_, new_B2581_, new_B2582_, new_B2583_,
    new_B2584_, new_B2585_, new_B2586_, new_B2587_, new_B2588_, new_B2589_,
    new_B2590_, new_B2591_, new_B2592_, new_B2593_, new_B2594_, new_B2595_,
    new_B2596_, new_B2597_, new_B2598_, new_B2599_, new_B2600_, new_B2601_,
    new_B2602_, new_B2603_, new_B2604_, new_B2605_, new_B2606_, new_B2607_,
    new_B2608_, new_B2609_, new_B2610_, new_B2611_, new_B2612_, new_B2613_,
    new_B2614_, new_B2615_, new_B2616_, new_B2617_, new_B2618_, new_B2619_,
    new_B2620_, new_B2621_, new_B2622_, new_B2623_, new_B2624_, new_B2625_,
    new_B2626_, new_B2627_, new_B2628_, new_B2629_, new_B2630_, new_B2631_,
    new_B2632_, new_B2633_, new_B2634_, new_B2635_, new_B2636_, new_B2637_,
    new_B2638_, new_B2639_, new_B2640_, new_B2641_, new_B2642_, new_B2643_,
    new_B2644_, new_B2645_, new_B2646_, new_B2647_, new_B2648_, new_B2649_,
    new_B2650_, new_B2651_, new_B2652_, new_B2653_, new_B2654_, new_B2655_,
    new_B2656_, new_B2657_, new_B2658_, new_B2659_, new_B2660_, new_B2661_,
    new_B2662_, new_B2663_, new_B2664_, new_B2665_, new_B2666_, new_B2667_,
    new_B2668_, new_B2669_, new_B2670_, new_B2671_, new_B2672_, new_B2673_,
    new_B2674_, new_B2675_, new_B2676_, new_B2677_, new_B2678_, new_B2679_,
    new_B2680_, new_B2681_, new_B2682_, new_B2683_, new_B2684_, new_B2685_,
    new_B2686_, new_B2687_, new_B2688_, new_B2689_, new_B2690_, new_B2691_,
    new_B2692_, new_B2693_, new_B2694_, new_B2695_, new_B2696_, new_B2697_,
    new_B2698_, new_B2699_, new_B2700_, new_B2701_, new_B2702_, new_B2703_,
    new_B2704_, new_B2705_, new_B2706_, new_B2707_, new_B2708_, new_B2709_,
    new_B2710_, new_B2711_, new_B2712_, new_B2713_, new_B2714_, new_B2715_,
    new_B2716_, new_B2717_, new_B2718_, new_B2719_, new_B2720_, new_B2721_,
    new_B2722_, new_B2723_, new_B2724_, new_B2725_, new_B2726_, new_B2727_,
    new_B2728_, new_B2729_, new_B2730_, new_B2731_, new_B2732_, new_B2733_,
    new_B2734_, new_B2735_, new_B2736_, new_B2737_, new_B2738_, new_B2739_,
    new_B2740_, new_B2741_, new_B2742_, new_B2743_, new_B2744_, new_B2745_,
    new_B2746_, new_B2747_, new_B2748_, new_B2749_, new_B2750_, new_B2751_,
    new_B2752_, new_B2753_, new_B2754_, new_B2755_, new_B2756_, new_B2757_,
    new_B2758_, new_B2759_, new_B2760_, new_B2761_, new_B2762_, new_B2763_,
    new_B2764_, new_B2765_, new_B2766_, new_B2767_, new_B2768_, new_B2769_,
    new_B2770_, new_B2771_, new_B2772_, new_B2773_, new_B2774_, new_B2775_,
    new_B2776_, new_B2777_, new_B2778_, new_B2779_, new_B2780_, new_B2781_,
    new_B2782_, new_B2783_, new_B2784_, new_B2785_, new_B2786_, new_B2787_,
    new_B2788_, new_B2789_, new_B2790_, new_B2791_, new_B2792_, new_B2793_,
    new_B2794_, new_B2795_, new_B2796_, new_B2797_, new_B2798_, new_B2799_,
    new_B2800_, new_B2801_, new_B2802_, new_B2803_, new_B2804_, new_B2805_,
    new_B2806_, new_B2807_, new_B2808_, new_B2809_, new_B2810_, new_B2811_,
    new_B2812_, new_B2813_, new_B2814_, new_B2815_, new_B2816_, new_B2817_,
    new_B2818_, new_B2819_, new_B2820_, new_B2821_, new_B2822_, new_B2823_,
    new_B2824_, new_B2825_, new_B2826_, new_B2827_, new_B2828_, new_B2829_,
    new_B2830_, new_B2831_, new_B2832_, new_B2833_, new_B2834_, new_B2835_,
    new_B2836_, new_B2837_, new_B2838_, new_B2839_, new_B2840_, new_B2841_,
    new_B2842_, new_B2843_, new_B2844_, new_B2845_, new_B2846_, new_B2847_,
    new_B2848_, new_B2849_, new_B2850_, new_B2851_, new_B2852_, new_B2853_,
    new_B2854_, new_B2855_, new_B2856_, new_B2857_, new_B2858_, new_B2859_,
    new_B2860_, new_B2861_, new_B2862_, new_B2863_, new_B2864_, new_B2865_,
    new_B2866_, new_B2867_, new_B2868_, new_B2869_, new_B2870_, new_B2871_,
    new_B2872_, new_B2873_, new_B2874_, new_B2875_, new_B2876_, new_B2877_,
    new_B2878_, new_B2879_, new_B2880_, new_B2881_, new_B2882_, new_B2883_,
    new_B2884_, new_B2885_, new_B2886_, new_B2887_, new_B2888_, new_B2889_,
    new_B2890_, new_B2891_, new_B2892_, new_B2893_, new_B2894_, new_B2895_,
    new_B2896_, new_B2897_, new_B2898_, new_B2899_, new_B2900_, new_B2901_,
    new_B2902_, new_B2903_, new_B2904_, new_B2905_, new_B2906_, new_B2907_,
    new_B2908_, new_B2909_, new_B2910_, new_B2911_, new_B2912_, new_B2913_,
    new_B2914_, new_B2915_, new_B2916_, new_B2917_, new_B2918_, new_B2919_,
    new_B2920_, new_B2921_, new_B2922_, new_B2923_, new_B2924_, new_B2925_,
    new_B2926_, new_B2927_, new_B2928_, new_B2929_, new_B2930_, new_B2931_,
    new_B2932_, new_B2933_, new_B2934_, new_B2935_, new_B2936_, new_B2937_,
    new_B2938_, new_B2939_, new_B2940_, new_B2941_, new_B2942_, new_B2943_,
    new_B2944_, new_B2945_, new_B2946_, new_B2947_, new_B2948_, new_B2949_,
    new_B2950_, new_B2951_, new_B2952_, new_B2953_, new_B2954_, new_B2955_,
    new_B2956_, new_B2957_, new_B2958_, new_B2959_, new_B2960_, new_B2961_,
    new_B2962_, new_B2963_, new_B2964_, new_B2965_, new_B2966_, new_B2967_,
    new_B2968_, new_B2969_, new_B2970_, new_B2971_, new_B2972_, new_B2973_,
    new_B2974_, new_B2975_, new_B2976_, new_B2977_, new_B2978_, new_B2979_,
    new_B2980_, new_B2981_, new_B2982_, new_B2983_, new_B2984_, new_B2985_,
    new_B2986_, new_B2987_, new_B2988_, new_B2989_, new_B2990_, new_B2991_,
    new_B2992_, new_B2993_, new_B2994_, new_B2995_, new_B2996_, new_B2997_,
    new_B2998_, new_B2999_, new_B3000_, new_B3001_, new_B3002_, new_B3003_,
    new_B3004_, new_B3005_, new_B3006_, new_B3007_, new_B3008_, new_B3009_,
    new_B3010_, new_B3011_, new_B3012_, new_B3013_, new_B3014_, new_B3015_,
    new_B3016_, new_B3017_, new_B3018_, new_B3019_, new_B3020_, new_B3021_,
    new_B3022_, new_B3023_, new_B3024_, new_B3025_, new_B3026_, new_B3027_,
    new_B3028_, new_B3029_, new_B3030_, new_B3031_, new_B3032_, new_B3033_,
    new_B3034_, new_B3035_, new_B3036_, new_B3037_, new_B3038_, new_B3039_,
    new_B3040_, new_B3041_, new_B3042_, new_B3043_, new_B3044_, new_B3045_,
    new_B3046_, new_B3047_, new_B3048_, new_B3049_, new_B3050_, new_B3051_,
    new_B3052_, new_B3053_, new_B3054_, new_B3055_, new_B3056_, new_B3057_,
    new_B3058_, new_B3059_, new_B3060_, new_B3061_, new_B3062_, new_B3063_,
    new_B3064_, new_B3065_, new_B3066_, new_B3067_, new_B3068_, new_B3069_,
    new_B3070_, new_B3071_, new_B3072_, new_B3073_, new_B3074_, new_B3075_,
    new_B3076_, new_B3077_, new_B3078_, new_B3079_, new_B3080_, new_B3081_,
    new_B3082_, new_B3083_, new_B3084_, new_B3085_, new_B3086_, new_B3087_,
    new_B3088_, new_B3089_, new_B3090_, new_B3091_, new_B3092_, new_B3093_,
    new_B3094_, new_B3095_, new_B3096_, new_B3097_, new_B3098_, new_B3099_,
    new_B3100_, new_B3101_, new_B3102_, new_B3103_, new_B3104_, new_B3105_,
    new_B3106_, new_B3107_, new_B3108_, new_B3109_, new_B3110_, new_B3111_,
    new_B3112_, new_B3113_, new_B3114_, new_B3115_, new_B3116_, new_B3117_,
    new_B3118_, new_B3119_, new_B3120_, new_B3121_, new_B3122_, new_B3123_,
    new_B3124_, new_B3125_, new_B3126_, new_B3127_, new_B3128_, new_B3129_,
    new_B3130_, new_B3131_, new_B3132_, new_B3133_, new_B3134_, new_B3135_,
    new_B3136_, new_B3137_, new_B3138_, new_B3139_, new_B3140_, new_B3141_,
    new_B3142_, new_B3143_, new_B3144_, new_B3145_, new_B3146_, new_B3147_,
    new_B3148_, new_B3149_, new_B3150_, new_B3151_, new_B3152_, new_B3153_,
    new_B3154_, new_B3155_, new_B3156_, new_B3157_, new_B3158_, new_B3159_,
    new_B3160_, new_B3161_, new_B3162_, new_B3163_, new_B3164_, new_B3165_,
    new_B3166_, new_B3167_, new_B3168_, new_B3169_, new_B3170_, new_B3171_,
    new_B3172_, new_B3173_, new_B3174_, new_B3175_, new_B3176_, new_B3177_,
    new_B3178_, new_B3179_, new_B3180_, new_B3181_, new_B3182_, new_B3183_,
    new_B3184_, new_B3185_, new_B3186_, new_B3187_, new_B3188_, new_B3189_,
    new_B3190_, new_B3191_, new_B3192_, new_B3193_, new_B3194_, new_B3195_,
    new_B3196_, new_B3197_, new_B3198_, new_B3199_, new_B3200_, new_B3201_,
    new_B3202_, new_B3203_, new_B3204_, new_B3205_, new_B3206_, new_B3207_,
    new_B3208_, new_B3209_, new_B3210_, new_B3211_, new_B3212_, new_B3213_,
    new_B3214_, new_B3215_, new_B3216_, new_B3217_, new_B3218_, new_B3219_,
    new_B3220_, new_B3221_, new_B3222_, new_B3223_, new_B3224_, new_B3225_,
    new_B3226_, new_B3227_, new_B3228_, new_B3229_, new_B3230_, new_B3231_,
    new_B3232_, new_B3233_, new_B3234_, new_B3235_, new_B3236_, new_B3237_,
    new_B3238_, new_B3239_, new_B3240_, new_B3241_, new_B3242_, new_B3243_,
    new_B3244_, new_B3245_, new_B3246_, new_B3247_, new_B3248_, new_B3249_,
    new_B3250_, new_B3251_, new_B3252_, new_B3253_, new_B3254_, new_B3255_,
    new_B3256_, new_B3257_, new_B3258_, new_B3259_, new_B3260_, new_B3261_,
    new_B3262_, new_B3263_, new_B3264_, new_B3265_, new_B3266_, new_B3267_,
    new_B3268_, new_B3269_, new_B3270_, new_B3271_, new_B3272_, new_B3273_,
    new_B3274_, new_B3275_, new_B3276_, new_B3277_, new_B3278_, new_B3279_,
    new_B3280_, new_B3281_, new_B3282_, new_B3283_, new_B3284_, new_B3285_,
    new_B3286_, new_B3287_, new_B3288_, new_B3289_, new_B3290_, new_B3291_,
    new_B3292_, new_B3293_, new_B3294_, new_B3295_, new_B3296_, new_B3297_,
    new_B3298_, new_B3299_, new_B3300_, new_B3301_, new_B3302_, new_B3303_,
    new_B3304_, new_B3305_, new_B3306_, new_B3307_, new_B3308_, new_B3309_,
    new_B3310_, new_B3311_, new_B3312_, new_B3313_, new_B3314_, new_B3315_,
    new_B3316_, new_B3317_, new_B3318_, new_B3319_, new_B3320_, new_B3321_,
    new_B3322_, new_B3323_, new_B3324_, new_B3325_, new_B3326_, new_B3327_,
    new_B3328_, new_B3329_, new_B3330_, new_B3331_, new_B3332_, new_B3333_,
    new_B3334_, new_B3335_, new_B3336_, new_B3337_, new_B3338_, new_B3339_,
    new_B3340_, new_B3341_, new_B3342_, new_B3343_, new_B3344_, new_B3345_,
    new_B3346_, new_B3347_, new_B3348_, new_B3349_, new_B3350_, new_B3351_,
    new_B3352_, new_B3353_, new_B3354_, new_B3355_, new_B3356_, new_B3357_,
    new_B3358_, new_B3359_, new_B3360_, new_B3361_, new_B3362_, new_B3363_,
    new_B3364_, new_B3365_, new_B3366_, new_B3367_, new_B3368_, new_B3369_,
    new_B3370_, new_B3371_, new_B3372_, new_B3373_, new_B3374_, new_B3375_,
    new_B3376_, new_B3377_, new_B3378_, new_B3379_, new_B3380_, new_B3381_,
    new_B3382_, new_B3383_, new_B3384_, new_B3385_, new_B3386_, new_B3387_,
    new_B3388_, new_B3389_, new_B3390_, new_B3391_, new_B3392_, new_B3393_,
    new_B3394_, new_B3395_, new_B3396_, new_B3397_, new_B3398_, new_B3399_,
    new_B3400_, new_B3401_, new_B3402_, new_B3403_, new_B3404_, new_B3405_,
    new_B3406_, new_B3407_, new_B3408_, new_B3409_, new_B3410_, new_B3411_,
    new_B3412_, new_B3413_, new_B3414_, new_B3415_, new_B3416_, new_B3417_,
    new_B3418_, new_B3419_, new_B3420_, new_B3421_, new_B3422_, new_B3423_,
    new_B3424_, new_B3425_, new_B3426_, new_B3427_, new_B3428_, new_B3429_,
    new_B3430_, new_B3431_, new_B3432_, new_B3433_, new_B3434_, new_B3435_,
    new_B3436_, new_B3437_, new_B3438_, new_B3439_, new_B3440_, new_B3441_,
    new_B3442_, new_B3443_, new_B3444_, new_B3445_, new_B3446_, new_B3447_,
    new_B3448_, new_B3449_, new_B3450_, new_B3451_, new_B3452_, new_B3453_,
    new_B3454_, new_B3455_, new_B3456_, new_B3457_, new_B3458_, new_B3459_,
    new_B3460_, new_B3461_, new_B3462_, new_B3463_, new_B3464_, new_B3465_,
    new_B3466_, new_B3467_, new_B3468_, new_B3469_, new_B3470_, new_B3471_,
    new_B3472_, new_B3473_, new_B3474_, new_B3475_, new_B3476_, new_B3477_,
    new_B3478_, new_B3479_, new_B3480_, new_B3481_, new_B3482_, new_B3483_,
    new_B3484_, new_B3485_, new_B3486_, new_B3487_, new_B3488_, new_B3489_,
    new_B3490_, new_B3491_, new_B3492_, new_B3493_, new_B3494_, new_B3495_,
    new_B3496_, new_B3497_, new_B3498_, new_B3499_, new_B3500_, new_B3501_,
    new_B3502_, new_B3503_, new_B3504_, new_B3505_, new_B3506_, new_B3507_,
    new_B3508_, new_B3509_, new_B3510_, new_B3511_, new_B3512_, new_B3513_,
    new_B3514_, new_B3515_, new_B3516_, new_B3517_, new_B3518_, new_B3519_,
    new_B3520_, new_B3521_, new_B3522_, new_B3523_, new_B3524_, new_B3525_,
    new_B3526_, new_B3527_, new_B3528_, new_B3529_, new_B3530_, new_B3531_,
    new_B3532_, new_B3533_, new_B3534_, new_B3535_, new_B3536_, new_B3537_,
    new_B3538_, new_B3539_, new_B3540_, new_B3541_, new_B3542_, new_B3543_,
    new_B3544_, new_B3545_, new_B3546_, new_B3547_, new_B3548_, new_B3549_,
    new_B3550_, new_B3551_, new_B3552_, new_B3553_, new_B3554_, new_B3555_,
    new_B3556_, new_B3557_, new_B3558_, new_B3559_, new_B3560_, new_B3561_,
    new_B3562_, new_B3563_, new_B3564_, new_B3565_, new_B3566_, new_B3567_,
    new_B3568_, new_B3569_, new_B3570_, new_B3571_, new_B3572_, new_B3573_,
    new_B3574_, new_B3575_, new_B3576_, new_B3577_, new_B3578_, new_B3579_,
    new_B3580_, new_B3581_, new_B3582_, new_B3583_, new_B3584_, new_B3585_,
    new_B3586_, new_B3587_, new_B3588_, new_B3589_, new_B3590_, new_B3591_,
    new_B3592_, new_B3593_, new_B3594_, new_B3595_, new_B3596_, new_B3597_,
    new_B3598_, new_B3599_, new_B3600_, new_B3601_, new_B3602_, new_B3603_,
    new_B3604_, new_B3605_, new_B3606_, new_B3607_, new_B3608_, new_B3609_,
    new_B3610_, new_B3611_, new_B3612_, new_B3613_, new_B3614_, new_B3615_,
    new_B3616_, new_B3617_, new_B3618_, new_B3619_, new_B3620_, new_B3621_,
    new_B3622_, new_B3623_, new_B3624_, new_B3625_, new_B3626_, new_B3627_,
    new_B3628_, new_B3629_, new_B3630_, new_B3631_, new_B3632_, new_B3633_,
    new_B3634_, new_B3635_, new_B3636_, new_B3637_, new_B3638_, new_B3639_,
    new_B3640_, new_B3641_, new_B3642_, new_B3643_, new_B3644_, new_B3645_,
    new_B3646_, new_B3647_, new_B3648_, new_B3649_, new_B3650_, new_B3651_,
    new_B3652_, new_B3653_, new_B3654_, new_B3655_, new_B3656_, new_B3657_,
    new_B3658_, new_B3659_, new_B3660_, new_B3661_, new_B3662_, new_B3663_,
    new_B3664_, new_B3665_, new_B3666_, new_B3667_, new_B3668_, new_B3669_,
    new_B3670_, new_B3671_, new_B3672_, new_B3673_, new_B3674_, new_B3675_,
    new_B3676_, new_B3677_, new_B3678_, new_B3679_, new_B3680_, new_B3681_,
    new_B3682_, new_B3683_, new_B3684_, new_B3685_, new_B3686_, new_B3687_,
    new_B3688_, new_B3689_, new_B3690_, new_B3691_, new_B3692_, new_B3693_,
    new_B3694_, new_B3695_, new_B3696_, new_B3697_, new_B3698_, new_B3699_,
    new_B3700_, new_B3701_, new_B3702_, new_B3703_, new_B3704_, new_B3705_,
    new_B3706_, new_B3707_, new_B3708_, new_B3709_, new_B3710_, new_B3711_,
    new_B3712_, new_B3713_, new_B3714_, new_B3715_, new_B3716_, new_B3717_,
    new_B3718_, new_B3719_, new_B3720_, new_B3721_, new_B3722_, new_B3723_,
    new_B3724_, new_B3725_, new_B3726_, new_B3727_, new_B3728_, new_B3729_,
    new_B3730_, new_B3731_, new_B3732_, new_B3733_, new_B3734_, new_B3735_,
    new_B3736_, new_B3737_, new_B3738_, new_B3739_, new_B3740_, new_B3741_,
    new_B3742_, new_B3743_, new_B3744_, new_B3745_, new_B3746_, new_B3747_,
    new_B3748_, new_B3749_, new_B3750_, new_B3751_, new_B3752_, new_B3753_,
    new_B3754_, new_B3755_, new_B3756_, new_B3757_, new_B3758_, new_B3759_,
    new_B3760_, new_B3761_, new_B3762_, new_B3763_, new_B3764_, new_B3765_,
    new_B3766_, new_B3767_, new_B3768_, new_B3769_, new_B3770_, new_B3771_,
    new_B3772_, new_B3773_, new_B3774_, new_B3775_, new_B3776_, new_B3777_,
    new_B3778_, new_B3779_, new_B3780_, new_B3781_, new_B3782_, new_B3783_,
    new_B3784_, new_B3785_, new_B3786_, new_B3787_, new_B3788_, new_B3789_,
    new_B3790_, new_B3791_, new_B3792_, new_B3793_, new_B3794_, new_B3795_,
    new_B3796_, new_B3797_, new_B3798_, new_B3799_, new_B3800_, new_B3801_,
    new_B3802_, new_B3803_, new_B3804_, new_B3805_, new_B3806_, new_B3807_,
    new_B3808_, new_B3809_, new_B3810_, new_B3811_, new_B3812_, new_B3813_,
    new_B3814_, new_B3815_, new_B3816_, new_B3817_, new_B3818_, new_B3819_,
    new_B3820_, new_B3821_, new_B3822_, new_B3823_, new_B3824_, new_B3825_,
    new_B3826_, new_B3827_, new_B3828_, new_B3829_, new_B3830_, new_B3831_,
    new_B3832_, new_B3833_, new_B3834_, new_B3835_, new_B3836_, new_B3837_,
    new_B3838_, new_B3839_, new_B3840_, new_B3841_, new_B3842_, new_B3843_,
    new_B3844_, new_B3845_, new_B3846_, new_B3847_, new_B3848_, new_B3849_,
    new_B3850_, new_B3851_, new_B3852_, new_B3853_, new_B3854_, new_B3855_,
    new_B3856_, new_B3857_, new_B3858_, new_B3859_, new_B3860_, new_B3861_,
    new_B3862_, new_B3863_, new_B3864_, new_B3865_, new_B3866_, new_B3867_,
    new_B3868_, new_B3869_, new_B3870_, new_B3871_, new_B3872_, new_B3873_,
    new_B3874_, new_B3875_, new_B3876_, new_B3877_, new_B3878_, new_B3879_,
    new_B3880_, new_B3881_, new_B3882_, new_B3883_, new_B3884_, new_B3885_,
    new_B3886_, new_B3887_, new_B3888_, new_B3889_, new_B3890_, new_B3891_,
    new_B3892_, new_B3893_, new_B3894_, new_B3895_, new_B3896_, new_B3897_,
    new_B3898_, new_B3899_, new_B3900_, new_B3901_, new_B3902_, new_B3903_,
    new_B3904_, new_B3905_, new_B3906_, new_B3907_, new_B3908_, new_B3909_,
    new_B3910_, new_B3911_, new_B3912_, new_B3913_, new_B3914_, new_B3915_,
    new_B3916_, new_B3917_, new_B3918_, new_B3919_, new_B3920_, new_B3921_,
    new_B3922_, new_B3923_, new_B3924_, new_B3925_, new_B3926_, new_B3927_,
    new_B3928_, new_B3929_, new_B3930_, new_B3931_, new_B3932_, new_B3933_,
    new_B3934_, new_B3935_, new_B3936_, new_B3937_, new_B3938_, new_B3939_,
    new_B3940_, new_B3941_, new_B3942_, new_B3943_, new_B3944_, new_B3945_,
    new_B3946_, new_B3947_, new_B3948_, new_B3949_, new_B3950_, new_B3951_,
    new_B3952_, new_B3953_, new_B3954_, new_B3955_, new_B3956_, new_B3957_,
    new_B3958_, new_B3959_, new_B3960_, new_B3961_, new_B3962_, new_B3963_,
    new_B3964_, new_B3965_, new_B3966_, new_B3967_, new_B3968_, new_B3969_,
    new_B3970_, new_B3971_, new_B3972_, new_B3973_, new_B3974_, new_B3975_,
    new_B3976_, new_B3977_, new_B3978_, new_B3979_, new_B3980_, new_B3981_,
    new_B3982_, new_B3983_, new_B3984_, new_B3985_, new_B3986_, new_B3987_,
    new_B3988_, new_B3989_, new_B3990_, new_B3991_, new_B3992_, new_B3993_,
    new_B3994_, new_B3995_, new_B3996_, new_B3997_, new_B3998_, new_B3999_,
    new_B4000_, new_B4001_, new_B4002_, new_B4003_, new_B4004_, new_B4005_,
    new_B4006_, new_B4007_, new_B4008_, new_B4009_, new_B4010_, new_B4011_,
    new_B4012_, new_B4013_, new_B4014_, new_B4015_, new_B4016_, new_B4017_,
    new_B4018_, new_B4019_, new_B4020_, new_B4021_, new_B4022_, new_B4023_,
    new_B4024_, new_B4025_, new_B4026_, new_B4027_, new_B4028_, new_B4029_,
    new_B4030_, new_B4031_, new_B4032_, new_B4033_, new_B4034_, new_B4035_,
    new_B4036_, new_B4037_, new_B4038_, new_B4039_, new_B4040_, new_B4041_,
    new_B4042_, new_B4043_, new_B4044_, new_B4045_, new_B4046_, new_B4047_,
    new_B4048_, new_B4049_, new_B4050_, new_B4051_, new_B4052_, new_B4053_,
    new_B4054_, new_B4055_, new_B4056_, new_B4057_, new_B4058_, new_B4059_,
    new_B4060_, new_B4061_, new_B4062_, new_B4063_, new_B4064_, new_B4065_,
    new_B4066_, new_B4067_, new_B4068_, new_B4069_, new_B4070_, new_B4071_,
    new_B4072_, new_B4073_, new_B4074_, new_B4075_, new_B4076_, new_B4077_,
    new_B4078_, new_B4079_, new_B4080_, new_B4081_, new_B4082_, new_B4083_,
    new_B4084_, new_B4085_, new_B4086_, new_B4087_, new_B4088_, new_B4089_,
    new_B4090_, new_B4091_, new_B4092_, new_B4093_, new_B4094_, new_B4095_,
    new_B4096_, new_B4097_, new_B4098_, new_B4099_, new_B4100_, new_B4101_,
    new_B4102_, new_B4103_, new_B4104_, new_B4105_, new_B4106_, new_B4107_,
    new_B4108_, new_B4109_, new_B4110_, new_B4111_, new_B4112_, new_B4113_,
    new_B4114_, new_B4115_, new_B4116_, new_B4117_, new_B4118_, new_B4119_,
    new_B4120_, new_B4121_, new_B4122_, new_B4123_, new_B4124_, new_B4125_,
    new_B4126_, new_B4127_, new_B4128_, new_B4129_, new_B4130_, new_B4131_,
    new_B4132_, new_B4133_, new_B4134_, new_B4135_, new_B4136_, new_B4137_,
    new_B4138_, new_B4139_, new_B4140_, new_B4141_, new_B4142_, new_B4143_,
    new_B4144_, new_B4145_, new_B4146_, new_B4147_, new_B4148_, new_B4149_,
    new_B4150_, new_B4151_, new_B4152_, new_B4153_, new_B4154_, new_B4155_,
    new_B4156_, new_B4157_, new_B4158_, new_B4159_, new_B4160_, new_B4161_,
    new_B4162_, new_B4163_, new_B4164_, new_B4165_, new_B4166_, new_B4167_,
    new_B4168_, new_B4169_, new_B4170_, new_B4171_, new_B4172_, new_B4173_,
    new_B4174_, new_B4175_, new_B4176_, new_B4177_, new_B4178_, new_B4179_,
    new_B4180_, new_B4181_, new_B4182_, new_B4183_, new_B4184_, new_B4185_,
    new_B4186_, new_B4187_, new_B4188_, new_B4189_, new_B4190_, new_B4191_,
    new_B4192_, new_B4193_, new_B4194_, new_B4195_, new_B4196_, new_B4197_,
    new_B4198_, new_B4199_, new_B4200_, new_B4201_, new_B4202_, new_B4203_,
    new_B4204_, new_B4205_, new_B4206_, new_B4207_, new_B4208_, new_B4209_,
    new_B4210_, new_B4211_, new_B4212_, new_B4213_, new_B4214_, new_B4215_,
    new_B4216_, new_B4217_, new_B4218_, new_B4219_, new_B4220_, new_B4221_,
    new_B4222_, new_B4223_, new_B4224_, new_B4225_, new_B4226_, new_B4227_,
    new_B4228_, new_B4229_, new_B4230_, new_B4231_, new_B4232_, new_B4233_,
    new_B4234_, new_B4235_, new_B4236_, new_B4237_, new_B4238_, new_B4239_,
    new_B4240_, new_B4241_, new_B4242_, new_B4243_, new_B4244_, new_B4245_,
    new_B4246_, new_B4247_, new_B4248_, new_B4249_, new_B4250_, new_B4251_,
    new_B4252_, new_B4253_, new_B4254_, new_B4255_, new_B4256_, new_B4257_,
    new_B4258_, new_B4259_, new_B4260_, new_B4261_, new_B4262_, new_B4263_,
    new_B4264_, new_B4265_, new_B4266_, new_B4267_, new_B4268_, new_B4269_,
    new_B4270_, new_B4271_, new_B4272_, new_B4273_, new_B4274_, new_B4275_,
    new_B4276_, new_B4277_, new_B4278_, new_B4279_, new_B4280_, new_B4281_,
    new_B4282_, new_B4283_, new_B4284_, new_B4285_, new_B4286_, new_B4287_,
    new_B4288_, new_B4289_, new_B4290_, new_B4291_, new_B4292_, new_B4293_,
    new_B4294_, new_B4295_, new_B4296_, new_B4297_, new_B4298_, new_B4299_,
    new_B4300_, new_B4301_, new_B4302_, new_B4303_, new_B4304_, new_B4305_,
    new_B4306_, new_B4307_, new_B4308_, new_B4309_, new_B4310_, new_B4311_,
    new_B4312_, new_B4313_, new_B4314_, new_B4315_, new_B4316_, new_B4317_,
    new_B4318_, new_B4319_, new_B4320_, new_B4321_, new_B4322_, new_B4323_,
    new_B4324_, new_B4325_, new_B4326_, new_B4327_, new_B4328_, new_B4329_,
    new_B4330_, new_B4331_, new_B4332_, new_B4333_, new_B4334_, new_B4335_,
    new_B4336_, new_B4337_, new_B4338_, new_B4339_, new_B4340_, new_B4341_,
    new_B4342_, new_B4343_, new_B4344_, new_B4345_, new_B4346_, new_B4347_,
    new_B4348_, new_B4349_, new_B4350_, new_B4351_, new_B4352_, new_B4353_,
    new_B4354_, new_B4355_, new_B4356_, new_B4357_, new_B4358_, new_B4359_,
    new_B4360_, new_B4361_, new_B4362_, new_B4363_, new_B4364_, new_B4365_,
    new_B4366_, new_B4367_, new_B4368_, new_B4369_, new_B4370_, new_B4371_,
    new_B4372_, new_B4373_, new_B4374_, new_B4375_, new_B4376_, new_B4377_,
    new_B4378_, new_B4379_, new_B4380_, new_B4381_, new_B4382_, new_B4383_,
    new_B4384_, new_B4385_, new_B4386_, new_B4387_, new_B4388_, new_B4389_,
    new_B4390_, new_B4391_, new_B4392_, new_B4393_, new_B4394_, new_B4395_,
    new_B4396_, new_B4397_, new_B4398_, new_B4399_, new_B4400_, new_B4401_,
    new_B4402_, new_B4403_, new_B4404_, new_B4405_, new_B4406_, new_B4407_,
    new_B4408_, new_B4409_, new_B4410_, new_B4411_, new_B4412_, new_B4413_,
    new_B4414_, new_B4415_, new_B4416_, new_B4417_, new_B4418_, new_B4419_,
    new_B4420_, new_B4421_, new_B4422_, new_B4423_, new_B4424_, new_B4425_,
    new_B4426_, new_B4427_, new_B4428_, new_B4429_, new_B4430_, new_B4431_,
    new_B4432_, new_B4433_, new_B4434_, new_B4435_, new_B4436_, new_B4437_,
    new_B4438_, new_B4439_, new_B4440_, new_B4441_, new_B4442_, new_B4443_,
    new_B4444_, new_B4445_, new_B4446_, new_B4447_, new_B4448_, new_B4449_,
    new_B4450_, new_B4451_, new_B4452_, new_B4453_, new_B4454_, new_B4455_,
    new_B4456_, new_B4457_, new_B4458_, new_B4459_, new_B4460_, new_B4461_,
    new_B4462_, new_B4463_, new_B4464_, new_B4465_, new_B4466_, new_B4467_,
    new_B4468_, new_B4469_, new_B4470_, new_B4471_, new_B4472_, new_B4473_,
    new_B4474_, new_B4475_, new_B4476_, new_B4477_, new_B4478_, new_B4479_,
    new_B4480_, new_B4481_, new_B4482_, new_B4483_, new_B4484_, new_B4485_,
    new_B4486_, new_B4487_, new_B4488_, new_B4489_, new_B4490_, new_B4491_,
    new_B4492_, new_B4493_, new_B4494_, new_B4495_, new_B4496_, new_B4497_,
    new_B4498_, new_B4499_, new_B4500_, new_B4501_, new_B4502_, new_B4503_,
    new_B4504_, new_B4505_, new_B4506_, new_B4507_, new_B4508_, new_B4509_,
    new_B4510_, new_B4511_, new_B4512_, new_B4513_, new_B4514_, new_B4515_,
    new_B4516_, new_B4517_, new_B4518_, new_B4519_, new_B4520_, new_B4521_,
    new_B4522_, new_B4523_, new_B4524_, new_B4525_, new_B4526_, new_B4527_,
    new_B4528_, new_B4529_, new_B4530_, new_B4531_, new_B4532_, new_B4533_,
    new_B4534_, new_B4535_, new_B4536_, new_B4537_, new_B4538_, new_B4539_,
    new_B4540_, new_B4541_, new_B4542_, new_B4543_, new_B4544_, new_B4545_,
    new_B4546_, new_B4547_, new_B4548_, new_B4549_, new_B4550_, new_B4551_,
    new_B4552_, new_B4553_, new_B4554_, new_B4555_, new_B4556_, new_B4557_,
    new_B4558_, new_B4559_, new_B4560_, new_B4561_, new_B4562_, new_B4563_,
    new_B4564_, new_B4565_, new_B4566_, new_B4567_, new_B4568_, new_B4569_,
    new_B4570_, new_B4571_, new_B4572_, new_B4573_, new_B4574_, new_B4575_,
    new_B4576_, new_B4577_, new_B4578_, new_B4579_, new_B4580_, new_B4581_,
    new_B4582_, new_B4583_, new_B4584_, new_B4585_, new_B4586_, new_B4587_,
    new_B4588_, new_B4589_, new_B4590_, new_B4591_, new_B4592_, new_B4593_,
    new_B4594_, new_B4595_, new_B4596_, new_B4597_, new_B4598_, new_B4599_,
    new_B4600_, new_B4601_, new_B4602_, new_B4603_, new_B4604_, new_B4605_,
    new_B4606_, new_B4607_, new_B4608_, new_B4609_, new_B4610_, new_B4611_,
    new_B4612_, new_B4613_, new_B4614_, new_B4615_, new_B4616_, new_B4617_,
    new_B4618_, new_B4619_, new_B4620_, new_B4621_, new_B4622_, new_B4623_,
    new_B4624_, new_B4625_, new_B4626_, new_B4627_, new_B4628_, new_B4629_,
    new_B4630_, new_B4631_, new_B4632_, new_B4633_, new_B4634_, new_B4635_,
    new_B4636_, new_B4637_, new_B4638_, new_B4639_, new_B4640_, new_B4641_,
    new_B4642_, new_B4643_, new_B4644_, new_B4645_, new_B4646_, new_B4647_,
    new_B4648_, new_B4649_, new_B4650_, new_B4651_, new_B4652_, new_B4653_,
    new_B4654_, new_B4655_, new_B4656_, new_B4657_, new_B4658_, new_B4659_,
    new_B4660_, new_B4661_, new_B4662_, new_B4663_, new_B4664_, new_B4665_,
    new_B4666_, new_B4667_, new_B4668_, new_B4669_, new_B4670_, new_B4671_,
    new_B4672_, new_B4673_, new_B4674_, new_B4675_, new_B4676_, new_B4677_,
    new_B4678_, new_B4679_, new_B4680_, new_B4681_, new_B4682_, new_B4683_,
    new_B4684_, new_B4685_, new_B4686_, new_B4687_, new_B4688_, new_B4689_,
    new_B4690_, new_B4691_, new_B4692_, new_B4693_, new_B4694_, new_B4695_,
    new_B4696_, new_B4697_, new_B4698_, new_B4699_, new_B4700_, new_B4701_,
    new_B4702_, new_B4703_, new_B4704_, new_B4705_, new_B4706_, new_B4707_,
    new_B4708_, new_B4709_, new_B4710_, new_B4711_, new_B4712_, new_B4713_,
    new_B4714_, new_B4715_, new_B4716_, new_B4717_, new_B4718_, new_B4719_,
    new_B4720_, new_B4721_, new_B4722_, new_B4723_, new_B4724_, new_B4725_,
    new_B4726_, new_B4727_, new_B4728_, new_B4729_, new_B4730_, new_B4731_,
    new_B4732_, new_B4733_, new_B4734_, new_B4735_, new_B4736_, new_B4737_,
    new_B4738_, new_B4739_, new_B4740_, new_B4741_, new_B4742_, new_B4743_,
    new_B4744_, new_B4745_, new_B4746_, new_B4747_, new_B4748_, new_B4749_,
    new_B4750_, new_B4751_, new_B4752_, new_B4753_, new_B4754_, new_B4755_,
    new_B4756_, new_B4757_, new_B4758_, new_B4759_, new_B4760_, new_B4761_,
    new_B4762_, new_B4763_, new_B4764_, new_B4765_, new_B4766_, new_B4767_,
    new_B4768_, new_B4769_, new_B4770_, new_B4771_, new_B4772_, new_B4773_,
    new_B4774_, new_B4775_, new_B4776_, new_B4777_, new_B4778_, new_B4779_,
    new_B4780_, new_B4781_, new_B4782_, new_B4783_, new_B4784_, new_B4785_,
    new_B4786_, new_B4787_, new_B4788_, new_B4789_, new_B4790_, new_B4791_,
    new_B4792_, new_B4793_, new_B4794_, new_B4795_, new_B4796_, new_B4797_,
    new_B4798_, new_B4799_, new_B4800_, new_B4801_, new_B4802_, new_B4803_,
    new_B4804_, new_B4805_, new_B4806_, new_B4807_, new_B4808_, new_B4809_,
    new_B4810_, new_B4811_, new_B4812_, new_B4813_, new_B4814_, new_B4815_,
    new_B4816_, new_B4817_, new_B4818_, new_B4819_, new_B4820_, new_B4821_,
    new_B4822_, new_B4823_, new_B4824_, new_B4825_, new_B4826_, new_B4827_,
    new_B4828_, new_B4829_, new_B4830_, new_B4831_, new_B4832_, new_B4833_,
    new_B4834_, new_B4835_, new_B4836_, new_B4837_, new_B4838_, new_B4839_,
    new_B4840_, new_B4841_, new_B4842_, new_B4843_, new_B4844_, new_B4845_,
    new_B4846_, new_B4847_, new_B4848_, new_B4849_, new_B4850_, new_B4851_,
    new_B4852_, new_B4853_, new_B4854_, new_B4855_, new_B4856_, new_B4857_,
    new_B4858_, new_B4859_, new_B4860_, new_B4861_, new_B4862_, new_B4863_,
    new_B4864_, new_B4865_, new_B4866_, new_B4867_, new_B4868_, new_B4869_,
    new_B4870_, new_B4871_, new_B4872_, new_B4873_, new_B4874_, new_B4875_,
    new_B4876_, new_B4877_, new_B4878_, new_B4879_, new_B4880_, new_B4881_,
    new_B4882_, new_B4883_, new_B4884_, new_B4885_, new_B4886_, new_B4887_,
    new_B4888_, new_B4889_, new_B4890_, new_B4891_, new_B4892_, new_B4893_,
    new_B4894_, new_B4895_, new_B4896_, new_B4897_, new_B4898_, new_B4899_,
    new_B4900_, new_B4901_, new_B4902_, new_B4903_, new_B4904_, new_B4905_,
    new_B4906_, new_B4907_, new_B4908_, new_B4909_, new_B4910_, new_B4911_,
    new_B4912_, new_B4913_, new_B4914_, new_B4915_, new_B4916_, new_B4917_,
    new_B4918_, new_B4919_, new_B4920_, new_B4921_, new_B4922_, new_B4923_,
    new_B4924_, new_B4925_, new_B4926_, new_B4927_, new_B4928_, new_B4929_,
    new_B4930_, new_B4931_, new_B4932_, new_B4933_, new_B4934_, new_B4935_,
    new_B4936_, new_B4937_, new_B4938_, new_B4939_, new_B4940_, new_B4941_,
    new_B4942_, new_B4943_, new_B4944_, new_B4945_, new_B4946_, new_B4947_,
    new_B4948_, new_B4949_, new_B4950_, new_B4951_, new_B4952_, new_B4953_,
    new_B4954_, new_B4955_, new_B4956_, new_B4957_, new_B4958_, new_B4959_,
    new_B4960_, new_B4961_, new_B4962_, new_B4963_, new_B4964_, new_B4965_,
    new_B4966_, new_B4967_, new_B4968_, new_B4969_, new_B4970_, new_B4971_,
    new_B4972_, new_B4973_, new_B4974_, new_B4975_, new_B4976_, new_B4977_,
    new_B4978_, new_B4979_, new_B4980_, new_B4981_, new_B4982_, new_B4983_,
    new_B4984_, new_B4985_, new_B4986_, new_B4987_, new_B4988_, new_B4989_,
    new_B4990_, new_B4991_, new_B4992_, new_B4993_, new_B4994_, new_B4995_,
    new_B4996_, new_B4997_, new_B4998_, new_B4999_, new_B5000_, new_B5001_,
    new_B5002_, new_B5003_, new_B5004_, new_B5005_, new_B5006_, new_B5007_,
    new_B5008_, new_B5009_, new_B5010_, new_B5011_, new_B5012_, new_B5013_,
    new_B5014_, new_B5015_, new_B5016_, new_B5017_, new_B5018_, new_B5019_,
    new_B5020_, new_B5021_, new_B5022_, new_B5023_, new_B5024_, new_B5025_,
    new_B5026_, new_B5027_, new_B5028_, new_B5029_, new_B5030_, new_B5031_,
    new_B5032_, new_B5033_, new_B5034_, new_B5035_, new_B5036_, new_B5037_,
    new_B5038_, new_B5039_, new_B5040_, new_B5041_, new_B5042_, new_B5043_,
    new_B5044_, new_B5045_, new_B5046_, new_B5047_, new_B5048_, new_B5049_,
    new_B5050_, new_B5051_, new_B5052_, new_B5053_, new_B5054_, new_B5055_,
    new_B5056_, new_B5057_, new_B5058_, new_B5059_, new_B5060_, new_B5061_,
    new_B5062_, new_B5063_, new_B5064_, new_B5065_, new_B5066_, new_B5067_,
    new_B5068_, new_B5069_, new_B5070_, new_B5071_, new_B5072_, new_B5073_,
    new_B5074_, new_B5075_, new_B5076_, new_B5077_, new_B5078_, new_B5079_,
    new_B5080_, new_B5081_, new_B5082_, new_B5083_, new_B5084_, new_B5085_,
    new_B5086_, new_B5087_, new_B5088_, new_B5089_, new_B5090_, new_B5091_,
    new_B5092_, new_B5093_, new_B5094_, new_B5095_, new_B5096_, new_B5097_,
    new_B5098_, new_B5099_, new_B5100_, new_B5101_, new_B5102_, new_B5103_,
    new_B5104_, new_B5105_, new_B5106_, new_B5107_, new_B5108_, new_B5109_,
    new_B5110_, new_B5111_, new_B5112_, new_B5113_, new_B5114_, new_B5115_,
    new_B5116_, new_B5117_, new_B5118_, new_B5119_, new_B5120_, new_B5121_,
    new_B5122_, new_B5123_, new_B5124_, new_B5125_, new_B5126_, new_B5127_,
    new_B5128_, new_B5129_, new_B5130_, new_B5131_, new_B5132_, new_B5133_,
    new_B5134_, new_B5135_, new_B5136_, new_B5137_, new_B5138_, new_B5139_,
    new_B5140_, new_B5141_, new_B5142_, new_B5143_, new_B5144_, new_B5145_,
    new_B5146_, new_B5147_, new_B5148_, new_B5149_, new_B5150_, new_B5151_,
    new_B5152_, new_B5153_, new_B5154_, new_B5155_, new_B5156_, new_B5157_,
    new_B5158_, new_B5159_, new_B5160_, new_B5161_, new_B5162_, new_B5163_,
    new_B5164_, new_B5165_, new_B5166_, new_B5167_, new_B5168_, new_B5169_,
    new_B5170_, new_B5171_, new_B5172_, new_B5173_, new_B5174_, new_B5175_,
    new_B5176_, new_B5177_, new_B5178_, new_B5179_, new_B5180_, new_B5181_,
    new_A6963_, new_A6962_, new_A6961_, new_A6960_, new_A6959_, new_A6958_,
    new_A6957_, new_A6956_, new_A6955_, new_A6954_, new_A6953_, new_A6952_,
    new_A6951_, new_A6950_, new_A6949_, new_A6948_, new_A6947_, new_A6946_,
    new_A6945_, new_A6944_, new_A6943_, new_A6942_, new_A6941_, new_A6940_,
    new_A6939_, new_A6938_, new_A6937_, new_A6936_, new_A6935_, new_A6934_,
    new_A6933_, new_A6932_, new_A6931_, new_A6964_, new_A6965_, new_A6966_,
    new_A6967_, new_A6968_, new_A6969_, new_A6970_, new_A6971_, new_A6972_,
    new_A6973_, new_A6974_, new_A6975_, new_A6976_, new_A6977_, new_A6978_,
    new_A6979_, new_A6980_, new_A6981_, new_A6982_, new_A6983_, new_A6984_,
    new_A6985_, new_A6986_, new_A6987_, new_A6988_, new_A6989_, new_A6990_,
    new_A6991_, new_A6992_, new_A6993_, new_A6994_, new_A6995_, new_A6996_,
    new_A6997_, new_A6998_, new_A6999_, new_A7000_, new_A7001_, new_A7002_,
    new_A7003_, new_A7004_, new_A7005_, new_A7006_, new_A7007_, new_A7008_,
    new_A7009_, new_A7010_, new_A7011_, new_A7012_, new_A7013_, new_A7014_,
    new_A7015_, new_A7016_, new_A7017_, new_A7018_, new_A7019_, new_A7020_,
    new_A7021_, new_A7022_, new_A7023_, new_A7024_, new_A7025_, new_A7026_,
    new_A7027_, new_A7028_, new_A7029_, new_A7030_, new_A7031_, new_A7032_,
    new_A7033_, new_A7034_, new_A7035_, new_A7036_, new_A7037_, new_A7038_,
    new_A7039_, new_A7040_, new_A7041_, new_A7042_, new_A7043_, new_A7044_,
    new_A7045_, new_A7046_, new_A7047_, new_A7048_, new_A7049_, new_A7050_,
    new_A7051_, new_A7052_, new_A7053_, new_A7054_, new_A7055_, new_A7056_,
    new_A7057_, new_A7058_, new_A7059_, new_A7060_, new_A7061_, new_A7062_,
    new_A7063_, new_A7064_, new_A7065_, new_A7066_, new_A7067_, new_A7068_,
    new_A7069_, new_A7070_, new_A7071_, new_A7072_, new_A7073_, new_A7074_,
    new_A7075_, new_A7076_, new_A7077_, new_A7078_, new_A7079_, new_A7080_,
    new_A7081_, new_A7082_, new_A7083_, new_A7084_, new_A7085_, new_A7086_,
    new_A7087_, new_A7088_, new_A7089_, new_A7090_, new_A7091_, new_A7092_,
    new_A7093_, new_A7094_, new_A7095_, new_A7096_, new_A7097_, new_A7098_,
    new_A7099_, new_A7100_, new_A7101_, new_A7102_, new_A7103_, new_A7104_,
    new_A7105_, new_A7106_, new_A7107_, new_A7108_, new_A7109_, new_A7110_,
    new_A7111_, new_A7112_, new_A7113_, new_A7114_, new_A7115_, new_A7116_,
    new_A7117_, new_A7118_, new_A7119_, new_A7120_, new_A7121_, new_A7122_,
    new_A7123_, new_A7124_, new_A7125_, new_A7126_, new_A7127_, new_A7128_,
    new_A7129_, new_A7130_, new_A7131_, new_A7132_, new_A7133_, new_A7134_,
    new_A7135_, new_A7136_, new_A7137_, new_A7138_, new_A7139_, new_A7140_,
    new_A7141_, new_A7142_, new_A7143_, new_A7144_, new_A7145_, new_A7146_,
    new_A7147_, new_A7148_, new_A7149_, new_A7150_, new_A7151_, new_A7152_,
    new_A7153_, new_A7154_, new_A7155_, new_A7156_, new_A7157_, new_A7158_,
    new_A7159_, new_A7160_, new_A7161_, new_A7162_, new_A7163_, new_A7164_,
    new_A7165_, new_A7166_, new_A7167_, new_A7168_, new_A7169_, new_A7170_,
    new_A7171_, new_A7172_, new_A7173_, new_A7174_, new_A7175_, new_A7176_,
    new_A7177_, new_A7178_, new_A7179_, new_A7180_, new_A7181_, new_A7182_,
    new_A7183_, new_A7184_, new_A7185_, new_A7186_, new_A7187_, new_A7188_,
    new_A7189_, new_A7190_, new_A7191_, new_A7192_, new_A7193_, new_A7194_,
    new_A7195_, new_A7196_, new_A7197_, new_A7198_, new_A7199_, new_A7200_,
    new_A7201_, new_A7202_, new_A7203_, new_A7204_, new_A7205_, new_A7206_,
    new_A7207_, new_A7208_, new_A7209_, new_A7210_, new_A7211_, new_A7212_,
    new_A7213_, new_A7214_, new_A7215_, new_A7216_, new_A7217_, new_A7218_,
    new_A7219_, new_A7220_, new_A7221_, new_A7222_, new_A7223_, new_A7224_,
    new_A7225_, new_A7226_, new_A7227_, new_A7228_, new_A7229_, new_A7230_,
    new_A7231_, new_A7232_, new_A7233_, new_A7234_, new_A7235_, new_A7236_,
    new_A7237_, new_A7238_, new_A7239_, new_A7240_, new_A7241_, new_A7242_,
    new_A7243_, new_A7244_, new_A7245_, new_A7246_, new_A7247_, new_A7248_,
    new_A7249_, new_A7250_, new_A7251_, new_A7252_, new_A7253_, new_A7254_,
    new_A7255_, new_A7256_, new_A7257_, new_A7258_, new_A7259_, new_A7260_,
    new_A7261_, new_A7262_, new_A7263_, new_A7264_, new_A7265_, new_A7266_,
    new_A7267_, new_A7268_, new_A7269_, new_A7270_, new_A7271_, new_A7272_,
    new_A7273_, new_A7274_, new_A7275_, new_A7276_, new_A7277_, new_A7278_,
    new_A7279_, new_A7280_, new_A7281_, new_A7282_, new_A7283_, new_A7284_,
    new_A7285_, new_A7286_, new_A7287_, new_A7288_, new_A7289_, new_A7290_,
    new_A7291_, new_A7292_, new_A7293_, new_A7294_, new_A7295_, new_A7296_,
    new_A7297_, new_A7298_, new_A7299_, new_A7300_, new_A7301_, new_A7302_,
    new_A7303_, new_A7304_, new_A7305_, new_A7306_, new_A7307_, new_A7308_,
    new_A7309_, new_A7310_, new_A7311_, new_A7312_, new_A7313_, new_A7314_,
    new_A7315_, new_A7316_, new_A7317_, new_A7318_, new_A7319_, new_A7320_,
    new_A7321_, new_A7322_, new_A7323_, new_A7324_, new_A7325_, new_A7326_,
    new_A7327_, new_A7328_, new_A7329_, new_A7330_, new_A7331_, new_A7332_,
    new_A7333_, new_A7334_, new_A7335_, new_A7336_, new_A7337_, new_A7338_,
    new_A7339_, new_A7340_, new_A7341_, new_A7342_, new_A7343_, new_A7344_,
    new_A7345_, new_A7346_, new_A7347_, new_A7348_, new_A7349_, new_A7350_,
    new_A7351_, new_A7352_, new_A7353_, new_A7354_, new_A7355_, new_A7356_,
    new_A7357_, new_A7358_, new_A7359_, new_A7360_, new_A7361_, new_A7362_,
    new_A7363_, new_A7364_, new_A7365_, new_A7366_, new_A7367_, new_A7368_,
    new_A7369_, new_A7370_, new_A7371_, new_A7372_, new_A7373_, new_A7374_,
    new_A7375_, new_A7376_, new_A7377_, new_A7378_, new_A7379_, new_A7380_,
    new_A7381_, new_A7382_, new_A7383_, new_A7384_, new_A7385_, new_A7386_,
    new_A7387_, new_A7388_, new_A7389_, new_A7390_, new_A7391_, new_A7392_,
    new_A7393_, new_A7394_, new_A7395_, new_A7396_, new_A7397_, new_A7398_,
    new_A7399_, new_A7400_, new_A7401_, new_A7402_, new_A7403_, new_A7404_,
    new_A7405_, new_A7406_, new_A7407_, new_A7408_, new_A7409_, new_A7410_,
    new_A7411_, new_A7412_, new_A7413_, new_A7414_, new_A7415_, new_A7416_,
    new_A7417_, new_A7418_, new_A7419_, new_A7420_, new_A7421_, new_A7422_,
    new_A7423_, new_A7424_, new_A7425_, new_A7426_, new_A7427_, new_A7428_,
    new_A7429_, new_A7430_, new_A7431_, new_A7432_, new_A7433_, new_A7434_,
    new_A7435_, new_A7436_, new_A7437_, new_A7438_, new_A7439_, new_A7440_,
    new_A7441_, new_A7442_, new_A7443_, new_A7444_, new_A7445_, new_A7446_,
    new_A7447_, new_A7448_, new_A7449_, new_A7450_, new_A7451_, new_A7452_,
    new_A7453_, new_A7454_, new_A7455_, new_A7456_, new_A7457_, new_A7458_,
    new_A7459_, new_A7460_, new_A7461_, new_A7462_, new_A7463_, new_A7464_,
    new_A7465_, new_A7466_, new_A7467_, new_A7468_, new_A7469_, new_A7470_,
    new_A7471_, new_A7472_, new_A7473_, new_A7474_, new_A7475_, new_A7476_,
    new_A7477_, new_A7478_, new_A7479_, new_A7480_, new_A7481_, new_A7482_,
    new_A7483_, new_A7484_, new_A7485_, new_A7486_, new_A7487_, new_A7488_,
    new_A7489_, new_A7490_, new_A7491_, new_A7492_, new_A7493_, new_A7494_,
    new_A7495_, new_A7496_, new_A7497_, new_A7498_, new_A7499_, new_A7500_,
    new_A7501_, new_A7502_, new_A7503_, new_A7504_, new_A7505_, new_A7506_,
    new_A7507_, new_A7508_, new_A7509_, new_A7510_, new_A7511_, new_A7512_,
    new_A7513_, new_A7514_, new_A7515_, new_A7516_, new_A7517_, new_A7518_,
    new_A7519_, new_A7520_, new_A7521_, new_A7522_, new_A7523_, new_A7524_,
    new_A7525_, new_A7526_, new_A7527_, new_A7528_, new_A7529_, new_A7530_,
    new_A7531_, new_A7532_, new_A7533_, new_A7534_, new_A7535_, new_A7536_,
    new_A7537_, new_A7538_, new_A7539_, new_A7540_, new_A7541_, new_A7542_,
    new_A7543_, new_A7544_, new_A7545_, new_A7546_, new_A7547_, new_A7548_,
    new_A7549_, new_A7550_, new_A7551_, new_A7552_, new_A7553_, new_A7554_,
    new_A7555_, new_A7556_, new_A7557_, new_A7558_, new_A7559_, new_A7560_,
    new_A7561_, new_A7562_, new_A7563_, new_A7564_, new_A7565_, new_A7566_,
    new_A7567_, new_A7568_, new_A7569_, new_A7570_, new_A7571_, new_A7572_,
    new_A7573_, new_A7574_, new_A7575_, new_A7576_, new_A7577_, new_A7578_,
    new_A7579_, new_A7580_, new_A7581_, new_A7582_, new_A7583_, new_A7584_,
    new_A7585_, new_A7586_, new_A7587_, new_A7588_, new_A7589_, new_A7590_,
    new_A7591_, new_A7592_, new_A7593_, new_A7594_, new_A7595_, new_A7596_,
    new_A7597_, new_A7598_, new_A7599_, new_A7600_, new_A7601_, new_A7602_,
    new_A7603_, new_A7604_, new_A7605_, new_A7606_, new_A7607_, new_A7608_,
    new_A7609_, new_A7610_, new_A7611_, new_A7612_, new_A7613_, new_A7614_,
    new_A7615_, new_A7616_, new_A7617_, new_A7618_, new_A7619_, new_A7620_,
    new_A7621_, new_A7622_, new_A7623_, new_A7624_, new_A7625_, new_A7626_,
    new_A7627_, new_A7628_, new_A7629_, new_A7630_, new_A7631_, new_A7632_,
    new_A7633_, new_A7634_, new_A7635_, new_A7636_, new_A7637_, new_A7638_,
    new_A7639_, new_A7640_, new_A7641_, new_A7642_, new_A7643_, new_A7644_,
    new_A7645_, new_A7646_, new_A7647_, new_A7648_, new_A7649_, new_A7650_,
    new_A7651_, new_A7652_, new_A7653_, new_A7654_, new_A7655_, new_A7656_,
    new_A7657_, new_A7658_, new_A7659_, new_A7660_, new_A7661_, new_A7662_,
    new_A7663_, new_A7664_, new_A7665_, new_A7666_, new_A7667_, new_A7668_,
    new_A7669_, new_A7670_, new_A7671_, new_A7672_, new_A7673_, new_A7674_,
    new_A7675_, new_A7676_, new_A7677_, new_A7678_, new_A7679_, new_A7680_,
    new_A7681_, new_A7682_, new_A7683_, new_A7684_, new_A7685_, new_A7686_,
    new_A7687_, new_A7688_, new_A7689_, new_A7690_, new_A7691_, new_A7692_,
    new_A7693_, new_A7694_, new_A7695_, new_A7696_, new_A7697_, new_A7698_,
    new_A7699_, new_A7700_, new_A7701_, new_A7702_, new_A7703_, new_A7704_,
    new_A7705_, new_A7706_, new_A7707_, new_A7708_, new_A7709_, new_A7710_,
    new_A7711_, new_A7712_, new_A7713_, new_A7714_, new_A7715_, new_A7716_,
    new_A7717_, new_A7718_, new_A7719_, new_A7720_, new_A7721_, new_A7722_,
    new_A7723_, new_A7724_, new_A7725_, new_A7726_, new_A7727_, new_A7728_,
    new_A7729_, new_A7730_, new_A7731_, new_A7732_, new_A7733_, new_A7734_,
    new_A7735_, new_A7736_, new_A7737_, new_A7738_, new_A7739_, new_A7740_,
    new_A7741_, new_A7742_, new_A7743_, new_A7744_, new_A7745_, new_A7746_,
    new_A7747_, new_A7748_, new_A7749_, new_A7750_, new_A7751_, new_A7752_,
    new_A7753_, new_A7754_, new_A7755_, new_A7756_, new_A7757_, new_A7758_,
    new_A7759_, new_A7760_, new_A7761_, new_A7762_, new_A7763_, new_A7764_,
    new_A7765_, new_A7766_, new_A7767_, new_A7768_, new_A7769_, new_A7770_,
    new_A7771_, new_A7772_, new_A7773_, new_A7774_, new_A7775_, new_A7776_,
    new_A7777_, new_A7778_, new_A7779_, new_A7780_, new_A7781_, new_A7782_,
    new_A7783_, new_A7784_, new_A7785_, new_A7786_, new_A7787_, new_A7788_,
    new_A7789_, new_A7790_, new_A7791_, new_A7792_, new_A7793_, new_A7794_,
    new_A7795_, new_A7796_, new_A7797_, new_A7798_, new_A7799_, new_A7800_,
    new_A7801_, new_A7802_, new_A7803_, new_A7804_, new_A7805_, new_A7806_,
    new_A7807_, new_A7808_, new_A7809_, new_A7810_, new_A7811_, new_A7812_,
    new_A7813_, new_A7814_, new_A7815_, new_A7816_, new_A7817_, new_A7818_,
    new_A7819_, new_A7820_, new_A7821_, new_A7822_, new_A7823_, new_A7824_,
    new_A7825_, new_A7826_, new_A7827_, new_A7828_, new_A7829_, new_A7830_,
    new_A7831_, new_A7832_, new_A7833_, new_A7834_, new_A7835_, new_A7836_,
    new_A7837_, new_A7838_, new_A7839_, new_A7840_, new_A7841_, new_A7842_,
    new_A7843_, new_A7844_, new_A7845_, new_A7846_, new_A7847_, new_A7848_,
    new_A7849_, new_A7850_, new_A7851_, new_A7852_, new_A7853_, new_A7854_,
    new_A7855_, new_A7856_, new_A7857_, new_A7858_, new_A7859_, new_A7860_,
    new_A7861_, new_A7862_, new_A7863_, new_A7864_, new_A7865_, new_A7866_,
    new_A7867_, new_A7868_, new_A7869_, new_A7870_, new_A7871_, new_A7872_,
    new_A7873_, new_A7874_, new_A7875_, new_A7876_, new_A7877_, new_A7878_,
    new_A7879_, new_A7880_, new_A7881_, new_A7882_, new_A7883_, new_A7884_,
    new_A7885_, new_A7886_, new_A7887_, new_A7888_, new_A7889_, new_A7890_,
    new_A7891_, new_A7892_, new_A7893_, new_A7894_, new_A7895_, new_A7896_,
    new_A7897_, new_A7898_, new_A7899_, new_A7900_, new_A7901_, new_A7902_,
    new_A7903_, new_A7904_, new_A7905_, new_A7906_, new_A7907_, new_A7908_,
    new_A7909_, new_A7910_, new_A7911_, new_A7912_, new_A7913_, new_A7914_,
    new_A7915_, new_A7916_, new_A7917_, new_A7918_, new_A7919_, new_A7920_,
    new_A7921_, new_A7922_, new_A7923_, new_A7924_, new_A7925_, new_A7926_,
    new_A7927_, new_A7928_, new_A7929_, new_A7930_, new_A7931_, new_A7932_,
    new_A7933_, new_A7934_, new_A7935_, new_A7936_, new_A7937_, new_A7938_,
    new_A7939_, new_A7940_, new_A7941_, new_A7942_, new_A7943_, new_A7944_,
    new_A7945_, new_A7946_, new_A7947_, new_A7948_, new_A7949_, new_A7950_,
    new_A7951_, new_A7952_, new_A7953_, new_A7954_, new_A7955_, new_A7956_,
    new_A7957_, new_A7958_, new_A7959_, new_A7960_, new_A7961_, new_A7962_,
    new_A7963_, new_A7964_, new_A7965_, new_A7966_, new_A7967_, new_A7968_,
    new_A7969_, new_A7970_, new_A7971_, new_A7972_, new_A7973_, new_A7974_,
    new_A7975_, new_A7976_, new_A7977_, new_A7978_, new_A7979_, new_A7980_,
    new_A7981_, new_A7982_, new_A7983_, new_A7984_, new_A7985_, new_A7986_,
    new_A7987_, new_A7988_, new_A7989_, new_A7990_, new_A7991_, new_A7992_,
    new_A7993_, new_A7994_, new_A7995_, new_A7996_, new_A7997_, new_A7998_,
    new_A7999_, new_A8000_, new_A8001_, new_A8002_, new_A8003_, new_A8004_,
    new_A8005_, new_A8006_, new_A8007_, new_A8008_, new_A8009_, new_A8010_,
    new_A8011_, new_A8012_, new_A8013_, new_A8014_, new_A8015_, new_A8016_,
    new_A8017_, new_A8018_, new_A8019_, new_A8020_, new_A8021_, new_A8022_,
    new_A8023_, new_A8024_, new_A8025_, new_A8026_, new_A8027_, new_A8028_,
    new_A8029_, new_A8030_, new_A8031_, new_A8032_, new_A8033_, new_A8034_,
    new_A8035_, new_A8036_, new_A8037_, new_A8038_, new_A8039_, new_A8040_,
    new_A8041_, new_A8042_, new_A8043_, new_A8044_, new_A8045_, new_A8046_,
    new_A8047_, new_A8048_, new_A8049_, new_A8050_, new_A8051_, new_A8052_,
    new_A8053_, new_A8054_, new_A8055_, new_A8056_, new_A8057_, new_A8058_,
    new_A8059_, new_A8060_, new_A8061_, new_A8062_, new_A8063_, new_A8064_,
    new_A8065_, new_A8066_, new_A8067_, new_A8068_, new_A8069_, new_A8070_,
    new_A8071_, new_A8072_, new_A8073_, new_A8074_, new_A8075_, new_A8076_,
    new_A8077_, new_A8078_, new_A8079_, new_A8080_, new_A8081_, new_A8082_,
    new_A8083_, new_A8084_, new_A8085_, new_A8086_, new_A8087_, new_A8088_,
    new_A8089_, new_A8090_, new_A8091_, new_A8092_, new_A8093_, new_A8094_,
    new_A8095_, new_A8096_, new_A8097_, new_A8098_, new_A8099_, new_A8100_,
    new_A8101_, new_A8102_, new_A8103_, new_A8104_, new_A8105_, new_A8106_,
    new_A8107_, new_A8108_, new_A8109_, new_A8110_, new_A8111_, new_A8112_,
    new_A8113_, new_A8114_, new_A8115_, new_A8116_, new_A8117_, new_A8118_,
    new_A8119_, new_A8120_, new_A8121_, new_A8122_, new_A8123_, new_A8124_,
    new_A8125_, new_A8126_, new_A8127_, new_A8128_, new_A8129_, new_A8130_,
    new_A8131_, new_A8132_, new_A8133_, new_A8134_, new_A8135_, new_A8136_,
    new_A8137_, new_A8138_, new_A8139_, new_A8140_, new_A8141_, new_A8142_,
    new_A8143_, new_A8144_, new_A8145_, new_A8146_, new_A8147_, new_A8148_,
    new_A8149_, new_A8150_, new_A8151_, new_A8152_, new_A8153_, new_A8154_,
    new_A8155_, new_A8156_, new_A8157_, new_A8158_, new_A8159_, new_A8160_,
    new_A8161_, new_A8162_, new_A8163_, new_A8164_, new_A8165_, new_A8166_,
    new_A8167_, new_A8168_, new_A8169_, new_A8170_, new_A8171_, new_A8172_,
    new_A8173_, new_A8174_, new_A8175_, new_A8176_, new_A8177_, new_A8178_,
    new_A8179_, new_A8180_, new_A8181_, new_A8182_, new_A8183_, new_A8184_,
    new_A8185_, new_A8186_, new_A8187_, new_A8188_, new_A8189_, new_A8190_,
    new_A8191_, new_A8192_, new_A8193_, new_A8194_, new_A8195_, new_A8196_,
    new_A8197_, new_A8198_, new_A8199_, new_A8200_, new_A8201_, new_A8202_,
    new_A8203_, new_A8204_, new_A8205_, new_A8206_, new_A8207_, new_A8208_,
    new_A8209_, new_A8210_, new_A8211_, new_A8212_, new_A8213_, new_A8214_,
    new_A8215_, new_A8216_, new_A8217_, new_A8218_, new_A8219_, new_A8220_,
    new_A8221_, new_A8222_, new_A8223_, new_A8224_, new_A8225_, new_A8226_,
    new_A8227_, new_A8228_, new_A8229_, new_A8230_, new_A8231_, new_A8232_,
    new_A8233_, new_A8234_, new_A8235_, new_A8236_, new_A8237_, new_A8238_,
    new_A8239_, new_A8240_, new_A8241_, new_A8242_, new_A8243_, new_A8244_,
    new_A8245_, new_A8246_, new_A8247_, new_A8248_, new_A8249_, new_A8250_,
    new_A8251_, new_A8252_, new_A8253_, new_A8254_, new_A8255_, new_A8256_,
    new_A8257_, new_A8258_, new_A8259_, new_A8260_, new_A8261_, new_A8262_,
    new_A8263_, new_A8264_, new_A8265_, new_A8266_, new_A8267_, new_A8268_,
    new_A8269_, new_A8270_, new_A8271_, new_A8272_, new_A8273_, new_A8274_,
    new_A8275_, new_A8276_, new_A8277_, new_A8278_, new_A8279_, new_A8280_,
    new_A8281_, new_A8282_, new_A8283_, new_A8284_, new_A8285_, new_A8286_,
    new_A8287_, new_A8288_, new_A8289_, new_A8290_, new_A8291_, new_A8292_,
    new_A8293_, new_A8294_, new_A8295_, new_A8296_, new_A8297_, new_A8298_,
    new_A8299_, new_A8300_, new_A8301_, new_A8302_, new_A8303_, new_A8304_,
    new_A8305_, new_A8306_, new_A8307_, new_A8308_, new_A8309_, new_A8310_,
    new_A8311_, new_A8312_, new_A8313_, new_A8314_, new_A8315_, new_A8316_,
    new_A8317_, new_A8318_, new_A8319_, new_A8320_, new_A8321_, new_A8322_,
    new_A8323_, new_A8324_, new_A8325_, new_A8326_, new_A8327_, new_A8328_,
    new_A8329_, new_A8330_, new_A8331_, new_A8332_, new_A8333_, new_A8334_,
    new_A8335_, new_A8336_, new_A8337_, new_A8338_, new_A8339_, new_A8340_,
    new_A8341_, new_A8342_, new_A8343_, new_A8344_, new_A8345_, new_A8346_,
    new_A8347_, new_A8348_, new_A8349_, new_A8350_, new_A8351_, new_A8352_,
    new_A8353_, new_A8354_, new_A8355_, new_A8356_, new_A8357_, new_A8358_,
    new_A8359_, new_A8360_, new_A8361_, new_A8362_, new_A8363_, new_A8364_,
    new_A8365_, new_A8366_, new_A8367_, new_A8368_, new_A8369_, new_A8370_,
    new_A8371_, new_A8372_, new_A8373_, new_A8374_, new_A8375_, new_A8376_,
    new_A8377_, new_A8378_, new_A8379_, new_A8380_, new_A8381_, new_A8382_,
    new_A8383_, new_A8384_, new_A8385_, new_A8386_, new_A8387_, new_A8388_,
    new_A8389_, new_A8390_, new_A8391_, new_A8392_, new_A8393_, new_A8394_,
    new_A8395_, new_A8396_, new_A8397_, new_A8398_, new_A8399_, new_A8400_,
    new_A8401_, new_A8402_, new_A8403_, new_A8404_, new_A8405_, new_A8406_,
    new_A8407_, new_A8408_, new_A8409_, new_A8410_, new_A8411_, new_A8412_,
    new_A8413_, new_A8414_, new_A8415_, new_A8416_, new_A8417_, new_A8418_,
    new_A8419_, new_A8420_, new_A8421_, new_A8422_, new_A8423_, new_A8424_,
    new_A8425_, new_A8426_, new_A8427_, new_A8428_, new_A8429_, new_A8430_,
    new_A8431_, new_A8432_, new_A8433_, new_A8434_, new_A8435_, new_A8436_,
    new_A8437_, new_A8438_, new_A8439_, new_A8440_, new_A8441_, new_A8442_,
    new_A8443_, new_A8444_, new_A8445_, new_A8446_, new_A8447_, new_A8448_,
    new_A8449_, new_A8450_, new_A8451_, new_A8452_, new_A8453_, new_A8454_,
    new_A8455_, new_A8456_, new_A8457_, new_A8458_, new_A8459_, new_A8460_,
    new_A8461_, new_A8462_, new_A8463_, new_A8464_, new_A8465_, new_A8466_,
    new_A8467_, new_A8468_, new_A8469_, new_A8470_, new_A8471_, new_A8472_,
    new_A8473_, new_A8474_, new_A8475_, new_A8476_, new_A8477_, new_A8478_,
    new_A8479_, new_A8480_, new_A8481_, new_A8482_, new_A8483_, new_A8484_,
    new_A8485_, new_A8486_, new_A8487_, new_A8488_, new_A8489_, new_A8490_,
    new_A8491_, new_A8492_, new_A8493_, new_A8494_, new_A8495_, new_A8496_,
    new_A8497_, new_A8498_, new_A8499_, new_A8500_, new_A8501_, new_A8502_,
    new_A8503_, new_A8504_, new_A8505_, new_A8506_, new_A8507_, new_A8508_,
    new_A8509_, new_A8510_, new_A8511_, new_A8512_, new_A8513_, new_A8514_,
    new_A8515_, new_A8516_, new_A8517_, new_A8518_, new_A8519_, new_A8520_,
    new_A8521_, new_A8522_, new_A8523_, new_A8524_, new_A8525_, new_A8526_,
    new_A8527_, new_A8528_, new_A8529_, new_A8530_, new_A8531_, new_A8532_,
    new_A8533_, new_A8534_, new_A8535_, new_A8536_, new_A8537_, new_A8538_,
    new_A8539_, new_A8540_, new_A8541_, new_A8542_, new_A8543_, new_A8544_,
    new_A8545_, new_A8546_, new_A8547_, new_A8548_, new_A8549_, new_A8550_,
    new_A8551_, new_A8552_, new_A8553_, new_A8554_, new_A8555_, new_A8556_,
    new_A8557_, new_A8558_, new_A8559_, new_A8560_, new_A8561_, new_A8562_,
    new_A8563_, new_A8564_, new_A8565_, new_A8566_, new_A8567_, new_A8568_,
    new_A8569_, new_A8570_, new_A8571_, new_A8572_, new_A8573_, new_A8574_,
    new_A8575_, new_A8576_, new_A8577_, new_A8578_, new_A8579_, new_A8580_,
    new_A8581_, new_A8582_, new_A8583_, new_A8584_, new_A8585_, new_A8586_,
    new_A8587_, new_A8588_, new_A8589_, new_A8590_, new_A8591_, new_A8592_,
    new_A8593_, new_A8594_, new_A8595_, new_A8596_, new_A8597_, new_A8598_,
    new_A8599_, new_A8600_, new_A8601_, new_A8602_, new_A8603_, new_A8604_,
    new_A8605_, new_A8606_, new_A8607_, new_A8608_, new_A8609_, new_A8610_,
    new_A8611_, new_A8612_, new_A8613_, new_A8614_, new_A8615_, new_A8616_,
    new_A8617_, new_A8618_, new_A8619_, new_A8620_, new_A8621_, new_A8622_,
    new_A8623_, new_A8624_, new_A8625_, new_A8626_, new_A8627_, new_A8628_,
    new_A8629_, new_A8630_, new_A8631_, new_A8632_, new_A8633_, new_A8634_,
    new_A8635_, new_A8636_, new_A8637_, new_A8638_, new_A8639_, new_A8640_,
    new_A8641_, new_A8642_, new_A8643_, new_A8644_, new_A8645_, new_A8646_,
    new_A8647_, new_A8648_, new_A8649_, new_A8650_, new_A8651_, new_A8652_,
    new_A8653_, new_A8654_, new_A8655_, new_A8656_, new_A8657_, new_A8658_,
    new_A8659_, new_A8660_, new_A8661_, new_A8662_, new_A8663_, new_A8664_,
    new_A8665_, new_A8666_, new_A8667_, new_A8668_, new_A8669_, new_A8670_,
    new_A8671_, new_A8672_, new_A8673_, new_A8674_, new_A8675_, new_A8676_,
    new_A8677_, new_A8678_, new_A8679_, new_A8680_, new_A8681_, new_A8682_,
    new_A8683_, new_A8684_, new_A8685_, new_A8686_, new_A8687_, new_A8688_,
    new_A8689_, new_A8690_, new_A8691_, new_A8692_, new_A8693_, new_A8694_,
    new_A8695_, new_A8696_, new_A8697_, new_A8698_, new_A8699_, new_A8700_,
    new_A8701_, new_A8702_, new_A8703_, new_A8704_, new_A8705_, new_A8706_,
    new_A8707_, new_A8708_, new_A8709_, new_A8710_, new_A8711_, new_A8712_,
    new_A8713_, new_A8714_, new_A8715_, new_A8716_, new_A8717_, new_A8718_,
    new_A8719_, new_A8720_, new_A8721_, new_A8722_, new_A8723_, new_A8724_,
    new_A8725_, new_A8726_, new_A8727_, new_A8728_, new_A8729_, new_A8730_,
    new_A8731_, new_A8732_, new_A8733_, new_A8734_, new_A8735_, new_A8736_,
    new_A8737_, new_A8738_, new_A8739_, new_A8740_, new_A8741_, new_A8742_,
    new_A8743_, new_A8744_, new_A8745_, new_A8746_, new_A8747_, new_A8748_,
    new_A8749_, new_A8750_, new_A8751_, new_A8752_, new_A8753_, new_A8754_,
    new_A8755_, new_A8756_, new_A8757_, new_A8758_, new_A8759_, new_A8760_,
    new_A8761_, new_A8762_, new_A8763_, new_A8764_, new_A8765_, new_A8766_,
    new_A8767_, new_A8768_, new_A8769_, new_A8770_, new_A8771_, new_A8772_,
    new_A8773_, new_A8774_, new_A8775_, new_A8776_, new_A8777_, new_A8778_,
    new_A8779_, new_A8780_, new_A8781_, new_A8782_, new_A8783_, new_A8784_,
    new_A8785_, new_A8786_, new_A8787_, new_A8788_, new_A8789_, new_A8790_,
    new_A8791_, new_A8792_, new_A8793_, new_A8794_, new_A8795_, new_A8796_,
    new_A8797_, new_A8798_, new_A8799_, new_A8800_, new_A8801_, new_A8802_,
    new_A8803_, new_A8804_, new_A8805_, new_A8806_, new_A8807_, new_A8808_,
    new_A8809_, new_A8810_, new_A8811_, new_A8812_, new_A8813_, new_A8814_,
    new_A8815_, new_A8816_, new_A8817_, new_A8818_, new_A8819_, new_A8820_,
    new_A8821_, new_A8822_, new_A8823_, new_A8824_, new_A8825_, new_A8826_,
    new_A8827_, new_A8828_, new_A8829_, new_A8830_, new_A8831_, new_A8832_,
    new_A8833_, new_A8834_, new_A8835_, new_A8836_, new_A8837_, new_A8838_,
    new_A8839_, new_A8840_, new_A8841_, new_A8842_, new_A8843_, new_A8844_,
    new_A8845_, new_A8846_, new_A8847_, new_A8848_, new_A8849_, new_A8850_,
    new_A8851_, new_A8852_, new_A8853_, new_A8854_, new_A8855_, new_A8856_,
    new_A8857_, new_A8858_, new_A8859_, new_A8860_, new_A8861_, new_A8862_,
    new_A8863_, new_A8864_, new_A8865_, new_A8866_, new_A8867_, new_A8868_,
    new_A8869_, new_A8870_, new_A8871_, new_A8872_, new_A8873_, new_A8874_,
    new_A8875_, new_A8876_, new_A8877_, new_A8878_, new_A8879_, new_A8880_,
    new_A8881_, new_A8882_, new_A8883_, new_A8884_, new_A8885_, new_A8886_,
    new_A8887_, new_A8888_, new_A8889_, new_A8890_, new_A8891_, new_A8892_,
    new_A8893_, new_A8894_, new_A8895_, new_A8896_, new_A8897_, new_A8898_,
    new_A8899_, new_A8900_, new_A8901_, new_A8902_, new_A8903_, new_A8904_,
    new_A8905_, new_A8906_, new_A8907_, new_A8908_, new_A8909_, new_A8910_,
    new_A8911_, new_A8912_, new_A8913_, new_A8914_, new_A8915_, new_A8916_,
    new_A8917_, new_A8918_, new_A8919_, new_A8920_, new_A8921_, new_A8922_,
    new_A8923_, new_A8924_, new_A8925_, new_A8926_, new_A8927_, new_A8928_,
    new_A8929_, new_A8930_, new_A8931_, new_A8932_, new_A8933_, new_A8934_,
    new_A8935_, new_A8936_, new_A8937_, new_A8938_, new_A8939_, new_A8940_,
    new_A8941_, new_A8942_, new_A8943_, new_A8944_, new_A8945_, new_A8946_,
    new_A8947_, new_A8948_, new_A8949_, new_A8950_, new_A8951_, new_A8952_,
    new_A8953_, new_A8954_, new_A8955_, new_A8956_, new_A8957_, new_A8958_,
    new_A8959_, new_A8960_, new_A8961_, new_A8962_, new_A8963_, new_A8964_,
    new_A8965_, new_A8966_, new_A8967_, new_A8968_, new_A8969_, new_A8970_,
    new_A8971_, new_A8972_, new_A8973_, new_A8974_, new_A8975_, new_A8976_,
    new_A8977_, new_A8978_, new_A8979_, new_A8980_, new_A8981_, new_A8982_,
    new_A8983_, new_A8984_, new_A8985_, new_A8986_, new_A8987_, new_A8988_,
    new_A8989_, new_A8990_, new_A8991_, new_A8992_, new_A8993_, new_A8994_,
    new_A8995_, new_A8996_, new_A8997_, new_A8998_, new_A8999_, new_A9000_,
    new_A9001_, new_A9002_, new_A9003_, new_A9004_, new_A9005_, new_A9006_,
    new_A9007_, new_A9008_, new_A9009_, new_A9010_, new_A9011_, new_A9012_,
    new_A9013_, new_A9014_, new_A9015_, new_A9016_, new_A9017_, new_A9018_,
    new_A9019_, new_A9020_, new_A9021_, new_A9022_, new_A9023_, new_A9024_,
    new_A9025_, new_A9026_, new_A9027_, new_A9028_, new_A9029_, new_A9030_,
    new_A9031_, new_A9032_, new_A9033_, new_A9034_, new_A9035_, new_A9036_,
    new_A9037_, new_A9038_, new_A9039_, new_A9040_, new_A9041_, new_A9042_,
    new_A9043_, new_A9044_, new_A9045_, new_A9046_, new_A9047_, new_A9048_,
    new_A9049_, new_A9050_, new_A9051_, new_A9052_, new_A9053_, new_A9054_,
    new_A9055_, new_A9056_, new_A9057_, new_A9058_, new_A9059_, new_A9060_,
    new_A9061_, new_A9062_, new_A9063_, new_A9064_, new_A9065_, new_A9066_,
    new_A9067_, new_A9068_, new_A9069_, new_A9070_, new_A9071_, new_A9072_,
    new_A9073_, new_A9074_, new_A9075_, new_A9076_, new_A9077_, new_A9078_,
    new_A9079_, new_A9080_, new_A9081_, new_A9082_, new_A9083_, new_A9084_,
    new_A9085_, new_A9086_, new_A9087_, new_A9088_, new_A9089_, new_A9090_,
    new_A9091_, new_A9092_, new_A9093_, new_A9094_, new_A9095_, new_A9096_,
    new_A9097_, new_A9098_, new_A9099_, new_A9100_, new_A9101_, new_A9102_,
    new_A9103_, new_A9104_, new_A9105_, new_A9106_, new_A9107_, new_A9108_,
    new_A9109_, new_A9110_, new_A9111_, new_A9112_, new_A9113_, new_A9114_,
    new_A9115_, new_A9116_, new_A9117_, new_A9118_, new_A9119_, new_A9120_,
    new_A9121_, new_A9122_, new_A9123_, new_A9124_, new_A9125_, new_A9126_,
    new_A9127_, new_A9128_, new_A9129_, new_A9130_, new_A9131_, new_A9132_,
    new_A9133_, new_A9134_, new_A9135_, new_A9136_, new_A9137_, new_A9138_,
    new_A9139_, new_A9140_, new_A9141_, new_A9142_, new_A9143_, new_A9144_,
    new_A9145_, new_A9146_, new_A9147_, new_A9148_, new_A9149_, new_A9150_,
    new_A9151_, new_A9152_, new_A9153_, new_A9154_, new_A9155_, new_A9156_,
    new_A9157_, new_A9158_, new_A9159_, new_A9160_, new_A9161_, new_A9162_,
    new_A9163_, new_A9164_, new_A9165_, new_A9166_, new_A9167_, new_A9168_,
    new_A9169_, new_A9170_, new_A9171_, new_A9172_, new_A9173_, new_A9174_,
    new_A9175_, new_A9176_, new_A9177_, new_A9178_, new_A9179_, new_A9180_,
    new_A9181_, new_A9182_, new_A9183_, new_A9184_, new_A9185_, new_A9186_,
    new_A9187_, new_A9188_, new_A9189_, new_A9190_, new_A9191_, new_A9192_,
    new_A9193_, new_A9194_, new_A9195_, new_A9196_, new_A9197_, new_A9198_,
    new_A9199_, new_A9200_, new_A9201_, new_A9202_, new_A9203_, new_A9204_,
    new_A9205_, new_A9206_, new_A9207_, new_A9208_, new_A9209_, new_A9210_,
    new_A9211_, new_A9212_, new_A9213_, new_A9214_, new_A9215_, new_A9216_,
    new_A9217_, new_A9218_, new_A9219_, new_A9220_, new_A9221_, new_A9222_,
    new_A9223_, new_A9224_, new_A9225_, new_A9226_, new_A9227_, new_A9228_,
    new_A9229_, new_A9230_, new_A9231_, new_A9232_, new_A9233_, new_A9234_,
    new_A9235_, new_A9236_, new_A9237_, new_A9238_, new_A9239_, new_A9240_,
    new_A9241_, new_A9242_, new_A9243_, new_A9244_, new_A9245_, new_A9246_,
    new_A9247_, new_A9248_, new_A9249_, new_A9250_, new_A9251_, new_A9252_,
    new_A9253_, new_A9254_, new_A9255_, new_A9256_, new_A9257_, new_A9258_,
    new_A9259_, new_A9260_, new_A9261_, new_A9262_, new_A9263_, new_A9264_,
    new_A9265_, new_A9266_, new_A9267_, new_A9268_, new_A9269_, new_A9270_,
    new_A9271_, new_A9272_, new_A9273_, new_A9274_, new_A9275_, new_A9276_,
    new_A9277_, new_A9278_, new_A9279_, new_A9280_, new_A9281_, new_A9282_,
    new_A9283_, new_A9284_, new_A9285_, new_A9286_, new_A9287_, new_A9288_,
    new_A9289_, new_A9290_, new_A9291_, new_A9292_, new_A9293_, new_A9294_,
    new_A9295_, new_A9296_, new_A9297_, new_A9298_, new_A9299_, new_A9300_,
    new_A9301_, new_A9302_, new_A9303_, new_A9304_, new_A9305_, new_A9306_,
    new_A9307_, new_A9308_, new_A9309_, new_A9310_, new_A9311_, new_A9312_,
    new_A9313_, new_A9314_, new_A9315_, new_A9316_, new_A9317_, new_A9318_,
    new_A9319_, new_A9320_, new_A9321_, new_A9322_, new_A9323_, new_A9324_,
    new_A9325_, new_A9326_, new_A9327_, new_A9328_, new_A9329_, new_A9330_,
    new_A9331_, new_A9332_, new_A9333_, new_A9334_, new_A9335_, new_A9336_,
    new_A9337_, new_A9338_, new_A9339_, new_A9340_, new_A9341_, new_A9342_,
    new_A9343_, new_A9344_, new_A9345_, new_A9346_, new_A9347_, new_A9348_,
    new_A9349_, new_A9350_, new_A9351_, new_A9352_, new_A9353_, new_A9354_,
    new_A9355_, new_A9356_, new_A9357_, new_A9358_, new_A9359_, new_A9360_,
    new_A9361_, new_A9362_, new_A9363_, new_A9364_, new_A9365_, new_A9366_,
    new_A9367_, new_A9368_, new_A9369_, new_A9370_, new_A9371_, new_A9372_,
    new_A9373_, new_A9374_, new_A9375_, new_A9376_, new_A9377_, new_A9378_,
    new_A9379_, new_A9380_, new_A9381_, new_A9382_, new_A9383_, new_A9384_,
    new_A9385_, new_A9386_, new_A9387_, new_A9388_, new_A9389_, new_A9390_,
    new_A9391_, new_A9392_, new_A9393_, new_A9394_, new_A9395_, new_A9396_,
    new_A9397_, new_A9398_, new_A9399_, new_A9400_, new_A9401_, new_A9402_,
    new_A9403_, new_A9404_, new_A9405_, new_A9406_, new_A9407_, new_A9408_,
    new_A9409_, new_A9410_, new_A9411_, new_A9412_, new_A9413_, new_A9414_,
    new_A9415_, new_A9416_, new_A9417_, new_A9418_, new_A9419_, new_A9420_,
    new_A9421_, new_A9422_, new_A9423_, new_A9424_, new_A9425_, new_A9426_,
    new_A9427_, new_A9428_, new_A9429_, new_A9430_, new_A9431_, new_A9432_,
    new_A9433_, new_A9434_, new_A9435_, new_A9436_, new_A9437_, new_A9438_,
    new_A9439_, new_A9440_, new_A9441_, new_A9442_, new_A9443_, new_A9444_,
    new_A9445_, new_A9446_, new_A9447_, new_A9448_, new_A9449_, new_A9450_,
    new_A9451_, new_A9452_, new_A9453_, new_A9454_, new_A9455_, new_A9456_,
    new_A9457_, new_A9458_, new_A9459_, new_A9460_, new_A9461_, new_A9462_,
    new_A9463_, new_A9464_, new_A9465_, new_A9466_, new_A9467_, new_A9468_,
    new_A9469_, new_A9470_, new_A9471_, new_A9472_, new_A9473_, new_A9474_,
    new_A9475_, new_A9476_, new_A9477_, new_A9478_, new_A9479_, new_A9480_,
    new_A9481_, new_A9482_, new_A9483_, new_A9484_, new_A9485_, new_A9486_,
    new_A9487_, new_A9488_, new_A9489_, new_A9490_, new_A9491_, new_A9492_,
    new_A9493_, new_A9494_, new_A9495_, new_A9496_, new_A9497_, new_A9498_,
    new_A9499_, new_A9500_, new_A9501_, new_A9502_, new_A9503_, new_A9504_,
    new_A9505_, new_A9506_, new_A9507_, new_A9508_, new_A9509_, new_A9510_,
    new_A9511_, new_A9512_, new_A9513_, new_A9514_, new_A9515_, new_A9516_,
    new_A9517_, new_A9518_, new_A9519_, new_A9520_, new_A9521_, new_A9522_,
    new_A9523_, new_A9524_, new_A9525_, new_A9526_, new_A9527_, new_A9528_,
    new_A9529_, new_A9530_, new_A9531_, new_A9532_, new_A9533_, new_A9534_,
    new_A9535_, new_A9536_, new_A9537_, new_A9538_, new_A9539_, new_A9540_,
    new_A9541_, new_A9542_, new_A9543_, new_A9544_, new_A9545_, new_A9546_,
    new_A9547_, new_A9548_, new_A9549_, new_A9550_, new_A9551_, new_A9552_,
    new_A9553_, new_A9554_, new_A9555_, new_A9556_, new_A9557_, new_A9558_,
    new_A9559_, new_A9560_, new_A9561_, new_A9562_, new_A9563_, new_A9564_,
    new_A9565_, new_A9566_, new_A9567_, new_A9568_, new_A9569_, new_A9570_,
    new_A9571_, new_A9572_, new_A9573_, new_A9574_, new_A9575_, new_A9576_,
    new_A9577_, new_A9578_, new_A9579_, new_A9580_, new_A9581_, new_A9582_,
    new_A9583_, new_A9584_, new_A9585_, new_A9586_, new_A9587_, new_A9588_,
    new_A9589_, new_A9590_, new_A9591_, new_A9592_, new_A9593_, new_A9594_,
    new_A9595_, new_A9596_, new_A9597_, new_A9598_, new_A9599_, new_A9600_,
    new_A9601_, new_A9602_, new_A9603_, new_A9604_, new_A9605_, new_A9606_,
    new_A9607_, new_A9608_, new_A9609_, new_A9610_, new_A9611_, new_A9612_,
    new_A9613_, new_A9614_, new_A9615_, new_A9616_, new_A9617_, new_A9618_,
    new_A9619_, new_A9620_, new_A9621_, new_A9622_, new_A9623_, new_A9624_,
    new_A9625_, new_A9626_, new_A9627_, new_A9628_, new_A9629_, new_A9630_,
    new_A9631_, new_A9632_, new_A9633_, new_A9634_, new_A9635_, new_A9636_,
    new_A9637_, new_A9638_, new_A9639_, new_A9640_, new_A9641_, new_A9642_,
    new_A9643_, new_A9644_, new_A9645_, new_A9646_, new_A9647_, new_A9648_,
    new_A9649_, new_A9650_, new_A9651_, new_A9652_, new_A9653_, new_A9654_,
    new_A9655_, new_A9656_, new_A9657_, new_A9658_, new_A9659_, new_A9660_,
    new_A9661_, new_A9662_, new_A9663_, new_A9664_, new_A9665_, new_A9666_,
    new_A9667_, new_A9668_, new_A9669_, new_A9670_, new_A9671_, new_A9672_,
    new_A9673_, new_A9674_, new_A9675_, new_A9676_, new_A9677_, new_A9678_,
    new_A9679_, new_A9680_, new_A9681_, new_A9682_, new_A9683_, new_A9684_,
    new_A9685_, new_A9686_, new_A9687_, new_A9688_, new_A9689_, new_A9690_,
    new_A9691_, new_A9692_, new_A9693_, new_A9694_, new_A9695_, new_A9696_,
    new_A9697_, new_A9698_, new_A9699_, new_A9700_, new_A9701_, new_A9702_,
    new_A9703_, new_A9704_, new_A9705_, new_A9706_, new_A9707_, new_A9708_,
    new_A9709_, new_A9710_, new_A9711_, new_A9712_, new_A9713_, new_A9714_,
    new_A9715_, new_A9716_, new_A9717_, new_A9718_, new_A9719_, new_A9720_,
    new_A9721_, new_A9722_, new_A9723_, new_A9724_, new_A9725_, new_A9726_,
    new_A9727_, new_A9728_, new_A9729_, new_A9730_, new_A9731_, new_A9732_,
    new_A9733_, new_A9734_, new_A9735_, new_A9736_, new_A9737_, new_A9738_,
    new_A9739_, new_A9740_, new_A9741_, new_A9742_, new_A9743_, new_A9744_,
    new_A9745_, new_A9746_, new_A9747_, new_A9748_, new_A9749_, new_A9750_,
    new_A9751_, new_A9752_, new_A9753_, new_A9754_, new_A9755_, new_A9756_,
    new_A9757_, new_A9758_, new_A9759_, new_A9760_, new_A9761_, new_A9762_,
    new_A9763_, new_A9764_, new_A9765_, new_A9766_, new_A9767_, new_A9768_,
    new_A9769_, new_A9770_, new_A9771_, new_A9772_, new_A9773_, new_A9774_,
    new_A9775_, new_A9776_, new_A9777_, new_A9778_, new_A9779_, new_A9780_,
    new_A9781_, new_A9782_, new_A9783_, new_A9784_, new_A9785_, new_A9786_,
    new_A9787_, new_A9788_, new_A9789_, new_A9790_, new_A9791_, new_A9792_,
    new_A9793_, new_A9794_, new_A9795_, new_A9796_, new_A9797_, new_A9798_,
    new_A9799_, new_A9800_, new_A9801_, new_A9802_, new_A9803_, new_A9804_,
    new_A9805_, new_A9806_, new_A9807_, new_A9808_, new_A9809_, new_A9810_,
    new_A9811_, new_A9812_, new_A9813_, new_A9814_, new_A9815_, new_A9816_,
    new_A9817_, new_A9818_, new_A9819_, new_A9820_, new_A9821_, new_A9822_,
    new_A9823_, new_A9824_, new_A9825_, new_A9826_, new_A9827_, new_A9828_,
    new_A9829_, new_A9830_, new_A9831_, new_A9832_, new_A9833_, new_A9834_,
    new_A9835_, new_A9836_, new_A9837_, new_A9838_, new_A9839_, new_A9840_,
    new_A9841_, new_A9842_, new_A9843_, new_A9844_, new_A9845_, new_A9846_,
    new_A9847_, new_A9848_, new_A9849_, new_A9850_, new_A9851_, new_A9852_,
    new_A9853_, new_A9854_, new_A9855_, new_A9856_, new_A9857_, new_A9858_,
    new_A9859_, new_A9860_, new_A9861_, new_A9862_, new_A9863_, new_A9864_,
    new_A9865_, new_A9866_, new_A9867_, new_A9868_, new_A9869_, new_A9870_,
    new_A9871_, new_A9872_, new_A9873_, new_A9874_, new_A9875_, new_A9876_,
    new_A9877_, new_A9878_, new_A9879_, new_A9880_, new_A9881_, new_A9882_,
    new_A9883_, new_A9884_, new_A9885_, new_A9886_, new_A9887_, new_A9888_,
    new_A9889_, new_A9890_, new_A9891_, new_A9892_, new_A9893_, new_A9894_,
    new_A9895_, new_A9896_, new_A9897_, new_A9898_, new_A9899_, new_A9900_,
    new_A9901_, new_A9902_, new_A9903_, new_A9904_, new_A9905_, new_A9906_,
    new_A9907_, new_A9908_, new_A9909_, new_A9910_, new_A9911_, new_A9912_,
    new_A9913_, new_A9914_, new_A9915_, new_A9916_, new_A9917_, new_A9918_,
    new_A9919_, new_A9920_, new_A9921_, new_A9922_, new_A9923_, new_A9924_,
    new_A9925_, new_A9926_, new_A9927_, new_A9928_, new_A9929_, new_A9930_,
    new_A9931_, new_A9932_, new_A9933_, new_A9934_, new_A9935_, new_A9936_,
    new_A9937_, new_A9938_, new_A9939_, new_A9940_, new_A9941_, new_A9942_,
    new_A9943_, new_A9944_, new_A9945_, new_A9946_, new_A9947_, new_A9948_,
    new_A9949_, new_A9950_, new_A9951_, new_A9952_, new_A9953_, new_A9954_,
    new_A9955_, new_A9956_, new_A9957_, new_A9958_, new_A9959_, new_A9960_,
    new_A9961_, new_A9962_, new_A9963_, new_A9964_, new_A9965_, new_A9966_,
    new_A9967_, new_A9968_, new_A9969_, new_A9970_, new_A9971_, new_A9972_,
    new_A9973_, new_A9974_, new_A9975_, new_A9976_, new_A9977_, new_A9978_,
    new_A9979_, new_A9980_, new_A9981_, new_A9982_, new_A9983_, new_A9984_,
    new_A9985_, new_A9986_, new_A9987_, new_A9988_, new_A9989_, new_A9990_,
    new_A9991_, new_A9992_, new_A9993_, new_A9994_, new_A9995_, new_A9996_,
    new_A9997_, new_A9998_, new_A9999_, new_B1_, new_B2_, new_B3_, new_B4_,
    new_B5_, new_B6_, new_B7_, new_B8_, new_B9_, new_B10_, new_B11_,
    new_B12_, new_B13_, new_B14_, new_B15_, new_B16_, new_B17_, new_B18_,
    new_B19_, new_B20_, new_B21_, new_B22_, new_B23_, new_B24_, new_B25_,
    new_B26_, new_B27_, new_B28_, new_B29_, new_B30_, new_B31_, new_B32_,
    new_B33_, new_B34_, new_B35_, new_B36_, new_B37_, new_B38_, new_B39_,
    new_B40_, new_B41_, new_B42_, new_B43_, new_B44_, new_B45_, new_B46_,
    new_B47_, new_B48_, new_B49_, new_B50_, new_B51_, new_B52_, new_B53_,
    new_B54_, new_B55_, new_B56_, new_B57_, new_B58_, new_B59_, new_B60_,
    new_B61_, new_B62_, new_B63_, new_B64_, new_B65_, new_B66_, new_B67_,
    new_B68_, new_B69_, new_B70_, new_B71_, new_B72_, new_B73_, new_B74_,
    new_B75_, new_B76_, new_B77_, new_B78_, new_B79_, new_B80_, new_B81_,
    new_B82_, new_B83_, new_B84_, new_B85_, new_B86_, new_B87_, new_B88_,
    new_B89_, new_B90_, new_B91_, new_B92_, new_B93_, new_B94_, new_B95_,
    new_B96_, new_B97_, new_B98_, new_B99_, new_B100_, new_B101_,
    new_B102_, new_B103_, new_B104_, new_B105_, new_B106_, new_B107_,
    new_B108_, new_B109_, new_B110_, new_B111_, new_B112_, new_B113_,
    new_B114_, new_B115_, new_B116_, new_B117_, new_B118_, new_B119_,
    new_B120_, new_B121_, new_B122_, new_B123_, new_B124_, new_B125_,
    new_B126_, new_B127_, new_B128_, new_B129_, new_B130_, new_B131_,
    new_B132_, new_B133_, new_B134_, new_B135_, new_B136_, new_B137_,
    new_B138_, new_B139_, new_B140_, new_B141_, new_B142_, new_B143_,
    new_B144_, new_B145_, new_B146_, new_B147_, new_B148_, new_B149_,
    new_B150_, new_B151_, new_B152_, new_B153_, new_B154_, new_B155_,
    new_B156_, new_B157_, new_B158_, new_B159_, new_B160_, new_B161_,
    new_B162_, new_B163_, new_B164_, new_B165_, new_B166_, new_B167_,
    new_B168_, new_B169_, new_B170_, new_B171_, new_B172_, new_B173_,
    new_B174_, new_B175_, new_B176_, new_B177_, new_B178_, new_B179_,
    new_B180_, new_B181_, new_B182_, new_B183_, new_B184_, new_B185_,
    new_B186_, new_B187_, new_B188_, new_B189_, new_B190_, new_B191_,
    new_B192_, new_B193_, new_B194_, new_B195_, new_B196_, new_B197_,
    new_B198_, new_B199_, new_B200_, new_B201_, new_B202_, new_B203_,
    new_B204_, new_B205_, new_B206_, new_B207_, new_B208_, new_B209_,
    new_B210_, new_B211_, new_B212_, new_B213_, new_B214_, new_B215_,
    new_B216_, new_B217_, new_B218_, new_B219_, new_B220_, new_B221_,
    new_B222_, new_B223_, new_B224_, new_B225_, new_B226_, new_B227_,
    new_B228_, new_B229_, new_B230_, new_B231_, new_B232_, new_B233_,
    new_B234_, new_B235_, new_B236_, new_B237_, new_B238_, new_B239_,
    new_B240_, new_B241_, new_B242_, new_B243_, new_B244_, new_B245_,
    new_B246_, new_B247_, new_B248_, new_B249_, new_B250_, new_B251_,
    new_B252_, new_B253_, new_B254_, new_B255_, new_B256_, new_B257_,
    new_B258_, new_B259_, new_B260_, new_B261_, new_B262_, new_B263_,
    new_B264_, new_B265_, new_B266_, new_B267_, new_B268_, new_B269_,
    new_B270_, new_B271_, new_B272_, new_B273_, new_B274_, new_B275_,
    new_B276_, new_B277_, new_B278_, new_B279_, new_B280_, new_B281_,
    new_B282_, new_B283_, new_B284_, new_B285_, new_B286_, new_B287_,
    new_B288_, new_B289_, new_B290_, new_B291_, new_B292_, new_B293_,
    new_B294_, new_B295_, new_B296_, new_B297_, new_B298_, new_B299_,
    new_B300_, new_B301_, new_B302_, new_B303_, new_B304_, new_B305_,
    new_B306_, new_B307_, new_B308_, new_B309_, new_B310_, new_B311_,
    new_B312_, new_B313_, new_B314_, new_B315_, new_B316_, new_B317_,
    new_B318_, new_B319_, new_B320_, new_B321_, new_B322_, new_B323_,
    new_B324_, new_B325_, new_B326_, new_B327_, new_B328_, new_B329_,
    new_B330_, new_B331_, new_B332_, new_B333_, new_B334_, new_B335_,
    new_B336_, new_B337_, new_B338_, new_B339_, new_B340_, new_B341_,
    new_B342_, new_B343_, new_B344_, new_B345_, new_B346_, new_B347_,
    new_B348_, new_B349_, new_B350_, new_B351_, new_B352_, new_B353_,
    new_B354_, new_B355_, new_B356_, new_B357_, new_B358_, new_B359_,
    new_B360_, new_B361_, new_B362_, new_B363_, new_B364_, new_B365_,
    new_B366_, new_B367_, new_B368_, new_B369_, new_B370_, new_B371_,
    new_B372_, new_B373_, new_B374_, new_B375_, new_B376_, new_B377_,
    new_B378_, new_B379_, new_B380_, new_B381_, new_B382_, new_B383_,
    new_B384_, new_B385_, new_B386_, new_B387_, new_B388_, new_B389_,
    new_B390_, new_B391_, new_B392_, new_B393_, new_B394_, new_B395_,
    new_B396_, new_B397_, new_B398_, new_B399_, new_B400_, new_B401_,
    new_B402_, new_B403_, new_B404_, new_B405_, new_B406_, new_B407_,
    new_B408_, new_B409_, new_B410_, new_B411_, new_B412_, new_B413_,
    new_B414_, new_B415_, new_B416_, new_B417_, new_B418_, new_B419_,
    new_B420_, new_B421_, new_B422_, new_B423_, new_B424_, new_B425_,
    new_B426_, new_B427_, new_B428_, new_B429_, new_B430_, new_B431_,
    new_B432_, new_B433_, new_B434_, new_B435_, new_B436_, new_B437_,
    new_B438_, new_B439_, new_B440_, new_B441_, new_B442_, new_B443_,
    new_B444_, new_B445_, new_B446_, new_B447_, new_B448_, new_B449_,
    new_B450_, new_B451_, new_B452_, new_B453_, new_B454_, new_B455_,
    new_B456_, new_B457_, new_B458_, new_B459_, new_B460_, new_B461_,
    new_B462_, new_B463_, new_B464_, new_B465_, new_B466_, new_B467_,
    new_B468_, new_B469_, new_B470_, new_B471_, new_B472_, new_B473_,
    new_B474_, new_B475_, new_B476_, new_B477_, new_B478_, new_B479_,
    new_B480_, new_B481_, new_B482_, new_B483_, new_B484_, new_B485_,
    new_B486_, new_B487_, new_B488_, new_B489_, new_B490_, new_B491_,
    new_B492_, new_B493_, new_B494_, new_B495_, new_B496_, new_B497_,
    new_B498_, new_B499_, new_B500_, new_B501_, new_B502_, new_B503_,
    new_B504_, new_B505_, new_B506_, new_B507_, new_B508_, new_B509_,
    new_B510_, new_B511_, new_B512_, new_B513_, new_B514_, new_B515_,
    new_B516_, new_B517_, new_B518_, new_B519_, new_B520_, new_B521_,
    new_B522_, new_B523_, new_B524_, new_B525_, new_B526_, new_B527_,
    new_B528_, new_B529_, new_B530_, new_B531_, new_B532_, new_B533_,
    new_B534_, new_B535_, new_B536_, new_B537_, new_B538_, new_B539_,
    new_B540_, new_B541_, new_B542_, new_B543_, new_B544_, new_B545_,
    new_B546_, new_B547_, new_B548_, new_B549_, new_B550_, new_B551_,
    new_B552_, new_B553_, new_B554_, new_B555_, new_B556_, new_B557_,
    new_B558_, new_B559_, new_B560_, new_B561_, new_B562_, new_B563_,
    new_B564_, new_B565_, new_B566_, new_B567_, new_B568_, new_B569_,
    new_B570_, new_B571_, new_B572_, new_B573_, new_B574_, new_B575_,
    new_B576_, new_B577_, new_B578_, new_B579_, new_B580_, new_B581_,
    new_B582_, new_B583_, new_B584_, new_B585_, new_B586_, new_B587_,
    new_B588_, new_B589_, new_B590_, new_B591_, new_B592_, new_B593_,
    new_B594_, new_B595_, new_B596_, new_B597_, new_B598_, new_B599_,
    new_B600_, new_B601_, new_B602_, new_B603_, new_B604_, new_B605_,
    new_B606_, new_B607_, new_B608_, new_B609_, new_B610_, new_B611_,
    new_B612_, new_B613_, new_B614_, new_B615_, new_B616_, new_B617_,
    new_B618_, new_B619_, new_B620_, new_B621_, new_B622_, new_B623_,
    new_B624_, new_B625_, new_B626_, new_B627_, new_B628_, new_B629_,
    new_B630_, new_B631_, new_B632_, new_B633_, new_B634_, new_B635_,
    new_B636_, new_B637_, new_B638_, new_B639_, new_B640_, new_B641_,
    new_B642_, new_B643_, new_B644_, new_B645_, new_B646_, new_B647_,
    new_B648_, new_B649_, new_B650_, new_B651_, new_B652_, new_B653_,
    new_B654_, new_B655_, new_B656_, new_B657_, new_B658_, new_B659_,
    new_B660_, new_B661_, new_B662_, new_B663_, new_B664_, new_B665_,
    new_B666_, new_B667_, new_B668_, new_B669_, new_B670_, new_B671_,
    new_B672_, new_B673_, new_B674_, new_B675_, new_B676_, new_B677_,
    new_B678_, new_B679_, new_B680_, new_B681_, new_B682_, new_B683_,
    new_B684_, new_B685_, new_B686_, new_B687_, new_B688_, new_B689_,
    new_B690_, new_B691_, new_B692_, new_B693_, new_B694_, new_B695_,
    new_B696_, new_B697_, new_B698_, new_B699_, new_B700_, new_B701_,
    new_B702_, new_B703_, new_B704_, new_B705_, new_B706_, new_B707_,
    new_B708_, new_B709_, new_B710_, new_B711_, new_B712_, new_B713_,
    new_B714_, new_B715_, new_B716_, new_B717_, new_B718_, new_B719_,
    new_B720_, new_B721_, new_B722_, new_B723_, new_B724_, new_B725_,
    new_B726_, new_B727_, new_B728_, new_B729_, new_B730_, new_B731_,
    new_B732_, new_B733_, new_B734_, new_B735_, new_B736_, new_B737_,
    new_B738_, new_B739_, new_B740_, new_B741_, new_B742_, new_B743_,
    new_B744_, new_B745_, new_B746_, new_B747_, new_B748_, new_B749_,
    new_B750_, new_B751_, new_B752_, new_B753_, new_B754_, new_B755_,
    new_B756_, new_B757_, new_B758_, new_B759_, new_B760_, new_B761_,
    new_B762_, new_B763_, new_B764_, new_B765_, new_B766_, new_B767_,
    new_B768_, new_B769_, new_B770_, new_B771_, new_B772_, new_B773_,
    new_B774_, new_B775_, new_B776_, new_B777_, new_B778_, new_B779_,
    new_B780_, new_B781_, new_B782_, new_B783_, new_B784_, new_B785_,
    new_B786_, new_B787_, new_B788_, new_B789_, new_B790_, new_B791_,
    new_B792_, new_B793_, new_B794_, new_B795_, new_B796_, new_B797_,
    new_B798_, new_B799_, new_B800_, new_B801_, new_B802_, new_B803_,
    new_B804_, new_B805_, new_B806_, new_B807_, new_B808_, new_B809_,
    new_B810_, new_B811_, new_B812_, new_B813_, new_B814_, new_B815_,
    new_B816_, new_B817_, new_B818_, new_B819_, new_B820_, new_B821_,
    new_B822_, new_B823_, new_B824_, new_B825_, new_B826_, new_B827_,
    new_B828_, new_B829_, new_B830_, new_B831_, new_B832_, new_B833_,
    new_B834_, new_B835_, new_B836_, new_B837_, new_B838_, new_B839_,
    new_B840_, new_B841_, new_B842_, new_B843_, new_B844_, new_B845_,
    new_B846_, new_B847_, new_B848_, new_B849_, new_B850_, new_B851_,
    new_B852_, new_B853_, new_B854_, new_B855_, new_B856_, new_B857_,
    new_B858_, new_B859_, new_B860_, new_B861_, new_B862_, new_B863_,
    new_B864_, new_B865_, new_B866_, new_B867_, new_B868_, new_B869_,
    new_B870_, new_B871_, new_B872_, new_B873_, new_B874_, new_B875_,
    new_B876_, new_B877_, new_B878_, new_B879_, new_B880_, new_B881_,
    new_B882_, new_B883_, new_B884_, new_B885_, new_B886_, new_B887_,
    new_B888_, new_B889_, new_B890_, new_B891_, new_B892_, new_B893_,
    new_B894_, new_B895_, new_B896_, new_B897_, new_B898_, new_B899_,
    new_B900_, new_B901_, new_B902_, new_B903_, new_B904_, new_B905_,
    new_B906_, new_B907_, new_B908_, new_B909_, new_B910_, new_B911_,
    new_B912_, new_B913_, new_B914_, new_B915_, new_B916_, new_B917_,
    new_B918_, new_B919_, new_B920_, new_B921_, new_B922_, new_B923_,
    new_B924_, new_B925_, new_B926_, new_B927_, new_B928_, new_B929_,
    new_B930_, new_B931_, new_B932_, new_B933_, new_B934_, new_B935_,
    new_B936_, new_B937_, new_B938_, new_B939_, new_B940_, new_B941_,
    new_B942_, new_B943_, new_B944_, new_B945_, new_B946_, new_B947_,
    new_B948_, new_B949_, new_B950_, new_B951_, new_B952_, new_B953_,
    new_B954_, new_B955_, new_B956_, new_B957_, new_B958_, new_B959_,
    new_B960_, new_B961_, new_B962_, new_B963_, new_B964_, new_B965_,
    new_B966_, new_B967_, new_B968_, new_B969_, new_B970_, new_B971_,
    new_B972_, new_B973_, new_B974_, new_B975_, new_B976_, new_B977_,
    new_B978_, new_B979_, new_B980_, new_B981_, new_B982_, new_B983_,
    new_B984_, new_B985_, new_B986_, new_B987_, new_B988_, new_B989_,
    new_B990_, new_B991_, new_B992_, new_B993_, new_B994_, new_B995_,
    new_B996_, new_B997_, new_B998_, new_B999_, new_B1000_, new_B1001_,
    new_B1002_, new_B1003_, new_B1004_, new_B1005_, new_B1006_, new_B1007_,
    new_B1008_, new_B1009_, new_B1010_, new_B1011_, new_B1012_, new_B1013_,
    new_B1014_, new_B1015_, new_B1016_, new_B1017_, new_B1018_, new_B1019_,
    new_B1020_, new_B1021_, new_B1022_, new_B1023_, new_B1024_, new_B1025_,
    new_B1026_, new_B1027_, new_B1028_, new_B1029_, new_B1030_, new_B1031_,
    new_B1032_, new_B1033_, new_B1034_, new_B1035_, new_B1036_, new_B1037_,
    new_B1038_, new_B1039_, new_B1040_, new_B1041_, new_B1042_, new_B1043_,
    new_B1044_, new_B1045_, new_B1046_, new_B1047_, new_B1048_, new_B1049_,
    new_B1050_, new_B1051_, new_B1052_, new_B1053_, new_B1054_, new_B1055_,
    new_B1056_, new_A6930_, new_A6929_, new_A6928_, new_A6927_, new_A6926_,
    new_A6925_, new_A6924_, new_A6923_, new_A6922_, new_A6921_, new_A6920_,
    new_A6919_, new_A6918_, new_A6917_, new_A6916_, new_A6915_, new_A6914_,
    new_A6913_, new_A6912_, new_A6911_, new_A6910_, new_A6909_, new_A6908_,
    new_A6902_, new_A6901_, new_A6900_, new_A6899_, new_A6898_, new_A6897_,
    new_A6896_, new_A6895_, new_A6894_, new_A6893_, new_A6892_, new_A6891_,
    new_A6890_, new_A6889_, new_A6888_, new_A6887_, new_A6886_, new_A6885_,
    new_A6884_, new_A6883_, new_A6882_, new_A6881_, new_A6880_, new_A6879_,
    new_A6878_, new_A6877_, new_A6876_, new_A6875_, new_A6869_, new_A6868_,
    new_A6867_, new_A6866_, new_A6865_, new_A6864_, new_A6863_, new_A6862_,
    new_A6861_, new_A6860_, new_A6859_, new_A6858_, new_A6857_, new_A6856_,
    new_A6855_, new_A6854_, new_A6853_, new_A6852_, new_A6851_, new_A6850_,
    new_A6849_, new_A6848_, new_A6847_, new_A6846_, new_A6845_, new_A6844_,
    new_A6843_, new_A6842_, new_A6836_, new_A6835_, new_A6834_, new_A6833_,
    new_A6832_, new_A6831_, new_A6830_, new_A6829_, new_A6828_, new_A6827_,
    new_A6826_, new_A6825_, new_A6824_, new_A6823_, new_A6822_, new_A6821_,
    new_A6820_, new_A6819_, new_A6818_, new_A6817_, new_A6816_, new_A6815_,
    new_A6814_, new_A6813_, new_A6812_, new_A6811_, new_A6810_, new_A6809_,
    new_A6803_, new_A6802_, new_A6801_, new_A6800_, new_A6799_, new_A6798_,
    new_A6797_, new_A6796_, new_A6795_, new_A6794_, new_A6793_, new_A6792_,
    new_A6791_, new_A6790_, new_A6789_, new_A6788_, new_A6787_, new_A6786_,
    new_A6785_, new_A6784_, new_A6783_, new_A6782_, new_A6781_, new_A6780_,
    new_A6779_, new_A6778_, new_A6777_, new_A6776_, new_A6770_, new_A6769_,
    new_A6768_, new_A6767_, new_A6766_, new_A6765_, new_A6764_, new_A6763_,
    new_A6762_, new_A6761_, new_A6760_, new_A6759_, new_A6758_, new_A6757_,
    new_A6756_, new_A6755_, new_A6754_, new_A6753_, new_A6752_, new_A6751_,
    new_A6750_, new_A6749_, new_A6748_, new_A6747_, new_A6746_, new_A6745_,
    new_A6744_, new_A6743_, new_A6737_, new_A6736_, new_A6735_, new_A6734_,
    new_A6733_, new_A6732_, new_A6731_, new_A6730_, new_A6729_, new_A6728_,
    new_A6727_, new_A6726_, new_A6725_, new_A6724_, new_A6723_, new_A6722_,
    new_A6721_, new_A6720_, new_A6719_, new_A6718_, new_A6717_, new_A6716_,
    new_A6715_, new_A6714_, new_A6713_, new_A6712_, new_A6711_, new_A6710_,
    new_A6704_, new_A6703_, new_A6702_, new_A6701_, new_A6700_, new_A6699_,
    new_A6698_, new_A6697_, new_A6696_, new_A6695_, new_A6694_, new_A6693_,
    new_A6692_, new_A6691_, new_A6690_, new_A6689_, new_A6688_, new_A6687_,
    new_A6686_, new_A6685_, new_A6684_, new_A6683_, new_A6682_, new_A6681_,
    new_A6680_, new_A6679_, new_A6678_, new_A6677_, new_A6671_, new_A6670_,
    new_A6669_, new_A6668_, new_A6667_, new_A6666_, new_A6665_, new_A6664_,
    new_A6663_, new_A6662_, new_A6661_, new_A6660_, new_A6659_, new_A6658_,
    new_A6657_, new_A6656_, new_A6655_, new_A6654_, new_A6653_, new_A6652_,
    new_A6651_, new_A6650_, new_A6649_, new_A6648_, new_A6647_, new_A6646_,
    new_A6645_, new_A6644_, new_A6638_, new_A6637_, new_A6636_, new_A6635_,
    new_A6634_, new_A6633_, new_A6632_, new_A6631_, new_A6630_, new_A6629_,
    new_A6628_, new_A6627_, new_A6626_, new_A6625_, new_A6624_, new_A6623_,
    new_A6622_, new_A6621_, new_A6620_, new_A6619_, new_A6618_, new_A6617_,
    new_A6616_, new_A6615_, new_A6614_, new_A6613_, new_A6612_, new_A6611_,
    new_A6605_, new_A6604_, new_A6603_, new_A6602_, new_A6601_, new_A6600_,
    new_A6599_, new_A6598_, new_A6597_, new_A6596_, new_A6595_, new_A6594_,
    new_A6593_, new_A6592_, new_A6591_, new_A6590_, new_A6589_, new_A6588_,
    new_A6587_, new_A6586_, new_A6585_, new_A6584_, new_A6583_, new_A6582_,
    new_A6581_, new_A6580_, new_A6579_, new_A6578_, new_A6572_, new_A6571_,
    new_A6570_, new_A6569_, new_A6568_, new_A6567_, new_A6566_, new_A6565_,
    new_A6564_, new_A6563_, new_A6562_, new_A6561_, new_A6560_, new_A6559_,
    new_A6558_, new_A6557_, new_A6556_, new_A6555_, new_A6554_, new_A6553_,
    new_A6552_, new_A6551_, new_A6550_, new_A6549_, new_A6548_, new_A6547_,
    new_A6546_, new_A6545_, new_A6539_, new_A6538_, new_A6537_, new_A6536_,
    new_A6535_, new_A6534_, new_A6533_, new_A6532_, new_A6531_, new_A6530_,
    new_A6529_, new_A6528_, new_A6527_, new_A6526_, new_A6525_, new_A6524_,
    new_A6523_, new_A6522_, new_A6521_, new_A6520_, new_A6519_, new_A6518_,
    new_A6517_, new_A6516_, new_A6515_, new_A6514_, new_A6513_, new_A6512_,
    new_A6506_, new_A6505_, new_A6504_, new_A6503_, new_A6502_, new_A6501_,
    new_A6500_, new_A6499_, new_A6498_, new_A6497_, new_A6496_, new_A6495_,
    new_A6494_, new_A6493_, new_A6492_, new_A6491_, new_A6490_, new_A6489_,
    new_A6488_, new_A6487_, new_A6486_, new_A6485_, new_A6484_, new_A6483_,
    new_A6482_, new_A6481_, new_A6480_, new_A6479_, new_A6473_, new_A6472_,
    new_A6471_, new_A6470_, new_A6469_, new_A6468_, new_A6467_, new_A6466_,
    new_A6465_, new_A6464_, new_A6463_, new_A6462_, new_A6461_, new_A6460_,
    new_A6459_, new_A6458_, new_A6457_, new_A6456_, new_A6455_, new_A6454_,
    new_A6453_, new_A6452_, new_A6451_, new_A6450_, new_A6449_, new_A6448_,
    new_A6447_, new_A6446_, new_A6440_, new_A6439_, new_A6438_, new_A6437_,
    new_A6436_, new_A6435_, new_A6434_, new_A6433_, new_A6432_, new_A6431_,
    new_A6430_, new_A6429_, new_A6428_, new_A6427_, new_A6426_, new_A6425_,
    new_A6424_, new_A6423_, new_A6422_, new_A6421_, new_A6420_, new_A6419_,
    new_A6418_, new_A6417_, new_A6416_, new_A6415_, new_A6414_, new_A6413_,
    new_A6407_, new_A6406_, new_A6405_, new_A6404_, new_A6403_, new_A6402_,
    new_A6401_, new_A6400_, new_A6399_, new_A6398_, new_A6397_, new_A6396_,
    new_A6395_, new_A6394_, new_A6393_, new_A6392_, new_A6391_, new_A6390_,
    new_A6389_, new_A6388_, new_A6387_, new_A6386_, new_A6385_, new_A6384_,
    new_A6383_, new_A6382_, new_A6381_, new_A6380_, new_A6374_, new_A6373_,
    new_A6372_, new_A6371_, new_A6370_, new_A6369_, new_A6368_, new_A6367_,
    new_A6366_, new_A6365_, new_A6364_, new_A6363_, new_A6362_, new_A6361_,
    new_A6360_, new_A6359_, new_A6358_, new_A6357_, new_A6356_, new_A6355_,
    new_A6354_, new_A6353_, new_A6352_, new_A6351_, new_A6350_, new_A6349_,
    new_A6348_, new_A6347_, new_A6341_, new_A6340_, new_A6339_, new_A6338_,
    new_A6337_, new_A6336_, new_A6335_, new_A6334_, new_A6333_, new_A6332_,
    new_A6331_, new_A6330_, new_A6329_, new_A6328_, new_A6327_, new_A6326_,
    new_A6325_, new_A6324_, new_A6323_, new_A6322_, new_A6321_, new_A6320_,
    new_A6319_, new_A6318_, new_A6317_, new_A6316_, new_A6315_, new_A6314_,
    new_A6308_, new_A6307_, new_A6306_, new_A6305_, new_A6304_, new_A6303_,
    new_A6302_, new_A6301_, new_A6300_, new_A6299_, new_A6298_, new_A6297_,
    new_A6296_, new_A6295_, new_A6294_, new_A6293_, new_A6292_, new_A6291_,
    new_A6290_, new_A6289_, new_A6288_, new_A6287_, new_A6286_, new_A6285_,
    new_A6284_, new_A6283_, new_A6282_, new_A6281_, new_A6275_, new_A6274_,
    new_A6273_, new_A6272_, new_A6271_, new_A6270_, new_A6269_, new_A6268_,
    new_A6267_, new_A6266_, new_A6265_, new_A6264_, new_A6263_, new_A6262_,
    new_A6261_, new_A6260_, new_A6259_, new_A6258_, new_A6257_, new_A6256_,
    new_A6255_, new_A6254_, new_A6253_, new_A6252_, new_A6251_, new_A6250_,
    new_A6249_, new_A6248_, new_A6242_, new_A6241_, new_A6240_, new_A6239_,
    new_A6238_, new_A6237_, new_A6236_, new_A6235_, new_A6234_, new_A6233_,
    new_A6232_, new_A6231_, new_A6230_, new_A6229_, new_A6228_, new_A6227_,
    new_A6226_, new_A6225_, new_A6224_, new_A6223_, new_A6222_, new_A6221_,
    new_A6220_, new_A6219_, new_A6218_, new_A6217_, new_A6216_, new_A6215_,
    new_A6209_, new_A6208_, new_A6207_, new_A6206_, new_A6205_, new_A6204_,
    new_A6203_, new_A6202_, new_A6201_, new_A6200_, new_A6199_, new_A6198_,
    new_A6197_, new_A6196_, new_A6195_, new_A6194_, new_A6193_, new_A6192_,
    new_A6191_, new_A6190_, new_A6189_, new_A6188_, new_A6187_, new_A6186_,
    new_A6185_, new_A6184_, new_A6183_, new_A6182_, new_A6176_, new_A6175_,
    new_A6174_, new_A6173_, new_A6172_, new_A6171_, new_A6170_, new_A6169_,
    new_A6168_, new_A6167_, new_A6166_, new_A6165_, new_A6164_, new_A6163_,
    new_A6162_, new_A6161_, new_A6160_, new_A6159_, new_A6158_, new_A6157_,
    new_A6156_, new_A6155_, new_A6154_, new_A6153_, new_A6152_, new_A6151_,
    new_A6150_, new_A6149_, new_A6143_, new_A6142_, new_A6141_, new_A6140_,
    new_A6139_, new_A6138_, new_A6137_, new_A6136_, new_A6135_, new_A6134_,
    new_A6133_, new_A6132_, new_A6131_, new_A6130_, new_A6129_, new_A6128_,
    new_A6127_, new_A6126_, new_A6125_, new_A6124_, new_A6123_, new_A6122_,
    new_A6121_, new_A6120_, new_A6119_, new_A6118_, new_A6117_, new_A6116_,
    new_A6110_, new_A6109_, new_A6108_, new_A6107_, new_A6106_, new_A6105_,
    new_A6104_, new_A6103_, new_A6102_, new_A6101_, new_A6100_, new_A6099_,
    new_A6098_, new_A6097_, new_A6096_, new_A6095_, new_A6094_, new_A6093_,
    new_A6092_, new_A6091_, new_A6090_, new_A6089_, new_A6088_, new_A6087_,
    new_A6086_, new_A6085_, new_A6084_, new_A6083_, new_A6077_, new_A6076_,
    new_A6075_, new_A6074_, new_A6073_, new_A6072_, new_A6071_, new_A6070_,
    new_A6069_, new_A6068_, new_A6067_, new_A6066_, new_A6065_, new_A6064_,
    new_A6063_, new_A6062_, new_A6061_, new_A6060_, new_A6059_, new_A6058_,
    new_A6057_, new_A6056_, new_A6055_, new_A6054_, new_A6053_, new_A6052_,
    new_A6051_, new_A6050_, new_A6044_, new_A6043_, new_A6042_, new_A6041_,
    new_A6040_, new_A6039_, new_A6038_, new_A6037_, new_A6036_, new_A6035_,
    new_A6034_, new_A6033_, new_A6032_, new_A6031_, new_A6030_, new_A6029_,
    new_A6028_, new_A6027_, new_A6026_, new_A6025_, new_A6024_, new_A6023_,
    new_A6022_, new_A6021_, new_A6020_, new_A6019_, new_A6018_, new_A6017_,
    new_A6011_, new_A6010_, new_A6009_, new_A6008_, new_A6007_, new_A6006_,
    new_A6005_, new_A6004_, new_A6003_, new_A6002_, new_A6001_, new_A6000_,
    new_A5999_, new_A5998_, new_A5997_, new_A5996_, new_A5995_, new_A5994_,
    new_A5993_, new_A5992_, new_A5991_, new_A5990_, new_A5989_, new_A5988_,
    new_A5987_, new_A5986_, new_A5985_, new_A5984_, new_A5978_, new_A5977_,
    new_A5976_, new_A5975_, new_A5974_, new_A5973_, new_A5972_, new_A5971_,
    new_A5970_, new_A5969_, new_A5968_, new_A5967_, new_A5966_, new_A5965_,
    new_A5964_, new_A5963_, new_A5962_, new_A5961_, new_A5960_, new_A5959_,
    new_A5958_, new_A5957_, new_A5956_, new_A5955_, new_A5954_, new_A5953_,
    new_A5952_, new_A5951_, new_A5945_, new_A5944_, new_A5943_, new_A5942_,
    new_A5941_, new_A5940_, new_A5939_, new_A5938_, new_A5937_, new_A5936_,
    new_A5935_, new_A5934_, new_A5933_, new_A5932_, new_A5931_, new_A5930_,
    new_A5929_, new_A5928_, new_A5927_, new_A5926_, new_A5925_, new_A5924_,
    new_A5923_, new_A5922_, new_A5921_, new_A5920_, new_A5919_, new_A5918_,
    new_A5912_, new_A5911_, new_A5910_, new_A5909_, new_A5908_, new_A5907_,
    new_A5906_, new_A5905_, new_A5904_, new_A5903_, new_A5902_, new_A5901_,
    new_A5900_, new_A5899_, new_A5898_, new_A5897_, new_A5896_, new_A5895_,
    new_A5894_, new_A5893_, new_A5892_, new_A5891_, new_A5890_, new_A5889_,
    new_A5888_, new_A5887_, new_A5886_, new_A5885_, new_A5879_, new_A5878_,
    new_A5877_, new_A5876_, new_A5875_, new_A5874_, new_A5873_, new_A5872_,
    new_A5871_, new_A5870_, new_A5869_, new_A5868_, new_A5867_, new_A5866_,
    new_A5865_, new_A5864_, new_A5863_, new_A5862_, new_A5861_, new_A5860_,
    new_A5859_, new_A5858_, new_A5857_, new_A5856_, new_A5855_, new_A5854_,
    new_A5853_, new_A5852_, new_A5846_, new_A5845_, new_A5844_, new_A5843_,
    new_A5842_, new_A5841_, new_A5840_, new_A5839_, new_A5838_, new_A5837_,
    new_A5836_, new_A5835_, new_A5834_, new_A5833_, new_A5832_, new_A5831_,
    new_A5830_, new_A5829_, new_A5828_, new_A5827_, new_A5826_, new_A5825_,
    new_A5824_, new_A5823_, new_A5822_, new_A5821_, new_A5820_, new_A5819_,
    new_A5813_, new_A5812_, new_A5811_, new_A5810_, new_A5809_, new_A5808_,
    new_A5807_, new_A5806_, new_A5805_, new_A5804_, new_A5803_, new_A5802_,
    new_A5801_, new_A5800_, new_A5799_, new_A5798_, new_A5797_, new_A5796_,
    new_A5795_, new_A5794_, new_A5793_, new_A5792_, new_A5791_, new_A5790_,
    new_A5789_, new_A5788_, new_A5787_, new_A5786_, new_A5780_, new_A5779_,
    new_A5778_, new_A5777_, new_A5776_, new_A5775_, new_A5774_, new_A5773_,
    new_A5772_, new_A5771_, new_A5770_, new_A5769_, new_A5768_, new_A5767_,
    new_A5766_, new_A5765_, new_A5764_, new_A5763_, new_A5762_, new_A5761_,
    new_A5760_, new_A5759_, new_A5758_, new_A5757_, new_A5756_, new_A5755_,
    new_A5754_, new_A5753_, new_A5747_, new_A5746_, new_A5745_, new_A5744_,
    new_A5743_, new_A5742_, new_A5741_, new_A5740_, new_A5739_, new_A5738_,
    new_A5737_, new_A5736_, new_A5735_, new_A5734_, new_A5733_, new_A5732_,
    new_A5731_, new_A5730_, new_A5729_, new_A5728_, new_A5727_, new_A5726_,
    new_A5725_, new_A5724_, new_A5723_, new_A5722_, new_A5721_, new_A5720_,
    new_A5714_, new_A5713_, new_A5712_, new_A5711_, new_A5710_, new_A5709_,
    new_A5708_, new_A5707_, new_A5706_, new_A5705_, new_A5704_, new_A5703_,
    new_A5702_, new_A5701_, new_A5700_, new_A5699_, new_A5698_, new_A5697_,
    new_A5696_, new_A5695_, new_A5694_, new_A5693_, new_A5692_, new_A5691_,
    new_A5690_, new_A5689_, new_A5688_, new_A5687_, new_A5681_, new_A5680_,
    new_A5679_, new_A5678_, new_A5677_, new_A5676_, new_A5675_, new_A5674_,
    new_A5673_, new_A5672_, new_A5671_, new_A5670_, new_A5669_, new_A5668_,
    new_A5667_, new_A5666_, new_A5665_, new_A5664_, new_A5663_, new_A5662_,
    new_A5661_, new_A5660_, new_A5659_, new_A5658_, new_A5657_, new_A5656_,
    new_A5655_, new_A5654_, new_A5648_, new_A5647_, new_A5646_, new_A5645_,
    new_A5644_, new_A5643_, new_A5642_, new_A5641_, new_A5640_, new_A5639_,
    new_A5638_, new_A5637_, new_A5636_, new_A5635_, new_A5634_, new_A5633_,
    new_A5632_, new_A5631_, new_A5630_, new_A5629_, new_A5628_, new_A5627_,
    new_A5626_, new_A5625_, new_A5624_, new_A5623_, new_A5622_, new_A5621_,
    new_A5615_, new_A5614_, new_A5613_, new_A5612_, new_A5611_, new_A5610_,
    new_A5609_, new_A5608_, new_A5607_, new_A5606_, new_A5605_, new_A5604_,
    new_A5603_, new_A5602_, new_A5601_, new_A5600_, new_A5599_, new_A5598_,
    new_A5597_, new_A5596_, new_A5595_, new_A5594_, new_A5593_, new_A5592_,
    new_A5591_, new_A5590_, new_A5589_, new_A5588_, new_A5582_, new_A5581_,
    new_A5580_, new_A5579_, new_A5578_, new_A5577_, new_A5576_, new_A5575_,
    new_A5574_, new_A5573_, new_A5572_, new_A5571_, new_A5570_, new_A5569_,
    new_A5568_, new_A5567_, new_A5566_, new_A5565_, new_A5564_, new_A5563_,
    new_A5562_, new_A5561_, new_A5560_, new_A5559_, new_A5558_, new_A5557_,
    new_A5556_, new_A5555_, new_A5549_, new_A5548_, new_A5547_, new_A5546_,
    new_A5545_, new_A5544_, new_A5543_, new_A5542_, new_A5541_, new_A5540_,
    new_A5539_, new_A5538_, new_A5537_, new_A5536_, new_A5535_, new_A5534_,
    new_A5533_, new_A5532_, new_A5531_, new_A5530_, new_A5529_, new_A5528_,
    new_A5527_, new_A5526_, new_A5525_, new_A5524_, new_A5523_, new_A5522_,
    new_A5516_, new_A5515_, new_A5514_, new_A5513_, new_A5512_, new_A5511_,
    new_A5510_, new_A5509_, new_A5508_, new_A5507_, new_A5506_, new_A5505_,
    new_A5504_, new_A5503_, new_A5502_, new_A5501_, new_A5500_, new_A5499_,
    new_A5498_, new_A5497_, new_A5496_, new_A5495_, new_A5494_, new_A5493_,
    new_A5492_, new_A5491_, new_A5490_, new_A5489_, new_A5483_, new_A5482_,
    new_A5481_, new_A5480_, new_A5479_, new_A5478_, new_A5477_, new_A5476_,
    new_A5475_, new_A5474_, new_A5473_, new_A5472_, new_A5471_, new_A5470_,
    new_A5469_, new_A5468_, new_A5467_, new_A5466_, new_A5465_, new_A5464_,
    new_A5463_, new_A5462_, new_A5461_, new_A5460_, new_A5459_, new_A5458_,
    new_A5457_, new_A5456_, new_A5450_, new_A5449_, new_A5448_, new_A5447_,
    new_A5446_, new_A5445_, new_A5444_, new_A5443_, new_A5442_, new_A5441_,
    new_A5440_, new_A5439_, new_A5438_, new_A5437_, new_A5436_, new_A5435_,
    new_A5434_, new_A5433_, new_A5432_, new_A5431_, new_A5430_, new_A5429_,
    new_A5428_, new_A5427_, new_A5426_, new_A5425_, new_A5424_, new_A5423_,
    new_A5417_, new_A5416_, new_A5415_, new_A5414_, new_A5413_, new_A5412_,
    new_A5411_, new_A5410_, new_A5409_, new_A5408_, new_A5407_, new_A5406_,
    new_A5405_, new_A5404_, new_A5403_, new_A5402_, new_A5401_, new_A5400_,
    new_A5399_, new_A5398_, new_A5397_, new_A5396_, new_A5395_, new_A5394_,
    new_A5393_, new_A5392_, new_A5391_, new_A5390_, new_A5384_, new_A5383_,
    new_A5382_, new_A5381_, new_A5380_, new_A5379_, new_A5378_, new_A5377_,
    new_A5376_, new_A5375_, new_A5374_, new_A5373_, new_A5372_, new_A5371_,
    new_A5370_, new_A5369_, new_A5368_, new_A5367_, new_A5366_, new_A5365_,
    new_A5364_, new_A5363_, new_A5362_, new_A5361_, new_A5360_, new_A5359_,
    new_A5358_, new_A5357_, new_A5351_, new_A5350_, new_A5349_, new_A5348_,
    new_A5347_, new_A5346_, new_A5345_, new_A5344_, new_A5343_, new_A5342_,
    new_A5341_, new_A5340_, new_A5339_, new_A5338_, new_A5337_, new_A5336_,
    new_A5335_, new_A5334_, new_A5333_, new_A5332_, new_A5331_, new_A5330_,
    new_A5329_, new_A5328_, new_A5327_, new_A5326_, new_A5325_, new_A5324_,
    new_A5318_, new_A5317_, new_A5316_, new_A5315_, new_A5314_, new_A5313_,
    new_A5312_, new_A5311_, new_A5310_, new_A5309_, new_A5308_, new_A5307_,
    new_A5306_, new_A5305_, new_A5304_, new_A5303_, new_A5302_, new_A5301_,
    new_A5300_, new_A5299_, new_A5298_, new_A5297_, new_A5296_, new_A5295_,
    new_A5294_, new_A5293_, new_A5292_, new_A5291_, new_A5285_, new_A5284_,
    new_A5283_, new_A5282_, new_A5281_, new_A5280_, new_A5279_, new_A5278_,
    new_A5277_, new_A5276_, new_A5275_, new_A5274_, new_A5273_, new_A5272_,
    new_A5271_, new_A5270_, new_A5269_, new_A5268_, new_A5267_, new_A5266_,
    new_A5265_, new_A5264_, new_A5263_, new_A5262_, new_A5261_, new_A5260_,
    new_A5259_, new_A5258_, new_A5252_, new_A5251_, new_A5250_, new_A5249_,
    new_A5248_, new_A5247_, new_A5246_, new_A5245_, new_A5244_, new_A5243_,
    new_A5242_, new_A5241_, new_A5240_, new_A5239_, new_A5238_, new_A5237_,
    new_A5236_, new_A5235_, new_A5234_, new_A5233_, new_A5232_, new_A5231_,
    new_A5230_, new_A5229_, new_A5228_, new_A5227_, new_A5226_, new_A5225_,
    new_A5219_, new_A5218_, new_A5217_, new_A5216_, new_A5215_, new_A5214_,
    new_A5213_, new_A5212_, new_A5211_, new_A5210_, new_A5209_, new_A5208_,
    new_A5207_, new_A5206_, new_A5205_, new_A5204_, new_A5203_, new_A5202_,
    new_A5201_, new_A5200_, new_A5199_, new_A5198_, new_A5197_, new_A5196_,
    new_A5195_, new_A5194_, new_A5193_, new_A5192_, new_A5186_, new_A5185_,
    new_A5184_, new_A5183_, new_A5182_, new_A5181_, new_A5180_, new_A5179_,
    new_A5178_, new_A5177_, new_A5176_, new_A5175_, new_A5174_, new_A5173_,
    new_A5172_, new_A5171_, new_A5170_, new_A5169_, new_A5168_, new_A5167_,
    new_A5166_, new_A5165_, new_A5164_, new_A5163_, new_A5162_, new_A5161_,
    new_A5160_, new_A5159_, new_A5153_, new_A5152_, new_A5151_, new_A5150_,
    new_A5149_, new_A5148_, new_A5147_, new_A5146_, new_A5145_, new_A5144_,
    new_A5143_, new_A5142_, new_A5141_, new_A5140_, new_A5139_, new_A5138_,
    new_A5137_, new_A5136_, new_A5135_, new_A5134_, new_A5133_, new_A5132_,
    new_A5131_, new_A5130_, new_A5129_, new_A5128_, new_A5127_, new_A5126_,
    new_A5120_, new_A5119_, new_A5118_, new_A5117_, new_A5116_, new_A5115_,
    new_A5114_, new_A5113_, new_A5112_, new_A5111_, new_A5110_, new_A5109_,
    new_A5108_, new_A5107_, new_A5106_, new_A5105_, new_A5104_, new_A5103_,
    new_A5102_, new_A5101_, new_A5100_, new_A5099_, new_A5098_, new_A5097_,
    new_A5096_, new_A5095_, new_A5094_, new_A5093_, new_A5087_, new_A5086_,
    new_A5085_, new_A5084_, new_A5083_, new_A5082_, new_A5081_, new_A5080_,
    new_A5079_, new_A5078_, new_A5077_, new_A5076_, new_A5075_, new_A5074_,
    new_A5073_, new_A5072_, new_A5071_, new_A5070_, new_A5069_, new_A5068_,
    new_A5067_, new_A5066_, new_A5065_, new_A5064_, new_A5063_, new_A5062_,
    new_A5061_, new_A5060_, new_A5054_, new_A5053_, new_A5052_, new_A5051_,
    new_A5050_, new_A5049_, new_A5048_, new_A5047_, new_A5046_, new_A5045_,
    new_A5044_, new_A5043_, new_A5042_, new_A5041_, new_A5040_, new_A5039_,
    new_A5038_, new_A5037_, new_A5036_, new_A5035_, new_A5034_, new_A5033_,
    new_A5032_, new_A5031_, new_A5030_, new_A5029_, new_A5028_, new_A5027_,
    new_A5021_, new_A5020_, new_A5019_, new_A5018_, new_A5017_, new_A5016_,
    new_A5015_, new_A5014_, new_A5013_, new_A5012_, new_A5011_, new_A5010_,
    new_A5009_, new_A5008_, new_A5007_, new_A5006_, new_A5005_, new_A5004_,
    new_A5003_, new_A5002_, new_A5001_, new_A5000_, new_A4999_, new_A4998_,
    new_A4997_, new_A4996_, new_A4995_, new_A4994_, new_A4988_, new_A4987_,
    new_A4986_, new_A4985_, new_A4984_, new_A4983_, new_A4982_, new_A4981_,
    new_A4980_, new_A4979_, new_A4978_, new_A4977_, new_A4976_, new_A4975_,
    new_A4974_, new_A4973_, new_A4972_, new_A4971_, new_A4970_, new_A4969_,
    new_A4968_, new_A4967_, new_A4966_, new_A4965_, new_A4964_, new_A4963_,
    new_A4962_, new_A4961_, new_A4955_, new_A4954_, new_A4953_, new_A4952_,
    new_A4951_, new_A4950_, new_A4949_, new_A4948_, new_A4947_, new_A4946_,
    new_A4945_, new_A4944_, new_A4943_, new_A4942_, new_A4941_, new_A4940_,
    new_A4939_, new_A4938_, new_A4937_, new_A4936_, new_A4935_, new_A4934_,
    new_A4933_, new_A4932_, new_A4931_, new_A4930_, new_A4929_, new_A4928_,
    new_A4922_, new_A4921_, new_A4920_, new_A4919_, new_A4918_, new_A4917_,
    new_A4916_, new_A4915_, new_A4914_, new_A4913_, new_A4912_, new_A4911_,
    new_A4910_, new_A4909_, new_A4908_, new_A4907_, new_A4906_, new_A4905_,
    new_A4904_, new_A4903_, new_A4902_, new_A4901_, new_A4900_, new_A4899_,
    new_A4898_, new_A4897_, new_A4896_, new_A4895_, new_A4889_, new_A4888_,
    new_A4887_, new_A4886_, new_A4885_, new_A4884_, new_A4883_, new_A4882_,
    new_A4881_, new_A4880_, new_A4879_, new_A4878_, new_A4877_, new_A4876_,
    new_A4875_, new_A4874_, new_A4873_, new_A4872_, new_A4871_, new_A4870_,
    new_A4869_, new_A4868_, new_A4867_, new_A4866_, new_A4865_, new_A4864_,
    new_A4863_, new_A4862_, new_A4856_, new_A4855_, new_A4854_, new_A4853_,
    new_A4852_, new_A4851_, new_A4850_, new_A4849_, new_A4848_, new_A4847_,
    new_A4846_, new_A4845_, new_A4844_, new_A4843_, new_A4842_, new_A4841_,
    new_A4840_, new_A4839_, new_A4838_, new_A4837_, new_A4836_, new_A4835_,
    new_A4834_, new_A4833_, new_A4832_, new_A4831_, new_A4830_, new_A4829_,
    new_A4823_, new_A4822_, new_A4821_, new_A4820_, new_A4819_, new_A4818_,
    new_A4817_, new_A4816_, new_A4815_, new_A4814_, new_A4813_, new_A4812_,
    new_A4811_, new_A4810_, new_A4809_, new_A4808_, new_A4807_, new_A4806_,
    new_A4805_, new_A4804_, new_A4803_, new_A4802_, new_A4801_, new_A4800_,
    new_A4799_, new_A4798_, new_A4797_, new_A4796_, new_A4790_, new_A4789_,
    new_A4788_, new_A4787_, new_A4786_, new_A4785_, new_A4784_, new_A4783_,
    new_A4782_, new_A4781_, new_A4780_, new_A4779_, new_A4778_, new_A4777_,
    new_A4776_, new_A4775_, new_A4774_, new_A4773_, new_A4772_, new_A4771_,
    new_A4770_, new_A4769_, new_A4768_, new_A4767_, new_A4766_, new_A4765_,
    new_A4764_, new_A4763_, new_A4757_, new_A4756_, new_A4755_, new_A4754_,
    new_A4753_, new_A4752_, new_A4751_, new_A4750_, new_A4749_, new_A4748_,
    new_A4747_, new_A4746_, new_A4745_, new_A4744_, new_A4743_, new_A4742_,
    new_A4741_, new_A4740_, new_A4739_, new_A4738_, new_A4737_, new_A4736_,
    new_A4735_, new_A4734_, new_A4733_, new_A4732_, new_A4731_, new_A4730_,
    new_A4724_, new_A4723_, new_A4722_, new_A4721_, new_A4720_, new_A4719_,
    new_A4718_, new_A4717_, new_A4716_, new_A4715_, new_A4714_, new_A4713_,
    new_A4712_, new_A4711_, new_A4710_, new_A4709_, new_A4708_, new_A4707_,
    new_A4706_, new_A4705_, new_A4704_, new_A4703_, new_A4702_, new_A4701_,
    new_A4700_, new_A4699_, new_A4698_, new_A4697_, new_A4691_, new_A4690_,
    new_A4689_, new_A4688_, new_A4687_, new_A4686_, new_A4685_, new_A4684_,
    new_A4683_, new_A4682_, new_A4681_, new_A4680_, new_A4679_, new_A4678_,
    new_A4677_, new_A4676_, new_A4675_, new_A4674_, new_A4673_, new_A4672_,
    new_A4671_, new_A4670_, new_A4669_, new_A4668_, new_A4667_, new_A4666_,
    new_A4665_, new_A4664_, new_A4658_, new_A4657_, new_A4656_, new_A4655_,
    new_A4654_, new_A4653_, new_A4652_, new_A4651_, new_A4650_, new_A4649_,
    new_A4648_, new_A4647_, new_A4646_, new_A4645_, new_A4644_, new_A4643_,
    new_A4642_, new_A4641_, new_A4640_, new_A4639_, new_A4638_, new_A4637_,
    new_A4636_, new_A4635_, new_A4634_, new_A4633_, new_A4632_, new_A4631_,
    new_A4625_, new_A4624_, new_A4623_, new_A4622_, new_A4621_, new_A4620_,
    new_A4619_, new_A4618_, new_A4617_, new_A4616_, new_A4615_, new_A4614_,
    new_A4613_, new_A4612_, new_A4611_, new_A4610_, new_A4609_, new_A4608_,
    new_A4607_, new_A4606_, new_A4605_, new_A4604_, new_A4603_, new_A4602_,
    new_A4601_, new_A4600_, new_A4599_, new_A4598_, new_A4592_, new_A4591_,
    new_A4590_, new_A4589_, new_A4588_, new_A4587_, new_A4586_, new_A4585_,
    new_A4584_, new_A4583_, new_A4582_, new_A4581_, new_A4580_, new_A4579_,
    new_A4578_, new_A4577_, new_A4576_, new_A4575_, new_A4574_, new_A4573_,
    new_A4572_, new_A4571_, new_A4570_, new_A4569_, new_A4568_, new_A4567_,
    new_A4566_, new_A4565_, new_A4559_, new_A4558_, new_A4557_, new_A4556_,
    new_A4555_, new_A4554_, new_A4553_, new_A4552_, new_A4551_, new_A4550_,
    new_A4549_, new_A4548_, new_A4547_, new_A4546_, new_A4545_, new_A4544_,
    new_A4543_, new_A4542_, new_A4541_, new_A4540_, new_A4539_, new_A4538_,
    new_A4537_, new_A4536_, new_A4535_, new_A4534_, new_A4533_, new_A4532_,
    new_A4526_, new_A4525_, new_A4524_, new_A4523_, new_A4522_, new_A4521_,
    new_A4520_, new_A4519_, new_A4518_, new_A4517_, new_A4516_, new_A4515_,
    new_A4514_, new_A4513_, new_A4512_, new_A4511_, new_A4510_, new_A4509_,
    new_A4508_, new_A4507_, new_A4506_, new_A4505_, new_A4504_, new_A4503_,
    new_A4502_, new_A4501_, new_A4500_, new_A4499_, new_A4493_, new_A4492_,
    new_A4491_, new_A4490_, new_A4489_, new_A4488_, new_A4487_, new_A4486_,
    new_A4485_, new_A4484_, new_A4483_, new_A4482_, new_A4481_, new_A4480_,
    new_A4479_, new_A4478_, new_A4477_, new_A4476_, new_A4475_, new_A4474_,
    new_A4473_, new_A4472_, new_A4471_, new_A4470_, new_A4469_, new_A4468_,
    new_A4467_, new_A4466_, new_A4460_, new_A4459_, new_A4458_, new_A4457_,
    new_A4456_, new_A4455_, new_A4454_, new_A4453_, new_A4452_, new_A4451_,
    new_A4450_, new_A4449_, new_A4448_, new_A4447_, new_A4446_, new_A4445_,
    new_A4444_, new_A4443_, new_A4442_, new_A4441_, new_A4440_, new_A4439_,
    new_A4438_, new_A4437_, new_A4436_, new_A4435_, new_A4434_, new_A4433_,
    new_A4427_, new_A4426_, new_A4425_, new_A4424_, new_A4423_, new_A4422_,
    new_A4421_, new_A4420_, new_A4419_, new_A4418_, new_A4417_, new_A4416_,
    new_A4415_, new_A4414_, new_A4413_, new_A4412_, new_A4411_, new_A4410_,
    new_A4409_, new_A4408_, new_A4407_, new_A4406_, new_A4405_, new_A4404_,
    new_A4403_, new_A4402_, new_A4401_, new_A4400_, new_A4394_, new_A4393_,
    new_A4392_, new_A4391_, new_A4390_, new_A4389_, new_A4388_, new_A4387_,
    new_A4386_, new_A4385_, new_A4384_, new_A4383_, new_A4382_, new_A4381_,
    new_A4380_, new_A4379_, new_A4378_, new_A4377_, new_A4376_, new_A4375_,
    new_A4374_, new_A4373_, new_A4372_, new_A4371_, new_A4370_, new_A4369_,
    new_A4368_, new_A4367_, new_A4361_, new_A4360_, new_A4359_, new_A4358_,
    new_A4357_, new_A4356_, new_A4355_, new_A4354_, new_A4353_, new_A4352_,
    new_A4351_, new_A4350_, new_A4349_, new_A4348_, new_A4347_, new_A4346_,
    new_A4345_, new_A4344_, new_A4343_, new_A4342_, new_A4341_, new_A4340_,
    new_A4339_, new_A4338_, new_A4337_, new_A4336_, new_A4335_, new_A4334_,
    new_A4328_, new_A4327_, new_A4326_, new_A4325_, new_A4324_, new_A4323_,
    new_A4322_, new_A4321_, new_A4320_, new_A4319_, new_A4318_, new_A4317_,
    new_A4316_, new_A4315_, new_A4314_, new_A4313_, new_A4312_, new_A4311_,
    new_A4310_, new_A4309_, new_A4308_, new_A4307_, new_A4306_, new_A4305_,
    new_A4304_, new_A4303_, new_A4302_, new_A4301_, new_A4295_, new_A4294_,
    new_A4293_, new_A4292_, new_A4291_, new_A4290_, new_A4289_, new_A4288_,
    new_A4287_, new_A4286_, new_A4285_, new_A4284_, new_A4283_, new_A4282_,
    new_A4281_, new_A4280_, new_A4279_, new_A4278_, new_A4277_, new_A4276_,
    new_A4275_, new_A4274_, new_A4273_, new_A4272_, new_A4271_, new_A4270_,
    new_A4269_, new_A4268_, new_A4262_, new_A4261_, new_A4260_, new_A4259_,
    new_A4258_, new_A4257_, new_A4256_, new_A4255_, new_A4254_, new_A4253_,
    new_A4252_, new_A4251_, new_A4250_, new_A4249_, new_A4248_, new_A4247_,
    new_A4246_, new_A4245_, new_A4244_, new_A4243_, new_A4242_, new_A4241_,
    new_A4240_, new_A4239_, new_A4238_, new_A4237_, new_A4236_, new_A4235_,
    new_A4229_, new_A4228_, new_A4227_, new_A4226_, new_A4225_, new_A4224_,
    new_A4223_, new_A4222_, new_A4221_, new_A4220_, new_A4219_, new_A4218_,
    new_A4217_, new_A4216_, new_A4215_, new_A4214_, new_A4213_, new_A4212_,
    new_A4211_, new_A4210_, new_A4209_, new_A4208_, new_A4207_, new_A4206_,
    new_A4205_, new_A4204_, new_A4203_, new_A4202_, new_A4196_, new_A4195_,
    new_A4194_, new_A4193_, new_A4192_, new_A4191_, new_A4190_, new_A4189_,
    new_A4188_, new_A4187_, new_A4186_, new_A4185_, new_A4184_, new_A4183_,
    new_A4182_, new_A4181_, new_A4180_, new_A4179_, new_A4178_, new_A4177_,
    new_A4176_, new_A4175_, new_A4174_, new_A4173_, new_A4172_, new_A4171_,
    new_A4170_, new_A4169_, new_A4163_, new_A4162_, new_A4161_, new_A4160_,
    new_A4159_, new_A4158_, new_A4157_, new_A4156_, new_A4155_, new_A4154_,
    new_A4153_, new_A4152_, new_A4151_, new_A4150_, new_A4149_, new_A4148_,
    new_A4147_, new_A4146_, new_A4145_, new_A4144_, new_A4143_, new_A4142_,
    new_A4141_, new_A4140_, new_A4139_, new_A4138_, new_A4137_, new_A4136_,
    new_A4130_, new_A4129_, new_A4128_, new_A4127_, new_A4126_, new_A4125_,
    new_A4124_, new_A4123_, new_A4122_, new_A4121_, new_A4120_, new_A4119_,
    new_A4118_, new_A4117_, new_A4116_, new_A4115_, new_A4114_, new_A4113_,
    new_A4112_, new_A4111_, new_A4110_, new_A4109_, new_A4108_, new_A4107_,
    new_A4106_, new_A4105_, new_A4104_, new_A4103_, new_A4097_, new_A4096_,
    new_A4095_, new_A4094_, new_A4093_, new_A4092_, new_A4091_, new_A4090_,
    new_A4089_, new_A4088_, new_A4087_, new_A4086_, new_A4085_, new_A4084_,
    new_A4083_, new_A4082_, new_A4081_, new_A4080_, new_A4079_, new_A4078_,
    new_A4077_, new_A4076_, new_A4075_, new_A4074_, new_A4073_, new_A4072_,
    new_A4071_, new_A4070_, new_A4064_, new_A4063_, new_A4062_, new_A4061_,
    new_A4060_, new_A4059_, new_A4058_, new_A4057_, new_A4056_, new_A4055_,
    new_A4054_, new_A4053_, new_A4052_, new_A4051_, new_A4050_, new_A4049_,
    new_A4048_, new_A4047_, new_A4046_, new_A4045_, new_A4044_, new_A4043_,
    new_A4042_, new_A4041_, new_A4040_, new_A4039_, new_A4038_, new_A4037_,
    new_A4031_, new_A4030_, new_A4029_, new_A4028_, new_A4027_, new_A4026_,
    new_A4025_, new_A4024_, new_A4023_, new_A4022_, new_A4021_, new_A4020_,
    new_A4019_, new_A4018_, new_A4017_, new_A4016_, new_A4015_, new_A4014_,
    new_A4013_, new_A4012_, new_A4011_, new_A4010_, new_A4009_, new_A4008_,
    new_A4007_, new_A4006_, new_A4005_, new_A4004_, new_A3998_, new_A3997_,
    new_A3996_, new_A3995_, new_A3994_, new_A3993_, new_A3992_, new_A3991_,
    new_A3990_, new_A3989_, new_A3988_, new_A3987_, new_A3986_, new_A3985_,
    new_A3984_, new_A3983_, new_A3982_, new_A3981_, new_A3980_, new_A3979_,
    new_A3978_, new_A3977_, new_A3976_, new_A3975_, new_A3974_, new_A3973_,
    new_A3972_, new_A3971_, new_A3965_, new_A3964_, new_A3963_, new_A3962_,
    new_A3961_, new_A3960_, new_A3959_, new_A3958_, new_A3957_, new_A3956_,
    new_A3955_, new_A3954_, new_A3953_, new_A3952_, new_A3951_, new_A3950_,
    new_A3949_, new_A3948_, new_A3947_, new_A3946_, new_A3945_, new_A3944_,
    new_A3943_, new_A3942_, new_A3941_, new_A3940_, new_A3939_, new_A3938_,
    new_A3932_, new_A3931_, new_A3930_, new_A3929_, new_A3928_, new_A3927_,
    new_A3926_, new_A3925_, new_A3924_, new_A3923_, new_A3922_, new_A3921_,
    new_A3920_, new_A3919_, new_A3918_, new_A3917_, new_A3916_, new_A3915_,
    new_A3914_, new_A3913_, new_A3912_, new_A3911_, new_A3910_, new_A3909_,
    new_A3908_, new_A3907_, new_A3906_, new_A3905_, new_A3899_, new_A3898_,
    new_A3897_, new_A3896_, new_A3895_, new_A3894_, new_A3893_, new_A3892_,
    new_A3891_, new_A3890_, new_A3889_, new_A3888_, new_A3887_, new_A3886_,
    new_A3885_, new_A3884_, new_A3883_, new_A3882_, new_A3881_, new_A3880_,
    new_A3879_, new_A3878_, new_A3877_, new_A3876_, new_A3875_, new_A3874_,
    new_A3873_, new_A3872_, new_A3866_, new_A3865_, new_A3864_, new_A3863_,
    new_A3862_, new_A3861_, new_A3860_, new_A3859_, new_A3858_, new_A3857_,
    new_A3856_, new_A3855_, new_A3854_, new_A3853_, new_A3852_, new_A3851_,
    new_A3850_, new_A3849_, new_A3848_, new_A3847_, new_A3846_, new_A3845_,
    new_A3844_, new_A3843_, new_A3842_, new_A3841_, new_A3840_, new_A3839_,
    new_A3833_, new_A3832_, new_A3831_, new_A3830_, new_A3829_, new_A3828_,
    new_A3827_, new_A3826_, new_A3825_, new_A3824_, new_A3823_, new_A3822_,
    new_A3821_, new_A3820_, new_A3819_, new_A3818_, new_A3817_, new_A3816_,
    new_A3815_, new_A3814_, new_A3813_, new_A3812_, new_A3811_, new_A3810_,
    new_A3809_, new_A3808_, new_A3807_, new_A3806_, new_A3800_, new_A3799_,
    new_A3798_, new_A3797_, new_A3796_, new_A3795_, new_A3794_, new_A3793_,
    new_A3792_, new_A3791_, new_A3790_, new_A3789_, new_A3788_, new_A3787_,
    new_A3786_, new_A3785_, new_A3784_, new_A3783_, new_A3782_, new_A3781_,
    new_A3780_, new_A3779_, new_A3778_, new_A3777_, new_A3776_, new_A3775_,
    new_A3774_, new_A3773_, new_A3767_, new_A3766_, new_A3765_, new_A3764_,
    new_A3763_, new_A3762_, new_A3761_, new_A3760_, new_A3759_, new_A3758_,
    new_A3757_, new_A3756_, new_A3755_, new_A3754_, new_A3753_, new_A3752_,
    new_A3751_, new_A3750_, new_A3749_, new_A3748_, new_A3747_, new_A3746_,
    new_A3745_, new_A3744_, new_A3743_, new_A3742_, new_A3741_, new_A3740_,
    new_A3734_, new_A3733_, new_A3732_, new_A3731_, new_A3730_, new_A3729_,
    new_A3728_, new_A3727_, new_A3726_, new_A3725_, new_A3724_, new_A3723_,
    new_A3722_, new_A3721_, new_A3720_, new_A3719_, new_A3718_, new_A3717_,
    new_A3716_, new_A3715_, new_A3714_, new_A3713_, new_A3712_, new_A3711_,
    new_A3710_, new_A3709_, new_A3708_, new_A3707_, new_A3701_, new_A3700_,
    new_A3699_, new_A3698_, new_A3697_, new_A3696_, new_A3695_, new_A3694_,
    new_A3693_, new_A3692_, new_A3691_, new_A3690_, new_A3689_, new_A3688_,
    new_A3687_, new_A3686_, new_A3685_, new_A3684_, new_A3683_, new_A3682_,
    new_A3681_, new_A3680_, new_A3679_, new_A3678_, new_A3677_, new_A3676_,
    new_A3675_, new_A3674_, new_A3668_, new_A3667_, new_A3666_, new_A3665_,
    new_A3664_, new_A3663_, new_A3662_, new_A3661_, new_A3660_, new_A3659_,
    new_A3658_, new_A3657_, new_A3656_, new_A3655_, new_A3654_, new_A3653_,
    new_A3652_, new_A3651_, new_A3650_, new_A3649_, new_A3648_, new_A3647_,
    new_A3646_, new_A3645_, new_A3644_, new_A3643_, new_A3642_, new_A3641_,
    new_A3635_, new_A3634_, new_A3633_, new_A3632_, new_A3631_, new_A3630_,
    new_A3629_, new_A3628_, new_A3627_, new_A3626_, new_A3625_, new_A3624_,
    new_A3623_, new_A3622_, new_A3621_, new_A3620_, new_A3619_, new_A3618_,
    new_A3617_, new_A3616_, new_A3615_, new_A3614_, new_A3613_, new_A3612_,
    new_A3611_, new_A3610_, new_A3609_, new_A3608_, new_A3602_, new_A3601_,
    new_A3600_, new_A3599_, new_A3598_, new_A3597_, new_A3596_, new_A3595_,
    new_A3594_, new_A3593_, new_A3592_, new_A3591_, new_A3590_, new_A3589_,
    new_A3588_, new_A3587_, new_A3586_, new_A3585_, new_A3584_, new_A3583_,
    new_A3582_, new_A3581_, new_A3580_, new_A3579_, new_A3578_, new_A3577_,
    new_A3576_, new_A3575_, new_A3569_, new_A3568_, new_A3567_, new_A3566_,
    new_A3565_, new_A3564_, new_A3563_, new_A3562_, new_A3561_, new_A3560_,
    new_A3559_, new_A3558_, new_A3557_, new_A3556_, new_A3555_, new_A3554_,
    new_A3553_, new_A3552_, new_A3551_, new_A3550_, new_A3549_, new_A3548_,
    new_A3547_, new_A3546_, new_A3545_, new_A3544_, new_A3543_, new_A3542_,
    new_A3536_, new_A3535_, new_A3534_, new_A3533_, new_A3532_, new_A3531_,
    new_A3530_, new_A3529_, new_A3528_, new_A3527_, new_A3526_, new_A3525_,
    new_A3524_, new_A3523_, new_A3522_, new_A3521_, new_A3520_, new_A3519_,
    new_A3518_, new_A3517_, new_A3516_, new_A3515_, new_A3514_, new_A3513_,
    new_A3512_, new_A3511_, new_A3510_, new_A3509_, new_A3503_, new_A3502_,
    new_A3501_, new_A3500_, new_A3499_, new_A3498_, new_A3497_, new_A3496_,
    new_A3495_, new_A3494_, new_A3493_, new_A3492_, new_A3491_, new_A3490_,
    new_A3489_, new_A3488_, new_A3487_, new_A3486_, new_A3485_, new_A3484_,
    new_A3483_, new_A3482_, new_A3481_, new_A3480_, new_A3479_, new_A3478_,
    new_A3477_, new_A3476_, new_A3470_, new_A3469_, new_A3468_, new_A3467_,
    new_A3466_, new_A3465_, new_A3464_, new_A3463_, new_A3462_, new_A3461_,
    new_A3460_, new_A3459_, new_A3458_, new_A3457_, new_A3456_, new_A3455_,
    new_A3454_, new_A3453_, new_A3452_, new_A3451_, new_A3450_, new_A3449_,
    new_A3448_, new_A3447_, new_A3446_, new_A3445_, new_A3444_, new_A3443_,
    new_A3437_, new_A3436_, new_A3435_, new_A3434_, new_A3433_, new_A3432_,
    new_A3431_, new_A3430_, new_A3429_, new_A3428_, new_A3427_, new_A3426_,
    new_A3425_, new_A3424_, new_A3423_, new_A3422_, new_A3421_, new_A3420_,
    new_A3419_, new_A3418_, new_A3417_, new_A3416_, new_A3415_, new_A3414_,
    new_A3413_, new_A3412_, new_A3411_, new_A3410_, new_A3404_, new_A3403_,
    new_A3402_, new_A3401_, new_A3400_, new_A3399_, new_A3398_, new_A3397_,
    new_A3396_, new_A3395_, new_A3394_, new_A3393_, new_A3392_, new_A3391_,
    new_A3390_, new_A3389_, new_A3388_, new_A3387_, new_A3386_, new_A3385_,
    new_A3384_, new_A3383_, new_A3382_, new_A3381_, new_A3380_, new_A3379_,
    new_A3378_, new_A3377_, new_A3371_, new_A3370_, new_A3369_, new_A3368_,
    new_A3367_, new_A3366_, new_A3365_, new_A3364_, new_A3363_, new_A3362_,
    new_A3361_, new_A3360_, new_A3359_, new_A3358_, new_A3357_, new_A3356_,
    new_A3355_, new_A3354_, new_A3353_, new_A3352_, new_A3351_, new_A3350_,
    new_A3349_, new_A3348_, new_A3347_, new_A3346_, new_A3345_, new_A3344_,
    new_A3338_, new_A3337_, new_A3336_, new_A3335_, new_A3334_, new_A3333_,
    new_A3332_, new_A3331_, new_A3330_, new_A3329_, new_A3328_, new_A3327_,
    new_A3326_, new_A3325_, new_A3324_, new_A3323_, new_A3322_, new_A3321_,
    new_A3320_, new_A3319_, new_A3318_, new_A3317_, new_A3316_, new_A3315_,
    new_A3314_, new_A3313_, new_A3312_, new_A3311_, new_A3305_, new_A3304_,
    new_A3303_, new_A3302_, new_A3301_, new_A3300_, new_A3299_, new_A3298_,
    new_A3297_, new_A3296_, new_A3295_, new_A3294_, new_A3293_, new_A3292_,
    new_A3291_, new_A3290_, new_A3289_, new_A3288_, new_A3287_, new_A3286_,
    new_A3285_, new_A3284_, new_A3283_, new_A3282_, new_A3281_, new_A3280_,
    new_A3279_, new_A3278_, new_A3272_, new_A3271_, new_A3270_, new_A3269_,
    new_A3268_, new_A3267_, new_A3266_, new_A3265_, new_A3264_, new_A3263_,
    new_A3262_, new_A3261_, new_A3260_, new_A3259_, new_A3258_, new_A3257_,
    new_A3256_, new_A3255_, new_A3254_, new_A3253_, new_A3252_, new_A3251_,
    new_A3250_, new_A3249_, new_A3248_, new_A3247_, new_A3246_, new_A3245_,
    new_A3239_, new_A3238_, new_A3237_, new_A3236_, new_A3235_, new_A3234_,
    new_A3233_, new_A3232_, new_A3231_, new_A3230_, new_A3229_, new_A3228_,
    new_A3227_, new_A3226_, new_A3225_, new_A3224_, new_A3223_, new_A3222_,
    new_A3221_, new_A3220_, new_A3219_, new_A3218_, new_A3217_, new_A3216_,
    new_A3215_, new_A3214_, new_A3213_, new_A3212_, new_A3206_, new_A3205_,
    new_A3204_, new_A3203_, new_A3202_, new_A3201_, new_A3200_, new_A3199_,
    new_A3198_, new_A3197_, new_A3196_, new_A3195_, new_A3194_, new_A3193_,
    new_A3192_, new_A3191_, new_A3190_, new_A3189_, new_A3188_, new_A3187_,
    new_A3186_, new_A3185_, new_A3184_, new_A3183_, new_A3182_, new_A3181_,
    new_A3180_, new_A3179_, new_A3173_, new_A3172_, new_A3171_, new_A3170_,
    new_A3169_, new_A3168_, new_A3167_, new_A3166_, new_A3165_, new_A3164_,
    new_A3163_, new_A3162_, new_A3161_, new_A3160_, new_A3159_, new_A3158_,
    new_A3157_, new_A3156_, new_A3155_, new_A3154_, new_A3153_, new_A3152_,
    new_A3151_, new_A3150_, new_A3149_, new_A3148_, new_A3147_, new_A3146_,
    new_A3140_, new_A3139_, new_A3138_, new_A3137_, new_A3136_, new_A3135_,
    new_A3134_, new_A3133_, new_A3132_, new_A3131_, new_A3130_, new_A3129_,
    new_A3128_, new_A3127_, new_A3126_, new_A3125_, new_A3124_, new_A3123_,
    new_A3122_, new_A3121_, new_A3120_, new_A3119_, new_A3118_, new_A3117_,
    new_A3116_, new_A3115_, new_A3114_, new_A3113_, new_A3107_, new_A3106_,
    new_A3105_, new_A3104_, new_A3103_, new_A3102_, new_A3101_, new_A3100_,
    new_A3099_, new_A3098_, new_A3097_, new_A3096_, new_A3095_, new_A3094_,
    new_A3093_, new_A3092_, new_A3091_, new_A3090_, new_A3089_, new_A3088_,
    new_A3087_, new_A3086_, new_A3085_, new_A3084_, new_A3083_, new_A3082_,
    new_A3081_, new_A3080_, new_A3074_, new_A3073_, new_A3072_, new_A3071_,
    new_A3070_, new_A3069_, new_A3068_, new_A3067_, new_A3066_, new_A3065_,
    new_A3064_, new_A3063_, new_A3062_, new_A3061_, new_A3060_, new_A3059_,
    new_A3058_, new_A3057_, new_A3056_, new_A3055_, new_A3054_, new_A3053_,
    new_A3052_, new_A3051_, new_A3050_, new_A3049_, new_A3048_, new_A3047_,
    new_A3041_, new_A3040_, new_A3039_, new_A3038_, new_A3037_, new_A3036_,
    new_A3035_, new_A3034_, new_A3033_, new_A3032_, new_A3031_, new_A3030_,
    new_A3029_, new_A3028_, new_A3027_, new_A3026_, new_A3025_, new_A3024_,
    new_A3023_, new_A3022_, new_A3021_, new_A3020_, new_A3019_, new_A3018_,
    new_A3017_, new_A3016_, new_A3015_, new_A3014_, new_A3008_, new_A3007_,
    new_A3006_, new_A3005_, new_A3004_, new_A3003_, new_A3002_, new_A3001_,
    new_A3000_, new_A2999_, new_A2998_, new_A2997_, new_A2996_, new_A2995_,
    new_A2994_, new_A2993_, new_A2992_, new_A2991_, new_A2990_, new_A2989_,
    new_A2988_, new_A2987_, new_A2986_, new_A2985_, new_A2984_, new_A2983_,
    new_A2982_, new_A2981_, new_A2975_, new_A2974_, new_A2973_, new_A2972_,
    new_A2971_, new_A2970_, new_A2969_, new_A2968_, new_A2967_, new_A2966_,
    new_A2965_, new_A2964_, new_A2963_, new_A2962_, new_A2961_, new_A2960_,
    new_A2959_, new_A2958_, new_A2957_, new_A2956_, new_A2955_, new_A2954_,
    new_A2953_, new_A2952_, new_A2951_, new_A2950_, new_A2949_, new_A2948_,
    new_A2942_, new_A2941_, new_A2940_, new_A2939_, new_A2938_, new_A2937_,
    new_A2936_, new_A2935_, new_A2934_, new_A2933_, new_A2932_, new_A2931_,
    new_A2930_, new_A2929_, new_A2928_, new_A2927_, new_A2926_, new_A2925_,
    new_A2924_, new_A2923_, new_A2922_, new_A2921_, new_A2920_, new_A2919_,
    new_A2918_, new_A2917_, new_A2916_, new_A2915_, new_A2909_, new_A2908_,
    new_A2907_, new_A2906_, new_A2905_, new_A2904_, new_A2903_, new_A2902_,
    new_A2901_, new_A2900_, new_A2899_, new_A2898_, new_A2897_, new_A2896_,
    new_A2895_, new_A2894_, new_A2893_, new_A2892_, new_A2891_, new_A2890_,
    new_A2889_, new_A2888_, new_A2887_, new_A2886_, new_A2885_, new_A2884_,
    new_A2883_, new_A2882_, new_A2876_, new_A2875_, new_A2874_, new_A2873_,
    new_A2872_, new_A2871_, new_A2870_, new_A2869_, new_A2868_, new_A2867_,
    new_A2866_, new_A2865_, new_A2864_, new_A2863_, new_A2862_, new_A2861_,
    new_A2860_, new_A2859_, new_A2858_, new_A2857_, new_A2856_, new_A2855_,
    new_A2854_, new_A2853_, new_A2852_, new_A2851_, new_A2850_, new_A2849_,
    new_A2843_, new_A2842_, new_A2841_, new_A2840_, new_A2839_, new_A2806_,
    new_A2807_, new_A2808_, new_A2809_, new_A2810_, new_A2816_, new_A2817_,
    new_A2818_, new_A2819_, new_A2820_, new_A2821_, new_A2822_, new_A2823_,
    new_A2824_, new_A2825_, new_A2826_, new_A2827_, new_A2828_, new_A2829_,
    new_A2830_, new_A2831_, new_A2832_, new_A2833_, new_A2834_, new_A2835_,
    new_A2836_, new_A2837_, new_A2838_;
  assign new_B5214_ = new_B5192_ & new_B5207_;
  assign new_B5213_ = ~new_B5192_ & ~new_B5214_;
  assign new_B5212_ = new_B5192_ | new_B5207_;
  assign new_B5211_ = ~B5185 | ~B5186;
  assign new_B5210_ = new_B5192_ | new_B5207_;
  assign new_B5209_ = ~new_B5208_ & ~new_B5192_;
  assign new_B5208_ = new_B5192_ & new_B5207_;
  assign new_B5207_ = ~B5183 | ~B5184;
  assign new_B5206_ = B5184 & new_B5196_;
  assign new_B5205_ = B5185 | new_B5192_;
  assign new_B5204_ = B5185 | B5186;
  assign new_B5203_ = ~new_B5213_ | ~new_B5212_;
  assign new_B5202_ = new_B5211_ & new_B5204_;
  assign new_B5201_ = B5185 ^ new_B5192_;
  assign new_B5200_ = ~new_B5209_ | ~new_B5210_;
  assign new_B5199_ = ~B5184 ^ new_B5196_;
  assign new_B5198_ = new_B5206_ | B5183;
  assign new_B5197_ = new_B5203_ & B5184;
  assign new_B5196_ = new_B5205_ & new_B5204_;
  assign new_B5195_ = new_B5200_ & B5184;
  assign new_B5194_ = new_B5202_ & new_B5201_;
  assign new_B5193_ = new_B5194_ ^ B5184;
  assign new_B5192_ = B5182 ^ B5183;
  assign new_B5191_ = new_B5192_ & new_B5199_;
  assign new_B5190_ = new_B5192_ & new_B5198_;
  assign new_B5189_ = new_B5197_ | new_B5196_;
  assign new_B5188_ = new_B5195_ | new_B5194_;
  assign new_B5187_ = new_B5193_ & new_B5192_;
  assign new_B5220_ = new_B5226_ & new_B5225_;
  assign new_B5221_ = new_B5228_ | new_B5227_;
  assign new_B5222_ = new_B5230_ | new_B5229_;
  assign new_B5223_ = new_B5225_ & new_B5231_;
  assign new_B5224_ = new_B5225_ & new_B5232_;
  assign new_B5225_ = B5215 ^ B5216;
  assign new_B5226_ = new_B5227_ ^ B5217;
  assign new_B5227_ = new_B5235_ & new_B5234_;
  assign new_B5228_ = new_B5233_ & B5217;
  assign new_B5229_ = new_B5238_ & new_B5237_;
  assign new_B5230_ = new_B5236_ & B5217;
  assign new_B5231_ = new_B5239_ | B5216;
  assign new_B5232_ = ~B5217 ^ new_B5229_;
  assign new_B5233_ = ~new_B5242_ | ~new_B5243_;
  assign new_B5234_ = B5218 ^ new_B5225_;
  assign new_B5235_ = new_B5244_ & new_B5237_;
  assign new_B5236_ = ~new_B5246_ | ~new_B5245_;
  assign new_B5237_ = B5218 | B5219;
  assign new_B5238_ = B5218 | new_B5225_;
  assign new_B5239_ = B5217 & new_B5229_;
  assign new_B5240_ = ~B5216 | ~B5217;
  assign new_B5241_ = new_B5225_ & new_B5240_;
  assign new_B5242_ = ~new_B5241_ & ~new_B5225_;
  assign new_B5243_ = new_B5225_ | new_B5240_;
  assign new_B5244_ = ~B5218 | ~B5219;
  assign new_B5245_ = new_B5225_ | new_B5240_;
  assign new_B5246_ = ~new_B5225_ & ~new_B5247_;
  assign new_B5247_ = new_B5225_ & new_B5240_;
  assign new_B5253_ = new_B5259_ & new_B5258_;
  assign new_B5254_ = new_B5261_ | new_B5260_;
  assign new_B5255_ = new_B5263_ | new_B5262_;
  assign new_B5256_ = new_B5258_ & new_B5264_;
  assign new_B5257_ = new_B5258_ & new_B5265_;
  assign new_B5258_ = B5248 ^ B5249;
  assign new_B5259_ = new_B5260_ ^ B5250;
  assign new_B5260_ = new_B5268_ & new_B5267_;
  assign new_B5261_ = new_B5266_ & B5250;
  assign new_B5262_ = new_B5271_ & new_B5270_;
  assign new_B5263_ = new_B5269_ & B5250;
  assign new_B5264_ = new_B5272_ | B5249;
  assign new_B5265_ = ~B5250 ^ new_B5262_;
  assign new_B5266_ = ~new_B5275_ | ~new_B5276_;
  assign new_B5267_ = B5251 ^ new_B5258_;
  assign new_B5268_ = new_B5277_ & new_B5270_;
  assign new_B5269_ = ~new_B5279_ | ~new_B5278_;
  assign new_B5270_ = B5251 | B5252;
  assign new_B5271_ = B5251 | new_B5258_;
  assign new_B5272_ = B5250 & new_B5262_;
  assign new_B5273_ = ~B5249 | ~B5250;
  assign new_B5274_ = new_B5258_ & new_B5273_;
  assign new_B5275_ = ~new_B5274_ & ~new_B5258_;
  assign new_B5276_ = new_B5258_ | new_B5273_;
  assign new_B5277_ = ~B5251 | ~B5252;
  assign new_B5278_ = new_B5258_ | new_B5273_;
  assign new_B5279_ = ~new_B5258_ & ~new_B5280_;
  assign new_B5280_ = new_B5258_ & new_B5273_;
  assign new_B5286_ = new_B5292_ & new_B5291_;
  assign new_B5287_ = new_B5294_ | new_B5293_;
  assign new_B5288_ = new_B5296_ | new_B5295_;
  assign new_B5289_ = new_B5291_ & new_B5297_;
  assign new_B5290_ = new_B5291_ & new_B5298_;
  assign new_B5291_ = B5281 ^ B5282;
  assign new_B5292_ = new_B5293_ ^ B5283;
  assign new_B5293_ = new_B5301_ & new_B5300_;
  assign new_B5294_ = new_B5299_ & B5283;
  assign new_B5295_ = new_B5304_ & new_B5303_;
  assign new_B5296_ = new_B5302_ & B5283;
  assign new_B5297_ = new_B5305_ | B5282;
  assign new_B5298_ = ~B5283 ^ new_B5295_;
  assign new_B5299_ = ~new_B5308_ | ~new_B5309_;
  assign new_B5300_ = B5284 ^ new_B5291_;
  assign new_B5301_ = new_B5310_ & new_B5303_;
  assign new_B5302_ = ~new_B5312_ | ~new_B5311_;
  assign new_B5303_ = B5284 | B5285;
  assign new_B5304_ = B5284 | new_B5291_;
  assign new_B5305_ = B5283 & new_B5295_;
  assign new_B5306_ = ~B5282 | ~B5283;
  assign new_B5307_ = new_B5291_ & new_B5306_;
  assign new_B5308_ = ~new_B5307_ & ~new_B5291_;
  assign new_B5309_ = new_B5291_ | new_B5306_;
  assign new_B5310_ = ~B5284 | ~B5285;
  assign new_B5311_ = new_B5291_ | new_B5306_;
  assign new_B5312_ = ~new_B5291_ & ~new_B5313_;
  assign new_B5313_ = new_B5291_ & new_B5306_;
  assign new_B5319_ = new_B5325_ & new_B5324_;
  assign new_B5320_ = new_B5327_ | new_B5326_;
  assign new_B5321_ = new_B5329_ | new_B5328_;
  assign new_B5322_ = new_B5324_ & new_B5330_;
  assign new_B5323_ = new_B5324_ & new_B5331_;
  assign new_B5324_ = B5314 ^ B5315;
  assign new_B5325_ = new_B5326_ ^ B5316;
  assign new_B5326_ = new_B5334_ & new_B5333_;
  assign new_B5327_ = new_B5332_ & B5316;
  assign new_B5328_ = new_B5337_ & new_B5336_;
  assign new_B5329_ = new_B5335_ & B5316;
  assign new_B5330_ = new_B5338_ | B5315;
  assign new_B5331_ = ~B5316 ^ new_B5328_;
  assign new_B5332_ = ~new_B5341_ | ~new_B5342_;
  assign new_B5333_ = B5317 ^ new_B5324_;
  assign new_B5334_ = new_B5343_ & new_B5336_;
  assign new_B5335_ = ~new_B5345_ | ~new_B5344_;
  assign new_B5336_ = B5317 | B5318;
  assign new_B5337_ = B5317 | new_B5324_;
  assign new_B5338_ = B5316 & new_B5328_;
  assign new_B5339_ = ~B5315 | ~B5316;
  assign new_B5340_ = new_B5324_ & new_B5339_;
  assign new_B5341_ = ~new_B5340_ & ~new_B5324_;
  assign new_B5342_ = new_B5324_ | new_B5339_;
  assign new_B5343_ = ~B5317 | ~B5318;
  assign new_B5344_ = new_B5324_ | new_B5339_;
  assign new_B5345_ = ~new_B5324_ & ~new_B5346_;
  assign new_B5346_ = new_B5324_ & new_B5339_;
  assign new_B5352_ = new_B5358_ & new_B5357_;
  assign new_B5353_ = new_B5360_ | new_B5359_;
  assign new_B5354_ = new_B5362_ | new_B5361_;
  assign new_B5355_ = new_B5357_ & new_B5363_;
  assign new_B5356_ = new_B5357_ & new_B5364_;
  assign new_B5357_ = B5347 ^ B5348;
  assign new_B5358_ = new_B5359_ ^ B5349;
  assign new_B5359_ = new_B5367_ & new_B5366_;
  assign new_B5360_ = new_B5365_ & B5349;
  assign new_B5361_ = new_B5370_ & new_B5369_;
  assign new_B5362_ = new_B5368_ & B5349;
  assign new_B5363_ = new_B5371_ | B5348;
  assign new_B5364_ = ~B5349 ^ new_B5361_;
  assign new_B5365_ = ~new_B5374_ | ~new_B5375_;
  assign new_B5366_ = B5350 ^ new_B5357_;
  assign new_B5367_ = new_B5376_ & new_B5369_;
  assign new_B5368_ = ~new_B5378_ | ~new_B5377_;
  assign new_B5369_ = B5350 | B5351;
  assign new_B5370_ = B5350 | new_B5357_;
  assign new_B5371_ = B5349 & new_B5361_;
  assign new_B5372_ = ~B5348 | ~B5349;
  assign new_B5373_ = new_B5357_ & new_B5372_;
  assign new_B5374_ = ~new_B5373_ & ~new_B5357_;
  assign new_B5375_ = new_B5357_ | new_B5372_;
  assign new_B5376_ = ~B5350 | ~B5351;
  assign new_B5377_ = new_B5357_ | new_B5372_;
  assign new_B5378_ = ~new_B5357_ & ~new_B5379_;
  assign new_B5379_ = new_B5357_ & new_B5372_;
  assign new_B5385_ = new_B5391_ & new_B5390_;
  assign new_B5386_ = new_B5393_ | new_B5392_;
  assign new_B5387_ = new_B5395_ | new_B5394_;
  assign new_B5388_ = new_B5390_ & new_B5396_;
  assign new_B5389_ = new_B5390_ & new_B5397_;
  assign new_B5390_ = B5380 ^ B5381;
  assign new_B5391_ = new_B5392_ ^ B5382;
  assign new_B5392_ = new_B5400_ & new_B5399_;
  assign new_B5393_ = new_B5398_ & B5382;
  assign new_B5394_ = new_B5403_ & new_B5402_;
  assign new_B5395_ = new_B5401_ & B5382;
  assign new_B5396_ = new_B5404_ | B5381;
  assign new_B5397_ = ~B5382 ^ new_B5394_;
  assign new_B5398_ = ~new_B5407_ | ~new_B5408_;
  assign new_B5399_ = B5383 ^ new_B5390_;
  assign new_B5400_ = new_B5409_ & new_B5402_;
  assign new_B5401_ = ~new_B5411_ | ~new_B5410_;
  assign new_B5402_ = B5383 | B5384;
  assign new_B5403_ = B5383 | new_B5390_;
  assign new_B5404_ = B5382 & new_B5394_;
  assign new_B5405_ = ~B5381 | ~B5382;
  assign new_B5406_ = new_B5390_ & new_B5405_;
  assign new_B5407_ = ~new_B5406_ & ~new_B5390_;
  assign new_B5408_ = new_B5390_ | new_B5405_;
  assign new_B5409_ = ~B5383 | ~B5384;
  assign new_B5410_ = new_B5390_ | new_B5405_;
  assign new_B5411_ = ~new_B5390_ & ~new_B5412_;
  assign new_B5412_ = new_B5390_ & new_B5405_;
  assign new_B5418_ = new_B5424_ & new_B5423_;
  assign new_B5419_ = new_B5426_ | new_B5425_;
  assign new_B5420_ = new_B5428_ | new_B5427_;
  assign new_B5421_ = new_B5423_ & new_B5429_;
  assign new_B5422_ = new_B5423_ & new_B5430_;
  assign new_B5423_ = B5413 ^ B5414;
  assign new_B5424_ = new_B5425_ ^ B5415;
  assign new_B5425_ = new_B5433_ & new_B5432_;
  assign new_B5426_ = new_B5431_ & B5415;
  assign new_B5427_ = new_B5436_ & new_B5435_;
  assign new_B5428_ = new_B5434_ & B5415;
  assign new_B5429_ = new_B5437_ | B5414;
  assign new_B5430_ = ~B5415 ^ new_B5427_;
  assign new_B5431_ = ~new_B5440_ | ~new_B5441_;
  assign new_B5432_ = B5416 ^ new_B5423_;
  assign new_B5433_ = new_B5442_ & new_B5435_;
  assign new_B5434_ = ~new_B5444_ | ~new_B5443_;
  assign new_B5435_ = B5416 | B5417;
  assign new_B5436_ = B5416 | new_B5423_;
  assign new_B5437_ = B5415 & new_B5427_;
  assign new_B5438_ = ~B5414 | ~B5415;
  assign new_B5439_ = new_B5423_ & new_B5438_;
  assign new_B5440_ = ~new_B5439_ & ~new_B5423_;
  assign new_B5441_ = new_B5423_ | new_B5438_;
  assign new_B5442_ = ~B5416 | ~B5417;
  assign new_B5443_ = new_B5423_ | new_B5438_;
  assign new_B5444_ = ~new_B5423_ & ~new_B5445_;
  assign new_B5445_ = new_B5423_ & new_B5438_;
  assign new_B5451_ = new_B5457_ & new_B5456_;
  assign new_B5452_ = new_B5459_ | new_B5458_;
  assign new_B5453_ = new_B5461_ | new_B5460_;
  assign new_B5454_ = new_B5456_ & new_B5462_;
  assign new_B5455_ = new_B5456_ & new_B5463_;
  assign new_B5456_ = B5446 ^ B5447;
  assign new_B5457_ = new_B5458_ ^ B5448;
  assign new_B5458_ = new_B5466_ & new_B5465_;
  assign new_B5459_ = new_B5464_ & B5448;
  assign new_B5460_ = new_B5469_ & new_B5468_;
  assign new_B5461_ = new_B5467_ & B5448;
  assign new_B5462_ = new_B5470_ | B5447;
  assign new_B5463_ = ~B5448 ^ new_B5460_;
  assign new_B5464_ = ~new_B5473_ | ~new_B5474_;
  assign new_B5465_ = B5449 ^ new_B5456_;
  assign new_B5466_ = new_B5475_ & new_B5468_;
  assign new_B5467_ = ~new_B5477_ | ~new_B5476_;
  assign new_B5468_ = B5449 | B5450;
  assign new_B5469_ = B5449 | new_B5456_;
  assign new_B5470_ = B5448 & new_B5460_;
  assign new_B5471_ = ~B5447 | ~B5448;
  assign new_B5472_ = new_B5456_ & new_B5471_;
  assign new_B5473_ = ~new_B5472_ & ~new_B5456_;
  assign new_B5474_ = new_B5456_ | new_B5471_;
  assign new_B5475_ = ~B5449 | ~B5450;
  assign new_B5476_ = new_B5456_ | new_B5471_;
  assign new_B5477_ = ~new_B5456_ & ~new_B5478_;
  assign new_B5478_ = new_B5456_ & new_B5471_;
  assign new_B5484_ = new_B5490_ & new_B5489_;
  assign new_B5485_ = new_B5492_ | new_B5491_;
  assign new_B5486_ = new_B5494_ | new_B5493_;
  assign new_B5487_ = new_B5489_ & new_B5495_;
  assign new_B5488_ = new_B5489_ & new_B5496_;
  assign new_B5489_ = B5479 ^ B5480;
  assign new_B5490_ = new_B5491_ ^ B5481;
  assign new_B5491_ = new_B5499_ & new_B5498_;
  assign new_B5492_ = new_B5497_ & B5481;
  assign new_B5493_ = new_B5502_ & new_B5501_;
  assign new_B5494_ = new_B5500_ & B5481;
  assign new_B5495_ = new_B5503_ | B5480;
  assign new_B5496_ = ~B5481 ^ new_B5493_;
  assign new_B5497_ = ~new_B5506_ | ~new_B5507_;
  assign new_B5498_ = B5482 ^ new_B5489_;
  assign new_B5499_ = new_B5508_ & new_B5501_;
  assign new_B5500_ = ~new_B5510_ | ~new_B5509_;
  assign new_B5501_ = B5482 | B5483;
  assign new_B5502_ = B5482 | new_B5489_;
  assign new_B5503_ = B5481 & new_B5493_;
  assign new_B5504_ = ~B5480 | ~B5481;
  assign new_B5505_ = new_B5489_ & new_B5504_;
  assign new_B5506_ = ~new_B5505_ & ~new_B5489_;
  assign new_B5507_ = new_B5489_ | new_B5504_;
  assign new_B5508_ = ~B5482 | ~B5483;
  assign new_B5509_ = new_B5489_ | new_B5504_;
  assign new_B5510_ = ~new_B5489_ & ~new_B5511_;
  assign new_B5511_ = new_B5489_ & new_B5504_;
  assign new_B5517_ = new_B5523_ & new_B5522_;
  assign new_B5518_ = new_B5525_ | new_B5524_;
  assign new_B5519_ = new_B5527_ | new_B5526_;
  assign new_B5520_ = new_B5522_ & new_B5528_;
  assign new_B5521_ = new_B5522_ & new_B5529_;
  assign new_B5522_ = B5512 ^ B5513;
  assign new_B5523_ = new_B5524_ ^ B5514;
  assign new_B5524_ = new_B5532_ & new_B5531_;
  assign new_B5525_ = new_B5530_ & B5514;
  assign new_B5526_ = new_B5535_ & new_B5534_;
  assign new_B5527_ = new_B5533_ & B5514;
  assign new_B5528_ = new_B5536_ | B5513;
  assign new_B5529_ = ~B5514 ^ new_B5526_;
  assign new_B5530_ = ~new_B5539_ | ~new_B5540_;
  assign new_B5531_ = B5515 ^ new_B5522_;
  assign new_B5532_ = new_B5541_ & new_B5534_;
  assign new_B5533_ = ~new_B5543_ | ~new_B5542_;
  assign new_B5534_ = B5515 | B5516;
  assign new_B5535_ = B5515 | new_B5522_;
  assign new_B5536_ = B5514 & new_B5526_;
  assign new_B5537_ = ~B5513 | ~B5514;
  assign new_B5538_ = new_B5522_ & new_B5537_;
  assign new_B5539_ = ~new_B5538_ & ~new_B5522_;
  assign new_B5540_ = new_B5522_ | new_B5537_;
  assign new_B5541_ = ~B5515 | ~B5516;
  assign new_B5542_ = new_B5522_ | new_B5537_;
  assign new_B5543_ = ~new_B5522_ & ~new_B5544_;
  assign new_B5544_ = new_B5522_ & new_B5537_;
  assign new_B5550_ = new_B5556_ & new_B5555_;
  assign new_B5551_ = new_B5558_ | new_B5557_;
  assign new_B5552_ = new_B5560_ | new_B5559_;
  assign new_B5553_ = new_B5555_ & new_B5561_;
  assign new_B5554_ = new_B5555_ & new_B5562_;
  assign new_B5555_ = B5545 ^ B5546;
  assign new_B5556_ = new_B5557_ ^ B5547;
  assign new_B5557_ = new_B5565_ & new_B5564_;
  assign new_B5558_ = new_B5563_ & B5547;
  assign new_B5559_ = new_B5568_ & new_B5567_;
  assign new_B5560_ = new_B5566_ & B5547;
  assign new_B5561_ = new_B5569_ | B5546;
  assign new_B5562_ = ~B5547 ^ new_B5559_;
  assign new_B5563_ = ~new_B5572_ | ~new_B5573_;
  assign new_B5564_ = B5548 ^ new_B5555_;
  assign new_B5565_ = new_B5574_ & new_B5567_;
  assign new_B5566_ = ~new_B5576_ | ~new_B5575_;
  assign new_B5567_ = B5548 | B5549;
  assign new_B5568_ = B5548 | new_B5555_;
  assign new_B5569_ = B5547 & new_B5559_;
  assign new_B5570_ = ~B5546 | ~B5547;
  assign new_B5571_ = new_B5555_ & new_B5570_;
  assign new_B5572_ = ~new_B5571_ & ~new_B5555_;
  assign new_B5573_ = new_B5555_ | new_B5570_;
  assign new_B5574_ = ~B5548 | ~B5549;
  assign new_B5575_ = new_B5555_ | new_B5570_;
  assign new_B5576_ = ~new_B5555_ & ~new_B5577_;
  assign new_B5577_ = new_B5555_ & new_B5570_;
  assign new_B5583_ = new_B5589_ & new_B5588_;
  assign new_B5584_ = new_B5591_ | new_B5590_;
  assign new_B5585_ = new_B5593_ | new_B5592_;
  assign new_B5586_ = new_B5588_ & new_B5594_;
  assign new_B5587_ = new_B5588_ & new_B5595_;
  assign new_B5588_ = B5578 ^ B5579;
  assign new_B5589_ = new_B5590_ ^ B5580;
  assign new_B5590_ = new_B5598_ & new_B5597_;
  assign new_B5591_ = new_B5596_ & B5580;
  assign new_B5592_ = new_B5601_ & new_B5600_;
  assign new_B5593_ = new_B5599_ & B5580;
  assign new_B5594_ = new_B5602_ | B5579;
  assign new_B5595_ = ~B5580 ^ new_B5592_;
  assign new_B5596_ = ~new_B5605_ | ~new_B5606_;
  assign new_B5597_ = B5581 ^ new_B5588_;
  assign new_B5598_ = new_B5607_ & new_B5600_;
  assign new_B5599_ = ~new_B5609_ | ~new_B5608_;
  assign new_B5600_ = B5581 | B5582;
  assign new_B5601_ = B5581 | new_B5588_;
  assign new_B5602_ = B5580 & new_B5592_;
  assign new_B5603_ = ~B5579 | ~B5580;
  assign new_B5604_ = new_B5588_ & new_B5603_;
  assign new_B5605_ = ~new_B5604_ & ~new_B5588_;
  assign new_B5606_ = new_B5588_ | new_B5603_;
  assign new_B5607_ = ~B5581 | ~B5582;
  assign new_B5608_ = new_B5588_ | new_B5603_;
  assign new_B5609_ = ~new_B5588_ & ~new_B5610_;
  assign new_B5610_ = new_B5588_ & new_B5603_;
  assign new_B5616_ = new_B5622_ & new_B5621_;
  assign new_B5617_ = new_B5624_ | new_B5623_;
  assign new_B5618_ = new_B5626_ | new_B5625_;
  assign new_B5619_ = new_B5621_ & new_B5627_;
  assign new_B5620_ = new_B5621_ & new_B5628_;
  assign new_B5621_ = B5611 ^ B5612;
  assign new_B5622_ = new_B5623_ ^ B5613;
  assign new_B5623_ = new_B5631_ & new_B5630_;
  assign new_B5624_ = new_B5629_ & B5613;
  assign new_B5625_ = new_B5634_ & new_B5633_;
  assign new_B5626_ = new_B5632_ & B5613;
  assign new_B5627_ = new_B5635_ | B5612;
  assign new_B5628_ = ~B5613 ^ new_B5625_;
  assign new_B5629_ = ~new_B5638_ | ~new_B5639_;
  assign new_B5630_ = B5614 ^ new_B5621_;
  assign new_B5631_ = new_B5640_ & new_B5633_;
  assign new_B5632_ = ~new_B5642_ | ~new_B5641_;
  assign new_B5633_ = B5614 | B5615;
  assign new_B5634_ = B5614 | new_B5621_;
  assign new_B5635_ = B5613 & new_B5625_;
  assign new_B5636_ = ~B5612 | ~B5613;
  assign new_B5637_ = new_B5621_ & new_B5636_;
  assign new_B5638_ = ~new_B5637_ & ~new_B5621_;
  assign new_B5639_ = new_B5621_ | new_B5636_;
  assign new_B5640_ = ~B5614 | ~B5615;
  assign new_B5641_ = new_B5621_ | new_B5636_;
  assign new_B5642_ = ~new_B5621_ & ~new_B5643_;
  assign new_B5643_ = new_B5621_ & new_B5636_;
  assign new_B5649_ = new_B5655_ & new_B5654_;
  assign new_B5650_ = new_B5657_ | new_B5656_;
  assign new_B5651_ = new_B5659_ | new_B5658_;
  assign new_B5652_ = new_B5654_ & new_B5660_;
  assign new_B5653_ = new_B5654_ & new_B5661_;
  assign new_B5654_ = B5644 ^ B5645;
  assign new_B5655_ = new_B5656_ ^ B5646;
  assign new_B5656_ = new_B5664_ & new_B5663_;
  assign new_B5657_ = new_B5662_ & B5646;
  assign new_B5658_ = new_B5667_ & new_B5666_;
  assign new_B5659_ = new_B5665_ & B5646;
  assign new_B5660_ = new_B5668_ | B5645;
  assign new_B5661_ = ~B5646 ^ new_B5658_;
  assign new_B5662_ = ~new_B5671_ | ~new_B5672_;
  assign new_B5663_ = B5647 ^ new_B5654_;
  assign new_B5664_ = new_B5673_ & new_B5666_;
  assign new_B5665_ = ~new_B5675_ | ~new_B5674_;
  assign new_B5666_ = B5647 | B5648;
  assign new_B5667_ = B5647 | new_B5654_;
  assign new_B5668_ = B5646 & new_B5658_;
  assign new_B5669_ = ~B5645 | ~B5646;
  assign new_B5670_ = new_B5654_ & new_B5669_;
  assign new_B5671_ = ~new_B5670_ & ~new_B5654_;
  assign new_B5672_ = new_B5654_ | new_B5669_;
  assign new_B5673_ = ~B5647 | ~B5648;
  assign new_B5674_ = new_B5654_ | new_B5669_;
  assign new_B5675_ = ~new_B5654_ & ~new_B5676_;
  assign new_B5676_ = new_B5654_ & new_B5669_;
  assign new_B5682_ = new_B5688_ & new_B5687_;
  assign new_B5683_ = new_B5690_ | new_B5689_;
  assign new_B5684_ = new_B5692_ | new_B5691_;
  assign new_B5685_ = new_B5687_ & new_B5693_;
  assign new_B5686_ = new_B5687_ & new_B5694_;
  assign new_B5687_ = B5677 ^ B5678;
  assign new_B5688_ = new_B5689_ ^ B5679;
  assign new_B5689_ = new_B5697_ & new_B5696_;
  assign new_B5690_ = new_B5695_ & B5679;
  assign new_B5691_ = new_B5700_ & new_B5699_;
  assign new_B5692_ = new_B5698_ & B5679;
  assign new_B5693_ = new_B5701_ | B5678;
  assign new_B5694_ = ~B5679 ^ new_B5691_;
  assign new_B5695_ = ~new_B5704_ | ~new_B5705_;
  assign new_B5696_ = B5680 ^ new_B5687_;
  assign new_B5697_ = new_B5706_ & new_B5699_;
  assign new_B5698_ = ~new_B5708_ | ~new_B5707_;
  assign new_B5699_ = B5680 | B5681;
  assign new_B5700_ = B5680 | new_B5687_;
  assign new_B5701_ = B5679 & new_B5691_;
  assign new_B5702_ = ~B5678 | ~B5679;
  assign new_B5703_ = new_B5687_ & new_B5702_;
  assign new_B5704_ = ~new_B5703_ & ~new_B5687_;
  assign new_B5705_ = new_B5687_ | new_B5702_;
  assign new_B5706_ = ~B5680 | ~B5681;
  assign new_B5707_ = new_B5687_ | new_B5702_;
  assign new_B5708_ = ~new_B5687_ & ~new_B5709_;
  assign new_B5709_ = new_B5687_ & new_B5702_;
  assign new_B5715_ = new_B5721_ & new_B5720_;
  assign new_B5716_ = new_B5723_ | new_B5722_;
  assign new_B5717_ = new_B5725_ | new_B5724_;
  assign new_B5718_ = new_B5720_ & new_B5726_;
  assign new_B5719_ = new_B5720_ & new_B5727_;
  assign new_B5720_ = B5710 ^ B5711;
  assign new_B5721_ = new_B5722_ ^ B5712;
  assign new_B5722_ = new_B5730_ & new_B5729_;
  assign new_B5723_ = new_B5728_ & B5712;
  assign new_B5724_ = new_B5733_ & new_B5732_;
  assign new_B5725_ = new_B5731_ & B5712;
  assign new_B5726_ = new_B5734_ | B5711;
  assign new_B5727_ = ~B5712 ^ new_B5724_;
  assign new_B5728_ = ~new_B5737_ | ~new_B5738_;
  assign new_B5729_ = B5713 ^ new_B5720_;
  assign new_B5730_ = new_B5739_ & new_B5732_;
  assign new_B5731_ = ~new_B5741_ | ~new_B5740_;
  assign new_B5732_ = B5713 | B5714;
  assign new_B5733_ = B5713 | new_B5720_;
  assign new_B5734_ = B5712 & new_B5724_;
  assign new_B5735_ = ~B5711 | ~B5712;
  assign new_B5736_ = new_B5720_ & new_B5735_;
  assign new_B5737_ = ~new_B5736_ & ~new_B5720_;
  assign new_B5738_ = new_B5720_ | new_B5735_;
  assign new_B5739_ = ~B5713 | ~B5714;
  assign new_B5740_ = new_B5720_ | new_B5735_;
  assign new_B5741_ = ~new_B5720_ & ~new_B5742_;
  assign new_B5742_ = new_B5720_ & new_B5735_;
  assign new_B5748_ = new_B5754_ & new_B5753_;
  assign new_B5749_ = new_B5756_ | new_B5755_;
  assign new_B5750_ = new_B5758_ | new_B5757_;
  assign new_B5751_ = new_B5753_ & new_B5759_;
  assign new_B5752_ = new_B5753_ & new_B5760_;
  assign new_B5753_ = B5743 ^ B5744;
  assign new_B5754_ = new_B5755_ ^ B5745;
  assign new_B5755_ = new_B5763_ & new_B5762_;
  assign new_B5756_ = new_B5761_ & B5745;
  assign new_B5757_ = new_B5766_ & new_B5765_;
  assign new_B5758_ = new_B5764_ & B5745;
  assign new_B5759_ = new_B5767_ | B5744;
  assign new_B5760_ = ~B5745 ^ new_B5757_;
  assign new_B5761_ = ~new_B5770_ | ~new_B5771_;
  assign new_B5762_ = B5746 ^ new_B5753_;
  assign new_B5763_ = new_B5772_ & new_B5765_;
  assign new_B5764_ = ~new_B5774_ | ~new_B5773_;
  assign new_B5765_ = B5746 | B5747;
  assign new_B5766_ = B5746 | new_B5753_;
  assign new_B5767_ = B5745 & new_B5757_;
  assign new_B5768_ = ~B5744 | ~B5745;
  assign new_B5769_ = new_B5753_ & new_B5768_;
  assign new_B5770_ = ~new_B5769_ & ~new_B5753_;
  assign new_B5771_ = new_B5753_ | new_B5768_;
  assign new_B5772_ = ~B5746 | ~B5747;
  assign new_B5773_ = new_B5753_ | new_B5768_;
  assign new_B5774_ = ~new_B5753_ & ~new_B5775_;
  assign new_B5775_ = new_B5753_ & new_B5768_;
  assign new_B5781_ = new_B5787_ & new_B5786_;
  assign new_B5782_ = new_B5789_ | new_B5788_;
  assign new_B5783_ = new_B5791_ | new_B5790_;
  assign new_B5784_ = new_B5786_ & new_B5792_;
  assign new_B5785_ = new_B5786_ & new_B5793_;
  assign new_B5786_ = B5776 ^ B5777;
  assign new_B5787_ = new_B5788_ ^ B5778;
  assign new_B5788_ = new_B5796_ & new_B5795_;
  assign new_B5789_ = new_B5794_ & B5778;
  assign new_B5790_ = new_B5799_ & new_B5798_;
  assign new_B5791_ = new_B5797_ & B5778;
  assign new_B5792_ = new_B5800_ | B5777;
  assign new_B5793_ = ~B5778 ^ new_B5790_;
  assign new_B5794_ = ~new_B5803_ | ~new_B5804_;
  assign new_B5795_ = B5779 ^ new_B5786_;
  assign new_B5796_ = new_B5805_ & new_B5798_;
  assign new_B5797_ = ~new_B5807_ | ~new_B5806_;
  assign new_B5798_ = B5779 | B5780;
  assign new_B5799_ = B5779 | new_B5786_;
  assign new_B5800_ = B5778 & new_B5790_;
  assign new_B5801_ = ~B5777 | ~B5778;
  assign new_B5802_ = new_B5786_ & new_B5801_;
  assign new_B5803_ = ~new_B5802_ & ~new_B5786_;
  assign new_B5804_ = new_B5786_ | new_B5801_;
  assign new_B5805_ = ~B5779 | ~B5780;
  assign new_B5806_ = new_B5786_ | new_B5801_;
  assign new_B5807_ = ~new_B5786_ & ~new_B5808_;
  assign new_B5808_ = new_B5786_ & new_B5801_;
  assign new_B5814_ = new_B5820_ & new_B5819_;
  assign new_B5815_ = new_B5822_ | new_B5821_;
  assign new_B5816_ = new_B5824_ | new_B5823_;
  assign new_B5817_ = new_B5819_ & new_B5825_;
  assign new_B5818_ = new_B5819_ & new_B5826_;
  assign new_B5819_ = B5809 ^ B5810;
  assign new_B5820_ = new_B5821_ ^ B5811;
  assign new_B5821_ = new_B5829_ & new_B5828_;
  assign new_B5822_ = new_B5827_ & B5811;
  assign new_B5823_ = new_B5832_ & new_B5831_;
  assign new_B5824_ = new_B5830_ & B5811;
  assign new_B5825_ = new_B5833_ | B5810;
  assign new_B5826_ = ~B5811 ^ new_B5823_;
  assign new_B5827_ = ~new_B5836_ | ~new_B5837_;
  assign new_B5828_ = B5812 ^ new_B5819_;
  assign new_B5829_ = new_B5838_ & new_B5831_;
  assign new_B5830_ = ~new_B5840_ | ~new_B5839_;
  assign new_B5831_ = B5812 | B5813;
  assign new_B5832_ = B5812 | new_B5819_;
  assign new_B5833_ = B5811 & new_B5823_;
  assign new_B5834_ = ~B5810 | ~B5811;
  assign new_B5835_ = new_B5819_ & new_B5834_;
  assign new_B5836_ = ~new_B5835_ & ~new_B5819_;
  assign new_B5837_ = new_B5819_ | new_B5834_;
  assign new_B5838_ = ~B5812 | ~B5813;
  assign new_B5839_ = new_B5819_ | new_B5834_;
  assign new_B5840_ = ~new_B5819_ & ~new_B5841_;
  assign new_B5841_ = new_B5819_ & new_B5834_;
  assign new_B5847_ = new_B5853_ & new_B5852_;
  assign new_B5848_ = new_B5855_ | new_B5854_;
  assign new_B5849_ = new_B5857_ | new_B5856_;
  assign new_B5850_ = new_B5852_ & new_B5858_;
  assign new_B5851_ = new_B5852_ & new_B5859_;
  assign new_B5852_ = B5842 ^ B5843;
  assign new_B5853_ = new_B5854_ ^ B5844;
  assign new_B5854_ = new_B5862_ & new_B5861_;
  assign new_B5855_ = new_B5860_ & B5844;
  assign new_B5856_ = new_B5865_ & new_B5864_;
  assign new_B5857_ = new_B5863_ & B5844;
  assign new_B5858_ = new_B5866_ | B5843;
  assign new_B5859_ = ~B5844 ^ new_B5856_;
  assign new_B5860_ = ~new_B5869_ | ~new_B5870_;
  assign new_B5861_ = B5845 ^ new_B5852_;
  assign new_B5862_ = new_B5871_ & new_B5864_;
  assign new_B5863_ = ~new_B5873_ | ~new_B5872_;
  assign new_B5864_ = B5845 | B5846;
  assign new_B5865_ = B5845 | new_B5852_;
  assign new_B5866_ = B5844 & new_B5856_;
  assign new_B5867_ = ~B5843 | ~B5844;
  assign new_B5868_ = new_B5852_ & new_B5867_;
  assign new_B5869_ = ~new_B5868_ & ~new_B5852_;
  assign new_B5870_ = new_B5852_ | new_B5867_;
  assign new_B5871_ = ~B5845 | ~B5846;
  assign new_B5872_ = new_B5852_ | new_B5867_;
  assign new_B5873_ = ~new_B5852_ & ~new_B5874_;
  assign new_B5874_ = new_B5852_ & new_B5867_;
  assign new_B5880_ = new_B5886_ & new_B5885_;
  assign new_B5881_ = new_B5888_ | new_B5887_;
  assign new_B5882_ = new_B5890_ | new_B5889_;
  assign new_B5883_ = new_B5885_ & new_B5891_;
  assign new_B5884_ = new_B5885_ & new_B5892_;
  assign new_B5885_ = B5875 ^ B5876;
  assign new_B5886_ = new_B5887_ ^ B5877;
  assign new_B5887_ = new_B5895_ & new_B5894_;
  assign new_B5888_ = new_B5893_ & B5877;
  assign new_B5889_ = new_B5898_ & new_B5897_;
  assign new_B5890_ = new_B5896_ & B5877;
  assign new_B5891_ = new_B5899_ | B5876;
  assign new_B5892_ = ~B5877 ^ new_B5889_;
  assign new_B5893_ = ~new_B5902_ | ~new_B5903_;
  assign new_B5894_ = B5878 ^ new_B5885_;
  assign new_B5895_ = new_B5904_ & new_B5897_;
  assign new_B5896_ = ~new_B5906_ | ~new_B5905_;
  assign new_B5897_ = B5878 | B5879;
  assign new_B5898_ = B5878 | new_B5885_;
  assign new_B5899_ = B5877 & new_B5889_;
  assign new_B5900_ = ~B5876 | ~B5877;
  assign new_B5901_ = new_B5885_ & new_B5900_;
  assign new_B5902_ = ~new_B5901_ & ~new_B5885_;
  assign new_B5903_ = new_B5885_ | new_B5900_;
  assign new_B5904_ = ~B5878 | ~B5879;
  assign new_B5905_ = new_B5885_ | new_B5900_;
  assign new_B5906_ = ~new_B5885_ & ~new_B5907_;
  assign new_B5907_ = new_B5885_ & new_B5900_;
  assign new_B5913_ = new_B5919_ & new_B5918_;
  assign new_B5914_ = new_B5921_ | new_B5920_;
  assign new_B5915_ = new_B5923_ | new_B5922_;
  assign new_B5916_ = new_B5918_ & new_B5924_;
  assign new_B5917_ = new_B5918_ & new_B5925_;
  assign new_B5918_ = B5908 ^ B5909;
  assign new_B5919_ = new_B5920_ ^ B5910;
  assign new_B5920_ = new_B5928_ & new_B5927_;
  assign new_B5921_ = new_B5926_ & B5910;
  assign new_B5922_ = new_B5931_ & new_B5930_;
  assign new_B5923_ = new_B5929_ & B5910;
  assign new_B5924_ = new_B5932_ | B5909;
  assign new_B5925_ = ~B5910 ^ new_B5922_;
  assign new_B5926_ = ~new_B5935_ | ~new_B5936_;
  assign new_B5927_ = B5911 ^ new_B5918_;
  assign new_B5928_ = new_B5937_ & new_B5930_;
  assign new_B5929_ = ~new_B5939_ | ~new_B5938_;
  assign new_B5930_ = B5911 | B5912;
  assign new_B5931_ = B5911 | new_B5918_;
  assign new_B5932_ = B5910 & new_B5922_;
  assign new_B5933_ = ~B5909 | ~B5910;
  assign new_B5934_ = new_B5918_ & new_B5933_;
  assign new_B5935_ = ~new_B5934_ & ~new_B5918_;
  assign new_B5936_ = new_B5918_ | new_B5933_;
  assign new_B5937_ = ~B5911 | ~B5912;
  assign new_B5938_ = new_B5918_ | new_B5933_;
  assign new_B5939_ = ~new_B5918_ & ~new_B5940_;
  assign new_B5940_ = new_B5918_ & new_B5933_;
  assign new_B5946_ = new_B5952_ & new_B5951_;
  assign new_B5947_ = new_B5954_ | new_B5953_;
  assign new_B5948_ = new_B5956_ | new_B5955_;
  assign new_B5949_ = new_B5951_ & new_B5957_;
  assign new_B5950_ = new_B5951_ & new_B5958_;
  assign new_B5951_ = B5941 ^ B5942;
  assign new_B5952_ = new_B5953_ ^ B5943;
  assign new_B5953_ = new_B5961_ & new_B5960_;
  assign new_B5954_ = new_B5959_ & B5943;
  assign new_B5955_ = new_B5964_ & new_B5963_;
  assign new_B5956_ = new_B5962_ & B5943;
  assign new_B5957_ = new_B5965_ | B5942;
  assign new_B5958_ = ~B5943 ^ new_B5955_;
  assign new_B5959_ = ~new_B5968_ | ~new_B5969_;
  assign new_B5960_ = B5944 ^ new_B5951_;
  assign new_B5961_ = new_B5970_ & new_B5963_;
  assign new_B5962_ = ~new_B5972_ | ~new_B5971_;
  assign new_B5963_ = B5944 | B5945;
  assign new_B5964_ = B5944 | new_B5951_;
  assign new_B5965_ = B5943 & new_B5955_;
  assign new_B5966_ = ~B5942 | ~B5943;
  assign new_B5967_ = new_B5951_ & new_B5966_;
  assign new_B5968_ = ~new_B5967_ & ~new_B5951_;
  assign new_B5969_ = new_B5951_ | new_B5966_;
  assign new_B5970_ = ~B5944 | ~B5945;
  assign new_B5971_ = new_B5951_ | new_B5966_;
  assign new_B5972_ = ~new_B5951_ & ~new_B5973_;
  assign new_B5973_ = new_B5951_ & new_B5966_;
  assign new_B5979_ = new_B5985_ & new_B5984_;
  assign new_B5980_ = new_B5987_ | new_B5986_;
  assign new_B5981_ = new_B5989_ | new_B5988_;
  assign new_B5982_ = new_B5984_ & new_B5990_;
  assign new_B5983_ = new_B5984_ & new_B5991_;
  assign new_B5984_ = B5974 ^ B5975;
  assign new_B5985_ = new_B5986_ ^ B5976;
  assign new_B5986_ = new_B5994_ & new_B5993_;
  assign new_B5987_ = new_B5992_ & B5976;
  assign new_B5988_ = new_B5997_ & new_B5996_;
  assign new_B5989_ = new_B5995_ & B5976;
  assign new_B5990_ = new_B5998_ | B5975;
  assign new_B5991_ = ~B5976 ^ new_B5988_;
  assign new_B5992_ = ~new_B6001_ | ~new_B6002_;
  assign new_B5993_ = B5977 ^ new_B5984_;
  assign new_B5994_ = new_B6003_ & new_B5996_;
  assign new_B5995_ = ~new_B6005_ | ~new_B6004_;
  assign new_B5996_ = B5977 | B5978;
  assign new_B5997_ = B5977 | new_B5984_;
  assign new_B5998_ = B5976 & new_B5988_;
  assign new_B5999_ = ~B5975 | ~B5976;
  assign new_B6000_ = new_B5984_ & new_B5999_;
  assign new_B6001_ = ~new_B6000_ & ~new_B5984_;
  assign new_B6002_ = new_B5984_ | new_B5999_;
  assign new_B6003_ = ~B5977 | ~B5978;
  assign new_B6004_ = new_B5984_ | new_B5999_;
  assign new_B6005_ = ~new_B5984_ & ~new_B6006_;
  assign new_B6006_ = new_B5984_ & new_B5999_;
  assign new_B6012_ = new_B6018_ & new_B6017_;
  assign new_B6013_ = new_B6020_ | new_B6019_;
  assign new_B6014_ = new_B6022_ | new_B6021_;
  assign new_B6015_ = new_B6017_ & new_B6023_;
  assign new_B6016_ = new_B6017_ & new_B6024_;
  assign new_B6017_ = B6007 ^ B6008;
  assign new_B6018_ = new_B6019_ ^ B6009;
  assign new_B6019_ = new_B6027_ & new_B6026_;
  assign new_B6020_ = new_B6025_ & B6009;
  assign new_B6021_ = new_B6030_ & new_B6029_;
  assign new_B6022_ = new_B6028_ & B6009;
  assign new_B6023_ = new_B6031_ | B6008;
  assign new_B6024_ = ~B6009 ^ new_B6021_;
  assign new_B6025_ = ~new_B6034_ | ~new_B6035_;
  assign new_B6026_ = B6010 ^ new_B6017_;
  assign new_B6027_ = new_B6036_ & new_B6029_;
  assign new_B6028_ = ~new_B6038_ | ~new_B6037_;
  assign new_B6029_ = B6010 | B6011;
  assign new_B6030_ = B6010 | new_B6017_;
  assign new_B6031_ = B6009 & new_B6021_;
  assign new_B6032_ = ~B6008 | ~B6009;
  assign new_B6033_ = new_B6017_ & new_B6032_;
  assign new_B6034_ = ~new_B6033_ & ~new_B6017_;
  assign new_B6035_ = new_B6017_ | new_B6032_;
  assign new_B6036_ = ~B6010 | ~B6011;
  assign new_B6037_ = new_B6017_ | new_B6032_;
  assign new_B6038_ = ~new_B6017_ & ~new_B6039_;
  assign new_B6039_ = new_B6017_ & new_B6032_;
  assign new_B6045_ = new_B6051_ & new_B6050_;
  assign new_B6046_ = new_B6053_ | new_B6052_;
  assign new_B6047_ = new_B6055_ | new_B6054_;
  assign new_B6048_ = new_B6050_ & new_B6056_;
  assign new_B6049_ = new_B6050_ & new_B6057_;
  assign new_B6050_ = B6040 ^ B6041;
  assign new_B6051_ = new_B6052_ ^ B6042;
  assign new_B6052_ = new_B6060_ & new_B6059_;
  assign new_B6053_ = new_B6058_ & B6042;
  assign new_B6054_ = new_B6063_ & new_B6062_;
  assign new_B6055_ = new_B6061_ & B6042;
  assign new_B6056_ = new_B6064_ | B6041;
  assign new_B6057_ = ~B6042 ^ new_B6054_;
  assign new_B6058_ = ~new_B6067_ | ~new_B6068_;
  assign new_B6059_ = B6043 ^ new_B6050_;
  assign new_B6060_ = new_B6069_ & new_B6062_;
  assign new_B6061_ = ~new_B6071_ | ~new_B6070_;
  assign new_B6062_ = B6043 | B6044;
  assign new_B6063_ = B6043 | new_B6050_;
  assign new_B6064_ = B6042 & new_B6054_;
  assign new_B6065_ = ~B6041 | ~B6042;
  assign new_B6066_ = new_B6050_ & new_B6065_;
  assign new_B6067_ = ~new_B6066_ & ~new_B6050_;
  assign new_B6068_ = new_B6050_ | new_B6065_;
  assign new_B6069_ = ~B6043 | ~B6044;
  assign new_B6070_ = new_B6050_ | new_B6065_;
  assign new_B6071_ = ~new_B6050_ & ~new_B6072_;
  assign new_B6072_ = new_B6050_ & new_B6065_;
  assign new_B6078_ = new_B6084_ & new_B6083_;
  assign new_B6079_ = new_B6086_ | new_B6085_;
  assign new_B6080_ = new_B6088_ | new_B6087_;
  assign new_B6081_ = new_B6083_ & new_B6089_;
  assign new_B6082_ = new_B6083_ & new_B6090_;
  assign new_B6083_ = B6073 ^ B6074;
  assign new_B6084_ = new_B6085_ ^ B6075;
  assign new_B6085_ = new_B6093_ & new_B6092_;
  assign new_B6086_ = new_B6091_ & B6075;
  assign new_B6087_ = new_B6096_ & new_B6095_;
  assign new_B6088_ = new_B6094_ & B6075;
  assign new_B6089_ = new_B6097_ | B6074;
  assign new_B6090_ = ~B6075 ^ new_B6087_;
  assign new_B6091_ = ~new_B6100_ | ~new_B6101_;
  assign new_B6092_ = B6076 ^ new_B6083_;
  assign new_B6093_ = new_B6102_ & new_B6095_;
  assign new_B6094_ = ~new_B6104_ | ~new_B6103_;
  assign new_B6095_ = B6076 | B6077;
  assign new_B6096_ = B6076 | new_B6083_;
  assign new_B6097_ = B6075 & new_B6087_;
  assign new_B6098_ = ~B6074 | ~B6075;
  assign new_B6099_ = new_B6083_ & new_B6098_;
  assign new_B6100_ = ~new_B6099_ & ~new_B6083_;
  assign new_B6101_ = new_B6083_ | new_B6098_;
  assign new_B6102_ = ~B6076 | ~B6077;
  assign new_B6103_ = new_B6083_ | new_B6098_;
  assign new_B6104_ = ~new_B6083_ & ~new_B6105_;
  assign new_B6105_ = new_B6083_ & new_B6098_;
  assign new_B6111_ = new_B6117_ & new_B6116_;
  assign new_B6112_ = new_B6119_ | new_B6118_;
  assign new_B6113_ = new_B6121_ | new_B6120_;
  assign new_B6114_ = new_B6116_ & new_B6122_;
  assign new_B6115_ = new_B6116_ & new_B6123_;
  assign new_B6116_ = B6106 ^ B6107;
  assign new_B6117_ = new_B6118_ ^ B6108;
  assign new_B6118_ = new_B6126_ & new_B6125_;
  assign new_B6119_ = new_B6124_ & B6108;
  assign new_B6120_ = new_B6129_ & new_B6128_;
  assign new_B6121_ = new_B6127_ & B6108;
  assign new_B6122_ = new_B6130_ | B6107;
  assign new_B6123_ = ~B6108 ^ new_B6120_;
  assign new_B6124_ = ~new_B6133_ | ~new_B6134_;
  assign new_B6125_ = B6109 ^ new_B6116_;
  assign new_B6126_ = new_B6135_ & new_B6128_;
  assign new_B6127_ = ~new_B6137_ | ~new_B6136_;
  assign new_B6128_ = B6109 | B6110;
  assign new_B6129_ = B6109 | new_B6116_;
  assign new_B6130_ = B6108 & new_B6120_;
  assign new_B6131_ = ~B6107 | ~B6108;
  assign new_B6132_ = new_B6116_ & new_B6131_;
  assign new_B6133_ = ~new_B6132_ & ~new_B6116_;
  assign new_B6134_ = new_B6116_ | new_B6131_;
  assign new_B6135_ = ~B6109 | ~B6110;
  assign new_B6136_ = new_B6116_ | new_B6131_;
  assign new_B6137_ = ~new_B6116_ & ~new_B6138_;
  assign new_B6138_ = new_B6116_ & new_B6131_;
  assign new_B6144_ = new_B6150_ & new_B6149_;
  assign new_B6145_ = new_B6152_ | new_B6151_;
  assign new_B6146_ = new_B6154_ | new_B6153_;
  assign new_B6147_ = new_B6149_ & new_B6155_;
  assign new_B6148_ = new_B6149_ & new_B6156_;
  assign new_B6149_ = B6139 ^ B6140;
  assign new_B6150_ = new_B6151_ ^ B6141;
  assign new_B6151_ = new_B6159_ & new_B6158_;
  assign new_B6152_ = new_B6157_ & B6141;
  assign new_B6153_ = new_B6162_ & new_B6161_;
  assign new_B6154_ = new_B6160_ & B6141;
  assign new_B6155_ = new_B6163_ | B6140;
  assign new_B6156_ = ~B6141 ^ new_B6153_;
  assign new_B6157_ = ~new_B6166_ | ~new_B6167_;
  assign new_B6158_ = B6142 ^ new_B6149_;
  assign new_B6159_ = new_B6168_ & new_B6161_;
  assign new_B6160_ = ~new_B6170_ | ~new_B6169_;
  assign new_B6161_ = B6142 | B6143;
  assign new_B6162_ = B6142 | new_B6149_;
  assign new_B6163_ = B6141 & new_B6153_;
  assign new_B6164_ = ~B6140 | ~B6141;
  assign new_B6165_ = new_B6149_ & new_B6164_;
  assign new_B6166_ = ~new_B6165_ & ~new_B6149_;
  assign new_B6167_ = new_B6149_ | new_B6164_;
  assign new_B6168_ = ~B6142 | ~B6143;
  assign new_B6169_ = new_B6149_ | new_B6164_;
  assign new_B6170_ = ~new_B6149_ & ~new_B6171_;
  assign new_B6171_ = new_B6149_ & new_B6164_;
  assign new_B6177_ = new_B6183_ & new_B6182_;
  assign new_B6178_ = new_B6185_ | new_B6184_;
  assign new_B6179_ = new_B6187_ | new_B6186_;
  assign new_B6180_ = new_B6182_ & new_B6188_;
  assign new_B6181_ = new_B6182_ & new_B6189_;
  assign new_B6182_ = B6172 ^ B6173;
  assign new_B6183_ = new_B6184_ ^ B6174;
  assign new_B6184_ = new_B6192_ & new_B6191_;
  assign new_B6185_ = new_B6190_ & B6174;
  assign new_B6186_ = new_B6195_ & new_B6194_;
  assign new_B6187_ = new_B6193_ & B6174;
  assign new_B6188_ = new_B6196_ | B6173;
  assign new_B6189_ = ~B6174 ^ new_B6186_;
  assign new_B6190_ = ~new_B6199_ | ~new_B6200_;
  assign new_B6191_ = B6175 ^ new_B6182_;
  assign new_B6192_ = new_B6201_ & new_B6194_;
  assign new_B6193_ = ~new_B6203_ | ~new_B6202_;
  assign new_B6194_ = B6175 | B6176;
  assign new_B6195_ = B6175 | new_B6182_;
  assign new_B6196_ = B6174 & new_B6186_;
  assign new_B6197_ = ~B6173 | ~B6174;
  assign new_B6198_ = new_B6182_ & new_B6197_;
  assign new_B6199_ = ~new_B6198_ & ~new_B6182_;
  assign new_B6200_ = new_B6182_ | new_B6197_;
  assign new_B6201_ = ~B6175 | ~B6176;
  assign new_B6202_ = new_B6182_ | new_B6197_;
  assign new_B6203_ = ~new_B6182_ & ~new_B6204_;
  assign new_B6204_ = new_B6182_ & new_B6197_;
  assign new_B6210_ = new_B6216_ & new_B6215_;
  assign new_B6211_ = new_B6218_ | new_B6217_;
  assign new_B6212_ = new_B6220_ | new_B6219_;
  assign new_B6213_ = new_B6215_ & new_B6221_;
  assign new_B6214_ = new_B6215_ & new_B6222_;
  assign new_B6215_ = B6205 ^ B6206;
  assign new_B6216_ = new_B6217_ ^ B6207;
  assign new_B6217_ = new_B6225_ & new_B6224_;
  assign new_B6218_ = new_B6223_ & B6207;
  assign new_B6219_ = new_B6228_ & new_B6227_;
  assign new_B6220_ = new_B6226_ & B6207;
  assign new_B6221_ = new_B6229_ | B6206;
  assign new_B6222_ = ~B6207 ^ new_B6219_;
  assign new_B6223_ = ~new_B6232_ | ~new_B6233_;
  assign new_B6224_ = B6208 ^ new_B6215_;
  assign new_B6225_ = new_B6234_ & new_B6227_;
  assign new_B6226_ = ~new_B6236_ | ~new_B6235_;
  assign new_B6227_ = B6208 | B6209;
  assign new_B6228_ = B6208 | new_B6215_;
  assign new_B6229_ = B6207 & new_B6219_;
  assign new_B6230_ = ~B6206 | ~B6207;
  assign new_B6231_ = new_B6215_ & new_B6230_;
  assign new_B6232_ = ~new_B6231_ & ~new_B6215_;
  assign new_B6233_ = new_B6215_ | new_B6230_;
  assign new_B6234_ = ~B6208 | ~B6209;
  assign new_B6235_ = new_B6215_ | new_B6230_;
  assign new_B6236_ = ~new_B6215_ & ~new_B6237_;
  assign new_B6237_ = new_B6215_ & new_B6230_;
  assign new_B6243_ = new_B6249_ & new_B6248_;
  assign new_B6244_ = new_B6251_ | new_B6250_;
  assign new_B6245_ = new_B6253_ | new_B6252_;
  assign new_B6246_ = new_B6248_ & new_B6254_;
  assign new_B6247_ = new_B6248_ & new_B6255_;
  assign new_B6248_ = B6238 ^ B6239;
  assign new_B6249_ = new_B6250_ ^ B6240;
  assign new_B6250_ = new_B6258_ & new_B6257_;
  assign new_B6251_ = new_B6256_ & B6240;
  assign new_B6252_ = new_B6261_ & new_B6260_;
  assign new_B6253_ = new_B6259_ & B6240;
  assign new_B6254_ = new_B6262_ | B6239;
  assign new_B6255_ = ~B6240 ^ new_B6252_;
  assign new_B6256_ = ~new_B6265_ | ~new_B6266_;
  assign new_B6257_ = B6241 ^ new_B6248_;
  assign new_B6258_ = new_B6267_ & new_B6260_;
  assign new_B6259_ = ~new_B6269_ | ~new_B6268_;
  assign new_B6260_ = B6241 | B6242;
  assign new_B6261_ = B6241 | new_B6248_;
  assign new_B6262_ = B6240 & new_B6252_;
  assign new_B6263_ = ~B6239 | ~B6240;
  assign new_B6264_ = new_B6248_ & new_B6263_;
  assign new_B6265_ = ~new_B6264_ & ~new_B6248_;
  assign new_B6266_ = new_B6248_ | new_B6263_;
  assign new_B6267_ = ~B6241 | ~B6242;
  assign new_B6268_ = new_B6248_ | new_B6263_;
  assign new_B6269_ = ~new_B6248_ & ~new_B6270_;
  assign new_B6270_ = new_B6248_ & new_B6263_;
  assign new_B6276_ = new_B6282_ & new_B6281_;
  assign new_B6277_ = new_B6284_ | new_B6283_;
  assign new_B6278_ = new_B6286_ | new_B6285_;
  assign new_B6279_ = new_B6281_ & new_B6287_;
  assign new_B6280_ = new_B6281_ & new_B6288_;
  assign new_B6281_ = B6271 ^ B6272;
  assign new_B6282_ = new_B6283_ ^ B6273;
  assign new_B6283_ = new_B6291_ & new_B6290_;
  assign new_B6284_ = new_B6289_ & B6273;
  assign new_B6285_ = new_B6294_ & new_B6293_;
  assign new_B6286_ = new_B6292_ & B6273;
  assign new_B6287_ = new_B6295_ | B6272;
  assign new_B6288_ = ~B6273 ^ new_B6285_;
  assign new_B6289_ = ~new_B6298_ | ~new_B6299_;
  assign new_B6290_ = B6274 ^ new_B6281_;
  assign new_B6291_ = new_B6300_ & new_B6293_;
  assign new_B6292_ = ~new_B6302_ | ~new_B6301_;
  assign new_B6293_ = B6274 | B6275;
  assign new_B6294_ = B6274 | new_B6281_;
  assign new_B6295_ = B6273 & new_B6285_;
  assign new_B6296_ = ~B6272 | ~B6273;
  assign new_B6297_ = new_B6281_ & new_B6296_;
  assign new_B6298_ = ~new_B6297_ & ~new_B6281_;
  assign new_B6299_ = new_B6281_ | new_B6296_;
  assign new_B6300_ = ~B6274 | ~B6275;
  assign new_B6301_ = new_B6281_ | new_B6296_;
  assign new_B6302_ = ~new_B6281_ & ~new_B6303_;
  assign new_B6303_ = new_B6281_ & new_B6296_;
  assign new_B6309_ = new_B6315_ & new_B6314_;
  assign new_B6310_ = new_B6317_ | new_B6316_;
  assign new_B6311_ = new_B6319_ | new_B6318_;
  assign new_B6312_ = new_B6314_ & new_B6320_;
  assign new_B6313_ = new_B6314_ & new_B6321_;
  assign new_B6314_ = B6304 ^ B6305;
  assign new_B6315_ = new_B6316_ ^ B6306;
  assign new_B6316_ = new_B6324_ & new_B6323_;
  assign new_B6317_ = new_B6322_ & B6306;
  assign new_B6318_ = new_B6327_ & new_B6326_;
  assign new_B6319_ = new_B6325_ & B6306;
  assign new_B6320_ = new_B6328_ | B6305;
  assign new_B6321_ = ~B6306 ^ new_B6318_;
  assign new_B6322_ = ~new_B6331_ | ~new_B6332_;
  assign new_B6323_ = B6307 ^ new_B6314_;
  assign new_B6324_ = new_B6333_ & new_B6326_;
  assign new_B6325_ = ~new_B6335_ | ~new_B6334_;
  assign new_B6326_ = B6307 | B6308;
  assign new_B6327_ = B6307 | new_B6314_;
  assign new_B6328_ = B6306 & new_B6318_;
  assign new_B6329_ = ~B6305 | ~B6306;
  assign new_B6330_ = new_B6314_ & new_B6329_;
  assign new_B6331_ = ~new_B6330_ & ~new_B6314_;
  assign new_B6332_ = new_B6314_ | new_B6329_;
  assign new_B6333_ = ~B6307 | ~B6308;
  assign new_B6334_ = new_B6314_ | new_B6329_;
  assign new_B6335_ = ~new_B6314_ & ~new_B6336_;
  assign new_B6336_ = new_B6314_ & new_B6329_;
  assign new_B6342_ = new_B6348_ & new_B6347_;
  assign new_B6343_ = new_B6350_ | new_B6349_;
  assign new_B6344_ = new_B6352_ | new_B6351_;
  assign new_B6345_ = new_B6347_ & new_B6353_;
  assign new_B6346_ = new_B6347_ & new_B6354_;
  assign new_B6347_ = B6337 ^ B6338;
  assign new_B6348_ = new_B6349_ ^ B6339;
  assign new_B6349_ = new_B6357_ & new_B6356_;
  assign new_B6350_ = new_B6355_ & B6339;
  assign new_B6351_ = new_B6360_ & new_B6359_;
  assign new_B6352_ = new_B6358_ & B6339;
  assign new_B6353_ = new_B6361_ | B6338;
  assign new_B6354_ = ~B6339 ^ new_B6351_;
  assign new_B6355_ = ~new_B6364_ | ~new_B6365_;
  assign new_B6356_ = B6340 ^ new_B6347_;
  assign new_B6357_ = new_B6366_ & new_B6359_;
  assign new_B6358_ = ~new_B6368_ | ~new_B6367_;
  assign new_B6359_ = B6340 | B6341;
  assign new_B6360_ = B6340 | new_B6347_;
  assign new_B6361_ = B6339 & new_B6351_;
  assign new_B6362_ = ~B6338 | ~B6339;
  assign new_B6363_ = new_B6347_ & new_B6362_;
  assign new_B6364_ = ~new_B6363_ & ~new_B6347_;
  assign new_B6365_ = new_B6347_ | new_B6362_;
  assign new_B6366_ = ~B6340 | ~B6341;
  assign new_B6367_ = new_B6347_ | new_B6362_;
  assign new_B6368_ = ~new_B6347_ & ~new_B6369_;
  assign new_B6369_ = new_B6347_ & new_B6362_;
  assign new_B6375_ = new_B6381_ & new_B6380_;
  assign new_B6376_ = new_B6383_ | new_B6382_;
  assign new_B6377_ = new_B6385_ | new_B6384_;
  assign new_B6378_ = new_B6380_ & new_B6386_;
  assign new_B6379_ = new_B6380_ & new_B6387_;
  assign new_B6380_ = B6370 ^ B6371;
  assign new_B6381_ = new_B6382_ ^ B6372;
  assign new_B6382_ = new_B6390_ & new_B6389_;
  assign new_B6383_ = new_B6388_ & B6372;
  assign new_B6384_ = new_B6393_ & new_B6392_;
  assign new_B6385_ = new_B6391_ & B6372;
  assign new_B6386_ = new_B6394_ | B6371;
  assign new_B6387_ = ~B6372 ^ new_B6384_;
  assign new_B6388_ = ~new_B6397_ | ~new_B6398_;
  assign new_B6389_ = B6373 ^ new_B6380_;
  assign new_B6390_ = new_B6399_ & new_B6392_;
  assign new_B6391_ = ~new_B6401_ | ~new_B6400_;
  assign new_B6392_ = B6373 | B6374;
  assign new_B6393_ = B6373 | new_B6380_;
  assign new_B6394_ = B6372 & new_B6384_;
  assign new_B6395_ = ~B6371 | ~B6372;
  assign new_B6396_ = new_B6380_ & new_B6395_;
  assign new_B6397_ = ~new_B6396_ & ~new_B6380_;
  assign new_B6398_ = new_B6380_ | new_B6395_;
  assign new_B6399_ = ~B6373 | ~B6374;
  assign new_B6400_ = new_B6380_ | new_B6395_;
  assign new_B6401_ = ~new_B6380_ & ~new_B6402_;
  assign new_B6402_ = new_B6380_ & new_B6395_;
  assign new_B6408_ = new_B6414_ & new_B6413_;
  assign new_B6409_ = new_B6416_ | new_B6415_;
  assign new_B6410_ = new_B6418_ | new_B6417_;
  assign new_B6411_ = new_B6413_ & new_B6419_;
  assign new_B6412_ = new_B6413_ & new_B6420_;
  assign new_B6413_ = B6403 ^ B6404;
  assign new_B6414_ = new_B6415_ ^ B6405;
  assign new_B6415_ = new_B6423_ & new_B6422_;
  assign new_B6416_ = new_B6421_ & B6405;
  assign new_B6417_ = new_B6426_ & new_B6425_;
  assign new_B6418_ = new_B6424_ & B6405;
  assign new_B6419_ = new_B6427_ | B6404;
  assign new_B6420_ = ~B6405 ^ new_B6417_;
  assign new_B6421_ = ~new_B6430_ | ~new_B6431_;
  assign new_B6422_ = B6406 ^ new_B6413_;
  assign new_B6423_ = new_B6432_ & new_B6425_;
  assign new_B6424_ = ~new_B6434_ | ~new_B6433_;
  assign new_B6425_ = B6406 | B6407;
  assign new_B6426_ = B6406 | new_B6413_;
  assign new_B6427_ = B6405 & new_B6417_;
  assign new_B6428_ = ~B6404 | ~B6405;
  assign new_B6429_ = new_B6413_ & new_B6428_;
  assign new_B6430_ = ~new_B6429_ & ~new_B6413_;
  assign new_B6431_ = new_B6413_ | new_B6428_;
  assign new_B6432_ = ~B6406 | ~B6407;
  assign new_B6433_ = new_B6413_ | new_B6428_;
  assign new_B6434_ = ~new_B6413_ & ~new_B6435_;
  assign new_B6435_ = new_B6413_ & new_B6428_;
  assign new_B6441_ = new_B6447_ & new_B6446_;
  assign new_B6442_ = new_B6449_ | new_B6448_;
  assign new_B6443_ = new_B6451_ | new_B6450_;
  assign new_B6444_ = new_B6446_ & new_B6452_;
  assign new_B6445_ = new_B6446_ & new_B6453_;
  assign new_B6446_ = B6436 ^ B6437;
  assign new_B6447_ = new_B6448_ ^ B6438;
  assign new_B6448_ = new_B6456_ & new_B6455_;
  assign new_B6449_ = new_B6454_ & B6438;
  assign new_B6450_ = new_B6459_ & new_B6458_;
  assign new_B6451_ = new_B6457_ & B6438;
  assign new_B6452_ = new_B6460_ | B6437;
  assign new_B6453_ = ~B6438 ^ new_B6450_;
  assign new_B6454_ = ~new_B6463_ | ~new_B6464_;
  assign new_B6455_ = B6439 ^ new_B6446_;
  assign new_B6456_ = new_B6465_ & new_B6458_;
  assign new_B6457_ = ~new_B6467_ | ~new_B6466_;
  assign new_B6458_ = B6439 | B6440;
  assign new_B6459_ = B6439 | new_B6446_;
  assign new_B6460_ = B6438 & new_B6450_;
  assign new_B6461_ = ~B6437 | ~B6438;
  assign new_B6462_ = new_B6446_ & new_B6461_;
  assign new_B6463_ = ~new_B6462_ & ~new_B6446_;
  assign new_B6464_ = new_B6446_ | new_B6461_;
  assign new_B6465_ = ~B6439 | ~B6440;
  assign new_B6466_ = new_B6446_ | new_B6461_;
  assign new_B6467_ = ~new_B6446_ & ~new_B6468_;
  assign new_B6468_ = new_B6446_ & new_B6461_;
  assign new_B6474_ = new_B6480_ & new_B6479_;
  assign new_B6475_ = new_B6482_ | new_B6481_;
  assign new_B6476_ = new_B6484_ | new_B6483_;
  assign new_B6477_ = new_B6479_ & new_B6485_;
  assign new_B6478_ = new_B6479_ & new_B6486_;
  assign new_B6479_ = B6469 ^ B6470;
  assign new_B6480_ = new_B6481_ ^ B6471;
  assign new_B6481_ = new_B6489_ & new_B6488_;
  assign new_B6482_ = new_B6487_ & B6471;
  assign new_B6483_ = new_B6492_ & new_B6491_;
  assign new_B6484_ = new_B6490_ & B6471;
  assign new_B6485_ = new_B6493_ | B6470;
  assign new_B6486_ = ~B6471 ^ new_B6483_;
  assign new_B6487_ = ~new_B6496_ | ~new_B6497_;
  assign new_B6488_ = B6472 ^ new_B6479_;
  assign new_B6489_ = new_B6498_ & new_B6491_;
  assign new_B6490_ = ~new_B6500_ | ~new_B6499_;
  assign new_B6491_ = B6472 | B6473;
  assign new_B6492_ = B6472 | new_B6479_;
  assign new_B6493_ = B6471 & new_B6483_;
  assign new_B6494_ = ~B6470 | ~B6471;
  assign new_B6495_ = new_B6479_ & new_B6494_;
  assign new_B6496_ = ~new_B6495_ & ~new_B6479_;
  assign new_B6497_ = new_B6479_ | new_B6494_;
  assign new_B6498_ = ~B6472 | ~B6473;
  assign new_B6499_ = new_B6479_ | new_B6494_;
  assign new_B6500_ = ~new_B6479_ & ~new_B6501_;
  assign new_B6501_ = new_B6479_ & new_B6494_;
  assign new_B6507_ = new_B6513_ & new_B6512_;
  assign new_B6508_ = new_B6515_ | new_B6514_;
  assign new_B6509_ = new_B6517_ | new_B6516_;
  assign new_B6510_ = new_B6512_ & new_B6518_;
  assign new_B6511_ = new_B6512_ & new_B6519_;
  assign new_B6512_ = B6502 ^ B6503;
  assign new_B6513_ = new_B6514_ ^ B6504;
  assign new_B6514_ = new_B6522_ & new_B6521_;
  assign new_B6515_ = new_B6520_ & B6504;
  assign new_B6516_ = new_B6525_ & new_B6524_;
  assign new_B6517_ = new_B6523_ & B6504;
  assign new_B6518_ = new_B6526_ | B6503;
  assign new_B6519_ = ~B6504 ^ new_B6516_;
  assign new_B6520_ = ~new_B6529_ | ~new_B6530_;
  assign new_B6521_ = B6505 ^ new_B6512_;
  assign new_B6522_ = new_B6531_ & new_B6524_;
  assign new_B6523_ = ~new_B6533_ | ~new_B6532_;
  assign new_B6524_ = B6505 | B6506;
  assign new_B6525_ = B6505 | new_B6512_;
  assign new_B6526_ = B6504 & new_B6516_;
  assign new_B6527_ = ~B6503 | ~B6504;
  assign new_B6528_ = new_B6512_ & new_B6527_;
  assign new_B6529_ = ~new_B6528_ & ~new_B6512_;
  assign new_B6530_ = new_B6512_ | new_B6527_;
  assign new_B6531_ = ~B6505 | ~B6506;
  assign new_B6532_ = new_B6512_ | new_B6527_;
  assign new_B6533_ = ~new_B6512_ & ~new_B6534_;
  assign new_B6534_ = new_B6512_ & new_B6527_;
  assign new_B6540_ = new_B6546_ & new_B6545_;
  assign new_B6541_ = new_B6548_ | new_B6547_;
  assign new_B6542_ = new_B6550_ | new_B6549_;
  assign new_B6543_ = new_B6545_ & new_B6551_;
  assign new_B6544_ = new_B6545_ & new_B6552_;
  assign new_B6545_ = B6535 ^ B6536;
  assign new_B6546_ = new_B6547_ ^ B6537;
  assign new_B6547_ = new_B6555_ & new_B6554_;
  assign new_B6548_ = new_B6553_ & B6537;
  assign new_B6549_ = new_B6558_ & new_B6557_;
  assign new_B6550_ = new_B6556_ & B6537;
  assign new_B6551_ = new_B6559_ | B6536;
  assign new_B6552_ = ~B6537 ^ new_B6549_;
  assign new_B6553_ = ~new_B6562_ | ~new_B6563_;
  assign new_B6554_ = B6538 ^ new_B6545_;
  assign new_B6555_ = new_B6564_ & new_B6557_;
  assign new_B6556_ = ~new_B6566_ | ~new_B6565_;
  assign new_B6557_ = B6538 | B6539;
  assign new_B6558_ = B6538 | new_B6545_;
  assign new_B6559_ = B6537 & new_B6549_;
  assign new_B6560_ = ~B6536 | ~B6537;
  assign new_B6561_ = new_B6545_ & new_B6560_;
  assign new_B6562_ = ~new_B6561_ & ~new_B6545_;
  assign new_B6563_ = new_B6545_ | new_B6560_;
  assign new_B6564_ = ~B6538 | ~B6539;
  assign new_B6565_ = new_B6545_ | new_B6560_;
  assign new_B6566_ = ~new_B6545_ & ~new_B6567_;
  assign new_B6567_ = new_B6545_ & new_B6560_;
  assign new_B6573_ = new_B6579_ & new_B6578_;
  assign new_B6574_ = new_B6581_ | new_B6580_;
  assign new_B6575_ = new_B6583_ | new_B6582_;
  assign new_B6576_ = new_B6578_ & new_B6584_;
  assign new_B6577_ = new_B6578_ & new_B6585_;
  assign new_B6578_ = B6568 ^ B6569;
  assign new_B6579_ = new_B6580_ ^ B6570;
  assign new_B6580_ = new_B6588_ & new_B6587_;
  assign new_B6581_ = new_B6586_ & B6570;
  assign new_B6582_ = new_B6591_ & new_B6590_;
  assign new_B6583_ = new_B6589_ & B6570;
  assign new_B6584_ = new_B6592_ | B6569;
  assign new_B6585_ = ~B6570 ^ new_B6582_;
  assign new_B6586_ = ~new_B6595_ | ~new_B6596_;
  assign new_B6587_ = B6571 ^ new_B6578_;
  assign new_B6588_ = new_B6597_ & new_B6590_;
  assign new_B6589_ = ~new_B6599_ | ~new_B6598_;
  assign new_B6590_ = B6571 | B6572;
  assign new_B6591_ = B6571 | new_B6578_;
  assign new_B6592_ = B6570 & new_B6582_;
  assign new_B6593_ = ~B6569 | ~B6570;
  assign new_B6594_ = new_B6578_ & new_B6593_;
  assign new_B6595_ = ~new_B6594_ & ~new_B6578_;
  assign new_B6596_ = new_B6578_ | new_B6593_;
  assign new_B6597_ = ~B6571 | ~B6572;
  assign new_B6598_ = new_B6578_ | new_B6593_;
  assign new_B6599_ = ~new_B6578_ & ~new_B6600_;
  assign new_B6600_ = new_B6578_ & new_B6593_;
  assign new_B6606_ = new_B6612_ & new_B6611_;
  assign new_B6607_ = new_B6614_ | new_B6613_;
  assign new_B6608_ = new_B6616_ | new_B6615_;
  assign new_B6609_ = new_B6611_ & new_B6617_;
  assign new_B6610_ = new_B6611_ & new_B6618_;
  assign new_B6611_ = B6601 ^ B6602;
  assign new_B6612_ = new_B6613_ ^ B6603;
  assign new_B6613_ = new_B6621_ & new_B6620_;
  assign new_B6614_ = new_B6619_ & B6603;
  assign new_B6615_ = new_B6624_ & new_B6623_;
  assign new_B6616_ = new_B6622_ & B6603;
  assign new_B6617_ = new_B6625_ | B6602;
  assign new_B6618_ = ~B6603 ^ new_B6615_;
  assign new_B6619_ = ~new_B6628_ | ~new_B6629_;
  assign new_B6620_ = B6604 ^ new_B6611_;
  assign new_B6621_ = new_B6630_ & new_B6623_;
  assign new_B6622_ = ~new_B6632_ | ~new_B6631_;
  assign new_B6623_ = B6604 | B6605;
  assign new_B6624_ = B6604 | new_B6611_;
  assign new_B6625_ = B6603 & new_B6615_;
  assign new_B6626_ = ~B6602 | ~B6603;
  assign new_B6627_ = new_B6611_ & new_B6626_;
  assign new_B6628_ = ~new_B6627_ & ~new_B6611_;
  assign new_B6629_ = new_B6611_ | new_B6626_;
  assign new_B6630_ = ~B6604 | ~B6605;
  assign new_B6631_ = new_B6611_ | new_B6626_;
  assign new_B6632_ = ~new_B6611_ & ~new_B6633_;
  assign new_B6633_ = new_B6611_ & new_B6626_;
  assign new_B6639_ = new_B6645_ & new_B6644_;
  assign new_B6640_ = new_B6647_ | new_B6646_;
  assign new_B6641_ = new_B6649_ | new_B6648_;
  assign new_B6642_ = new_B6644_ & new_B6650_;
  assign new_B6643_ = new_B6644_ & new_B6651_;
  assign new_B6644_ = B6634 ^ B6635;
  assign new_B6645_ = new_B6646_ ^ B6636;
  assign new_B6646_ = new_B6654_ & new_B6653_;
  assign new_B6647_ = new_B6652_ & B6636;
  assign new_B6648_ = new_B6657_ & new_B6656_;
  assign new_B6649_ = new_B6655_ & B6636;
  assign new_B6650_ = new_B6658_ | B6635;
  assign new_B6651_ = ~B6636 ^ new_B6648_;
  assign new_B6652_ = ~new_B6661_ | ~new_B6662_;
  assign new_B6653_ = B6637 ^ new_B6644_;
  assign new_B6654_ = new_B6663_ & new_B6656_;
  assign new_B6655_ = ~new_B6665_ | ~new_B6664_;
  assign new_B6656_ = B6637 | B6638;
  assign new_B6657_ = B6637 | new_B6644_;
  assign new_B6658_ = B6636 & new_B6648_;
  assign new_B6659_ = ~B6635 | ~B6636;
  assign new_B6660_ = new_B6644_ & new_B6659_;
  assign new_B6661_ = ~new_B6660_ & ~new_B6644_;
  assign new_B6662_ = new_B6644_ | new_B6659_;
  assign new_B6663_ = ~B6637 | ~B6638;
  assign new_B6664_ = new_B6644_ | new_B6659_;
  assign new_B6665_ = ~new_B6644_ & ~new_B6666_;
  assign new_B6666_ = new_B6644_ & new_B6659_;
  assign new_B6672_ = new_B6678_ & new_B6677_;
  assign new_B6673_ = new_B6680_ | new_B6679_;
  assign new_B6674_ = new_B6682_ | new_B6681_;
  assign new_B6675_ = new_B6677_ & new_B6683_;
  assign new_B6676_ = new_B6677_ & new_B6684_;
  assign new_B6677_ = B6667 ^ B6668;
  assign new_B6678_ = new_B6679_ ^ B6669;
  assign new_B6679_ = new_B6687_ & new_B6686_;
  assign new_B6680_ = new_B6685_ & B6669;
  assign new_B6681_ = new_B6690_ & new_B6689_;
  assign new_B6682_ = new_B6688_ & B6669;
  assign new_B6683_ = new_B6691_ | B6668;
  assign new_B6684_ = ~B6669 ^ new_B6681_;
  assign new_B6685_ = ~new_B6694_ | ~new_B6695_;
  assign new_B6686_ = B6670 ^ new_B6677_;
  assign new_B6687_ = new_B6696_ & new_B6689_;
  assign new_B6688_ = ~new_B6698_ | ~new_B6697_;
  assign new_B6689_ = B6670 | B6671;
  assign new_B6690_ = B6670 | new_B6677_;
  assign new_B6691_ = B6669 & new_B6681_;
  assign new_B6692_ = ~B6668 | ~B6669;
  assign new_B6693_ = new_B6677_ & new_B6692_;
  assign new_B6694_ = ~new_B6693_ & ~new_B6677_;
  assign new_B6695_ = new_B6677_ | new_B6692_;
  assign new_B6696_ = ~B6670 | ~B6671;
  assign new_B6697_ = new_B6677_ | new_B6692_;
  assign new_B6698_ = ~new_B6677_ & ~new_B6699_;
  assign new_B6699_ = new_B6677_ & new_B6692_;
  assign new_B6705_ = new_B6711_ & new_B6710_;
  assign new_B6706_ = new_B6713_ | new_B6712_;
  assign new_B6707_ = new_B6715_ | new_B6714_;
  assign new_B6708_ = new_B6710_ & new_B6716_;
  assign new_B6709_ = new_B6710_ & new_B6717_;
  assign new_B6710_ = B6700 ^ B6701;
  assign new_B6711_ = new_B6712_ ^ B6702;
  assign new_B6712_ = new_B6720_ & new_B6719_;
  assign new_B6713_ = new_B6718_ & B6702;
  assign new_B6714_ = new_B6723_ & new_B6722_;
  assign new_B6715_ = new_B6721_ & B6702;
  assign new_B6716_ = new_B6724_ | B6701;
  assign new_B6717_ = ~B6702 ^ new_B6714_;
  assign new_B6718_ = ~new_B6727_ | ~new_B6728_;
  assign new_B6719_ = B6703 ^ new_B6710_;
  assign new_B6720_ = new_B6729_ & new_B6722_;
  assign new_B6721_ = ~new_B6731_ | ~new_B6730_;
  assign new_B6722_ = B6703 | B6704;
  assign new_B6723_ = B6703 | new_B6710_;
  assign new_B6724_ = B6702 & new_B6714_;
  assign new_B6725_ = ~B6701 | ~B6702;
  assign new_B6726_ = new_B6710_ & new_B6725_;
  assign new_B6727_ = ~new_B6726_ & ~new_B6710_;
  assign new_B6728_ = new_B6710_ | new_B6725_;
  assign new_B6729_ = ~B6703 | ~B6704;
  assign new_B6730_ = new_B6710_ | new_B6725_;
  assign new_B6731_ = ~new_B6710_ & ~new_B6732_;
  assign new_B6732_ = new_B6710_ & new_B6725_;
  assign new_B6738_ = new_B6744_ & new_B6743_;
  assign new_B6739_ = new_B6746_ | new_B6745_;
  assign new_B6740_ = new_B6748_ | new_B6747_;
  assign new_B6741_ = new_B6743_ & new_B6749_;
  assign new_B6742_ = new_B6743_ & new_B6750_;
  assign new_B6743_ = B6733 ^ B6734;
  assign new_B6744_ = new_B6745_ ^ B6735;
  assign new_B6745_ = new_B6753_ & new_B6752_;
  assign new_B6746_ = new_B6751_ & B6735;
  assign new_B6747_ = new_B6756_ & new_B6755_;
  assign new_B6748_ = new_B6754_ & B6735;
  assign new_B6749_ = new_B6757_ | B6734;
  assign new_B6750_ = ~B6735 ^ new_B6747_;
  assign new_B6751_ = ~new_B6760_ | ~new_B6761_;
  assign new_B6752_ = B6736 ^ new_B6743_;
  assign new_B6753_ = new_B6762_ & new_B6755_;
  assign new_B6754_ = ~new_B6764_ | ~new_B6763_;
  assign new_B6755_ = B6736 | B6737;
  assign new_B6756_ = B6736 | new_B6743_;
  assign new_B6757_ = B6735 & new_B6747_;
  assign new_B6758_ = ~B6734 | ~B6735;
  assign new_B6759_ = new_B6743_ & new_B6758_;
  assign new_B6760_ = ~new_B6759_ & ~new_B6743_;
  assign new_B6761_ = new_B6743_ | new_B6758_;
  assign new_B6762_ = ~B6736 | ~B6737;
  assign new_B6763_ = new_B6743_ | new_B6758_;
  assign new_B6764_ = ~new_B6743_ & ~new_B6765_;
  assign new_B6765_ = new_B6743_ & new_B6758_;
  assign new_B6771_ = new_B6777_ & new_B6776_;
  assign new_B6772_ = new_B6779_ | new_B6778_;
  assign new_B6773_ = new_B6781_ | new_B6780_;
  assign new_B6774_ = new_B6776_ & new_B6782_;
  assign new_B6775_ = new_B6776_ & new_B6783_;
  assign new_B6776_ = B6766 ^ B6767;
  assign new_B6777_ = new_B6778_ ^ B6768;
  assign new_B6778_ = new_B6786_ & new_B6785_;
  assign new_B6779_ = new_B6784_ & B6768;
  assign new_B6780_ = new_B6789_ & new_B6788_;
  assign new_B6781_ = new_B6787_ & B6768;
  assign new_B6782_ = new_B6790_ | B6767;
  assign new_B6783_ = ~B6768 ^ new_B6780_;
  assign new_B6784_ = ~new_B6793_ | ~new_B6794_;
  assign new_B6785_ = B6769 ^ new_B6776_;
  assign new_B6786_ = new_B6795_ & new_B6788_;
  assign new_B6787_ = ~new_B6797_ | ~new_B6796_;
  assign new_B6788_ = B6769 | B6770;
  assign new_B6789_ = B6769 | new_B6776_;
  assign new_B6790_ = B6768 & new_B6780_;
  assign new_B6791_ = ~B6767 | ~B6768;
  assign new_B6792_ = new_B6776_ & new_B6791_;
  assign new_B6793_ = ~new_B6792_ & ~new_B6776_;
  assign new_B6794_ = new_B6776_ | new_B6791_;
  assign new_B6795_ = ~B6769 | ~B6770;
  assign new_B6796_ = new_B6776_ | new_B6791_;
  assign new_B6797_ = ~new_B6776_ & ~new_B6798_;
  assign new_B6798_ = new_B6776_ & new_B6791_;
  assign new_B6804_ = new_B6810_ & new_B6809_;
  assign new_B6805_ = new_B6812_ | new_B6811_;
  assign new_B6806_ = new_B6814_ | new_B6813_;
  assign new_B6807_ = new_B6809_ & new_B6815_;
  assign new_B6808_ = new_B6809_ & new_B6816_;
  assign new_B6809_ = B6799 ^ B6800;
  assign new_B6810_ = new_B6811_ ^ B6801;
  assign new_B6811_ = new_B6819_ & new_B6818_;
  assign new_B6812_ = new_B6817_ & B6801;
  assign new_B6813_ = new_B6822_ & new_B6821_;
  assign new_B6814_ = new_B6820_ & B6801;
  assign new_B6815_ = new_B6823_ | B6800;
  assign new_B6816_ = ~B6801 ^ new_B6813_;
  assign new_B6817_ = ~new_B6826_ | ~new_B6827_;
  assign new_B6818_ = B6802 ^ new_B6809_;
  assign new_B6819_ = new_B6828_ & new_B6821_;
  assign new_B6820_ = ~new_B6830_ | ~new_B6829_;
  assign new_B6821_ = B6802 | B6803;
  assign new_B6822_ = B6802 | new_B6809_;
  assign new_B6823_ = B6801 & new_B6813_;
  assign new_B6824_ = ~B6800 | ~B6801;
  assign new_B6825_ = new_B6809_ & new_B6824_;
  assign new_B6826_ = ~new_B6825_ & ~new_B6809_;
  assign new_B6827_ = new_B6809_ | new_B6824_;
  assign new_B6828_ = ~B6802 | ~B6803;
  assign new_B6829_ = new_B6809_ | new_B6824_;
  assign new_B6830_ = ~new_B6809_ & ~new_B6831_;
  assign new_B6831_ = new_B6809_ & new_B6824_;
  assign new_B6837_ = new_B6843_ & new_B6842_;
  assign new_B6838_ = new_B6845_ | new_B6844_;
  assign new_B6839_ = new_B6847_ | new_B6846_;
  assign new_B6840_ = new_B6842_ & new_B6848_;
  assign new_B6841_ = new_B6842_ & new_B6849_;
  assign new_B6842_ = B6832 ^ B6833;
  assign new_B6843_ = new_B6844_ ^ B6834;
  assign new_B6844_ = new_B6852_ & new_B6851_;
  assign new_B6845_ = new_B6850_ & B6834;
  assign new_B6846_ = new_B6855_ & new_B6854_;
  assign new_B6847_ = new_B6853_ & B6834;
  assign new_B6848_ = new_B6856_ | B6833;
  assign new_B6849_ = ~B6834 ^ new_B6846_;
  assign new_B6850_ = ~new_B6859_ | ~new_B6860_;
  assign new_B6851_ = B6835 ^ new_B6842_;
  assign new_B6852_ = new_B6861_ & new_B6854_;
  assign new_B6853_ = ~new_B6863_ | ~new_B6862_;
  assign new_B6854_ = B6835 | B6836;
  assign new_B6855_ = B6835 | new_B6842_;
  assign new_B6856_ = B6834 & new_B6846_;
  assign new_B6857_ = ~B6833 | ~B6834;
  assign new_B6858_ = new_B6842_ & new_B6857_;
  assign new_B6859_ = ~new_B6858_ & ~new_B6842_;
  assign new_B6860_ = new_B6842_ | new_B6857_;
  assign new_B6861_ = ~B6835 | ~B6836;
  assign new_B6862_ = new_B6842_ | new_B6857_;
  assign new_B6863_ = ~new_B6842_ & ~new_B6864_;
  assign new_B6864_ = new_B6842_ & new_B6857_;
  assign new_B6870_ = new_B6876_ & new_B6875_;
  assign new_B6871_ = new_B6878_ | new_B6877_;
  assign new_B6872_ = new_B6880_ | new_B6879_;
  assign new_B6873_ = new_B6875_ & new_B6881_;
  assign new_B6874_ = new_B6875_ & new_B6882_;
  assign new_B6875_ = B6865 ^ B6866;
  assign new_B6876_ = new_B6877_ ^ B6867;
  assign new_B6877_ = new_B6885_ & new_B6884_;
  assign new_B6878_ = new_B6883_ & B6867;
  assign new_B6879_ = new_B6888_ & new_B6887_;
  assign new_B6880_ = new_B6886_ & B6867;
  assign new_B6881_ = new_B6889_ | B6866;
  assign new_B6882_ = ~B6867 ^ new_B6879_;
  assign new_B6883_ = ~new_B6892_ | ~new_B6893_;
  assign new_B6884_ = B6868 ^ new_B6875_;
  assign new_B6885_ = new_B6894_ & new_B6887_;
  assign new_B6886_ = ~new_B6896_ | ~new_B6895_;
  assign new_B6887_ = B6868 | B6869;
  assign new_B6888_ = B6868 | new_B6875_;
  assign new_B6889_ = B6867 & new_B6879_;
  assign new_B6890_ = ~B6866 | ~B6867;
  assign new_B6891_ = new_B6875_ & new_B6890_;
  assign new_B6892_ = ~new_B6891_ & ~new_B6875_;
  assign new_B6893_ = new_B6875_ | new_B6890_;
  assign new_B6894_ = ~B6868 | ~B6869;
  assign new_B6895_ = new_B6875_ | new_B6890_;
  assign new_B6896_ = ~new_B6875_ & ~new_B6897_;
  assign new_B6897_ = new_B6875_ & new_B6890_;
  assign new_B6903_ = new_B6909_ & new_B6908_;
  assign new_B6904_ = new_B6911_ | new_B6910_;
  assign new_B6905_ = new_B6913_ | new_B6912_;
  assign new_B6906_ = new_B6908_ & new_B6914_;
  assign new_B6907_ = new_B6908_ & new_B6915_;
  assign new_B6908_ = B6898 ^ B6899;
  assign new_B6909_ = new_B6910_ ^ B6900;
  assign new_B6910_ = new_B6918_ & new_B6917_;
  assign new_B6911_ = new_B6916_ & B6900;
  assign new_B6912_ = new_B6921_ & new_B6920_;
  assign new_B6913_ = new_B6919_ & B6900;
  assign new_B6914_ = new_B6922_ | B6899;
  assign new_B6915_ = ~B6900 ^ new_B6912_;
  assign new_B6916_ = ~new_B6925_ | ~new_B6926_;
  assign new_B6917_ = B6901 ^ new_B6908_;
  assign new_B6918_ = new_B6927_ & new_B6920_;
  assign new_B6919_ = ~new_B6929_ | ~new_B6928_;
  assign new_B6920_ = B6901 | B6902;
  assign new_B6921_ = B6901 | new_B6908_;
  assign new_B6922_ = B6900 & new_B6912_;
  assign new_B6923_ = ~B6899 | ~B6900;
  assign new_B6924_ = new_B6908_ & new_B6923_;
  assign new_B6925_ = ~new_B6924_ & ~new_B6908_;
  assign new_B6926_ = new_B6908_ | new_B6923_;
  assign new_B6927_ = ~B6901 | ~B6902;
  assign new_B6928_ = new_B6908_ | new_B6923_;
  assign new_B6929_ = ~new_B6908_ & ~new_B6930_;
  assign new_B6930_ = new_B6908_ & new_B6923_;
  assign new_B6936_ = new_B6942_ & new_B6941_;
  assign new_B6937_ = new_B6944_ | new_B6943_;
  assign new_B6938_ = new_B6946_ | new_B6945_;
  assign new_B6939_ = new_B6941_ & new_B6947_;
  assign new_B6940_ = new_B6941_ & new_B6948_;
  assign new_B6941_ = B6931 ^ B6932;
  assign new_B6942_ = new_B6943_ ^ B6933;
  assign new_B6943_ = new_B6951_ & new_B6950_;
  assign new_B6944_ = new_B6949_ & B6933;
  assign new_B6945_ = new_B6954_ & new_B6953_;
  assign new_B6946_ = new_B6952_ & B6933;
  assign new_B6947_ = new_B6955_ | B6932;
  assign new_B6948_ = ~B6933 ^ new_B6945_;
  assign new_B6949_ = ~new_B6958_ | ~new_B6959_;
  assign new_B6950_ = B6934 ^ new_B6941_;
  assign new_B6951_ = new_B6960_ & new_B6953_;
  assign new_B6952_ = ~new_B6962_ | ~new_B6961_;
  assign new_B6953_ = B6934 | B6935;
  assign new_B6954_ = B6934 | new_B6941_;
  assign new_B6955_ = B6933 & new_B6945_;
  assign new_B6956_ = ~B6932 | ~B6933;
  assign new_B6957_ = new_B6941_ & new_B6956_;
  assign new_B6958_ = ~new_B6957_ & ~new_B6941_;
  assign new_B6959_ = new_B6941_ | new_B6956_;
  assign new_B6960_ = ~B6934 | ~B6935;
  assign new_B6961_ = new_B6941_ | new_B6956_;
  assign new_B6962_ = ~new_B6941_ & ~new_B6963_;
  assign new_B6963_ = new_B6941_ & new_B6956_;
  assign new_B6969_ = new_B6975_ & new_B6974_;
  assign new_B6970_ = new_B6977_ | new_B6976_;
  assign new_B6971_ = new_B6979_ | new_B6978_;
  assign new_B6972_ = new_B6974_ & new_B6980_;
  assign new_B6973_ = new_B6974_ & new_B6981_;
  assign new_B6974_ = B6964 ^ B6965;
  assign new_B6975_ = new_B6976_ ^ B6966;
  assign new_B6976_ = new_B6984_ & new_B6983_;
  assign new_B6977_ = new_B6982_ & B6966;
  assign new_B6978_ = new_B6987_ & new_B6986_;
  assign new_B6979_ = new_B6985_ & B6966;
  assign new_B6980_ = new_B6988_ | B6965;
  assign new_B6981_ = ~B6966 ^ new_B6978_;
  assign new_B6982_ = ~new_B6991_ | ~new_B6992_;
  assign new_B6983_ = B6967 ^ new_B6974_;
  assign new_B6984_ = new_B6993_ & new_B6986_;
  assign new_B6985_ = ~new_B6995_ | ~new_B6994_;
  assign new_B6986_ = B6967 | B6968;
  assign new_B6987_ = B6967 | new_B6974_;
  assign new_B6988_ = B6966 & new_B6978_;
  assign new_B6989_ = ~B6965 | ~B6966;
  assign new_B6990_ = new_B6974_ & new_B6989_;
  assign new_B6991_ = ~new_B6990_ & ~new_B6974_;
  assign new_B6992_ = new_B6974_ | new_B6989_;
  assign new_B6993_ = ~B6967 | ~B6968;
  assign new_B6994_ = new_B6974_ | new_B6989_;
  assign new_B6995_ = ~new_B6974_ & ~new_B6996_;
  assign new_B6996_ = new_B6974_ & new_B6989_;
  assign new_B7002_ = new_B7008_ & new_B7007_;
  assign new_B7003_ = new_B7010_ | new_B7009_;
  assign new_B7004_ = new_B7012_ | new_B7011_;
  assign new_B7005_ = new_B7007_ & new_B7013_;
  assign new_B7006_ = new_B7007_ & new_B7014_;
  assign new_B7007_ = B6997 ^ B6998;
  assign new_B7008_ = new_B7009_ ^ B6999;
  assign new_B7009_ = new_B7017_ & new_B7016_;
  assign new_B7010_ = new_B7015_ & B6999;
  assign new_B7011_ = new_B7020_ & new_B7019_;
  assign new_B7012_ = new_B7018_ & B6999;
  assign new_B7013_ = new_B7021_ | B6998;
  assign new_B7014_ = ~B6999 ^ new_B7011_;
  assign new_B7015_ = ~new_B7024_ | ~new_B7025_;
  assign new_B7016_ = B7000 ^ new_B7007_;
  assign new_B7017_ = new_B7026_ & new_B7019_;
  assign new_B7018_ = ~new_B7028_ | ~new_B7027_;
  assign new_B7019_ = B7000 | B7001;
  assign new_B7020_ = B7000 | new_B7007_;
  assign new_B7021_ = B6999 & new_B7011_;
  assign new_B7022_ = ~B6998 | ~B6999;
  assign new_B7023_ = new_B7007_ & new_B7022_;
  assign new_B7024_ = ~new_B7023_ & ~new_B7007_;
  assign new_B7025_ = new_B7007_ | new_B7022_;
  assign new_B7026_ = ~B7000 | ~B7001;
  assign new_B7027_ = new_B7007_ | new_B7022_;
  assign new_B7028_ = ~new_B7007_ & ~new_B7029_;
  assign new_B7029_ = new_B7007_ & new_B7022_;
  assign new_B7035_ = new_B7041_ & new_B7040_;
  assign new_B7036_ = new_B7043_ | new_B7042_;
  assign new_B7037_ = new_B7045_ | new_B7044_;
  assign new_B7038_ = new_B7040_ & new_B7046_;
  assign new_B7039_ = new_B7040_ & new_B7047_;
  assign new_B7040_ = B7030 ^ B7031;
  assign new_B7041_ = new_B7042_ ^ B7032;
  assign new_B7042_ = new_B7050_ & new_B7049_;
  assign new_B7043_ = new_B7048_ & B7032;
  assign new_B7044_ = new_B7053_ & new_B7052_;
  assign new_B7045_ = new_B7051_ & B7032;
  assign new_B7046_ = new_B7054_ | B7031;
  assign new_B7047_ = ~B7032 ^ new_B7044_;
  assign new_B7048_ = ~new_B7057_ | ~new_B7058_;
  assign new_B7049_ = B7033 ^ new_B7040_;
  assign new_B7050_ = new_B7059_ & new_B7052_;
  assign new_B7051_ = ~new_B7061_ | ~new_B7060_;
  assign new_B7052_ = B7033 | B7034;
  assign new_B7053_ = B7033 | new_B7040_;
  assign new_B7054_ = B7032 & new_B7044_;
  assign new_B7055_ = ~B7031 | ~B7032;
  assign new_B7056_ = new_B7040_ & new_B7055_;
  assign new_B7057_ = ~new_B7056_ & ~new_B7040_;
  assign new_B7058_ = new_B7040_ | new_B7055_;
  assign new_B7059_ = ~B7033 | ~B7034;
  assign new_B7060_ = new_B7040_ | new_B7055_;
  assign new_B7061_ = ~new_B7040_ & ~new_B7062_;
  assign new_B7062_ = new_B7040_ & new_B7055_;
  assign new_B7068_ = new_B7074_ & new_B7073_;
  assign new_B7069_ = new_B7076_ | new_B7075_;
  assign new_B7070_ = new_B7078_ | new_B7077_;
  assign new_B7071_ = new_B7073_ & new_B7079_;
  assign new_B7072_ = new_B7073_ & new_B7080_;
  assign new_B7073_ = B7063 ^ B7064;
  assign new_B7074_ = new_B7075_ ^ B7065;
  assign new_B7075_ = new_B7083_ & new_B7082_;
  assign new_B7076_ = new_B7081_ & B7065;
  assign new_B7077_ = new_B7086_ & new_B7085_;
  assign new_B7078_ = new_B7084_ & B7065;
  assign new_B7079_ = new_B7087_ | B7064;
  assign new_B7080_ = ~B7065 ^ new_B7077_;
  assign new_B7081_ = ~new_B7090_ | ~new_B7091_;
  assign new_B7082_ = B7066 ^ new_B7073_;
  assign new_B7083_ = new_B7092_ & new_B7085_;
  assign new_B7084_ = ~new_B7094_ | ~new_B7093_;
  assign new_B7085_ = B7066 | B7067;
  assign new_B7086_ = B7066 | new_B7073_;
  assign new_B7087_ = B7065 & new_B7077_;
  assign new_B7088_ = ~B7064 | ~B7065;
  assign new_B7089_ = new_B7073_ & new_B7088_;
  assign new_B7090_ = ~new_B7089_ & ~new_B7073_;
  assign new_B7091_ = new_B7073_ | new_B7088_;
  assign new_B7092_ = ~B7066 | ~B7067;
  assign new_B7093_ = new_B7073_ | new_B7088_;
  assign new_B7094_ = ~new_B7073_ & ~new_B7095_;
  assign new_B7095_ = new_B7073_ & new_B7088_;
  assign new_B7101_ = new_B7107_ & new_B7106_;
  assign new_B7102_ = new_B7109_ | new_B7108_;
  assign new_B7103_ = new_B7111_ | new_B7110_;
  assign new_B7104_ = new_B7106_ & new_B7112_;
  assign new_B7105_ = new_B7106_ & new_B7113_;
  assign new_B7106_ = B7096 ^ B7097;
  assign new_B7107_ = new_B7108_ ^ B7098;
  assign new_B7108_ = new_B7116_ & new_B7115_;
  assign new_B7109_ = new_B7114_ & B7098;
  assign new_B7110_ = new_B7119_ & new_B7118_;
  assign new_B7111_ = new_B7117_ & B7098;
  assign new_B7112_ = new_B7120_ | B7097;
  assign new_B7113_ = ~B7098 ^ new_B7110_;
  assign new_B7114_ = ~new_B7123_ | ~new_B7124_;
  assign new_B7115_ = B7099 ^ new_B7106_;
  assign new_B7116_ = new_B7125_ & new_B7118_;
  assign new_B7117_ = ~new_B7127_ | ~new_B7126_;
  assign new_B7118_ = B7099 | B7100;
  assign new_B7119_ = B7099 | new_B7106_;
  assign new_B7120_ = B7098 & new_B7110_;
  assign new_B7121_ = ~B7097 | ~B7098;
  assign new_B7122_ = new_B7106_ & new_B7121_;
  assign new_B7123_ = ~new_B7122_ & ~new_B7106_;
  assign new_B7124_ = new_B7106_ | new_B7121_;
  assign new_B7125_ = ~B7099 | ~B7100;
  assign new_B7126_ = new_B7106_ | new_B7121_;
  assign new_B7127_ = ~new_B7106_ & ~new_B7128_;
  assign new_B7128_ = new_B7106_ & new_B7121_;
  assign new_B7134_ = new_B7140_ & new_B7139_;
  assign new_B7135_ = new_B7142_ | new_B7141_;
  assign new_B7136_ = new_B7144_ | new_B7143_;
  assign new_B7137_ = new_B7139_ & new_B7145_;
  assign new_B7138_ = new_B7139_ & new_B7146_;
  assign new_B7139_ = B7129 ^ B7130;
  assign new_B7140_ = new_B7141_ ^ B7131;
  assign new_B7141_ = new_B7149_ & new_B7148_;
  assign new_B7142_ = new_B7147_ & B7131;
  assign new_B7143_ = new_B7152_ & new_B7151_;
  assign new_B7144_ = new_B7150_ & B7131;
  assign new_B7145_ = new_B7153_ | B7130;
  assign new_B7146_ = ~B7131 ^ new_B7143_;
  assign new_B7147_ = ~new_B7156_ | ~new_B7157_;
  assign new_B7148_ = B7132 ^ new_B7139_;
  assign new_B7149_ = new_B7158_ & new_B7151_;
  assign new_B7150_ = ~new_B7160_ | ~new_B7159_;
  assign new_B7151_ = B7132 | B7133;
  assign new_B7152_ = B7132 | new_B7139_;
  assign new_B7153_ = B7131 & new_B7143_;
  assign new_B7154_ = ~B7130 | ~B7131;
  assign new_B7155_ = new_B7139_ & new_B7154_;
  assign new_B7156_ = ~new_B7155_ & ~new_B7139_;
  assign new_B7157_ = new_B7139_ | new_B7154_;
  assign new_B7158_ = ~B7132 | ~B7133;
  assign new_B7159_ = new_B7139_ | new_B7154_;
  assign new_B7160_ = ~new_B7139_ & ~new_B7161_;
  assign new_B7161_ = new_B7139_ & new_B7154_;
  assign new_B7167_ = new_B7173_ & new_B7172_;
  assign new_B7168_ = new_B7175_ | new_B7174_;
  assign new_B7169_ = new_B7177_ | new_B7176_;
  assign new_B7170_ = new_B7172_ & new_B7178_;
  assign new_B7171_ = new_B7172_ & new_B7179_;
  assign new_B7172_ = B7162 ^ B7163;
  assign new_B7173_ = new_B7174_ ^ B7164;
  assign new_B7174_ = new_B7182_ & new_B7181_;
  assign new_B7175_ = new_B7180_ & B7164;
  assign new_B7176_ = new_B7185_ & new_B7184_;
  assign new_B7177_ = new_B7183_ & B7164;
  assign new_B7178_ = new_B7186_ | B7163;
  assign new_B7179_ = ~B7164 ^ new_B7176_;
  assign new_B7180_ = ~new_B7189_ | ~new_B7190_;
  assign new_B7181_ = B7165 ^ new_B7172_;
  assign new_B7182_ = new_B7191_ & new_B7184_;
  assign new_B7183_ = ~new_B7193_ | ~new_B7192_;
  assign new_B7184_ = B7165 | B7166;
  assign new_B7185_ = B7165 | new_B7172_;
  assign new_B7186_ = B7164 & new_B7176_;
  assign new_B7187_ = ~B7163 | ~B7164;
  assign new_B7188_ = new_B7172_ & new_B7187_;
  assign new_B7189_ = ~new_B7188_ & ~new_B7172_;
  assign new_B7190_ = new_B7172_ | new_B7187_;
  assign new_B7191_ = ~B7165 | ~B7166;
  assign new_B7192_ = new_B7172_ | new_B7187_;
  assign new_B7193_ = ~new_B7172_ & ~new_B7194_;
  assign new_B7194_ = new_B7172_ & new_B7187_;
  assign new_B7200_ = new_B7206_ & new_B7205_;
  assign new_B7201_ = new_B7208_ | new_B7207_;
  assign new_B7202_ = new_B7210_ | new_B7209_;
  assign new_B7203_ = new_B7205_ & new_B7211_;
  assign new_B7204_ = new_B7205_ & new_B7212_;
  assign new_B7205_ = B7195 ^ B7196;
  assign new_B7206_ = new_B7207_ ^ B7197;
  assign new_B7207_ = new_B7215_ & new_B7214_;
  assign new_B7208_ = new_B7213_ & B7197;
  assign new_B7209_ = new_B7218_ & new_B7217_;
  assign new_B7210_ = new_B7216_ & B7197;
  assign new_B7211_ = new_B7219_ | B7196;
  assign new_B7212_ = ~B7197 ^ new_B7209_;
  assign new_B7213_ = ~new_B7222_ | ~new_B7223_;
  assign new_B7214_ = B7198 ^ new_B7205_;
  assign new_B7215_ = new_B7224_ & new_B7217_;
  assign new_B7216_ = ~new_B7226_ | ~new_B7225_;
  assign new_B7217_ = B7198 | B7199;
  assign new_B7218_ = B7198 | new_B7205_;
  assign new_B7219_ = B7197 & new_B7209_;
  assign new_B7220_ = ~B7196 | ~B7197;
  assign new_B7221_ = new_B7205_ & new_B7220_;
  assign new_B7222_ = ~new_B7221_ & ~new_B7205_;
  assign new_B7223_ = new_B7205_ | new_B7220_;
  assign new_B7224_ = ~B7198 | ~B7199;
  assign new_B7225_ = new_B7205_ | new_B7220_;
  assign new_B7226_ = ~new_B7205_ & ~new_B7227_;
  assign new_B7227_ = new_B7205_ & new_B7220_;
  assign new_B7233_ = new_B7239_ & new_B7238_;
  assign new_B7234_ = new_B7241_ | new_B7240_;
  assign new_B7235_ = new_B7243_ | new_B7242_;
  assign new_B7236_ = new_B7238_ & new_B7244_;
  assign new_B7237_ = new_B7238_ & new_B7245_;
  assign new_B7238_ = B7228 ^ B7229;
  assign new_B7239_ = new_B7240_ ^ B7230;
  assign new_B7240_ = new_B7248_ & new_B7247_;
  assign new_B7241_ = new_B7246_ & B7230;
  assign new_B7242_ = new_B7251_ & new_B7250_;
  assign new_B7243_ = new_B7249_ & B7230;
  assign new_B7244_ = new_B7252_ | B7229;
  assign new_B7245_ = ~B7230 ^ new_B7242_;
  assign new_B7246_ = ~new_B7255_ | ~new_B7256_;
  assign new_B7247_ = B7231 ^ new_B7238_;
  assign new_B7248_ = new_B7257_ & new_B7250_;
  assign new_B7249_ = ~new_B7259_ | ~new_B7258_;
  assign new_B7250_ = B7231 | B7232;
  assign new_B7251_ = B7231 | new_B7238_;
  assign new_B7252_ = B7230 & new_B7242_;
  assign new_B7253_ = ~B7229 | ~B7230;
  assign new_B7254_ = new_B7238_ & new_B7253_;
  assign new_B7255_ = ~new_B7254_ & ~new_B7238_;
  assign new_B7256_ = new_B7238_ | new_B7253_;
  assign new_B7257_ = ~B7231 | ~B7232;
  assign new_B7258_ = new_B7238_ | new_B7253_;
  assign new_B7259_ = ~new_B7238_ & ~new_B7260_;
  assign new_B7260_ = new_B7238_ & new_B7253_;
  assign new_B7266_ = new_B7272_ & new_B7271_;
  assign new_B7267_ = new_B7274_ | new_B7273_;
  assign new_B7268_ = new_B7276_ | new_B7275_;
  assign new_B7269_ = new_B7271_ & new_B7277_;
  assign new_B7270_ = new_B7271_ & new_B7278_;
  assign new_B7271_ = B7261 ^ B7262;
  assign new_B7272_ = new_B7273_ ^ B7263;
  assign new_B7273_ = new_B7281_ & new_B7280_;
  assign new_B7274_ = new_B7279_ & B7263;
  assign new_B7275_ = new_B7284_ & new_B7283_;
  assign new_B7276_ = new_B7282_ & B7263;
  assign new_B7277_ = new_B7285_ | B7262;
  assign new_B7278_ = ~B7263 ^ new_B7275_;
  assign new_B7279_ = ~new_B7288_ | ~new_B7289_;
  assign new_B7280_ = B7264 ^ new_B7271_;
  assign new_B7281_ = new_B7290_ & new_B7283_;
  assign new_B7282_ = ~new_B7292_ | ~new_B7291_;
  assign new_B7283_ = B7264 | B7265;
  assign new_B7284_ = B7264 | new_B7271_;
  assign new_B7285_ = B7263 & new_B7275_;
  assign new_B7286_ = ~B7262 | ~B7263;
  assign new_B7287_ = new_B7271_ & new_B7286_;
  assign new_B7288_ = ~new_B7287_ & ~new_B7271_;
  assign new_B7289_ = new_B7271_ | new_B7286_;
  assign new_B7290_ = ~B7264 | ~B7265;
  assign new_B7291_ = new_B7271_ | new_B7286_;
  assign new_B7292_ = ~new_B7271_ & ~new_B7293_;
  assign new_B7293_ = new_B7271_ & new_B7286_;
  assign new_B7299_ = new_B7305_ & new_B7304_;
  assign new_B7300_ = new_B7307_ | new_B7306_;
  assign new_B7301_ = new_B7309_ | new_B7308_;
  assign new_B7302_ = new_B7304_ & new_B7310_;
  assign new_B7303_ = new_B7304_ & new_B7311_;
  assign new_B7304_ = B7294 ^ B7295;
  assign new_B7305_ = new_B7306_ ^ B7296;
  assign new_B7306_ = new_B7314_ & new_B7313_;
  assign new_B7307_ = new_B7312_ & B7296;
  assign new_B7308_ = new_B7317_ & new_B7316_;
  assign new_B7309_ = new_B7315_ & B7296;
  assign new_B7310_ = new_B7318_ | B7295;
  assign new_B7311_ = ~B7296 ^ new_B7308_;
  assign new_B7312_ = ~new_B7321_ | ~new_B7322_;
  assign new_B7313_ = B7297 ^ new_B7304_;
  assign new_B7314_ = new_B7323_ & new_B7316_;
  assign new_B7315_ = ~new_B7325_ | ~new_B7324_;
  assign new_B7316_ = B7297 | B7298;
  assign new_B7317_ = B7297 | new_B7304_;
  assign new_B7318_ = B7296 & new_B7308_;
  assign new_B7319_ = ~B7295 | ~B7296;
  assign new_B7320_ = new_B7304_ & new_B7319_;
  assign new_B7321_ = ~new_B7320_ & ~new_B7304_;
  assign new_B7322_ = new_B7304_ | new_B7319_;
  assign new_B7323_ = ~B7297 | ~B7298;
  assign new_B7324_ = new_B7304_ | new_B7319_;
  assign new_B7325_ = ~new_B7304_ & ~new_B7326_;
  assign new_B7326_ = new_B7304_ & new_B7319_;
  assign new_B7332_ = new_B7338_ & new_B7337_;
  assign new_B7333_ = new_B7340_ | new_B7339_;
  assign new_B7334_ = new_B7342_ | new_B7341_;
  assign new_B7335_ = new_B7337_ & new_B7343_;
  assign new_B7336_ = new_B7337_ & new_B7344_;
  assign new_B7337_ = B7327 ^ B7328;
  assign new_B7338_ = new_B7339_ ^ B7329;
  assign new_B7339_ = new_B7347_ & new_B7346_;
  assign new_B7340_ = new_B7345_ & B7329;
  assign new_B7341_ = new_B7350_ & new_B7349_;
  assign new_B7342_ = new_B7348_ & B7329;
  assign new_B7343_ = new_B7351_ | B7328;
  assign new_B7344_ = ~B7329 ^ new_B7341_;
  assign new_B7345_ = ~new_B7354_ | ~new_B7355_;
  assign new_B7346_ = B7330 ^ new_B7337_;
  assign new_B7347_ = new_B7356_ & new_B7349_;
  assign new_B7348_ = ~new_B7358_ | ~new_B7357_;
  assign new_B7349_ = B7330 | B7331;
  assign new_B7350_ = B7330 | new_B7337_;
  assign new_B7351_ = B7329 & new_B7341_;
  assign new_B7352_ = ~B7328 | ~B7329;
  assign new_B7353_ = new_B7337_ & new_B7352_;
  assign new_B7354_ = ~new_B7353_ & ~new_B7337_;
  assign new_B7355_ = new_B7337_ | new_B7352_;
  assign new_B7356_ = ~B7330 | ~B7331;
  assign new_B7357_ = new_B7337_ | new_B7352_;
  assign new_B7358_ = ~new_B7337_ & ~new_B7359_;
  assign new_B7359_ = new_B7337_ & new_B7352_;
  assign new_B7365_ = new_B7371_ & new_B7370_;
  assign new_B7366_ = new_B7373_ | new_B7372_;
  assign new_B7367_ = new_B7375_ | new_B7374_;
  assign new_B7368_ = new_B7370_ & new_B7376_;
  assign new_B7369_ = new_B7370_ & new_B7377_;
  assign new_B7370_ = B7360 ^ B7361;
  assign new_B7371_ = new_B7372_ ^ B7362;
  assign new_B7372_ = new_B7380_ & new_B7379_;
  assign new_B7373_ = new_B7378_ & B7362;
  assign new_B7374_ = new_B7383_ & new_B7382_;
  assign new_B7375_ = new_B7381_ & B7362;
  assign new_B7376_ = new_B7384_ | B7361;
  assign new_B7377_ = ~B7362 ^ new_B7374_;
  assign new_B7378_ = ~new_B7387_ | ~new_B7388_;
  assign new_B7379_ = B7363 ^ new_B7370_;
  assign new_B7380_ = new_B7389_ & new_B7382_;
  assign new_B7381_ = ~new_B7391_ | ~new_B7390_;
  assign new_B7382_ = B7363 | B7364;
  assign new_B7383_ = B7363 | new_B7370_;
  assign new_B7384_ = B7362 & new_B7374_;
  assign new_B7385_ = ~B7361 | ~B7362;
  assign new_B7386_ = new_B7370_ & new_B7385_;
  assign new_B7387_ = ~new_B7386_ & ~new_B7370_;
  assign new_B7388_ = new_B7370_ | new_B7385_;
  assign new_B7389_ = ~B7363 | ~B7364;
  assign new_B7390_ = new_B7370_ | new_B7385_;
  assign new_B7391_ = ~new_B7370_ & ~new_B7392_;
  assign new_B7392_ = new_B7370_ & new_B7385_;
  assign new_B7398_ = new_B7404_ & new_B7403_;
  assign new_B7399_ = new_B7406_ | new_B7405_;
  assign new_B7400_ = new_B7408_ | new_B7407_;
  assign new_B7401_ = new_B7403_ & new_B7409_;
  assign new_B7402_ = new_B7403_ & new_B7410_;
  assign new_B7403_ = B7393 ^ B7394;
  assign new_B7404_ = new_B7405_ ^ B7395;
  assign new_B7405_ = new_B7413_ & new_B7412_;
  assign new_B7406_ = new_B7411_ & B7395;
  assign new_B7407_ = new_B7416_ & new_B7415_;
  assign new_B7408_ = new_B7414_ & B7395;
  assign new_B7409_ = new_B7417_ | B7394;
  assign new_B7410_ = ~B7395 ^ new_B7407_;
  assign new_B7411_ = ~new_B7420_ | ~new_B7421_;
  assign new_B7412_ = B7396 ^ new_B7403_;
  assign new_B7413_ = new_B7422_ & new_B7415_;
  assign new_B7414_ = ~new_B7424_ | ~new_B7423_;
  assign new_B7415_ = B7396 | B7397;
  assign new_B7416_ = B7396 | new_B7403_;
  assign new_B7417_ = B7395 & new_B7407_;
  assign new_B7418_ = ~B7394 | ~B7395;
  assign new_B7419_ = new_B7403_ & new_B7418_;
  assign new_B7420_ = ~new_B7419_ & ~new_B7403_;
  assign new_B7421_ = new_B7403_ | new_B7418_;
  assign new_B7422_ = ~B7396 | ~B7397;
  assign new_B7423_ = new_B7403_ | new_B7418_;
  assign new_B7424_ = ~new_B7403_ & ~new_B7425_;
  assign new_B7425_ = new_B7403_ & new_B7418_;
  assign new_B7431_ = new_B7437_ & new_B7436_;
  assign new_B7432_ = new_B7439_ | new_B7438_;
  assign new_B7433_ = new_B7441_ | new_B7440_;
  assign new_B7434_ = new_B7436_ & new_B7442_;
  assign new_B7435_ = new_B7436_ & new_B7443_;
  assign new_B7436_ = B7426 ^ B7427;
  assign new_B7437_ = new_B7438_ ^ B7428;
  assign new_B7438_ = new_B7446_ & new_B7445_;
  assign new_B7439_ = new_B7444_ & B7428;
  assign new_B7440_ = new_B7449_ & new_B7448_;
  assign new_B7441_ = new_B7447_ & B7428;
  assign new_B7442_ = new_B7450_ | B7427;
  assign new_B7443_ = ~B7428 ^ new_B7440_;
  assign new_B7444_ = ~new_B7453_ | ~new_B7454_;
  assign new_B7445_ = B7429 ^ new_B7436_;
  assign new_B7446_ = new_B7455_ & new_B7448_;
  assign new_B7447_ = ~new_B7457_ | ~new_B7456_;
  assign new_B7448_ = B7429 | B7430;
  assign new_B7449_ = B7429 | new_B7436_;
  assign new_B7450_ = B7428 & new_B7440_;
  assign new_B7451_ = ~B7427 | ~B7428;
  assign new_B7452_ = new_B7436_ & new_B7451_;
  assign new_B7453_ = ~new_B7452_ & ~new_B7436_;
  assign new_B7454_ = new_B7436_ | new_B7451_;
  assign new_B7455_ = ~B7429 | ~B7430;
  assign new_B7456_ = new_B7436_ | new_B7451_;
  assign new_B7457_ = ~new_B7436_ & ~new_B7458_;
  assign new_B7458_ = new_B7436_ & new_B7451_;
  assign new_B7464_ = new_B7470_ & new_B7469_;
  assign new_B7465_ = new_B7472_ | new_B7471_;
  assign new_B7466_ = new_B7474_ | new_B7473_;
  assign new_B7467_ = new_B7469_ & new_B7475_;
  assign new_B7468_ = new_B7469_ & new_B7476_;
  assign new_B7469_ = B7459 ^ B7460;
  assign new_B7470_ = new_B7471_ ^ B7461;
  assign new_B7471_ = new_B7479_ & new_B7478_;
  assign new_B7472_ = new_B7477_ & B7461;
  assign new_B7473_ = new_B7482_ & new_B7481_;
  assign new_B7474_ = new_B7480_ & B7461;
  assign new_B7475_ = new_B7483_ | B7460;
  assign new_B7476_ = ~B7461 ^ new_B7473_;
  assign new_B7477_ = ~new_B7486_ | ~new_B7487_;
  assign new_B7478_ = B7462 ^ new_B7469_;
  assign new_B7479_ = new_B7488_ & new_B7481_;
  assign new_B7480_ = ~new_B7490_ | ~new_B7489_;
  assign new_B7481_ = B7462 | B7463;
  assign new_B7482_ = B7462 | new_B7469_;
  assign new_B7483_ = B7461 & new_B7473_;
  assign new_B7484_ = ~B7460 | ~B7461;
  assign new_B7485_ = new_B7469_ & new_B7484_;
  assign new_B7486_ = ~new_B7485_ & ~new_B7469_;
  assign new_B7487_ = new_B7469_ | new_B7484_;
  assign new_B7488_ = ~B7462 | ~B7463;
  assign new_B7489_ = new_B7469_ | new_B7484_;
  assign new_B7490_ = ~new_B7469_ & ~new_B7491_;
  assign new_B7491_ = new_B7469_ & new_B7484_;
  assign new_B7497_ = new_B7503_ & new_B7502_;
  assign new_B7498_ = new_B7505_ | new_B7504_;
  assign new_B7499_ = new_B7507_ | new_B7506_;
  assign new_B7500_ = new_B7502_ & new_B7508_;
  assign new_B7501_ = new_B7502_ & new_B7509_;
  assign new_B7502_ = B7492 ^ B7493;
  assign new_B7503_ = new_B7504_ ^ B7494;
  assign new_B7504_ = new_B7512_ & new_B7511_;
  assign new_B7505_ = new_B7510_ & B7494;
  assign new_B7506_ = new_B7515_ & new_B7514_;
  assign new_B7507_ = new_B7513_ & B7494;
  assign new_B7508_ = new_B7516_ | B7493;
  assign new_B7509_ = ~B7494 ^ new_B7506_;
  assign new_B7510_ = ~new_B7519_ | ~new_B7520_;
  assign new_B7511_ = B7495 ^ new_B7502_;
  assign new_B7512_ = new_B7521_ & new_B7514_;
  assign new_B7513_ = ~new_B7523_ | ~new_B7522_;
  assign new_B7514_ = B7495 | B7496;
  assign new_B7515_ = B7495 | new_B7502_;
  assign new_B7516_ = B7494 & new_B7506_;
  assign new_B7517_ = ~B7493 | ~B7494;
  assign new_B7518_ = new_B7502_ & new_B7517_;
  assign new_B7519_ = ~new_B7518_ & ~new_B7502_;
  assign new_B7520_ = new_B7502_ | new_B7517_;
  assign new_B7521_ = ~B7495 | ~B7496;
  assign new_B7522_ = new_B7502_ | new_B7517_;
  assign new_B7523_ = ~new_B7502_ & ~new_B7524_;
  assign new_B7524_ = new_B7502_ & new_B7517_;
  assign new_B7530_ = new_B7536_ & new_B7535_;
  assign new_B7531_ = new_B7538_ | new_B7537_;
  assign new_B7532_ = new_B7540_ | new_B7539_;
  assign new_B7533_ = new_B7535_ & new_B7541_;
  assign new_B7534_ = new_B7535_ & new_B7542_;
  assign new_B7535_ = B7525 ^ B7526;
  assign new_B7536_ = new_B7537_ ^ B7527;
  assign new_B7537_ = new_B7545_ & new_B7544_;
  assign new_B7538_ = new_B7543_ & B7527;
  assign new_B7539_ = new_B7548_ & new_B7547_;
  assign new_B7540_ = new_B7546_ & B7527;
  assign new_B7541_ = new_B7549_ | B7526;
  assign new_B7542_ = ~B7527 ^ new_B7539_;
  assign new_B7543_ = ~new_B7552_ | ~new_B7553_;
  assign new_B7544_ = B7528 ^ new_B7535_;
  assign new_B7545_ = new_B7554_ & new_B7547_;
  assign new_B7546_ = ~new_B7556_ | ~new_B7555_;
  assign new_B7547_ = B7528 | B7529;
  assign new_B7548_ = B7528 | new_B7535_;
  assign new_B7549_ = B7527 & new_B7539_;
  assign new_B7550_ = ~B7526 | ~B7527;
  assign new_B7551_ = new_B7535_ & new_B7550_;
  assign new_B7552_ = ~new_B7551_ & ~new_B7535_;
  assign new_B7553_ = new_B7535_ | new_B7550_;
  assign new_B7554_ = ~B7528 | ~B7529;
  assign new_B7555_ = new_B7535_ | new_B7550_;
  assign new_B7556_ = ~new_B7535_ & ~new_B7557_;
  assign new_B7557_ = new_B7535_ & new_B7550_;
  assign new_B7563_ = new_B7569_ & new_B7568_;
  assign new_B7564_ = new_B7571_ | new_B7570_;
  assign new_B7565_ = new_B7573_ | new_B7572_;
  assign new_B7566_ = new_B7568_ & new_B7574_;
  assign new_B7567_ = new_B7568_ & new_B7575_;
  assign new_B7568_ = B7558 ^ B7559;
  assign new_B7569_ = new_B7570_ ^ B7560;
  assign new_B7570_ = new_B7578_ & new_B7577_;
  assign new_B7571_ = new_B7576_ & B7560;
  assign new_B7572_ = new_B7581_ & new_B7580_;
  assign new_B7573_ = new_B7579_ & B7560;
  assign new_B7574_ = new_B7582_ | B7559;
  assign new_B7575_ = ~B7560 ^ new_B7572_;
  assign new_B7576_ = ~new_B7585_ | ~new_B7586_;
  assign new_B7577_ = B7561 ^ new_B7568_;
  assign new_B7578_ = new_B7587_ & new_B7580_;
  assign new_B7579_ = ~new_B7589_ | ~new_B7588_;
  assign new_B7580_ = B7561 | B7562;
  assign new_B7581_ = B7561 | new_B7568_;
  assign new_B7582_ = B7560 & new_B7572_;
  assign new_B7583_ = ~B7559 | ~B7560;
  assign new_B7584_ = new_B7568_ & new_B7583_;
  assign new_B7585_ = ~new_B7584_ & ~new_B7568_;
  assign new_B7586_ = new_B7568_ | new_B7583_;
  assign new_B7587_ = ~B7561 | ~B7562;
  assign new_B7588_ = new_B7568_ | new_B7583_;
  assign new_B7589_ = ~new_B7568_ & ~new_B7590_;
  assign new_B7590_ = new_B7568_ & new_B7583_;
  assign new_B7596_ = new_B7602_ & new_B7601_;
  assign new_B7597_ = new_B7604_ | new_B7603_;
  assign new_B7598_ = new_B7606_ | new_B7605_;
  assign new_B7599_ = new_B7601_ & new_B7607_;
  assign new_B7600_ = new_B7601_ & new_B7608_;
  assign new_B7601_ = B7591 ^ B7592;
  assign new_B7602_ = new_B7603_ ^ B7593;
  assign new_B7603_ = new_B7611_ & new_B7610_;
  assign new_B7604_ = new_B7609_ & B7593;
  assign new_B7605_ = new_B7614_ & new_B7613_;
  assign new_B7606_ = new_B7612_ & B7593;
  assign new_B7607_ = new_B7615_ | B7592;
  assign new_B7608_ = ~B7593 ^ new_B7605_;
  assign new_B7609_ = ~new_B7618_ | ~new_B7619_;
  assign new_B7610_ = B7594 ^ new_B7601_;
  assign new_B7611_ = new_B7620_ & new_B7613_;
  assign new_B7612_ = ~new_B7622_ | ~new_B7621_;
  assign new_B7613_ = B7594 | B7595;
  assign new_B7614_ = B7594 | new_B7601_;
  assign new_B7615_ = B7593 & new_B7605_;
  assign new_B7616_ = ~B7592 | ~B7593;
  assign new_B7617_ = new_B7601_ & new_B7616_;
  assign new_B7618_ = ~new_B7617_ & ~new_B7601_;
  assign new_B7619_ = new_B7601_ | new_B7616_;
  assign new_B7620_ = ~B7594 | ~B7595;
  assign new_B7621_ = new_B7601_ | new_B7616_;
  assign new_B7622_ = ~new_B7601_ & ~new_B7623_;
  assign new_B7623_ = new_B7601_ & new_B7616_;
  assign new_B7629_ = new_B7635_ & new_B7634_;
  assign new_B7630_ = new_B7637_ | new_B7636_;
  assign new_B7631_ = new_B7639_ | new_B7638_;
  assign new_B7632_ = new_B7634_ & new_B7640_;
  assign new_B7633_ = new_B7634_ & new_B7641_;
  assign new_B7634_ = B7624 ^ B7625;
  assign new_B7635_ = new_B7636_ ^ B7626;
  assign new_B7636_ = new_B7644_ & new_B7643_;
  assign new_B7637_ = new_B7642_ & B7626;
  assign new_B7638_ = new_B7647_ & new_B7646_;
  assign new_B7639_ = new_B7645_ & B7626;
  assign new_B7640_ = new_B7648_ | B7625;
  assign new_B7641_ = ~B7626 ^ new_B7638_;
  assign new_B7642_ = ~new_B7651_ | ~new_B7652_;
  assign new_B7643_ = B7627 ^ new_B7634_;
  assign new_B7644_ = new_B7653_ & new_B7646_;
  assign new_B7645_ = ~new_B7655_ | ~new_B7654_;
  assign new_B7646_ = B7627 | B7628;
  assign new_B7647_ = B7627 | new_B7634_;
  assign new_B7648_ = B7626 & new_B7638_;
  assign new_B7649_ = ~B7625 | ~B7626;
  assign new_B7650_ = new_B7634_ & new_B7649_;
  assign new_B7651_ = ~new_B7650_ & ~new_B7634_;
  assign new_B7652_ = new_B7634_ | new_B7649_;
  assign new_B7653_ = ~B7627 | ~B7628;
  assign new_B7654_ = new_B7634_ | new_B7649_;
  assign new_B7655_ = ~new_B7634_ & ~new_B7656_;
  assign new_B7656_ = new_B7634_ & new_B7649_;
  assign new_B7662_ = new_B7668_ & new_B7667_;
  assign new_B7663_ = new_B7670_ | new_B7669_;
  assign new_B7664_ = new_B7672_ | new_B7671_;
  assign new_B7665_ = new_B7667_ & new_B7673_;
  assign new_B7666_ = new_B7667_ & new_B7674_;
  assign new_B7667_ = B7657 ^ B7658;
  assign new_B7668_ = new_B7669_ ^ B7659;
  assign new_B7669_ = new_B7677_ & new_B7676_;
  assign new_B7670_ = new_B7675_ & B7659;
  assign new_B7671_ = new_B7680_ & new_B7679_;
  assign new_B7672_ = new_B7678_ & B7659;
  assign new_B7673_ = new_B7681_ | B7658;
  assign new_B7674_ = ~B7659 ^ new_B7671_;
  assign new_B7675_ = ~new_B7684_ | ~new_B7685_;
  assign new_B7676_ = B7660 ^ new_B7667_;
  assign new_B7677_ = new_B7686_ & new_B7679_;
  assign new_B7678_ = ~new_B7688_ | ~new_B7687_;
  assign new_B7679_ = B7660 | B7661;
  assign new_B7680_ = B7660 | new_B7667_;
  assign new_B7681_ = B7659 & new_B7671_;
  assign new_B7682_ = ~B7658 | ~B7659;
  assign new_B7683_ = new_B7667_ & new_B7682_;
  assign new_B7684_ = ~new_B7683_ & ~new_B7667_;
  assign new_B7685_ = new_B7667_ | new_B7682_;
  assign new_B7686_ = ~B7660 | ~B7661;
  assign new_B7687_ = new_B7667_ | new_B7682_;
  assign new_B7688_ = ~new_B7667_ & ~new_B7689_;
  assign new_B7689_ = new_B7667_ & new_B7682_;
  assign new_B7695_ = new_B7701_ & new_B7700_;
  assign new_B7696_ = new_B7703_ | new_B7702_;
  assign new_B7697_ = new_B7705_ | new_B7704_;
  assign new_B7698_ = new_B7700_ & new_B7706_;
  assign new_B7699_ = new_B7700_ & new_B7707_;
  assign new_B7700_ = B7690 ^ B7691;
  assign new_B7701_ = new_B7702_ ^ B7692;
  assign new_B7702_ = new_B7710_ & new_B7709_;
  assign new_B7703_ = new_B7708_ & B7692;
  assign new_B7704_ = new_B7713_ & new_B7712_;
  assign new_B7705_ = new_B7711_ & B7692;
  assign new_B7706_ = new_B7714_ | B7691;
  assign new_B7707_ = ~B7692 ^ new_B7704_;
  assign new_B7708_ = ~new_B7717_ | ~new_B7718_;
  assign new_B7709_ = B7693 ^ new_B7700_;
  assign new_B7710_ = new_B7719_ & new_B7712_;
  assign new_B7711_ = ~new_B7721_ | ~new_B7720_;
  assign new_B7712_ = B7693 | B7694;
  assign new_B7713_ = B7693 | new_B7700_;
  assign new_B7714_ = B7692 & new_B7704_;
  assign new_B7715_ = ~B7691 | ~B7692;
  assign new_B7716_ = new_B7700_ & new_B7715_;
  assign new_B7717_ = ~new_B7716_ & ~new_B7700_;
  assign new_B7718_ = new_B7700_ | new_B7715_;
  assign new_B7719_ = ~B7693 | ~B7694;
  assign new_B7720_ = new_B7700_ | new_B7715_;
  assign new_B7721_ = ~new_B7700_ & ~new_B7722_;
  assign new_B7722_ = new_B7700_ & new_B7715_;
  assign new_B7728_ = new_B7734_ & new_B7733_;
  assign new_B7729_ = new_B7736_ | new_B7735_;
  assign new_B7730_ = new_B7738_ | new_B7737_;
  assign new_B7731_ = new_B7733_ & new_B7739_;
  assign new_B7732_ = new_B7733_ & new_B7740_;
  assign new_B7733_ = B7723 ^ B7724;
  assign new_B7734_ = new_B7735_ ^ B7725;
  assign new_B7735_ = new_B7743_ & new_B7742_;
  assign new_B7736_ = new_B7741_ & B7725;
  assign new_B7737_ = new_B7746_ & new_B7745_;
  assign new_B7738_ = new_B7744_ & B7725;
  assign new_B7739_ = new_B7747_ | B7724;
  assign new_B7740_ = ~B7725 ^ new_B7737_;
  assign new_B7741_ = ~new_B7750_ | ~new_B7751_;
  assign new_B7742_ = B7726 ^ new_B7733_;
  assign new_B7743_ = new_B7752_ & new_B7745_;
  assign new_B7744_ = ~new_B7754_ | ~new_B7753_;
  assign new_B7745_ = B7726 | B7727;
  assign new_B7746_ = B7726 | new_B7733_;
  assign new_B7747_ = B7725 & new_B7737_;
  assign new_B7748_ = ~B7724 | ~B7725;
  assign new_B7749_ = new_B7733_ & new_B7748_;
  assign new_B7750_ = ~new_B7749_ & ~new_B7733_;
  assign new_B7751_ = new_B7733_ | new_B7748_;
  assign new_B7752_ = ~B7726 | ~B7727;
  assign new_B7753_ = new_B7733_ | new_B7748_;
  assign new_B7754_ = ~new_B7733_ & ~new_B7755_;
  assign new_B7755_ = new_B7733_ & new_B7748_;
  assign new_B7761_ = new_B7767_ & new_B7766_;
  assign new_B7762_ = new_B7769_ | new_B7768_;
  assign new_B7763_ = new_B7771_ | new_B7770_;
  assign new_B7764_ = new_B7766_ & new_B7772_;
  assign new_B7765_ = new_B7766_ & new_B7773_;
  assign new_B7766_ = B7756 ^ B7757;
  assign new_B7767_ = new_B7768_ ^ B7758;
  assign new_B7768_ = new_B7776_ & new_B7775_;
  assign new_B7769_ = new_B7774_ & B7758;
  assign new_B7770_ = new_B7779_ & new_B7778_;
  assign new_B7771_ = new_B7777_ & B7758;
  assign new_B7772_ = new_B7780_ | B7757;
  assign new_B7773_ = ~B7758 ^ new_B7770_;
  assign new_B7774_ = ~new_B7783_ | ~new_B7784_;
  assign new_B7775_ = B7759 ^ new_B7766_;
  assign new_B7776_ = new_B7785_ & new_B7778_;
  assign new_B7777_ = ~new_B7787_ | ~new_B7786_;
  assign new_B7778_ = B7759 | B7760;
  assign new_B7779_ = B7759 | new_B7766_;
  assign new_B7780_ = B7758 & new_B7770_;
  assign new_B7781_ = ~B7757 | ~B7758;
  assign new_B7782_ = new_B7766_ & new_B7781_;
  assign new_B7783_ = ~new_B7782_ & ~new_B7766_;
  assign new_B7784_ = new_B7766_ | new_B7781_;
  assign new_B7785_ = ~B7759 | ~B7760;
  assign new_B7786_ = new_B7766_ | new_B7781_;
  assign new_B7787_ = ~new_B7766_ & ~new_B7788_;
  assign new_B7788_ = new_B7766_ & new_B7781_;
  assign new_B7794_ = new_B7800_ & new_B7799_;
  assign new_B7795_ = new_B7802_ | new_B7801_;
  assign new_B7796_ = new_B7804_ | new_B7803_;
  assign new_B7797_ = new_B7799_ & new_B7805_;
  assign new_B7798_ = new_B7799_ & new_B7806_;
  assign new_B7799_ = B7789 ^ B7790;
  assign new_B7800_ = new_B7801_ ^ B7791;
  assign new_B7801_ = new_B7809_ & new_B7808_;
  assign new_B7802_ = new_B7807_ & B7791;
  assign new_B7803_ = new_B7812_ & new_B7811_;
  assign new_B7804_ = new_B7810_ & B7791;
  assign new_B7805_ = new_B7813_ | B7790;
  assign new_B7806_ = ~B7791 ^ new_B7803_;
  assign new_B7807_ = ~new_B7816_ | ~new_B7817_;
  assign new_B7808_ = B7792 ^ new_B7799_;
  assign new_B7809_ = new_B7818_ & new_B7811_;
  assign new_B7810_ = ~new_B7820_ | ~new_B7819_;
  assign new_B7811_ = B7792 | B7793;
  assign new_B7812_ = B7792 | new_B7799_;
  assign new_B7813_ = B7791 & new_B7803_;
  assign new_B7814_ = ~B7790 | ~B7791;
  assign new_B7815_ = new_B7799_ & new_B7814_;
  assign new_B7816_ = ~new_B7815_ & ~new_B7799_;
  assign new_B7817_ = new_B7799_ | new_B7814_;
  assign new_B7818_ = ~B7792 | ~B7793;
  assign new_B7819_ = new_B7799_ | new_B7814_;
  assign new_B7820_ = ~new_B7799_ & ~new_B7821_;
  assign new_B7821_ = new_B7799_ & new_B7814_;
  assign new_B7827_ = new_B7833_ & new_B7832_;
  assign new_B7828_ = new_B7835_ | new_B7834_;
  assign new_B7829_ = new_B7837_ | new_B7836_;
  assign new_B7830_ = new_B7832_ & new_B7838_;
  assign new_B7831_ = new_B7832_ & new_B7839_;
  assign new_B7832_ = B7822 ^ B7823;
  assign new_B7833_ = new_B7834_ ^ B7824;
  assign new_B7834_ = new_B7842_ & new_B7841_;
  assign new_B7835_ = new_B7840_ & B7824;
  assign new_B7836_ = new_B7845_ & new_B7844_;
  assign new_B7837_ = new_B7843_ & B7824;
  assign new_B7838_ = new_B7846_ | B7823;
  assign new_B7839_ = ~B7824 ^ new_B7836_;
  assign new_B7840_ = ~new_B7849_ | ~new_B7850_;
  assign new_B7841_ = B7825 ^ new_B7832_;
  assign new_B7842_ = new_B7851_ & new_B7844_;
  assign new_B7843_ = ~new_B7853_ | ~new_B7852_;
  assign new_B7844_ = B7825 | B7826;
  assign new_B7845_ = B7825 | new_B7832_;
  assign new_B7846_ = B7824 & new_B7836_;
  assign new_B7847_ = ~B7823 | ~B7824;
  assign new_B7848_ = new_B7832_ & new_B7847_;
  assign new_B7849_ = ~new_B7848_ & ~new_B7832_;
  assign new_B7850_ = new_B7832_ | new_B7847_;
  assign new_B7851_ = ~B7825 | ~B7826;
  assign new_B7852_ = new_B7832_ | new_B7847_;
  assign new_B7853_ = ~new_B7832_ & ~new_B7854_;
  assign new_B7854_ = new_B7832_ & new_B7847_;
  assign new_B7860_ = new_B7866_ & new_B7865_;
  assign new_B7861_ = new_B7868_ | new_B7867_;
  assign new_B7862_ = new_B7870_ | new_B7869_;
  assign new_B7863_ = new_B7865_ & new_B7871_;
  assign new_B7864_ = new_B7865_ & new_B7872_;
  assign new_B7865_ = B7855 ^ B7856;
  assign new_B7866_ = new_B7867_ ^ B7857;
  assign new_B7867_ = new_B7875_ & new_B7874_;
  assign new_B7868_ = new_B7873_ & B7857;
  assign new_B7869_ = new_B7878_ & new_B7877_;
  assign new_B7870_ = new_B7876_ & B7857;
  assign new_B7871_ = new_B7879_ | B7856;
  assign new_B7872_ = ~B7857 ^ new_B7869_;
  assign new_B7873_ = ~new_B7882_ | ~new_B7883_;
  assign new_B7874_ = B7858 ^ new_B7865_;
  assign new_B7875_ = new_B7884_ & new_B7877_;
  assign new_B7876_ = ~new_B7886_ | ~new_B7885_;
  assign new_B7877_ = B7858 | B7859;
  assign new_B7878_ = B7858 | new_B7865_;
  assign new_B7879_ = B7857 & new_B7869_;
  assign new_B7880_ = ~B7856 | ~B7857;
  assign new_B7881_ = new_B7865_ & new_B7880_;
  assign new_B7882_ = ~new_B7881_ & ~new_B7865_;
  assign new_B7883_ = new_B7865_ | new_B7880_;
  assign new_B7884_ = ~B7858 | ~B7859;
  assign new_B7885_ = new_B7865_ | new_B7880_;
  assign new_B7886_ = ~new_B7865_ & ~new_B7887_;
  assign new_B7887_ = new_B7865_ & new_B7880_;
  assign new_B7893_ = new_B7899_ & new_B7898_;
  assign new_B7894_ = new_B7901_ | new_B7900_;
  assign new_B7895_ = new_B7903_ | new_B7902_;
  assign new_B7896_ = new_B7898_ & new_B7904_;
  assign new_B7897_ = new_B7898_ & new_B7905_;
  assign new_B7898_ = B7888 ^ B7889;
  assign new_B7899_ = new_B7900_ ^ B7890;
  assign new_B7900_ = new_B7908_ & new_B7907_;
  assign new_B7901_ = new_B7906_ & B7890;
  assign new_B7902_ = new_B7911_ & new_B7910_;
  assign new_B7903_ = new_B7909_ & B7890;
  assign new_B7904_ = new_B7912_ | B7889;
  assign new_B7905_ = ~B7890 ^ new_B7902_;
  assign new_B7906_ = ~new_B7915_ | ~new_B7916_;
  assign new_B7907_ = B7891 ^ new_B7898_;
  assign new_B7908_ = new_B7917_ & new_B7910_;
  assign new_B7909_ = ~new_B7919_ | ~new_B7918_;
  assign new_B7910_ = B7891 | B7892;
  assign new_B7911_ = B7891 | new_B7898_;
  assign new_B7912_ = B7890 & new_B7902_;
  assign new_B7913_ = ~B7889 | ~B7890;
  assign new_B7914_ = new_B7898_ & new_B7913_;
  assign new_B7915_ = ~new_B7914_ & ~new_B7898_;
  assign new_B7916_ = new_B7898_ | new_B7913_;
  assign new_B7917_ = ~B7891 | ~B7892;
  assign new_B7918_ = new_B7898_ | new_B7913_;
  assign new_B7919_ = ~new_B7898_ & ~new_B7920_;
  assign new_B7920_ = new_B7898_ & new_B7913_;
  assign new_B7926_ = new_B7932_ & new_B7931_;
  assign new_B7927_ = new_B7934_ | new_B7933_;
  assign new_B7928_ = new_B7936_ | new_B7935_;
  assign new_B7929_ = new_B7931_ & new_B7937_;
  assign new_B7930_ = new_B7931_ & new_B7938_;
  assign new_B7931_ = B7921 ^ B7922;
  assign new_B7932_ = new_B7933_ ^ B7923;
  assign new_B7933_ = new_B7941_ & new_B7940_;
  assign new_B7934_ = new_B7939_ & B7923;
  assign new_B7935_ = new_B7944_ & new_B7943_;
  assign new_B7936_ = new_B7942_ & B7923;
  assign new_B7937_ = new_B7945_ | B7922;
  assign new_B7938_ = ~B7923 ^ new_B7935_;
  assign new_B7939_ = ~new_B7948_ | ~new_B7949_;
  assign new_B7940_ = B7924 ^ new_B7931_;
  assign new_B7941_ = new_B7950_ & new_B7943_;
  assign new_B7942_ = ~new_B7952_ | ~new_B7951_;
  assign new_B7943_ = B7924 | B7925;
  assign new_B7944_ = B7924 | new_B7931_;
  assign new_B7945_ = B7923 & new_B7935_;
  assign new_B7946_ = ~B7922 | ~B7923;
  assign new_B7947_ = new_B7931_ & new_B7946_;
  assign new_B7948_ = ~new_B7947_ & ~new_B7931_;
  assign new_B7949_ = new_B7931_ | new_B7946_;
  assign new_B7950_ = ~B7924 | ~B7925;
  assign new_B7951_ = new_B7931_ | new_B7946_;
  assign new_B7952_ = ~new_B7931_ & ~new_B7953_;
  assign new_B7953_ = new_B7931_ & new_B7946_;
  assign new_B7959_ = new_B7965_ & new_B7964_;
  assign new_B7960_ = new_B7967_ | new_B7966_;
  assign new_B7961_ = new_B7969_ | new_B7968_;
  assign new_B7962_ = new_B7964_ & new_B7970_;
  assign new_B7963_ = new_B7964_ & new_B7971_;
  assign new_B7964_ = B7954 ^ B7955;
  assign new_B7965_ = new_B7966_ ^ B7956;
  assign new_B7966_ = new_B7974_ & new_B7973_;
  assign new_B7967_ = new_B7972_ & B7956;
  assign new_B7968_ = new_B7977_ & new_B7976_;
  assign new_B7969_ = new_B7975_ & B7956;
  assign new_B7970_ = new_B7978_ | B7955;
  assign new_B7971_ = ~B7956 ^ new_B7968_;
  assign new_B7972_ = ~new_B7981_ | ~new_B7982_;
  assign new_B7973_ = B7957 ^ new_B7964_;
  assign new_B7974_ = new_B7983_ & new_B7976_;
  assign new_B7975_ = ~new_B7985_ | ~new_B7984_;
  assign new_B7976_ = B7957 | B7958;
  assign new_B7977_ = B7957 | new_B7964_;
  assign new_B7978_ = B7956 & new_B7968_;
  assign new_B7979_ = ~B7955 | ~B7956;
  assign new_B7980_ = new_B7964_ & new_B7979_;
  assign new_B7981_ = ~new_B7980_ & ~new_B7964_;
  assign new_B7982_ = new_B7964_ | new_B7979_;
  assign new_B7983_ = ~B7957 | ~B7958;
  assign new_B7984_ = new_B7964_ | new_B7979_;
  assign new_B7985_ = ~new_B7964_ & ~new_B7986_;
  assign new_B7986_ = new_B7964_ & new_B7979_;
  assign new_B7992_ = new_B7998_ & new_B7997_;
  assign new_B7993_ = new_B8000_ | new_B7999_;
  assign new_B7994_ = new_B8002_ | new_B8001_;
  assign new_B7995_ = new_B7997_ & new_B8003_;
  assign new_B7996_ = new_B7997_ & new_B8004_;
  assign new_B7997_ = B7987 ^ B7988;
  assign new_B7998_ = new_B7999_ ^ B7989;
  assign new_B7999_ = new_B8007_ & new_B8006_;
  assign new_B8000_ = new_B8005_ & B7989;
  assign new_B8001_ = new_B8010_ & new_B8009_;
  assign new_B8002_ = new_B8008_ & B7989;
  assign new_B8003_ = new_B8011_ | B7988;
  assign new_B8004_ = ~B7989 ^ new_B8001_;
  assign new_B8005_ = ~new_B8014_ | ~new_B8015_;
  assign new_B8006_ = B7990 ^ new_B7997_;
  assign new_B8007_ = new_B8016_ & new_B8009_;
  assign new_B8008_ = ~new_B8018_ | ~new_B8017_;
  assign new_B8009_ = B7990 | B7991;
  assign new_B8010_ = B7990 | new_B7997_;
  assign new_B8011_ = B7989 & new_B8001_;
  assign new_B8012_ = ~B7988 | ~B7989;
  assign new_B8013_ = new_B7997_ & new_B8012_;
  assign new_B8014_ = ~new_B8013_ & ~new_B7997_;
  assign new_B8015_ = new_B7997_ | new_B8012_;
  assign new_B8016_ = ~B7990 | ~B7991;
  assign new_B8017_ = new_B7997_ | new_B8012_;
  assign new_B8018_ = ~new_B7997_ & ~new_B8019_;
  assign new_B8019_ = new_B7997_ & new_B8012_;
  assign new_B8025_ = new_B8031_ & new_B8030_;
  assign new_B8026_ = new_B8033_ | new_B8032_;
  assign new_B8027_ = new_B8035_ | new_B8034_;
  assign new_B8028_ = new_B8030_ & new_B8036_;
  assign new_B8029_ = new_B8030_ & new_B8037_;
  assign new_B8030_ = B8020 ^ B8021;
  assign new_B8031_ = new_B8032_ ^ B8022;
  assign new_B8032_ = new_B8040_ & new_B8039_;
  assign new_B8033_ = new_B8038_ & B8022;
  assign new_B8034_ = new_B8043_ & new_B8042_;
  assign new_B8035_ = new_B8041_ & B8022;
  assign new_B8036_ = new_B8044_ | B8021;
  assign new_B8037_ = ~B8022 ^ new_B8034_;
  assign new_B8038_ = ~new_B8047_ | ~new_B8048_;
  assign new_B8039_ = B8023 ^ new_B8030_;
  assign new_B8040_ = new_B8049_ & new_B8042_;
  assign new_B8041_ = ~new_B8051_ | ~new_B8050_;
  assign new_B8042_ = B8023 | B8024;
  assign new_B8043_ = B8023 | new_B8030_;
  assign new_B8044_ = B8022 & new_B8034_;
  assign new_B8045_ = ~B8021 | ~B8022;
  assign new_B8046_ = new_B8030_ & new_B8045_;
  assign new_B8047_ = ~new_B8046_ & ~new_B8030_;
  assign new_B8048_ = new_B8030_ | new_B8045_;
  assign new_B8049_ = ~B8023 | ~B8024;
  assign new_B8050_ = new_B8030_ | new_B8045_;
  assign new_B8051_ = ~new_B8030_ & ~new_B8052_;
  assign new_B8052_ = new_B8030_ & new_B8045_;
  assign new_B8058_ = new_B8064_ & new_B8063_;
  assign new_B8059_ = new_B8066_ | new_B8065_;
  assign new_B8060_ = new_B8068_ | new_B8067_;
  assign new_B8061_ = new_B8063_ & new_B8069_;
  assign new_B8062_ = new_B8063_ & new_B8070_;
  assign new_B8063_ = B8053 ^ B8054;
  assign new_B8064_ = new_B8065_ ^ B8055;
  assign new_B8065_ = new_B8073_ & new_B8072_;
  assign new_B8066_ = new_B8071_ & B8055;
  assign new_B8067_ = new_B8076_ & new_B8075_;
  assign new_B8068_ = new_B8074_ & B8055;
  assign new_B8069_ = new_B8077_ | B8054;
  assign new_B8070_ = ~B8055 ^ new_B8067_;
  assign new_B8071_ = ~new_B8080_ | ~new_B8081_;
  assign new_B8072_ = B8056 ^ new_B8063_;
  assign new_B8073_ = new_B8082_ & new_B8075_;
  assign new_B8074_ = ~new_B8084_ | ~new_B8083_;
  assign new_B8075_ = B8056 | B8057;
  assign new_B8076_ = B8056 | new_B8063_;
  assign new_B8077_ = B8055 & new_B8067_;
  assign new_B8078_ = ~B8054 | ~B8055;
  assign new_B8079_ = new_B8063_ & new_B8078_;
  assign new_B8080_ = ~new_B8079_ & ~new_B8063_;
  assign new_B8081_ = new_B8063_ | new_B8078_;
  assign new_B8082_ = ~B8056 | ~B8057;
  assign new_B8083_ = new_B8063_ | new_B8078_;
  assign new_B8084_ = ~new_B8063_ & ~new_B8085_;
  assign new_B8085_ = new_B8063_ & new_B8078_;
  assign new_B8091_ = new_B8097_ & new_B8096_;
  assign new_B8092_ = new_B8099_ | new_B8098_;
  assign new_B8093_ = new_B8101_ | new_B8100_;
  assign new_B8094_ = new_B8096_ & new_B8102_;
  assign new_B8095_ = new_B8096_ & new_B8103_;
  assign new_B8096_ = B8086 ^ B8087;
  assign new_B8097_ = new_B8098_ ^ B8088;
  assign new_B8098_ = new_B8106_ & new_B8105_;
  assign new_B8099_ = new_B8104_ & B8088;
  assign new_B8100_ = new_B8109_ & new_B8108_;
  assign new_B8101_ = new_B8107_ & B8088;
  assign new_B8102_ = new_B8110_ | B8087;
  assign new_B8103_ = ~B8088 ^ new_B8100_;
  assign new_B8104_ = ~new_B8113_ | ~new_B8114_;
  assign new_B8105_ = B8089 ^ new_B8096_;
  assign new_B8106_ = new_B8115_ & new_B8108_;
  assign new_B8107_ = ~new_B8117_ | ~new_B8116_;
  assign new_B8108_ = B8089 | B8090;
  assign new_B8109_ = B8089 | new_B8096_;
  assign new_B8110_ = B8088 & new_B8100_;
  assign new_B8111_ = ~B8087 | ~B8088;
  assign new_B8112_ = new_B8096_ & new_B8111_;
  assign new_B8113_ = ~new_B8112_ & ~new_B8096_;
  assign new_B8114_ = new_B8096_ | new_B8111_;
  assign new_B8115_ = ~B8089 | ~B8090;
  assign new_B8116_ = new_B8096_ | new_B8111_;
  assign new_B8117_ = ~new_B8096_ & ~new_B8118_;
  assign new_B8118_ = new_B8096_ & new_B8111_;
  assign new_B8124_ = new_B8130_ & new_B8129_;
  assign new_B8125_ = new_B8132_ | new_B8131_;
  assign new_B8126_ = new_B8134_ | new_B8133_;
  assign new_B8127_ = new_B8129_ & new_B8135_;
  assign new_B8128_ = new_B8129_ & new_B8136_;
  assign new_B8129_ = B8119 ^ B8120;
  assign new_B8130_ = new_B8131_ ^ B8121;
  assign new_B8131_ = new_B8139_ & new_B8138_;
  assign new_B8132_ = new_B8137_ & B8121;
  assign new_B8133_ = new_B8142_ & new_B8141_;
  assign new_B8134_ = new_B8140_ & B8121;
  assign new_B8135_ = new_B8143_ | B8120;
  assign new_B8136_ = ~B8121 ^ new_B8133_;
  assign new_B8137_ = ~new_B8146_ | ~new_B8147_;
  assign new_B8138_ = B8122 ^ new_B8129_;
  assign new_B8139_ = new_B8148_ & new_B8141_;
  assign new_B8140_ = ~new_B8150_ | ~new_B8149_;
  assign new_B8141_ = B8122 | B8123;
  assign new_B8142_ = B8122 | new_B8129_;
  assign new_B8143_ = B8121 & new_B8133_;
  assign new_B8144_ = ~B8120 | ~B8121;
  assign new_B8145_ = new_B8129_ & new_B8144_;
  assign new_B8146_ = ~new_B8145_ & ~new_B8129_;
  assign new_B8147_ = new_B8129_ | new_B8144_;
  assign new_B8148_ = ~B8122 | ~B8123;
  assign new_B8149_ = new_B8129_ | new_B8144_;
  assign new_B8150_ = ~new_B8129_ & ~new_B8151_;
  assign new_B8151_ = new_B8129_ & new_B8144_;
  assign new_B8157_ = new_B8163_ & new_B8162_;
  assign new_B8158_ = new_B8165_ | new_B8164_;
  assign new_B8159_ = new_B8167_ | new_B8166_;
  assign new_B8160_ = new_B8162_ & new_B8168_;
  assign new_B8161_ = new_B8162_ & new_B8169_;
  assign new_B8162_ = B8152 ^ B8153;
  assign new_B8163_ = new_B8164_ ^ B8154;
  assign new_B8164_ = new_B8172_ & new_B8171_;
  assign new_B8165_ = new_B8170_ & B8154;
  assign new_B8166_ = new_B8175_ & new_B8174_;
  assign new_B8167_ = new_B8173_ & B8154;
  assign new_B8168_ = new_B8176_ | B8153;
  assign new_B8169_ = ~B8154 ^ new_B8166_;
  assign new_B8170_ = ~new_B8179_ | ~new_B8180_;
  assign new_B8171_ = B8155 ^ new_B8162_;
  assign new_B8172_ = new_B8181_ & new_B8174_;
  assign new_B8173_ = ~new_B8183_ | ~new_B8182_;
  assign new_B8174_ = B8155 | B8156;
  assign new_B8175_ = B8155 | new_B8162_;
  assign new_B8176_ = B8154 & new_B8166_;
  assign new_B8177_ = ~B8153 | ~B8154;
  assign new_B8178_ = new_B8162_ & new_B8177_;
  assign new_B8179_ = ~new_B8178_ & ~new_B8162_;
  assign new_B8180_ = new_B8162_ | new_B8177_;
  assign new_B8181_ = ~B8155 | ~B8156;
  assign new_B8182_ = new_B8162_ | new_B8177_;
  assign new_B8183_ = ~new_B8162_ & ~new_B8184_;
  assign new_B8184_ = new_B8162_ & new_B8177_;
  assign new_B8190_ = new_B8196_ & new_B8195_;
  assign new_B8191_ = new_B8198_ | new_B8197_;
  assign new_B8192_ = new_B8200_ | new_B8199_;
  assign new_B8193_ = new_B8195_ & new_B8201_;
  assign new_B8194_ = new_B8195_ & new_B8202_;
  assign new_B8195_ = B8185 ^ B8186;
  assign new_B8196_ = new_B8197_ ^ B8187;
  assign new_B8197_ = new_B8205_ & new_B8204_;
  assign new_B8198_ = new_B8203_ & B8187;
  assign new_B8199_ = new_B8208_ & new_B8207_;
  assign new_B8200_ = new_B8206_ & B8187;
  assign new_B8201_ = new_B8209_ | B8186;
  assign new_B8202_ = ~B8187 ^ new_B8199_;
  assign new_B8203_ = ~new_B8212_ | ~new_B8213_;
  assign new_B8204_ = B8188 ^ new_B8195_;
  assign new_B8205_ = new_B8214_ & new_B8207_;
  assign new_B8206_ = ~new_B8216_ | ~new_B8215_;
  assign new_B8207_ = B8188 | B8189;
  assign new_B8208_ = B8188 | new_B8195_;
  assign new_B8209_ = B8187 & new_B8199_;
  assign new_B8210_ = ~B8186 | ~B8187;
  assign new_B8211_ = new_B8195_ & new_B8210_;
  assign new_B8212_ = ~new_B8211_ & ~new_B8195_;
  assign new_B8213_ = new_B8195_ | new_B8210_;
  assign new_B8214_ = ~B8188 | ~B8189;
  assign new_B8215_ = new_B8195_ | new_B8210_;
  assign new_B8216_ = ~new_B8195_ & ~new_B8217_;
  assign new_B8217_ = new_B8195_ & new_B8210_;
  assign new_B8223_ = new_B8229_ & new_B8228_;
  assign new_B8224_ = new_B8231_ | new_B8230_;
  assign new_B8225_ = new_B8233_ | new_B8232_;
  assign new_B8226_ = new_B8228_ & new_B8234_;
  assign new_B8227_ = new_B8228_ & new_B8235_;
  assign new_B8228_ = B8218 ^ B8219;
  assign new_B8229_ = new_B8230_ ^ B8220;
  assign new_B8230_ = new_B8238_ & new_B8237_;
  assign new_B8231_ = new_B8236_ & B8220;
  assign new_B8232_ = new_B8241_ & new_B8240_;
  assign new_B8233_ = new_B8239_ & B8220;
  assign new_B8234_ = new_B8242_ | B8219;
  assign new_B8235_ = ~B8220 ^ new_B8232_;
  assign new_B8236_ = ~new_B8245_ | ~new_B8246_;
  assign new_B8237_ = B8221 ^ new_B8228_;
  assign new_B8238_ = new_B8247_ & new_B8240_;
  assign new_B8239_ = ~new_B8249_ | ~new_B8248_;
  assign new_B8240_ = B8221 | B8222;
  assign new_B8241_ = B8221 | new_B8228_;
  assign new_B8242_ = B8220 & new_B8232_;
  assign new_B8243_ = ~B8219 | ~B8220;
  assign new_B8244_ = new_B8228_ & new_B8243_;
  assign new_B8245_ = ~new_B8244_ & ~new_B8228_;
  assign new_B8246_ = new_B8228_ | new_B8243_;
  assign new_B8247_ = ~B8221 | ~B8222;
  assign new_B8248_ = new_B8228_ | new_B8243_;
  assign new_B8249_ = ~new_B8228_ & ~new_B8250_;
  assign new_B8250_ = new_B8228_ & new_B8243_;
  assign new_B8256_ = new_B8262_ & new_B8261_;
  assign new_B8257_ = new_B8264_ | new_B8263_;
  assign new_B8258_ = new_B8266_ | new_B8265_;
  assign new_B8259_ = new_B8261_ & new_B8267_;
  assign new_B8260_ = new_B8261_ & new_B8268_;
  assign new_B8261_ = B8251 ^ B8252;
  assign new_B8262_ = new_B8263_ ^ B8253;
  assign new_B8263_ = new_B8271_ & new_B8270_;
  assign new_B8264_ = new_B8269_ & B8253;
  assign new_B8265_ = new_B8274_ & new_B8273_;
  assign new_B8266_ = new_B8272_ & B8253;
  assign new_B8267_ = new_B8275_ | B8252;
  assign new_B8268_ = ~B8253 ^ new_B8265_;
  assign new_B8269_ = ~new_B8278_ | ~new_B8279_;
  assign new_B8270_ = B8254 ^ new_B8261_;
  assign new_B8271_ = new_B8280_ & new_B8273_;
  assign new_B8272_ = ~new_B8282_ | ~new_B8281_;
  assign new_B8273_ = B8254 | B8255;
  assign new_B8274_ = B8254 | new_B8261_;
  assign new_B8275_ = B8253 & new_B8265_;
  assign new_B8276_ = ~B8252 | ~B8253;
  assign new_B8277_ = new_B8261_ & new_B8276_;
  assign new_B8278_ = ~new_B8277_ & ~new_B8261_;
  assign new_B8279_ = new_B8261_ | new_B8276_;
  assign new_B8280_ = ~B8254 | ~B8255;
  assign new_B8281_ = new_B8261_ | new_B8276_;
  assign new_B8282_ = ~new_B8261_ & ~new_B8283_;
  assign new_B8283_ = new_B8261_ & new_B8276_;
  assign new_B8289_ = new_B8295_ & new_B8294_;
  assign new_B8290_ = new_B8297_ | new_B8296_;
  assign new_B8291_ = new_B8299_ | new_B8298_;
  assign new_B8292_ = new_B8294_ & new_B8300_;
  assign new_B8293_ = new_B8294_ & new_B8301_;
  assign new_B8294_ = B8284 ^ B8285;
  assign new_B8295_ = new_B8296_ ^ B8286;
  assign new_B8296_ = new_B8304_ & new_B8303_;
  assign new_B8297_ = new_B8302_ & B8286;
  assign new_B8298_ = new_B8307_ & new_B8306_;
  assign new_B8299_ = new_B8305_ & B8286;
  assign new_B8300_ = new_B8308_ | B8285;
  assign new_B8301_ = ~B8286 ^ new_B8298_;
  assign new_B8302_ = ~new_B8311_ | ~new_B8312_;
  assign new_B8303_ = B8287 ^ new_B8294_;
  assign new_B8304_ = new_B8313_ & new_B8306_;
  assign new_B8305_ = ~new_B8315_ | ~new_B8314_;
  assign new_B8306_ = B8287 | B8288;
  assign new_B8307_ = B8287 | new_B8294_;
  assign new_B8308_ = B8286 & new_B8298_;
  assign new_B8309_ = ~B8285 | ~B8286;
  assign new_B8310_ = new_B8294_ & new_B8309_;
  assign new_B8311_ = ~new_B8310_ & ~new_B8294_;
  assign new_B8312_ = new_B8294_ | new_B8309_;
  assign new_B8313_ = ~B8287 | ~B8288;
  assign new_B8314_ = new_B8294_ | new_B8309_;
  assign new_B8315_ = ~new_B8294_ & ~new_B8316_;
  assign new_B8316_ = new_B8294_ & new_B8309_;
  assign new_B8322_ = new_B8328_ & new_B8327_;
  assign new_B8323_ = new_B8330_ | new_B8329_;
  assign new_B8324_ = new_B8332_ | new_B8331_;
  assign new_B8325_ = new_B8327_ & new_B8333_;
  assign new_B8326_ = new_B8327_ & new_B8334_;
  assign new_B8327_ = B8317 ^ B8318;
  assign new_B8328_ = new_B8329_ ^ B8319;
  assign new_B8329_ = new_B8337_ & new_B8336_;
  assign new_B8330_ = new_B8335_ & B8319;
  assign new_B8331_ = new_B8340_ & new_B8339_;
  assign new_B8332_ = new_B8338_ & B8319;
  assign new_B8333_ = new_B8341_ | B8318;
  assign new_B8334_ = ~B8319 ^ new_B8331_;
  assign new_B8335_ = ~new_B8344_ | ~new_B8345_;
  assign new_B8336_ = B8320 ^ new_B8327_;
  assign new_B8337_ = new_B8346_ & new_B8339_;
  assign new_B8338_ = ~new_B8348_ | ~new_B8347_;
  assign new_B8339_ = B8320 | B8321;
  assign new_B8340_ = B8320 | new_B8327_;
  assign new_B8341_ = B8319 & new_B8331_;
  assign new_B8342_ = ~B8318 | ~B8319;
  assign new_B8343_ = new_B8327_ & new_B8342_;
  assign new_B8344_ = ~new_B8343_ & ~new_B8327_;
  assign new_B8345_ = new_B8327_ | new_B8342_;
  assign new_B8346_ = ~B8320 | ~B8321;
  assign new_B8347_ = new_B8327_ | new_B8342_;
  assign new_B8348_ = ~new_B8327_ & ~new_B8349_;
  assign new_B8349_ = new_B8327_ & new_B8342_;
  assign new_B8355_ = new_B8361_ & new_B8360_;
  assign new_B8356_ = new_B8363_ | new_B8362_;
  assign new_B8357_ = new_B8365_ | new_B8364_;
  assign new_B8358_ = new_B8360_ & new_B8366_;
  assign new_B8359_ = new_B8360_ & new_B8367_;
  assign new_B8360_ = B8350 ^ B8351;
  assign new_B8361_ = new_B8362_ ^ B8352;
  assign new_B8362_ = new_B8370_ & new_B8369_;
  assign new_B8363_ = new_B8368_ & B8352;
  assign new_B8364_ = new_B8373_ & new_B8372_;
  assign new_B8365_ = new_B8371_ & B8352;
  assign new_B8366_ = new_B8374_ | B8351;
  assign new_B8367_ = ~B8352 ^ new_B8364_;
  assign new_B8368_ = ~new_B8377_ | ~new_B8378_;
  assign new_B8369_ = B8353 ^ new_B8360_;
  assign new_B8370_ = new_B8379_ & new_B8372_;
  assign new_B8371_ = ~new_B8381_ | ~new_B8380_;
  assign new_B8372_ = B8353 | B8354;
  assign new_B8373_ = B8353 | new_B8360_;
  assign new_B8374_ = B8352 & new_B8364_;
  assign new_B8375_ = ~B8351 | ~B8352;
  assign new_B8376_ = new_B8360_ & new_B8375_;
  assign new_B8377_ = ~new_B8376_ & ~new_B8360_;
  assign new_B8378_ = new_B8360_ | new_B8375_;
  assign new_B8379_ = ~B8353 | ~B8354;
  assign new_B8380_ = new_B8360_ | new_B8375_;
  assign new_B8381_ = ~new_B8360_ & ~new_B8382_;
  assign new_B8382_ = new_B8360_ & new_B8375_;
  assign new_B8388_ = new_B8394_ & new_B8393_;
  assign new_B8389_ = new_B8396_ | new_B8395_;
  assign new_B8390_ = new_B8398_ | new_B8397_;
  assign new_B8391_ = new_B8393_ & new_B8399_;
  assign new_B8392_ = new_B8393_ & new_B8400_;
  assign new_B8393_ = B8383 ^ B8384;
  assign new_B8394_ = new_B8395_ ^ B8385;
  assign new_B8395_ = new_B8403_ & new_B8402_;
  assign new_B8396_ = new_B8401_ & B8385;
  assign new_B8397_ = new_B8406_ & new_B8405_;
  assign new_B8398_ = new_B8404_ & B8385;
  assign new_B8399_ = new_B8407_ | B8384;
  assign new_B8400_ = ~B8385 ^ new_B8397_;
  assign new_B8401_ = ~new_B8410_ | ~new_B8411_;
  assign new_B8402_ = B8386 ^ new_B8393_;
  assign new_B8403_ = new_B8412_ & new_B8405_;
  assign new_B8404_ = ~new_B8414_ | ~new_B8413_;
  assign new_B8405_ = B8386 | B8387;
  assign new_B8406_ = B8386 | new_B8393_;
  assign new_B8407_ = B8385 & new_B8397_;
  assign new_B8408_ = ~B8384 | ~B8385;
  assign new_B8409_ = new_B8393_ & new_B8408_;
  assign new_B8410_ = ~new_B8409_ & ~new_B8393_;
  assign new_B8411_ = new_B8393_ | new_B8408_;
  assign new_B8412_ = ~B8386 | ~B8387;
  assign new_B8413_ = new_B8393_ | new_B8408_;
  assign new_B8414_ = ~new_B8393_ & ~new_B8415_;
  assign new_B8415_ = new_B8393_ & new_B8408_;
  assign new_B8421_ = new_B8427_ & new_B8426_;
  assign new_B8422_ = new_B8429_ | new_B8428_;
  assign new_B8423_ = new_B8431_ | new_B8430_;
  assign new_B8424_ = new_B8426_ & new_B8432_;
  assign new_B8425_ = new_B8426_ & new_B8433_;
  assign new_B8426_ = B8416 ^ B8417;
  assign new_B8427_ = new_B8428_ ^ B8418;
  assign new_B8428_ = new_B8436_ & new_B8435_;
  assign new_B8429_ = new_B8434_ & B8418;
  assign new_B8430_ = new_B8439_ & new_B8438_;
  assign new_B8431_ = new_B8437_ & B8418;
  assign new_B8432_ = new_B8440_ | B8417;
  assign new_B8433_ = ~B8418 ^ new_B8430_;
  assign new_B8434_ = ~new_B8443_ | ~new_B8444_;
  assign new_B8435_ = B8419 ^ new_B8426_;
  assign new_B8436_ = new_B8445_ & new_B8438_;
  assign new_B8437_ = ~new_B8447_ | ~new_B8446_;
  assign new_B8438_ = B8419 | B8420;
  assign new_B8439_ = B8419 | new_B8426_;
  assign new_B8440_ = B8418 & new_B8430_;
  assign new_B8441_ = ~B8417 | ~B8418;
  assign new_B8442_ = new_B8426_ & new_B8441_;
  assign new_B8443_ = ~new_B8442_ & ~new_B8426_;
  assign new_B8444_ = new_B8426_ | new_B8441_;
  assign new_B8445_ = ~B8419 | ~B8420;
  assign new_B8446_ = new_B8426_ | new_B8441_;
  assign new_B8447_ = ~new_B8426_ & ~new_B8448_;
  assign new_B8448_ = new_B8426_ & new_B8441_;
  assign new_B8454_ = new_B8460_ & new_B8459_;
  assign new_B8455_ = new_B8462_ | new_B8461_;
  assign new_B8456_ = new_B8464_ | new_B8463_;
  assign new_B8457_ = new_B8459_ & new_B8465_;
  assign new_B8458_ = new_B8459_ & new_B8466_;
  assign new_B8459_ = B8449 ^ B8450;
  assign new_B8460_ = new_B8461_ ^ B8451;
  assign new_B8461_ = new_B8469_ & new_B8468_;
  assign new_B8462_ = new_B8467_ & B8451;
  assign new_B8463_ = new_B8472_ & new_B8471_;
  assign new_B8464_ = new_B8470_ & B8451;
  assign new_B8465_ = new_B8473_ | B8450;
  assign new_B8466_ = ~B8451 ^ new_B8463_;
  assign new_B8467_ = ~new_B8476_ | ~new_B8477_;
  assign new_B8468_ = B8452 ^ new_B8459_;
  assign new_B8469_ = new_B8478_ & new_B8471_;
  assign new_B8470_ = ~new_B8480_ | ~new_B8479_;
  assign new_B8471_ = B8452 | B8453;
  assign new_B8472_ = B8452 | new_B8459_;
  assign new_B8473_ = B8451 & new_B8463_;
  assign new_B8474_ = ~B8450 | ~B8451;
  assign new_B8475_ = new_B8459_ & new_B8474_;
  assign new_B8476_ = ~new_B8475_ & ~new_B8459_;
  assign new_B8477_ = new_B8459_ | new_B8474_;
  assign new_B8478_ = ~B8452 | ~B8453;
  assign new_B8479_ = new_B8459_ | new_B8474_;
  assign new_B8480_ = ~new_B8459_ & ~new_B8481_;
  assign new_B8481_ = new_B8459_ & new_B8474_;
  assign new_B8487_ = new_B8493_ & new_B8492_;
  assign new_B8488_ = new_B8495_ | new_B8494_;
  assign new_B8489_ = new_B8497_ | new_B8496_;
  assign new_B8490_ = new_B8492_ & new_B8498_;
  assign new_B8491_ = new_B8492_ & new_B8499_;
  assign new_B8492_ = B8482 ^ B8483;
  assign new_B8493_ = new_B8494_ ^ B8484;
  assign new_B8494_ = new_B8502_ & new_B8501_;
  assign new_B8495_ = new_B8500_ & B8484;
  assign new_B8496_ = new_B8505_ & new_B8504_;
  assign new_B8497_ = new_B8503_ & B8484;
  assign new_B8498_ = new_B8506_ | B8483;
  assign new_B8499_ = ~B8484 ^ new_B8496_;
  assign new_B8500_ = ~new_B8509_ | ~new_B8510_;
  assign new_B8501_ = B8485 ^ new_B8492_;
  assign new_B8502_ = new_B8511_ & new_B8504_;
  assign new_B8503_ = ~new_B8513_ | ~new_B8512_;
  assign new_B8504_ = B8485 | B8486;
  assign new_B8505_ = B8485 | new_B8492_;
  assign new_B8506_ = B8484 & new_B8496_;
  assign new_B8507_ = ~B8483 | ~B8484;
  assign new_B8508_ = new_B8492_ & new_B8507_;
  assign new_B8509_ = ~new_B8508_ & ~new_B8492_;
  assign new_B8510_ = new_B8492_ | new_B8507_;
  assign new_B8511_ = ~B8485 | ~B8486;
  assign new_B8512_ = new_B8492_ | new_B8507_;
  assign new_B8513_ = ~new_B8492_ & ~new_B8514_;
  assign new_B8514_ = new_B8492_ & new_B8507_;
  assign new_B8520_ = new_B8526_ & new_B8525_;
  assign new_B8521_ = new_B8528_ | new_B8527_;
  assign new_B8522_ = new_B8530_ | new_B8529_;
  assign new_B8523_ = new_B8525_ & new_B8531_;
  assign new_B8524_ = new_B8525_ & new_B8532_;
  assign new_B8525_ = B8515 ^ B8516;
  assign new_B8526_ = new_B8527_ ^ B8517;
  assign new_B8527_ = new_B8535_ & new_B8534_;
  assign new_B8528_ = new_B8533_ & B8517;
  assign new_B8529_ = new_B8538_ & new_B8537_;
  assign new_B8530_ = new_B8536_ & B8517;
  assign new_B8531_ = new_B8539_ | B8516;
  assign new_B8532_ = ~B8517 ^ new_B8529_;
  assign new_B8533_ = ~new_B8542_ | ~new_B8543_;
  assign new_B8534_ = B8518 ^ new_B8525_;
  assign new_B8535_ = new_B8544_ & new_B8537_;
  assign new_B8536_ = ~new_B8546_ | ~new_B8545_;
  assign new_B8537_ = B8518 | B8519;
  assign new_B8538_ = B8518 | new_B8525_;
  assign new_B8539_ = B8517 & new_B8529_;
  assign new_B8540_ = ~B8516 | ~B8517;
  assign new_B8541_ = new_B8525_ & new_B8540_;
  assign new_B8542_ = ~new_B8541_ & ~new_B8525_;
  assign new_B8543_ = new_B8525_ | new_B8540_;
  assign new_B8544_ = ~B8518 | ~B8519;
  assign new_B8545_ = new_B8525_ | new_B8540_;
  assign new_B8546_ = ~new_B8525_ & ~new_B8547_;
  assign new_B8547_ = new_B8525_ & new_B8540_;
  assign new_B8553_ = new_B8559_ & new_B8558_;
  assign new_B8554_ = new_B8561_ | new_B8560_;
  assign new_B8555_ = new_B8563_ | new_B8562_;
  assign new_B8556_ = new_B8558_ & new_B8564_;
  assign new_B8557_ = new_B8558_ & new_B8565_;
  assign new_B8558_ = B8548 ^ B8549;
  assign new_B8559_ = new_B8560_ ^ B8550;
  assign new_B8560_ = new_B8568_ & new_B8567_;
  assign new_B8561_ = new_B8566_ & B8550;
  assign new_B8562_ = new_B8571_ & new_B8570_;
  assign new_B8563_ = new_B8569_ & B8550;
  assign new_B8564_ = new_B8572_ | B8549;
  assign new_B8565_ = ~B8550 ^ new_B8562_;
  assign new_B8566_ = ~new_B8575_ | ~new_B8576_;
  assign new_B8567_ = B8551 ^ new_B8558_;
  assign new_B8568_ = new_B8577_ & new_B8570_;
  assign new_B8569_ = ~new_B8579_ | ~new_B8578_;
  assign new_B8570_ = B8551 | B8552;
  assign new_B8571_ = B8551 | new_B8558_;
  assign new_B8572_ = B8550 & new_B8562_;
  assign new_B8573_ = ~B8549 | ~B8550;
  assign new_B8574_ = new_B8558_ & new_B8573_;
  assign new_B8575_ = ~new_B8574_ & ~new_B8558_;
  assign new_B8576_ = new_B8558_ | new_B8573_;
  assign new_B8577_ = ~B8551 | ~B8552;
  assign new_B8578_ = new_B8558_ | new_B8573_;
  assign new_B8579_ = ~new_B8558_ & ~new_B8580_;
  assign new_B8580_ = new_B8558_ & new_B8573_;
  assign new_B8586_ = new_B8592_ & new_B8591_;
  assign new_B8587_ = new_B8594_ | new_B8593_;
  assign new_B8588_ = new_B8596_ | new_B8595_;
  assign new_B8589_ = new_B8591_ & new_B8597_;
  assign new_B8590_ = new_B8591_ & new_B8598_;
  assign new_B8591_ = B8581 ^ B8582;
  assign new_B8592_ = new_B8593_ ^ B8583;
  assign new_B8593_ = new_B8601_ & new_B8600_;
  assign new_B8594_ = new_B8599_ & B8583;
  assign new_B8595_ = new_B8604_ & new_B8603_;
  assign new_B8596_ = new_B8602_ & B8583;
  assign new_B8597_ = new_B8605_ | B8582;
  assign new_B8598_ = ~B8583 ^ new_B8595_;
  assign new_B8599_ = ~new_B8608_ | ~new_B8609_;
  assign new_B8600_ = B8584 ^ new_B8591_;
  assign new_B8601_ = new_B8610_ & new_B8603_;
  assign new_B8602_ = ~new_B8612_ | ~new_B8611_;
  assign new_B8603_ = B8584 | B8585;
  assign new_B8604_ = B8584 | new_B8591_;
  assign new_B8605_ = B8583 & new_B8595_;
  assign new_B8606_ = ~B8582 | ~B8583;
  assign new_B8607_ = new_B8591_ & new_B8606_;
  assign new_B8608_ = ~new_B8607_ & ~new_B8591_;
  assign new_B8609_ = new_B8591_ | new_B8606_;
  assign new_B8610_ = ~B8584 | ~B8585;
  assign new_B8611_ = new_B8591_ | new_B8606_;
  assign new_B8612_ = ~new_B8591_ & ~new_B8613_;
  assign new_B8613_ = new_B8591_ & new_B8606_;
  assign new_B8619_ = new_B8625_ & new_B8624_;
  assign new_B8620_ = new_B8627_ | new_B8626_;
  assign new_B8621_ = new_B8629_ | new_B8628_;
  assign new_B8622_ = new_B8624_ & new_B8630_;
  assign new_B8623_ = new_B8624_ & new_B8631_;
  assign new_B8624_ = B8614 ^ B8615;
  assign new_B8625_ = new_B8626_ ^ B8616;
  assign new_B8626_ = new_B8634_ & new_B8633_;
  assign new_B8627_ = new_B8632_ & B8616;
  assign new_B8628_ = new_B8637_ & new_B8636_;
  assign new_B8629_ = new_B8635_ & B8616;
  assign new_B8630_ = new_B8638_ | B8615;
  assign new_B8631_ = ~B8616 ^ new_B8628_;
  assign new_B8632_ = ~new_B8641_ | ~new_B8642_;
  assign new_B8633_ = B8617 ^ new_B8624_;
  assign new_B8634_ = new_B8643_ & new_B8636_;
  assign new_B8635_ = ~new_B8645_ | ~new_B8644_;
  assign new_B8636_ = B8617 | B8618;
  assign new_B8637_ = B8617 | new_B8624_;
  assign new_B8638_ = B8616 & new_B8628_;
  assign new_B8639_ = ~B8615 | ~B8616;
  assign new_B8640_ = new_B8624_ & new_B8639_;
  assign new_B8641_ = ~new_B8640_ & ~new_B8624_;
  assign new_B8642_ = new_B8624_ | new_B8639_;
  assign new_B8643_ = ~B8617 | ~B8618;
  assign new_B8644_ = new_B8624_ | new_B8639_;
  assign new_B8645_ = ~new_B8624_ & ~new_B8646_;
  assign new_B8646_ = new_B8624_ & new_B8639_;
  assign new_B8652_ = new_B8658_ & new_B8657_;
  assign new_B8653_ = new_B8660_ | new_B8659_;
  assign new_B8654_ = new_B8662_ | new_B8661_;
  assign new_B8655_ = new_B8657_ & new_B8663_;
  assign new_B8656_ = new_B8657_ & new_B8664_;
  assign new_B8657_ = B8647 ^ B8648;
  assign new_B8658_ = new_B8659_ ^ B8649;
  assign new_B8659_ = new_B8667_ & new_B8666_;
  assign new_B8660_ = new_B8665_ & B8649;
  assign new_B8661_ = new_B8670_ & new_B8669_;
  assign new_B8662_ = new_B8668_ & B8649;
  assign new_B8663_ = new_B8671_ | B8648;
  assign new_B8664_ = ~B8649 ^ new_B8661_;
  assign new_B8665_ = ~new_B8674_ | ~new_B8675_;
  assign new_B8666_ = B8650 ^ new_B8657_;
  assign new_B8667_ = new_B8676_ & new_B8669_;
  assign new_B8668_ = ~new_B8678_ | ~new_B8677_;
  assign new_B8669_ = B8650 | B8651;
  assign new_B8670_ = B8650 | new_B8657_;
  assign new_B8671_ = B8649 & new_B8661_;
  assign new_B8672_ = ~B8648 | ~B8649;
  assign new_B8673_ = new_B8657_ & new_B8672_;
  assign new_B8674_ = ~new_B8673_ & ~new_B8657_;
  assign new_B8675_ = new_B8657_ | new_B8672_;
  assign new_B8676_ = ~B8650 | ~B8651;
  assign new_B8677_ = new_B8657_ | new_B8672_;
  assign new_B8678_ = ~new_B8657_ & ~new_B8679_;
  assign new_B8679_ = new_B8657_ & new_B8672_;
  assign new_B8685_ = new_B8691_ & new_B8690_;
  assign new_B8686_ = new_B8693_ | new_B8692_;
  assign new_B8687_ = new_B8695_ | new_B8694_;
  assign new_B8688_ = new_B8690_ & new_B8696_;
  assign new_B8689_ = new_B8690_ & new_B8697_;
  assign new_B8690_ = B8680 ^ B8681;
  assign new_B8691_ = new_B8692_ ^ B8682;
  assign new_B8692_ = new_B8700_ & new_B8699_;
  assign new_B8693_ = new_B8698_ & B8682;
  assign new_B8694_ = new_B8703_ & new_B8702_;
  assign new_B8695_ = new_B8701_ & B8682;
  assign new_B8696_ = new_B8704_ | B8681;
  assign new_B8697_ = ~B8682 ^ new_B8694_;
  assign new_B8698_ = ~new_B8707_ | ~new_B8708_;
  assign new_B8699_ = B8683 ^ new_B8690_;
  assign new_B8700_ = new_B8709_ & new_B8702_;
  assign new_B8701_ = ~new_B8711_ | ~new_B8710_;
  assign new_B8702_ = B8683 | B8684;
  assign new_B8703_ = B8683 | new_B8690_;
  assign new_B8704_ = B8682 & new_B8694_;
  assign new_B8705_ = ~B8681 | ~B8682;
  assign new_B8706_ = new_B8690_ & new_B8705_;
  assign new_B8707_ = ~new_B8706_ & ~new_B8690_;
  assign new_B8708_ = new_B8690_ | new_B8705_;
  assign new_B8709_ = ~B8683 | ~B8684;
  assign new_B8710_ = new_B8690_ | new_B8705_;
  assign new_B8711_ = ~new_B8690_ & ~new_B8712_;
  assign new_B8712_ = new_B8690_ & new_B8705_;
  assign new_B8718_ = new_B8724_ & new_B8723_;
  assign new_B8719_ = new_B8726_ | new_B8725_;
  assign new_B8720_ = new_B8728_ | new_B8727_;
  assign new_B8721_ = new_B8723_ & new_B8729_;
  assign new_B8722_ = new_B8723_ & new_B8730_;
  assign new_B8723_ = B8713 ^ B8714;
  assign new_B8724_ = new_B8725_ ^ B8715;
  assign new_B8725_ = new_B8733_ & new_B8732_;
  assign new_B8726_ = new_B8731_ & B8715;
  assign new_B8727_ = new_B8736_ & new_B8735_;
  assign new_B8728_ = new_B8734_ & B8715;
  assign new_B8729_ = new_B8737_ | B8714;
  assign new_B8730_ = ~B8715 ^ new_B8727_;
  assign new_B8731_ = ~new_B8740_ | ~new_B8741_;
  assign new_B8732_ = B8716 ^ new_B8723_;
  assign new_B8733_ = new_B8742_ & new_B8735_;
  assign new_B8734_ = ~new_B8744_ | ~new_B8743_;
  assign new_B8735_ = B8716 | B8717;
  assign new_B8736_ = B8716 | new_B8723_;
  assign new_B8737_ = B8715 & new_B8727_;
  assign new_B8738_ = ~B8714 | ~B8715;
  assign new_B8739_ = new_B8723_ & new_B8738_;
  assign new_B8740_ = ~new_B8739_ & ~new_B8723_;
  assign new_B8741_ = new_B8723_ | new_B8738_;
  assign new_B8742_ = ~B8716 | ~B8717;
  assign new_B8743_ = new_B8723_ | new_B8738_;
  assign new_B8744_ = ~new_B8723_ & ~new_B8745_;
  assign new_B8745_ = new_B8723_ & new_B8738_;
  assign new_B8751_ = new_B8757_ & new_B8756_;
  assign new_B8752_ = new_B8759_ | new_B8758_;
  assign new_B8753_ = new_B8761_ | new_B8760_;
  assign new_B8754_ = new_B8756_ & new_B8762_;
  assign new_B8755_ = new_B8756_ & new_B8763_;
  assign new_B8756_ = B8746 ^ B8747;
  assign new_B8757_ = new_B8758_ ^ B8748;
  assign new_B8758_ = new_B8766_ & new_B8765_;
  assign new_B8759_ = new_B8764_ & B8748;
  assign new_B8760_ = new_B8769_ & new_B8768_;
  assign new_B8761_ = new_B8767_ & B8748;
  assign new_B8762_ = new_B8770_ | B8747;
  assign new_B8763_ = ~B8748 ^ new_B8760_;
  assign new_B8764_ = ~new_B8773_ | ~new_B8774_;
  assign new_B8765_ = B8749 ^ new_B8756_;
  assign new_B8766_ = new_B8775_ & new_B8768_;
  assign new_B8767_ = ~new_B8777_ | ~new_B8776_;
  assign new_B8768_ = B8749 | B8750;
  assign new_B8769_ = B8749 | new_B8756_;
  assign new_B8770_ = B8748 & new_B8760_;
  assign new_B8771_ = ~B8747 | ~B8748;
  assign new_B8772_ = new_B8756_ & new_B8771_;
  assign new_B8773_ = ~new_B8772_ & ~new_B8756_;
  assign new_B8774_ = new_B8756_ | new_B8771_;
  assign new_B8775_ = ~B8749 | ~B8750;
  assign new_B8776_ = new_B8756_ | new_B8771_;
  assign new_B8777_ = ~new_B8756_ & ~new_B8778_;
  assign new_B8778_ = new_B8756_ & new_B8771_;
  assign new_B8784_ = new_B8790_ & new_B8789_;
  assign new_B8785_ = new_B8792_ | new_B8791_;
  assign new_B8786_ = new_B8794_ | new_B8793_;
  assign new_B8787_ = new_B8789_ & new_B8795_;
  assign new_B8788_ = new_B8789_ & new_B8796_;
  assign new_B8789_ = B8779 ^ B8780;
  assign new_B8790_ = new_B8791_ ^ B8781;
  assign new_B8791_ = new_B8799_ & new_B8798_;
  assign new_B8792_ = new_B8797_ & B8781;
  assign new_B8793_ = new_B8802_ & new_B8801_;
  assign new_B8794_ = new_B8800_ & B8781;
  assign new_B8795_ = new_B8803_ | B8780;
  assign new_B8796_ = ~B8781 ^ new_B8793_;
  assign new_B8797_ = ~new_B8806_ | ~new_B8807_;
  assign new_B8798_ = B8782 ^ new_B8789_;
  assign new_B8799_ = new_B8808_ & new_B8801_;
  assign new_B8800_ = ~new_B8810_ | ~new_B8809_;
  assign new_B8801_ = B8782 | B8783;
  assign new_B8802_ = B8782 | new_B8789_;
  assign new_B8803_ = B8781 & new_B8793_;
  assign new_B8804_ = ~B8780 | ~B8781;
  assign new_B8805_ = new_B8789_ & new_B8804_;
  assign new_B8806_ = ~new_B8805_ & ~new_B8789_;
  assign new_B8807_ = new_B8789_ | new_B8804_;
  assign new_B8808_ = ~B8782 | ~B8783;
  assign new_B8809_ = new_B8789_ | new_B8804_;
  assign new_B8810_ = ~new_B8789_ & ~new_B8811_;
  assign new_B8811_ = new_B8789_ & new_B8804_;
  assign new_B8817_ = new_B8823_ & new_B8822_;
  assign new_B8818_ = new_B8825_ | new_B8824_;
  assign new_B8819_ = new_B8827_ | new_B8826_;
  assign new_B8820_ = new_B8822_ & new_B8828_;
  assign new_B8821_ = new_B8822_ & new_B8829_;
  assign new_B8822_ = B8812 ^ B8813;
  assign new_B8823_ = new_B8824_ ^ B8814;
  assign new_B8824_ = new_B8832_ & new_B8831_;
  assign new_B8825_ = new_B8830_ & B8814;
  assign new_B8826_ = new_B8835_ & new_B8834_;
  assign new_B8827_ = new_B8833_ & B8814;
  assign new_B8828_ = new_B8836_ | B8813;
  assign new_B8829_ = ~B8814 ^ new_B8826_;
  assign new_B8830_ = ~new_B8839_ | ~new_B8840_;
  assign new_B8831_ = B8815 ^ new_B8822_;
  assign new_B8832_ = new_B8841_ & new_B8834_;
  assign new_B8833_ = ~new_B8843_ | ~new_B8842_;
  assign new_B8834_ = B8815 | B8816;
  assign new_B8835_ = B8815 | new_B8822_;
  assign new_B8836_ = B8814 & new_B8826_;
  assign new_B8837_ = ~B8813 | ~B8814;
  assign new_B8838_ = new_B8822_ & new_B8837_;
  assign new_B8839_ = ~new_B8838_ & ~new_B8822_;
  assign new_B8840_ = new_B8822_ | new_B8837_;
  assign new_B8841_ = ~B8815 | ~B8816;
  assign new_B8842_ = new_B8822_ | new_B8837_;
  assign new_B8843_ = ~new_B8822_ & ~new_B8844_;
  assign new_B8844_ = new_B8822_ & new_B8837_;
  assign new_B8850_ = new_B8856_ & new_B8855_;
  assign new_B8851_ = new_B8858_ | new_B8857_;
  assign new_B8852_ = new_B8860_ | new_B8859_;
  assign new_B8853_ = new_B8855_ & new_B8861_;
  assign new_B8854_ = new_B8855_ & new_B8862_;
  assign new_B8855_ = B8845 ^ B8846;
  assign new_B8856_ = new_B8857_ ^ B8847;
  assign new_B8857_ = new_B8865_ & new_B8864_;
  assign new_B8858_ = new_B8863_ & B8847;
  assign new_B8859_ = new_B8868_ & new_B8867_;
  assign new_B8860_ = new_B8866_ & B8847;
  assign new_B8861_ = new_B8869_ | B8846;
  assign new_B8862_ = ~B8847 ^ new_B8859_;
  assign new_B8863_ = ~new_B8872_ | ~new_B8873_;
  assign new_B8864_ = B8848 ^ new_B8855_;
  assign new_B8865_ = new_B8874_ & new_B8867_;
  assign new_B8866_ = ~new_B8876_ | ~new_B8875_;
  assign new_B8867_ = B8848 | B8849;
  assign new_B8868_ = B8848 | new_B8855_;
  assign new_B8869_ = B8847 & new_B8859_;
  assign new_B8870_ = ~B8846 | ~B8847;
  assign new_B8871_ = new_B8855_ & new_B8870_;
  assign new_B8872_ = ~new_B8871_ & ~new_B8855_;
  assign new_B8873_ = new_B8855_ | new_B8870_;
  assign new_B8874_ = ~B8848 | ~B8849;
  assign new_B8875_ = new_B8855_ | new_B8870_;
  assign new_B8876_ = ~new_B8855_ & ~new_B8877_;
  assign new_B8877_ = new_B8855_ & new_B8870_;
  assign new_B8883_ = new_B8889_ & new_B8888_;
  assign new_B8884_ = new_B8891_ | new_B8890_;
  assign new_B8885_ = new_B8893_ | new_B8892_;
  assign new_B8886_ = new_B8888_ & new_B8894_;
  assign new_B8887_ = new_B8888_ & new_B8895_;
  assign new_B8888_ = B8878 ^ B8879;
  assign new_B8889_ = new_B8890_ ^ B8880;
  assign new_B8890_ = new_B8898_ & new_B8897_;
  assign new_B8891_ = new_B8896_ & B8880;
  assign new_B8892_ = new_B8901_ & new_B8900_;
  assign new_B8893_ = new_B8899_ & B8880;
  assign new_B8894_ = new_B8902_ | B8879;
  assign new_B8895_ = ~B8880 ^ new_B8892_;
  assign new_B8896_ = ~new_B8905_ | ~new_B8906_;
  assign new_B8897_ = B8881 ^ new_B8888_;
  assign new_B8898_ = new_B8907_ & new_B8900_;
  assign new_B8899_ = ~new_B8909_ | ~new_B8908_;
  assign new_B8900_ = B8881 | B8882;
  assign new_B8901_ = B8881 | new_B8888_;
  assign new_B8902_ = B8880 & new_B8892_;
  assign new_B8903_ = ~B8879 | ~B8880;
  assign new_B8904_ = new_B8888_ & new_B8903_;
  assign new_B8905_ = ~new_B8904_ & ~new_B8888_;
  assign new_B8906_ = new_B8888_ | new_B8903_;
  assign new_B8907_ = ~B8881 | ~B8882;
  assign new_B8908_ = new_B8888_ | new_B8903_;
  assign new_B8909_ = ~new_B8888_ & ~new_B8910_;
  assign new_B8910_ = new_B8888_ & new_B8903_;
  assign new_B8916_ = new_B8922_ & new_B8921_;
  assign new_B8917_ = new_B8924_ | new_B8923_;
  assign new_B8918_ = new_B8926_ | new_B8925_;
  assign new_B8919_ = new_B8921_ & new_B8927_;
  assign new_B8920_ = new_B8921_ & new_B8928_;
  assign new_B8921_ = B8911 ^ B8912;
  assign new_B8922_ = new_B8923_ ^ B8913;
  assign new_B8923_ = new_B8931_ & new_B8930_;
  assign new_B8924_ = new_B8929_ & B8913;
  assign new_B8925_ = new_B8934_ & new_B8933_;
  assign new_B8926_ = new_B8932_ & B8913;
  assign new_B8927_ = new_B8935_ | B8912;
  assign new_B8928_ = ~B8913 ^ new_B8925_;
  assign new_B8929_ = ~new_B8938_ | ~new_B8939_;
  assign new_B8930_ = B8914 ^ new_B8921_;
  assign new_B8931_ = new_B8940_ & new_B8933_;
  assign new_B8932_ = ~new_B8942_ | ~new_B8941_;
  assign new_B8933_ = B8914 | B8915;
  assign new_B8934_ = B8914 | new_B8921_;
  assign new_B8935_ = B8913 & new_B8925_;
  assign new_B8936_ = ~B8912 | ~B8913;
  assign new_B8937_ = new_B8921_ & new_B8936_;
  assign new_B8938_ = ~new_B8937_ & ~new_B8921_;
  assign new_B8939_ = new_B8921_ | new_B8936_;
  assign new_B8940_ = ~B8914 | ~B8915;
  assign new_B8941_ = new_B8921_ | new_B8936_;
  assign new_B8942_ = ~new_B8921_ & ~new_B8943_;
  assign new_B8943_ = new_B8921_ & new_B8936_;
  assign new_B8949_ = new_B8955_ & new_B8954_;
  assign new_B8950_ = new_B8957_ | new_B8956_;
  assign new_B8951_ = new_B8959_ | new_B8958_;
  assign new_B8952_ = new_B8954_ & new_B8960_;
  assign new_B8953_ = new_B8954_ & new_B8961_;
  assign new_B8954_ = B8944 ^ B8945;
  assign new_B8955_ = new_B8956_ ^ B8946;
  assign new_B8956_ = new_B8964_ & new_B8963_;
  assign new_B8957_ = new_B8962_ & B8946;
  assign new_B8958_ = new_B8967_ & new_B8966_;
  assign new_B8959_ = new_B8965_ & B8946;
  assign new_B8960_ = new_B8968_ | B8945;
  assign new_B8961_ = ~B8946 ^ new_B8958_;
  assign new_B8962_ = ~new_B8971_ | ~new_B8972_;
  assign new_B8963_ = B8947 ^ new_B8954_;
  assign new_B8964_ = new_B8973_ & new_B8966_;
  assign new_B8965_ = ~new_B8975_ | ~new_B8974_;
  assign new_B8966_ = B8947 | B8948;
  assign new_B8967_ = B8947 | new_B8954_;
  assign new_B8968_ = B8946 & new_B8958_;
  assign new_B8969_ = ~B8945 | ~B8946;
  assign new_B8970_ = new_B8954_ & new_B8969_;
  assign new_B8971_ = ~new_B8970_ & ~new_B8954_;
  assign new_B8972_ = new_B8954_ | new_B8969_;
  assign new_B8973_ = ~B8947 | ~B8948;
  assign new_B8974_ = new_B8954_ | new_B8969_;
  assign new_B8975_ = ~new_B8954_ & ~new_B8976_;
  assign new_B8976_ = new_B8954_ & new_B8969_;
  assign new_B8982_ = new_B8988_ & new_B8987_;
  assign new_B8983_ = new_B8990_ | new_B8989_;
  assign new_B8984_ = new_B8992_ | new_B8991_;
  assign new_B8985_ = new_B8987_ & new_B8993_;
  assign new_B8986_ = new_B8987_ & new_B8994_;
  assign new_B8987_ = B8977 ^ B8978;
  assign new_B8988_ = new_B8989_ ^ B8979;
  assign new_B8989_ = new_B8997_ & new_B8996_;
  assign new_B8990_ = new_B8995_ & B8979;
  assign new_B8991_ = new_B9000_ & new_B8999_;
  assign new_B8992_ = new_B8998_ & B8979;
  assign new_B8993_ = new_B9001_ | B8978;
  assign new_B8994_ = ~B8979 ^ new_B8991_;
  assign new_B8995_ = ~new_B9004_ | ~new_B9005_;
  assign new_B8996_ = B8980 ^ new_B8987_;
  assign new_B8997_ = new_B9006_ & new_B8999_;
  assign new_B8998_ = ~new_B9008_ | ~new_B9007_;
  assign new_B8999_ = B8980 | B8981;
  assign new_B9000_ = B8980 | new_B8987_;
  assign new_B9001_ = B8979 & new_B8991_;
  assign new_B9002_ = ~B8978 | ~B8979;
  assign new_B9003_ = new_B8987_ & new_B9002_;
  assign new_B9004_ = ~new_B9003_ & ~new_B8987_;
  assign new_B9005_ = new_B8987_ | new_B9002_;
  assign new_B9006_ = ~B8980 | ~B8981;
  assign new_B9007_ = new_B8987_ | new_B9002_;
  assign new_B9008_ = ~new_B8987_ & ~new_B9009_;
  assign new_B9009_ = new_B8987_ & new_B9002_;
  assign new_B9015_ = new_B9021_ & new_B9020_;
  assign new_B9016_ = new_B9023_ | new_B9022_;
  assign new_B9017_ = new_B9025_ | new_B9024_;
  assign new_B9018_ = new_B9020_ & new_B9026_;
  assign new_B9019_ = new_B9020_ & new_B9027_;
  assign new_B9020_ = B9010 ^ B9011;
  assign new_B9021_ = new_B9022_ ^ B9012;
  assign new_B9022_ = new_B9030_ & new_B9029_;
  assign new_B9023_ = new_B9028_ & B9012;
  assign new_B9024_ = new_B9033_ & new_B9032_;
  assign new_B9025_ = new_B9031_ & B9012;
  assign new_B9026_ = new_B9034_ | B9011;
  assign new_B9027_ = ~B9012 ^ new_B9024_;
  assign new_B9028_ = ~new_B9037_ | ~new_B9038_;
  assign new_B9029_ = B9013 ^ new_B9020_;
  assign new_B9030_ = new_B9039_ & new_B9032_;
  assign new_B9031_ = ~new_B9041_ | ~new_B9040_;
  assign new_B9032_ = B9013 | B9014;
  assign new_B9033_ = B9013 | new_B9020_;
  assign new_B9034_ = B9012 & new_B9024_;
  assign new_B9035_ = ~B9011 | ~B9012;
  assign new_B9036_ = new_B9020_ & new_B9035_;
  assign new_B9037_ = ~new_B9036_ & ~new_B9020_;
  assign new_B9038_ = new_B9020_ | new_B9035_;
  assign new_B9039_ = ~B9013 | ~B9014;
  assign new_B9040_ = new_B9020_ | new_B9035_;
  assign new_B9041_ = ~new_B9020_ & ~new_B9042_;
  assign new_B9042_ = new_B9020_ & new_B9035_;
  assign new_B9048_ = new_B9054_ & new_B9053_;
  assign new_B9049_ = new_B9056_ | new_B9055_;
  assign new_B9050_ = new_B9058_ | new_B9057_;
  assign new_B9051_ = new_B9053_ & new_B9059_;
  assign new_B9052_ = new_B9053_ & new_B9060_;
  assign new_B9053_ = B9043 ^ B9044;
  assign new_B9054_ = new_B9055_ ^ B9045;
  assign new_B9055_ = new_B9063_ & new_B9062_;
  assign new_B9056_ = new_B9061_ & B9045;
  assign new_B9057_ = new_B9066_ & new_B9065_;
  assign new_B9058_ = new_B9064_ & B9045;
  assign new_B9059_ = new_B9067_ | B9044;
  assign new_B9060_ = ~B9045 ^ new_B9057_;
  assign new_B9061_ = ~new_B9070_ | ~new_B9071_;
  assign new_B9062_ = B9046 ^ new_B9053_;
  assign new_B9063_ = new_B9072_ & new_B9065_;
  assign new_B9064_ = ~new_B9074_ | ~new_B9073_;
  assign new_B9065_ = B9046 | B9047;
  assign new_B9066_ = B9046 | new_B9053_;
  assign new_B9067_ = B9045 & new_B9057_;
  assign new_B9068_ = ~B9044 | ~B9045;
  assign new_B9069_ = new_B9053_ & new_B9068_;
  assign new_B9070_ = ~new_B9069_ & ~new_B9053_;
  assign new_B9071_ = new_B9053_ | new_B9068_;
  assign new_B9072_ = ~B9046 | ~B9047;
  assign new_B9073_ = new_B9053_ | new_B9068_;
  assign new_B9074_ = ~new_B9053_ & ~new_B9075_;
  assign new_B9075_ = new_B9053_ & new_B9068_;
  assign new_B9081_ = new_B9087_ & new_B9086_;
  assign new_B9082_ = new_B9089_ | new_B9088_;
  assign new_B9083_ = new_B9091_ | new_B9090_;
  assign new_B9084_ = new_B9086_ & new_B9092_;
  assign new_B9085_ = new_B9086_ & new_B9093_;
  assign new_B9086_ = B9076 ^ B9077;
  assign new_B9087_ = new_B9088_ ^ B9078;
  assign new_B9088_ = new_B9096_ & new_B9095_;
  assign new_B9089_ = new_B9094_ & B9078;
  assign new_B9090_ = new_B9099_ & new_B9098_;
  assign new_B9091_ = new_B9097_ & B9078;
  assign new_B9092_ = new_B9100_ | B9077;
  assign new_B9093_ = ~B9078 ^ new_B9090_;
  assign new_B9094_ = ~new_B9103_ | ~new_B9104_;
  assign new_B9095_ = B9079 ^ new_B9086_;
  assign new_B9096_ = new_B9105_ & new_B9098_;
  assign new_B9097_ = ~new_B9107_ | ~new_B9106_;
  assign new_B9098_ = B9079 | B9080;
  assign new_B9099_ = B9079 | new_B9086_;
  assign new_B9100_ = B9078 & new_B9090_;
  assign new_B9101_ = ~B9077 | ~B9078;
  assign new_B9102_ = new_B9086_ & new_B9101_;
  assign new_B9103_ = ~new_B9102_ & ~new_B9086_;
  assign new_B9104_ = new_B9086_ | new_B9101_;
  assign new_B9105_ = ~B9079 | ~B9080;
  assign new_B9106_ = new_B9086_ | new_B9101_;
  assign new_B9107_ = ~new_B9086_ & ~new_B9108_;
  assign new_B9108_ = new_B9086_ & new_B9101_;
  assign new_B9114_ = new_B9120_ & new_B9119_;
  assign new_B9115_ = new_B9122_ | new_B9121_;
  assign new_B9116_ = new_B9124_ | new_B9123_;
  assign new_B9117_ = new_B9119_ & new_B9125_;
  assign new_B9118_ = new_B9119_ & new_B9126_;
  assign new_B9119_ = B9109 ^ B9110;
  assign new_B9120_ = new_B9121_ ^ B9111;
  assign new_B9121_ = new_B9129_ & new_B9128_;
  assign new_B9122_ = new_B9127_ & B9111;
  assign new_B9123_ = new_B9132_ & new_B9131_;
  assign new_B9124_ = new_B9130_ & B9111;
  assign new_B9125_ = new_B9133_ | B9110;
  assign new_B9126_ = ~B9111 ^ new_B9123_;
  assign new_B9127_ = ~new_B9136_ | ~new_B9137_;
  assign new_B9128_ = B9112 ^ new_B9119_;
  assign new_B9129_ = new_B9138_ & new_B9131_;
  assign new_B9130_ = ~new_B9140_ | ~new_B9139_;
  assign new_B9131_ = B9112 | B9113;
  assign new_B9132_ = B9112 | new_B9119_;
  assign new_B9133_ = B9111 & new_B9123_;
  assign new_B9134_ = ~B9110 | ~B9111;
  assign new_B9135_ = new_B9119_ & new_B9134_;
  assign new_B9136_ = ~new_B9135_ & ~new_B9119_;
  assign new_B9137_ = new_B9119_ | new_B9134_;
  assign new_B9138_ = ~B9112 | ~B9113;
  assign new_B9139_ = new_B9119_ | new_B9134_;
  assign new_B9140_ = ~new_B9119_ & ~new_B9141_;
  assign new_B9141_ = new_B9119_ & new_B9134_;
  assign new_B9147_ = new_B9153_ & new_B9152_;
  assign new_B9148_ = new_B9155_ | new_B9154_;
  assign new_B9149_ = new_B9157_ | new_B9156_;
  assign new_B9150_ = new_B9152_ & new_B9158_;
  assign new_B9151_ = new_B9152_ & new_B9159_;
  assign new_B9152_ = B9142 ^ B9143;
  assign new_B9153_ = new_B9154_ ^ B9144;
  assign new_B9154_ = new_B9162_ & new_B9161_;
  assign new_B9155_ = new_B9160_ & B9144;
  assign new_B9156_ = new_B9165_ & new_B9164_;
  assign new_B9157_ = new_B9163_ & B9144;
  assign new_B9158_ = new_B9166_ | B9143;
  assign new_B9159_ = ~B9144 ^ new_B9156_;
  assign new_B9160_ = ~new_B9169_ | ~new_B9170_;
  assign new_B9161_ = B9145 ^ new_B9152_;
  assign new_B9162_ = new_B9171_ & new_B9164_;
  assign new_B9163_ = ~new_B9173_ | ~new_B9172_;
  assign new_B9164_ = B9145 | B9146;
  assign new_B9165_ = B9145 | new_B9152_;
  assign new_B9166_ = B9144 & new_B9156_;
  assign new_B9167_ = ~B9143 | ~B9144;
  assign new_B9168_ = new_B9152_ & new_B9167_;
  assign new_B9169_ = ~new_B9168_ & ~new_B9152_;
  assign new_B9170_ = new_B9152_ | new_B9167_;
  assign new_B9171_ = ~B9145 | ~B9146;
  assign new_B9172_ = new_B9152_ | new_B9167_;
  assign new_B9173_ = ~new_B9152_ & ~new_B9174_;
  assign new_B9174_ = new_B9152_ & new_B9167_;
  assign new_B9180_ = new_B9186_ & new_B9185_;
  assign new_B9181_ = new_B9188_ | new_B9187_;
  assign new_B9182_ = new_B9190_ | new_B9189_;
  assign new_B9183_ = new_B9185_ & new_B9191_;
  assign new_B9184_ = new_B9185_ & new_B9192_;
  assign new_B9185_ = B9175 ^ B9176;
  assign new_B9186_ = new_B9187_ ^ B9177;
  assign new_B9187_ = new_B9195_ & new_B9194_;
  assign new_B9188_ = new_B9193_ & B9177;
  assign new_B9189_ = new_B9198_ & new_B9197_;
  assign new_B9190_ = new_B9196_ & B9177;
  assign new_B9191_ = new_B9199_ | B9176;
  assign new_B9192_ = ~B9177 ^ new_B9189_;
  assign new_B9193_ = ~new_B9202_ | ~new_B9203_;
  assign new_B9194_ = B9178 ^ new_B9185_;
  assign new_B9195_ = new_B9204_ & new_B9197_;
  assign new_B9196_ = ~new_B9206_ | ~new_B9205_;
  assign new_B9197_ = B9178 | B9179;
  assign new_B9198_ = B9178 | new_B9185_;
  assign new_B9199_ = B9177 & new_B9189_;
  assign new_B9200_ = ~B9176 | ~B9177;
  assign new_B9201_ = new_B9185_ & new_B9200_;
  assign new_B9202_ = ~new_B9201_ & ~new_B9185_;
  assign new_B9203_ = new_B9185_ | new_B9200_;
  assign new_B9204_ = ~B9178 | ~B9179;
  assign new_B9205_ = new_B9185_ | new_B9200_;
  assign new_B9206_ = ~new_B9185_ & ~new_B9207_;
  assign new_B9207_ = new_B9185_ & new_B9200_;
  assign new_B9213_ = new_B9219_ & new_B9218_;
  assign new_B9214_ = new_B9221_ | new_B9220_;
  assign new_B9215_ = new_B9223_ | new_B9222_;
  assign new_B9216_ = new_B9218_ & new_B9224_;
  assign new_B9217_ = new_B9218_ & new_B9225_;
  assign new_B9218_ = B9208 ^ B9209;
  assign new_B9219_ = new_B9220_ ^ B9210;
  assign new_B9220_ = new_B9228_ & new_B9227_;
  assign new_B9221_ = new_B9226_ & B9210;
  assign new_B9222_ = new_B9231_ & new_B9230_;
  assign new_B9223_ = new_B9229_ & B9210;
  assign new_B9224_ = new_B9232_ | B9209;
  assign new_B9225_ = ~B9210 ^ new_B9222_;
  assign new_B9226_ = ~new_B9235_ | ~new_B9236_;
  assign new_B9227_ = B9211 ^ new_B9218_;
  assign new_B9228_ = new_B9237_ & new_B9230_;
  assign new_B9229_ = ~new_B9239_ | ~new_B9238_;
  assign new_B9230_ = B9211 | B9212;
  assign new_B9231_ = B9211 | new_B9218_;
  assign new_B9232_ = B9210 & new_B9222_;
  assign new_B9233_ = ~B9209 | ~B9210;
  assign new_B9234_ = new_B9218_ & new_B9233_;
  assign new_B9235_ = ~new_B9234_ & ~new_B9218_;
  assign new_B9236_ = new_B9218_ | new_B9233_;
  assign new_B9237_ = ~B9211 | ~B9212;
  assign new_B9238_ = new_B9218_ | new_B9233_;
  assign new_B9239_ = ~new_B9218_ & ~new_B9240_;
  assign new_B9240_ = new_B9218_ & new_B9233_;
  assign new_B9246_ = new_B9252_ & new_B9251_;
  assign new_B9247_ = new_B9254_ | new_B9253_;
  assign new_B9248_ = new_B9256_ | new_B9255_;
  assign new_B9249_ = new_B9251_ & new_B9257_;
  assign new_B9250_ = new_B9251_ & new_B9258_;
  assign new_B9251_ = B9241 ^ B9242;
  assign new_B9252_ = new_B9253_ ^ B9243;
  assign new_B9253_ = new_B9261_ & new_B9260_;
  assign new_B9254_ = new_B9259_ & B9243;
  assign new_B9255_ = new_B9264_ & new_B9263_;
  assign new_B9256_ = new_B9262_ & B9243;
  assign new_B9257_ = new_B9265_ | B9242;
  assign new_B9258_ = ~B9243 ^ new_B9255_;
  assign new_B9259_ = ~new_B9268_ | ~new_B9269_;
  assign new_B9260_ = B9244 ^ new_B9251_;
  assign new_B9261_ = new_B9270_ & new_B9263_;
  assign new_B9262_ = ~new_B9272_ | ~new_B9271_;
  assign new_B9263_ = B9244 | B9245;
  assign new_B9264_ = B9244 | new_B9251_;
  assign new_B9265_ = B9243 & new_B9255_;
  assign new_B9266_ = ~B9242 | ~B9243;
  assign new_B9267_ = new_B9251_ & new_B9266_;
  assign new_B9268_ = ~new_B9267_ & ~new_B9251_;
  assign new_B9269_ = new_B9251_ | new_B9266_;
  assign new_B9270_ = ~B9244 | ~B9245;
  assign new_B9271_ = new_B9251_ | new_B9266_;
  assign new_B9272_ = ~new_B9251_ & ~new_B9273_;
  assign new_B9273_ = new_B9251_ & new_B9266_;
  assign new_B9279_ = new_B9285_ & new_B9284_;
  assign new_B9280_ = new_B9287_ | new_B9286_;
  assign new_B9281_ = new_B9289_ | new_B9288_;
  assign new_B9282_ = new_B9284_ & new_B9290_;
  assign new_B9283_ = new_B9284_ & new_B9291_;
  assign new_B9284_ = B9274 ^ B9275;
  assign new_B9285_ = new_B9286_ ^ B9276;
  assign new_B9286_ = new_B9294_ & new_B9293_;
  assign new_B9287_ = new_B9292_ & B9276;
  assign new_B9288_ = new_B9297_ & new_B9296_;
  assign new_B9289_ = new_B9295_ & B9276;
  assign new_B9290_ = new_B9298_ | B9275;
  assign new_B9291_ = ~B9276 ^ new_B9288_;
  assign new_B9292_ = ~new_B9301_ | ~new_B9302_;
  assign new_B9293_ = B9277 ^ new_B9284_;
  assign new_B9294_ = new_B9303_ & new_B9296_;
  assign new_B9295_ = ~new_B9305_ | ~new_B9304_;
  assign new_B9296_ = B9277 | B9278;
  assign new_B9297_ = B9277 | new_B9284_;
  assign new_B9298_ = B9276 & new_B9288_;
  assign new_B9299_ = ~B9275 | ~B9276;
  assign new_B9300_ = new_B9284_ & new_B9299_;
  assign new_B9301_ = ~new_B9300_ & ~new_B9284_;
  assign new_B9302_ = new_B9284_ | new_B9299_;
  assign new_B9303_ = ~B9277 | ~B9278;
  assign new_B9304_ = new_B9284_ | new_B9299_;
  assign new_B9305_ = ~new_B9284_ & ~new_B9306_;
  assign new_B9306_ = new_B9284_ & new_B9299_;
  assign new_B1089_ = new_B1067_ & new_B1082_;
  assign new_B1088_ = ~new_B1067_ & ~new_B1089_;
  assign new_B1087_ = new_B1067_ | new_B1082_;
  assign new_B1086_ = ~new_B1060_ | ~new_B1061_;
  assign new_B1085_ = new_B1067_ | new_B1082_;
  assign new_B1084_ = ~new_B1083_ & ~new_B1067_;
  assign new_B1083_ = new_B1067_ & new_B1082_;
  assign new_B1082_ = ~new_B1058_ | ~new_B1059_;
  assign new_B1081_ = new_B1059_ & new_B1071_;
  assign new_B1080_ = new_B1060_ | new_B1067_;
  assign new_B1079_ = new_B1060_ | new_B1061_;
  assign new_B1078_ = ~new_B1088_ | ~new_B1087_;
  assign new_B1077_ = new_B1086_ & new_B1079_;
  assign new_B1076_ = new_B1060_ ^ new_B1067_;
  assign new_B1075_ = ~new_B1084_ | ~new_B1085_;
  assign new_B1074_ = ~new_B1059_ ^ new_B1071_;
  assign new_B1073_ = new_B1081_ | new_B1058_;
  assign new_B1072_ = new_B1078_ & new_B1059_;
  assign new_B1071_ = new_B1080_ & new_B1079_;
  assign new_B1070_ = new_B1075_ & new_B1059_;
  assign new_B1069_ = new_B1077_ & new_B1076_;
  assign new_B1068_ = new_B1069_ ^ new_B1059_;
  assign new_B1067_ = new_B1057_ ^ new_B1058_;
  assign new_B1066_ = new_B1067_ & new_B1074_;
  assign new_B1065_ = new_B1067_ & new_B1073_;
  assign new_B1064_ = new_B1072_ | new_B1071_;
  assign new_B1063_ = new_B1070_ | new_B1069_;
  assign new_B1062_ = new_B1068_ & new_B1067_;
  assign new_B1061_ = new_B5191_;
  assign new_B1060_ = new_B5220_;
  assign new_B1059_ = new_B5253_;
  assign new_B1058_ = new_B5286_;
  assign new_B1057_ = new_B5319_;
  assign new_B1090_ = new_B5352_;
  assign new_B1091_ = new_B5385_;
  assign new_B1092_ = new_B5418_;
  assign new_B1093_ = new_B5451_;
  assign new_B1094_ = new_B5484_;
  assign new_B1095_ = new_B1101_ & new_B1100_;
  assign new_B1096_ = new_B1103_ | new_B1102_;
  assign new_B1097_ = new_B1105_ | new_B1104_;
  assign new_B1098_ = new_B1100_ & new_B1106_;
  assign new_B1099_ = new_B1100_ & new_B1107_;
  assign new_B1100_ = new_B1090_ ^ new_B1091_;
  assign new_B1101_ = new_B1102_ ^ new_B1092_;
  assign new_B1102_ = new_B1110_ & new_B1109_;
  assign new_B1103_ = new_B1108_ & new_B1092_;
  assign new_B1104_ = new_B1113_ & new_B1112_;
  assign new_B1105_ = new_B1111_ & new_B1092_;
  assign new_B1106_ = new_B1114_ | new_B1091_;
  assign new_B1107_ = ~new_B1092_ ^ new_B1104_;
  assign new_B1108_ = ~new_B1117_ | ~new_B1118_;
  assign new_B1109_ = new_B1093_ ^ new_B1100_;
  assign new_B1110_ = new_B1119_ & new_B1112_;
  assign new_B1111_ = ~new_B1121_ | ~new_B1120_;
  assign new_B1112_ = new_B1093_ | new_B1094_;
  assign new_B1113_ = new_B1093_ | new_B1100_;
  assign new_B1114_ = new_B1092_ & new_B1104_;
  assign new_B1115_ = ~new_B1091_ | ~new_B1092_;
  assign new_B1116_ = new_B1100_ & new_B1115_;
  assign new_B1117_ = ~new_B1116_ & ~new_B1100_;
  assign new_B1118_ = new_B1100_ | new_B1115_;
  assign new_B1119_ = ~new_B1093_ | ~new_B1094_;
  assign new_B1120_ = new_B1100_ | new_B1115_;
  assign new_B1121_ = ~new_B1100_ & ~new_B1122_;
  assign new_B1122_ = new_B1100_ & new_B1115_;
  assign new_B1123_ = new_B5517_;
  assign new_B1124_ = new_B5550_;
  assign new_B1125_ = new_B5583_;
  assign new_B1126_ = new_B5616_;
  assign new_B1127_ = new_B5649_;
  assign new_B1128_ = new_B1134_ & new_B1133_;
  assign new_B1129_ = new_B1136_ | new_B1135_;
  assign new_B1130_ = new_B1138_ | new_B1137_;
  assign new_B1131_ = new_B1133_ & new_B1139_;
  assign new_B1132_ = new_B1133_ & new_B1140_;
  assign new_B1133_ = new_B1123_ ^ new_B1124_;
  assign new_B1134_ = new_B1135_ ^ new_B1125_;
  assign new_B1135_ = new_B1143_ & new_B1142_;
  assign new_B1136_ = new_B1141_ & new_B1125_;
  assign new_B1137_ = new_B1146_ & new_B1145_;
  assign new_B1138_ = new_B1144_ & new_B1125_;
  assign new_B1139_ = new_B1147_ | new_B1124_;
  assign new_B1140_ = ~new_B1125_ ^ new_B1137_;
  assign new_B1141_ = ~new_B1150_ | ~new_B1151_;
  assign new_B1142_ = new_B1126_ ^ new_B1133_;
  assign new_B1143_ = new_B1152_ & new_B1145_;
  assign new_B1144_ = ~new_B1154_ | ~new_B1153_;
  assign new_B1145_ = new_B1126_ | new_B1127_;
  assign new_B1146_ = new_B1126_ | new_B1133_;
  assign new_B1147_ = new_B1125_ & new_B1137_;
  assign new_B1148_ = ~new_B1124_ | ~new_B1125_;
  assign new_B1149_ = new_B1133_ & new_B1148_;
  assign new_B1150_ = ~new_B1149_ & ~new_B1133_;
  assign new_B1151_ = new_B1133_ | new_B1148_;
  assign new_B1152_ = ~new_B1126_ | ~new_B1127_;
  assign new_B1153_ = new_B1133_ | new_B1148_;
  assign new_B1154_ = ~new_B1133_ & ~new_B1155_;
  assign new_B1155_ = new_B1133_ & new_B1148_;
  assign new_B1156_ = new_B5682_;
  assign new_B1157_ = new_B5715_;
  assign new_B1158_ = new_B5748_;
  assign new_B1159_ = new_B5781_;
  assign new_B1160_ = new_B5814_;
  assign new_B1161_ = new_B1167_ & new_B1166_;
  assign new_B1162_ = new_B1169_ | new_B1168_;
  assign new_B1163_ = new_B1171_ | new_B1170_;
  assign new_B1164_ = new_B1166_ & new_B1172_;
  assign new_B1165_ = new_B1166_ & new_B1173_;
  assign new_B1166_ = new_B1156_ ^ new_B1157_;
  assign new_B1167_ = new_B1168_ ^ new_B1158_;
  assign new_B1168_ = new_B1176_ & new_B1175_;
  assign new_B1169_ = new_B1174_ & new_B1158_;
  assign new_B1170_ = new_B1179_ & new_B1178_;
  assign new_B1171_ = new_B1177_ & new_B1158_;
  assign new_B1172_ = new_B1180_ | new_B1157_;
  assign new_B1173_ = ~new_B1158_ ^ new_B1170_;
  assign new_B1174_ = ~new_B1183_ | ~new_B1184_;
  assign new_B1175_ = new_B1159_ ^ new_B1166_;
  assign new_B1176_ = new_B1185_ & new_B1178_;
  assign new_B1177_ = ~new_B1187_ | ~new_B1186_;
  assign new_B1178_ = new_B1159_ | new_B1160_;
  assign new_B1179_ = new_B1159_ | new_B1166_;
  assign new_B1180_ = new_B1158_ & new_B1170_;
  assign new_B1181_ = ~new_B1157_ | ~new_B1158_;
  assign new_B1182_ = new_B1166_ & new_B1181_;
  assign new_B1183_ = ~new_B1182_ & ~new_B1166_;
  assign new_B1184_ = new_B1166_ | new_B1181_;
  assign new_B1185_ = ~new_B1159_ | ~new_B1160_;
  assign new_B1186_ = new_B1166_ | new_B1181_;
  assign new_B1187_ = ~new_B1166_ & ~new_B1188_;
  assign new_B1188_ = new_B1166_ & new_B1181_;
  assign new_B1189_ = new_B5847_;
  assign new_B1190_ = new_B5880_;
  assign new_B1191_ = new_B5913_;
  assign new_B1192_ = new_B5946_;
  assign new_B1193_ = new_B5979_;
  assign new_B1194_ = new_B1200_ & new_B1199_;
  assign new_B1195_ = new_B1202_ | new_B1201_;
  assign new_B1196_ = new_B1204_ | new_B1203_;
  assign new_B1197_ = new_B1199_ & new_B1205_;
  assign new_B1198_ = new_B1199_ & new_B1206_;
  assign new_B1199_ = new_B1189_ ^ new_B1190_;
  assign new_B1200_ = new_B1201_ ^ new_B1191_;
  assign new_B1201_ = new_B1209_ & new_B1208_;
  assign new_B1202_ = new_B1207_ & new_B1191_;
  assign new_B1203_ = new_B1212_ & new_B1211_;
  assign new_B1204_ = new_B1210_ & new_B1191_;
  assign new_B1205_ = new_B1213_ | new_B1190_;
  assign new_B1206_ = ~new_B1191_ ^ new_B1203_;
  assign new_B1207_ = ~new_B1216_ | ~new_B1217_;
  assign new_B1208_ = new_B1192_ ^ new_B1199_;
  assign new_B1209_ = new_B1218_ & new_B1211_;
  assign new_B1210_ = ~new_B1220_ | ~new_B1219_;
  assign new_B1211_ = new_B1192_ | new_B1193_;
  assign new_B1212_ = new_B1192_ | new_B1199_;
  assign new_B1213_ = new_B1191_ & new_B1203_;
  assign new_B1214_ = ~new_B1190_ | ~new_B1191_;
  assign new_B1215_ = new_B1199_ & new_B1214_;
  assign new_B1216_ = ~new_B1215_ & ~new_B1199_;
  assign new_B1217_ = new_B1199_ | new_B1214_;
  assign new_B1218_ = ~new_B1192_ | ~new_B1193_;
  assign new_B1219_ = new_B1199_ | new_B1214_;
  assign new_B1220_ = ~new_B1199_ & ~new_B1221_;
  assign new_B1221_ = new_B1199_ & new_B1214_;
  assign new_B1222_ = new_B6012_;
  assign new_B1223_ = new_B6045_;
  assign new_B1224_ = new_B6078_;
  assign new_B1225_ = new_B6111_;
  assign new_B1226_ = new_B6144_;
  assign new_B1227_ = new_B1233_ & new_B1232_;
  assign new_B1228_ = new_B1235_ | new_B1234_;
  assign new_B1229_ = new_B1237_ | new_B1236_;
  assign new_B1230_ = new_B1232_ & new_B1238_;
  assign new_B1231_ = new_B1232_ & new_B1239_;
  assign new_B1232_ = new_B1222_ ^ new_B1223_;
  assign new_B1233_ = new_B1234_ ^ new_B1224_;
  assign new_B1234_ = new_B1242_ & new_B1241_;
  assign new_B1235_ = new_B1240_ & new_B1224_;
  assign new_B1236_ = new_B1245_ & new_B1244_;
  assign new_B1237_ = new_B1243_ & new_B1224_;
  assign new_B1238_ = new_B1246_ | new_B1223_;
  assign new_B1239_ = ~new_B1224_ ^ new_B1236_;
  assign new_B1240_ = ~new_B1249_ | ~new_B1250_;
  assign new_B1241_ = new_B1225_ ^ new_B1232_;
  assign new_B1242_ = new_B1251_ & new_B1244_;
  assign new_B1243_ = ~new_B1253_ | ~new_B1252_;
  assign new_B1244_ = new_B1225_ | new_B1226_;
  assign new_B1245_ = new_B1225_ | new_B1232_;
  assign new_B1246_ = new_B1224_ & new_B1236_;
  assign new_B1247_ = ~new_B1223_ | ~new_B1224_;
  assign new_B1248_ = new_B1232_ & new_B1247_;
  assign new_B1249_ = ~new_B1248_ & ~new_B1232_;
  assign new_B1250_ = new_B1232_ | new_B1247_;
  assign new_B1251_ = ~new_B1225_ | ~new_B1226_;
  assign new_B1252_ = new_B1232_ | new_B1247_;
  assign new_B1253_ = ~new_B1232_ & ~new_B1254_;
  assign new_B1254_ = new_B1232_ & new_B1247_;
  assign new_B1255_ = new_B6177_;
  assign new_B1256_ = new_B6210_;
  assign new_B1257_ = new_B6243_;
  assign new_B1258_ = new_B6276_;
  assign new_B1259_ = new_B6309_;
  assign new_B1260_ = new_B1266_ & new_B1265_;
  assign new_B1261_ = new_B1268_ | new_B1267_;
  assign new_B1262_ = new_B1270_ | new_B1269_;
  assign new_B1263_ = new_B1265_ & new_B1271_;
  assign new_B1264_ = new_B1265_ & new_B1272_;
  assign new_B1265_ = new_B1255_ ^ new_B1256_;
  assign new_B1266_ = new_B1267_ ^ new_B1257_;
  assign new_B1267_ = new_B1275_ & new_B1274_;
  assign new_B1268_ = new_B1273_ & new_B1257_;
  assign new_B1269_ = new_B1278_ & new_B1277_;
  assign new_B1270_ = new_B1276_ & new_B1257_;
  assign new_B1271_ = new_B1279_ | new_B1256_;
  assign new_B1272_ = ~new_B1257_ ^ new_B1269_;
  assign new_B1273_ = ~new_B1282_ | ~new_B1283_;
  assign new_B1274_ = new_B1258_ ^ new_B1265_;
  assign new_B1275_ = new_B1284_ & new_B1277_;
  assign new_B1276_ = ~new_B1286_ | ~new_B1285_;
  assign new_B1277_ = new_B1258_ | new_B1259_;
  assign new_B1278_ = new_B1258_ | new_B1265_;
  assign new_B1279_ = new_B1257_ & new_B1269_;
  assign new_B1280_ = ~new_B1256_ | ~new_B1257_;
  assign new_B1281_ = new_B1265_ & new_B1280_;
  assign new_B1282_ = ~new_B1281_ & ~new_B1265_;
  assign new_B1283_ = new_B1265_ | new_B1280_;
  assign new_B1284_ = ~new_B1258_ | ~new_B1259_;
  assign new_B1285_ = new_B1265_ | new_B1280_;
  assign new_B1286_ = ~new_B1265_ & ~new_B1287_;
  assign new_B1287_ = new_B1265_ & new_B1280_;
  assign new_B1288_ = new_B6342_;
  assign new_B1289_ = new_B6375_;
  assign new_B1290_ = new_B6408_;
  assign new_B1291_ = new_B6441_;
  assign new_B1292_ = new_B6474_;
  assign new_B1293_ = new_B1299_ & new_B1298_;
  assign new_B1294_ = new_B1301_ | new_B1300_;
  assign new_B1295_ = new_B1303_ | new_B1302_;
  assign new_B1296_ = new_B1298_ & new_B1304_;
  assign new_B1297_ = new_B1298_ & new_B1305_;
  assign new_B1298_ = new_B1288_ ^ new_B1289_;
  assign new_B1299_ = new_B1300_ ^ new_B1290_;
  assign new_B1300_ = new_B1308_ & new_B1307_;
  assign new_B1301_ = new_B1306_ & new_B1290_;
  assign new_B1302_ = new_B1311_ & new_B1310_;
  assign new_B1303_ = new_B1309_ & new_B1290_;
  assign new_B1304_ = new_B1312_ | new_B1289_;
  assign new_B1305_ = ~new_B1290_ ^ new_B1302_;
  assign new_B1306_ = ~new_B1315_ | ~new_B1316_;
  assign new_B1307_ = new_B1291_ ^ new_B1298_;
  assign new_B1308_ = new_B1317_ & new_B1310_;
  assign new_B1309_ = ~new_B1319_ | ~new_B1318_;
  assign new_B1310_ = new_B1291_ | new_B1292_;
  assign new_B1311_ = new_B1291_ | new_B1298_;
  assign new_B1312_ = new_B1290_ & new_B1302_;
  assign new_B1313_ = ~new_B1289_ | ~new_B1290_;
  assign new_B1314_ = new_B1298_ & new_B1313_;
  assign new_B1315_ = ~new_B1314_ & ~new_B1298_;
  assign new_B1316_ = new_B1298_ | new_B1313_;
  assign new_B1317_ = ~new_B1291_ | ~new_B1292_;
  assign new_B1318_ = new_B1298_ | new_B1313_;
  assign new_B1319_ = ~new_B1298_ & ~new_B1320_;
  assign new_B1320_ = new_B1298_ & new_B1313_;
  assign new_B1321_ = new_B6507_;
  assign new_B1322_ = new_B6540_;
  assign new_B1323_ = new_B6573_;
  assign new_B1324_ = new_B6606_;
  assign new_B1325_ = new_B6639_;
  assign new_B1326_ = new_B1332_ & new_B1331_;
  assign new_B1327_ = new_B1334_ | new_B1333_;
  assign new_B1328_ = new_B1336_ | new_B1335_;
  assign new_B1329_ = new_B1331_ & new_B1337_;
  assign new_B1330_ = new_B1331_ & new_B1338_;
  assign new_B1331_ = new_B1321_ ^ new_B1322_;
  assign new_B1332_ = new_B1333_ ^ new_B1323_;
  assign new_B1333_ = new_B1341_ & new_B1340_;
  assign new_B1334_ = new_B1339_ & new_B1323_;
  assign new_B1335_ = new_B1344_ & new_B1343_;
  assign new_B1336_ = new_B1342_ & new_B1323_;
  assign new_B1337_ = new_B1345_ | new_B1322_;
  assign new_B1338_ = ~new_B1323_ ^ new_B1335_;
  assign new_B1339_ = ~new_B1348_ | ~new_B1349_;
  assign new_B1340_ = new_B1324_ ^ new_B1331_;
  assign new_B1341_ = new_B1350_ & new_B1343_;
  assign new_B1342_ = ~new_B1352_ | ~new_B1351_;
  assign new_B1343_ = new_B1324_ | new_B1325_;
  assign new_B1344_ = new_B1324_ | new_B1331_;
  assign new_B1345_ = new_B1323_ & new_B1335_;
  assign new_B1346_ = ~new_B1322_ | ~new_B1323_;
  assign new_B1347_ = new_B1331_ & new_B1346_;
  assign new_B1348_ = ~new_B1347_ & ~new_B1331_;
  assign new_B1349_ = new_B1331_ | new_B1346_;
  assign new_B1350_ = ~new_B1324_ | ~new_B1325_;
  assign new_B1351_ = new_B1331_ | new_B1346_;
  assign new_B1352_ = ~new_B1331_ & ~new_B1353_;
  assign new_B1353_ = new_B1331_ & new_B1346_;
  assign new_B1354_ = new_B6672_;
  assign new_B1355_ = new_B6705_;
  assign new_B1356_ = new_B6738_;
  assign new_B1357_ = new_B6771_;
  assign new_B1358_ = new_B6804_;
  assign new_B1359_ = new_B1365_ & new_B1364_;
  assign new_B1360_ = new_B1367_ | new_B1366_;
  assign new_B1361_ = new_B1369_ | new_B1368_;
  assign new_B1362_ = new_B1364_ & new_B1370_;
  assign new_B1363_ = new_B1364_ & new_B1371_;
  assign new_B1364_ = new_B1354_ ^ new_B1355_;
  assign new_B1365_ = new_B1366_ ^ new_B1356_;
  assign new_B1366_ = new_B1374_ & new_B1373_;
  assign new_B1367_ = new_B1372_ & new_B1356_;
  assign new_B1368_ = new_B1377_ & new_B1376_;
  assign new_B1369_ = new_B1375_ & new_B1356_;
  assign new_B1370_ = new_B1378_ | new_B1355_;
  assign new_B1371_ = ~new_B1356_ ^ new_B1368_;
  assign new_B1372_ = ~new_B1381_ | ~new_B1382_;
  assign new_B1373_ = new_B1357_ ^ new_B1364_;
  assign new_B1374_ = new_B1383_ & new_B1376_;
  assign new_B1375_ = ~new_B1385_ | ~new_B1384_;
  assign new_B1376_ = new_B1357_ | new_B1358_;
  assign new_B1377_ = new_B1357_ | new_B1364_;
  assign new_B1378_ = new_B1356_ & new_B1368_;
  assign new_B1379_ = ~new_B1355_ | ~new_B1356_;
  assign new_B1380_ = new_B1364_ & new_B1379_;
  assign new_B1381_ = ~new_B1380_ & ~new_B1364_;
  assign new_B1382_ = new_B1364_ | new_B1379_;
  assign new_B1383_ = ~new_B1357_ | ~new_B1358_;
  assign new_B1384_ = new_B1364_ | new_B1379_;
  assign new_B1385_ = ~new_B1364_ & ~new_B1386_;
  assign new_B1386_ = new_B1364_ & new_B1379_;
  assign new_B1387_ = new_B6837_;
  assign new_B1388_ = new_B6870_;
  assign new_B1389_ = new_B6903_;
  assign new_B1390_ = new_B6936_;
  assign new_B1391_ = new_B6969_;
  assign new_B1392_ = new_B1398_ & new_B1397_;
  assign new_B1393_ = new_B1400_ | new_B1399_;
  assign new_B1394_ = new_B1402_ | new_B1401_;
  assign new_B1395_ = new_B1397_ & new_B1403_;
  assign new_B1396_ = new_B1397_ & new_B1404_;
  assign new_B1397_ = new_B1387_ ^ new_B1388_;
  assign new_B1398_ = new_B1399_ ^ new_B1389_;
  assign new_B1399_ = new_B1407_ & new_B1406_;
  assign new_B1400_ = new_B1405_ & new_B1389_;
  assign new_B1401_ = new_B1410_ & new_B1409_;
  assign new_B1402_ = new_B1408_ & new_B1389_;
  assign new_B1403_ = new_B1411_ | new_B1388_;
  assign new_B1404_ = ~new_B1389_ ^ new_B1401_;
  assign new_B1405_ = ~new_B1414_ | ~new_B1415_;
  assign new_B1406_ = new_B1390_ ^ new_B1397_;
  assign new_B1407_ = new_B1416_ & new_B1409_;
  assign new_B1408_ = ~new_B1418_ | ~new_B1417_;
  assign new_B1409_ = new_B1390_ | new_B1391_;
  assign new_B1410_ = new_B1390_ | new_B1397_;
  assign new_B1411_ = new_B1389_ & new_B1401_;
  assign new_B1412_ = ~new_B1388_ | ~new_B1389_;
  assign new_B1413_ = new_B1397_ & new_B1412_;
  assign new_B1414_ = ~new_B1413_ & ~new_B1397_;
  assign new_B1415_ = new_B1397_ | new_B1412_;
  assign new_B1416_ = ~new_B1390_ | ~new_B1391_;
  assign new_B1417_ = new_B1397_ | new_B1412_;
  assign new_B1418_ = ~new_B1397_ & ~new_B1419_;
  assign new_B1419_ = new_B1397_ & new_B1412_;
  assign new_B1420_ = new_B7002_;
  assign new_B1421_ = new_B7035_;
  assign new_B1422_ = new_B7068_;
  assign new_B1423_ = new_B7101_;
  assign new_B1424_ = new_B7134_;
  assign new_B1425_ = new_B1431_ & new_B1430_;
  assign new_B1426_ = new_B1433_ | new_B1432_;
  assign new_B1427_ = new_B1435_ | new_B1434_;
  assign new_B1428_ = new_B1430_ & new_B1436_;
  assign new_B1429_ = new_B1430_ & new_B1437_;
  assign new_B1430_ = new_B1420_ ^ new_B1421_;
  assign new_B1431_ = new_B1432_ ^ new_B1422_;
  assign new_B1432_ = new_B1440_ & new_B1439_;
  assign new_B1433_ = new_B1438_ & new_B1422_;
  assign new_B1434_ = new_B1443_ & new_B1442_;
  assign new_B1435_ = new_B1441_ & new_B1422_;
  assign new_B1436_ = new_B1444_ | new_B1421_;
  assign new_B1437_ = ~new_B1422_ ^ new_B1434_;
  assign new_B1438_ = ~new_B1447_ | ~new_B1448_;
  assign new_B1439_ = new_B1423_ ^ new_B1430_;
  assign new_B1440_ = new_B1449_ & new_B1442_;
  assign new_B1441_ = ~new_B1451_ | ~new_B1450_;
  assign new_B1442_ = new_B1423_ | new_B1424_;
  assign new_B1443_ = new_B1423_ | new_B1430_;
  assign new_B1444_ = new_B1422_ & new_B1434_;
  assign new_B1445_ = ~new_B1421_ | ~new_B1422_;
  assign new_B1446_ = new_B1430_ & new_B1445_;
  assign new_B1447_ = ~new_B1446_ & ~new_B1430_;
  assign new_B1448_ = new_B1430_ | new_B1445_;
  assign new_B1449_ = ~new_B1423_ | ~new_B1424_;
  assign new_B1450_ = new_B1430_ | new_B1445_;
  assign new_B1451_ = ~new_B1430_ & ~new_B1452_;
  assign new_B1452_ = new_B1430_ & new_B1445_;
  assign new_B1453_ = new_B7167_;
  assign new_B1454_ = new_B7200_;
  assign new_B1455_ = new_B7233_;
  assign new_B1456_ = new_B7266_;
  assign new_B1457_ = new_B7299_;
  assign new_B1458_ = new_B1464_ & new_B1463_;
  assign new_B1459_ = new_B1466_ | new_B1465_;
  assign new_B1460_ = new_B1468_ | new_B1467_;
  assign new_B1461_ = new_B1463_ & new_B1469_;
  assign new_B1462_ = new_B1463_ & new_B1470_;
  assign new_B1463_ = new_B1453_ ^ new_B1454_;
  assign new_B1464_ = new_B1465_ ^ new_B1455_;
  assign new_B1465_ = new_B1473_ & new_B1472_;
  assign new_B1466_ = new_B1471_ & new_B1455_;
  assign new_B1467_ = new_B1476_ & new_B1475_;
  assign new_B1468_ = new_B1474_ & new_B1455_;
  assign new_B1469_ = new_B1477_ | new_B1454_;
  assign new_B1470_ = ~new_B1455_ ^ new_B1467_;
  assign new_B1471_ = ~new_B1480_ | ~new_B1481_;
  assign new_B1472_ = new_B1456_ ^ new_B1463_;
  assign new_B1473_ = new_B1482_ & new_B1475_;
  assign new_B1474_ = ~new_B1484_ | ~new_B1483_;
  assign new_B1475_ = new_B1456_ | new_B1457_;
  assign new_B1476_ = new_B1456_ | new_B1463_;
  assign new_B1477_ = new_B1455_ & new_B1467_;
  assign new_B1478_ = ~new_B1454_ | ~new_B1455_;
  assign new_B1479_ = new_B1463_ & new_B1478_;
  assign new_B1480_ = ~new_B1479_ & ~new_B1463_;
  assign new_B1481_ = new_B1463_ | new_B1478_;
  assign new_B1482_ = ~new_B1456_ | ~new_B1457_;
  assign new_B1483_ = new_B1463_ | new_B1478_;
  assign new_B1484_ = ~new_B1463_ & ~new_B1485_;
  assign new_B1485_ = new_B1463_ & new_B1478_;
  assign new_B1486_ = new_B7332_;
  assign new_B1487_ = new_B7365_;
  assign new_B1488_ = new_B7398_;
  assign new_B1489_ = new_B7431_;
  assign new_B1490_ = new_B7464_;
  assign new_B1491_ = new_B1497_ & new_B1496_;
  assign new_B1492_ = new_B1499_ | new_B1498_;
  assign new_B1493_ = new_B1501_ | new_B1500_;
  assign new_B1494_ = new_B1496_ & new_B1502_;
  assign new_B1495_ = new_B1496_ & new_B1503_;
  assign new_B1496_ = new_B1486_ ^ new_B1487_;
  assign new_B1497_ = new_B1498_ ^ new_B1488_;
  assign new_B1498_ = new_B1506_ & new_B1505_;
  assign new_B1499_ = new_B1504_ & new_B1488_;
  assign new_B1500_ = new_B1509_ & new_B1508_;
  assign new_B1501_ = new_B1507_ & new_B1488_;
  assign new_B1502_ = new_B1510_ | new_B1487_;
  assign new_B1503_ = ~new_B1488_ ^ new_B1500_;
  assign new_B1504_ = ~new_B1513_ | ~new_B1514_;
  assign new_B1505_ = new_B1489_ ^ new_B1496_;
  assign new_B1506_ = new_B1515_ & new_B1508_;
  assign new_B1507_ = ~new_B1517_ | ~new_B1516_;
  assign new_B1508_ = new_B1489_ | new_B1490_;
  assign new_B1509_ = new_B1489_ | new_B1496_;
  assign new_B1510_ = new_B1488_ & new_B1500_;
  assign new_B1511_ = ~new_B1487_ | ~new_B1488_;
  assign new_B1512_ = new_B1496_ & new_B1511_;
  assign new_B1513_ = ~new_B1512_ & ~new_B1496_;
  assign new_B1514_ = new_B1496_ | new_B1511_;
  assign new_B1515_ = ~new_B1489_ | ~new_B1490_;
  assign new_B1516_ = new_B1496_ | new_B1511_;
  assign new_B1517_ = ~new_B1496_ & ~new_B1518_;
  assign new_B1518_ = new_B1496_ & new_B1511_;
  assign new_B1519_ = new_B7497_;
  assign new_B1520_ = new_B7530_;
  assign new_B1521_ = new_B7563_;
  assign new_B1522_ = new_B7596_;
  assign new_B1523_ = new_B7629_;
  assign new_B1524_ = new_B1530_ & new_B1529_;
  assign new_B1525_ = new_B1532_ | new_B1531_;
  assign new_B1526_ = new_B1534_ | new_B1533_;
  assign new_B1527_ = new_B1529_ & new_B1535_;
  assign new_B1528_ = new_B1529_ & new_B1536_;
  assign new_B1529_ = new_B1519_ ^ new_B1520_;
  assign new_B1530_ = new_B1531_ ^ new_B1521_;
  assign new_B1531_ = new_B1539_ & new_B1538_;
  assign new_B1532_ = new_B1537_ & new_B1521_;
  assign new_B1533_ = new_B1542_ & new_B1541_;
  assign new_B1534_ = new_B1540_ & new_B1521_;
  assign new_B1535_ = new_B1543_ | new_B1520_;
  assign new_B1536_ = ~new_B1521_ ^ new_B1533_;
  assign new_B1537_ = ~new_B1546_ | ~new_B1547_;
  assign new_B1538_ = new_B1522_ ^ new_B1529_;
  assign new_B1539_ = new_B1548_ & new_B1541_;
  assign new_B1540_ = ~new_B1550_ | ~new_B1549_;
  assign new_B1541_ = new_B1522_ | new_B1523_;
  assign new_B1542_ = new_B1522_ | new_B1529_;
  assign new_B1543_ = new_B1521_ & new_B1533_;
  assign new_B1544_ = ~new_B1520_ | ~new_B1521_;
  assign new_B1545_ = new_B1529_ & new_B1544_;
  assign new_B1546_ = ~new_B1545_ & ~new_B1529_;
  assign new_B1547_ = new_B1529_ | new_B1544_;
  assign new_B1548_ = ~new_B1522_ | ~new_B1523_;
  assign new_B1549_ = new_B1529_ | new_B1544_;
  assign new_B1550_ = ~new_B1529_ & ~new_B1551_;
  assign new_B1551_ = new_B1529_ & new_B1544_;
  assign new_B1552_ = new_B7662_;
  assign new_B1553_ = new_B7695_;
  assign new_B1554_ = new_B7728_;
  assign new_B1555_ = new_B7761_;
  assign new_B1556_ = new_B7794_;
  assign new_B1557_ = new_B1563_ & new_B1562_;
  assign new_B1558_ = new_B1565_ | new_B1564_;
  assign new_B1559_ = new_B1567_ | new_B1566_;
  assign new_B1560_ = new_B1562_ & new_B1568_;
  assign new_B1561_ = new_B1562_ & new_B1569_;
  assign new_B1562_ = new_B1552_ ^ new_B1553_;
  assign new_B1563_ = new_B1564_ ^ new_B1554_;
  assign new_B1564_ = new_B1572_ & new_B1571_;
  assign new_B1565_ = new_B1570_ & new_B1554_;
  assign new_B1566_ = new_B1575_ & new_B1574_;
  assign new_B1567_ = new_B1573_ & new_B1554_;
  assign new_B1568_ = new_B1576_ | new_B1553_;
  assign new_B1569_ = ~new_B1554_ ^ new_B1566_;
  assign new_B1570_ = ~new_B1579_ | ~new_B1580_;
  assign new_B1571_ = new_B1555_ ^ new_B1562_;
  assign new_B1572_ = new_B1581_ & new_B1574_;
  assign new_B1573_ = ~new_B1583_ | ~new_B1582_;
  assign new_B1574_ = new_B1555_ | new_B1556_;
  assign new_B1575_ = new_B1555_ | new_B1562_;
  assign new_B1576_ = new_B1554_ & new_B1566_;
  assign new_B1577_ = ~new_B1553_ | ~new_B1554_;
  assign new_B1578_ = new_B1562_ & new_B1577_;
  assign new_B1579_ = ~new_B1578_ & ~new_B1562_;
  assign new_B1580_ = new_B1562_ | new_B1577_;
  assign new_B1581_ = ~new_B1555_ | ~new_B1556_;
  assign new_B1582_ = new_B1562_ | new_B1577_;
  assign new_B1583_ = ~new_B1562_ & ~new_B1584_;
  assign new_B1584_ = new_B1562_ & new_B1577_;
  assign new_B1585_ = new_B7827_;
  assign new_B1586_ = new_B7860_;
  assign new_B1587_ = new_B7893_;
  assign new_B1588_ = new_B7926_;
  assign new_B1589_ = new_B7959_;
  assign new_B1590_ = new_B1596_ & new_B1595_;
  assign new_B1591_ = new_B1598_ | new_B1597_;
  assign new_B1592_ = new_B1600_ | new_B1599_;
  assign new_B1593_ = new_B1595_ & new_B1601_;
  assign new_B1594_ = new_B1595_ & new_B1602_;
  assign new_B1595_ = new_B1585_ ^ new_B1586_;
  assign new_B1596_ = new_B1597_ ^ new_B1587_;
  assign new_B1597_ = new_B1605_ & new_B1604_;
  assign new_B1598_ = new_B1603_ & new_B1587_;
  assign new_B1599_ = new_B1608_ & new_B1607_;
  assign new_B1600_ = new_B1606_ & new_B1587_;
  assign new_B1601_ = new_B1609_ | new_B1586_;
  assign new_B1602_ = ~new_B1587_ ^ new_B1599_;
  assign new_B1603_ = ~new_B1612_ | ~new_B1613_;
  assign new_B1604_ = new_B1588_ ^ new_B1595_;
  assign new_B1605_ = new_B1614_ & new_B1607_;
  assign new_B1606_ = ~new_B1616_ | ~new_B1615_;
  assign new_B1607_ = new_B1588_ | new_B1589_;
  assign new_B1608_ = new_B1588_ | new_B1595_;
  assign new_B1609_ = new_B1587_ & new_B1599_;
  assign new_B1610_ = ~new_B1586_ | ~new_B1587_;
  assign new_B1611_ = new_B1595_ & new_B1610_;
  assign new_B1612_ = ~new_B1611_ & ~new_B1595_;
  assign new_B1613_ = new_B1595_ | new_B1610_;
  assign new_B1614_ = ~new_B1588_ | ~new_B1589_;
  assign new_B1615_ = new_B1595_ | new_B1610_;
  assign new_B1616_ = ~new_B1595_ & ~new_B1617_;
  assign new_B1617_ = new_B1595_ & new_B1610_;
  assign new_B1618_ = new_B7992_;
  assign new_B1619_ = new_B8025_;
  assign new_B1620_ = new_B8058_;
  assign new_B1621_ = new_B8091_;
  assign new_B1622_ = new_B8124_;
  assign new_B1623_ = new_B1629_ & new_B1628_;
  assign new_B1624_ = new_B1631_ | new_B1630_;
  assign new_B1625_ = new_B1633_ | new_B1632_;
  assign new_B1626_ = new_B1628_ & new_B1634_;
  assign new_B1627_ = new_B1628_ & new_B1635_;
  assign new_B1628_ = new_B1618_ ^ new_B1619_;
  assign new_B1629_ = new_B1630_ ^ new_B1620_;
  assign new_B1630_ = new_B1638_ & new_B1637_;
  assign new_B1631_ = new_B1636_ & new_B1620_;
  assign new_B1632_ = new_B1641_ & new_B1640_;
  assign new_B1633_ = new_B1639_ & new_B1620_;
  assign new_B1634_ = new_B1642_ | new_B1619_;
  assign new_B1635_ = ~new_B1620_ ^ new_B1632_;
  assign new_B1636_ = ~new_B1645_ | ~new_B1646_;
  assign new_B1637_ = new_B1621_ ^ new_B1628_;
  assign new_B1638_ = new_B1647_ & new_B1640_;
  assign new_B1639_ = ~new_B1649_ | ~new_B1648_;
  assign new_B1640_ = new_B1621_ | new_B1622_;
  assign new_B1641_ = new_B1621_ | new_B1628_;
  assign new_B1642_ = new_B1620_ & new_B1632_;
  assign new_B1643_ = ~new_B1619_ | ~new_B1620_;
  assign new_B1644_ = new_B1628_ & new_B1643_;
  assign new_B1645_ = ~new_B1644_ & ~new_B1628_;
  assign new_B1646_ = new_B1628_ | new_B1643_;
  assign new_B1647_ = ~new_B1621_ | ~new_B1622_;
  assign new_B1648_ = new_B1628_ | new_B1643_;
  assign new_B1649_ = ~new_B1628_ & ~new_B1650_;
  assign new_B1650_ = new_B1628_ & new_B1643_;
  assign new_B1651_ = new_B8157_;
  assign new_B1652_ = new_B8190_;
  assign new_B1653_ = new_B8223_;
  assign new_B1654_ = new_B8256_;
  assign new_B1655_ = new_B8289_;
  assign new_B1656_ = new_B1662_ & new_B1661_;
  assign new_B1657_ = new_B1664_ | new_B1663_;
  assign new_B1658_ = new_B1666_ | new_B1665_;
  assign new_B1659_ = new_B1661_ & new_B1667_;
  assign new_B1660_ = new_B1661_ & new_B1668_;
  assign new_B1661_ = new_B1651_ ^ new_B1652_;
  assign new_B1662_ = new_B1663_ ^ new_B1653_;
  assign new_B1663_ = new_B1671_ & new_B1670_;
  assign new_B1664_ = new_B1669_ & new_B1653_;
  assign new_B1665_ = new_B1674_ & new_B1673_;
  assign new_B1666_ = new_B1672_ & new_B1653_;
  assign new_B1667_ = new_B1675_ | new_B1652_;
  assign new_B1668_ = ~new_B1653_ ^ new_B1665_;
  assign new_B1669_ = ~new_B1678_ | ~new_B1679_;
  assign new_B1670_ = new_B1654_ ^ new_B1661_;
  assign new_B1671_ = new_B1680_ & new_B1673_;
  assign new_B1672_ = ~new_B1682_ | ~new_B1681_;
  assign new_B1673_ = new_B1654_ | new_B1655_;
  assign new_B1674_ = new_B1654_ | new_B1661_;
  assign new_B1675_ = new_B1653_ & new_B1665_;
  assign new_B1676_ = ~new_B1652_ | ~new_B1653_;
  assign new_B1677_ = new_B1661_ & new_B1676_;
  assign new_B1678_ = ~new_B1677_ & ~new_B1661_;
  assign new_B1679_ = new_B1661_ | new_B1676_;
  assign new_B1680_ = ~new_B1654_ | ~new_B1655_;
  assign new_B1681_ = new_B1661_ | new_B1676_;
  assign new_B1682_ = ~new_B1661_ & ~new_B1683_;
  assign new_B1683_ = new_B1661_ & new_B1676_;
  assign new_B1684_ = new_B8322_;
  assign new_B1685_ = new_B8355_;
  assign new_B1686_ = new_B8388_;
  assign new_B1687_ = new_B8421_;
  assign new_B1688_ = new_B8454_;
  assign new_B1689_ = new_B1695_ & new_B1694_;
  assign new_B1690_ = new_B1697_ | new_B1696_;
  assign new_B1691_ = new_B1699_ | new_B1698_;
  assign new_B1692_ = new_B1694_ & new_B1700_;
  assign new_B1693_ = new_B1694_ & new_B1701_;
  assign new_B1694_ = new_B1684_ ^ new_B1685_;
  assign new_B1695_ = new_B1696_ ^ new_B1686_;
  assign new_B1696_ = new_B1704_ & new_B1703_;
  assign new_B1697_ = new_B1702_ & new_B1686_;
  assign new_B1698_ = new_B1707_ & new_B1706_;
  assign new_B1699_ = new_B1705_ & new_B1686_;
  assign new_B1700_ = new_B1708_ | new_B1685_;
  assign new_B1701_ = ~new_B1686_ ^ new_B1698_;
  assign new_B1702_ = ~new_B1711_ | ~new_B1712_;
  assign new_B1703_ = new_B1687_ ^ new_B1694_;
  assign new_B1704_ = new_B1713_ & new_B1706_;
  assign new_B1705_ = ~new_B1715_ | ~new_B1714_;
  assign new_B1706_ = new_B1687_ | new_B1688_;
  assign new_B1707_ = new_B1687_ | new_B1694_;
  assign new_B1708_ = new_B1686_ & new_B1698_;
  assign new_B1709_ = ~new_B1685_ | ~new_B1686_;
  assign new_B1710_ = new_B1694_ & new_B1709_;
  assign new_B1711_ = ~new_B1710_ & ~new_B1694_;
  assign new_B1712_ = new_B1694_ | new_B1709_;
  assign new_B1713_ = ~new_B1687_ | ~new_B1688_;
  assign new_B1714_ = new_B1694_ | new_B1709_;
  assign new_B1715_ = ~new_B1694_ & ~new_B1716_;
  assign new_B1716_ = new_B1694_ & new_B1709_;
  assign new_B1717_ = new_B8487_;
  assign new_B1718_ = new_B8520_;
  assign new_B1719_ = new_B8553_;
  assign new_B1720_ = new_B8586_;
  assign new_B1721_ = new_B8619_;
  assign new_B1722_ = new_B1728_ & new_B1727_;
  assign new_B1723_ = new_B1730_ | new_B1729_;
  assign new_B1724_ = new_B1732_ | new_B1731_;
  assign new_B1725_ = new_B1727_ & new_B1733_;
  assign new_B1726_ = new_B1727_ & new_B1734_;
  assign new_B1727_ = new_B1717_ ^ new_B1718_;
  assign new_B1728_ = new_B1729_ ^ new_B1719_;
  assign new_B1729_ = new_B1737_ & new_B1736_;
  assign new_B1730_ = new_B1735_ & new_B1719_;
  assign new_B1731_ = new_B1740_ & new_B1739_;
  assign new_B1732_ = new_B1738_ & new_B1719_;
  assign new_B1733_ = new_B1741_ | new_B1718_;
  assign new_B1734_ = ~new_B1719_ ^ new_B1731_;
  assign new_B1735_ = ~new_B1744_ | ~new_B1745_;
  assign new_B1736_ = new_B1720_ ^ new_B1727_;
  assign new_B1737_ = new_B1746_ & new_B1739_;
  assign new_B1738_ = ~new_B1748_ | ~new_B1747_;
  assign new_B1739_ = new_B1720_ | new_B1721_;
  assign new_B1740_ = new_B1720_ | new_B1727_;
  assign new_B1741_ = new_B1719_ & new_B1731_;
  assign new_B1742_ = ~new_B1718_ | ~new_B1719_;
  assign new_B1743_ = new_B1727_ & new_B1742_;
  assign new_B1744_ = ~new_B1743_ & ~new_B1727_;
  assign new_B1745_ = new_B1727_ | new_B1742_;
  assign new_B1746_ = ~new_B1720_ | ~new_B1721_;
  assign new_B1747_ = new_B1727_ | new_B1742_;
  assign new_B1748_ = ~new_B1727_ & ~new_B1749_;
  assign new_B1749_ = new_B1727_ & new_B1742_;
  assign new_B1750_ = new_B8652_;
  assign new_B1751_ = new_B8685_;
  assign new_B1752_ = new_B8718_;
  assign new_B1753_ = new_B8751_;
  assign new_B1754_ = new_B8784_;
  assign new_B1755_ = new_B1761_ & new_B1760_;
  assign new_B1756_ = new_B1763_ | new_B1762_;
  assign new_B1757_ = new_B1765_ | new_B1764_;
  assign new_B1758_ = new_B1760_ & new_B1766_;
  assign new_B1759_ = new_B1760_ & new_B1767_;
  assign new_B1760_ = new_B1750_ ^ new_B1751_;
  assign new_B1761_ = new_B1762_ ^ new_B1752_;
  assign new_B1762_ = new_B1770_ & new_B1769_;
  assign new_B1763_ = new_B1768_ & new_B1752_;
  assign new_B1764_ = new_B1773_ & new_B1772_;
  assign new_B1765_ = new_B1771_ & new_B1752_;
  assign new_B1766_ = new_B1774_ | new_B1751_;
  assign new_B1767_ = ~new_B1752_ ^ new_B1764_;
  assign new_B1768_ = ~new_B1777_ | ~new_B1778_;
  assign new_B1769_ = new_B1753_ ^ new_B1760_;
  assign new_B1770_ = new_B1779_ & new_B1772_;
  assign new_B1771_ = ~new_B1781_ | ~new_B1780_;
  assign new_B1772_ = new_B1753_ | new_B1754_;
  assign new_B1773_ = new_B1753_ | new_B1760_;
  assign new_B1774_ = new_B1752_ & new_B1764_;
  assign new_B1775_ = ~new_B1751_ | ~new_B1752_;
  assign new_B1776_ = new_B1760_ & new_B1775_;
  assign new_B1777_ = ~new_B1776_ & ~new_B1760_;
  assign new_B1778_ = new_B1760_ | new_B1775_;
  assign new_B1779_ = ~new_B1753_ | ~new_B1754_;
  assign new_B1780_ = new_B1760_ | new_B1775_;
  assign new_B1781_ = ~new_B1760_ & ~new_B1782_;
  assign new_B1782_ = new_B1760_ & new_B1775_;
  assign new_B1783_ = new_B8817_;
  assign new_B1784_ = new_B8850_;
  assign new_B1785_ = new_B8883_;
  assign new_B1786_ = new_B8916_;
  assign new_B1787_ = new_B8949_;
  assign new_B1788_ = new_B1794_ & new_B1793_;
  assign new_B1789_ = new_B1796_ | new_B1795_;
  assign new_B1790_ = new_B1798_ | new_B1797_;
  assign new_B1791_ = new_B1793_ & new_B1799_;
  assign new_B1792_ = new_B1793_ & new_B1800_;
  assign new_B1793_ = new_B1783_ ^ new_B1784_;
  assign new_B1794_ = new_B1795_ ^ new_B1785_;
  assign new_B1795_ = new_B1803_ & new_B1802_;
  assign new_B1796_ = new_B1801_ & new_B1785_;
  assign new_B1797_ = new_B1806_ & new_B1805_;
  assign new_B1798_ = new_B1804_ & new_B1785_;
  assign new_B1799_ = new_B1807_ | new_B1784_;
  assign new_B1800_ = ~new_B1785_ ^ new_B1797_;
  assign new_B1801_ = ~new_B1810_ | ~new_B1811_;
  assign new_B1802_ = new_B1786_ ^ new_B1793_;
  assign new_B1803_ = new_B1812_ & new_B1805_;
  assign new_B1804_ = ~new_B1814_ | ~new_B1813_;
  assign new_B1805_ = new_B1786_ | new_B1787_;
  assign new_B1806_ = new_B1786_ | new_B1793_;
  assign new_B1807_ = new_B1785_ & new_B1797_;
  assign new_B1808_ = ~new_B1784_ | ~new_B1785_;
  assign new_B1809_ = new_B1793_ & new_B1808_;
  assign new_B1810_ = ~new_B1809_ & ~new_B1793_;
  assign new_B1811_ = new_B1793_ | new_B1808_;
  assign new_B1812_ = ~new_B1786_ | ~new_B1787_;
  assign new_B1813_ = new_B1793_ | new_B1808_;
  assign new_B1814_ = ~new_B1793_ & ~new_B1815_;
  assign new_B1815_ = new_B1793_ & new_B1808_;
  assign new_B1816_ = new_B8982_;
  assign new_B1817_ = new_B9015_;
  assign new_B1818_ = new_B9048_;
  assign new_B1819_ = new_B9081_;
  assign new_B1820_ = new_B9114_;
  assign new_B1821_ = new_B1827_ & new_B1826_;
  assign new_B1822_ = new_B1829_ | new_B1828_;
  assign new_B1823_ = new_B1831_ | new_B1830_;
  assign new_B1824_ = new_B1826_ & new_B1832_;
  assign new_B1825_ = new_B1826_ & new_B1833_;
  assign new_B1826_ = new_B1816_ ^ new_B1817_;
  assign new_B1827_ = new_B1828_ ^ new_B1818_;
  assign new_B1828_ = new_B1836_ & new_B1835_;
  assign new_B1829_ = new_B1834_ & new_B1818_;
  assign new_B1830_ = new_B1839_ & new_B1838_;
  assign new_B1831_ = new_B1837_ & new_B1818_;
  assign new_B1832_ = new_B1840_ | new_B1817_;
  assign new_B1833_ = ~new_B1818_ ^ new_B1830_;
  assign new_B1834_ = ~new_B1843_ | ~new_B1844_;
  assign new_B1835_ = new_B1819_ ^ new_B1826_;
  assign new_B1836_ = new_B1845_ & new_B1838_;
  assign new_B1837_ = ~new_B1847_ | ~new_B1846_;
  assign new_B1838_ = new_B1819_ | new_B1820_;
  assign new_B1839_ = new_B1819_ | new_B1826_;
  assign new_B1840_ = new_B1818_ & new_B1830_;
  assign new_B1841_ = ~new_B1817_ | ~new_B1818_;
  assign new_B1842_ = new_B1826_ & new_B1841_;
  assign new_B1843_ = ~new_B1842_ & ~new_B1826_;
  assign new_B1844_ = new_B1826_ | new_B1841_;
  assign new_B1845_ = ~new_B1819_ | ~new_B1820_;
  assign new_B1846_ = new_B1826_ | new_B1841_;
  assign new_B1847_ = ~new_B1826_ & ~new_B1848_;
  assign new_B1848_ = new_B1826_ & new_B1841_;
  assign new_B1849_ = new_B9147_;
  assign new_B1850_ = new_B9180_;
  assign new_B1851_ = new_B9213_;
  assign new_B1852_ = new_B9246_;
  assign new_B1853_ = new_B9279_;
  assign new_B1854_ = new_B1860_ & new_B1859_;
  assign new_B1855_ = new_B1862_ | new_B1861_;
  assign new_B1856_ = new_B1864_ | new_B1863_;
  assign new_B1857_ = new_B1859_ & new_B1865_;
  assign new_B1858_ = new_B1859_ & new_B1866_;
  assign new_B1859_ = new_B1849_ ^ new_B1850_;
  assign new_B1860_ = new_B1861_ ^ new_B1851_;
  assign new_B1861_ = new_B1869_ & new_B1868_;
  assign new_B1862_ = new_B1867_ & new_B1851_;
  assign new_B1863_ = new_B1872_ & new_B1871_;
  assign new_B1864_ = new_B1870_ & new_B1851_;
  assign new_B1865_ = new_B1873_ | new_B1850_;
  assign new_B1866_ = ~new_B1851_ ^ new_B1863_;
  assign new_B1867_ = ~new_B1876_ | ~new_B1877_;
  assign new_B1868_ = new_B1852_ ^ new_B1859_;
  assign new_B1869_ = new_B1878_ & new_B1871_;
  assign new_B1870_ = ~new_B1880_ | ~new_B1879_;
  assign new_B1871_ = new_B1852_ | new_B1853_;
  assign new_B1872_ = new_B1852_ | new_B1859_;
  assign new_B1873_ = new_B1851_ & new_B1863_;
  assign new_B1874_ = ~new_B1850_ | ~new_B1851_;
  assign new_B1875_ = new_B1859_ & new_B1874_;
  assign new_B1876_ = ~new_B1875_ & ~new_B1859_;
  assign new_B1877_ = new_B1859_ | new_B1874_;
  assign new_B1878_ = ~new_B1852_ | ~new_B1853_;
  assign new_B1879_ = new_B1859_ | new_B1874_;
  assign new_B1880_ = ~new_B1859_ & ~new_B1881_;
  assign new_B1881_ = new_B1859_ & new_B1874_;
  assign new_B1882_ = new_B5190_;
  assign new_B1883_ = new_B5221_;
  assign new_B1884_ = new_B5254_;
  assign new_B1885_ = new_B5287_;
  assign new_B1886_ = new_B5320_;
  assign new_B1887_ = new_B1893_ & new_B1892_;
  assign new_B1888_ = new_B1895_ | new_B1894_;
  assign new_B1889_ = new_B1897_ | new_B1896_;
  assign new_B1890_ = new_B1892_ & new_B1898_;
  assign new_B1891_ = new_B1892_ & new_B1899_;
  assign new_B1892_ = new_B1882_ ^ new_B1883_;
  assign new_B1893_ = new_B1894_ ^ new_B1884_;
  assign new_B1894_ = new_B1902_ & new_B1901_;
  assign new_B1895_ = new_B1900_ & new_B1884_;
  assign new_B1896_ = new_B1905_ & new_B1904_;
  assign new_B1897_ = new_B1903_ & new_B1884_;
  assign new_B1898_ = new_B1906_ | new_B1883_;
  assign new_B1899_ = ~new_B1884_ ^ new_B1896_;
  assign new_B1900_ = ~new_B1909_ | ~new_B1910_;
  assign new_B1901_ = new_B1885_ ^ new_B1892_;
  assign new_B1902_ = new_B1911_ & new_B1904_;
  assign new_B1903_ = ~new_B1913_ | ~new_B1912_;
  assign new_B1904_ = new_B1885_ | new_B1886_;
  assign new_B1905_ = new_B1885_ | new_B1892_;
  assign new_B1906_ = new_B1884_ & new_B1896_;
  assign new_B1907_ = ~new_B1883_ | ~new_B1884_;
  assign new_B1908_ = new_B1892_ & new_B1907_;
  assign new_B1909_ = ~new_B1908_ & ~new_B1892_;
  assign new_B1910_ = new_B1892_ | new_B1907_;
  assign new_B1911_ = ~new_B1885_ | ~new_B1886_;
  assign new_B1912_ = new_B1892_ | new_B1907_;
  assign new_B1913_ = ~new_B1892_ & ~new_B1914_;
  assign new_B1914_ = new_B1892_ & new_B1907_;
  assign new_B1915_ = new_B5353_;
  assign new_B1916_ = new_B5386_;
  assign new_B1917_ = new_B5419_;
  assign new_B1918_ = new_B5452_;
  assign new_B1919_ = new_B5485_;
  assign new_B1920_ = new_B1926_ & new_B1925_;
  assign new_B1921_ = new_B1928_ | new_B1927_;
  assign new_B1922_ = new_B1930_ | new_B1929_;
  assign new_B1923_ = new_B1925_ & new_B1931_;
  assign new_B1924_ = new_B1925_ & new_B1932_;
  assign new_B1925_ = new_B1915_ ^ new_B1916_;
  assign new_B1926_ = new_B1927_ ^ new_B1917_;
  assign new_B1927_ = new_B1935_ & new_B1934_;
  assign new_B1928_ = new_B1933_ & new_B1917_;
  assign new_B1929_ = new_B1938_ & new_B1937_;
  assign new_B1930_ = new_B1936_ & new_B1917_;
  assign new_B1931_ = new_B1939_ | new_B1916_;
  assign new_B1932_ = ~new_B1917_ ^ new_B1929_;
  assign new_B1933_ = ~new_B1942_ | ~new_B1943_;
  assign new_B1934_ = new_B1918_ ^ new_B1925_;
  assign new_B1935_ = new_B1944_ & new_B1937_;
  assign new_B1936_ = ~new_B1946_ | ~new_B1945_;
  assign new_B1937_ = new_B1918_ | new_B1919_;
  assign new_B1938_ = new_B1918_ | new_B1925_;
  assign new_B1939_ = new_B1917_ & new_B1929_;
  assign new_B1940_ = ~new_B1916_ | ~new_B1917_;
  assign new_B1941_ = new_B1925_ & new_B1940_;
  assign new_B1942_ = ~new_B1941_ & ~new_B1925_;
  assign new_B1943_ = new_B1925_ | new_B1940_;
  assign new_B1944_ = ~new_B1918_ | ~new_B1919_;
  assign new_B1945_ = new_B1925_ | new_B1940_;
  assign new_B1946_ = ~new_B1925_ & ~new_B1947_;
  assign new_B1947_ = new_B1925_ & new_B1940_;
  assign new_B1948_ = new_B5518_;
  assign new_B1949_ = new_B5551_;
  assign new_B1950_ = new_B5584_;
  assign new_B1951_ = new_B5617_;
  assign new_B1952_ = new_B5650_;
  assign new_B1953_ = new_B1959_ & new_B1958_;
  assign new_B1954_ = new_B1961_ | new_B1960_;
  assign new_B1955_ = new_B1963_ | new_B1962_;
  assign new_B1956_ = new_B1958_ & new_B1964_;
  assign new_B1957_ = new_B1958_ & new_B1965_;
  assign new_B1958_ = new_B1948_ ^ new_B1949_;
  assign new_B1959_ = new_B1960_ ^ new_B1950_;
  assign new_B1960_ = new_B1968_ & new_B1967_;
  assign new_B1961_ = new_B1966_ & new_B1950_;
  assign new_B1962_ = new_B1971_ & new_B1970_;
  assign new_B1963_ = new_B1969_ & new_B1950_;
  assign new_B1964_ = new_B1972_ | new_B1949_;
  assign new_B1965_ = ~new_B1950_ ^ new_B1962_;
  assign new_B1966_ = ~new_B1975_ | ~new_B1976_;
  assign new_B1967_ = new_B1951_ ^ new_B1958_;
  assign new_B1968_ = new_B1977_ & new_B1970_;
  assign new_B1969_ = ~new_B1979_ | ~new_B1978_;
  assign new_B1970_ = new_B1951_ | new_B1952_;
  assign new_B1971_ = new_B1951_ | new_B1958_;
  assign new_B1972_ = new_B1950_ & new_B1962_;
  assign new_B1973_ = ~new_B1949_ | ~new_B1950_;
  assign new_B1974_ = new_B1958_ & new_B1973_;
  assign new_B1975_ = ~new_B1974_ & ~new_B1958_;
  assign new_B1976_ = new_B1958_ | new_B1973_;
  assign new_B1977_ = ~new_B1951_ | ~new_B1952_;
  assign new_B1978_ = new_B1958_ | new_B1973_;
  assign new_B1979_ = ~new_B1958_ & ~new_B1980_;
  assign new_B1980_ = new_B1958_ & new_B1973_;
  assign new_B1981_ = new_B5683_;
  assign new_B1982_ = new_B5716_;
  assign new_B1983_ = new_B5749_;
  assign new_B1984_ = new_B5782_;
  assign new_B1985_ = new_B5815_;
  assign new_B1986_ = new_B1992_ & new_B1991_;
  assign new_B1987_ = new_B1994_ | new_B1993_;
  assign new_B1988_ = new_B1996_ | new_B1995_;
  assign new_B1989_ = new_B1991_ & new_B1997_;
  assign new_B1990_ = new_B1991_ & new_B1998_;
  assign new_B1991_ = new_B1981_ ^ new_B1982_;
  assign new_B1992_ = new_B1993_ ^ new_B1983_;
  assign new_B1993_ = new_B2001_ & new_B2000_;
  assign new_B1994_ = new_B1999_ & new_B1983_;
  assign new_B1995_ = new_B2004_ & new_B2003_;
  assign new_B1996_ = new_B2002_ & new_B1983_;
  assign new_B1997_ = new_B2005_ | new_B1982_;
  assign new_B1998_ = ~new_B1983_ ^ new_B1995_;
  assign new_B1999_ = ~new_B2008_ | ~new_B2009_;
  assign new_B2000_ = new_B1984_ ^ new_B1991_;
  assign new_B2001_ = new_B2010_ & new_B2003_;
  assign new_B2002_ = ~new_B2012_ | ~new_B2011_;
  assign new_B2003_ = new_B1984_ | new_B1985_;
  assign new_B2004_ = new_B1984_ | new_B1991_;
  assign new_B2005_ = new_B1983_ & new_B1995_;
  assign new_B2006_ = ~new_B1982_ | ~new_B1983_;
  assign new_B2007_ = new_B1991_ & new_B2006_;
  assign new_B2008_ = ~new_B2007_ & ~new_B1991_;
  assign new_B2009_ = new_B1991_ | new_B2006_;
  assign new_B2010_ = ~new_B1984_ | ~new_B1985_;
  assign new_B2011_ = new_B1991_ | new_B2006_;
  assign new_B2012_ = ~new_B1991_ & ~new_B2013_;
  assign new_B2013_ = new_B1991_ & new_B2006_;
  assign new_B2014_ = new_B5848_;
  assign new_B2015_ = new_B5881_;
  assign new_B2016_ = new_B5914_;
  assign new_B2017_ = new_B5947_;
  assign new_B2018_ = new_B5980_;
  assign new_B2019_ = new_B2025_ & new_B2024_;
  assign new_B2020_ = new_B2027_ | new_B2026_;
  assign new_B2021_ = new_B2029_ | new_B2028_;
  assign new_B2022_ = new_B2024_ & new_B2030_;
  assign new_B2023_ = new_B2024_ & new_B2031_;
  assign new_B2024_ = new_B2014_ ^ new_B2015_;
  assign new_B2025_ = new_B2026_ ^ new_B2016_;
  assign new_B2026_ = new_B2034_ & new_B2033_;
  assign new_B2027_ = new_B2032_ & new_B2016_;
  assign new_B2028_ = new_B2037_ & new_B2036_;
  assign new_B2029_ = new_B2035_ & new_B2016_;
  assign new_B2030_ = new_B2038_ | new_B2015_;
  assign new_B2031_ = ~new_B2016_ ^ new_B2028_;
  assign new_B2032_ = ~new_B2041_ | ~new_B2042_;
  assign new_B2033_ = new_B2017_ ^ new_B2024_;
  assign new_B2034_ = new_B2043_ & new_B2036_;
  assign new_B2035_ = ~new_B2045_ | ~new_B2044_;
  assign new_B2036_ = new_B2017_ | new_B2018_;
  assign new_B2037_ = new_B2017_ | new_B2024_;
  assign new_B2038_ = new_B2016_ & new_B2028_;
  assign new_B2039_ = ~new_B2015_ | ~new_B2016_;
  assign new_B2040_ = new_B2024_ & new_B2039_;
  assign new_B2041_ = ~new_B2040_ & ~new_B2024_;
  assign new_B2042_ = new_B2024_ | new_B2039_;
  assign new_B2043_ = ~new_B2017_ | ~new_B2018_;
  assign new_B2044_ = new_B2024_ | new_B2039_;
  assign new_B2045_ = ~new_B2024_ & ~new_B2046_;
  assign new_B2046_ = new_B2024_ & new_B2039_;
  assign new_B2047_ = new_B6013_;
  assign new_B2048_ = new_B6046_;
  assign new_B2049_ = new_B6079_;
  assign new_B2050_ = new_B6112_;
  assign new_B2051_ = new_B6145_;
  assign new_B2052_ = new_B2058_ & new_B2057_;
  assign new_B2053_ = new_B2060_ | new_B2059_;
  assign new_B2054_ = new_B2062_ | new_B2061_;
  assign new_B2055_ = new_B2057_ & new_B2063_;
  assign new_B2056_ = new_B2057_ & new_B2064_;
  assign new_B2057_ = new_B2047_ ^ new_B2048_;
  assign new_B2058_ = new_B2059_ ^ new_B2049_;
  assign new_B2059_ = new_B2067_ & new_B2066_;
  assign new_B2060_ = new_B2065_ & new_B2049_;
  assign new_B2061_ = new_B2070_ & new_B2069_;
  assign new_B2062_ = new_B2068_ & new_B2049_;
  assign new_B2063_ = new_B2071_ | new_B2048_;
  assign new_B2064_ = ~new_B2049_ ^ new_B2061_;
  assign new_B2065_ = ~new_B2074_ | ~new_B2075_;
  assign new_B2066_ = new_B2050_ ^ new_B2057_;
  assign new_B2067_ = new_B2076_ & new_B2069_;
  assign new_B2068_ = ~new_B2078_ | ~new_B2077_;
  assign new_B2069_ = new_B2050_ | new_B2051_;
  assign new_B2070_ = new_B2050_ | new_B2057_;
  assign new_B2071_ = new_B2049_ & new_B2061_;
  assign new_B2072_ = ~new_B2048_ | ~new_B2049_;
  assign new_B2073_ = new_B2057_ & new_B2072_;
  assign new_B2074_ = ~new_B2073_ & ~new_B2057_;
  assign new_B2075_ = new_B2057_ | new_B2072_;
  assign new_B2076_ = ~new_B2050_ | ~new_B2051_;
  assign new_B2077_ = new_B2057_ | new_B2072_;
  assign new_B2078_ = ~new_B2057_ & ~new_B2079_;
  assign new_B2079_ = new_B2057_ & new_B2072_;
  assign new_B2080_ = new_B6178_;
  assign new_B2081_ = new_B6211_;
  assign new_B2082_ = new_B6244_;
  assign new_B2083_ = new_B6277_;
  assign new_B2084_ = new_B6310_;
  assign new_B2085_ = new_B2091_ & new_B2090_;
  assign new_B2086_ = new_B2093_ | new_B2092_;
  assign new_B2087_ = new_B2095_ | new_B2094_;
  assign new_B2088_ = new_B2090_ & new_B2096_;
  assign new_B2089_ = new_B2090_ & new_B2097_;
  assign new_B2090_ = new_B2080_ ^ new_B2081_;
  assign new_B2091_ = new_B2092_ ^ new_B2082_;
  assign new_B2092_ = new_B2100_ & new_B2099_;
  assign new_B2093_ = new_B2098_ & new_B2082_;
  assign new_B2094_ = new_B2103_ & new_B2102_;
  assign new_B2095_ = new_B2101_ & new_B2082_;
  assign new_B2096_ = new_B2104_ | new_B2081_;
  assign new_B2097_ = ~new_B2082_ ^ new_B2094_;
  assign new_B2098_ = ~new_B2107_ | ~new_B2108_;
  assign new_B2099_ = new_B2083_ ^ new_B2090_;
  assign new_B2100_ = new_B2109_ & new_B2102_;
  assign new_B2101_ = ~new_B2111_ | ~new_B2110_;
  assign new_B2102_ = new_B2083_ | new_B2084_;
  assign new_B2103_ = new_B2083_ | new_B2090_;
  assign new_B2104_ = new_B2082_ & new_B2094_;
  assign new_B2105_ = ~new_B2081_ | ~new_B2082_;
  assign new_B2106_ = new_B2090_ & new_B2105_;
  assign new_B2107_ = ~new_B2106_ & ~new_B2090_;
  assign new_B2108_ = new_B2090_ | new_B2105_;
  assign new_B2109_ = ~new_B2083_ | ~new_B2084_;
  assign new_B2110_ = new_B2090_ | new_B2105_;
  assign new_B2111_ = ~new_B2090_ & ~new_B2112_;
  assign new_B2112_ = new_B2090_ & new_B2105_;
  assign new_B2113_ = new_B6343_;
  assign new_B2114_ = new_B6376_;
  assign new_B2115_ = new_B6409_;
  assign new_B2116_ = new_B6442_;
  assign new_B2117_ = new_B6475_;
  assign new_B2118_ = new_B2124_ & new_B2123_;
  assign new_B2119_ = new_B2126_ | new_B2125_;
  assign new_B2120_ = new_B2128_ | new_B2127_;
  assign new_B2121_ = new_B2123_ & new_B2129_;
  assign new_B2122_ = new_B2123_ & new_B2130_;
  assign new_B2123_ = new_B2113_ ^ new_B2114_;
  assign new_B2124_ = new_B2125_ ^ new_B2115_;
  assign new_B2125_ = new_B2133_ & new_B2132_;
  assign new_B2126_ = new_B2131_ & new_B2115_;
  assign new_B2127_ = new_B2136_ & new_B2135_;
  assign new_B2128_ = new_B2134_ & new_B2115_;
  assign new_B2129_ = new_B2137_ | new_B2114_;
  assign new_B2130_ = ~new_B2115_ ^ new_B2127_;
  assign new_B2131_ = ~new_B2140_ | ~new_B2141_;
  assign new_B2132_ = new_B2116_ ^ new_B2123_;
  assign new_B2133_ = new_B2142_ & new_B2135_;
  assign new_B2134_ = ~new_B2144_ | ~new_B2143_;
  assign new_B2135_ = new_B2116_ | new_B2117_;
  assign new_B2136_ = new_B2116_ | new_B2123_;
  assign new_B2137_ = new_B2115_ & new_B2127_;
  assign new_B2138_ = ~new_B2114_ | ~new_B2115_;
  assign new_B2139_ = new_B2123_ & new_B2138_;
  assign new_B2140_ = ~new_B2139_ & ~new_B2123_;
  assign new_B2141_ = new_B2123_ | new_B2138_;
  assign new_B2142_ = ~new_B2116_ | ~new_B2117_;
  assign new_B2143_ = new_B2123_ | new_B2138_;
  assign new_B2144_ = ~new_B2123_ & ~new_B2145_;
  assign new_B2145_ = new_B2123_ & new_B2138_;
  assign new_B2146_ = new_B6508_;
  assign new_B2147_ = new_B6541_;
  assign new_B2148_ = new_B6574_;
  assign new_B2149_ = new_B6607_;
  assign new_B2150_ = new_B6640_;
  assign new_B2151_ = new_B2157_ & new_B2156_;
  assign new_B2152_ = new_B2159_ | new_B2158_;
  assign new_B2153_ = new_B2161_ | new_B2160_;
  assign new_B2154_ = new_B2156_ & new_B2162_;
  assign new_B2155_ = new_B2156_ & new_B2163_;
  assign new_B2156_ = new_B2146_ ^ new_B2147_;
  assign new_B2157_ = new_B2158_ ^ new_B2148_;
  assign new_B2158_ = new_B2166_ & new_B2165_;
  assign new_B2159_ = new_B2164_ & new_B2148_;
  assign new_B2160_ = new_B2169_ & new_B2168_;
  assign new_B2161_ = new_B2167_ & new_B2148_;
  assign new_B2162_ = new_B2170_ | new_B2147_;
  assign new_B2163_ = ~new_B2148_ ^ new_B2160_;
  assign new_B2164_ = ~new_B2173_ | ~new_B2174_;
  assign new_B2165_ = new_B2149_ ^ new_B2156_;
  assign new_B2166_ = new_B2175_ & new_B2168_;
  assign new_B2167_ = ~new_B2177_ | ~new_B2176_;
  assign new_B2168_ = new_B2149_ | new_B2150_;
  assign new_B2169_ = new_B2149_ | new_B2156_;
  assign new_B2170_ = new_B2148_ & new_B2160_;
  assign new_B2171_ = ~new_B2147_ | ~new_B2148_;
  assign new_B2172_ = new_B2156_ & new_B2171_;
  assign new_B2173_ = ~new_B2172_ & ~new_B2156_;
  assign new_B2174_ = new_B2156_ | new_B2171_;
  assign new_B2175_ = ~new_B2149_ | ~new_B2150_;
  assign new_B2176_ = new_B2156_ | new_B2171_;
  assign new_B2177_ = ~new_B2156_ & ~new_B2178_;
  assign new_B2178_ = new_B2156_ & new_B2171_;
  assign new_B2179_ = new_B6673_;
  assign new_B2180_ = new_B6706_;
  assign new_B2181_ = new_B6739_;
  assign new_B2182_ = new_B6772_;
  assign new_B2183_ = new_B6805_;
  assign new_B2184_ = new_B2190_ & new_B2189_;
  assign new_B2185_ = new_B2192_ | new_B2191_;
  assign new_B2186_ = new_B2194_ | new_B2193_;
  assign new_B2187_ = new_B2189_ & new_B2195_;
  assign new_B2188_ = new_B2189_ & new_B2196_;
  assign new_B2189_ = new_B2179_ ^ new_B2180_;
  assign new_B2190_ = new_B2191_ ^ new_B2181_;
  assign new_B2191_ = new_B2199_ & new_B2198_;
  assign new_B2192_ = new_B2197_ & new_B2181_;
  assign new_B2193_ = new_B2202_ & new_B2201_;
  assign new_B2194_ = new_B2200_ & new_B2181_;
  assign new_B2195_ = new_B2203_ | new_B2180_;
  assign new_B2196_ = ~new_B2181_ ^ new_B2193_;
  assign new_B2197_ = ~new_B2206_ | ~new_B2207_;
  assign new_B2198_ = new_B2182_ ^ new_B2189_;
  assign new_B2199_ = new_B2208_ & new_B2201_;
  assign new_B2200_ = ~new_B2210_ | ~new_B2209_;
  assign new_B2201_ = new_B2182_ | new_B2183_;
  assign new_B2202_ = new_B2182_ | new_B2189_;
  assign new_B2203_ = new_B2181_ & new_B2193_;
  assign new_B2204_ = ~new_B2180_ | ~new_B2181_;
  assign new_B2205_ = new_B2189_ & new_B2204_;
  assign new_B2206_ = ~new_B2205_ & ~new_B2189_;
  assign new_B2207_ = new_B2189_ | new_B2204_;
  assign new_B2208_ = ~new_B2182_ | ~new_B2183_;
  assign new_B2209_ = new_B2189_ | new_B2204_;
  assign new_B2210_ = ~new_B2189_ & ~new_B2211_;
  assign new_B2211_ = new_B2189_ & new_B2204_;
  assign new_B2212_ = new_B6838_;
  assign new_B2213_ = new_B6871_;
  assign new_B2214_ = new_B6904_;
  assign new_B2215_ = new_B6937_;
  assign new_B2216_ = new_B6970_;
  assign new_B2217_ = new_B2223_ & new_B2222_;
  assign new_B2218_ = new_B2225_ | new_B2224_;
  assign new_B2219_ = new_B2227_ | new_B2226_;
  assign new_B2220_ = new_B2222_ & new_B2228_;
  assign new_B2221_ = new_B2222_ & new_B2229_;
  assign new_B2222_ = new_B2212_ ^ new_B2213_;
  assign new_B2223_ = new_B2224_ ^ new_B2214_;
  assign new_B2224_ = new_B2232_ & new_B2231_;
  assign new_B2225_ = new_B2230_ & new_B2214_;
  assign new_B2226_ = new_B2235_ & new_B2234_;
  assign new_B2227_ = new_B2233_ & new_B2214_;
  assign new_B2228_ = new_B2236_ | new_B2213_;
  assign new_B2229_ = ~new_B2214_ ^ new_B2226_;
  assign new_B2230_ = ~new_B2239_ | ~new_B2240_;
  assign new_B2231_ = new_B2215_ ^ new_B2222_;
  assign new_B2232_ = new_B2241_ & new_B2234_;
  assign new_B2233_ = ~new_B2243_ | ~new_B2242_;
  assign new_B2234_ = new_B2215_ | new_B2216_;
  assign new_B2235_ = new_B2215_ | new_B2222_;
  assign new_B2236_ = new_B2214_ & new_B2226_;
  assign new_B2237_ = ~new_B2213_ | ~new_B2214_;
  assign new_B2238_ = new_B2222_ & new_B2237_;
  assign new_B2239_ = ~new_B2238_ & ~new_B2222_;
  assign new_B2240_ = new_B2222_ | new_B2237_;
  assign new_B2241_ = ~new_B2215_ | ~new_B2216_;
  assign new_B2242_ = new_B2222_ | new_B2237_;
  assign new_B2243_ = ~new_B2222_ & ~new_B2244_;
  assign new_B2244_ = new_B2222_ & new_B2237_;
  assign new_B2245_ = new_B7003_;
  assign new_B2246_ = new_B7036_;
  assign new_B2247_ = new_B7069_;
  assign new_B2248_ = new_B7102_;
  assign new_B2249_ = new_B7135_;
  assign new_B2250_ = new_B2256_ & new_B2255_;
  assign new_B2251_ = new_B2258_ | new_B2257_;
  assign new_B2252_ = new_B2260_ | new_B2259_;
  assign new_B2253_ = new_B2255_ & new_B2261_;
  assign new_B2254_ = new_B2255_ & new_B2262_;
  assign new_B2255_ = new_B2245_ ^ new_B2246_;
  assign new_B2256_ = new_B2257_ ^ new_B2247_;
  assign new_B2257_ = new_B2265_ & new_B2264_;
  assign new_B2258_ = new_B2263_ & new_B2247_;
  assign new_B2259_ = new_B2268_ & new_B2267_;
  assign new_B2260_ = new_B2266_ & new_B2247_;
  assign new_B2261_ = new_B2269_ | new_B2246_;
  assign new_B2262_ = ~new_B2247_ ^ new_B2259_;
  assign new_B2263_ = ~new_B2272_ | ~new_B2273_;
  assign new_B2264_ = new_B2248_ ^ new_B2255_;
  assign new_B2265_ = new_B2274_ & new_B2267_;
  assign new_B2266_ = ~new_B2276_ | ~new_B2275_;
  assign new_B2267_ = new_B2248_ | new_B2249_;
  assign new_B2268_ = new_B2248_ | new_B2255_;
  assign new_B2269_ = new_B2247_ & new_B2259_;
  assign new_B2270_ = ~new_B2246_ | ~new_B2247_;
  assign new_B2271_ = new_B2255_ & new_B2270_;
  assign new_B2272_ = ~new_B2271_ & ~new_B2255_;
  assign new_B2273_ = new_B2255_ | new_B2270_;
  assign new_B2274_ = ~new_B2248_ | ~new_B2249_;
  assign new_B2275_ = new_B2255_ | new_B2270_;
  assign new_B2276_ = ~new_B2255_ & ~new_B2277_;
  assign new_B2277_ = new_B2255_ & new_B2270_;
  assign new_B2278_ = new_B7168_;
  assign new_B2279_ = new_B7201_;
  assign new_B2280_ = new_B7234_;
  assign new_B2281_ = new_B7267_;
  assign new_B2282_ = new_B7300_;
  assign new_B2283_ = new_B2289_ & new_B2288_;
  assign new_B2284_ = new_B2291_ | new_B2290_;
  assign new_B2285_ = new_B2293_ | new_B2292_;
  assign new_B2286_ = new_B2288_ & new_B2294_;
  assign new_B2287_ = new_B2288_ & new_B2295_;
  assign new_B2288_ = new_B2278_ ^ new_B2279_;
  assign new_B2289_ = new_B2290_ ^ new_B2280_;
  assign new_B2290_ = new_B2298_ & new_B2297_;
  assign new_B2291_ = new_B2296_ & new_B2280_;
  assign new_B2292_ = new_B2301_ & new_B2300_;
  assign new_B2293_ = new_B2299_ & new_B2280_;
  assign new_B2294_ = new_B2302_ | new_B2279_;
  assign new_B2295_ = ~new_B2280_ ^ new_B2292_;
  assign new_B2296_ = ~new_B2305_ | ~new_B2306_;
  assign new_B2297_ = new_B2281_ ^ new_B2288_;
  assign new_B2298_ = new_B2307_ & new_B2300_;
  assign new_B2299_ = ~new_B2309_ | ~new_B2308_;
  assign new_B2300_ = new_B2281_ | new_B2282_;
  assign new_B2301_ = new_B2281_ | new_B2288_;
  assign new_B2302_ = new_B2280_ & new_B2292_;
  assign new_B2303_ = ~new_B2279_ | ~new_B2280_;
  assign new_B2304_ = new_B2288_ & new_B2303_;
  assign new_B2305_ = ~new_B2304_ & ~new_B2288_;
  assign new_B2306_ = new_B2288_ | new_B2303_;
  assign new_B2307_ = ~new_B2281_ | ~new_B2282_;
  assign new_B2308_ = new_B2288_ | new_B2303_;
  assign new_B2309_ = ~new_B2288_ & ~new_B2310_;
  assign new_B2310_ = new_B2288_ & new_B2303_;
  assign new_B2311_ = new_B7333_;
  assign new_B2312_ = new_B7366_;
  assign new_B2313_ = new_B7399_;
  assign new_B2314_ = new_B7432_;
  assign new_B2315_ = new_B7465_;
  assign new_B2316_ = new_B2322_ & new_B2321_;
  assign new_B2317_ = new_B2324_ | new_B2323_;
  assign new_B2318_ = new_B2326_ | new_B2325_;
  assign new_B2319_ = new_B2321_ & new_B2327_;
  assign new_B2320_ = new_B2321_ & new_B2328_;
  assign new_B2321_ = new_B2311_ ^ new_B2312_;
  assign new_B2322_ = new_B2323_ ^ new_B2313_;
  assign new_B2323_ = new_B2331_ & new_B2330_;
  assign new_B2324_ = new_B2329_ & new_B2313_;
  assign new_B2325_ = new_B2334_ & new_B2333_;
  assign new_B2326_ = new_B2332_ & new_B2313_;
  assign new_B2327_ = new_B2335_ | new_B2312_;
  assign new_B2328_ = ~new_B2313_ ^ new_B2325_;
  assign new_B2329_ = ~new_B2338_ | ~new_B2339_;
  assign new_B2330_ = new_B2314_ ^ new_B2321_;
  assign new_B2331_ = new_B2340_ & new_B2333_;
  assign new_B2332_ = ~new_B2342_ | ~new_B2341_;
  assign new_B2333_ = new_B2314_ | new_B2315_;
  assign new_B2334_ = new_B2314_ | new_B2321_;
  assign new_B2335_ = new_B2313_ & new_B2325_;
  assign new_B2336_ = ~new_B2312_ | ~new_B2313_;
  assign new_B2337_ = new_B2321_ & new_B2336_;
  assign new_B2338_ = ~new_B2337_ & ~new_B2321_;
  assign new_B2339_ = new_B2321_ | new_B2336_;
  assign new_B2340_ = ~new_B2314_ | ~new_B2315_;
  assign new_B2341_ = new_B2321_ | new_B2336_;
  assign new_B2342_ = ~new_B2321_ & ~new_B2343_;
  assign new_B2343_ = new_B2321_ & new_B2336_;
  assign new_B2344_ = new_B7498_;
  assign new_B2345_ = new_B7531_;
  assign new_B2346_ = new_B7564_;
  assign new_B2347_ = new_B7597_;
  assign new_B2348_ = new_B7630_;
  assign new_B2349_ = new_B2355_ & new_B2354_;
  assign new_B2350_ = new_B2357_ | new_B2356_;
  assign new_B2351_ = new_B2359_ | new_B2358_;
  assign new_B2352_ = new_B2354_ & new_B2360_;
  assign new_B2353_ = new_B2354_ & new_B2361_;
  assign new_B2354_ = new_B2344_ ^ new_B2345_;
  assign new_B2355_ = new_B2356_ ^ new_B2346_;
  assign new_B2356_ = new_B2364_ & new_B2363_;
  assign new_B2357_ = new_B2362_ & new_B2346_;
  assign new_B2358_ = new_B2367_ & new_B2366_;
  assign new_B2359_ = new_B2365_ & new_B2346_;
  assign new_B2360_ = new_B2368_ | new_B2345_;
  assign new_B2361_ = ~new_B2346_ ^ new_B2358_;
  assign new_B2362_ = ~new_B2371_ | ~new_B2372_;
  assign new_B2363_ = new_B2347_ ^ new_B2354_;
  assign new_B2364_ = new_B2373_ & new_B2366_;
  assign new_B2365_ = ~new_B2375_ | ~new_B2374_;
  assign new_B2366_ = new_B2347_ | new_B2348_;
  assign new_B2367_ = new_B2347_ | new_B2354_;
  assign new_B2368_ = new_B2346_ & new_B2358_;
  assign new_B2369_ = ~new_B2345_ | ~new_B2346_;
  assign new_B2370_ = new_B2354_ & new_B2369_;
  assign new_B2371_ = ~new_B2370_ & ~new_B2354_;
  assign new_B2372_ = new_B2354_ | new_B2369_;
  assign new_B2373_ = ~new_B2347_ | ~new_B2348_;
  assign new_B2374_ = new_B2354_ | new_B2369_;
  assign new_B2375_ = ~new_B2354_ & ~new_B2376_;
  assign new_B2376_ = new_B2354_ & new_B2369_;
  assign new_B2377_ = new_B7663_;
  assign new_B2378_ = new_B7696_;
  assign new_B2379_ = new_B7729_;
  assign new_B2380_ = new_B7762_;
  assign new_B2381_ = new_B7795_;
  assign new_B2382_ = new_B2388_ & new_B2387_;
  assign new_B2383_ = new_B2390_ | new_B2389_;
  assign new_B2384_ = new_B2392_ | new_B2391_;
  assign new_B2385_ = new_B2387_ & new_B2393_;
  assign new_B2386_ = new_B2387_ & new_B2394_;
  assign new_B2387_ = new_B2377_ ^ new_B2378_;
  assign new_B2388_ = new_B2389_ ^ new_B2379_;
  assign new_B2389_ = new_B2397_ & new_B2396_;
  assign new_B2390_ = new_B2395_ & new_B2379_;
  assign new_B2391_ = new_B2400_ & new_B2399_;
  assign new_B2392_ = new_B2398_ & new_B2379_;
  assign new_B2393_ = new_B2401_ | new_B2378_;
  assign new_B2394_ = ~new_B2379_ ^ new_B2391_;
  assign new_B2395_ = ~new_B2404_ | ~new_B2405_;
  assign new_B2396_ = new_B2380_ ^ new_B2387_;
  assign new_B2397_ = new_B2406_ & new_B2399_;
  assign new_B2398_ = ~new_B2408_ | ~new_B2407_;
  assign new_B2399_ = new_B2380_ | new_B2381_;
  assign new_B2400_ = new_B2380_ | new_B2387_;
  assign new_B2401_ = new_B2379_ & new_B2391_;
  assign new_B2402_ = ~new_B2378_ | ~new_B2379_;
  assign new_B2403_ = new_B2387_ & new_B2402_;
  assign new_B2404_ = ~new_B2403_ & ~new_B2387_;
  assign new_B2405_ = new_B2387_ | new_B2402_;
  assign new_B2406_ = ~new_B2380_ | ~new_B2381_;
  assign new_B2407_ = new_B2387_ | new_B2402_;
  assign new_B2408_ = ~new_B2387_ & ~new_B2409_;
  assign new_B2409_ = new_B2387_ & new_B2402_;
  assign new_B2410_ = new_B7828_;
  assign new_B2411_ = new_B7861_;
  assign new_B2412_ = new_B7894_;
  assign new_B2413_ = new_B7927_;
  assign new_B2414_ = new_B7960_;
  assign new_B2415_ = new_B2421_ & new_B2420_;
  assign new_B2416_ = new_B2423_ | new_B2422_;
  assign new_B2417_ = new_B2425_ | new_B2424_;
  assign new_B2418_ = new_B2420_ & new_B2426_;
  assign new_B2419_ = new_B2420_ & new_B2427_;
  assign new_B2420_ = new_B2410_ ^ new_B2411_;
  assign new_B2421_ = new_B2422_ ^ new_B2412_;
  assign new_B2422_ = new_B2430_ & new_B2429_;
  assign new_B2423_ = new_B2428_ & new_B2412_;
  assign new_B2424_ = new_B2433_ & new_B2432_;
  assign new_B2425_ = new_B2431_ & new_B2412_;
  assign new_B2426_ = new_B2434_ | new_B2411_;
  assign new_B2427_ = ~new_B2412_ ^ new_B2424_;
  assign new_B2428_ = ~new_B2437_ | ~new_B2438_;
  assign new_B2429_ = new_B2413_ ^ new_B2420_;
  assign new_B2430_ = new_B2439_ & new_B2432_;
  assign new_B2431_ = ~new_B2441_ | ~new_B2440_;
  assign new_B2432_ = new_B2413_ | new_B2414_;
  assign new_B2433_ = new_B2413_ | new_B2420_;
  assign new_B2434_ = new_B2412_ & new_B2424_;
  assign new_B2435_ = ~new_B2411_ | ~new_B2412_;
  assign new_B2436_ = new_B2420_ & new_B2435_;
  assign new_B2437_ = ~new_B2436_ & ~new_B2420_;
  assign new_B2438_ = new_B2420_ | new_B2435_;
  assign new_B2439_ = ~new_B2413_ | ~new_B2414_;
  assign new_B2440_ = new_B2420_ | new_B2435_;
  assign new_B2441_ = ~new_B2420_ & ~new_B2442_;
  assign new_B2442_ = new_B2420_ & new_B2435_;
  assign new_B2443_ = new_B7993_;
  assign new_B2444_ = new_B8026_;
  assign new_B2445_ = new_B8059_;
  assign new_B2446_ = new_B8092_;
  assign new_B2447_ = new_B8125_;
  assign new_B2448_ = new_B2454_ & new_B2453_;
  assign new_B2449_ = new_B2456_ | new_B2455_;
  assign new_B2450_ = new_B2458_ | new_B2457_;
  assign new_B2451_ = new_B2453_ & new_B2459_;
  assign new_B2452_ = new_B2453_ & new_B2460_;
  assign new_B2453_ = new_B2443_ ^ new_B2444_;
  assign new_B2454_ = new_B2455_ ^ new_B2445_;
  assign new_B2455_ = new_B2463_ & new_B2462_;
  assign new_B2456_ = new_B2461_ & new_B2445_;
  assign new_B2457_ = new_B2466_ & new_B2465_;
  assign new_B2458_ = new_B2464_ & new_B2445_;
  assign new_B2459_ = new_B2467_ | new_B2444_;
  assign new_B2460_ = ~new_B2445_ ^ new_B2457_;
  assign new_B2461_ = ~new_B2470_ | ~new_B2471_;
  assign new_B2462_ = new_B2446_ ^ new_B2453_;
  assign new_B2463_ = new_B2472_ & new_B2465_;
  assign new_B2464_ = ~new_B2474_ | ~new_B2473_;
  assign new_B2465_ = new_B2446_ | new_B2447_;
  assign new_B2466_ = new_B2446_ | new_B2453_;
  assign new_B2467_ = new_B2445_ & new_B2457_;
  assign new_B2468_ = ~new_B2444_ | ~new_B2445_;
  assign new_B2469_ = new_B2453_ & new_B2468_;
  assign new_B2470_ = ~new_B2469_ & ~new_B2453_;
  assign new_B2471_ = new_B2453_ | new_B2468_;
  assign new_B2472_ = ~new_B2446_ | ~new_B2447_;
  assign new_B2473_ = new_B2453_ | new_B2468_;
  assign new_B2474_ = ~new_B2453_ & ~new_B2475_;
  assign new_B2475_ = new_B2453_ & new_B2468_;
  assign new_B2476_ = new_B8158_;
  assign new_B2477_ = new_B8191_;
  assign new_B2478_ = new_B8224_;
  assign new_B2479_ = new_B8257_;
  assign new_B2480_ = new_B8290_;
  assign new_B2481_ = new_B2487_ & new_B2486_;
  assign new_B2482_ = new_B2489_ | new_B2488_;
  assign new_B2483_ = new_B2491_ | new_B2490_;
  assign new_B2484_ = new_B2486_ & new_B2492_;
  assign new_B2485_ = new_B2486_ & new_B2493_;
  assign new_B2486_ = new_B2476_ ^ new_B2477_;
  assign new_B2487_ = new_B2488_ ^ new_B2478_;
  assign new_B2488_ = new_B2496_ & new_B2495_;
  assign new_B2489_ = new_B2494_ & new_B2478_;
  assign new_B2490_ = new_B2499_ & new_B2498_;
  assign new_B2491_ = new_B2497_ & new_B2478_;
  assign new_B2492_ = new_B2500_ | new_B2477_;
  assign new_B2493_ = ~new_B2478_ ^ new_B2490_;
  assign new_B2494_ = ~new_B2503_ | ~new_B2504_;
  assign new_B2495_ = new_B2479_ ^ new_B2486_;
  assign new_B2496_ = new_B2505_ & new_B2498_;
  assign new_B2497_ = ~new_B2507_ | ~new_B2506_;
  assign new_B2498_ = new_B2479_ | new_B2480_;
  assign new_B2499_ = new_B2479_ | new_B2486_;
  assign new_B2500_ = new_B2478_ & new_B2490_;
  assign new_B2501_ = ~new_B2477_ | ~new_B2478_;
  assign new_B2502_ = new_B2486_ & new_B2501_;
  assign new_B2503_ = ~new_B2502_ & ~new_B2486_;
  assign new_B2504_ = new_B2486_ | new_B2501_;
  assign new_B2505_ = ~new_B2479_ | ~new_B2480_;
  assign new_B2506_ = new_B2486_ | new_B2501_;
  assign new_B2507_ = ~new_B2486_ & ~new_B2508_;
  assign new_B2508_ = new_B2486_ & new_B2501_;
  assign new_B2509_ = new_B8323_;
  assign new_B2510_ = new_B8356_;
  assign new_B2511_ = new_B8389_;
  assign new_B2512_ = new_B8422_;
  assign new_B2513_ = new_B8455_;
  assign new_B2514_ = new_B2520_ & new_B2519_;
  assign new_B2515_ = new_B2522_ | new_B2521_;
  assign new_B2516_ = new_B2524_ | new_B2523_;
  assign new_B2517_ = new_B2519_ & new_B2525_;
  assign new_B2518_ = new_B2519_ & new_B2526_;
  assign new_B2519_ = new_B2509_ ^ new_B2510_;
  assign new_B2520_ = new_B2521_ ^ new_B2511_;
  assign new_B2521_ = new_B2529_ & new_B2528_;
  assign new_B2522_ = new_B2527_ & new_B2511_;
  assign new_B2523_ = new_B2532_ & new_B2531_;
  assign new_B2524_ = new_B2530_ & new_B2511_;
  assign new_B2525_ = new_B2533_ | new_B2510_;
  assign new_B2526_ = ~new_B2511_ ^ new_B2523_;
  assign new_B2527_ = ~new_B2536_ | ~new_B2537_;
  assign new_B2528_ = new_B2512_ ^ new_B2519_;
  assign new_B2529_ = new_B2538_ & new_B2531_;
  assign new_B2530_ = ~new_B2540_ | ~new_B2539_;
  assign new_B2531_ = new_B2512_ | new_B2513_;
  assign new_B2532_ = new_B2512_ | new_B2519_;
  assign new_B2533_ = new_B2511_ & new_B2523_;
  assign new_B2534_ = ~new_B2510_ | ~new_B2511_;
  assign new_B2535_ = new_B2519_ & new_B2534_;
  assign new_B2536_ = ~new_B2535_ & ~new_B2519_;
  assign new_B2537_ = new_B2519_ | new_B2534_;
  assign new_B2538_ = ~new_B2512_ | ~new_B2513_;
  assign new_B2539_ = new_B2519_ | new_B2534_;
  assign new_B2540_ = ~new_B2519_ & ~new_B2541_;
  assign new_B2541_ = new_B2519_ & new_B2534_;
  assign new_B2542_ = new_B8488_;
  assign new_B2543_ = new_B8521_;
  assign new_B2544_ = new_B8554_;
  assign new_B2545_ = new_B8587_;
  assign new_B2546_ = new_B8620_;
  assign new_B2547_ = new_B2553_ & new_B2552_;
  assign new_B2548_ = new_B2555_ | new_B2554_;
  assign new_B2549_ = new_B2557_ | new_B2556_;
  assign new_B2550_ = new_B2552_ & new_B2558_;
  assign new_B2551_ = new_B2552_ & new_B2559_;
  assign new_B2552_ = new_B2542_ ^ new_B2543_;
  assign new_B2553_ = new_B2554_ ^ new_B2544_;
  assign new_B2554_ = new_B2562_ & new_B2561_;
  assign new_B2555_ = new_B2560_ & new_B2544_;
  assign new_B2556_ = new_B2565_ & new_B2564_;
  assign new_B2557_ = new_B2563_ & new_B2544_;
  assign new_B2558_ = new_B2566_ | new_B2543_;
  assign new_B2559_ = ~new_B2544_ ^ new_B2556_;
  assign new_B2560_ = ~new_B2569_ | ~new_B2570_;
  assign new_B2561_ = new_B2545_ ^ new_B2552_;
  assign new_B2562_ = new_B2571_ & new_B2564_;
  assign new_B2563_ = ~new_B2573_ | ~new_B2572_;
  assign new_B2564_ = new_B2545_ | new_B2546_;
  assign new_B2565_ = new_B2545_ | new_B2552_;
  assign new_B2566_ = new_B2544_ & new_B2556_;
  assign new_B2567_ = ~new_B2543_ | ~new_B2544_;
  assign new_B2568_ = new_B2552_ & new_B2567_;
  assign new_B2569_ = ~new_B2568_ & ~new_B2552_;
  assign new_B2570_ = new_B2552_ | new_B2567_;
  assign new_B2571_ = ~new_B2545_ | ~new_B2546_;
  assign new_B2572_ = new_B2552_ | new_B2567_;
  assign new_B2573_ = ~new_B2552_ & ~new_B2574_;
  assign new_B2574_ = new_B2552_ & new_B2567_;
  assign new_B2575_ = new_B8653_;
  assign new_B2576_ = new_B8686_;
  assign new_B2577_ = new_B8719_;
  assign new_B2578_ = new_B8752_;
  assign new_B2579_ = new_B8785_;
  assign new_B2580_ = new_B2586_ & new_B2585_;
  assign new_B2581_ = new_B2588_ | new_B2587_;
  assign new_B2582_ = new_B2590_ | new_B2589_;
  assign new_B2583_ = new_B2585_ & new_B2591_;
  assign new_B2584_ = new_B2585_ & new_B2592_;
  assign new_B2585_ = new_B2575_ ^ new_B2576_;
  assign new_B2586_ = new_B2587_ ^ new_B2577_;
  assign new_B2587_ = new_B2595_ & new_B2594_;
  assign new_B2588_ = new_B2593_ & new_B2577_;
  assign new_B2589_ = new_B2598_ & new_B2597_;
  assign new_B2590_ = new_B2596_ & new_B2577_;
  assign new_B2591_ = new_B2599_ | new_B2576_;
  assign new_B2592_ = ~new_B2577_ ^ new_B2589_;
  assign new_B2593_ = ~new_B2602_ | ~new_B2603_;
  assign new_B2594_ = new_B2578_ ^ new_B2585_;
  assign new_B2595_ = new_B2604_ & new_B2597_;
  assign new_B2596_ = ~new_B2606_ | ~new_B2605_;
  assign new_B2597_ = new_B2578_ | new_B2579_;
  assign new_B2598_ = new_B2578_ | new_B2585_;
  assign new_B2599_ = new_B2577_ & new_B2589_;
  assign new_B2600_ = ~new_B2576_ | ~new_B2577_;
  assign new_B2601_ = new_B2585_ & new_B2600_;
  assign new_B2602_ = ~new_B2601_ & ~new_B2585_;
  assign new_B2603_ = new_B2585_ | new_B2600_;
  assign new_B2604_ = ~new_B2578_ | ~new_B2579_;
  assign new_B2605_ = new_B2585_ | new_B2600_;
  assign new_B2606_ = ~new_B2585_ & ~new_B2607_;
  assign new_B2607_ = new_B2585_ & new_B2600_;
  assign new_B2608_ = new_B8818_;
  assign new_B2609_ = new_B8851_;
  assign new_B2610_ = new_B8884_;
  assign new_B2611_ = new_B8917_;
  assign new_B2612_ = new_B8950_;
  assign new_B2613_ = new_B2619_ & new_B2618_;
  assign new_B2614_ = new_B2621_ | new_B2620_;
  assign new_B2615_ = new_B2623_ | new_B2622_;
  assign new_B2616_ = new_B2618_ & new_B2624_;
  assign new_B2617_ = new_B2618_ & new_B2625_;
  assign new_B2618_ = new_B2608_ ^ new_B2609_;
  assign new_B2619_ = new_B2620_ ^ new_B2610_;
  assign new_B2620_ = new_B2628_ & new_B2627_;
  assign new_B2621_ = new_B2626_ & new_B2610_;
  assign new_B2622_ = new_B2631_ & new_B2630_;
  assign new_B2623_ = new_B2629_ & new_B2610_;
  assign new_B2624_ = new_B2632_ | new_B2609_;
  assign new_B2625_ = ~new_B2610_ ^ new_B2622_;
  assign new_B2626_ = ~new_B2635_ | ~new_B2636_;
  assign new_B2627_ = new_B2611_ ^ new_B2618_;
  assign new_B2628_ = new_B2637_ & new_B2630_;
  assign new_B2629_ = ~new_B2639_ | ~new_B2638_;
  assign new_B2630_ = new_B2611_ | new_B2612_;
  assign new_B2631_ = new_B2611_ | new_B2618_;
  assign new_B2632_ = new_B2610_ & new_B2622_;
  assign new_B2633_ = ~new_B2609_ | ~new_B2610_;
  assign new_B2634_ = new_B2618_ & new_B2633_;
  assign new_B2635_ = ~new_B2634_ & ~new_B2618_;
  assign new_B2636_ = new_B2618_ | new_B2633_;
  assign new_B2637_ = ~new_B2611_ | ~new_B2612_;
  assign new_B2638_ = new_B2618_ | new_B2633_;
  assign new_B2639_ = ~new_B2618_ & ~new_B2640_;
  assign new_B2640_ = new_B2618_ & new_B2633_;
  assign new_B2641_ = new_B8983_;
  assign new_B2642_ = new_B9016_;
  assign new_B2643_ = new_B9049_;
  assign new_B2644_ = new_B9082_;
  assign new_B2645_ = new_B9115_;
  assign new_B2646_ = new_B2652_ & new_B2651_;
  assign new_B2647_ = new_B2654_ | new_B2653_;
  assign new_B2648_ = new_B2656_ | new_B2655_;
  assign new_B2649_ = new_B2651_ & new_B2657_;
  assign new_B2650_ = new_B2651_ & new_B2658_;
  assign new_B2651_ = new_B2641_ ^ new_B2642_;
  assign new_B2652_ = new_B2653_ ^ new_B2643_;
  assign new_B2653_ = new_B2661_ & new_B2660_;
  assign new_B2654_ = new_B2659_ & new_B2643_;
  assign new_B2655_ = new_B2664_ & new_B2663_;
  assign new_B2656_ = new_B2662_ & new_B2643_;
  assign new_B2657_ = new_B2665_ | new_B2642_;
  assign new_B2658_ = ~new_B2643_ ^ new_B2655_;
  assign new_B2659_ = ~new_B2668_ | ~new_B2669_;
  assign new_B2660_ = new_B2644_ ^ new_B2651_;
  assign new_B2661_ = new_B2670_ & new_B2663_;
  assign new_B2662_ = ~new_B2672_ | ~new_B2671_;
  assign new_B2663_ = new_B2644_ | new_B2645_;
  assign new_B2664_ = new_B2644_ | new_B2651_;
  assign new_B2665_ = new_B2643_ & new_B2655_;
  assign new_B2666_ = ~new_B2642_ | ~new_B2643_;
  assign new_B2667_ = new_B2651_ & new_B2666_;
  assign new_B2668_ = ~new_B2667_ & ~new_B2651_;
  assign new_B2669_ = new_B2651_ | new_B2666_;
  assign new_B2670_ = ~new_B2644_ | ~new_B2645_;
  assign new_B2671_ = new_B2651_ | new_B2666_;
  assign new_B2672_ = ~new_B2651_ & ~new_B2673_;
  assign new_B2673_ = new_B2651_ & new_B2666_;
  assign new_B2674_ = new_B9148_;
  assign new_B2675_ = new_B9181_;
  assign new_B2676_ = new_B9214_;
  assign new_B2677_ = new_B9247_;
  assign new_B2678_ = new_B9280_;
  assign new_B2679_ = new_B2685_ & new_B2684_;
  assign new_B2680_ = new_B2687_ | new_B2686_;
  assign new_B2681_ = new_B2689_ | new_B2688_;
  assign new_B2682_ = new_B2684_ & new_B2690_;
  assign new_B2683_ = new_B2684_ & new_B2691_;
  assign new_B2684_ = new_B2674_ ^ new_B2675_;
  assign new_B2685_ = new_B2686_ ^ new_B2676_;
  assign new_B2686_ = new_B2694_ & new_B2693_;
  assign new_B2687_ = new_B2692_ & new_B2676_;
  assign new_B2688_ = new_B2697_ & new_B2696_;
  assign new_B2689_ = new_B2695_ & new_B2676_;
  assign new_B2690_ = new_B2698_ | new_B2675_;
  assign new_B2691_ = ~new_B2676_ ^ new_B2688_;
  assign new_B2692_ = ~new_B2701_ | ~new_B2702_;
  assign new_B2693_ = new_B2677_ ^ new_B2684_;
  assign new_B2694_ = new_B2703_ & new_B2696_;
  assign new_B2695_ = ~new_B2705_ | ~new_B2704_;
  assign new_B2696_ = new_B2677_ | new_B2678_;
  assign new_B2697_ = new_B2677_ | new_B2684_;
  assign new_B2698_ = new_B2676_ & new_B2688_;
  assign new_B2699_ = ~new_B2675_ | ~new_B2676_;
  assign new_B2700_ = new_B2684_ & new_B2699_;
  assign new_B2701_ = ~new_B2700_ & ~new_B2684_;
  assign new_B2702_ = new_B2684_ | new_B2699_;
  assign new_B2703_ = ~new_B2677_ | ~new_B2678_;
  assign new_B2704_ = new_B2684_ | new_B2699_;
  assign new_B2705_ = ~new_B2684_ & ~new_B2706_;
  assign new_B2706_ = new_B2684_ & new_B2699_;
  assign new_B2707_ = new_B5189_;
  assign new_B2708_ = new_B5222_;
  assign new_B2709_ = new_B5255_;
  assign new_B2710_ = new_B5288_;
  assign new_B2711_ = new_B5321_;
  assign new_B2712_ = new_B2718_ & new_B2717_;
  assign new_B2713_ = new_B2720_ | new_B2719_;
  assign new_B2714_ = new_B2722_ | new_B2721_;
  assign new_B2715_ = new_B2717_ & new_B2723_;
  assign new_B2716_ = new_B2717_ & new_B2724_;
  assign new_B2717_ = new_B2707_ ^ new_B2708_;
  assign new_B2718_ = new_B2719_ ^ new_B2709_;
  assign new_B2719_ = new_B2727_ & new_B2726_;
  assign new_B2720_ = new_B2725_ & new_B2709_;
  assign new_B2721_ = new_B2730_ & new_B2729_;
  assign new_B2722_ = new_B2728_ & new_B2709_;
  assign new_B2723_ = new_B2731_ | new_B2708_;
  assign new_B2724_ = ~new_B2709_ ^ new_B2721_;
  assign new_B2725_ = ~new_B2734_ | ~new_B2735_;
  assign new_B2726_ = new_B2710_ ^ new_B2717_;
  assign new_B2727_ = new_B2736_ & new_B2729_;
  assign new_B2728_ = ~new_B2738_ | ~new_B2737_;
  assign new_B2729_ = new_B2710_ | new_B2711_;
  assign new_B2730_ = new_B2710_ | new_B2717_;
  assign new_B2731_ = new_B2709_ & new_B2721_;
  assign new_B2732_ = ~new_B2708_ | ~new_B2709_;
  assign new_B2733_ = new_B2717_ & new_B2732_;
  assign new_B2734_ = ~new_B2733_ & ~new_B2717_;
  assign new_B2735_ = new_B2717_ | new_B2732_;
  assign new_B2736_ = ~new_B2710_ | ~new_B2711_;
  assign new_B2737_ = new_B2717_ | new_B2732_;
  assign new_B2738_ = ~new_B2717_ & ~new_B2739_;
  assign new_B2739_ = new_B2717_ & new_B2732_;
  assign new_B2740_ = new_B5354_;
  assign new_B2741_ = new_B5387_;
  assign new_B2742_ = new_B5420_;
  assign new_B2743_ = new_B5453_;
  assign new_B2744_ = new_B5486_;
  assign new_B2745_ = new_B2751_ & new_B2750_;
  assign new_B2746_ = new_B2753_ | new_B2752_;
  assign new_B2747_ = new_B2755_ | new_B2754_;
  assign new_B2748_ = new_B2750_ & new_B2756_;
  assign new_B2749_ = new_B2750_ & new_B2757_;
  assign new_B2750_ = new_B2740_ ^ new_B2741_;
  assign new_B2751_ = new_B2752_ ^ new_B2742_;
  assign new_B2752_ = new_B2760_ & new_B2759_;
  assign new_B2753_ = new_B2758_ & new_B2742_;
  assign new_B2754_ = new_B2763_ & new_B2762_;
  assign new_B2755_ = new_B2761_ & new_B2742_;
  assign new_B2756_ = new_B2764_ | new_B2741_;
  assign new_B2757_ = ~new_B2742_ ^ new_B2754_;
  assign new_B2758_ = ~new_B2767_ | ~new_B2768_;
  assign new_B2759_ = new_B2743_ ^ new_B2750_;
  assign new_B2760_ = new_B2769_ & new_B2762_;
  assign new_B2761_ = ~new_B2771_ | ~new_B2770_;
  assign new_B2762_ = new_B2743_ | new_B2744_;
  assign new_B2763_ = new_B2743_ | new_B2750_;
  assign new_B2764_ = new_B2742_ & new_B2754_;
  assign new_B2765_ = ~new_B2741_ | ~new_B2742_;
  assign new_B2766_ = new_B2750_ & new_B2765_;
  assign new_B2767_ = ~new_B2766_ & ~new_B2750_;
  assign new_B2768_ = new_B2750_ | new_B2765_;
  assign new_B2769_ = ~new_B2743_ | ~new_B2744_;
  assign new_B2770_ = new_B2750_ | new_B2765_;
  assign new_B2771_ = ~new_B2750_ & ~new_B2772_;
  assign new_B2772_ = new_B2750_ & new_B2765_;
  assign new_B2773_ = new_B5519_;
  assign new_B2774_ = new_B5552_;
  assign new_B2775_ = new_B5585_;
  assign new_B2776_ = new_B5618_;
  assign new_B2777_ = new_B5651_;
  assign new_B2778_ = new_B2784_ & new_B2783_;
  assign new_B2779_ = new_B2786_ | new_B2785_;
  assign new_B2780_ = new_B2788_ | new_B2787_;
  assign new_B2781_ = new_B2783_ & new_B2789_;
  assign new_B2782_ = new_B2783_ & new_B2790_;
  assign new_B2783_ = new_B2773_ ^ new_B2774_;
  assign new_B2784_ = new_B2785_ ^ new_B2775_;
  assign new_B2785_ = new_B2793_ & new_B2792_;
  assign new_B2786_ = new_B2791_ & new_B2775_;
  assign new_B2787_ = new_B2796_ & new_B2795_;
  assign new_B2788_ = new_B2794_ & new_B2775_;
  assign new_B2789_ = new_B2797_ | new_B2774_;
  assign new_B2790_ = ~new_B2775_ ^ new_B2787_;
  assign new_B2791_ = ~new_B2800_ | ~new_B2801_;
  assign new_B2792_ = new_B2776_ ^ new_B2783_;
  assign new_B2793_ = new_B2802_ & new_B2795_;
  assign new_B2794_ = ~new_B2804_ | ~new_B2803_;
  assign new_B2795_ = new_B2776_ | new_B2777_;
  assign new_B2796_ = new_B2776_ | new_B2783_;
  assign new_B2797_ = new_B2775_ & new_B2787_;
  assign new_B2798_ = ~new_B2774_ | ~new_B2775_;
  assign new_B2799_ = new_B2783_ & new_B2798_;
  assign new_B2800_ = ~new_B2799_ & ~new_B2783_;
  assign new_B2801_ = new_B2783_ | new_B2798_;
  assign new_B2802_ = ~new_B2776_ | ~new_B2777_;
  assign new_B2803_ = new_B2783_ | new_B2798_;
  assign new_B2804_ = ~new_B2783_ & ~new_B2805_;
  assign new_B2805_ = new_B2783_ & new_B2798_;
  assign new_B2806_ = new_B5684_;
  assign new_B2807_ = new_B5717_;
  assign new_B2808_ = new_B5750_;
  assign new_B2809_ = new_B5783_;
  assign new_B2810_ = new_B5816_;
  assign new_B2811_ = new_B2817_ & new_B2816_;
  assign new_B2812_ = new_B2819_ | new_B2818_;
  assign new_B2813_ = new_B2821_ | new_B2820_;
  assign new_B2814_ = new_B2816_ & new_B2822_;
  assign new_B2815_ = new_B2816_ & new_B2823_;
  assign new_B2816_ = new_B2806_ ^ new_B2807_;
  assign new_B2817_ = new_B2818_ ^ new_B2808_;
  assign new_B2818_ = new_B2826_ & new_B2825_;
  assign new_B2819_ = new_B2824_ & new_B2808_;
  assign new_B2820_ = new_B2829_ & new_B2828_;
  assign new_B2821_ = new_B2827_ & new_B2808_;
  assign new_B2822_ = new_B2830_ | new_B2807_;
  assign new_B2823_ = ~new_B2808_ ^ new_B2820_;
  assign new_B2824_ = ~new_B2833_ | ~new_B2834_;
  assign new_B2825_ = new_B2809_ ^ new_B2816_;
  assign new_B2826_ = new_B2835_ & new_B2828_;
  assign new_B2827_ = ~new_B2837_ | ~new_B2836_;
  assign new_B2828_ = new_B2809_ | new_B2810_;
  assign new_B2829_ = new_B2809_ | new_B2816_;
  assign new_B2830_ = new_B2808_ & new_B2820_;
  assign new_B2831_ = ~new_B2807_ | ~new_B2808_;
  assign new_B2832_ = new_B2816_ & new_B2831_;
  assign new_B2833_ = ~new_B2832_ & ~new_B2816_;
  assign new_B2834_ = new_B2816_ | new_B2831_;
  assign new_B2835_ = ~new_B2809_ | ~new_B2810_;
  assign new_B2836_ = new_B2816_ | new_B2831_;
  assign new_B2837_ = ~new_B2816_ & ~new_B2838_;
  assign new_B2838_ = new_B2816_ & new_B2831_;
  assign new_B2839_ = new_B5849_;
  assign new_B2840_ = new_B5882_;
  assign new_B2841_ = new_B5915_;
  assign new_B2842_ = new_B5948_;
  assign new_B2843_ = new_B5981_;
  assign new_B2844_ = new_B2850_ & new_B2849_;
  assign new_B2845_ = new_B2852_ | new_B2851_;
  assign new_B2846_ = new_B2854_ | new_B2853_;
  assign new_B2847_ = new_B2849_ & new_B2855_;
  assign new_B2848_ = new_B2849_ & new_B2856_;
  assign new_B2849_ = new_B2839_ ^ new_B2840_;
  assign new_B2850_ = new_B2851_ ^ new_B2841_;
  assign new_B2851_ = new_B2859_ & new_B2858_;
  assign new_B2852_ = new_B2857_ & new_B2841_;
  assign new_B2853_ = new_B2862_ & new_B2861_;
  assign new_B2854_ = new_B2860_ & new_B2841_;
  assign new_B2855_ = new_B2863_ | new_B2840_;
  assign new_B2856_ = ~new_B2841_ ^ new_B2853_;
  assign new_B2857_ = ~new_B2866_ | ~new_B2867_;
  assign new_B2858_ = new_B2842_ ^ new_B2849_;
  assign new_B2859_ = new_B2868_ & new_B2861_;
  assign new_B2860_ = ~new_B2870_ | ~new_B2869_;
  assign new_B2861_ = new_B2842_ | new_B2843_;
  assign new_B2862_ = new_B2842_ | new_B2849_;
  assign new_B2863_ = new_B2841_ & new_B2853_;
  assign new_B2864_ = ~new_B2840_ | ~new_B2841_;
  assign new_B2865_ = new_B2849_ & new_B2864_;
  assign new_B2866_ = ~new_B2865_ & ~new_B2849_;
  assign new_B2867_ = new_B2849_ | new_B2864_;
  assign new_B2868_ = ~new_B2842_ | ~new_B2843_;
  assign new_B2869_ = new_B2849_ | new_B2864_;
  assign new_B2870_ = ~new_B2849_ & ~new_B2871_;
  assign new_B2871_ = new_B2849_ & new_B2864_;
  assign new_B2872_ = new_B6014_;
  assign new_B2873_ = new_B6047_;
  assign new_B2874_ = new_B6080_;
  assign new_B2875_ = new_B6113_;
  assign new_B2876_ = new_B6146_;
  assign new_B2877_ = new_B2883_ & new_B2882_;
  assign new_B2878_ = new_B2885_ | new_B2884_;
  assign new_B2879_ = new_B2887_ | new_B2886_;
  assign new_B2880_ = new_B2882_ & new_B2888_;
  assign new_B2881_ = new_B2882_ & new_B2889_;
  assign new_B2882_ = new_B2872_ ^ new_B2873_;
  assign new_B2883_ = new_B2884_ ^ new_B2874_;
  assign new_B2884_ = new_B2892_ & new_B2891_;
  assign new_B2885_ = new_B2890_ & new_B2874_;
  assign new_B2886_ = new_B2895_ & new_B2894_;
  assign new_B2887_ = new_B2893_ & new_B2874_;
  assign new_B2888_ = new_B2896_ | new_B2873_;
  assign new_B2889_ = ~new_B2874_ ^ new_B2886_;
  assign new_B2890_ = ~new_B2899_ | ~new_B2900_;
  assign new_B2891_ = new_B2875_ ^ new_B2882_;
  assign new_B2892_ = new_B2901_ & new_B2894_;
  assign new_B2893_ = ~new_B2903_ | ~new_B2902_;
  assign new_B2894_ = new_B2875_ | new_B2876_;
  assign new_B2895_ = new_B2875_ | new_B2882_;
  assign new_B2896_ = new_B2874_ & new_B2886_;
  assign new_B2897_ = ~new_B2873_ | ~new_B2874_;
  assign new_B2898_ = new_B2882_ & new_B2897_;
  assign new_B2899_ = ~new_B2898_ & ~new_B2882_;
  assign new_B2900_ = new_B2882_ | new_B2897_;
  assign new_B2901_ = ~new_B2875_ | ~new_B2876_;
  assign new_B2902_ = new_B2882_ | new_B2897_;
  assign new_B2903_ = ~new_B2882_ & ~new_B2904_;
  assign new_B2904_ = new_B2882_ & new_B2897_;
  assign new_B2905_ = new_B6179_;
  assign new_B2906_ = new_B6212_;
  assign new_B2907_ = new_B6245_;
  assign new_B2908_ = new_B6278_;
  assign new_B2909_ = new_B6311_;
  assign new_B2910_ = new_B2916_ & new_B2915_;
  assign new_B2911_ = new_B2918_ | new_B2917_;
  assign new_B2912_ = new_B2920_ | new_B2919_;
  assign new_B2913_ = new_B2915_ & new_B2921_;
  assign new_B2914_ = new_B2915_ & new_B2922_;
  assign new_B2915_ = new_B2905_ ^ new_B2906_;
  assign new_B2916_ = new_B2917_ ^ new_B2907_;
  assign new_B2917_ = new_B2925_ & new_B2924_;
  assign new_B2918_ = new_B2923_ & new_B2907_;
  assign new_B2919_ = new_B2928_ & new_B2927_;
  assign new_B2920_ = new_B2926_ & new_B2907_;
  assign new_B2921_ = new_B2929_ | new_B2906_;
  assign new_B2922_ = ~new_B2907_ ^ new_B2919_;
  assign new_B2923_ = ~new_B2932_ | ~new_B2933_;
  assign new_B2924_ = new_B2908_ ^ new_B2915_;
  assign new_B2925_ = new_B2934_ & new_B2927_;
  assign new_B2926_ = ~new_B2936_ | ~new_B2935_;
  assign new_B2927_ = new_B2908_ | new_B2909_;
  assign new_B2928_ = new_B2908_ | new_B2915_;
  assign new_B2929_ = new_B2907_ & new_B2919_;
  assign new_B2930_ = ~new_B2906_ | ~new_B2907_;
  assign new_B2931_ = new_B2915_ & new_B2930_;
  assign new_B2932_ = ~new_B2931_ & ~new_B2915_;
  assign new_B2933_ = new_B2915_ | new_B2930_;
  assign new_B2934_ = ~new_B2908_ | ~new_B2909_;
  assign new_B2935_ = new_B2915_ | new_B2930_;
  assign new_B2936_ = ~new_B2915_ & ~new_B2937_;
  assign new_B2937_ = new_B2915_ & new_B2930_;
  assign new_B2938_ = new_B6344_;
  assign new_B2939_ = new_B6377_;
  assign new_B2940_ = new_B6410_;
  assign new_B2941_ = new_B6443_;
  assign new_B2942_ = new_B6476_;
  assign new_B2943_ = new_B2949_ & new_B2948_;
  assign new_B2944_ = new_B2951_ | new_B2950_;
  assign new_B2945_ = new_B2953_ | new_B2952_;
  assign new_B2946_ = new_B2948_ & new_B2954_;
  assign new_B2947_ = new_B2948_ & new_B2955_;
  assign new_B2948_ = new_B2938_ ^ new_B2939_;
  assign new_B2949_ = new_B2950_ ^ new_B2940_;
  assign new_B2950_ = new_B2958_ & new_B2957_;
  assign new_B2951_ = new_B2956_ & new_B2940_;
  assign new_B2952_ = new_B2961_ & new_B2960_;
  assign new_B2953_ = new_B2959_ & new_B2940_;
  assign new_B2954_ = new_B2962_ | new_B2939_;
  assign new_B2955_ = ~new_B2940_ ^ new_B2952_;
  assign new_B2956_ = ~new_B2965_ | ~new_B2966_;
  assign new_B2957_ = new_B2941_ ^ new_B2948_;
  assign new_B2958_ = new_B2967_ & new_B2960_;
  assign new_B2959_ = ~new_B2969_ | ~new_B2968_;
  assign new_B2960_ = new_B2941_ | new_B2942_;
  assign new_B2961_ = new_B2941_ | new_B2948_;
  assign new_B2962_ = new_B2940_ & new_B2952_;
  assign new_B2963_ = ~new_B2939_ | ~new_B2940_;
  assign new_B2964_ = new_B2948_ & new_B2963_;
  assign new_B2965_ = ~new_B2964_ & ~new_B2948_;
  assign new_B2966_ = new_B2948_ | new_B2963_;
  assign new_B2967_ = ~new_B2941_ | ~new_B2942_;
  assign new_B2968_ = new_B2948_ | new_B2963_;
  assign new_B2969_ = ~new_B2948_ & ~new_B2970_;
  assign new_B2970_ = new_B2948_ & new_B2963_;
  assign new_B2971_ = new_B6509_;
  assign new_B2972_ = new_B6542_;
  assign new_B2973_ = new_B6575_;
  assign new_B2974_ = new_B6608_;
  assign new_B2975_ = new_B6641_;
  assign new_B2976_ = new_B2982_ & new_B2981_;
  assign new_B2977_ = new_B2984_ | new_B2983_;
  assign new_B2978_ = new_B2986_ | new_B2985_;
  assign new_B2979_ = new_B2981_ & new_B2987_;
  assign new_B2980_ = new_B2981_ & new_B2988_;
  assign new_B2981_ = new_B2971_ ^ new_B2972_;
  assign new_B2982_ = new_B2983_ ^ new_B2973_;
  assign new_B2983_ = new_B2991_ & new_B2990_;
  assign new_B2984_ = new_B2989_ & new_B2973_;
  assign new_B2985_ = new_B2994_ & new_B2993_;
  assign new_B2986_ = new_B2992_ & new_B2973_;
  assign new_B2987_ = new_B2995_ | new_B2972_;
  assign new_B2988_ = ~new_B2973_ ^ new_B2985_;
  assign new_B2989_ = ~new_B2998_ | ~new_B2999_;
  assign new_B2990_ = new_B2974_ ^ new_B2981_;
  assign new_B2991_ = new_B3000_ & new_B2993_;
  assign new_B2992_ = ~new_B3002_ | ~new_B3001_;
  assign new_B2993_ = new_B2974_ | new_B2975_;
  assign new_B2994_ = new_B2974_ | new_B2981_;
  assign new_B2995_ = new_B2973_ & new_B2985_;
  assign new_B2996_ = ~new_B2972_ | ~new_B2973_;
  assign new_B2997_ = new_B2981_ & new_B2996_;
  assign new_B2998_ = ~new_B2997_ & ~new_B2981_;
  assign new_B2999_ = new_B2981_ | new_B2996_;
  assign new_B3000_ = ~new_B2974_ | ~new_B2975_;
  assign new_B3001_ = new_B2981_ | new_B2996_;
  assign new_B3002_ = ~new_B2981_ & ~new_B3003_;
  assign new_B3003_ = new_B2981_ & new_B2996_;
  assign new_B3004_ = new_B6674_;
  assign new_B3005_ = new_B6707_;
  assign new_B3006_ = new_B6740_;
  assign new_B3007_ = new_B6773_;
  assign new_B3008_ = new_B6806_;
  assign new_B3009_ = new_B3015_ & new_B3014_;
  assign new_B3010_ = new_B3017_ | new_B3016_;
  assign new_B3011_ = new_B3019_ | new_B3018_;
  assign new_B3012_ = new_B3014_ & new_B3020_;
  assign new_B3013_ = new_B3014_ & new_B3021_;
  assign new_B3014_ = new_B3004_ ^ new_B3005_;
  assign new_B3015_ = new_B3016_ ^ new_B3006_;
  assign new_B3016_ = new_B3024_ & new_B3023_;
  assign new_B3017_ = new_B3022_ & new_B3006_;
  assign new_B3018_ = new_B3027_ & new_B3026_;
  assign new_B3019_ = new_B3025_ & new_B3006_;
  assign new_B3020_ = new_B3028_ | new_B3005_;
  assign new_B3021_ = ~new_B3006_ ^ new_B3018_;
  assign new_B3022_ = ~new_B3031_ | ~new_B3032_;
  assign new_B3023_ = new_B3007_ ^ new_B3014_;
  assign new_B3024_ = new_B3033_ & new_B3026_;
  assign new_B3025_ = ~new_B3035_ | ~new_B3034_;
  assign new_B3026_ = new_B3007_ | new_B3008_;
  assign new_B3027_ = new_B3007_ | new_B3014_;
  assign new_B3028_ = new_B3006_ & new_B3018_;
  assign new_B3029_ = ~new_B3005_ | ~new_B3006_;
  assign new_B3030_ = new_B3014_ & new_B3029_;
  assign new_B3031_ = ~new_B3030_ & ~new_B3014_;
  assign new_B3032_ = new_B3014_ | new_B3029_;
  assign new_B3033_ = ~new_B3007_ | ~new_B3008_;
  assign new_B3034_ = new_B3014_ | new_B3029_;
  assign new_B3035_ = ~new_B3014_ & ~new_B3036_;
  assign new_B3036_ = new_B3014_ & new_B3029_;
  assign new_B3037_ = new_B6839_;
  assign new_B3038_ = new_B6872_;
  assign new_B3039_ = new_B6905_;
  assign new_B3040_ = new_B6938_;
  assign new_B3041_ = new_B6971_;
  assign new_B3042_ = new_B3048_ & new_B3047_;
  assign new_B3043_ = new_B3050_ | new_B3049_;
  assign new_B3044_ = new_B3052_ | new_B3051_;
  assign new_B3045_ = new_B3047_ & new_B3053_;
  assign new_B3046_ = new_B3047_ & new_B3054_;
  assign new_B3047_ = new_B3037_ ^ new_B3038_;
  assign new_B3048_ = new_B3049_ ^ new_B3039_;
  assign new_B3049_ = new_B3057_ & new_B3056_;
  assign new_B3050_ = new_B3055_ & new_B3039_;
  assign new_B3051_ = new_B3060_ & new_B3059_;
  assign new_B3052_ = new_B3058_ & new_B3039_;
  assign new_B3053_ = new_B3061_ | new_B3038_;
  assign new_B3054_ = ~new_B3039_ ^ new_B3051_;
  assign new_B3055_ = ~new_B3064_ | ~new_B3065_;
  assign new_B3056_ = new_B3040_ ^ new_B3047_;
  assign new_B3057_ = new_B3066_ & new_B3059_;
  assign new_B3058_ = ~new_B3068_ | ~new_B3067_;
  assign new_B3059_ = new_B3040_ | new_B3041_;
  assign new_B3060_ = new_B3040_ | new_B3047_;
  assign new_B3061_ = new_B3039_ & new_B3051_;
  assign new_B3062_ = ~new_B3038_ | ~new_B3039_;
  assign new_B3063_ = new_B3047_ & new_B3062_;
  assign new_B3064_ = ~new_B3063_ & ~new_B3047_;
  assign new_B3065_ = new_B3047_ | new_B3062_;
  assign new_B3066_ = ~new_B3040_ | ~new_B3041_;
  assign new_B3067_ = new_B3047_ | new_B3062_;
  assign new_B3068_ = ~new_B3047_ & ~new_B3069_;
  assign new_B3069_ = new_B3047_ & new_B3062_;
  assign new_B3070_ = new_B7004_;
  assign new_B3071_ = new_B7037_;
  assign new_B3072_ = new_B7070_;
  assign new_B3073_ = new_B7103_;
  assign new_B3074_ = new_B7136_;
  assign new_B3075_ = new_B3081_ & new_B3080_;
  assign new_B3076_ = new_B3083_ | new_B3082_;
  assign new_B3077_ = new_B3085_ | new_B3084_;
  assign new_B3078_ = new_B3080_ & new_B3086_;
  assign new_B3079_ = new_B3080_ & new_B3087_;
  assign new_B3080_ = new_B3070_ ^ new_B3071_;
  assign new_B3081_ = new_B3082_ ^ new_B3072_;
  assign new_B3082_ = new_B3090_ & new_B3089_;
  assign new_B3083_ = new_B3088_ & new_B3072_;
  assign new_B3084_ = new_B3093_ & new_B3092_;
  assign new_B3085_ = new_B3091_ & new_B3072_;
  assign new_B3086_ = new_B3094_ | new_B3071_;
  assign new_B3087_ = ~new_B3072_ ^ new_B3084_;
  assign new_B3088_ = ~new_B3097_ | ~new_B3098_;
  assign new_B3089_ = new_B3073_ ^ new_B3080_;
  assign new_B3090_ = new_B3099_ & new_B3092_;
  assign new_B3091_ = ~new_B3101_ | ~new_B3100_;
  assign new_B3092_ = new_B3073_ | new_B3074_;
  assign new_B3093_ = new_B3073_ | new_B3080_;
  assign new_B3094_ = new_B3072_ & new_B3084_;
  assign new_B3095_ = ~new_B3071_ | ~new_B3072_;
  assign new_B3096_ = new_B3080_ & new_B3095_;
  assign new_B3097_ = ~new_B3096_ & ~new_B3080_;
  assign new_B3098_ = new_B3080_ | new_B3095_;
  assign new_B3099_ = ~new_B3073_ | ~new_B3074_;
  assign new_B3100_ = new_B3080_ | new_B3095_;
  assign new_B3101_ = ~new_B3080_ & ~new_B3102_;
  assign new_B3102_ = new_B3080_ & new_B3095_;
  assign new_B3103_ = new_B7169_;
  assign new_B3104_ = new_B7202_;
  assign new_B3105_ = new_B7235_;
  assign new_B3106_ = new_B7268_;
  assign new_B3107_ = new_B7301_;
  assign new_B3108_ = new_B3114_ & new_B3113_;
  assign new_B3109_ = new_B3116_ | new_B3115_;
  assign new_B3110_ = new_B3118_ | new_B3117_;
  assign new_B3111_ = new_B3113_ & new_B3119_;
  assign new_B3112_ = new_B3113_ & new_B3120_;
  assign new_B3113_ = new_B3103_ ^ new_B3104_;
  assign new_B3114_ = new_B3115_ ^ new_B3105_;
  assign new_B3115_ = new_B3123_ & new_B3122_;
  assign new_B3116_ = new_B3121_ & new_B3105_;
  assign new_B3117_ = new_B3126_ & new_B3125_;
  assign new_B3118_ = new_B3124_ & new_B3105_;
  assign new_B3119_ = new_B3127_ | new_B3104_;
  assign new_B3120_ = ~new_B3105_ ^ new_B3117_;
  assign new_B3121_ = ~new_B3130_ | ~new_B3131_;
  assign new_B3122_ = new_B3106_ ^ new_B3113_;
  assign new_B3123_ = new_B3132_ & new_B3125_;
  assign new_B3124_ = ~new_B3134_ | ~new_B3133_;
  assign new_B3125_ = new_B3106_ | new_B3107_;
  assign new_B3126_ = new_B3106_ | new_B3113_;
  assign new_B3127_ = new_B3105_ & new_B3117_;
  assign new_B3128_ = ~new_B3104_ | ~new_B3105_;
  assign new_B3129_ = new_B3113_ & new_B3128_;
  assign new_B3130_ = ~new_B3129_ & ~new_B3113_;
  assign new_B3131_ = new_B3113_ | new_B3128_;
  assign new_B3132_ = ~new_B3106_ | ~new_B3107_;
  assign new_B3133_ = new_B3113_ | new_B3128_;
  assign new_B3134_ = ~new_B3113_ & ~new_B3135_;
  assign new_B3135_ = new_B3113_ & new_B3128_;
  assign new_B3136_ = new_B7334_;
  assign new_B3137_ = new_B7367_;
  assign new_B3138_ = new_B7400_;
  assign new_B3139_ = new_B7433_;
  assign new_B3140_ = new_B7466_;
  assign new_B3141_ = new_B3147_ & new_B3146_;
  assign new_B3142_ = new_B3149_ | new_B3148_;
  assign new_B3143_ = new_B3151_ | new_B3150_;
  assign new_B3144_ = new_B3146_ & new_B3152_;
  assign new_B3145_ = new_B3146_ & new_B3153_;
  assign new_B3146_ = new_B3136_ ^ new_B3137_;
  assign new_B3147_ = new_B3148_ ^ new_B3138_;
  assign new_B3148_ = new_B3156_ & new_B3155_;
  assign new_B3149_ = new_B3154_ & new_B3138_;
  assign new_B3150_ = new_B3159_ & new_B3158_;
  assign new_B3151_ = new_B3157_ & new_B3138_;
  assign new_B3152_ = new_B3160_ | new_B3137_;
  assign new_B3153_ = ~new_B3138_ ^ new_B3150_;
  assign new_B3154_ = ~new_B3163_ | ~new_B3164_;
  assign new_B3155_ = new_B3139_ ^ new_B3146_;
  assign new_B3156_ = new_B3165_ & new_B3158_;
  assign new_B3157_ = ~new_B3167_ | ~new_B3166_;
  assign new_B3158_ = new_B3139_ | new_B3140_;
  assign new_B3159_ = new_B3139_ | new_B3146_;
  assign new_B3160_ = new_B3138_ & new_B3150_;
  assign new_B3161_ = ~new_B3137_ | ~new_B3138_;
  assign new_B3162_ = new_B3146_ & new_B3161_;
  assign new_B3163_ = ~new_B3162_ & ~new_B3146_;
  assign new_B3164_ = new_B3146_ | new_B3161_;
  assign new_B3165_ = ~new_B3139_ | ~new_B3140_;
  assign new_B3166_ = new_B3146_ | new_B3161_;
  assign new_B3167_ = ~new_B3146_ & ~new_B3168_;
  assign new_B3168_ = new_B3146_ & new_B3161_;
  assign new_B3169_ = new_B7499_;
  assign new_B3170_ = new_B7532_;
  assign new_B3171_ = new_B7565_;
  assign new_B3172_ = new_B7598_;
  assign new_B3173_ = new_B7631_;
  assign new_B3174_ = new_B3180_ & new_B3179_;
  assign new_B3175_ = new_B3182_ | new_B3181_;
  assign new_B3176_ = new_B3184_ | new_B3183_;
  assign new_B3177_ = new_B3179_ & new_B3185_;
  assign new_B3178_ = new_B3179_ & new_B3186_;
  assign new_B3179_ = new_B3169_ ^ new_B3170_;
  assign new_B3180_ = new_B3181_ ^ new_B3171_;
  assign new_B3181_ = new_B3189_ & new_B3188_;
  assign new_B3182_ = new_B3187_ & new_B3171_;
  assign new_B3183_ = new_B3192_ & new_B3191_;
  assign new_B3184_ = new_B3190_ & new_B3171_;
  assign new_B3185_ = new_B3193_ | new_B3170_;
  assign new_B3186_ = ~new_B3171_ ^ new_B3183_;
  assign new_B3187_ = ~new_B3196_ | ~new_B3197_;
  assign new_B3188_ = new_B3172_ ^ new_B3179_;
  assign new_B3189_ = new_B3198_ & new_B3191_;
  assign new_B3190_ = ~new_B3200_ | ~new_B3199_;
  assign new_B3191_ = new_B3172_ | new_B3173_;
  assign new_B3192_ = new_B3172_ | new_B3179_;
  assign new_B3193_ = new_B3171_ & new_B3183_;
  assign new_B3194_ = ~new_B3170_ | ~new_B3171_;
  assign new_B3195_ = new_B3179_ & new_B3194_;
  assign new_B3196_ = ~new_B3195_ & ~new_B3179_;
  assign new_B3197_ = new_B3179_ | new_B3194_;
  assign new_B3198_ = ~new_B3172_ | ~new_B3173_;
  assign new_B3199_ = new_B3179_ | new_B3194_;
  assign new_B3200_ = ~new_B3179_ & ~new_B3201_;
  assign new_B3201_ = new_B3179_ & new_B3194_;
  assign new_B3202_ = new_B7664_;
  assign new_B3203_ = new_B7697_;
  assign new_B3204_ = new_B7730_;
  assign new_B3205_ = new_B7763_;
  assign new_B3206_ = new_B7796_;
  assign new_B3207_ = new_B3213_ & new_B3212_;
  assign new_B3208_ = new_B3215_ | new_B3214_;
  assign new_B3209_ = new_B3217_ | new_B3216_;
  assign new_B3210_ = new_B3212_ & new_B3218_;
  assign new_B3211_ = new_B3212_ & new_B3219_;
  assign new_B3212_ = new_B3202_ ^ new_B3203_;
  assign new_B3213_ = new_B3214_ ^ new_B3204_;
  assign new_B3214_ = new_B3222_ & new_B3221_;
  assign new_B3215_ = new_B3220_ & new_B3204_;
  assign new_B3216_ = new_B3225_ & new_B3224_;
  assign new_B3217_ = new_B3223_ & new_B3204_;
  assign new_B3218_ = new_B3226_ | new_B3203_;
  assign new_B3219_ = ~new_B3204_ ^ new_B3216_;
  assign new_B3220_ = ~new_B3229_ | ~new_B3230_;
  assign new_B3221_ = new_B3205_ ^ new_B3212_;
  assign new_B3222_ = new_B3231_ & new_B3224_;
  assign new_B3223_ = ~new_B3233_ | ~new_B3232_;
  assign new_B3224_ = new_B3205_ | new_B3206_;
  assign new_B3225_ = new_B3205_ | new_B3212_;
  assign new_B3226_ = new_B3204_ & new_B3216_;
  assign new_B3227_ = ~new_B3203_ | ~new_B3204_;
  assign new_B3228_ = new_B3212_ & new_B3227_;
  assign new_B3229_ = ~new_B3228_ & ~new_B3212_;
  assign new_B3230_ = new_B3212_ | new_B3227_;
  assign new_B3231_ = ~new_B3205_ | ~new_B3206_;
  assign new_B3232_ = new_B3212_ | new_B3227_;
  assign new_B3233_ = ~new_B3212_ & ~new_B3234_;
  assign new_B3234_ = new_B3212_ & new_B3227_;
  assign new_B3235_ = new_B7829_;
  assign new_B3236_ = new_B7862_;
  assign new_B3237_ = new_B7895_;
  assign new_B3238_ = new_B7928_;
  assign new_B3239_ = new_B7961_;
  assign new_B3240_ = new_B3246_ & new_B3245_;
  assign new_B3241_ = new_B3248_ | new_B3247_;
  assign new_B3242_ = new_B3250_ | new_B3249_;
  assign new_B3243_ = new_B3245_ & new_B3251_;
  assign new_B3244_ = new_B3245_ & new_B3252_;
  assign new_B3245_ = new_B3235_ ^ new_B3236_;
  assign new_B3246_ = new_B3247_ ^ new_B3237_;
  assign new_B3247_ = new_B3255_ & new_B3254_;
  assign new_B3248_ = new_B3253_ & new_B3237_;
  assign new_B3249_ = new_B3258_ & new_B3257_;
  assign new_B3250_ = new_B3256_ & new_B3237_;
  assign new_B3251_ = new_B3259_ | new_B3236_;
  assign new_B3252_ = ~new_B3237_ ^ new_B3249_;
  assign new_B3253_ = ~new_B3262_ | ~new_B3263_;
  assign new_B3254_ = new_B3238_ ^ new_B3245_;
  assign new_B3255_ = new_B3264_ & new_B3257_;
  assign new_B3256_ = ~new_B3266_ | ~new_B3265_;
  assign new_B3257_ = new_B3238_ | new_B3239_;
  assign new_B3258_ = new_B3238_ | new_B3245_;
  assign new_B3259_ = new_B3237_ & new_B3249_;
  assign new_B3260_ = ~new_B3236_ | ~new_B3237_;
  assign new_B3261_ = new_B3245_ & new_B3260_;
  assign new_B3262_ = ~new_B3261_ & ~new_B3245_;
  assign new_B3263_ = new_B3245_ | new_B3260_;
  assign new_B3264_ = ~new_B3238_ | ~new_B3239_;
  assign new_B3265_ = new_B3245_ | new_B3260_;
  assign new_B3266_ = ~new_B3245_ & ~new_B3267_;
  assign new_B3267_ = new_B3245_ & new_B3260_;
  assign new_B3268_ = new_B7994_;
  assign new_B3269_ = new_B8027_;
  assign new_B3270_ = new_B8060_;
  assign new_B3271_ = new_B8093_;
  assign new_B3272_ = new_B8126_;
  assign new_B3273_ = new_B3279_ & new_B3278_;
  assign new_B3274_ = new_B3281_ | new_B3280_;
  assign new_B3275_ = new_B3283_ | new_B3282_;
  assign new_B3276_ = new_B3278_ & new_B3284_;
  assign new_B3277_ = new_B3278_ & new_B3285_;
  assign new_B3278_ = new_B3268_ ^ new_B3269_;
  assign new_B3279_ = new_B3280_ ^ new_B3270_;
  assign new_B3280_ = new_B3288_ & new_B3287_;
  assign new_B3281_ = new_B3286_ & new_B3270_;
  assign new_B3282_ = new_B3291_ & new_B3290_;
  assign new_B3283_ = new_B3289_ & new_B3270_;
  assign new_B3284_ = new_B3292_ | new_B3269_;
  assign new_B3285_ = ~new_B3270_ ^ new_B3282_;
  assign new_B3286_ = ~new_B3295_ | ~new_B3296_;
  assign new_B3287_ = new_B3271_ ^ new_B3278_;
  assign new_B3288_ = new_B3297_ & new_B3290_;
  assign new_B3289_ = ~new_B3299_ | ~new_B3298_;
  assign new_B3290_ = new_B3271_ | new_B3272_;
  assign new_B3291_ = new_B3271_ | new_B3278_;
  assign new_B3292_ = new_B3270_ & new_B3282_;
  assign new_B3293_ = ~new_B3269_ | ~new_B3270_;
  assign new_B3294_ = new_B3278_ & new_B3293_;
  assign new_B3295_ = ~new_B3294_ & ~new_B3278_;
  assign new_B3296_ = new_B3278_ | new_B3293_;
  assign new_B3297_ = ~new_B3271_ | ~new_B3272_;
  assign new_B3298_ = new_B3278_ | new_B3293_;
  assign new_B3299_ = ~new_B3278_ & ~new_B3300_;
  assign new_B3300_ = new_B3278_ & new_B3293_;
  assign new_B3301_ = new_B8159_;
  assign new_B3302_ = new_B8192_;
  assign new_B3303_ = new_B8225_;
  assign new_B3304_ = new_B8258_;
  assign new_B3305_ = new_B8291_;
  assign new_B3306_ = new_B3312_ & new_B3311_;
  assign new_B3307_ = new_B3314_ | new_B3313_;
  assign new_B3308_ = new_B3316_ | new_B3315_;
  assign new_B3309_ = new_B3311_ & new_B3317_;
  assign new_B3310_ = new_B3311_ & new_B3318_;
  assign new_B3311_ = new_B3301_ ^ new_B3302_;
  assign new_B3312_ = new_B3313_ ^ new_B3303_;
  assign new_B3313_ = new_B3321_ & new_B3320_;
  assign new_B3314_ = new_B3319_ & new_B3303_;
  assign new_B3315_ = new_B3324_ & new_B3323_;
  assign new_B3316_ = new_B3322_ & new_B3303_;
  assign new_B3317_ = new_B3325_ | new_B3302_;
  assign new_B3318_ = ~new_B3303_ ^ new_B3315_;
  assign new_B3319_ = ~new_B3328_ | ~new_B3329_;
  assign new_B3320_ = new_B3304_ ^ new_B3311_;
  assign new_B3321_ = new_B3330_ & new_B3323_;
  assign new_B3322_ = ~new_B3332_ | ~new_B3331_;
  assign new_B3323_ = new_B3304_ | new_B3305_;
  assign new_B3324_ = new_B3304_ | new_B3311_;
  assign new_B3325_ = new_B3303_ & new_B3315_;
  assign new_B3326_ = ~new_B3302_ | ~new_B3303_;
  assign new_B3327_ = new_B3311_ & new_B3326_;
  assign new_B3328_ = ~new_B3327_ & ~new_B3311_;
  assign new_B3329_ = new_B3311_ | new_B3326_;
  assign new_B3330_ = ~new_B3304_ | ~new_B3305_;
  assign new_B3331_ = new_B3311_ | new_B3326_;
  assign new_B3332_ = ~new_B3311_ & ~new_B3333_;
  assign new_B3333_ = new_B3311_ & new_B3326_;
  assign new_B3334_ = new_B8324_;
  assign new_B3335_ = new_B8357_;
  assign new_B3336_ = new_B8390_;
  assign new_B3337_ = new_B8423_;
  assign new_B3338_ = new_B8456_;
  assign new_B3339_ = new_B3345_ & new_B3344_;
  assign new_B3340_ = new_B3347_ | new_B3346_;
  assign new_B3341_ = new_B3349_ | new_B3348_;
  assign new_B3342_ = new_B3344_ & new_B3350_;
  assign new_B3343_ = new_B3344_ & new_B3351_;
  assign new_B3344_ = new_B3334_ ^ new_B3335_;
  assign new_B3345_ = new_B3346_ ^ new_B3336_;
  assign new_B3346_ = new_B3354_ & new_B3353_;
  assign new_B3347_ = new_B3352_ & new_B3336_;
  assign new_B3348_ = new_B3357_ & new_B3356_;
  assign new_B3349_ = new_B3355_ & new_B3336_;
  assign new_B3350_ = new_B3358_ | new_B3335_;
  assign new_B3351_ = ~new_B3336_ ^ new_B3348_;
  assign new_B3352_ = ~new_B3361_ | ~new_B3362_;
  assign new_B3353_ = new_B3337_ ^ new_B3344_;
  assign new_B3354_ = new_B3363_ & new_B3356_;
  assign new_B3355_ = ~new_B3365_ | ~new_B3364_;
  assign new_B3356_ = new_B3337_ | new_B3338_;
  assign new_B3357_ = new_B3337_ | new_B3344_;
  assign new_B3358_ = new_B3336_ & new_B3348_;
  assign new_B3359_ = ~new_B3335_ | ~new_B3336_;
  assign new_B3360_ = new_B3344_ & new_B3359_;
  assign new_B3361_ = ~new_B3360_ & ~new_B3344_;
  assign new_B3362_ = new_B3344_ | new_B3359_;
  assign new_B3363_ = ~new_B3337_ | ~new_B3338_;
  assign new_B3364_ = new_B3344_ | new_B3359_;
  assign new_B3365_ = ~new_B3344_ & ~new_B3366_;
  assign new_B3366_ = new_B3344_ & new_B3359_;
  assign new_B3367_ = new_B8489_;
  assign new_B3368_ = new_B8522_;
  assign new_B3369_ = new_B8555_;
  assign new_B3370_ = new_B8588_;
  assign new_B3371_ = new_B8621_;
  assign new_B3372_ = new_B3378_ & new_B3377_;
  assign new_B3373_ = new_B3380_ | new_B3379_;
  assign new_B3374_ = new_B3382_ | new_B3381_;
  assign new_B3375_ = new_B3377_ & new_B3383_;
  assign new_B3376_ = new_B3377_ & new_B3384_;
  assign new_B3377_ = new_B3367_ ^ new_B3368_;
  assign new_B3378_ = new_B3379_ ^ new_B3369_;
  assign new_B3379_ = new_B3387_ & new_B3386_;
  assign new_B3380_ = new_B3385_ & new_B3369_;
  assign new_B3381_ = new_B3390_ & new_B3389_;
  assign new_B3382_ = new_B3388_ & new_B3369_;
  assign new_B3383_ = new_B3391_ | new_B3368_;
  assign new_B3384_ = ~new_B3369_ ^ new_B3381_;
  assign new_B3385_ = ~new_B3394_ | ~new_B3395_;
  assign new_B3386_ = new_B3370_ ^ new_B3377_;
  assign new_B3387_ = new_B3396_ & new_B3389_;
  assign new_B3388_ = ~new_B3398_ | ~new_B3397_;
  assign new_B3389_ = new_B3370_ | new_B3371_;
  assign new_B3390_ = new_B3370_ | new_B3377_;
  assign new_B3391_ = new_B3369_ & new_B3381_;
  assign new_B3392_ = ~new_B3368_ | ~new_B3369_;
  assign new_B3393_ = new_B3377_ & new_B3392_;
  assign new_B3394_ = ~new_B3393_ & ~new_B3377_;
  assign new_B3395_ = new_B3377_ | new_B3392_;
  assign new_B3396_ = ~new_B3370_ | ~new_B3371_;
  assign new_B3397_ = new_B3377_ | new_B3392_;
  assign new_B3398_ = ~new_B3377_ & ~new_B3399_;
  assign new_B3399_ = new_B3377_ & new_B3392_;
  assign new_B3400_ = new_B8654_;
  assign new_B3401_ = new_B8687_;
  assign new_B3402_ = new_B8720_;
  assign new_B3403_ = new_B8753_;
  assign new_B3404_ = new_B8786_;
  assign new_B3405_ = new_B3411_ & new_B3410_;
  assign new_B3406_ = new_B3413_ | new_B3412_;
  assign new_B3407_ = new_B3415_ | new_B3414_;
  assign new_B3408_ = new_B3410_ & new_B3416_;
  assign new_B3409_ = new_B3410_ & new_B3417_;
  assign new_B3410_ = new_B3400_ ^ new_B3401_;
  assign new_B3411_ = new_B3412_ ^ new_B3402_;
  assign new_B3412_ = new_B3420_ & new_B3419_;
  assign new_B3413_ = new_B3418_ & new_B3402_;
  assign new_B3414_ = new_B3423_ & new_B3422_;
  assign new_B3415_ = new_B3421_ & new_B3402_;
  assign new_B3416_ = new_B3424_ | new_B3401_;
  assign new_B3417_ = ~new_B3402_ ^ new_B3414_;
  assign new_B3418_ = ~new_B3427_ | ~new_B3428_;
  assign new_B3419_ = new_B3403_ ^ new_B3410_;
  assign new_B3420_ = new_B3429_ & new_B3422_;
  assign new_B3421_ = ~new_B3431_ | ~new_B3430_;
  assign new_B3422_ = new_B3403_ | new_B3404_;
  assign new_B3423_ = new_B3403_ | new_B3410_;
  assign new_B3424_ = new_B3402_ & new_B3414_;
  assign new_B3425_ = ~new_B3401_ | ~new_B3402_;
  assign new_B3426_ = new_B3410_ & new_B3425_;
  assign new_B3427_ = ~new_B3426_ & ~new_B3410_;
  assign new_B3428_ = new_B3410_ | new_B3425_;
  assign new_B3429_ = ~new_B3403_ | ~new_B3404_;
  assign new_B3430_ = new_B3410_ | new_B3425_;
  assign new_B3431_ = ~new_B3410_ & ~new_B3432_;
  assign new_B3432_ = new_B3410_ & new_B3425_;
  assign new_B3433_ = new_B8819_;
  assign new_B3434_ = new_B8852_;
  assign new_B3435_ = new_B8885_;
  assign new_B3436_ = new_B8918_;
  assign new_B3437_ = new_B8951_;
  assign new_B3438_ = new_B3444_ & new_B3443_;
  assign new_B3439_ = new_B3446_ | new_B3445_;
  assign new_B3440_ = new_B3448_ | new_B3447_;
  assign new_B3441_ = new_B3443_ & new_B3449_;
  assign new_B3442_ = new_B3443_ & new_B3450_;
  assign new_B3443_ = new_B3433_ ^ new_B3434_;
  assign new_B3444_ = new_B3445_ ^ new_B3435_;
  assign new_B3445_ = new_B3453_ & new_B3452_;
  assign new_B3446_ = new_B3451_ & new_B3435_;
  assign new_B3447_ = new_B3456_ & new_B3455_;
  assign new_B3448_ = new_B3454_ & new_B3435_;
  assign new_B3449_ = new_B3457_ | new_B3434_;
  assign new_B3450_ = ~new_B3435_ ^ new_B3447_;
  assign new_B3451_ = ~new_B3460_ | ~new_B3461_;
  assign new_B3452_ = new_B3436_ ^ new_B3443_;
  assign new_B3453_ = new_B3462_ & new_B3455_;
  assign new_B3454_ = ~new_B3464_ | ~new_B3463_;
  assign new_B3455_ = new_B3436_ | new_B3437_;
  assign new_B3456_ = new_B3436_ | new_B3443_;
  assign new_B3457_ = new_B3435_ & new_B3447_;
  assign new_B3458_ = ~new_B3434_ | ~new_B3435_;
  assign new_B3459_ = new_B3443_ & new_B3458_;
  assign new_B3460_ = ~new_B3459_ & ~new_B3443_;
  assign new_B3461_ = new_B3443_ | new_B3458_;
  assign new_B3462_ = ~new_B3436_ | ~new_B3437_;
  assign new_B3463_ = new_B3443_ | new_B3458_;
  assign new_B3464_ = ~new_B3443_ & ~new_B3465_;
  assign new_B3465_ = new_B3443_ & new_B3458_;
  assign new_B3466_ = new_B8984_;
  assign new_B3467_ = new_B9017_;
  assign new_B3468_ = new_B9050_;
  assign new_B3469_ = new_B9083_;
  assign new_B3470_ = new_B9116_;
  assign new_B3471_ = new_B3477_ & new_B3476_;
  assign new_B3472_ = new_B3479_ | new_B3478_;
  assign new_B3473_ = new_B3481_ | new_B3480_;
  assign new_B3474_ = new_B3476_ & new_B3482_;
  assign new_B3475_ = new_B3476_ & new_B3483_;
  assign new_B3476_ = new_B3466_ ^ new_B3467_;
  assign new_B3477_ = new_B3478_ ^ new_B3468_;
  assign new_B3478_ = new_B3486_ & new_B3485_;
  assign new_B3479_ = new_B3484_ & new_B3468_;
  assign new_B3480_ = new_B3489_ & new_B3488_;
  assign new_B3481_ = new_B3487_ & new_B3468_;
  assign new_B3482_ = new_B3490_ | new_B3467_;
  assign new_B3483_ = ~new_B3468_ ^ new_B3480_;
  assign new_B3484_ = ~new_B3493_ | ~new_B3494_;
  assign new_B3485_ = new_B3469_ ^ new_B3476_;
  assign new_B3486_ = new_B3495_ & new_B3488_;
  assign new_B3487_ = ~new_B3497_ | ~new_B3496_;
  assign new_B3488_ = new_B3469_ | new_B3470_;
  assign new_B3489_ = new_B3469_ | new_B3476_;
  assign new_B3490_ = new_B3468_ & new_B3480_;
  assign new_B3491_ = ~new_B3467_ | ~new_B3468_;
  assign new_B3492_ = new_B3476_ & new_B3491_;
  assign new_B3493_ = ~new_B3492_ & ~new_B3476_;
  assign new_B3494_ = new_B3476_ | new_B3491_;
  assign new_B3495_ = ~new_B3469_ | ~new_B3470_;
  assign new_B3496_ = new_B3476_ | new_B3491_;
  assign new_B3497_ = ~new_B3476_ & ~new_B3498_;
  assign new_B3498_ = new_B3476_ & new_B3491_;
  assign new_B3499_ = new_B9149_;
  assign new_B3500_ = new_B9182_;
  assign new_B3501_ = new_B9215_;
  assign new_B3502_ = new_B9248_;
  assign new_B3503_ = new_B9281_;
  assign new_B3504_ = new_B3510_ & new_B3509_;
  assign new_B3505_ = new_B3512_ | new_B3511_;
  assign new_B3506_ = new_B3514_ | new_B3513_;
  assign new_B3507_ = new_B3509_ & new_B3515_;
  assign new_B3508_ = new_B3509_ & new_B3516_;
  assign new_B3509_ = new_B3499_ ^ new_B3500_;
  assign new_B3510_ = new_B3511_ ^ new_B3501_;
  assign new_B3511_ = new_B3519_ & new_B3518_;
  assign new_B3512_ = new_B3517_ & new_B3501_;
  assign new_B3513_ = new_B3522_ & new_B3521_;
  assign new_B3514_ = new_B3520_ & new_B3501_;
  assign new_B3515_ = new_B3523_ | new_B3500_;
  assign new_B3516_ = ~new_B3501_ ^ new_B3513_;
  assign new_B3517_ = ~new_B3526_ | ~new_B3527_;
  assign new_B3518_ = new_B3502_ ^ new_B3509_;
  assign new_B3519_ = new_B3528_ & new_B3521_;
  assign new_B3520_ = ~new_B3530_ | ~new_B3529_;
  assign new_B3521_ = new_B3502_ | new_B3503_;
  assign new_B3522_ = new_B3502_ | new_B3509_;
  assign new_B3523_ = new_B3501_ & new_B3513_;
  assign new_B3524_ = ~new_B3500_ | ~new_B3501_;
  assign new_B3525_ = new_B3509_ & new_B3524_;
  assign new_B3526_ = ~new_B3525_ & ~new_B3509_;
  assign new_B3527_ = new_B3509_ | new_B3524_;
  assign new_B3528_ = ~new_B3502_ | ~new_B3503_;
  assign new_B3529_ = new_B3509_ | new_B3524_;
  assign new_B3530_ = ~new_B3509_ & ~new_B3531_;
  assign new_B3531_ = new_B3509_ & new_B3524_;
  assign new_B3532_ = new_B5188_;
  assign new_B3533_ = new_B5223_;
  assign new_B3534_ = new_B5256_;
  assign new_B3535_ = new_B5289_;
  assign new_B3536_ = new_B5322_;
  assign new_B3537_ = new_B3543_ & new_B3542_;
  assign new_B3538_ = new_B3545_ | new_B3544_;
  assign new_B3539_ = new_B3547_ | new_B3546_;
  assign new_B3540_ = new_B3542_ & new_B3548_;
  assign new_B3541_ = new_B3542_ & new_B3549_;
  assign new_B3542_ = new_B3532_ ^ new_B3533_;
  assign new_B3543_ = new_B3544_ ^ new_B3534_;
  assign new_B3544_ = new_B3552_ & new_B3551_;
  assign new_B3545_ = new_B3550_ & new_B3534_;
  assign new_B3546_ = new_B3555_ & new_B3554_;
  assign new_B3547_ = new_B3553_ & new_B3534_;
  assign new_B3548_ = new_B3556_ | new_B3533_;
  assign new_B3549_ = ~new_B3534_ ^ new_B3546_;
  assign new_B3550_ = ~new_B3559_ | ~new_B3560_;
  assign new_B3551_ = new_B3535_ ^ new_B3542_;
  assign new_B3552_ = new_B3561_ & new_B3554_;
  assign new_B3553_ = ~new_B3563_ | ~new_B3562_;
  assign new_B3554_ = new_B3535_ | new_B3536_;
  assign new_B3555_ = new_B3535_ | new_B3542_;
  assign new_B3556_ = new_B3534_ & new_B3546_;
  assign new_B3557_ = ~new_B3533_ | ~new_B3534_;
  assign new_B3558_ = new_B3542_ & new_B3557_;
  assign new_B3559_ = ~new_B3558_ & ~new_B3542_;
  assign new_B3560_ = new_B3542_ | new_B3557_;
  assign new_B3561_ = ~new_B3535_ | ~new_B3536_;
  assign new_B3562_ = new_B3542_ | new_B3557_;
  assign new_B3563_ = ~new_B3542_ & ~new_B3564_;
  assign new_B3564_ = new_B3542_ & new_B3557_;
  assign new_B3565_ = new_B5355_;
  assign new_B3566_ = new_B5388_;
  assign new_B3567_ = new_B5421_;
  assign new_B3568_ = new_B5454_;
  assign new_B3569_ = new_B5487_;
  assign new_B3570_ = new_B3576_ & new_B3575_;
  assign new_B3571_ = new_B3578_ | new_B3577_;
  assign new_B3572_ = new_B3580_ | new_B3579_;
  assign new_B3573_ = new_B3575_ & new_B3581_;
  assign new_B3574_ = new_B3575_ & new_B3582_;
  assign new_B3575_ = new_B3565_ ^ new_B3566_;
  assign new_B3576_ = new_B3577_ ^ new_B3567_;
  assign new_B3577_ = new_B3585_ & new_B3584_;
  assign new_B3578_ = new_B3583_ & new_B3567_;
  assign new_B3579_ = new_B3588_ & new_B3587_;
  assign new_B3580_ = new_B3586_ & new_B3567_;
  assign new_B3581_ = new_B3589_ | new_B3566_;
  assign new_B3582_ = ~new_B3567_ ^ new_B3579_;
  assign new_B3583_ = ~new_B3592_ | ~new_B3593_;
  assign new_B3584_ = new_B3568_ ^ new_B3575_;
  assign new_B3585_ = new_B3594_ & new_B3587_;
  assign new_B3586_ = ~new_B3596_ | ~new_B3595_;
  assign new_B3587_ = new_B3568_ | new_B3569_;
  assign new_B3588_ = new_B3568_ | new_B3575_;
  assign new_B3589_ = new_B3567_ & new_B3579_;
  assign new_B3590_ = ~new_B3566_ | ~new_B3567_;
  assign new_B3591_ = new_B3575_ & new_B3590_;
  assign new_B3592_ = ~new_B3591_ & ~new_B3575_;
  assign new_B3593_ = new_B3575_ | new_B3590_;
  assign new_B3594_ = ~new_B3568_ | ~new_B3569_;
  assign new_B3595_ = new_B3575_ | new_B3590_;
  assign new_B3596_ = ~new_B3575_ & ~new_B3597_;
  assign new_B3597_ = new_B3575_ & new_B3590_;
  assign new_B3598_ = new_B5520_;
  assign new_B3599_ = new_B5553_;
  assign new_B3600_ = new_B5586_;
  assign new_B3601_ = new_B5619_;
  assign new_B3602_ = new_B5652_;
  assign new_B3603_ = new_B3609_ & new_B3608_;
  assign new_B3604_ = new_B3611_ | new_B3610_;
  assign new_B3605_ = new_B3613_ | new_B3612_;
  assign new_B3606_ = new_B3608_ & new_B3614_;
  assign new_B3607_ = new_B3608_ & new_B3615_;
  assign new_B3608_ = new_B3598_ ^ new_B3599_;
  assign new_B3609_ = new_B3610_ ^ new_B3600_;
  assign new_B3610_ = new_B3618_ & new_B3617_;
  assign new_B3611_ = new_B3616_ & new_B3600_;
  assign new_B3612_ = new_B3621_ & new_B3620_;
  assign new_B3613_ = new_B3619_ & new_B3600_;
  assign new_B3614_ = new_B3622_ | new_B3599_;
  assign new_B3615_ = ~new_B3600_ ^ new_B3612_;
  assign new_B3616_ = ~new_B3625_ | ~new_B3626_;
  assign new_B3617_ = new_B3601_ ^ new_B3608_;
  assign new_B3618_ = new_B3627_ & new_B3620_;
  assign new_B3619_ = ~new_B3629_ | ~new_B3628_;
  assign new_B3620_ = new_B3601_ | new_B3602_;
  assign new_B3621_ = new_B3601_ | new_B3608_;
  assign new_B3622_ = new_B3600_ & new_B3612_;
  assign new_B3623_ = ~new_B3599_ | ~new_B3600_;
  assign new_B3624_ = new_B3608_ & new_B3623_;
  assign new_B3625_ = ~new_B3624_ & ~new_B3608_;
  assign new_B3626_ = new_B3608_ | new_B3623_;
  assign new_B3627_ = ~new_B3601_ | ~new_B3602_;
  assign new_B3628_ = new_B3608_ | new_B3623_;
  assign new_B3629_ = ~new_B3608_ & ~new_B3630_;
  assign new_B3630_ = new_B3608_ & new_B3623_;
  assign new_B3631_ = new_B5685_;
  assign new_B3632_ = new_B5718_;
  assign new_B3633_ = new_B5751_;
  assign new_B3634_ = new_B5784_;
  assign new_B3635_ = new_B5817_;
  assign new_B3636_ = new_B3642_ & new_B3641_;
  assign new_B3637_ = new_B3644_ | new_B3643_;
  assign new_B3638_ = new_B3646_ | new_B3645_;
  assign new_B3639_ = new_B3641_ & new_B3647_;
  assign new_B3640_ = new_B3641_ & new_B3648_;
  assign new_B3641_ = new_B3631_ ^ new_B3632_;
  assign new_B3642_ = new_B3643_ ^ new_B3633_;
  assign new_B3643_ = new_B3651_ & new_B3650_;
  assign new_B3644_ = new_B3649_ & new_B3633_;
  assign new_B3645_ = new_B3654_ & new_B3653_;
  assign new_B3646_ = new_B3652_ & new_B3633_;
  assign new_B3647_ = new_B3655_ | new_B3632_;
  assign new_B3648_ = ~new_B3633_ ^ new_B3645_;
  assign new_B3649_ = ~new_B3658_ | ~new_B3659_;
  assign new_B3650_ = new_B3634_ ^ new_B3641_;
  assign new_B3651_ = new_B3660_ & new_B3653_;
  assign new_B3652_ = ~new_B3662_ | ~new_B3661_;
  assign new_B3653_ = new_B3634_ | new_B3635_;
  assign new_B3654_ = new_B3634_ | new_B3641_;
  assign new_B3655_ = new_B3633_ & new_B3645_;
  assign new_B3656_ = ~new_B3632_ | ~new_B3633_;
  assign new_B3657_ = new_B3641_ & new_B3656_;
  assign new_B3658_ = ~new_B3657_ & ~new_B3641_;
  assign new_B3659_ = new_B3641_ | new_B3656_;
  assign new_B3660_ = ~new_B3634_ | ~new_B3635_;
  assign new_B3661_ = new_B3641_ | new_B3656_;
  assign new_B3662_ = ~new_B3641_ & ~new_B3663_;
  assign new_B3663_ = new_B3641_ & new_B3656_;
  assign new_B3664_ = new_B5850_;
  assign new_B3665_ = new_B5883_;
  assign new_B3666_ = new_B5916_;
  assign new_B3667_ = new_B5949_;
  assign new_B3668_ = new_B5982_;
  assign new_B3669_ = new_B3675_ & new_B3674_;
  assign new_B3670_ = new_B3677_ | new_B3676_;
  assign new_B3671_ = new_B3679_ | new_B3678_;
  assign new_B3672_ = new_B3674_ & new_B3680_;
  assign new_B3673_ = new_B3674_ & new_B3681_;
  assign new_B3674_ = new_B3664_ ^ new_B3665_;
  assign new_B3675_ = new_B3676_ ^ new_B3666_;
  assign new_B3676_ = new_B3684_ & new_B3683_;
  assign new_B3677_ = new_B3682_ & new_B3666_;
  assign new_B3678_ = new_B3687_ & new_B3686_;
  assign new_B3679_ = new_B3685_ & new_B3666_;
  assign new_B3680_ = new_B3688_ | new_B3665_;
  assign new_B3681_ = ~new_B3666_ ^ new_B3678_;
  assign new_B3682_ = ~new_B3691_ | ~new_B3692_;
  assign new_B3683_ = new_B3667_ ^ new_B3674_;
  assign new_B3684_ = new_B3693_ & new_B3686_;
  assign new_B3685_ = ~new_B3695_ | ~new_B3694_;
  assign new_B3686_ = new_B3667_ | new_B3668_;
  assign new_B3687_ = new_B3667_ | new_B3674_;
  assign new_B3688_ = new_B3666_ & new_B3678_;
  assign new_B3689_ = ~new_B3665_ | ~new_B3666_;
  assign new_B3690_ = new_B3674_ & new_B3689_;
  assign new_B3691_ = ~new_B3690_ & ~new_B3674_;
  assign new_B3692_ = new_B3674_ | new_B3689_;
  assign new_B3693_ = ~new_B3667_ | ~new_B3668_;
  assign new_B3694_ = new_B3674_ | new_B3689_;
  assign new_B3695_ = ~new_B3674_ & ~new_B3696_;
  assign new_B3696_ = new_B3674_ & new_B3689_;
  assign new_B3697_ = new_B6015_;
  assign new_B3698_ = new_B6048_;
  assign new_B3699_ = new_B6081_;
  assign new_B3700_ = new_B6114_;
  assign new_B3701_ = new_B6147_;
  assign new_B3702_ = new_B3708_ & new_B3707_;
  assign new_B3703_ = new_B3710_ | new_B3709_;
  assign new_B3704_ = new_B3712_ | new_B3711_;
  assign new_B3705_ = new_B3707_ & new_B3713_;
  assign new_B3706_ = new_B3707_ & new_B3714_;
  assign new_B3707_ = new_B3697_ ^ new_B3698_;
  assign new_B3708_ = new_B3709_ ^ new_B3699_;
  assign new_B3709_ = new_B3717_ & new_B3716_;
  assign new_B3710_ = new_B3715_ & new_B3699_;
  assign new_B3711_ = new_B3720_ & new_B3719_;
  assign new_B3712_ = new_B3718_ & new_B3699_;
  assign new_B3713_ = new_B3721_ | new_B3698_;
  assign new_B3714_ = ~new_B3699_ ^ new_B3711_;
  assign new_B3715_ = ~new_B3724_ | ~new_B3725_;
  assign new_B3716_ = new_B3700_ ^ new_B3707_;
  assign new_B3717_ = new_B3726_ & new_B3719_;
  assign new_B3718_ = ~new_B3728_ | ~new_B3727_;
  assign new_B3719_ = new_B3700_ | new_B3701_;
  assign new_B3720_ = new_B3700_ | new_B3707_;
  assign new_B3721_ = new_B3699_ & new_B3711_;
  assign new_B3722_ = ~new_B3698_ | ~new_B3699_;
  assign new_B3723_ = new_B3707_ & new_B3722_;
  assign new_B3724_ = ~new_B3723_ & ~new_B3707_;
  assign new_B3725_ = new_B3707_ | new_B3722_;
  assign new_B3726_ = ~new_B3700_ | ~new_B3701_;
  assign new_B3727_ = new_B3707_ | new_B3722_;
  assign new_B3728_ = ~new_B3707_ & ~new_B3729_;
  assign new_B3729_ = new_B3707_ & new_B3722_;
  assign new_B3730_ = new_B6180_;
  assign new_B3731_ = new_B6213_;
  assign new_B3732_ = new_B6246_;
  assign new_B3733_ = new_B6279_;
  assign new_B3734_ = new_B6312_;
  assign new_B3735_ = new_B3741_ & new_B3740_;
  assign new_B3736_ = new_B3743_ | new_B3742_;
  assign new_B3737_ = new_B3745_ | new_B3744_;
  assign new_B3738_ = new_B3740_ & new_B3746_;
  assign new_B3739_ = new_B3740_ & new_B3747_;
  assign new_B3740_ = new_B3730_ ^ new_B3731_;
  assign new_B3741_ = new_B3742_ ^ new_B3732_;
  assign new_B3742_ = new_B3750_ & new_B3749_;
  assign new_B3743_ = new_B3748_ & new_B3732_;
  assign new_B3744_ = new_B3753_ & new_B3752_;
  assign new_B3745_ = new_B3751_ & new_B3732_;
  assign new_B3746_ = new_B3754_ | new_B3731_;
  assign new_B3747_ = ~new_B3732_ ^ new_B3744_;
  assign new_B3748_ = ~new_B3757_ | ~new_B3758_;
  assign new_B3749_ = new_B3733_ ^ new_B3740_;
  assign new_B3750_ = new_B3759_ & new_B3752_;
  assign new_B3751_ = ~new_B3761_ | ~new_B3760_;
  assign new_B3752_ = new_B3733_ | new_B3734_;
  assign new_B3753_ = new_B3733_ | new_B3740_;
  assign new_B3754_ = new_B3732_ & new_B3744_;
  assign new_B3755_ = ~new_B3731_ | ~new_B3732_;
  assign new_B3756_ = new_B3740_ & new_B3755_;
  assign new_B3757_ = ~new_B3756_ & ~new_B3740_;
  assign new_B3758_ = new_B3740_ | new_B3755_;
  assign new_B3759_ = ~new_B3733_ | ~new_B3734_;
  assign new_B3760_ = new_B3740_ | new_B3755_;
  assign new_B3761_ = ~new_B3740_ & ~new_B3762_;
  assign new_B3762_ = new_B3740_ & new_B3755_;
  assign new_B3763_ = new_B6345_;
  assign new_B3764_ = new_B6378_;
  assign new_B3765_ = new_B6411_;
  assign new_B3766_ = new_B6444_;
  assign new_B3767_ = new_B6477_;
  assign new_B3768_ = new_B3774_ & new_B3773_;
  assign new_B3769_ = new_B3776_ | new_B3775_;
  assign new_B3770_ = new_B3778_ | new_B3777_;
  assign new_B3771_ = new_B3773_ & new_B3779_;
  assign new_B3772_ = new_B3773_ & new_B3780_;
  assign new_B3773_ = new_B3763_ ^ new_B3764_;
  assign new_B3774_ = new_B3775_ ^ new_B3765_;
  assign new_B3775_ = new_B3783_ & new_B3782_;
  assign new_B3776_ = new_B3781_ & new_B3765_;
  assign new_B3777_ = new_B3786_ & new_B3785_;
  assign new_B3778_ = new_B3784_ & new_B3765_;
  assign new_B3779_ = new_B3787_ | new_B3764_;
  assign new_B3780_ = ~new_B3765_ ^ new_B3777_;
  assign new_B3781_ = ~new_B3790_ | ~new_B3791_;
  assign new_B3782_ = new_B3766_ ^ new_B3773_;
  assign new_B3783_ = new_B3792_ & new_B3785_;
  assign new_B3784_ = ~new_B3794_ | ~new_B3793_;
  assign new_B3785_ = new_B3766_ | new_B3767_;
  assign new_B3786_ = new_B3766_ | new_B3773_;
  assign new_B3787_ = new_B3765_ & new_B3777_;
  assign new_B3788_ = ~new_B3764_ | ~new_B3765_;
  assign new_B3789_ = new_B3773_ & new_B3788_;
  assign new_B3790_ = ~new_B3789_ & ~new_B3773_;
  assign new_B3791_ = new_B3773_ | new_B3788_;
  assign new_B3792_ = ~new_B3766_ | ~new_B3767_;
  assign new_B3793_ = new_B3773_ | new_B3788_;
  assign new_B3794_ = ~new_B3773_ & ~new_B3795_;
  assign new_B3795_ = new_B3773_ & new_B3788_;
  assign new_B3796_ = new_B6510_;
  assign new_B3797_ = new_B6543_;
  assign new_B3798_ = new_B6576_;
  assign new_B3799_ = new_B6609_;
  assign new_B3800_ = new_B6642_;
  assign new_B3801_ = new_B3807_ & new_B3806_;
  assign new_B3802_ = new_B3809_ | new_B3808_;
  assign new_B3803_ = new_B3811_ | new_B3810_;
  assign new_B3804_ = new_B3806_ & new_B3812_;
  assign new_B3805_ = new_B3806_ & new_B3813_;
  assign new_B3806_ = new_B3796_ ^ new_B3797_;
  assign new_B3807_ = new_B3808_ ^ new_B3798_;
  assign new_B3808_ = new_B3816_ & new_B3815_;
  assign new_B3809_ = new_B3814_ & new_B3798_;
  assign new_B3810_ = new_B3819_ & new_B3818_;
  assign new_B3811_ = new_B3817_ & new_B3798_;
  assign new_B3812_ = new_B3820_ | new_B3797_;
  assign new_B3813_ = ~new_B3798_ ^ new_B3810_;
  assign new_B3814_ = ~new_B3823_ | ~new_B3824_;
  assign new_B3815_ = new_B3799_ ^ new_B3806_;
  assign new_B3816_ = new_B3825_ & new_B3818_;
  assign new_B3817_ = ~new_B3827_ | ~new_B3826_;
  assign new_B3818_ = new_B3799_ | new_B3800_;
  assign new_B3819_ = new_B3799_ | new_B3806_;
  assign new_B3820_ = new_B3798_ & new_B3810_;
  assign new_B3821_ = ~new_B3797_ | ~new_B3798_;
  assign new_B3822_ = new_B3806_ & new_B3821_;
  assign new_B3823_ = ~new_B3822_ & ~new_B3806_;
  assign new_B3824_ = new_B3806_ | new_B3821_;
  assign new_B3825_ = ~new_B3799_ | ~new_B3800_;
  assign new_B3826_ = new_B3806_ | new_B3821_;
  assign new_B3827_ = ~new_B3806_ & ~new_B3828_;
  assign new_B3828_ = new_B3806_ & new_B3821_;
  assign new_B3829_ = new_B6675_;
  assign new_B3830_ = new_B6708_;
  assign new_B3831_ = new_B6741_;
  assign new_B3832_ = new_B6774_;
  assign new_B3833_ = new_B6807_;
  assign new_B3834_ = new_B3840_ & new_B3839_;
  assign new_B3835_ = new_B3842_ | new_B3841_;
  assign new_B3836_ = new_B3844_ | new_B3843_;
  assign new_B3837_ = new_B3839_ & new_B3845_;
  assign new_B3838_ = new_B3839_ & new_B3846_;
  assign new_B3839_ = new_B3829_ ^ new_B3830_;
  assign new_B3840_ = new_B3841_ ^ new_B3831_;
  assign new_B3841_ = new_B3849_ & new_B3848_;
  assign new_B3842_ = new_B3847_ & new_B3831_;
  assign new_B3843_ = new_B3852_ & new_B3851_;
  assign new_B3844_ = new_B3850_ & new_B3831_;
  assign new_B3845_ = new_B3853_ | new_B3830_;
  assign new_B3846_ = ~new_B3831_ ^ new_B3843_;
  assign new_B3847_ = ~new_B3856_ | ~new_B3857_;
  assign new_B3848_ = new_B3832_ ^ new_B3839_;
  assign new_B3849_ = new_B3858_ & new_B3851_;
  assign new_B3850_ = ~new_B3860_ | ~new_B3859_;
  assign new_B3851_ = new_B3832_ | new_B3833_;
  assign new_B3852_ = new_B3832_ | new_B3839_;
  assign new_B3853_ = new_B3831_ & new_B3843_;
  assign new_B3854_ = ~new_B3830_ | ~new_B3831_;
  assign new_B3855_ = new_B3839_ & new_B3854_;
  assign new_B3856_ = ~new_B3855_ & ~new_B3839_;
  assign new_B3857_ = new_B3839_ | new_B3854_;
  assign new_B3858_ = ~new_B3832_ | ~new_B3833_;
  assign new_B3859_ = new_B3839_ | new_B3854_;
  assign new_B3860_ = ~new_B3839_ & ~new_B3861_;
  assign new_B3861_ = new_B3839_ & new_B3854_;
  assign new_B3862_ = new_B6840_;
  assign new_B3863_ = new_B6873_;
  assign new_B3864_ = new_B6906_;
  assign new_B3865_ = new_B6939_;
  assign new_B3866_ = new_B6972_;
  assign new_B3867_ = new_B3873_ & new_B3872_;
  assign new_B3868_ = new_B3875_ | new_B3874_;
  assign new_B3869_ = new_B3877_ | new_B3876_;
  assign new_B3870_ = new_B3872_ & new_B3878_;
  assign new_B3871_ = new_B3872_ & new_B3879_;
  assign new_B3872_ = new_B3862_ ^ new_B3863_;
  assign new_B3873_ = new_B3874_ ^ new_B3864_;
  assign new_B3874_ = new_B3882_ & new_B3881_;
  assign new_B3875_ = new_B3880_ & new_B3864_;
  assign new_B3876_ = new_B3885_ & new_B3884_;
  assign new_B3877_ = new_B3883_ & new_B3864_;
  assign new_B3878_ = new_B3886_ | new_B3863_;
  assign new_B3879_ = ~new_B3864_ ^ new_B3876_;
  assign new_B3880_ = ~new_B3889_ | ~new_B3890_;
  assign new_B3881_ = new_B3865_ ^ new_B3872_;
  assign new_B3882_ = new_B3891_ & new_B3884_;
  assign new_B3883_ = ~new_B3893_ | ~new_B3892_;
  assign new_B3884_ = new_B3865_ | new_B3866_;
  assign new_B3885_ = new_B3865_ | new_B3872_;
  assign new_B3886_ = new_B3864_ & new_B3876_;
  assign new_B3887_ = ~new_B3863_ | ~new_B3864_;
  assign new_B3888_ = new_B3872_ & new_B3887_;
  assign new_B3889_ = ~new_B3888_ & ~new_B3872_;
  assign new_B3890_ = new_B3872_ | new_B3887_;
  assign new_B3891_ = ~new_B3865_ | ~new_B3866_;
  assign new_B3892_ = new_B3872_ | new_B3887_;
  assign new_B3893_ = ~new_B3872_ & ~new_B3894_;
  assign new_B3894_ = new_B3872_ & new_B3887_;
  assign new_B3895_ = new_B7005_;
  assign new_B3896_ = new_B7038_;
  assign new_B3897_ = new_B7071_;
  assign new_B3898_ = new_B7104_;
  assign new_B3899_ = new_B7137_;
  assign new_B3900_ = new_B3906_ & new_B3905_;
  assign new_B3901_ = new_B3908_ | new_B3907_;
  assign new_B3902_ = new_B3910_ | new_B3909_;
  assign new_B3903_ = new_B3905_ & new_B3911_;
  assign new_B3904_ = new_B3905_ & new_B3912_;
  assign new_B3905_ = new_B3895_ ^ new_B3896_;
  assign new_B3906_ = new_B3907_ ^ new_B3897_;
  assign new_B3907_ = new_B3915_ & new_B3914_;
  assign new_B3908_ = new_B3913_ & new_B3897_;
  assign new_B3909_ = new_B3918_ & new_B3917_;
  assign new_B3910_ = new_B3916_ & new_B3897_;
  assign new_B3911_ = new_B3919_ | new_B3896_;
  assign new_B3912_ = ~new_B3897_ ^ new_B3909_;
  assign new_B3913_ = ~new_B3922_ | ~new_B3923_;
  assign new_B3914_ = new_B3898_ ^ new_B3905_;
  assign new_B3915_ = new_B3924_ & new_B3917_;
  assign new_B3916_ = ~new_B3926_ | ~new_B3925_;
  assign new_B3917_ = new_B3898_ | new_B3899_;
  assign new_B3918_ = new_B3898_ | new_B3905_;
  assign new_B3919_ = new_B3897_ & new_B3909_;
  assign new_B3920_ = ~new_B3896_ | ~new_B3897_;
  assign new_B3921_ = new_B3905_ & new_B3920_;
  assign new_B3922_ = ~new_B3921_ & ~new_B3905_;
  assign new_B3923_ = new_B3905_ | new_B3920_;
  assign new_B3924_ = ~new_B3898_ | ~new_B3899_;
  assign new_B3925_ = new_B3905_ | new_B3920_;
  assign new_B3926_ = ~new_B3905_ & ~new_B3927_;
  assign new_B3927_ = new_B3905_ & new_B3920_;
  assign new_B3928_ = new_B7170_;
  assign new_B3929_ = new_B7203_;
  assign new_B3930_ = new_B7236_;
  assign new_B3931_ = new_B7269_;
  assign new_B3932_ = new_B7302_;
  assign new_B3933_ = new_B3939_ & new_B3938_;
  assign new_B3934_ = new_B3941_ | new_B3940_;
  assign new_B3935_ = new_B3943_ | new_B3942_;
  assign new_B3936_ = new_B3938_ & new_B3944_;
  assign new_B3937_ = new_B3938_ & new_B3945_;
  assign new_B3938_ = new_B3928_ ^ new_B3929_;
  assign new_B3939_ = new_B3940_ ^ new_B3930_;
  assign new_B3940_ = new_B3948_ & new_B3947_;
  assign new_B3941_ = new_B3946_ & new_B3930_;
  assign new_B3942_ = new_B3951_ & new_B3950_;
  assign new_B3943_ = new_B3949_ & new_B3930_;
  assign new_B3944_ = new_B3952_ | new_B3929_;
  assign new_B3945_ = ~new_B3930_ ^ new_B3942_;
  assign new_B3946_ = ~new_B3955_ | ~new_B3956_;
  assign new_B3947_ = new_B3931_ ^ new_B3938_;
  assign new_B3948_ = new_B3957_ & new_B3950_;
  assign new_B3949_ = ~new_B3959_ | ~new_B3958_;
  assign new_B3950_ = new_B3931_ | new_B3932_;
  assign new_B3951_ = new_B3931_ | new_B3938_;
  assign new_B3952_ = new_B3930_ & new_B3942_;
  assign new_B3953_ = ~new_B3929_ | ~new_B3930_;
  assign new_B3954_ = new_B3938_ & new_B3953_;
  assign new_B3955_ = ~new_B3954_ & ~new_B3938_;
  assign new_B3956_ = new_B3938_ | new_B3953_;
  assign new_B3957_ = ~new_B3931_ | ~new_B3932_;
  assign new_B3958_ = new_B3938_ | new_B3953_;
  assign new_B3959_ = ~new_B3938_ & ~new_B3960_;
  assign new_B3960_ = new_B3938_ & new_B3953_;
  assign new_B3961_ = new_B7335_;
  assign new_B3962_ = new_B7368_;
  assign new_B3963_ = new_B7401_;
  assign new_B3964_ = new_B7434_;
  assign new_B3965_ = new_B7467_;
  assign new_B3966_ = new_B3972_ & new_B3971_;
  assign new_B3967_ = new_B3974_ | new_B3973_;
  assign new_B3968_ = new_B3976_ | new_B3975_;
  assign new_B3969_ = new_B3971_ & new_B3977_;
  assign new_B3970_ = new_B3971_ & new_B3978_;
  assign new_B3971_ = new_B3961_ ^ new_B3962_;
  assign new_B3972_ = new_B3973_ ^ new_B3963_;
  assign new_B3973_ = new_B3981_ & new_B3980_;
  assign new_B3974_ = new_B3979_ & new_B3963_;
  assign new_B3975_ = new_B3984_ & new_B3983_;
  assign new_B3976_ = new_B3982_ & new_B3963_;
  assign new_B3977_ = new_B3985_ | new_B3962_;
  assign new_B3978_ = ~new_B3963_ ^ new_B3975_;
  assign new_B3979_ = ~new_B3988_ | ~new_B3989_;
  assign new_B3980_ = new_B3964_ ^ new_B3971_;
  assign new_B3981_ = new_B3990_ & new_B3983_;
  assign new_B3982_ = ~new_B3992_ | ~new_B3991_;
  assign new_B3983_ = new_B3964_ | new_B3965_;
  assign new_B3984_ = new_B3964_ | new_B3971_;
  assign new_B3985_ = new_B3963_ & new_B3975_;
  assign new_B3986_ = ~new_B3962_ | ~new_B3963_;
  assign new_B3987_ = new_B3971_ & new_B3986_;
  assign new_B3988_ = ~new_B3987_ & ~new_B3971_;
  assign new_B3989_ = new_B3971_ | new_B3986_;
  assign new_B3990_ = ~new_B3964_ | ~new_B3965_;
  assign new_B3991_ = new_B3971_ | new_B3986_;
  assign new_B3992_ = ~new_B3971_ & ~new_B3993_;
  assign new_B3993_ = new_B3971_ & new_B3986_;
  assign new_B3994_ = new_B7500_;
  assign new_B3995_ = new_B7533_;
  assign new_B3996_ = new_B7566_;
  assign new_B3997_ = new_B7599_;
  assign new_B3998_ = new_B7632_;
  assign new_B3999_ = new_B4005_ & new_B4004_;
  assign new_B4000_ = new_B4007_ | new_B4006_;
  assign new_B4001_ = new_B4009_ | new_B4008_;
  assign new_B4002_ = new_B4004_ & new_B4010_;
  assign new_B4003_ = new_B4004_ & new_B4011_;
  assign new_B4004_ = new_B3994_ ^ new_B3995_;
  assign new_B4005_ = new_B4006_ ^ new_B3996_;
  assign new_B4006_ = new_B4014_ & new_B4013_;
  assign new_B4007_ = new_B4012_ & new_B3996_;
  assign new_B4008_ = new_B4017_ & new_B4016_;
  assign new_B4009_ = new_B4015_ & new_B3996_;
  assign new_B4010_ = new_B4018_ | new_B3995_;
  assign new_B4011_ = ~new_B3996_ ^ new_B4008_;
  assign new_B4012_ = ~new_B4021_ | ~new_B4022_;
  assign new_B4013_ = new_B3997_ ^ new_B4004_;
  assign new_B4014_ = new_B4023_ & new_B4016_;
  assign new_B4015_ = ~new_B4025_ | ~new_B4024_;
  assign new_B4016_ = new_B3997_ | new_B3998_;
  assign new_B4017_ = new_B3997_ | new_B4004_;
  assign new_B4018_ = new_B3996_ & new_B4008_;
  assign new_B4019_ = ~new_B3995_ | ~new_B3996_;
  assign new_B4020_ = new_B4004_ & new_B4019_;
  assign new_B4021_ = ~new_B4020_ & ~new_B4004_;
  assign new_B4022_ = new_B4004_ | new_B4019_;
  assign new_B4023_ = ~new_B3997_ | ~new_B3998_;
  assign new_B4024_ = new_B4004_ | new_B4019_;
  assign new_B4025_ = ~new_B4004_ & ~new_B4026_;
  assign new_B4026_ = new_B4004_ & new_B4019_;
  assign new_B4027_ = new_B7665_;
  assign new_B4028_ = new_B7698_;
  assign new_B4029_ = new_B7731_;
  assign new_B4030_ = new_B7764_;
  assign new_B4031_ = new_B7797_;
  assign new_B4032_ = new_B4038_ & new_B4037_;
  assign new_B4033_ = new_B4040_ | new_B4039_;
  assign new_B4034_ = new_B4042_ | new_B4041_;
  assign new_B4035_ = new_B4037_ & new_B4043_;
  assign new_B4036_ = new_B4037_ & new_B4044_;
  assign new_B4037_ = new_B4027_ ^ new_B4028_;
  assign new_B4038_ = new_B4039_ ^ new_B4029_;
  assign new_B4039_ = new_B4047_ & new_B4046_;
  assign new_B4040_ = new_B4045_ & new_B4029_;
  assign new_B4041_ = new_B4050_ & new_B4049_;
  assign new_B4042_ = new_B4048_ & new_B4029_;
  assign new_B4043_ = new_B4051_ | new_B4028_;
  assign new_B4044_ = ~new_B4029_ ^ new_B4041_;
  assign new_B4045_ = ~new_B4054_ | ~new_B4055_;
  assign new_B4046_ = new_B4030_ ^ new_B4037_;
  assign new_B4047_ = new_B4056_ & new_B4049_;
  assign new_B4048_ = ~new_B4058_ | ~new_B4057_;
  assign new_B4049_ = new_B4030_ | new_B4031_;
  assign new_B4050_ = new_B4030_ | new_B4037_;
  assign new_B4051_ = new_B4029_ & new_B4041_;
  assign new_B4052_ = ~new_B4028_ | ~new_B4029_;
  assign new_B4053_ = new_B4037_ & new_B4052_;
  assign new_B4054_ = ~new_B4053_ & ~new_B4037_;
  assign new_B4055_ = new_B4037_ | new_B4052_;
  assign new_B4056_ = ~new_B4030_ | ~new_B4031_;
  assign new_B4057_ = new_B4037_ | new_B4052_;
  assign new_B4058_ = ~new_B4037_ & ~new_B4059_;
  assign new_B4059_ = new_B4037_ & new_B4052_;
  assign new_B4060_ = new_B7830_;
  assign new_B4061_ = new_B7863_;
  assign new_B4062_ = new_B7896_;
  assign new_B4063_ = new_B7929_;
  assign new_B4064_ = new_B7962_;
  assign new_B4065_ = new_B4071_ & new_B4070_;
  assign new_B4066_ = new_B4073_ | new_B4072_;
  assign new_B4067_ = new_B4075_ | new_B4074_;
  assign new_B4068_ = new_B4070_ & new_B4076_;
  assign new_B4069_ = new_B4070_ & new_B4077_;
  assign new_B4070_ = new_B4060_ ^ new_B4061_;
  assign new_B4071_ = new_B4072_ ^ new_B4062_;
  assign new_B4072_ = new_B4080_ & new_B4079_;
  assign new_B4073_ = new_B4078_ & new_B4062_;
  assign new_B4074_ = new_B4083_ & new_B4082_;
  assign new_B4075_ = new_B4081_ & new_B4062_;
  assign new_B4076_ = new_B4084_ | new_B4061_;
  assign new_B4077_ = ~new_B4062_ ^ new_B4074_;
  assign new_B4078_ = ~new_B4087_ | ~new_B4088_;
  assign new_B4079_ = new_B4063_ ^ new_B4070_;
  assign new_B4080_ = new_B4089_ & new_B4082_;
  assign new_B4081_ = ~new_B4091_ | ~new_B4090_;
  assign new_B4082_ = new_B4063_ | new_B4064_;
  assign new_B4083_ = new_B4063_ | new_B4070_;
  assign new_B4084_ = new_B4062_ & new_B4074_;
  assign new_B4085_ = ~new_B4061_ | ~new_B4062_;
  assign new_B4086_ = new_B4070_ & new_B4085_;
  assign new_B4087_ = ~new_B4086_ & ~new_B4070_;
  assign new_B4088_ = new_B4070_ | new_B4085_;
  assign new_B4089_ = ~new_B4063_ | ~new_B4064_;
  assign new_B4090_ = new_B4070_ | new_B4085_;
  assign new_B4091_ = ~new_B4070_ & ~new_B4092_;
  assign new_B4092_ = new_B4070_ & new_B4085_;
  assign new_B4093_ = new_B7995_;
  assign new_B4094_ = new_B8028_;
  assign new_B4095_ = new_B8061_;
  assign new_B4096_ = new_B8094_;
  assign new_B4097_ = new_B8127_;
  assign new_B4098_ = new_B4104_ & new_B4103_;
  assign new_B4099_ = new_B4106_ | new_B4105_;
  assign new_B4100_ = new_B4108_ | new_B4107_;
  assign new_B4101_ = new_B4103_ & new_B4109_;
  assign new_B4102_ = new_B4103_ & new_B4110_;
  assign new_B4103_ = new_B4093_ ^ new_B4094_;
  assign new_B4104_ = new_B4105_ ^ new_B4095_;
  assign new_B4105_ = new_B4113_ & new_B4112_;
  assign new_B4106_ = new_B4111_ & new_B4095_;
  assign new_B4107_ = new_B4116_ & new_B4115_;
  assign new_B4108_ = new_B4114_ & new_B4095_;
  assign new_B4109_ = new_B4117_ | new_B4094_;
  assign new_B4110_ = ~new_B4095_ ^ new_B4107_;
  assign new_B4111_ = ~new_B4120_ | ~new_B4121_;
  assign new_B4112_ = new_B4096_ ^ new_B4103_;
  assign new_B4113_ = new_B4122_ & new_B4115_;
  assign new_B4114_ = ~new_B4124_ | ~new_B4123_;
  assign new_B4115_ = new_B4096_ | new_B4097_;
  assign new_B4116_ = new_B4096_ | new_B4103_;
  assign new_B4117_ = new_B4095_ & new_B4107_;
  assign new_B4118_ = ~new_B4094_ | ~new_B4095_;
  assign new_B4119_ = new_B4103_ & new_B4118_;
  assign new_B4120_ = ~new_B4119_ & ~new_B4103_;
  assign new_B4121_ = new_B4103_ | new_B4118_;
  assign new_B4122_ = ~new_B4096_ | ~new_B4097_;
  assign new_B4123_ = new_B4103_ | new_B4118_;
  assign new_B4124_ = ~new_B4103_ & ~new_B4125_;
  assign new_B4125_ = new_B4103_ & new_B4118_;
  assign new_B4126_ = new_B8160_;
  assign new_B4127_ = new_B8193_;
  assign new_B4128_ = new_B8226_;
  assign new_B4129_ = new_B8259_;
  assign new_B4130_ = new_B8292_;
  assign new_B4131_ = new_B4137_ & new_B4136_;
  assign new_B4132_ = new_B4139_ | new_B4138_;
  assign new_B4133_ = new_B4141_ | new_B4140_;
  assign new_B4134_ = new_B4136_ & new_B4142_;
  assign new_B4135_ = new_B4136_ & new_B4143_;
  assign new_B4136_ = new_B4126_ ^ new_B4127_;
  assign new_B4137_ = new_B4138_ ^ new_B4128_;
  assign new_B4138_ = new_B4146_ & new_B4145_;
  assign new_B4139_ = new_B4144_ & new_B4128_;
  assign new_B4140_ = new_B4149_ & new_B4148_;
  assign new_B4141_ = new_B4147_ & new_B4128_;
  assign new_B4142_ = new_B4150_ | new_B4127_;
  assign new_B4143_ = ~new_B4128_ ^ new_B4140_;
  assign new_B4144_ = ~new_B4153_ | ~new_B4154_;
  assign new_B4145_ = new_B4129_ ^ new_B4136_;
  assign new_B4146_ = new_B4155_ & new_B4148_;
  assign new_B4147_ = ~new_B4157_ | ~new_B4156_;
  assign new_B4148_ = new_B4129_ | new_B4130_;
  assign new_B4149_ = new_B4129_ | new_B4136_;
  assign new_B4150_ = new_B4128_ & new_B4140_;
  assign new_B4151_ = ~new_B4127_ | ~new_B4128_;
  assign new_B4152_ = new_B4136_ & new_B4151_;
  assign new_B4153_ = ~new_B4152_ & ~new_B4136_;
  assign new_B4154_ = new_B4136_ | new_B4151_;
  assign new_B4155_ = ~new_B4129_ | ~new_B4130_;
  assign new_B4156_ = new_B4136_ | new_B4151_;
  assign new_B4157_ = ~new_B4136_ & ~new_B4158_;
  assign new_B4158_ = new_B4136_ & new_B4151_;
  assign new_B4159_ = new_B8325_;
  assign new_B4160_ = new_B8358_;
  assign new_B4161_ = new_B8391_;
  assign new_B4162_ = new_B8424_;
  assign new_B4163_ = new_B8457_;
  assign new_B4164_ = new_B4170_ & new_B4169_;
  assign new_B4165_ = new_B4172_ | new_B4171_;
  assign new_B4166_ = new_B4174_ | new_B4173_;
  assign new_B4167_ = new_B4169_ & new_B4175_;
  assign new_B4168_ = new_B4169_ & new_B4176_;
  assign new_B4169_ = new_B4159_ ^ new_B4160_;
  assign new_B4170_ = new_B4171_ ^ new_B4161_;
  assign new_B4171_ = new_B4179_ & new_B4178_;
  assign new_B4172_ = new_B4177_ & new_B4161_;
  assign new_B4173_ = new_B4182_ & new_B4181_;
  assign new_B4174_ = new_B4180_ & new_B4161_;
  assign new_B4175_ = new_B4183_ | new_B4160_;
  assign new_B4176_ = ~new_B4161_ ^ new_B4173_;
  assign new_B4177_ = ~new_B4186_ | ~new_B4187_;
  assign new_B4178_ = new_B4162_ ^ new_B4169_;
  assign new_B4179_ = new_B4188_ & new_B4181_;
  assign new_B4180_ = ~new_B4190_ | ~new_B4189_;
  assign new_B4181_ = new_B4162_ | new_B4163_;
  assign new_B4182_ = new_B4162_ | new_B4169_;
  assign new_B4183_ = new_B4161_ & new_B4173_;
  assign new_B4184_ = ~new_B4160_ | ~new_B4161_;
  assign new_B4185_ = new_B4169_ & new_B4184_;
  assign new_B4186_ = ~new_B4185_ & ~new_B4169_;
  assign new_B4187_ = new_B4169_ | new_B4184_;
  assign new_B4188_ = ~new_B4162_ | ~new_B4163_;
  assign new_B4189_ = new_B4169_ | new_B4184_;
  assign new_B4190_ = ~new_B4169_ & ~new_B4191_;
  assign new_B4191_ = new_B4169_ & new_B4184_;
  assign new_B4192_ = new_B8490_;
  assign new_B4193_ = new_B8523_;
  assign new_B4194_ = new_B8556_;
  assign new_B4195_ = new_B8589_;
  assign new_B4196_ = new_B8622_;
  assign new_B4197_ = new_B4203_ & new_B4202_;
  assign new_B4198_ = new_B4205_ | new_B4204_;
  assign new_B4199_ = new_B4207_ | new_B4206_;
  assign new_B4200_ = new_B4202_ & new_B4208_;
  assign new_B4201_ = new_B4202_ & new_B4209_;
  assign new_B4202_ = new_B4192_ ^ new_B4193_;
  assign new_B4203_ = new_B4204_ ^ new_B4194_;
  assign new_B4204_ = new_B4212_ & new_B4211_;
  assign new_B4205_ = new_B4210_ & new_B4194_;
  assign new_B4206_ = new_B4215_ & new_B4214_;
  assign new_B4207_ = new_B4213_ & new_B4194_;
  assign new_B4208_ = new_B4216_ | new_B4193_;
  assign new_B4209_ = ~new_B4194_ ^ new_B4206_;
  assign new_B4210_ = ~new_B4219_ | ~new_B4220_;
  assign new_B4211_ = new_B4195_ ^ new_B4202_;
  assign new_B4212_ = new_B4221_ & new_B4214_;
  assign new_B4213_ = ~new_B4223_ | ~new_B4222_;
  assign new_B4214_ = new_B4195_ | new_B4196_;
  assign new_B4215_ = new_B4195_ | new_B4202_;
  assign new_B4216_ = new_B4194_ & new_B4206_;
  assign new_B4217_ = ~new_B4193_ | ~new_B4194_;
  assign new_B4218_ = new_B4202_ & new_B4217_;
  assign new_B4219_ = ~new_B4218_ & ~new_B4202_;
  assign new_B4220_ = new_B4202_ | new_B4217_;
  assign new_B4221_ = ~new_B4195_ | ~new_B4196_;
  assign new_B4222_ = new_B4202_ | new_B4217_;
  assign new_B4223_ = ~new_B4202_ & ~new_B4224_;
  assign new_B4224_ = new_B4202_ & new_B4217_;
  assign new_B4225_ = new_B8655_;
  assign new_B4226_ = new_B8688_;
  assign new_B4227_ = new_B8721_;
  assign new_B4228_ = new_B8754_;
  assign new_B4229_ = new_B8787_;
  assign new_B4230_ = new_B4236_ & new_B4235_;
  assign new_B4231_ = new_B4238_ | new_B4237_;
  assign new_B4232_ = new_B4240_ | new_B4239_;
  assign new_B4233_ = new_B4235_ & new_B4241_;
  assign new_B4234_ = new_B4235_ & new_B4242_;
  assign new_B4235_ = new_B4225_ ^ new_B4226_;
  assign new_B4236_ = new_B4237_ ^ new_B4227_;
  assign new_B4237_ = new_B4245_ & new_B4244_;
  assign new_B4238_ = new_B4243_ & new_B4227_;
  assign new_B4239_ = new_B4248_ & new_B4247_;
  assign new_B4240_ = new_B4246_ & new_B4227_;
  assign new_B4241_ = new_B4249_ | new_B4226_;
  assign new_B4242_ = ~new_B4227_ ^ new_B4239_;
  assign new_B4243_ = ~new_B4252_ | ~new_B4253_;
  assign new_B4244_ = new_B4228_ ^ new_B4235_;
  assign new_B4245_ = new_B4254_ & new_B4247_;
  assign new_B4246_ = ~new_B4256_ | ~new_B4255_;
  assign new_B4247_ = new_B4228_ | new_B4229_;
  assign new_B4248_ = new_B4228_ | new_B4235_;
  assign new_B4249_ = new_B4227_ & new_B4239_;
  assign new_B4250_ = ~new_B4226_ | ~new_B4227_;
  assign new_B4251_ = new_B4235_ & new_B4250_;
  assign new_B4252_ = ~new_B4251_ & ~new_B4235_;
  assign new_B4253_ = new_B4235_ | new_B4250_;
  assign new_B4254_ = ~new_B4228_ | ~new_B4229_;
  assign new_B4255_ = new_B4235_ | new_B4250_;
  assign new_B4256_ = ~new_B4235_ & ~new_B4257_;
  assign new_B4257_ = new_B4235_ & new_B4250_;
  assign new_B4258_ = new_B8820_;
  assign new_B4259_ = new_B8853_;
  assign new_B4260_ = new_B8886_;
  assign new_B4261_ = new_B8919_;
  assign new_B4262_ = new_B8952_;
  assign new_B4263_ = new_B4269_ & new_B4268_;
  assign new_B4264_ = new_B4271_ | new_B4270_;
  assign new_B4265_ = new_B4273_ | new_B4272_;
  assign new_B4266_ = new_B4268_ & new_B4274_;
  assign new_B4267_ = new_B4268_ & new_B4275_;
  assign new_B4268_ = new_B4258_ ^ new_B4259_;
  assign new_B4269_ = new_B4270_ ^ new_B4260_;
  assign new_B4270_ = new_B4278_ & new_B4277_;
  assign new_B4271_ = new_B4276_ & new_B4260_;
  assign new_B4272_ = new_B4281_ & new_B4280_;
  assign new_B4273_ = new_B4279_ & new_B4260_;
  assign new_B4274_ = new_B4282_ | new_B4259_;
  assign new_B4275_ = ~new_B4260_ ^ new_B4272_;
  assign new_B4276_ = ~new_B4285_ | ~new_B4286_;
  assign new_B4277_ = new_B4261_ ^ new_B4268_;
  assign new_B4278_ = new_B4287_ & new_B4280_;
  assign new_B4279_ = ~new_B4289_ | ~new_B4288_;
  assign new_B4280_ = new_B4261_ | new_B4262_;
  assign new_B4281_ = new_B4261_ | new_B4268_;
  assign new_B4282_ = new_B4260_ & new_B4272_;
  assign new_B4283_ = ~new_B4259_ | ~new_B4260_;
  assign new_B4284_ = new_B4268_ & new_B4283_;
  assign new_B4285_ = ~new_B4284_ & ~new_B4268_;
  assign new_B4286_ = new_B4268_ | new_B4283_;
  assign new_B4287_ = ~new_B4261_ | ~new_B4262_;
  assign new_B4288_ = new_B4268_ | new_B4283_;
  assign new_B4289_ = ~new_B4268_ & ~new_B4290_;
  assign new_B4290_ = new_B4268_ & new_B4283_;
  assign new_B4291_ = new_B8985_;
  assign new_B4292_ = new_B9018_;
  assign new_B4293_ = new_B9051_;
  assign new_B4294_ = new_B9084_;
  assign new_B4295_ = new_B9117_;
  assign new_B4296_ = new_B4302_ & new_B4301_;
  assign new_B4297_ = new_B4304_ | new_B4303_;
  assign new_B4298_ = new_B4306_ | new_B4305_;
  assign new_B4299_ = new_B4301_ & new_B4307_;
  assign new_B4300_ = new_B4301_ & new_B4308_;
  assign new_B4301_ = new_B4291_ ^ new_B4292_;
  assign new_B4302_ = new_B4303_ ^ new_B4293_;
  assign new_B4303_ = new_B4311_ & new_B4310_;
  assign new_B4304_ = new_B4309_ & new_B4293_;
  assign new_B4305_ = new_B4314_ & new_B4313_;
  assign new_B4306_ = new_B4312_ & new_B4293_;
  assign new_B4307_ = new_B4315_ | new_B4292_;
  assign new_B4308_ = ~new_B4293_ ^ new_B4305_;
  assign new_B4309_ = ~new_B4318_ | ~new_B4319_;
  assign new_B4310_ = new_B4294_ ^ new_B4301_;
  assign new_B4311_ = new_B4320_ & new_B4313_;
  assign new_B4312_ = ~new_B4322_ | ~new_B4321_;
  assign new_B4313_ = new_B4294_ | new_B4295_;
  assign new_B4314_ = new_B4294_ | new_B4301_;
  assign new_B4315_ = new_B4293_ & new_B4305_;
  assign new_B4316_ = ~new_B4292_ | ~new_B4293_;
  assign new_B4317_ = new_B4301_ & new_B4316_;
  assign new_B4318_ = ~new_B4317_ & ~new_B4301_;
  assign new_B4319_ = new_B4301_ | new_B4316_;
  assign new_B4320_ = ~new_B4294_ | ~new_B4295_;
  assign new_B4321_ = new_B4301_ | new_B4316_;
  assign new_B4322_ = ~new_B4301_ & ~new_B4323_;
  assign new_B4323_ = new_B4301_ & new_B4316_;
  assign new_B4324_ = new_B9150_;
  assign new_B4325_ = new_B9183_;
  assign new_B4326_ = new_B9216_;
  assign new_B4327_ = new_B9249_;
  assign new_B4328_ = new_B9282_;
  assign new_B4329_ = new_B4335_ & new_B4334_;
  assign new_B4330_ = new_B4337_ | new_B4336_;
  assign new_B4331_ = new_B4339_ | new_B4338_;
  assign new_B4332_ = new_B4334_ & new_B4340_;
  assign new_B4333_ = new_B4334_ & new_B4341_;
  assign new_B4334_ = new_B4324_ ^ new_B4325_;
  assign new_B4335_ = new_B4336_ ^ new_B4326_;
  assign new_B4336_ = new_B4344_ & new_B4343_;
  assign new_B4337_ = new_B4342_ & new_B4326_;
  assign new_B4338_ = new_B4347_ & new_B4346_;
  assign new_B4339_ = new_B4345_ & new_B4326_;
  assign new_B4340_ = new_B4348_ | new_B4325_;
  assign new_B4341_ = ~new_B4326_ ^ new_B4338_;
  assign new_B4342_ = ~new_B4351_ | ~new_B4352_;
  assign new_B4343_ = new_B4327_ ^ new_B4334_;
  assign new_B4344_ = new_B4353_ & new_B4346_;
  assign new_B4345_ = ~new_B4355_ | ~new_B4354_;
  assign new_B4346_ = new_B4327_ | new_B4328_;
  assign new_B4347_ = new_B4327_ | new_B4334_;
  assign new_B4348_ = new_B4326_ & new_B4338_;
  assign new_B4349_ = ~new_B4325_ | ~new_B4326_;
  assign new_B4350_ = new_B4334_ & new_B4349_;
  assign new_B4351_ = ~new_B4350_ & ~new_B4334_;
  assign new_B4352_ = new_B4334_ | new_B4349_;
  assign new_B4353_ = ~new_B4327_ | ~new_B4328_;
  assign new_B4354_ = new_B4334_ | new_B4349_;
  assign new_B4355_ = ~new_B4334_ & ~new_B4356_;
  assign new_B4356_ = new_B4334_ & new_B4349_;
  assign new_B4357_ = new_B5187_;
  assign new_B4358_ = new_B5224_;
  assign new_B4359_ = new_B5257_;
  assign new_B4360_ = new_B5290_;
  assign new_B4361_ = new_B5323_;
  assign new_B4362_ = new_B4368_ & new_B4367_;
  assign new_B4363_ = new_B4370_ | new_B4369_;
  assign new_B4364_ = new_B4372_ | new_B4371_;
  assign new_B4365_ = new_B4367_ & new_B4373_;
  assign new_B4366_ = new_B4367_ & new_B4374_;
  assign new_B4367_ = new_B4357_ ^ new_B4358_;
  assign new_B4368_ = new_B4369_ ^ new_B4359_;
  assign new_B4369_ = new_B4377_ & new_B4376_;
  assign new_B4370_ = new_B4375_ & new_B4359_;
  assign new_B4371_ = new_B4380_ & new_B4379_;
  assign new_B4372_ = new_B4378_ & new_B4359_;
  assign new_B4373_ = new_B4381_ | new_B4358_;
  assign new_B4374_ = ~new_B4359_ ^ new_B4371_;
  assign new_B4375_ = ~new_B4384_ | ~new_B4385_;
  assign new_B4376_ = new_B4360_ ^ new_B4367_;
  assign new_B4377_ = new_B4386_ & new_B4379_;
  assign new_B4378_ = ~new_B4388_ | ~new_B4387_;
  assign new_B4379_ = new_B4360_ | new_B4361_;
  assign new_B4380_ = new_B4360_ | new_B4367_;
  assign new_B4381_ = new_B4359_ & new_B4371_;
  assign new_B4382_ = ~new_B4358_ | ~new_B4359_;
  assign new_B4383_ = new_B4367_ & new_B4382_;
  assign new_B4384_ = ~new_B4383_ & ~new_B4367_;
  assign new_B4385_ = new_B4367_ | new_B4382_;
  assign new_B4386_ = ~new_B4360_ | ~new_B4361_;
  assign new_B4387_ = new_B4367_ | new_B4382_;
  assign new_B4388_ = ~new_B4367_ & ~new_B4389_;
  assign new_B4389_ = new_B4367_ & new_B4382_;
  assign new_B4390_ = new_B5356_;
  assign new_B4391_ = new_B5389_;
  assign new_B4392_ = new_B5422_;
  assign new_B4393_ = new_B5455_;
  assign new_B4394_ = new_B5488_;
  assign new_B4395_ = new_B4401_ & new_B4400_;
  assign new_B4396_ = new_B4403_ | new_B4402_;
  assign new_B4397_ = new_B4405_ | new_B4404_;
  assign new_B4398_ = new_B4400_ & new_B4406_;
  assign new_B4399_ = new_B4400_ & new_B4407_;
  assign new_B4400_ = new_B4390_ ^ new_B4391_;
  assign new_B4401_ = new_B4402_ ^ new_B4392_;
  assign new_B4402_ = new_B4410_ & new_B4409_;
  assign new_B4403_ = new_B4408_ & new_B4392_;
  assign new_B4404_ = new_B4413_ & new_B4412_;
  assign new_B4405_ = new_B4411_ & new_B4392_;
  assign new_B4406_ = new_B4414_ | new_B4391_;
  assign new_B4407_ = ~new_B4392_ ^ new_B4404_;
  assign new_B4408_ = ~new_B4417_ | ~new_B4418_;
  assign new_B4409_ = new_B4393_ ^ new_B4400_;
  assign new_B4410_ = new_B4419_ & new_B4412_;
  assign new_B4411_ = ~new_B4421_ | ~new_B4420_;
  assign new_B4412_ = new_B4393_ | new_B4394_;
  assign new_B4413_ = new_B4393_ | new_B4400_;
  assign new_B4414_ = new_B4392_ & new_B4404_;
  assign new_B4415_ = ~new_B4391_ | ~new_B4392_;
  assign new_B4416_ = new_B4400_ & new_B4415_;
  assign new_B4417_ = ~new_B4416_ & ~new_B4400_;
  assign new_B4418_ = new_B4400_ | new_B4415_;
  assign new_B4419_ = ~new_B4393_ | ~new_B4394_;
  assign new_B4420_ = new_B4400_ | new_B4415_;
  assign new_B4421_ = ~new_B4400_ & ~new_B4422_;
  assign new_B4422_ = new_B4400_ & new_B4415_;
  assign new_B4423_ = new_B5521_;
  assign new_B4424_ = new_B5554_;
  assign new_B4425_ = new_B5587_;
  assign new_B4426_ = new_B5620_;
  assign new_B4427_ = new_B5653_;
  assign new_B4428_ = new_B4434_ & new_B4433_;
  assign new_B4429_ = new_B4436_ | new_B4435_;
  assign new_B4430_ = new_B4438_ | new_B4437_;
  assign new_B4431_ = new_B4433_ & new_B4439_;
  assign new_B4432_ = new_B4433_ & new_B4440_;
  assign new_B4433_ = new_B4423_ ^ new_B4424_;
  assign new_B4434_ = new_B4435_ ^ new_B4425_;
  assign new_B4435_ = new_B4443_ & new_B4442_;
  assign new_B4436_ = new_B4441_ & new_B4425_;
  assign new_B4437_ = new_B4446_ & new_B4445_;
  assign new_B4438_ = new_B4444_ & new_B4425_;
  assign new_B4439_ = new_B4447_ | new_B4424_;
  assign new_B4440_ = ~new_B4425_ ^ new_B4437_;
  assign new_B4441_ = ~new_B4450_ | ~new_B4451_;
  assign new_B4442_ = new_B4426_ ^ new_B4433_;
  assign new_B4443_ = new_B4452_ & new_B4445_;
  assign new_B4444_ = ~new_B4454_ | ~new_B4453_;
  assign new_B4445_ = new_B4426_ | new_B4427_;
  assign new_B4446_ = new_B4426_ | new_B4433_;
  assign new_B4447_ = new_B4425_ & new_B4437_;
  assign new_B4448_ = ~new_B4424_ | ~new_B4425_;
  assign new_B4449_ = new_B4433_ & new_B4448_;
  assign new_B4450_ = ~new_B4449_ & ~new_B4433_;
  assign new_B4451_ = new_B4433_ | new_B4448_;
  assign new_B4452_ = ~new_B4426_ | ~new_B4427_;
  assign new_B4453_ = new_B4433_ | new_B4448_;
  assign new_B4454_ = ~new_B4433_ & ~new_B4455_;
  assign new_B4455_ = new_B4433_ & new_B4448_;
  assign new_B4456_ = new_B5686_;
  assign new_B4457_ = new_B5719_;
  assign new_B4458_ = new_B5752_;
  assign new_B4459_ = new_B5785_;
  assign new_B4460_ = new_B5818_;
  assign new_B4461_ = new_B4467_ & new_B4466_;
  assign new_B4462_ = new_B4469_ | new_B4468_;
  assign new_B4463_ = new_B4471_ | new_B4470_;
  assign new_B4464_ = new_B4466_ & new_B4472_;
  assign new_B4465_ = new_B4466_ & new_B4473_;
  assign new_B4466_ = new_B4456_ ^ new_B4457_;
  assign new_B4467_ = new_B4468_ ^ new_B4458_;
  assign new_B4468_ = new_B4476_ & new_B4475_;
  assign new_B4469_ = new_B4474_ & new_B4458_;
  assign new_B4470_ = new_B4479_ & new_B4478_;
  assign new_B4471_ = new_B4477_ & new_B4458_;
  assign new_B4472_ = new_B4480_ | new_B4457_;
  assign new_B4473_ = ~new_B4458_ ^ new_B4470_;
  assign new_B4474_ = ~new_B4483_ | ~new_B4484_;
  assign new_B4475_ = new_B4459_ ^ new_B4466_;
  assign new_B4476_ = new_B4485_ & new_B4478_;
  assign new_B4477_ = ~new_B4487_ | ~new_B4486_;
  assign new_B4478_ = new_B4459_ | new_B4460_;
  assign new_B4479_ = new_B4459_ | new_B4466_;
  assign new_B4480_ = new_B4458_ & new_B4470_;
  assign new_B4481_ = ~new_B4457_ | ~new_B4458_;
  assign new_B4482_ = new_B4466_ & new_B4481_;
  assign new_B4483_ = ~new_B4482_ & ~new_B4466_;
  assign new_B4484_ = new_B4466_ | new_B4481_;
  assign new_B4485_ = ~new_B4459_ | ~new_B4460_;
  assign new_B4486_ = new_B4466_ | new_B4481_;
  assign new_B4487_ = ~new_B4466_ & ~new_B4488_;
  assign new_B4488_ = new_B4466_ & new_B4481_;
  assign new_B4489_ = new_B5851_;
  assign new_B4490_ = new_B5884_;
  assign new_B4491_ = new_B5917_;
  assign new_B4492_ = new_B5950_;
  assign new_B4493_ = new_B5983_;
  assign new_B4494_ = new_B4500_ & new_B4499_;
  assign new_B4495_ = new_B4502_ | new_B4501_;
  assign new_B4496_ = new_B4504_ | new_B4503_;
  assign new_B4497_ = new_B4499_ & new_B4505_;
  assign new_B4498_ = new_B4499_ & new_B4506_;
  assign new_B4499_ = new_B4489_ ^ new_B4490_;
  assign new_B4500_ = new_B4501_ ^ new_B4491_;
  assign new_B4501_ = new_B4509_ & new_B4508_;
  assign new_B4502_ = new_B4507_ & new_B4491_;
  assign new_B4503_ = new_B4512_ & new_B4511_;
  assign new_B4504_ = new_B4510_ & new_B4491_;
  assign new_B4505_ = new_B4513_ | new_B4490_;
  assign new_B4506_ = ~new_B4491_ ^ new_B4503_;
  assign new_B4507_ = ~new_B4516_ | ~new_B4517_;
  assign new_B4508_ = new_B4492_ ^ new_B4499_;
  assign new_B4509_ = new_B4518_ & new_B4511_;
  assign new_B4510_ = ~new_B4520_ | ~new_B4519_;
  assign new_B4511_ = new_B4492_ | new_B4493_;
  assign new_B4512_ = new_B4492_ | new_B4499_;
  assign new_B4513_ = new_B4491_ & new_B4503_;
  assign new_B4514_ = ~new_B4490_ | ~new_B4491_;
  assign new_B4515_ = new_B4499_ & new_B4514_;
  assign new_B4516_ = ~new_B4515_ & ~new_B4499_;
  assign new_B4517_ = new_B4499_ | new_B4514_;
  assign new_B4518_ = ~new_B4492_ | ~new_B4493_;
  assign new_B4519_ = new_B4499_ | new_B4514_;
  assign new_B4520_ = ~new_B4499_ & ~new_B4521_;
  assign new_B4521_ = new_B4499_ & new_B4514_;
  assign new_B4522_ = new_B6016_;
  assign new_B4523_ = new_B6049_;
  assign new_B4524_ = new_B6082_;
  assign new_B4525_ = new_B6115_;
  assign new_B4526_ = new_B6148_;
  assign new_B4527_ = new_B4533_ & new_B4532_;
  assign new_B4528_ = new_B4535_ | new_B4534_;
  assign new_B4529_ = new_B4537_ | new_B4536_;
  assign new_B4530_ = new_B4532_ & new_B4538_;
  assign new_B4531_ = new_B4532_ & new_B4539_;
  assign new_B4532_ = new_B4522_ ^ new_B4523_;
  assign new_B4533_ = new_B4534_ ^ new_B4524_;
  assign new_B4534_ = new_B4542_ & new_B4541_;
  assign new_B4535_ = new_B4540_ & new_B4524_;
  assign new_B4536_ = new_B4545_ & new_B4544_;
  assign new_B4537_ = new_B4543_ & new_B4524_;
  assign new_B4538_ = new_B4546_ | new_B4523_;
  assign new_B4539_ = ~new_B4524_ ^ new_B4536_;
  assign new_B4540_ = ~new_B4549_ | ~new_B4550_;
  assign new_B4541_ = new_B4525_ ^ new_B4532_;
  assign new_B4542_ = new_B4551_ & new_B4544_;
  assign new_B4543_ = ~new_B4553_ | ~new_B4552_;
  assign new_B4544_ = new_B4525_ | new_B4526_;
  assign new_B4545_ = new_B4525_ | new_B4532_;
  assign new_B4546_ = new_B4524_ & new_B4536_;
  assign new_B4547_ = ~new_B4523_ | ~new_B4524_;
  assign new_B4548_ = new_B4532_ & new_B4547_;
  assign new_B4549_ = ~new_B4548_ & ~new_B4532_;
  assign new_B4550_ = new_B4532_ | new_B4547_;
  assign new_B4551_ = ~new_B4525_ | ~new_B4526_;
  assign new_B4552_ = new_B4532_ | new_B4547_;
  assign new_B4553_ = ~new_B4532_ & ~new_B4554_;
  assign new_B4554_ = new_B4532_ & new_B4547_;
  assign new_B4555_ = new_B6181_;
  assign new_B4556_ = new_B6214_;
  assign new_B4557_ = new_B6247_;
  assign new_B4558_ = new_B6280_;
  assign new_B4559_ = new_B6313_;
  assign new_B4560_ = new_B4566_ & new_B4565_;
  assign new_B4561_ = new_B4568_ | new_B4567_;
  assign new_B4562_ = new_B4570_ | new_B4569_;
  assign new_B4563_ = new_B4565_ & new_B4571_;
  assign new_B4564_ = new_B4565_ & new_B4572_;
  assign new_B4565_ = new_B4555_ ^ new_B4556_;
  assign new_B4566_ = new_B4567_ ^ new_B4557_;
  assign new_B4567_ = new_B4575_ & new_B4574_;
  assign new_B4568_ = new_B4573_ & new_B4557_;
  assign new_B4569_ = new_B4578_ & new_B4577_;
  assign new_B4570_ = new_B4576_ & new_B4557_;
  assign new_B4571_ = new_B4579_ | new_B4556_;
  assign new_B4572_ = ~new_B4557_ ^ new_B4569_;
  assign new_B4573_ = ~new_B4582_ | ~new_B4583_;
  assign new_B4574_ = new_B4558_ ^ new_B4565_;
  assign new_B4575_ = new_B4584_ & new_B4577_;
  assign new_B4576_ = ~new_B4586_ | ~new_B4585_;
  assign new_B4577_ = new_B4558_ | new_B4559_;
  assign new_B4578_ = new_B4558_ | new_B4565_;
  assign new_B4579_ = new_B4557_ & new_B4569_;
  assign new_B4580_ = ~new_B4556_ | ~new_B4557_;
  assign new_B4581_ = new_B4565_ & new_B4580_;
  assign new_B4582_ = ~new_B4581_ & ~new_B4565_;
  assign new_B4583_ = new_B4565_ | new_B4580_;
  assign new_B4584_ = ~new_B4558_ | ~new_B4559_;
  assign new_B4585_ = new_B4565_ | new_B4580_;
  assign new_B4586_ = ~new_B4565_ & ~new_B4587_;
  assign new_B4587_ = new_B4565_ & new_B4580_;
  assign new_B4588_ = new_B6346_;
  assign new_B4589_ = new_B6379_;
  assign new_B4590_ = new_B6412_;
  assign new_B4591_ = new_B6445_;
  assign new_B4592_ = new_B6478_;
  assign new_B4593_ = new_B4599_ & new_B4598_;
  assign new_B4594_ = new_B4601_ | new_B4600_;
  assign new_B4595_ = new_B4603_ | new_B4602_;
  assign new_B4596_ = new_B4598_ & new_B4604_;
  assign new_B4597_ = new_B4598_ & new_B4605_;
  assign new_B4598_ = new_B4588_ ^ new_B4589_;
  assign new_B4599_ = new_B4600_ ^ new_B4590_;
  assign new_B4600_ = new_B4608_ & new_B4607_;
  assign new_B4601_ = new_B4606_ & new_B4590_;
  assign new_B4602_ = new_B4611_ & new_B4610_;
  assign new_B4603_ = new_B4609_ & new_B4590_;
  assign new_B4604_ = new_B4612_ | new_B4589_;
  assign new_B4605_ = ~new_B4590_ ^ new_B4602_;
  assign new_B4606_ = ~new_B4615_ | ~new_B4616_;
  assign new_B4607_ = new_B4591_ ^ new_B4598_;
  assign new_B4608_ = new_B4617_ & new_B4610_;
  assign new_B4609_ = ~new_B4619_ | ~new_B4618_;
  assign new_B4610_ = new_B4591_ | new_B4592_;
  assign new_B4611_ = new_B4591_ | new_B4598_;
  assign new_B4612_ = new_B4590_ & new_B4602_;
  assign new_B4613_ = ~new_B4589_ | ~new_B4590_;
  assign new_B4614_ = new_B4598_ & new_B4613_;
  assign new_B4615_ = ~new_B4614_ & ~new_B4598_;
  assign new_B4616_ = new_B4598_ | new_B4613_;
  assign new_B4617_ = ~new_B4591_ | ~new_B4592_;
  assign new_B4618_ = new_B4598_ | new_B4613_;
  assign new_B4619_ = ~new_B4598_ & ~new_B4620_;
  assign new_B4620_ = new_B4598_ & new_B4613_;
  assign new_B4621_ = new_B6511_;
  assign new_B4622_ = new_B6544_;
  assign new_B4623_ = new_B6577_;
  assign new_B4624_ = new_B6610_;
  assign new_B4625_ = new_B6643_;
  assign new_B4626_ = new_B4632_ & new_B4631_;
  assign new_B4627_ = new_B4634_ | new_B4633_;
  assign new_B4628_ = new_B4636_ | new_B4635_;
  assign new_B4629_ = new_B4631_ & new_B4637_;
  assign new_B4630_ = new_B4631_ & new_B4638_;
  assign new_B4631_ = new_B4621_ ^ new_B4622_;
  assign new_B4632_ = new_B4633_ ^ new_B4623_;
  assign new_B4633_ = new_B4641_ & new_B4640_;
  assign new_B4634_ = new_B4639_ & new_B4623_;
  assign new_B4635_ = new_B4644_ & new_B4643_;
  assign new_B4636_ = new_B4642_ & new_B4623_;
  assign new_B4637_ = new_B4645_ | new_B4622_;
  assign new_B4638_ = ~new_B4623_ ^ new_B4635_;
  assign new_B4639_ = ~new_B4648_ | ~new_B4649_;
  assign new_B4640_ = new_B4624_ ^ new_B4631_;
  assign new_B4641_ = new_B4650_ & new_B4643_;
  assign new_B4642_ = ~new_B4652_ | ~new_B4651_;
  assign new_B4643_ = new_B4624_ | new_B4625_;
  assign new_B4644_ = new_B4624_ | new_B4631_;
  assign new_B4645_ = new_B4623_ & new_B4635_;
  assign new_B4646_ = ~new_B4622_ | ~new_B4623_;
  assign new_B4647_ = new_B4631_ & new_B4646_;
  assign new_B4648_ = ~new_B4647_ & ~new_B4631_;
  assign new_B4649_ = new_B4631_ | new_B4646_;
  assign new_B4650_ = ~new_B4624_ | ~new_B4625_;
  assign new_B4651_ = new_B4631_ | new_B4646_;
  assign new_B4652_ = ~new_B4631_ & ~new_B4653_;
  assign new_B4653_ = new_B4631_ & new_B4646_;
  assign new_B4654_ = new_B6676_;
  assign new_B4655_ = new_B6709_;
  assign new_B4656_ = new_B6742_;
  assign new_B4657_ = new_B6775_;
  assign new_B4658_ = new_B6808_;
  assign new_B4659_ = new_B4665_ & new_B4664_;
  assign new_B4660_ = new_B4667_ | new_B4666_;
  assign new_B4661_ = new_B4669_ | new_B4668_;
  assign new_B4662_ = new_B4664_ & new_B4670_;
  assign new_B4663_ = new_B4664_ & new_B4671_;
  assign new_B4664_ = new_B4654_ ^ new_B4655_;
  assign new_B4665_ = new_B4666_ ^ new_B4656_;
  assign new_B4666_ = new_B4674_ & new_B4673_;
  assign new_B4667_ = new_B4672_ & new_B4656_;
  assign new_B4668_ = new_B4677_ & new_B4676_;
  assign new_B4669_ = new_B4675_ & new_B4656_;
  assign new_B4670_ = new_B4678_ | new_B4655_;
  assign new_B4671_ = ~new_B4656_ ^ new_B4668_;
  assign new_B4672_ = ~new_B4681_ | ~new_B4682_;
  assign new_B4673_ = new_B4657_ ^ new_B4664_;
  assign new_B4674_ = new_B4683_ & new_B4676_;
  assign new_B4675_ = ~new_B4685_ | ~new_B4684_;
  assign new_B4676_ = new_B4657_ | new_B4658_;
  assign new_B4677_ = new_B4657_ | new_B4664_;
  assign new_B4678_ = new_B4656_ & new_B4668_;
  assign new_B4679_ = ~new_B4655_ | ~new_B4656_;
  assign new_B4680_ = new_B4664_ & new_B4679_;
  assign new_B4681_ = ~new_B4680_ & ~new_B4664_;
  assign new_B4682_ = new_B4664_ | new_B4679_;
  assign new_B4683_ = ~new_B4657_ | ~new_B4658_;
  assign new_B4684_ = new_B4664_ | new_B4679_;
  assign new_B4685_ = ~new_B4664_ & ~new_B4686_;
  assign new_B4686_ = new_B4664_ & new_B4679_;
  assign new_B4687_ = new_B6841_;
  assign new_B4688_ = new_B6874_;
  assign new_B4689_ = new_B6907_;
  assign new_B4690_ = new_B6940_;
  assign new_B4691_ = new_B6973_;
  assign new_B4692_ = new_B4698_ & new_B4697_;
  assign new_B4693_ = new_B4700_ | new_B4699_;
  assign new_B4694_ = new_B4702_ | new_B4701_;
  assign new_B4695_ = new_B4697_ & new_B4703_;
  assign new_B4696_ = new_B4697_ & new_B4704_;
  assign new_B4697_ = new_B4687_ ^ new_B4688_;
  assign new_B4698_ = new_B4699_ ^ new_B4689_;
  assign new_B4699_ = new_B4707_ & new_B4706_;
  assign new_B4700_ = new_B4705_ & new_B4689_;
  assign new_B4701_ = new_B4710_ & new_B4709_;
  assign new_B4702_ = new_B4708_ & new_B4689_;
  assign new_B4703_ = new_B4711_ | new_B4688_;
  assign new_B4704_ = ~new_B4689_ ^ new_B4701_;
  assign new_B4705_ = ~new_B4714_ | ~new_B4715_;
  assign new_B4706_ = new_B4690_ ^ new_B4697_;
  assign new_B4707_ = new_B4716_ & new_B4709_;
  assign new_B4708_ = ~new_B4718_ | ~new_B4717_;
  assign new_B4709_ = new_B4690_ | new_B4691_;
  assign new_B4710_ = new_B4690_ | new_B4697_;
  assign new_B4711_ = new_B4689_ & new_B4701_;
  assign new_B4712_ = ~new_B4688_ | ~new_B4689_;
  assign new_B4713_ = new_B4697_ & new_B4712_;
  assign new_B4714_ = ~new_B4713_ & ~new_B4697_;
  assign new_B4715_ = new_B4697_ | new_B4712_;
  assign new_B4716_ = ~new_B4690_ | ~new_B4691_;
  assign new_B4717_ = new_B4697_ | new_B4712_;
  assign new_B4718_ = ~new_B4697_ & ~new_B4719_;
  assign new_B4719_ = new_B4697_ & new_B4712_;
  assign new_B4720_ = new_B7006_;
  assign new_B4721_ = new_B7039_;
  assign new_B4722_ = new_B7072_;
  assign new_B4723_ = new_B7105_;
  assign new_B4724_ = new_B7138_;
  assign new_B4725_ = new_B4731_ & new_B4730_;
  assign new_B4726_ = new_B4733_ | new_B4732_;
  assign new_B4727_ = new_B4735_ | new_B4734_;
  assign new_B4728_ = new_B4730_ & new_B4736_;
  assign new_B4729_ = new_B4730_ & new_B4737_;
  assign new_B4730_ = new_B4720_ ^ new_B4721_;
  assign new_B4731_ = new_B4732_ ^ new_B4722_;
  assign new_B4732_ = new_B4740_ & new_B4739_;
  assign new_B4733_ = new_B4738_ & new_B4722_;
  assign new_B4734_ = new_B4743_ & new_B4742_;
  assign new_B4735_ = new_B4741_ & new_B4722_;
  assign new_B4736_ = new_B4744_ | new_B4721_;
  assign new_B4737_ = ~new_B4722_ ^ new_B4734_;
  assign new_B4738_ = ~new_B4747_ | ~new_B4748_;
  assign new_B4739_ = new_B4723_ ^ new_B4730_;
  assign new_B4740_ = new_B4749_ & new_B4742_;
  assign new_B4741_ = ~new_B4751_ | ~new_B4750_;
  assign new_B4742_ = new_B4723_ | new_B4724_;
  assign new_B4743_ = new_B4723_ | new_B4730_;
  assign new_B4744_ = new_B4722_ & new_B4734_;
  assign new_B4745_ = ~new_B4721_ | ~new_B4722_;
  assign new_B4746_ = new_B4730_ & new_B4745_;
  assign new_B4747_ = ~new_B4746_ & ~new_B4730_;
  assign new_B4748_ = new_B4730_ | new_B4745_;
  assign new_B4749_ = ~new_B4723_ | ~new_B4724_;
  assign new_B4750_ = new_B4730_ | new_B4745_;
  assign new_B4751_ = ~new_B4730_ & ~new_B4752_;
  assign new_B4752_ = new_B4730_ & new_B4745_;
  assign new_B4753_ = new_B7171_;
  assign new_B4754_ = new_B7204_;
  assign new_B4755_ = new_B7237_;
  assign new_B4756_ = new_B7270_;
  assign new_B4757_ = new_B7303_;
  assign new_B4758_ = new_B4764_ & new_B4763_;
  assign new_B4759_ = new_B4766_ | new_B4765_;
  assign new_B4760_ = new_B4768_ | new_B4767_;
  assign new_B4761_ = new_B4763_ & new_B4769_;
  assign new_B4762_ = new_B4763_ & new_B4770_;
  assign new_B4763_ = new_B4753_ ^ new_B4754_;
  assign new_B4764_ = new_B4765_ ^ new_B4755_;
  assign new_B4765_ = new_B4773_ & new_B4772_;
  assign new_B4766_ = new_B4771_ & new_B4755_;
  assign new_B4767_ = new_B4776_ & new_B4775_;
  assign new_B4768_ = new_B4774_ & new_B4755_;
  assign new_B4769_ = new_B4777_ | new_B4754_;
  assign new_B4770_ = ~new_B4755_ ^ new_B4767_;
  assign new_B4771_ = ~new_B4780_ | ~new_B4781_;
  assign new_B4772_ = new_B4756_ ^ new_B4763_;
  assign new_B4773_ = new_B4782_ & new_B4775_;
  assign new_B4774_ = ~new_B4784_ | ~new_B4783_;
  assign new_B4775_ = new_B4756_ | new_B4757_;
  assign new_B4776_ = new_B4756_ | new_B4763_;
  assign new_B4777_ = new_B4755_ & new_B4767_;
  assign new_B4778_ = ~new_B4754_ | ~new_B4755_;
  assign new_B4779_ = new_B4763_ & new_B4778_;
  assign new_B4780_ = ~new_B4779_ & ~new_B4763_;
  assign new_B4781_ = new_B4763_ | new_B4778_;
  assign new_B4782_ = ~new_B4756_ | ~new_B4757_;
  assign new_B4783_ = new_B4763_ | new_B4778_;
  assign new_B4784_ = ~new_B4763_ & ~new_B4785_;
  assign new_B4785_ = new_B4763_ & new_B4778_;
  assign new_B4786_ = new_B7336_;
  assign new_B4787_ = new_B7369_;
  assign new_B4788_ = new_B7402_;
  assign new_B4789_ = new_B7435_;
  assign new_B4790_ = new_B7468_;
  assign new_B4791_ = new_B4797_ & new_B4796_;
  assign new_B4792_ = new_B4799_ | new_B4798_;
  assign new_B4793_ = new_B4801_ | new_B4800_;
  assign new_B4794_ = new_B4796_ & new_B4802_;
  assign new_B4795_ = new_B4796_ & new_B4803_;
  assign new_B4796_ = new_B4786_ ^ new_B4787_;
  assign new_B4797_ = new_B4798_ ^ new_B4788_;
  assign new_B4798_ = new_B4806_ & new_B4805_;
  assign new_B4799_ = new_B4804_ & new_B4788_;
  assign new_B4800_ = new_B4809_ & new_B4808_;
  assign new_B4801_ = new_B4807_ & new_B4788_;
  assign new_B4802_ = new_B4810_ | new_B4787_;
  assign new_B4803_ = ~new_B4788_ ^ new_B4800_;
  assign new_B4804_ = ~new_B4813_ | ~new_B4814_;
  assign new_B4805_ = new_B4789_ ^ new_B4796_;
  assign new_B4806_ = new_B4815_ & new_B4808_;
  assign new_B4807_ = ~new_B4817_ | ~new_B4816_;
  assign new_B4808_ = new_B4789_ | new_B4790_;
  assign new_B4809_ = new_B4789_ | new_B4796_;
  assign new_B4810_ = new_B4788_ & new_B4800_;
  assign new_B4811_ = ~new_B4787_ | ~new_B4788_;
  assign new_B4812_ = new_B4796_ & new_B4811_;
  assign new_B4813_ = ~new_B4812_ & ~new_B4796_;
  assign new_B4814_ = new_B4796_ | new_B4811_;
  assign new_B4815_ = ~new_B4789_ | ~new_B4790_;
  assign new_B4816_ = new_B4796_ | new_B4811_;
  assign new_B4817_ = ~new_B4796_ & ~new_B4818_;
  assign new_B4818_ = new_B4796_ & new_B4811_;
  assign new_B4819_ = new_B7501_;
  assign new_B4820_ = new_B7534_;
  assign new_B4821_ = new_B7567_;
  assign new_B4822_ = new_B7600_;
  assign new_B4823_ = new_B7633_;
  assign new_B4824_ = new_B4830_ & new_B4829_;
  assign new_B4825_ = new_B4832_ | new_B4831_;
  assign new_B4826_ = new_B4834_ | new_B4833_;
  assign new_B4827_ = new_B4829_ & new_B4835_;
  assign new_B4828_ = new_B4829_ & new_B4836_;
  assign new_B4829_ = new_B4819_ ^ new_B4820_;
  assign new_B4830_ = new_B4831_ ^ new_B4821_;
  assign new_B4831_ = new_B4839_ & new_B4838_;
  assign new_B4832_ = new_B4837_ & new_B4821_;
  assign new_B4833_ = new_B4842_ & new_B4841_;
  assign new_B4834_ = new_B4840_ & new_B4821_;
  assign new_B4835_ = new_B4843_ | new_B4820_;
  assign new_B4836_ = ~new_B4821_ ^ new_B4833_;
  assign new_B4837_ = ~new_B4846_ | ~new_B4847_;
  assign new_B4838_ = new_B4822_ ^ new_B4829_;
  assign new_B4839_ = new_B4848_ & new_B4841_;
  assign new_B4840_ = ~new_B4850_ | ~new_B4849_;
  assign new_B4841_ = new_B4822_ | new_B4823_;
  assign new_B4842_ = new_B4822_ | new_B4829_;
  assign new_B4843_ = new_B4821_ & new_B4833_;
  assign new_B4844_ = ~new_B4820_ | ~new_B4821_;
  assign new_B4845_ = new_B4829_ & new_B4844_;
  assign new_B4846_ = ~new_B4845_ & ~new_B4829_;
  assign new_B4847_ = new_B4829_ | new_B4844_;
  assign new_B4848_ = ~new_B4822_ | ~new_B4823_;
  assign new_B4849_ = new_B4829_ | new_B4844_;
  assign new_B4850_ = ~new_B4829_ & ~new_B4851_;
  assign new_B4851_ = new_B4829_ & new_B4844_;
  assign new_B4852_ = new_B7666_;
  assign new_B4853_ = new_B7699_;
  assign new_B4854_ = new_B7732_;
  assign new_B4855_ = new_B7765_;
  assign new_B4856_ = new_B7798_;
  assign new_B4857_ = new_B4863_ & new_B4862_;
  assign new_B4858_ = new_B4865_ | new_B4864_;
  assign new_B4859_ = new_B4867_ | new_B4866_;
  assign new_B4860_ = new_B4862_ & new_B4868_;
  assign new_B4861_ = new_B4862_ & new_B4869_;
  assign new_B4862_ = new_B4852_ ^ new_B4853_;
  assign new_B4863_ = new_B4864_ ^ new_B4854_;
  assign new_B4864_ = new_B4872_ & new_B4871_;
  assign new_B4865_ = new_B4870_ & new_B4854_;
  assign new_B4866_ = new_B4875_ & new_B4874_;
  assign new_B4867_ = new_B4873_ & new_B4854_;
  assign new_B4868_ = new_B4876_ | new_B4853_;
  assign new_B4869_ = ~new_B4854_ ^ new_B4866_;
  assign new_B4870_ = ~new_B4879_ | ~new_B4880_;
  assign new_B4871_ = new_B4855_ ^ new_B4862_;
  assign new_B4872_ = new_B4881_ & new_B4874_;
  assign new_B4873_ = ~new_B4883_ | ~new_B4882_;
  assign new_B4874_ = new_B4855_ | new_B4856_;
  assign new_B4875_ = new_B4855_ | new_B4862_;
  assign new_B4876_ = new_B4854_ & new_B4866_;
  assign new_B4877_ = ~new_B4853_ | ~new_B4854_;
  assign new_B4878_ = new_B4862_ & new_B4877_;
  assign new_B4879_ = ~new_B4878_ & ~new_B4862_;
  assign new_B4880_ = new_B4862_ | new_B4877_;
  assign new_B4881_ = ~new_B4855_ | ~new_B4856_;
  assign new_B4882_ = new_B4862_ | new_B4877_;
  assign new_B4883_ = ~new_B4862_ & ~new_B4884_;
  assign new_B4884_ = new_B4862_ & new_B4877_;
  assign new_B4885_ = new_B7831_;
  assign new_B4886_ = new_B7864_;
  assign new_B4887_ = new_B7897_;
  assign new_B4888_ = new_B7930_;
  assign new_B4889_ = new_B7963_;
  assign new_B4890_ = new_B4896_ & new_B4895_;
  assign new_B4891_ = new_B4898_ | new_B4897_;
  assign new_B4892_ = new_B4900_ | new_B4899_;
  assign new_B4893_ = new_B4895_ & new_B4901_;
  assign new_B4894_ = new_B4895_ & new_B4902_;
  assign new_B4895_ = new_B4885_ ^ new_B4886_;
  assign new_B4896_ = new_B4897_ ^ new_B4887_;
  assign new_B4897_ = new_B4905_ & new_B4904_;
  assign new_B4898_ = new_B4903_ & new_B4887_;
  assign new_B4899_ = new_B4908_ & new_B4907_;
  assign new_B4900_ = new_B4906_ & new_B4887_;
  assign new_B4901_ = new_B4909_ | new_B4886_;
  assign new_B4902_ = ~new_B4887_ ^ new_B4899_;
  assign new_B4903_ = ~new_B4912_ | ~new_B4913_;
  assign new_B4904_ = new_B4888_ ^ new_B4895_;
  assign new_B4905_ = new_B4914_ & new_B4907_;
  assign new_B4906_ = ~new_B4916_ | ~new_B4915_;
  assign new_B4907_ = new_B4888_ | new_B4889_;
  assign new_B4908_ = new_B4888_ | new_B4895_;
  assign new_B4909_ = new_B4887_ & new_B4899_;
  assign new_B4910_ = ~new_B4886_ | ~new_B4887_;
  assign new_B4911_ = new_B4895_ & new_B4910_;
  assign new_B4912_ = ~new_B4911_ & ~new_B4895_;
  assign new_B4913_ = new_B4895_ | new_B4910_;
  assign new_B4914_ = ~new_B4888_ | ~new_B4889_;
  assign new_B4915_ = new_B4895_ | new_B4910_;
  assign new_B4916_ = ~new_B4895_ & ~new_B4917_;
  assign new_B4917_ = new_B4895_ & new_B4910_;
  assign new_B4918_ = new_B7996_;
  assign new_B4919_ = new_B8029_;
  assign new_B4920_ = new_B8062_;
  assign new_B4921_ = new_B8095_;
  assign new_B4922_ = new_B8128_;
  assign new_B4923_ = new_B4929_ & new_B4928_;
  assign new_B4924_ = new_B4931_ | new_B4930_;
  assign new_B4925_ = new_B4933_ | new_B4932_;
  assign new_B4926_ = new_B4928_ & new_B4934_;
  assign new_B4927_ = new_B4928_ & new_B4935_;
  assign new_B4928_ = new_B4918_ ^ new_B4919_;
  assign new_B4929_ = new_B4930_ ^ new_B4920_;
  assign new_B4930_ = new_B4938_ & new_B4937_;
  assign new_B4931_ = new_B4936_ & new_B4920_;
  assign new_B4932_ = new_B4941_ & new_B4940_;
  assign new_B4933_ = new_B4939_ & new_B4920_;
  assign new_B4934_ = new_B4942_ | new_B4919_;
  assign new_B4935_ = ~new_B4920_ ^ new_B4932_;
  assign new_B4936_ = ~new_B4945_ | ~new_B4946_;
  assign new_B4937_ = new_B4921_ ^ new_B4928_;
  assign new_B4938_ = new_B4947_ & new_B4940_;
  assign new_B4939_ = ~new_B4949_ | ~new_B4948_;
  assign new_B4940_ = new_B4921_ | new_B4922_;
  assign new_B4941_ = new_B4921_ | new_B4928_;
  assign new_B4942_ = new_B4920_ & new_B4932_;
  assign new_B4943_ = ~new_B4919_ | ~new_B4920_;
  assign new_B4944_ = new_B4928_ & new_B4943_;
  assign new_B4945_ = ~new_B4944_ & ~new_B4928_;
  assign new_B4946_ = new_B4928_ | new_B4943_;
  assign new_B4947_ = ~new_B4921_ | ~new_B4922_;
  assign new_B4948_ = new_B4928_ | new_B4943_;
  assign new_B4949_ = ~new_B4928_ & ~new_B4950_;
  assign new_B4950_ = new_B4928_ & new_B4943_;
  assign new_B4951_ = new_B8161_;
  assign new_B4952_ = new_B8194_;
  assign new_B4953_ = new_B8227_;
  assign new_B4954_ = new_B8260_;
  assign new_B4955_ = new_B8293_;
  assign new_B4956_ = new_B4962_ & new_B4961_;
  assign new_B4957_ = new_B4964_ | new_B4963_;
  assign new_B4958_ = new_B4966_ | new_B4965_;
  assign new_B4959_ = new_B4961_ & new_B4967_;
  assign new_B4960_ = new_B4961_ & new_B4968_;
  assign new_B4961_ = new_B4951_ ^ new_B4952_;
  assign new_B4962_ = new_B4963_ ^ new_B4953_;
  assign new_B4963_ = new_B4971_ & new_B4970_;
  assign new_B4964_ = new_B4969_ & new_B4953_;
  assign new_B4965_ = new_B4974_ & new_B4973_;
  assign new_B4966_ = new_B4972_ & new_B4953_;
  assign new_B4967_ = new_B4975_ | new_B4952_;
  assign new_B4968_ = ~new_B4953_ ^ new_B4965_;
  assign new_B4969_ = ~new_B4978_ | ~new_B4979_;
  assign new_B4970_ = new_B4954_ ^ new_B4961_;
  assign new_B4971_ = new_B4980_ & new_B4973_;
  assign new_B4972_ = ~new_B4982_ | ~new_B4981_;
  assign new_B4973_ = new_B4954_ | new_B4955_;
  assign new_B4974_ = new_B4954_ | new_B4961_;
  assign new_B4975_ = new_B4953_ & new_B4965_;
  assign new_B4976_ = ~new_B4952_ | ~new_B4953_;
  assign new_B4977_ = new_B4961_ & new_B4976_;
  assign new_B4978_ = ~new_B4977_ & ~new_B4961_;
  assign new_B4979_ = new_B4961_ | new_B4976_;
  assign new_B4980_ = ~new_B4954_ | ~new_B4955_;
  assign new_B4981_ = new_B4961_ | new_B4976_;
  assign new_B4982_ = ~new_B4961_ & ~new_B4983_;
  assign new_B4983_ = new_B4961_ & new_B4976_;
  assign new_B4984_ = new_B8326_;
  assign new_B4985_ = new_B8359_;
  assign new_B4986_ = new_B8392_;
  assign new_B4987_ = new_B8425_;
  assign new_B4988_ = new_B8458_;
  assign new_B4989_ = new_B4995_ & new_B4994_;
  assign new_B4990_ = new_B4997_ | new_B4996_;
  assign new_B4991_ = new_B4999_ | new_B4998_;
  assign new_B4992_ = new_B4994_ & new_B5000_;
  assign new_B4993_ = new_B4994_ & new_B5001_;
  assign new_B4994_ = new_B4984_ ^ new_B4985_;
  assign new_B4995_ = new_B4996_ ^ new_B4986_;
  assign new_B4996_ = new_B5004_ & new_B5003_;
  assign new_B4997_ = new_B5002_ & new_B4986_;
  assign new_B4998_ = new_B5007_ & new_B5006_;
  assign new_B4999_ = new_B5005_ & new_B4986_;
  assign new_B5000_ = new_B5008_ | new_B4985_;
  assign new_B5001_ = ~new_B4986_ ^ new_B4998_;
  assign new_B5002_ = ~new_B5011_ | ~new_B5012_;
  assign new_B5003_ = new_B4987_ ^ new_B4994_;
  assign new_B5004_ = new_B5013_ & new_B5006_;
  assign new_B5005_ = ~new_B5015_ | ~new_B5014_;
  assign new_B5006_ = new_B4987_ | new_B4988_;
  assign new_B5007_ = new_B4987_ | new_B4994_;
  assign new_B5008_ = new_B4986_ & new_B4998_;
  assign new_B5009_ = ~new_B4985_ | ~new_B4986_;
  assign new_B5010_ = new_B4994_ & new_B5009_;
  assign new_B5011_ = ~new_B5010_ & ~new_B4994_;
  assign new_B5012_ = new_B4994_ | new_B5009_;
  assign new_B5013_ = ~new_B4987_ | ~new_B4988_;
  assign new_B5014_ = new_B4994_ | new_B5009_;
  assign new_B5015_ = ~new_B4994_ & ~new_B5016_;
  assign new_B5016_ = new_B4994_ & new_B5009_;
  assign new_B5017_ = new_B8491_;
  assign new_B5018_ = new_B8524_;
  assign new_B5019_ = new_B8557_;
  assign new_B5020_ = new_B8590_;
  assign new_B5021_ = new_B8623_;
  assign new_B5022_ = new_B5028_ & new_B5027_;
  assign new_B5023_ = new_B5030_ | new_B5029_;
  assign new_B5024_ = new_B5032_ | new_B5031_;
  assign new_B5025_ = new_B5027_ & new_B5033_;
  assign new_B5026_ = new_B5027_ & new_B5034_;
  assign new_B5027_ = new_B5017_ ^ new_B5018_;
  assign new_B5028_ = new_B5029_ ^ new_B5019_;
  assign new_B5029_ = new_B5037_ & new_B5036_;
  assign new_B5030_ = new_B5035_ & new_B5019_;
  assign new_B5031_ = new_B5040_ & new_B5039_;
  assign new_B5032_ = new_B5038_ & new_B5019_;
  assign new_B5033_ = new_B5041_ | new_B5018_;
  assign new_B5034_ = ~new_B5019_ ^ new_B5031_;
  assign new_B5035_ = ~new_B5044_ | ~new_B5045_;
  assign new_B5036_ = new_B5020_ ^ new_B5027_;
  assign new_B5037_ = new_B5046_ & new_B5039_;
  assign new_B5038_ = ~new_B5048_ | ~new_B5047_;
  assign new_B5039_ = new_B5020_ | new_B5021_;
  assign new_B5040_ = new_B5020_ | new_B5027_;
  assign new_B5041_ = new_B5019_ & new_B5031_;
  assign new_B5042_ = ~new_B5018_ | ~new_B5019_;
  assign new_B5043_ = new_B5027_ & new_B5042_;
  assign new_B5044_ = ~new_B5043_ & ~new_B5027_;
  assign new_B5045_ = new_B5027_ | new_B5042_;
  assign new_B5046_ = ~new_B5020_ | ~new_B5021_;
  assign new_B5047_ = new_B5027_ | new_B5042_;
  assign new_B5048_ = ~new_B5027_ & ~new_B5049_;
  assign new_B5049_ = new_B5027_ & new_B5042_;
  assign new_B5050_ = new_B8656_;
  assign new_B5051_ = new_B8689_;
  assign new_B5052_ = new_B8722_;
  assign new_B5053_ = new_B8755_;
  assign new_B5054_ = new_B8788_;
  assign new_B5055_ = new_B5061_ & new_B5060_;
  assign new_B5056_ = new_B5063_ | new_B5062_;
  assign new_B5057_ = new_B5065_ | new_B5064_;
  assign new_B5058_ = new_B5060_ & new_B5066_;
  assign new_B5059_ = new_B5060_ & new_B5067_;
  assign new_B5060_ = new_B5050_ ^ new_B5051_;
  assign new_B5061_ = new_B5062_ ^ new_B5052_;
  assign new_B5062_ = new_B5070_ & new_B5069_;
  assign new_B5063_ = new_B5068_ & new_B5052_;
  assign new_B5064_ = new_B5073_ & new_B5072_;
  assign new_B5065_ = new_B5071_ & new_B5052_;
  assign new_B5066_ = new_B5074_ | new_B5051_;
  assign new_B5067_ = ~new_B5052_ ^ new_B5064_;
  assign new_B5068_ = ~new_B5077_ | ~new_B5078_;
  assign new_B5069_ = new_B5053_ ^ new_B5060_;
  assign new_B5070_ = new_B5079_ & new_B5072_;
  assign new_B5071_ = ~new_B5081_ | ~new_B5080_;
  assign new_B5072_ = new_B5053_ | new_B5054_;
  assign new_B5073_ = new_B5053_ | new_B5060_;
  assign new_B5074_ = new_B5052_ & new_B5064_;
  assign new_B5075_ = ~new_B5051_ | ~new_B5052_;
  assign new_B5076_ = new_B5060_ & new_B5075_;
  assign new_B5077_ = ~new_B5076_ & ~new_B5060_;
  assign new_B5078_ = new_B5060_ | new_B5075_;
  assign new_B5079_ = ~new_B5053_ | ~new_B5054_;
  assign new_B5080_ = new_B5060_ | new_B5075_;
  assign new_B5081_ = ~new_B5060_ & ~new_B5082_;
  assign new_B5082_ = new_B5060_ & new_B5075_;
  assign new_B5083_ = new_B8821_;
  assign new_B5084_ = new_B8854_;
  assign new_B5085_ = new_B8887_;
  assign new_B5086_ = new_B8920_;
  assign new_B5087_ = new_B8953_;
  assign new_B5088_ = new_B5094_ & new_B5093_;
  assign new_B5089_ = new_B5096_ | new_B5095_;
  assign new_B5090_ = new_B5098_ | new_B5097_;
  assign new_B5091_ = new_B5093_ & new_B5099_;
  assign new_B5092_ = new_B5093_ & new_B5100_;
  assign new_B5093_ = new_B5083_ ^ new_B5084_;
  assign new_B5094_ = new_B5095_ ^ new_B5085_;
  assign new_B5095_ = new_B5103_ & new_B5102_;
  assign new_B5096_ = new_B5101_ & new_B5085_;
  assign new_B5097_ = new_B5106_ & new_B5105_;
  assign new_B5098_ = new_B5104_ & new_B5085_;
  assign new_B5099_ = new_B5107_ | new_B5084_;
  assign new_B5100_ = ~new_B5085_ ^ new_B5097_;
  assign new_B5101_ = ~new_B5110_ | ~new_B5111_;
  assign new_B5102_ = new_B5086_ ^ new_B5093_;
  assign new_B5103_ = new_B5112_ & new_B5105_;
  assign new_B5104_ = ~new_B5114_ | ~new_B5113_;
  assign new_B5105_ = new_B5086_ | new_B5087_;
  assign new_B5106_ = new_B5086_ | new_B5093_;
  assign new_B5107_ = new_B5085_ & new_B5097_;
  assign new_B5108_ = ~new_B5084_ | ~new_B5085_;
  assign new_B5109_ = new_B5093_ & new_B5108_;
  assign new_B5110_ = ~new_B5109_ & ~new_B5093_;
  assign new_B5111_ = new_B5093_ | new_B5108_;
  assign new_B5112_ = ~new_B5086_ | ~new_B5087_;
  assign new_B5113_ = new_B5093_ | new_B5108_;
  assign new_B5114_ = ~new_B5093_ & ~new_B5115_;
  assign new_B5115_ = new_B5093_ & new_B5108_;
  assign new_B5116_ = new_B8986_;
  assign new_B5117_ = new_B9019_;
  assign new_B5118_ = new_B9052_;
  assign new_B5119_ = new_B9085_;
  assign new_B5120_ = new_B9118_;
  assign new_B5121_ = new_B5127_ & new_B5126_;
  assign new_B5122_ = new_B5129_ | new_B5128_;
  assign new_B5123_ = new_B5131_ | new_B5130_;
  assign new_B5124_ = new_B5126_ & new_B5132_;
  assign new_B5125_ = new_B5126_ & new_B5133_;
  assign new_B5126_ = new_B5116_ ^ new_B5117_;
  assign new_B5127_ = new_B5128_ ^ new_B5118_;
  assign new_B5128_ = new_B5136_ & new_B5135_;
  assign new_B5129_ = new_B5134_ & new_B5118_;
  assign new_B5130_ = new_B5139_ & new_B5138_;
  assign new_B5131_ = new_B5137_ & new_B5118_;
  assign new_B5132_ = new_B5140_ | new_B5117_;
  assign new_B5133_ = ~new_B5118_ ^ new_B5130_;
  assign new_B5134_ = ~new_B5143_ | ~new_B5144_;
  assign new_B5135_ = new_B5119_ ^ new_B5126_;
  assign new_B5136_ = new_B5145_ & new_B5138_;
  assign new_B5137_ = ~new_B5147_ | ~new_B5146_;
  assign new_B5138_ = new_B5119_ | new_B5120_;
  assign new_B5139_ = new_B5119_ | new_B5126_;
  assign new_B5140_ = new_B5118_ & new_B5130_;
  assign new_B5141_ = ~new_B5117_ | ~new_B5118_;
  assign new_B5142_ = new_B5126_ & new_B5141_;
  assign new_B5143_ = ~new_B5142_ & ~new_B5126_;
  assign new_B5144_ = new_B5126_ | new_B5141_;
  assign new_B5145_ = ~new_B5119_ | ~new_B5120_;
  assign new_B5146_ = new_B5126_ | new_B5141_;
  assign new_B5147_ = ~new_B5126_ & ~new_B5148_;
  assign new_B5148_ = new_B5126_ & new_B5141_;
  assign new_B5149_ = new_B9151_;
  assign new_B5150_ = new_B9184_;
  assign new_B5151_ = new_B9217_;
  assign new_B5152_ = new_B9250_;
  assign new_B5153_ = new_B9283_;
  assign new_B5154_ = new_B5160_ & new_B5159_;
  assign new_B5155_ = new_B5162_ | new_B5161_;
  assign new_B5156_ = new_B5164_ | new_B5163_;
  assign new_B5157_ = new_B5159_ & new_B5165_;
  assign new_B5158_ = new_B5159_ & new_B5166_;
  assign new_B5159_ = new_B5149_ ^ new_B5150_;
  assign new_B5160_ = new_B5161_ ^ new_B5151_;
  assign new_B5161_ = new_B5169_ & new_B5168_;
  assign new_B5162_ = new_B5167_ & new_B5151_;
  assign new_B5163_ = new_B5172_ & new_B5171_;
  assign new_B5164_ = new_B5170_ & new_B5151_;
  assign new_B5165_ = new_B5173_ | new_B5150_;
  assign new_B5166_ = ~new_B5151_ ^ new_B5163_;
  assign new_B5167_ = ~new_B5176_ | ~new_B5177_;
  assign new_B5168_ = new_B5152_ ^ new_B5159_;
  assign new_B5169_ = new_B5178_ & new_B5171_;
  assign new_B5170_ = ~new_B5180_ | ~new_B5179_;
  assign new_B5171_ = new_B5152_ | new_B5153_;
  assign new_B5172_ = new_B5152_ | new_B5159_;
  assign new_B5173_ = new_B5151_ & new_B5163_;
  assign new_B5174_ = ~new_B5150_ | ~new_B5151_;
  assign new_B5175_ = new_B5159_ & new_B5174_;
  assign new_B5176_ = ~new_B5175_ & ~new_B5159_;
  assign new_B5177_ = new_B5159_ | new_B5174_;
  assign new_B5178_ = ~new_B5152_ | ~new_B5153_;
  assign new_B5179_ = new_B5159_ | new_B5174_;
  assign new_B5180_ = ~new_B5159_ & ~new_B5181_;
  assign new_B5181_ = new_B5159_ & new_B5174_;
  assign new_A6963_ = new_A6941_ & new_A6956_;
  assign new_A6962_ = ~new_A6941_ & ~new_A6963_;
  assign new_A6961_ = new_A6941_ | new_A6956_;
  assign new_A6960_ = ~new_A6934_ | ~new_A6935_;
  assign new_A6959_ = new_A6941_ | new_A6956_;
  assign new_A6958_ = ~new_A6957_ & ~new_A6941_;
  assign new_A6957_ = new_A6941_ & new_A6956_;
  assign new_A6956_ = ~new_A6932_ | ~new_A6933_;
  assign new_A6955_ = new_A6933_ & new_A6945_;
  assign new_A6954_ = new_A6934_ | new_A6941_;
  assign new_A6953_ = new_A6934_ | new_A6935_;
  assign new_A6952_ = ~new_A6962_ | ~new_A6961_;
  assign new_A6951_ = new_A6960_ & new_A6953_;
  assign new_A6950_ = new_A6934_ ^ new_A6941_;
  assign new_A6949_ = ~new_A6958_ | ~new_A6959_;
  assign new_A6948_ = ~new_A6933_ ^ new_A6945_;
  assign new_A6947_ = new_A6955_ | new_A6932_;
  assign new_A6946_ = new_A6952_ & new_A6933_;
  assign new_A6945_ = new_A6954_ & new_A6953_;
  assign new_A6944_ = new_A6949_ & new_A6933_;
  assign new_A6943_ = new_A6951_ & new_A6950_;
  assign new_A6942_ = new_A6943_ ^ new_A6933_;
  assign new_A6941_ = new_A6931_ ^ new_A6932_;
  assign new_A6940_ = new_A6941_ & new_A6948_;
  assign new_A6939_ = new_A6941_ & new_A6947_;
  assign new_A6938_ = new_A6946_ | new_A6945_;
  assign new_A6937_ = new_A6944_ | new_A6943_;
  assign new_A6936_ = new_A6942_ & new_A6941_;
  assign new_A6935_ = new_B1066_;
  assign new_A6934_ = new_B1095_;
  assign new_A6933_ = new_B1128_;
  assign new_A6932_ = new_B1161_;
  assign new_A6931_ = new_B1194_;
  assign new_A6964_ = new_B1227_;
  assign new_A6965_ = new_B1260_;
  assign new_A6966_ = new_B1293_;
  assign new_A6967_ = new_B1326_;
  assign new_A6968_ = new_B1359_;
  assign new_A6969_ = new_A6975_ & new_A6974_;
  assign new_A6970_ = new_A6977_ | new_A6976_;
  assign new_A6971_ = new_A6979_ | new_A6978_;
  assign new_A6972_ = new_A6974_ & new_A6980_;
  assign new_A6973_ = new_A6974_ & new_A6981_;
  assign new_A6974_ = new_A6964_ ^ new_A6965_;
  assign new_A6975_ = new_A6976_ ^ new_A6966_;
  assign new_A6976_ = new_A6984_ & new_A6983_;
  assign new_A6977_ = new_A6982_ & new_A6966_;
  assign new_A6978_ = new_A6987_ & new_A6986_;
  assign new_A6979_ = new_A6985_ & new_A6966_;
  assign new_A6980_ = new_A6988_ | new_A6965_;
  assign new_A6981_ = ~new_A6966_ ^ new_A6978_;
  assign new_A6982_ = ~new_A6991_ | ~new_A6992_;
  assign new_A6983_ = new_A6967_ ^ new_A6974_;
  assign new_A6984_ = new_A6993_ & new_A6986_;
  assign new_A6985_ = ~new_A6995_ | ~new_A6994_;
  assign new_A6986_ = new_A6967_ | new_A6968_;
  assign new_A6987_ = new_A6967_ | new_A6974_;
  assign new_A6988_ = new_A6966_ & new_A6978_;
  assign new_A6989_ = ~new_A6965_ | ~new_A6966_;
  assign new_A6990_ = new_A6974_ & new_A6989_;
  assign new_A6991_ = ~new_A6990_ & ~new_A6974_;
  assign new_A6992_ = new_A6974_ | new_A6989_;
  assign new_A6993_ = ~new_A6967_ | ~new_A6968_;
  assign new_A6994_ = new_A6974_ | new_A6989_;
  assign new_A6995_ = ~new_A6974_ & ~new_A6996_;
  assign new_A6996_ = new_A6974_ & new_A6989_;
  assign new_A6997_ = new_B1392_;
  assign new_A6998_ = new_B1425_;
  assign new_A6999_ = new_B1458_;
  assign new_A7000_ = new_B1491_;
  assign new_A7001_ = new_B1524_;
  assign new_A7002_ = new_A7008_ & new_A7007_;
  assign new_A7003_ = new_A7010_ | new_A7009_;
  assign new_A7004_ = new_A7012_ | new_A7011_;
  assign new_A7005_ = new_A7007_ & new_A7013_;
  assign new_A7006_ = new_A7007_ & new_A7014_;
  assign new_A7007_ = new_A6997_ ^ new_A6998_;
  assign new_A7008_ = new_A7009_ ^ new_A6999_;
  assign new_A7009_ = new_A7017_ & new_A7016_;
  assign new_A7010_ = new_A7015_ & new_A6999_;
  assign new_A7011_ = new_A7020_ & new_A7019_;
  assign new_A7012_ = new_A7018_ & new_A6999_;
  assign new_A7013_ = new_A7021_ | new_A6998_;
  assign new_A7014_ = ~new_A6999_ ^ new_A7011_;
  assign new_A7015_ = ~new_A7024_ | ~new_A7025_;
  assign new_A7016_ = new_A7000_ ^ new_A7007_;
  assign new_A7017_ = new_A7026_ & new_A7019_;
  assign new_A7018_ = ~new_A7028_ | ~new_A7027_;
  assign new_A7019_ = new_A7000_ | new_A7001_;
  assign new_A7020_ = new_A7000_ | new_A7007_;
  assign new_A7021_ = new_A6999_ & new_A7011_;
  assign new_A7022_ = ~new_A6998_ | ~new_A6999_;
  assign new_A7023_ = new_A7007_ & new_A7022_;
  assign new_A7024_ = ~new_A7023_ & ~new_A7007_;
  assign new_A7025_ = new_A7007_ | new_A7022_;
  assign new_A7026_ = ~new_A7000_ | ~new_A7001_;
  assign new_A7027_ = new_A7007_ | new_A7022_;
  assign new_A7028_ = ~new_A7007_ & ~new_A7029_;
  assign new_A7029_ = new_A7007_ & new_A7022_;
  assign new_A7030_ = new_B1557_;
  assign new_A7031_ = new_B1590_;
  assign new_A7032_ = new_B1623_;
  assign new_A7033_ = new_B1656_;
  assign new_A7034_ = new_B1689_;
  assign new_A7035_ = new_A7041_ & new_A7040_;
  assign new_A7036_ = new_A7043_ | new_A7042_;
  assign new_A7037_ = new_A7045_ | new_A7044_;
  assign new_A7038_ = new_A7040_ & new_A7046_;
  assign new_A7039_ = new_A7040_ & new_A7047_;
  assign new_A7040_ = new_A7030_ ^ new_A7031_;
  assign new_A7041_ = new_A7042_ ^ new_A7032_;
  assign new_A7042_ = new_A7050_ & new_A7049_;
  assign new_A7043_ = new_A7048_ & new_A7032_;
  assign new_A7044_ = new_A7053_ & new_A7052_;
  assign new_A7045_ = new_A7051_ & new_A7032_;
  assign new_A7046_ = new_A7054_ | new_A7031_;
  assign new_A7047_ = ~new_A7032_ ^ new_A7044_;
  assign new_A7048_ = ~new_A7057_ | ~new_A7058_;
  assign new_A7049_ = new_A7033_ ^ new_A7040_;
  assign new_A7050_ = new_A7059_ & new_A7052_;
  assign new_A7051_ = ~new_A7061_ | ~new_A7060_;
  assign new_A7052_ = new_A7033_ | new_A7034_;
  assign new_A7053_ = new_A7033_ | new_A7040_;
  assign new_A7054_ = new_A7032_ & new_A7044_;
  assign new_A7055_ = ~new_A7031_ | ~new_A7032_;
  assign new_A7056_ = new_A7040_ & new_A7055_;
  assign new_A7057_ = ~new_A7056_ & ~new_A7040_;
  assign new_A7058_ = new_A7040_ | new_A7055_;
  assign new_A7059_ = ~new_A7033_ | ~new_A7034_;
  assign new_A7060_ = new_A7040_ | new_A7055_;
  assign new_A7061_ = ~new_A7040_ & ~new_A7062_;
  assign new_A7062_ = new_A7040_ & new_A7055_;
  assign new_A7063_ = new_B1722_;
  assign new_A7064_ = new_B1755_;
  assign new_A7065_ = new_B1788_;
  assign new_A7066_ = new_B1821_;
  assign new_A7067_ = new_B1854_;
  assign new_A7068_ = new_A7074_ & new_A7073_;
  assign new_A7069_ = new_A7076_ | new_A7075_;
  assign new_A7070_ = new_A7078_ | new_A7077_;
  assign new_A7071_ = new_A7073_ & new_A7079_;
  assign new_A7072_ = new_A7073_ & new_A7080_;
  assign new_A7073_ = new_A7063_ ^ new_A7064_;
  assign new_A7074_ = new_A7075_ ^ new_A7065_;
  assign new_A7075_ = new_A7083_ & new_A7082_;
  assign new_A7076_ = new_A7081_ & new_A7065_;
  assign new_A7077_ = new_A7086_ & new_A7085_;
  assign new_A7078_ = new_A7084_ & new_A7065_;
  assign new_A7079_ = new_A7087_ | new_A7064_;
  assign new_A7080_ = ~new_A7065_ ^ new_A7077_;
  assign new_A7081_ = ~new_A7090_ | ~new_A7091_;
  assign new_A7082_ = new_A7066_ ^ new_A7073_;
  assign new_A7083_ = new_A7092_ & new_A7085_;
  assign new_A7084_ = ~new_A7094_ | ~new_A7093_;
  assign new_A7085_ = new_A7066_ | new_A7067_;
  assign new_A7086_ = new_A7066_ | new_A7073_;
  assign new_A7087_ = new_A7065_ & new_A7077_;
  assign new_A7088_ = ~new_A7064_ | ~new_A7065_;
  assign new_A7089_ = new_A7073_ & new_A7088_;
  assign new_A7090_ = ~new_A7089_ & ~new_A7073_;
  assign new_A7091_ = new_A7073_ | new_A7088_;
  assign new_A7092_ = ~new_A7066_ | ~new_A7067_;
  assign new_A7093_ = new_A7073_ | new_A7088_;
  assign new_A7094_ = ~new_A7073_ & ~new_A7095_;
  assign new_A7095_ = new_A7073_ & new_A7088_;
  assign new_A7096_ = new_B1887_;
  assign new_A7097_ = new_B1920_;
  assign new_A7098_ = new_B1953_;
  assign new_A7099_ = new_B1986_;
  assign new_A7100_ = new_B2019_;
  assign new_A7101_ = new_A7107_ & new_A7106_;
  assign new_A7102_ = new_A7109_ | new_A7108_;
  assign new_A7103_ = new_A7111_ | new_A7110_;
  assign new_A7104_ = new_A7106_ & new_A7112_;
  assign new_A7105_ = new_A7106_ & new_A7113_;
  assign new_A7106_ = new_A7096_ ^ new_A7097_;
  assign new_A7107_ = new_A7108_ ^ new_A7098_;
  assign new_A7108_ = new_A7116_ & new_A7115_;
  assign new_A7109_ = new_A7114_ & new_A7098_;
  assign new_A7110_ = new_A7119_ & new_A7118_;
  assign new_A7111_ = new_A7117_ & new_A7098_;
  assign new_A7112_ = new_A7120_ | new_A7097_;
  assign new_A7113_ = ~new_A7098_ ^ new_A7110_;
  assign new_A7114_ = ~new_A7123_ | ~new_A7124_;
  assign new_A7115_ = new_A7099_ ^ new_A7106_;
  assign new_A7116_ = new_A7125_ & new_A7118_;
  assign new_A7117_ = ~new_A7127_ | ~new_A7126_;
  assign new_A7118_ = new_A7099_ | new_A7100_;
  assign new_A7119_ = new_A7099_ | new_A7106_;
  assign new_A7120_ = new_A7098_ & new_A7110_;
  assign new_A7121_ = ~new_A7097_ | ~new_A7098_;
  assign new_A7122_ = new_A7106_ & new_A7121_;
  assign new_A7123_ = ~new_A7122_ & ~new_A7106_;
  assign new_A7124_ = new_A7106_ | new_A7121_;
  assign new_A7125_ = ~new_A7099_ | ~new_A7100_;
  assign new_A7126_ = new_A7106_ | new_A7121_;
  assign new_A7127_ = ~new_A7106_ & ~new_A7128_;
  assign new_A7128_ = new_A7106_ & new_A7121_;
  assign new_A7129_ = new_B2052_;
  assign new_A7130_ = new_B2085_;
  assign new_A7131_ = new_B2118_;
  assign new_A7132_ = new_B2151_;
  assign new_A7133_ = new_B2184_;
  assign new_A7134_ = new_A7140_ & new_A7139_;
  assign new_A7135_ = new_A7142_ | new_A7141_;
  assign new_A7136_ = new_A7144_ | new_A7143_;
  assign new_A7137_ = new_A7139_ & new_A7145_;
  assign new_A7138_ = new_A7139_ & new_A7146_;
  assign new_A7139_ = new_A7129_ ^ new_A7130_;
  assign new_A7140_ = new_A7141_ ^ new_A7131_;
  assign new_A7141_ = new_A7149_ & new_A7148_;
  assign new_A7142_ = new_A7147_ & new_A7131_;
  assign new_A7143_ = new_A7152_ & new_A7151_;
  assign new_A7144_ = new_A7150_ & new_A7131_;
  assign new_A7145_ = new_A7153_ | new_A7130_;
  assign new_A7146_ = ~new_A7131_ ^ new_A7143_;
  assign new_A7147_ = ~new_A7156_ | ~new_A7157_;
  assign new_A7148_ = new_A7132_ ^ new_A7139_;
  assign new_A7149_ = new_A7158_ & new_A7151_;
  assign new_A7150_ = ~new_A7160_ | ~new_A7159_;
  assign new_A7151_ = new_A7132_ | new_A7133_;
  assign new_A7152_ = new_A7132_ | new_A7139_;
  assign new_A7153_ = new_A7131_ & new_A7143_;
  assign new_A7154_ = ~new_A7130_ | ~new_A7131_;
  assign new_A7155_ = new_A7139_ & new_A7154_;
  assign new_A7156_ = ~new_A7155_ & ~new_A7139_;
  assign new_A7157_ = new_A7139_ | new_A7154_;
  assign new_A7158_ = ~new_A7132_ | ~new_A7133_;
  assign new_A7159_ = new_A7139_ | new_A7154_;
  assign new_A7160_ = ~new_A7139_ & ~new_A7161_;
  assign new_A7161_ = new_A7139_ & new_A7154_;
  assign new_A7162_ = new_B2217_;
  assign new_A7163_ = new_B2250_;
  assign new_A7164_ = new_B2283_;
  assign new_A7165_ = new_B2316_;
  assign new_A7166_ = new_B2349_;
  assign new_A7167_ = new_A7173_ & new_A7172_;
  assign new_A7168_ = new_A7175_ | new_A7174_;
  assign new_A7169_ = new_A7177_ | new_A7176_;
  assign new_A7170_ = new_A7172_ & new_A7178_;
  assign new_A7171_ = new_A7172_ & new_A7179_;
  assign new_A7172_ = new_A7162_ ^ new_A7163_;
  assign new_A7173_ = new_A7174_ ^ new_A7164_;
  assign new_A7174_ = new_A7182_ & new_A7181_;
  assign new_A7175_ = new_A7180_ & new_A7164_;
  assign new_A7176_ = new_A7185_ & new_A7184_;
  assign new_A7177_ = new_A7183_ & new_A7164_;
  assign new_A7178_ = new_A7186_ | new_A7163_;
  assign new_A7179_ = ~new_A7164_ ^ new_A7176_;
  assign new_A7180_ = ~new_A7189_ | ~new_A7190_;
  assign new_A7181_ = new_A7165_ ^ new_A7172_;
  assign new_A7182_ = new_A7191_ & new_A7184_;
  assign new_A7183_ = ~new_A7193_ | ~new_A7192_;
  assign new_A7184_ = new_A7165_ | new_A7166_;
  assign new_A7185_ = new_A7165_ | new_A7172_;
  assign new_A7186_ = new_A7164_ & new_A7176_;
  assign new_A7187_ = ~new_A7163_ | ~new_A7164_;
  assign new_A7188_ = new_A7172_ & new_A7187_;
  assign new_A7189_ = ~new_A7188_ & ~new_A7172_;
  assign new_A7190_ = new_A7172_ | new_A7187_;
  assign new_A7191_ = ~new_A7165_ | ~new_A7166_;
  assign new_A7192_ = new_A7172_ | new_A7187_;
  assign new_A7193_ = ~new_A7172_ & ~new_A7194_;
  assign new_A7194_ = new_A7172_ & new_A7187_;
  assign new_A7195_ = new_B2382_;
  assign new_A7196_ = new_B2415_;
  assign new_A7197_ = new_B2448_;
  assign new_A7198_ = new_B2481_;
  assign new_A7199_ = new_B2514_;
  assign new_A7200_ = new_A7206_ & new_A7205_;
  assign new_A7201_ = new_A7208_ | new_A7207_;
  assign new_A7202_ = new_A7210_ | new_A7209_;
  assign new_A7203_ = new_A7205_ & new_A7211_;
  assign new_A7204_ = new_A7205_ & new_A7212_;
  assign new_A7205_ = new_A7195_ ^ new_A7196_;
  assign new_A7206_ = new_A7207_ ^ new_A7197_;
  assign new_A7207_ = new_A7215_ & new_A7214_;
  assign new_A7208_ = new_A7213_ & new_A7197_;
  assign new_A7209_ = new_A7218_ & new_A7217_;
  assign new_A7210_ = new_A7216_ & new_A7197_;
  assign new_A7211_ = new_A7219_ | new_A7196_;
  assign new_A7212_ = ~new_A7197_ ^ new_A7209_;
  assign new_A7213_ = ~new_A7222_ | ~new_A7223_;
  assign new_A7214_ = new_A7198_ ^ new_A7205_;
  assign new_A7215_ = new_A7224_ & new_A7217_;
  assign new_A7216_ = ~new_A7226_ | ~new_A7225_;
  assign new_A7217_ = new_A7198_ | new_A7199_;
  assign new_A7218_ = new_A7198_ | new_A7205_;
  assign new_A7219_ = new_A7197_ & new_A7209_;
  assign new_A7220_ = ~new_A7196_ | ~new_A7197_;
  assign new_A7221_ = new_A7205_ & new_A7220_;
  assign new_A7222_ = ~new_A7221_ & ~new_A7205_;
  assign new_A7223_ = new_A7205_ | new_A7220_;
  assign new_A7224_ = ~new_A7198_ | ~new_A7199_;
  assign new_A7225_ = new_A7205_ | new_A7220_;
  assign new_A7226_ = ~new_A7205_ & ~new_A7227_;
  assign new_A7227_ = new_A7205_ & new_A7220_;
  assign new_A7228_ = new_B2547_;
  assign new_A7229_ = new_B2580_;
  assign new_A7230_ = new_B2613_;
  assign new_A7231_ = new_B2646_;
  assign new_A7232_ = new_B2679_;
  assign new_A7233_ = new_A7239_ & new_A7238_;
  assign new_A7234_ = new_A7241_ | new_A7240_;
  assign new_A7235_ = new_A7243_ | new_A7242_;
  assign new_A7236_ = new_A7238_ & new_A7244_;
  assign new_A7237_ = new_A7238_ & new_A7245_;
  assign new_A7238_ = new_A7228_ ^ new_A7229_;
  assign new_A7239_ = new_A7240_ ^ new_A7230_;
  assign new_A7240_ = new_A7248_ & new_A7247_;
  assign new_A7241_ = new_A7246_ & new_A7230_;
  assign new_A7242_ = new_A7251_ & new_A7250_;
  assign new_A7243_ = new_A7249_ & new_A7230_;
  assign new_A7244_ = new_A7252_ | new_A7229_;
  assign new_A7245_ = ~new_A7230_ ^ new_A7242_;
  assign new_A7246_ = ~new_A7255_ | ~new_A7256_;
  assign new_A7247_ = new_A7231_ ^ new_A7238_;
  assign new_A7248_ = new_A7257_ & new_A7250_;
  assign new_A7249_ = ~new_A7259_ | ~new_A7258_;
  assign new_A7250_ = new_A7231_ | new_A7232_;
  assign new_A7251_ = new_A7231_ | new_A7238_;
  assign new_A7252_ = new_A7230_ & new_A7242_;
  assign new_A7253_ = ~new_A7229_ | ~new_A7230_;
  assign new_A7254_ = new_A7238_ & new_A7253_;
  assign new_A7255_ = ~new_A7254_ & ~new_A7238_;
  assign new_A7256_ = new_A7238_ | new_A7253_;
  assign new_A7257_ = ~new_A7231_ | ~new_A7232_;
  assign new_A7258_ = new_A7238_ | new_A7253_;
  assign new_A7259_ = ~new_A7238_ & ~new_A7260_;
  assign new_A7260_ = new_A7238_ & new_A7253_;
  assign new_A7261_ = new_B2712_;
  assign new_A7262_ = new_B2745_;
  assign new_A7263_ = new_B2778_;
  assign new_A7264_ = new_B2811_;
  assign new_A7265_ = new_B2844_;
  assign new_A7266_ = new_A7272_ & new_A7271_;
  assign new_A7267_ = new_A7274_ | new_A7273_;
  assign new_A7268_ = new_A7276_ | new_A7275_;
  assign new_A7269_ = new_A7271_ & new_A7277_;
  assign new_A7270_ = new_A7271_ & new_A7278_;
  assign new_A7271_ = new_A7261_ ^ new_A7262_;
  assign new_A7272_ = new_A7273_ ^ new_A7263_;
  assign new_A7273_ = new_A7281_ & new_A7280_;
  assign new_A7274_ = new_A7279_ & new_A7263_;
  assign new_A7275_ = new_A7284_ & new_A7283_;
  assign new_A7276_ = new_A7282_ & new_A7263_;
  assign new_A7277_ = new_A7285_ | new_A7262_;
  assign new_A7278_ = ~new_A7263_ ^ new_A7275_;
  assign new_A7279_ = ~new_A7288_ | ~new_A7289_;
  assign new_A7280_ = new_A7264_ ^ new_A7271_;
  assign new_A7281_ = new_A7290_ & new_A7283_;
  assign new_A7282_ = ~new_A7292_ | ~new_A7291_;
  assign new_A7283_ = new_A7264_ | new_A7265_;
  assign new_A7284_ = new_A7264_ | new_A7271_;
  assign new_A7285_ = new_A7263_ & new_A7275_;
  assign new_A7286_ = ~new_A7262_ | ~new_A7263_;
  assign new_A7287_ = new_A7271_ & new_A7286_;
  assign new_A7288_ = ~new_A7287_ & ~new_A7271_;
  assign new_A7289_ = new_A7271_ | new_A7286_;
  assign new_A7290_ = ~new_A7264_ | ~new_A7265_;
  assign new_A7291_ = new_A7271_ | new_A7286_;
  assign new_A7292_ = ~new_A7271_ & ~new_A7293_;
  assign new_A7293_ = new_A7271_ & new_A7286_;
  assign new_A7294_ = new_B2877_;
  assign new_A7295_ = new_B2910_;
  assign new_A7296_ = new_B2943_;
  assign new_A7297_ = new_B2976_;
  assign new_A7298_ = new_B3009_;
  assign new_A7299_ = new_A7305_ & new_A7304_;
  assign new_A7300_ = new_A7307_ | new_A7306_;
  assign new_A7301_ = new_A7309_ | new_A7308_;
  assign new_A7302_ = new_A7304_ & new_A7310_;
  assign new_A7303_ = new_A7304_ & new_A7311_;
  assign new_A7304_ = new_A7294_ ^ new_A7295_;
  assign new_A7305_ = new_A7306_ ^ new_A7296_;
  assign new_A7306_ = new_A7314_ & new_A7313_;
  assign new_A7307_ = new_A7312_ & new_A7296_;
  assign new_A7308_ = new_A7317_ & new_A7316_;
  assign new_A7309_ = new_A7315_ & new_A7296_;
  assign new_A7310_ = new_A7318_ | new_A7295_;
  assign new_A7311_ = ~new_A7296_ ^ new_A7308_;
  assign new_A7312_ = ~new_A7321_ | ~new_A7322_;
  assign new_A7313_ = new_A7297_ ^ new_A7304_;
  assign new_A7314_ = new_A7323_ & new_A7316_;
  assign new_A7315_ = ~new_A7325_ | ~new_A7324_;
  assign new_A7316_ = new_A7297_ | new_A7298_;
  assign new_A7317_ = new_A7297_ | new_A7304_;
  assign new_A7318_ = new_A7296_ & new_A7308_;
  assign new_A7319_ = ~new_A7295_ | ~new_A7296_;
  assign new_A7320_ = new_A7304_ & new_A7319_;
  assign new_A7321_ = ~new_A7320_ & ~new_A7304_;
  assign new_A7322_ = new_A7304_ | new_A7319_;
  assign new_A7323_ = ~new_A7297_ | ~new_A7298_;
  assign new_A7324_ = new_A7304_ | new_A7319_;
  assign new_A7325_ = ~new_A7304_ & ~new_A7326_;
  assign new_A7326_ = new_A7304_ & new_A7319_;
  assign new_A7327_ = new_B3042_;
  assign new_A7328_ = new_B3075_;
  assign new_A7329_ = new_B3108_;
  assign new_A7330_ = new_B3141_;
  assign new_A7331_ = new_B3174_;
  assign new_A7332_ = new_A7338_ & new_A7337_;
  assign new_A7333_ = new_A7340_ | new_A7339_;
  assign new_A7334_ = new_A7342_ | new_A7341_;
  assign new_A7335_ = new_A7337_ & new_A7343_;
  assign new_A7336_ = new_A7337_ & new_A7344_;
  assign new_A7337_ = new_A7327_ ^ new_A7328_;
  assign new_A7338_ = new_A7339_ ^ new_A7329_;
  assign new_A7339_ = new_A7347_ & new_A7346_;
  assign new_A7340_ = new_A7345_ & new_A7329_;
  assign new_A7341_ = new_A7350_ & new_A7349_;
  assign new_A7342_ = new_A7348_ & new_A7329_;
  assign new_A7343_ = new_A7351_ | new_A7328_;
  assign new_A7344_ = ~new_A7329_ ^ new_A7341_;
  assign new_A7345_ = ~new_A7354_ | ~new_A7355_;
  assign new_A7346_ = new_A7330_ ^ new_A7337_;
  assign new_A7347_ = new_A7356_ & new_A7349_;
  assign new_A7348_ = ~new_A7358_ | ~new_A7357_;
  assign new_A7349_ = new_A7330_ | new_A7331_;
  assign new_A7350_ = new_A7330_ | new_A7337_;
  assign new_A7351_ = new_A7329_ & new_A7341_;
  assign new_A7352_ = ~new_A7328_ | ~new_A7329_;
  assign new_A7353_ = new_A7337_ & new_A7352_;
  assign new_A7354_ = ~new_A7353_ & ~new_A7337_;
  assign new_A7355_ = new_A7337_ | new_A7352_;
  assign new_A7356_ = ~new_A7330_ | ~new_A7331_;
  assign new_A7357_ = new_A7337_ | new_A7352_;
  assign new_A7358_ = ~new_A7337_ & ~new_A7359_;
  assign new_A7359_ = new_A7337_ & new_A7352_;
  assign new_A7360_ = new_B3207_;
  assign new_A7361_ = new_B3240_;
  assign new_A7362_ = new_B3273_;
  assign new_A7363_ = new_B3306_;
  assign new_A7364_ = new_B3339_;
  assign new_A7365_ = new_A7371_ & new_A7370_;
  assign new_A7366_ = new_A7373_ | new_A7372_;
  assign new_A7367_ = new_A7375_ | new_A7374_;
  assign new_A7368_ = new_A7370_ & new_A7376_;
  assign new_A7369_ = new_A7370_ & new_A7377_;
  assign new_A7370_ = new_A7360_ ^ new_A7361_;
  assign new_A7371_ = new_A7372_ ^ new_A7362_;
  assign new_A7372_ = new_A7380_ & new_A7379_;
  assign new_A7373_ = new_A7378_ & new_A7362_;
  assign new_A7374_ = new_A7383_ & new_A7382_;
  assign new_A7375_ = new_A7381_ & new_A7362_;
  assign new_A7376_ = new_A7384_ | new_A7361_;
  assign new_A7377_ = ~new_A7362_ ^ new_A7374_;
  assign new_A7378_ = ~new_A7387_ | ~new_A7388_;
  assign new_A7379_ = new_A7363_ ^ new_A7370_;
  assign new_A7380_ = new_A7389_ & new_A7382_;
  assign new_A7381_ = ~new_A7391_ | ~new_A7390_;
  assign new_A7382_ = new_A7363_ | new_A7364_;
  assign new_A7383_ = new_A7363_ | new_A7370_;
  assign new_A7384_ = new_A7362_ & new_A7374_;
  assign new_A7385_ = ~new_A7361_ | ~new_A7362_;
  assign new_A7386_ = new_A7370_ & new_A7385_;
  assign new_A7387_ = ~new_A7386_ & ~new_A7370_;
  assign new_A7388_ = new_A7370_ | new_A7385_;
  assign new_A7389_ = ~new_A7363_ | ~new_A7364_;
  assign new_A7390_ = new_A7370_ | new_A7385_;
  assign new_A7391_ = ~new_A7370_ & ~new_A7392_;
  assign new_A7392_ = new_A7370_ & new_A7385_;
  assign new_A7393_ = new_B3372_;
  assign new_A7394_ = new_B3405_;
  assign new_A7395_ = new_B3438_;
  assign new_A7396_ = new_B3471_;
  assign new_A7397_ = new_B3504_;
  assign new_A7398_ = new_A7404_ & new_A7403_;
  assign new_A7399_ = new_A7406_ | new_A7405_;
  assign new_A7400_ = new_A7408_ | new_A7407_;
  assign new_A7401_ = new_A7403_ & new_A7409_;
  assign new_A7402_ = new_A7403_ & new_A7410_;
  assign new_A7403_ = new_A7393_ ^ new_A7394_;
  assign new_A7404_ = new_A7405_ ^ new_A7395_;
  assign new_A7405_ = new_A7413_ & new_A7412_;
  assign new_A7406_ = new_A7411_ & new_A7395_;
  assign new_A7407_ = new_A7416_ & new_A7415_;
  assign new_A7408_ = new_A7414_ & new_A7395_;
  assign new_A7409_ = new_A7417_ | new_A7394_;
  assign new_A7410_ = ~new_A7395_ ^ new_A7407_;
  assign new_A7411_ = ~new_A7420_ | ~new_A7421_;
  assign new_A7412_ = new_A7396_ ^ new_A7403_;
  assign new_A7413_ = new_A7422_ & new_A7415_;
  assign new_A7414_ = ~new_A7424_ | ~new_A7423_;
  assign new_A7415_ = new_A7396_ | new_A7397_;
  assign new_A7416_ = new_A7396_ | new_A7403_;
  assign new_A7417_ = new_A7395_ & new_A7407_;
  assign new_A7418_ = ~new_A7394_ | ~new_A7395_;
  assign new_A7419_ = new_A7403_ & new_A7418_;
  assign new_A7420_ = ~new_A7419_ & ~new_A7403_;
  assign new_A7421_ = new_A7403_ | new_A7418_;
  assign new_A7422_ = ~new_A7396_ | ~new_A7397_;
  assign new_A7423_ = new_A7403_ | new_A7418_;
  assign new_A7424_ = ~new_A7403_ & ~new_A7425_;
  assign new_A7425_ = new_A7403_ & new_A7418_;
  assign new_A7426_ = new_B3537_;
  assign new_A7427_ = new_B3570_;
  assign new_A7428_ = new_B3603_;
  assign new_A7429_ = new_B3636_;
  assign new_A7430_ = new_B3669_;
  assign new_A7431_ = new_A7437_ & new_A7436_;
  assign new_A7432_ = new_A7439_ | new_A7438_;
  assign new_A7433_ = new_A7441_ | new_A7440_;
  assign new_A7434_ = new_A7436_ & new_A7442_;
  assign new_A7435_ = new_A7436_ & new_A7443_;
  assign new_A7436_ = new_A7426_ ^ new_A7427_;
  assign new_A7437_ = new_A7438_ ^ new_A7428_;
  assign new_A7438_ = new_A7446_ & new_A7445_;
  assign new_A7439_ = new_A7444_ & new_A7428_;
  assign new_A7440_ = new_A7449_ & new_A7448_;
  assign new_A7441_ = new_A7447_ & new_A7428_;
  assign new_A7442_ = new_A7450_ | new_A7427_;
  assign new_A7443_ = ~new_A7428_ ^ new_A7440_;
  assign new_A7444_ = ~new_A7453_ | ~new_A7454_;
  assign new_A7445_ = new_A7429_ ^ new_A7436_;
  assign new_A7446_ = new_A7455_ & new_A7448_;
  assign new_A7447_ = ~new_A7457_ | ~new_A7456_;
  assign new_A7448_ = new_A7429_ | new_A7430_;
  assign new_A7449_ = new_A7429_ | new_A7436_;
  assign new_A7450_ = new_A7428_ & new_A7440_;
  assign new_A7451_ = ~new_A7427_ | ~new_A7428_;
  assign new_A7452_ = new_A7436_ & new_A7451_;
  assign new_A7453_ = ~new_A7452_ & ~new_A7436_;
  assign new_A7454_ = new_A7436_ | new_A7451_;
  assign new_A7455_ = ~new_A7429_ | ~new_A7430_;
  assign new_A7456_ = new_A7436_ | new_A7451_;
  assign new_A7457_ = ~new_A7436_ & ~new_A7458_;
  assign new_A7458_ = new_A7436_ & new_A7451_;
  assign new_A7459_ = new_B3702_;
  assign new_A7460_ = new_B3735_;
  assign new_A7461_ = new_B3768_;
  assign new_A7462_ = new_B3801_;
  assign new_A7463_ = new_B3834_;
  assign new_A7464_ = new_A7470_ & new_A7469_;
  assign new_A7465_ = new_A7472_ | new_A7471_;
  assign new_A7466_ = new_A7474_ | new_A7473_;
  assign new_A7467_ = new_A7469_ & new_A7475_;
  assign new_A7468_ = new_A7469_ & new_A7476_;
  assign new_A7469_ = new_A7459_ ^ new_A7460_;
  assign new_A7470_ = new_A7471_ ^ new_A7461_;
  assign new_A7471_ = new_A7479_ & new_A7478_;
  assign new_A7472_ = new_A7477_ & new_A7461_;
  assign new_A7473_ = new_A7482_ & new_A7481_;
  assign new_A7474_ = new_A7480_ & new_A7461_;
  assign new_A7475_ = new_A7483_ | new_A7460_;
  assign new_A7476_ = ~new_A7461_ ^ new_A7473_;
  assign new_A7477_ = ~new_A7486_ | ~new_A7487_;
  assign new_A7478_ = new_A7462_ ^ new_A7469_;
  assign new_A7479_ = new_A7488_ & new_A7481_;
  assign new_A7480_ = ~new_A7490_ | ~new_A7489_;
  assign new_A7481_ = new_A7462_ | new_A7463_;
  assign new_A7482_ = new_A7462_ | new_A7469_;
  assign new_A7483_ = new_A7461_ & new_A7473_;
  assign new_A7484_ = ~new_A7460_ | ~new_A7461_;
  assign new_A7485_ = new_A7469_ & new_A7484_;
  assign new_A7486_ = ~new_A7485_ & ~new_A7469_;
  assign new_A7487_ = new_A7469_ | new_A7484_;
  assign new_A7488_ = ~new_A7462_ | ~new_A7463_;
  assign new_A7489_ = new_A7469_ | new_A7484_;
  assign new_A7490_ = ~new_A7469_ & ~new_A7491_;
  assign new_A7491_ = new_A7469_ & new_A7484_;
  assign new_A7492_ = new_B3867_;
  assign new_A7493_ = new_B3900_;
  assign new_A7494_ = new_B3933_;
  assign new_A7495_ = new_B3966_;
  assign new_A7496_ = new_B3999_;
  assign new_A7497_ = new_A7503_ & new_A7502_;
  assign new_A7498_ = new_A7505_ | new_A7504_;
  assign new_A7499_ = new_A7507_ | new_A7506_;
  assign new_A7500_ = new_A7502_ & new_A7508_;
  assign new_A7501_ = new_A7502_ & new_A7509_;
  assign new_A7502_ = new_A7492_ ^ new_A7493_;
  assign new_A7503_ = new_A7504_ ^ new_A7494_;
  assign new_A7504_ = new_A7512_ & new_A7511_;
  assign new_A7505_ = new_A7510_ & new_A7494_;
  assign new_A7506_ = new_A7515_ & new_A7514_;
  assign new_A7507_ = new_A7513_ & new_A7494_;
  assign new_A7508_ = new_A7516_ | new_A7493_;
  assign new_A7509_ = ~new_A7494_ ^ new_A7506_;
  assign new_A7510_ = ~new_A7519_ | ~new_A7520_;
  assign new_A7511_ = new_A7495_ ^ new_A7502_;
  assign new_A7512_ = new_A7521_ & new_A7514_;
  assign new_A7513_ = ~new_A7523_ | ~new_A7522_;
  assign new_A7514_ = new_A7495_ | new_A7496_;
  assign new_A7515_ = new_A7495_ | new_A7502_;
  assign new_A7516_ = new_A7494_ & new_A7506_;
  assign new_A7517_ = ~new_A7493_ | ~new_A7494_;
  assign new_A7518_ = new_A7502_ & new_A7517_;
  assign new_A7519_ = ~new_A7518_ & ~new_A7502_;
  assign new_A7520_ = new_A7502_ | new_A7517_;
  assign new_A7521_ = ~new_A7495_ | ~new_A7496_;
  assign new_A7522_ = new_A7502_ | new_A7517_;
  assign new_A7523_ = ~new_A7502_ & ~new_A7524_;
  assign new_A7524_ = new_A7502_ & new_A7517_;
  assign new_A7525_ = new_B4032_;
  assign new_A7526_ = new_B4065_;
  assign new_A7527_ = new_B4098_;
  assign new_A7528_ = new_B4131_;
  assign new_A7529_ = new_B4164_;
  assign new_A7530_ = new_A7536_ & new_A7535_;
  assign new_A7531_ = new_A7538_ | new_A7537_;
  assign new_A7532_ = new_A7540_ | new_A7539_;
  assign new_A7533_ = new_A7535_ & new_A7541_;
  assign new_A7534_ = new_A7535_ & new_A7542_;
  assign new_A7535_ = new_A7525_ ^ new_A7526_;
  assign new_A7536_ = new_A7537_ ^ new_A7527_;
  assign new_A7537_ = new_A7545_ & new_A7544_;
  assign new_A7538_ = new_A7543_ & new_A7527_;
  assign new_A7539_ = new_A7548_ & new_A7547_;
  assign new_A7540_ = new_A7546_ & new_A7527_;
  assign new_A7541_ = new_A7549_ | new_A7526_;
  assign new_A7542_ = ~new_A7527_ ^ new_A7539_;
  assign new_A7543_ = ~new_A7552_ | ~new_A7553_;
  assign new_A7544_ = new_A7528_ ^ new_A7535_;
  assign new_A7545_ = new_A7554_ & new_A7547_;
  assign new_A7546_ = ~new_A7556_ | ~new_A7555_;
  assign new_A7547_ = new_A7528_ | new_A7529_;
  assign new_A7548_ = new_A7528_ | new_A7535_;
  assign new_A7549_ = new_A7527_ & new_A7539_;
  assign new_A7550_ = ~new_A7526_ | ~new_A7527_;
  assign new_A7551_ = new_A7535_ & new_A7550_;
  assign new_A7552_ = ~new_A7551_ & ~new_A7535_;
  assign new_A7553_ = new_A7535_ | new_A7550_;
  assign new_A7554_ = ~new_A7528_ | ~new_A7529_;
  assign new_A7555_ = new_A7535_ | new_A7550_;
  assign new_A7556_ = ~new_A7535_ & ~new_A7557_;
  assign new_A7557_ = new_A7535_ & new_A7550_;
  assign new_A7558_ = new_B4197_;
  assign new_A7559_ = new_B4230_;
  assign new_A7560_ = new_B4263_;
  assign new_A7561_ = new_B4296_;
  assign new_A7562_ = new_B4329_;
  assign new_A7563_ = new_A7569_ & new_A7568_;
  assign new_A7564_ = new_A7571_ | new_A7570_;
  assign new_A7565_ = new_A7573_ | new_A7572_;
  assign new_A7566_ = new_A7568_ & new_A7574_;
  assign new_A7567_ = new_A7568_ & new_A7575_;
  assign new_A7568_ = new_A7558_ ^ new_A7559_;
  assign new_A7569_ = new_A7570_ ^ new_A7560_;
  assign new_A7570_ = new_A7578_ & new_A7577_;
  assign new_A7571_ = new_A7576_ & new_A7560_;
  assign new_A7572_ = new_A7581_ & new_A7580_;
  assign new_A7573_ = new_A7579_ & new_A7560_;
  assign new_A7574_ = new_A7582_ | new_A7559_;
  assign new_A7575_ = ~new_A7560_ ^ new_A7572_;
  assign new_A7576_ = ~new_A7585_ | ~new_A7586_;
  assign new_A7577_ = new_A7561_ ^ new_A7568_;
  assign new_A7578_ = new_A7587_ & new_A7580_;
  assign new_A7579_ = ~new_A7589_ | ~new_A7588_;
  assign new_A7580_ = new_A7561_ | new_A7562_;
  assign new_A7581_ = new_A7561_ | new_A7568_;
  assign new_A7582_ = new_A7560_ & new_A7572_;
  assign new_A7583_ = ~new_A7559_ | ~new_A7560_;
  assign new_A7584_ = new_A7568_ & new_A7583_;
  assign new_A7585_ = ~new_A7584_ & ~new_A7568_;
  assign new_A7586_ = new_A7568_ | new_A7583_;
  assign new_A7587_ = ~new_A7561_ | ~new_A7562_;
  assign new_A7588_ = new_A7568_ | new_A7583_;
  assign new_A7589_ = ~new_A7568_ & ~new_A7590_;
  assign new_A7590_ = new_A7568_ & new_A7583_;
  assign new_A7591_ = new_B4362_;
  assign new_A7592_ = new_B4395_;
  assign new_A7593_ = new_B4428_;
  assign new_A7594_ = new_B4461_;
  assign new_A7595_ = new_B4494_;
  assign new_A7596_ = new_A7602_ & new_A7601_;
  assign new_A7597_ = new_A7604_ | new_A7603_;
  assign new_A7598_ = new_A7606_ | new_A7605_;
  assign new_A7599_ = new_A7601_ & new_A7607_;
  assign new_A7600_ = new_A7601_ & new_A7608_;
  assign new_A7601_ = new_A7591_ ^ new_A7592_;
  assign new_A7602_ = new_A7603_ ^ new_A7593_;
  assign new_A7603_ = new_A7611_ & new_A7610_;
  assign new_A7604_ = new_A7609_ & new_A7593_;
  assign new_A7605_ = new_A7614_ & new_A7613_;
  assign new_A7606_ = new_A7612_ & new_A7593_;
  assign new_A7607_ = new_A7615_ | new_A7592_;
  assign new_A7608_ = ~new_A7593_ ^ new_A7605_;
  assign new_A7609_ = ~new_A7618_ | ~new_A7619_;
  assign new_A7610_ = new_A7594_ ^ new_A7601_;
  assign new_A7611_ = new_A7620_ & new_A7613_;
  assign new_A7612_ = ~new_A7622_ | ~new_A7621_;
  assign new_A7613_ = new_A7594_ | new_A7595_;
  assign new_A7614_ = new_A7594_ | new_A7601_;
  assign new_A7615_ = new_A7593_ & new_A7605_;
  assign new_A7616_ = ~new_A7592_ | ~new_A7593_;
  assign new_A7617_ = new_A7601_ & new_A7616_;
  assign new_A7618_ = ~new_A7617_ & ~new_A7601_;
  assign new_A7619_ = new_A7601_ | new_A7616_;
  assign new_A7620_ = ~new_A7594_ | ~new_A7595_;
  assign new_A7621_ = new_A7601_ | new_A7616_;
  assign new_A7622_ = ~new_A7601_ & ~new_A7623_;
  assign new_A7623_ = new_A7601_ & new_A7616_;
  assign new_A7624_ = new_B4527_;
  assign new_A7625_ = new_B4560_;
  assign new_A7626_ = new_B4593_;
  assign new_A7627_ = new_B4626_;
  assign new_A7628_ = new_B4659_;
  assign new_A7629_ = new_A7635_ & new_A7634_;
  assign new_A7630_ = new_A7637_ | new_A7636_;
  assign new_A7631_ = new_A7639_ | new_A7638_;
  assign new_A7632_ = new_A7634_ & new_A7640_;
  assign new_A7633_ = new_A7634_ & new_A7641_;
  assign new_A7634_ = new_A7624_ ^ new_A7625_;
  assign new_A7635_ = new_A7636_ ^ new_A7626_;
  assign new_A7636_ = new_A7644_ & new_A7643_;
  assign new_A7637_ = new_A7642_ & new_A7626_;
  assign new_A7638_ = new_A7647_ & new_A7646_;
  assign new_A7639_ = new_A7645_ & new_A7626_;
  assign new_A7640_ = new_A7648_ | new_A7625_;
  assign new_A7641_ = ~new_A7626_ ^ new_A7638_;
  assign new_A7642_ = ~new_A7651_ | ~new_A7652_;
  assign new_A7643_ = new_A7627_ ^ new_A7634_;
  assign new_A7644_ = new_A7653_ & new_A7646_;
  assign new_A7645_ = ~new_A7655_ | ~new_A7654_;
  assign new_A7646_ = new_A7627_ | new_A7628_;
  assign new_A7647_ = new_A7627_ | new_A7634_;
  assign new_A7648_ = new_A7626_ & new_A7638_;
  assign new_A7649_ = ~new_A7625_ | ~new_A7626_;
  assign new_A7650_ = new_A7634_ & new_A7649_;
  assign new_A7651_ = ~new_A7650_ & ~new_A7634_;
  assign new_A7652_ = new_A7634_ | new_A7649_;
  assign new_A7653_ = ~new_A7627_ | ~new_A7628_;
  assign new_A7654_ = new_A7634_ | new_A7649_;
  assign new_A7655_ = ~new_A7634_ & ~new_A7656_;
  assign new_A7656_ = new_A7634_ & new_A7649_;
  assign new_A7657_ = new_B4692_;
  assign new_A7658_ = new_B4725_;
  assign new_A7659_ = new_B4758_;
  assign new_A7660_ = new_B4791_;
  assign new_A7661_ = new_B4824_;
  assign new_A7662_ = new_A7668_ & new_A7667_;
  assign new_A7663_ = new_A7670_ | new_A7669_;
  assign new_A7664_ = new_A7672_ | new_A7671_;
  assign new_A7665_ = new_A7667_ & new_A7673_;
  assign new_A7666_ = new_A7667_ & new_A7674_;
  assign new_A7667_ = new_A7657_ ^ new_A7658_;
  assign new_A7668_ = new_A7669_ ^ new_A7659_;
  assign new_A7669_ = new_A7677_ & new_A7676_;
  assign new_A7670_ = new_A7675_ & new_A7659_;
  assign new_A7671_ = new_A7680_ & new_A7679_;
  assign new_A7672_ = new_A7678_ & new_A7659_;
  assign new_A7673_ = new_A7681_ | new_A7658_;
  assign new_A7674_ = ~new_A7659_ ^ new_A7671_;
  assign new_A7675_ = ~new_A7684_ | ~new_A7685_;
  assign new_A7676_ = new_A7660_ ^ new_A7667_;
  assign new_A7677_ = new_A7686_ & new_A7679_;
  assign new_A7678_ = ~new_A7688_ | ~new_A7687_;
  assign new_A7679_ = new_A7660_ | new_A7661_;
  assign new_A7680_ = new_A7660_ | new_A7667_;
  assign new_A7681_ = new_A7659_ & new_A7671_;
  assign new_A7682_ = ~new_A7658_ | ~new_A7659_;
  assign new_A7683_ = new_A7667_ & new_A7682_;
  assign new_A7684_ = ~new_A7683_ & ~new_A7667_;
  assign new_A7685_ = new_A7667_ | new_A7682_;
  assign new_A7686_ = ~new_A7660_ | ~new_A7661_;
  assign new_A7687_ = new_A7667_ | new_A7682_;
  assign new_A7688_ = ~new_A7667_ & ~new_A7689_;
  assign new_A7689_ = new_A7667_ & new_A7682_;
  assign new_A7690_ = new_B4857_;
  assign new_A7691_ = new_B4890_;
  assign new_A7692_ = new_B4923_;
  assign new_A7693_ = new_B4956_;
  assign new_A7694_ = new_B4989_;
  assign new_A7695_ = new_A7701_ & new_A7700_;
  assign new_A7696_ = new_A7703_ | new_A7702_;
  assign new_A7697_ = new_A7705_ | new_A7704_;
  assign new_A7698_ = new_A7700_ & new_A7706_;
  assign new_A7699_ = new_A7700_ & new_A7707_;
  assign new_A7700_ = new_A7690_ ^ new_A7691_;
  assign new_A7701_ = new_A7702_ ^ new_A7692_;
  assign new_A7702_ = new_A7710_ & new_A7709_;
  assign new_A7703_ = new_A7708_ & new_A7692_;
  assign new_A7704_ = new_A7713_ & new_A7712_;
  assign new_A7705_ = new_A7711_ & new_A7692_;
  assign new_A7706_ = new_A7714_ | new_A7691_;
  assign new_A7707_ = ~new_A7692_ ^ new_A7704_;
  assign new_A7708_ = ~new_A7717_ | ~new_A7718_;
  assign new_A7709_ = new_A7693_ ^ new_A7700_;
  assign new_A7710_ = new_A7719_ & new_A7712_;
  assign new_A7711_ = ~new_A7721_ | ~new_A7720_;
  assign new_A7712_ = new_A7693_ | new_A7694_;
  assign new_A7713_ = new_A7693_ | new_A7700_;
  assign new_A7714_ = new_A7692_ & new_A7704_;
  assign new_A7715_ = ~new_A7691_ | ~new_A7692_;
  assign new_A7716_ = new_A7700_ & new_A7715_;
  assign new_A7717_ = ~new_A7716_ & ~new_A7700_;
  assign new_A7718_ = new_A7700_ | new_A7715_;
  assign new_A7719_ = ~new_A7693_ | ~new_A7694_;
  assign new_A7720_ = new_A7700_ | new_A7715_;
  assign new_A7721_ = ~new_A7700_ & ~new_A7722_;
  assign new_A7722_ = new_A7700_ & new_A7715_;
  assign new_A7723_ = new_B5022_;
  assign new_A7724_ = new_B5055_;
  assign new_A7725_ = new_B5088_;
  assign new_A7726_ = new_B5121_;
  assign new_A7727_ = new_B5154_;
  assign new_A7728_ = new_A7734_ & new_A7733_;
  assign new_A7729_ = new_A7736_ | new_A7735_;
  assign new_A7730_ = new_A7738_ | new_A7737_;
  assign new_A7731_ = new_A7733_ & new_A7739_;
  assign new_A7732_ = new_A7733_ & new_A7740_;
  assign new_A7733_ = new_A7723_ ^ new_A7724_;
  assign new_A7734_ = new_A7735_ ^ new_A7725_;
  assign new_A7735_ = new_A7743_ & new_A7742_;
  assign new_A7736_ = new_A7741_ & new_A7725_;
  assign new_A7737_ = new_A7746_ & new_A7745_;
  assign new_A7738_ = new_A7744_ & new_A7725_;
  assign new_A7739_ = new_A7747_ | new_A7724_;
  assign new_A7740_ = ~new_A7725_ ^ new_A7737_;
  assign new_A7741_ = ~new_A7750_ | ~new_A7751_;
  assign new_A7742_ = new_A7726_ ^ new_A7733_;
  assign new_A7743_ = new_A7752_ & new_A7745_;
  assign new_A7744_ = ~new_A7754_ | ~new_A7753_;
  assign new_A7745_ = new_A7726_ | new_A7727_;
  assign new_A7746_ = new_A7726_ | new_A7733_;
  assign new_A7747_ = new_A7725_ & new_A7737_;
  assign new_A7748_ = ~new_A7724_ | ~new_A7725_;
  assign new_A7749_ = new_A7733_ & new_A7748_;
  assign new_A7750_ = ~new_A7749_ & ~new_A7733_;
  assign new_A7751_ = new_A7733_ | new_A7748_;
  assign new_A7752_ = ~new_A7726_ | ~new_A7727_;
  assign new_A7753_ = new_A7733_ | new_A7748_;
  assign new_A7754_ = ~new_A7733_ & ~new_A7755_;
  assign new_A7755_ = new_A7733_ & new_A7748_;
  assign new_A7756_ = new_B1065_;
  assign new_A7757_ = new_B1096_;
  assign new_A7758_ = new_B1129_;
  assign new_A7759_ = new_B1162_;
  assign new_A7760_ = new_B1195_;
  assign new_A7761_ = new_A7767_ & new_A7766_;
  assign new_A7762_ = new_A7769_ | new_A7768_;
  assign new_A7763_ = new_A7771_ | new_A7770_;
  assign new_A7764_ = new_A7766_ & new_A7772_;
  assign new_A7765_ = new_A7766_ & new_A7773_;
  assign new_A7766_ = new_A7756_ ^ new_A7757_;
  assign new_A7767_ = new_A7768_ ^ new_A7758_;
  assign new_A7768_ = new_A7776_ & new_A7775_;
  assign new_A7769_ = new_A7774_ & new_A7758_;
  assign new_A7770_ = new_A7779_ & new_A7778_;
  assign new_A7771_ = new_A7777_ & new_A7758_;
  assign new_A7772_ = new_A7780_ | new_A7757_;
  assign new_A7773_ = ~new_A7758_ ^ new_A7770_;
  assign new_A7774_ = ~new_A7783_ | ~new_A7784_;
  assign new_A7775_ = new_A7759_ ^ new_A7766_;
  assign new_A7776_ = new_A7785_ & new_A7778_;
  assign new_A7777_ = ~new_A7787_ | ~new_A7786_;
  assign new_A7778_ = new_A7759_ | new_A7760_;
  assign new_A7779_ = new_A7759_ | new_A7766_;
  assign new_A7780_ = new_A7758_ & new_A7770_;
  assign new_A7781_ = ~new_A7757_ | ~new_A7758_;
  assign new_A7782_ = new_A7766_ & new_A7781_;
  assign new_A7783_ = ~new_A7782_ & ~new_A7766_;
  assign new_A7784_ = new_A7766_ | new_A7781_;
  assign new_A7785_ = ~new_A7759_ | ~new_A7760_;
  assign new_A7786_ = new_A7766_ | new_A7781_;
  assign new_A7787_ = ~new_A7766_ & ~new_A7788_;
  assign new_A7788_ = new_A7766_ & new_A7781_;
  assign new_A7789_ = new_B1228_;
  assign new_A7790_ = new_B1261_;
  assign new_A7791_ = new_B1294_;
  assign new_A7792_ = new_B1327_;
  assign new_A7793_ = new_B1360_;
  assign new_A7794_ = new_A7800_ & new_A7799_;
  assign new_A7795_ = new_A7802_ | new_A7801_;
  assign new_A7796_ = new_A7804_ | new_A7803_;
  assign new_A7797_ = new_A7799_ & new_A7805_;
  assign new_A7798_ = new_A7799_ & new_A7806_;
  assign new_A7799_ = new_A7789_ ^ new_A7790_;
  assign new_A7800_ = new_A7801_ ^ new_A7791_;
  assign new_A7801_ = new_A7809_ & new_A7808_;
  assign new_A7802_ = new_A7807_ & new_A7791_;
  assign new_A7803_ = new_A7812_ & new_A7811_;
  assign new_A7804_ = new_A7810_ & new_A7791_;
  assign new_A7805_ = new_A7813_ | new_A7790_;
  assign new_A7806_ = ~new_A7791_ ^ new_A7803_;
  assign new_A7807_ = ~new_A7816_ | ~new_A7817_;
  assign new_A7808_ = new_A7792_ ^ new_A7799_;
  assign new_A7809_ = new_A7818_ & new_A7811_;
  assign new_A7810_ = ~new_A7820_ | ~new_A7819_;
  assign new_A7811_ = new_A7792_ | new_A7793_;
  assign new_A7812_ = new_A7792_ | new_A7799_;
  assign new_A7813_ = new_A7791_ & new_A7803_;
  assign new_A7814_ = ~new_A7790_ | ~new_A7791_;
  assign new_A7815_ = new_A7799_ & new_A7814_;
  assign new_A7816_ = ~new_A7815_ & ~new_A7799_;
  assign new_A7817_ = new_A7799_ | new_A7814_;
  assign new_A7818_ = ~new_A7792_ | ~new_A7793_;
  assign new_A7819_ = new_A7799_ | new_A7814_;
  assign new_A7820_ = ~new_A7799_ & ~new_A7821_;
  assign new_A7821_ = new_A7799_ & new_A7814_;
  assign new_A7822_ = new_B1393_;
  assign new_A7823_ = new_B1426_;
  assign new_A7824_ = new_B1459_;
  assign new_A7825_ = new_B1492_;
  assign new_A7826_ = new_B1525_;
  assign new_A7827_ = new_A7833_ & new_A7832_;
  assign new_A7828_ = new_A7835_ | new_A7834_;
  assign new_A7829_ = new_A7837_ | new_A7836_;
  assign new_A7830_ = new_A7832_ & new_A7838_;
  assign new_A7831_ = new_A7832_ & new_A7839_;
  assign new_A7832_ = new_A7822_ ^ new_A7823_;
  assign new_A7833_ = new_A7834_ ^ new_A7824_;
  assign new_A7834_ = new_A7842_ & new_A7841_;
  assign new_A7835_ = new_A7840_ & new_A7824_;
  assign new_A7836_ = new_A7845_ & new_A7844_;
  assign new_A7837_ = new_A7843_ & new_A7824_;
  assign new_A7838_ = new_A7846_ | new_A7823_;
  assign new_A7839_ = ~new_A7824_ ^ new_A7836_;
  assign new_A7840_ = ~new_A7849_ | ~new_A7850_;
  assign new_A7841_ = new_A7825_ ^ new_A7832_;
  assign new_A7842_ = new_A7851_ & new_A7844_;
  assign new_A7843_ = ~new_A7853_ | ~new_A7852_;
  assign new_A7844_ = new_A7825_ | new_A7826_;
  assign new_A7845_ = new_A7825_ | new_A7832_;
  assign new_A7846_ = new_A7824_ & new_A7836_;
  assign new_A7847_ = ~new_A7823_ | ~new_A7824_;
  assign new_A7848_ = new_A7832_ & new_A7847_;
  assign new_A7849_ = ~new_A7848_ & ~new_A7832_;
  assign new_A7850_ = new_A7832_ | new_A7847_;
  assign new_A7851_ = ~new_A7825_ | ~new_A7826_;
  assign new_A7852_ = new_A7832_ | new_A7847_;
  assign new_A7853_ = ~new_A7832_ & ~new_A7854_;
  assign new_A7854_ = new_A7832_ & new_A7847_;
  assign new_A7855_ = new_B1558_;
  assign new_A7856_ = new_B1591_;
  assign new_A7857_ = new_B1624_;
  assign new_A7858_ = new_B1657_;
  assign new_A7859_ = new_B1690_;
  assign new_A7860_ = new_A7866_ & new_A7865_;
  assign new_A7861_ = new_A7868_ | new_A7867_;
  assign new_A7862_ = new_A7870_ | new_A7869_;
  assign new_A7863_ = new_A7865_ & new_A7871_;
  assign new_A7864_ = new_A7865_ & new_A7872_;
  assign new_A7865_ = new_A7855_ ^ new_A7856_;
  assign new_A7866_ = new_A7867_ ^ new_A7857_;
  assign new_A7867_ = new_A7875_ & new_A7874_;
  assign new_A7868_ = new_A7873_ & new_A7857_;
  assign new_A7869_ = new_A7878_ & new_A7877_;
  assign new_A7870_ = new_A7876_ & new_A7857_;
  assign new_A7871_ = new_A7879_ | new_A7856_;
  assign new_A7872_ = ~new_A7857_ ^ new_A7869_;
  assign new_A7873_ = ~new_A7882_ | ~new_A7883_;
  assign new_A7874_ = new_A7858_ ^ new_A7865_;
  assign new_A7875_ = new_A7884_ & new_A7877_;
  assign new_A7876_ = ~new_A7886_ | ~new_A7885_;
  assign new_A7877_ = new_A7858_ | new_A7859_;
  assign new_A7878_ = new_A7858_ | new_A7865_;
  assign new_A7879_ = new_A7857_ & new_A7869_;
  assign new_A7880_ = ~new_A7856_ | ~new_A7857_;
  assign new_A7881_ = new_A7865_ & new_A7880_;
  assign new_A7882_ = ~new_A7881_ & ~new_A7865_;
  assign new_A7883_ = new_A7865_ | new_A7880_;
  assign new_A7884_ = ~new_A7858_ | ~new_A7859_;
  assign new_A7885_ = new_A7865_ | new_A7880_;
  assign new_A7886_ = ~new_A7865_ & ~new_A7887_;
  assign new_A7887_ = new_A7865_ & new_A7880_;
  assign new_A7888_ = new_B1723_;
  assign new_A7889_ = new_B1756_;
  assign new_A7890_ = new_B1789_;
  assign new_A7891_ = new_B1822_;
  assign new_A7892_ = new_B1855_;
  assign new_A7893_ = new_A7899_ & new_A7898_;
  assign new_A7894_ = new_A7901_ | new_A7900_;
  assign new_A7895_ = new_A7903_ | new_A7902_;
  assign new_A7896_ = new_A7898_ & new_A7904_;
  assign new_A7897_ = new_A7898_ & new_A7905_;
  assign new_A7898_ = new_A7888_ ^ new_A7889_;
  assign new_A7899_ = new_A7900_ ^ new_A7890_;
  assign new_A7900_ = new_A7908_ & new_A7907_;
  assign new_A7901_ = new_A7906_ & new_A7890_;
  assign new_A7902_ = new_A7911_ & new_A7910_;
  assign new_A7903_ = new_A7909_ & new_A7890_;
  assign new_A7904_ = new_A7912_ | new_A7889_;
  assign new_A7905_ = ~new_A7890_ ^ new_A7902_;
  assign new_A7906_ = ~new_A7915_ | ~new_A7916_;
  assign new_A7907_ = new_A7891_ ^ new_A7898_;
  assign new_A7908_ = new_A7917_ & new_A7910_;
  assign new_A7909_ = ~new_A7919_ | ~new_A7918_;
  assign new_A7910_ = new_A7891_ | new_A7892_;
  assign new_A7911_ = new_A7891_ | new_A7898_;
  assign new_A7912_ = new_A7890_ & new_A7902_;
  assign new_A7913_ = ~new_A7889_ | ~new_A7890_;
  assign new_A7914_ = new_A7898_ & new_A7913_;
  assign new_A7915_ = ~new_A7914_ & ~new_A7898_;
  assign new_A7916_ = new_A7898_ | new_A7913_;
  assign new_A7917_ = ~new_A7891_ | ~new_A7892_;
  assign new_A7918_ = new_A7898_ | new_A7913_;
  assign new_A7919_ = ~new_A7898_ & ~new_A7920_;
  assign new_A7920_ = new_A7898_ & new_A7913_;
  assign new_A7921_ = new_B1888_;
  assign new_A7922_ = new_B1921_;
  assign new_A7923_ = new_B1954_;
  assign new_A7924_ = new_B1987_;
  assign new_A7925_ = new_B2020_;
  assign new_A7926_ = new_A7932_ & new_A7931_;
  assign new_A7927_ = new_A7934_ | new_A7933_;
  assign new_A7928_ = new_A7936_ | new_A7935_;
  assign new_A7929_ = new_A7931_ & new_A7937_;
  assign new_A7930_ = new_A7931_ & new_A7938_;
  assign new_A7931_ = new_A7921_ ^ new_A7922_;
  assign new_A7932_ = new_A7933_ ^ new_A7923_;
  assign new_A7933_ = new_A7941_ & new_A7940_;
  assign new_A7934_ = new_A7939_ & new_A7923_;
  assign new_A7935_ = new_A7944_ & new_A7943_;
  assign new_A7936_ = new_A7942_ & new_A7923_;
  assign new_A7937_ = new_A7945_ | new_A7922_;
  assign new_A7938_ = ~new_A7923_ ^ new_A7935_;
  assign new_A7939_ = ~new_A7948_ | ~new_A7949_;
  assign new_A7940_ = new_A7924_ ^ new_A7931_;
  assign new_A7941_ = new_A7950_ & new_A7943_;
  assign new_A7942_ = ~new_A7952_ | ~new_A7951_;
  assign new_A7943_ = new_A7924_ | new_A7925_;
  assign new_A7944_ = new_A7924_ | new_A7931_;
  assign new_A7945_ = new_A7923_ & new_A7935_;
  assign new_A7946_ = ~new_A7922_ | ~new_A7923_;
  assign new_A7947_ = new_A7931_ & new_A7946_;
  assign new_A7948_ = ~new_A7947_ & ~new_A7931_;
  assign new_A7949_ = new_A7931_ | new_A7946_;
  assign new_A7950_ = ~new_A7924_ | ~new_A7925_;
  assign new_A7951_ = new_A7931_ | new_A7946_;
  assign new_A7952_ = ~new_A7931_ & ~new_A7953_;
  assign new_A7953_ = new_A7931_ & new_A7946_;
  assign new_A7954_ = new_B2053_;
  assign new_A7955_ = new_B2086_;
  assign new_A7956_ = new_B2119_;
  assign new_A7957_ = new_B2152_;
  assign new_A7958_ = new_B2185_;
  assign new_A7959_ = new_A7965_ & new_A7964_;
  assign new_A7960_ = new_A7967_ | new_A7966_;
  assign new_A7961_ = new_A7969_ | new_A7968_;
  assign new_A7962_ = new_A7964_ & new_A7970_;
  assign new_A7963_ = new_A7964_ & new_A7971_;
  assign new_A7964_ = new_A7954_ ^ new_A7955_;
  assign new_A7965_ = new_A7966_ ^ new_A7956_;
  assign new_A7966_ = new_A7974_ & new_A7973_;
  assign new_A7967_ = new_A7972_ & new_A7956_;
  assign new_A7968_ = new_A7977_ & new_A7976_;
  assign new_A7969_ = new_A7975_ & new_A7956_;
  assign new_A7970_ = new_A7978_ | new_A7955_;
  assign new_A7971_ = ~new_A7956_ ^ new_A7968_;
  assign new_A7972_ = ~new_A7981_ | ~new_A7982_;
  assign new_A7973_ = new_A7957_ ^ new_A7964_;
  assign new_A7974_ = new_A7983_ & new_A7976_;
  assign new_A7975_ = ~new_A7985_ | ~new_A7984_;
  assign new_A7976_ = new_A7957_ | new_A7958_;
  assign new_A7977_ = new_A7957_ | new_A7964_;
  assign new_A7978_ = new_A7956_ & new_A7968_;
  assign new_A7979_ = ~new_A7955_ | ~new_A7956_;
  assign new_A7980_ = new_A7964_ & new_A7979_;
  assign new_A7981_ = ~new_A7980_ & ~new_A7964_;
  assign new_A7982_ = new_A7964_ | new_A7979_;
  assign new_A7983_ = ~new_A7957_ | ~new_A7958_;
  assign new_A7984_ = new_A7964_ | new_A7979_;
  assign new_A7985_ = ~new_A7964_ & ~new_A7986_;
  assign new_A7986_ = new_A7964_ & new_A7979_;
  assign new_A7987_ = new_B2218_;
  assign new_A7988_ = new_B2251_;
  assign new_A7989_ = new_B2284_;
  assign new_A7990_ = new_B2317_;
  assign new_A7991_ = new_B2350_;
  assign new_A7992_ = new_A7998_ & new_A7997_;
  assign new_A7993_ = new_A8000_ | new_A7999_;
  assign new_A7994_ = new_A8002_ | new_A8001_;
  assign new_A7995_ = new_A7997_ & new_A8003_;
  assign new_A7996_ = new_A7997_ & new_A8004_;
  assign new_A7997_ = new_A7987_ ^ new_A7988_;
  assign new_A7998_ = new_A7999_ ^ new_A7989_;
  assign new_A7999_ = new_A8007_ & new_A8006_;
  assign new_A8000_ = new_A8005_ & new_A7989_;
  assign new_A8001_ = new_A8010_ & new_A8009_;
  assign new_A8002_ = new_A8008_ & new_A7989_;
  assign new_A8003_ = new_A8011_ | new_A7988_;
  assign new_A8004_ = ~new_A7989_ ^ new_A8001_;
  assign new_A8005_ = ~new_A8014_ | ~new_A8015_;
  assign new_A8006_ = new_A7990_ ^ new_A7997_;
  assign new_A8007_ = new_A8016_ & new_A8009_;
  assign new_A8008_ = ~new_A8018_ | ~new_A8017_;
  assign new_A8009_ = new_A7990_ | new_A7991_;
  assign new_A8010_ = new_A7990_ | new_A7997_;
  assign new_A8011_ = new_A7989_ & new_A8001_;
  assign new_A8012_ = ~new_A7988_ | ~new_A7989_;
  assign new_A8013_ = new_A7997_ & new_A8012_;
  assign new_A8014_ = ~new_A8013_ & ~new_A7997_;
  assign new_A8015_ = new_A7997_ | new_A8012_;
  assign new_A8016_ = ~new_A7990_ | ~new_A7991_;
  assign new_A8017_ = new_A7997_ | new_A8012_;
  assign new_A8018_ = ~new_A7997_ & ~new_A8019_;
  assign new_A8019_ = new_A7997_ & new_A8012_;
  assign new_A8020_ = new_B2383_;
  assign new_A8021_ = new_B2416_;
  assign new_A8022_ = new_B2449_;
  assign new_A8023_ = new_B2482_;
  assign new_A8024_ = new_B2515_;
  assign new_A8025_ = new_A8031_ & new_A8030_;
  assign new_A8026_ = new_A8033_ | new_A8032_;
  assign new_A8027_ = new_A8035_ | new_A8034_;
  assign new_A8028_ = new_A8030_ & new_A8036_;
  assign new_A8029_ = new_A8030_ & new_A8037_;
  assign new_A8030_ = new_A8020_ ^ new_A8021_;
  assign new_A8031_ = new_A8032_ ^ new_A8022_;
  assign new_A8032_ = new_A8040_ & new_A8039_;
  assign new_A8033_ = new_A8038_ & new_A8022_;
  assign new_A8034_ = new_A8043_ & new_A8042_;
  assign new_A8035_ = new_A8041_ & new_A8022_;
  assign new_A8036_ = new_A8044_ | new_A8021_;
  assign new_A8037_ = ~new_A8022_ ^ new_A8034_;
  assign new_A8038_ = ~new_A8047_ | ~new_A8048_;
  assign new_A8039_ = new_A8023_ ^ new_A8030_;
  assign new_A8040_ = new_A8049_ & new_A8042_;
  assign new_A8041_ = ~new_A8051_ | ~new_A8050_;
  assign new_A8042_ = new_A8023_ | new_A8024_;
  assign new_A8043_ = new_A8023_ | new_A8030_;
  assign new_A8044_ = new_A8022_ & new_A8034_;
  assign new_A8045_ = ~new_A8021_ | ~new_A8022_;
  assign new_A8046_ = new_A8030_ & new_A8045_;
  assign new_A8047_ = ~new_A8046_ & ~new_A8030_;
  assign new_A8048_ = new_A8030_ | new_A8045_;
  assign new_A8049_ = ~new_A8023_ | ~new_A8024_;
  assign new_A8050_ = new_A8030_ | new_A8045_;
  assign new_A8051_ = ~new_A8030_ & ~new_A8052_;
  assign new_A8052_ = new_A8030_ & new_A8045_;
  assign new_A8053_ = new_B2548_;
  assign new_A8054_ = new_B2581_;
  assign new_A8055_ = new_B2614_;
  assign new_A8056_ = new_B2647_;
  assign new_A8057_ = new_B2680_;
  assign new_A8058_ = new_A8064_ & new_A8063_;
  assign new_A8059_ = new_A8066_ | new_A8065_;
  assign new_A8060_ = new_A8068_ | new_A8067_;
  assign new_A8061_ = new_A8063_ & new_A8069_;
  assign new_A8062_ = new_A8063_ & new_A8070_;
  assign new_A8063_ = new_A8053_ ^ new_A8054_;
  assign new_A8064_ = new_A8065_ ^ new_A8055_;
  assign new_A8065_ = new_A8073_ & new_A8072_;
  assign new_A8066_ = new_A8071_ & new_A8055_;
  assign new_A8067_ = new_A8076_ & new_A8075_;
  assign new_A8068_ = new_A8074_ & new_A8055_;
  assign new_A8069_ = new_A8077_ | new_A8054_;
  assign new_A8070_ = ~new_A8055_ ^ new_A8067_;
  assign new_A8071_ = ~new_A8080_ | ~new_A8081_;
  assign new_A8072_ = new_A8056_ ^ new_A8063_;
  assign new_A8073_ = new_A8082_ & new_A8075_;
  assign new_A8074_ = ~new_A8084_ | ~new_A8083_;
  assign new_A8075_ = new_A8056_ | new_A8057_;
  assign new_A8076_ = new_A8056_ | new_A8063_;
  assign new_A8077_ = new_A8055_ & new_A8067_;
  assign new_A8078_ = ~new_A8054_ | ~new_A8055_;
  assign new_A8079_ = new_A8063_ & new_A8078_;
  assign new_A8080_ = ~new_A8079_ & ~new_A8063_;
  assign new_A8081_ = new_A8063_ | new_A8078_;
  assign new_A8082_ = ~new_A8056_ | ~new_A8057_;
  assign new_A8083_ = new_A8063_ | new_A8078_;
  assign new_A8084_ = ~new_A8063_ & ~new_A8085_;
  assign new_A8085_ = new_A8063_ & new_A8078_;
  assign new_A8086_ = new_B2713_;
  assign new_A8087_ = new_B2746_;
  assign new_A8088_ = new_B2779_;
  assign new_A8089_ = new_B2812_;
  assign new_A8090_ = new_B2845_;
  assign new_A8091_ = new_A8097_ & new_A8096_;
  assign new_A8092_ = new_A8099_ | new_A8098_;
  assign new_A8093_ = new_A8101_ | new_A8100_;
  assign new_A8094_ = new_A8096_ & new_A8102_;
  assign new_A8095_ = new_A8096_ & new_A8103_;
  assign new_A8096_ = new_A8086_ ^ new_A8087_;
  assign new_A8097_ = new_A8098_ ^ new_A8088_;
  assign new_A8098_ = new_A8106_ & new_A8105_;
  assign new_A8099_ = new_A8104_ & new_A8088_;
  assign new_A8100_ = new_A8109_ & new_A8108_;
  assign new_A8101_ = new_A8107_ & new_A8088_;
  assign new_A8102_ = new_A8110_ | new_A8087_;
  assign new_A8103_ = ~new_A8088_ ^ new_A8100_;
  assign new_A8104_ = ~new_A8113_ | ~new_A8114_;
  assign new_A8105_ = new_A8089_ ^ new_A8096_;
  assign new_A8106_ = new_A8115_ & new_A8108_;
  assign new_A8107_ = ~new_A8117_ | ~new_A8116_;
  assign new_A8108_ = new_A8089_ | new_A8090_;
  assign new_A8109_ = new_A8089_ | new_A8096_;
  assign new_A8110_ = new_A8088_ & new_A8100_;
  assign new_A8111_ = ~new_A8087_ | ~new_A8088_;
  assign new_A8112_ = new_A8096_ & new_A8111_;
  assign new_A8113_ = ~new_A8112_ & ~new_A8096_;
  assign new_A8114_ = new_A8096_ | new_A8111_;
  assign new_A8115_ = ~new_A8089_ | ~new_A8090_;
  assign new_A8116_ = new_A8096_ | new_A8111_;
  assign new_A8117_ = ~new_A8096_ & ~new_A8118_;
  assign new_A8118_ = new_A8096_ & new_A8111_;
  assign new_A8119_ = new_B2878_;
  assign new_A8120_ = new_B2911_;
  assign new_A8121_ = new_B2944_;
  assign new_A8122_ = new_B2977_;
  assign new_A8123_ = new_B3010_;
  assign new_A8124_ = new_A8130_ & new_A8129_;
  assign new_A8125_ = new_A8132_ | new_A8131_;
  assign new_A8126_ = new_A8134_ | new_A8133_;
  assign new_A8127_ = new_A8129_ & new_A8135_;
  assign new_A8128_ = new_A8129_ & new_A8136_;
  assign new_A8129_ = new_A8119_ ^ new_A8120_;
  assign new_A8130_ = new_A8131_ ^ new_A8121_;
  assign new_A8131_ = new_A8139_ & new_A8138_;
  assign new_A8132_ = new_A8137_ & new_A8121_;
  assign new_A8133_ = new_A8142_ & new_A8141_;
  assign new_A8134_ = new_A8140_ & new_A8121_;
  assign new_A8135_ = new_A8143_ | new_A8120_;
  assign new_A8136_ = ~new_A8121_ ^ new_A8133_;
  assign new_A8137_ = ~new_A8146_ | ~new_A8147_;
  assign new_A8138_ = new_A8122_ ^ new_A8129_;
  assign new_A8139_ = new_A8148_ & new_A8141_;
  assign new_A8140_ = ~new_A8150_ | ~new_A8149_;
  assign new_A8141_ = new_A8122_ | new_A8123_;
  assign new_A8142_ = new_A8122_ | new_A8129_;
  assign new_A8143_ = new_A8121_ & new_A8133_;
  assign new_A8144_ = ~new_A8120_ | ~new_A8121_;
  assign new_A8145_ = new_A8129_ & new_A8144_;
  assign new_A8146_ = ~new_A8145_ & ~new_A8129_;
  assign new_A8147_ = new_A8129_ | new_A8144_;
  assign new_A8148_ = ~new_A8122_ | ~new_A8123_;
  assign new_A8149_ = new_A8129_ | new_A8144_;
  assign new_A8150_ = ~new_A8129_ & ~new_A8151_;
  assign new_A8151_ = new_A8129_ & new_A8144_;
  assign new_A8152_ = new_B3043_;
  assign new_A8153_ = new_B3076_;
  assign new_A8154_ = new_B3109_;
  assign new_A8155_ = new_B3142_;
  assign new_A8156_ = new_B3175_;
  assign new_A8157_ = new_A8163_ & new_A8162_;
  assign new_A8158_ = new_A8165_ | new_A8164_;
  assign new_A8159_ = new_A8167_ | new_A8166_;
  assign new_A8160_ = new_A8162_ & new_A8168_;
  assign new_A8161_ = new_A8162_ & new_A8169_;
  assign new_A8162_ = new_A8152_ ^ new_A8153_;
  assign new_A8163_ = new_A8164_ ^ new_A8154_;
  assign new_A8164_ = new_A8172_ & new_A8171_;
  assign new_A8165_ = new_A8170_ & new_A8154_;
  assign new_A8166_ = new_A8175_ & new_A8174_;
  assign new_A8167_ = new_A8173_ & new_A8154_;
  assign new_A8168_ = new_A8176_ | new_A8153_;
  assign new_A8169_ = ~new_A8154_ ^ new_A8166_;
  assign new_A8170_ = ~new_A8179_ | ~new_A8180_;
  assign new_A8171_ = new_A8155_ ^ new_A8162_;
  assign new_A8172_ = new_A8181_ & new_A8174_;
  assign new_A8173_ = ~new_A8183_ | ~new_A8182_;
  assign new_A8174_ = new_A8155_ | new_A8156_;
  assign new_A8175_ = new_A8155_ | new_A8162_;
  assign new_A8176_ = new_A8154_ & new_A8166_;
  assign new_A8177_ = ~new_A8153_ | ~new_A8154_;
  assign new_A8178_ = new_A8162_ & new_A8177_;
  assign new_A8179_ = ~new_A8178_ & ~new_A8162_;
  assign new_A8180_ = new_A8162_ | new_A8177_;
  assign new_A8181_ = ~new_A8155_ | ~new_A8156_;
  assign new_A8182_ = new_A8162_ | new_A8177_;
  assign new_A8183_ = ~new_A8162_ & ~new_A8184_;
  assign new_A8184_ = new_A8162_ & new_A8177_;
  assign new_A8185_ = new_B3208_;
  assign new_A8186_ = new_B3241_;
  assign new_A8187_ = new_B3274_;
  assign new_A8188_ = new_B3307_;
  assign new_A8189_ = new_B3340_;
  assign new_A8190_ = new_A8196_ & new_A8195_;
  assign new_A8191_ = new_A8198_ | new_A8197_;
  assign new_A8192_ = new_A8200_ | new_A8199_;
  assign new_A8193_ = new_A8195_ & new_A8201_;
  assign new_A8194_ = new_A8195_ & new_A8202_;
  assign new_A8195_ = new_A8185_ ^ new_A8186_;
  assign new_A8196_ = new_A8197_ ^ new_A8187_;
  assign new_A8197_ = new_A8205_ & new_A8204_;
  assign new_A8198_ = new_A8203_ & new_A8187_;
  assign new_A8199_ = new_A8208_ & new_A8207_;
  assign new_A8200_ = new_A8206_ & new_A8187_;
  assign new_A8201_ = new_A8209_ | new_A8186_;
  assign new_A8202_ = ~new_A8187_ ^ new_A8199_;
  assign new_A8203_ = ~new_A8212_ | ~new_A8213_;
  assign new_A8204_ = new_A8188_ ^ new_A8195_;
  assign new_A8205_ = new_A8214_ & new_A8207_;
  assign new_A8206_ = ~new_A8216_ | ~new_A8215_;
  assign new_A8207_ = new_A8188_ | new_A8189_;
  assign new_A8208_ = new_A8188_ | new_A8195_;
  assign new_A8209_ = new_A8187_ & new_A8199_;
  assign new_A8210_ = ~new_A8186_ | ~new_A8187_;
  assign new_A8211_ = new_A8195_ & new_A8210_;
  assign new_A8212_ = ~new_A8211_ & ~new_A8195_;
  assign new_A8213_ = new_A8195_ | new_A8210_;
  assign new_A8214_ = ~new_A8188_ | ~new_A8189_;
  assign new_A8215_ = new_A8195_ | new_A8210_;
  assign new_A8216_ = ~new_A8195_ & ~new_A8217_;
  assign new_A8217_ = new_A8195_ & new_A8210_;
  assign new_A8218_ = new_B3373_;
  assign new_A8219_ = new_B3406_;
  assign new_A8220_ = new_B3439_;
  assign new_A8221_ = new_B3472_;
  assign new_A8222_ = new_B3505_;
  assign new_A8223_ = new_A8229_ & new_A8228_;
  assign new_A8224_ = new_A8231_ | new_A8230_;
  assign new_A8225_ = new_A8233_ | new_A8232_;
  assign new_A8226_ = new_A8228_ & new_A8234_;
  assign new_A8227_ = new_A8228_ & new_A8235_;
  assign new_A8228_ = new_A8218_ ^ new_A8219_;
  assign new_A8229_ = new_A8230_ ^ new_A8220_;
  assign new_A8230_ = new_A8238_ & new_A8237_;
  assign new_A8231_ = new_A8236_ & new_A8220_;
  assign new_A8232_ = new_A8241_ & new_A8240_;
  assign new_A8233_ = new_A8239_ & new_A8220_;
  assign new_A8234_ = new_A8242_ | new_A8219_;
  assign new_A8235_ = ~new_A8220_ ^ new_A8232_;
  assign new_A8236_ = ~new_A8245_ | ~new_A8246_;
  assign new_A8237_ = new_A8221_ ^ new_A8228_;
  assign new_A8238_ = new_A8247_ & new_A8240_;
  assign new_A8239_ = ~new_A8249_ | ~new_A8248_;
  assign new_A8240_ = new_A8221_ | new_A8222_;
  assign new_A8241_ = new_A8221_ | new_A8228_;
  assign new_A8242_ = new_A8220_ & new_A8232_;
  assign new_A8243_ = ~new_A8219_ | ~new_A8220_;
  assign new_A8244_ = new_A8228_ & new_A8243_;
  assign new_A8245_ = ~new_A8244_ & ~new_A8228_;
  assign new_A8246_ = new_A8228_ | new_A8243_;
  assign new_A8247_ = ~new_A8221_ | ~new_A8222_;
  assign new_A8248_ = new_A8228_ | new_A8243_;
  assign new_A8249_ = ~new_A8228_ & ~new_A8250_;
  assign new_A8250_ = new_A8228_ & new_A8243_;
  assign new_A8251_ = new_B3538_;
  assign new_A8252_ = new_B3571_;
  assign new_A8253_ = new_B3604_;
  assign new_A8254_ = new_B3637_;
  assign new_A8255_ = new_B3670_;
  assign new_A8256_ = new_A8262_ & new_A8261_;
  assign new_A8257_ = new_A8264_ | new_A8263_;
  assign new_A8258_ = new_A8266_ | new_A8265_;
  assign new_A8259_ = new_A8261_ & new_A8267_;
  assign new_A8260_ = new_A8261_ & new_A8268_;
  assign new_A8261_ = new_A8251_ ^ new_A8252_;
  assign new_A8262_ = new_A8263_ ^ new_A8253_;
  assign new_A8263_ = new_A8271_ & new_A8270_;
  assign new_A8264_ = new_A8269_ & new_A8253_;
  assign new_A8265_ = new_A8274_ & new_A8273_;
  assign new_A8266_ = new_A8272_ & new_A8253_;
  assign new_A8267_ = new_A8275_ | new_A8252_;
  assign new_A8268_ = ~new_A8253_ ^ new_A8265_;
  assign new_A8269_ = ~new_A8278_ | ~new_A8279_;
  assign new_A8270_ = new_A8254_ ^ new_A8261_;
  assign new_A8271_ = new_A8280_ & new_A8273_;
  assign new_A8272_ = ~new_A8282_ | ~new_A8281_;
  assign new_A8273_ = new_A8254_ | new_A8255_;
  assign new_A8274_ = new_A8254_ | new_A8261_;
  assign new_A8275_ = new_A8253_ & new_A8265_;
  assign new_A8276_ = ~new_A8252_ | ~new_A8253_;
  assign new_A8277_ = new_A8261_ & new_A8276_;
  assign new_A8278_ = ~new_A8277_ & ~new_A8261_;
  assign new_A8279_ = new_A8261_ | new_A8276_;
  assign new_A8280_ = ~new_A8254_ | ~new_A8255_;
  assign new_A8281_ = new_A8261_ | new_A8276_;
  assign new_A8282_ = ~new_A8261_ & ~new_A8283_;
  assign new_A8283_ = new_A8261_ & new_A8276_;
  assign new_A8284_ = new_B3703_;
  assign new_A8285_ = new_B3736_;
  assign new_A8286_ = new_B3769_;
  assign new_A8287_ = new_B3802_;
  assign new_A8288_ = new_B3835_;
  assign new_A8289_ = new_A8295_ & new_A8294_;
  assign new_A8290_ = new_A8297_ | new_A8296_;
  assign new_A8291_ = new_A8299_ | new_A8298_;
  assign new_A8292_ = new_A8294_ & new_A8300_;
  assign new_A8293_ = new_A8294_ & new_A8301_;
  assign new_A8294_ = new_A8284_ ^ new_A8285_;
  assign new_A8295_ = new_A8296_ ^ new_A8286_;
  assign new_A8296_ = new_A8304_ & new_A8303_;
  assign new_A8297_ = new_A8302_ & new_A8286_;
  assign new_A8298_ = new_A8307_ & new_A8306_;
  assign new_A8299_ = new_A8305_ & new_A8286_;
  assign new_A8300_ = new_A8308_ | new_A8285_;
  assign new_A8301_ = ~new_A8286_ ^ new_A8298_;
  assign new_A8302_ = ~new_A8311_ | ~new_A8312_;
  assign new_A8303_ = new_A8287_ ^ new_A8294_;
  assign new_A8304_ = new_A8313_ & new_A8306_;
  assign new_A8305_ = ~new_A8315_ | ~new_A8314_;
  assign new_A8306_ = new_A8287_ | new_A8288_;
  assign new_A8307_ = new_A8287_ | new_A8294_;
  assign new_A8308_ = new_A8286_ & new_A8298_;
  assign new_A8309_ = ~new_A8285_ | ~new_A8286_;
  assign new_A8310_ = new_A8294_ & new_A8309_;
  assign new_A8311_ = ~new_A8310_ & ~new_A8294_;
  assign new_A8312_ = new_A8294_ | new_A8309_;
  assign new_A8313_ = ~new_A8287_ | ~new_A8288_;
  assign new_A8314_ = new_A8294_ | new_A8309_;
  assign new_A8315_ = ~new_A8294_ & ~new_A8316_;
  assign new_A8316_ = new_A8294_ & new_A8309_;
  assign new_A8317_ = new_B3868_;
  assign new_A8318_ = new_B3901_;
  assign new_A8319_ = new_B3934_;
  assign new_A8320_ = new_B3967_;
  assign new_A8321_ = new_B4000_;
  assign new_A8322_ = new_A8328_ & new_A8327_;
  assign new_A8323_ = new_A8330_ | new_A8329_;
  assign new_A8324_ = new_A8332_ | new_A8331_;
  assign new_A8325_ = new_A8327_ & new_A8333_;
  assign new_A8326_ = new_A8327_ & new_A8334_;
  assign new_A8327_ = new_A8317_ ^ new_A8318_;
  assign new_A8328_ = new_A8329_ ^ new_A8319_;
  assign new_A8329_ = new_A8337_ & new_A8336_;
  assign new_A8330_ = new_A8335_ & new_A8319_;
  assign new_A8331_ = new_A8340_ & new_A8339_;
  assign new_A8332_ = new_A8338_ & new_A8319_;
  assign new_A8333_ = new_A8341_ | new_A8318_;
  assign new_A8334_ = ~new_A8319_ ^ new_A8331_;
  assign new_A8335_ = ~new_A8344_ | ~new_A8345_;
  assign new_A8336_ = new_A8320_ ^ new_A8327_;
  assign new_A8337_ = new_A8346_ & new_A8339_;
  assign new_A8338_ = ~new_A8348_ | ~new_A8347_;
  assign new_A8339_ = new_A8320_ | new_A8321_;
  assign new_A8340_ = new_A8320_ | new_A8327_;
  assign new_A8341_ = new_A8319_ & new_A8331_;
  assign new_A8342_ = ~new_A8318_ | ~new_A8319_;
  assign new_A8343_ = new_A8327_ & new_A8342_;
  assign new_A8344_ = ~new_A8343_ & ~new_A8327_;
  assign new_A8345_ = new_A8327_ | new_A8342_;
  assign new_A8346_ = ~new_A8320_ | ~new_A8321_;
  assign new_A8347_ = new_A8327_ | new_A8342_;
  assign new_A8348_ = ~new_A8327_ & ~new_A8349_;
  assign new_A8349_ = new_A8327_ & new_A8342_;
  assign new_A8350_ = new_B4033_;
  assign new_A8351_ = new_B4066_;
  assign new_A8352_ = new_B4099_;
  assign new_A8353_ = new_B4132_;
  assign new_A8354_ = new_B4165_;
  assign new_A8355_ = new_A8361_ & new_A8360_;
  assign new_A8356_ = new_A8363_ | new_A8362_;
  assign new_A8357_ = new_A8365_ | new_A8364_;
  assign new_A8358_ = new_A8360_ & new_A8366_;
  assign new_A8359_ = new_A8360_ & new_A8367_;
  assign new_A8360_ = new_A8350_ ^ new_A8351_;
  assign new_A8361_ = new_A8362_ ^ new_A8352_;
  assign new_A8362_ = new_A8370_ & new_A8369_;
  assign new_A8363_ = new_A8368_ & new_A8352_;
  assign new_A8364_ = new_A8373_ & new_A8372_;
  assign new_A8365_ = new_A8371_ & new_A8352_;
  assign new_A8366_ = new_A8374_ | new_A8351_;
  assign new_A8367_ = ~new_A8352_ ^ new_A8364_;
  assign new_A8368_ = ~new_A8377_ | ~new_A8378_;
  assign new_A8369_ = new_A8353_ ^ new_A8360_;
  assign new_A8370_ = new_A8379_ & new_A8372_;
  assign new_A8371_ = ~new_A8381_ | ~new_A8380_;
  assign new_A8372_ = new_A8353_ | new_A8354_;
  assign new_A8373_ = new_A8353_ | new_A8360_;
  assign new_A8374_ = new_A8352_ & new_A8364_;
  assign new_A8375_ = ~new_A8351_ | ~new_A8352_;
  assign new_A8376_ = new_A8360_ & new_A8375_;
  assign new_A8377_ = ~new_A8376_ & ~new_A8360_;
  assign new_A8378_ = new_A8360_ | new_A8375_;
  assign new_A8379_ = ~new_A8353_ | ~new_A8354_;
  assign new_A8380_ = new_A8360_ | new_A8375_;
  assign new_A8381_ = ~new_A8360_ & ~new_A8382_;
  assign new_A8382_ = new_A8360_ & new_A8375_;
  assign new_A8383_ = new_B4198_;
  assign new_A8384_ = new_B4231_;
  assign new_A8385_ = new_B4264_;
  assign new_A8386_ = new_B4297_;
  assign new_A8387_ = new_B4330_;
  assign new_A8388_ = new_A8394_ & new_A8393_;
  assign new_A8389_ = new_A8396_ | new_A8395_;
  assign new_A8390_ = new_A8398_ | new_A8397_;
  assign new_A8391_ = new_A8393_ & new_A8399_;
  assign new_A8392_ = new_A8393_ & new_A8400_;
  assign new_A8393_ = new_A8383_ ^ new_A8384_;
  assign new_A8394_ = new_A8395_ ^ new_A8385_;
  assign new_A8395_ = new_A8403_ & new_A8402_;
  assign new_A8396_ = new_A8401_ & new_A8385_;
  assign new_A8397_ = new_A8406_ & new_A8405_;
  assign new_A8398_ = new_A8404_ & new_A8385_;
  assign new_A8399_ = new_A8407_ | new_A8384_;
  assign new_A8400_ = ~new_A8385_ ^ new_A8397_;
  assign new_A8401_ = ~new_A8410_ | ~new_A8411_;
  assign new_A8402_ = new_A8386_ ^ new_A8393_;
  assign new_A8403_ = new_A8412_ & new_A8405_;
  assign new_A8404_ = ~new_A8414_ | ~new_A8413_;
  assign new_A8405_ = new_A8386_ | new_A8387_;
  assign new_A8406_ = new_A8386_ | new_A8393_;
  assign new_A8407_ = new_A8385_ & new_A8397_;
  assign new_A8408_ = ~new_A8384_ | ~new_A8385_;
  assign new_A8409_ = new_A8393_ & new_A8408_;
  assign new_A8410_ = ~new_A8409_ & ~new_A8393_;
  assign new_A8411_ = new_A8393_ | new_A8408_;
  assign new_A8412_ = ~new_A8386_ | ~new_A8387_;
  assign new_A8413_ = new_A8393_ | new_A8408_;
  assign new_A8414_ = ~new_A8393_ & ~new_A8415_;
  assign new_A8415_ = new_A8393_ & new_A8408_;
  assign new_A8416_ = new_B4363_;
  assign new_A8417_ = new_B4396_;
  assign new_A8418_ = new_B4429_;
  assign new_A8419_ = new_B4462_;
  assign new_A8420_ = new_B4495_;
  assign new_A8421_ = new_A8427_ & new_A8426_;
  assign new_A8422_ = new_A8429_ | new_A8428_;
  assign new_A8423_ = new_A8431_ | new_A8430_;
  assign new_A8424_ = new_A8426_ & new_A8432_;
  assign new_A8425_ = new_A8426_ & new_A8433_;
  assign new_A8426_ = new_A8416_ ^ new_A8417_;
  assign new_A8427_ = new_A8428_ ^ new_A8418_;
  assign new_A8428_ = new_A8436_ & new_A8435_;
  assign new_A8429_ = new_A8434_ & new_A8418_;
  assign new_A8430_ = new_A8439_ & new_A8438_;
  assign new_A8431_ = new_A8437_ & new_A8418_;
  assign new_A8432_ = new_A8440_ | new_A8417_;
  assign new_A8433_ = ~new_A8418_ ^ new_A8430_;
  assign new_A8434_ = ~new_A8443_ | ~new_A8444_;
  assign new_A8435_ = new_A8419_ ^ new_A8426_;
  assign new_A8436_ = new_A8445_ & new_A8438_;
  assign new_A8437_ = ~new_A8447_ | ~new_A8446_;
  assign new_A8438_ = new_A8419_ | new_A8420_;
  assign new_A8439_ = new_A8419_ | new_A8426_;
  assign new_A8440_ = new_A8418_ & new_A8430_;
  assign new_A8441_ = ~new_A8417_ | ~new_A8418_;
  assign new_A8442_ = new_A8426_ & new_A8441_;
  assign new_A8443_ = ~new_A8442_ & ~new_A8426_;
  assign new_A8444_ = new_A8426_ | new_A8441_;
  assign new_A8445_ = ~new_A8419_ | ~new_A8420_;
  assign new_A8446_ = new_A8426_ | new_A8441_;
  assign new_A8447_ = ~new_A8426_ & ~new_A8448_;
  assign new_A8448_ = new_A8426_ & new_A8441_;
  assign new_A8449_ = new_B4528_;
  assign new_A8450_ = new_B4561_;
  assign new_A8451_ = new_B4594_;
  assign new_A8452_ = new_B4627_;
  assign new_A8453_ = new_B4660_;
  assign new_A8454_ = new_A8460_ & new_A8459_;
  assign new_A8455_ = new_A8462_ | new_A8461_;
  assign new_A8456_ = new_A8464_ | new_A8463_;
  assign new_A8457_ = new_A8459_ & new_A8465_;
  assign new_A8458_ = new_A8459_ & new_A8466_;
  assign new_A8459_ = new_A8449_ ^ new_A8450_;
  assign new_A8460_ = new_A8461_ ^ new_A8451_;
  assign new_A8461_ = new_A8469_ & new_A8468_;
  assign new_A8462_ = new_A8467_ & new_A8451_;
  assign new_A8463_ = new_A8472_ & new_A8471_;
  assign new_A8464_ = new_A8470_ & new_A8451_;
  assign new_A8465_ = new_A8473_ | new_A8450_;
  assign new_A8466_ = ~new_A8451_ ^ new_A8463_;
  assign new_A8467_ = ~new_A8476_ | ~new_A8477_;
  assign new_A8468_ = new_A8452_ ^ new_A8459_;
  assign new_A8469_ = new_A8478_ & new_A8471_;
  assign new_A8470_ = ~new_A8480_ | ~new_A8479_;
  assign new_A8471_ = new_A8452_ | new_A8453_;
  assign new_A8472_ = new_A8452_ | new_A8459_;
  assign new_A8473_ = new_A8451_ & new_A8463_;
  assign new_A8474_ = ~new_A8450_ | ~new_A8451_;
  assign new_A8475_ = new_A8459_ & new_A8474_;
  assign new_A8476_ = ~new_A8475_ & ~new_A8459_;
  assign new_A8477_ = new_A8459_ | new_A8474_;
  assign new_A8478_ = ~new_A8452_ | ~new_A8453_;
  assign new_A8479_ = new_A8459_ | new_A8474_;
  assign new_A8480_ = ~new_A8459_ & ~new_A8481_;
  assign new_A8481_ = new_A8459_ & new_A8474_;
  assign new_A8482_ = new_B4693_;
  assign new_A8483_ = new_B4726_;
  assign new_A8484_ = new_B4759_;
  assign new_A8485_ = new_B4792_;
  assign new_A8486_ = new_B4825_;
  assign new_A8487_ = new_A8493_ & new_A8492_;
  assign new_A8488_ = new_A8495_ | new_A8494_;
  assign new_A8489_ = new_A8497_ | new_A8496_;
  assign new_A8490_ = new_A8492_ & new_A8498_;
  assign new_A8491_ = new_A8492_ & new_A8499_;
  assign new_A8492_ = new_A8482_ ^ new_A8483_;
  assign new_A8493_ = new_A8494_ ^ new_A8484_;
  assign new_A8494_ = new_A8502_ & new_A8501_;
  assign new_A8495_ = new_A8500_ & new_A8484_;
  assign new_A8496_ = new_A8505_ & new_A8504_;
  assign new_A8497_ = new_A8503_ & new_A8484_;
  assign new_A8498_ = new_A8506_ | new_A8483_;
  assign new_A8499_ = ~new_A8484_ ^ new_A8496_;
  assign new_A8500_ = ~new_A8509_ | ~new_A8510_;
  assign new_A8501_ = new_A8485_ ^ new_A8492_;
  assign new_A8502_ = new_A8511_ & new_A8504_;
  assign new_A8503_ = ~new_A8513_ | ~new_A8512_;
  assign new_A8504_ = new_A8485_ | new_A8486_;
  assign new_A8505_ = new_A8485_ | new_A8492_;
  assign new_A8506_ = new_A8484_ & new_A8496_;
  assign new_A8507_ = ~new_A8483_ | ~new_A8484_;
  assign new_A8508_ = new_A8492_ & new_A8507_;
  assign new_A8509_ = ~new_A8508_ & ~new_A8492_;
  assign new_A8510_ = new_A8492_ | new_A8507_;
  assign new_A8511_ = ~new_A8485_ | ~new_A8486_;
  assign new_A8512_ = new_A8492_ | new_A8507_;
  assign new_A8513_ = ~new_A8492_ & ~new_A8514_;
  assign new_A8514_ = new_A8492_ & new_A8507_;
  assign new_A8515_ = new_B4858_;
  assign new_A8516_ = new_B4891_;
  assign new_A8517_ = new_B4924_;
  assign new_A8518_ = new_B4957_;
  assign new_A8519_ = new_B4990_;
  assign new_A8520_ = new_A8526_ & new_A8525_;
  assign new_A8521_ = new_A8528_ | new_A8527_;
  assign new_A8522_ = new_A8530_ | new_A8529_;
  assign new_A8523_ = new_A8525_ & new_A8531_;
  assign new_A8524_ = new_A8525_ & new_A8532_;
  assign new_A8525_ = new_A8515_ ^ new_A8516_;
  assign new_A8526_ = new_A8527_ ^ new_A8517_;
  assign new_A8527_ = new_A8535_ & new_A8534_;
  assign new_A8528_ = new_A8533_ & new_A8517_;
  assign new_A8529_ = new_A8538_ & new_A8537_;
  assign new_A8530_ = new_A8536_ & new_A8517_;
  assign new_A8531_ = new_A8539_ | new_A8516_;
  assign new_A8532_ = ~new_A8517_ ^ new_A8529_;
  assign new_A8533_ = ~new_A8542_ | ~new_A8543_;
  assign new_A8534_ = new_A8518_ ^ new_A8525_;
  assign new_A8535_ = new_A8544_ & new_A8537_;
  assign new_A8536_ = ~new_A8546_ | ~new_A8545_;
  assign new_A8537_ = new_A8518_ | new_A8519_;
  assign new_A8538_ = new_A8518_ | new_A8525_;
  assign new_A8539_ = new_A8517_ & new_A8529_;
  assign new_A8540_ = ~new_A8516_ | ~new_A8517_;
  assign new_A8541_ = new_A8525_ & new_A8540_;
  assign new_A8542_ = ~new_A8541_ & ~new_A8525_;
  assign new_A8543_ = new_A8525_ | new_A8540_;
  assign new_A8544_ = ~new_A8518_ | ~new_A8519_;
  assign new_A8545_ = new_A8525_ | new_A8540_;
  assign new_A8546_ = ~new_A8525_ & ~new_A8547_;
  assign new_A8547_ = new_A8525_ & new_A8540_;
  assign new_A8548_ = new_B5023_;
  assign new_A8549_ = new_B5056_;
  assign new_A8550_ = new_B5089_;
  assign new_A8551_ = new_B5122_;
  assign new_A8552_ = new_B5155_;
  assign new_A8553_ = new_A8559_ & new_A8558_;
  assign new_A8554_ = new_A8561_ | new_A8560_;
  assign new_A8555_ = new_A8563_ | new_A8562_;
  assign new_A8556_ = new_A8558_ & new_A8564_;
  assign new_A8557_ = new_A8558_ & new_A8565_;
  assign new_A8558_ = new_A8548_ ^ new_A8549_;
  assign new_A8559_ = new_A8560_ ^ new_A8550_;
  assign new_A8560_ = new_A8568_ & new_A8567_;
  assign new_A8561_ = new_A8566_ & new_A8550_;
  assign new_A8562_ = new_A8571_ & new_A8570_;
  assign new_A8563_ = new_A8569_ & new_A8550_;
  assign new_A8564_ = new_A8572_ | new_A8549_;
  assign new_A8565_ = ~new_A8550_ ^ new_A8562_;
  assign new_A8566_ = ~new_A8575_ | ~new_A8576_;
  assign new_A8567_ = new_A8551_ ^ new_A8558_;
  assign new_A8568_ = new_A8577_ & new_A8570_;
  assign new_A8569_ = ~new_A8579_ | ~new_A8578_;
  assign new_A8570_ = new_A8551_ | new_A8552_;
  assign new_A8571_ = new_A8551_ | new_A8558_;
  assign new_A8572_ = new_A8550_ & new_A8562_;
  assign new_A8573_ = ~new_A8549_ | ~new_A8550_;
  assign new_A8574_ = new_A8558_ & new_A8573_;
  assign new_A8575_ = ~new_A8574_ & ~new_A8558_;
  assign new_A8576_ = new_A8558_ | new_A8573_;
  assign new_A8577_ = ~new_A8551_ | ~new_A8552_;
  assign new_A8578_ = new_A8558_ | new_A8573_;
  assign new_A8579_ = ~new_A8558_ & ~new_A8580_;
  assign new_A8580_ = new_A8558_ & new_A8573_;
  assign new_A8581_ = new_B1064_;
  assign new_A8582_ = new_B1097_;
  assign new_A8583_ = new_B1130_;
  assign new_A8584_ = new_B1163_;
  assign new_A8585_ = new_B1196_;
  assign new_A8586_ = new_A8592_ & new_A8591_;
  assign new_A8587_ = new_A8594_ | new_A8593_;
  assign new_A8588_ = new_A8596_ | new_A8595_;
  assign new_A8589_ = new_A8591_ & new_A8597_;
  assign new_A8590_ = new_A8591_ & new_A8598_;
  assign new_A8591_ = new_A8581_ ^ new_A8582_;
  assign new_A8592_ = new_A8593_ ^ new_A8583_;
  assign new_A8593_ = new_A8601_ & new_A8600_;
  assign new_A8594_ = new_A8599_ & new_A8583_;
  assign new_A8595_ = new_A8604_ & new_A8603_;
  assign new_A8596_ = new_A8602_ & new_A8583_;
  assign new_A8597_ = new_A8605_ | new_A8582_;
  assign new_A8598_ = ~new_A8583_ ^ new_A8595_;
  assign new_A8599_ = ~new_A8608_ | ~new_A8609_;
  assign new_A8600_ = new_A8584_ ^ new_A8591_;
  assign new_A8601_ = new_A8610_ & new_A8603_;
  assign new_A8602_ = ~new_A8612_ | ~new_A8611_;
  assign new_A8603_ = new_A8584_ | new_A8585_;
  assign new_A8604_ = new_A8584_ | new_A8591_;
  assign new_A8605_ = new_A8583_ & new_A8595_;
  assign new_A8606_ = ~new_A8582_ | ~new_A8583_;
  assign new_A8607_ = new_A8591_ & new_A8606_;
  assign new_A8608_ = ~new_A8607_ & ~new_A8591_;
  assign new_A8609_ = new_A8591_ | new_A8606_;
  assign new_A8610_ = ~new_A8584_ | ~new_A8585_;
  assign new_A8611_ = new_A8591_ | new_A8606_;
  assign new_A8612_ = ~new_A8591_ & ~new_A8613_;
  assign new_A8613_ = new_A8591_ & new_A8606_;
  assign new_A8614_ = new_B1229_;
  assign new_A8615_ = new_B1262_;
  assign new_A8616_ = new_B1295_;
  assign new_A8617_ = new_B1328_;
  assign new_A8618_ = new_B1361_;
  assign new_A8619_ = new_A8625_ & new_A8624_;
  assign new_A8620_ = new_A8627_ | new_A8626_;
  assign new_A8621_ = new_A8629_ | new_A8628_;
  assign new_A8622_ = new_A8624_ & new_A8630_;
  assign new_A8623_ = new_A8624_ & new_A8631_;
  assign new_A8624_ = new_A8614_ ^ new_A8615_;
  assign new_A8625_ = new_A8626_ ^ new_A8616_;
  assign new_A8626_ = new_A8634_ & new_A8633_;
  assign new_A8627_ = new_A8632_ & new_A8616_;
  assign new_A8628_ = new_A8637_ & new_A8636_;
  assign new_A8629_ = new_A8635_ & new_A8616_;
  assign new_A8630_ = new_A8638_ | new_A8615_;
  assign new_A8631_ = ~new_A8616_ ^ new_A8628_;
  assign new_A8632_ = ~new_A8641_ | ~new_A8642_;
  assign new_A8633_ = new_A8617_ ^ new_A8624_;
  assign new_A8634_ = new_A8643_ & new_A8636_;
  assign new_A8635_ = ~new_A8645_ | ~new_A8644_;
  assign new_A8636_ = new_A8617_ | new_A8618_;
  assign new_A8637_ = new_A8617_ | new_A8624_;
  assign new_A8638_ = new_A8616_ & new_A8628_;
  assign new_A8639_ = ~new_A8615_ | ~new_A8616_;
  assign new_A8640_ = new_A8624_ & new_A8639_;
  assign new_A8641_ = ~new_A8640_ & ~new_A8624_;
  assign new_A8642_ = new_A8624_ | new_A8639_;
  assign new_A8643_ = ~new_A8617_ | ~new_A8618_;
  assign new_A8644_ = new_A8624_ | new_A8639_;
  assign new_A8645_ = ~new_A8624_ & ~new_A8646_;
  assign new_A8646_ = new_A8624_ & new_A8639_;
  assign new_A8647_ = new_B1394_;
  assign new_A8648_ = new_B1427_;
  assign new_A8649_ = new_B1460_;
  assign new_A8650_ = new_B1493_;
  assign new_A8651_ = new_B1526_;
  assign new_A8652_ = new_A8658_ & new_A8657_;
  assign new_A8653_ = new_A8660_ | new_A8659_;
  assign new_A8654_ = new_A8662_ | new_A8661_;
  assign new_A8655_ = new_A8657_ & new_A8663_;
  assign new_A8656_ = new_A8657_ & new_A8664_;
  assign new_A8657_ = new_A8647_ ^ new_A8648_;
  assign new_A8658_ = new_A8659_ ^ new_A8649_;
  assign new_A8659_ = new_A8667_ & new_A8666_;
  assign new_A8660_ = new_A8665_ & new_A8649_;
  assign new_A8661_ = new_A8670_ & new_A8669_;
  assign new_A8662_ = new_A8668_ & new_A8649_;
  assign new_A8663_ = new_A8671_ | new_A8648_;
  assign new_A8664_ = ~new_A8649_ ^ new_A8661_;
  assign new_A8665_ = ~new_A8674_ | ~new_A8675_;
  assign new_A8666_ = new_A8650_ ^ new_A8657_;
  assign new_A8667_ = new_A8676_ & new_A8669_;
  assign new_A8668_ = ~new_A8678_ | ~new_A8677_;
  assign new_A8669_ = new_A8650_ | new_A8651_;
  assign new_A8670_ = new_A8650_ | new_A8657_;
  assign new_A8671_ = new_A8649_ & new_A8661_;
  assign new_A8672_ = ~new_A8648_ | ~new_A8649_;
  assign new_A8673_ = new_A8657_ & new_A8672_;
  assign new_A8674_ = ~new_A8673_ & ~new_A8657_;
  assign new_A8675_ = new_A8657_ | new_A8672_;
  assign new_A8676_ = ~new_A8650_ | ~new_A8651_;
  assign new_A8677_ = new_A8657_ | new_A8672_;
  assign new_A8678_ = ~new_A8657_ & ~new_A8679_;
  assign new_A8679_ = new_A8657_ & new_A8672_;
  assign new_A8680_ = new_B1559_;
  assign new_A8681_ = new_B1592_;
  assign new_A8682_ = new_B1625_;
  assign new_A8683_ = new_B1658_;
  assign new_A8684_ = new_B1691_;
  assign new_A8685_ = new_A8691_ & new_A8690_;
  assign new_A8686_ = new_A8693_ | new_A8692_;
  assign new_A8687_ = new_A8695_ | new_A8694_;
  assign new_A8688_ = new_A8690_ & new_A8696_;
  assign new_A8689_ = new_A8690_ & new_A8697_;
  assign new_A8690_ = new_A8680_ ^ new_A8681_;
  assign new_A8691_ = new_A8692_ ^ new_A8682_;
  assign new_A8692_ = new_A8700_ & new_A8699_;
  assign new_A8693_ = new_A8698_ & new_A8682_;
  assign new_A8694_ = new_A8703_ & new_A8702_;
  assign new_A8695_ = new_A8701_ & new_A8682_;
  assign new_A8696_ = new_A8704_ | new_A8681_;
  assign new_A8697_ = ~new_A8682_ ^ new_A8694_;
  assign new_A8698_ = ~new_A8707_ | ~new_A8708_;
  assign new_A8699_ = new_A8683_ ^ new_A8690_;
  assign new_A8700_ = new_A8709_ & new_A8702_;
  assign new_A8701_ = ~new_A8711_ | ~new_A8710_;
  assign new_A8702_ = new_A8683_ | new_A8684_;
  assign new_A8703_ = new_A8683_ | new_A8690_;
  assign new_A8704_ = new_A8682_ & new_A8694_;
  assign new_A8705_ = ~new_A8681_ | ~new_A8682_;
  assign new_A8706_ = new_A8690_ & new_A8705_;
  assign new_A8707_ = ~new_A8706_ & ~new_A8690_;
  assign new_A8708_ = new_A8690_ | new_A8705_;
  assign new_A8709_ = ~new_A8683_ | ~new_A8684_;
  assign new_A8710_ = new_A8690_ | new_A8705_;
  assign new_A8711_ = ~new_A8690_ & ~new_A8712_;
  assign new_A8712_ = new_A8690_ & new_A8705_;
  assign new_A8713_ = new_B1724_;
  assign new_A8714_ = new_B1757_;
  assign new_A8715_ = new_B1790_;
  assign new_A8716_ = new_B1823_;
  assign new_A8717_ = new_B1856_;
  assign new_A8718_ = new_A8724_ & new_A8723_;
  assign new_A8719_ = new_A8726_ | new_A8725_;
  assign new_A8720_ = new_A8728_ | new_A8727_;
  assign new_A8721_ = new_A8723_ & new_A8729_;
  assign new_A8722_ = new_A8723_ & new_A8730_;
  assign new_A8723_ = new_A8713_ ^ new_A8714_;
  assign new_A8724_ = new_A8725_ ^ new_A8715_;
  assign new_A8725_ = new_A8733_ & new_A8732_;
  assign new_A8726_ = new_A8731_ & new_A8715_;
  assign new_A8727_ = new_A8736_ & new_A8735_;
  assign new_A8728_ = new_A8734_ & new_A8715_;
  assign new_A8729_ = new_A8737_ | new_A8714_;
  assign new_A8730_ = ~new_A8715_ ^ new_A8727_;
  assign new_A8731_ = ~new_A8740_ | ~new_A8741_;
  assign new_A8732_ = new_A8716_ ^ new_A8723_;
  assign new_A8733_ = new_A8742_ & new_A8735_;
  assign new_A8734_ = ~new_A8744_ | ~new_A8743_;
  assign new_A8735_ = new_A8716_ | new_A8717_;
  assign new_A8736_ = new_A8716_ | new_A8723_;
  assign new_A8737_ = new_A8715_ & new_A8727_;
  assign new_A8738_ = ~new_A8714_ | ~new_A8715_;
  assign new_A8739_ = new_A8723_ & new_A8738_;
  assign new_A8740_ = ~new_A8739_ & ~new_A8723_;
  assign new_A8741_ = new_A8723_ | new_A8738_;
  assign new_A8742_ = ~new_A8716_ | ~new_A8717_;
  assign new_A8743_ = new_A8723_ | new_A8738_;
  assign new_A8744_ = ~new_A8723_ & ~new_A8745_;
  assign new_A8745_ = new_A8723_ & new_A8738_;
  assign new_A8746_ = new_B1889_;
  assign new_A8747_ = new_B1922_;
  assign new_A8748_ = new_B1955_;
  assign new_A8749_ = new_B1988_;
  assign new_A8750_ = new_B2021_;
  assign new_A8751_ = new_A8757_ & new_A8756_;
  assign new_A8752_ = new_A8759_ | new_A8758_;
  assign new_A8753_ = new_A8761_ | new_A8760_;
  assign new_A8754_ = new_A8756_ & new_A8762_;
  assign new_A8755_ = new_A8756_ & new_A8763_;
  assign new_A8756_ = new_A8746_ ^ new_A8747_;
  assign new_A8757_ = new_A8758_ ^ new_A8748_;
  assign new_A8758_ = new_A8766_ & new_A8765_;
  assign new_A8759_ = new_A8764_ & new_A8748_;
  assign new_A8760_ = new_A8769_ & new_A8768_;
  assign new_A8761_ = new_A8767_ & new_A8748_;
  assign new_A8762_ = new_A8770_ | new_A8747_;
  assign new_A8763_ = ~new_A8748_ ^ new_A8760_;
  assign new_A8764_ = ~new_A8773_ | ~new_A8774_;
  assign new_A8765_ = new_A8749_ ^ new_A8756_;
  assign new_A8766_ = new_A8775_ & new_A8768_;
  assign new_A8767_ = ~new_A8777_ | ~new_A8776_;
  assign new_A8768_ = new_A8749_ | new_A8750_;
  assign new_A8769_ = new_A8749_ | new_A8756_;
  assign new_A8770_ = new_A8748_ & new_A8760_;
  assign new_A8771_ = ~new_A8747_ | ~new_A8748_;
  assign new_A8772_ = new_A8756_ & new_A8771_;
  assign new_A8773_ = ~new_A8772_ & ~new_A8756_;
  assign new_A8774_ = new_A8756_ | new_A8771_;
  assign new_A8775_ = ~new_A8749_ | ~new_A8750_;
  assign new_A8776_ = new_A8756_ | new_A8771_;
  assign new_A8777_ = ~new_A8756_ & ~new_A8778_;
  assign new_A8778_ = new_A8756_ & new_A8771_;
  assign new_A8779_ = new_B2054_;
  assign new_A8780_ = new_B2087_;
  assign new_A8781_ = new_B2120_;
  assign new_A8782_ = new_B2153_;
  assign new_A8783_ = new_B2186_;
  assign new_A8784_ = new_A8790_ & new_A8789_;
  assign new_A8785_ = new_A8792_ | new_A8791_;
  assign new_A8786_ = new_A8794_ | new_A8793_;
  assign new_A8787_ = new_A8789_ & new_A8795_;
  assign new_A8788_ = new_A8789_ & new_A8796_;
  assign new_A8789_ = new_A8779_ ^ new_A8780_;
  assign new_A8790_ = new_A8791_ ^ new_A8781_;
  assign new_A8791_ = new_A8799_ & new_A8798_;
  assign new_A8792_ = new_A8797_ & new_A8781_;
  assign new_A8793_ = new_A8802_ & new_A8801_;
  assign new_A8794_ = new_A8800_ & new_A8781_;
  assign new_A8795_ = new_A8803_ | new_A8780_;
  assign new_A8796_ = ~new_A8781_ ^ new_A8793_;
  assign new_A8797_ = ~new_A8806_ | ~new_A8807_;
  assign new_A8798_ = new_A8782_ ^ new_A8789_;
  assign new_A8799_ = new_A8808_ & new_A8801_;
  assign new_A8800_ = ~new_A8810_ | ~new_A8809_;
  assign new_A8801_ = new_A8782_ | new_A8783_;
  assign new_A8802_ = new_A8782_ | new_A8789_;
  assign new_A8803_ = new_A8781_ & new_A8793_;
  assign new_A8804_ = ~new_A8780_ | ~new_A8781_;
  assign new_A8805_ = new_A8789_ & new_A8804_;
  assign new_A8806_ = ~new_A8805_ & ~new_A8789_;
  assign new_A8807_ = new_A8789_ | new_A8804_;
  assign new_A8808_ = ~new_A8782_ | ~new_A8783_;
  assign new_A8809_ = new_A8789_ | new_A8804_;
  assign new_A8810_ = ~new_A8789_ & ~new_A8811_;
  assign new_A8811_ = new_A8789_ & new_A8804_;
  assign new_A8812_ = new_B2219_;
  assign new_A8813_ = new_B2252_;
  assign new_A8814_ = new_B2285_;
  assign new_A8815_ = new_B2318_;
  assign new_A8816_ = new_B2351_;
  assign new_A8817_ = new_A8823_ & new_A8822_;
  assign new_A8818_ = new_A8825_ | new_A8824_;
  assign new_A8819_ = new_A8827_ | new_A8826_;
  assign new_A8820_ = new_A8822_ & new_A8828_;
  assign new_A8821_ = new_A8822_ & new_A8829_;
  assign new_A8822_ = new_A8812_ ^ new_A8813_;
  assign new_A8823_ = new_A8824_ ^ new_A8814_;
  assign new_A8824_ = new_A8832_ & new_A8831_;
  assign new_A8825_ = new_A8830_ & new_A8814_;
  assign new_A8826_ = new_A8835_ & new_A8834_;
  assign new_A8827_ = new_A8833_ & new_A8814_;
  assign new_A8828_ = new_A8836_ | new_A8813_;
  assign new_A8829_ = ~new_A8814_ ^ new_A8826_;
  assign new_A8830_ = ~new_A8839_ | ~new_A8840_;
  assign new_A8831_ = new_A8815_ ^ new_A8822_;
  assign new_A8832_ = new_A8841_ & new_A8834_;
  assign new_A8833_ = ~new_A8843_ | ~new_A8842_;
  assign new_A8834_ = new_A8815_ | new_A8816_;
  assign new_A8835_ = new_A8815_ | new_A8822_;
  assign new_A8836_ = new_A8814_ & new_A8826_;
  assign new_A8837_ = ~new_A8813_ | ~new_A8814_;
  assign new_A8838_ = new_A8822_ & new_A8837_;
  assign new_A8839_ = ~new_A8838_ & ~new_A8822_;
  assign new_A8840_ = new_A8822_ | new_A8837_;
  assign new_A8841_ = ~new_A8815_ | ~new_A8816_;
  assign new_A8842_ = new_A8822_ | new_A8837_;
  assign new_A8843_ = ~new_A8822_ & ~new_A8844_;
  assign new_A8844_ = new_A8822_ & new_A8837_;
  assign new_A8845_ = new_B2384_;
  assign new_A8846_ = new_B2417_;
  assign new_A8847_ = new_B2450_;
  assign new_A8848_ = new_B2483_;
  assign new_A8849_ = new_B2516_;
  assign new_A8850_ = new_A8856_ & new_A8855_;
  assign new_A8851_ = new_A8858_ | new_A8857_;
  assign new_A8852_ = new_A8860_ | new_A8859_;
  assign new_A8853_ = new_A8855_ & new_A8861_;
  assign new_A8854_ = new_A8855_ & new_A8862_;
  assign new_A8855_ = new_A8845_ ^ new_A8846_;
  assign new_A8856_ = new_A8857_ ^ new_A8847_;
  assign new_A8857_ = new_A8865_ & new_A8864_;
  assign new_A8858_ = new_A8863_ & new_A8847_;
  assign new_A8859_ = new_A8868_ & new_A8867_;
  assign new_A8860_ = new_A8866_ & new_A8847_;
  assign new_A8861_ = new_A8869_ | new_A8846_;
  assign new_A8862_ = ~new_A8847_ ^ new_A8859_;
  assign new_A8863_ = ~new_A8872_ | ~new_A8873_;
  assign new_A8864_ = new_A8848_ ^ new_A8855_;
  assign new_A8865_ = new_A8874_ & new_A8867_;
  assign new_A8866_ = ~new_A8876_ | ~new_A8875_;
  assign new_A8867_ = new_A8848_ | new_A8849_;
  assign new_A8868_ = new_A8848_ | new_A8855_;
  assign new_A8869_ = new_A8847_ & new_A8859_;
  assign new_A8870_ = ~new_A8846_ | ~new_A8847_;
  assign new_A8871_ = new_A8855_ & new_A8870_;
  assign new_A8872_ = ~new_A8871_ & ~new_A8855_;
  assign new_A8873_ = new_A8855_ | new_A8870_;
  assign new_A8874_ = ~new_A8848_ | ~new_A8849_;
  assign new_A8875_ = new_A8855_ | new_A8870_;
  assign new_A8876_ = ~new_A8855_ & ~new_A8877_;
  assign new_A8877_ = new_A8855_ & new_A8870_;
  assign new_A8878_ = new_B2549_;
  assign new_A8879_ = new_B2582_;
  assign new_A8880_ = new_B2615_;
  assign new_A8881_ = new_B2648_;
  assign new_A8882_ = new_B2681_;
  assign new_A8883_ = new_A8889_ & new_A8888_;
  assign new_A8884_ = new_A8891_ | new_A8890_;
  assign new_A8885_ = new_A8893_ | new_A8892_;
  assign new_A8886_ = new_A8888_ & new_A8894_;
  assign new_A8887_ = new_A8888_ & new_A8895_;
  assign new_A8888_ = new_A8878_ ^ new_A8879_;
  assign new_A8889_ = new_A8890_ ^ new_A8880_;
  assign new_A8890_ = new_A8898_ & new_A8897_;
  assign new_A8891_ = new_A8896_ & new_A8880_;
  assign new_A8892_ = new_A8901_ & new_A8900_;
  assign new_A8893_ = new_A8899_ & new_A8880_;
  assign new_A8894_ = new_A8902_ | new_A8879_;
  assign new_A8895_ = ~new_A8880_ ^ new_A8892_;
  assign new_A8896_ = ~new_A8905_ | ~new_A8906_;
  assign new_A8897_ = new_A8881_ ^ new_A8888_;
  assign new_A8898_ = new_A8907_ & new_A8900_;
  assign new_A8899_ = ~new_A8909_ | ~new_A8908_;
  assign new_A8900_ = new_A8881_ | new_A8882_;
  assign new_A8901_ = new_A8881_ | new_A8888_;
  assign new_A8902_ = new_A8880_ & new_A8892_;
  assign new_A8903_ = ~new_A8879_ | ~new_A8880_;
  assign new_A8904_ = new_A8888_ & new_A8903_;
  assign new_A8905_ = ~new_A8904_ & ~new_A8888_;
  assign new_A8906_ = new_A8888_ | new_A8903_;
  assign new_A8907_ = ~new_A8881_ | ~new_A8882_;
  assign new_A8908_ = new_A8888_ | new_A8903_;
  assign new_A8909_ = ~new_A8888_ & ~new_A8910_;
  assign new_A8910_ = new_A8888_ & new_A8903_;
  assign new_A8911_ = new_B2714_;
  assign new_A8912_ = new_B2747_;
  assign new_A8913_ = new_B2780_;
  assign new_A8914_ = new_B2813_;
  assign new_A8915_ = new_B2846_;
  assign new_A8916_ = new_A8922_ & new_A8921_;
  assign new_A8917_ = new_A8924_ | new_A8923_;
  assign new_A8918_ = new_A8926_ | new_A8925_;
  assign new_A8919_ = new_A8921_ & new_A8927_;
  assign new_A8920_ = new_A8921_ & new_A8928_;
  assign new_A8921_ = new_A8911_ ^ new_A8912_;
  assign new_A8922_ = new_A8923_ ^ new_A8913_;
  assign new_A8923_ = new_A8931_ & new_A8930_;
  assign new_A8924_ = new_A8929_ & new_A8913_;
  assign new_A8925_ = new_A8934_ & new_A8933_;
  assign new_A8926_ = new_A8932_ & new_A8913_;
  assign new_A8927_ = new_A8935_ | new_A8912_;
  assign new_A8928_ = ~new_A8913_ ^ new_A8925_;
  assign new_A8929_ = ~new_A8938_ | ~new_A8939_;
  assign new_A8930_ = new_A8914_ ^ new_A8921_;
  assign new_A8931_ = new_A8940_ & new_A8933_;
  assign new_A8932_ = ~new_A8942_ | ~new_A8941_;
  assign new_A8933_ = new_A8914_ | new_A8915_;
  assign new_A8934_ = new_A8914_ | new_A8921_;
  assign new_A8935_ = new_A8913_ & new_A8925_;
  assign new_A8936_ = ~new_A8912_ | ~new_A8913_;
  assign new_A8937_ = new_A8921_ & new_A8936_;
  assign new_A8938_ = ~new_A8937_ & ~new_A8921_;
  assign new_A8939_ = new_A8921_ | new_A8936_;
  assign new_A8940_ = ~new_A8914_ | ~new_A8915_;
  assign new_A8941_ = new_A8921_ | new_A8936_;
  assign new_A8942_ = ~new_A8921_ & ~new_A8943_;
  assign new_A8943_ = new_A8921_ & new_A8936_;
  assign new_A8944_ = new_B2879_;
  assign new_A8945_ = new_B2912_;
  assign new_A8946_ = new_B2945_;
  assign new_A8947_ = new_B2978_;
  assign new_A8948_ = new_B3011_;
  assign new_A8949_ = new_A8955_ & new_A8954_;
  assign new_A8950_ = new_A8957_ | new_A8956_;
  assign new_A8951_ = new_A8959_ | new_A8958_;
  assign new_A8952_ = new_A8954_ & new_A8960_;
  assign new_A8953_ = new_A8954_ & new_A8961_;
  assign new_A8954_ = new_A8944_ ^ new_A8945_;
  assign new_A8955_ = new_A8956_ ^ new_A8946_;
  assign new_A8956_ = new_A8964_ & new_A8963_;
  assign new_A8957_ = new_A8962_ & new_A8946_;
  assign new_A8958_ = new_A8967_ & new_A8966_;
  assign new_A8959_ = new_A8965_ & new_A8946_;
  assign new_A8960_ = new_A8968_ | new_A8945_;
  assign new_A8961_ = ~new_A8946_ ^ new_A8958_;
  assign new_A8962_ = ~new_A8971_ | ~new_A8972_;
  assign new_A8963_ = new_A8947_ ^ new_A8954_;
  assign new_A8964_ = new_A8973_ & new_A8966_;
  assign new_A8965_ = ~new_A8975_ | ~new_A8974_;
  assign new_A8966_ = new_A8947_ | new_A8948_;
  assign new_A8967_ = new_A8947_ | new_A8954_;
  assign new_A8968_ = new_A8946_ & new_A8958_;
  assign new_A8969_ = ~new_A8945_ | ~new_A8946_;
  assign new_A8970_ = new_A8954_ & new_A8969_;
  assign new_A8971_ = ~new_A8970_ & ~new_A8954_;
  assign new_A8972_ = new_A8954_ | new_A8969_;
  assign new_A8973_ = ~new_A8947_ | ~new_A8948_;
  assign new_A8974_ = new_A8954_ | new_A8969_;
  assign new_A8975_ = ~new_A8954_ & ~new_A8976_;
  assign new_A8976_ = new_A8954_ & new_A8969_;
  assign new_A8977_ = new_B3044_;
  assign new_A8978_ = new_B3077_;
  assign new_A8979_ = new_B3110_;
  assign new_A8980_ = new_B3143_;
  assign new_A8981_ = new_B3176_;
  assign new_A8982_ = new_A8988_ & new_A8987_;
  assign new_A8983_ = new_A8990_ | new_A8989_;
  assign new_A8984_ = new_A8992_ | new_A8991_;
  assign new_A8985_ = new_A8987_ & new_A8993_;
  assign new_A8986_ = new_A8987_ & new_A8994_;
  assign new_A8987_ = new_A8977_ ^ new_A8978_;
  assign new_A8988_ = new_A8989_ ^ new_A8979_;
  assign new_A8989_ = new_A8997_ & new_A8996_;
  assign new_A8990_ = new_A8995_ & new_A8979_;
  assign new_A8991_ = new_A9000_ & new_A8999_;
  assign new_A8992_ = new_A8998_ & new_A8979_;
  assign new_A8993_ = new_A9001_ | new_A8978_;
  assign new_A8994_ = ~new_A8979_ ^ new_A8991_;
  assign new_A8995_ = ~new_A9004_ | ~new_A9005_;
  assign new_A8996_ = new_A8980_ ^ new_A8987_;
  assign new_A8997_ = new_A9006_ & new_A8999_;
  assign new_A8998_ = ~new_A9008_ | ~new_A9007_;
  assign new_A8999_ = new_A8980_ | new_A8981_;
  assign new_A9000_ = new_A8980_ | new_A8987_;
  assign new_A9001_ = new_A8979_ & new_A8991_;
  assign new_A9002_ = ~new_A8978_ | ~new_A8979_;
  assign new_A9003_ = new_A8987_ & new_A9002_;
  assign new_A9004_ = ~new_A9003_ & ~new_A8987_;
  assign new_A9005_ = new_A8987_ | new_A9002_;
  assign new_A9006_ = ~new_A8980_ | ~new_A8981_;
  assign new_A9007_ = new_A8987_ | new_A9002_;
  assign new_A9008_ = ~new_A8987_ & ~new_A9009_;
  assign new_A9009_ = new_A8987_ & new_A9002_;
  assign new_A9010_ = new_B3209_;
  assign new_A9011_ = new_B3242_;
  assign new_A9012_ = new_B3275_;
  assign new_A9013_ = new_B3308_;
  assign new_A9014_ = new_B3341_;
  assign new_A9015_ = new_A9021_ & new_A9020_;
  assign new_A9016_ = new_A9023_ | new_A9022_;
  assign new_A9017_ = new_A9025_ | new_A9024_;
  assign new_A9018_ = new_A9020_ & new_A9026_;
  assign new_A9019_ = new_A9020_ & new_A9027_;
  assign new_A9020_ = new_A9010_ ^ new_A9011_;
  assign new_A9021_ = new_A9022_ ^ new_A9012_;
  assign new_A9022_ = new_A9030_ & new_A9029_;
  assign new_A9023_ = new_A9028_ & new_A9012_;
  assign new_A9024_ = new_A9033_ & new_A9032_;
  assign new_A9025_ = new_A9031_ & new_A9012_;
  assign new_A9026_ = new_A9034_ | new_A9011_;
  assign new_A9027_ = ~new_A9012_ ^ new_A9024_;
  assign new_A9028_ = ~new_A9037_ | ~new_A9038_;
  assign new_A9029_ = new_A9013_ ^ new_A9020_;
  assign new_A9030_ = new_A9039_ & new_A9032_;
  assign new_A9031_ = ~new_A9041_ | ~new_A9040_;
  assign new_A9032_ = new_A9013_ | new_A9014_;
  assign new_A9033_ = new_A9013_ | new_A9020_;
  assign new_A9034_ = new_A9012_ & new_A9024_;
  assign new_A9035_ = ~new_A9011_ | ~new_A9012_;
  assign new_A9036_ = new_A9020_ & new_A9035_;
  assign new_A9037_ = ~new_A9036_ & ~new_A9020_;
  assign new_A9038_ = new_A9020_ | new_A9035_;
  assign new_A9039_ = ~new_A9013_ | ~new_A9014_;
  assign new_A9040_ = new_A9020_ | new_A9035_;
  assign new_A9041_ = ~new_A9020_ & ~new_A9042_;
  assign new_A9042_ = new_A9020_ & new_A9035_;
  assign new_A9043_ = new_B3374_;
  assign new_A9044_ = new_B3407_;
  assign new_A9045_ = new_B3440_;
  assign new_A9046_ = new_B3473_;
  assign new_A9047_ = new_B3506_;
  assign new_A9048_ = new_A9054_ & new_A9053_;
  assign new_A9049_ = new_A9056_ | new_A9055_;
  assign new_A9050_ = new_A9058_ | new_A9057_;
  assign new_A9051_ = new_A9053_ & new_A9059_;
  assign new_A9052_ = new_A9053_ & new_A9060_;
  assign new_A9053_ = new_A9043_ ^ new_A9044_;
  assign new_A9054_ = new_A9055_ ^ new_A9045_;
  assign new_A9055_ = new_A9063_ & new_A9062_;
  assign new_A9056_ = new_A9061_ & new_A9045_;
  assign new_A9057_ = new_A9066_ & new_A9065_;
  assign new_A9058_ = new_A9064_ & new_A9045_;
  assign new_A9059_ = new_A9067_ | new_A9044_;
  assign new_A9060_ = ~new_A9045_ ^ new_A9057_;
  assign new_A9061_ = ~new_A9070_ | ~new_A9071_;
  assign new_A9062_ = new_A9046_ ^ new_A9053_;
  assign new_A9063_ = new_A9072_ & new_A9065_;
  assign new_A9064_ = ~new_A9074_ | ~new_A9073_;
  assign new_A9065_ = new_A9046_ | new_A9047_;
  assign new_A9066_ = new_A9046_ | new_A9053_;
  assign new_A9067_ = new_A9045_ & new_A9057_;
  assign new_A9068_ = ~new_A9044_ | ~new_A9045_;
  assign new_A9069_ = new_A9053_ & new_A9068_;
  assign new_A9070_ = ~new_A9069_ & ~new_A9053_;
  assign new_A9071_ = new_A9053_ | new_A9068_;
  assign new_A9072_ = ~new_A9046_ | ~new_A9047_;
  assign new_A9073_ = new_A9053_ | new_A9068_;
  assign new_A9074_ = ~new_A9053_ & ~new_A9075_;
  assign new_A9075_ = new_A9053_ & new_A9068_;
  assign new_A9076_ = new_B3539_;
  assign new_A9077_ = new_B3572_;
  assign new_A9078_ = new_B3605_;
  assign new_A9079_ = new_B3638_;
  assign new_A9080_ = new_B3671_;
  assign new_A9081_ = new_A9087_ & new_A9086_;
  assign new_A9082_ = new_A9089_ | new_A9088_;
  assign new_A9083_ = new_A9091_ | new_A9090_;
  assign new_A9084_ = new_A9086_ & new_A9092_;
  assign new_A9085_ = new_A9086_ & new_A9093_;
  assign new_A9086_ = new_A9076_ ^ new_A9077_;
  assign new_A9087_ = new_A9088_ ^ new_A9078_;
  assign new_A9088_ = new_A9096_ & new_A9095_;
  assign new_A9089_ = new_A9094_ & new_A9078_;
  assign new_A9090_ = new_A9099_ & new_A9098_;
  assign new_A9091_ = new_A9097_ & new_A9078_;
  assign new_A9092_ = new_A9100_ | new_A9077_;
  assign new_A9093_ = ~new_A9078_ ^ new_A9090_;
  assign new_A9094_ = ~new_A9103_ | ~new_A9104_;
  assign new_A9095_ = new_A9079_ ^ new_A9086_;
  assign new_A9096_ = new_A9105_ & new_A9098_;
  assign new_A9097_ = ~new_A9107_ | ~new_A9106_;
  assign new_A9098_ = new_A9079_ | new_A9080_;
  assign new_A9099_ = new_A9079_ | new_A9086_;
  assign new_A9100_ = new_A9078_ & new_A9090_;
  assign new_A9101_ = ~new_A9077_ | ~new_A9078_;
  assign new_A9102_ = new_A9086_ & new_A9101_;
  assign new_A9103_ = ~new_A9102_ & ~new_A9086_;
  assign new_A9104_ = new_A9086_ | new_A9101_;
  assign new_A9105_ = ~new_A9079_ | ~new_A9080_;
  assign new_A9106_ = new_A9086_ | new_A9101_;
  assign new_A9107_ = ~new_A9086_ & ~new_A9108_;
  assign new_A9108_ = new_A9086_ & new_A9101_;
  assign new_A9109_ = new_B3704_;
  assign new_A9110_ = new_B3737_;
  assign new_A9111_ = new_B3770_;
  assign new_A9112_ = new_B3803_;
  assign new_A9113_ = new_B3836_;
  assign new_A9114_ = new_A9120_ & new_A9119_;
  assign new_A9115_ = new_A9122_ | new_A9121_;
  assign new_A9116_ = new_A9124_ | new_A9123_;
  assign new_A9117_ = new_A9119_ & new_A9125_;
  assign new_A9118_ = new_A9119_ & new_A9126_;
  assign new_A9119_ = new_A9109_ ^ new_A9110_;
  assign new_A9120_ = new_A9121_ ^ new_A9111_;
  assign new_A9121_ = new_A9129_ & new_A9128_;
  assign new_A9122_ = new_A9127_ & new_A9111_;
  assign new_A9123_ = new_A9132_ & new_A9131_;
  assign new_A9124_ = new_A9130_ & new_A9111_;
  assign new_A9125_ = new_A9133_ | new_A9110_;
  assign new_A9126_ = ~new_A9111_ ^ new_A9123_;
  assign new_A9127_ = ~new_A9136_ | ~new_A9137_;
  assign new_A9128_ = new_A9112_ ^ new_A9119_;
  assign new_A9129_ = new_A9138_ & new_A9131_;
  assign new_A9130_ = ~new_A9140_ | ~new_A9139_;
  assign new_A9131_ = new_A9112_ | new_A9113_;
  assign new_A9132_ = new_A9112_ | new_A9119_;
  assign new_A9133_ = new_A9111_ & new_A9123_;
  assign new_A9134_ = ~new_A9110_ | ~new_A9111_;
  assign new_A9135_ = new_A9119_ & new_A9134_;
  assign new_A9136_ = ~new_A9135_ & ~new_A9119_;
  assign new_A9137_ = new_A9119_ | new_A9134_;
  assign new_A9138_ = ~new_A9112_ | ~new_A9113_;
  assign new_A9139_ = new_A9119_ | new_A9134_;
  assign new_A9140_ = ~new_A9119_ & ~new_A9141_;
  assign new_A9141_ = new_A9119_ & new_A9134_;
  assign new_A9142_ = new_B3869_;
  assign new_A9143_ = new_B3902_;
  assign new_A9144_ = new_B3935_;
  assign new_A9145_ = new_B3968_;
  assign new_A9146_ = new_B4001_;
  assign new_A9147_ = new_A9153_ & new_A9152_;
  assign new_A9148_ = new_A9155_ | new_A9154_;
  assign new_A9149_ = new_A9157_ | new_A9156_;
  assign new_A9150_ = new_A9152_ & new_A9158_;
  assign new_A9151_ = new_A9152_ & new_A9159_;
  assign new_A9152_ = new_A9142_ ^ new_A9143_;
  assign new_A9153_ = new_A9154_ ^ new_A9144_;
  assign new_A9154_ = new_A9162_ & new_A9161_;
  assign new_A9155_ = new_A9160_ & new_A9144_;
  assign new_A9156_ = new_A9165_ & new_A9164_;
  assign new_A9157_ = new_A9163_ & new_A9144_;
  assign new_A9158_ = new_A9166_ | new_A9143_;
  assign new_A9159_ = ~new_A9144_ ^ new_A9156_;
  assign new_A9160_ = ~new_A9169_ | ~new_A9170_;
  assign new_A9161_ = new_A9145_ ^ new_A9152_;
  assign new_A9162_ = new_A9171_ & new_A9164_;
  assign new_A9163_ = ~new_A9173_ | ~new_A9172_;
  assign new_A9164_ = new_A9145_ | new_A9146_;
  assign new_A9165_ = new_A9145_ | new_A9152_;
  assign new_A9166_ = new_A9144_ & new_A9156_;
  assign new_A9167_ = ~new_A9143_ | ~new_A9144_;
  assign new_A9168_ = new_A9152_ & new_A9167_;
  assign new_A9169_ = ~new_A9168_ & ~new_A9152_;
  assign new_A9170_ = new_A9152_ | new_A9167_;
  assign new_A9171_ = ~new_A9145_ | ~new_A9146_;
  assign new_A9172_ = new_A9152_ | new_A9167_;
  assign new_A9173_ = ~new_A9152_ & ~new_A9174_;
  assign new_A9174_ = new_A9152_ & new_A9167_;
  assign new_A9175_ = new_B4034_;
  assign new_A9176_ = new_B4067_;
  assign new_A9177_ = new_B4100_;
  assign new_A9178_ = new_B4133_;
  assign new_A9179_ = new_B4166_;
  assign new_A9180_ = new_A9186_ & new_A9185_;
  assign new_A9181_ = new_A9188_ | new_A9187_;
  assign new_A9182_ = new_A9190_ | new_A9189_;
  assign new_A9183_ = new_A9185_ & new_A9191_;
  assign new_A9184_ = new_A9185_ & new_A9192_;
  assign new_A9185_ = new_A9175_ ^ new_A9176_;
  assign new_A9186_ = new_A9187_ ^ new_A9177_;
  assign new_A9187_ = new_A9195_ & new_A9194_;
  assign new_A9188_ = new_A9193_ & new_A9177_;
  assign new_A9189_ = new_A9198_ & new_A9197_;
  assign new_A9190_ = new_A9196_ & new_A9177_;
  assign new_A9191_ = new_A9199_ | new_A9176_;
  assign new_A9192_ = ~new_A9177_ ^ new_A9189_;
  assign new_A9193_ = ~new_A9202_ | ~new_A9203_;
  assign new_A9194_ = new_A9178_ ^ new_A9185_;
  assign new_A9195_ = new_A9204_ & new_A9197_;
  assign new_A9196_ = ~new_A9206_ | ~new_A9205_;
  assign new_A9197_ = new_A9178_ | new_A9179_;
  assign new_A9198_ = new_A9178_ | new_A9185_;
  assign new_A9199_ = new_A9177_ & new_A9189_;
  assign new_A9200_ = ~new_A9176_ | ~new_A9177_;
  assign new_A9201_ = new_A9185_ & new_A9200_;
  assign new_A9202_ = ~new_A9201_ & ~new_A9185_;
  assign new_A9203_ = new_A9185_ | new_A9200_;
  assign new_A9204_ = ~new_A9178_ | ~new_A9179_;
  assign new_A9205_ = new_A9185_ | new_A9200_;
  assign new_A9206_ = ~new_A9185_ & ~new_A9207_;
  assign new_A9207_ = new_A9185_ & new_A9200_;
  assign new_A9208_ = new_B4199_;
  assign new_A9209_ = new_B4232_;
  assign new_A9210_ = new_B4265_;
  assign new_A9211_ = new_B4298_;
  assign new_A9212_ = new_B4331_;
  assign new_A9213_ = new_A9219_ & new_A9218_;
  assign new_A9214_ = new_A9221_ | new_A9220_;
  assign new_A9215_ = new_A9223_ | new_A9222_;
  assign new_A9216_ = new_A9218_ & new_A9224_;
  assign new_A9217_ = new_A9218_ & new_A9225_;
  assign new_A9218_ = new_A9208_ ^ new_A9209_;
  assign new_A9219_ = new_A9220_ ^ new_A9210_;
  assign new_A9220_ = new_A9228_ & new_A9227_;
  assign new_A9221_ = new_A9226_ & new_A9210_;
  assign new_A9222_ = new_A9231_ & new_A9230_;
  assign new_A9223_ = new_A9229_ & new_A9210_;
  assign new_A9224_ = new_A9232_ | new_A9209_;
  assign new_A9225_ = ~new_A9210_ ^ new_A9222_;
  assign new_A9226_ = ~new_A9235_ | ~new_A9236_;
  assign new_A9227_ = new_A9211_ ^ new_A9218_;
  assign new_A9228_ = new_A9237_ & new_A9230_;
  assign new_A9229_ = ~new_A9239_ | ~new_A9238_;
  assign new_A9230_ = new_A9211_ | new_A9212_;
  assign new_A9231_ = new_A9211_ | new_A9218_;
  assign new_A9232_ = new_A9210_ & new_A9222_;
  assign new_A9233_ = ~new_A9209_ | ~new_A9210_;
  assign new_A9234_ = new_A9218_ & new_A9233_;
  assign new_A9235_ = ~new_A9234_ & ~new_A9218_;
  assign new_A9236_ = new_A9218_ | new_A9233_;
  assign new_A9237_ = ~new_A9211_ | ~new_A9212_;
  assign new_A9238_ = new_A9218_ | new_A9233_;
  assign new_A9239_ = ~new_A9218_ & ~new_A9240_;
  assign new_A9240_ = new_A9218_ & new_A9233_;
  assign new_A9241_ = new_B4364_;
  assign new_A9242_ = new_B4397_;
  assign new_A9243_ = new_B4430_;
  assign new_A9244_ = new_B4463_;
  assign new_A9245_ = new_B4496_;
  assign new_A9246_ = new_A9252_ & new_A9251_;
  assign new_A9247_ = new_A9254_ | new_A9253_;
  assign new_A9248_ = new_A9256_ | new_A9255_;
  assign new_A9249_ = new_A9251_ & new_A9257_;
  assign new_A9250_ = new_A9251_ & new_A9258_;
  assign new_A9251_ = new_A9241_ ^ new_A9242_;
  assign new_A9252_ = new_A9253_ ^ new_A9243_;
  assign new_A9253_ = new_A9261_ & new_A9260_;
  assign new_A9254_ = new_A9259_ & new_A9243_;
  assign new_A9255_ = new_A9264_ & new_A9263_;
  assign new_A9256_ = new_A9262_ & new_A9243_;
  assign new_A9257_ = new_A9265_ | new_A9242_;
  assign new_A9258_ = ~new_A9243_ ^ new_A9255_;
  assign new_A9259_ = ~new_A9268_ | ~new_A9269_;
  assign new_A9260_ = new_A9244_ ^ new_A9251_;
  assign new_A9261_ = new_A9270_ & new_A9263_;
  assign new_A9262_ = ~new_A9272_ | ~new_A9271_;
  assign new_A9263_ = new_A9244_ | new_A9245_;
  assign new_A9264_ = new_A9244_ | new_A9251_;
  assign new_A9265_ = new_A9243_ & new_A9255_;
  assign new_A9266_ = ~new_A9242_ | ~new_A9243_;
  assign new_A9267_ = new_A9251_ & new_A9266_;
  assign new_A9268_ = ~new_A9267_ & ~new_A9251_;
  assign new_A9269_ = new_A9251_ | new_A9266_;
  assign new_A9270_ = ~new_A9244_ | ~new_A9245_;
  assign new_A9271_ = new_A9251_ | new_A9266_;
  assign new_A9272_ = ~new_A9251_ & ~new_A9273_;
  assign new_A9273_ = new_A9251_ & new_A9266_;
  assign new_A9274_ = new_B4529_;
  assign new_A9275_ = new_B4562_;
  assign new_A9276_ = new_B4595_;
  assign new_A9277_ = new_B4628_;
  assign new_A9278_ = new_B4661_;
  assign new_A9279_ = new_A9285_ & new_A9284_;
  assign new_A9280_ = new_A9287_ | new_A9286_;
  assign new_A9281_ = new_A9289_ | new_A9288_;
  assign new_A9282_ = new_A9284_ & new_A9290_;
  assign new_A9283_ = new_A9284_ & new_A9291_;
  assign new_A9284_ = new_A9274_ ^ new_A9275_;
  assign new_A9285_ = new_A9286_ ^ new_A9276_;
  assign new_A9286_ = new_A9294_ & new_A9293_;
  assign new_A9287_ = new_A9292_ & new_A9276_;
  assign new_A9288_ = new_A9297_ & new_A9296_;
  assign new_A9289_ = new_A9295_ & new_A9276_;
  assign new_A9290_ = new_A9298_ | new_A9275_;
  assign new_A9291_ = ~new_A9276_ ^ new_A9288_;
  assign new_A9292_ = ~new_A9301_ | ~new_A9302_;
  assign new_A9293_ = new_A9277_ ^ new_A9284_;
  assign new_A9294_ = new_A9303_ & new_A9296_;
  assign new_A9295_ = ~new_A9305_ | ~new_A9304_;
  assign new_A9296_ = new_A9277_ | new_A9278_;
  assign new_A9297_ = new_A9277_ | new_A9284_;
  assign new_A9298_ = new_A9276_ & new_A9288_;
  assign new_A9299_ = ~new_A9275_ | ~new_A9276_;
  assign new_A9300_ = new_A9284_ & new_A9299_;
  assign new_A9301_ = ~new_A9300_ & ~new_A9284_;
  assign new_A9302_ = new_A9284_ | new_A9299_;
  assign new_A9303_ = ~new_A9277_ | ~new_A9278_;
  assign new_A9304_ = new_A9284_ | new_A9299_;
  assign new_A9305_ = ~new_A9284_ & ~new_A9306_;
  assign new_A9306_ = new_A9284_ & new_A9299_;
  assign new_A9307_ = new_B4694_;
  assign new_A9308_ = new_B4727_;
  assign new_A9309_ = new_B4760_;
  assign new_A9310_ = new_B4793_;
  assign new_A9311_ = new_B4826_;
  assign new_A9312_ = new_A9318_ & new_A9317_;
  assign new_A9313_ = new_A9320_ | new_A9319_;
  assign new_A9314_ = new_A9322_ | new_A9321_;
  assign new_A9315_ = new_A9317_ & new_A9323_;
  assign new_A9316_ = new_A9317_ & new_A9324_;
  assign new_A9317_ = new_A9307_ ^ new_A9308_;
  assign new_A9318_ = new_A9319_ ^ new_A9309_;
  assign new_A9319_ = new_A9327_ & new_A9326_;
  assign new_A9320_ = new_A9325_ & new_A9309_;
  assign new_A9321_ = new_A9330_ & new_A9329_;
  assign new_A9322_ = new_A9328_ & new_A9309_;
  assign new_A9323_ = new_A9331_ | new_A9308_;
  assign new_A9324_ = ~new_A9309_ ^ new_A9321_;
  assign new_A9325_ = ~new_A9334_ | ~new_A9335_;
  assign new_A9326_ = new_A9310_ ^ new_A9317_;
  assign new_A9327_ = new_A9336_ & new_A9329_;
  assign new_A9328_ = ~new_A9338_ | ~new_A9337_;
  assign new_A9329_ = new_A9310_ | new_A9311_;
  assign new_A9330_ = new_A9310_ | new_A9317_;
  assign new_A9331_ = new_A9309_ & new_A9321_;
  assign new_A9332_ = ~new_A9308_ | ~new_A9309_;
  assign new_A9333_ = new_A9317_ & new_A9332_;
  assign new_A9334_ = ~new_A9333_ & ~new_A9317_;
  assign new_A9335_ = new_A9317_ | new_A9332_;
  assign new_A9336_ = ~new_A9310_ | ~new_A9311_;
  assign new_A9337_ = new_A9317_ | new_A9332_;
  assign new_A9338_ = ~new_A9317_ & ~new_A9339_;
  assign new_A9339_ = new_A9317_ & new_A9332_;
  assign new_A9340_ = new_B4859_;
  assign new_A9341_ = new_B4892_;
  assign new_A9342_ = new_B4925_;
  assign new_A9343_ = new_B4958_;
  assign new_A9344_ = new_B4991_;
  assign new_A9345_ = new_A9351_ & new_A9350_;
  assign new_A9346_ = new_A9353_ | new_A9352_;
  assign new_A9347_ = new_A9355_ | new_A9354_;
  assign new_A9348_ = new_A9350_ & new_A9356_;
  assign new_A9349_ = new_A9350_ & new_A9357_;
  assign new_A9350_ = new_A9340_ ^ new_A9341_;
  assign new_A9351_ = new_A9352_ ^ new_A9342_;
  assign new_A9352_ = new_A9360_ & new_A9359_;
  assign new_A9353_ = new_A9358_ & new_A9342_;
  assign new_A9354_ = new_A9363_ & new_A9362_;
  assign new_A9355_ = new_A9361_ & new_A9342_;
  assign new_A9356_ = new_A9364_ | new_A9341_;
  assign new_A9357_ = ~new_A9342_ ^ new_A9354_;
  assign new_A9358_ = ~new_A9367_ | ~new_A9368_;
  assign new_A9359_ = new_A9343_ ^ new_A9350_;
  assign new_A9360_ = new_A9369_ & new_A9362_;
  assign new_A9361_ = ~new_A9371_ | ~new_A9370_;
  assign new_A9362_ = new_A9343_ | new_A9344_;
  assign new_A9363_ = new_A9343_ | new_A9350_;
  assign new_A9364_ = new_A9342_ & new_A9354_;
  assign new_A9365_ = ~new_A9341_ | ~new_A9342_;
  assign new_A9366_ = new_A9350_ & new_A9365_;
  assign new_A9367_ = ~new_A9366_ & ~new_A9350_;
  assign new_A9368_ = new_A9350_ | new_A9365_;
  assign new_A9369_ = ~new_A9343_ | ~new_A9344_;
  assign new_A9370_ = new_A9350_ | new_A9365_;
  assign new_A9371_ = ~new_A9350_ & ~new_A9372_;
  assign new_A9372_ = new_A9350_ & new_A9365_;
  assign new_A9373_ = new_B5024_;
  assign new_A9374_ = new_B5057_;
  assign new_A9375_ = new_B5090_;
  assign new_A9376_ = new_B5123_;
  assign new_A9377_ = new_B5156_;
  assign new_A9378_ = new_A9384_ & new_A9383_;
  assign new_A9379_ = new_A9386_ | new_A9385_;
  assign new_A9380_ = new_A9388_ | new_A9387_;
  assign new_A9381_ = new_A9383_ & new_A9389_;
  assign new_A9382_ = new_A9383_ & new_A9390_;
  assign new_A9383_ = new_A9373_ ^ new_A9374_;
  assign new_A9384_ = new_A9385_ ^ new_A9375_;
  assign new_A9385_ = new_A9393_ & new_A9392_;
  assign new_A9386_ = new_A9391_ & new_A9375_;
  assign new_A9387_ = new_A9396_ & new_A9395_;
  assign new_A9388_ = new_A9394_ & new_A9375_;
  assign new_A9389_ = new_A9397_ | new_A9374_;
  assign new_A9390_ = ~new_A9375_ ^ new_A9387_;
  assign new_A9391_ = ~new_A9400_ | ~new_A9401_;
  assign new_A9392_ = new_A9376_ ^ new_A9383_;
  assign new_A9393_ = new_A9402_ & new_A9395_;
  assign new_A9394_ = ~new_A9404_ | ~new_A9403_;
  assign new_A9395_ = new_A9376_ | new_A9377_;
  assign new_A9396_ = new_A9376_ | new_A9383_;
  assign new_A9397_ = new_A9375_ & new_A9387_;
  assign new_A9398_ = ~new_A9374_ | ~new_A9375_;
  assign new_A9399_ = new_A9383_ & new_A9398_;
  assign new_A9400_ = ~new_A9399_ & ~new_A9383_;
  assign new_A9401_ = new_A9383_ | new_A9398_;
  assign new_A9402_ = ~new_A9376_ | ~new_A9377_;
  assign new_A9403_ = new_A9383_ | new_A9398_;
  assign new_A9404_ = ~new_A9383_ & ~new_A9405_;
  assign new_A9405_ = new_A9383_ & new_A9398_;
  assign new_A9406_ = new_B1063_;
  assign new_A9407_ = new_B1098_;
  assign new_A9408_ = new_B1131_;
  assign new_A9409_ = new_B1164_;
  assign new_A9410_ = new_B1197_;
  assign new_A9411_ = new_A9417_ & new_A9416_;
  assign new_A9412_ = new_A9419_ | new_A9418_;
  assign new_A9413_ = new_A9421_ | new_A9420_;
  assign new_A9414_ = new_A9416_ & new_A9422_;
  assign new_A9415_ = new_A9416_ & new_A9423_;
  assign new_A9416_ = new_A9406_ ^ new_A9407_;
  assign new_A9417_ = new_A9418_ ^ new_A9408_;
  assign new_A9418_ = new_A9426_ & new_A9425_;
  assign new_A9419_ = new_A9424_ & new_A9408_;
  assign new_A9420_ = new_A9429_ & new_A9428_;
  assign new_A9421_ = new_A9427_ & new_A9408_;
  assign new_A9422_ = new_A9430_ | new_A9407_;
  assign new_A9423_ = ~new_A9408_ ^ new_A9420_;
  assign new_A9424_ = ~new_A9433_ | ~new_A9434_;
  assign new_A9425_ = new_A9409_ ^ new_A9416_;
  assign new_A9426_ = new_A9435_ & new_A9428_;
  assign new_A9427_ = ~new_A9437_ | ~new_A9436_;
  assign new_A9428_ = new_A9409_ | new_A9410_;
  assign new_A9429_ = new_A9409_ | new_A9416_;
  assign new_A9430_ = new_A9408_ & new_A9420_;
  assign new_A9431_ = ~new_A9407_ | ~new_A9408_;
  assign new_A9432_ = new_A9416_ & new_A9431_;
  assign new_A9433_ = ~new_A9432_ & ~new_A9416_;
  assign new_A9434_ = new_A9416_ | new_A9431_;
  assign new_A9435_ = ~new_A9409_ | ~new_A9410_;
  assign new_A9436_ = new_A9416_ | new_A9431_;
  assign new_A9437_ = ~new_A9416_ & ~new_A9438_;
  assign new_A9438_ = new_A9416_ & new_A9431_;
  assign new_A9439_ = new_B1230_;
  assign new_A9440_ = new_B1263_;
  assign new_A9441_ = new_B1296_;
  assign new_A9442_ = new_B1329_;
  assign new_A9443_ = new_B1362_;
  assign new_A9444_ = new_A9450_ & new_A9449_;
  assign new_A9445_ = new_A9452_ | new_A9451_;
  assign new_A9446_ = new_A9454_ | new_A9453_;
  assign new_A9447_ = new_A9449_ & new_A9455_;
  assign new_A9448_ = new_A9449_ & new_A9456_;
  assign new_A9449_ = new_A9439_ ^ new_A9440_;
  assign new_A9450_ = new_A9451_ ^ new_A9441_;
  assign new_A9451_ = new_A9459_ & new_A9458_;
  assign new_A9452_ = new_A9457_ & new_A9441_;
  assign new_A9453_ = new_A9462_ & new_A9461_;
  assign new_A9454_ = new_A9460_ & new_A9441_;
  assign new_A9455_ = new_A9463_ | new_A9440_;
  assign new_A9456_ = ~new_A9441_ ^ new_A9453_;
  assign new_A9457_ = ~new_A9466_ | ~new_A9467_;
  assign new_A9458_ = new_A9442_ ^ new_A9449_;
  assign new_A9459_ = new_A9468_ & new_A9461_;
  assign new_A9460_ = ~new_A9470_ | ~new_A9469_;
  assign new_A9461_ = new_A9442_ | new_A9443_;
  assign new_A9462_ = new_A9442_ | new_A9449_;
  assign new_A9463_ = new_A9441_ & new_A9453_;
  assign new_A9464_ = ~new_A9440_ | ~new_A9441_;
  assign new_A9465_ = new_A9449_ & new_A9464_;
  assign new_A9466_ = ~new_A9465_ & ~new_A9449_;
  assign new_A9467_ = new_A9449_ | new_A9464_;
  assign new_A9468_ = ~new_A9442_ | ~new_A9443_;
  assign new_A9469_ = new_A9449_ | new_A9464_;
  assign new_A9470_ = ~new_A9449_ & ~new_A9471_;
  assign new_A9471_ = new_A9449_ & new_A9464_;
  assign new_A9472_ = new_B1395_;
  assign new_A9473_ = new_B1428_;
  assign new_A9474_ = new_B1461_;
  assign new_A9475_ = new_B1494_;
  assign new_A9476_ = new_B1527_;
  assign new_A9477_ = new_A9483_ & new_A9482_;
  assign new_A9478_ = new_A9485_ | new_A9484_;
  assign new_A9479_ = new_A9487_ | new_A9486_;
  assign new_A9480_ = new_A9482_ & new_A9488_;
  assign new_A9481_ = new_A9482_ & new_A9489_;
  assign new_A9482_ = new_A9472_ ^ new_A9473_;
  assign new_A9483_ = new_A9484_ ^ new_A9474_;
  assign new_A9484_ = new_A9492_ & new_A9491_;
  assign new_A9485_ = new_A9490_ & new_A9474_;
  assign new_A9486_ = new_A9495_ & new_A9494_;
  assign new_A9487_ = new_A9493_ & new_A9474_;
  assign new_A9488_ = new_A9496_ | new_A9473_;
  assign new_A9489_ = ~new_A9474_ ^ new_A9486_;
  assign new_A9490_ = ~new_A9499_ | ~new_A9500_;
  assign new_A9491_ = new_A9475_ ^ new_A9482_;
  assign new_A9492_ = new_A9501_ & new_A9494_;
  assign new_A9493_ = ~new_A9503_ | ~new_A9502_;
  assign new_A9494_ = new_A9475_ | new_A9476_;
  assign new_A9495_ = new_A9475_ | new_A9482_;
  assign new_A9496_ = new_A9474_ & new_A9486_;
  assign new_A9497_ = ~new_A9473_ | ~new_A9474_;
  assign new_A9498_ = new_A9482_ & new_A9497_;
  assign new_A9499_ = ~new_A9498_ & ~new_A9482_;
  assign new_A9500_ = new_A9482_ | new_A9497_;
  assign new_A9501_ = ~new_A9475_ | ~new_A9476_;
  assign new_A9502_ = new_A9482_ | new_A9497_;
  assign new_A9503_ = ~new_A9482_ & ~new_A9504_;
  assign new_A9504_ = new_A9482_ & new_A9497_;
  assign new_A9505_ = new_B1560_;
  assign new_A9506_ = new_B1593_;
  assign new_A9507_ = new_B1626_;
  assign new_A9508_ = new_B1659_;
  assign new_A9509_ = new_B1692_;
  assign new_A9510_ = new_A9516_ & new_A9515_;
  assign new_A9511_ = new_A9518_ | new_A9517_;
  assign new_A9512_ = new_A9520_ | new_A9519_;
  assign new_A9513_ = new_A9515_ & new_A9521_;
  assign new_A9514_ = new_A9515_ & new_A9522_;
  assign new_A9515_ = new_A9505_ ^ new_A9506_;
  assign new_A9516_ = new_A9517_ ^ new_A9507_;
  assign new_A9517_ = new_A9525_ & new_A9524_;
  assign new_A9518_ = new_A9523_ & new_A9507_;
  assign new_A9519_ = new_A9528_ & new_A9527_;
  assign new_A9520_ = new_A9526_ & new_A9507_;
  assign new_A9521_ = new_A9529_ | new_A9506_;
  assign new_A9522_ = ~new_A9507_ ^ new_A9519_;
  assign new_A9523_ = ~new_A9532_ | ~new_A9533_;
  assign new_A9524_ = new_A9508_ ^ new_A9515_;
  assign new_A9525_ = new_A9534_ & new_A9527_;
  assign new_A9526_ = ~new_A9536_ | ~new_A9535_;
  assign new_A9527_ = new_A9508_ | new_A9509_;
  assign new_A9528_ = new_A9508_ | new_A9515_;
  assign new_A9529_ = new_A9507_ & new_A9519_;
  assign new_A9530_ = ~new_A9506_ | ~new_A9507_;
  assign new_A9531_ = new_A9515_ & new_A9530_;
  assign new_A9532_ = ~new_A9531_ & ~new_A9515_;
  assign new_A9533_ = new_A9515_ | new_A9530_;
  assign new_A9534_ = ~new_A9508_ | ~new_A9509_;
  assign new_A9535_ = new_A9515_ | new_A9530_;
  assign new_A9536_ = ~new_A9515_ & ~new_A9537_;
  assign new_A9537_ = new_A9515_ & new_A9530_;
  assign new_A9538_ = new_B1725_;
  assign new_A9539_ = new_B1758_;
  assign new_A9540_ = new_B1791_;
  assign new_A9541_ = new_B1824_;
  assign new_A9542_ = new_B1857_;
  assign new_A9543_ = new_A9549_ & new_A9548_;
  assign new_A9544_ = new_A9551_ | new_A9550_;
  assign new_A9545_ = new_A9553_ | new_A9552_;
  assign new_A9546_ = new_A9548_ & new_A9554_;
  assign new_A9547_ = new_A9548_ & new_A9555_;
  assign new_A9548_ = new_A9538_ ^ new_A9539_;
  assign new_A9549_ = new_A9550_ ^ new_A9540_;
  assign new_A9550_ = new_A9558_ & new_A9557_;
  assign new_A9551_ = new_A9556_ & new_A9540_;
  assign new_A9552_ = new_A9561_ & new_A9560_;
  assign new_A9553_ = new_A9559_ & new_A9540_;
  assign new_A9554_ = new_A9562_ | new_A9539_;
  assign new_A9555_ = ~new_A9540_ ^ new_A9552_;
  assign new_A9556_ = ~new_A9565_ | ~new_A9566_;
  assign new_A9557_ = new_A9541_ ^ new_A9548_;
  assign new_A9558_ = new_A9567_ & new_A9560_;
  assign new_A9559_ = ~new_A9569_ | ~new_A9568_;
  assign new_A9560_ = new_A9541_ | new_A9542_;
  assign new_A9561_ = new_A9541_ | new_A9548_;
  assign new_A9562_ = new_A9540_ & new_A9552_;
  assign new_A9563_ = ~new_A9539_ | ~new_A9540_;
  assign new_A9564_ = new_A9548_ & new_A9563_;
  assign new_A9565_ = ~new_A9564_ & ~new_A9548_;
  assign new_A9566_ = new_A9548_ | new_A9563_;
  assign new_A9567_ = ~new_A9541_ | ~new_A9542_;
  assign new_A9568_ = new_A9548_ | new_A9563_;
  assign new_A9569_ = ~new_A9548_ & ~new_A9570_;
  assign new_A9570_ = new_A9548_ & new_A9563_;
  assign new_A9571_ = new_B1890_;
  assign new_A9572_ = new_B1923_;
  assign new_A9573_ = new_B1956_;
  assign new_A9574_ = new_B1989_;
  assign new_A9575_ = new_B2022_;
  assign new_A9576_ = new_A9582_ & new_A9581_;
  assign new_A9577_ = new_A9584_ | new_A9583_;
  assign new_A9578_ = new_A9586_ | new_A9585_;
  assign new_A9579_ = new_A9581_ & new_A9587_;
  assign new_A9580_ = new_A9581_ & new_A9588_;
  assign new_A9581_ = new_A9571_ ^ new_A9572_;
  assign new_A9582_ = new_A9583_ ^ new_A9573_;
  assign new_A9583_ = new_A9591_ & new_A9590_;
  assign new_A9584_ = new_A9589_ & new_A9573_;
  assign new_A9585_ = new_A9594_ & new_A9593_;
  assign new_A9586_ = new_A9592_ & new_A9573_;
  assign new_A9587_ = new_A9595_ | new_A9572_;
  assign new_A9588_ = ~new_A9573_ ^ new_A9585_;
  assign new_A9589_ = ~new_A9598_ | ~new_A9599_;
  assign new_A9590_ = new_A9574_ ^ new_A9581_;
  assign new_A9591_ = new_A9600_ & new_A9593_;
  assign new_A9592_ = ~new_A9602_ | ~new_A9601_;
  assign new_A9593_ = new_A9574_ | new_A9575_;
  assign new_A9594_ = new_A9574_ | new_A9581_;
  assign new_A9595_ = new_A9573_ & new_A9585_;
  assign new_A9596_ = ~new_A9572_ | ~new_A9573_;
  assign new_A9597_ = new_A9581_ & new_A9596_;
  assign new_A9598_ = ~new_A9597_ & ~new_A9581_;
  assign new_A9599_ = new_A9581_ | new_A9596_;
  assign new_A9600_ = ~new_A9574_ | ~new_A9575_;
  assign new_A9601_ = new_A9581_ | new_A9596_;
  assign new_A9602_ = ~new_A9581_ & ~new_A9603_;
  assign new_A9603_ = new_A9581_ & new_A9596_;
  assign new_A9604_ = new_B2055_;
  assign new_A9605_ = new_B2088_;
  assign new_A9606_ = new_B2121_;
  assign new_A9607_ = new_B2154_;
  assign new_A9608_ = new_B2187_;
  assign new_A9609_ = new_A9615_ & new_A9614_;
  assign new_A9610_ = new_A9617_ | new_A9616_;
  assign new_A9611_ = new_A9619_ | new_A9618_;
  assign new_A9612_ = new_A9614_ & new_A9620_;
  assign new_A9613_ = new_A9614_ & new_A9621_;
  assign new_A9614_ = new_A9604_ ^ new_A9605_;
  assign new_A9615_ = new_A9616_ ^ new_A9606_;
  assign new_A9616_ = new_A9624_ & new_A9623_;
  assign new_A9617_ = new_A9622_ & new_A9606_;
  assign new_A9618_ = new_A9627_ & new_A9626_;
  assign new_A9619_ = new_A9625_ & new_A9606_;
  assign new_A9620_ = new_A9628_ | new_A9605_;
  assign new_A9621_ = ~new_A9606_ ^ new_A9618_;
  assign new_A9622_ = ~new_A9631_ | ~new_A9632_;
  assign new_A9623_ = new_A9607_ ^ new_A9614_;
  assign new_A9624_ = new_A9633_ & new_A9626_;
  assign new_A9625_ = ~new_A9635_ | ~new_A9634_;
  assign new_A9626_ = new_A9607_ | new_A9608_;
  assign new_A9627_ = new_A9607_ | new_A9614_;
  assign new_A9628_ = new_A9606_ & new_A9618_;
  assign new_A9629_ = ~new_A9605_ | ~new_A9606_;
  assign new_A9630_ = new_A9614_ & new_A9629_;
  assign new_A9631_ = ~new_A9630_ & ~new_A9614_;
  assign new_A9632_ = new_A9614_ | new_A9629_;
  assign new_A9633_ = ~new_A9607_ | ~new_A9608_;
  assign new_A9634_ = new_A9614_ | new_A9629_;
  assign new_A9635_ = ~new_A9614_ & ~new_A9636_;
  assign new_A9636_ = new_A9614_ & new_A9629_;
  assign new_A9637_ = new_B2220_;
  assign new_A9638_ = new_B2253_;
  assign new_A9639_ = new_B2286_;
  assign new_A9640_ = new_B2319_;
  assign new_A9641_ = new_B2352_;
  assign new_A9642_ = new_A9648_ & new_A9647_;
  assign new_A9643_ = new_A9650_ | new_A9649_;
  assign new_A9644_ = new_A9652_ | new_A9651_;
  assign new_A9645_ = new_A9647_ & new_A9653_;
  assign new_A9646_ = new_A9647_ & new_A9654_;
  assign new_A9647_ = new_A9637_ ^ new_A9638_;
  assign new_A9648_ = new_A9649_ ^ new_A9639_;
  assign new_A9649_ = new_A9657_ & new_A9656_;
  assign new_A9650_ = new_A9655_ & new_A9639_;
  assign new_A9651_ = new_A9660_ & new_A9659_;
  assign new_A9652_ = new_A9658_ & new_A9639_;
  assign new_A9653_ = new_A9661_ | new_A9638_;
  assign new_A9654_ = ~new_A9639_ ^ new_A9651_;
  assign new_A9655_ = ~new_A9664_ | ~new_A9665_;
  assign new_A9656_ = new_A9640_ ^ new_A9647_;
  assign new_A9657_ = new_A9666_ & new_A9659_;
  assign new_A9658_ = ~new_A9668_ | ~new_A9667_;
  assign new_A9659_ = new_A9640_ | new_A9641_;
  assign new_A9660_ = new_A9640_ | new_A9647_;
  assign new_A9661_ = new_A9639_ & new_A9651_;
  assign new_A9662_ = ~new_A9638_ | ~new_A9639_;
  assign new_A9663_ = new_A9647_ & new_A9662_;
  assign new_A9664_ = ~new_A9663_ & ~new_A9647_;
  assign new_A9665_ = new_A9647_ | new_A9662_;
  assign new_A9666_ = ~new_A9640_ | ~new_A9641_;
  assign new_A9667_ = new_A9647_ | new_A9662_;
  assign new_A9668_ = ~new_A9647_ & ~new_A9669_;
  assign new_A9669_ = new_A9647_ & new_A9662_;
  assign new_A9670_ = new_B2385_;
  assign new_A9671_ = new_B2418_;
  assign new_A9672_ = new_B2451_;
  assign new_A9673_ = new_B2484_;
  assign new_A9674_ = new_B2517_;
  assign new_A9675_ = new_A9681_ & new_A9680_;
  assign new_A9676_ = new_A9683_ | new_A9682_;
  assign new_A9677_ = new_A9685_ | new_A9684_;
  assign new_A9678_ = new_A9680_ & new_A9686_;
  assign new_A9679_ = new_A9680_ & new_A9687_;
  assign new_A9680_ = new_A9670_ ^ new_A9671_;
  assign new_A9681_ = new_A9682_ ^ new_A9672_;
  assign new_A9682_ = new_A9690_ & new_A9689_;
  assign new_A9683_ = new_A9688_ & new_A9672_;
  assign new_A9684_ = new_A9693_ & new_A9692_;
  assign new_A9685_ = new_A9691_ & new_A9672_;
  assign new_A9686_ = new_A9694_ | new_A9671_;
  assign new_A9687_ = ~new_A9672_ ^ new_A9684_;
  assign new_A9688_ = ~new_A9697_ | ~new_A9698_;
  assign new_A9689_ = new_A9673_ ^ new_A9680_;
  assign new_A9690_ = new_A9699_ & new_A9692_;
  assign new_A9691_ = ~new_A9701_ | ~new_A9700_;
  assign new_A9692_ = new_A9673_ | new_A9674_;
  assign new_A9693_ = new_A9673_ | new_A9680_;
  assign new_A9694_ = new_A9672_ & new_A9684_;
  assign new_A9695_ = ~new_A9671_ | ~new_A9672_;
  assign new_A9696_ = new_A9680_ & new_A9695_;
  assign new_A9697_ = ~new_A9696_ & ~new_A9680_;
  assign new_A9698_ = new_A9680_ | new_A9695_;
  assign new_A9699_ = ~new_A9673_ | ~new_A9674_;
  assign new_A9700_ = new_A9680_ | new_A9695_;
  assign new_A9701_ = ~new_A9680_ & ~new_A9702_;
  assign new_A9702_ = new_A9680_ & new_A9695_;
  assign new_A9703_ = new_B2550_;
  assign new_A9704_ = new_B2583_;
  assign new_A9705_ = new_B2616_;
  assign new_A9706_ = new_B2649_;
  assign new_A9707_ = new_B2682_;
  assign new_A9708_ = new_A9714_ & new_A9713_;
  assign new_A9709_ = new_A9716_ | new_A9715_;
  assign new_A9710_ = new_A9718_ | new_A9717_;
  assign new_A9711_ = new_A9713_ & new_A9719_;
  assign new_A9712_ = new_A9713_ & new_A9720_;
  assign new_A9713_ = new_A9703_ ^ new_A9704_;
  assign new_A9714_ = new_A9715_ ^ new_A9705_;
  assign new_A9715_ = new_A9723_ & new_A9722_;
  assign new_A9716_ = new_A9721_ & new_A9705_;
  assign new_A9717_ = new_A9726_ & new_A9725_;
  assign new_A9718_ = new_A9724_ & new_A9705_;
  assign new_A9719_ = new_A9727_ | new_A9704_;
  assign new_A9720_ = ~new_A9705_ ^ new_A9717_;
  assign new_A9721_ = ~new_A9730_ | ~new_A9731_;
  assign new_A9722_ = new_A9706_ ^ new_A9713_;
  assign new_A9723_ = new_A9732_ & new_A9725_;
  assign new_A9724_ = ~new_A9734_ | ~new_A9733_;
  assign new_A9725_ = new_A9706_ | new_A9707_;
  assign new_A9726_ = new_A9706_ | new_A9713_;
  assign new_A9727_ = new_A9705_ & new_A9717_;
  assign new_A9728_ = ~new_A9704_ | ~new_A9705_;
  assign new_A9729_ = new_A9713_ & new_A9728_;
  assign new_A9730_ = ~new_A9729_ & ~new_A9713_;
  assign new_A9731_ = new_A9713_ | new_A9728_;
  assign new_A9732_ = ~new_A9706_ | ~new_A9707_;
  assign new_A9733_ = new_A9713_ | new_A9728_;
  assign new_A9734_ = ~new_A9713_ & ~new_A9735_;
  assign new_A9735_ = new_A9713_ & new_A9728_;
  assign new_A9736_ = new_B2715_;
  assign new_A9737_ = new_B2748_;
  assign new_A9738_ = new_B2781_;
  assign new_A9739_ = new_B2814_;
  assign new_A9740_ = new_B2847_;
  assign new_A9741_ = new_A9747_ & new_A9746_;
  assign new_A9742_ = new_A9749_ | new_A9748_;
  assign new_A9743_ = new_A9751_ | new_A9750_;
  assign new_A9744_ = new_A9746_ & new_A9752_;
  assign new_A9745_ = new_A9746_ & new_A9753_;
  assign new_A9746_ = new_A9736_ ^ new_A9737_;
  assign new_A9747_ = new_A9748_ ^ new_A9738_;
  assign new_A9748_ = new_A9756_ & new_A9755_;
  assign new_A9749_ = new_A9754_ & new_A9738_;
  assign new_A9750_ = new_A9759_ & new_A9758_;
  assign new_A9751_ = new_A9757_ & new_A9738_;
  assign new_A9752_ = new_A9760_ | new_A9737_;
  assign new_A9753_ = ~new_A9738_ ^ new_A9750_;
  assign new_A9754_ = ~new_A9763_ | ~new_A9764_;
  assign new_A9755_ = new_A9739_ ^ new_A9746_;
  assign new_A9756_ = new_A9765_ & new_A9758_;
  assign new_A9757_ = ~new_A9767_ | ~new_A9766_;
  assign new_A9758_ = new_A9739_ | new_A9740_;
  assign new_A9759_ = new_A9739_ | new_A9746_;
  assign new_A9760_ = new_A9738_ & new_A9750_;
  assign new_A9761_ = ~new_A9737_ | ~new_A9738_;
  assign new_A9762_ = new_A9746_ & new_A9761_;
  assign new_A9763_ = ~new_A9762_ & ~new_A9746_;
  assign new_A9764_ = new_A9746_ | new_A9761_;
  assign new_A9765_ = ~new_A9739_ | ~new_A9740_;
  assign new_A9766_ = new_A9746_ | new_A9761_;
  assign new_A9767_ = ~new_A9746_ & ~new_A9768_;
  assign new_A9768_ = new_A9746_ & new_A9761_;
  assign new_A9769_ = new_B2880_;
  assign new_A9770_ = new_B2913_;
  assign new_A9771_ = new_B2946_;
  assign new_A9772_ = new_B2979_;
  assign new_A9773_ = new_B3012_;
  assign new_A9774_ = new_A9780_ & new_A9779_;
  assign new_A9775_ = new_A9782_ | new_A9781_;
  assign new_A9776_ = new_A9784_ | new_A9783_;
  assign new_A9777_ = new_A9779_ & new_A9785_;
  assign new_A9778_ = new_A9779_ & new_A9786_;
  assign new_A9779_ = new_A9769_ ^ new_A9770_;
  assign new_A9780_ = new_A9781_ ^ new_A9771_;
  assign new_A9781_ = new_A9789_ & new_A9788_;
  assign new_A9782_ = new_A9787_ & new_A9771_;
  assign new_A9783_ = new_A9792_ & new_A9791_;
  assign new_A9784_ = new_A9790_ & new_A9771_;
  assign new_A9785_ = new_A9793_ | new_A9770_;
  assign new_A9786_ = ~new_A9771_ ^ new_A9783_;
  assign new_A9787_ = ~new_A9796_ | ~new_A9797_;
  assign new_A9788_ = new_A9772_ ^ new_A9779_;
  assign new_A9789_ = new_A9798_ & new_A9791_;
  assign new_A9790_ = ~new_A9800_ | ~new_A9799_;
  assign new_A9791_ = new_A9772_ | new_A9773_;
  assign new_A9792_ = new_A9772_ | new_A9779_;
  assign new_A9793_ = new_A9771_ & new_A9783_;
  assign new_A9794_ = ~new_A9770_ | ~new_A9771_;
  assign new_A9795_ = new_A9779_ & new_A9794_;
  assign new_A9796_ = ~new_A9795_ & ~new_A9779_;
  assign new_A9797_ = new_A9779_ | new_A9794_;
  assign new_A9798_ = ~new_A9772_ | ~new_A9773_;
  assign new_A9799_ = new_A9779_ | new_A9794_;
  assign new_A9800_ = ~new_A9779_ & ~new_A9801_;
  assign new_A9801_ = new_A9779_ & new_A9794_;
  assign new_A9802_ = new_B3045_;
  assign new_A9803_ = new_B3078_;
  assign new_A9804_ = new_B3111_;
  assign new_A9805_ = new_B3144_;
  assign new_A9806_ = new_B3177_;
  assign new_A9807_ = new_A9813_ & new_A9812_;
  assign new_A9808_ = new_A9815_ | new_A9814_;
  assign new_A9809_ = new_A9817_ | new_A9816_;
  assign new_A9810_ = new_A9812_ & new_A9818_;
  assign new_A9811_ = new_A9812_ & new_A9819_;
  assign new_A9812_ = new_A9802_ ^ new_A9803_;
  assign new_A9813_ = new_A9814_ ^ new_A9804_;
  assign new_A9814_ = new_A9822_ & new_A9821_;
  assign new_A9815_ = new_A9820_ & new_A9804_;
  assign new_A9816_ = new_A9825_ & new_A9824_;
  assign new_A9817_ = new_A9823_ & new_A9804_;
  assign new_A9818_ = new_A9826_ | new_A9803_;
  assign new_A9819_ = ~new_A9804_ ^ new_A9816_;
  assign new_A9820_ = ~new_A9829_ | ~new_A9830_;
  assign new_A9821_ = new_A9805_ ^ new_A9812_;
  assign new_A9822_ = new_A9831_ & new_A9824_;
  assign new_A9823_ = ~new_A9833_ | ~new_A9832_;
  assign new_A9824_ = new_A9805_ | new_A9806_;
  assign new_A9825_ = new_A9805_ | new_A9812_;
  assign new_A9826_ = new_A9804_ & new_A9816_;
  assign new_A9827_ = ~new_A9803_ | ~new_A9804_;
  assign new_A9828_ = new_A9812_ & new_A9827_;
  assign new_A9829_ = ~new_A9828_ & ~new_A9812_;
  assign new_A9830_ = new_A9812_ | new_A9827_;
  assign new_A9831_ = ~new_A9805_ | ~new_A9806_;
  assign new_A9832_ = new_A9812_ | new_A9827_;
  assign new_A9833_ = ~new_A9812_ & ~new_A9834_;
  assign new_A9834_ = new_A9812_ & new_A9827_;
  assign new_A9835_ = new_B3210_;
  assign new_A9836_ = new_B3243_;
  assign new_A9837_ = new_B3276_;
  assign new_A9838_ = new_B3309_;
  assign new_A9839_ = new_B3342_;
  assign new_A9840_ = new_A9846_ & new_A9845_;
  assign new_A9841_ = new_A9848_ | new_A9847_;
  assign new_A9842_ = new_A9850_ | new_A9849_;
  assign new_A9843_ = new_A9845_ & new_A9851_;
  assign new_A9844_ = new_A9845_ & new_A9852_;
  assign new_A9845_ = new_A9835_ ^ new_A9836_;
  assign new_A9846_ = new_A9847_ ^ new_A9837_;
  assign new_A9847_ = new_A9855_ & new_A9854_;
  assign new_A9848_ = new_A9853_ & new_A9837_;
  assign new_A9849_ = new_A9858_ & new_A9857_;
  assign new_A9850_ = new_A9856_ & new_A9837_;
  assign new_A9851_ = new_A9859_ | new_A9836_;
  assign new_A9852_ = ~new_A9837_ ^ new_A9849_;
  assign new_A9853_ = ~new_A9862_ | ~new_A9863_;
  assign new_A9854_ = new_A9838_ ^ new_A9845_;
  assign new_A9855_ = new_A9864_ & new_A9857_;
  assign new_A9856_ = ~new_A9866_ | ~new_A9865_;
  assign new_A9857_ = new_A9838_ | new_A9839_;
  assign new_A9858_ = new_A9838_ | new_A9845_;
  assign new_A9859_ = new_A9837_ & new_A9849_;
  assign new_A9860_ = ~new_A9836_ | ~new_A9837_;
  assign new_A9861_ = new_A9845_ & new_A9860_;
  assign new_A9862_ = ~new_A9861_ & ~new_A9845_;
  assign new_A9863_ = new_A9845_ | new_A9860_;
  assign new_A9864_ = ~new_A9838_ | ~new_A9839_;
  assign new_A9865_ = new_A9845_ | new_A9860_;
  assign new_A9866_ = ~new_A9845_ & ~new_A9867_;
  assign new_A9867_ = new_A9845_ & new_A9860_;
  assign new_A9868_ = new_B3375_;
  assign new_A9869_ = new_B3408_;
  assign new_A9870_ = new_B3441_;
  assign new_A9871_ = new_B3474_;
  assign new_A9872_ = new_B3507_;
  assign new_A9873_ = new_A9879_ & new_A9878_;
  assign new_A9874_ = new_A9881_ | new_A9880_;
  assign new_A9875_ = new_A9883_ | new_A9882_;
  assign new_A9876_ = new_A9878_ & new_A9884_;
  assign new_A9877_ = new_A9878_ & new_A9885_;
  assign new_A9878_ = new_A9868_ ^ new_A9869_;
  assign new_A9879_ = new_A9880_ ^ new_A9870_;
  assign new_A9880_ = new_A9888_ & new_A9887_;
  assign new_A9881_ = new_A9886_ & new_A9870_;
  assign new_A9882_ = new_A9891_ & new_A9890_;
  assign new_A9883_ = new_A9889_ & new_A9870_;
  assign new_A9884_ = new_A9892_ | new_A9869_;
  assign new_A9885_ = ~new_A9870_ ^ new_A9882_;
  assign new_A9886_ = ~new_A9895_ | ~new_A9896_;
  assign new_A9887_ = new_A9871_ ^ new_A9878_;
  assign new_A9888_ = new_A9897_ & new_A9890_;
  assign new_A9889_ = ~new_A9899_ | ~new_A9898_;
  assign new_A9890_ = new_A9871_ | new_A9872_;
  assign new_A9891_ = new_A9871_ | new_A9878_;
  assign new_A9892_ = new_A9870_ & new_A9882_;
  assign new_A9893_ = ~new_A9869_ | ~new_A9870_;
  assign new_A9894_ = new_A9878_ & new_A9893_;
  assign new_A9895_ = ~new_A9894_ & ~new_A9878_;
  assign new_A9896_ = new_A9878_ | new_A9893_;
  assign new_A9897_ = ~new_A9871_ | ~new_A9872_;
  assign new_A9898_ = new_A9878_ | new_A9893_;
  assign new_A9899_ = ~new_A9878_ & ~new_A9900_;
  assign new_A9900_ = new_A9878_ & new_A9893_;
  assign new_A9901_ = new_B3540_;
  assign new_A9902_ = new_B3573_;
  assign new_A9903_ = new_B3606_;
  assign new_A9904_ = new_B3639_;
  assign new_A9905_ = new_B3672_;
  assign new_A9906_ = new_A9912_ & new_A9911_;
  assign new_A9907_ = new_A9914_ | new_A9913_;
  assign new_A9908_ = new_A9916_ | new_A9915_;
  assign new_A9909_ = new_A9911_ & new_A9917_;
  assign new_A9910_ = new_A9911_ & new_A9918_;
  assign new_A9911_ = new_A9901_ ^ new_A9902_;
  assign new_A9912_ = new_A9913_ ^ new_A9903_;
  assign new_A9913_ = new_A9921_ & new_A9920_;
  assign new_A9914_ = new_A9919_ & new_A9903_;
  assign new_A9915_ = new_A9924_ & new_A9923_;
  assign new_A9916_ = new_A9922_ & new_A9903_;
  assign new_A9917_ = new_A9925_ | new_A9902_;
  assign new_A9918_ = ~new_A9903_ ^ new_A9915_;
  assign new_A9919_ = ~new_A9928_ | ~new_A9929_;
  assign new_A9920_ = new_A9904_ ^ new_A9911_;
  assign new_A9921_ = new_A9930_ & new_A9923_;
  assign new_A9922_ = ~new_A9932_ | ~new_A9931_;
  assign new_A9923_ = new_A9904_ | new_A9905_;
  assign new_A9924_ = new_A9904_ | new_A9911_;
  assign new_A9925_ = new_A9903_ & new_A9915_;
  assign new_A9926_ = ~new_A9902_ | ~new_A9903_;
  assign new_A9927_ = new_A9911_ & new_A9926_;
  assign new_A9928_ = ~new_A9927_ & ~new_A9911_;
  assign new_A9929_ = new_A9911_ | new_A9926_;
  assign new_A9930_ = ~new_A9904_ | ~new_A9905_;
  assign new_A9931_ = new_A9911_ | new_A9926_;
  assign new_A9932_ = ~new_A9911_ & ~new_A9933_;
  assign new_A9933_ = new_A9911_ & new_A9926_;
  assign new_A9934_ = new_B3705_;
  assign new_A9935_ = new_B3738_;
  assign new_A9936_ = new_B3771_;
  assign new_A9937_ = new_B3804_;
  assign new_A9938_ = new_B3837_;
  assign new_A9939_ = new_A9945_ & new_A9944_;
  assign new_A9940_ = new_A9947_ | new_A9946_;
  assign new_A9941_ = new_A9949_ | new_A9948_;
  assign new_A9942_ = new_A9944_ & new_A9950_;
  assign new_A9943_ = new_A9944_ & new_A9951_;
  assign new_A9944_ = new_A9934_ ^ new_A9935_;
  assign new_A9945_ = new_A9946_ ^ new_A9936_;
  assign new_A9946_ = new_A9954_ & new_A9953_;
  assign new_A9947_ = new_A9952_ & new_A9936_;
  assign new_A9948_ = new_A9957_ & new_A9956_;
  assign new_A9949_ = new_A9955_ & new_A9936_;
  assign new_A9950_ = new_A9958_ | new_A9935_;
  assign new_A9951_ = ~new_A9936_ ^ new_A9948_;
  assign new_A9952_ = ~new_A9961_ | ~new_A9962_;
  assign new_A9953_ = new_A9937_ ^ new_A9944_;
  assign new_A9954_ = new_A9963_ & new_A9956_;
  assign new_A9955_ = ~new_A9965_ | ~new_A9964_;
  assign new_A9956_ = new_A9937_ | new_A9938_;
  assign new_A9957_ = new_A9937_ | new_A9944_;
  assign new_A9958_ = new_A9936_ & new_A9948_;
  assign new_A9959_ = ~new_A9935_ | ~new_A9936_;
  assign new_A9960_ = new_A9944_ & new_A9959_;
  assign new_A9961_ = ~new_A9960_ & ~new_A9944_;
  assign new_A9962_ = new_A9944_ | new_A9959_;
  assign new_A9963_ = ~new_A9937_ | ~new_A9938_;
  assign new_A9964_ = new_A9944_ | new_A9959_;
  assign new_A9965_ = ~new_A9944_ & ~new_A9966_;
  assign new_A9966_ = new_A9944_ & new_A9959_;
  assign new_A9967_ = new_B3870_;
  assign new_A9968_ = new_B3903_;
  assign new_A9969_ = new_B3936_;
  assign new_A9970_ = new_B3969_;
  assign new_A9971_ = new_B4002_;
  assign new_A9972_ = new_A9978_ & new_A9977_;
  assign new_A9973_ = new_A9980_ | new_A9979_;
  assign new_A9974_ = new_A9982_ | new_A9981_;
  assign new_A9975_ = new_A9977_ & new_A9983_;
  assign new_A9976_ = new_A9977_ & new_A9984_;
  assign new_A9977_ = new_A9967_ ^ new_A9968_;
  assign new_A9978_ = new_A9979_ ^ new_A9969_;
  assign new_A9979_ = new_A9987_ & new_A9986_;
  assign new_A9980_ = new_A9985_ & new_A9969_;
  assign new_A9981_ = new_A9990_ & new_A9989_;
  assign new_A9982_ = new_A9988_ & new_A9969_;
  assign new_A9983_ = new_A9991_ | new_A9968_;
  assign new_A9984_ = ~new_A9969_ ^ new_A9981_;
  assign new_A9985_ = ~new_A9994_ | ~new_A9995_;
  assign new_A9986_ = new_A9970_ ^ new_A9977_;
  assign new_A9987_ = new_A9996_ & new_A9989_;
  assign new_A9988_ = ~new_A9998_ | ~new_A9997_;
  assign new_A9989_ = new_A9970_ | new_A9971_;
  assign new_A9990_ = new_A9970_ | new_A9977_;
  assign new_A9991_ = new_A9969_ & new_A9981_;
  assign new_A9992_ = ~new_A9968_ | ~new_A9969_;
  assign new_A9993_ = new_A9977_ & new_A9992_;
  assign new_A9994_ = ~new_A9993_ & ~new_A9977_;
  assign new_A9995_ = new_A9977_ | new_A9992_;
  assign new_A9996_ = ~new_A9970_ | ~new_A9971_;
  assign new_A9997_ = new_A9977_ | new_A9992_;
  assign new_A9998_ = ~new_A9977_ & ~new_A9999_;
  assign new_A9999_ = new_A9977_ & new_A9992_;
  assign new_B1_ = new_B4035_;
  assign new_B2_ = new_B4068_;
  assign new_B3_ = new_B4101_;
  assign new_B4_ = new_B4134_;
  assign new_B5_ = new_B4167_;
  assign new_B6_ = new_B12_ & new_B11_;
  assign new_B7_ = new_B14_ | new_B13_;
  assign new_B8_ = new_B16_ | new_B15_;
  assign new_B9_ = new_B11_ & new_B17_;
  assign new_B10_ = new_B11_ & new_B18_;
  assign new_B11_ = new_B1_ ^ new_B2_;
  assign new_B12_ = new_B13_ ^ new_B3_;
  assign new_B13_ = new_B21_ & new_B20_;
  assign new_B14_ = new_B19_ & new_B3_;
  assign new_B15_ = new_B24_ & new_B23_;
  assign new_B16_ = new_B22_ & new_B3_;
  assign new_B17_ = new_B25_ | new_B2_;
  assign new_B18_ = ~new_B3_ ^ new_B15_;
  assign new_B19_ = ~new_B28_ | ~new_B29_;
  assign new_B20_ = new_B4_ ^ new_B11_;
  assign new_B21_ = new_B30_ & new_B23_;
  assign new_B22_ = ~new_B32_ | ~new_B31_;
  assign new_B23_ = new_B4_ | new_B5_;
  assign new_B24_ = new_B4_ | new_B11_;
  assign new_B25_ = new_B3_ & new_B15_;
  assign new_B26_ = ~new_B2_ | ~new_B3_;
  assign new_B27_ = new_B11_ & new_B26_;
  assign new_B28_ = ~new_B27_ & ~new_B11_;
  assign new_B29_ = new_B11_ | new_B26_;
  assign new_B30_ = ~new_B4_ | ~new_B5_;
  assign new_B31_ = new_B11_ | new_B26_;
  assign new_B32_ = ~new_B11_ & ~new_B33_;
  assign new_B33_ = new_B11_ & new_B26_;
  assign new_B34_ = new_B4200_;
  assign new_B35_ = new_B4233_;
  assign new_B36_ = new_B4266_;
  assign new_B37_ = new_B4299_;
  assign new_B38_ = new_B4332_;
  assign new_B39_ = new_B45_ & new_B44_;
  assign new_B40_ = new_B47_ | new_B46_;
  assign new_B41_ = new_B49_ | new_B48_;
  assign new_B42_ = new_B44_ & new_B50_;
  assign new_B43_ = new_B44_ & new_B51_;
  assign new_B44_ = new_B34_ ^ new_B35_;
  assign new_B45_ = new_B46_ ^ new_B36_;
  assign new_B46_ = new_B54_ & new_B53_;
  assign new_B47_ = new_B52_ & new_B36_;
  assign new_B48_ = new_B57_ & new_B56_;
  assign new_B49_ = new_B55_ & new_B36_;
  assign new_B50_ = new_B58_ | new_B35_;
  assign new_B51_ = ~new_B36_ ^ new_B48_;
  assign new_B52_ = ~new_B61_ | ~new_B62_;
  assign new_B53_ = new_B37_ ^ new_B44_;
  assign new_B54_ = new_B63_ & new_B56_;
  assign new_B55_ = ~new_B65_ | ~new_B64_;
  assign new_B56_ = new_B37_ | new_B38_;
  assign new_B57_ = new_B37_ | new_B44_;
  assign new_B58_ = new_B36_ & new_B48_;
  assign new_B59_ = ~new_B35_ | ~new_B36_;
  assign new_B60_ = new_B44_ & new_B59_;
  assign new_B61_ = ~new_B60_ & ~new_B44_;
  assign new_B62_ = new_B44_ | new_B59_;
  assign new_B63_ = ~new_B37_ | ~new_B38_;
  assign new_B64_ = new_B44_ | new_B59_;
  assign new_B65_ = ~new_B44_ & ~new_B66_;
  assign new_B66_ = new_B44_ & new_B59_;
  assign new_B67_ = new_B4365_;
  assign new_B68_ = new_B4398_;
  assign new_B69_ = new_B4431_;
  assign new_B70_ = new_B4464_;
  assign new_B71_ = new_B4497_;
  assign new_B72_ = new_B78_ & new_B77_;
  assign new_B73_ = new_B80_ | new_B79_;
  assign new_B74_ = new_B82_ | new_B81_;
  assign new_B75_ = new_B77_ & new_B83_;
  assign new_B76_ = new_B77_ & new_B84_;
  assign new_B77_ = new_B67_ ^ new_B68_;
  assign new_B78_ = new_B79_ ^ new_B69_;
  assign new_B79_ = new_B87_ & new_B86_;
  assign new_B80_ = new_B85_ & new_B69_;
  assign new_B81_ = new_B90_ & new_B89_;
  assign new_B82_ = new_B88_ & new_B69_;
  assign new_B83_ = new_B91_ | new_B68_;
  assign new_B84_ = ~new_B69_ ^ new_B81_;
  assign new_B85_ = ~new_B94_ | ~new_B95_;
  assign new_B86_ = new_B70_ ^ new_B77_;
  assign new_B87_ = new_B96_ & new_B89_;
  assign new_B88_ = ~new_B98_ | ~new_B97_;
  assign new_B89_ = new_B70_ | new_B71_;
  assign new_B90_ = new_B70_ | new_B77_;
  assign new_B91_ = new_B69_ & new_B81_;
  assign new_B92_ = ~new_B68_ | ~new_B69_;
  assign new_B93_ = new_B77_ & new_B92_;
  assign new_B94_ = ~new_B93_ & ~new_B77_;
  assign new_B95_ = new_B77_ | new_B92_;
  assign new_B96_ = ~new_B70_ | ~new_B71_;
  assign new_B97_ = new_B77_ | new_B92_;
  assign new_B98_ = ~new_B77_ & ~new_B99_;
  assign new_B99_ = new_B77_ & new_B92_;
  assign new_B100_ = new_B4530_;
  assign new_B101_ = new_B4563_;
  assign new_B102_ = new_B4596_;
  assign new_B103_ = new_B4629_;
  assign new_B104_ = new_B4662_;
  assign new_B105_ = new_B111_ & new_B110_;
  assign new_B106_ = new_B113_ | new_B112_;
  assign new_B107_ = new_B115_ | new_B114_;
  assign new_B108_ = new_B110_ & new_B116_;
  assign new_B109_ = new_B110_ & new_B117_;
  assign new_B110_ = new_B100_ ^ new_B101_;
  assign new_B111_ = new_B112_ ^ new_B102_;
  assign new_B112_ = new_B120_ & new_B119_;
  assign new_B113_ = new_B118_ & new_B102_;
  assign new_B114_ = new_B123_ & new_B122_;
  assign new_B115_ = new_B121_ & new_B102_;
  assign new_B116_ = new_B124_ | new_B101_;
  assign new_B117_ = ~new_B102_ ^ new_B114_;
  assign new_B118_ = ~new_B127_ | ~new_B128_;
  assign new_B119_ = new_B103_ ^ new_B110_;
  assign new_B120_ = new_B129_ & new_B122_;
  assign new_B121_ = ~new_B131_ | ~new_B130_;
  assign new_B122_ = new_B103_ | new_B104_;
  assign new_B123_ = new_B103_ | new_B110_;
  assign new_B124_ = new_B102_ & new_B114_;
  assign new_B125_ = ~new_B101_ | ~new_B102_;
  assign new_B126_ = new_B110_ & new_B125_;
  assign new_B127_ = ~new_B126_ & ~new_B110_;
  assign new_B128_ = new_B110_ | new_B125_;
  assign new_B129_ = ~new_B103_ | ~new_B104_;
  assign new_B130_ = new_B110_ | new_B125_;
  assign new_B131_ = ~new_B110_ & ~new_B132_;
  assign new_B132_ = new_B110_ & new_B125_;
  assign new_B133_ = new_B4695_;
  assign new_B134_ = new_B4728_;
  assign new_B135_ = new_B4761_;
  assign new_B136_ = new_B4794_;
  assign new_B137_ = new_B4827_;
  assign new_B138_ = new_B144_ & new_B143_;
  assign new_B139_ = new_B146_ | new_B145_;
  assign new_B140_ = new_B148_ | new_B147_;
  assign new_B141_ = new_B143_ & new_B149_;
  assign new_B142_ = new_B143_ & new_B150_;
  assign new_B143_ = new_B133_ ^ new_B134_;
  assign new_B144_ = new_B145_ ^ new_B135_;
  assign new_B145_ = new_B153_ & new_B152_;
  assign new_B146_ = new_B151_ & new_B135_;
  assign new_B147_ = new_B156_ & new_B155_;
  assign new_B148_ = new_B154_ & new_B135_;
  assign new_B149_ = new_B157_ | new_B134_;
  assign new_B150_ = ~new_B135_ ^ new_B147_;
  assign new_B151_ = ~new_B160_ | ~new_B161_;
  assign new_B152_ = new_B136_ ^ new_B143_;
  assign new_B153_ = new_B162_ & new_B155_;
  assign new_B154_ = ~new_B164_ | ~new_B163_;
  assign new_B155_ = new_B136_ | new_B137_;
  assign new_B156_ = new_B136_ | new_B143_;
  assign new_B157_ = new_B135_ & new_B147_;
  assign new_B158_ = ~new_B134_ | ~new_B135_;
  assign new_B159_ = new_B143_ & new_B158_;
  assign new_B160_ = ~new_B159_ & ~new_B143_;
  assign new_B161_ = new_B143_ | new_B158_;
  assign new_B162_ = ~new_B136_ | ~new_B137_;
  assign new_B163_ = new_B143_ | new_B158_;
  assign new_B164_ = ~new_B143_ & ~new_B165_;
  assign new_B165_ = new_B143_ & new_B158_;
  assign new_B166_ = new_B4860_;
  assign new_B167_ = new_B4893_;
  assign new_B168_ = new_B4926_;
  assign new_B169_ = new_B4959_;
  assign new_B170_ = new_B4992_;
  assign new_B171_ = new_B177_ & new_B176_;
  assign new_B172_ = new_B179_ | new_B178_;
  assign new_B173_ = new_B181_ | new_B180_;
  assign new_B174_ = new_B176_ & new_B182_;
  assign new_B175_ = new_B176_ & new_B183_;
  assign new_B176_ = new_B166_ ^ new_B167_;
  assign new_B177_ = new_B178_ ^ new_B168_;
  assign new_B178_ = new_B186_ & new_B185_;
  assign new_B179_ = new_B184_ & new_B168_;
  assign new_B180_ = new_B189_ & new_B188_;
  assign new_B181_ = new_B187_ & new_B168_;
  assign new_B182_ = new_B190_ | new_B167_;
  assign new_B183_ = ~new_B168_ ^ new_B180_;
  assign new_B184_ = ~new_B193_ | ~new_B194_;
  assign new_B185_ = new_B169_ ^ new_B176_;
  assign new_B186_ = new_B195_ & new_B188_;
  assign new_B187_ = ~new_B197_ | ~new_B196_;
  assign new_B188_ = new_B169_ | new_B170_;
  assign new_B189_ = new_B169_ | new_B176_;
  assign new_B190_ = new_B168_ & new_B180_;
  assign new_B191_ = ~new_B167_ | ~new_B168_;
  assign new_B192_ = new_B176_ & new_B191_;
  assign new_B193_ = ~new_B192_ & ~new_B176_;
  assign new_B194_ = new_B176_ | new_B191_;
  assign new_B195_ = ~new_B169_ | ~new_B170_;
  assign new_B196_ = new_B176_ | new_B191_;
  assign new_B197_ = ~new_B176_ & ~new_B198_;
  assign new_B198_ = new_B176_ & new_B191_;
  assign new_B199_ = new_B5025_;
  assign new_B200_ = new_B5058_;
  assign new_B201_ = new_B5091_;
  assign new_B202_ = new_B5124_;
  assign new_B203_ = new_B5157_;
  assign new_B204_ = new_B210_ & new_B209_;
  assign new_B205_ = new_B212_ | new_B211_;
  assign new_B206_ = new_B214_ | new_B213_;
  assign new_B207_ = new_B209_ & new_B215_;
  assign new_B208_ = new_B209_ & new_B216_;
  assign new_B209_ = new_B199_ ^ new_B200_;
  assign new_B210_ = new_B211_ ^ new_B201_;
  assign new_B211_ = new_B219_ & new_B218_;
  assign new_B212_ = new_B217_ & new_B201_;
  assign new_B213_ = new_B222_ & new_B221_;
  assign new_B214_ = new_B220_ & new_B201_;
  assign new_B215_ = new_B223_ | new_B200_;
  assign new_B216_ = ~new_B201_ ^ new_B213_;
  assign new_B217_ = ~new_B226_ | ~new_B227_;
  assign new_B218_ = new_B202_ ^ new_B209_;
  assign new_B219_ = new_B228_ & new_B221_;
  assign new_B220_ = ~new_B230_ | ~new_B229_;
  assign new_B221_ = new_B202_ | new_B203_;
  assign new_B222_ = new_B202_ | new_B209_;
  assign new_B223_ = new_B201_ & new_B213_;
  assign new_B224_ = ~new_B200_ | ~new_B201_;
  assign new_B225_ = new_B209_ & new_B224_;
  assign new_B226_ = ~new_B225_ & ~new_B209_;
  assign new_B227_ = new_B209_ | new_B224_;
  assign new_B228_ = ~new_B202_ | ~new_B203_;
  assign new_B229_ = new_B209_ | new_B224_;
  assign new_B230_ = ~new_B209_ & ~new_B231_;
  assign new_B231_ = new_B209_ & new_B224_;
  assign new_B232_ = new_B1062_;
  assign new_B233_ = new_B1099_;
  assign new_B234_ = new_B1132_;
  assign new_B235_ = new_B1165_;
  assign new_B236_ = new_B1198_;
  assign new_B237_ = new_B243_ & new_B242_;
  assign new_B238_ = new_B245_ | new_B244_;
  assign new_B239_ = new_B247_ | new_B246_;
  assign new_B240_ = new_B242_ & new_B248_;
  assign new_B241_ = new_B242_ & new_B249_;
  assign new_B242_ = new_B232_ ^ new_B233_;
  assign new_B243_ = new_B244_ ^ new_B234_;
  assign new_B244_ = new_B252_ & new_B251_;
  assign new_B245_ = new_B250_ & new_B234_;
  assign new_B246_ = new_B255_ & new_B254_;
  assign new_B247_ = new_B253_ & new_B234_;
  assign new_B248_ = new_B256_ | new_B233_;
  assign new_B249_ = ~new_B234_ ^ new_B246_;
  assign new_B250_ = ~new_B259_ | ~new_B260_;
  assign new_B251_ = new_B235_ ^ new_B242_;
  assign new_B252_ = new_B261_ & new_B254_;
  assign new_B253_ = ~new_B263_ | ~new_B262_;
  assign new_B254_ = new_B235_ | new_B236_;
  assign new_B255_ = new_B235_ | new_B242_;
  assign new_B256_ = new_B234_ & new_B246_;
  assign new_B257_ = ~new_B233_ | ~new_B234_;
  assign new_B258_ = new_B242_ & new_B257_;
  assign new_B259_ = ~new_B258_ & ~new_B242_;
  assign new_B260_ = new_B242_ | new_B257_;
  assign new_B261_ = ~new_B235_ | ~new_B236_;
  assign new_B262_ = new_B242_ | new_B257_;
  assign new_B263_ = ~new_B242_ & ~new_B264_;
  assign new_B264_ = new_B242_ & new_B257_;
  assign new_B265_ = new_B1231_;
  assign new_B266_ = new_B1264_;
  assign new_B267_ = new_B1297_;
  assign new_B268_ = new_B1330_;
  assign new_B269_ = new_B1363_;
  assign new_B270_ = new_B276_ & new_B275_;
  assign new_B271_ = new_B278_ | new_B277_;
  assign new_B272_ = new_B280_ | new_B279_;
  assign new_B273_ = new_B275_ & new_B281_;
  assign new_B274_ = new_B275_ & new_B282_;
  assign new_B275_ = new_B265_ ^ new_B266_;
  assign new_B276_ = new_B277_ ^ new_B267_;
  assign new_B277_ = new_B285_ & new_B284_;
  assign new_B278_ = new_B283_ & new_B267_;
  assign new_B279_ = new_B288_ & new_B287_;
  assign new_B280_ = new_B286_ & new_B267_;
  assign new_B281_ = new_B289_ | new_B266_;
  assign new_B282_ = ~new_B267_ ^ new_B279_;
  assign new_B283_ = ~new_B292_ | ~new_B293_;
  assign new_B284_ = new_B268_ ^ new_B275_;
  assign new_B285_ = new_B294_ & new_B287_;
  assign new_B286_ = ~new_B296_ | ~new_B295_;
  assign new_B287_ = new_B268_ | new_B269_;
  assign new_B288_ = new_B268_ | new_B275_;
  assign new_B289_ = new_B267_ & new_B279_;
  assign new_B290_ = ~new_B266_ | ~new_B267_;
  assign new_B291_ = new_B275_ & new_B290_;
  assign new_B292_ = ~new_B291_ & ~new_B275_;
  assign new_B293_ = new_B275_ | new_B290_;
  assign new_B294_ = ~new_B268_ | ~new_B269_;
  assign new_B295_ = new_B275_ | new_B290_;
  assign new_B296_ = ~new_B275_ & ~new_B297_;
  assign new_B297_ = new_B275_ & new_B290_;
  assign new_B298_ = new_B1396_;
  assign new_B299_ = new_B1429_;
  assign new_B300_ = new_B1462_;
  assign new_B301_ = new_B1495_;
  assign new_B302_ = new_B1528_;
  assign new_B303_ = new_B309_ & new_B308_;
  assign new_B304_ = new_B311_ | new_B310_;
  assign new_B305_ = new_B313_ | new_B312_;
  assign new_B306_ = new_B308_ & new_B314_;
  assign new_B307_ = new_B308_ & new_B315_;
  assign new_B308_ = new_B298_ ^ new_B299_;
  assign new_B309_ = new_B310_ ^ new_B300_;
  assign new_B310_ = new_B318_ & new_B317_;
  assign new_B311_ = new_B316_ & new_B300_;
  assign new_B312_ = new_B321_ & new_B320_;
  assign new_B313_ = new_B319_ & new_B300_;
  assign new_B314_ = new_B322_ | new_B299_;
  assign new_B315_ = ~new_B300_ ^ new_B312_;
  assign new_B316_ = ~new_B325_ | ~new_B326_;
  assign new_B317_ = new_B301_ ^ new_B308_;
  assign new_B318_ = new_B327_ & new_B320_;
  assign new_B319_ = ~new_B329_ | ~new_B328_;
  assign new_B320_ = new_B301_ | new_B302_;
  assign new_B321_ = new_B301_ | new_B308_;
  assign new_B322_ = new_B300_ & new_B312_;
  assign new_B323_ = ~new_B299_ | ~new_B300_;
  assign new_B324_ = new_B308_ & new_B323_;
  assign new_B325_ = ~new_B324_ & ~new_B308_;
  assign new_B326_ = new_B308_ | new_B323_;
  assign new_B327_ = ~new_B301_ | ~new_B302_;
  assign new_B328_ = new_B308_ | new_B323_;
  assign new_B329_ = ~new_B308_ & ~new_B330_;
  assign new_B330_ = new_B308_ & new_B323_;
  assign new_B331_ = new_B1561_;
  assign new_B332_ = new_B1594_;
  assign new_B333_ = new_B1627_;
  assign new_B334_ = new_B1660_;
  assign new_B335_ = new_B1693_;
  assign new_B336_ = new_B342_ & new_B341_;
  assign new_B337_ = new_B344_ | new_B343_;
  assign new_B338_ = new_B346_ | new_B345_;
  assign new_B339_ = new_B341_ & new_B347_;
  assign new_B340_ = new_B341_ & new_B348_;
  assign new_B341_ = new_B331_ ^ new_B332_;
  assign new_B342_ = new_B343_ ^ new_B333_;
  assign new_B343_ = new_B351_ & new_B350_;
  assign new_B344_ = new_B349_ & new_B333_;
  assign new_B345_ = new_B354_ & new_B353_;
  assign new_B346_ = new_B352_ & new_B333_;
  assign new_B347_ = new_B355_ | new_B332_;
  assign new_B348_ = ~new_B333_ ^ new_B345_;
  assign new_B349_ = ~new_B358_ | ~new_B359_;
  assign new_B350_ = new_B334_ ^ new_B341_;
  assign new_B351_ = new_B360_ & new_B353_;
  assign new_B352_ = ~new_B362_ | ~new_B361_;
  assign new_B353_ = new_B334_ | new_B335_;
  assign new_B354_ = new_B334_ | new_B341_;
  assign new_B355_ = new_B333_ & new_B345_;
  assign new_B356_ = ~new_B332_ | ~new_B333_;
  assign new_B357_ = new_B341_ & new_B356_;
  assign new_B358_ = ~new_B357_ & ~new_B341_;
  assign new_B359_ = new_B341_ | new_B356_;
  assign new_B360_ = ~new_B334_ | ~new_B335_;
  assign new_B361_ = new_B341_ | new_B356_;
  assign new_B362_ = ~new_B341_ & ~new_B363_;
  assign new_B363_ = new_B341_ & new_B356_;
  assign new_B364_ = new_B1726_;
  assign new_B365_ = new_B1759_;
  assign new_B366_ = new_B1792_;
  assign new_B367_ = new_B1825_;
  assign new_B368_ = new_B1858_;
  assign new_B369_ = new_B375_ & new_B374_;
  assign new_B370_ = new_B377_ | new_B376_;
  assign new_B371_ = new_B379_ | new_B378_;
  assign new_B372_ = new_B374_ & new_B380_;
  assign new_B373_ = new_B374_ & new_B381_;
  assign new_B374_ = new_B364_ ^ new_B365_;
  assign new_B375_ = new_B376_ ^ new_B366_;
  assign new_B376_ = new_B384_ & new_B383_;
  assign new_B377_ = new_B382_ & new_B366_;
  assign new_B378_ = new_B387_ & new_B386_;
  assign new_B379_ = new_B385_ & new_B366_;
  assign new_B380_ = new_B388_ | new_B365_;
  assign new_B381_ = ~new_B366_ ^ new_B378_;
  assign new_B382_ = ~new_B391_ | ~new_B392_;
  assign new_B383_ = new_B367_ ^ new_B374_;
  assign new_B384_ = new_B393_ & new_B386_;
  assign new_B385_ = ~new_B395_ | ~new_B394_;
  assign new_B386_ = new_B367_ | new_B368_;
  assign new_B387_ = new_B367_ | new_B374_;
  assign new_B388_ = new_B366_ & new_B378_;
  assign new_B389_ = ~new_B365_ | ~new_B366_;
  assign new_B390_ = new_B374_ & new_B389_;
  assign new_B391_ = ~new_B390_ & ~new_B374_;
  assign new_B392_ = new_B374_ | new_B389_;
  assign new_B393_ = ~new_B367_ | ~new_B368_;
  assign new_B394_ = new_B374_ | new_B389_;
  assign new_B395_ = ~new_B374_ & ~new_B396_;
  assign new_B396_ = new_B374_ & new_B389_;
  assign new_B397_ = new_B1891_;
  assign new_B398_ = new_B1924_;
  assign new_B399_ = new_B1957_;
  assign new_B400_ = new_B1990_;
  assign new_B401_ = new_B2023_;
  assign new_B402_ = new_B408_ & new_B407_;
  assign new_B403_ = new_B410_ | new_B409_;
  assign new_B404_ = new_B412_ | new_B411_;
  assign new_B405_ = new_B407_ & new_B413_;
  assign new_B406_ = new_B407_ & new_B414_;
  assign new_B407_ = new_B397_ ^ new_B398_;
  assign new_B408_ = new_B409_ ^ new_B399_;
  assign new_B409_ = new_B417_ & new_B416_;
  assign new_B410_ = new_B415_ & new_B399_;
  assign new_B411_ = new_B420_ & new_B419_;
  assign new_B412_ = new_B418_ & new_B399_;
  assign new_B413_ = new_B421_ | new_B398_;
  assign new_B414_ = ~new_B399_ ^ new_B411_;
  assign new_B415_ = ~new_B424_ | ~new_B425_;
  assign new_B416_ = new_B400_ ^ new_B407_;
  assign new_B417_ = new_B426_ & new_B419_;
  assign new_B418_ = ~new_B428_ | ~new_B427_;
  assign new_B419_ = new_B400_ | new_B401_;
  assign new_B420_ = new_B400_ | new_B407_;
  assign new_B421_ = new_B399_ & new_B411_;
  assign new_B422_ = ~new_B398_ | ~new_B399_;
  assign new_B423_ = new_B407_ & new_B422_;
  assign new_B424_ = ~new_B423_ & ~new_B407_;
  assign new_B425_ = new_B407_ | new_B422_;
  assign new_B426_ = ~new_B400_ | ~new_B401_;
  assign new_B427_ = new_B407_ | new_B422_;
  assign new_B428_ = ~new_B407_ & ~new_B429_;
  assign new_B429_ = new_B407_ & new_B422_;
  assign new_B430_ = new_B2056_;
  assign new_B431_ = new_B2089_;
  assign new_B432_ = new_B2122_;
  assign new_B433_ = new_B2155_;
  assign new_B434_ = new_B2188_;
  assign new_B435_ = new_B441_ & new_B440_;
  assign new_B436_ = new_B443_ | new_B442_;
  assign new_B437_ = new_B445_ | new_B444_;
  assign new_B438_ = new_B440_ & new_B446_;
  assign new_B439_ = new_B440_ & new_B447_;
  assign new_B440_ = new_B430_ ^ new_B431_;
  assign new_B441_ = new_B442_ ^ new_B432_;
  assign new_B442_ = new_B450_ & new_B449_;
  assign new_B443_ = new_B448_ & new_B432_;
  assign new_B444_ = new_B453_ & new_B452_;
  assign new_B445_ = new_B451_ & new_B432_;
  assign new_B446_ = new_B454_ | new_B431_;
  assign new_B447_ = ~new_B432_ ^ new_B444_;
  assign new_B448_ = ~new_B457_ | ~new_B458_;
  assign new_B449_ = new_B433_ ^ new_B440_;
  assign new_B450_ = new_B459_ & new_B452_;
  assign new_B451_ = ~new_B461_ | ~new_B460_;
  assign new_B452_ = new_B433_ | new_B434_;
  assign new_B453_ = new_B433_ | new_B440_;
  assign new_B454_ = new_B432_ & new_B444_;
  assign new_B455_ = ~new_B431_ | ~new_B432_;
  assign new_B456_ = new_B440_ & new_B455_;
  assign new_B457_ = ~new_B456_ & ~new_B440_;
  assign new_B458_ = new_B440_ | new_B455_;
  assign new_B459_ = ~new_B433_ | ~new_B434_;
  assign new_B460_ = new_B440_ | new_B455_;
  assign new_B461_ = ~new_B440_ & ~new_B462_;
  assign new_B462_ = new_B440_ & new_B455_;
  assign new_B463_ = new_B2221_;
  assign new_B464_ = new_B2254_;
  assign new_B465_ = new_B2287_;
  assign new_B466_ = new_B2320_;
  assign new_B467_ = new_B2353_;
  assign new_B468_ = new_B474_ & new_B473_;
  assign new_B469_ = new_B476_ | new_B475_;
  assign new_B470_ = new_B478_ | new_B477_;
  assign new_B471_ = new_B473_ & new_B479_;
  assign new_B472_ = new_B473_ & new_B480_;
  assign new_B473_ = new_B463_ ^ new_B464_;
  assign new_B474_ = new_B475_ ^ new_B465_;
  assign new_B475_ = new_B483_ & new_B482_;
  assign new_B476_ = new_B481_ & new_B465_;
  assign new_B477_ = new_B486_ & new_B485_;
  assign new_B478_ = new_B484_ & new_B465_;
  assign new_B479_ = new_B487_ | new_B464_;
  assign new_B480_ = ~new_B465_ ^ new_B477_;
  assign new_B481_ = ~new_B490_ | ~new_B491_;
  assign new_B482_ = new_B466_ ^ new_B473_;
  assign new_B483_ = new_B492_ & new_B485_;
  assign new_B484_ = ~new_B494_ | ~new_B493_;
  assign new_B485_ = new_B466_ | new_B467_;
  assign new_B486_ = new_B466_ | new_B473_;
  assign new_B487_ = new_B465_ & new_B477_;
  assign new_B488_ = ~new_B464_ | ~new_B465_;
  assign new_B489_ = new_B473_ & new_B488_;
  assign new_B490_ = ~new_B489_ & ~new_B473_;
  assign new_B491_ = new_B473_ | new_B488_;
  assign new_B492_ = ~new_B466_ | ~new_B467_;
  assign new_B493_ = new_B473_ | new_B488_;
  assign new_B494_ = ~new_B473_ & ~new_B495_;
  assign new_B495_ = new_B473_ & new_B488_;
  assign new_B496_ = new_B2386_;
  assign new_B497_ = new_B2419_;
  assign new_B498_ = new_B2452_;
  assign new_B499_ = new_B2485_;
  assign new_B500_ = new_B2518_;
  assign new_B501_ = new_B507_ & new_B506_;
  assign new_B502_ = new_B509_ | new_B508_;
  assign new_B503_ = new_B511_ | new_B510_;
  assign new_B504_ = new_B506_ & new_B512_;
  assign new_B505_ = new_B506_ & new_B513_;
  assign new_B506_ = new_B496_ ^ new_B497_;
  assign new_B507_ = new_B508_ ^ new_B498_;
  assign new_B508_ = new_B516_ & new_B515_;
  assign new_B509_ = new_B514_ & new_B498_;
  assign new_B510_ = new_B519_ & new_B518_;
  assign new_B511_ = new_B517_ & new_B498_;
  assign new_B512_ = new_B520_ | new_B497_;
  assign new_B513_ = ~new_B498_ ^ new_B510_;
  assign new_B514_ = ~new_B523_ | ~new_B524_;
  assign new_B515_ = new_B499_ ^ new_B506_;
  assign new_B516_ = new_B525_ & new_B518_;
  assign new_B517_ = ~new_B527_ | ~new_B526_;
  assign new_B518_ = new_B499_ | new_B500_;
  assign new_B519_ = new_B499_ | new_B506_;
  assign new_B520_ = new_B498_ & new_B510_;
  assign new_B521_ = ~new_B497_ | ~new_B498_;
  assign new_B522_ = new_B506_ & new_B521_;
  assign new_B523_ = ~new_B522_ & ~new_B506_;
  assign new_B524_ = new_B506_ | new_B521_;
  assign new_B525_ = ~new_B499_ | ~new_B500_;
  assign new_B526_ = new_B506_ | new_B521_;
  assign new_B527_ = ~new_B506_ & ~new_B528_;
  assign new_B528_ = new_B506_ & new_B521_;
  assign new_B529_ = new_B2551_;
  assign new_B530_ = new_B2584_;
  assign new_B531_ = new_B2617_;
  assign new_B532_ = new_B2650_;
  assign new_B533_ = new_B2683_;
  assign new_B534_ = new_B540_ & new_B539_;
  assign new_B535_ = new_B542_ | new_B541_;
  assign new_B536_ = new_B544_ | new_B543_;
  assign new_B537_ = new_B539_ & new_B545_;
  assign new_B538_ = new_B539_ & new_B546_;
  assign new_B539_ = new_B529_ ^ new_B530_;
  assign new_B540_ = new_B541_ ^ new_B531_;
  assign new_B541_ = new_B549_ & new_B548_;
  assign new_B542_ = new_B547_ & new_B531_;
  assign new_B543_ = new_B552_ & new_B551_;
  assign new_B544_ = new_B550_ & new_B531_;
  assign new_B545_ = new_B553_ | new_B530_;
  assign new_B546_ = ~new_B531_ ^ new_B543_;
  assign new_B547_ = ~new_B556_ | ~new_B557_;
  assign new_B548_ = new_B532_ ^ new_B539_;
  assign new_B549_ = new_B558_ & new_B551_;
  assign new_B550_ = ~new_B560_ | ~new_B559_;
  assign new_B551_ = new_B532_ | new_B533_;
  assign new_B552_ = new_B532_ | new_B539_;
  assign new_B553_ = new_B531_ & new_B543_;
  assign new_B554_ = ~new_B530_ | ~new_B531_;
  assign new_B555_ = new_B539_ & new_B554_;
  assign new_B556_ = ~new_B555_ & ~new_B539_;
  assign new_B557_ = new_B539_ | new_B554_;
  assign new_B558_ = ~new_B532_ | ~new_B533_;
  assign new_B559_ = new_B539_ | new_B554_;
  assign new_B560_ = ~new_B539_ & ~new_B561_;
  assign new_B561_ = new_B539_ & new_B554_;
  assign new_B562_ = new_B2716_;
  assign new_B563_ = new_B2749_;
  assign new_B564_ = new_B2782_;
  assign new_B565_ = new_B2815_;
  assign new_B566_ = new_B2848_;
  assign new_B567_ = new_B573_ & new_B572_;
  assign new_B568_ = new_B575_ | new_B574_;
  assign new_B569_ = new_B577_ | new_B576_;
  assign new_B570_ = new_B572_ & new_B578_;
  assign new_B571_ = new_B572_ & new_B579_;
  assign new_B572_ = new_B562_ ^ new_B563_;
  assign new_B573_ = new_B574_ ^ new_B564_;
  assign new_B574_ = new_B582_ & new_B581_;
  assign new_B575_ = new_B580_ & new_B564_;
  assign new_B576_ = new_B585_ & new_B584_;
  assign new_B577_ = new_B583_ & new_B564_;
  assign new_B578_ = new_B586_ | new_B563_;
  assign new_B579_ = ~new_B564_ ^ new_B576_;
  assign new_B580_ = ~new_B589_ | ~new_B590_;
  assign new_B581_ = new_B565_ ^ new_B572_;
  assign new_B582_ = new_B591_ & new_B584_;
  assign new_B583_ = ~new_B593_ | ~new_B592_;
  assign new_B584_ = new_B565_ | new_B566_;
  assign new_B585_ = new_B565_ | new_B572_;
  assign new_B586_ = new_B564_ & new_B576_;
  assign new_B587_ = ~new_B563_ | ~new_B564_;
  assign new_B588_ = new_B572_ & new_B587_;
  assign new_B589_ = ~new_B588_ & ~new_B572_;
  assign new_B590_ = new_B572_ | new_B587_;
  assign new_B591_ = ~new_B565_ | ~new_B566_;
  assign new_B592_ = new_B572_ | new_B587_;
  assign new_B593_ = ~new_B572_ & ~new_B594_;
  assign new_B594_ = new_B572_ & new_B587_;
  assign new_B595_ = new_B2881_;
  assign new_B596_ = new_B2914_;
  assign new_B597_ = new_B2947_;
  assign new_B598_ = new_B2980_;
  assign new_B599_ = new_B3013_;
  assign new_B600_ = new_B606_ & new_B605_;
  assign new_B601_ = new_B608_ | new_B607_;
  assign new_B602_ = new_B610_ | new_B609_;
  assign new_B603_ = new_B605_ & new_B611_;
  assign new_B604_ = new_B605_ & new_B612_;
  assign new_B605_ = new_B595_ ^ new_B596_;
  assign new_B606_ = new_B607_ ^ new_B597_;
  assign new_B607_ = new_B615_ & new_B614_;
  assign new_B608_ = new_B613_ & new_B597_;
  assign new_B609_ = new_B618_ & new_B617_;
  assign new_B610_ = new_B616_ & new_B597_;
  assign new_B611_ = new_B619_ | new_B596_;
  assign new_B612_ = ~new_B597_ ^ new_B609_;
  assign new_B613_ = ~new_B622_ | ~new_B623_;
  assign new_B614_ = new_B598_ ^ new_B605_;
  assign new_B615_ = new_B624_ & new_B617_;
  assign new_B616_ = ~new_B626_ | ~new_B625_;
  assign new_B617_ = new_B598_ | new_B599_;
  assign new_B618_ = new_B598_ | new_B605_;
  assign new_B619_ = new_B597_ & new_B609_;
  assign new_B620_ = ~new_B596_ | ~new_B597_;
  assign new_B621_ = new_B605_ & new_B620_;
  assign new_B622_ = ~new_B621_ & ~new_B605_;
  assign new_B623_ = new_B605_ | new_B620_;
  assign new_B624_ = ~new_B598_ | ~new_B599_;
  assign new_B625_ = new_B605_ | new_B620_;
  assign new_B626_ = ~new_B605_ & ~new_B627_;
  assign new_B627_ = new_B605_ & new_B620_;
  assign new_B628_ = new_B3046_;
  assign new_B629_ = new_B3079_;
  assign new_B630_ = new_B3112_;
  assign new_B631_ = new_B3145_;
  assign new_B632_ = new_B3178_;
  assign new_B633_ = new_B639_ & new_B638_;
  assign new_B634_ = new_B641_ | new_B640_;
  assign new_B635_ = new_B643_ | new_B642_;
  assign new_B636_ = new_B638_ & new_B644_;
  assign new_B637_ = new_B638_ & new_B645_;
  assign new_B638_ = new_B628_ ^ new_B629_;
  assign new_B639_ = new_B640_ ^ new_B630_;
  assign new_B640_ = new_B648_ & new_B647_;
  assign new_B641_ = new_B646_ & new_B630_;
  assign new_B642_ = new_B651_ & new_B650_;
  assign new_B643_ = new_B649_ & new_B630_;
  assign new_B644_ = new_B652_ | new_B629_;
  assign new_B645_ = ~new_B630_ ^ new_B642_;
  assign new_B646_ = ~new_B655_ | ~new_B656_;
  assign new_B647_ = new_B631_ ^ new_B638_;
  assign new_B648_ = new_B657_ & new_B650_;
  assign new_B649_ = ~new_B659_ | ~new_B658_;
  assign new_B650_ = new_B631_ | new_B632_;
  assign new_B651_ = new_B631_ | new_B638_;
  assign new_B652_ = new_B630_ & new_B642_;
  assign new_B653_ = ~new_B629_ | ~new_B630_;
  assign new_B654_ = new_B638_ & new_B653_;
  assign new_B655_ = ~new_B654_ & ~new_B638_;
  assign new_B656_ = new_B638_ | new_B653_;
  assign new_B657_ = ~new_B631_ | ~new_B632_;
  assign new_B658_ = new_B638_ | new_B653_;
  assign new_B659_ = ~new_B638_ & ~new_B660_;
  assign new_B660_ = new_B638_ & new_B653_;
  assign new_B661_ = new_B3211_;
  assign new_B662_ = new_B3244_;
  assign new_B663_ = new_B3277_;
  assign new_B664_ = new_B3310_;
  assign new_B665_ = new_B3343_;
  assign new_B666_ = new_B672_ & new_B671_;
  assign new_B667_ = new_B674_ | new_B673_;
  assign new_B668_ = new_B676_ | new_B675_;
  assign new_B669_ = new_B671_ & new_B677_;
  assign new_B670_ = new_B671_ & new_B678_;
  assign new_B671_ = new_B661_ ^ new_B662_;
  assign new_B672_ = new_B673_ ^ new_B663_;
  assign new_B673_ = new_B681_ & new_B680_;
  assign new_B674_ = new_B679_ & new_B663_;
  assign new_B675_ = new_B684_ & new_B683_;
  assign new_B676_ = new_B682_ & new_B663_;
  assign new_B677_ = new_B685_ | new_B662_;
  assign new_B678_ = ~new_B663_ ^ new_B675_;
  assign new_B679_ = ~new_B688_ | ~new_B689_;
  assign new_B680_ = new_B664_ ^ new_B671_;
  assign new_B681_ = new_B690_ & new_B683_;
  assign new_B682_ = ~new_B692_ | ~new_B691_;
  assign new_B683_ = new_B664_ | new_B665_;
  assign new_B684_ = new_B664_ | new_B671_;
  assign new_B685_ = new_B663_ & new_B675_;
  assign new_B686_ = ~new_B662_ | ~new_B663_;
  assign new_B687_ = new_B671_ & new_B686_;
  assign new_B688_ = ~new_B687_ & ~new_B671_;
  assign new_B689_ = new_B671_ | new_B686_;
  assign new_B690_ = ~new_B664_ | ~new_B665_;
  assign new_B691_ = new_B671_ | new_B686_;
  assign new_B692_ = ~new_B671_ & ~new_B693_;
  assign new_B693_ = new_B671_ & new_B686_;
  assign new_B694_ = new_B3376_;
  assign new_B695_ = new_B3409_;
  assign new_B696_ = new_B3442_;
  assign new_B697_ = new_B3475_;
  assign new_B698_ = new_B3508_;
  assign new_B699_ = new_B705_ & new_B704_;
  assign new_B700_ = new_B707_ | new_B706_;
  assign new_B701_ = new_B709_ | new_B708_;
  assign new_B702_ = new_B704_ & new_B710_;
  assign new_B703_ = new_B704_ & new_B711_;
  assign new_B704_ = new_B694_ ^ new_B695_;
  assign new_B705_ = new_B706_ ^ new_B696_;
  assign new_B706_ = new_B714_ & new_B713_;
  assign new_B707_ = new_B712_ & new_B696_;
  assign new_B708_ = new_B717_ & new_B716_;
  assign new_B709_ = new_B715_ & new_B696_;
  assign new_B710_ = new_B718_ | new_B695_;
  assign new_B711_ = ~new_B696_ ^ new_B708_;
  assign new_B712_ = ~new_B721_ | ~new_B722_;
  assign new_B713_ = new_B697_ ^ new_B704_;
  assign new_B714_ = new_B723_ & new_B716_;
  assign new_B715_ = ~new_B725_ | ~new_B724_;
  assign new_B716_ = new_B697_ | new_B698_;
  assign new_B717_ = new_B697_ | new_B704_;
  assign new_B718_ = new_B696_ & new_B708_;
  assign new_B719_ = ~new_B695_ | ~new_B696_;
  assign new_B720_ = new_B704_ & new_B719_;
  assign new_B721_ = ~new_B720_ & ~new_B704_;
  assign new_B722_ = new_B704_ | new_B719_;
  assign new_B723_ = ~new_B697_ | ~new_B698_;
  assign new_B724_ = new_B704_ | new_B719_;
  assign new_B725_ = ~new_B704_ & ~new_B726_;
  assign new_B726_ = new_B704_ & new_B719_;
  assign new_B727_ = new_B3541_;
  assign new_B728_ = new_B3574_;
  assign new_B729_ = new_B3607_;
  assign new_B730_ = new_B3640_;
  assign new_B731_ = new_B3673_;
  assign new_B732_ = new_B738_ & new_B737_;
  assign new_B733_ = new_B740_ | new_B739_;
  assign new_B734_ = new_B742_ | new_B741_;
  assign new_B735_ = new_B737_ & new_B743_;
  assign new_B736_ = new_B737_ & new_B744_;
  assign new_B737_ = new_B727_ ^ new_B728_;
  assign new_B738_ = new_B739_ ^ new_B729_;
  assign new_B739_ = new_B747_ & new_B746_;
  assign new_B740_ = new_B745_ & new_B729_;
  assign new_B741_ = new_B750_ & new_B749_;
  assign new_B742_ = new_B748_ & new_B729_;
  assign new_B743_ = new_B751_ | new_B728_;
  assign new_B744_ = ~new_B729_ ^ new_B741_;
  assign new_B745_ = ~new_B754_ | ~new_B755_;
  assign new_B746_ = new_B730_ ^ new_B737_;
  assign new_B747_ = new_B756_ & new_B749_;
  assign new_B748_ = ~new_B758_ | ~new_B757_;
  assign new_B749_ = new_B730_ | new_B731_;
  assign new_B750_ = new_B730_ | new_B737_;
  assign new_B751_ = new_B729_ & new_B741_;
  assign new_B752_ = ~new_B728_ | ~new_B729_;
  assign new_B753_ = new_B737_ & new_B752_;
  assign new_B754_ = ~new_B753_ & ~new_B737_;
  assign new_B755_ = new_B737_ | new_B752_;
  assign new_B756_ = ~new_B730_ | ~new_B731_;
  assign new_B757_ = new_B737_ | new_B752_;
  assign new_B758_ = ~new_B737_ & ~new_B759_;
  assign new_B759_ = new_B737_ & new_B752_;
  assign new_B760_ = new_B3706_;
  assign new_B761_ = new_B3739_;
  assign new_B762_ = new_B3772_;
  assign new_B763_ = new_B3805_;
  assign new_B764_ = new_B3838_;
  assign new_B765_ = new_B771_ & new_B770_;
  assign new_B766_ = new_B773_ | new_B772_;
  assign new_B767_ = new_B775_ | new_B774_;
  assign new_B768_ = new_B770_ & new_B776_;
  assign new_B769_ = new_B770_ & new_B777_;
  assign new_B770_ = new_B760_ ^ new_B761_;
  assign new_B771_ = new_B772_ ^ new_B762_;
  assign new_B772_ = new_B780_ & new_B779_;
  assign new_B773_ = new_B778_ & new_B762_;
  assign new_B774_ = new_B783_ & new_B782_;
  assign new_B775_ = new_B781_ & new_B762_;
  assign new_B776_ = new_B784_ | new_B761_;
  assign new_B777_ = ~new_B762_ ^ new_B774_;
  assign new_B778_ = ~new_B787_ | ~new_B788_;
  assign new_B779_ = new_B763_ ^ new_B770_;
  assign new_B780_ = new_B789_ & new_B782_;
  assign new_B781_ = ~new_B791_ | ~new_B790_;
  assign new_B782_ = new_B763_ | new_B764_;
  assign new_B783_ = new_B763_ | new_B770_;
  assign new_B784_ = new_B762_ & new_B774_;
  assign new_B785_ = ~new_B761_ | ~new_B762_;
  assign new_B786_ = new_B770_ & new_B785_;
  assign new_B787_ = ~new_B786_ & ~new_B770_;
  assign new_B788_ = new_B770_ | new_B785_;
  assign new_B789_ = ~new_B763_ | ~new_B764_;
  assign new_B790_ = new_B770_ | new_B785_;
  assign new_B791_ = ~new_B770_ & ~new_B792_;
  assign new_B792_ = new_B770_ & new_B785_;
  assign new_B793_ = new_B3871_;
  assign new_B794_ = new_B3904_;
  assign new_B795_ = new_B3937_;
  assign new_B796_ = new_B3970_;
  assign new_B797_ = new_B4003_;
  assign new_B798_ = new_B804_ & new_B803_;
  assign new_B799_ = new_B806_ | new_B805_;
  assign new_B800_ = new_B808_ | new_B807_;
  assign new_B801_ = new_B803_ & new_B809_;
  assign new_B802_ = new_B803_ & new_B810_;
  assign new_B803_ = new_B793_ ^ new_B794_;
  assign new_B804_ = new_B805_ ^ new_B795_;
  assign new_B805_ = new_B813_ & new_B812_;
  assign new_B806_ = new_B811_ & new_B795_;
  assign new_B807_ = new_B816_ & new_B815_;
  assign new_B808_ = new_B814_ & new_B795_;
  assign new_B809_ = new_B817_ | new_B794_;
  assign new_B810_ = ~new_B795_ ^ new_B807_;
  assign new_B811_ = ~new_B820_ | ~new_B821_;
  assign new_B812_ = new_B796_ ^ new_B803_;
  assign new_B813_ = new_B822_ & new_B815_;
  assign new_B814_ = ~new_B824_ | ~new_B823_;
  assign new_B815_ = new_B796_ | new_B797_;
  assign new_B816_ = new_B796_ | new_B803_;
  assign new_B817_ = new_B795_ & new_B807_;
  assign new_B818_ = ~new_B794_ | ~new_B795_;
  assign new_B819_ = new_B803_ & new_B818_;
  assign new_B820_ = ~new_B819_ & ~new_B803_;
  assign new_B821_ = new_B803_ | new_B818_;
  assign new_B822_ = ~new_B796_ | ~new_B797_;
  assign new_B823_ = new_B803_ | new_B818_;
  assign new_B824_ = ~new_B803_ & ~new_B825_;
  assign new_B825_ = new_B803_ & new_B818_;
  assign new_B826_ = new_B4036_;
  assign new_B827_ = new_B4069_;
  assign new_B828_ = new_B4102_;
  assign new_B829_ = new_B4135_;
  assign new_B830_ = new_B4168_;
  assign new_B831_ = new_B837_ & new_B836_;
  assign new_B832_ = new_B839_ | new_B838_;
  assign new_B833_ = new_B841_ | new_B840_;
  assign new_B834_ = new_B836_ & new_B842_;
  assign new_B835_ = new_B836_ & new_B843_;
  assign new_B836_ = new_B826_ ^ new_B827_;
  assign new_B837_ = new_B838_ ^ new_B828_;
  assign new_B838_ = new_B846_ & new_B845_;
  assign new_B839_ = new_B844_ & new_B828_;
  assign new_B840_ = new_B849_ & new_B848_;
  assign new_B841_ = new_B847_ & new_B828_;
  assign new_B842_ = new_B850_ | new_B827_;
  assign new_B843_ = ~new_B828_ ^ new_B840_;
  assign new_B844_ = ~new_B853_ | ~new_B854_;
  assign new_B845_ = new_B829_ ^ new_B836_;
  assign new_B846_ = new_B855_ & new_B848_;
  assign new_B847_ = ~new_B857_ | ~new_B856_;
  assign new_B848_ = new_B829_ | new_B830_;
  assign new_B849_ = new_B829_ | new_B836_;
  assign new_B850_ = new_B828_ & new_B840_;
  assign new_B851_ = ~new_B827_ | ~new_B828_;
  assign new_B852_ = new_B836_ & new_B851_;
  assign new_B853_ = ~new_B852_ & ~new_B836_;
  assign new_B854_ = new_B836_ | new_B851_;
  assign new_B855_ = ~new_B829_ | ~new_B830_;
  assign new_B856_ = new_B836_ | new_B851_;
  assign new_B857_ = ~new_B836_ & ~new_B858_;
  assign new_B858_ = new_B836_ & new_B851_;
  assign new_B859_ = new_B4201_;
  assign new_B860_ = new_B4234_;
  assign new_B861_ = new_B4267_;
  assign new_B862_ = new_B4300_;
  assign new_B863_ = new_B4333_;
  assign new_B864_ = new_B870_ & new_B869_;
  assign new_B865_ = new_B872_ | new_B871_;
  assign new_B866_ = new_B874_ | new_B873_;
  assign new_B867_ = new_B869_ & new_B875_;
  assign new_B868_ = new_B869_ & new_B876_;
  assign new_B869_ = new_B859_ ^ new_B860_;
  assign new_B870_ = new_B871_ ^ new_B861_;
  assign new_B871_ = new_B879_ & new_B878_;
  assign new_B872_ = new_B877_ & new_B861_;
  assign new_B873_ = new_B882_ & new_B881_;
  assign new_B874_ = new_B880_ & new_B861_;
  assign new_B875_ = new_B883_ | new_B860_;
  assign new_B876_ = ~new_B861_ ^ new_B873_;
  assign new_B877_ = ~new_B886_ | ~new_B887_;
  assign new_B878_ = new_B862_ ^ new_B869_;
  assign new_B879_ = new_B888_ & new_B881_;
  assign new_B880_ = ~new_B890_ | ~new_B889_;
  assign new_B881_ = new_B862_ | new_B863_;
  assign new_B882_ = new_B862_ | new_B869_;
  assign new_B883_ = new_B861_ & new_B873_;
  assign new_B884_ = ~new_B860_ | ~new_B861_;
  assign new_B885_ = new_B869_ & new_B884_;
  assign new_B886_ = ~new_B885_ & ~new_B869_;
  assign new_B887_ = new_B869_ | new_B884_;
  assign new_B888_ = ~new_B862_ | ~new_B863_;
  assign new_B889_ = new_B869_ | new_B884_;
  assign new_B890_ = ~new_B869_ & ~new_B891_;
  assign new_B891_ = new_B869_ & new_B884_;
  assign new_B892_ = new_B4366_;
  assign new_B893_ = new_B4399_;
  assign new_B894_ = new_B4432_;
  assign new_B895_ = new_B4465_;
  assign new_B896_ = new_B4498_;
  assign new_B897_ = new_B903_ & new_B902_;
  assign new_B898_ = new_B905_ | new_B904_;
  assign new_B899_ = new_B907_ | new_B906_;
  assign new_B900_ = new_B902_ & new_B908_;
  assign new_B901_ = new_B902_ & new_B909_;
  assign new_B902_ = new_B892_ ^ new_B893_;
  assign new_B903_ = new_B904_ ^ new_B894_;
  assign new_B904_ = new_B912_ & new_B911_;
  assign new_B905_ = new_B910_ & new_B894_;
  assign new_B906_ = new_B915_ & new_B914_;
  assign new_B907_ = new_B913_ & new_B894_;
  assign new_B908_ = new_B916_ | new_B893_;
  assign new_B909_ = ~new_B894_ ^ new_B906_;
  assign new_B910_ = ~new_B919_ | ~new_B920_;
  assign new_B911_ = new_B895_ ^ new_B902_;
  assign new_B912_ = new_B921_ & new_B914_;
  assign new_B913_ = ~new_B923_ | ~new_B922_;
  assign new_B914_ = new_B895_ | new_B896_;
  assign new_B915_ = new_B895_ | new_B902_;
  assign new_B916_ = new_B894_ & new_B906_;
  assign new_B917_ = ~new_B893_ | ~new_B894_;
  assign new_B918_ = new_B902_ & new_B917_;
  assign new_B919_ = ~new_B918_ & ~new_B902_;
  assign new_B920_ = new_B902_ | new_B917_;
  assign new_B921_ = ~new_B895_ | ~new_B896_;
  assign new_B922_ = new_B902_ | new_B917_;
  assign new_B923_ = ~new_B902_ & ~new_B924_;
  assign new_B924_ = new_B902_ & new_B917_;
  assign new_B925_ = new_B4531_;
  assign new_B926_ = new_B4564_;
  assign new_B927_ = new_B4597_;
  assign new_B928_ = new_B4630_;
  assign new_B929_ = new_B4663_;
  assign new_B930_ = new_B936_ & new_B935_;
  assign new_B931_ = new_B938_ | new_B937_;
  assign new_B932_ = new_B940_ | new_B939_;
  assign new_B933_ = new_B935_ & new_B941_;
  assign new_B934_ = new_B935_ & new_B942_;
  assign new_B935_ = new_B925_ ^ new_B926_;
  assign new_B936_ = new_B937_ ^ new_B927_;
  assign new_B937_ = new_B945_ & new_B944_;
  assign new_B938_ = new_B943_ & new_B927_;
  assign new_B939_ = new_B948_ & new_B947_;
  assign new_B940_ = new_B946_ & new_B927_;
  assign new_B941_ = new_B949_ | new_B926_;
  assign new_B942_ = ~new_B927_ ^ new_B939_;
  assign new_B943_ = ~new_B952_ | ~new_B953_;
  assign new_B944_ = new_B928_ ^ new_B935_;
  assign new_B945_ = new_B954_ & new_B947_;
  assign new_B946_ = ~new_B956_ | ~new_B955_;
  assign new_B947_ = new_B928_ | new_B929_;
  assign new_B948_ = new_B928_ | new_B935_;
  assign new_B949_ = new_B927_ & new_B939_;
  assign new_B950_ = ~new_B926_ | ~new_B927_;
  assign new_B951_ = new_B935_ & new_B950_;
  assign new_B952_ = ~new_B951_ & ~new_B935_;
  assign new_B953_ = new_B935_ | new_B950_;
  assign new_B954_ = ~new_B928_ | ~new_B929_;
  assign new_B955_ = new_B935_ | new_B950_;
  assign new_B956_ = ~new_B935_ & ~new_B957_;
  assign new_B957_ = new_B935_ & new_B950_;
  assign new_B958_ = new_B4696_;
  assign new_B959_ = new_B4729_;
  assign new_B960_ = new_B4762_;
  assign new_B961_ = new_B4795_;
  assign new_B962_ = new_B4828_;
  assign new_B963_ = new_B969_ & new_B968_;
  assign new_B964_ = new_B971_ | new_B970_;
  assign new_B965_ = new_B973_ | new_B972_;
  assign new_B966_ = new_B968_ & new_B974_;
  assign new_B967_ = new_B968_ & new_B975_;
  assign new_B968_ = new_B958_ ^ new_B959_;
  assign new_B969_ = new_B970_ ^ new_B960_;
  assign new_B970_ = new_B978_ & new_B977_;
  assign new_B971_ = new_B976_ & new_B960_;
  assign new_B972_ = new_B981_ & new_B980_;
  assign new_B973_ = new_B979_ & new_B960_;
  assign new_B974_ = new_B982_ | new_B959_;
  assign new_B975_ = ~new_B960_ ^ new_B972_;
  assign new_B976_ = ~new_B985_ | ~new_B986_;
  assign new_B977_ = new_B961_ ^ new_B968_;
  assign new_B978_ = new_B987_ & new_B980_;
  assign new_B979_ = ~new_B989_ | ~new_B988_;
  assign new_B980_ = new_B961_ | new_B962_;
  assign new_B981_ = new_B961_ | new_B968_;
  assign new_B982_ = new_B960_ & new_B972_;
  assign new_B983_ = ~new_B959_ | ~new_B960_;
  assign new_B984_ = new_B968_ & new_B983_;
  assign new_B985_ = ~new_B984_ & ~new_B968_;
  assign new_B986_ = new_B968_ | new_B983_;
  assign new_B987_ = ~new_B961_ | ~new_B962_;
  assign new_B988_ = new_B968_ | new_B983_;
  assign new_B989_ = ~new_B968_ & ~new_B990_;
  assign new_B990_ = new_B968_ & new_B983_;
  assign new_B991_ = new_B4861_;
  assign new_B992_ = new_B4894_;
  assign new_B993_ = new_B4927_;
  assign new_B994_ = new_B4960_;
  assign new_B995_ = new_B4993_;
  assign new_B996_ = new_B1002_ & new_B1001_;
  assign new_B997_ = new_B1004_ | new_B1003_;
  assign new_B998_ = new_B1006_ | new_B1005_;
  assign new_B999_ = new_B1001_ & new_B1007_;
  assign new_B1000_ = new_B1001_ & new_B1008_;
  assign new_B1001_ = new_B991_ ^ new_B992_;
  assign new_B1002_ = new_B1003_ ^ new_B993_;
  assign new_B1003_ = new_B1011_ & new_B1010_;
  assign new_B1004_ = new_B1009_ & new_B993_;
  assign new_B1005_ = new_B1014_ & new_B1013_;
  assign new_B1006_ = new_B1012_ & new_B993_;
  assign new_B1007_ = new_B1015_ | new_B992_;
  assign new_B1008_ = ~new_B993_ ^ new_B1005_;
  assign new_B1009_ = ~new_B1018_ | ~new_B1019_;
  assign new_B1010_ = new_B994_ ^ new_B1001_;
  assign new_B1011_ = new_B1020_ & new_B1013_;
  assign new_B1012_ = ~new_B1022_ | ~new_B1021_;
  assign new_B1013_ = new_B994_ | new_B995_;
  assign new_B1014_ = new_B994_ | new_B1001_;
  assign new_B1015_ = new_B993_ & new_B1005_;
  assign new_B1016_ = ~new_B992_ | ~new_B993_;
  assign new_B1017_ = new_B1001_ & new_B1016_;
  assign new_B1018_ = ~new_B1017_ & ~new_B1001_;
  assign new_B1019_ = new_B1001_ | new_B1016_;
  assign new_B1020_ = ~new_B994_ | ~new_B995_;
  assign new_B1021_ = new_B1001_ | new_B1016_;
  assign new_B1022_ = ~new_B1001_ & ~new_B1023_;
  assign new_B1023_ = new_B1001_ & new_B1016_;
  assign new_B1024_ = new_B5026_;
  assign new_B1025_ = new_B5059_;
  assign new_B1026_ = new_B5092_;
  assign new_B1027_ = new_B5125_;
  assign new_B1028_ = new_B5158_;
  assign new_B1029_ = new_B1035_ & new_B1034_;
  assign new_B1030_ = new_B1037_ | new_B1036_;
  assign new_B1031_ = new_B1039_ | new_B1038_;
  assign new_B1032_ = new_B1034_ & new_B1040_;
  assign new_B1033_ = new_B1034_ & new_B1041_;
  assign new_B1034_ = new_B1024_ ^ new_B1025_;
  assign new_B1035_ = new_B1036_ ^ new_B1026_;
  assign new_B1036_ = new_B1044_ & new_B1043_;
  assign new_B1037_ = new_B1042_ & new_B1026_;
  assign new_B1038_ = new_B1047_ & new_B1046_;
  assign new_B1039_ = new_B1045_ & new_B1026_;
  assign new_B1040_ = new_B1048_ | new_B1025_;
  assign new_B1041_ = ~new_B1026_ ^ new_B1038_;
  assign new_B1042_ = ~new_B1051_ | ~new_B1052_;
  assign new_B1043_ = new_B1027_ ^ new_B1034_;
  assign new_B1044_ = new_B1053_ & new_B1046_;
  assign new_B1045_ = ~new_B1055_ | ~new_B1054_;
  assign new_B1046_ = new_B1027_ | new_B1028_;
  assign new_B1047_ = new_B1027_ | new_B1034_;
  assign new_B1048_ = new_B1026_ & new_B1038_;
  assign new_B1049_ = ~new_B1025_ | ~new_B1026_;
  assign new_B1050_ = new_B1034_ & new_B1049_;
  assign new_B1051_ = ~new_B1050_ & ~new_B1034_;
  assign new_B1052_ = new_B1034_ | new_B1049_;
  assign new_B1053_ = ~new_B1027_ | ~new_B1028_;
  assign new_B1054_ = new_B1034_ | new_B1049_;
  assign new_B1055_ = ~new_B1034_ & ~new_B1056_;
  assign new_B1056_ = new_B1034_ & new_B1049_;
  assign new_A6930_ = new_A6908_ & new_A6923_;
  assign new_A6929_ = ~new_A6908_ & ~new_A6930_;
  assign new_A6928_ = new_A6908_ | new_A6923_;
  assign new_A6927_ = ~new_A6901_ | ~new_A6902_;
  assign new_A6926_ = new_A6908_ | new_A6923_;
  assign new_A6925_ = ~new_A6924_ & ~new_A6908_;
  assign new_A6924_ = new_A6908_ & new_A6923_;
  assign new_A6923_ = ~new_A6899_ | ~new_A6900_;
  assign new_A6922_ = new_A6900_ & new_A6912_;
  assign new_A6921_ = new_A6901_ | new_A6908_;
  assign new_A6920_ = new_A6901_ | new_A6902_;
  assign new_A6919_ = ~new_A6929_ | ~new_A6928_;
  assign new_A6918_ = new_A6927_ & new_A6920_;
  assign new_A6917_ = new_A6901_ ^ new_A6908_;
  assign new_A6916_ = ~new_A6925_ | ~new_A6926_;
  assign new_A6915_ = ~new_A6900_ ^ new_A6912_;
  assign new_A6914_ = new_A6922_ | new_A6899_;
  assign new_A6913_ = new_A6919_ & new_A6900_;
  assign new_A6912_ = new_A6921_ & new_A6920_;
  assign new_A6911_ = new_A6916_ & new_A6900_;
  assign new_A6910_ = new_A6918_ & new_A6917_;
  assign new_A6909_ = new_A6910_ ^ new_A6900_;
  assign new_A6908_ = new_A6898_ ^ new_A6899_;
  assign A6907 = new_A6908_ & new_A6915_;
  assign A6906 = new_A6908_ & new_A6914_;
  assign A6905 = new_A6913_ | new_A6912_;
  assign A6904 = new_A6911_ | new_A6910_;
  assign A6903 = new_A6909_ & new_A6908_;
  assign new_A6902_ = new_B1033_;
  assign new_A6901_ = new_B1000_;
  assign new_A6900_ = new_B967_;
  assign new_A6899_ = new_B934_;
  assign new_A6898_ = new_B901_;
  assign new_A6897_ = new_A6875_ & new_A6890_;
  assign new_A6896_ = ~new_A6875_ & ~new_A6897_;
  assign new_A6895_ = new_A6875_ | new_A6890_;
  assign new_A6894_ = ~new_A6868_ | ~new_A6869_;
  assign new_A6893_ = new_A6875_ | new_A6890_;
  assign new_A6892_ = ~new_A6891_ & ~new_A6875_;
  assign new_A6891_ = new_A6875_ & new_A6890_;
  assign new_A6890_ = ~new_A6866_ | ~new_A6867_;
  assign new_A6889_ = new_A6867_ & new_A6879_;
  assign new_A6888_ = new_A6868_ | new_A6875_;
  assign new_A6887_ = new_A6868_ | new_A6869_;
  assign new_A6886_ = ~new_A6896_ | ~new_A6895_;
  assign new_A6885_ = new_A6894_ & new_A6887_;
  assign new_A6884_ = new_A6868_ ^ new_A6875_;
  assign new_A6883_ = ~new_A6892_ | ~new_A6893_;
  assign new_A6882_ = ~new_A6867_ ^ new_A6879_;
  assign new_A6881_ = new_A6889_ | new_A6866_;
  assign new_A6880_ = new_A6886_ & new_A6867_;
  assign new_A6879_ = new_A6888_ & new_A6887_;
  assign new_A6878_ = new_A6883_ & new_A6867_;
  assign new_A6877_ = new_A6885_ & new_A6884_;
  assign new_A6876_ = new_A6877_ ^ new_A6867_;
  assign new_A6875_ = new_A6865_ ^ new_A6866_;
  assign A6874 = new_A6875_ & new_A6882_;
  assign A6873 = new_A6875_ & new_A6881_;
  assign A6872 = new_A6880_ | new_A6879_;
  assign A6871 = new_A6878_ | new_A6877_;
  assign A6870 = new_A6876_ & new_A6875_;
  assign new_A6869_ = new_B868_;
  assign new_A6868_ = new_B835_;
  assign new_A6867_ = new_B802_;
  assign new_A6866_ = new_B769_;
  assign new_A6865_ = new_B736_;
  assign new_A6864_ = new_A6842_ & new_A6857_;
  assign new_A6863_ = ~new_A6842_ & ~new_A6864_;
  assign new_A6862_ = new_A6842_ | new_A6857_;
  assign new_A6861_ = ~new_A6835_ | ~new_A6836_;
  assign new_A6860_ = new_A6842_ | new_A6857_;
  assign new_A6859_ = ~new_A6858_ & ~new_A6842_;
  assign new_A6858_ = new_A6842_ & new_A6857_;
  assign new_A6857_ = ~new_A6833_ | ~new_A6834_;
  assign new_A6856_ = new_A6834_ & new_A6846_;
  assign new_A6855_ = new_A6835_ | new_A6842_;
  assign new_A6854_ = new_A6835_ | new_A6836_;
  assign new_A6853_ = ~new_A6863_ | ~new_A6862_;
  assign new_A6852_ = new_A6861_ & new_A6854_;
  assign new_A6851_ = new_A6835_ ^ new_A6842_;
  assign new_A6850_ = ~new_A6859_ | ~new_A6860_;
  assign new_A6849_ = ~new_A6834_ ^ new_A6846_;
  assign new_A6848_ = new_A6856_ | new_A6833_;
  assign new_A6847_ = new_A6853_ & new_A6834_;
  assign new_A6846_ = new_A6855_ & new_A6854_;
  assign new_A6845_ = new_A6850_ & new_A6834_;
  assign new_A6844_ = new_A6852_ & new_A6851_;
  assign new_A6843_ = new_A6844_ ^ new_A6834_;
  assign new_A6842_ = new_A6832_ ^ new_A6833_;
  assign A6841 = new_A6842_ & new_A6849_;
  assign A6840 = new_A6842_ & new_A6848_;
  assign A6839 = new_A6847_ | new_A6846_;
  assign A6838 = new_A6845_ | new_A6844_;
  assign A6837 = new_A6843_ & new_A6842_;
  assign new_A6836_ = new_B703_;
  assign new_A6835_ = new_B670_;
  assign new_A6834_ = new_B637_;
  assign new_A6833_ = new_B604_;
  assign new_A6832_ = new_B571_;
  assign new_A6831_ = new_A6809_ & new_A6824_;
  assign new_A6830_ = ~new_A6809_ & ~new_A6831_;
  assign new_A6829_ = new_A6809_ | new_A6824_;
  assign new_A6828_ = ~new_A6802_ | ~new_A6803_;
  assign new_A6827_ = new_A6809_ | new_A6824_;
  assign new_A6826_ = ~new_A6825_ & ~new_A6809_;
  assign new_A6825_ = new_A6809_ & new_A6824_;
  assign new_A6824_ = ~new_A6800_ | ~new_A6801_;
  assign new_A6823_ = new_A6801_ & new_A6813_;
  assign new_A6822_ = new_A6802_ | new_A6809_;
  assign new_A6821_ = new_A6802_ | new_A6803_;
  assign new_A6820_ = ~new_A6830_ | ~new_A6829_;
  assign new_A6819_ = new_A6828_ & new_A6821_;
  assign new_A6818_ = new_A6802_ ^ new_A6809_;
  assign new_A6817_ = ~new_A6826_ | ~new_A6827_;
  assign new_A6816_ = ~new_A6801_ ^ new_A6813_;
  assign new_A6815_ = new_A6823_ | new_A6800_;
  assign new_A6814_ = new_A6820_ & new_A6801_;
  assign new_A6813_ = new_A6822_ & new_A6821_;
  assign new_A6812_ = new_A6817_ & new_A6801_;
  assign new_A6811_ = new_A6819_ & new_A6818_;
  assign new_A6810_ = new_A6811_ ^ new_A6801_;
  assign new_A6809_ = new_A6799_ ^ new_A6800_;
  assign A6808 = new_A6809_ & new_A6816_;
  assign A6807 = new_A6809_ & new_A6815_;
  assign A6806 = new_A6814_ | new_A6813_;
  assign A6805 = new_A6812_ | new_A6811_;
  assign A6804 = new_A6810_ & new_A6809_;
  assign new_A6803_ = new_B538_;
  assign new_A6802_ = new_B505_;
  assign new_A6801_ = new_B472_;
  assign new_A6800_ = new_B439_;
  assign new_A6799_ = new_B406_;
  assign new_A6798_ = new_A6776_ & new_A6791_;
  assign new_A6797_ = ~new_A6776_ & ~new_A6798_;
  assign new_A6796_ = new_A6776_ | new_A6791_;
  assign new_A6795_ = ~new_A6769_ | ~new_A6770_;
  assign new_A6794_ = new_A6776_ | new_A6791_;
  assign new_A6793_ = ~new_A6792_ & ~new_A6776_;
  assign new_A6792_ = new_A6776_ & new_A6791_;
  assign new_A6791_ = ~new_A6767_ | ~new_A6768_;
  assign new_A6790_ = new_A6768_ & new_A6780_;
  assign new_A6789_ = new_A6769_ | new_A6776_;
  assign new_A6788_ = new_A6769_ | new_A6770_;
  assign new_A6787_ = ~new_A6797_ | ~new_A6796_;
  assign new_A6786_ = new_A6795_ & new_A6788_;
  assign new_A6785_ = new_A6769_ ^ new_A6776_;
  assign new_A6784_ = ~new_A6793_ | ~new_A6794_;
  assign new_A6783_ = ~new_A6768_ ^ new_A6780_;
  assign new_A6782_ = new_A6790_ | new_A6767_;
  assign new_A6781_ = new_A6787_ & new_A6768_;
  assign new_A6780_ = new_A6789_ & new_A6788_;
  assign new_A6779_ = new_A6784_ & new_A6768_;
  assign new_A6778_ = new_A6786_ & new_A6785_;
  assign new_A6777_ = new_A6778_ ^ new_A6768_;
  assign new_A6776_ = new_A6766_ ^ new_A6767_;
  assign A6775 = new_A6776_ & new_A6783_;
  assign A6774 = new_A6776_ & new_A6782_;
  assign A6773 = new_A6781_ | new_A6780_;
  assign A6772 = new_A6779_ | new_A6778_;
  assign A6771 = new_A6777_ & new_A6776_;
  assign new_A6770_ = new_B373_;
  assign new_A6769_ = new_B340_;
  assign new_A6768_ = new_B307_;
  assign new_A6767_ = new_B274_;
  assign new_A6766_ = new_B241_;
  assign new_A6765_ = new_A6743_ & new_A6758_;
  assign new_A6764_ = ~new_A6743_ & ~new_A6765_;
  assign new_A6763_ = new_A6743_ | new_A6758_;
  assign new_A6762_ = ~new_A6736_ | ~new_A6737_;
  assign new_A6761_ = new_A6743_ | new_A6758_;
  assign new_A6760_ = ~new_A6759_ & ~new_A6743_;
  assign new_A6759_ = new_A6743_ & new_A6758_;
  assign new_A6758_ = ~new_A6734_ | ~new_A6735_;
  assign new_A6757_ = new_A6735_ & new_A6747_;
  assign new_A6756_ = new_A6736_ | new_A6743_;
  assign new_A6755_ = new_A6736_ | new_A6737_;
  assign new_A6754_ = ~new_A6764_ | ~new_A6763_;
  assign new_A6753_ = new_A6762_ & new_A6755_;
  assign new_A6752_ = new_A6736_ ^ new_A6743_;
  assign new_A6751_ = ~new_A6760_ | ~new_A6761_;
  assign new_A6750_ = ~new_A6735_ ^ new_A6747_;
  assign new_A6749_ = new_A6757_ | new_A6734_;
  assign new_A6748_ = new_A6754_ & new_A6735_;
  assign new_A6747_ = new_A6756_ & new_A6755_;
  assign new_A6746_ = new_A6751_ & new_A6735_;
  assign new_A6745_ = new_A6753_ & new_A6752_;
  assign new_A6744_ = new_A6745_ ^ new_A6735_;
  assign new_A6743_ = new_A6733_ ^ new_A6734_;
  assign A6742 = new_A6743_ & new_A6750_;
  assign A6741 = new_A6743_ & new_A6749_;
  assign A6740 = new_A6748_ | new_A6747_;
  assign A6739 = new_A6746_ | new_A6745_;
  assign A6738 = new_A6744_ & new_A6743_;
  assign new_A6737_ = new_B208_;
  assign new_A6736_ = new_B175_;
  assign new_A6735_ = new_B142_;
  assign new_A6734_ = new_B109_;
  assign new_A6733_ = new_B76_;
  assign new_A6732_ = new_A6710_ & new_A6725_;
  assign new_A6731_ = ~new_A6710_ & ~new_A6732_;
  assign new_A6730_ = new_A6710_ | new_A6725_;
  assign new_A6729_ = ~new_A6703_ | ~new_A6704_;
  assign new_A6728_ = new_A6710_ | new_A6725_;
  assign new_A6727_ = ~new_A6726_ & ~new_A6710_;
  assign new_A6726_ = new_A6710_ & new_A6725_;
  assign new_A6725_ = ~new_A6701_ | ~new_A6702_;
  assign new_A6724_ = new_A6702_ & new_A6714_;
  assign new_A6723_ = new_A6703_ | new_A6710_;
  assign new_A6722_ = new_A6703_ | new_A6704_;
  assign new_A6721_ = ~new_A6731_ | ~new_A6730_;
  assign new_A6720_ = new_A6729_ & new_A6722_;
  assign new_A6719_ = new_A6703_ ^ new_A6710_;
  assign new_A6718_ = ~new_A6727_ | ~new_A6728_;
  assign new_A6717_ = ~new_A6702_ ^ new_A6714_;
  assign new_A6716_ = new_A6724_ | new_A6701_;
  assign new_A6715_ = new_A6721_ & new_A6702_;
  assign new_A6714_ = new_A6723_ & new_A6722_;
  assign new_A6713_ = new_A6718_ & new_A6702_;
  assign new_A6712_ = new_A6720_ & new_A6719_;
  assign new_A6711_ = new_A6712_ ^ new_A6702_;
  assign new_A6710_ = new_A6700_ ^ new_A6701_;
  assign A6709 = new_A6710_ & new_A6717_;
  assign A6708 = new_A6710_ & new_A6716_;
  assign A6707 = new_A6715_ | new_A6714_;
  assign A6706 = new_A6713_ | new_A6712_;
  assign A6705 = new_A6711_ & new_A6710_;
  assign new_A6704_ = new_B43_;
  assign new_A6703_ = new_B10_;
  assign new_A6702_ = new_A9976_;
  assign new_A6701_ = new_A9943_;
  assign new_A6700_ = new_A9910_;
  assign new_A6699_ = new_A6677_ & new_A6692_;
  assign new_A6698_ = ~new_A6677_ & ~new_A6699_;
  assign new_A6697_ = new_A6677_ | new_A6692_;
  assign new_A6696_ = ~new_A6670_ | ~new_A6671_;
  assign new_A6695_ = new_A6677_ | new_A6692_;
  assign new_A6694_ = ~new_A6693_ & ~new_A6677_;
  assign new_A6693_ = new_A6677_ & new_A6692_;
  assign new_A6692_ = ~new_A6668_ | ~new_A6669_;
  assign new_A6691_ = new_A6669_ & new_A6681_;
  assign new_A6690_ = new_A6670_ | new_A6677_;
  assign new_A6689_ = new_A6670_ | new_A6671_;
  assign new_A6688_ = ~new_A6698_ | ~new_A6697_;
  assign new_A6687_ = new_A6696_ & new_A6689_;
  assign new_A6686_ = new_A6670_ ^ new_A6677_;
  assign new_A6685_ = ~new_A6694_ | ~new_A6695_;
  assign new_A6684_ = ~new_A6669_ ^ new_A6681_;
  assign new_A6683_ = new_A6691_ | new_A6668_;
  assign new_A6682_ = new_A6688_ & new_A6669_;
  assign new_A6681_ = new_A6690_ & new_A6689_;
  assign new_A6680_ = new_A6685_ & new_A6669_;
  assign new_A6679_ = new_A6687_ & new_A6686_;
  assign new_A6678_ = new_A6679_ ^ new_A6669_;
  assign new_A6677_ = new_A6667_ ^ new_A6668_;
  assign A6676 = new_A6677_ & new_A6684_;
  assign A6675 = new_A6677_ & new_A6683_;
  assign A6674 = new_A6682_ | new_A6681_;
  assign A6673 = new_A6680_ | new_A6679_;
  assign A6672 = new_A6678_ & new_A6677_;
  assign new_A6671_ = new_A9877_;
  assign new_A6670_ = new_A9844_;
  assign new_A6669_ = new_A9811_;
  assign new_A6668_ = new_A9778_;
  assign new_A6667_ = new_A9745_;
  assign new_A6666_ = new_A6644_ & new_A6659_;
  assign new_A6665_ = ~new_A6644_ & ~new_A6666_;
  assign new_A6664_ = new_A6644_ | new_A6659_;
  assign new_A6663_ = ~new_A6637_ | ~new_A6638_;
  assign new_A6662_ = new_A6644_ | new_A6659_;
  assign new_A6661_ = ~new_A6660_ & ~new_A6644_;
  assign new_A6660_ = new_A6644_ & new_A6659_;
  assign new_A6659_ = ~new_A6635_ | ~new_A6636_;
  assign new_A6658_ = new_A6636_ & new_A6648_;
  assign new_A6657_ = new_A6637_ | new_A6644_;
  assign new_A6656_ = new_A6637_ | new_A6638_;
  assign new_A6655_ = ~new_A6665_ | ~new_A6664_;
  assign new_A6654_ = new_A6663_ & new_A6656_;
  assign new_A6653_ = new_A6637_ ^ new_A6644_;
  assign new_A6652_ = ~new_A6661_ | ~new_A6662_;
  assign new_A6651_ = ~new_A6636_ ^ new_A6648_;
  assign new_A6650_ = new_A6658_ | new_A6635_;
  assign new_A6649_ = new_A6655_ & new_A6636_;
  assign new_A6648_ = new_A6657_ & new_A6656_;
  assign new_A6647_ = new_A6652_ & new_A6636_;
  assign new_A6646_ = new_A6654_ & new_A6653_;
  assign new_A6645_ = new_A6646_ ^ new_A6636_;
  assign new_A6644_ = new_A6634_ ^ new_A6635_;
  assign A6643 = new_A6644_ & new_A6651_;
  assign A6642 = new_A6644_ & new_A6650_;
  assign A6641 = new_A6649_ | new_A6648_;
  assign A6640 = new_A6647_ | new_A6646_;
  assign A6639 = new_A6645_ & new_A6644_;
  assign new_A6638_ = new_A9712_;
  assign new_A6637_ = new_A9679_;
  assign new_A6636_ = new_A9646_;
  assign new_A6635_ = new_A9613_;
  assign new_A6634_ = new_A9580_;
  assign new_A6633_ = new_A6611_ & new_A6626_;
  assign new_A6632_ = ~new_A6611_ & ~new_A6633_;
  assign new_A6631_ = new_A6611_ | new_A6626_;
  assign new_A6630_ = ~new_A6604_ | ~new_A6605_;
  assign new_A6629_ = new_A6611_ | new_A6626_;
  assign new_A6628_ = ~new_A6627_ & ~new_A6611_;
  assign new_A6627_ = new_A6611_ & new_A6626_;
  assign new_A6626_ = ~new_A6602_ | ~new_A6603_;
  assign new_A6625_ = new_A6603_ & new_A6615_;
  assign new_A6624_ = new_A6604_ | new_A6611_;
  assign new_A6623_ = new_A6604_ | new_A6605_;
  assign new_A6622_ = ~new_A6632_ | ~new_A6631_;
  assign new_A6621_ = new_A6630_ & new_A6623_;
  assign new_A6620_ = new_A6604_ ^ new_A6611_;
  assign new_A6619_ = ~new_A6628_ | ~new_A6629_;
  assign new_A6618_ = ~new_A6603_ ^ new_A6615_;
  assign new_A6617_ = new_A6625_ | new_A6602_;
  assign new_A6616_ = new_A6622_ & new_A6603_;
  assign new_A6615_ = new_A6624_ & new_A6623_;
  assign new_A6614_ = new_A6619_ & new_A6603_;
  assign new_A6613_ = new_A6621_ & new_A6620_;
  assign new_A6612_ = new_A6613_ ^ new_A6603_;
  assign new_A6611_ = new_A6601_ ^ new_A6602_;
  assign A6610 = new_A6611_ & new_A6618_;
  assign A6609 = new_A6611_ & new_A6617_;
  assign A6608 = new_A6616_ | new_A6615_;
  assign A6607 = new_A6614_ | new_A6613_;
  assign A6606 = new_A6612_ & new_A6611_;
  assign new_A6605_ = new_A9547_;
  assign new_A6604_ = new_A9514_;
  assign new_A6603_ = new_A9481_;
  assign new_A6602_ = new_A9448_;
  assign new_A6601_ = new_A9415_;
  assign new_A6600_ = new_A6578_ & new_A6593_;
  assign new_A6599_ = ~new_A6578_ & ~new_A6600_;
  assign new_A6598_ = new_A6578_ | new_A6593_;
  assign new_A6597_ = ~new_A6571_ | ~new_A6572_;
  assign new_A6596_ = new_A6578_ | new_A6593_;
  assign new_A6595_ = ~new_A6594_ & ~new_A6578_;
  assign new_A6594_ = new_A6578_ & new_A6593_;
  assign new_A6593_ = ~new_A6569_ | ~new_A6570_;
  assign new_A6592_ = new_A6570_ & new_A6582_;
  assign new_A6591_ = new_A6571_ | new_A6578_;
  assign new_A6590_ = new_A6571_ | new_A6572_;
  assign new_A6589_ = ~new_A6599_ | ~new_A6598_;
  assign new_A6588_ = new_A6597_ & new_A6590_;
  assign new_A6587_ = new_A6571_ ^ new_A6578_;
  assign new_A6586_ = ~new_A6595_ | ~new_A6596_;
  assign new_A6585_ = ~new_A6570_ ^ new_A6582_;
  assign new_A6584_ = new_A6592_ | new_A6569_;
  assign new_A6583_ = new_A6589_ & new_A6570_;
  assign new_A6582_ = new_A6591_ & new_A6590_;
  assign new_A6581_ = new_A6586_ & new_A6570_;
  assign new_A6580_ = new_A6588_ & new_A6587_;
  assign new_A6579_ = new_A6580_ ^ new_A6570_;
  assign new_A6578_ = new_A6568_ ^ new_A6569_;
  assign A6577 = new_A6578_ & new_A6585_;
  assign A6576 = new_A6578_ & new_A6584_;
  assign A6575 = new_A6583_ | new_A6582_;
  assign A6574 = new_A6581_ | new_A6580_;
  assign A6573 = new_A6579_ & new_A6578_;
  assign new_A6572_ = new_A9382_;
  assign new_A6571_ = new_A9349_;
  assign new_A6570_ = new_A9316_;
  assign new_A6569_ = new_A9283_;
  assign new_A6568_ = new_A9250_;
  assign new_A6567_ = new_A6545_ & new_A6560_;
  assign new_A6566_ = ~new_A6545_ & ~new_A6567_;
  assign new_A6565_ = new_A6545_ | new_A6560_;
  assign new_A6564_ = ~new_A6538_ | ~new_A6539_;
  assign new_A6563_ = new_A6545_ | new_A6560_;
  assign new_A6562_ = ~new_A6561_ & ~new_A6545_;
  assign new_A6561_ = new_A6545_ & new_A6560_;
  assign new_A6560_ = ~new_A6536_ | ~new_A6537_;
  assign new_A6559_ = new_A6537_ & new_A6549_;
  assign new_A6558_ = new_A6538_ | new_A6545_;
  assign new_A6557_ = new_A6538_ | new_A6539_;
  assign new_A6556_ = ~new_A6566_ | ~new_A6565_;
  assign new_A6555_ = new_A6564_ & new_A6557_;
  assign new_A6554_ = new_A6538_ ^ new_A6545_;
  assign new_A6553_ = ~new_A6562_ | ~new_A6563_;
  assign new_A6552_ = ~new_A6537_ ^ new_A6549_;
  assign new_A6551_ = new_A6559_ | new_A6536_;
  assign new_A6550_ = new_A6556_ & new_A6537_;
  assign new_A6549_ = new_A6558_ & new_A6557_;
  assign new_A6548_ = new_A6553_ & new_A6537_;
  assign new_A6547_ = new_A6555_ & new_A6554_;
  assign new_A6546_ = new_A6547_ ^ new_A6537_;
  assign new_A6545_ = new_A6535_ ^ new_A6536_;
  assign A6544 = new_A6545_ & new_A6552_;
  assign A6543 = new_A6545_ & new_A6551_;
  assign A6542 = new_A6550_ | new_A6549_;
  assign A6541 = new_A6548_ | new_A6547_;
  assign A6540 = new_A6546_ & new_A6545_;
  assign new_A6539_ = new_A9217_;
  assign new_A6538_ = new_A9184_;
  assign new_A6537_ = new_A9151_;
  assign new_A6536_ = new_A9118_;
  assign new_A6535_ = new_A9085_;
  assign new_A6534_ = new_A6512_ & new_A6527_;
  assign new_A6533_ = ~new_A6512_ & ~new_A6534_;
  assign new_A6532_ = new_A6512_ | new_A6527_;
  assign new_A6531_ = ~new_A6505_ | ~new_A6506_;
  assign new_A6530_ = new_A6512_ | new_A6527_;
  assign new_A6529_ = ~new_A6528_ & ~new_A6512_;
  assign new_A6528_ = new_A6512_ & new_A6527_;
  assign new_A6527_ = ~new_A6503_ | ~new_A6504_;
  assign new_A6526_ = new_A6504_ & new_A6516_;
  assign new_A6525_ = new_A6505_ | new_A6512_;
  assign new_A6524_ = new_A6505_ | new_A6506_;
  assign new_A6523_ = ~new_A6533_ | ~new_A6532_;
  assign new_A6522_ = new_A6531_ & new_A6524_;
  assign new_A6521_ = new_A6505_ ^ new_A6512_;
  assign new_A6520_ = ~new_A6529_ | ~new_A6530_;
  assign new_A6519_ = ~new_A6504_ ^ new_A6516_;
  assign new_A6518_ = new_A6526_ | new_A6503_;
  assign new_A6517_ = new_A6523_ & new_A6504_;
  assign new_A6516_ = new_A6525_ & new_A6524_;
  assign new_A6515_ = new_A6520_ & new_A6504_;
  assign new_A6514_ = new_A6522_ & new_A6521_;
  assign new_A6513_ = new_A6514_ ^ new_A6504_;
  assign new_A6512_ = new_A6502_ ^ new_A6503_;
  assign A6511 = new_A6512_ & new_A6519_;
  assign A6510 = new_A6512_ & new_A6518_;
  assign A6509 = new_A6517_ | new_A6516_;
  assign A6508 = new_A6515_ | new_A6514_;
  assign A6507 = new_A6513_ & new_A6512_;
  assign new_A6506_ = new_A9052_;
  assign new_A6505_ = new_A9019_;
  assign new_A6504_ = new_A8986_;
  assign new_A6503_ = new_A8953_;
  assign new_A6502_ = new_A8920_;
  assign new_A6501_ = new_A6479_ & new_A6494_;
  assign new_A6500_ = ~new_A6479_ & ~new_A6501_;
  assign new_A6499_ = new_A6479_ | new_A6494_;
  assign new_A6498_ = ~new_A6472_ | ~new_A6473_;
  assign new_A6497_ = new_A6479_ | new_A6494_;
  assign new_A6496_ = ~new_A6495_ & ~new_A6479_;
  assign new_A6495_ = new_A6479_ & new_A6494_;
  assign new_A6494_ = ~new_A6470_ | ~new_A6471_;
  assign new_A6493_ = new_A6471_ & new_A6483_;
  assign new_A6492_ = new_A6472_ | new_A6479_;
  assign new_A6491_ = new_A6472_ | new_A6473_;
  assign new_A6490_ = ~new_A6500_ | ~new_A6499_;
  assign new_A6489_ = new_A6498_ & new_A6491_;
  assign new_A6488_ = new_A6472_ ^ new_A6479_;
  assign new_A6487_ = ~new_A6496_ | ~new_A6497_;
  assign new_A6486_ = ~new_A6471_ ^ new_A6483_;
  assign new_A6485_ = new_A6493_ | new_A6470_;
  assign new_A6484_ = new_A6490_ & new_A6471_;
  assign new_A6483_ = new_A6492_ & new_A6491_;
  assign new_A6482_ = new_A6487_ & new_A6471_;
  assign new_A6481_ = new_A6489_ & new_A6488_;
  assign new_A6480_ = new_A6481_ ^ new_A6471_;
  assign new_A6479_ = new_A6469_ ^ new_A6470_;
  assign A6478 = new_A6479_ & new_A6486_;
  assign A6477 = new_A6479_ & new_A6485_;
  assign A6476 = new_A6484_ | new_A6483_;
  assign A6475 = new_A6482_ | new_A6481_;
  assign A6474 = new_A6480_ & new_A6479_;
  assign new_A6473_ = new_A8887_;
  assign new_A6472_ = new_A8854_;
  assign new_A6471_ = new_A8821_;
  assign new_A6470_ = new_A8788_;
  assign new_A6469_ = new_A8755_;
  assign new_A6468_ = new_A6446_ & new_A6461_;
  assign new_A6467_ = ~new_A6446_ & ~new_A6468_;
  assign new_A6466_ = new_A6446_ | new_A6461_;
  assign new_A6465_ = ~new_A6439_ | ~new_A6440_;
  assign new_A6464_ = new_A6446_ | new_A6461_;
  assign new_A6463_ = ~new_A6462_ & ~new_A6446_;
  assign new_A6462_ = new_A6446_ & new_A6461_;
  assign new_A6461_ = ~new_A6437_ | ~new_A6438_;
  assign new_A6460_ = new_A6438_ & new_A6450_;
  assign new_A6459_ = new_A6439_ | new_A6446_;
  assign new_A6458_ = new_A6439_ | new_A6440_;
  assign new_A6457_ = ~new_A6467_ | ~new_A6466_;
  assign new_A6456_ = new_A6465_ & new_A6458_;
  assign new_A6455_ = new_A6439_ ^ new_A6446_;
  assign new_A6454_ = ~new_A6463_ | ~new_A6464_;
  assign new_A6453_ = ~new_A6438_ ^ new_A6450_;
  assign new_A6452_ = new_A6460_ | new_A6437_;
  assign new_A6451_ = new_A6457_ & new_A6438_;
  assign new_A6450_ = new_A6459_ & new_A6458_;
  assign new_A6449_ = new_A6454_ & new_A6438_;
  assign new_A6448_ = new_A6456_ & new_A6455_;
  assign new_A6447_ = new_A6448_ ^ new_A6438_;
  assign new_A6446_ = new_A6436_ ^ new_A6437_;
  assign A6445 = new_A6446_ & new_A6453_;
  assign A6444 = new_A6446_ & new_A6452_;
  assign A6443 = new_A6451_ | new_A6450_;
  assign A6442 = new_A6449_ | new_A6448_;
  assign A6441 = new_A6447_ & new_A6446_;
  assign new_A6440_ = new_A8722_;
  assign new_A6439_ = new_A8689_;
  assign new_A6438_ = new_A8656_;
  assign new_A6437_ = new_A8623_;
  assign new_A6436_ = new_A8590_;
  assign new_A6435_ = new_A6413_ & new_A6428_;
  assign new_A6434_ = ~new_A6413_ & ~new_A6435_;
  assign new_A6433_ = new_A6413_ | new_A6428_;
  assign new_A6432_ = ~new_A6406_ | ~new_A6407_;
  assign new_A6431_ = new_A6413_ | new_A6428_;
  assign new_A6430_ = ~new_A6429_ & ~new_A6413_;
  assign new_A6429_ = new_A6413_ & new_A6428_;
  assign new_A6428_ = ~new_A6404_ | ~new_A6405_;
  assign new_A6427_ = new_A6405_ & new_A6417_;
  assign new_A6426_ = new_A6406_ | new_A6413_;
  assign new_A6425_ = new_A6406_ | new_A6407_;
  assign new_A6424_ = ~new_A6434_ | ~new_A6433_;
  assign new_A6423_ = new_A6432_ & new_A6425_;
  assign new_A6422_ = new_A6406_ ^ new_A6413_;
  assign new_A6421_ = ~new_A6430_ | ~new_A6431_;
  assign new_A6420_ = ~new_A6405_ ^ new_A6417_;
  assign new_A6419_ = new_A6427_ | new_A6404_;
  assign new_A6418_ = new_A6424_ & new_A6405_;
  assign new_A6417_ = new_A6426_ & new_A6425_;
  assign new_A6416_ = new_A6421_ & new_A6405_;
  assign new_A6415_ = new_A6423_ & new_A6422_;
  assign new_A6414_ = new_A6415_ ^ new_A6405_;
  assign new_A6413_ = new_A6403_ ^ new_A6404_;
  assign A6412 = new_A6413_ & new_A6420_;
  assign A6411 = new_A6413_ & new_A6419_;
  assign A6410 = new_A6418_ | new_A6417_;
  assign A6409 = new_A6416_ | new_A6415_;
  assign A6408 = new_A6414_ & new_A6413_;
  assign new_A6407_ = new_A8557_;
  assign new_A6406_ = new_A8524_;
  assign new_A6405_ = new_A8491_;
  assign new_A6404_ = new_A8458_;
  assign new_A6403_ = new_A8425_;
  assign new_A6402_ = new_A6380_ & new_A6395_;
  assign new_A6401_ = ~new_A6380_ & ~new_A6402_;
  assign new_A6400_ = new_A6380_ | new_A6395_;
  assign new_A6399_ = ~new_A6373_ | ~new_A6374_;
  assign new_A6398_ = new_A6380_ | new_A6395_;
  assign new_A6397_ = ~new_A6396_ & ~new_A6380_;
  assign new_A6396_ = new_A6380_ & new_A6395_;
  assign new_A6395_ = ~new_A6371_ | ~new_A6372_;
  assign new_A6394_ = new_A6372_ & new_A6384_;
  assign new_A6393_ = new_A6373_ | new_A6380_;
  assign new_A6392_ = new_A6373_ | new_A6374_;
  assign new_A6391_ = ~new_A6401_ | ~new_A6400_;
  assign new_A6390_ = new_A6399_ & new_A6392_;
  assign new_A6389_ = new_A6373_ ^ new_A6380_;
  assign new_A6388_ = ~new_A6397_ | ~new_A6398_;
  assign new_A6387_ = ~new_A6372_ ^ new_A6384_;
  assign new_A6386_ = new_A6394_ | new_A6371_;
  assign new_A6385_ = new_A6391_ & new_A6372_;
  assign new_A6384_ = new_A6393_ & new_A6392_;
  assign new_A6383_ = new_A6388_ & new_A6372_;
  assign new_A6382_ = new_A6390_ & new_A6389_;
  assign new_A6381_ = new_A6382_ ^ new_A6372_;
  assign new_A6380_ = new_A6370_ ^ new_A6371_;
  assign A6379 = new_A6380_ & new_A6387_;
  assign A6378 = new_A6380_ & new_A6386_;
  assign A6377 = new_A6385_ | new_A6384_;
  assign A6376 = new_A6383_ | new_A6382_;
  assign A6375 = new_A6381_ & new_A6380_;
  assign new_A6374_ = new_A8392_;
  assign new_A6373_ = new_A8359_;
  assign new_A6372_ = new_A8326_;
  assign new_A6371_ = new_A8293_;
  assign new_A6370_ = new_A8260_;
  assign new_A6369_ = new_A6347_ & new_A6362_;
  assign new_A6368_ = ~new_A6347_ & ~new_A6369_;
  assign new_A6367_ = new_A6347_ | new_A6362_;
  assign new_A6366_ = ~new_A6340_ | ~new_A6341_;
  assign new_A6365_ = new_A6347_ | new_A6362_;
  assign new_A6364_ = ~new_A6363_ & ~new_A6347_;
  assign new_A6363_ = new_A6347_ & new_A6362_;
  assign new_A6362_ = ~new_A6338_ | ~new_A6339_;
  assign new_A6361_ = new_A6339_ & new_A6351_;
  assign new_A6360_ = new_A6340_ | new_A6347_;
  assign new_A6359_ = new_A6340_ | new_A6341_;
  assign new_A6358_ = ~new_A6368_ | ~new_A6367_;
  assign new_A6357_ = new_A6366_ & new_A6359_;
  assign new_A6356_ = new_A6340_ ^ new_A6347_;
  assign new_A6355_ = ~new_A6364_ | ~new_A6365_;
  assign new_A6354_ = ~new_A6339_ ^ new_A6351_;
  assign new_A6353_ = new_A6361_ | new_A6338_;
  assign new_A6352_ = new_A6358_ & new_A6339_;
  assign new_A6351_ = new_A6360_ & new_A6359_;
  assign new_A6350_ = new_A6355_ & new_A6339_;
  assign new_A6349_ = new_A6357_ & new_A6356_;
  assign new_A6348_ = new_A6349_ ^ new_A6339_;
  assign new_A6347_ = new_A6337_ ^ new_A6338_;
  assign A6346 = new_A6347_ & new_A6354_;
  assign A6345 = new_A6347_ & new_A6353_;
  assign A6344 = new_A6352_ | new_A6351_;
  assign A6343 = new_A6350_ | new_A6349_;
  assign A6342 = new_A6348_ & new_A6347_;
  assign new_A6341_ = new_A8227_;
  assign new_A6340_ = new_A8194_;
  assign new_A6339_ = new_A8161_;
  assign new_A6338_ = new_A8128_;
  assign new_A6337_ = new_A8095_;
  assign new_A6336_ = new_A6314_ & new_A6329_;
  assign new_A6335_ = ~new_A6314_ & ~new_A6336_;
  assign new_A6334_ = new_A6314_ | new_A6329_;
  assign new_A6333_ = ~new_A6307_ | ~new_A6308_;
  assign new_A6332_ = new_A6314_ | new_A6329_;
  assign new_A6331_ = ~new_A6330_ & ~new_A6314_;
  assign new_A6330_ = new_A6314_ & new_A6329_;
  assign new_A6329_ = ~new_A6305_ | ~new_A6306_;
  assign new_A6328_ = new_A6306_ & new_A6318_;
  assign new_A6327_ = new_A6307_ | new_A6314_;
  assign new_A6326_ = new_A6307_ | new_A6308_;
  assign new_A6325_ = ~new_A6335_ | ~new_A6334_;
  assign new_A6324_ = new_A6333_ & new_A6326_;
  assign new_A6323_ = new_A6307_ ^ new_A6314_;
  assign new_A6322_ = ~new_A6331_ | ~new_A6332_;
  assign new_A6321_ = ~new_A6306_ ^ new_A6318_;
  assign new_A6320_ = new_A6328_ | new_A6305_;
  assign new_A6319_ = new_A6325_ & new_A6306_;
  assign new_A6318_ = new_A6327_ & new_A6326_;
  assign new_A6317_ = new_A6322_ & new_A6306_;
  assign new_A6316_ = new_A6324_ & new_A6323_;
  assign new_A6315_ = new_A6316_ ^ new_A6306_;
  assign new_A6314_ = new_A6304_ ^ new_A6305_;
  assign A6313 = new_A6314_ & new_A6321_;
  assign A6312 = new_A6314_ & new_A6320_;
  assign A6311 = new_A6319_ | new_A6318_;
  assign A6310 = new_A6317_ | new_A6316_;
  assign A6309 = new_A6315_ & new_A6314_;
  assign new_A6308_ = new_A8062_;
  assign new_A6307_ = new_A8029_;
  assign new_A6306_ = new_A7996_;
  assign new_A6305_ = new_A7963_;
  assign new_A6304_ = new_A7930_;
  assign new_A6303_ = new_A6281_ & new_A6296_;
  assign new_A6302_ = ~new_A6281_ & ~new_A6303_;
  assign new_A6301_ = new_A6281_ | new_A6296_;
  assign new_A6300_ = ~new_A6274_ | ~new_A6275_;
  assign new_A6299_ = new_A6281_ | new_A6296_;
  assign new_A6298_ = ~new_A6297_ & ~new_A6281_;
  assign new_A6297_ = new_A6281_ & new_A6296_;
  assign new_A6296_ = ~new_A6272_ | ~new_A6273_;
  assign new_A6295_ = new_A6273_ & new_A6285_;
  assign new_A6294_ = new_A6274_ | new_A6281_;
  assign new_A6293_ = new_A6274_ | new_A6275_;
  assign new_A6292_ = ~new_A6302_ | ~new_A6301_;
  assign new_A6291_ = new_A6300_ & new_A6293_;
  assign new_A6290_ = new_A6274_ ^ new_A6281_;
  assign new_A6289_ = ~new_A6298_ | ~new_A6299_;
  assign new_A6288_ = ~new_A6273_ ^ new_A6285_;
  assign new_A6287_ = new_A6295_ | new_A6272_;
  assign new_A6286_ = new_A6292_ & new_A6273_;
  assign new_A6285_ = new_A6294_ & new_A6293_;
  assign new_A6284_ = new_A6289_ & new_A6273_;
  assign new_A6283_ = new_A6291_ & new_A6290_;
  assign new_A6282_ = new_A6283_ ^ new_A6273_;
  assign new_A6281_ = new_A6271_ ^ new_A6272_;
  assign A6280 = new_A6281_ & new_A6288_;
  assign A6279 = new_A6281_ & new_A6287_;
  assign A6278 = new_A6286_ | new_A6285_;
  assign A6277 = new_A6284_ | new_A6283_;
  assign A6276 = new_A6282_ & new_A6281_;
  assign new_A6275_ = new_A7897_;
  assign new_A6274_ = new_A7864_;
  assign new_A6273_ = new_A7831_;
  assign new_A6272_ = new_A7798_;
  assign new_A6271_ = new_A7765_;
  assign new_A6270_ = new_A6248_ & new_A6263_;
  assign new_A6269_ = ~new_A6248_ & ~new_A6270_;
  assign new_A6268_ = new_A6248_ | new_A6263_;
  assign new_A6267_ = ~new_A6241_ | ~new_A6242_;
  assign new_A6266_ = new_A6248_ | new_A6263_;
  assign new_A6265_ = ~new_A6264_ & ~new_A6248_;
  assign new_A6264_ = new_A6248_ & new_A6263_;
  assign new_A6263_ = ~new_A6239_ | ~new_A6240_;
  assign new_A6262_ = new_A6240_ & new_A6252_;
  assign new_A6261_ = new_A6241_ | new_A6248_;
  assign new_A6260_ = new_A6241_ | new_A6242_;
  assign new_A6259_ = ~new_A6269_ | ~new_A6268_;
  assign new_A6258_ = new_A6267_ & new_A6260_;
  assign new_A6257_ = new_A6241_ ^ new_A6248_;
  assign new_A6256_ = ~new_A6265_ | ~new_A6266_;
  assign new_A6255_ = ~new_A6240_ ^ new_A6252_;
  assign new_A6254_ = new_A6262_ | new_A6239_;
  assign new_A6253_ = new_A6259_ & new_A6240_;
  assign new_A6252_ = new_A6261_ & new_A6260_;
  assign new_A6251_ = new_A6256_ & new_A6240_;
  assign new_A6250_ = new_A6258_ & new_A6257_;
  assign new_A6249_ = new_A6250_ ^ new_A6240_;
  assign new_A6248_ = new_A6238_ ^ new_A6239_;
  assign A6247 = new_A6248_ & new_A6255_;
  assign A6246 = new_A6248_ & new_A6254_;
  assign A6245 = new_A6253_ | new_A6252_;
  assign A6244 = new_A6251_ | new_A6250_;
  assign A6243 = new_A6249_ & new_A6248_;
  assign new_A6242_ = new_A7732_;
  assign new_A6241_ = new_A7699_;
  assign new_A6240_ = new_A7666_;
  assign new_A6239_ = new_A7633_;
  assign new_A6238_ = new_A7600_;
  assign new_A6237_ = new_A6215_ & new_A6230_;
  assign new_A6236_ = ~new_A6215_ & ~new_A6237_;
  assign new_A6235_ = new_A6215_ | new_A6230_;
  assign new_A6234_ = ~new_A6208_ | ~new_A6209_;
  assign new_A6233_ = new_A6215_ | new_A6230_;
  assign new_A6232_ = ~new_A6231_ & ~new_A6215_;
  assign new_A6231_ = new_A6215_ & new_A6230_;
  assign new_A6230_ = ~new_A6206_ | ~new_A6207_;
  assign new_A6229_ = new_A6207_ & new_A6219_;
  assign new_A6228_ = new_A6208_ | new_A6215_;
  assign new_A6227_ = new_A6208_ | new_A6209_;
  assign new_A6226_ = ~new_A6236_ | ~new_A6235_;
  assign new_A6225_ = new_A6234_ & new_A6227_;
  assign new_A6224_ = new_A6208_ ^ new_A6215_;
  assign new_A6223_ = ~new_A6232_ | ~new_A6233_;
  assign new_A6222_ = ~new_A6207_ ^ new_A6219_;
  assign new_A6221_ = new_A6229_ | new_A6206_;
  assign new_A6220_ = new_A6226_ & new_A6207_;
  assign new_A6219_ = new_A6228_ & new_A6227_;
  assign new_A6218_ = new_A6223_ & new_A6207_;
  assign new_A6217_ = new_A6225_ & new_A6224_;
  assign new_A6216_ = new_A6217_ ^ new_A6207_;
  assign new_A6215_ = new_A6205_ ^ new_A6206_;
  assign A6214 = new_A6215_ & new_A6222_;
  assign A6213 = new_A6215_ & new_A6221_;
  assign A6212 = new_A6220_ | new_A6219_;
  assign A6211 = new_A6218_ | new_A6217_;
  assign A6210 = new_A6216_ & new_A6215_;
  assign new_A6209_ = new_A7567_;
  assign new_A6208_ = new_A7534_;
  assign new_A6207_ = new_A7501_;
  assign new_A6206_ = new_A7468_;
  assign new_A6205_ = new_A7435_;
  assign new_A6204_ = new_A6182_ & new_A6197_;
  assign new_A6203_ = ~new_A6182_ & ~new_A6204_;
  assign new_A6202_ = new_A6182_ | new_A6197_;
  assign new_A6201_ = ~new_A6175_ | ~new_A6176_;
  assign new_A6200_ = new_A6182_ | new_A6197_;
  assign new_A6199_ = ~new_A6198_ & ~new_A6182_;
  assign new_A6198_ = new_A6182_ & new_A6197_;
  assign new_A6197_ = ~new_A6173_ | ~new_A6174_;
  assign new_A6196_ = new_A6174_ & new_A6186_;
  assign new_A6195_ = new_A6175_ | new_A6182_;
  assign new_A6194_ = new_A6175_ | new_A6176_;
  assign new_A6193_ = ~new_A6203_ | ~new_A6202_;
  assign new_A6192_ = new_A6201_ & new_A6194_;
  assign new_A6191_ = new_A6175_ ^ new_A6182_;
  assign new_A6190_ = ~new_A6199_ | ~new_A6200_;
  assign new_A6189_ = ~new_A6174_ ^ new_A6186_;
  assign new_A6188_ = new_A6196_ | new_A6173_;
  assign new_A6187_ = new_A6193_ & new_A6174_;
  assign new_A6186_ = new_A6195_ & new_A6194_;
  assign new_A6185_ = new_A6190_ & new_A6174_;
  assign new_A6184_ = new_A6192_ & new_A6191_;
  assign new_A6183_ = new_A6184_ ^ new_A6174_;
  assign new_A6182_ = new_A6172_ ^ new_A6173_;
  assign A6181 = new_A6182_ & new_A6189_;
  assign A6180 = new_A6182_ & new_A6188_;
  assign A6179 = new_A6187_ | new_A6186_;
  assign A6178 = new_A6185_ | new_A6184_;
  assign A6177 = new_A6183_ & new_A6182_;
  assign new_A6176_ = new_A7402_;
  assign new_A6175_ = new_A7369_;
  assign new_A6174_ = new_A7336_;
  assign new_A6173_ = new_A7303_;
  assign new_A6172_ = new_A7270_;
  assign new_A6171_ = new_A6149_ & new_A6164_;
  assign new_A6170_ = ~new_A6149_ & ~new_A6171_;
  assign new_A6169_ = new_A6149_ | new_A6164_;
  assign new_A6168_ = ~new_A6142_ | ~new_A6143_;
  assign new_A6167_ = new_A6149_ | new_A6164_;
  assign new_A6166_ = ~new_A6165_ & ~new_A6149_;
  assign new_A6165_ = new_A6149_ & new_A6164_;
  assign new_A6164_ = ~new_A6140_ | ~new_A6141_;
  assign new_A6163_ = new_A6141_ & new_A6153_;
  assign new_A6162_ = new_A6142_ | new_A6149_;
  assign new_A6161_ = new_A6142_ | new_A6143_;
  assign new_A6160_ = ~new_A6170_ | ~new_A6169_;
  assign new_A6159_ = new_A6168_ & new_A6161_;
  assign new_A6158_ = new_A6142_ ^ new_A6149_;
  assign new_A6157_ = ~new_A6166_ | ~new_A6167_;
  assign new_A6156_ = ~new_A6141_ ^ new_A6153_;
  assign new_A6155_ = new_A6163_ | new_A6140_;
  assign new_A6154_ = new_A6160_ & new_A6141_;
  assign new_A6153_ = new_A6162_ & new_A6161_;
  assign new_A6152_ = new_A6157_ & new_A6141_;
  assign new_A6151_ = new_A6159_ & new_A6158_;
  assign new_A6150_ = new_A6151_ ^ new_A6141_;
  assign new_A6149_ = new_A6139_ ^ new_A6140_;
  assign A6148 = new_A6149_ & new_A6156_;
  assign A6147 = new_A6149_ & new_A6155_;
  assign A6146 = new_A6154_ | new_A6153_;
  assign A6145 = new_A6152_ | new_A6151_;
  assign A6144 = new_A6150_ & new_A6149_;
  assign new_A6143_ = new_A7237_;
  assign new_A6142_ = new_A7204_;
  assign new_A6141_ = new_A7171_;
  assign new_A6140_ = new_A7138_;
  assign new_A6139_ = new_A7105_;
  assign new_A6138_ = new_A6116_ & new_A6131_;
  assign new_A6137_ = ~new_A6116_ & ~new_A6138_;
  assign new_A6136_ = new_A6116_ | new_A6131_;
  assign new_A6135_ = ~new_A6109_ | ~new_A6110_;
  assign new_A6134_ = new_A6116_ | new_A6131_;
  assign new_A6133_ = ~new_A6132_ & ~new_A6116_;
  assign new_A6132_ = new_A6116_ & new_A6131_;
  assign new_A6131_ = ~new_A6107_ | ~new_A6108_;
  assign new_A6130_ = new_A6108_ & new_A6120_;
  assign new_A6129_ = new_A6109_ | new_A6116_;
  assign new_A6128_ = new_A6109_ | new_A6110_;
  assign new_A6127_ = ~new_A6137_ | ~new_A6136_;
  assign new_A6126_ = new_A6135_ & new_A6128_;
  assign new_A6125_ = new_A6109_ ^ new_A6116_;
  assign new_A6124_ = ~new_A6133_ | ~new_A6134_;
  assign new_A6123_ = ~new_A6108_ ^ new_A6120_;
  assign new_A6122_ = new_A6130_ | new_A6107_;
  assign new_A6121_ = new_A6127_ & new_A6108_;
  assign new_A6120_ = new_A6129_ & new_A6128_;
  assign new_A6119_ = new_A6124_ & new_A6108_;
  assign new_A6118_ = new_A6126_ & new_A6125_;
  assign new_A6117_ = new_A6118_ ^ new_A6108_;
  assign new_A6116_ = new_A6106_ ^ new_A6107_;
  assign A6115 = new_A6116_ & new_A6123_;
  assign A6114 = new_A6116_ & new_A6122_;
  assign A6113 = new_A6121_ | new_A6120_;
  assign A6112 = new_A6119_ | new_A6118_;
  assign A6111 = new_A6117_ & new_A6116_;
  assign new_A6110_ = new_A7072_;
  assign new_A6109_ = new_A7039_;
  assign new_A6108_ = new_A7006_;
  assign new_A6107_ = new_A6973_;
  assign new_A6106_ = new_A6936_;
  assign new_A6105_ = new_A6083_ & new_A6098_;
  assign new_A6104_ = ~new_A6083_ & ~new_A6105_;
  assign new_A6103_ = new_A6083_ | new_A6098_;
  assign new_A6102_ = ~new_A6076_ | ~new_A6077_;
  assign new_A6101_ = new_A6083_ | new_A6098_;
  assign new_A6100_ = ~new_A6099_ & ~new_A6083_;
  assign new_A6099_ = new_A6083_ & new_A6098_;
  assign new_A6098_ = ~new_A6074_ | ~new_A6075_;
  assign new_A6097_ = new_A6075_ & new_A6087_;
  assign new_A6096_ = new_A6076_ | new_A6083_;
  assign new_A6095_ = new_A6076_ | new_A6077_;
  assign new_A6094_ = ~new_A6104_ | ~new_A6103_;
  assign new_A6093_ = new_A6102_ & new_A6095_;
  assign new_A6092_ = new_A6076_ ^ new_A6083_;
  assign new_A6091_ = ~new_A6100_ | ~new_A6101_;
  assign new_A6090_ = ~new_A6075_ ^ new_A6087_;
  assign new_A6089_ = new_A6097_ | new_A6074_;
  assign new_A6088_ = new_A6094_ & new_A6075_;
  assign new_A6087_ = new_A6096_ & new_A6095_;
  assign new_A6086_ = new_A6091_ & new_A6075_;
  assign new_A6085_ = new_A6093_ & new_A6092_;
  assign new_A6084_ = new_A6085_ ^ new_A6075_;
  assign new_A6083_ = new_A6073_ ^ new_A6074_;
  assign A6082 = new_A6083_ & new_A6090_;
  assign A6081 = new_A6083_ & new_A6089_;
  assign A6080 = new_A6088_ | new_A6087_;
  assign A6079 = new_A6086_ | new_A6085_;
  assign A6078 = new_A6084_ & new_A6083_;
  assign new_A6077_ = new_B1032_;
  assign new_A6076_ = new_B999_;
  assign new_A6075_ = new_B966_;
  assign new_A6074_ = new_B933_;
  assign new_A6073_ = new_B900_;
  assign new_A6072_ = new_A6050_ & new_A6065_;
  assign new_A6071_ = ~new_A6050_ & ~new_A6072_;
  assign new_A6070_ = new_A6050_ | new_A6065_;
  assign new_A6069_ = ~new_A6043_ | ~new_A6044_;
  assign new_A6068_ = new_A6050_ | new_A6065_;
  assign new_A6067_ = ~new_A6066_ & ~new_A6050_;
  assign new_A6066_ = new_A6050_ & new_A6065_;
  assign new_A6065_ = ~new_A6041_ | ~new_A6042_;
  assign new_A6064_ = new_A6042_ & new_A6054_;
  assign new_A6063_ = new_A6043_ | new_A6050_;
  assign new_A6062_ = new_A6043_ | new_A6044_;
  assign new_A6061_ = ~new_A6071_ | ~new_A6070_;
  assign new_A6060_ = new_A6069_ & new_A6062_;
  assign new_A6059_ = new_A6043_ ^ new_A6050_;
  assign new_A6058_ = ~new_A6067_ | ~new_A6068_;
  assign new_A6057_ = ~new_A6042_ ^ new_A6054_;
  assign new_A6056_ = new_A6064_ | new_A6041_;
  assign new_A6055_ = new_A6061_ & new_A6042_;
  assign new_A6054_ = new_A6063_ & new_A6062_;
  assign new_A6053_ = new_A6058_ & new_A6042_;
  assign new_A6052_ = new_A6060_ & new_A6059_;
  assign new_A6051_ = new_A6052_ ^ new_A6042_;
  assign new_A6050_ = new_A6040_ ^ new_A6041_;
  assign A6049 = new_A6050_ & new_A6057_;
  assign A6048 = new_A6050_ & new_A6056_;
  assign A6047 = new_A6055_ | new_A6054_;
  assign A6046 = new_A6053_ | new_A6052_;
  assign A6045 = new_A6051_ & new_A6050_;
  assign new_A6044_ = new_B867_;
  assign new_A6043_ = new_B834_;
  assign new_A6042_ = new_B801_;
  assign new_A6041_ = new_B768_;
  assign new_A6040_ = new_B735_;
  assign new_A6039_ = new_A6017_ & new_A6032_;
  assign new_A6038_ = ~new_A6017_ & ~new_A6039_;
  assign new_A6037_ = new_A6017_ | new_A6032_;
  assign new_A6036_ = ~new_A6010_ | ~new_A6011_;
  assign new_A6035_ = new_A6017_ | new_A6032_;
  assign new_A6034_ = ~new_A6033_ & ~new_A6017_;
  assign new_A6033_ = new_A6017_ & new_A6032_;
  assign new_A6032_ = ~new_A6008_ | ~new_A6009_;
  assign new_A6031_ = new_A6009_ & new_A6021_;
  assign new_A6030_ = new_A6010_ | new_A6017_;
  assign new_A6029_ = new_A6010_ | new_A6011_;
  assign new_A6028_ = ~new_A6038_ | ~new_A6037_;
  assign new_A6027_ = new_A6036_ & new_A6029_;
  assign new_A6026_ = new_A6010_ ^ new_A6017_;
  assign new_A6025_ = ~new_A6034_ | ~new_A6035_;
  assign new_A6024_ = ~new_A6009_ ^ new_A6021_;
  assign new_A6023_ = new_A6031_ | new_A6008_;
  assign new_A6022_ = new_A6028_ & new_A6009_;
  assign new_A6021_ = new_A6030_ & new_A6029_;
  assign new_A6020_ = new_A6025_ & new_A6009_;
  assign new_A6019_ = new_A6027_ & new_A6026_;
  assign new_A6018_ = new_A6019_ ^ new_A6009_;
  assign new_A6017_ = new_A6007_ ^ new_A6008_;
  assign A6016 = new_A6017_ & new_A6024_;
  assign A6015 = new_A6017_ & new_A6023_;
  assign A6014 = new_A6022_ | new_A6021_;
  assign A6013 = new_A6020_ | new_A6019_;
  assign A6012 = new_A6018_ & new_A6017_;
  assign new_A6011_ = new_B702_;
  assign new_A6010_ = new_B669_;
  assign new_A6009_ = new_B636_;
  assign new_A6008_ = new_B603_;
  assign new_A6007_ = new_B570_;
  assign new_A6006_ = new_A5984_ & new_A5999_;
  assign new_A6005_ = ~new_A5984_ & ~new_A6006_;
  assign new_A6004_ = new_A5984_ | new_A5999_;
  assign new_A6003_ = ~new_A5977_ | ~new_A5978_;
  assign new_A6002_ = new_A5984_ | new_A5999_;
  assign new_A6001_ = ~new_A6000_ & ~new_A5984_;
  assign new_A6000_ = new_A5984_ & new_A5999_;
  assign new_A5999_ = ~new_A5975_ | ~new_A5976_;
  assign new_A5998_ = new_A5976_ & new_A5988_;
  assign new_A5997_ = new_A5977_ | new_A5984_;
  assign new_A5996_ = new_A5977_ | new_A5978_;
  assign new_A5995_ = ~new_A6005_ | ~new_A6004_;
  assign new_A5994_ = new_A6003_ & new_A5996_;
  assign new_A5993_ = new_A5977_ ^ new_A5984_;
  assign new_A5992_ = ~new_A6001_ | ~new_A6002_;
  assign new_A5991_ = ~new_A5976_ ^ new_A5988_;
  assign new_A5990_ = new_A5998_ | new_A5975_;
  assign new_A5989_ = new_A5995_ & new_A5976_;
  assign new_A5988_ = new_A5997_ & new_A5996_;
  assign new_A5987_ = new_A5992_ & new_A5976_;
  assign new_A5986_ = new_A5994_ & new_A5993_;
  assign new_A5985_ = new_A5986_ ^ new_A5976_;
  assign new_A5984_ = new_A5974_ ^ new_A5975_;
  assign A5983 = new_A5984_ & new_A5991_;
  assign A5982 = new_A5984_ & new_A5990_;
  assign A5981 = new_A5989_ | new_A5988_;
  assign A5980 = new_A5987_ | new_A5986_;
  assign A5979 = new_A5985_ & new_A5984_;
  assign new_A5978_ = new_B537_;
  assign new_A5977_ = new_B504_;
  assign new_A5976_ = new_B471_;
  assign new_A5975_ = new_B438_;
  assign new_A5974_ = new_B405_;
  assign new_A5973_ = new_A5951_ & new_A5966_;
  assign new_A5972_ = ~new_A5951_ & ~new_A5973_;
  assign new_A5971_ = new_A5951_ | new_A5966_;
  assign new_A5970_ = ~new_A5944_ | ~new_A5945_;
  assign new_A5969_ = new_A5951_ | new_A5966_;
  assign new_A5968_ = ~new_A5967_ & ~new_A5951_;
  assign new_A5967_ = new_A5951_ & new_A5966_;
  assign new_A5966_ = ~new_A5942_ | ~new_A5943_;
  assign new_A5965_ = new_A5943_ & new_A5955_;
  assign new_A5964_ = new_A5944_ | new_A5951_;
  assign new_A5963_ = new_A5944_ | new_A5945_;
  assign new_A5962_ = ~new_A5972_ | ~new_A5971_;
  assign new_A5961_ = new_A5970_ & new_A5963_;
  assign new_A5960_ = new_A5944_ ^ new_A5951_;
  assign new_A5959_ = ~new_A5968_ | ~new_A5969_;
  assign new_A5958_ = ~new_A5943_ ^ new_A5955_;
  assign new_A5957_ = new_A5965_ | new_A5942_;
  assign new_A5956_ = new_A5962_ & new_A5943_;
  assign new_A5955_ = new_A5964_ & new_A5963_;
  assign new_A5954_ = new_A5959_ & new_A5943_;
  assign new_A5953_ = new_A5961_ & new_A5960_;
  assign new_A5952_ = new_A5953_ ^ new_A5943_;
  assign new_A5951_ = new_A5941_ ^ new_A5942_;
  assign A5950 = new_A5951_ & new_A5958_;
  assign A5949 = new_A5951_ & new_A5957_;
  assign A5948 = new_A5956_ | new_A5955_;
  assign A5947 = new_A5954_ | new_A5953_;
  assign A5946 = new_A5952_ & new_A5951_;
  assign new_A5945_ = new_B372_;
  assign new_A5944_ = new_B339_;
  assign new_A5943_ = new_B306_;
  assign new_A5942_ = new_B273_;
  assign new_A5941_ = new_B240_;
  assign new_A5940_ = new_A5918_ & new_A5933_;
  assign new_A5939_ = ~new_A5918_ & ~new_A5940_;
  assign new_A5938_ = new_A5918_ | new_A5933_;
  assign new_A5937_ = ~new_A5911_ | ~new_A5912_;
  assign new_A5936_ = new_A5918_ | new_A5933_;
  assign new_A5935_ = ~new_A5934_ & ~new_A5918_;
  assign new_A5934_ = new_A5918_ & new_A5933_;
  assign new_A5933_ = ~new_A5909_ | ~new_A5910_;
  assign new_A5932_ = new_A5910_ & new_A5922_;
  assign new_A5931_ = new_A5911_ | new_A5918_;
  assign new_A5930_ = new_A5911_ | new_A5912_;
  assign new_A5929_ = ~new_A5939_ | ~new_A5938_;
  assign new_A5928_ = new_A5937_ & new_A5930_;
  assign new_A5927_ = new_A5911_ ^ new_A5918_;
  assign new_A5926_ = ~new_A5935_ | ~new_A5936_;
  assign new_A5925_ = ~new_A5910_ ^ new_A5922_;
  assign new_A5924_ = new_A5932_ | new_A5909_;
  assign new_A5923_ = new_A5929_ & new_A5910_;
  assign new_A5922_ = new_A5931_ & new_A5930_;
  assign new_A5921_ = new_A5926_ & new_A5910_;
  assign new_A5920_ = new_A5928_ & new_A5927_;
  assign new_A5919_ = new_A5920_ ^ new_A5910_;
  assign new_A5918_ = new_A5908_ ^ new_A5909_;
  assign A5917 = new_A5918_ & new_A5925_;
  assign A5916 = new_A5918_ & new_A5924_;
  assign A5915 = new_A5923_ | new_A5922_;
  assign A5914 = new_A5921_ | new_A5920_;
  assign A5913 = new_A5919_ & new_A5918_;
  assign new_A5912_ = new_B207_;
  assign new_A5911_ = new_B174_;
  assign new_A5910_ = new_B141_;
  assign new_A5909_ = new_B108_;
  assign new_A5908_ = new_B75_;
  assign new_A5907_ = new_A5885_ & new_A5900_;
  assign new_A5906_ = ~new_A5885_ & ~new_A5907_;
  assign new_A5905_ = new_A5885_ | new_A5900_;
  assign new_A5904_ = ~new_A5878_ | ~new_A5879_;
  assign new_A5903_ = new_A5885_ | new_A5900_;
  assign new_A5902_ = ~new_A5901_ & ~new_A5885_;
  assign new_A5901_ = new_A5885_ & new_A5900_;
  assign new_A5900_ = ~new_A5876_ | ~new_A5877_;
  assign new_A5899_ = new_A5877_ & new_A5889_;
  assign new_A5898_ = new_A5878_ | new_A5885_;
  assign new_A5897_ = new_A5878_ | new_A5879_;
  assign new_A5896_ = ~new_A5906_ | ~new_A5905_;
  assign new_A5895_ = new_A5904_ & new_A5897_;
  assign new_A5894_ = new_A5878_ ^ new_A5885_;
  assign new_A5893_ = ~new_A5902_ | ~new_A5903_;
  assign new_A5892_ = ~new_A5877_ ^ new_A5889_;
  assign new_A5891_ = new_A5899_ | new_A5876_;
  assign new_A5890_ = new_A5896_ & new_A5877_;
  assign new_A5889_ = new_A5898_ & new_A5897_;
  assign new_A5888_ = new_A5893_ & new_A5877_;
  assign new_A5887_ = new_A5895_ & new_A5894_;
  assign new_A5886_ = new_A5887_ ^ new_A5877_;
  assign new_A5885_ = new_A5875_ ^ new_A5876_;
  assign A5884 = new_A5885_ & new_A5892_;
  assign A5883 = new_A5885_ & new_A5891_;
  assign A5882 = new_A5890_ | new_A5889_;
  assign A5881 = new_A5888_ | new_A5887_;
  assign A5880 = new_A5886_ & new_A5885_;
  assign new_A5879_ = new_B42_;
  assign new_A5878_ = new_B9_;
  assign new_A5877_ = new_A9975_;
  assign new_A5876_ = new_A9942_;
  assign new_A5875_ = new_A9909_;
  assign new_A5874_ = new_A5852_ & new_A5867_;
  assign new_A5873_ = ~new_A5852_ & ~new_A5874_;
  assign new_A5872_ = new_A5852_ | new_A5867_;
  assign new_A5871_ = ~new_A5845_ | ~new_A5846_;
  assign new_A5870_ = new_A5852_ | new_A5867_;
  assign new_A5869_ = ~new_A5868_ & ~new_A5852_;
  assign new_A5868_ = new_A5852_ & new_A5867_;
  assign new_A5867_ = ~new_A5843_ | ~new_A5844_;
  assign new_A5866_ = new_A5844_ & new_A5856_;
  assign new_A5865_ = new_A5845_ | new_A5852_;
  assign new_A5864_ = new_A5845_ | new_A5846_;
  assign new_A5863_ = ~new_A5873_ | ~new_A5872_;
  assign new_A5862_ = new_A5871_ & new_A5864_;
  assign new_A5861_ = new_A5845_ ^ new_A5852_;
  assign new_A5860_ = ~new_A5869_ | ~new_A5870_;
  assign new_A5859_ = ~new_A5844_ ^ new_A5856_;
  assign new_A5858_ = new_A5866_ | new_A5843_;
  assign new_A5857_ = new_A5863_ & new_A5844_;
  assign new_A5856_ = new_A5865_ & new_A5864_;
  assign new_A5855_ = new_A5860_ & new_A5844_;
  assign new_A5854_ = new_A5862_ & new_A5861_;
  assign new_A5853_ = new_A5854_ ^ new_A5844_;
  assign new_A5852_ = new_A5842_ ^ new_A5843_;
  assign A5851 = new_A5852_ & new_A5859_;
  assign A5850 = new_A5852_ & new_A5858_;
  assign A5849 = new_A5857_ | new_A5856_;
  assign A5848 = new_A5855_ | new_A5854_;
  assign A5847 = new_A5853_ & new_A5852_;
  assign new_A5846_ = new_A9876_;
  assign new_A5845_ = new_A9843_;
  assign new_A5844_ = new_A9810_;
  assign new_A5843_ = new_A9777_;
  assign new_A5842_ = new_A9744_;
  assign new_A5841_ = new_A5819_ & new_A5834_;
  assign new_A5840_ = ~new_A5819_ & ~new_A5841_;
  assign new_A5839_ = new_A5819_ | new_A5834_;
  assign new_A5838_ = ~new_A5812_ | ~new_A5813_;
  assign new_A5837_ = new_A5819_ | new_A5834_;
  assign new_A5836_ = ~new_A5835_ & ~new_A5819_;
  assign new_A5835_ = new_A5819_ & new_A5834_;
  assign new_A5834_ = ~new_A5810_ | ~new_A5811_;
  assign new_A5833_ = new_A5811_ & new_A5823_;
  assign new_A5832_ = new_A5812_ | new_A5819_;
  assign new_A5831_ = new_A5812_ | new_A5813_;
  assign new_A5830_ = ~new_A5840_ | ~new_A5839_;
  assign new_A5829_ = new_A5838_ & new_A5831_;
  assign new_A5828_ = new_A5812_ ^ new_A5819_;
  assign new_A5827_ = ~new_A5836_ | ~new_A5837_;
  assign new_A5826_ = ~new_A5811_ ^ new_A5823_;
  assign new_A5825_ = new_A5833_ | new_A5810_;
  assign new_A5824_ = new_A5830_ & new_A5811_;
  assign new_A5823_ = new_A5832_ & new_A5831_;
  assign new_A5822_ = new_A5827_ & new_A5811_;
  assign new_A5821_ = new_A5829_ & new_A5828_;
  assign new_A5820_ = new_A5821_ ^ new_A5811_;
  assign new_A5819_ = new_A5809_ ^ new_A5810_;
  assign A5818 = new_A5819_ & new_A5826_;
  assign A5817 = new_A5819_ & new_A5825_;
  assign A5816 = new_A5824_ | new_A5823_;
  assign A5815 = new_A5822_ | new_A5821_;
  assign A5814 = new_A5820_ & new_A5819_;
  assign new_A5813_ = new_A9711_;
  assign new_A5812_ = new_A9678_;
  assign new_A5811_ = new_A9645_;
  assign new_A5810_ = new_A9612_;
  assign new_A5809_ = new_A9579_;
  assign new_A5808_ = new_A5786_ & new_A5801_;
  assign new_A5807_ = ~new_A5786_ & ~new_A5808_;
  assign new_A5806_ = new_A5786_ | new_A5801_;
  assign new_A5805_ = ~new_A5779_ | ~new_A5780_;
  assign new_A5804_ = new_A5786_ | new_A5801_;
  assign new_A5803_ = ~new_A5802_ & ~new_A5786_;
  assign new_A5802_ = new_A5786_ & new_A5801_;
  assign new_A5801_ = ~new_A5777_ | ~new_A5778_;
  assign new_A5800_ = new_A5778_ & new_A5790_;
  assign new_A5799_ = new_A5779_ | new_A5786_;
  assign new_A5798_ = new_A5779_ | new_A5780_;
  assign new_A5797_ = ~new_A5807_ | ~new_A5806_;
  assign new_A5796_ = new_A5805_ & new_A5798_;
  assign new_A5795_ = new_A5779_ ^ new_A5786_;
  assign new_A5794_ = ~new_A5803_ | ~new_A5804_;
  assign new_A5793_ = ~new_A5778_ ^ new_A5790_;
  assign new_A5792_ = new_A5800_ | new_A5777_;
  assign new_A5791_ = new_A5797_ & new_A5778_;
  assign new_A5790_ = new_A5799_ & new_A5798_;
  assign new_A5789_ = new_A5794_ & new_A5778_;
  assign new_A5788_ = new_A5796_ & new_A5795_;
  assign new_A5787_ = new_A5788_ ^ new_A5778_;
  assign new_A5786_ = new_A5776_ ^ new_A5777_;
  assign A5785 = new_A5786_ & new_A5793_;
  assign A5784 = new_A5786_ & new_A5792_;
  assign A5783 = new_A5791_ | new_A5790_;
  assign A5782 = new_A5789_ | new_A5788_;
  assign A5781 = new_A5787_ & new_A5786_;
  assign new_A5780_ = new_A9546_;
  assign new_A5779_ = new_A9513_;
  assign new_A5778_ = new_A9480_;
  assign new_A5777_ = new_A9447_;
  assign new_A5776_ = new_A9414_;
  assign new_A5775_ = new_A5753_ & new_A5768_;
  assign new_A5774_ = ~new_A5753_ & ~new_A5775_;
  assign new_A5773_ = new_A5753_ | new_A5768_;
  assign new_A5772_ = ~new_A5746_ | ~new_A5747_;
  assign new_A5771_ = new_A5753_ | new_A5768_;
  assign new_A5770_ = ~new_A5769_ & ~new_A5753_;
  assign new_A5769_ = new_A5753_ & new_A5768_;
  assign new_A5768_ = ~new_A5744_ | ~new_A5745_;
  assign new_A5767_ = new_A5745_ & new_A5757_;
  assign new_A5766_ = new_A5746_ | new_A5753_;
  assign new_A5765_ = new_A5746_ | new_A5747_;
  assign new_A5764_ = ~new_A5774_ | ~new_A5773_;
  assign new_A5763_ = new_A5772_ & new_A5765_;
  assign new_A5762_ = new_A5746_ ^ new_A5753_;
  assign new_A5761_ = ~new_A5770_ | ~new_A5771_;
  assign new_A5760_ = ~new_A5745_ ^ new_A5757_;
  assign new_A5759_ = new_A5767_ | new_A5744_;
  assign new_A5758_ = new_A5764_ & new_A5745_;
  assign new_A5757_ = new_A5766_ & new_A5765_;
  assign new_A5756_ = new_A5761_ & new_A5745_;
  assign new_A5755_ = new_A5763_ & new_A5762_;
  assign new_A5754_ = new_A5755_ ^ new_A5745_;
  assign new_A5753_ = new_A5743_ ^ new_A5744_;
  assign A5752 = new_A5753_ & new_A5760_;
  assign A5751 = new_A5753_ & new_A5759_;
  assign A5750 = new_A5758_ | new_A5757_;
  assign A5749 = new_A5756_ | new_A5755_;
  assign A5748 = new_A5754_ & new_A5753_;
  assign new_A5747_ = new_A9381_;
  assign new_A5746_ = new_A9348_;
  assign new_A5745_ = new_A9315_;
  assign new_A5744_ = new_A9282_;
  assign new_A5743_ = new_A9249_;
  assign new_A5742_ = new_A5720_ & new_A5735_;
  assign new_A5741_ = ~new_A5720_ & ~new_A5742_;
  assign new_A5740_ = new_A5720_ | new_A5735_;
  assign new_A5739_ = ~new_A5713_ | ~new_A5714_;
  assign new_A5738_ = new_A5720_ | new_A5735_;
  assign new_A5737_ = ~new_A5736_ & ~new_A5720_;
  assign new_A5736_ = new_A5720_ & new_A5735_;
  assign new_A5735_ = ~new_A5711_ | ~new_A5712_;
  assign new_A5734_ = new_A5712_ & new_A5724_;
  assign new_A5733_ = new_A5713_ | new_A5720_;
  assign new_A5732_ = new_A5713_ | new_A5714_;
  assign new_A5731_ = ~new_A5741_ | ~new_A5740_;
  assign new_A5730_ = new_A5739_ & new_A5732_;
  assign new_A5729_ = new_A5713_ ^ new_A5720_;
  assign new_A5728_ = ~new_A5737_ | ~new_A5738_;
  assign new_A5727_ = ~new_A5712_ ^ new_A5724_;
  assign new_A5726_ = new_A5734_ | new_A5711_;
  assign new_A5725_ = new_A5731_ & new_A5712_;
  assign new_A5724_ = new_A5733_ & new_A5732_;
  assign new_A5723_ = new_A5728_ & new_A5712_;
  assign new_A5722_ = new_A5730_ & new_A5729_;
  assign new_A5721_ = new_A5722_ ^ new_A5712_;
  assign new_A5720_ = new_A5710_ ^ new_A5711_;
  assign A5719 = new_A5720_ & new_A5727_;
  assign A5718 = new_A5720_ & new_A5726_;
  assign A5717 = new_A5725_ | new_A5724_;
  assign A5716 = new_A5723_ | new_A5722_;
  assign A5715 = new_A5721_ & new_A5720_;
  assign new_A5714_ = new_A9216_;
  assign new_A5713_ = new_A9183_;
  assign new_A5712_ = new_A9150_;
  assign new_A5711_ = new_A9117_;
  assign new_A5710_ = new_A9084_;
  assign new_A5709_ = new_A5687_ & new_A5702_;
  assign new_A5708_ = ~new_A5687_ & ~new_A5709_;
  assign new_A5707_ = new_A5687_ | new_A5702_;
  assign new_A5706_ = ~new_A5680_ | ~new_A5681_;
  assign new_A5705_ = new_A5687_ | new_A5702_;
  assign new_A5704_ = ~new_A5703_ & ~new_A5687_;
  assign new_A5703_ = new_A5687_ & new_A5702_;
  assign new_A5702_ = ~new_A5678_ | ~new_A5679_;
  assign new_A5701_ = new_A5679_ & new_A5691_;
  assign new_A5700_ = new_A5680_ | new_A5687_;
  assign new_A5699_ = new_A5680_ | new_A5681_;
  assign new_A5698_ = ~new_A5708_ | ~new_A5707_;
  assign new_A5697_ = new_A5706_ & new_A5699_;
  assign new_A5696_ = new_A5680_ ^ new_A5687_;
  assign new_A5695_ = ~new_A5704_ | ~new_A5705_;
  assign new_A5694_ = ~new_A5679_ ^ new_A5691_;
  assign new_A5693_ = new_A5701_ | new_A5678_;
  assign new_A5692_ = new_A5698_ & new_A5679_;
  assign new_A5691_ = new_A5700_ & new_A5699_;
  assign new_A5690_ = new_A5695_ & new_A5679_;
  assign new_A5689_ = new_A5697_ & new_A5696_;
  assign new_A5688_ = new_A5689_ ^ new_A5679_;
  assign new_A5687_ = new_A5677_ ^ new_A5678_;
  assign A5686 = new_A5687_ & new_A5694_;
  assign A5685 = new_A5687_ & new_A5693_;
  assign A5684 = new_A5692_ | new_A5691_;
  assign A5683 = new_A5690_ | new_A5689_;
  assign A5682 = new_A5688_ & new_A5687_;
  assign new_A5681_ = new_A9051_;
  assign new_A5680_ = new_A9018_;
  assign new_A5679_ = new_A8985_;
  assign new_A5678_ = new_A8952_;
  assign new_A5677_ = new_A8919_;
  assign new_A5676_ = new_A5654_ & new_A5669_;
  assign new_A5675_ = ~new_A5654_ & ~new_A5676_;
  assign new_A5674_ = new_A5654_ | new_A5669_;
  assign new_A5673_ = ~new_A5647_ | ~new_A5648_;
  assign new_A5672_ = new_A5654_ | new_A5669_;
  assign new_A5671_ = ~new_A5670_ & ~new_A5654_;
  assign new_A5670_ = new_A5654_ & new_A5669_;
  assign new_A5669_ = ~new_A5645_ | ~new_A5646_;
  assign new_A5668_ = new_A5646_ & new_A5658_;
  assign new_A5667_ = new_A5647_ | new_A5654_;
  assign new_A5666_ = new_A5647_ | new_A5648_;
  assign new_A5665_ = ~new_A5675_ | ~new_A5674_;
  assign new_A5664_ = new_A5673_ & new_A5666_;
  assign new_A5663_ = new_A5647_ ^ new_A5654_;
  assign new_A5662_ = ~new_A5671_ | ~new_A5672_;
  assign new_A5661_ = ~new_A5646_ ^ new_A5658_;
  assign new_A5660_ = new_A5668_ | new_A5645_;
  assign new_A5659_ = new_A5665_ & new_A5646_;
  assign new_A5658_ = new_A5667_ & new_A5666_;
  assign new_A5657_ = new_A5662_ & new_A5646_;
  assign new_A5656_ = new_A5664_ & new_A5663_;
  assign new_A5655_ = new_A5656_ ^ new_A5646_;
  assign new_A5654_ = new_A5644_ ^ new_A5645_;
  assign A5653 = new_A5654_ & new_A5661_;
  assign A5652 = new_A5654_ & new_A5660_;
  assign A5651 = new_A5659_ | new_A5658_;
  assign A5650 = new_A5657_ | new_A5656_;
  assign A5649 = new_A5655_ & new_A5654_;
  assign new_A5648_ = new_A8886_;
  assign new_A5647_ = new_A8853_;
  assign new_A5646_ = new_A8820_;
  assign new_A5645_ = new_A8787_;
  assign new_A5644_ = new_A8754_;
  assign new_A5643_ = new_A5621_ & new_A5636_;
  assign new_A5642_ = ~new_A5621_ & ~new_A5643_;
  assign new_A5641_ = new_A5621_ | new_A5636_;
  assign new_A5640_ = ~new_A5614_ | ~new_A5615_;
  assign new_A5639_ = new_A5621_ | new_A5636_;
  assign new_A5638_ = ~new_A5637_ & ~new_A5621_;
  assign new_A5637_ = new_A5621_ & new_A5636_;
  assign new_A5636_ = ~new_A5612_ | ~new_A5613_;
  assign new_A5635_ = new_A5613_ & new_A5625_;
  assign new_A5634_ = new_A5614_ | new_A5621_;
  assign new_A5633_ = new_A5614_ | new_A5615_;
  assign new_A5632_ = ~new_A5642_ | ~new_A5641_;
  assign new_A5631_ = new_A5640_ & new_A5633_;
  assign new_A5630_ = new_A5614_ ^ new_A5621_;
  assign new_A5629_ = ~new_A5638_ | ~new_A5639_;
  assign new_A5628_ = ~new_A5613_ ^ new_A5625_;
  assign new_A5627_ = new_A5635_ | new_A5612_;
  assign new_A5626_ = new_A5632_ & new_A5613_;
  assign new_A5625_ = new_A5634_ & new_A5633_;
  assign new_A5624_ = new_A5629_ & new_A5613_;
  assign new_A5623_ = new_A5631_ & new_A5630_;
  assign new_A5622_ = new_A5623_ ^ new_A5613_;
  assign new_A5621_ = new_A5611_ ^ new_A5612_;
  assign A5620 = new_A5621_ & new_A5628_;
  assign A5619 = new_A5621_ & new_A5627_;
  assign A5618 = new_A5626_ | new_A5625_;
  assign A5617 = new_A5624_ | new_A5623_;
  assign A5616 = new_A5622_ & new_A5621_;
  assign new_A5615_ = new_A8721_;
  assign new_A5614_ = new_A8688_;
  assign new_A5613_ = new_A8655_;
  assign new_A5612_ = new_A8622_;
  assign new_A5611_ = new_A8589_;
  assign new_A5610_ = new_A5588_ & new_A5603_;
  assign new_A5609_ = ~new_A5588_ & ~new_A5610_;
  assign new_A5608_ = new_A5588_ | new_A5603_;
  assign new_A5607_ = ~new_A5581_ | ~new_A5582_;
  assign new_A5606_ = new_A5588_ | new_A5603_;
  assign new_A5605_ = ~new_A5604_ & ~new_A5588_;
  assign new_A5604_ = new_A5588_ & new_A5603_;
  assign new_A5603_ = ~new_A5579_ | ~new_A5580_;
  assign new_A5602_ = new_A5580_ & new_A5592_;
  assign new_A5601_ = new_A5581_ | new_A5588_;
  assign new_A5600_ = new_A5581_ | new_A5582_;
  assign new_A5599_ = ~new_A5609_ | ~new_A5608_;
  assign new_A5598_ = new_A5607_ & new_A5600_;
  assign new_A5597_ = new_A5581_ ^ new_A5588_;
  assign new_A5596_ = ~new_A5605_ | ~new_A5606_;
  assign new_A5595_ = ~new_A5580_ ^ new_A5592_;
  assign new_A5594_ = new_A5602_ | new_A5579_;
  assign new_A5593_ = new_A5599_ & new_A5580_;
  assign new_A5592_ = new_A5601_ & new_A5600_;
  assign new_A5591_ = new_A5596_ & new_A5580_;
  assign new_A5590_ = new_A5598_ & new_A5597_;
  assign new_A5589_ = new_A5590_ ^ new_A5580_;
  assign new_A5588_ = new_A5578_ ^ new_A5579_;
  assign A5587 = new_A5588_ & new_A5595_;
  assign A5586 = new_A5588_ & new_A5594_;
  assign A5585 = new_A5593_ | new_A5592_;
  assign A5584 = new_A5591_ | new_A5590_;
  assign A5583 = new_A5589_ & new_A5588_;
  assign new_A5582_ = new_A8556_;
  assign new_A5581_ = new_A8523_;
  assign new_A5580_ = new_A8490_;
  assign new_A5579_ = new_A8457_;
  assign new_A5578_ = new_A8424_;
  assign new_A5577_ = new_A5555_ & new_A5570_;
  assign new_A5576_ = ~new_A5555_ & ~new_A5577_;
  assign new_A5575_ = new_A5555_ | new_A5570_;
  assign new_A5574_ = ~new_A5548_ | ~new_A5549_;
  assign new_A5573_ = new_A5555_ | new_A5570_;
  assign new_A5572_ = ~new_A5571_ & ~new_A5555_;
  assign new_A5571_ = new_A5555_ & new_A5570_;
  assign new_A5570_ = ~new_A5546_ | ~new_A5547_;
  assign new_A5569_ = new_A5547_ & new_A5559_;
  assign new_A5568_ = new_A5548_ | new_A5555_;
  assign new_A5567_ = new_A5548_ | new_A5549_;
  assign new_A5566_ = ~new_A5576_ | ~new_A5575_;
  assign new_A5565_ = new_A5574_ & new_A5567_;
  assign new_A5564_ = new_A5548_ ^ new_A5555_;
  assign new_A5563_ = ~new_A5572_ | ~new_A5573_;
  assign new_A5562_ = ~new_A5547_ ^ new_A5559_;
  assign new_A5561_ = new_A5569_ | new_A5546_;
  assign new_A5560_ = new_A5566_ & new_A5547_;
  assign new_A5559_ = new_A5568_ & new_A5567_;
  assign new_A5558_ = new_A5563_ & new_A5547_;
  assign new_A5557_ = new_A5565_ & new_A5564_;
  assign new_A5556_ = new_A5557_ ^ new_A5547_;
  assign new_A5555_ = new_A5545_ ^ new_A5546_;
  assign A5554 = new_A5555_ & new_A5562_;
  assign A5553 = new_A5555_ & new_A5561_;
  assign A5552 = new_A5560_ | new_A5559_;
  assign A5551 = new_A5558_ | new_A5557_;
  assign A5550 = new_A5556_ & new_A5555_;
  assign new_A5549_ = new_A8391_;
  assign new_A5548_ = new_A8358_;
  assign new_A5547_ = new_A8325_;
  assign new_A5546_ = new_A8292_;
  assign new_A5545_ = new_A8259_;
  assign new_A5544_ = new_A5522_ & new_A5537_;
  assign new_A5543_ = ~new_A5522_ & ~new_A5544_;
  assign new_A5542_ = new_A5522_ | new_A5537_;
  assign new_A5541_ = ~new_A5515_ | ~new_A5516_;
  assign new_A5540_ = new_A5522_ | new_A5537_;
  assign new_A5539_ = ~new_A5538_ & ~new_A5522_;
  assign new_A5538_ = new_A5522_ & new_A5537_;
  assign new_A5537_ = ~new_A5513_ | ~new_A5514_;
  assign new_A5536_ = new_A5514_ & new_A5526_;
  assign new_A5535_ = new_A5515_ | new_A5522_;
  assign new_A5534_ = new_A5515_ | new_A5516_;
  assign new_A5533_ = ~new_A5543_ | ~new_A5542_;
  assign new_A5532_ = new_A5541_ & new_A5534_;
  assign new_A5531_ = new_A5515_ ^ new_A5522_;
  assign new_A5530_ = ~new_A5539_ | ~new_A5540_;
  assign new_A5529_ = ~new_A5514_ ^ new_A5526_;
  assign new_A5528_ = new_A5536_ | new_A5513_;
  assign new_A5527_ = new_A5533_ & new_A5514_;
  assign new_A5526_ = new_A5535_ & new_A5534_;
  assign new_A5525_ = new_A5530_ & new_A5514_;
  assign new_A5524_ = new_A5532_ & new_A5531_;
  assign new_A5523_ = new_A5524_ ^ new_A5514_;
  assign new_A5522_ = new_A5512_ ^ new_A5513_;
  assign A5521 = new_A5522_ & new_A5529_;
  assign A5520 = new_A5522_ & new_A5528_;
  assign A5519 = new_A5527_ | new_A5526_;
  assign A5518 = new_A5525_ | new_A5524_;
  assign A5517 = new_A5523_ & new_A5522_;
  assign new_A5516_ = new_A8226_;
  assign new_A5515_ = new_A8193_;
  assign new_A5514_ = new_A8160_;
  assign new_A5513_ = new_A8127_;
  assign new_A5512_ = new_A8094_;
  assign new_A5511_ = new_A5489_ & new_A5504_;
  assign new_A5510_ = ~new_A5489_ & ~new_A5511_;
  assign new_A5509_ = new_A5489_ | new_A5504_;
  assign new_A5508_ = ~new_A5482_ | ~new_A5483_;
  assign new_A5507_ = new_A5489_ | new_A5504_;
  assign new_A5506_ = ~new_A5505_ & ~new_A5489_;
  assign new_A5505_ = new_A5489_ & new_A5504_;
  assign new_A5504_ = ~new_A5480_ | ~new_A5481_;
  assign new_A5503_ = new_A5481_ & new_A5493_;
  assign new_A5502_ = new_A5482_ | new_A5489_;
  assign new_A5501_ = new_A5482_ | new_A5483_;
  assign new_A5500_ = ~new_A5510_ | ~new_A5509_;
  assign new_A5499_ = new_A5508_ & new_A5501_;
  assign new_A5498_ = new_A5482_ ^ new_A5489_;
  assign new_A5497_ = ~new_A5506_ | ~new_A5507_;
  assign new_A5496_ = ~new_A5481_ ^ new_A5493_;
  assign new_A5495_ = new_A5503_ | new_A5480_;
  assign new_A5494_ = new_A5500_ & new_A5481_;
  assign new_A5493_ = new_A5502_ & new_A5501_;
  assign new_A5492_ = new_A5497_ & new_A5481_;
  assign new_A5491_ = new_A5499_ & new_A5498_;
  assign new_A5490_ = new_A5491_ ^ new_A5481_;
  assign new_A5489_ = new_A5479_ ^ new_A5480_;
  assign A5488 = new_A5489_ & new_A5496_;
  assign A5487 = new_A5489_ & new_A5495_;
  assign A5486 = new_A5494_ | new_A5493_;
  assign A5485 = new_A5492_ | new_A5491_;
  assign A5484 = new_A5490_ & new_A5489_;
  assign new_A5483_ = new_A8061_;
  assign new_A5482_ = new_A8028_;
  assign new_A5481_ = new_A7995_;
  assign new_A5480_ = new_A7962_;
  assign new_A5479_ = new_A7929_;
  assign new_A5478_ = new_A5456_ & new_A5471_;
  assign new_A5477_ = ~new_A5456_ & ~new_A5478_;
  assign new_A5476_ = new_A5456_ | new_A5471_;
  assign new_A5475_ = ~new_A5449_ | ~new_A5450_;
  assign new_A5474_ = new_A5456_ | new_A5471_;
  assign new_A5473_ = ~new_A5472_ & ~new_A5456_;
  assign new_A5472_ = new_A5456_ & new_A5471_;
  assign new_A5471_ = ~new_A5447_ | ~new_A5448_;
  assign new_A5470_ = new_A5448_ & new_A5460_;
  assign new_A5469_ = new_A5449_ | new_A5456_;
  assign new_A5468_ = new_A5449_ | new_A5450_;
  assign new_A5467_ = ~new_A5477_ | ~new_A5476_;
  assign new_A5466_ = new_A5475_ & new_A5468_;
  assign new_A5465_ = new_A5449_ ^ new_A5456_;
  assign new_A5464_ = ~new_A5473_ | ~new_A5474_;
  assign new_A5463_ = ~new_A5448_ ^ new_A5460_;
  assign new_A5462_ = new_A5470_ | new_A5447_;
  assign new_A5461_ = new_A5467_ & new_A5448_;
  assign new_A5460_ = new_A5469_ & new_A5468_;
  assign new_A5459_ = new_A5464_ & new_A5448_;
  assign new_A5458_ = new_A5466_ & new_A5465_;
  assign new_A5457_ = new_A5458_ ^ new_A5448_;
  assign new_A5456_ = new_A5446_ ^ new_A5447_;
  assign A5455 = new_A5456_ & new_A5463_;
  assign A5454 = new_A5456_ & new_A5462_;
  assign A5453 = new_A5461_ | new_A5460_;
  assign A5452 = new_A5459_ | new_A5458_;
  assign A5451 = new_A5457_ & new_A5456_;
  assign new_A5450_ = new_A7896_;
  assign new_A5449_ = new_A7863_;
  assign new_A5448_ = new_A7830_;
  assign new_A5447_ = new_A7797_;
  assign new_A5446_ = new_A7764_;
  assign new_A5445_ = new_A5423_ & new_A5438_;
  assign new_A5444_ = ~new_A5423_ & ~new_A5445_;
  assign new_A5443_ = new_A5423_ | new_A5438_;
  assign new_A5442_ = ~new_A5416_ | ~new_A5417_;
  assign new_A5441_ = new_A5423_ | new_A5438_;
  assign new_A5440_ = ~new_A5439_ & ~new_A5423_;
  assign new_A5439_ = new_A5423_ & new_A5438_;
  assign new_A5438_ = ~new_A5414_ | ~new_A5415_;
  assign new_A5437_ = new_A5415_ & new_A5427_;
  assign new_A5436_ = new_A5416_ | new_A5423_;
  assign new_A5435_ = new_A5416_ | new_A5417_;
  assign new_A5434_ = ~new_A5444_ | ~new_A5443_;
  assign new_A5433_ = new_A5442_ & new_A5435_;
  assign new_A5432_ = new_A5416_ ^ new_A5423_;
  assign new_A5431_ = ~new_A5440_ | ~new_A5441_;
  assign new_A5430_ = ~new_A5415_ ^ new_A5427_;
  assign new_A5429_ = new_A5437_ | new_A5414_;
  assign new_A5428_ = new_A5434_ & new_A5415_;
  assign new_A5427_ = new_A5436_ & new_A5435_;
  assign new_A5426_ = new_A5431_ & new_A5415_;
  assign new_A5425_ = new_A5433_ & new_A5432_;
  assign new_A5424_ = new_A5425_ ^ new_A5415_;
  assign new_A5423_ = new_A5413_ ^ new_A5414_;
  assign A5422 = new_A5423_ & new_A5430_;
  assign A5421 = new_A5423_ & new_A5429_;
  assign A5420 = new_A5428_ | new_A5427_;
  assign A5419 = new_A5426_ | new_A5425_;
  assign A5418 = new_A5424_ & new_A5423_;
  assign new_A5417_ = new_A7731_;
  assign new_A5416_ = new_A7698_;
  assign new_A5415_ = new_A7665_;
  assign new_A5414_ = new_A7632_;
  assign new_A5413_ = new_A7599_;
  assign new_A5412_ = new_A5390_ & new_A5405_;
  assign new_A5411_ = ~new_A5390_ & ~new_A5412_;
  assign new_A5410_ = new_A5390_ | new_A5405_;
  assign new_A5409_ = ~new_A5383_ | ~new_A5384_;
  assign new_A5408_ = new_A5390_ | new_A5405_;
  assign new_A5407_ = ~new_A5406_ & ~new_A5390_;
  assign new_A5406_ = new_A5390_ & new_A5405_;
  assign new_A5405_ = ~new_A5381_ | ~new_A5382_;
  assign new_A5404_ = new_A5382_ & new_A5394_;
  assign new_A5403_ = new_A5383_ | new_A5390_;
  assign new_A5402_ = new_A5383_ | new_A5384_;
  assign new_A5401_ = ~new_A5411_ | ~new_A5410_;
  assign new_A5400_ = new_A5409_ & new_A5402_;
  assign new_A5399_ = new_A5383_ ^ new_A5390_;
  assign new_A5398_ = ~new_A5407_ | ~new_A5408_;
  assign new_A5397_ = ~new_A5382_ ^ new_A5394_;
  assign new_A5396_ = new_A5404_ | new_A5381_;
  assign new_A5395_ = new_A5401_ & new_A5382_;
  assign new_A5394_ = new_A5403_ & new_A5402_;
  assign new_A5393_ = new_A5398_ & new_A5382_;
  assign new_A5392_ = new_A5400_ & new_A5399_;
  assign new_A5391_ = new_A5392_ ^ new_A5382_;
  assign new_A5390_ = new_A5380_ ^ new_A5381_;
  assign A5389 = new_A5390_ & new_A5397_;
  assign A5388 = new_A5390_ & new_A5396_;
  assign A5387 = new_A5395_ | new_A5394_;
  assign A5386 = new_A5393_ | new_A5392_;
  assign A5385 = new_A5391_ & new_A5390_;
  assign new_A5384_ = new_A7566_;
  assign new_A5383_ = new_A7533_;
  assign new_A5382_ = new_A7500_;
  assign new_A5381_ = new_A7467_;
  assign new_A5380_ = new_A7434_;
  assign new_A5379_ = new_A5357_ & new_A5372_;
  assign new_A5378_ = ~new_A5357_ & ~new_A5379_;
  assign new_A5377_ = new_A5357_ | new_A5372_;
  assign new_A5376_ = ~new_A5350_ | ~new_A5351_;
  assign new_A5375_ = new_A5357_ | new_A5372_;
  assign new_A5374_ = ~new_A5373_ & ~new_A5357_;
  assign new_A5373_ = new_A5357_ & new_A5372_;
  assign new_A5372_ = ~new_A5348_ | ~new_A5349_;
  assign new_A5371_ = new_A5349_ & new_A5361_;
  assign new_A5370_ = new_A5350_ | new_A5357_;
  assign new_A5369_ = new_A5350_ | new_A5351_;
  assign new_A5368_ = ~new_A5378_ | ~new_A5377_;
  assign new_A5367_ = new_A5376_ & new_A5369_;
  assign new_A5366_ = new_A5350_ ^ new_A5357_;
  assign new_A5365_ = ~new_A5374_ | ~new_A5375_;
  assign new_A5364_ = ~new_A5349_ ^ new_A5361_;
  assign new_A5363_ = new_A5371_ | new_A5348_;
  assign new_A5362_ = new_A5368_ & new_A5349_;
  assign new_A5361_ = new_A5370_ & new_A5369_;
  assign new_A5360_ = new_A5365_ & new_A5349_;
  assign new_A5359_ = new_A5367_ & new_A5366_;
  assign new_A5358_ = new_A5359_ ^ new_A5349_;
  assign new_A5357_ = new_A5347_ ^ new_A5348_;
  assign A5356 = new_A5357_ & new_A5364_;
  assign A5355 = new_A5357_ & new_A5363_;
  assign A5354 = new_A5362_ | new_A5361_;
  assign A5353 = new_A5360_ | new_A5359_;
  assign A5352 = new_A5358_ & new_A5357_;
  assign new_A5351_ = new_A7401_;
  assign new_A5350_ = new_A7368_;
  assign new_A5349_ = new_A7335_;
  assign new_A5348_ = new_A7302_;
  assign new_A5347_ = new_A7269_;
  assign new_A5346_ = new_A5324_ & new_A5339_;
  assign new_A5345_ = ~new_A5324_ & ~new_A5346_;
  assign new_A5344_ = new_A5324_ | new_A5339_;
  assign new_A5343_ = ~new_A5317_ | ~new_A5318_;
  assign new_A5342_ = new_A5324_ | new_A5339_;
  assign new_A5341_ = ~new_A5340_ & ~new_A5324_;
  assign new_A5340_ = new_A5324_ & new_A5339_;
  assign new_A5339_ = ~new_A5315_ | ~new_A5316_;
  assign new_A5338_ = new_A5316_ & new_A5328_;
  assign new_A5337_ = new_A5317_ | new_A5324_;
  assign new_A5336_ = new_A5317_ | new_A5318_;
  assign new_A5335_ = ~new_A5345_ | ~new_A5344_;
  assign new_A5334_ = new_A5343_ & new_A5336_;
  assign new_A5333_ = new_A5317_ ^ new_A5324_;
  assign new_A5332_ = ~new_A5341_ | ~new_A5342_;
  assign new_A5331_ = ~new_A5316_ ^ new_A5328_;
  assign new_A5330_ = new_A5338_ | new_A5315_;
  assign new_A5329_ = new_A5335_ & new_A5316_;
  assign new_A5328_ = new_A5337_ & new_A5336_;
  assign new_A5327_ = new_A5332_ & new_A5316_;
  assign new_A5326_ = new_A5334_ & new_A5333_;
  assign new_A5325_ = new_A5326_ ^ new_A5316_;
  assign new_A5324_ = new_A5314_ ^ new_A5315_;
  assign A5323 = new_A5324_ & new_A5331_;
  assign A5322 = new_A5324_ & new_A5330_;
  assign A5321 = new_A5329_ | new_A5328_;
  assign A5320 = new_A5327_ | new_A5326_;
  assign A5319 = new_A5325_ & new_A5324_;
  assign new_A5318_ = new_A7236_;
  assign new_A5317_ = new_A7203_;
  assign new_A5316_ = new_A7170_;
  assign new_A5315_ = new_A7137_;
  assign new_A5314_ = new_A7104_;
  assign new_A5313_ = new_A5291_ & new_A5306_;
  assign new_A5312_ = ~new_A5291_ & ~new_A5313_;
  assign new_A5311_ = new_A5291_ | new_A5306_;
  assign new_A5310_ = ~new_A5284_ | ~new_A5285_;
  assign new_A5309_ = new_A5291_ | new_A5306_;
  assign new_A5308_ = ~new_A5307_ & ~new_A5291_;
  assign new_A5307_ = new_A5291_ & new_A5306_;
  assign new_A5306_ = ~new_A5282_ | ~new_A5283_;
  assign new_A5305_ = new_A5283_ & new_A5295_;
  assign new_A5304_ = new_A5284_ | new_A5291_;
  assign new_A5303_ = new_A5284_ | new_A5285_;
  assign new_A5302_ = ~new_A5312_ | ~new_A5311_;
  assign new_A5301_ = new_A5310_ & new_A5303_;
  assign new_A5300_ = new_A5284_ ^ new_A5291_;
  assign new_A5299_ = ~new_A5308_ | ~new_A5309_;
  assign new_A5298_ = ~new_A5283_ ^ new_A5295_;
  assign new_A5297_ = new_A5305_ | new_A5282_;
  assign new_A5296_ = new_A5302_ & new_A5283_;
  assign new_A5295_ = new_A5304_ & new_A5303_;
  assign new_A5294_ = new_A5299_ & new_A5283_;
  assign new_A5293_ = new_A5301_ & new_A5300_;
  assign new_A5292_ = new_A5293_ ^ new_A5283_;
  assign new_A5291_ = new_A5281_ ^ new_A5282_;
  assign A5290 = new_A5291_ & new_A5298_;
  assign A5289 = new_A5291_ & new_A5297_;
  assign A5288 = new_A5296_ | new_A5295_;
  assign A5287 = new_A5294_ | new_A5293_;
  assign A5286 = new_A5292_ & new_A5291_;
  assign new_A5285_ = new_A7071_;
  assign new_A5284_ = new_A7038_;
  assign new_A5283_ = new_A7005_;
  assign new_A5282_ = new_A6972_;
  assign new_A5281_ = new_A6937_;
  assign new_A5280_ = new_A5258_ & new_A5273_;
  assign new_A5279_ = ~new_A5258_ & ~new_A5280_;
  assign new_A5278_ = new_A5258_ | new_A5273_;
  assign new_A5277_ = ~new_A5251_ | ~new_A5252_;
  assign new_A5276_ = new_A5258_ | new_A5273_;
  assign new_A5275_ = ~new_A5274_ & ~new_A5258_;
  assign new_A5274_ = new_A5258_ & new_A5273_;
  assign new_A5273_ = ~new_A5249_ | ~new_A5250_;
  assign new_A5272_ = new_A5250_ & new_A5262_;
  assign new_A5271_ = new_A5251_ | new_A5258_;
  assign new_A5270_ = new_A5251_ | new_A5252_;
  assign new_A5269_ = ~new_A5279_ | ~new_A5278_;
  assign new_A5268_ = new_A5277_ & new_A5270_;
  assign new_A5267_ = new_A5251_ ^ new_A5258_;
  assign new_A5266_ = ~new_A5275_ | ~new_A5276_;
  assign new_A5265_ = ~new_A5250_ ^ new_A5262_;
  assign new_A5264_ = new_A5272_ | new_A5249_;
  assign new_A5263_ = new_A5269_ & new_A5250_;
  assign new_A5262_ = new_A5271_ & new_A5270_;
  assign new_A5261_ = new_A5266_ & new_A5250_;
  assign new_A5260_ = new_A5268_ & new_A5267_;
  assign new_A5259_ = new_A5260_ ^ new_A5250_;
  assign new_A5258_ = new_A5248_ ^ new_A5249_;
  assign A5257 = new_A5258_ & new_A5265_;
  assign A5256 = new_A5258_ & new_A5264_;
  assign A5255 = new_A5263_ | new_A5262_;
  assign A5254 = new_A5261_ | new_A5260_;
  assign A5253 = new_A5259_ & new_A5258_;
  assign new_A5252_ = new_B1031_;
  assign new_A5251_ = new_B998_;
  assign new_A5250_ = new_B965_;
  assign new_A5249_ = new_B932_;
  assign new_A5248_ = new_B899_;
  assign new_A5247_ = new_A5225_ & new_A5240_;
  assign new_A5246_ = ~new_A5225_ & ~new_A5247_;
  assign new_A5245_ = new_A5225_ | new_A5240_;
  assign new_A5244_ = ~new_A5218_ | ~new_A5219_;
  assign new_A5243_ = new_A5225_ | new_A5240_;
  assign new_A5242_ = ~new_A5241_ & ~new_A5225_;
  assign new_A5241_ = new_A5225_ & new_A5240_;
  assign new_A5240_ = ~new_A5216_ | ~new_A5217_;
  assign new_A5239_ = new_A5217_ & new_A5229_;
  assign new_A5238_ = new_A5218_ | new_A5225_;
  assign new_A5237_ = new_A5218_ | new_A5219_;
  assign new_A5236_ = ~new_A5246_ | ~new_A5245_;
  assign new_A5235_ = new_A5244_ & new_A5237_;
  assign new_A5234_ = new_A5218_ ^ new_A5225_;
  assign new_A5233_ = ~new_A5242_ | ~new_A5243_;
  assign new_A5232_ = ~new_A5217_ ^ new_A5229_;
  assign new_A5231_ = new_A5239_ | new_A5216_;
  assign new_A5230_ = new_A5236_ & new_A5217_;
  assign new_A5229_ = new_A5238_ & new_A5237_;
  assign new_A5228_ = new_A5233_ & new_A5217_;
  assign new_A5227_ = new_A5235_ & new_A5234_;
  assign new_A5226_ = new_A5227_ ^ new_A5217_;
  assign new_A5225_ = new_A5215_ ^ new_A5216_;
  assign A5224 = new_A5225_ & new_A5232_;
  assign A5223 = new_A5225_ & new_A5231_;
  assign A5222 = new_A5230_ | new_A5229_;
  assign A5221 = new_A5228_ | new_A5227_;
  assign A5220 = new_A5226_ & new_A5225_;
  assign new_A5219_ = new_B866_;
  assign new_A5218_ = new_B833_;
  assign new_A5217_ = new_B800_;
  assign new_A5216_ = new_B767_;
  assign new_A5215_ = new_B734_;
  assign new_A5214_ = new_A5192_ & new_A5207_;
  assign new_A5213_ = ~new_A5192_ & ~new_A5214_;
  assign new_A5212_ = new_A5192_ | new_A5207_;
  assign new_A5211_ = ~new_A5185_ | ~new_A5186_;
  assign new_A5210_ = new_A5192_ | new_A5207_;
  assign new_A5209_ = ~new_A5208_ & ~new_A5192_;
  assign new_A5208_ = new_A5192_ & new_A5207_;
  assign new_A5207_ = ~new_A5183_ | ~new_A5184_;
  assign new_A5206_ = new_A5184_ & new_A5196_;
  assign new_A5205_ = new_A5185_ | new_A5192_;
  assign new_A5204_ = new_A5185_ | new_A5186_;
  assign new_A5203_ = ~new_A5213_ | ~new_A5212_;
  assign new_A5202_ = new_A5211_ & new_A5204_;
  assign new_A5201_ = new_A5185_ ^ new_A5192_;
  assign new_A5200_ = ~new_A5209_ | ~new_A5210_;
  assign new_A5199_ = ~new_A5184_ ^ new_A5196_;
  assign new_A5198_ = new_A5206_ | new_A5183_;
  assign new_A5197_ = new_A5203_ & new_A5184_;
  assign new_A5196_ = new_A5205_ & new_A5204_;
  assign new_A5195_ = new_A5200_ & new_A5184_;
  assign new_A5194_ = new_A5202_ & new_A5201_;
  assign new_A5193_ = new_A5194_ ^ new_A5184_;
  assign new_A5192_ = new_A5182_ ^ new_A5183_;
  assign A5191 = new_A5192_ & new_A5199_;
  assign A5190 = new_A5192_ & new_A5198_;
  assign A5189 = new_A5197_ | new_A5196_;
  assign A5188 = new_A5195_ | new_A5194_;
  assign A5187 = new_A5193_ & new_A5192_;
  assign new_A5186_ = new_B701_;
  assign new_A5185_ = new_B668_;
  assign new_A5184_ = new_B635_;
  assign new_A5183_ = new_B602_;
  assign new_A5182_ = new_B569_;
  assign new_A5181_ = new_A5159_ & new_A5174_;
  assign new_A5180_ = ~new_A5159_ & ~new_A5181_;
  assign new_A5179_ = new_A5159_ | new_A5174_;
  assign new_A5178_ = ~new_A5152_ | ~new_A5153_;
  assign new_A5177_ = new_A5159_ | new_A5174_;
  assign new_A5176_ = ~new_A5175_ & ~new_A5159_;
  assign new_A5175_ = new_A5159_ & new_A5174_;
  assign new_A5174_ = ~new_A5150_ | ~new_A5151_;
  assign new_A5173_ = new_A5151_ & new_A5163_;
  assign new_A5172_ = new_A5152_ | new_A5159_;
  assign new_A5171_ = new_A5152_ | new_A5153_;
  assign new_A5170_ = ~new_A5180_ | ~new_A5179_;
  assign new_A5169_ = new_A5178_ & new_A5171_;
  assign new_A5168_ = new_A5152_ ^ new_A5159_;
  assign new_A5167_ = ~new_A5176_ | ~new_A5177_;
  assign new_A5166_ = ~new_A5151_ ^ new_A5163_;
  assign new_A5165_ = new_A5173_ | new_A5150_;
  assign new_A5164_ = new_A5170_ & new_A5151_;
  assign new_A5163_ = new_A5172_ & new_A5171_;
  assign new_A5162_ = new_A5167_ & new_A5151_;
  assign new_A5161_ = new_A5169_ & new_A5168_;
  assign new_A5160_ = new_A5161_ ^ new_A5151_;
  assign new_A5159_ = new_A5149_ ^ new_A5150_;
  assign A5158 = new_A5159_ & new_A5166_;
  assign A5157 = new_A5159_ & new_A5165_;
  assign A5156 = new_A5164_ | new_A5163_;
  assign A5155 = new_A5162_ | new_A5161_;
  assign A5154 = new_A5160_ & new_A5159_;
  assign new_A5153_ = new_B536_;
  assign new_A5152_ = new_B503_;
  assign new_A5151_ = new_B470_;
  assign new_A5150_ = new_B437_;
  assign new_A5149_ = new_B404_;
  assign new_A5148_ = new_A5126_ & new_A5141_;
  assign new_A5147_ = ~new_A5126_ & ~new_A5148_;
  assign new_A5146_ = new_A5126_ | new_A5141_;
  assign new_A5145_ = ~new_A5119_ | ~new_A5120_;
  assign new_A5144_ = new_A5126_ | new_A5141_;
  assign new_A5143_ = ~new_A5142_ & ~new_A5126_;
  assign new_A5142_ = new_A5126_ & new_A5141_;
  assign new_A5141_ = ~new_A5117_ | ~new_A5118_;
  assign new_A5140_ = new_A5118_ & new_A5130_;
  assign new_A5139_ = new_A5119_ | new_A5126_;
  assign new_A5138_ = new_A5119_ | new_A5120_;
  assign new_A5137_ = ~new_A5147_ | ~new_A5146_;
  assign new_A5136_ = new_A5145_ & new_A5138_;
  assign new_A5135_ = new_A5119_ ^ new_A5126_;
  assign new_A5134_ = ~new_A5143_ | ~new_A5144_;
  assign new_A5133_ = ~new_A5118_ ^ new_A5130_;
  assign new_A5132_ = new_A5140_ | new_A5117_;
  assign new_A5131_ = new_A5137_ & new_A5118_;
  assign new_A5130_ = new_A5139_ & new_A5138_;
  assign new_A5129_ = new_A5134_ & new_A5118_;
  assign new_A5128_ = new_A5136_ & new_A5135_;
  assign new_A5127_ = new_A5128_ ^ new_A5118_;
  assign new_A5126_ = new_A5116_ ^ new_A5117_;
  assign A5125 = new_A5126_ & new_A5133_;
  assign A5124 = new_A5126_ & new_A5132_;
  assign A5123 = new_A5131_ | new_A5130_;
  assign A5122 = new_A5129_ | new_A5128_;
  assign A5121 = new_A5127_ & new_A5126_;
  assign new_A5120_ = new_B371_;
  assign new_A5119_ = new_B338_;
  assign new_A5118_ = new_B305_;
  assign new_A5117_ = new_B272_;
  assign new_A5116_ = new_B239_;
  assign new_A5115_ = new_A5093_ & new_A5108_;
  assign new_A5114_ = ~new_A5093_ & ~new_A5115_;
  assign new_A5113_ = new_A5093_ | new_A5108_;
  assign new_A5112_ = ~new_A5086_ | ~new_A5087_;
  assign new_A5111_ = new_A5093_ | new_A5108_;
  assign new_A5110_ = ~new_A5109_ & ~new_A5093_;
  assign new_A5109_ = new_A5093_ & new_A5108_;
  assign new_A5108_ = ~new_A5084_ | ~new_A5085_;
  assign new_A5107_ = new_A5085_ & new_A5097_;
  assign new_A5106_ = new_A5086_ | new_A5093_;
  assign new_A5105_ = new_A5086_ | new_A5087_;
  assign new_A5104_ = ~new_A5114_ | ~new_A5113_;
  assign new_A5103_ = new_A5112_ & new_A5105_;
  assign new_A5102_ = new_A5086_ ^ new_A5093_;
  assign new_A5101_ = ~new_A5110_ | ~new_A5111_;
  assign new_A5100_ = ~new_A5085_ ^ new_A5097_;
  assign new_A5099_ = new_A5107_ | new_A5084_;
  assign new_A5098_ = new_A5104_ & new_A5085_;
  assign new_A5097_ = new_A5106_ & new_A5105_;
  assign new_A5096_ = new_A5101_ & new_A5085_;
  assign new_A5095_ = new_A5103_ & new_A5102_;
  assign new_A5094_ = new_A5095_ ^ new_A5085_;
  assign new_A5093_ = new_A5083_ ^ new_A5084_;
  assign A5092 = new_A5093_ & new_A5100_;
  assign A5091 = new_A5093_ & new_A5099_;
  assign A5090 = new_A5098_ | new_A5097_;
  assign A5089 = new_A5096_ | new_A5095_;
  assign A5088 = new_A5094_ & new_A5093_;
  assign new_A5087_ = new_B206_;
  assign new_A5086_ = new_B173_;
  assign new_A5085_ = new_B140_;
  assign new_A5084_ = new_B107_;
  assign new_A5083_ = new_B74_;
  assign new_A5082_ = new_A5060_ & new_A5075_;
  assign new_A5081_ = ~new_A5060_ & ~new_A5082_;
  assign new_A5080_ = new_A5060_ | new_A5075_;
  assign new_A5079_ = ~new_A5053_ | ~new_A5054_;
  assign new_A5078_ = new_A5060_ | new_A5075_;
  assign new_A5077_ = ~new_A5076_ & ~new_A5060_;
  assign new_A5076_ = new_A5060_ & new_A5075_;
  assign new_A5075_ = ~new_A5051_ | ~new_A5052_;
  assign new_A5074_ = new_A5052_ & new_A5064_;
  assign new_A5073_ = new_A5053_ | new_A5060_;
  assign new_A5072_ = new_A5053_ | new_A5054_;
  assign new_A5071_ = ~new_A5081_ | ~new_A5080_;
  assign new_A5070_ = new_A5079_ & new_A5072_;
  assign new_A5069_ = new_A5053_ ^ new_A5060_;
  assign new_A5068_ = ~new_A5077_ | ~new_A5078_;
  assign new_A5067_ = ~new_A5052_ ^ new_A5064_;
  assign new_A5066_ = new_A5074_ | new_A5051_;
  assign new_A5065_ = new_A5071_ & new_A5052_;
  assign new_A5064_ = new_A5073_ & new_A5072_;
  assign new_A5063_ = new_A5068_ & new_A5052_;
  assign new_A5062_ = new_A5070_ & new_A5069_;
  assign new_A5061_ = new_A5062_ ^ new_A5052_;
  assign new_A5060_ = new_A5050_ ^ new_A5051_;
  assign A5059 = new_A5060_ & new_A5067_;
  assign A5058 = new_A5060_ & new_A5066_;
  assign A5057 = new_A5065_ | new_A5064_;
  assign A5056 = new_A5063_ | new_A5062_;
  assign A5055 = new_A5061_ & new_A5060_;
  assign new_A5054_ = new_B41_;
  assign new_A5053_ = new_B8_;
  assign new_A5052_ = new_A9974_;
  assign new_A5051_ = new_A9941_;
  assign new_A5050_ = new_A9908_;
  assign new_A5049_ = new_A5027_ & new_A5042_;
  assign new_A5048_ = ~new_A5027_ & ~new_A5049_;
  assign new_A5047_ = new_A5027_ | new_A5042_;
  assign new_A5046_ = ~new_A5020_ | ~new_A5021_;
  assign new_A5045_ = new_A5027_ | new_A5042_;
  assign new_A5044_ = ~new_A5043_ & ~new_A5027_;
  assign new_A5043_ = new_A5027_ & new_A5042_;
  assign new_A5042_ = ~new_A5018_ | ~new_A5019_;
  assign new_A5041_ = new_A5019_ & new_A5031_;
  assign new_A5040_ = new_A5020_ | new_A5027_;
  assign new_A5039_ = new_A5020_ | new_A5021_;
  assign new_A5038_ = ~new_A5048_ | ~new_A5047_;
  assign new_A5037_ = new_A5046_ & new_A5039_;
  assign new_A5036_ = new_A5020_ ^ new_A5027_;
  assign new_A5035_ = ~new_A5044_ | ~new_A5045_;
  assign new_A5034_ = ~new_A5019_ ^ new_A5031_;
  assign new_A5033_ = new_A5041_ | new_A5018_;
  assign new_A5032_ = new_A5038_ & new_A5019_;
  assign new_A5031_ = new_A5040_ & new_A5039_;
  assign new_A5030_ = new_A5035_ & new_A5019_;
  assign new_A5029_ = new_A5037_ & new_A5036_;
  assign new_A5028_ = new_A5029_ ^ new_A5019_;
  assign new_A5027_ = new_A5017_ ^ new_A5018_;
  assign A5026 = new_A5027_ & new_A5034_;
  assign A5025 = new_A5027_ & new_A5033_;
  assign A5024 = new_A5032_ | new_A5031_;
  assign A5023 = new_A5030_ | new_A5029_;
  assign A5022 = new_A5028_ & new_A5027_;
  assign new_A5021_ = new_A9875_;
  assign new_A5020_ = new_A9842_;
  assign new_A5019_ = new_A9809_;
  assign new_A5018_ = new_A9776_;
  assign new_A5017_ = new_A9743_;
  assign new_A5016_ = new_A4994_ & new_A5009_;
  assign new_A5015_ = ~new_A4994_ & ~new_A5016_;
  assign new_A5014_ = new_A4994_ | new_A5009_;
  assign new_A5013_ = ~new_A4987_ | ~new_A4988_;
  assign new_A5012_ = new_A4994_ | new_A5009_;
  assign new_A5011_ = ~new_A5010_ & ~new_A4994_;
  assign new_A5010_ = new_A4994_ & new_A5009_;
  assign new_A5009_ = ~new_A4985_ | ~new_A4986_;
  assign new_A5008_ = new_A4986_ & new_A4998_;
  assign new_A5007_ = new_A4987_ | new_A4994_;
  assign new_A5006_ = new_A4987_ | new_A4988_;
  assign new_A5005_ = ~new_A5015_ | ~new_A5014_;
  assign new_A5004_ = new_A5013_ & new_A5006_;
  assign new_A5003_ = new_A4987_ ^ new_A4994_;
  assign new_A5002_ = ~new_A5011_ | ~new_A5012_;
  assign new_A5001_ = ~new_A4986_ ^ new_A4998_;
  assign new_A5000_ = new_A5008_ | new_A4985_;
  assign new_A4999_ = new_A5005_ & new_A4986_;
  assign new_A4998_ = new_A5007_ & new_A5006_;
  assign new_A4997_ = new_A5002_ & new_A4986_;
  assign new_A4996_ = new_A5004_ & new_A5003_;
  assign new_A4995_ = new_A4996_ ^ new_A4986_;
  assign new_A4994_ = new_A4984_ ^ new_A4985_;
  assign A4993 = new_A4994_ & new_A5001_;
  assign A4992 = new_A4994_ & new_A5000_;
  assign A4991 = new_A4999_ | new_A4998_;
  assign A4990 = new_A4997_ | new_A4996_;
  assign A4989 = new_A4995_ & new_A4994_;
  assign new_A4988_ = new_A9710_;
  assign new_A4987_ = new_A9677_;
  assign new_A4986_ = new_A9644_;
  assign new_A4985_ = new_A9611_;
  assign new_A4984_ = new_A9578_;
  assign new_A4983_ = new_A4961_ & new_A4976_;
  assign new_A4982_ = ~new_A4961_ & ~new_A4983_;
  assign new_A4981_ = new_A4961_ | new_A4976_;
  assign new_A4980_ = ~new_A4954_ | ~new_A4955_;
  assign new_A4979_ = new_A4961_ | new_A4976_;
  assign new_A4978_ = ~new_A4977_ & ~new_A4961_;
  assign new_A4977_ = new_A4961_ & new_A4976_;
  assign new_A4976_ = ~new_A4952_ | ~new_A4953_;
  assign new_A4975_ = new_A4953_ & new_A4965_;
  assign new_A4974_ = new_A4954_ | new_A4961_;
  assign new_A4973_ = new_A4954_ | new_A4955_;
  assign new_A4972_ = ~new_A4982_ | ~new_A4981_;
  assign new_A4971_ = new_A4980_ & new_A4973_;
  assign new_A4970_ = new_A4954_ ^ new_A4961_;
  assign new_A4969_ = ~new_A4978_ | ~new_A4979_;
  assign new_A4968_ = ~new_A4953_ ^ new_A4965_;
  assign new_A4967_ = new_A4975_ | new_A4952_;
  assign new_A4966_ = new_A4972_ & new_A4953_;
  assign new_A4965_ = new_A4974_ & new_A4973_;
  assign new_A4964_ = new_A4969_ & new_A4953_;
  assign new_A4963_ = new_A4971_ & new_A4970_;
  assign new_A4962_ = new_A4963_ ^ new_A4953_;
  assign new_A4961_ = new_A4951_ ^ new_A4952_;
  assign A4960 = new_A4961_ & new_A4968_;
  assign A4959 = new_A4961_ & new_A4967_;
  assign A4958 = new_A4966_ | new_A4965_;
  assign A4957 = new_A4964_ | new_A4963_;
  assign A4956 = new_A4962_ & new_A4961_;
  assign new_A4955_ = new_A9545_;
  assign new_A4954_ = new_A9512_;
  assign new_A4953_ = new_A9479_;
  assign new_A4952_ = new_A9446_;
  assign new_A4951_ = new_A9413_;
  assign new_A4950_ = new_A4928_ & new_A4943_;
  assign new_A4949_ = ~new_A4928_ & ~new_A4950_;
  assign new_A4948_ = new_A4928_ | new_A4943_;
  assign new_A4947_ = ~new_A4921_ | ~new_A4922_;
  assign new_A4946_ = new_A4928_ | new_A4943_;
  assign new_A4945_ = ~new_A4944_ & ~new_A4928_;
  assign new_A4944_ = new_A4928_ & new_A4943_;
  assign new_A4943_ = ~new_A4919_ | ~new_A4920_;
  assign new_A4942_ = new_A4920_ & new_A4932_;
  assign new_A4941_ = new_A4921_ | new_A4928_;
  assign new_A4940_ = new_A4921_ | new_A4922_;
  assign new_A4939_ = ~new_A4949_ | ~new_A4948_;
  assign new_A4938_ = new_A4947_ & new_A4940_;
  assign new_A4937_ = new_A4921_ ^ new_A4928_;
  assign new_A4936_ = ~new_A4945_ | ~new_A4946_;
  assign new_A4935_ = ~new_A4920_ ^ new_A4932_;
  assign new_A4934_ = new_A4942_ | new_A4919_;
  assign new_A4933_ = new_A4939_ & new_A4920_;
  assign new_A4932_ = new_A4941_ & new_A4940_;
  assign new_A4931_ = new_A4936_ & new_A4920_;
  assign new_A4930_ = new_A4938_ & new_A4937_;
  assign new_A4929_ = new_A4930_ ^ new_A4920_;
  assign new_A4928_ = new_A4918_ ^ new_A4919_;
  assign A4927 = new_A4928_ & new_A4935_;
  assign A4926 = new_A4928_ & new_A4934_;
  assign A4925 = new_A4933_ | new_A4932_;
  assign A4924 = new_A4931_ | new_A4930_;
  assign A4923 = new_A4929_ & new_A4928_;
  assign new_A4922_ = new_A9380_;
  assign new_A4921_ = new_A9347_;
  assign new_A4920_ = new_A9314_;
  assign new_A4919_ = new_A9281_;
  assign new_A4918_ = new_A9248_;
  assign new_A4917_ = new_A4895_ & new_A4910_;
  assign new_A4916_ = ~new_A4895_ & ~new_A4917_;
  assign new_A4915_ = new_A4895_ | new_A4910_;
  assign new_A4914_ = ~new_A4888_ | ~new_A4889_;
  assign new_A4913_ = new_A4895_ | new_A4910_;
  assign new_A4912_ = ~new_A4911_ & ~new_A4895_;
  assign new_A4911_ = new_A4895_ & new_A4910_;
  assign new_A4910_ = ~new_A4886_ | ~new_A4887_;
  assign new_A4909_ = new_A4887_ & new_A4899_;
  assign new_A4908_ = new_A4888_ | new_A4895_;
  assign new_A4907_ = new_A4888_ | new_A4889_;
  assign new_A4906_ = ~new_A4916_ | ~new_A4915_;
  assign new_A4905_ = new_A4914_ & new_A4907_;
  assign new_A4904_ = new_A4888_ ^ new_A4895_;
  assign new_A4903_ = ~new_A4912_ | ~new_A4913_;
  assign new_A4902_ = ~new_A4887_ ^ new_A4899_;
  assign new_A4901_ = new_A4909_ | new_A4886_;
  assign new_A4900_ = new_A4906_ & new_A4887_;
  assign new_A4899_ = new_A4908_ & new_A4907_;
  assign new_A4898_ = new_A4903_ & new_A4887_;
  assign new_A4897_ = new_A4905_ & new_A4904_;
  assign new_A4896_ = new_A4897_ ^ new_A4887_;
  assign new_A4895_ = new_A4885_ ^ new_A4886_;
  assign A4894 = new_A4895_ & new_A4902_;
  assign A4893 = new_A4895_ & new_A4901_;
  assign A4892 = new_A4900_ | new_A4899_;
  assign A4891 = new_A4898_ | new_A4897_;
  assign A4890 = new_A4896_ & new_A4895_;
  assign new_A4889_ = new_A9215_;
  assign new_A4888_ = new_A9182_;
  assign new_A4887_ = new_A9149_;
  assign new_A4886_ = new_A9116_;
  assign new_A4885_ = new_A9083_;
  assign new_A4884_ = new_A4862_ & new_A4877_;
  assign new_A4883_ = ~new_A4862_ & ~new_A4884_;
  assign new_A4882_ = new_A4862_ | new_A4877_;
  assign new_A4881_ = ~new_A4855_ | ~new_A4856_;
  assign new_A4880_ = new_A4862_ | new_A4877_;
  assign new_A4879_ = ~new_A4878_ & ~new_A4862_;
  assign new_A4878_ = new_A4862_ & new_A4877_;
  assign new_A4877_ = ~new_A4853_ | ~new_A4854_;
  assign new_A4876_ = new_A4854_ & new_A4866_;
  assign new_A4875_ = new_A4855_ | new_A4862_;
  assign new_A4874_ = new_A4855_ | new_A4856_;
  assign new_A4873_ = ~new_A4883_ | ~new_A4882_;
  assign new_A4872_ = new_A4881_ & new_A4874_;
  assign new_A4871_ = new_A4855_ ^ new_A4862_;
  assign new_A4870_ = ~new_A4879_ | ~new_A4880_;
  assign new_A4869_ = ~new_A4854_ ^ new_A4866_;
  assign new_A4868_ = new_A4876_ | new_A4853_;
  assign new_A4867_ = new_A4873_ & new_A4854_;
  assign new_A4866_ = new_A4875_ & new_A4874_;
  assign new_A4865_ = new_A4870_ & new_A4854_;
  assign new_A4864_ = new_A4872_ & new_A4871_;
  assign new_A4863_ = new_A4864_ ^ new_A4854_;
  assign new_A4862_ = new_A4852_ ^ new_A4853_;
  assign A4861 = new_A4862_ & new_A4869_;
  assign A4860 = new_A4862_ & new_A4868_;
  assign A4859 = new_A4867_ | new_A4866_;
  assign A4858 = new_A4865_ | new_A4864_;
  assign A4857 = new_A4863_ & new_A4862_;
  assign new_A4856_ = new_A9050_;
  assign new_A4855_ = new_A9017_;
  assign new_A4854_ = new_A8984_;
  assign new_A4853_ = new_A8951_;
  assign new_A4852_ = new_A8918_;
  assign new_A4851_ = new_A4829_ & new_A4844_;
  assign new_A4850_ = ~new_A4829_ & ~new_A4851_;
  assign new_A4849_ = new_A4829_ | new_A4844_;
  assign new_A4848_ = ~new_A4822_ | ~new_A4823_;
  assign new_A4847_ = new_A4829_ | new_A4844_;
  assign new_A4846_ = ~new_A4845_ & ~new_A4829_;
  assign new_A4845_ = new_A4829_ & new_A4844_;
  assign new_A4844_ = ~new_A4820_ | ~new_A4821_;
  assign new_A4843_ = new_A4821_ & new_A4833_;
  assign new_A4842_ = new_A4822_ | new_A4829_;
  assign new_A4841_ = new_A4822_ | new_A4823_;
  assign new_A4840_ = ~new_A4850_ | ~new_A4849_;
  assign new_A4839_ = new_A4848_ & new_A4841_;
  assign new_A4838_ = new_A4822_ ^ new_A4829_;
  assign new_A4837_ = ~new_A4846_ | ~new_A4847_;
  assign new_A4836_ = ~new_A4821_ ^ new_A4833_;
  assign new_A4835_ = new_A4843_ | new_A4820_;
  assign new_A4834_ = new_A4840_ & new_A4821_;
  assign new_A4833_ = new_A4842_ & new_A4841_;
  assign new_A4832_ = new_A4837_ & new_A4821_;
  assign new_A4831_ = new_A4839_ & new_A4838_;
  assign new_A4830_ = new_A4831_ ^ new_A4821_;
  assign new_A4829_ = new_A4819_ ^ new_A4820_;
  assign A4828 = new_A4829_ & new_A4836_;
  assign A4827 = new_A4829_ & new_A4835_;
  assign A4826 = new_A4834_ | new_A4833_;
  assign A4825 = new_A4832_ | new_A4831_;
  assign A4824 = new_A4830_ & new_A4829_;
  assign new_A4823_ = new_A8885_;
  assign new_A4822_ = new_A8852_;
  assign new_A4821_ = new_A8819_;
  assign new_A4820_ = new_A8786_;
  assign new_A4819_ = new_A8753_;
  assign new_A4818_ = new_A4796_ & new_A4811_;
  assign new_A4817_ = ~new_A4796_ & ~new_A4818_;
  assign new_A4816_ = new_A4796_ | new_A4811_;
  assign new_A4815_ = ~new_A4789_ | ~new_A4790_;
  assign new_A4814_ = new_A4796_ | new_A4811_;
  assign new_A4813_ = ~new_A4812_ & ~new_A4796_;
  assign new_A4812_ = new_A4796_ & new_A4811_;
  assign new_A4811_ = ~new_A4787_ | ~new_A4788_;
  assign new_A4810_ = new_A4788_ & new_A4800_;
  assign new_A4809_ = new_A4789_ | new_A4796_;
  assign new_A4808_ = new_A4789_ | new_A4790_;
  assign new_A4807_ = ~new_A4817_ | ~new_A4816_;
  assign new_A4806_ = new_A4815_ & new_A4808_;
  assign new_A4805_ = new_A4789_ ^ new_A4796_;
  assign new_A4804_ = ~new_A4813_ | ~new_A4814_;
  assign new_A4803_ = ~new_A4788_ ^ new_A4800_;
  assign new_A4802_ = new_A4810_ | new_A4787_;
  assign new_A4801_ = new_A4807_ & new_A4788_;
  assign new_A4800_ = new_A4809_ & new_A4808_;
  assign new_A4799_ = new_A4804_ & new_A4788_;
  assign new_A4798_ = new_A4806_ & new_A4805_;
  assign new_A4797_ = new_A4798_ ^ new_A4788_;
  assign new_A4796_ = new_A4786_ ^ new_A4787_;
  assign A4795 = new_A4796_ & new_A4803_;
  assign A4794 = new_A4796_ & new_A4802_;
  assign A4793 = new_A4801_ | new_A4800_;
  assign A4792 = new_A4799_ | new_A4798_;
  assign A4791 = new_A4797_ & new_A4796_;
  assign new_A4790_ = new_A8720_;
  assign new_A4789_ = new_A8687_;
  assign new_A4788_ = new_A8654_;
  assign new_A4787_ = new_A8621_;
  assign new_A4786_ = new_A8588_;
  assign new_A4785_ = new_A4763_ & new_A4778_;
  assign new_A4784_ = ~new_A4763_ & ~new_A4785_;
  assign new_A4783_ = new_A4763_ | new_A4778_;
  assign new_A4782_ = ~new_A4756_ | ~new_A4757_;
  assign new_A4781_ = new_A4763_ | new_A4778_;
  assign new_A4780_ = ~new_A4779_ & ~new_A4763_;
  assign new_A4779_ = new_A4763_ & new_A4778_;
  assign new_A4778_ = ~new_A4754_ | ~new_A4755_;
  assign new_A4777_ = new_A4755_ & new_A4767_;
  assign new_A4776_ = new_A4756_ | new_A4763_;
  assign new_A4775_ = new_A4756_ | new_A4757_;
  assign new_A4774_ = ~new_A4784_ | ~new_A4783_;
  assign new_A4773_ = new_A4782_ & new_A4775_;
  assign new_A4772_ = new_A4756_ ^ new_A4763_;
  assign new_A4771_ = ~new_A4780_ | ~new_A4781_;
  assign new_A4770_ = ~new_A4755_ ^ new_A4767_;
  assign new_A4769_ = new_A4777_ | new_A4754_;
  assign new_A4768_ = new_A4774_ & new_A4755_;
  assign new_A4767_ = new_A4776_ & new_A4775_;
  assign new_A4766_ = new_A4771_ & new_A4755_;
  assign new_A4765_ = new_A4773_ & new_A4772_;
  assign new_A4764_ = new_A4765_ ^ new_A4755_;
  assign new_A4763_ = new_A4753_ ^ new_A4754_;
  assign A4762 = new_A4763_ & new_A4770_;
  assign A4761 = new_A4763_ & new_A4769_;
  assign A4760 = new_A4768_ | new_A4767_;
  assign A4759 = new_A4766_ | new_A4765_;
  assign A4758 = new_A4764_ & new_A4763_;
  assign new_A4757_ = new_A8555_;
  assign new_A4756_ = new_A8522_;
  assign new_A4755_ = new_A8489_;
  assign new_A4754_ = new_A8456_;
  assign new_A4753_ = new_A8423_;
  assign new_A4752_ = new_A4730_ & new_A4745_;
  assign new_A4751_ = ~new_A4730_ & ~new_A4752_;
  assign new_A4750_ = new_A4730_ | new_A4745_;
  assign new_A4749_ = ~new_A4723_ | ~new_A4724_;
  assign new_A4748_ = new_A4730_ | new_A4745_;
  assign new_A4747_ = ~new_A4746_ & ~new_A4730_;
  assign new_A4746_ = new_A4730_ & new_A4745_;
  assign new_A4745_ = ~new_A4721_ | ~new_A4722_;
  assign new_A4744_ = new_A4722_ & new_A4734_;
  assign new_A4743_ = new_A4723_ | new_A4730_;
  assign new_A4742_ = new_A4723_ | new_A4724_;
  assign new_A4741_ = ~new_A4751_ | ~new_A4750_;
  assign new_A4740_ = new_A4749_ & new_A4742_;
  assign new_A4739_ = new_A4723_ ^ new_A4730_;
  assign new_A4738_ = ~new_A4747_ | ~new_A4748_;
  assign new_A4737_ = ~new_A4722_ ^ new_A4734_;
  assign new_A4736_ = new_A4744_ | new_A4721_;
  assign new_A4735_ = new_A4741_ & new_A4722_;
  assign new_A4734_ = new_A4743_ & new_A4742_;
  assign new_A4733_ = new_A4738_ & new_A4722_;
  assign new_A4732_ = new_A4740_ & new_A4739_;
  assign new_A4731_ = new_A4732_ ^ new_A4722_;
  assign new_A4730_ = new_A4720_ ^ new_A4721_;
  assign A4729 = new_A4730_ & new_A4737_;
  assign A4728 = new_A4730_ & new_A4736_;
  assign A4727 = new_A4735_ | new_A4734_;
  assign A4726 = new_A4733_ | new_A4732_;
  assign A4725 = new_A4731_ & new_A4730_;
  assign new_A4724_ = new_A8390_;
  assign new_A4723_ = new_A8357_;
  assign new_A4722_ = new_A8324_;
  assign new_A4721_ = new_A8291_;
  assign new_A4720_ = new_A8258_;
  assign new_A4719_ = new_A4697_ & new_A4712_;
  assign new_A4718_ = ~new_A4697_ & ~new_A4719_;
  assign new_A4717_ = new_A4697_ | new_A4712_;
  assign new_A4716_ = ~new_A4690_ | ~new_A4691_;
  assign new_A4715_ = new_A4697_ | new_A4712_;
  assign new_A4714_ = ~new_A4713_ & ~new_A4697_;
  assign new_A4713_ = new_A4697_ & new_A4712_;
  assign new_A4712_ = ~new_A4688_ | ~new_A4689_;
  assign new_A4711_ = new_A4689_ & new_A4701_;
  assign new_A4710_ = new_A4690_ | new_A4697_;
  assign new_A4709_ = new_A4690_ | new_A4691_;
  assign new_A4708_ = ~new_A4718_ | ~new_A4717_;
  assign new_A4707_ = new_A4716_ & new_A4709_;
  assign new_A4706_ = new_A4690_ ^ new_A4697_;
  assign new_A4705_ = ~new_A4714_ | ~new_A4715_;
  assign new_A4704_ = ~new_A4689_ ^ new_A4701_;
  assign new_A4703_ = new_A4711_ | new_A4688_;
  assign new_A4702_ = new_A4708_ & new_A4689_;
  assign new_A4701_ = new_A4710_ & new_A4709_;
  assign new_A4700_ = new_A4705_ & new_A4689_;
  assign new_A4699_ = new_A4707_ & new_A4706_;
  assign new_A4698_ = new_A4699_ ^ new_A4689_;
  assign new_A4697_ = new_A4687_ ^ new_A4688_;
  assign A4696 = new_A4697_ & new_A4704_;
  assign A4695 = new_A4697_ & new_A4703_;
  assign A4694 = new_A4702_ | new_A4701_;
  assign A4693 = new_A4700_ | new_A4699_;
  assign A4692 = new_A4698_ & new_A4697_;
  assign new_A4691_ = new_A8225_;
  assign new_A4690_ = new_A8192_;
  assign new_A4689_ = new_A8159_;
  assign new_A4688_ = new_A8126_;
  assign new_A4687_ = new_A8093_;
  assign new_A4686_ = new_A4664_ & new_A4679_;
  assign new_A4685_ = ~new_A4664_ & ~new_A4686_;
  assign new_A4684_ = new_A4664_ | new_A4679_;
  assign new_A4683_ = ~new_A4657_ | ~new_A4658_;
  assign new_A4682_ = new_A4664_ | new_A4679_;
  assign new_A4681_ = ~new_A4680_ & ~new_A4664_;
  assign new_A4680_ = new_A4664_ & new_A4679_;
  assign new_A4679_ = ~new_A4655_ | ~new_A4656_;
  assign new_A4678_ = new_A4656_ & new_A4668_;
  assign new_A4677_ = new_A4657_ | new_A4664_;
  assign new_A4676_ = new_A4657_ | new_A4658_;
  assign new_A4675_ = ~new_A4685_ | ~new_A4684_;
  assign new_A4674_ = new_A4683_ & new_A4676_;
  assign new_A4673_ = new_A4657_ ^ new_A4664_;
  assign new_A4672_ = ~new_A4681_ | ~new_A4682_;
  assign new_A4671_ = ~new_A4656_ ^ new_A4668_;
  assign new_A4670_ = new_A4678_ | new_A4655_;
  assign new_A4669_ = new_A4675_ & new_A4656_;
  assign new_A4668_ = new_A4677_ & new_A4676_;
  assign new_A4667_ = new_A4672_ & new_A4656_;
  assign new_A4666_ = new_A4674_ & new_A4673_;
  assign new_A4665_ = new_A4666_ ^ new_A4656_;
  assign new_A4664_ = new_A4654_ ^ new_A4655_;
  assign A4663 = new_A4664_ & new_A4671_;
  assign A4662 = new_A4664_ & new_A4670_;
  assign A4661 = new_A4669_ | new_A4668_;
  assign A4660 = new_A4667_ | new_A4666_;
  assign A4659 = new_A4665_ & new_A4664_;
  assign new_A4658_ = new_A8060_;
  assign new_A4657_ = new_A8027_;
  assign new_A4656_ = new_A7994_;
  assign new_A4655_ = new_A7961_;
  assign new_A4654_ = new_A7928_;
  assign new_A4653_ = new_A4631_ & new_A4646_;
  assign new_A4652_ = ~new_A4631_ & ~new_A4653_;
  assign new_A4651_ = new_A4631_ | new_A4646_;
  assign new_A4650_ = ~new_A4624_ | ~new_A4625_;
  assign new_A4649_ = new_A4631_ | new_A4646_;
  assign new_A4648_ = ~new_A4647_ & ~new_A4631_;
  assign new_A4647_ = new_A4631_ & new_A4646_;
  assign new_A4646_ = ~new_A4622_ | ~new_A4623_;
  assign new_A4645_ = new_A4623_ & new_A4635_;
  assign new_A4644_ = new_A4624_ | new_A4631_;
  assign new_A4643_ = new_A4624_ | new_A4625_;
  assign new_A4642_ = ~new_A4652_ | ~new_A4651_;
  assign new_A4641_ = new_A4650_ & new_A4643_;
  assign new_A4640_ = new_A4624_ ^ new_A4631_;
  assign new_A4639_ = ~new_A4648_ | ~new_A4649_;
  assign new_A4638_ = ~new_A4623_ ^ new_A4635_;
  assign new_A4637_ = new_A4645_ | new_A4622_;
  assign new_A4636_ = new_A4642_ & new_A4623_;
  assign new_A4635_ = new_A4644_ & new_A4643_;
  assign new_A4634_ = new_A4639_ & new_A4623_;
  assign new_A4633_ = new_A4641_ & new_A4640_;
  assign new_A4632_ = new_A4633_ ^ new_A4623_;
  assign new_A4631_ = new_A4621_ ^ new_A4622_;
  assign A4630 = new_A4631_ & new_A4638_;
  assign A4629 = new_A4631_ & new_A4637_;
  assign A4628 = new_A4636_ | new_A4635_;
  assign A4627 = new_A4634_ | new_A4633_;
  assign A4626 = new_A4632_ & new_A4631_;
  assign new_A4625_ = new_A7895_;
  assign new_A4624_ = new_A7862_;
  assign new_A4623_ = new_A7829_;
  assign new_A4622_ = new_A7796_;
  assign new_A4621_ = new_A7763_;
  assign new_A4620_ = new_A4598_ & new_A4613_;
  assign new_A4619_ = ~new_A4598_ & ~new_A4620_;
  assign new_A4618_ = new_A4598_ | new_A4613_;
  assign new_A4617_ = ~new_A4591_ | ~new_A4592_;
  assign new_A4616_ = new_A4598_ | new_A4613_;
  assign new_A4615_ = ~new_A4614_ & ~new_A4598_;
  assign new_A4614_ = new_A4598_ & new_A4613_;
  assign new_A4613_ = ~new_A4589_ | ~new_A4590_;
  assign new_A4612_ = new_A4590_ & new_A4602_;
  assign new_A4611_ = new_A4591_ | new_A4598_;
  assign new_A4610_ = new_A4591_ | new_A4592_;
  assign new_A4609_ = ~new_A4619_ | ~new_A4618_;
  assign new_A4608_ = new_A4617_ & new_A4610_;
  assign new_A4607_ = new_A4591_ ^ new_A4598_;
  assign new_A4606_ = ~new_A4615_ | ~new_A4616_;
  assign new_A4605_ = ~new_A4590_ ^ new_A4602_;
  assign new_A4604_ = new_A4612_ | new_A4589_;
  assign new_A4603_ = new_A4609_ & new_A4590_;
  assign new_A4602_ = new_A4611_ & new_A4610_;
  assign new_A4601_ = new_A4606_ & new_A4590_;
  assign new_A4600_ = new_A4608_ & new_A4607_;
  assign new_A4599_ = new_A4600_ ^ new_A4590_;
  assign new_A4598_ = new_A4588_ ^ new_A4589_;
  assign A4597 = new_A4598_ & new_A4605_;
  assign A4596 = new_A4598_ & new_A4604_;
  assign A4595 = new_A4603_ | new_A4602_;
  assign A4594 = new_A4601_ | new_A4600_;
  assign A4593 = new_A4599_ & new_A4598_;
  assign new_A4592_ = new_A7730_;
  assign new_A4591_ = new_A7697_;
  assign new_A4590_ = new_A7664_;
  assign new_A4589_ = new_A7631_;
  assign new_A4588_ = new_A7598_;
  assign new_A4587_ = new_A4565_ & new_A4580_;
  assign new_A4586_ = ~new_A4565_ & ~new_A4587_;
  assign new_A4585_ = new_A4565_ | new_A4580_;
  assign new_A4584_ = ~new_A4558_ | ~new_A4559_;
  assign new_A4583_ = new_A4565_ | new_A4580_;
  assign new_A4582_ = ~new_A4581_ & ~new_A4565_;
  assign new_A4581_ = new_A4565_ & new_A4580_;
  assign new_A4580_ = ~new_A4556_ | ~new_A4557_;
  assign new_A4579_ = new_A4557_ & new_A4569_;
  assign new_A4578_ = new_A4558_ | new_A4565_;
  assign new_A4577_ = new_A4558_ | new_A4559_;
  assign new_A4576_ = ~new_A4586_ | ~new_A4585_;
  assign new_A4575_ = new_A4584_ & new_A4577_;
  assign new_A4574_ = new_A4558_ ^ new_A4565_;
  assign new_A4573_ = ~new_A4582_ | ~new_A4583_;
  assign new_A4572_ = ~new_A4557_ ^ new_A4569_;
  assign new_A4571_ = new_A4579_ | new_A4556_;
  assign new_A4570_ = new_A4576_ & new_A4557_;
  assign new_A4569_ = new_A4578_ & new_A4577_;
  assign new_A4568_ = new_A4573_ & new_A4557_;
  assign new_A4567_ = new_A4575_ & new_A4574_;
  assign new_A4566_ = new_A4567_ ^ new_A4557_;
  assign new_A4565_ = new_A4555_ ^ new_A4556_;
  assign A4564 = new_A4565_ & new_A4572_;
  assign A4563 = new_A4565_ & new_A4571_;
  assign A4562 = new_A4570_ | new_A4569_;
  assign A4561 = new_A4568_ | new_A4567_;
  assign A4560 = new_A4566_ & new_A4565_;
  assign new_A4559_ = new_A7565_;
  assign new_A4558_ = new_A7532_;
  assign new_A4557_ = new_A7499_;
  assign new_A4556_ = new_A7466_;
  assign new_A4555_ = new_A7433_;
  assign new_A4554_ = new_A4532_ & new_A4547_;
  assign new_A4553_ = ~new_A4532_ & ~new_A4554_;
  assign new_A4552_ = new_A4532_ | new_A4547_;
  assign new_A4551_ = ~new_A4525_ | ~new_A4526_;
  assign new_A4550_ = new_A4532_ | new_A4547_;
  assign new_A4549_ = ~new_A4548_ & ~new_A4532_;
  assign new_A4548_ = new_A4532_ & new_A4547_;
  assign new_A4547_ = ~new_A4523_ | ~new_A4524_;
  assign new_A4546_ = new_A4524_ & new_A4536_;
  assign new_A4545_ = new_A4525_ | new_A4532_;
  assign new_A4544_ = new_A4525_ | new_A4526_;
  assign new_A4543_ = ~new_A4553_ | ~new_A4552_;
  assign new_A4542_ = new_A4551_ & new_A4544_;
  assign new_A4541_ = new_A4525_ ^ new_A4532_;
  assign new_A4540_ = ~new_A4549_ | ~new_A4550_;
  assign new_A4539_ = ~new_A4524_ ^ new_A4536_;
  assign new_A4538_ = new_A4546_ | new_A4523_;
  assign new_A4537_ = new_A4543_ & new_A4524_;
  assign new_A4536_ = new_A4545_ & new_A4544_;
  assign new_A4535_ = new_A4540_ & new_A4524_;
  assign new_A4534_ = new_A4542_ & new_A4541_;
  assign new_A4533_ = new_A4534_ ^ new_A4524_;
  assign new_A4532_ = new_A4522_ ^ new_A4523_;
  assign A4531 = new_A4532_ & new_A4539_;
  assign A4530 = new_A4532_ & new_A4538_;
  assign A4529 = new_A4537_ | new_A4536_;
  assign A4528 = new_A4535_ | new_A4534_;
  assign A4527 = new_A4533_ & new_A4532_;
  assign new_A4526_ = new_A7400_;
  assign new_A4525_ = new_A7367_;
  assign new_A4524_ = new_A7334_;
  assign new_A4523_ = new_A7301_;
  assign new_A4522_ = new_A7268_;
  assign new_A4521_ = new_A4499_ & new_A4514_;
  assign new_A4520_ = ~new_A4499_ & ~new_A4521_;
  assign new_A4519_ = new_A4499_ | new_A4514_;
  assign new_A4518_ = ~new_A4492_ | ~new_A4493_;
  assign new_A4517_ = new_A4499_ | new_A4514_;
  assign new_A4516_ = ~new_A4515_ & ~new_A4499_;
  assign new_A4515_ = new_A4499_ & new_A4514_;
  assign new_A4514_ = ~new_A4490_ | ~new_A4491_;
  assign new_A4513_ = new_A4491_ & new_A4503_;
  assign new_A4512_ = new_A4492_ | new_A4499_;
  assign new_A4511_ = new_A4492_ | new_A4493_;
  assign new_A4510_ = ~new_A4520_ | ~new_A4519_;
  assign new_A4509_ = new_A4518_ & new_A4511_;
  assign new_A4508_ = new_A4492_ ^ new_A4499_;
  assign new_A4507_ = ~new_A4516_ | ~new_A4517_;
  assign new_A4506_ = ~new_A4491_ ^ new_A4503_;
  assign new_A4505_ = new_A4513_ | new_A4490_;
  assign new_A4504_ = new_A4510_ & new_A4491_;
  assign new_A4503_ = new_A4512_ & new_A4511_;
  assign new_A4502_ = new_A4507_ & new_A4491_;
  assign new_A4501_ = new_A4509_ & new_A4508_;
  assign new_A4500_ = new_A4501_ ^ new_A4491_;
  assign new_A4499_ = new_A4489_ ^ new_A4490_;
  assign A4498 = new_A4499_ & new_A4506_;
  assign A4497 = new_A4499_ & new_A4505_;
  assign A4496 = new_A4504_ | new_A4503_;
  assign A4495 = new_A4502_ | new_A4501_;
  assign A4494 = new_A4500_ & new_A4499_;
  assign new_A4493_ = new_A7235_;
  assign new_A4492_ = new_A7202_;
  assign new_A4491_ = new_A7169_;
  assign new_A4490_ = new_A7136_;
  assign new_A4489_ = new_A7103_;
  assign new_A4488_ = new_A4466_ & new_A4481_;
  assign new_A4487_ = ~new_A4466_ & ~new_A4488_;
  assign new_A4486_ = new_A4466_ | new_A4481_;
  assign new_A4485_ = ~new_A4459_ | ~new_A4460_;
  assign new_A4484_ = new_A4466_ | new_A4481_;
  assign new_A4483_ = ~new_A4482_ & ~new_A4466_;
  assign new_A4482_ = new_A4466_ & new_A4481_;
  assign new_A4481_ = ~new_A4457_ | ~new_A4458_;
  assign new_A4480_ = new_A4458_ & new_A4470_;
  assign new_A4479_ = new_A4459_ | new_A4466_;
  assign new_A4478_ = new_A4459_ | new_A4460_;
  assign new_A4477_ = ~new_A4487_ | ~new_A4486_;
  assign new_A4476_ = new_A4485_ & new_A4478_;
  assign new_A4475_ = new_A4459_ ^ new_A4466_;
  assign new_A4474_ = ~new_A4483_ | ~new_A4484_;
  assign new_A4473_ = ~new_A4458_ ^ new_A4470_;
  assign new_A4472_ = new_A4480_ | new_A4457_;
  assign new_A4471_ = new_A4477_ & new_A4458_;
  assign new_A4470_ = new_A4479_ & new_A4478_;
  assign new_A4469_ = new_A4474_ & new_A4458_;
  assign new_A4468_ = new_A4476_ & new_A4475_;
  assign new_A4467_ = new_A4468_ ^ new_A4458_;
  assign new_A4466_ = new_A4456_ ^ new_A4457_;
  assign A4465 = new_A4466_ & new_A4473_;
  assign A4464 = new_A4466_ & new_A4472_;
  assign A4463 = new_A4471_ | new_A4470_;
  assign A4462 = new_A4469_ | new_A4468_;
  assign A4461 = new_A4467_ & new_A4466_;
  assign new_A4460_ = new_A7070_;
  assign new_A4459_ = new_A7037_;
  assign new_A4458_ = new_A7004_;
  assign new_A4457_ = new_A6971_;
  assign new_A4456_ = new_A6938_;
  assign new_A4455_ = new_A4433_ & new_A4448_;
  assign new_A4454_ = ~new_A4433_ & ~new_A4455_;
  assign new_A4453_ = new_A4433_ | new_A4448_;
  assign new_A4452_ = ~new_A4426_ | ~new_A4427_;
  assign new_A4451_ = new_A4433_ | new_A4448_;
  assign new_A4450_ = ~new_A4449_ & ~new_A4433_;
  assign new_A4449_ = new_A4433_ & new_A4448_;
  assign new_A4448_ = ~new_A4424_ | ~new_A4425_;
  assign new_A4447_ = new_A4425_ & new_A4437_;
  assign new_A4446_ = new_A4426_ | new_A4433_;
  assign new_A4445_ = new_A4426_ | new_A4427_;
  assign new_A4444_ = ~new_A4454_ | ~new_A4453_;
  assign new_A4443_ = new_A4452_ & new_A4445_;
  assign new_A4442_ = new_A4426_ ^ new_A4433_;
  assign new_A4441_ = ~new_A4450_ | ~new_A4451_;
  assign new_A4440_ = ~new_A4425_ ^ new_A4437_;
  assign new_A4439_ = new_A4447_ | new_A4424_;
  assign new_A4438_ = new_A4444_ & new_A4425_;
  assign new_A4437_ = new_A4446_ & new_A4445_;
  assign new_A4436_ = new_A4441_ & new_A4425_;
  assign new_A4435_ = new_A4443_ & new_A4442_;
  assign new_A4434_ = new_A4435_ ^ new_A4425_;
  assign new_A4433_ = new_A4423_ ^ new_A4424_;
  assign A4432 = new_A4433_ & new_A4440_;
  assign A4431 = new_A4433_ & new_A4439_;
  assign A4430 = new_A4438_ | new_A4437_;
  assign A4429 = new_A4436_ | new_A4435_;
  assign A4428 = new_A4434_ & new_A4433_;
  assign new_A4427_ = new_B1030_;
  assign new_A4426_ = new_B997_;
  assign new_A4425_ = new_B964_;
  assign new_A4424_ = new_B931_;
  assign new_A4423_ = new_B898_;
  assign new_A4422_ = new_A4400_ & new_A4415_;
  assign new_A4421_ = ~new_A4400_ & ~new_A4422_;
  assign new_A4420_ = new_A4400_ | new_A4415_;
  assign new_A4419_ = ~new_A4393_ | ~new_A4394_;
  assign new_A4418_ = new_A4400_ | new_A4415_;
  assign new_A4417_ = ~new_A4416_ & ~new_A4400_;
  assign new_A4416_ = new_A4400_ & new_A4415_;
  assign new_A4415_ = ~new_A4391_ | ~new_A4392_;
  assign new_A4414_ = new_A4392_ & new_A4404_;
  assign new_A4413_ = new_A4393_ | new_A4400_;
  assign new_A4412_ = new_A4393_ | new_A4394_;
  assign new_A4411_ = ~new_A4421_ | ~new_A4420_;
  assign new_A4410_ = new_A4419_ & new_A4412_;
  assign new_A4409_ = new_A4393_ ^ new_A4400_;
  assign new_A4408_ = ~new_A4417_ | ~new_A4418_;
  assign new_A4407_ = ~new_A4392_ ^ new_A4404_;
  assign new_A4406_ = new_A4414_ | new_A4391_;
  assign new_A4405_ = new_A4411_ & new_A4392_;
  assign new_A4404_ = new_A4413_ & new_A4412_;
  assign new_A4403_ = new_A4408_ & new_A4392_;
  assign new_A4402_ = new_A4410_ & new_A4409_;
  assign new_A4401_ = new_A4402_ ^ new_A4392_;
  assign new_A4400_ = new_A4390_ ^ new_A4391_;
  assign A4399 = new_A4400_ & new_A4407_;
  assign A4398 = new_A4400_ & new_A4406_;
  assign A4397 = new_A4405_ | new_A4404_;
  assign A4396 = new_A4403_ | new_A4402_;
  assign A4395 = new_A4401_ & new_A4400_;
  assign new_A4394_ = new_B865_;
  assign new_A4393_ = new_B832_;
  assign new_A4392_ = new_B799_;
  assign new_A4391_ = new_B766_;
  assign new_A4390_ = new_B733_;
  assign new_A4389_ = new_A4367_ & new_A4382_;
  assign new_A4388_ = ~new_A4367_ & ~new_A4389_;
  assign new_A4387_ = new_A4367_ | new_A4382_;
  assign new_A4386_ = ~new_A4360_ | ~new_A4361_;
  assign new_A4385_ = new_A4367_ | new_A4382_;
  assign new_A4384_ = ~new_A4383_ & ~new_A4367_;
  assign new_A4383_ = new_A4367_ & new_A4382_;
  assign new_A4382_ = ~new_A4358_ | ~new_A4359_;
  assign new_A4381_ = new_A4359_ & new_A4371_;
  assign new_A4380_ = new_A4360_ | new_A4367_;
  assign new_A4379_ = new_A4360_ | new_A4361_;
  assign new_A4378_ = ~new_A4388_ | ~new_A4387_;
  assign new_A4377_ = new_A4386_ & new_A4379_;
  assign new_A4376_ = new_A4360_ ^ new_A4367_;
  assign new_A4375_ = ~new_A4384_ | ~new_A4385_;
  assign new_A4374_ = ~new_A4359_ ^ new_A4371_;
  assign new_A4373_ = new_A4381_ | new_A4358_;
  assign new_A4372_ = new_A4378_ & new_A4359_;
  assign new_A4371_ = new_A4380_ & new_A4379_;
  assign new_A4370_ = new_A4375_ & new_A4359_;
  assign new_A4369_ = new_A4377_ & new_A4376_;
  assign new_A4368_ = new_A4369_ ^ new_A4359_;
  assign new_A4367_ = new_A4357_ ^ new_A4358_;
  assign A4366 = new_A4367_ & new_A4374_;
  assign A4365 = new_A4367_ & new_A4373_;
  assign A4364 = new_A4372_ | new_A4371_;
  assign A4363 = new_A4370_ | new_A4369_;
  assign A4362 = new_A4368_ & new_A4367_;
  assign new_A4361_ = new_B700_;
  assign new_A4360_ = new_B667_;
  assign new_A4359_ = new_B634_;
  assign new_A4358_ = new_B601_;
  assign new_A4357_ = new_B568_;
  assign new_A4356_ = new_A4334_ & new_A4349_;
  assign new_A4355_ = ~new_A4334_ & ~new_A4356_;
  assign new_A4354_ = new_A4334_ | new_A4349_;
  assign new_A4353_ = ~new_A4327_ | ~new_A4328_;
  assign new_A4352_ = new_A4334_ | new_A4349_;
  assign new_A4351_ = ~new_A4350_ & ~new_A4334_;
  assign new_A4350_ = new_A4334_ & new_A4349_;
  assign new_A4349_ = ~new_A4325_ | ~new_A4326_;
  assign new_A4348_ = new_A4326_ & new_A4338_;
  assign new_A4347_ = new_A4327_ | new_A4334_;
  assign new_A4346_ = new_A4327_ | new_A4328_;
  assign new_A4345_ = ~new_A4355_ | ~new_A4354_;
  assign new_A4344_ = new_A4353_ & new_A4346_;
  assign new_A4343_ = new_A4327_ ^ new_A4334_;
  assign new_A4342_ = ~new_A4351_ | ~new_A4352_;
  assign new_A4341_ = ~new_A4326_ ^ new_A4338_;
  assign new_A4340_ = new_A4348_ | new_A4325_;
  assign new_A4339_ = new_A4345_ & new_A4326_;
  assign new_A4338_ = new_A4347_ & new_A4346_;
  assign new_A4337_ = new_A4342_ & new_A4326_;
  assign new_A4336_ = new_A4344_ & new_A4343_;
  assign new_A4335_ = new_A4336_ ^ new_A4326_;
  assign new_A4334_ = new_A4324_ ^ new_A4325_;
  assign A4333 = new_A4334_ & new_A4341_;
  assign A4332 = new_A4334_ & new_A4340_;
  assign A4331 = new_A4339_ | new_A4338_;
  assign A4330 = new_A4337_ | new_A4336_;
  assign A4329 = new_A4335_ & new_A4334_;
  assign new_A4328_ = new_B535_;
  assign new_A4327_ = new_B502_;
  assign new_A4326_ = new_B469_;
  assign new_A4325_ = new_B436_;
  assign new_A4324_ = new_B403_;
  assign new_A4323_ = new_A4301_ & new_A4316_;
  assign new_A4322_ = ~new_A4301_ & ~new_A4323_;
  assign new_A4321_ = new_A4301_ | new_A4316_;
  assign new_A4320_ = ~new_A4294_ | ~new_A4295_;
  assign new_A4319_ = new_A4301_ | new_A4316_;
  assign new_A4318_ = ~new_A4317_ & ~new_A4301_;
  assign new_A4317_ = new_A4301_ & new_A4316_;
  assign new_A4316_ = ~new_A4292_ | ~new_A4293_;
  assign new_A4315_ = new_A4293_ & new_A4305_;
  assign new_A4314_ = new_A4294_ | new_A4301_;
  assign new_A4313_ = new_A4294_ | new_A4295_;
  assign new_A4312_ = ~new_A4322_ | ~new_A4321_;
  assign new_A4311_ = new_A4320_ & new_A4313_;
  assign new_A4310_ = new_A4294_ ^ new_A4301_;
  assign new_A4309_ = ~new_A4318_ | ~new_A4319_;
  assign new_A4308_ = ~new_A4293_ ^ new_A4305_;
  assign new_A4307_ = new_A4315_ | new_A4292_;
  assign new_A4306_ = new_A4312_ & new_A4293_;
  assign new_A4305_ = new_A4314_ & new_A4313_;
  assign new_A4304_ = new_A4309_ & new_A4293_;
  assign new_A4303_ = new_A4311_ & new_A4310_;
  assign new_A4302_ = new_A4303_ ^ new_A4293_;
  assign new_A4301_ = new_A4291_ ^ new_A4292_;
  assign A4300 = new_A4301_ & new_A4308_;
  assign A4299 = new_A4301_ & new_A4307_;
  assign A4298 = new_A4306_ | new_A4305_;
  assign A4297 = new_A4304_ | new_A4303_;
  assign A4296 = new_A4302_ & new_A4301_;
  assign new_A4295_ = new_B370_;
  assign new_A4294_ = new_B337_;
  assign new_A4293_ = new_B304_;
  assign new_A4292_ = new_B271_;
  assign new_A4291_ = new_B238_;
  assign new_A4290_ = new_A4268_ & new_A4283_;
  assign new_A4289_ = ~new_A4268_ & ~new_A4290_;
  assign new_A4288_ = new_A4268_ | new_A4283_;
  assign new_A4287_ = ~new_A4261_ | ~new_A4262_;
  assign new_A4286_ = new_A4268_ | new_A4283_;
  assign new_A4285_ = ~new_A4284_ & ~new_A4268_;
  assign new_A4284_ = new_A4268_ & new_A4283_;
  assign new_A4283_ = ~new_A4259_ | ~new_A4260_;
  assign new_A4282_ = new_A4260_ & new_A4272_;
  assign new_A4281_ = new_A4261_ | new_A4268_;
  assign new_A4280_ = new_A4261_ | new_A4262_;
  assign new_A4279_ = ~new_A4289_ | ~new_A4288_;
  assign new_A4278_ = new_A4287_ & new_A4280_;
  assign new_A4277_ = new_A4261_ ^ new_A4268_;
  assign new_A4276_ = ~new_A4285_ | ~new_A4286_;
  assign new_A4275_ = ~new_A4260_ ^ new_A4272_;
  assign new_A4274_ = new_A4282_ | new_A4259_;
  assign new_A4273_ = new_A4279_ & new_A4260_;
  assign new_A4272_ = new_A4281_ & new_A4280_;
  assign new_A4271_ = new_A4276_ & new_A4260_;
  assign new_A4270_ = new_A4278_ & new_A4277_;
  assign new_A4269_ = new_A4270_ ^ new_A4260_;
  assign new_A4268_ = new_A4258_ ^ new_A4259_;
  assign A4267 = new_A4268_ & new_A4275_;
  assign A4266 = new_A4268_ & new_A4274_;
  assign A4265 = new_A4273_ | new_A4272_;
  assign A4264 = new_A4271_ | new_A4270_;
  assign A4263 = new_A4269_ & new_A4268_;
  assign new_A4262_ = new_B205_;
  assign new_A4261_ = new_B172_;
  assign new_A4260_ = new_B139_;
  assign new_A4259_ = new_B106_;
  assign new_A4258_ = new_B73_;
  assign new_A4257_ = new_A4235_ & new_A4250_;
  assign new_A4256_ = ~new_A4235_ & ~new_A4257_;
  assign new_A4255_ = new_A4235_ | new_A4250_;
  assign new_A4254_ = ~new_A4228_ | ~new_A4229_;
  assign new_A4253_ = new_A4235_ | new_A4250_;
  assign new_A4252_ = ~new_A4251_ & ~new_A4235_;
  assign new_A4251_ = new_A4235_ & new_A4250_;
  assign new_A4250_ = ~new_A4226_ | ~new_A4227_;
  assign new_A4249_ = new_A4227_ & new_A4239_;
  assign new_A4248_ = new_A4228_ | new_A4235_;
  assign new_A4247_ = new_A4228_ | new_A4229_;
  assign new_A4246_ = ~new_A4256_ | ~new_A4255_;
  assign new_A4245_ = new_A4254_ & new_A4247_;
  assign new_A4244_ = new_A4228_ ^ new_A4235_;
  assign new_A4243_ = ~new_A4252_ | ~new_A4253_;
  assign new_A4242_ = ~new_A4227_ ^ new_A4239_;
  assign new_A4241_ = new_A4249_ | new_A4226_;
  assign new_A4240_ = new_A4246_ & new_A4227_;
  assign new_A4239_ = new_A4248_ & new_A4247_;
  assign new_A4238_ = new_A4243_ & new_A4227_;
  assign new_A4237_ = new_A4245_ & new_A4244_;
  assign new_A4236_ = new_A4237_ ^ new_A4227_;
  assign new_A4235_ = new_A4225_ ^ new_A4226_;
  assign A4234 = new_A4235_ & new_A4242_;
  assign A4233 = new_A4235_ & new_A4241_;
  assign A4232 = new_A4240_ | new_A4239_;
  assign A4231 = new_A4238_ | new_A4237_;
  assign A4230 = new_A4236_ & new_A4235_;
  assign new_A4229_ = new_B40_;
  assign new_A4228_ = new_B7_;
  assign new_A4227_ = new_A9973_;
  assign new_A4226_ = new_A9940_;
  assign new_A4225_ = new_A9907_;
  assign new_A4224_ = new_A4202_ & new_A4217_;
  assign new_A4223_ = ~new_A4202_ & ~new_A4224_;
  assign new_A4222_ = new_A4202_ | new_A4217_;
  assign new_A4221_ = ~new_A4195_ | ~new_A4196_;
  assign new_A4220_ = new_A4202_ | new_A4217_;
  assign new_A4219_ = ~new_A4218_ & ~new_A4202_;
  assign new_A4218_ = new_A4202_ & new_A4217_;
  assign new_A4217_ = ~new_A4193_ | ~new_A4194_;
  assign new_A4216_ = new_A4194_ & new_A4206_;
  assign new_A4215_ = new_A4195_ | new_A4202_;
  assign new_A4214_ = new_A4195_ | new_A4196_;
  assign new_A4213_ = ~new_A4223_ | ~new_A4222_;
  assign new_A4212_ = new_A4221_ & new_A4214_;
  assign new_A4211_ = new_A4195_ ^ new_A4202_;
  assign new_A4210_ = ~new_A4219_ | ~new_A4220_;
  assign new_A4209_ = ~new_A4194_ ^ new_A4206_;
  assign new_A4208_ = new_A4216_ | new_A4193_;
  assign new_A4207_ = new_A4213_ & new_A4194_;
  assign new_A4206_ = new_A4215_ & new_A4214_;
  assign new_A4205_ = new_A4210_ & new_A4194_;
  assign new_A4204_ = new_A4212_ & new_A4211_;
  assign new_A4203_ = new_A4204_ ^ new_A4194_;
  assign new_A4202_ = new_A4192_ ^ new_A4193_;
  assign A4201 = new_A4202_ & new_A4209_;
  assign A4200 = new_A4202_ & new_A4208_;
  assign A4199 = new_A4207_ | new_A4206_;
  assign A4198 = new_A4205_ | new_A4204_;
  assign A4197 = new_A4203_ & new_A4202_;
  assign new_A4196_ = new_A9874_;
  assign new_A4195_ = new_A9841_;
  assign new_A4194_ = new_A9808_;
  assign new_A4193_ = new_A9775_;
  assign new_A4192_ = new_A9742_;
  assign new_A4191_ = new_A4169_ & new_A4184_;
  assign new_A4190_ = ~new_A4169_ & ~new_A4191_;
  assign new_A4189_ = new_A4169_ | new_A4184_;
  assign new_A4188_ = ~new_A4162_ | ~new_A4163_;
  assign new_A4187_ = new_A4169_ | new_A4184_;
  assign new_A4186_ = ~new_A4185_ & ~new_A4169_;
  assign new_A4185_ = new_A4169_ & new_A4184_;
  assign new_A4184_ = ~new_A4160_ | ~new_A4161_;
  assign new_A4183_ = new_A4161_ & new_A4173_;
  assign new_A4182_ = new_A4162_ | new_A4169_;
  assign new_A4181_ = new_A4162_ | new_A4163_;
  assign new_A4180_ = ~new_A4190_ | ~new_A4189_;
  assign new_A4179_ = new_A4188_ & new_A4181_;
  assign new_A4178_ = new_A4162_ ^ new_A4169_;
  assign new_A4177_ = ~new_A4186_ | ~new_A4187_;
  assign new_A4176_ = ~new_A4161_ ^ new_A4173_;
  assign new_A4175_ = new_A4183_ | new_A4160_;
  assign new_A4174_ = new_A4180_ & new_A4161_;
  assign new_A4173_ = new_A4182_ & new_A4181_;
  assign new_A4172_ = new_A4177_ & new_A4161_;
  assign new_A4171_ = new_A4179_ & new_A4178_;
  assign new_A4170_ = new_A4171_ ^ new_A4161_;
  assign new_A4169_ = new_A4159_ ^ new_A4160_;
  assign A4168 = new_A4169_ & new_A4176_;
  assign A4167 = new_A4169_ & new_A4175_;
  assign A4166 = new_A4174_ | new_A4173_;
  assign A4165 = new_A4172_ | new_A4171_;
  assign A4164 = new_A4170_ & new_A4169_;
  assign new_A4163_ = new_A9709_;
  assign new_A4162_ = new_A9676_;
  assign new_A4161_ = new_A9643_;
  assign new_A4160_ = new_A9610_;
  assign new_A4159_ = new_A9577_;
  assign new_A4158_ = new_A4136_ & new_A4151_;
  assign new_A4157_ = ~new_A4136_ & ~new_A4158_;
  assign new_A4156_ = new_A4136_ | new_A4151_;
  assign new_A4155_ = ~new_A4129_ | ~new_A4130_;
  assign new_A4154_ = new_A4136_ | new_A4151_;
  assign new_A4153_ = ~new_A4152_ & ~new_A4136_;
  assign new_A4152_ = new_A4136_ & new_A4151_;
  assign new_A4151_ = ~new_A4127_ | ~new_A4128_;
  assign new_A4150_ = new_A4128_ & new_A4140_;
  assign new_A4149_ = new_A4129_ | new_A4136_;
  assign new_A4148_ = new_A4129_ | new_A4130_;
  assign new_A4147_ = ~new_A4157_ | ~new_A4156_;
  assign new_A4146_ = new_A4155_ & new_A4148_;
  assign new_A4145_ = new_A4129_ ^ new_A4136_;
  assign new_A4144_ = ~new_A4153_ | ~new_A4154_;
  assign new_A4143_ = ~new_A4128_ ^ new_A4140_;
  assign new_A4142_ = new_A4150_ | new_A4127_;
  assign new_A4141_ = new_A4147_ & new_A4128_;
  assign new_A4140_ = new_A4149_ & new_A4148_;
  assign new_A4139_ = new_A4144_ & new_A4128_;
  assign new_A4138_ = new_A4146_ & new_A4145_;
  assign new_A4137_ = new_A4138_ ^ new_A4128_;
  assign new_A4136_ = new_A4126_ ^ new_A4127_;
  assign A4135 = new_A4136_ & new_A4143_;
  assign A4134 = new_A4136_ & new_A4142_;
  assign A4133 = new_A4141_ | new_A4140_;
  assign A4132 = new_A4139_ | new_A4138_;
  assign A4131 = new_A4137_ & new_A4136_;
  assign new_A4130_ = new_A9544_;
  assign new_A4129_ = new_A9511_;
  assign new_A4128_ = new_A9478_;
  assign new_A4127_ = new_A9445_;
  assign new_A4126_ = new_A9412_;
  assign new_A4125_ = new_A4103_ & new_A4118_;
  assign new_A4124_ = ~new_A4103_ & ~new_A4125_;
  assign new_A4123_ = new_A4103_ | new_A4118_;
  assign new_A4122_ = ~new_A4096_ | ~new_A4097_;
  assign new_A4121_ = new_A4103_ | new_A4118_;
  assign new_A4120_ = ~new_A4119_ & ~new_A4103_;
  assign new_A4119_ = new_A4103_ & new_A4118_;
  assign new_A4118_ = ~new_A4094_ | ~new_A4095_;
  assign new_A4117_ = new_A4095_ & new_A4107_;
  assign new_A4116_ = new_A4096_ | new_A4103_;
  assign new_A4115_ = new_A4096_ | new_A4097_;
  assign new_A4114_ = ~new_A4124_ | ~new_A4123_;
  assign new_A4113_ = new_A4122_ & new_A4115_;
  assign new_A4112_ = new_A4096_ ^ new_A4103_;
  assign new_A4111_ = ~new_A4120_ | ~new_A4121_;
  assign new_A4110_ = ~new_A4095_ ^ new_A4107_;
  assign new_A4109_ = new_A4117_ | new_A4094_;
  assign new_A4108_ = new_A4114_ & new_A4095_;
  assign new_A4107_ = new_A4116_ & new_A4115_;
  assign new_A4106_ = new_A4111_ & new_A4095_;
  assign new_A4105_ = new_A4113_ & new_A4112_;
  assign new_A4104_ = new_A4105_ ^ new_A4095_;
  assign new_A4103_ = new_A4093_ ^ new_A4094_;
  assign A4102 = new_A4103_ & new_A4110_;
  assign A4101 = new_A4103_ & new_A4109_;
  assign A4100 = new_A4108_ | new_A4107_;
  assign A4099 = new_A4106_ | new_A4105_;
  assign A4098 = new_A4104_ & new_A4103_;
  assign new_A4097_ = new_A9379_;
  assign new_A4096_ = new_A9346_;
  assign new_A4095_ = new_A9313_;
  assign new_A4094_ = new_A9280_;
  assign new_A4093_ = new_A9247_;
  assign new_A4092_ = new_A4070_ & new_A4085_;
  assign new_A4091_ = ~new_A4070_ & ~new_A4092_;
  assign new_A4090_ = new_A4070_ | new_A4085_;
  assign new_A4089_ = ~new_A4063_ | ~new_A4064_;
  assign new_A4088_ = new_A4070_ | new_A4085_;
  assign new_A4087_ = ~new_A4086_ & ~new_A4070_;
  assign new_A4086_ = new_A4070_ & new_A4085_;
  assign new_A4085_ = ~new_A4061_ | ~new_A4062_;
  assign new_A4084_ = new_A4062_ & new_A4074_;
  assign new_A4083_ = new_A4063_ | new_A4070_;
  assign new_A4082_ = new_A4063_ | new_A4064_;
  assign new_A4081_ = ~new_A4091_ | ~new_A4090_;
  assign new_A4080_ = new_A4089_ & new_A4082_;
  assign new_A4079_ = new_A4063_ ^ new_A4070_;
  assign new_A4078_ = ~new_A4087_ | ~new_A4088_;
  assign new_A4077_ = ~new_A4062_ ^ new_A4074_;
  assign new_A4076_ = new_A4084_ | new_A4061_;
  assign new_A4075_ = new_A4081_ & new_A4062_;
  assign new_A4074_ = new_A4083_ & new_A4082_;
  assign new_A4073_ = new_A4078_ & new_A4062_;
  assign new_A4072_ = new_A4080_ & new_A4079_;
  assign new_A4071_ = new_A4072_ ^ new_A4062_;
  assign new_A4070_ = new_A4060_ ^ new_A4061_;
  assign A4069 = new_A4070_ & new_A4077_;
  assign A4068 = new_A4070_ & new_A4076_;
  assign A4067 = new_A4075_ | new_A4074_;
  assign A4066 = new_A4073_ | new_A4072_;
  assign A4065 = new_A4071_ & new_A4070_;
  assign new_A4064_ = new_A9214_;
  assign new_A4063_ = new_A9181_;
  assign new_A4062_ = new_A9148_;
  assign new_A4061_ = new_A9115_;
  assign new_A4060_ = new_A9082_;
  assign new_A4059_ = new_A4037_ & new_A4052_;
  assign new_A4058_ = ~new_A4037_ & ~new_A4059_;
  assign new_A4057_ = new_A4037_ | new_A4052_;
  assign new_A4056_ = ~new_A4030_ | ~new_A4031_;
  assign new_A4055_ = new_A4037_ | new_A4052_;
  assign new_A4054_ = ~new_A4053_ & ~new_A4037_;
  assign new_A4053_ = new_A4037_ & new_A4052_;
  assign new_A4052_ = ~new_A4028_ | ~new_A4029_;
  assign new_A4051_ = new_A4029_ & new_A4041_;
  assign new_A4050_ = new_A4030_ | new_A4037_;
  assign new_A4049_ = new_A4030_ | new_A4031_;
  assign new_A4048_ = ~new_A4058_ | ~new_A4057_;
  assign new_A4047_ = new_A4056_ & new_A4049_;
  assign new_A4046_ = new_A4030_ ^ new_A4037_;
  assign new_A4045_ = ~new_A4054_ | ~new_A4055_;
  assign new_A4044_ = ~new_A4029_ ^ new_A4041_;
  assign new_A4043_ = new_A4051_ | new_A4028_;
  assign new_A4042_ = new_A4048_ & new_A4029_;
  assign new_A4041_ = new_A4050_ & new_A4049_;
  assign new_A4040_ = new_A4045_ & new_A4029_;
  assign new_A4039_ = new_A4047_ & new_A4046_;
  assign new_A4038_ = new_A4039_ ^ new_A4029_;
  assign new_A4037_ = new_A4027_ ^ new_A4028_;
  assign A4036 = new_A4037_ & new_A4044_;
  assign A4035 = new_A4037_ & new_A4043_;
  assign A4034 = new_A4042_ | new_A4041_;
  assign A4033 = new_A4040_ | new_A4039_;
  assign A4032 = new_A4038_ & new_A4037_;
  assign new_A4031_ = new_A9049_;
  assign new_A4030_ = new_A9016_;
  assign new_A4029_ = new_A8983_;
  assign new_A4028_ = new_A8950_;
  assign new_A4027_ = new_A8917_;
  assign new_A4026_ = new_A4004_ & new_A4019_;
  assign new_A4025_ = ~new_A4004_ & ~new_A4026_;
  assign new_A4024_ = new_A4004_ | new_A4019_;
  assign new_A4023_ = ~new_A3997_ | ~new_A3998_;
  assign new_A4022_ = new_A4004_ | new_A4019_;
  assign new_A4021_ = ~new_A4020_ & ~new_A4004_;
  assign new_A4020_ = new_A4004_ & new_A4019_;
  assign new_A4019_ = ~new_A3995_ | ~new_A3996_;
  assign new_A4018_ = new_A3996_ & new_A4008_;
  assign new_A4017_ = new_A3997_ | new_A4004_;
  assign new_A4016_ = new_A3997_ | new_A3998_;
  assign new_A4015_ = ~new_A4025_ | ~new_A4024_;
  assign new_A4014_ = new_A4023_ & new_A4016_;
  assign new_A4013_ = new_A3997_ ^ new_A4004_;
  assign new_A4012_ = ~new_A4021_ | ~new_A4022_;
  assign new_A4011_ = ~new_A3996_ ^ new_A4008_;
  assign new_A4010_ = new_A4018_ | new_A3995_;
  assign new_A4009_ = new_A4015_ & new_A3996_;
  assign new_A4008_ = new_A4017_ & new_A4016_;
  assign new_A4007_ = new_A4012_ & new_A3996_;
  assign new_A4006_ = new_A4014_ & new_A4013_;
  assign new_A4005_ = new_A4006_ ^ new_A3996_;
  assign new_A4004_ = new_A3994_ ^ new_A3995_;
  assign A4003 = new_A4004_ & new_A4011_;
  assign A4002 = new_A4004_ & new_A4010_;
  assign A4001 = new_A4009_ | new_A4008_;
  assign A4000 = new_A4007_ | new_A4006_;
  assign A3999 = new_A4005_ & new_A4004_;
  assign new_A3998_ = new_A8884_;
  assign new_A3997_ = new_A8851_;
  assign new_A3996_ = new_A8818_;
  assign new_A3995_ = new_A8785_;
  assign new_A3994_ = new_A8752_;
  assign new_A3993_ = new_A3971_ & new_A3986_;
  assign new_A3992_ = ~new_A3971_ & ~new_A3993_;
  assign new_A3991_ = new_A3971_ | new_A3986_;
  assign new_A3990_ = ~new_A3964_ | ~new_A3965_;
  assign new_A3989_ = new_A3971_ | new_A3986_;
  assign new_A3988_ = ~new_A3987_ & ~new_A3971_;
  assign new_A3987_ = new_A3971_ & new_A3986_;
  assign new_A3986_ = ~new_A3962_ | ~new_A3963_;
  assign new_A3985_ = new_A3963_ & new_A3975_;
  assign new_A3984_ = new_A3964_ | new_A3971_;
  assign new_A3983_ = new_A3964_ | new_A3965_;
  assign new_A3982_ = ~new_A3992_ | ~new_A3991_;
  assign new_A3981_ = new_A3990_ & new_A3983_;
  assign new_A3980_ = new_A3964_ ^ new_A3971_;
  assign new_A3979_ = ~new_A3988_ | ~new_A3989_;
  assign new_A3978_ = ~new_A3963_ ^ new_A3975_;
  assign new_A3977_ = new_A3985_ | new_A3962_;
  assign new_A3976_ = new_A3982_ & new_A3963_;
  assign new_A3975_ = new_A3984_ & new_A3983_;
  assign new_A3974_ = new_A3979_ & new_A3963_;
  assign new_A3973_ = new_A3981_ & new_A3980_;
  assign new_A3972_ = new_A3973_ ^ new_A3963_;
  assign new_A3971_ = new_A3961_ ^ new_A3962_;
  assign A3970 = new_A3971_ & new_A3978_;
  assign A3969 = new_A3971_ & new_A3977_;
  assign A3968 = new_A3976_ | new_A3975_;
  assign A3967 = new_A3974_ | new_A3973_;
  assign A3966 = new_A3972_ & new_A3971_;
  assign new_A3965_ = new_A8719_;
  assign new_A3964_ = new_A8686_;
  assign new_A3963_ = new_A8653_;
  assign new_A3962_ = new_A8620_;
  assign new_A3961_ = new_A8587_;
  assign new_A3960_ = new_A3938_ & new_A3953_;
  assign new_A3959_ = ~new_A3938_ & ~new_A3960_;
  assign new_A3958_ = new_A3938_ | new_A3953_;
  assign new_A3957_ = ~new_A3931_ | ~new_A3932_;
  assign new_A3956_ = new_A3938_ | new_A3953_;
  assign new_A3955_ = ~new_A3954_ & ~new_A3938_;
  assign new_A3954_ = new_A3938_ & new_A3953_;
  assign new_A3953_ = ~new_A3929_ | ~new_A3930_;
  assign new_A3952_ = new_A3930_ & new_A3942_;
  assign new_A3951_ = new_A3931_ | new_A3938_;
  assign new_A3950_ = new_A3931_ | new_A3932_;
  assign new_A3949_ = ~new_A3959_ | ~new_A3958_;
  assign new_A3948_ = new_A3957_ & new_A3950_;
  assign new_A3947_ = new_A3931_ ^ new_A3938_;
  assign new_A3946_ = ~new_A3955_ | ~new_A3956_;
  assign new_A3945_ = ~new_A3930_ ^ new_A3942_;
  assign new_A3944_ = new_A3952_ | new_A3929_;
  assign new_A3943_ = new_A3949_ & new_A3930_;
  assign new_A3942_ = new_A3951_ & new_A3950_;
  assign new_A3941_ = new_A3946_ & new_A3930_;
  assign new_A3940_ = new_A3948_ & new_A3947_;
  assign new_A3939_ = new_A3940_ ^ new_A3930_;
  assign new_A3938_ = new_A3928_ ^ new_A3929_;
  assign A3937 = new_A3938_ & new_A3945_;
  assign A3936 = new_A3938_ & new_A3944_;
  assign A3935 = new_A3943_ | new_A3942_;
  assign A3934 = new_A3941_ | new_A3940_;
  assign A3933 = new_A3939_ & new_A3938_;
  assign new_A3932_ = new_A8554_;
  assign new_A3931_ = new_A8521_;
  assign new_A3930_ = new_A8488_;
  assign new_A3929_ = new_A8455_;
  assign new_A3928_ = new_A8422_;
  assign new_A3927_ = new_A3905_ & new_A3920_;
  assign new_A3926_ = ~new_A3905_ & ~new_A3927_;
  assign new_A3925_ = new_A3905_ | new_A3920_;
  assign new_A3924_ = ~new_A3898_ | ~new_A3899_;
  assign new_A3923_ = new_A3905_ | new_A3920_;
  assign new_A3922_ = ~new_A3921_ & ~new_A3905_;
  assign new_A3921_ = new_A3905_ & new_A3920_;
  assign new_A3920_ = ~new_A3896_ | ~new_A3897_;
  assign new_A3919_ = new_A3897_ & new_A3909_;
  assign new_A3918_ = new_A3898_ | new_A3905_;
  assign new_A3917_ = new_A3898_ | new_A3899_;
  assign new_A3916_ = ~new_A3926_ | ~new_A3925_;
  assign new_A3915_ = new_A3924_ & new_A3917_;
  assign new_A3914_ = new_A3898_ ^ new_A3905_;
  assign new_A3913_ = ~new_A3922_ | ~new_A3923_;
  assign new_A3912_ = ~new_A3897_ ^ new_A3909_;
  assign new_A3911_ = new_A3919_ | new_A3896_;
  assign new_A3910_ = new_A3916_ & new_A3897_;
  assign new_A3909_ = new_A3918_ & new_A3917_;
  assign new_A3908_ = new_A3913_ & new_A3897_;
  assign new_A3907_ = new_A3915_ & new_A3914_;
  assign new_A3906_ = new_A3907_ ^ new_A3897_;
  assign new_A3905_ = new_A3895_ ^ new_A3896_;
  assign A3904 = new_A3905_ & new_A3912_;
  assign A3903 = new_A3905_ & new_A3911_;
  assign A3902 = new_A3910_ | new_A3909_;
  assign A3901 = new_A3908_ | new_A3907_;
  assign A3900 = new_A3906_ & new_A3905_;
  assign new_A3899_ = new_A8389_;
  assign new_A3898_ = new_A8356_;
  assign new_A3897_ = new_A8323_;
  assign new_A3896_ = new_A8290_;
  assign new_A3895_ = new_A8257_;
  assign new_A3894_ = new_A3872_ & new_A3887_;
  assign new_A3893_ = ~new_A3872_ & ~new_A3894_;
  assign new_A3892_ = new_A3872_ | new_A3887_;
  assign new_A3891_ = ~new_A3865_ | ~new_A3866_;
  assign new_A3890_ = new_A3872_ | new_A3887_;
  assign new_A3889_ = ~new_A3888_ & ~new_A3872_;
  assign new_A3888_ = new_A3872_ & new_A3887_;
  assign new_A3887_ = ~new_A3863_ | ~new_A3864_;
  assign new_A3886_ = new_A3864_ & new_A3876_;
  assign new_A3885_ = new_A3865_ | new_A3872_;
  assign new_A3884_ = new_A3865_ | new_A3866_;
  assign new_A3883_ = ~new_A3893_ | ~new_A3892_;
  assign new_A3882_ = new_A3891_ & new_A3884_;
  assign new_A3881_ = new_A3865_ ^ new_A3872_;
  assign new_A3880_ = ~new_A3889_ | ~new_A3890_;
  assign new_A3879_ = ~new_A3864_ ^ new_A3876_;
  assign new_A3878_ = new_A3886_ | new_A3863_;
  assign new_A3877_ = new_A3883_ & new_A3864_;
  assign new_A3876_ = new_A3885_ & new_A3884_;
  assign new_A3875_ = new_A3880_ & new_A3864_;
  assign new_A3874_ = new_A3882_ & new_A3881_;
  assign new_A3873_ = new_A3874_ ^ new_A3864_;
  assign new_A3872_ = new_A3862_ ^ new_A3863_;
  assign A3871 = new_A3872_ & new_A3879_;
  assign A3870 = new_A3872_ & new_A3878_;
  assign A3869 = new_A3877_ | new_A3876_;
  assign A3868 = new_A3875_ | new_A3874_;
  assign A3867 = new_A3873_ & new_A3872_;
  assign new_A3866_ = new_A8224_;
  assign new_A3865_ = new_A8191_;
  assign new_A3864_ = new_A8158_;
  assign new_A3863_ = new_A8125_;
  assign new_A3862_ = new_A8092_;
  assign new_A3861_ = new_A3839_ & new_A3854_;
  assign new_A3860_ = ~new_A3839_ & ~new_A3861_;
  assign new_A3859_ = new_A3839_ | new_A3854_;
  assign new_A3858_ = ~new_A3832_ | ~new_A3833_;
  assign new_A3857_ = new_A3839_ | new_A3854_;
  assign new_A3856_ = ~new_A3855_ & ~new_A3839_;
  assign new_A3855_ = new_A3839_ & new_A3854_;
  assign new_A3854_ = ~new_A3830_ | ~new_A3831_;
  assign new_A3853_ = new_A3831_ & new_A3843_;
  assign new_A3852_ = new_A3832_ | new_A3839_;
  assign new_A3851_ = new_A3832_ | new_A3833_;
  assign new_A3850_ = ~new_A3860_ | ~new_A3859_;
  assign new_A3849_ = new_A3858_ & new_A3851_;
  assign new_A3848_ = new_A3832_ ^ new_A3839_;
  assign new_A3847_ = ~new_A3856_ | ~new_A3857_;
  assign new_A3846_ = ~new_A3831_ ^ new_A3843_;
  assign new_A3845_ = new_A3853_ | new_A3830_;
  assign new_A3844_ = new_A3850_ & new_A3831_;
  assign new_A3843_ = new_A3852_ & new_A3851_;
  assign new_A3842_ = new_A3847_ & new_A3831_;
  assign new_A3841_ = new_A3849_ & new_A3848_;
  assign new_A3840_ = new_A3841_ ^ new_A3831_;
  assign new_A3839_ = new_A3829_ ^ new_A3830_;
  assign A3838 = new_A3839_ & new_A3846_;
  assign A3837 = new_A3839_ & new_A3845_;
  assign A3836 = new_A3844_ | new_A3843_;
  assign A3835 = new_A3842_ | new_A3841_;
  assign A3834 = new_A3840_ & new_A3839_;
  assign new_A3833_ = new_A8059_;
  assign new_A3832_ = new_A8026_;
  assign new_A3831_ = new_A7993_;
  assign new_A3830_ = new_A7960_;
  assign new_A3829_ = new_A7927_;
  assign new_A3828_ = new_A3806_ & new_A3821_;
  assign new_A3827_ = ~new_A3806_ & ~new_A3828_;
  assign new_A3826_ = new_A3806_ | new_A3821_;
  assign new_A3825_ = ~new_A3799_ | ~new_A3800_;
  assign new_A3824_ = new_A3806_ | new_A3821_;
  assign new_A3823_ = ~new_A3822_ & ~new_A3806_;
  assign new_A3822_ = new_A3806_ & new_A3821_;
  assign new_A3821_ = ~new_A3797_ | ~new_A3798_;
  assign new_A3820_ = new_A3798_ & new_A3810_;
  assign new_A3819_ = new_A3799_ | new_A3806_;
  assign new_A3818_ = new_A3799_ | new_A3800_;
  assign new_A3817_ = ~new_A3827_ | ~new_A3826_;
  assign new_A3816_ = new_A3825_ & new_A3818_;
  assign new_A3815_ = new_A3799_ ^ new_A3806_;
  assign new_A3814_ = ~new_A3823_ | ~new_A3824_;
  assign new_A3813_ = ~new_A3798_ ^ new_A3810_;
  assign new_A3812_ = new_A3820_ | new_A3797_;
  assign new_A3811_ = new_A3817_ & new_A3798_;
  assign new_A3810_ = new_A3819_ & new_A3818_;
  assign new_A3809_ = new_A3814_ & new_A3798_;
  assign new_A3808_ = new_A3816_ & new_A3815_;
  assign new_A3807_ = new_A3808_ ^ new_A3798_;
  assign new_A3806_ = new_A3796_ ^ new_A3797_;
  assign A3805 = new_A3806_ & new_A3813_;
  assign A3804 = new_A3806_ & new_A3812_;
  assign A3803 = new_A3811_ | new_A3810_;
  assign A3802 = new_A3809_ | new_A3808_;
  assign A3801 = new_A3807_ & new_A3806_;
  assign new_A3800_ = new_A7894_;
  assign new_A3799_ = new_A7861_;
  assign new_A3798_ = new_A7828_;
  assign new_A3797_ = new_A7795_;
  assign new_A3796_ = new_A7762_;
  assign new_A3795_ = new_A3773_ & new_A3788_;
  assign new_A3794_ = ~new_A3773_ & ~new_A3795_;
  assign new_A3793_ = new_A3773_ | new_A3788_;
  assign new_A3792_ = ~new_A3766_ | ~new_A3767_;
  assign new_A3791_ = new_A3773_ | new_A3788_;
  assign new_A3790_ = ~new_A3789_ & ~new_A3773_;
  assign new_A3789_ = new_A3773_ & new_A3788_;
  assign new_A3788_ = ~new_A3764_ | ~new_A3765_;
  assign new_A3787_ = new_A3765_ & new_A3777_;
  assign new_A3786_ = new_A3766_ | new_A3773_;
  assign new_A3785_ = new_A3766_ | new_A3767_;
  assign new_A3784_ = ~new_A3794_ | ~new_A3793_;
  assign new_A3783_ = new_A3792_ & new_A3785_;
  assign new_A3782_ = new_A3766_ ^ new_A3773_;
  assign new_A3781_ = ~new_A3790_ | ~new_A3791_;
  assign new_A3780_ = ~new_A3765_ ^ new_A3777_;
  assign new_A3779_ = new_A3787_ | new_A3764_;
  assign new_A3778_ = new_A3784_ & new_A3765_;
  assign new_A3777_ = new_A3786_ & new_A3785_;
  assign new_A3776_ = new_A3781_ & new_A3765_;
  assign new_A3775_ = new_A3783_ & new_A3782_;
  assign new_A3774_ = new_A3775_ ^ new_A3765_;
  assign new_A3773_ = new_A3763_ ^ new_A3764_;
  assign A3772 = new_A3773_ & new_A3780_;
  assign A3771 = new_A3773_ & new_A3779_;
  assign A3770 = new_A3778_ | new_A3777_;
  assign A3769 = new_A3776_ | new_A3775_;
  assign A3768 = new_A3774_ & new_A3773_;
  assign new_A3767_ = new_A7729_;
  assign new_A3766_ = new_A7696_;
  assign new_A3765_ = new_A7663_;
  assign new_A3764_ = new_A7630_;
  assign new_A3763_ = new_A7597_;
  assign new_A3762_ = new_A3740_ & new_A3755_;
  assign new_A3761_ = ~new_A3740_ & ~new_A3762_;
  assign new_A3760_ = new_A3740_ | new_A3755_;
  assign new_A3759_ = ~new_A3733_ | ~new_A3734_;
  assign new_A3758_ = new_A3740_ | new_A3755_;
  assign new_A3757_ = ~new_A3756_ & ~new_A3740_;
  assign new_A3756_ = new_A3740_ & new_A3755_;
  assign new_A3755_ = ~new_A3731_ | ~new_A3732_;
  assign new_A3754_ = new_A3732_ & new_A3744_;
  assign new_A3753_ = new_A3733_ | new_A3740_;
  assign new_A3752_ = new_A3733_ | new_A3734_;
  assign new_A3751_ = ~new_A3761_ | ~new_A3760_;
  assign new_A3750_ = new_A3759_ & new_A3752_;
  assign new_A3749_ = new_A3733_ ^ new_A3740_;
  assign new_A3748_ = ~new_A3757_ | ~new_A3758_;
  assign new_A3747_ = ~new_A3732_ ^ new_A3744_;
  assign new_A3746_ = new_A3754_ | new_A3731_;
  assign new_A3745_ = new_A3751_ & new_A3732_;
  assign new_A3744_ = new_A3753_ & new_A3752_;
  assign new_A3743_ = new_A3748_ & new_A3732_;
  assign new_A3742_ = new_A3750_ & new_A3749_;
  assign new_A3741_ = new_A3742_ ^ new_A3732_;
  assign new_A3740_ = new_A3730_ ^ new_A3731_;
  assign A3739 = new_A3740_ & new_A3747_;
  assign A3738 = new_A3740_ & new_A3746_;
  assign A3737 = new_A3745_ | new_A3744_;
  assign A3736 = new_A3743_ | new_A3742_;
  assign A3735 = new_A3741_ & new_A3740_;
  assign new_A3734_ = new_A7564_;
  assign new_A3733_ = new_A7531_;
  assign new_A3732_ = new_A7498_;
  assign new_A3731_ = new_A7465_;
  assign new_A3730_ = new_A7432_;
  assign new_A3729_ = new_A3707_ & new_A3722_;
  assign new_A3728_ = ~new_A3707_ & ~new_A3729_;
  assign new_A3727_ = new_A3707_ | new_A3722_;
  assign new_A3726_ = ~new_A3700_ | ~new_A3701_;
  assign new_A3725_ = new_A3707_ | new_A3722_;
  assign new_A3724_ = ~new_A3723_ & ~new_A3707_;
  assign new_A3723_ = new_A3707_ & new_A3722_;
  assign new_A3722_ = ~new_A3698_ | ~new_A3699_;
  assign new_A3721_ = new_A3699_ & new_A3711_;
  assign new_A3720_ = new_A3700_ | new_A3707_;
  assign new_A3719_ = new_A3700_ | new_A3701_;
  assign new_A3718_ = ~new_A3728_ | ~new_A3727_;
  assign new_A3717_ = new_A3726_ & new_A3719_;
  assign new_A3716_ = new_A3700_ ^ new_A3707_;
  assign new_A3715_ = ~new_A3724_ | ~new_A3725_;
  assign new_A3714_ = ~new_A3699_ ^ new_A3711_;
  assign new_A3713_ = new_A3721_ | new_A3698_;
  assign new_A3712_ = new_A3718_ & new_A3699_;
  assign new_A3711_ = new_A3720_ & new_A3719_;
  assign new_A3710_ = new_A3715_ & new_A3699_;
  assign new_A3709_ = new_A3717_ & new_A3716_;
  assign new_A3708_ = new_A3709_ ^ new_A3699_;
  assign new_A3707_ = new_A3697_ ^ new_A3698_;
  assign A3706 = new_A3707_ & new_A3714_;
  assign A3705 = new_A3707_ & new_A3713_;
  assign A3704 = new_A3712_ | new_A3711_;
  assign A3703 = new_A3710_ | new_A3709_;
  assign A3702 = new_A3708_ & new_A3707_;
  assign new_A3701_ = new_A7399_;
  assign new_A3700_ = new_A7366_;
  assign new_A3699_ = new_A7333_;
  assign new_A3698_ = new_A7300_;
  assign new_A3697_ = new_A7267_;
  assign new_A3696_ = new_A3674_ & new_A3689_;
  assign new_A3695_ = ~new_A3674_ & ~new_A3696_;
  assign new_A3694_ = new_A3674_ | new_A3689_;
  assign new_A3693_ = ~new_A3667_ | ~new_A3668_;
  assign new_A3692_ = new_A3674_ | new_A3689_;
  assign new_A3691_ = ~new_A3690_ & ~new_A3674_;
  assign new_A3690_ = new_A3674_ & new_A3689_;
  assign new_A3689_ = ~new_A3665_ | ~new_A3666_;
  assign new_A3688_ = new_A3666_ & new_A3678_;
  assign new_A3687_ = new_A3667_ | new_A3674_;
  assign new_A3686_ = new_A3667_ | new_A3668_;
  assign new_A3685_ = ~new_A3695_ | ~new_A3694_;
  assign new_A3684_ = new_A3693_ & new_A3686_;
  assign new_A3683_ = new_A3667_ ^ new_A3674_;
  assign new_A3682_ = ~new_A3691_ | ~new_A3692_;
  assign new_A3681_ = ~new_A3666_ ^ new_A3678_;
  assign new_A3680_ = new_A3688_ | new_A3665_;
  assign new_A3679_ = new_A3685_ & new_A3666_;
  assign new_A3678_ = new_A3687_ & new_A3686_;
  assign new_A3677_ = new_A3682_ & new_A3666_;
  assign new_A3676_ = new_A3684_ & new_A3683_;
  assign new_A3675_ = new_A3676_ ^ new_A3666_;
  assign new_A3674_ = new_A3664_ ^ new_A3665_;
  assign A3673 = new_A3674_ & new_A3681_;
  assign A3672 = new_A3674_ & new_A3680_;
  assign A3671 = new_A3679_ | new_A3678_;
  assign A3670 = new_A3677_ | new_A3676_;
  assign A3669 = new_A3675_ & new_A3674_;
  assign new_A3668_ = new_A7234_;
  assign new_A3667_ = new_A7201_;
  assign new_A3666_ = new_A7168_;
  assign new_A3665_ = new_A7135_;
  assign new_A3664_ = new_A7102_;
  assign new_A3663_ = new_A3641_ & new_A3656_;
  assign new_A3662_ = ~new_A3641_ & ~new_A3663_;
  assign new_A3661_ = new_A3641_ | new_A3656_;
  assign new_A3660_ = ~new_A3634_ | ~new_A3635_;
  assign new_A3659_ = new_A3641_ | new_A3656_;
  assign new_A3658_ = ~new_A3657_ & ~new_A3641_;
  assign new_A3657_ = new_A3641_ & new_A3656_;
  assign new_A3656_ = ~new_A3632_ | ~new_A3633_;
  assign new_A3655_ = new_A3633_ & new_A3645_;
  assign new_A3654_ = new_A3634_ | new_A3641_;
  assign new_A3653_ = new_A3634_ | new_A3635_;
  assign new_A3652_ = ~new_A3662_ | ~new_A3661_;
  assign new_A3651_ = new_A3660_ & new_A3653_;
  assign new_A3650_ = new_A3634_ ^ new_A3641_;
  assign new_A3649_ = ~new_A3658_ | ~new_A3659_;
  assign new_A3648_ = ~new_A3633_ ^ new_A3645_;
  assign new_A3647_ = new_A3655_ | new_A3632_;
  assign new_A3646_ = new_A3652_ & new_A3633_;
  assign new_A3645_ = new_A3654_ & new_A3653_;
  assign new_A3644_ = new_A3649_ & new_A3633_;
  assign new_A3643_ = new_A3651_ & new_A3650_;
  assign new_A3642_ = new_A3643_ ^ new_A3633_;
  assign new_A3641_ = new_A3631_ ^ new_A3632_;
  assign A3640 = new_A3641_ & new_A3648_;
  assign A3639 = new_A3641_ & new_A3647_;
  assign A3638 = new_A3646_ | new_A3645_;
  assign A3637 = new_A3644_ | new_A3643_;
  assign A3636 = new_A3642_ & new_A3641_;
  assign new_A3635_ = new_A7069_;
  assign new_A3634_ = new_A7036_;
  assign new_A3633_ = new_A7003_;
  assign new_A3632_ = new_A6970_;
  assign new_A3631_ = new_A6939_;
  assign new_A3630_ = new_A3608_ & new_A3623_;
  assign new_A3629_ = ~new_A3608_ & ~new_A3630_;
  assign new_A3628_ = new_A3608_ | new_A3623_;
  assign new_A3627_ = ~new_A3601_ | ~new_A3602_;
  assign new_A3626_ = new_A3608_ | new_A3623_;
  assign new_A3625_ = ~new_A3624_ & ~new_A3608_;
  assign new_A3624_ = new_A3608_ & new_A3623_;
  assign new_A3623_ = ~new_A3599_ | ~new_A3600_;
  assign new_A3622_ = new_A3600_ & new_A3612_;
  assign new_A3621_ = new_A3601_ | new_A3608_;
  assign new_A3620_ = new_A3601_ | new_A3602_;
  assign new_A3619_ = ~new_A3629_ | ~new_A3628_;
  assign new_A3618_ = new_A3627_ & new_A3620_;
  assign new_A3617_ = new_A3601_ ^ new_A3608_;
  assign new_A3616_ = ~new_A3625_ | ~new_A3626_;
  assign new_A3615_ = ~new_A3600_ ^ new_A3612_;
  assign new_A3614_ = new_A3622_ | new_A3599_;
  assign new_A3613_ = new_A3619_ & new_A3600_;
  assign new_A3612_ = new_A3621_ & new_A3620_;
  assign new_A3611_ = new_A3616_ & new_A3600_;
  assign new_A3610_ = new_A3618_ & new_A3617_;
  assign new_A3609_ = new_A3610_ ^ new_A3600_;
  assign new_A3608_ = new_A3598_ ^ new_A3599_;
  assign A3607 = new_A3608_ & new_A3615_;
  assign A3606 = new_A3608_ & new_A3614_;
  assign A3605 = new_A3613_ | new_A3612_;
  assign A3604 = new_A3611_ | new_A3610_;
  assign A3603 = new_A3609_ & new_A3608_;
  assign new_A3602_ = new_B1029_;
  assign new_A3601_ = new_B996_;
  assign new_A3600_ = new_B963_;
  assign new_A3599_ = new_B930_;
  assign new_A3598_ = new_B897_;
  assign new_A3597_ = new_A3575_ & new_A3590_;
  assign new_A3596_ = ~new_A3575_ & ~new_A3597_;
  assign new_A3595_ = new_A3575_ | new_A3590_;
  assign new_A3594_ = ~new_A3568_ | ~new_A3569_;
  assign new_A3593_ = new_A3575_ | new_A3590_;
  assign new_A3592_ = ~new_A3591_ & ~new_A3575_;
  assign new_A3591_ = new_A3575_ & new_A3590_;
  assign new_A3590_ = ~new_A3566_ | ~new_A3567_;
  assign new_A3589_ = new_A3567_ & new_A3579_;
  assign new_A3588_ = new_A3568_ | new_A3575_;
  assign new_A3587_ = new_A3568_ | new_A3569_;
  assign new_A3586_ = ~new_A3596_ | ~new_A3595_;
  assign new_A3585_ = new_A3594_ & new_A3587_;
  assign new_A3584_ = new_A3568_ ^ new_A3575_;
  assign new_A3583_ = ~new_A3592_ | ~new_A3593_;
  assign new_A3582_ = ~new_A3567_ ^ new_A3579_;
  assign new_A3581_ = new_A3589_ | new_A3566_;
  assign new_A3580_ = new_A3586_ & new_A3567_;
  assign new_A3579_ = new_A3588_ & new_A3587_;
  assign new_A3578_ = new_A3583_ & new_A3567_;
  assign new_A3577_ = new_A3585_ & new_A3584_;
  assign new_A3576_ = new_A3577_ ^ new_A3567_;
  assign new_A3575_ = new_A3565_ ^ new_A3566_;
  assign A3574 = new_A3575_ & new_A3582_;
  assign A3573 = new_A3575_ & new_A3581_;
  assign A3572 = new_A3580_ | new_A3579_;
  assign A3571 = new_A3578_ | new_A3577_;
  assign A3570 = new_A3576_ & new_A3575_;
  assign new_A3569_ = new_B864_;
  assign new_A3568_ = new_B831_;
  assign new_A3567_ = new_B798_;
  assign new_A3566_ = new_B765_;
  assign new_A3565_ = new_B732_;
  assign new_A3564_ = new_A3542_ & new_A3557_;
  assign new_A3563_ = ~new_A3542_ & ~new_A3564_;
  assign new_A3562_ = new_A3542_ | new_A3557_;
  assign new_A3561_ = ~new_A3535_ | ~new_A3536_;
  assign new_A3560_ = new_A3542_ | new_A3557_;
  assign new_A3559_ = ~new_A3558_ & ~new_A3542_;
  assign new_A3558_ = new_A3542_ & new_A3557_;
  assign new_A3557_ = ~new_A3533_ | ~new_A3534_;
  assign new_A3556_ = new_A3534_ & new_A3546_;
  assign new_A3555_ = new_A3535_ | new_A3542_;
  assign new_A3554_ = new_A3535_ | new_A3536_;
  assign new_A3553_ = ~new_A3563_ | ~new_A3562_;
  assign new_A3552_ = new_A3561_ & new_A3554_;
  assign new_A3551_ = new_A3535_ ^ new_A3542_;
  assign new_A3550_ = ~new_A3559_ | ~new_A3560_;
  assign new_A3549_ = ~new_A3534_ ^ new_A3546_;
  assign new_A3548_ = new_A3556_ | new_A3533_;
  assign new_A3547_ = new_A3553_ & new_A3534_;
  assign new_A3546_ = new_A3555_ & new_A3554_;
  assign new_A3545_ = new_A3550_ & new_A3534_;
  assign new_A3544_ = new_A3552_ & new_A3551_;
  assign new_A3543_ = new_A3544_ ^ new_A3534_;
  assign new_A3542_ = new_A3532_ ^ new_A3533_;
  assign A3541 = new_A3542_ & new_A3549_;
  assign A3540 = new_A3542_ & new_A3548_;
  assign A3539 = new_A3547_ | new_A3546_;
  assign A3538 = new_A3545_ | new_A3544_;
  assign A3537 = new_A3543_ & new_A3542_;
  assign new_A3536_ = new_B699_;
  assign new_A3535_ = new_B666_;
  assign new_A3534_ = new_B633_;
  assign new_A3533_ = new_B600_;
  assign new_A3532_ = new_B567_;
  assign new_A3531_ = new_A3509_ & new_A3524_;
  assign new_A3530_ = ~new_A3509_ & ~new_A3531_;
  assign new_A3529_ = new_A3509_ | new_A3524_;
  assign new_A3528_ = ~new_A3502_ | ~new_A3503_;
  assign new_A3527_ = new_A3509_ | new_A3524_;
  assign new_A3526_ = ~new_A3525_ & ~new_A3509_;
  assign new_A3525_ = new_A3509_ & new_A3524_;
  assign new_A3524_ = ~new_A3500_ | ~new_A3501_;
  assign new_A3523_ = new_A3501_ & new_A3513_;
  assign new_A3522_ = new_A3502_ | new_A3509_;
  assign new_A3521_ = new_A3502_ | new_A3503_;
  assign new_A3520_ = ~new_A3530_ | ~new_A3529_;
  assign new_A3519_ = new_A3528_ & new_A3521_;
  assign new_A3518_ = new_A3502_ ^ new_A3509_;
  assign new_A3517_ = ~new_A3526_ | ~new_A3527_;
  assign new_A3516_ = ~new_A3501_ ^ new_A3513_;
  assign new_A3515_ = new_A3523_ | new_A3500_;
  assign new_A3514_ = new_A3520_ & new_A3501_;
  assign new_A3513_ = new_A3522_ & new_A3521_;
  assign new_A3512_ = new_A3517_ & new_A3501_;
  assign new_A3511_ = new_A3519_ & new_A3518_;
  assign new_A3510_ = new_A3511_ ^ new_A3501_;
  assign new_A3509_ = new_A3499_ ^ new_A3500_;
  assign A3508 = new_A3509_ & new_A3516_;
  assign A3507 = new_A3509_ & new_A3515_;
  assign A3506 = new_A3514_ | new_A3513_;
  assign A3505 = new_A3512_ | new_A3511_;
  assign A3504 = new_A3510_ & new_A3509_;
  assign new_A3503_ = new_B534_;
  assign new_A3502_ = new_B501_;
  assign new_A3501_ = new_B468_;
  assign new_A3500_ = new_B435_;
  assign new_A3499_ = new_B402_;
  assign new_A3498_ = new_A3476_ & new_A3491_;
  assign new_A3497_ = ~new_A3476_ & ~new_A3498_;
  assign new_A3496_ = new_A3476_ | new_A3491_;
  assign new_A3495_ = ~new_A3469_ | ~new_A3470_;
  assign new_A3494_ = new_A3476_ | new_A3491_;
  assign new_A3493_ = ~new_A3492_ & ~new_A3476_;
  assign new_A3492_ = new_A3476_ & new_A3491_;
  assign new_A3491_ = ~new_A3467_ | ~new_A3468_;
  assign new_A3490_ = new_A3468_ & new_A3480_;
  assign new_A3489_ = new_A3469_ | new_A3476_;
  assign new_A3488_ = new_A3469_ | new_A3470_;
  assign new_A3487_ = ~new_A3497_ | ~new_A3496_;
  assign new_A3486_ = new_A3495_ & new_A3488_;
  assign new_A3485_ = new_A3469_ ^ new_A3476_;
  assign new_A3484_ = ~new_A3493_ | ~new_A3494_;
  assign new_A3483_ = ~new_A3468_ ^ new_A3480_;
  assign new_A3482_ = new_A3490_ | new_A3467_;
  assign new_A3481_ = new_A3487_ & new_A3468_;
  assign new_A3480_ = new_A3489_ & new_A3488_;
  assign new_A3479_ = new_A3484_ & new_A3468_;
  assign new_A3478_ = new_A3486_ & new_A3485_;
  assign new_A3477_ = new_A3478_ ^ new_A3468_;
  assign new_A3476_ = new_A3466_ ^ new_A3467_;
  assign A3475 = new_A3476_ & new_A3483_;
  assign A3474 = new_A3476_ & new_A3482_;
  assign A3473 = new_A3481_ | new_A3480_;
  assign A3472 = new_A3479_ | new_A3478_;
  assign A3471 = new_A3477_ & new_A3476_;
  assign new_A3470_ = new_B369_;
  assign new_A3469_ = new_B336_;
  assign new_A3468_ = new_B303_;
  assign new_A3467_ = new_B270_;
  assign new_A3466_ = new_B237_;
  assign new_A3465_ = new_A3443_ & new_A3458_;
  assign new_A3464_ = ~new_A3443_ & ~new_A3465_;
  assign new_A3463_ = new_A3443_ | new_A3458_;
  assign new_A3462_ = ~new_A3436_ | ~new_A3437_;
  assign new_A3461_ = new_A3443_ | new_A3458_;
  assign new_A3460_ = ~new_A3459_ & ~new_A3443_;
  assign new_A3459_ = new_A3443_ & new_A3458_;
  assign new_A3458_ = ~new_A3434_ | ~new_A3435_;
  assign new_A3457_ = new_A3435_ & new_A3447_;
  assign new_A3456_ = new_A3436_ | new_A3443_;
  assign new_A3455_ = new_A3436_ | new_A3437_;
  assign new_A3454_ = ~new_A3464_ | ~new_A3463_;
  assign new_A3453_ = new_A3462_ & new_A3455_;
  assign new_A3452_ = new_A3436_ ^ new_A3443_;
  assign new_A3451_ = ~new_A3460_ | ~new_A3461_;
  assign new_A3450_ = ~new_A3435_ ^ new_A3447_;
  assign new_A3449_ = new_A3457_ | new_A3434_;
  assign new_A3448_ = new_A3454_ & new_A3435_;
  assign new_A3447_ = new_A3456_ & new_A3455_;
  assign new_A3446_ = new_A3451_ & new_A3435_;
  assign new_A3445_ = new_A3453_ & new_A3452_;
  assign new_A3444_ = new_A3445_ ^ new_A3435_;
  assign new_A3443_ = new_A3433_ ^ new_A3434_;
  assign A3442 = new_A3443_ & new_A3450_;
  assign A3441 = new_A3443_ & new_A3449_;
  assign A3440 = new_A3448_ | new_A3447_;
  assign A3439 = new_A3446_ | new_A3445_;
  assign A3438 = new_A3444_ & new_A3443_;
  assign new_A3437_ = new_B204_;
  assign new_A3436_ = new_B171_;
  assign new_A3435_ = new_B138_;
  assign new_A3434_ = new_B105_;
  assign new_A3433_ = new_B72_;
  assign new_A3432_ = new_A3410_ & new_A3425_;
  assign new_A3431_ = ~new_A3410_ & ~new_A3432_;
  assign new_A3430_ = new_A3410_ | new_A3425_;
  assign new_A3429_ = ~new_A3403_ | ~new_A3404_;
  assign new_A3428_ = new_A3410_ | new_A3425_;
  assign new_A3427_ = ~new_A3426_ & ~new_A3410_;
  assign new_A3426_ = new_A3410_ & new_A3425_;
  assign new_A3425_ = ~new_A3401_ | ~new_A3402_;
  assign new_A3424_ = new_A3402_ & new_A3414_;
  assign new_A3423_ = new_A3403_ | new_A3410_;
  assign new_A3422_ = new_A3403_ | new_A3404_;
  assign new_A3421_ = ~new_A3431_ | ~new_A3430_;
  assign new_A3420_ = new_A3429_ & new_A3422_;
  assign new_A3419_ = new_A3403_ ^ new_A3410_;
  assign new_A3418_ = ~new_A3427_ | ~new_A3428_;
  assign new_A3417_ = ~new_A3402_ ^ new_A3414_;
  assign new_A3416_ = new_A3424_ | new_A3401_;
  assign new_A3415_ = new_A3421_ & new_A3402_;
  assign new_A3414_ = new_A3423_ & new_A3422_;
  assign new_A3413_ = new_A3418_ & new_A3402_;
  assign new_A3412_ = new_A3420_ & new_A3419_;
  assign new_A3411_ = new_A3412_ ^ new_A3402_;
  assign new_A3410_ = new_A3400_ ^ new_A3401_;
  assign A3409 = new_A3410_ & new_A3417_;
  assign A3408 = new_A3410_ & new_A3416_;
  assign A3407 = new_A3415_ | new_A3414_;
  assign A3406 = new_A3413_ | new_A3412_;
  assign A3405 = new_A3411_ & new_A3410_;
  assign new_A3404_ = new_B39_;
  assign new_A3403_ = new_B6_;
  assign new_A3402_ = new_A9972_;
  assign new_A3401_ = new_A9939_;
  assign new_A3400_ = new_A9906_;
  assign new_A3399_ = new_A3377_ & new_A3392_;
  assign new_A3398_ = ~new_A3377_ & ~new_A3399_;
  assign new_A3397_ = new_A3377_ | new_A3392_;
  assign new_A3396_ = ~new_A3370_ | ~new_A3371_;
  assign new_A3395_ = new_A3377_ | new_A3392_;
  assign new_A3394_ = ~new_A3393_ & ~new_A3377_;
  assign new_A3393_ = new_A3377_ & new_A3392_;
  assign new_A3392_ = ~new_A3368_ | ~new_A3369_;
  assign new_A3391_ = new_A3369_ & new_A3381_;
  assign new_A3390_ = new_A3370_ | new_A3377_;
  assign new_A3389_ = new_A3370_ | new_A3371_;
  assign new_A3388_ = ~new_A3398_ | ~new_A3397_;
  assign new_A3387_ = new_A3396_ & new_A3389_;
  assign new_A3386_ = new_A3370_ ^ new_A3377_;
  assign new_A3385_ = ~new_A3394_ | ~new_A3395_;
  assign new_A3384_ = ~new_A3369_ ^ new_A3381_;
  assign new_A3383_ = new_A3391_ | new_A3368_;
  assign new_A3382_ = new_A3388_ & new_A3369_;
  assign new_A3381_ = new_A3390_ & new_A3389_;
  assign new_A3380_ = new_A3385_ & new_A3369_;
  assign new_A3379_ = new_A3387_ & new_A3386_;
  assign new_A3378_ = new_A3379_ ^ new_A3369_;
  assign new_A3377_ = new_A3367_ ^ new_A3368_;
  assign A3376 = new_A3377_ & new_A3384_;
  assign A3375 = new_A3377_ & new_A3383_;
  assign A3374 = new_A3382_ | new_A3381_;
  assign A3373 = new_A3380_ | new_A3379_;
  assign A3372 = new_A3378_ & new_A3377_;
  assign new_A3371_ = new_A9873_;
  assign new_A3370_ = new_A9840_;
  assign new_A3369_ = new_A9807_;
  assign new_A3368_ = new_A9774_;
  assign new_A3367_ = new_A9741_;
  assign new_A3366_ = new_A3344_ & new_A3359_;
  assign new_A3365_ = ~new_A3344_ & ~new_A3366_;
  assign new_A3364_ = new_A3344_ | new_A3359_;
  assign new_A3363_ = ~new_A3337_ | ~new_A3338_;
  assign new_A3362_ = new_A3344_ | new_A3359_;
  assign new_A3361_ = ~new_A3360_ & ~new_A3344_;
  assign new_A3360_ = new_A3344_ & new_A3359_;
  assign new_A3359_ = ~new_A3335_ | ~new_A3336_;
  assign new_A3358_ = new_A3336_ & new_A3348_;
  assign new_A3357_ = new_A3337_ | new_A3344_;
  assign new_A3356_ = new_A3337_ | new_A3338_;
  assign new_A3355_ = ~new_A3365_ | ~new_A3364_;
  assign new_A3354_ = new_A3363_ & new_A3356_;
  assign new_A3353_ = new_A3337_ ^ new_A3344_;
  assign new_A3352_ = ~new_A3361_ | ~new_A3362_;
  assign new_A3351_ = ~new_A3336_ ^ new_A3348_;
  assign new_A3350_ = new_A3358_ | new_A3335_;
  assign new_A3349_ = new_A3355_ & new_A3336_;
  assign new_A3348_ = new_A3357_ & new_A3356_;
  assign new_A3347_ = new_A3352_ & new_A3336_;
  assign new_A3346_ = new_A3354_ & new_A3353_;
  assign new_A3345_ = new_A3346_ ^ new_A3336_;
  assign new_A3344_ = new_A3334_ ^ new_A3335_;
  assign A3343 = new_A3344_ & new_A3351_;
  assign A3342 = new_A3344_ & new_A3350_;
  assign A3341 = new_A3349_ | new_A3348_;
  assign A3340 = new_A3347_ | new_A3346_;
  assign A3339 = new_A3345_ & new_A3344_;
  assign new_A3338_ = new_A9708_;
  assign new_A3337_ = new_A9675_;
  assign new_A3336_ = new_A9642_;
  assign new_A3335_ = new_A9609_;
  assign new_A3334_ = new_A9576_;
  assign new_A3333_ = new_A3311_ & new_A3326_;
  assign new_A3332_ = ~new_A3311_ & ~new_A3333_;
  assign new_A3331_ = new_A3311_ | new_A3326_;
  assign new_A3330_ = ~new_A3304_ | ~new_A3305_;
  assign new_A3329_ = new_A3311_ | new_A3326_;
  assign new_A3328_ = ~new_A3327_ & ~new_A3311_;
  assign new_A3327_ = new_A3311_ & new_A3326_;
  assign new_A3326_ = ~new_A3302_ | ~new_A3303_;
  assign new_A3325_ = new_A3303_ & new_A3315_;
  assign new_A3324_ = new_A3304_ | new_A3311_;
  assign new_A3323_ = new_A3304_ | new_A3305_;
  assign new_A3322_ = ~new_A3332_ | ~new_A3331_;
  assign new_A3321_ = new_A3330_ & new_A3323_;
  assign new_A3320_ = new_A3304_ ^ new_A3311_;
  assign new_A3319_ = ~new_A3328_ | ~new_A3329_;
  assign new_A3318_ = ~new_A3303_ ^ new_A3315_;
  assign new_A3317_ = new_A3325_ | new_A3302_;
  assign new_A3316_ = new_A3322_ & new_A3303_;
  assign new_A3315_ = new_A3324_ & new_A3323_;
  assign new_A3314_ = new_A3319_ & new_A3303_;
  assign new_A3313_ = new_A3321_ & new_A3320_;
  assign new_A3312_ = new_A3313_ ^ new_A3303_;
  assign new_A3311_ = new_A3301_ ^ new_A3302_;
  assign A3310 = new_A3311_ & new_A3318_;
  assign A3309 = new_A3311_ & new_A3317_;
  assign A3308 = new_A3316_ | new_A3315_;
  assign A3307 = new_A3314_ | new_A3313_;
  assign A3306 = new_A3312_ & new_A3311_;
  assign new_A3305_ = new_A9543_;
  assign new_A3304_ = new_A9510_;
  assign new_A3303_ = new_A9477_;
  assign new_A3302_ = new_A9444_;
  assign new_A3301_ = new_A9411_;
  assign new_A3300_ = new_A3278_ & new_A3293_;
  assign new_A3299_ = ~new_A3278_ & ~new_A3300_;
  assign new_A3298_ = new_A3278_ | new_A3293_;
  assign new_A3297_ = ~new_A3271_ | ~new_A3272_;
  assign new_A3296_ = new_A3278_ | new_A3293_;
  assign new_A3295_ = ~new_A3294_ & ~new_A3278_;
  assign new_A3294_ = new_A3278_ & new_A3293_;
  assign new_A3293_ = ~new_A3269_ | ~new_A3270_;
  assign new_A3292_ = new_A3270_ & new_A3282_;
  assign new_A3291_ = new_A3271_ | new_A3278_;
  assign new_A3290_ = new_A3271_ | new_A3272_;
  assign new_A3289_ = ~new_A3299_ | ~new_A3298_;
  assign new_A3288_ = new_A3297_ & new_A3290_;
  assign new_A3287_ = new_A3271_ ^ new_A3278_;
  assign new_A3286_ = ~new_A3295_ | ~new_A3296_;
  assign new_A3285_ = ~new_A3270_ ^ new_A3282_;
  assign new_A3284_ = new_A3292_ | new_A3269_;
  assign new_A3283_ = new_A3289_ & new_A3270_;
  assign new_A3282_ = new_A3291_ & new_A3290_;
  assign new_A3281_ = new_A3286_ & new_A3270_;
  assign new_A3280_ = new_A3288_ & new_A3287_;
  assign new_A3279_ = new_A3280_ ^ new_A3270_;
  assign new_A3278_ = new_A3268_ ^ new_A3269_;
  assign A3277 = new_A3278_ & new_A3285_;
  assign A3276 = new_A3278_ & new_A3284_;
  assign A3275 = new_A3283_ | new_A3282_;
  assign A3274 = new_A3281_ | new_A3280_;
  assign A3273 = new_A3279_ & new_A3278_;
  assign new_A3272_ = new_A9378_;
  assign new_A3271_ = new_A9345_;
  assign new_A3270_ = new_A9312_;
  assign new_A3269_ = new_A9279_;
  assign new_A3268_ = new_A9246_;
  assign new_A3267_ = new_A3245_ & new_A3260_;
  assign new_A3266_ = ~new_A3245_ & ~new_A3267_;
  assign new_A3265_ = new_A3245_ | new_A3260_;
  assign new_A3264_ = ~new_A3238_ | ~new_A3239_;
  assign new_A3263_ = new_A3245_ | new_A3260_;
  assign new_A3262_ = ~new_A3261_ & ~new_A3245_;
  assign new_A3261_ = new_A3245_ & new_A3260_;
  assign new_A3260_ = ~new_A3236_ | ~new_A3237_;
  assign new_A3259_ = new_A3237_ & new_A3249_;
  assign new_A3258_ = new_A3238_ | new_A3245_;
  assign new_A3257_ = new_A3238_ | new_A3239_;
  assign new_A3256_ = ~new_A3266_ | ~new_A3265_;
  assign new_A3255_ = new_A3264_ & new_A3257_;
  assign new_A3254_ = new_A3238_ ^ new_A3245_;
  assign new_A3253_ = ~new_A3262_ | ~new_A3263_;
  assign new_A3252_ = ~new_A3237_ ^ new_A3249_;
  assign new_A3251_ = new_A3259_ | new_A3236_;
  assign new_A3250_ = new_A3256_ & new_A3237_;
  assign new_A3249_ = new_A3258_ & new_A3257_;
  assign new_A3248_ = new_A3253_ & new_A3237_;
  assign new_A3247_ = new_A3255_ & new_A3254_;
  assign new_A3246_ = new_A3247_ ^ new_A3237_;
  assign new_A3245_ = new_A3235_ ^ new_A3236_;
  assign A3244 = new_A3245_ & new_A3252_;
  assign A3243 = new_A3245_ & new_A3251_;
  assign A3242 = new_A3250_ | new_A3249_;
  assign A3241 = new_A3248_ | new_A3247_;
  assign A3240 = new_A3246_ & new_A3245_;
  assign new_A3239_ = new_A9213_;
  assign new_A3238_ = new_A9180_;
  assign new_A3237_ = new_A9147_;
  assign new_A3236_ = new_A9114_;
  assign new_A3235_ = new_A9081_;
  assign new_A3234_ = new_A3212_ & new_A3227_;
  assign new_A3233_ = ~new_A3212_ & ~new_A3234_;
  assign new_A3232_ = new_A3212_ | new_A3227_;
  assign new_A3231_ = ~new_A3205_ | ~new_A3206_;
  assign new_A3230_ = new_A3212_ | new_A3227_;
  assign new_A3229_ = ~new_A3228_ & ~new_A3212_;
  assign new_A3228_ = new_A3212_ & new_A3227_;
  assign new_A3227_ = ~new_A3203_ | ~new_A3204_;
  assign new_A3226_ = new_A3204_ & new_A3216_;
  assign new_A3225_ = new_A3205_ | new_A3212_;
  assign new_A3224_ = new_A3205_ | new_A3206_;
  assign new_A3223_ = ~new_A3233_ | ~new_A3232_;
  assign new_A3222_ = new_A3231_ & new_A3224_;
  assign new_A3221_ = new_A3205_ ^ new_A3212_;
  assign new_A3220_ = ~new_A3229_ | ~new_A3230_;
  assign new_A3219_ = ~new_A3204_ ^ new_A3216_;
  assign new_A3218_ = new_A3226_ | new_A3203_;
  assign new_A3217_ = new_A3223_ & new_A3204_;
  assign new_A3216_ = new_A3225_ & new_A3224_;
  assign new_A3215_ = new_A3220_ & new_A3204_;
  assign new_A3214_ = new_A3222_ & new_A3221_;
  assign new_A3213_ = new_A3214_ ^ new_A3204_;
  assign new_A3212_ = new_A3202_ ^ new_A3203_;
  assign A3211 = new_A3212_ & new_A3219_;
  assign A3210 = new_A3212_ & new_A3218_;
  assign A3209 = new_A3217_ | new_A3216_;
  assign A3208 = new_A3215_ | new_A3214_;
  assign A3207 = new_A3213_ & new_A3212_;
  assign new_A3206_ = new_A9048_;
  assign new_A3205_ = new_A9015_;
  assign new_A3204_ = new_A8982_;
  assign new_A3203_ = new_A8949_;
  assign new_A3202_ = new_A8916_;
  assign new_A3201_ = new_A3179_ & new_A3194_;
  assign new_A3200_ = ~new_A3179_ & ~new_A3201_;
  assign new_A3199_ = new_A3179_ | new_A3194_;
  assign new_A3198_ = ~new_A3172_ | ~new_A3173_;
  assign new_A3197_ = new_A3179_ | new_A3194_;
  assign new_A3196_ = ~new_A3195_ & ~new_A3179_;
  assign new_A3195_ = new_A3179_ & new_A3194_;
  assign new_A3194_ = ~new_A3170_ | ~new_A3171_;
  assign new_A3193_ = new_A3171_ & new_A3183_;
  assign new_A3192_ = new_A3172_ | new_A3179_;
  assign new_A3191_ = new_A3172_ | new_A3173_;
  assign new_A3190_ = ~new_A3200_ | ~new_A3199_;
  assign new_A3189_ = new_A3198_ & new_A3191_;
  assign new_A3188_ = new_A3172_ ^ new_A3179_;
  assign new_A3187_ = ~new_A3196_ | ~new_A3197_;
  assign new_A3186_ = ~new_A3171_ ^ new_A3183_;
  assign new_A3185_ = new_A3193_ | new_A3170_;
  assign new_A3184_ = new_A3190_ & new_A3171_;
  assign new_A3183_ = new_A3192_ & new_A3191_;
  assign new_A3182_ = new_A3187_ & new_A3171_;
  assign new_A3181_ = new_A3189_ & new_A3188_;
  assign new_A3180_ = new_A3181_ ^ new_A3171_;
  assign new_A3179_ = new_A3169_ ^ new_A3170_;
  assign A3178 = new_A3179_ & new_A3186_;
  assign A3177 = new_A3179_ & new_A3185_;
  assign A3176 = new_A3184_ | new_A3183_;
  assign A3175 = new_A3182_ | new_A3181_;
  assign A3174 = new_A3180_ & new_A3179_;
  assign new_A3173_ = new_A8883_;
  assign new_A3172_ = new_A8850_;
  assign new_A3171_ = new_A8817_;
  assign new_A3170_ = new_A8784_;
  assign new_A3169_ = new_A8751_;
  assign new_A3168_ = new_A3146_ & new_A3161_;
  assign new_A3167_ = ~new_A3146_ & ~new_A3168_;
  assign new_A3166_ = new_A3146_ | new_A3161_;
  assign new_A3165_ = ~new_A3139_ | ~new_A3140_;
  assign new_A3164_ = new_A3146_ | new_A3161_;
  assign new_A3163_ = ~new_A3162_ & ~new_A3146_;
  assign new_A3162_ = new_A3146_ & new_A3161_;
  assign new_A3161_ = ~new_A3137_ | ~new_A3138_;
  assign new_A3160_ = new_A3138_ & new_A3150_;
  assign new_A3159_ = new_A3139_ | new_A3146_;
  assign new_A3158_ = new_A3139_ | new_A3140_;
  assign new_A3157_ = ~new_A3167_ | ~new_A3166_;
  assign new_A3156_ = new_A3165_ & new_A3158_;
  assign new_A3155_ = new_A3139_ ^ new_A3146_;
  assign new_A3154_ = ~new_A3163_ | ~new_A3164_;
  assign new_A3153_ = ~new_A3138_ ^ new_A3150_;
  assign new_A3152_ = new_A3160_ | new_A3137_;
  assign new_A3151_ = new_A3157_ & new_A3138_;
  assign new_A3150_ = new_A3159_ & new_A3158_;
  assign new_A3149_ = new_A3154_ & new_A3138_;
  assign new_A3148_ = new_A3156_ & new_A3155_;
  assign new_A3147_ = new_A3148_ ^ new_A3138_;
  assign new_A3146_ = new_A3136_ ^ new_A3137_;
  assign A3145 = new_A3146_ & new_A3153_;
  assign A3144 = new_A3146_ & new_A3152_;
  assign A3143 = new_A3151_ | new_A3150_;
  assign A3142 = new_A3149_ | new_A3148_;
  assign A3141 = new_A3147_ & new_A3146_;
  assign new_A3140_ = new_A8718_;
  assign new_A3139_ = new_A8685_;
  assign new_A3138_ = new_A8652_;
  assign new_A3137_ = new_A8619_;
  assign new_A3136_ = new_A8586_;
  assign new_A3135_ = new_A3113_ & new_A3128_;
  assign new_A3134_ = ~new_A3113_ & ~new_A3135_;
  assign new_A3133_ = new_A3113_ | new_A3128_;
  assign new_A3132_ = ~new_A3106_ | ~new_A3107_;
  assign new_A3131_ = new_A3113_ | new_A3128_;
  assign new_A3130_ = ~new_A3129_ & ~new_A3113_;
  assign new_A3129_ = new_A3113_ & new_A3128_;
  assign new_A3128_ = ~new_A3104_ | ~new_A3105_;
  assign new_A3127_ = new_A3105_ & new_A3117_;
  assign new_A3126_ = new_A3106_ | new_A3113_;
  assign new_A3125_ = new_A3106_ | new_A3107_;
  assign new_A3124_ = ~new_A3134_ | ~new_A3133_;
  assign new_A3123_ = new_A3132_ & new_A3125_;
  assign new_A3122_ = new_A3106_ ^ new_A3113_;
  assign new_A3121_ = ~new_A3130_ | ~new_A3131_;
  assign new_A3120_ = ~new_A3105_ ^ new_A3117_;
  assign new_A3119_ = new_A3127_ | new_A3104_;
  assign new_A3118_ = new_A3124_ & new_A3105_;
  assign new_A3117_ = new_A3126_ & new_A3125_;
  assign new_A3116_ = new_A3121_ & new_A3105_;
  assign new_A3115_ = new_A3123_ & new_A3122_;
  assign new_A3114_ = new_A3115_ ^ new_A3105_;
  assign new_A3113_ = new_A3103_ ^ new_A3104_;
  assign A3112 = new_A3113_ & new_A3120_;
  assign A3111 = new_A3113_ & new_A3119_;
  assign A3110 = new_A3118_ | new_A3117_;
  assign A3109 = new_A3116_ | new_A3115_;
  assign A3108 = new_A3114_ & new_A3113_;
  assign new_A3107_ = new_A8553_;
  assign new_A3106_ = new_A8520_;
  assign new_A3105_ = new_A8487_;
  assign new_A3104_ = new_A8454_;
  assign new_A3103_ = new_A8421_;
  assign new_A3102_ = new_A3080_ & new_A3095_;
  assign new_A3101_ = ~new_A3080_ & ~new_A3102_;
  assign new_A3100_ = new_A3080_ | new_A3095_;
  assign new_A3099_ = ~new_A3073_ | ~new_A3074_;
  assign new_A3098_ = new_A3080_ | new_A3095_;
  assign new_A3097_ = ~new_A3096_ & ~new_A3080_;
  assign new_A3096_ = new_A3080_ & new_A3095_;
  assign new_A3095_ = ~new_A3071_ | ~new_A3072_;
  assign new_A3094_ = new_A3072_ & new_A3084_;
  assign new_A3093_ = new_A3073_ | new_A3080_;
  assign new_A3092_ = new_A3073_ | new_A3074_;
  assign new_A3091_ = ~new_A3101_ | ~new_A3100_;
  assign new_A3090_ = new_A3099_ & new_A3092_;
  assign new_A3089_ = new_A3073_ ^ new_A3080_;
  assign new_A3088_ = ~new_A3097_ | ~new_A3098_;
  assign new_A3087_ = ~new_A3072_ ^ new_A3084_;
  assign new_A3086_ = new_A3094_ | new_A3071_;
  assign new_A3085_ = new_A3091_ & new_A3072_;
  assign new_A3084_ = new_A3093_ & new_A3092_;
  assign new_A3083_ = new_A3088_ & new_A3072_;
  assign new_A3082_ = new_A3090_ & new_A3089_;
  assign new_A3081_ = new_A3082_ ^ new_A3072_;
  assign new_A3080_ = new_A3070_ ^ new_A3071_;
  assign A3079 = new_A3080_ & new_A3087_;
  assign A3078 = new_A3080_ & new_A3086_;
  assign A3077 = new_A3085_ | new_A3084_;
  assign A3076 = new_A3083_ | new_A3082_;
  assign A3075 = new_A3081_ & new_A3080_;
  assign new_A3074_ = new_A8388_;
  assign new_A3073_ = new_A8355_;
  assign new_A3072_ = new_A8322_;
  assign new_A3071_ = new_A8289_;
  assign new_A3070_ = new_A8256_;
  assign new_A3069_ = new_A3047_ & new_A3062_;
  assign new_A3068_ = ~new_A3047_ & ~new_A3069_;
  assign new_A3067_ = new_A3047_ | new_A3062_;
  assign new_A3066_ = ~new_A3040_ | ~new_A3041_;
  assign new_A3065_ = new_A3047_ | new_A3062_;
  assign new_A3064_ = ~new_A3063_ & ~new_A3047_;
  assign new_A3063_ = new_A3047_ & new_A3062_;
  assign new_A3062_ = ~new_A3038_ | ~new_A3039_;
  assign new_A3061_ = new_A3039_ & new_A3051_;
  assign new_A3060_ = new_A3040_ | new_A3047_;
  assign new_A3059_ = new_A3040_ | new_A3041_;
  assign new_A3058_ = ~new_A3068_ | ~new_A3067_;
  assign new_A3057_ = new_A3066_ & new_A3059_;
  assign new_A3056_ = new_A3040_ ^ new_A3047_;
  assign new_A3055_ = ~new_A3064_ | ~new_A3065_;
  assign new_A3054_ = ~new_A3039_ ^ new_A3051_;
  assign new_A3053_ = new_A3061_ | new_A3038_;
  assign new_A3052_ = new_A3058_ & new_A3039_;
  assign new_A3051_ = new_A3060_ & new_A3059_;
  assign new_A3050_ = new_A3055_ & new_A3039_;
  assign new_A3049_ = new_A3057_ & new_A3056_;
  assign new_A3048_ = new_A3049_ ^ new_A3039_;
  assign new_A3047_ = new_A3037_ ^ new_A3038_;
  assign A3046 = new_A3047_ & new_A3054_;
  assign A3045 = new_A3047_ & new_A3053_;
  assign A3044 = new_A3052_ | new_A3051_;
  assign A3043 = new_A3050_ | new_A3049_;
  assign A3042 = new_A3048_ & new_A3047_;
  assign new_A3041_ = new_A8223_;
  assign new_A3040_ = new_A8190_;
  assign new_A3039_ = new_A8157_;
  assign new_A3038_ = new_A8124_;
  assign new_A3037_ = new_A8091_;
  assign new_A3036_ = new_A3014_ & new_A3029_;
  assign new_A3035_ = ~new_A3014_ & ~new_A3036_;
  assign new_A3034_ = new_A3014_ | new_A3029_;
  assign new_A3033_ = ~new_A3007_ | ~new_A3008_;
  assign new_A3032_ = new_A3014_ | new_A3029_;
  assign new_A3031_ = ~new_A3030_ & ~new_A3014_;
  assign new_A3030_ = new_A3014_ & new_A3029_;
  assign new_A3029_ = ~new_A3005_ | ~new_A3006_;
  assign new_A3028_ = new_A3006_ & new_A3018_;
  assign new_A3027_ = new_A3007_ | new_A3014_;
  assign new_A3026_ = new_A3007_ | new_A3008_;
  assign new_A3025_ = ~new_A3035_ | ~new_A3034_;
  assign new_A3024_ = new_A3033_ & new_A3026_;
  assign new_A3023_ = new_A3007_ ^ new_A3014_;
  assign new_A3022_ = ~new_A3031_ | ~new_A3032_;
  assign new_A3021_ = ~new_A3006_ ^ new_A3018_;
  assign new_A3020_ = new_A3028_ | new_A3005_;
  assign new_A3019_ = new_A3025_ & new_A3006_;
  assign new_A3018_ = new_A3027_ & new_A3026_;
  assign new_A3017_ = new_A3022_ & new_A3006_;
  assign new_A3016_ = new_A3024_ & new_A3023_;
  assign new_A3015_ = new_A3016_ ^ new_A3006_;
  assign new_A3014_ = new_A3004_ ^ new_A3005_;
  assign A3013 = new_A3014_ & new_A3021_;
  assign A3012 = new_A3014_ & new_A3020_;
  assign A3011 = new_A3019_ | new_A3018_;
  assign A3010 = new_A3017_ | new_A3016_;
  assign A3009 = new_A3015_ & new_A3014_;
  assign new_A3008_ = new_A8058_;
  assign new_A3007_ = new_A8025_;
  assign new_A3006_ = new_A7992_;
  assign new_A3005_ = new_A7959_;
  assign new_A3004_ = new_A7926_;
  assign new_A3003_ = new_A2981_ & new_A2996_;
  assign new_A3002_ = ~new_A2981_ & ~new_A3003_;
  assign new_A3001_ = new_A2981_ | new_A2996_;
  assign new_A3000_ = ~new_A2974_ | ~new_A2975_;
  assign new_A2999_ = new_A2981_ | new_A2996_;
  assign new_A2998_ = ~new_A2997_ & ~new_A2981_;
  assign new_A2997_ = new_A2981_ & new_A2996_;
  assign new_A2996_ = ~new_A2972_ | ~new_A2973_;
  assign new_A2995_ = new_A2973_ & new_A2985_;
  assign new_A2994_ = new_A2974_ | new_A2981_;
  assign new_A2993_ = new_A2974_ | new_A2975_;
  assign new_A2992_ = ~new_A3002_ | ~new_A3001_;
  assign new_A2991_ = new_A3000_ & new_A2993_;
  assign new_A2990_ = new_A2974_ ^ new_A2981_;
  assign new_A2989_ = ~new_A2998_ | ~new_A2999_;
  assign new_A2988_ = ~new_A2973_ ^ new_A2985_;
  assign new_A2987_ = new_A2995_ | new_A2972_;
  assign new_A2986_ = new_A2992_ & new_A2973_;
  assign new_A2985_ = new_A2994_ & new_A2993_;
  assign new_A2984_ = new_A2989_ & new_A2973_;
  assign new_A2983_ = new_A2991_ & new_A2990_;
  assign new_A2982_ = new_A2983_ ^ new_A2973_;
  assign new_A2981_ = new_A2971_ ^ new_A2972_;
  assign A2980 = new_A2981_ & new_A2988_;
  assign A2979 = new_A2981_ & new_A2987_;
  assign A2978 = new_A2986_ | new_A2985_;
  assign A2977 = new_A2984_ | new_A2983_;
  assign A2976 = new_A2982_ & new_A2981_;
  assign new_A2975_ = new_A7893_;
  assign new_A2974_ = new_A7860_;
  assign new_A2973_ = new_A7827_;
  assign new_A2972_ = new_A7794_;
  assign new_A2971_ = new_A7761_;
  assign new_A2970_ = new_A2948_ & new_A2963_;
  assign new_A2969_ = ~new_A2948_ & ~new_A2970_;
  assign new_A2968_ = new_A2948_ | new_A2963_;
  assign new_A2967_ = ~new_A2941_ | ~new_A2942_;
  assign new_A2966_ = new_A2948_ | new_A2963_;
  assign new_A2965_ = ~new_A2964_ & ~new_A2948_;
  assign new_A2964_ = new_A2948_ & new_A2963_;
  assign new_A2963_ = ~new_A2939_ | ~new_A2940_;
  assign new_A2962_ = new_A2940_ & new_A2952_;
  assign new_A2961_ = new_A2941_ | new_A2948_;
  assign new_A2960_ = new_A2941_ | new_A2942_;
  assign new_A2959_ = ~new_A2969_ | ~new_A2968_;
  assign new_A2958_ = new_A2967_ & new_A2960_;
  assign new_A2957_ = new_A2941_ ^ new_A2948_;
  assign new_A2956_ = ~new_A2965_ | ~new_A2966_;
  assign new_A2955_ = ~new_A2940_ ^ new_A2952_;
  assign new_A2954_ = new_A2962_ | new_A2939_;
  assign new_A2953_ = new_A2959_ & new_A2940_;
  assign new_A2952_ = new_A2961_ & new_A2960_;
  assign new_A2951_ = new_A2956_ & new_A2940_;
  assign new_A2950_ = new_A2958_ & new_A2957_;
  assign new_A2949_ = new_A2950_ ^ new_A2940_;
  assign new_A2948_ = new_A2938_ ^ new_A2939_;
  assign A2947 = new_A2948_ & new_A2955_;
  assign A2946 = new_A2948_ & new_A2954_;
  assign A2945 = new_A2953_ | new_A2952_;
  assign A2944 = new_A2951_ | new_A2950_;
  assign A2943 = new_A2949_ & new_A2948_;
  assign new_A2942_ = new_A7728_;
  assign new_A2941_ = new_A7695_;
  assign new_A2940_ = new_A7662_;
  assign new_A2939_ = new_A7629_;
  assign new_A2938_ = new_A7596_;
  assign new_A2937_ = new_A2915_ & new_A2930_;
  assign new_A2936_ = ~new_A2915_ & ~new_A2937_;
  assign new_A2935_ = new_A2915_ | new_A2930_;
  assign new_A2934_ = ~new_A2908_ | ~new_A2909_;
  assign new_A2933_ = new_A2915_ | new_A2930_;
  assign new_A2932_ = ~new_A2931_ & ~new_A2915_;
  assign new_A2931_ = new_A2915_ & new_A2930_;
  assign new_A2930_ = ~new_A2906_ | ~new_A2907_;
  assign new_A2929_ = new_A2907_ & new_A2919_;
  assign new_A2928_ = new_A2908_ | new_A2915_;
  assign new_A2927_ = new_A2908_ | new_A2909_;
  assign new_A2926_ = ~new_A2936_ | ~new_A2935_;
  assign new_A2925_ = new_A2934_ & new_A2927_;
  assign new_A2924_ = new_A2908_ ^ new_A2915_;
  assign new_A2923_ = ~new_A2932_ | ~new_A2933_;
  assign new_A2922_ = ~new_A2907_ ^ new_A2919_;
  assign new_A2921_ = new_A2929_ | new_A2906_;
  assign new_A2920_ = new_A2926_ & new_A2907_;
  assign new_A2919_ = new_A2928_ & new_A2927_;
  assign new_A2918_ = new_A2923_ & new_A2907_;
  assign new_A2917_ = new_A2925_ & new_A2924_;
  assign new_A2916_ = new_A2917_ ^ new_A2907_;
  assign new_A2915_ = new_A2905_ ^ new_A2906_;
  assign A2914 = new_A2915_ & new_A2922_;
  assign A2913 = new_A2915_ & new_A2921_;
  assign A2912 = new_A2920_ | new_A2919_;
  assign A2911 = new_A2918_ | new_A2917_;
  assign A2910 = new_A2916_ & new_A2915_;
  assign new_A2909_ = new_A7563_;
  assign new_A2908_ = new_A7530_;
  assign new_A2907_ = new_A7497_;
  assign new_A2906_ = new_A7464_;
  assign new_A2905_ = new_A7431_;
  assign new_A2904_ = new_A2882_ & new_A2897_;
  assign new_A2903_ = ~new_A2882_ & ~new_A2904_;
  assign new_A2902_ = new_A2882_ | new_A2897_;
  assign new_A2901_ = ~new_A2875_ | ~new_A2876_;
  assign new_A2900_ = new_A2882_ | new_A2897_;
  assign new_A2899_ = ~new_A2898_ & ~new_A2882_;
  assign new_A2898_ = new_A2882_ & new_A2897_;
  assign new_A2897_ = ~new_A2873_ | ~new_A2874_;
  assign new_A2896_ = new_A2874_ & new_A2886_;
  assign new_A2895_ = new_A2875_ | new_A2882_;
  assign new_A2894_ = new_A2875_ | new_A2876_;
  assign new_A2893_ = ~new_A2903_ | ~new_A2902_;
  assign new_A2892_ = new_A2901_ & new_A2894_;
  assign new_A2891_ = new_A2875_ ^ new_A2882_;
  assign new_A2890_ = ~new_A2899_ | ~new_A2900_;
  assign new_A2889_ = ~new_A2874_ ^ new_A2886_;
  assign new_A2888_ = new_A2896_ | new_A2873_;
  assign new_A2887_ = new_A2893_ & new_A2874_;
  assign new_A2886_ = new_A2895_ & new_A2894_;
  assign new_A2885_ = new_A2890_ & new_A2874_;
  assign new_A2884_ = new_A2892_ & new_A2891_;
  assign new_A2883_ = new_A2884_ ^ new_A2874_;
  assign new_A2882_ = new_A2872_ ^ new_A2873_;
  assign A2881 = new_A2882_ & new_A2889_;
  assign A2880 = new_A2882_ & new_A2888_;
  assign A2879 = new_A2887_ | new_A2886_;
  assign A2878 = new_A2885_ | new_A2884_;
  assign A2877 = new_A2883_ & new_A2882_;
  assign new_A2876_ = new_A7398_;
  assign new_A2875_ = new_A7365_;
  assign new_A2874_ = new_A7332_;
  assign new_A2873_ = new_A7299_;
  assign new_A2872_ = new_A7266_;
  assign new_A2871_ = new_A2849_ & new_A2864_;
  assign new_A2870_ = ~new_A2849_ & ~new_A2871_;
  assign new_A2869_ = new_A2849_ | new_A2864_;
  assign new_A2868_ = ~new_A2842_ | ~new_A2843_;
  assign new_A2867_ = new_A2849_ | new_A2864_;
  assign new_A2866_ = ~new_A2865_ & ~new_A2849_;
  assign new_A2865_ = new_A2849_ & new_A2864_;
  assign new_A2864_ = ~new_A2840_ | ~new_A2841_;
  assign new_A2863_ = new_A2841_ & new_A2853_;
  assign new_A2862_ = new_A2842_ | new_A2849_;
  assign new_A2861_ = new_A2842_ | new_A2843_;
  assign new_A2860_ = ~new_A2870_ | ~new_A2869_;
  assign new_A2859_ = new_A2868_ & new_A2861_;
  assign new_A2858_ = new_A2842_ ^ new_A2849_;
  assign new_A2857_ = ~new_A2866_ | ~new_A2867_;
  assign new_A2856_ = ~new_A2841_ ^ new_A2853_;
  assign new_A2855_ = new_A2863_ | new_A2840_;
  assign new_A2854_ = new_A2860_ & new_A2841_;
  assign new_A2853_ = new_A2862_ & new_A2861_;
  assign new_A2852_ = new_A2857_ & new_A2841_;
  assign new_A2851_ = new_A2859_ & new_A2858_;
  assign new_A2850_ = new_A2851_ ^ new_A2841_;
  assign new_A2849_ = new_A2839_ ^ new_A2840_;
  assign A2848 = new_A2849_ & new_A2856_;
  assign A2847 = new_A2849_ & new_A2855_;
  assign A2846 = new_A2854_ | new_A2853_;
  assign A2845 = new_A2852_ | new_A2851_;
  assign A2844 = new_A2850_ & new_A2849_;
  assign new_A2843_ = new_A7233_;
  assign new_A2842_ = new_A7200_;
  assign new_A2841_ = new_A7167_;
  assign new_A2840_ = new_A7134_;
  assign new_A2839_ = new_A7101_;
  assign new_A2806_ = new_A7068_;
  assign new_A2807_ = new_A7035_;
  assign new_A2808_ = new_A7002_;
  assign new_A2809_ = new_A6969_;
  assign new_A2810_ = new_A6940_;
  assign A2811 = new_A2817_ & new_A2816_;
  assign A2812 = new_A2819_ | new_A2818_;
  assign A2813 = new_A2821_ | new_A2820_;
  assign A2814 = new_A2816_ & new_A2822_;
  assign A2815 = new_A2816_ & new_A2823_;
  assign new_A2816_ = new_A2806_ ^ new_A2807_;
  assign new_A2817_ = new_A2818_ ^ new_A2808_;
  assign new_A2818_ = new_A2826_ & new_A2825_;
  assign new_A2819_ = new_A2824_ & new_A2808_;
  assign new_A2820_ = new_A2829_ & new_A2828_;
  assign new_A2821_ = new_A2827_ & new_A2808_;
  assign new_A2822_ = new_A2830_ | new_A2807_;
  assign new_A2823_ = ~new_A2808_ ^ new_A2820_;
  assign new_A2824_ = ~new_A2833_ | ~new_A2834_;
  assign new_A2825_ = new_A2809_ ^ new_A2816_;
  assign new_A2826_ = new_A2835_ & new_A2828_;
  assign new_A2827_ = ~new_A2837_ | ~new_A2836_;
  assign new_A2828_ = new_A2809_ | new_A2810_;
  assign new_A2829_ = new_A2809_ | new_A2816_;
  assign new_A2830_ = new_A2808_ & new_A2820_;
  assign new_A2831_ = ~new_A2807_ | ~new_A2808_;
  assign new_A2832_ = new_A2816_ & new_A2831_;
  assign new_A2833_ = ~new_A2832_ & ~new_A2816_;
  assign new_A2834_ = new_A2816_ | new_A2831_;
  assign new_A2835_ = ~new_A2809_ | ~new_A2810_;
  assign new_A2836_ = new_A2816_ | new_A2831_;
  assign new_A2837_ = ~new_A2816_ & ~new_A2838_;
  assign new_A2838_ = new_A2816_ & new_A2831_;
endmodule


